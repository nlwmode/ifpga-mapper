module top (\m0_addr_i[0]_pad , \m0_addr_i[10]_pad , \m0_addr_i[11]_pad , \m0_addr_i[12]_pad , \m0_addr_i[13]_pad , \m0_addr_i[14]_pad , \m0_addr_i[15]_pad , \m0_addr_i[16]_pad , \m0_addr_i[17]_pad , \m0_addr_i[18]_pad , \m0_addr_i[19]_pad , \m0_addr_i[1]_pad , \m0_addr_i[20]_pad , \m0_addr_i[21]_pad , \m0_addr_i[22]_pad , \m0_addr_i[23]_pad , \m0_addr_i[24]_pad , \m0_addr_i[25]_pad , \m0_addr_i[26]_pad , \m0_addr_i[27]_pad , \m0_addr_i[28]_pad , \m0_addr_i[29]_pad , \m0_addr_i[2]_pad , \m0_addr_i[30]_pad , \m0_addr_i[31]_pad , \m0_addr_i[3]_pad , \m0_addr_i[4]_pad , \m0_addr_i[5]_pad , \m0_addr_i[6]_pad , \m0_addr_i[7]_pad , \m0_addr_i[8]_pad , \m0_addr_i[9]_pad , \m0_cyc_i_pad , \m0_data_i[0]_pad , \m0_data_i[10]_pad , \m0_data_i[11]_pad , \m0_data_i[12]_pad , \m0_data_i[13]_pad , \m0_data_i[14]_pad , \m0_data_i[15]_pad , \m0_data_i[16]_pad , \m0_data_i[17]_pad , \m0_data_i[18]_pad , \m0_data_i[19]_pad , \m0_data_i[1]_pad , \m0_data_i[20]_pad , \m0_data_i[21]_pad , \m0_data_i[22]_pad , \m0_data_i[23]_pad , \m0_data_i[24]_pad , \m0_data_i[25]_pad , \m0_data_i[26]_pad , \m0_data_i[27]_pad , \m0_data_i[28]_pad , \m0_data_i[29]_pad , \m0_data_i[2]_pad , \m0_data_i[30]_pad , \m0_data_i[31]_pad , \m0_data_i[3]_pad , \m0_data_i[4]_pad , \m0_data_i[5]_pad , \m0_data_i[6]_pad , \m0_data_i[7]_pad , \m0_data_i[8]_pad , \m0_data_i[9]_pad , \m0_s0_cyc_o_reg/NET0131 , \m0_s10_cyc_o_reg/NET0131 , \m0_s11_cyc_o_reg/NET0131 , \m0_s12_cyc_o_reg/NET0131 , \m0_s13_cyc_o_reg/NET0131 , \m0_s14_cyc_o_reg/NET0131 , \m0_s15_cyc_o_reg/NET0131 , \m0_s1_cyc_o_reg/NET0131 , \m0_s2_cyc_o_reg/NET0131 , \m0_s3_cyc_o_reg/NET0131 , \m0_s4_cyc_o_reg/NET0131 , \m0_s5_cyc_o_reg/NET0131 , \m0_s6_cyc_o_reg/NET0131 , \m0_s7_cyc_o_reg/NET0131 , \m0_s8_cyc_o_reg/NET0131 , \m0_s9_cyc_o_reg/NET0131 , \m0_sel_i[0]_pad , \m0_sel_i[1]_pad , \m0_sel_i[2]_pad , \m0_sel_i[3]_pad , \m0_stb_i_pad , \m0_we_i_pad , \m1_addr_i[0]_pad , \m1_addr_i[10]_pad , \m1_addr_i[11]_pad , \m1_addr_i[12]_pad , \m1_addr_i[13]_pad , \m1_addr_i[14]_pad , \m1_addr_i[15]_pad , \m1_addr_i[16]_pad , \m1_addr_i[17]_pad , \m1_addr_i[18]_pad , \m1_addr_i[19]_pad , \m1_addr_i[1]_pad , \m1_addr_i[20]_pad , \m1_addr_i[21]_pad , \m1_addr_i[22]_pad , \m1_addr_i[23]_pad , \m1_addr_i[24]_pad , \m1_addr_i[25]_pad , \m1_addr_i[26]_pad , \m1_addr_i[27]_pad , \m1_addr_i[28]_pad , \m1_addr_i[29]_pad , \m1_addr_i[2]_pad , \m1_addr_i[30]_pad , \m1_addr_i[31]_pad , \m1_addr_i[3]_pad , \m1_addr_i[4]_pad , \m1_addr_i[5]_pad , \m1_addr_i[6]_pad , \m1_addr_i[7]_pad , \m1_addr_i[8]_pad , \m1_addr_i[9]_pad , \m1_cyc_i_pad , \m1_data_i[0]_pad , \m1_data_i[10]_pad , \m1_data_i[11]_pad , \m1_data_i[12]_pad , \m1_data_i[13]_pad , \m1_data_i[14]_pad , \m1_data_i[15]_pad , \m1_data_i[16]_pad , \m1_data_i[17]_pad , \m1_data_i[18]_pad , \m1_data_i[19]_pad , \m1_data_i[1]_pad , \m1_data_i[20]_pad , \m1_data_i[21]_pad , \m1_data_i[22]_pad , \m1_data_i[23]_pad , \m1_data_i[24]_pad , \m1_data_i[25]_pad , \m1_data_i[26]_pad , \m1_data_i[27]_pad , \m1_data_i[28]_pad , \m1_data_i[29]_pad , \m1_data_i[2]_pad , \m1_data_i[30]_pad , \m1_data_i[31]_pad , \m1_data_i[3]_pad , \m1_data_i[4]_pad , \m1_data_i[5]_pad , \m1_data_i[6]_pad , \m1_data_i[7]_pad , \m1_data_i[8]_pad , \m1_data_i[9]_pad , \m1_s0_cyc_o_reg/NET0131 , \m1_s10_cyc_o_reg/NET0131 , \m1_s11_cyc_o_reg/NET0131 , \m1_s12_cyc_o_reg/NET0131 , \m1_s13_cyc_o_reg/NET0131 , \m1_s14_cyc_o_reg/NET0131 , \m1_s15_cyc_o_reg/NET0131 , \m1_s1_cyc_o_reg/NET0131 , \m1_s2_cyc_o_reg/NET0131 , \m1_s3_cyc_o_reg/NET0131 , \m1_s4_cyc_o_reg/NET0131 , \m1_s5_cyc_o_reg/NET0131 , \m1_s6_cyc_o_reg/NET0131 , \m1_s7_cyc_o_reg/NET0131 , \m1_s8_cyc_o_reg/NET0131 , \m1_s9_cyc_o_reg/NET0131 , \m1_sel_i[0]_pad , \m1_sel_i[1]_pad , \m1_sel_i[2]_pad , \m1_sel_i[3]_pad , \m1_stb_i_pad , \m1_we_i_pad , \m2_addr_i[0]_pad , \m2_addr_i[10]_pad , \m2_addr_i[11]_pad , \m2_addr_i[12]_pad , \m2_addr_i[13]_pad , \m2_addr_i[14]_pad , \m2_addr_i[15]_pad , \m2_addr_i[16]_pad , \m2_addr_i[17]_pad , \m2_addr_i[18]_pad , \m2_addr_i[19]_pad , \m2_addr_i[1]_pad , \m2_addr_i[20]_pad , \m2_addr_i[21]_pad , \m2_addr_i[22]_pad , \m2_addr_i[23]_pad , \m2_addr_i[24]_pad , \m2_addr_i[25]_pad , \m2_addr_i[26]_pad , \m2_addr_i[27]_pad , \m2_addr_i[28]_pad , \m2_addr_i[29]_pad , \m2_addr_i[2]_pad , \m2_addr_i[30]_pad , \m2_addr_i[31]_pad , \m2_addr_i[3]_pad , \m2_addr_i[4]_pad , \m2_addr_i[5]_pad , \m2_addr_i[6]_pad , \m2_addr_i[7]_pad , \m2_addr_i[8]_pad , \m2_addr_i[9]_pad , \m2_cyc_i_pad , \m2_data_i[0]_pad , \m2_data_i[10]_pad , \m2_data_i[11]_pad , \m2_data_i[12]_pad , \m2_data_i[13]_pad , \m2_data_i[14]_pad , \m2_data_i[15]_pad , \m2_data_i[16]_pad , \m2_data_i[17]_pad , \m2_data_i[18]_pad , \m2_data_i[19]_pad , \m2_data_i[1]_pad , \m2_data_i[20]_pad , \m2_data_i[21]_pad , \m2_data_i[22]_pad , \m2_data_i[23]_pad , \m2_data_i[24]_pad , \m2_data_i[25]_pad , \m2_data_i[26]_pad , \m2_data_i[27]_pad , \m2_data_i[28]_pad , \m2_data_i[29]_pad , \m2_data_i[2]_pad , \m2_data_i[30]_pad , \m2_data_i[31]_pad , \m2_data_i[3]_pad , \m2_data_i[4]_pad , \m2_data_i[5]_pad , \m2_data_i[6]_pad , \m2_data_i[7]_pad , \m2_data_i[8]_pad , \m2_data_i[9]_pad , \m2_s0_cyc_o_reg/NET0131 , \m2_s10_cyc_o_reg/NET0131 , \m2_s11_cyc_o_reg/NET0131 , \m2_s12_cyc_o_reg/NET0131 , \m2_s13_cyc_o_reg/NET0131 , \m2_s14_cyc_o_reg/NET0131 , \m2_s15_cyc_o_reg/NET0131 , \m2_s1_cyc_o_reg/NET0131 , \m2_s2_cyc_o_reg/NET0131 , \m2_s3_cyc_o_reg/NET0131 , \m2_s4_cyc_o_reg/NET0131 , \m2_s5_cyc_o_reg/NET0131 , \m2_s6_cyc_o_reg/NET0131 , \m2_s7_cyc_o_reg/NET0131 , \m2_s8_cyc_o_reg/NET0131 , \m2_s9_cyc_o_reg/NET0131 , \m2_sel_i[0]_pad , \m2_sel_i[1]_pad , \m2_sel_i[2]_pad , \m2_sel_i[3]_pad , \m2_stb_i_pad , \m2_we_i_pad , \m3_addr_i[0]_pad , \m3_addr_i[10]_pad , \m3_addr_i[11]_pad , \m3_addr_i[12]_pad , \m3_addr_i[13]_pad , \m3_addr_i[14]_pad , \m3_addr_i[15]_pad , \m3_addr_i[16]_pad , \m3_addr_i[17]_pad , \m3_addr_i[18]_pad , \m3_addr_i[19]_pad , \m3_addr_i[1]_pad , \m3_addr_i[20]_pad , \m3_addr_i[21]_pad , \m3_addr_i[22]_pad , \m3_addr_i[23]_pad , \m3_addr_i[24]_pad , \m3_addr_i[25]_pad , \m3_addr_i[26]_pad , \m3_addr_i[27]_pad , \m3_addr_i[28]_pad , \m3_addr_i[29]_pad , \m3_addr_i[2]_pad , \m3_addr_i[30]_pad , \m3_addr_i[31]_pad , \m3_addr_i[3]_pad , \m3_addr_i[4]_pad , \m3_addr_i[5]_pad , \m3_addr_i[6]_pad , \m3_addr_i[7]_pad , \m3_addr_i[8]_pad , \m3_addr_i[9]_pad , \m3_cyc_i_pad , \m3_data_i[0]_pad , \m3_data_i[10]_pad , \m3_data_i[11]_pad , \m3_data_i[12]_pad , \m3_data_i[13]_pad , \m3_data_i[14]_pad , \m3_data_i[15]_pad , \m3_data_i[16]_pad , \m3_data_i[17]_pad , \m3_data_i[18]_pad , \m3_data_i[19]_pad , \m3_data_i[1]_pad , \m3_data_i[20]_pad , \m3_data_i[21]_pad , \m3_data_i[22]_pad , \m3_data_i[23]_pad , \m3_data_i[24]_pad , \m3_data_i[25]_pad , \m3_data_i[26]_pad , \m3_data_i[27]_pad , \m3_data_i[28]_pad , \m3_data_i[29]_pad , \m3_data_i[2]_pad , \m3_data_i[30]_pad , \m3_data_i[31]_pad , \m3_data_i[3]_pad , \m3_data_i[4]_pad , \m3_data_i[5]_pad , \m3_data_i[6]_pad , \m3_data_i[7]_pad , \m3_data_i[8]_pad , \m3_data_i[9]_pad , \m3_s0_cyc_o_reg/NET0131 , \m3_s10_cyc_o_reg/NET0131 , \m3_s11_cyc_o_reg/NET0131 , \m3_s12_cyc_o_reg/NET0131 , \m3_s13_cyc_o_reg/NET0131 , \m3_s14_cyc_o_reg/NET0131 , \m3_s15_cyc_o_reg/NET0131 , \m3_s1_cyc_o_reg/NET0131 , \m3_s2_cyc_o_reg/NET0131 , \m3_s3_cyc_o_reg/NET0131 , \m3_s4_cyc_o_reg/NET0131 , \m3_s5_cyc_o_reg/NET0131 , \m3_s6_cyc_o_reg/NET0131 , \m3_s7_cyc_o_reg/NET0131 , \m3_s8_cyc_o_reg/NET0131 , \m3_s9_cyc_o_reg/NET0131 , \m3_sel_i[0]_pad , \m3_sel_i[1]_pad , \m3_sel_i[2]_pad , \m3_sel_i[3]_pad , \m3_stb_i_pad , \m3_we_i_pad , \m4_addr_i[0]_pad , \m4_addr_i[10]_pad , \m4_addr_i[11]_pad , \m4_addr_i[12]_pad , \m4_addr_i[13]_pad , \m4_addr_i[14]_pad , \m4_addr_i[15]_pad , \m4_addr_i[16]_pad , \m4_addr_i[17]_pad , \m4_addr_i[18]_pad , \m4_addr_i[19]_pad , \m4_addr_i[1]_pad , \m4_addr_i[20]_pad , \m4_addr_i[21]_pad , \m4_addr_i[22]_pad , \m4_addr_i[23]_pad , \m4_addr_i[24]_pad , \m4_addr_i[25]_pad , \m4_addr_i[26]_pad , \m4_addr_i[27]_pad , \m4_addr_i[28]_pad , \m4_addr_i[29]_pad , \m4_addr_i[2]_pad , \m4_addr_i[30]_pad , \m4_addr_i[31]_pad , \m4_addr_i[3]_pad , \m4_addr_i[4]_pad , \m4_addr_i[5]_pad , \m4_addr_i[6]_pad , \m4_addr_i[7]_pad , \m4_addr_i[8]_pad , \m4_addr_i[9]_pad , \m4_cyc_i_pad , \m4_data_i[0]_pad , \m4_data_i[10]_pad , \m4_data_i[11]_pad , \m4_data_i[12]_pad , \m4_data_i[13]_pad , \m4_data_i[14]_pad , \m4_data_i[15]_pad , \m4_data_i[16]_pad , \m4_data_i[17]_pad , \m4_data_i[18]_pad , \m4_data_i[19]_pad , \m4_data_i[1]_pad , \m4_data_i[20]_pad , \m4_data_i[21]_pad , \m4_data_i[22]_pad , \m4_data_i[23]_pad , \m4_data_i[24]_pad , \m4_data_i[25]_pad , \m4_data_i[26]_pad , \m4_data_i[27]_pad , \m4_data_i[28]_pad , \m4_data_i[29]_pad , \m4_data_i[2]_pad , \m4_data_i[30]_pad , \m4_data_i[31]_pad , \m4_data_i[3]_pad , \m4_data_i[4]_pad , \m4_data_i[5]_pad , \m4_data_i[6]_pad , \m4_data_i[7]_pad , \m4_data_i[8]_pad , \m4_data_i[9]_pad , \m4_s0_cyc_o_reg/NET0131 , \m4_s10_cyc_o_reg/NET0131 , \m4_s11_cyc_o_reg/NET0131 , \m4_s12_cyc_o_reg/NET0131 , \m4_s13_cyc_o_reg/NET0131 , \m4_s14_cyc_o_reg/NET0131 , \m4_s15_cyc_o_reg/NET0131 , \m4_s1_cyc_o_reg/NET0131 , \m4_s2_cyc_o_reg/NET0131 , \m4_s3_cyc_o_reg/NET0131 , \m4_s4_cyc_o_reg/NET0131 , \m4_s5_cyc_o_reg/NET0131 , \m4_s6_cyc_o_reg/NET0131 , \m4_s7_cyc_o_reg/NET0131 , \m4_s8_cyc_o_reg/NET0131 , \m4_s9_cyc_o_reg/NET0131 , \m4_sel_i[0]_pad , \m4_sel_i[1]_pad , \m4_sel_i[2]_pad , \m4_sel_i[3]_pad , \m4_stb_i_pad , \m4_we_i_pad , \m5_addr_i[0]_pad , \m5_addr_i[10]_pad , \m5_addr_i[11]_pad , \m5_addr_i[12]_pad , \m5_addr_i[13]_pad , \m5_addr_i[14]_pad , \m5_addr_i[15]_pad , \m5_addr_i[16]_pad , \m5_addr_i[17]_pad , \m5_addr_i[18]_pad , \m5_addr_i[19]_pad , \m5_addr_i[1]_pad , \m5_addr_i[20]_pad , \m5_addr_i[21]_pad , \m5_addr_i[22]_pad , \m5_addr_i[23]_pad , \m5_addr_i[24]_pad , \m5_addr_i[25]_pad , \m5_addr_i[26]_pad , \m5_addr_i[27]_pad , \m5_addr_i[28]_pad , \m5_addr_i[29]_pad , \m5_addr_i[2]_pad , \m5_addr_i[30]_pad , \m5_addr_i[31]_pad , \m5_addr_i[3]_pad , \m5_addr_i[4]_pad , \m5_addr_i[5]_pad , \m5_addr_i[6]_pad , \m5_addr_i[7]_pad , \m5_addr_i[8]_pad , \m5_addr_i[9]_pad , \m5_cyc_i_pad , \m5_data_i[0]_pad , \m5_data_i[10]_pad , \m5_data_i[11]_pad , \m5_data_i[12]_pad , \m5_data_i[13]_pad , \m5_data_i[14]_pad , \m5_data_i[15]_pad , \m5_data_i[16]_pad , \m5_data_i[17]_pad , \m5_data_i[18]_pad , \m5_data_i[19]_pad , \m5_data_i[1]_pad , \m5_data_i[20]_pad , \m5_data_i[21]_pad , \m5_data_i[22]_pad , \m5_data_i[23]_pad , \m5_data_i[24]_pad , \m5_data_i[25]_pad , \m5_data_i[26]_pad , \m5_data_i[27]_pad , \m5_data_i[28]_pad , \m5_data_i[29]_pad , \m5_data_i[2]_pad , \m5_data_i[30]_pad , \m5_data_i[31]_pad , \m5_data_i[3]_pad , \m5_data_i[4]_pad , \m5_data_i[5]_pad , \m5_data_i[6]_pad , \m5_data_i[7]_pad , \m5_data_i[8]_pad , \m5_data_i[9]_pad , \m5_s0_cyc_o_reg/NET0131 , \m5_s10_cyc_o_reg/NET0131 , \m5_s11_cyc_o_reg/NET0131 , \m5_s12_cyc_o_reg/NET0131 , \m5_s13_cyc_o_reg/NET0131 , \m5_s14_cyc_o_reg/NET0131 , \m5_s15_cyc_o_reg/NET0131 , \m5_s1_cyc_o_reg/NET0131 , \m5_s2_cyc_o_reg/NET0131 , \m5_s3_cyc_o_reg/NET0131 , \m5_s4_cyc_o_reg/NET0131 , \m5_s5_cyc_o_reg/NET0131 , \m5_s6_cyc_o_reg/NET0131 , \m5_s7_cyc_o_reg/NET0131 , \m5_s8_cyc_o_reg/NET0131 , \m5_s9_cyc_o_reg/NET0131 , \m5_sel_i[0]_pad , \m5_sel_i[1]_pad , \m5_sel_i[2]_pad , \m5_sel_i[3]_pad , \m5_stb_i_pad , \m5_we_i_pad , \m6_addr_i[0]_pad , \m6_addr_i[10]_pad , \m6_addr_i[11]_pad , \m6_addr_i[12]_pad , \m6_addr_i[13]_pad , \m6_addr_i[14]_pad , \m6_addr_i[15]_pad , \m6_addr_i[16]_pad , \m6_addr_i[17]_pad , \m6_addr_i[18]_pad , \m6_addr_i[19]_pad , \m6_addr_i[1]_pad , \m6_addr_i[20]_pad , \m6_addr_i[21]_pad , \m6_addr_i[22]_pad , \m6_addr_i[23]_pad , \m6_addr_i[24]_pad , \m6_addr_i[25]_pad , \m6_addr_i[26]_pad , \m6_addr_i[27]_pad , \m6_addr_i[28]_pad , \m6_addr_i[29]_pad , \m6_addr_i[2]_pad , \m6_addr_i[30]_pad , \m6_addr_i[31]_pad , \m6_addr_i[3]_pad , \m6_addr_i[4]_pad , \m6_addr_i[5]_pad , \m6_addr_i[6]_pad , \m6_addr_i[7]_pad , \m6_addr_i[8]_pad , \m6_addr_i[9]_pad , \m6_cyc_i_pad , \m6_data_i[0]_pad , \m6_data_i[10]_pad , \m6_data_i[11]_pad , \m6_data_i[12]_pad , \m6_data_i[13]_pad , \m6_data_i[14]_pad , \m6_data_i[15]_pad , \m6_data_i[16]_pad , \m6_data_i[17]_pad , \m6_data_i[18]_pad , \m6_data_i[19]_pad , \m6_data_i[1]_pad , \m6_data_i[20]_pad , \m6_data_i[21]_pad , \m6_data_i[22]_pad , \m6_data_i[23]_pad , \m6_data_i[24]_pad , \m6_data_i[25]_pad , \m6_data_i[26]_pad , \m6_data_i[27]_pad , \m6_data_i[28]_pad , \m6_data_i[29]_pad , \m6_data_i[2]_pad , \m6_data_i[30]_pad , \m6_data_i[31]_pad , \m6_data_i[3]_pad , \m6_data_i[4]_pad , \m6_data_i[5]_pad , \m6_data_i[6]_pad , \m6_data_i[7]_pad , \m6_data_i[8]_pad , \m6_data_i[9]_pad , \m6_s0_cyc_o_reg/NET0131 , \m6_s10_cyc_o_reg/NET0131 , \m6_s11_cyc_o_reg/NET0131 , \m6_s12_cyc_o_reg/NET0131 , \m6_s13_cyc_o_reg/NET0131 , \m6_s14_cyc_o_reg/NET0131 , \m6_s15_cyc_o_reg/NET0131 , \m6_s1_cyc_o_reg/NET0131 , \m6_s2_cyc_o_reg/NET0131 , \m6_s3_cyc_o_reg/NET0131 , \m6_s4_cyc_o_reg/NET0131 , \m6_s5_cyc_o_reg/NET0131 , \m6_s6_cyc_o_reg/NET0131 , \m6_s7_cyc_o_reg/NET0131 , \m6_s8_cyc_o_reg/NET0131 , \m6_s9_cyc_o_reg/NET0131 , \m6_sel_i[0]_pad , \m6_sel_i[1]_pad , \m6_sel_i[2]_pad , \m6_sel_i[3]_pad , \m6_stb_i_pad , \m6_we_i_pad , \m7_addr_i[0]_pad , \m7_addr_i[10]_pad , \m7_addr_i[11]_pad , \m7_addr_i[12]_pad , \m7_addr_i[13]_pad , \m7_addr_i[14]_pad , \m7_addr_i[15]_pad , \m7_addr_i[16]_pad , \m7_addr_i[17]_pad , \m7_addr_i[18]_pad , \m7_addr_i[19]_pad , \m7_addr_i[1]_pad , \m7_addr_i[20]_pad , \m7_addr_i[21]_pad , \m7_addr_i[22]_pad , \m7_addr_i[23]_pad , \m7_addr_i[24]_pad , \m7_addr_i[25]_pad , \m7_addr_i[26]_pad , \m7_addr_i[27]_pad , \m7_addr_i[28]_pad , \m7_addr_i[29]_pad , \m7_addr_i[2]_pad , \m7_addr_i[30]_pad , \m7_addr_i[31]_pad , \m7_addr_i[3]_pad , \m7_addr_i[4]_pad , \m7_addr_i[5]_pad , \m7_addr_i[6]_pad , \m7_addr_i[7]_pad , \m7_addr_i[8]_pad , \m7_addr_i[9]_pad , \m7_cyc_i_pad , \m7_data_i[0]_pad , \m7_data_i[10]_pad , \m7_data_i[11]_pad , \m7_data_i[12]_pad , \m7_data_i[13]_pad , \m7_data_i[14]_pad , \m7_data_i[15]_pad , \m7_data_i[16]_pad , \m7_data_i[17]_pad , \m7_data_i[18]_pad , \m7_data_i[19]_pad , \m7_data_i[1]_pad , \m7_data_i[20]_pad , \m7_data_i[21]_pad , \m7_data_i[22]_pad , \m7_data_i[23]_pad , \m7_data_i[24]_pad , \m7_data_i[25]_pad , \m7_data_i[26]_pad , \m7_data_i[27]_pad , \m7_data_i[28]_pad , \m7_data_i[29]_pad , \m7_data_i[2]_pad , \m7_data_i[30]_pad , \m7_data_i[31]_pad , \m7_data_i[3]_pad , \m7_data_i[4]_pad , \m7_data_i[5]_pad , \m7_data_i[6]_pad , \m7_data_i[7]_pad , \m7_data_i[8]_pad , \m7_data_i[9]_pad , \m7_s0_cyc_o_reg/NET0131 , \m7_s10_cyc_o_reg/NET0131 , \m7_s11_cyc_o_reg/NET0131 , \m7_s12_cyc_o_reg/NET0131 , \m7_s13_cyc_o_reg/NET0131 , \m7_s14_cyc_o_reg/NET0131 , \m7_s15_cyc_o_reg/NET0131 , \m7_s1_cyc_o_reg/NET0131 , \m7_s2_cyc_o_reg/NET0131 , \m7_s3_cyc_o_reg/NET0131 , \m7_s4_cyc_o_reg/NET0131 , \m7_s5_cyc_o_reg/NET0131 , \m7_s6_cyc_o_reg/NET0131 , \m7_s7_cyc_o_reg/NET0131 , \m7_s8_cyc_o_reg/NET0131 , \m7_s9_cyc_o_reg/NET0131 , \m7_sel_i[0]_pad , \m7_sel_i[1]_pad , \m7_sel_i[2]_pad , \m7_sel_i[3]_pad , \m7_stb_i_pad , \m7_we_i_pad , \rf_conf0_reg[0]/NET0131 , \rf_conf0_reg[10]/NET0131 , \rf_conf0_reg[11]/NET0131 , \rf_conf0_reg[12]/NET0131 , \rf_conf0_reg[13]/NET0131 , \rf_conf0_reg[14]/NET0131 , \rf_conf0_reg[15]/NET0131 , \rf_conf0_reg[1]/NET0131 , \rf_conf0_reg[2]/NET0131 , \rf_conf0_reg[3]/NET0131 , \rf_conf0_reg[4]/NET0131 , \rf_conf0_reg[5]/NET0131 , \rf_conf0_reg[6]/NET0131 , \rf_conf0_reg[7]/NET0131 , \rf_conf0_reg[8]/NET0131 , \rf_conf0_reg[9]/NET0131 , \rf_conf10_reg[0]/NET0131 , \rf_conf10_reg[10]/NET0131 , \rf_conf10_reg[11]/NET0131 , \rf_conf10_reg[12]/NET0131 , \rf_conf10_reg[13]/NET0131 , \rf_conf10_reg[14]/NET0131 , \rf_conf10_reg[15]/NET0131 , \rf_conf10_reg[1]/NET0131 , \rf_conf10_reg[2]/NET0131 , \rf_conf10_reg[3]/NET0131 , \rf_conf10_reg[4]/NET0131 , \rf_conf10_reg[5]/NET0131 , \rf_conf10_reg[6]/NET0131 , \rf_conf10_reg[7]/NET0131 , \rf_conf10_reg[8]/NET0131 , \rf_conf10_reg[9]/NET0131 , \rf_conf11_reg[0]/NET0131 , \rf_conf11_reg[10]/NET0131 , \rf_conf11_reg[11]/NET0131 , \rf_conf11_reg[12]/NET0131 , \rf_conf11_reg[13]/NET0131 , \rf_conf11_reg[14]/NET0131 , \rf_conf11_reg[15]/NET0131 , \rf_conf11_reg[1]/NET0131 , \rf_conf11_reg[2]/NET0131 , \rf_conf11_reg[3]/NET0131 , \rf_conf11_reg[4]/NET0131 , \rf_conf11_reg[5]/NET0131 , \rf_conf11_reg[6]/NET0131 , \rf_conf11_reg[7]/NET0131 , \rf_conf11_reg[8]/NET0131 , \rf_conf11_reg[9]/NET0131 , \rf_conf12_reg[0]/NET0131 , \rf_conf12_reg[10]/NET0131 , \rf_conf12_reg[11]/NET0131 , \rf_conf12_reg[12]/NET0131 , \rf_conf12_reg[13]/NET0131 , \rf_conf12_reg[14]/NET0131 , \rf_conf12_reg[15]/NET0131 , \rf_conf12_reg[1]/NET0131 , \rf_conf12_reg[2]/NET0131 , \rf_conf12_reg[3]/NET0131 , \rf_conf12_reg[4]/NET0131 , \rf_conf12_reg[5]/NET0131 , \rf_conf12_reg[6]/NET0131 , \rf_conf12_reg[7]/NET0131 , \rf_conf12_reg[8]/NET0131 , \rf_conf12_reg[9]/NET0131 , \rf_conf13_reg[0]/NET0131 , \rf_conf13_reg[10]/NET0131 , \rf_conf13_reg[11]/NET0131 , \rf_conf13_reg[12]/NET0131 , \rf_conf13_reg[13]/NET0131 , \rf_conf13_reg[14]/NET0131 , \rf_conf13_reg[15]/NET0131 , \rf_conf13_reg[1]/NET0131 , \rf_conf13_reg[2]/NET0131 , \rf_conf13_reg[3]/NET0131 , \rf_conf13_reg[4]/NET0131 , \rf_conf13_reg[5]/NET0131 , \rf_conf13_reg[6]/NET0131 , \rf_conf13_reg[7]/NET0131 , \rf_conf13_reg[8]/NET0131 , \rf_conf13_reg[9]/NET0131 , \rf_conf14_reg[0]/NET0131 , \rf_conf14_reg[10]/NET0131 , \rf_conf14_reg[11]/NET0131 , \rf_conf14_reg[12]/NET0131 , \rf_conf14_reg[13]/NET0131 , \rf_conf14_reg[14]/NET0131 , \rf_conf14_reg[15]/NET0131 , \rf_conf14_reg[1]/NET0131 , \rf_conf14_reg[2]/NET0131 , \rf_conf14_reg[3]/NET0131 , \rf_conf14_reg[4]/NET0131 , \rf_conf14_reg[5]/NET0131 , \rf_conf14_reg[6]/NET0131 , \rf_conf14_reg[7]/NET0131 , \rf_conf14_reg[8]/NET0131 , \rf_conf14_reg[9]/NET0131 , \rf_conf15_reg[0]/NET0131 , \rf_conf15_reg[10]/NET0131 , \rf_conf15_reg[11]/NET0131 , \rf_conf15_reg[12]/NET0131 , \rf_conf15_reg[13]/NET0131 , \rf_conf15_reg[14]/NET0131 , \rf_conf15_reg[15]/NET0131 , \rf_conf15_reg[1]/NET0131 , \rf_conf15_reg[2]/NET0131 , \rf_conf15_reg[3]/NET0131 , \rf_conf15_reg[4]/NET0131 , \rf_conf15_reg[5]/NET0131 , \rf_conf15_reg[6]/NET0131 , \rf_conf15_reg[7]/NET0131 , \rf_conf15_reg[8]/NET0131 , \rf_conf15_reg[9]/NET0131 , \rf_conf1_reg[0]/NET0131 , \rf_conf1_reg[10]/NET0131 , \rf_conf1_reg[11]/NET0131 , \rf_conf1_reg[12]/NET0131 , \rf_conf1_reg[13]/NET0131 , \rf_conf1_reg[14]/NET0131 , \rf_conf1_reg[15]/NET0131 , \rf_conf1_reg[1]/NET0131 , \rf_conf1_reg[2]/NET0131 , \rf_conf1_reg[3]/NET0131 , \rf_conf1_reg[4]/NET0131 , \rf_conf1_reg[5]/NET0131 , \rf_conf1_reg[6]/NET0131 , \rf_conf1_reg[7]/NET0131 , \rf_conf1_reg[8]/NET0131 , \rf_conf1_reg[9]/NET0131 , \rf_conf2_reg[0]/NET0131 , \rf_conf2_reg[10]/NET0131 , \rf_conf2_reg[11]/NET0131 , \rf_conf2_reg[12]/NET0131 , \rf_conf2_reg[13]/NET0131 , \rf_conf2_reg[14]/NET0131 , \rf_conf2_reg[15]/NET0131 , \rf_conf2_reg[1]/NET0131 , \rf_conf2_reg[2]/NET0131 , \rf_conf2_reg[3]/NET0131 , \rf_conf2_reg[4]/NET0131 , \rf_conf2_reg[5]/NET0131 , \rf_conf2_reg[6]/NET0131 , \rf_conf2_reg[7]/NET0131 , \rf_conf2_reg[8]/NET0131 , \rf_conf2_reg[9]/NET0131 , \rf_conf3_reg[0]/NET0131 , \rf_conf3_reg[10]/NET0131 , \rf_conf3_reg[11]/NET0131 , \rf_conf3_reg[12]/NET0131 , \rf_conf3_reg[13]/NET0131 , \rf_conf3_reg[14]/NET0131 , \rf_conf3_reg[15]/NET0131 , \rf_conf3_reg[1]/NET0131 , \rf_conf3_reg[2]/NET0131 , \rf_conf3_reg[3]/NET0131 , \rf_conf3_reg[4]/NET0131 , \rf_conf3_reg[5]/NET0131 , \rf_conf3_reg[6]/NET0131 , \rf_conf3_reg[7]/NET0131 , \rf_conf3_reg[8]/NET0131 , \rf_conf3_reg[9]/NET0131 , \rf_conf4_reg[0]/NET0131 , \rf_conf4_reg[10]/NET0131 , \rf_conf4_reg[11]/NET0131 , \rf_conf4_reg[12]/NET0131 , \rf_conf4_reg[13]/NET0131 , \rf_conf4_reg[14]/NET0131 , \rf_conf4_reg[15]/NET0131 , \rf_conf4_reg[1]/NET0131 , \rf_conf4_reg[2]/NET0131 , \rf_conf4_reg[3]/NET0131 , \rf_conf4_reg[4]/NET0131 , \rf_conf4_reg[5]/NET0131 , \rf_conf4_reg[6]/NET0131 , \rf_conf4_reg[7]/NET0131 , \rf_conf4_reg[8]/NET0131 , \rf_conf4_reg[9]/NET0131 , \rf_conf5_reg[0]/NET0131 , \rf_conf5_reg[10]/NET0131 , \rf_conf5_reg[11]/NET0131 , \rf_conf5_reg[12]/NET0131 , \rf_conf5_reg[13]/NET0131 , \rf_conf5_reg[14]/NET0131 , \rf_conf5_reg[15]/NET0131 , \rf_conf5_reg[1]/NET0131 , \rf_conf5_reg[2]/NET0131 , \rf_conf5_reg[3]/NET0131 , \rf_conf5_reg[4]/NET0131 , \rf_conf5_reg[5]/NET0131 , \rf_conf5_reg[6]/NET0131 , \rf_conf5_reg[7]/NET0131 , \rf_conf5_reg[8]/NET0131 , \rf_conf5_reg[9]/NET0131 , \rf_conf6_reg[0]/NET0131 , \rf_conf6_reg[10]/NET0131 , \rf_conf6_reg[11]/NET0131 , \rf_conf6_reg[12]/NET0131 , \rf_conf6_reg[13]/NET0131 , \rf_conf6_reg[14]/NET0131 , \rf_conf6_reg[15]/NET0131 , \rf_conf6_reg[1]/NET0131 , \rf_conf6_reg[2]/NET0131 , \rf_conf6_reg[3]/NET0131 , \rf_conf6_reg[4]/NET0131 , \rf_conf6_reg[5]/NET0131 , \rf_conf6_reg[6]/NET0131 , \rf_conf6_reg[7]/NET0131 , \rf_conf6_reg[8]/NET0131 , \rf_conf6_reg[9]/NET0131 , \rf_conf7_reg[0]/NET0131 , \rf_conf7_reg[10]/NET0131 , \rf_conf7_reg[11]/NET0131 , \rf_conf7_reg[12]/NET0131 , \rf_conf7_reg[13]/NET0131 , \rf_conf7_reg[14]/NET0131 , \rf_conf7_reg[15]/NET0131 , \rf_conf7_reg[1]/NET0131 , \rf_conf7_reg[2]/NET0131 , \rf_conf7_reg[3]/NET0131 , \rf_conf7_reg[4]/NET0131 , \rf_conf7_reg[5]/NET0131 , \rf_conf7_reg[6]/NET0131 , \rf_conf7_reg[7]/NET0131 , \rf_conf7_reg[8]/NET0131 , \rf_conf7_reg[9]/NET0131 , \rf_conf8_reg[0]/NET0131 , \rf_conf8_reg[10]/NET0131 , \rf_conf8_reg[11]/NET0131 , \rf_conf8_reg[12]/NET0131 , \rf_conf8_reg[13]/NET0131 , \rf_conf8_reg[14]/NET0131 , \rf_conf8_reg[15]/NET0131 , \rf_conf8_reg[1]/NET0131 , \rf_conf8_reg[2]/NET0131 , \rf_conf8_reg[3]/NET0131 , \rf_conf8_reg[4]/NET0131 , \rf_conf8_reg[5]/NET0131 , \rf_conf8_reg[6]/NET0131 , \rf_conf8_reg[7]/NET0131 , \rf_conf8_reg[8]/NET0131 , \rf_conf8_reg[9]/NET0131 , \rf_conf9_reg[0]/NET0131 , \rf_conf9_reg[10]/NET0131 , \rf_conf9_reg[11]/NET0131 , \rf_conf9_reg[12]/NET0131 , \rf_conf9_reg[13]/NET0131 , \rf_conf9_reg[14]/NET0131 , \rf_conf9_reg[15]/NET0131 , \rf_conf9_reg[1]/NET0131 , \rf_conf9_reg[2]/NET0131 , \rf_conf9_reg[3]/NET0131 , \rf_conf9_reg[4]/NET0131 , \rf_conf9_reg[5]/NET0131 , \rf_conf9_reg[6]/NET0131 , \rf_conf9_reg[7]/NET0131 , \rf_conf9_reg[8]/NET0131 , \rf_conf9_reg[9]/NET0131 , \rf_rf_ack_reg/P0001 , \rf_rf_dout_reg[0]/P0001 , \rf_rf_dout_reg[10]/P0001 , \rf_rf_dout_reg[11]/P0001 , \rf_rf_dout_reg[12]/P0001 , \rf_rf_dout_reg[13]/P0001 , \rf_rf_dout_reg[14]/P0001 , \rf_rf_dout_reg[15]/P0001 , \rf_rf_dout_reg[1]/P0001 , \rf_rf_dout_reg[2]/P0001 , \rf_rf_dout_reg[3]/P0001 , \rf_rf_dout_reg[4]/P0001 , \rf_rf_dout_reg[5]/P0001 , \rf_rf_dout_reg[6]/P0001 , \rf_rf_dout_reg[7]/P0001 , \rf_rf_dout_reg[8]/P0001 , \rf_rf_dout_reg[9]/P0001 , \rf_rf_we_reg/P0001 , rst_i_pad, \s0_ack_i_pad , \s0_data_i[0]_pad , \s0_data_i[10]_pad , \s0_data_i[11]_pad , \s0_data_i[12]_pad , \s0_data_i[13]_pad , \s0_data_i[14]_pad , \s0_data_i[15]_pad , \s0_data_i[16]_pad , \s0_data_i[17]_pad , \s0_data_i[18]_pad , \s0_data_i[19]_pad , \s0_data_i[1]_pad , \s0_data_i[20]_pad , \s0_data_i[21]_pad , \s0_data_i[22]_pad , \s0_data_i[23]_pad , \s0_data_i[24]_pad , \s0_data_i[25]_pad , \s0_data_i[26]_pad , \s0_data_i[27]_pad , \s0_data_i[28]_pad , \s0_data_i[29]_pad , \s0_data_i[2]_pad , \s0_data_i[30]_pad , \s0_data_i[31]_pad , \s0_data_i[3]_pad , \s0_data_i[4]_pad , \s0_data_i[5]_pad , \s0_data_i[6]_pad , \s0_data_i[7]_pad , \s0_data_i[8]_pad , \s0_data_i[9]_pad , \s0_err_i_pad , \s0_m0_cyc_r_reg/P0001 , \s0_m1_cyc_r_reg/P0001 , \s0_m2_cyc_r_reg/P0001 , \s0_m3_cyc_r_reg/P0001 , \s0_m4_cyc_r_reg/P0001 , \s0_m5_cyc_r_reg/P0001 , \s0_m6_cyc_r_reg/P0001 , \s0_m7_cyc_r_reg/P0001 , \s0_msel_arb0_state_reg[0]/NET0131 , \s0_msel_arb0_state_reg[1]/NET0131 , \s0_msel_arb0_state_reg[2]/NET0131 , \s0_msel_arb1_state_reg[0]/NET0131 , \s0_msel_arb1_state_reg[1]/NET0131 , \s0_msel_arb1_state_reg[2]/NET0131 , \s0_msel_arb2_state_reg[0]/NET0131 , \s0_msel_arb2_state_reg[1]/NET0131 , \s0_msel_arb2_state_reg[2]/NET0131 , \s0_msel_arb3_state_reg[0]/NET0131 , \s0_msel_arb3_state_reg[1]/NET0131 , \s0_msel_arb3_state_reg[2]/NET0131 , \s0_msel_pri_out_reg[0]/NET0131 , \s0_msel_pri_out_reg[1]/NET0131 , \s0_next_reg/P0001 , \s0_rty_i_pad , \s10_ack_i_pad , \s10_data_i[0]_pad , \s10_data_i[10]_pad , \s10_data_i[11]_pad , \s10_data_i[12]_pad , \s10_data_i[13]_pad , \s10_data_i[14]_pad , \s10_data_i[15]_pad , \s10_data_i[16]_pad , \s10_data_i[17]_pad , \s10_data_i[18]_pad , \s10_data_i[19]_pad , \s10_data_i[1]_pad , \s10_data_i[20]_pad , \s10_data_i[21]_pad , \s10_data_i[22]_pad , \s10_data_i[23]_pad , \s10_data_i[24]_pad , \s10_data_i[25]_pad , \s10_data_i[26]_pad , \s10_data_i[27]_pad , \s10_data_i[28]_pad , \s10_data_i[29]_pad , \s10_data_i[2]_pad , \s10_data_i[30]_pad , \s10_data_i[31]_pad , \s10_data_i[3]_pad , \s10_data_i[4]_pad , \s10_data_i[5]_pad , \s10_data_i[6]_pad , \s10_data_i[7]_pad , \s10_data_i[8]_pad , \s10_data_i[9]_pad , \s10_err_i_pad , \s10_m0_cyc_r_reg/P0001 , \s10_m1_cyc_r_reg/P0001 , \s10_m2_cyc_r_reg/P0001 , \s10_m3_cyc_r_reg/P0001 , \s10_m4_cyc_r_reg/P0001 , \s10_m5_cyc_r_reg/P0001 , \s10_m6_cyc_r_reg/P0001 , \s10_m7_cyc_r_reg/P0001 , \s10_msel_arb0_state_reg[0]/NET0131 , \s10_msel_arb0_state_reg[1]/NET0131 , \s10_msel_arb0_state_reg[2]/NET0131 , \s10_msel_arb1_state_reg[0]/NET0131 , \s10_msel_arb1_state_reg[1]/NET0131 , \s10_msel_arb1_state_reg[2]/NET0131 , \s10_msel_arb2_state_reg[0]/NET0131 , \s10_msel_arb2_state_reg[1]/NET0131 , \s10_msel_arb2_state_reg[2]/NET0131 , \s10_msel_arb3_state_reg[0]/NET0131 , \s10_msel_arb3_state_reg[1]/NET0131 , \s10_msel_arb3_state_reg[2]/NET0131 , \s10_msel_pri_out_reg[0]/NET0131 , \s10_msel_pri_out_reg[1]/NET0131 , \s10_next_reg/P0001 , \s10_rty_i_pad , \s11_ack_i_pad , \s11_data_i[0]_pad , \s11_data_i[10]_pad , \s11_data_i[11]_pad , \s11_data_i[12]_pad , \s11_data_i[13]_pad , \s11_data_i[14]_pad , \s11_data_i[15]_pad , \s11_data_i[16]_pad , \s11_data_i[17]_pad , \s11_data_i[18]_pad , \s11_data_i[19]_pad , \s11_data_i[1]_pad , \s11_data_i[20]_pad , \s11_data_i[21]_pad , \s11_data_i[22]_pad , \s11_data_i[23]_pad , \s11_data_i[24]_pad , \s11_data_i[25]_pad , \s11_data_i[26]_pad , \s11_data_i[27]_pad , \s11_data_i[28]_pad , \s11_data_i[29]_pad , \s11_data_i[2]_pad , \s11_data_i[30]_pad , \s11_data_i[31]_pad , \s11_data_i[3]_pad , \s11_data_i[4]_pad , \s11_data_i[5]_pad , \s11_data_i[6]_pad , \s11_data_i[7]_pad , \s11_data_i[8]_pad , \s11_data_i[9]_pad , \s11_err_i_pad , \s11_m0_cyc_r_reg/P0001 , \s11_m1_cyc_r_reg/P0001 , \s11_m2_cyc_r_reg/P0001 , \s11_m3_cyc_r_reg/P0001 , \s11_m4_cyc_r_reg/P0001 , \s11_m5_cyc_r_reg/P0001 , \s11_m6_cyc_r_reg/P0001 , \s11_m7_cyc_r_reg/P0001 , \s11_msel_arb0_state_reg[0]/NET0131 , \s11_msel_arb0_state_reg[1]/NET0131 , \s11_msel_arb0_state_reg[2]/NET0131 , \s11_msel_arb1_state_reg[0]/NET0131 , \s11_msel_arb1_state_reg[1]/NET0131 , \s11_msel_arb1_state_reg[2]/NET0131 , \s11_msel_arb2_state_reg[0]/NET0131 , \s11_msel_arb2_state_reg[1]/NET0131 , \s11_msel_arb2_state_reg[2]/NET0131 , \s11_msel_arb3_state_reg[0]/NET0131 , \s11_msel_arb3_state_reg[1]/NET0131 , \s11_msel_arb3_state_reg[2]/NET0131 , \s11_msel_pri_out_reg[0]/NET0131 , \s11_msel_pri_out_reg[1]/NET0131 , \s11_next_reg/P0001 , \s11_rty_i_pad , \s12_ack_i_pad , \s12_data_i[0]_pad , \s12_data_i[10]_pad , \s12_data_i[11]_pad , \s12_data_i[12]_pad , \s12_data_i[13]_pad , \s12_data_i[14]_pad , \s12_data_i[15]_pad , \s12_data_i[16]_pad , \s12_data_i[17]_pad , \s12_data_i[18]_pad , \s12_data_i[19]_pad , \s12_data_i[1]_pad , \s12_data_i[20]_pad , \s12_data_i[21]_pad , \s12_data_i[22]_pad , \s12_data_i[23]_pad , \s12_data_i[24]_pad , \s12_data_i[25]_pad , \s12_data_i[26]_pad , \s12_data_i[27]_pad , \s12_data_i[28]_pad , \s12_data_i[29]_pad , \s12_data_i[2]_pad , \s12_data_i[30]_pad , \s12_data_i[31]_pad , \s12_data_i[3]_pad , \s12_data_i[4]_pad , \s12_data_i[5]_pad , \s12_data_i[6]_pad , \s12_data_i[7]_pad , \s12_data_i[8]_pad , \s12_data_i[9]_pad , \s12_err_i_pad , \s12_m0_cyc_r_reg/P0001 , \s12_m1_cyc_r_reg/P0001 , \s12_m2_cyc_r_reg/P0001 , \s12_m3_cyc_r_reg/P0001 , \s12_m4_cyc_r_reg/P0001 , \s12_m5_cyc_r_reg/P0001 , \s12_m6_cyc_r_reg/P0001 , \s12_m7_cyc_r_reg/P0001 , \s12_msel_arb0_state_reg[0]/NET0131 , \s12_msel_arb0_state_reg[1]/NET0131 , \s12_msel_arb0_state_reg[2]/NET0131 , \s12_msel_arb1_state_reg[0]/NET0131 , \s12_msel_arb1_state_reg[1]/NET0131 , \s12_msel_arb1_state_reg[2]/NET0131 , \s12_msel_arb2_state_reg[0]/NET0131 , \s12_msel_arb2_state_reg[1]/NET0131 , \s12_msel_arb2_state_reg[2]/NET0131 , \s12_msel_arb3_state_reg[0]/NET0131 , \s12_msel_arb3_state_reg[1]/NET0131 , \s12_msel_arb3_state_reg[2]/NET0131 , \s12_msel_pri_out_reg[0]/NET0131 , \s12_msel_pri_out_reg[1]/NET0131 , \s12_next_reg/P0001 , \s12_rty_i_pad , \s13_ack_i_pad , \s13_data_i[0]_pad , \s13_data_i[10]_pad , \s13_data_i[11]_pad , \s13_data_i[12]_pad , \s13_data_i[13]_pad , \s13_data_i[14]_pad , \s13_data_i[15]_pad , \s13_data_i[16]_pad , \s13_data_i[17]_pad , \s13_data_i[18]_pad , \s13_data_i[19]_pad , \s13_data_i[1]_pad , \s13_data_i[20]_pad , \s13_data_i[21]_pad , \s13_data_i[22]_pad , \s13_data_i[23]_pad , \s13_data_i[24]_pad , \s13_data_i[25]_pad , \s13_data_i[26]_pad , \s13_data_i[27]_pad , \s13_data_i[28]_pad , \s13_data_i[29]_pad , \s13_data_i[2]_pad , \s13_data_i[30]_pad , \s13_data_i[31]_pad , \s13_data_i[3]_pad , \s13_data_i[4]_pad , \s13_data_i[5]_pad , \s13_data_i[6]_pad , \s13_data_i[7]_pad , \s13_data_i[8]_pad , \s13_data_i[9]_pad , \s13_err_i_pad , \s13_m0_cyc_r_reg/P0001 , \s13_m1_cyc_r_reg/P0001 , \s13_m2_cyc_r_reg/P0001 , \s13_m3_cyc_r_reg/P0001 , \s13_m4_cyc_r_reg/P0001 , \s13_m5_cyc_r_reg/P0001 , \s13_m6_cyc_r_reg/P0001 , \s13_m7_cyc_r_reg/P0001 , \s13_msel_arb0_state_reg[0]/NET0131 , \s13_msel_arb0_state_reg[1]/NET0131 , \s13_msel_arb0_state_reg[2]/NET0131 , \s13_msel_arb1_state_reg[0]/NET0131 , \s13_msel_arb1_state_reg[1]/NET0131 , \s13_msel_arb1_state_reg[2]/NET0131 , \s13_msel_arb2_state_reg[0]/NET0131 , \s13_msel_arb2_state_reg[1]/NET0131 , \s13_msel_arb2_state_reg[2]/NET0131 , \s13_msel_arb3_state_reg[0]/NET0131 , \s13_msel_arb3_state_reg[1]/NET0131 , \s13_msel_arb3_state_reg[2]/NET0131 , \s13_msel_pri_out_reg[0]/NET0131 , \s13_msel_pri_out_reg[1]/NET0131 , \s13_next_reg/P0001 , \s13_rty_i_pad , \s14_ack_i_pad , \s14_data_i[0]_pad , \s14_data_i[10]_pad , \s14_data_i[11]_pad , \s14_data_i[12]_pad , \s14_data_i[13]_pad , \s14_data_i[14]_pad , \s14_data_i[15]_pad , \s14_data_i[16]_pad , \s14_data_i[17]_pad , \s14_data_i[18]_pad , \s14_data_i[19]_pad , \s14_data_i[1]_pad , \s14_data_i[20]_pad , \s14_data_i[21]_pad , \s14_data_i[22]_pad , \s14_data_i[23]_pad , \s14_data_i[24]_pad , \s14_data_i[25]_pad , \s14_data_i[26]_pad , \s14_data_i[27]_pad , \s14_data_i[28]_pad , \s14_data_i[29]_pad , \s14_data_i[2]_pad , \s14_data_i[30]_pad , \s14_data_i[31]_pad , \s14_data_i[3]_pad , \s14_data_i[4]_pad , \s14_data_i[5]_pad , \s14_data_i[6]_pad , \s14_data_i[7]_pad , \s14_data_i[8]_pad , \s14_data_i[9]_pad , \s14_err_i_pad , \s14_m0_cyc_r_reg/P0001 , \s14_m1_cyc_r_reg/P0001 , \s14_m2_cyc_r_reg/P0001 , \s14_m3_cyc_r_reg/P0001 , \s14_m4_cyc_r_reg/P0001 , \s14_m5_cyc_r_reg/P0001 , \s14_m6_cyc_r_reg/P0001 , \s14_m7_cyc_r_reg/P0001 , \s14_msel_arb0_state_reg[0]/NET0131 , \s14_msel_arb0_state_reg[1]/NET0131 , \s14_msel_arb0_state_reg[2]/NET0131 , \s14_msel_arb1_state_reg[0]/NET0131 , \s14_msel_arb1_state_reg[1]/NET0131 , \s14_msel_arb1_state_reg[2]/NET0131 , \s14_msel_arb2_state_reg[0]/NET0131 , \s14_msel_arb2_state_reg[1]/NET0131 , \s14_msel_arb2_state_reg[2]/NET0131 , \s14_msel_arb3_state_reg[0]/NET0131 , \s14_msel_arb3_state_reg[1]/NET0131 , \s14_msel_arb3_state_reg[2]/NET0131 , \s14_msel_pri_out_reg[0]/NET0131 , \s14_msel_pri_out_reg[1]/NET0131 , \s14_next_reg/P0001 , \s14_rty_i_pad , \s15_ack_i_pad , \s15_data_i[0]_pad , \s15_data_i[10]_pad , \s15_data_i[11]_pad , \s15_data_i[12]_pad , \s15_data_i[13]_pad , \s15_data_i[14]_pad , \s15_data_i[15]_pad , \s15_data_i[16]_pad , \s15_data_i[17]_pad , \s15_data_i[18]_pad , \s15_data_i[19]_pad , \s15_data_i[1]_pad , \s15_data_i[20]_pad , \s15_data_i[21]_pad , \s15_data_i[22]_pad , \s15_data_i[23]_pad , \s15_data_i[24]_pad , \s15_data_i[25]_pad , \s15_data_i[26]_pad , \s15_data_i[27]_pad , \s15_data_i[28]_pad , \s15_data_i[29]_pad , \s15_data_i[2]_pad , \s15_data_i[30]_pad , \s15_data_i[31]_pad , \s15_data_i[3]_pad , \s15_data_i[4]_pad , \s15_data_i[5]_pad , \s15_data_i[6]_pad , \s15_data_i[7]_pad , \s15_data_i[8]_pad , \s15_data_i[9]_pad , \s15_err_i_pad , \s15_m0_cyc_r_reg/P0001 , \s15_m1_cyc_r_reg/P0001 , \s15_m2_cyc_r_reg/P0001 , \s15_m3_cyc_r_reg/P0001 , \s15_m4_cyc_r_reg/P0001 , \s15_m5_cyc_r_reg/P0001 , \s15_m6_cyc_r_reg/P0001 , \s15_m7_cyc_r_reg/P0001 , \s15_msel_arb0_state_reg[0]/NET0131 , \s15_msel_arb0_state_reg[1]/NET0131 , \s15_msel_arb0_state_reg[2]/NET0131 , \s15_msel_arb1_state_reg[0]/NET0131 , \s15_msel_arb1_state_reg[1]/NET0131 , \s15_msel_arb1_state_reg[2]/NET0131 , \s15_msel_arb2_state_reg[0]/NET0131 , \s15_msel_arb2_state_reg[1]/NET0131 , \s15_msel_arb2_state_reg[2]/NET0131 , \s15_msel_arb3_state_reg[0]/NET0131 , \s15_msel_arb3_state_reg[1]/NET0131 , \s15_msel_arb3_state_reg[2]/NET0131 , \s15_msel_pri_out_reg[0]/NET0131 , \s15_msel_pri_out_reg[1]/NET0131 , \s15_next_reg/P0001 , \s15_rty_i_pad , \s1_ack_i_pad , \s1_data_i[0]_pad , \s1_data_i[10]_pad , \s1_data_i[11]_pad , \s1_data_i[12]_pad , \s1_data_i[13]_pad , \s1_data_i[14]_pad , \s1_data_i[15]_pad , \s1_data_i[16]_pad , \s1_data_i[17]_pad , \s1_data_i[18]_pad , \s1_data_i[19]_pad , \s1_data_i[1]_pad , \s1_data_i[20]_pad , \s1_data_i[21]_pad , \s1_data_i[22]_pad , \s1_data_i[23]_pad , \s1_data_i[24]_pad , \s1_data_i[25]_pad , \s1_data_i[26]_pad , \s1_data_i[27]_pad , \s1_data_i[28]_pad , \s1_data_i[29]_pad , \s1_data_i[2]_pad , \s1_data_i[30]_pad , \s1_data_i[31]_pad , \s1_data_i[3]_pad , \s1_data_i[4]_pad , \s1_data_i[5]_pad , \s1_data_i[6]_pad , \s1_data_i[7]_pad , \s1_data_i[8]_pad , \s1_data_i[9]_pad , \s1_err_i_pad , \s1_m0_cyc_r_reg/P0001 , \s1_m1_cyc_r_reg/P0001 , \s1_m2_cyc_r_reg/P0001 , \s1_m3_cyc_r_reg/P0001 , \s1_m4_cyc_r_reg/P0001 , \s1_m5_cyc_r_reg/P0001 , \s1_m6_cyc_r_reg/P0001 , \s1_m7_cyc_r_reg/P0001 , \s1_msel_arb0_state_reg[0]/NET0131 , \s1_msel_arb0_state_reg[1]/NET0131 , \s1_msel_arb0_state_reg[2]/NET0131 , \s1_msel_arb1_state_reg[0]/NET0131 , \s1_msel_arb1_state_reg[1]/NET0131 , \s1_msel_arb1_state_reg[2]/NET0131 , \s1_msel_arb2_state_reg[0]/NET0131 , \s1_msel_arb2_state_reg[1]/NET0131 , \s1_msel_arb2_state_reg[2]/NET0131 , \s1_msel_arb3_state_reg[0]/NET0131 , \s1_msel_arb3_state_reg[1]/NET0131 , \s1_msel_arb3_state_reg[2]/NET0131 , \s1_msel_pri_out_reg[0]/NET0131 , \s1_msel_pri_out_reg[1]/NET0131 , \s1_next_reg/P0001 , \s1_rty_i_pad , \s2_ack_i_pad , \s2_data_i[0]_pad , \s2_data_i[10]_pad , \s2_data_i[11]_pad , \s2_data_i[12]_pad , \s2_data_i[13]_pad , \s2_data_i[14]_pad , \s2_data_i[15]_pad , \s2_data_i[16]_pad , \s2_data_i[17]_pad , \s2_data_i[18]_pad , \s2_data_i[19]_pad , \s2_data_i[1]_pad , \s2_data_i[20]_pad , \s2_data_i[21]_pad , \s2_data_i[22]_pad , \s2_data_i[23]_pad , \s2_data_i[24]_pad , \s2_data_i[25]_pad , \s2_data_i[26]_pad , \s2_data_i[27]_pad , \s2_data_i[28]_pad , \s2_data_i[29]_pad , \s2_data_i[2]_pad , \s2_data_i[30]_pad , \s2_data_i[31]_pad , \s2_data_i[3]_pad , \s2_data_i[4]_pad , \s2_data_i[5]_pad , \s2_data_i[6]_pad , \s2_data_i[7]_pad , \s2_data_i[8]_pad , \s2_data_i[9]_pad , \s2_err_i_pad , \s2_m0_cyc_r_reg/P0001 , \s2_m1_cyc_r_reg/P0001 , \s2_m2_cyc_r_reg/P0001 , \s2_m3_cyc_r_reg/P0001 , \s2_m4_cyc_r_reg/P0001 , \s2_m5_cyc_r_reg/P0001 , \s2_m6_cyc_r_reg/P0001 , \s2_m7_cyc_r_reg/P0001 , \s2_msel_arb0_state_reg[0]/NET0131 , \s2_msel_arb0_state_reg[1]/NET0131 , \s2_msel_arb0_state_reg[2]/NET0131 , \s2_msel_arb1_state_reg[0]/NET0131 , \s2_msel_arb1_state_reg[1]/NET0131 , \s2_msel_arb1_state_reg[2]/NET0131 , \s2_msel_arb2_state_reg[0]/NET0131 , \s2_msel_arb2_state_reg[1]/NET0131 , \s2_msel_arb2_state_reg[2]/NET0131 , \s2_msel_arb3_state_reg[0]/NET0131 , \s2_msel_arb3_state_reg[1]/NET0131 , \s2_msel_arb3_state_reg[2]/NET0131 , \s2_msel_pri_out_reg[0]/NET0131 , \s2_msel_pri_out_reg[1]/NET0131 , \s2_next_reg/P0001 , \s2_rty_i_pad , \s3_ack_i_pad , \s3_data_i[0]_pad , \s3_data_i[10]_pad , \s3_data_i[11]_pad , \s3_data_i[12]_pad , \s3_data_i[13]_pad , \s3_data_i[14]_pad , \s3_data_i[15]_pad , \s3_data_i[16]_pad , \s3_data_i[17]_pad , \s3_data_i[18]_pad , \s3_data_i[19]_pad , \s3_data_i[1]_pad , \s3_data_i[20]_pad , \s3_data_i[21]_pad , \s3_data_i[22]_pad , \s3_data_i[23]_pad , \s3_data_i[24]_pad , \s3_data_i[25]_pad , \s3_data_i[26]_pad , \s3_data_i[27]_pad , \s3_data_i[28]_pad , \s3_data_i[29]_pad , \s3_data_i[2]_pad , \s3_data_i[30]_pad , \s3_data_i[31]_pad , \s3_data_i[3]_pad , \s3_data_i[4]_pad , \s3_data_i[5]_pad , \s3_data_i[6]_pad , \s3_data_i[7]_pad , \s3_data_i[8]_pad , \s3_data_i[9]_pad , \s3_err_i_pad , \s3_m0_cyc_r_reg/P0001 , \s3_m1_cyc_r_reg/P0001 , \s3_m2_cyc_r_reg/P0001 , \s3_m3_cyc_r_reg/P0001 , \s3_m4_cyc_r_reg/P0001 , \s3_m5_cyc_r_reg/P0001 , \s3_m6_cyc_r_reg/P0001 , \s3_m7_cyc_r_reg/P0001 , \s3_msel_arb0_state_reg[0]/NET0131 , \s3_msel_arb0_state_reg[1]/NET0131 , \s3_msel_arb0_state_reg[2]/NET0131 , \s3_msel_arb1_state_reg[0]/NET0131 , \s3_msel_arb1_state_reg[1]/NET0131 , \s3_msel_arb1_state_reg[2]/NET0131 , \s3_msel_arb2_state_reg[0]/NET0131 , \s3_msel_arb2_state_reg[1]/NET0131 , \s3_msel_arb2_state_reg[2]/NET0131 , \s3_msel_arb3_state_reg[0]/NET0131 , \s3_msel_arb3_state_reg[1]/NET0131 , \s3_msel_arb3_state_reg[2]/NET0131 , \s3_msel_pri_out_reg[0]/NET0131 , \s3_msel_pri_out_reg[1]/NET0131 , \s3_next_reg/P0001 , \s3_rty_i_pad , \s4_ack_i_pad , \s4_data_i[0]_pad , \s4_data_i[10]_pad , \s4_data_i[11]_pad , \s4_data_i[12]_pad , \s4_data_i[13]_pad , \s4_data_i[14]_pad , \s4_data_i[15]_pad , \s4_data_i[16]_pad , \s4_data_i[17]_pad , \s4_data_i[18]_pad , \s4_data_i[19]_pad , \s4_data_i[1]_pad , \s4_data_i[20]_pad , \s4_data_i[21]_pad , \s4_data_i[22]_pad , \s4_data_i[23]_pad , \s4_data_i[24]_pad , \s4_data_i[25]_pad , \s4_data_i[26]_pad , \s4_data_i[27]_pad , \s4_data_i[28]_pad , \s4_data_i[29]_pad , \s4_data_i[2]_pad , \s4_data_i[30]_pad , \s4_data_i[31]_pad , \s4_data_i[3]_pad , \s4_data_i[4]_pad , \s4_data_i[5]_pad , \s4_data_i[6]_pad , \s4_data_i[7]_pad , \s4_data_i[8]_pad , \s4_data_i[9]_pad , \s4_err_i_pad , \s4_m0_cyc_r_reg/P0001 , \s4_m1_cyc_r_reg/P0001 , \s4_m2_cyc_r_reg/P0001 , \s4_m3_cyc_r_reg/P0001 , \s4_m4_cyc_r_reg/P0001 , \s4_m5_cyc_r_reg/P0001 , \s4_m6_cyc_r_reg/P0001 , \s4_m7_cyc_r_reg/P0001 , \s4_msel_arb0_state_reg[0]/NET0131 , \s4_msel_arb0_state_reg[1]/NET0131 , \s4_msel_arb0_state_reg[2]/NET0131 , \s4_msel_arb1_state_reg[0]/NET0131 , \s4_msel_arb1_state_reg[1]/NET0131 , \s4_msel_arb1_state_reg[2]/NET0131 , \s4_msel_arb2_state_reg[0]/NET0131 , \s4_msel_arb2_state_reg[1]/NET0131 , \s4_msel_arb2_state_reg[2]/NET0131 , \s4_msel_arb3_state_reg[0]/NET0131 , \s4_msel_arb3_state_reg[1]/NET0131 , \s4_msel_arb3_state_reg[2]/NET0131 , \s4_msel_pri_out_reg[0]/NET0131 , \s4_msel_pri_out_reg[1]/NET0131 , \s4_next_reg/P0001 , \s4_rty_i_pad , \s5_ack_i_pad , \s5_data_i[0]_pad , \s5_data_i[10]_pad , \s5_data_i[11]_pad , \s5_data_i[12]_pad , \s5_data_i[13]_pad , \s5_data_i[14]_pad , \s5_data_i[15]_pad , \s5_data_i[16]_pad , \s5_data_i[17]_pad , \s5_data_i[18]_pad , \s5_data_i[19]_pad , \s5_data_i[1]_pad , \s5_data_i[20]_pad , \s5_data_i[21]_pad , \s5_data_i[22]_pad , \s5_data_i[23]_pad , \s5_data_i[24]_pad , \s5_data_i[25]_pad , \s5_data_i[26]_pad , \s5_data_i[27]_pad , \s5_data_i[28]_pad , \s5_data_i[29]_pad , \s5_data_i[2]_pad , \s5_data_i[30]_pad , \s5_data_i[31]_pad , \s5_data_i[3]_pad , \s5_data_i[4]_pad , \s5_data_i[5]_pad , \s5_data_i[6]_pad , \s5_data_i[7]_pad , \s5_data_i[8]_pad , \s5_data_i[9]_pad , \s5_err_i_pad , \s5_m0_cyc_r_reg/P0001 , \s5_m1_cyc_r_reg/P0001 , \s5_m2_cyc_r_reg/P0001 , \s5_m3_cyc_r_reg/P0001 , \s5_m4_cyc_r_reg/P0001 , \s5_m5_cyc_r_reg/P0001 , \s5_m6_cyc_r_reg/P0001 , \s5_m7_cyc_r_reg/P0001 , \s5_msel_arb0_state_reg[0]/NET0131 , \s5_msel_arb0_state_reg[1]/NET0131 , \s5_msel_arb0_state_reg[2]/NET0131 , \s5_msel_arb1_state_reg[0]/NET0131 , \s5_msel_arb1_state_reg[1]/NET0131 , \s5_msel_arb1_state_reg[2]/NET0131 , \s5_msel_arb2_state_reg[0]/NET0131 , \s5_msel_arb2_state_reg[1]/NET0131 , \s5_msel_arb2_state_reg[2]/NET0131 , \s5_msel_arb3_state_reg[0]/NET0131 , \s5_msel_arb3_state_reg[1]/NET0131 , \s5_msel_arb3_state_reg[2]/NET0131 , \s5_msel_pri_out_reg[0]/NET0131 , \s5_msel_pri_out_reg[1]/NET0131 , \s5_next_reg/P0001 , \s5_rty_i_pad , \s6_ack_i_pad , \s6_data_i[0]_pad , \s6_data_i[10]_pad , \s6_data_i[11]_pad , \s6_data_i[12]_pad , \s6_data_i[13]_pad , \s6_data_i[14]_pad , \s6_data_i[15]_pad , \s6_data_i[16]_pad , \s6_data_i[17]_pad , \s6_data_i[18]_pad , \s6_data_i[19]_pad , \s6_data_i[1]_pad , \s6_data_i[20]_pad , \s6_data_i[21]_pad , \s6_data_i[22]_pad , \s6_data_i[23]_pad , \s6_data_i[24]_pad , \s6_data_i[25]_pad , \s6_data_i[26]_pad , \s6_data_i[27]_pad , \s6_data_i[28]_pad , \s6_data_i[29]_pad , \s6_data_i[2]_pad , \s6_data_i[30]_pad , \s6_data_i[31]_pad , \s6_data_i[3]_pad , \s6_data_i[4]_pad , \s6_data_i[5]_pad , \s6_data_i[6]_pad , \s6_data_i[7]_pad , \s6_data_i[8]_pad , \s6_data_i[9]_pad , \s6_err_i_pad , \s6_m0_cyc_r_reg/P0001 , \s6_m1_cyc_r_reg/P0001 , \s6_m2_cyc_r_reg/P0001 , \s6_m3_cyc_r_reg/P0001 , \s6_m4_cyc_r_reg/P0001 , \s6_m5_cyc_r_reg/P0001 , \s6_m6_cyc_r_reg/P0001 , \s6_m7_cyc_r_reg/P0001 , \s6_msel_arb0_state_reg[0]/NET0131 , \s6_msel_arb0_state_reg[1]/NET0131 , \s6_msel_arb0_state_reg[2]/NET0131 , \s6_msel_arb1_state_reg[0]/NET0131 , \s6_msel_arb1_state_reg[1]/NET0131 , \s6_msel_arb1_state_reg[2]/NET0131 , \s6_msel_arb2_state_reg[0]/NET0131 , \s6_msel_arb2_state_reg[1]/NET0131 , \s6_msel_arb2_state_reg[2]/NET0131 , \s6_msel_arb3_state_reg[0]/NET0131 , \s6_msel_arb3_state_reg[1]/NET0131 , \s6_msel_arb3_state_reg[2]/NET0131 , \s6_msel_pri_out_reg[0]/NET0131 , \s6_msel_pri_out_reg[1]/NET0131 , \s6_next_reg/P0001 , \s6_rty_i_pad , \s7_ack_i_pad , \s7_data_i[0]_pad , \s7_data_i[10]_pad , \s7_data_i[11]_pad , \s7_data_i[12]_pad , \s7_data_i[13]_pad , \s7_data_i[14]_pad , \s7_data_i[15]_pad , \s7_data_i[16]_pad , \s7_data_i[17]_pad , \s7_data_i[18]_pad , \s7_data_i[19]_pad , \s7_data_i[1]_pad , \s7_data_i[20]_pad , \s7_data_i[21]_pad , \s7_data_i[22]_pad , \s7_data_i[23]_pad , \s7_data_i[24]_pad , \s7_data_i[25]_pad , \s7_data_i[26]_pad , \s7_data_i[27]_pad , \s7_data_i[28]_pad , \s7_data_i[29]_pad , \s7_data_i[2]_pad , \s7_data_i[30]_pad , \s7_data_i[31]_pad , \s7_data_i[3]_pad , \s7_data_i[4]_pad , \s7_data_i[5]_pad , \s7_data_i[6]_pad , \s7_data_i[7]_pad , \s7_data_i[8]_pad , \s7_data_i[9]_pad , \s7_err_i_pad , \s7_m0_cyc_r_reg/P0001 , \s7_m1_cyc_r_reg/P0001 , \s7_m2_cyc_r_reg/P0001 , \s7_m3_cyc_r_reg/P0001 , \s7_m4_cyc_r_reg/P0001 , \s7_m5_cyc_r_reg/P0001 , \s7_m6_cyc_r_reg/P0001 , \s7_m7_cyc_r_reg/P0001 , \s7_msel_arb0_state_reg[0]/NET0131 , \s7_msel_arb0_state_reg[1]/NET0131 , \s7_msel_arb0_state_reg[2]/NET0131 , \s7_msel_arb1_state_reg[0]/NET0131 , \s7_msel_arb1_state_reg[1]/NET0131 , \s7_msel_arb1_state_reg[2]/NET0131 , \s7_msel_arb2_state_reg[0]/NET0131 , \s7_msel_arb2_state_reg[1]/NET0131 , \s7_msel_arb2_state_reg[2]/NET0131 , \s7_msel_arb3_state_reg[0]/NET0131 , \s7_msel_arb3_state_reg[1]/NET0131 , \s7_msel_arb3_state_reg[2]/NET0131 , \s7_msel_pri_out_reg[0]/NET0131 , \s7_msel_pri_out_reg[1]/NET0131 , \s7_next_reg/P0001 , \s7_rty_i_pad , \s8_ack_i_pad , \s8_data_i[0]_pad , \s8_data_i[10]_pad , \s8_data_i[11]_pad , \s8_data_i[12]_pad , \s8_data_i[13]_pad , \s8_data_i[14]_pad , \s8_data_i[15]_pad , \s8_data_i[16]_pad , \s8_data_i[17]_pad , \s8_data_i[18]_pad , \s8_data_i[19]_pad , \s8_data_i[1]_pad , \s8_data_i[20]_pad , \s8_data_i[21]_pad , \s8_data_i[22]_pad , \s8_data_i[23]_pad , \s8_data_i[24]_pad , \s8_data_i[25]_pad , \s8_data_i[26]_pad , \s8_data_i[27]_pad , \s8_data_i[28]_pad , \s8_data_i[29]_pad , \s8_data_i[2]_pad , \s8_data_i[30]_pad , \s8_data_i[31]_pad , \s8_data_i[3]_pad , \s8_data_i[4]_pad , \s8_data_i[5]_pad , \s8_data_i[6]_pad , \s8_data_i[7]_pad , \s8_data_i[8]_pad , \s8_data_i[9]_pad , \s8_err_i_pad , \s8_m0_cyc_r_reg/P0001 , \s8_m1_cyc_r_reg/P0001 , \s8_m2_cyc_r_reg/P0001 , \s8_m3_cyc_r_reg/P0001 , \s8_m4_cyc_r_reg/P0001 , \s8_m5_cyc_r_reg/P0001 , \s8_m6_cyc_r_reg/P0001 , \s8_m7_cyc_r_reg/P0001 , \s8_msel_arb0_state_reg[0]/NET0131 , \s8_msel_arb0_state_reg[1]/NET0131 , \s8_msel_arb0_state_reg[2]/NET0131 , \s8_msel_arb1_state_reg[0]/NET0131 , \s8_msel_arb1_state_reg[1]/NET0131 , \s8_msel_arb1_state_reg[2]/NET0131 , \s8_msel_arb2_state_reg[0]/NET0131 , \s8_msel_arb2_state_reg[1]/NET0131 , \s8_msel_arb2_state_reg[2]/NET0131 , \s8_msel_arb3_state_reg[0]/NET0131 , \s8_msel_arb3_state_reg[1]/NET0131 , \s8_msel_arb3_state_reg[2]/NET0131 , \s8_msel_pri_out_reg[0]/NET0131 , \s8_msel_pri_out_reg[1]/NET0131 , \s8_next_reg/P0001 , \s8_rty_i_pad , \s9_ack_i_pad , \s9_data_i[0]_pad , \s9_data_i[10]_pad , \s9_data_i[11]_pad , \s9_data_i[12]_pad , \s9_data_i[13]_pad , \s9_data_i[14]_pad , \s9_data_i[15]_pad , \s9_data_i[16]_pad , \s9_data_i[17]_pad , \s9_data_i[18]_pad , \s9_data_i[19]_pad , \s9_data_i[1]_pad , \s9_data_i[20]_pad , \s9_data_i[21]_pad , \s9_data_i[22]_pad , \s9_data_i[23]_pad , \s9_data_i[24]_pad , \s9_data_i[25]_pad , \s9_data_i[26]_pad , \s9_data_i[27]_pad , \s9_data_i[28]_pad , \s9_data_i[29]_pad , \s9_data_i[2]_pad , \s9_data_i[30]_pad , \s9_data_i[31]_pad , \s9_data_i[3]_pad , \s9_data_i[4]_pad , \s9_data_i[5]_pad , \s9_data_i[6]_pad , \s9_data_i[7]_pad , \s9_data_i[8]_pad , \s9_data_i[9]_pad , \s9_err_i_pad , \s9_m0_cyc_r_reg/P0001 , \s9_m1_cyc_r_reg/P0001 , \s9_m2_cyc_r_reg/P0001 , \s9_m3_cyc_r_reg/P0001 , \s9_m4_cyc_r_reg/P0001 , \s9_m5_cyc_r_reg/P0001 , \s9_m6_cyc_r_reg/P0001 , \s9_m7_cyc_r_reg/P0001 , \s9_msel_arb0_state_reg[0]/NET0131 , \s9_msel_arb0_state_reg[1]/NET0131 , \s9_msel_arb0_state_reg[2]/NET0131 , \s9_msel_arb1_state_reg[0]/NET0131 , \s9_msel_arb1_state_reg[1]/NET0131 , \s9_msel_arb1_state_reg[2]/NET0131 , \s9_msel_arb2_state_reg[0]/NET0131 , \s9_msel_arb2_state_reg[1]/NET0131 , \s9_msel_arb2_state_reg[2]/NET0131 , \s9_msel_arb3_state_reg[0]/NET0131 , \s9_msel_arb3_state_reg[1]/NET0131 , \s9_msel_arb3_state_reg[2]/NET0131 , \s9_msel_pri_out_reg[0]/NET0131 , \s9_msel_pri_out_reg[1]/NET0131 , \s9_next_reg/P0001 , \s9_rty_i_pad , \_al_n0 , \_al_n1 , \g106655/_1_ , \g106703/_1_ , \g69412/_0_ , \g69413/_0_ , \g69417/_1_ , \g69418/_0_ , \g69420/_1_ , \g69421/_0_ , \g69423/_1_ , \g69424/_0_ , \g69426/_1_ , \g69428/_1_ , \g69430/_1_ , \g69432/_1_ , \g69434/_1_ , \g69436/_1_ , \g69438/_1_ , \g69757/_2_ , \g69758/_2_ , \g69759/_2_ , \g69760/_2_ , \g69761/_0_ , \g69762/_2_ , \g69763/_2_ , \g69764/_2_ , \g69765/_2_ , \g69766/_2_ , \g69767/_0_ , \g69768/_0_ , \g69769/_0_ , \g69770/_0_ , \g69771/_0_ , \g69772/_0_ , \g70206/_0_ , \g70392/_0_ , \g70393/_0_ , \g70394/_0_ , \g70395/_0_ , \g70396/_0_ , \g70397/_0_ , \g70398/_0_ , \g70399/_0_ , \g70400/_0_ , \g70401/_0_ , \g70402/_0_ , \g70403/_0_ , \g70404/_0_ , \g70405/_0_ , \g70406/_0_ , \g70407/_0_ , \g70408/_0_ , \g70409/_0_ , \g70410/_0_ , \g70411/_0_ , \g70412/_0_ , \g70413/_0_ , \g70414/_0_ , \g70415/_0_ , \g70416/_0_ , \g70417/_0_ , \g70418/_0_ , \g70419/_0_ , \g70420/_0_ , \g70421/_0_ , \g70422/_0_ , \g70423/_0_ , \g70424/_0_ , \g70425/_0_ , \g70426/_0_ , \g70427/_0_ , \g70428/_0_ , \g70429/_0_ , \g70430/_0_ , \g70431/_0_ , \g70432/_0_ , \g70433/_0_ , \g70434/_0_ , \g70435/_0_ , \g70436/_0_ , \g70437/_0_ , \g70438/_0_ , \g70439/_0_ , \g70440/_0_ , \g70441/_0_ , \g70442/_0_ , \g70443/_0_ , \g70444/_0_ , \g70445/_0_ , \g70446/_0_ , \g70447/_0_ , \g70448/_0_ , \g70449/_0_ , \g70450/_0_ , \g70451/_0_ , \g70452/_0_ , \g70453/_0_ , \g70454/_0_ , \g70455/_0_ , \g70456/_0_ , \g70457/_0_ , \g70458/_0_ , \g70459/_0_ , \g70460/_0_ , \g70461/_0_ , \g70462/_0_ , \g70463/_0_ , \g70464/_0_ , \g70465/_0_ , \g70466/_0_ , \g70467/_0_ , \g70468/_0_ , \g70469/_0_ , \g70470/_0_ , \g70471/_0_ , \g70472/_0_ , \g70473/_0_ , \g70474/_0_ , \g70475/_0_ , \g70476/_0_ , \g70477/_0_ , \g70478/_0_ , \g70479/_0_ , \g70480/_0_ , \g70481/_0_ , \g70482/_0_ , \g70483/_0_ , \g70484/_0_ , \g70485/_0_ , \g70486/_0_ , \g70487/_0_ , \g70488/_0_ , \g70489/_0_ , \g70490/_0_ , \g70491/_0_ , \g70492/_0_ , \g70493/_0_ , \g70494/_0_ , \g70495/_0_ , \g70496/_0_ , \g70497/_0_ , \g70498/_0_ , \g70499/_0_ , \g70500/_0_ , \g70501/_0_ , \g70502/_0_ , \g70503/_0_ , \g70504/_0_ , \g70505/_0_ , \g70506/_0_ , \g70507/_0_ , \g70508/_0_ , \g70509/_0_ , \g70510/_0_ , \g70511/_0_ , \g70513/_0_ , \g70515/_0_ , \g70516/_0_ , \g70517/_0_ , \g70518/_0_ , \g70519/_0_ , \g70521/_0_ , \g70522/_0_ , \g70524/_0_ , \g70557/_0_ , \g70559/_0_ , \g70560/_0_ , \g70561/_0_ , \g70562/_0_ , \g70563/_0_ , \g70564/_0_ , \g70565/_0_ , \g70566/_0_ , \g70567/_0_ , \g70568/_0_ , \g70569/_0_ , \g70570/_0_ , \g70571/_0_ , \g70572/_0_ , \g70573/_0_ , \g70574/_0_ , \g70575/_0_ , \g70576/_0_ , \g70577/_0_ , \g70578/_0_ , \g70579/_0_ , \g70580/_0_ , \g70581/_0_ , \g70582/_0_ , \g70583/_0_ , \g70584/_0_ , \g70585/_0_ , \g70586/_0_ , \g70587/_0_ , \g70588/_0_ , \g70589/_0_ , \g70590/_0_ , \g70591/_0_ , \g70592/_0_ , \g70593/_0_ , \g70594/_0_ , \g70595/_0_ , \g70596/_0_ , \g70597/_0_ , \g70598/_0_ , \g70599/_0_ , \g70600/_0_ , \g70601/_0_ , \g70602/_0_ , \g70603/_0_ , \g70604/_0_ , \g70605/_0_ , \g70606/_0_ , \g70607/_0_ , \g70608/_0_ , \g70609/_0_ , \g70610/_0_ , \g70611/_0_ , \g70612/_0_ , \g70613/_0_ , \g70614/_0_ , \g70615/_0_ , \g70616/_0_ , \g70617/_0_ , \g70618/_0_ , \g70619/_0_ , \g70620/_0_ , \g70621/_0_ , \g70622/_0_ , \g70623/_0_ , \g70624/_0_ , \g70625/_0_ , \g70626/_0_ , \g70627/_0_ , \g70628/_0_ , \g70629/_0_ , \g70630/_0_ , \g70631/_0_ , \g70632/_0_ , \g70633/_0_ , \g70634/_0_ , \g70635/_0_ , \g70636/_0_ , \g70637/_0_ , \g70638/_0_ , \g70639/_0_ , \g70640/_0_ , \g70641/_0_ , \g70642/_0_ , \g70643/_0_ , \g70644/_0_ , \g70645/_0_ , \g70646/_0_ , \g70647/_0_ , \g70648/_0_ , \g70649/_0_ , \g70650/_0_ , \g70651/_0_ , \g70652/_0_ , \g70653/_0_ , \g70654/_0_ , \g70655/_0_ , \g70656/_0_ , \g70657/_0_ , \g70658/_0_ , \g70659/_0_ , \g70660/_0_ , \g70661/_0_ , \g70662/_0_ , \g70663/_0_ , \g70664/_0_ , \g70665/_0_ , \g70666/_0_ , \g70667/_0_ , \g70668/_0_ , \g70669/_0_ , \g70670/_0_ , \g70671/_0_ , \g70672/_0_ , \g70673/_0_ , \g70674/_0_ , \g70675/_0_ , \g70676/_0_ , \g70677/_0_ , \g70678/_0_ , \g70679/_0_ , \g70680/_0_ , \g70681/_0_ , \g70682/_0_ , \g70683/_0_ , \g70684/_0_ , \g70685/_0_ , \g70686/_0_ , \g70687/_0_ , \g70688/_0_ , \g70689/_0_ , \g70690/_0_ , \g70691/_0_ , \g70692/_0_ , \g70693/_0_ , \g70694/_0_ , \g70695/_0_ , \g70696/_0_ , \g70697/_0_ , \g70698/_0_ , \g70699/_0_ , \g70700/_0_ , \g70701/_0_ , \g70702/_0_ , \g70703/_0_ , \g70704/_0_ , \g70705/_0_ , \g70706/_0_ , \g70707/_0_ , \g70708/_0_ , \g70709/_0_ , \g70710/_0_ , \g70711/_0_ , \g70712/_0_ , \g70713/_0_ , \g70714/_0_ , \g70715/_0_ , \g70716/_0_ , \g70717/_0_ , \g70718/_0_ , \g70719/_0_ , \g70720/_0_ , \g70721/_0_ , \g70722/_0_ , \g70723/_0_ , \g70724/_0_ , \g70725/_0_ , \g70726/_0_ , \g70727/_0_ , \g70728/_0_ , \g70729/_0_ , \g70730/_0_ , \g70731/_0_ , \g70732/_0_ , \g70733/_0_ , \g70734/_0_ , \g70735/_0_ , \g70736/_0_ , \g70737/_0_ , \g70738/_0_ , \g70739/_0_ , \g70740/_0_ , \g70741/_0_ , \g70742/_0_ , \g70743/_0_ , \g70744/_0_ , \g70745/_0_ , \g70746/_0_ , \g70747/_0_ , \g70748/_0_ , \g70749/_0_ , \g70750/_0_ , \g70751/_0_ , \g70752/_0_ , \g70753/_0_ , \g70754/_0_ , \g70755/_0_ , \g70756/_0_ , \g70757/_0_ , \g70758/_0_ , \g70759/_0_ , \g70760/_0_ , \g70761/_0_ , \g70762/_0_ , \g70763/_0_ , \g70764/_0_ , \g70765/_0_ , \g70766/_0_ , \g70767/_0_ , \g70768/_0_ , \g70769/_0_ , \g70770/_0_ , \g70771/_0_ , \g70772/_0_ , \g70773/_0_ , \g70774/_0_ , \g70775/_0_ , \g70776/_0_ , \g70777/_0_ , \g70778/_0_ , \g70779/_0_ , \g70780/_0_ , \g70781/_0_ , \g70782/_0_ , \g70783/_0_ , \g70784/_0_ , \g70785/_0_ , \g70786/_0_ , \g70787/_0_ , \g70788/_0_ , \g70789/_0_ , \g70790/_0_ , \g70791/_0_ , \g70792/_0_ , \g70793/_0_ , \g70794/_0_ , \g70795/_0_ , \g70796/_0_ , \g70797/_0_ , \g70798/_0_ , \g70799/_0_ , \g70800/_0_ , \g70801/_0_ , \g70802/_0_ , \g70803/_0_ , \g70804/_0_ , \g70805/_0_ , \g70806/_0_ , \g70807/_0_ , \g70808/_0_ , \g70809/_0_ , \g70810/_0_ , \g70811/_0_ , \g70812/_0_ , \g70813/_0_ , \g70814/_0_ , \g70815/_0_ , \g70816/_0_ , \g70817/_0_ , \g70818/_0_ , \g70819/_0_ , \g70820/_0_ , \g70821/_0_ , \g70822/_0_ , \g70823/_0_ , \g70824/_0_ , \g70825/_0_ , \g70826/_0_ , \g70827/_0_ , \g70828/_0_ , \g70829/_0_ , \g70830/_0_ , \g70831/_0_ , \g70832/_0_ , \g70833/_0_ , \g70834/_0_ , \g70835/_0_ , \g70836/_0_ , \g70837/_0_ , \g70838/_0_ , \g70839/_0_ , \g70840/_0_ , \g70841/_0_ , \g70842/_0_ , \g70843/_0_ , \g70844/_0_ , \g70845/_0_ , \g70846/_0_ , \g70847/_0_ , \g70848/_0_ , \g70849/_0_ , \g70850/_0_ , \g70851/_0_ , \g70852/_0_ , \g70853/_0_ , \g70854/_0_ , \g70855/_0_ , \g70856/_0_ , \g70857/_0_ , \g70858/_0_ , \g70859/_0_ , \g70860/_0_ , \g70861/_0_ , \g71404/_0_ , \g71407/_0_ , \g72631/_0_ , \g72631/_1_ , \g72633/_0_ , \g72642/_0_ , \g72649/_0_ , \g72649/_1_ , \g72652/_0_ , \g72660/_0_ , \g72666/_0_ , \g72666/_1_ , \g72671/_0_ , \g72681/_0_ , \g72681/_1_ , \g72689/_0_ , \g72696/_0_ , \g72696/_1_ , \g72698/_0_ , \g72707/_0_ , \g72715/_0_ , \g72715/_1_ , \g72718/_0_ , \g72726/_0_ , \g72732/_0_ , \g72732/_1_ , \g72736/_0_ , \g72743/_0_ , \g72745/_0_ , \g72745/_1_ , \g72752/_0_ , \g72752/_1_ , \g72756/_0_ , \g72763/_0_ , \g72763/_1_ , \g72765/_0_ , \g72767/_0_ , \g72767/_1_ , \g72769/_0_ , \g72769/_1_ , \g72772/_0_ , \g72772/_1_ , \g72774/_0_ , \g72774/_1_ , \g72790/_0_ , \g72790/_1_ , \g72797/_0_ , \g73807/_0_ , \g73820/_0_ , \g73832/_0_ , \g73844/_0_ , \g73856/_0_ , \g73871/_0_ , \g73883/_0_ , \g73895/_0_ , \g73905/_3_ , \g73910/_0_ , \g73922/_0_ , \g73934/_0_ , \g73946/_0_ , \g73958/_0_ , \g73970/_0_ , \g73982/_0_ , \g87036/_0_ , \g87042/_0_ , \g87043/_0_ , \g87044/_0_ , \g87045/_0_ , \g87046/_0_ , \g87047/_0_ , \g87048/_0_ , \g87049/_0_ , \g87050/_0_ , \g87051/_0_ , \g87052/_0_ , \g87053/_0_ , \g87054/_0_ , \g87055/_0_ , \g87062/_0_ , \g88572/_0_ , \g88681/_0_ , \g88682/_0_ , \g88683/_0_ , \g88684/_0_ , \g88685/_0_ , \g88686/_0_ , \g88687/_0_ , \g88688/_0_ , \g88689/_0_ , \g88690/_0_ , \g88691/_0_ , \g88692/_0_ , \g88693/_0_ , \g88695/_0_ , \g88697/_0_ , \g88698/_0_ , \g88700/_0_ , \g88701/_0_ , \g88703/_0_ , \g88704/_0_ , \g88705/_0_ , \g88706/_0_ , \g88707/_0_ , \g88709/_0_ , \g88710/_0_ , \g88711/_0_ , \g88712/_0_ , \g88713/_0_ , \g88714/_0_ , \g88716/_0_ , \g88717/_0_ , \g88718/_0_ , \g88719/_0_ , \g88720/_0_ , \g88722/_0_ , \g88723/_0_ , \g88724/_0_ , \g88725/_0_ , \g88726/_0_ , \g88727/_0_ , \g88728/_0_ , \g88729/_0_ , \g88731/_0_ , \g88732/_0_ , \g88733/_0_ , \g88734/_0_ , \g88736/_0_ , \g88737/_0_ , \g88738/_0_ , \g88739/_0_ , \g88740/_0_ , \g88741/_0_ , \g88742/_0_ , \g88743/_0_ , \g88744/_0_ , \g88745/_0_ , \g88746/_0_ , \g88748/_0_ , \g88749/_0_ , \g88750/_0_ , \g88752/_0_ , \g88753/_0_ , \g88754/_0_ , \g88755/_0_ , \g88756/_0_ , \g88757/_0_ , \g88759/_0_ , \g88760/_0_ , \g88761/_0_ , \g88762/_0_ , \g88764/_0_ , \g88765/_0_ , \g88766/_0_ , \g88768/_0_ , \g88769/_0_ , \g88770/_0_ , \g88771/_0_ , \g88772/_0_ , \g88773/_0_ , \g88775/_0_ , \g88776/_0_ , \g88777/_0_ , \g88778/_0_ , \g88779/_0_ , \g88780/_0_ , \g88782/_0_ , \g88783/_0_ , \g88784/_0_ , \g88785/_0_ , \g88786/_0_ , \g88787/_0_ , \g88789/_0_ , \g88790/_0_ , \g88791/_0_ , \g88792/_0_ , \g88793/_0_ , \g88795/_0_ , \g88796/_0_ , \g88797/_0_ , \g88799/_0_ , \g88800/_0_ , \g88801/_0_ , \g88802/_0_ , \g88806/_0_ , \g88807/_0_ , \g88808/_0_ , \g88809/_0_ , \g88810/_0_ , \g88813/_0_ , \g88814/_0_ , \g88815/_0_ , \m0_ack_o_pad , \m0_data_o[0]_pad , \m0_data_o[10]_pad , \m0_data_o[11]_pad , \m0_data_o[12]_pad , \m0_data_o[13]_pad , \m0_data_o[14]_pad , \m0_data_o[15]_pad , \m0_data_o[16]_pad , \m0_data_o[17]_pad , \m0_data_o[18]_pad , \m0_data_o[19]_pad , \m0_data_o[1]_pad , \m0_data_o[20]_pad , \m0_data_o[21]_pad , \m0_data_o[22]_pad , \m0_data_o[23]_pad , \m0_data_o[24]_pad , \m0_data_o[25]_pad , \m0_data_o[26]_pad , \m0_data_o[27]_pad , \m0_data_o[28]_pad , \m0_data_o[29]_pad , \m0_data_o[2]_pad , \m0_data_o[30]_pad , \m0_data_o[31]_pad , \m0_data_o[3]_pad , \m0_data_o[4]_pad , \m0_data_o[5]_pad , \m0_data_o[6]_pad , \m0_data_o[7]_pad , \m0_data_o[8]_pad , \m0_data_o[9]_pad , \m0_err_o_pad , \m0_rty_o_pad , \m1_ack_o_pad , \m1_data_o[0]_pad , \m1_data_o[10]_pad , \m1_data_o[11]_pad , \m1_data_o[12]_pad , \m1_data_o[13]_pad , \m1_data_o[14]_pad , \m1_data_o[15]_pad , \m1_data_o[16]_pad , \m1_data_o[17]_pad , \m1_data_o[18]_pad , \m1_data_o[19]_pad , \m1_data_o[1]_pad , \m1_data_o[20]_pad , \m1_data_o[21]_pad , \m1_data_o[22]_pad , \m1_data_o[23]_pad , \m1_data_o[24]_pad , \m1_data_o[25]_pad , \m1_data_o[26]_pad , \m1_data_o[27]_pad , \m1_data_o[28]_pad , \m1_data_o[29]_pad , \m1_data_o[2]_pad , \m1_data_o[30]_pad , \m1_data_o[31]_pad , \m1_data_o[3]_pad , \m1_data_o[4]_pad , \m1_data_o[5]_pad , \m1_data_o[6]_pad , \m1_data_o[7]_pad , \m1_data_o[8]_pad , \m1_data_o[9]_pad , \m1_err_o_pad , \m1_rty_o_pad , \m2_ack_o_pad , \m2_data_o[0]_pad , \m2_data_o[10]_pad , \m2_data_o[11]_pad , \m2_data_o[12]_pad , \m2_data_o[13]_pad , \m2_data_o[14]_pad , \m2_data_o[15]_pad , \m2_data_o[16]_pad , \m2_data_o[17]_pad , \m2_data_o[18]_pad , \m2_data_o[19]_pad , \m2_data_o[1]_pad , \m2_data_o[20]_pad , \m2_data_o[21]_pad , \m2_data_o[22]_pad , \m2_data_o[23]_pad , \m2_data_o[24]_pad , \m2_data_o[25]_pad , \m2_data_o[26]_pad , \m2_data_o[27]_pad , \m2_data_o[28]_pad , \m2_data_o[29]_pad , \m2_data_o[2]_pad , \m2_data_o[30]_pad , \m2_data_o[31]_pad , \m2_data_o[3]_pad , \m2_data_o[4]_pad , \m2_data_o[5]_pad , \m2_data_o[6]_pad , \m2_data_o[7]_pad , \m2_data_o[8]_pad , \m2_data_o[9]_pad , \m2_err_o_pad , \m2_rty_o_pad , \m3_ack_o_pad , \m3_data_o[0]_pad , \m3_data_o[10]_pad , \m3_data_o[11]_pad , \m3_data_o[12]_pad , \m3_data_o[13]_pad , \m3_data_o[14]_pad , \m3_data_o[15]_pad , \m3_data_o[16]_pad , \m3_data_o[17]_pad , \m3_data_o[18]_pad , \m3_data_o[19]_pad , \m3_data_o[1]_pad , \m3_data_o[20]_pad , \m3_data_o[21]_pad , \m3_data_o[22]_pad , \m3_data_o[23]_pad , \m3_data_o[24]_pad , \m3_data_o[25]_pad , \m3_data_o[26]_pad , \m3_data_o[27]_pad , \m3_data_o[28]_pad , \m3_data_o[29]_pad , \m3_data_o[2]_pad , \m3_data_o[30]_pad , \m3_data_o[31]_pad , \m3_data_o[3]_pad , \m3_data_o[4]_pad , \m3_data_o[5]_pad , \m3_data_o[6]_pad , \m3_data_o[7]_pad , \m3_data_o[8]_pad , \m3_data_o[9]_pad , \m3_err_o_pad , \m3_rty_o_pad , \m4_ack_o_pad , \m4_data_o[0]_pad , \m4_data_o[10]_pad , \m4_data_o[11]_pad , \m4_data_o[12]_pad , \m4_data_o[13]_pad , \m4_data_o[14]_pad , \m4_data_o[15]_pad , \m4_data_o[16]_pad , \m4_data_o[17]_pad , \m4_data_o[18]_pad , \m4_data_o[19]_pad , \m4_data_o[1]_pad , \m4_data_o[20]_pad , \m4_data_o[21]_pad , \m4_data_o[22]_pad , \m4_data_o[23]_pad , \m4_data_o[24]_pad , \m4_data_o[25]_pad , \m4_data_o[26]_pad , \m4_data_o[27]_pad , \m4_data_o[28]_pad , \m4_data_o[29]_pad , \m4_data_o[2]_pad , \m4_data_o[30]_pad , \m4_data_o[31]_pad , \m4_data_o[3]_pad , \m4_data_o[4]_pad , \m4_data_o[5]_pad , \m4_data_o[6]_pad , \m4_data_o[7]_pad , \m4_data_o[8]_pad , \m4_data_o[9]_pad , \m4_err_o_pad , \m4_rty_o_pad , \m5_ack_o_pad , \m5_data_o[0]_pad , \m5_data_o[10]_pad , \m5_data_o[11]_pad , \m5_data_o[12]_pad , \m5_data_o[13]_pad , \m5_data_o[14]_pad , \m5_data_o[15]_pad , \m5_data_o[16]_pad , \m5_data_o[17]_pad , \m5_data_o[18]_pad , \m5_data_o[19]_pad , \m5_data_o[1]_pad , \m5_data_o[20]_pad , \m5_data_o[21]_pad , \m5_data_o[22]_pad , \m5_data_o[23]_pad , \m5_data_o[24]_pad , \m5_data_o[25]_pad , \m5_data_o[26]_pad , \m5_data_o[27]_pad , \m5_data_o[28]_pad , \m5_data_o[29]_pad , \m5_data_o[2]_pad , \m5_data_o[30]_pad , \m5_data_o[31]_pad , \m5_data_o[3]_pad , \m5_data_o[4]_pad , \m5_data_o[5]_pad , \m5_data_o[6]_pad , \m5_data_o[7]_pad , \m5_data_o[8]_pad , \m5_data_o[9]_pad , \m5_err_o_pad , \m5_rty_o_pad , \m6_ack_o_pad , \m6_data_o[0]_pad , \m6_data_o[10]_pad , \m6_data_o[11]_pad , \m6_data_o[12]_pad , \m6_data_o[13]_pad , \m6_data_o[14]_pad , \m6_data_o[15]_pad , \m6_data_o[16]_pad , \m6_data_o[17]_pad , \m6_data_o[18]_pad , \m6_data_o[19]_pad , \m6_data_o[1]_pad , \m6_data_o[20]_pad , \m6_data_o[21]_pad , \m6_data_o[22]_pad , \m6_data_o[23]_pad , \m6_data_o[24]_pad , \m6_data_o[25]_pad , \m6_data_o[26]_pad , \m6_data_o[27]_pad , \m6_data_o[28]_pad , \m6_data_o[29]_pad , \m6_data_o[2]_pad , \m6_data_o[30]_pad , \m6_data_o[31]_pad , \m6_data_o[3]_pad , \m6_data_o[4]_pad , \m6_data_o[5]_pad , \m6_data_o[6]_pad , \m6_data_o[7]_pad , \m6_data_o[8]_pad , \m6_data_o[9]_pad , \m6_err_o_pad , \m6_rty_o_pad , \m7_ack_o_pad , \m7_data_o[0]_pad , \m7_data_o[10]_pad , \m7_data_o[11]_pad , \m7_data_o[12]_pad , \m7_data_o[13]_pad , \m7_data_o[14]_pad , \m7_data_o[15]_pad , \m7_data_o[16]_pad , \m7_data_o[17]_pad , \m7_data_o[18]_pad , \m7_data_o[19]_pad , \m7_data_o[1]_pad , \m7_data_o[20]_pad , \m7_data_o[21]_pad , \m7_data_o[22]_pad , \m7_data_o[23]_pad , \m7_data_o[24]_pad , \m7_data_o[25]_pad , \m7_data_o[26]_pad , \m7_data_o[27]_pad , \m7_data_o[28]_pad , \m7_data_o[29]_pad , \m7_data_o[2]_pad , \m7_data_o[30]_pad , \m7_data_o[31]_pad , \m7_data_o[3]_pad , \m7_data_o[4]_pad , \m7_data_o[5]_pad , \m7_data_o[6]_pad , \m7_data_o[7]_pad , \m7_data_o[8]_pad , \m7_data_o[9]_pad , \m7_err_o_pad , \m7_rty_o_pad , \s0_addr_o[0]_pad , \s0_addr_o[10]_pad , \s0_addr_o[11]_pad , \s0_addr_o[12]_pad , \s0_addr_o[13]_pad , \s0_addr_o[14]_pad , \s0_addr_o[15]_pad , \s0_addr_o[16]_pad , \s0_addr_o[17]_pad , \s0_addr_o[18]_pad , \s0_addr_o[19]_pad , \s0_addr_o[1]_pad , \s0_addr_o[20]_pad , \s0_addr_o[21]_pad , \s0_addr_o[22]_pad , \s0_addr_o[23]_pad , \s0_addr_o[24]_pad , \s0_addr_o[25]_pad , \s0_addr_o[26]_pad , \s0_addr_o[27]_pad , \s0_addr_o[28]_pad , \s0_addr_o[29]_pad , \s0_addr_o[2]_pad , \s0_addr_o[30]_pad , \s0_addr_o[31]_pad , \s0_addr_o[3]_pad , \s0_addr_o[4]_pad , \s0_addr_o[5]_pad , \s0_addr_o[6]_pad , \s0_addr_o[7]_pad , \s0_addr_o[8]_pad , \s0_addr_o[9]_pad , \s0_data_o[0]_pad , \s0_data_o[10]_pad , \s0_data_o[11]_pad , \s0_data_o[12]_pad , \s0_data_o[13]_pad , \s0_data_o[14]_pad , \s0_data_o[15]_pad , \s0_data_o[16]_pad , \s0_data_o[17]_pad , \s0_data_o[18]_pad , \s0_data_o[19]_pad , \s0_data_o[1]_pad , \s0_data_o[20]_pad , \s0_data_o[21]_pad , \s0_data_o[22]_pad , \s0_data_o[23]_pad , \s0_data_o[24]_pad , \s0_data_o[25]_pad , \s0_data_o[26]_pad , \s0_data_o[27]_pad , \s0_data_o[28]_pad , \s0_data_o[29]_pad , \s0_data_o[2]_pad , \s0_data_o[30]_pad , \s0_data_o[31]_pad , \s0_data_o[3]_pad , \s0_data_o[4]_pad , \s0_data_o[5]_pad , \s0_data_o[6]_pad , \s0_data_o[7]_pad , \s0_data_o[8]_pad , \s0_data_o[9]_pad , \s0_sel_o[0]_pad , \s0_sel_o[1]_pad , \s0_sel_o[2]_pad , \s0_sel_o[3]_pad , \s0_stb_o_pad , \s0_we_o_pad , \s10_addr_o[0]_pad , \s10_addr_o[10]_pad , \s10_addr_o[11]_pad , \s10_addr_o[12]_pad , \s10_addr_o[13]_pad , \s10_addr_o[14]_pad , \s10_addr_o[15]_pad , \s10_addr_o[16]_pad , \s10_addr_o[17]_pad , \s10_addr_o[18]_pad , \s10_addr_o[19]_pad , \s10_addr_o[1]_pad , \s10_addr_o[20]_pad , \s10_addr_o[21]_pad , \s10_addr_o[22]_pad , \s10_addr_o[23]_pad , \s10_addr_o[24]_pad , \s10_addr_o[25]_pad , \s10_addr_o[26]_pad , \s10_addr_o[27]_pad , \s10_addr_o[28]_pad , \s10_addr_o[29]_pad , \s10_addr_o[2]_pad , \s10_addr_o[30]_pad , \s10_addr_o[31]_pad , \s10_addr_o[3]_pad , \s10_addr_o[4]_pad , \s10_addr_o[5]_pad , \s10_addr_o[6]_pad , \s10_addr_o[7]_pad , \s10_addr_o[8]_pad , \s10_addr_o[9]_pad , \s10_data_o[0]_pad , \s10_data_o[10]_pad , \s10_data_o[11]_pad , \s10_data_o[12]_pad , \s10_data_o[13]_pad , \s10_data_o[14]_pad , \s10_data_o[15]_pad , \s10_data_o[16]_pad , \s10_data_o[17]_pad , \s10_data_o[18]_pad , \s10_data_o[19]_pad , \s10_data_o[1]_pad , \s10_data_o[20]_pad , \s10_data_o[21]_pad , \s10_data_o[22]_pad , \s10_data_o[23]_pad , \s10_data_o[24]_pad , \s10_data_o[25]_pad , \s10_data_o[26]_pad , \s10_data_o[27]_pad , \s10_data_o[28]_pad , \s10_data_o[29]_pad , \s10_data_o[2]_pad , \s10_data_o[30]_pad , \s10_data_o[31]_pad , \s10_data_o[3]_pad , \s10_data_o[4]_pad , \s10_data_o[5]_pad , \s10_data_o[6]_pad , \s10_data_o[7]_pad , \s10_data_o[8]_pad , \s10_data_o[9]_pad , \s10_sel_o[0]_pad , \s10_sel_o[1]_pad , \s10_sel_o[2]_pad , \s10_sel_o[3]_pad , \s10_stb_o_pad , \s10_we_o_pad , \s11_addr_o[0]_pad , \s11_addr_o[10]_pad , \s11_addr_o[11]_pad , \s11_addr_o[12]_pad , \s11_addr_o[13]_pad , \s11_addr_o[14]_pad , \s11_addr_o[15]_pad , \s11_addr_o[16]_pad , \s11_addr_o[17]_pad , \s11_addr_o[18]_pad , \s11_addr_o[19]_pad , \s11_addr_o[1]_pad , \s11_addr_o[20]_pad , \s11_addr_o[21]_pad , \s11_addr_o[22]_pad , \s11_addr_o[23]_pad , \s11_addr_o[24]_pad , \s11_addr_o[25]_pad , \s11_addr_o[26]_pad , \s11_addr_o[27]_pad , \s11_addr_o[28]_pad , \s11_addr_o[29]_pad , \s11_addr_o[2]_pad , \s11_addr_o[30]_pad , \s11_addr_o[31]_pad , \s11_addr_o[3]_pad , \s11_addr_o[4]_pad , \s11_addr_o[5]_pad , \s11_addr_o[6]_pad , \s11_addr_o[7]_pad , \s11_addr_o[8]_pad , \s11_addr_o[9]_pad , \s11_data_o[0]_pad , \s11_data_o[10]_pad , \s11_data_o[11]_pad , \s11_data_o[12]_pad , \s11_data_o[13]_pad , \s11_data_o[14]_pad , \s11_data_o[15]_pad , \s11_data_o[16]_pad , \s11_data_o[17]_pad , \s11_data_o[18]_pad , \s11_data_o[19]_pad , \s11_data_o[1]_pad , \s11_data_o[20]_pad , \s11_data_o[21]_pad , \s11_data_o[22]_pad , \s11_data_o[23]_pad , \s11_data_o[24]_pad , \s11_data_o[25]_pad , \s11_data_o[26]_pad , \s11_data_o[27]_pad , \s11_data_o[28]_pad , \s11_data_o[29]_pad , \s11_data_o[2]_pad , \s11_data_o[30]_pad , \s11_data_o[31]_pad , \s11_data_o[3]_pad , \s11_data_o[4]_pad , \s11_data_o[5]_pad , \s11_data_o[6]_pad , \s11_data_o[7]_pad , \s11_data_o[8]_pad , \s11_data_o[9]_pad , \s11_sel_o[0]_pad , \s11_sel_o[1]_pad , \s11_sel_o[2]_pad , \s11_sel_o[3]_pad , \s11_stb_o_pad , \s11_we_o_pad , \s12_addr_o[0]_pad , \s12_addr_o[10]_pad , \s12_addr_o[11]_pad , \s12_addr_o[12]_pad , \s12_addr_o[13]_pad , \s12_addr_o[14]_pad , \s12_addr_o[15]_pad , \s12_addr_o[16]_pad , \s12_addr_o[17]_pad , \s12_addr_o[18]_pad , \s12_addr_o[19]_pad , \s12_addr_o[1]_pad , \s12_addr_o[20]_pad , \s12_addr_o[21]_pad , \s12_addr_o[22]_pad , \s12_addr_o[23]_pad , \s12_addr_o[24]_pad , \s12_addr_o[25]_pad , \s12_addr_o[26]_pad , \s12_addr_o[27]_pad , \s12_addr_o[28]_pad , \s12_addr_o[29]_pad , \s12_addr_o[2]_pad , \s12_addr_o[30]_pad , \s12_addr_o[31]_pad , \s12_addr_o[3]_pad , \s12_addr_o[4]_pad , \s12_addr_o[5]_pad , \s12_addr_o[6]_pad , \s12_addr_o[7]_pad , \s12_addr_o[8]_pad , \s12_addr_o[9]_pad , \s12_data_o[0]_pad , \s12_data_o[10]_pad , \s12_data_o[11]_pad , \s12_data_o[12]_pad , \s12_data_o[13]_pad , \s12_data_o[14]_pad , \s12_data_o[15]_pad , \s12_data_o[16]_pad , \s12_data_o[17]_pad , \s12_data_o[18]_pad , \s12_data_o[19]_pad , \s12_data_o[1]_pad , \s12_data_o[20]_pad , \s12_data_o[21]_pad , \s12_data_o[22]_pad , \s12_data_o[23]_pad , \s12_data_o[24]_pad , \s12_data_o[25]_pad , \s12_data_o[26]_pad , \s12_data_o[27]_pad , \s12_data_o[28]_pad , \s12_data_o[29]_pad , \s12_data_o[2]_pad , \s12_data_o[30]_pad , \s12_data_o[31]_pad , \s12_data_o[3]_pad , \s12_data_o[4]_pad , \s12_data_o[5]_pad , \s12_data_o[6]_pad , \s12_data_o[7]_pad , \s12_data_o[8]_pad , \s12_data_o[9]_pad , \s12_sel_o[0]_pad , \s12_sel_o[1]_pad , \s12_sel_o[2]_pad , \s12_sel_o[3]_pad , \s12_stb_o_pad , \s12_we_o_pad , \s13_addr_o[0]_pad , \s13_addr_o[10]_pad , \s13_addr_o[11]_pad , \s13_addr_o[12]_pad , \s13_addr_o[13]_pad , \s13_addr_o[14]_pad , \s13_addr_o[15]_pad , \s13_addr_o[16]_pad , \s13_addr_o[17]_pad , \s13_addr_o[18]_pad , \s13_addr_o[19]_pad , \s13_addr_o[1]_pad , \s13_addr_o[20]_pad , \s13_addr_o[21]_pad , \s13_addr_o[22]_pad , \s13_addr_o[23]_pad , \s13_addr_o[24]_pad , \s13_addr_o[25]_pad , \s13_addr_o[26]_pad , \s13_addr_o[27]_pad , \s13_addr_o[28]_pad , \s13_addr_o[29]_pad , \s13_addr_o[2]_pad , \s13_addr_o[30]_pad , \s13_addr_o[31]_pad , \s13_addr_o[3]_pad , \s13_addr_o[4]_pad , \s13_addr_o[5]_pad , \s13_addr_o[6]_pad , \s13_addr_o[7]_pad , \s13_addr_o[8]_pad , \s13_addr_o[9]_pad , \s13_data_o[0]_pad , \s13_data_o[10]_pad , \s13_data_o[11]_pad , \s13_data_o[12]_pad , \s13_data_o[13]_pad , \s13_data_o[14]_pad , \s13_data_o[15]_pad , \s13_data_o[16]_pad , \s13_data_o[17]_pad , \s13_data_o[18]_pad , \s13_data_o[19]_pad , \s13_data_o[1]_pad , \s13_data_o[20]_pad , \s13_data_o[21]_pad , \s13_data_o[22]_pad , \s13_data_o[23]_pad , \s13_data_o[24]_pad , \s13_data_o[25]_pad , \s13_data_o[26]_pad , \s13_data_o[27]_pad , \s13_data_o[28]_pad , \s13_data_o[29]_pad , \s13_data_o[2]_pad , \s13_data_o[30]_pad , \s13_data_o[31]_pad , \s13_data_o[3]_pad , \s13_data_o[4]_pad , \s13_data_o[5]_pad , \s13_data_o[6]_pad , \s13_data_o[7]_pad , \s13_data_o[8]_pad , \s13_data_o[9]_pad , \s13_sel_o[0]_pad , \s13_sel_o[1]_pad , \s13_sel_o[2]_pad , \s13_sel_o[3]_pad , \s13_stb_o_pad , \s13_we_o_pad , \s14_addr_o[0]_pad , \s14_addr_o[10]_pad , \s14_addr_o[11]_pad , \s14_addr_o[12]_pad , \s14_addr_o[13]_pad , \s14_addr_o[14]_pad , \s14_addr_o[15]_pad , \s14_addr_o[16]_pad , \s14_addr_o[17]_pad , \s14_addr_o[18]_pad , \s14_addr_o[19]_pad , \s14_addr_o[1]_pad , \s14_addr_o[20]_pad , \s14_addr_o[21]_pad , \s14_addr_o[22]_pad , \s14_addr_o[23]_pad , \s14_addr_o[24]_pad , \s14_addr_o[25]_pad , \s14_addr_o[26]_pad , \s14_addr_o[27]_pad , \s14_addr_o[28]_pad , \s14_addr_o[29]_pad , \s14_addr_o[2]_pad , \s14_addr_o[30]_pad , \s14_addr_o[31]_pad , \s14_addr_o[3]_pad , \s14_addr_o[4]_pad , \s14_addr_o[5]_pad , \s14_addr_o[6]_pad , \s14_addr_o[7]_pad , \s14_addr_o[8]_pad , \s14_addr_o[9]_pad , \s14_data_o[0]_pad , \s14_data_o[10]_pad , \s14_data_o[11]_pad , \s14_data_o[12]_pad , \s14_data_o[13]_pad , \s14_data_o[14]_pad , \s14_data_o[15]_pad , \s14_data_o[16]_pad , \s14_data_o[17]_pad , \s14_data_o[18]_pad , \s14_data_o[19]_pad , \s14_data_o[1]_pad , \s14_data_o[20]_pad , \s14_data_o[21]_pad , \s14_data_o[22]_pad , \s14_data_o[23]_pad , \s14_data_o[24]_pad , \s14_data_o[25]_pad , \s14_data_o[26]_pad , \s14_data_o[27]_pad , \s14_data_o[28]_pad , \s14_data_o[29]_pad , \s14_data_o[2]_pad , \s14_data_o[30]_pad , \s14_data_o[31]_pad , \s14_data_o[3]_pad , \s14_data_o[4]_pad , \s14_data_o[5]_pad , \s14_data_o[6]_pad , \s14_data_o[7]_pad , \s14_data_o[8]_pad , \s14_data_o[9]_pad , \s14_sel_o[0]_pad , \s14_sel_o[1]_pad , \s14_sel_o[2]_pad , \s14_sel_o[3]_pad , \s14_stb_o_pad , \s14_we_o_pad , \s15_addr_o[0]_pad , \s15_addr_o[10]_pad , \s15_addr_o[11]_pad , \s15_addr_o[12]_pad , \s15_addr_o[13]_pad , \s15_addr_o[14]_pad , \s15_addr_o[15]_pad , \s15_addr_o[16]_pad , \s15_addr_o[17]_pad , \s15_addr_o[18]_pad , \s15_addr_o[19]_pad , \s15_addr_o[1]_pad , \s15_addr_o[20]_pad , \s15_addr_o[21]_pad , \s15_addr_o[22]_pad , \s15_addr_o[23]_pad , \s15_addr_o[24]_pad , \s15_addr_o[25]_pad , \s15_addr_o[26]_pad , \s15_addr_o[27]_pad , \s15_addr_o[28]_pad , \s15_addr_o[29]_pad , \s15_addr_o[2]_pad , \s15_addr_o[30]_pad , \s15_addr_o[31]_pad , \s15_addr_o[3]_pad , \s15_addr_o[4]_pad , \s15_addr_o[6]_pad , \s15_addr_o[7]_pad , \s15_addr_o[8]_pad , \s15_addr_o[9]_pad , \s15_cyc_o_pad , \s15_data_o[0]_pad , \s15_data_o[10]_pad , \s15_data_o[11]_pad , \s15_data_o[12]_pad , \s15_data_o[13]_pad , \s15_data_o[14]_pad , \s15_data_o[15]_pad , \s15_data_o[16]_pad , \s15_data_o[17]_pad , \s15_data_o[18]_pad , \s15_data_o[19]_pad , \s15_data_o[1]_pad , \s15_data_o[20]_pad , \s15_data_o[21]_pad , \s15_data_o[22]_pad , \s15_data_o[23]_pad , \s15_data_o[24]_pad , \s15_data_o[25]_pad , \s15_data_o[26]_pad , \s15_data_o[27]_pad , \s15_data_o[28]_pad , \s15_data_o[29]_pad , \s15_data_o[2]_pad , \s15_data_o[30]_pad , \s15_data_o[31]_pad , \s15_data_o[3]_pad , \s15_data_o[4]_pad , \s15_data_o[5]_pad , \s15_data_o[6]_pad , \s15_data_o[7]_pad , \s15_data_o[8]_pad , \s15_data_o[9]_pad , \s15_sel_o[0]_pad , \s15_sel_o[1]_pad , \s15_sel_o[2]_pad , \s15_sel_o[3]_pad , \s15_stb_o_pad , \s15_we_o_pad , \s1_addr_o[0]_pad , \s1_addr_o[10]_pad , \s1_addr_o[11]_pad , \s1_addr_o[12]_pad , \s1_addr_o[13]_pad , \s1_addr_o[14]_pad , \s1_addr_o[15]_pad , \s1_addr_o[16]_pad , \s1_addr_o[17]_pad , \s1_addr_o[18]_pad , \s1_addr_o[19]_pad , \s1_addr_o[1]_pad , \s1_addr_o[20]_pad , \s1_addr_o[21]_pad , \s1_addr_o[22]_pad , \s1_addr_o[23]_pad , \s1_addr_o[24]_pad , \s1_addr_o[25]_pad , \s1_addr_o[26]_pad , \s1_addr_o[27]_pad , \s1_addr_o[28]_pad , \s1_addr_o[29]_pad , \s1_addr_o[2]_pad , \s1_addr_o[30]_pad , \s1_addr_o[31]_pad , \s1_addr_o[3]_pad , \s1_addr_o[4]_pad , \s1_addr_o[5]_pad , \s1_addr_o[6]_pad , \s1_addr_o[7]_pad , \s1_addr_o[8]_pad , \s1_addr_o[9]_pad , \s1_data_o[0]_pad , \s1_data_o[10]_pad , \s1_data_o[11]_pad , \s1_data_o[12]_pad , \s1_data_o[13]_pad , \s1_data_o[14]_pad , \s1_data_o[15]_pad , \s1_data_o[16]_pad , \s1_data_o[17]_pad , \s1_data_o[18]_pad , \s1_data_o[19]_pad , \s1_data_o[1]_pad , \s1_data_o[20]_pad , \s1_data_o[21]_pad , \s1_data_o[22]_pad , \s1_data_o[23]_pad , \s1_data_o[24]_pad , \s1_data_o[25]_pad , \s1_data_o[26]_pad , \s1_data_o[27]_pad , \s1_data_o[28]_pad , \s1_data_o[29]_pad , \s1_data_o[2]_pad , \s1_data_o[30]_pad , \s1_data_o[31]_pad , \s1_data_o[3]_pad , \s1_data_o[4]_pad , \s1_data_o[5]_pad , \s1_data_o[6]_pad , \s1_data_o[7]_pad , \s1_data_o[8]_pad , \s1_data_o[9]_pad , \s1_sel_o[0]_pad , \s1_sel_o[1]_pad , \s1_sel_o[2]_pad , \s1_sel_o[3]_pad , \s1_stb_o_pad , \s1_we_o_pad , \s2_addr_o[0]_pad , \s2_addr_o[10]_pad , \s2_addr_o[11]_pad , \s2_addr_o[12]_pad , \s2_addr_o[13]_pad , \s2_addr_o[14]_pad , \s2_addr_o[15]_pad , \s2_addr_o[16]_pad , \s2_addr_o[17]_pad , \s2_addr_o[18]_pad , \s2_addr_o[19]_pad , \s2_addr_o[1]_pad , \s2_addr_o[20]_pad , \s2_addr_o[21]_pad , \s2_addr_o[22]_pad , \s2_addr_o[23]_pad , \s2_addr_o[24]_pad , \s2_addr_o[25]_pad , \s2_addr_o[26]_pad , \s2_addr_o[27]_pad , \s2_addr_o[28]_pad , \s2_addr_o[29]_pad , \s2_addr_o[2]_pad , \s2_addr_o[30]_pad , \s2_addr_o[31]_pad , \s2_addr_o[3]_pad , \s2_addr_o[4]_pad , \s2_addr_o[5]_pad , \s2_addr_o[6]_pad , \s2_addr_o[7]_pad , \s2_addr_o[8]_pad , \s2_addr_o[9]_pad , \s2_data_o[0]_pad , \s2_data_o[10]_pad , \s2_data_o[11]_pad , \s2_data_o[12]_pad , \s2_data_o[13]_pad , \s2_data_o[14]_pad , \s2_data_o[15]_pad , \s2_data_o[16]_pad , \s2_data_o[17]_pad , \s2_data_o[18]_pad , \s2_data_o[19]_pad , \s2_data_o[1]_pad , \s2_data_o[20]_pad , \s2_data_o[21]_pad , \s2_data_o[22]_pad , \s2_data_o[23]_pad , \s2_data_o[24]_pad , \s2_data_o[25]_pad , \s2_data_o[26]_pad , \s2_data_o[27]_pad , \s2_data_o[28]_pad , \s2_data_o[29]_pad , \s2_data_o[2]_pad , \s2_data_o[30]_pad , \s2_data_o[31]_pad , \s2_data_o[3]_pad , \s2_data_o[4]_pad , \s2_data_o[5]_pad , \s2_data_o[6]_pad , \s2_data_o[7]_pad , \s2_data_o[8]_pad , \s2_data_o[9]_pad , \s2_sel_o[0]_pad , \s2_sel_o[1]_pad , \s2_sel_o[2]_pad , \s2_sel_o[3]_pad , \s2_stb_o_pad , \s2_we_o_pad , \s3_addr_o[0]_pad , \s3_addr_o[10]_pad , \s3_addr_o[11]_pad , \s3_addr_o[12]_pad , \s3_addr_o[13]_pad , \s3_addr_o[14]_pad , \s3_addr_o[15]_pad , \s3_addr_o[16]_pad , \s3_addr_o[17]_pad , \s3_addr_o[18]_pad , \s3_addr_o[19]_pad , \s3_addr_o[1]_pad , \s3_addr_o[20]_pad , \s3_addr_o[21]_pad , \s3_addr_o[22]_pad , \s3_addr_o[23]_pad , \s3_addr_o[24]_pad , \s3_addr_o[25]_pad , \s3_addr_o[26]_pad , \s3_addr_o[27]_pad , \s3_addr_o[28]_pad , \s3_addr_o[29]_pad , \s3_addr_o[2]_pad , \s3_addr_o[30]_pad , \s3_addr_o[31]_pad , \s3_addr_o[3]_pad , \s3_addr_o[4]_pad , \s3_addr_o[5]_pad , \s3_addr_o[6]_pad , \s3_addr_o[7]_pad , \s3_addr_o[8]_pad , \s3_addr_o[9]_pad , \s3_data_o[0]_pad , \s3_data_o[10]_pad , \s3_data_o[11]_pad , \s3_data_o[12]_pad , \s3_data_o[13]_pad , \s3_data_o[14]_pad , \s3_data_o[15]_pad , \s3_data_o[16]_pad , \s3_data_o[17]_pad , \s3_data_o[18]_pad , \s3_data_o[19]_pad , \s3_data_o[1]_pad , \s3_data_o[20]_pad , \s3_data_o[21]_pad , \s3_data_o[22]_pad , \s3_data_o[23]_pad , \s3_data_o[24]_pad , \s3_data_o[25]_pad , \s3_data_o[26]_pad , \s3_data_o[27]_pad , \s3_data_o[28]_pad , \s3_data_o[29]_pad , \s3_data_o[2]_pad , \s3_data_o[30]_pad , \s3_data_o[31]_pad , \s3_data_o[3]_pad , \s3_data_o[4]_pad , \s3_data_o[5]_pad , \s3_data_o[6]_pad , \s3_data_o[7]_pad , \s3_data_o[8]_pad , \s3_data_o[9]_pad , \s3_sel_o[0]_pad , \s3_sel_o[1]_pad , \s3_sel_o[2]_pad , \s3_sel_o[3]_pad , \s3_stb_o_pad , \s3_we_o_pad , \s4_addr_o[0]_pad , \s4_addr_o[10]_pad , \s4_addr_o[11]_pad , \s4_addr_o[12]_pad , \s4_addr_o[13]_pad , \s4_addr_o[14]_pad , \s4_addr_o[15]_pad , \s4_addr_o[16]_pad , \s4_addr_o[17]_pad , \s4_addr_o[18]_pad , \s4_addr_o[19]_pad , \s4_addr_o[1]_pad , \s4_addr_o[20]_pad , \s4_addr_o[21]_pad , \s4_addr_o[22]_pad , \s4_addr_o[23]_pad , \s4_addr_o[24]_pad , \s4_addr_o[25]_pad , \s4_addr_o[26]_pad , \s4_addr_o[27]_pad , \s4_addr_o[28]_pad , \s4_addr_o[29]_pad , \s4_addr_o[2]_pad , \s4_addr_o[30]_pad , \s4_addr_o[31]_pad , \s4_addr_o[3]_pad , \s4_addr_o[4]_pad , \s4_addr_o[5]_pad , \s4_addr_o[6]_pad , \s4_addr_o[7]_pad , \s4_addr_o[8]_pad , \s4_addr_o[9]_pad , \s4_data_o[0]_pad , \s4_data_o[10]_pad , \s4_data_o[11]_pad , \s4_data_o[12]_pad , \s4_data_o[13]_pad , \s4_data_o[14]_pad , \s4_data_o[15]_pad , \s4_data_o[16]_pad , \s4_data_o[17]_pad , \s4_data_o[18]_pad , \s4_data_o[19]_pad , \s4_data_o[1]_pad , \s4_data_o[20]_pad , \s4_data_o[21]_pad , \s4_data_o[22]_pad , \s4_data_o[23]_pad , \s4_data_o[24]_pad , \s4_data_o[25]_pad , \s4_data_o[26]_pad , \s4_data_o[27]_pad , \s4_data_o[28]_pad , \s4_data_o[29]_pad , \s4_data_o[2]_pad , \s4_data_o[30]_pad , \s4_data_o[31]_pad , \s4_data_o[3]_pad , \s4_data_o[4]_pad , \s4_data_o[5]_pad , \s4_data_o[6]_pad , \s4_data_o[7]_pad , \s4_data_o[8]_pad , \s4_data_o[9]_pad , \s4_sel_o[0]_pad , \s4_sel_o[1]_pad , \s4_sel_o[2]_pad , \s4_sel_o[3]_pad , \s4_stb_o_pad , \s4_we_o_pad , \s5_addr_o[0]_pad , \s5_addr_o[10]_pad , \s5_addr_o[11]_pad , \s5_addr_o[12]_pad , \s5_addr_o[13]_pad , \s5_addr_o[14]_pad , \s5_addr_o[15]_pad , \s5_addr_o[16]_pad , \s5_addr_o[17]_pad , \s5_addr_o[18]_pad , \s5_addr_o[19]_pad , \s5_addr_o[1]_pad , \s5_addr_o[20]_pad , \s5_addr_o[21]_pad , \s5_addr_o[22]_pad , \s5_addr_o[23]_pad , \s5_addr_o[24]_pad , \s5_addr_o[25]_pad , \s5_addr_o[26]_pad , \s5_addr_o[27]_pad , \s5_addr_o[28]_pad , \s5_addr_o[29]_pad , \s5_addr_o[2]_pad , \s5_addr_o[30]_pad , \s5_addr_o[31]_pad , \s5_addr_o[3]_pad , \s5_addr_o[4]_pad , \s5_addr_o[5]_pad , \s5_addr_o[6]_pad , \s5_addr_o[7]_pad , \s5_addr_o[8]_pad , \s5_addr_o[9]_pad , \s5_data_o[0]_pad , \s5_data_o[10]_pad , \s5_data_o[11]_pad , \s5_data_o[12]_pad , \s5_data_o[13]_pad , \s5_data_o[14]_pad , \s5_data_o[15]_pad , \s5_data_o[16]_pad , \s5_data_o[17]_pad , \s5_data_o[18]_pad , \s5_data_o[19]_pad , \s5_data_o[1]_pad , \s5_data_o[20]_pad , \s5_data_o[21]_pad , \s5_data_o[22]_pad , \s5_data_o[23]_pad , \s5_data_o[24]_pad , \s5_data_o[25]_pad , \s5_data_o[26]_pad , \s5_data_o[27]_pad , \s5_data_o[28]_pad , \s5_data_o[29]_pad , \s5_data_o[2]_pad , \s5_data_o[30]_pad , \s5_data_o[31]_pad , \s5_data_o[3]_pad , \s5_data_o[4]_pad , \s5_data_o[5]_pad , \s5_data_o[6]_pad , \s5_data_o[7]_pad , \s5_data_o[8]_pad , \s5_data_o[9]_pad , \s5_sel_o[0]_pad , \s5_sel_o[1]_pad , \s5_sel_o[2]_pad , \s5_sel_o[3]_pad , \s5_stb_o_pad , \s5_we_o_pad , \s6_addr_o[0]_pad , \s6_addr_o[10]_pad , \s6_addr_o[11]_pad , \s6_addr_o[12]_pad , \s6_addr_o[13]_pad , \s6_addr_o[14]_pad , \s6_addr_o[15]_pad , \s6_addr_o[16]_pad , \s6_addr_o[17]_pad , \s6_addr_o[18]_pad , \s6_addr_o[19]_pad , \s6_addr_o[1]_pad , \s6_addr_o[20]_pad , \s6_addr_o[21]_pad , \s6_addr_o[22]_pad , \s6_addr_o[23]_pad , \s6_addr_o[24]_pad , \s6_addr_o[25]_pad , \s6_addr_o[26]_pad , \s6_addr_o[27]_pad , \s6_addr_o[28]_pad , \s6_addr_o[29]_pad , \s6_addr_o[2]_pad , \s6_addr_o[30]_pad , \s6_addr_o[31]_pad , \s6_addr_o[3]_pad , \s6_addr_o[4]_pad , \s6_addr_o[5]_pad , \s6_addr_o[6]_pad , \s6_addr_o[7]_pad , \s6_addr_o[8]_pad , \s6_addr_o[9]_pad , \s6_data_o[0]_pad , \s6_data_o[10]_pad , \s6_data_o[11]_pad , \s6_data_o[12]_pad , \s6_data_o[13]_pad , \s6_data_o[14]_pad , \s6_data_o[15]_pad , \s6_data_o[16]_pad , \s6_data_o[17]_pad , \s6_data_o[18]_pad , \s6_data_o[19]_pad , \s6_data_o[1]_pad , \s6_data_o[20]_pad , \s6_data_o[21]_pad , \s6_data_o[22]_pad , \s6_data_o[23]_pad , \s6_data_o[24]_pad , \s6_data_o[25]_pad , \s6_data_o[26]_pad , \s6_data_o[27]_pad , \s6_data_o[28]_pad , \s6_data_o[29]_pad , \s6_data_o[2]_pad , \s6_data_o[30]_pad , \s6_data_o[31]_pad , \s6_data_o[3]_pad , \s6_data_o[4]_pad , \s6_data_o[5]_pad , \s6_data_o[6]_pad , \s6_data_o[7]_pad , \s6_data_o[8]_pad , \s6_data_o[9]_pad , \s6_sel_o[0]_pad , \s6_sel_o[1]_pad , \s6_sel_o[2]_pad , \s6_sel_o[3]_pad , \s6_stb_o_pad , \s6_we_o_pad , \s7_addr_o[0]_pad , \s7_addr_o[10]_pad , \s7_addr_o[11]_pad , \s7_addr_o[12]_pad , \s7_addr_o[13]_pad , \s7_addr_o[14]_pad , \s7_addr_o[15]_pad , \s7_addr_o[16]_pad , \s7_addr_o[17]_pad , \s7_addr_o[18]_pad , \s7_addr_o[19]_pad , \s7_addr_o[1]_pad , \s7_addr_o[20]_pad , \s7_addr_o[21]_pad , \s7_addr_o[22]_pad , \s7_addr_o[23]_pad , \s7_addr_o[24]_pad , \s7_addr_o[25]_pad , \s7_addr_o[26]_pad , \s7_addr_o[27]_pad , \s7_addr_o[28]_pad , \s7_addr_o[29]_pad , \s7_addr_o[2]_pad , \s7_addr_o[30]_pad , \s7_addr_o[31]_pad , \s7_addr_o[3]_pad , \s7_addr_o[4]_pad , \s7_addr_o[5]_pad , \s7_addr_o[6]_pad , \s7_addr_o[7]_pad , \s7_addr_o[8]_pad , \s7_addr_o[9]_pad , \s7_data_o[0]_pad , \s7_data_o[10]_pad , \s7_data_o[11]_pad , \s7_data_o[12]_pad , \s7_data_o[13]_pad , \s7_data_o[14]_pad , \s7_data_o[15]_pad , \s7_data_o[16]_pad , \s7_data_o[17]_pad , \s7_data_o[18]_pad , \s7_data_o[19]_pad , \s7_data_o[1]_pad , \s7_data_o[20]_pad , \s7_data_o[21]_pad , \s7_data_o[22]_pad , \s7_data_o[23]_pad , \s7_data_o[24]_pad , \s7_data_o[25]_pad , \s7_data_o[26]_pad , \s7_data_o[27]_pad , \s7_data_o[28]_pad , \s7_data_o[29]_pad , \s7_data_o[2]_pad , \s7_data_o[30]_pad , \s7_data_o[31]_pad , \s7_data_o[3]_pad , \s7_data_o[4]_pad , \s7_data_o[5]_pad , \s7_data_o[6]_pad , \s7_data_o[7]_pad , \s7_data_o[8]_pad , \s7_data_o[9]_pad , \s7_sel_o[0]_pad , \s7_sel_o[1]_pad , \s7_sel_o[2]_pad , \s7_sel_o[3]_pad , \s7_stb_o_pad , \s7_we_o_pad , \s8_addr_o[0]_pad , \s8_addr_o[10]_pad , \s8_addr_o[11]_pad , \s8_addr_o[12]_pad , \s8_addr_o[13]_pad , \s8_addr_o[14]_pad , \s8_addr_o[15]_pad , \s8_addr_o[16]_pad , \s8_addr_o[17]_pad , \s8_addr_o[18]_pad , \s8_addr_o[19]_pad , \s8_addr_o[1]_pad , \s8_addr_o[20]_pad , \s8_addr_o[21]_pad , \s8_addr_o[22]_pad , \s8_addr_o[23]_pad , \s8_addr_o[24]_pad , \s8_addr_o[25]_pad , \s8_addr_o[26]_pad , \s8_addr_o[27]_pad , \s8_addr_o[28]_pad , \s8_addr_o[29]_pad , \s8_addr_o[2]_pad , \s8_addr_o[30]_pad , \s8_addr_o[31]_pad , \s8_addr_o[3]_pad , \s8_addr_o[4]_pad , \s8_addr_o[5]_pad , \s8_addr_o[6]_pad , \s8_addr_o[7]_pad , \s8_addr_o[8]_pad , \s8_addr_o[9]_pad , \s8_data_o[0]_pad , \s8_data_o[10]_pad , \s8_data_o[11]_pad , \s8_data_o[12]_pad , \s8_data_o[13]_pad , \s8_data_o[14]_pad , \s8_data_o[15]_pad , \s8_data_o[16]_pad , \s8_data_o[17]_pad , \s8_data_o[18]_pad , \s8_data_o[19]_pad , \s8_data_o[1]_pad , \s8_data_o[20]_pad , \s8_data_o[21]_pad , \s8_data_o[22]_pad , \s8_data_o[23]_pad , \s8_data_o[24]_pad , \s8_data_o[25]_pad , \s8_data_o[26]_pad , \s8_data_o[27]_pad , \s8_data_o[28]_pad , \s8_data_o[29]_pad , \s8_data_o[2]_pad , \s8_data_o[30]_pad , \s8_data_o[31]_pad , \s8_data_o[3]_pad , \s8_data_o[4]_pad , \s8_data_o[5]_pad , \s8_data_o[6]_pad , \s8_data_o[7]_pad , \s8_data_o[8]_pad , \s8_data_o[9]_pad , \s8_sel_o[0]_pad , \s8_sel_o[1]_pad , \s8_sel_o[2]_pad , \s8_sel_o[3]_pad , \s8_stb_o_pad , \s8_we_o_pad , \s9_addr_o[0]_pad , \s9_addr_o[10]_pad , \s9_addr_o[11]_pad , \s9_addr_o[12]_pad , \s9_addr_o[13]_pad , \s9_addr_o[14]_pad , \s9_addr_o[15]_pad , \s9_addr_o[16]_pad , \s9_addr_o[17]_pad , \s9_addr_o[18]_pad , \s9_addr_o[19]_pad , \s9_addr_o[1]_pad , \s9_addr_o[20]_pad , \s9_addr_o[21]_pad , \s9_addr_o[22]_pad , \s9_addr_o[23]_pad , \s9_addr_o[24]_pad , \s9_addr_o[25]_pad , \s9_addr_o[26]_pad , \s9_addr_o[27]_pad , \s9_addr_o[28]_pad , \s9_addr_o[29]_pad , \s9_addr_o[2]_pad , \s9_addr_o[30]_pad , \s9_addr_o[31]_pad , \s9_addr_o[3]_pad , \s9_addr_o[4]_pad , \s9_addr_o[5]_pad , \s9_addr_o[6]_pad , \s9_addr_o[7]_pad , \s9_addr_o[8]_pad , \s9_addr_o[9]_pad , \s9_data_o[0]_pad , \s9_data_o[10]_pad , \s9_data_o[11]_pad , \s9_data_o[12]_pad , \s9_data_o[13]_pad , \s9_data_o[14]_pad , \s9_data_o[15]_pad , \s9_data_o[16]_pad , \s9_data_o[17]_pad , \s9_data_o[18]_pad , \s9_data_o[19]_pad , \s9_data_o[1]_pad , \s9_data_o[20]_pad , \s9_data_o[21]_pad , \s9_data_o[22]_pad , \s9_data_o[23]_pad , \s9_data_o[24]_pad , \s9_data_o[25]_pad , \s9_data_o[26]_pad , \s9_data_o[27]_pad , \s9_data_o[28]_pad , \s9_data_o[29]_pad , \s9_data_o[2]_pad , \s9_data_o[30]_pad , \s9_data_o[31]_pad , \s9_data_o[3]_pad , \s9_data_o[4]_pad , \s9_data_o[5]_pad , \s9_data_o[6]_pad , \s9_data_o[7]_pad , \s9_data_o[8]_pad , \s9_data_o[9]_pad , \s9_sel_o[0]_pad , \s9_sel_o[1]_pad , \s9_sel_o[2]_pad , \s9_sel_o[3]_pad , \s9_stb_o_pad , \s9_we_o_pad );
	input \m0_addr_i[0]_pad  ;
	input \m0_addr_i[10]_pad  ;
	input \m0_addr_i[11]_pad  ;
	input \m0_addr_i[12]_pad  ;
	input \m0_addr_i[13]_pad  ;
	input \m0_addr_i[14]_pad  ;
	input \m0_addr_i[15]_pad  ;
	input \m0_addr_i[16]_pad  ;
	input \m0_addr_i[17]_pad  ;
	input \m0_addr_i[18]_pad  ;
	input \m0_addr_i[19]_pad  ;
	input \m0_addr_i[1]_pad  ;
	input \m0_addr_i[20]_pad  ;
	input \m0_addr_i[21]_pad  ;
	input \m0_addr_i[22]_pad  ;
	input \m0_addr_i[23]_pad  ;
	input \m0_addr_i[24]_pad  ;
	input \m0_addr_i[25]_pad  ;
	input \m0_addr_i[26]_pad  ;
	input \m0_addr_i[27]_pad  ;
	input \m0_addr_i[28]_pad  ;
	input \m0_addr_i[29]_pad  ;
	input \m0_addr_i[2]_pad  ;
	input \m0_addr_i[30]_pad  ;
	input \m0_addr_i[31]_pad  ;
	input \m0_addr_i[3]_pad  ;
	input \m0_addr_i[4]_pad  ;
	input \m0_addr_i[5]_pad  ;
	input \m0_addr_i[6]_pad  ;
	input \m0_addr_i[7]_pad  ;
	input \m0_addr_i[8]_pad  ;
	input \m0_addr_i[9]_pad  ;
	input \m0_cyc_i_pad  ;
	input \m0_data_i[0]_pad  ;
	input \m0_data_i[10]_pad  ;
	input \m0_data_i[11]_pad  ;
	input \m0_data_i[12]_pad  ;
	input \m0_data_i[13]_pad  ;
	input \m0_data_i[14]_pad  ;
	input \m0_data_i[15]_pad  ;
	input \m0_data_i[16]_pad  ;
	input \m0_data_i[17]_pad  ;
	input \m0_data_i[18]_pad  ;
	input \m0_data_i[19]_pad  ;
	input \m0_data_i[1]_pad  ;
	input \m0_data_i[20]_pad  ;
	input \m0_data_i[21]_pad  ;
	input \m0_data_i[22]_pad  ;
	input \m0_data_i[23]_pad  ;
	input \m0_data_i[24]_pad  ;
	input \m0_data_i[25]_pad  ;
	input \m0_data_i[26]_pad  ;
	input \m0_data_i[27]_pad  ;
	input \m0_data_i[28]_pad  ;
	input \m0_data_i[29]_pad  ;
	input \m0_data_i[2]_pad  ;
	input \m0_data_i[30]_pad  ;
	input \m0_data_i[31]_pad  ;
	input \m0_data_i[3]_pad  ;
	input \m0_data_i[4]_pad  ;
	input \m0_data_i[5]_pad  ;
	input \m0_data_i[6]_pad  ;
	input \m0_data_i[7]_pad  ;
	input \m0_data_i[8]_pad  ;
	input \m0_data_i[9]_pad  ;
	input \m0_s0_cyc_o_reg/NET0131  ;
	input \m0_s10_cyc_o_reg/NET0131  ;
	input \m0_s11_cyc_o_reg/NET0131  ;
	input \m0_s12_cyc_o_reg/NET0131  ;
	input \m0_s13_cyc_o_reg/NET0131  ;
	input \m0_s14_cyc_o_reg/NET0131  ;
	input \m0_s15_cyc_o_reg/NET0131  ;
	input \m0_s1_cyc_o_reg/NET0131  ;
	input \m0_s2_cyc_o_reg/NET0131  ;
	input \m0_s3_cyc_o_reg/NET0131  ;
	input \m0_s4_cyc_o_reg/NET0131  ;
	input \m0_s5_cyc_o_reg/NET0131  ;
	input \m0_s6_cyc_o_reg/NET0131  ;
	input \m0_s7_cyc_o_reg/NET0131  ;
	input \m0_s8_cyc_o_reg/NET0131  ;
	input \m0_s9_cyc_o_reg/NET0131  ;
	input \m0_sel_i[0]_pad  ;
	input \m0_sel_i[1]_pad  ;
	input \m0_sel_i[2]_pad  ;
	input \m0_sel_i[3]_pad  ;
	input \m0_stb_i_pad  ;
	input \m0_we_i_pad  ;
	input \m1_addr_i[0]_pad  ;
	input \m1_addr_i[10]_pad  ;
	input \m1_addr_i[11]_pad  ;
	input \m1_addr_i[12]_pad  ;
	input \m1_addr_i[13]_pad  ;
	input \m1_addr_i[14]_pad  ;
	input \m1_addr_i[15]_pad  ;
	input \m1_addr_i[16]_pad  ;
	input \m1_addr_i[17]_pad  ;
	input \m1_addr_i[18]_pad  ;
	input \m1_addr_i[19]_pad  ;
	input \m1_addr_i[1]_pad  ;
	input \m1_addr_i[20]_pad  ;
	input \m1_addr_i[21]_pad  ;
	input \m1_addr_i[22]_pad  ;
	input \m1_addr_i[23]_pad  ;
	input \m1_addr_i[24]_pad  ;
	input \m1_addr_i[25]_pad  ;
	input \m1_addr_i[26]_pad  ;
	input \m1_addr_i[27]_pad  ;
	input \m1_addr_i[28]_pad  ;
	input \m1_addr_i[29]_pad  ;
	input \m1_addr_i[2]_pad  ;
	input \m1_addr_i[30]_pad  ;
	input \m1_addr_i[31]_pad  ;
	input \m1_addr_i[3]_pad  ;
	input \m1_addr_i[4]_pad  ;
	input \m1_addr_i[5]_pad  ;
	input \m1_addr_i[6]_pad  ;
	input \m1_addr_i[7]_pad  ;
	input \m1_addr_i[8]_pad  ;
	input \m1_addr_i[9]_pad  ;
	input \m1_cyc_i_pad  ;
	input \m1_data_i[0]_pad  ;
	input \m1_data_i[10]_pad  ;
	input \m1_data_i[11]_pad  ;
	input \m1_data_i[12]_pad  ;
	input \m1_data_i[13]_pad  ;
	input \m1_data_i[14]_pad  ;
	input \m1_data_i[15]_pad  ;
	input \m1_data_i[16]_pad  ;
	input \m1_data_i[17]_pad  ;
	input \m1_data_i[18]_pad  ;
	input \m1_data_i[19]_pad  ;
	input \m1_data_i[1]_pad  ;
	input \m1_data_i[20]_pad  ;
	input \m1_data_i[21]_pad  ;
	input \m1_data_i[22]_pad  ;
	input \m1_data_i[23]_pad  ;
	input \m1_data_i[24]_pad  ;
	input \m1_data_i[25]_pad  ;
	input \m1_data_i[26]_pad  ;
	input \m1_data_i[27]_pad  ;
	input \m1_data_i[28]_pad  ;
	input \m1_data_i[29]_pad  ;
	input \m1_data_i[2]_pad  ;
	input \m1_data_i[30]_pad  ;
	input \m1_data_i[31]_pad  ;
	input \m1_data_i[3]_pad  ;
	input \m1_data_i[4]_pad  ;
	input \m1_data_i[5]_pad  ;
	input \m1_data_i[6]_pad  ;
	input \m1_data_i[7]_pad  ;
	input \m1_data_i[8]_pad  ;
	input \m1_data_i[9]_pad  ;
	input \m1_s0_cyc_o_reg/NET0131  ;
	input \m1_s10_cyc_o_reg/NET0131  ;
	input \m1_s11_cyc_o_reg/NET0131  ;
	input \m1_s12_cyc_o_reg/NET0131  ;
	input \m1_s13_cyc_o_reg/NET0131  ;
	input \m1_s14_cyc_o_reg/NET0131  ;
	input \m1_s15_cyc_o_reg/NET0131  ;
	input \m1_s1_cyc_o_reg/NET0131  ;
	input \m1_s2_cyc_o_reg/NET0131  ;
	input \m1_s3_cyc_o_reg/NET0131  ;
	input \m1_s4_cyc_o_reg/NET0131  ;
	input \m1_s5_cyc_o_reg/NET0131  ;
	input \m1_s6_cyc_o_reg/NET0131  ;
	input \m1_s7_cyc_o_reg/NET0131  ;
	input \m1_s8_cyc_o_reg/NET0131  ;
	input \m1_s9_cyc_o_reg/NET0131  ;
	input \m1_sel_i[0]_pad  ;
	input \m1_sel_i[1]_pad  ;
	input \m1_sel_i[2]_pad  ;
	input \m1_sel_i[3]_pad  ;
	input \m1_stb_i_pad  ;
	input \m1_we_i_pad  ;
	input \m2_addr_i[0]_pad  ;
	input \m2_addr_i[10]_pad  ;
	input \m2_addr_i[11]_pad  ;
	input \m2_addr_i[12]_pad  ;
	input \m2_addr_i[13]_pad  ;
	input \m2_addr_i[14]_pad  ;
	input \m2_addr_i[15]_pad  ;
	input \m2_addr_i[16]_pad  ;
	input \m2_addr_i[17]_pad  ;
	input \m2_addr_i[18]_pad  ;
	input \m2_addr_i[19]_pad  ;
	input \m2_addr_i[1]_pad  ;
	input \m2_addr_i[20]_pad  ;
	input \m2_addr_i[21]_pad  ;
	input \m2_addr_i[22]_pad  ;
	input \m2_addr_i[23]_pad  ;
	input \m2_addr_i[24]_pad  ;
	input \m2_addr_i[25]_pad  ;
	input \m2_addr_i[26]_pad  ;
	input \m2_addr_i[27]_pad  ;
	input \m2_addr_i[28]_pad  ;
	input \m2_addr_i[29]_pad  ;
	input \m2_addr_i[2]_pad  ;
	input \m2_addr_i[30]_pad  ;
	input \m2_addr_i[31]_pad  ;
	input \m2_addr_i[3]_pad  ;
	input \m2_addr_i[4]_pad  ;
	input \m2_addr_i[5]_pad  ;
	input \m2_addr_i[6]_pad  ;
	input \m2_addr_i[7]_pad  ;
	input \m2_addr_i[8]_pad  ;
	input \m2_addr_i[9]_pad  ;
	input \m2_cyc_i_pad  ;
	input \m2_data_i[0]_pad  ;
	input \m2_data_i[10]_pad  ;
	input \m2_data_i[11]_pad  ;
	input \m2_data_i[12]_pad  ;
	input \m2_data_i[13]_pad  ;
	input \m2_data_i[14]_pad  ;
	input \m2_data_i[15]_pad  ;
	input \m2_data_i[16]_pad  ;
	input \m2_data_i[17]_pad  ;
	input \m2_data_i[18]_pad  ;
	input \m2_data_i[19]_pad  ;
	input \m2_data_i[1]_pad  ;
	input \m2_data_i[20]_pad  ;
	input \m2_data_i[21]_pad  ;
	input \m2_data_i[22]_pad  ;
	input \m2_data_i[23]_pad  ;
	input \m2_data_i[24]_pad  ;
	input \m2_data_i[25]_pad  ;
	input \m2_data_i[26]_pad  ;
	input \m2_data_i[27]_pad  ;
	input \m2_data_i[28]_pad  ;
	input \m2_data_i[29]_pad  ;
	input \m2_data_i[2]_pad  ;
	input \m2_data_i[30]_pad  ;
	input \m2_data_i[31]_pad  ;
	input \m2_data_i[3]_pad  ;
	input \m2_data_i[4]_pad  ;
	input \m2_data_i[5]_pad  ;
	input \m2_data_i[6]_pad  ;
	input \m2_data_i[7]_pad  ;
	input \m2_data_i[8]_pad  ;
	input \m2_data_i[9]_pad  ;
	input \m2_s0_cyc_o_reg/NET0131  ;
	input \m2_s10_cyc_o_reg/NET0131  ;
	input \m2_s11_cyc_o_reg/NET0131  ;
	input \m2_s12_cyc_o_reg/NET0131  ;
	input \m2_s13_cyc_o_reg/NET0131  ;
	input \m2_s14_cyc_o_reg/NET0131  ;
	input \m2_s15_cyc_o_reg/NET0131  ;
	input \m2_s1_cyc_o_reg/NET0131  ;
	input \m2_s2_cyc_o_reg/NET0131  ;
	input \m2_s3_cyc_o_reg/NET0131  ;
	input \m2_s4_cyc_o_reg/NET0131  ;
	input \m2_s5_cyc_o_reg/NET0131  ;
	input \m2_s6_cyc_o_reg/NET0131  ;
	input \m2_s7_cyc_o_reg/NET0131  ;
	input \m2_s8_cyc_o_reg/NET0131  ;
	input \m2_s9_cyc_o_reg/NET0131  ;
	input \m2_sel_i[0]_pad  ;
	input \m2_sel_i[1]_pad  ;
	input \m2_sel_i[2]_pad  ;
	input \m2_sel_i[3]_pad  ;
	input \m2_stb_i_pad  ;
	input \m2_we_i_pad  ;
	input \m3_addr_i[0]_pad  ;
	input \m3_addr_i[10]_pad  ;
	input \m3_addr_i[11]_pad  ;
	input \m3_addr_i[12]_pad  ;
	input \m3_addr_i[13]_pad  ;
	input \m3_addr_i[14]_pad  ;
	input \m3_addr_i[15]_pad  ;
	input \m3_addr_i[16]_pad  ;
	input \m3_addr_i[17]_pad  ;
	input \m3_addr_i[18]_pad  ;
	input \m3_addr_i[19]_pad  ;
	input \m3_addr_i[1]_pad  ;
	input \m3_addr_i[20]_pad  ;
	input \m3_addr_i[21]_pad  ;
	input \m3_addr_i[22]_pad  ;
	input \m3_addr_i[23]_pad  ;
	input \m3_addr_i[24]_pad  ;
	input \m3_addr_i[25]_pad  ;
	input \m3_addr_i[26]_pad  ;
	input \m3_addr_i[27]_pad  ;
	input \m3_addr_i[28]_pad  ;
	input \m3_addr_i[29]_pad  ;
	input \m3_addr_i[2]_pad  ;
	input \m3_addr_i[30]_pad  ;
	input \m3_addr_i[31]_pad  ;
	input \m3_addr_i[3]_pad  ;
	input \m3_addr_i[4]_pad  ;
	input \m3_addr_i[5]_pad  ;
	input \m3_addr_i[6]_pad  ;
	input \m3_addr_i[7]_pad  ;
	input \m3_addr_i[8]_pad  ;
	input \m3_addr_i[9]_pad  ;
	input \m3_cyc_i_pad  ;
	input \m3_data_i[0]_pad  ;
	input \m3_data_i[10]_pad  ;
	input \m3_data_i[11]_pad  ;
	input \m3_data_i[12]_pad  ;
	input \m3_data_i[13]_pad  ;
	input \m3_data_i[14]_pad  ;
	input \m3_data_i[15]_pad  ;
	input \m3_data_i[16]_pad  ;
	input \m3_data_i[17]_pad  ;
	input \m3_data_i[18]_pad  ;
	input \m3_data_i[19]_pad  ;
	input \m3_data_i[1]_pad  ;
	input \m3_data_i[20]_pad  ;
	input \m3_data_i[21]_pad  ;
	input \m3_data_i[22]_pad  ;
	input \m3_data_i[23]_pad  ;
	input \m3_data_i[24]_pad  ;
	input \m3_data_i[25]_pad  ;
	input \m3_data_i[26]_pad  ;
	input \m3_data_i[27]_pad  ;
	input \m3_data_i[28]_pad  ;
	input \m3_data_i[29]_pad  ;
	input \m3_data_i[2]_pad  ;
	input \m3_data_i[30]_pad  ;
	input \m3_data_i[31]_pad  ;
	input \m3_data_i[3]_pad  ;
	input \m3_data_i[4]_pad  ;
	input \m3_data_i[5]_pad  ;
	input \m3_data_i[6]_pad  ;
	input \m3_data_i[7]_pad  ;
	input \m3_data_i[8]_pad  ;
	input \m3_data_i[9]_pad  ;
	input \m3_s0_cyc_o_reg/NET0131  ;
	input \m3_s10_cyc_o_reg/NET0131  ;
	input \m3_s11_cyc_o_reg/NET0131  ;
	input \m3_s12_cyc_o_reg/NET0131  ;
	input \m3_s13_cyc_o_reg/NET0131  ;
	input \m3_s14_cyc_o_reg/NET0131  ;
	input \m3_s15_cyc_o_reg/NET0131  ;
	input \m3_s1_cyc_o_reg/NET0131  ;
	input \m3_s2_cyc_o_reg/NET0131  ;
	input \m3_s3_cyc_o_reg/NET0131  ;
	input \m3_s4_cyc_o_reg/NET0131  ;
	input \m3_s5_cyc_o_reg/NET0131  ;
	input \m3_s6_cyc_o_reg/NET0131  ;
	input \m3_s7_cyc_o_reg/NET0131  ;
	input \m3_s8_cyc_o_reg/NET0131  ;
	input \m3_s9_cyc_o_reg/NET0131  ;
	input \m3_sel_i[0]_pad  ;
	input \m3_sel_i[1]_pad  ;
	input \m3_sel_i[2]_pad  ;
	input \m3_sel_i[3]_pad  ;
	input \m3_stb_i_pad  ;
	input \m3_we_i_pad  ;
	input \m4_addr_i[0]_pad  ;
	input \m4_addr_i[10]_pad  ;
	input \m4_addr_i[11]_pad  ;
	input \m4_addr_i[12]_pad  ;
	input \m4_addr_i[13]_pad  ;
	input \m4_addr_i[14]_pad  ;
	input \m4_addr_i[15]_pad  ;
	input \m4_addr_i[16]_pad  ;
	input \m4_addr_i[17]_pad  ;
	input \m4_addr_i[18]_pad  ;
	input \m4_addr_i[19]_pad  ;
	input \m4_addr_i[1]_pad  ;
	input \m4_addr_i[20]_pad  ;
	input \m4_addr_i[21]_pad  ;
	input \m4_addr_i[22]_pad  ;
	input \m4_addr_i[23]_pad  ;
	input \m4_addr_i[24]_pad  ;
	input \m4_addr_i[25]_pad  ;
	input \m4_addr_i[26]_pad  ;
	input \m4_addr_i[27]_pad  ;
	input \m4_addr_i[28]_pad  ;
	input \m4_addr_i[29]_pad  ;
	input \m4_addr_i[2]_pad  ;
	input \m4_addr_i[30]_pad  ;
	input \m4_addr_i[31]_pad  ;
	input \m4_addr_i[3]_pad  ;
	input \m4_addr_i[4]_pad  ;
	input \m4_addr_i[5]_pad  ;
	input \m4_addr_i[6]_pad  ;
	input \m4_addr_i[7]_pad  ;
	input \m4_addr_i[8]_pad  ;
	input \m4_addr_i[9]_pad  ;
	input \m4_cyc_i_pad  ;
	input \m4_data_i[0]_pad  ;
	input \m4_data_i[10]_pad  ;
	input \m4_data_i[11]_pad  ;
	input \m4_data_i[12]_pad  ;
	input \m4_data_i[13]_pad  ;
	input \m4_data_i[14]_pad  ;
	input \m4_data_i[15]_pad  ;
	input \m4_data_i[16]_pad  ;
	input \m4_data_i[17]_pad  ;
	input \m4_data_i[18]_pad  ;
	input \m4_data_i[19]_pad  ;
	input \m4_data_i[1]_pad  ;
	input \m4_data_i[20]_pad  ;
	input \m4_data_i[21]_pad  ;
	input \m4_data_i[22]_pad  ;
	input \m4_data_i[23]_pad  ;
	input \m4_data_i[24]_pad  ;
	input \m4_data_i[25]_pad  ;
	input \m4_data_i[26]_pad  ;
	input \m4_data_i[27]_pad  ;
	input \m4_data_i[28]_pad  ;
	input \m4_data_i[29]_pad  ;
	input \m4_data_i[2]_pad  ;
	input \m4_data_i[30]_pad  ;
	input \m4_data_i[31]_pad  ;
	input \m4_data_i[3]_pad  ;
	input \m4_data_i[4]_pad  ;
	input \m4_data_i[5]_pad  ;
	input \m4_data_i[6]_pad  ;
	input \m4_data_i[7]_pad  ;
	input \m4_data_i[8]_pad  ;
	input \m4_data_i[9]_pad  ;
	input \m4_s0_cyc_o_reg/NET0131  ;
	input \m4_s10_cyc_o_reg/NET0131  ;
	input \m4_s11_cyc_o_reg/NET0131  ;
	input \m4_s12_cyc_o_reg/NET0131  ;
	input \m4_s13_cyc_o_reg/NET0131  ;
	input \m4_s14_cyc_o_reg/NET0131  ;
	input \m4_s15_cyc_o_reg/NET0131  ;
	input \m4_s1_cyc_o_reg/NET0131  ;
	input \m4_s2_cyc_o_reg/NET0131  ;
	input \m4_s3_cyc_o_reg/NET0131  ;
	input \m4_s4_cyc_o_reg/NET0131  ;
	input \m4_s5_cyc_o_reg/NET0131  ;
	input \m4_s6_cyc_o_reg/NET0131  ;
	input \m4_s7_cyc_o_reg/NET0131  ;
	input \m4_s8_cyc_o_reg/NET0131  ;
	input \m4_s9_cyc_o_reg/NET0131  ;
	input \m4_sel_i[0]_pad  ;
	input \m4_sel_i[1]_pad  ;
	input \m4_sel_i[2]_pad  ;
	input \m4_sel_i[3]_pad  ;
	input \m4_stb_i_pad  ;
	input \m4_we_i_pad  ;
	input \m5_addr_i[0]_pad  ;
	input \m5_addr_i[10]_pad  ;
	input \m5_addr_i[11]_pad  ;
	input \m5_addr_i[12]_pad  ;
	input \m5_addr_i[13]_pad  ;
	input \m5_addr_i[14]_pad  ;
	input \m5_addr_i[15]_pad  ;
	input \m5_addr_i[16]_pad  ;
	input \m5_addr_i[17]_pad  ;
	input \m5_addr_i[18]_pad  ;
	input \m5_addr_i[19]_pad  ;
	input \m5_addr_i[1]_pad  ;
	input \m5_addr_i[20]_pad  ;
	input \m5_addr_i[21]_pad  ;
	input \m5_addr_i[22]_pad  ;
	input \m5_addr_i[23]_pad  ;
	input \m5_addr_i[24]_pad  ;
	input \m5_addr_i[25]_pad  ;
	input \m5_addr_i[26]_pad  ;
	input \m5_addr_i[27]_pad  ;
	input \m5_addr_i[28]_pad  ;
	input \m5_addr_i[29]_pad  ;
	input \m5_addr_i[2]_pad  ;
	input \m5_addr_i[30]_pad  ;
	input \m5_addr_i[31]_pad  ;
	input \m5_addr_i[3]_pad  ;
	input \m5_addr_i[4]_pad  ;
	input \m5_addr_i[5]_pad  ;
	input \m5_addr_i[6]_pad  ;
	input \m5_addr_i[7]_pad  ;
	input \m5_addr_i[8]_pad  ;
	input \m5_addr_i[9]_pad  ;
	input \m5_cyc_i_pad  ;
	input \m5_data_i[0]_pad  ;
	input \m5_data_i[10]_pad  ;
	input \m5_data_i[11]_pad  ;
	input \m5_data_i[12]_pad  ;
	input \m5_data_i[13]_pad  ;
	input \m5_data_i[14]_pad  ;
	input \m5_data_i[15]_pad  ;
	input \m5_data_i[16]_pad  ;
	input \m5_data_i[17]_pad  ;
	input \m5_data_i[18]_pad  ;
	input \m5_data_i[19]_pad  ;
	input \m5_data_i[1]_pad  ;
	input \m5_data_i[20]_pad  ;
	input \m5_data_i[21]_pad  ;
	input \m5_data_i[22]_pad  ;
	input \m5_data_i[23]_pad  ;
	input \m5_data_i[24]_pad  ;
	input \m5_data_i[25]_pad  ;
	input \m5_data_i[26]_pad  ;
	input \m5_data_i[27]_pad  ;
	input \m5_data_i[28]_pad  ;
	input \m5_data_i[29]_pad  ;
	input \m5_data_i[2]_pad  ;
	input \m5_data_i[30]_pad  ;
	input \m5_data_i[31]_pad  ;
	input \m5_data_i[3]_pad  ;
	input \m5_data_i[4]_pad  ;
	input \m5_data_i[5]_pad  ;
	input \m5_data_i[6]_pad  ;
	input \m5_data_i[7]_pad  ;
	input \m5_data_i[8]_pad  ;
	input \m5_data_i[9]_pad  ;
	input \m5_s0_cyc_o_reg/NET0131  ;
	input \m5_s10_cyc_o_reg/NET0131  ;
	input \m5_s11_cyc_o_reg/NET0131  ;
	input \m5_s12_cyc_o_reg/NET0131  ;
	input \m5_s13_cyc_o_reg/NET0131  ;
	input \m5_s14_cyc_o_reg/NET0131  ;
	input \m5_s15_cyc_o_reg/NET0131  ;
	input \m5_s1_cyc_o_reg/NET0131  ;
	input \m5_s2_cyc_o_reg/NET0131  ;
	input \m5_s3_cyc_o_reg/NET0131  ;
	input \m5_s4_cyc_o_reg/NET0131  ;
	input \m5_s5_cyc_o_reg/NET0131  ;
	input \m5_s6_cyc_o_reg/NET0131  ;
	input \m5_s7_cyc_o_reg/NET0131  ;
	input \m5_s8_cyc_o_reg/NET0131  ;
	input \m5_s9_cyc_o_reg/NET0131  ;
	input \m5_sel_i[0]_pad  ;
	input \m5_sel_i[1]_pad  ;
	input \m5_sel_i[2]_pad  ;
	input \m5_sel_i[3]_pad  ;
	input \m5_stb_i_pad  ;
	input \m5_we_i_pad  ;
	input \m6_addr_i[0]_pad  ;
	input \m6_addr_i[10]_pad  ;
	input \m6_addr_i[11]_pad  ;
	input \m6_addr_i[12]_pad  ;
	input \m6_addr_i[13]_pad  ;
	input \m6_addr_i[14]_pad  ;
	input \m6_addr_i[15]_pad  ;
	input \m6_addr_i[16]_pad  ;
	input \m6_addr_i[17]_pad  ;
	input \m6_addr_i[18]_pad  ;
	input \m6_addr_i[19]_pad  ;
	input \m6_addr_i[1]_pad  ;
	input \m6_addr_i[20]_pad  ;
	input \m6_addr_i[21]_pad  ;
	input \m6_addr_i[22]_pad  ;
	input \m6_addr_i[23]_pad  ;
	input \m6_addr_i[24]_pad  ;
	input \m6_addr_i[25]_pad  ;
	input \m6_addr_i[26]_pad  ;
	input \m6_addr_i[27]_pad  ;
	input \m6_addr_i[28]_pad  ;
	input \m6_addr_i[29]_pad  ;
	input \m6_addr_i[2]_pad  ;
	input \m6_addr_i[30]_pad  ;
	input \m6_addr_i[31]_pad  ;
	input \m6_addr_i[3]_pad  ;
	input \m6_addr_i[4]_pad  ;
	input \m6_addr_i[5]_pad  ;
	input \m6_addr_i[6]_pad  ;
	input \m6_addr_i[7]_pad  ;
	input \m6_addr_i[8]_pad  ;
	input \m6_addr_i[9]_pad  ;
	input \m6_cyc_i_pad  ;
	input \m6_data_i[0]_pad  ;
	input \m6_data_i[10]_pad  ;
	input \m6_data_i[11]_pad  ;
	input \m6_data_i[12]_pad  ;
	input \m6_data_i[13]_pad  ;
	input \m6_data_i[14]_pad  ;
	input \m6_data_i[15]_pad  ;
	input \m6_data_i[16]_pad  ;
	input \m6_data_i[17]_pad  ;
	input \m6_data_i[18]_pad  ;
	input \m6_data_i[19]_pad  ;
	input \m6_data_i[1]_pad  ;
	input \m6_data_i[20]_pad  ;
	input \m6_data_i[21]_pad  ;
	input \m6_data_i[22]_pad  ;
	input \m6_data_i[23]_pad  ;
	input \m6_data_i[24]_pad  ;
	input \m6_data_i[25]_pad  ;
	input \m6_data_i[26]_pad  ;
	input \m6_data_i[27]_pad  ;
	input \m6_data_i[28]_pad  ;
	input \m6_data_i[29]_pad  ;
	input \m6_data_i[2]_pad  ;
	input \m6_data_i[30]_pad  ;
	input \m6_data_i[31]_pad  ;
	input \m6_data_i[3]_pad  ;
	input \m6_data_i[4]_pad  ;
	input \m6_data_i[5]_pad  ;
	input \m6_data_i[6]_pad  ;
	input \m6_data_i[7]_pad  ;
	input \m6_data_i[8]_pad  ;
	input \m6_data_i[9]_pad  ;
	input \m6_s0_cyc_o_reg/NET0131  ;
	input \m6_s10_cyc_o_reg/NET0131  ;
	input \m6_s11_cyc_o_reg/NET0131  ;
	input \m6_s12_cyc_o_reg/NET0131  ;
	input \m6_s13_cyc_o_reg/NET0131  ;
	input \m6_s14_cyc_o_reg/NET0131  ;
	input \m6_s15_cyc_o_reg/NET0131  ;
	input \m6_s1_cyc_o_reg/NET0131  ;
	input \m6_s2_cyc_o_reg/NET0131  ;
	input \m6_s3_cyc_o_reg/NET0131  ;
	input \m6_s4_cyc_o_reg/NET0131  ;
	input \m6_s5_cyc_o_reg/NET0131  ;
	input \m6_s6_cyc_o_reg/NET0131  ;
	input \m6_s7_cyc_o_reg/NET0131  ;
	input \m6_s8_cyc_o_reg/NET0131  ;
	input \m6_s9_cyc_o_reg/NET0131  ;
	input \m6_sel_i[0]_pad  ;
	input \m6_sel_i[1]_pad  ;
	input \m6_sel_i[2]_pad  ;
	input \m6_sel_i[3]_pad  ;
	input \m6_stb_i_pad  ;
	input \m6_we_i_pad  ;
	input \m7_addr_i[0]_pad  ;
	input \m7_addr_i[10]_pad  ;
	input \m7_addr_i[11]_pad  ;
	input \m7_addr_i[12]_pad  ;
	input \m7_addr_i[13]_pad  ;
	input \m7_addr_i[14]_pad  ;
	input \m7_addr_i[15]_pad  ;
	input \m7_addr_i[16]_pad  ;
	input \m7_addr_i[17]_pad  ;
	input \m7_addr_i[18]_pad  ;
	input \m7_addr_i[19]_pad  ;
	input \m7_addr_i[1]_pad  ;
	input \m7_addr_i[20]_pad  ;
	input \m7_addr_i[21]_pad  ;
	input \m7_addr_i[22]_pad  ;
	input \m7_addr_i[23]_pad  ;
	input \m7_addr_i[24]_pad  ;
	input \m7_addr_i[25]_pad  ;
	input \m7_addr_i[26]_pad  ;
	input \m7_addr_i[27]_pad  ;
	input \m7_addr_i[28]_pad  ;
	input \m7_addr_i[29]_pad  ;
	input \m7_addr_i[2]_pad  ;
	input \m7_addr_i[30]_pad  ;
	input \m7_addr_i[31]_pad  ;
	input \m7_addr_i[3]_pad  ;
	input \m7_addr_i[4]_pad  ;
	input \m7_addr_i[5]_pad  ;
	input \m7_addr_i[6]_pad  ;
	input \m7_addr_i[7]_pad  ;
	input \m7_addr_i[8]_pad  ;
	input \m7_addr_i[9]_pad  ;
	input \m7_cyc_i_pad  ;
	input \m7_data_i[0]_pad  ;
	input \m7_data_i[10]_pad  ;
	input \m7_data_i[11]_pad  ;
	input \m7_data_i[12]_pad  ;
	input \m7_data_i[13]_pad  ;
	input \m7_data_i[14]_pad  ;
	input \m7_data_i[15]_pad  ;
	input \m7_data_i[16]_pad  ;
	input \m7_data_i[17]_pad  ;
	input \m7_data_i[18]_pad  ;
	input \m7_data_i[19]_pad  ;
	input \m7_data_i[1]_pad  ;
	input \m7_data_i[20]_pad  ;
	input \m7_data_i[21]_pad  ;
	input \m7_data_i[22]_pad  ;
	input \m7_data_i[23]_pad  ;
	input \m7_data_i[24]_pad  ;
	input \m7_data_i[25]_pad  ;
	input \m7_data_i[26]_pad  ;
	input \m7_data_i[27]_pad  ;
	input \m7_data_i[28]_pad  ;
	input \m7_data_i[29]_pad  ;
	input \m7_data_i[2]_pad  ;
	input \m7_data_i[30]_pad  ;
	input \m7_data_i[31]_pad  ;
	input \m7_data_i[3]_pad  ;
	input \m7_data_i[4]_pad  ;
	input \m7_data_i[5]_pad  ;
	input \m7_data_i[6]_pad  ;
	input \m7_data_i[7]_pad  ;
	input \m7_data_i[8]_pad  ;
	input \m7_data_i[9]_pad  ;
	input \m7_s0_cyc_o_reg/NET0131  ;
	input \m7_s10_cyc_o_reg/NET0131  ;
	input \m7_s11_cyc_o_reg/NET0131  ;
	input \m7_s12_cyc_o_reg/NET0131  ;
	input \m7_s13_cyc_o_reg/NET0131  ;
	input \m7_s14_cyc_o_reg/NET0131  ;
	input \m7_s15_cyc_o_reg/NET0131  ;
	input \m7_s1_cyc_o_reg/NET0131  ;
	input \m7_s2_cyc_o_reg/NET0131  ;
	input \m7_s3_cyc_o_reg/NET0131  ;
	input \m7_s4_cyc_o_reg/NET0131  ;
	input \m7_s5_cyc_o_reg/NET0131  ;
	input \m7_s6_cyc_o_reg/NET0131  ;
	input \m7_s7_cyc_o_reg/NET0131  ;
	input \m7_s8_cyc_o_reg/NET0131  ;
	input \m7_s9_cyc_o_reg/NET0131  ;
	input \m7_sel_i[0]_pad  ;
	input \m7_sel_i[1]_pad  ;
	input \m7_sel_i[2]_pad  ;
	input \m7_sel_i[3]_pad  ;
	input \m7_stb_i_pad  ;
	input \m7_we_i_pad  ;
	input \rf_conf0_reg[0]/NET0131  ;
	input \rf_conf0_reg[10]/NET0131  ;
	input \rf_conf0_reg[11]/NET0131  ;
	input \rf_conf0_reg[12]/NET0131  ;
	input \rf_conf0_reg[13]/NET0131  ;
	input \rf_conf0_reg[14]/NET0131  ;
	input \rf_conf0_reg[15]/NET0131  ;
	input \rf_conf0_reg[1]/NET0131  ;
	input \rf_conf0_reg[2]/NET0131  ;
	input \rf_conf0_reg[3]/NET0131  ;
	input \rf_conf0_reg[4]/NET0131  ;
	input \rf_conf0_reg[5]/NET0131  ;
	input \rf_conf0_reg[6]/NET0131  ;
	input \rf_conf0_reg[7]/NET0131  ;
	input \rf_conf0_reg[8]/NET0131  ;
	input \rf_conf0_reg[9]/NET0131  ;
	input \rf_conf10_reg[0]/NET0131  ;
	input \rf_conf10_reg[10]/NET0131  ;
	input \rf_conf10_reg[11]/NET0131  ;
	input \rf_conf10_reg[12]/NET0131  ;
	input \rf_conf10_reg[13]/NET0131  ;
	input \rf_conf10_reg[14]/NET0131  ;
	input \rf_conf10_reg[15]/NET0131  ;
	input \rf_conf10_reg[1]/NET0131  ;
	input \rf_conf10_reg[2]/NET0131  ;
	input \rf_conf10_reg[3]/NET0131  ;
	input \rf_conf10_reg[4]/NET0131  ;
	input \rf_conf10_reg[5]/NET0131  ;
	input \rf_conf10_reg[6]/NET0131  ;
	input \rf_conf10_reg[7]/NET0131  ;
	input \rf_conf10_reg[8]/NET0131  ;
	input \rf_conf10_reg[9]/NET0131  ;
	input \rf_conf11_reg[0]/NET0131  ;
	input \rf_conf11_reg[10]/NET0131  ;
	input \rf_conf11_reg[11]/NET0131  ;
	input \rf_conf11_reg[12]/NET0131  ;
	input \rf_conf11_reg[13]/NET0131  ;
	input \rf_conf11_reg[14]/NET0131  ;
	input \rf_conf11_reg[15]/NET0131  ;
	input \rf_conf11_reg[1]/NET0131  ;
	input \rf_conf11_reg[2]/NET0131  ;
	input \rf_conf11_reg[3]/NET0131  ;
	input \rf_conf11_reg[4]/NET0131  ;
	input \rf_conf11_reg[5]/NET0131  ;
	input \rf_conf11_reg[6]/NET0131  ;
	input \rf_conf11_reg[7]/NET0131  ;
	input \rf_conf11_reg[8]/NET0131  ;
	input \rf_conf11_reg[9]/NET0131  ;
	input \rf_conf12_reg[0]/NET0131  ;
	input \rf_conf12_reg[10]/NET0131  ;
	input \rf_conf12_reg[11]/NET0131  ;
	input \rf_conf12_reg[12]/NET0131  ;
	input \rf_conf12_reg[13]/NET0131  ;
	input \rf_conf12_reg[14]/NET0131  ;
	input \rf_conf12_reg[15]/NET0131  ;
	input \rf_conf12_reg[1]/NET0131  ;
	input \rf_conf12_reg[2]/NET0131  ;
	input \rf_conf12_reg[3]/NET0131  ;
	input \rf_conf12_reg[4]/NET0131  ;
	input \rf_conf12_reg[5]/NET0131  ;
	input \rf_conf12_reg[6]/NET0131  ;
	input \rf_conf12_reg[7]/NET0131  ;
	input \rf_conf12_reg[8]/NET0131  ;
	input \rf_conf12_reg[9]/NET0131  ;
	input \rf_conf13_reg[0]/NET0131  ;
	input \rf_conf13_reg[10]/NET0131  ;
	input \rf_conf13_reg[11]/NET0131  ;
	input \rf_conf13_reg[12]/NET0131  ;
	input \rf_conf13_reg[13]/NET0131  ;
	input \rf_conf13_reg[14]/NET0131  ;
	input \rf_conf13_reg[15]/NET0131  ;
	input \rf_conf13_reg[1]/NET0131  ;
	input \rf_conf13_reg[2]/NET0131  ;
	input \rf_conf13_reg[3]/NET0131  ;
	input \rf_conf13_reg[4]/NET0131  ;
	input \rf_conf13_reg[5]/NET0131  ;
	input \rf_conf13_reg[6]/NET0131  ;
	input \rf_conf13_reg[7]/NET0131  ;
	input \rf_conf13_reg[8]/NET0131  ;
	input \rf_conf13_reg[9]/NET0131  ;
	input \rf_conf14_reg[0]/NET0131  ;
	input \rf_conf14_reg[10]/NET0131  ;
	input \rf_conf14_reg[11]/NET0131  ;
	input \rf_conf14_reg[12]/NET0131  ;
	input \rf_conf14_reg[13]/NET0131  ;
	input \rf_conf14_reg[14]/NET0131  ;
	input \rf_conf14_reg[15]/NET0131  ;
	input \rf_conf14_reg[1]/NET0131  ;
	input \rf_conf14_reg[2]/NET0131  ;
	input \rf_conf14_reg[3]/NET0131  ;
	input \rf_conf14_reg[4]/NET0131  ;
	input \rf_conf14_reg[5]/NET0131  ;
	input \rf_conf14_reg[6]/NET0131  ;
	input \rf_conf14_reg[7]/NET0131  ;
	input \rf_conf14_reg[8]/NET0131  ;
	input \rf_conf14_reg[9]/NET0131  ;
	input \rf_conf15_reg[0]/NET0131  ;
	input \rf_conf15_reg[10]/NET0131  ;
	input \rf_conf15_reg[11]/NET0131  ;
	input \rf_conf15_reg[12]/NET0131  ;
	input \rf_conf15_reg[13]/NET0131  ;
	input \rf_conf15_reg[14]/NET0131  ;
	input \rf_conf15_reg[15]/NET0131  ;
	input \rf_conf15_reg[1]/NET0131  ;
	input \rf_conf15_reg[2]/NET0131  ;
	input \rf_conf15_reg[3]/NET0131  ;
	input \rf_conf15_reg[4]/NET0131  ;
	input \rf_conf15_reg[5]/NET0131  ;
	input \rf_conf15_reg[6]/NET0131  ;
	input \rf_conf15_reg[7]/NET0131  ;
	input \rf_conf15_reg[8]/NET0131  ;
	input \rf_conf15_reg[9]/NET0131  ;
	input \rf_conf1_reg[0]/NET0131  ;
	input \rf_conf1_reg[10]/NET0131  ;
	input \rf_conf1_reg[11]/NET0131  ;
	input \rf_conf1_reg[12]/NET0131  ;
	input \rf_conf1_reg[13]/NET0131  ;
	input \rf_conf1_reg[14]/NET0131  ;
	input \rf_conf1_reg[15]/NET0131  ;
	input \rf_conf1_reg[1]/NET0131  ;
	input \rf_conf1_reg[2]/NET0131  ;
	input \rf_conf1_reg[3]/NET0131  ;
	input \rf_conf1_reg[4]/NET0131  ;
	input \rf_conf1_reg[5]/NET0131  ;
	input \rf_conf1_reg[6]/NET0131  ;
	input \rf_conf1_reg[7]/NET0131  ;
	input \rf_conf1_reg[8]/NET0131  ;
	input \rf_conf1_reg[9]/NET0131  ;
	input \rf_conf2_reg[0]/NET0131  ;
	input \rf_conf2_reg[10]/NET0131  ;
	input \rf_conf2_reg[11]/NET0131  ;
	input \rf_conf2_reg[12]/NET0131  ;
	input \rf_conf2_reg[13]/NET0131  ;
	input \rf_conf2_reg[14]/NET0131  ;
	input \rf_conf2_reg[15]/NET0131  ;
	input \rf_conf2_reg[1]/NET0131  ;
	input \rf_conf2_reg[2]/NET0131  ;
	input \rf_conf2_reg[3]/NET0131  ;
	input \rf_conf2_reg[4]/NET0131  ;
	input \rf_conf2_reg[5]/NET0131  ;
	input \rf_conf2_reg[6]/NET0131  ;
	input \rf_conf2_reg[7]/NET0131  ;
	input \rf_conf2_reg[8]/NET0131  ;
	input \rf_conf2_reg[9]/NET0131  ;
	input \rf_conf3_reg[0]/NET0131  ;
	input \rf_conf3_reg[10]/NET0131  ;
	input \rf_conf3_reg[11]/NET0131  ;
	input \rf_conf3_reg[12]/NET0131  ;
	input \rf_conf3_reg[13]/NET0131  ;
	input \rf_conf3_reg[14]/NET0131  ;
	input \rf_conf3_reg[15]/NET0131  ;
	input \rf_conf3_reg[1]/NET0131  ;
	input \rf_conf3_reg[2]/NET0131  ;
	input \rf_conf3_reg[3]/NET0131  ;
	input \rf_conf3_reg[4]/NET0131  ;
	input \rf_conf3_reg[5]/NET0131  ;
	input \rf_conf3_reg[6]/NET0131  ;
	input \rf_conf3_reg[7]/NET0131  ;
	input \rf_conf3_reg[8]/NET0131  ;
	input \rf_conf3_reg[9]/NET0131  ;
	input \rf_conf4_reg[0]/NET0131  ;
	input \rf_conf4_reg[10]/NET0131  ;
	input \rf_conf4_reg[11]/NET0131  ;
	input \rf_conf4_reg[12]/NET0131  ;
	input \rf_conf4_reg[13]/NET0131  ;
	input \rf_conf4_reg[14]/NET0131  ;
	input \rf_conf4_reg[15]/NET0131  ;
	input \rf_conf4_reg[1]/NET0131  ;
	input \rf_conf4_reg[2]/NET0131  ;
	input \rf_conf4_reg[3]/NET0131  ;
	input \rf_conf4_reg[4]/NET0131  ;
	input \rf_conf4_reg[5]/NET0131  ;
	input \rf_conf4_reg[6]/NET0131  ;
	input \rf_conf4_reg[7]/NET0131  ;
	input \rf_conf4_reg[8]/NET0131  ;
	input \rf_conf4_reg[9]/NET0131  ;
	input \rf_conf5_reg[0]/NET0131  ;
	input \rf_conf5_reg[10]/NET0131  ;
	input \rf_conf5_reg[11]/NET0131  ;
	input \rf_conf5_reg[12]/NET0131  ;
	input \rf_conf5_reg[13]/NET0131  ;
	input \rf_conf5_reg[14]/NET0131  ;
	input \rf_conf5_reg[15]/NET0131  ;
	input \rf_conf5_reg[1]/NET0131  ;
	input \rf_conf5_reg[2]/NET0131  ;
	input \rf_conf5_reg[3]/NET0131  ;
	input \rf_conf5_reg[4]/NET0131  ;
	input \rf_conf5_reg[5]/NET0131  ;
	input \rf_conf5_reg[6]/NET0131  ;
	input \rf_conf5_reg[7]/NET0131  ;
	input \rf_conf5_reg[8]/NET0131  ;
	input \rf_conf5_reg[9]/NET0131  ;
	input \rf_conf6_reg[0]/NET0131  ;
	input \rf_conf6_reg[10]/NET0131  ;
	input \rf_conf6_reg[11]/NET0131  ;
	input \rf_conf6_reg[12]/NET0131  ;
	input \rf_conf6_reg[13]/NET0131  ;
	input \rf_conf6_reg[14]/NET0131  ;
	input \rf_conf6_reg[15]/NET0131  ;
	input \rf_conf6_reg[1]/NET0131  ;
	input \rf_conf6_reg[2]/NET0131  ;
	input \rf_conf6_reg[3]/NET0131  ;
	input \rf_conf6_reg[4]/NET0131  ;
	input \rf_conf6_reg[5]/NET0131  ;
	input \rf_conf6_reg[6]/NET0131  ;
	input \rf_conf6_reg[7]/NET0131  ;
	input \rf_conf6_reg[8]/NET0131  ;
	input \rf_conf6_reg[9]/NET0131  ;
	input \rf_conf7_reg[0]/NET0131  ;
	input \rf_conf7_reg[10]/NET0131  ;
	input \rf_conf7_reg[11]/NET0131  ;
	input \rf_conf7_reg[12]/NET0131  ;
	input \rf_conf7_reg[13]/NET0131  ;
	input \rf_conf7_reg[14]/NET0131  ;
	input \rf_conf7_reg[15]/NET0131  ;
	input \rf_conf7_reg[1]/NET0131  ;
	input \rf_conf7_reg[2]/NET0131  ;
	input \rf_conf7_reg[3]/NET0131  ;
	input \rf_conf7_reg[4]/NET0131  ;
	input \rf_conf7_reg[5]/NET0131  ;
	input \rf_conf7_reg[6]/NET0131  ;
	input \rf_conf7_reg[7]/NET0131  ;
	input \rf_conf7_reg[8]/NET0131  ;
	input \rf_conf7_reg[9]/NET0131  ;
	input \rf_conf8_reg[0]/NET0131  ;
	input \rf_conf8_reg[10]/NET0131  ;
	input \rf_conf8_reg[11]/NET0131  ;
	input \rf_conf8_reg[12]/NET0131  ;
	input \rf_conf8_reg[13]/NET0131  ;
	input \rf_conf8_reg[14]/NET0131  ;
	input \rf_conf8_reg[15]/NET0131  ;
	input \rf_conf8_reg[1]/NET0131  ;
	input \rf_conf8_reg[2]/NET0131  ;
	input \rf_conf8_reg[3]/NET0131  ;
	input \rf_conf8_reg[4]/NET0131  ;
	input \rf_conf8_reg[5]/NET0131  ;
	input \rf_conf8_reg[6]/NET0131  ;
	input \rf_conf8_reg[7]/NET0131  ;
	input \rf_conf8_reg[8]/NET0131  ;
	input \rf_conf8_reg[9]/NET0131  ;
	input \rf_conf9_reg[0]/NET0131  ;
	input \rf_conf9_reg[10]/NET0131  ;
	input \rf_conf9_reg[11]/NET0131  ;
	input \rf_conf9_reg[12]/NET0131  ;
	input \rf_conf9_reg[13]/NET0131  ;
	input \rf_conf9_reg[14]/NET0131  ;
	input \rf_conf9_reg[15]/NET0131  ;
	input \rf_conf9_reg[1]/NET0131  ;
	input \rf_conf9_reg[2]/NET0131  ;
	input \rf_conf9_reg[3]/NET0131  ;
	input \rf_conf9_reg[4]/NET0131  ;
	input \rf_conf9_reg[5]/NET0131  ;
	input \rf_conf9_reg[6]/NET0131  ;
	input \rf_conf9_reg[7]/NET0131  ;
	input \rf_conf9_reg[8]/NET0131  ;
	input \rf_conf9_reg[9]/NET0131  ;
	input \rf_rf_ack_reg/P0001  ;
	input \rf_rf_dout_reg[0]/P0001  ;
	input \rf_rf_dout_reg[10]/P0001  ;
	input \rf_rf_dout_reg[11]/P0001  ;
	input \rf_rf_dout_reg[12]/P0001  ;
	input \rf_rf_dout_reg[13]/P0001  ;
	input \rf_rf_dout_reg[14]/P0001  ;
	input \rf_rf_dout_reg[15]/P0001  ;
	input \rf_rf_dout_reg[1]/P0001  ;
	input \rf_rf_dout_reg[2]/P0001  ;
	input \rf_rf_dout_reg[3]/P0001  ;
	input \rf_rf_dout_reg[4]/P0001  ;
	input \rf_rf_dout_reg[5]/P0001  ;
	input \rf_rf_dout_reg[6]/P0001  ;
	input \rf_rf_dout_reg[7]/P0001  ;
	input \rf_rf_dout_reg[8]/P0001  ;
	input \rf_rf_dout_reg[9]/P0001  ;
	input \rf_rf_we_reg/P0001  ;
	input rst_i_pad ;
	input \s0_ack_i_pad  ;
	input \s0_data_i[0]_pad  ;
	input \s0_data_i[10]_pad  ;
	input \s0_data_i[11]_pad  ;
	input \s0_data_i[12]_pad  ;
	input \s0_data_i[13]_pad  ;
	input \s0_data_i[14]_pad  ;
	input \s0_data_i[15]_pad  ;
	input \s0_data_i[16]_pad  ;
	input \s0_data_i[17]_pad  ;
	input \s0_data_i[18]_pad  ;
	input \s0_data_i[19]_pad  ;
	input \s0_data_i[1]_pad  ;
	input \s0_data_i[20]_pad  ;
	input \s0_data_i[21]_pad  ;
	input \s0_data_i[22]_pad  ;
	input \s0_data_i[23]_pad  ;
	input \s0_data_i[24]_pad  ;
	input \s0_data_i[25]_pad  ;
	input \s0_data_i[26]_pad  ;
	input \s0_data_i[27]_pad  ;
	input \s0_data_i[28]_pad  ;
	input \s0_data_i[29]_pad  ;
	input \s0_data_i[2]_pad  ;
	input \s0_data_i[30]_pad  ;
	input \s0_data_i[31]_pad  ;
	input \s0_data_i[3]_pad  ;
	input \s0_data_i[4]_pad  ;
	input \s0_data_i[5]_pad  ;
	input \s0_data_i[6]_pad  ;
	input \s0_data_i[7]_pad  ;
	input \s0_data_i[8]_pad  ;
	input \s0_data_i[9]_pad  ;
	input \s0_err_i_pad  ;
	input \s0_m0_cyc_r_reg/P0001  ;
	input \s0_m1_cyc_r_reg/P0001  ;
	input \s0_m2_cyc_r_reg/P0001  ;
	input \s0_m3_cyc_r_reg/P0001  ;
	input \s0_m4_cyc_r_reg/P0001  ;
	input \s0_m5_cyc_r_reg/P0001  ;
	input \s0_m6_cyc_r_reg/P0001  ;
	input \s0_m7_cyc_r_reg/P0001  ;
	input \s0_msel_arb0_state_reg[0]/NET0131  ;
	input \s0_msel_arb0_state_reg[1]/NET0131  ;
	input \s0_msel_arb0_state_reg[2]/NET0131  ;
	input \s0_msel_arb1_state_reg[0]/NET0131  ;
	input \s0_msel_arb1_state_reg[1]/NET0131  ;
	input \s0_msel_arb1_state_reg[2]/NET0131  ;
	input \s0_msel_arb2_state_reg[0]/NET0131  ;
	input \s0_msel_arb2_state_reg[1]/NET0131  ;
	input \s0_msel_arb2_state_reg[2]/NET0131  ;
	input \s0_msel_arb3_state_reg[0]/NET0131  ;
	input \s0_msel_arb3_state_reg[1]/NET0131  ;
	input \s0_msel_arb3_state_reg[2]/NET0131  ;
	input \s0_msel_pri_out_reg[0]/NET0131  ;
	input \s0_msel_pri_out_reg[1]/NET0131  ;
	input \s0_next_reg/P0001  ;
	input \s0_rty_i_pad  ;
	input \s10_ack_i_pad  ;
	input \s10_data_i[0]_pad  ;
	input \s10_data_i[10]_pad  ;
	input \s10_data_i[11]_pad  ;
	input \s10_data_i[12]_pad  ;
	input \s10_data_i[13]_pad  ;
	input \s10_data_i[14]_pad  ;
	input \s10_data_i[15]_pad  ;
	input \s10_data_i[16]_pad  ;
	input \s10_data_i[17]_pad  ;
	input \s10_data_i[18]_pad  ;
	input \s10_data_i[19]_pad  ;
	input \s10_data_i[1]_pad  ;
	input \s10_data_i[20]_pad  ;
	input \s10_data_i[21]_pad  ;
	input \s10_data_i[22]_pad  ;
	input \s10_data_i[23]_pad  ;
	input \s10_data_i[24]_pad  ;
	input \s10_data_i[25]_pad  ;
	input \s10_data_i[26]_pad  ;
	input \s10_data_i[27]_pad  ;
	input \s10_data_i[28]_pad  ;
	input \s10_data_i[29]_pad  ;
	input \s10_data_i[2]_pad  ;
	input \s10_data_i[30]_pad  ;
	input \s10_data_i[31]_pad  ;
	input \s10_data_i[3]_pad  ;
	input \s10_data_i[4]_pad  ;
	input \s10_data_i[5]_pad  ;
	input \s10_data_i[6]_pad  ;
	input \s10_data_i[7]_pad  ;
	input \s10_data_i[8]_pad  ;
	input \s10_data_i[9]_pad  ;
	input \s10_err_i_pad  ;
	input \s10_m0_cyc_r_reg/P0001  ;
	input \s10_m1_cyc_r_reg/P0001  ;
	input \s10_m2_cyc_r_reg/P0001  ;
	input \s10_m3_cyc_r_reg/P0001  ;
	input \s10_m4_cyc_r_reg/P0001  ;
	input \s10_m5_cyc_r_reg/P0001  ;
	input \s10_m6_cyc_r_reg/P0001  ;
	input \s10_m7_cyc_r_reg/P0001  ;
	input \s10_msel_arb0_state_reg[0]/NET0131  ;
	input \s10_msel_arb0_state_reg[1]/NET0131  ;
	input \s10_msel_arb0_state_reg[2]/NET0131  ;
	input \s10_msel_arb1_state_reg[0]/NET0131  ;
	input \s10_msel_arb1_state_reg[1]/NET0131  ;
	input \s10_msel_arb1_state_reg[2]/NET0131  ;
	input \s10_msel_arb2_state_reg[0]/NET0131  ;
	input \s10_msel_arb2_state_reg[1]/NET0131  ;
	input \s10_msel_arb2_state_reg[2]/NET0131  ;
	input \s10_msel_arb3_state_reg[0]/NET0131  ;
	input \s10_msel_arb3_state_reg[1]/NET0131  ;
	input \s10_msel_arb3_state_reg[2]/NET0131  ;
	input \s10_msel_pri_out_reg[0]/NET0131  ;
	input \s10_msel_pri_out_reg[1]/NET0131  ;
	input \s10_next_reg/P0001  ;
	input \s10_rty_i_pad  ;
	input \s11_ack_i_pad  ;
	input \s11_data_i[0]_pad  ;
	input \s11_data_i[10]_pad  ;
	input \s11_data_i[11]_pad  ;
	input \s11_data_i[12]_pad  ;
	input \s11_data_i[13]_pad  ;
	input \s11_data_i[14]_pad  ;
	input \s11_data_i[15]_pad  ;
	input \s11_data_i[16]_pad  ;
	input \s11_data_i[17]_pad  ;
	input \s11_data_i[18]_pad  ;
	input \s11_data_i[19]_pad  ;
	input \s11_data_i[1]_pad  ;
	input \s11_data_i[20]_pad  ;
	input \s11_data_i[21]_pad  ;
	input \s11_data_i[22]_pad  ;
	input \s11_data_i[23]_pad  ;
	input \s11_data_i[24]_pad  ;
	input \s11_data_i[25]_pad  ;
	input \s11_data_i[26]_pad  ;
	input \s11_data_i[27]_pad  ;
	input \s11_data_i[28]_pad  ;
	input \s11_data_i[29]_pad  ;
	input \s11_data_i[2]_pad  ;
	input \s11_data_i[30]_pad  ;
	input \s11_data_i[31]_pad  ;
	input \s11_data_i[3]_pad  ;
	input \s11_data_i[4]_pad  ;
	input \s11_data_i[5]_pad  ;
	input \s11_data_i[6]_pad  ;
	input \s11_data_i[7]_pad  ;
	input \s11_data_i[8]_pad  ;
	input \s11_data_i[9]_pad  ;
	input \s11_err_i_pad  ;
	input \s11_m0_cyc_r_reg/P0001  ;
	input \s11_m1_cyc_r_reg/P0001  ;
	input \s11_m2_cyc_r_reg/P0001  ;
	input \s11_m3_cyc_r_reg/P0001  ;
	input \s11_m4_cyc_r_reg/P0001  ;
	input \s11_m5_cyc_r_reg/P0001  ;
	input \s11_m6_cyc_r_reg/P0001  ;
	input \s11_m7_cyc_r_reg/P0001  ;
	input \s11_msel_arb0_state_reg[0]/NET0131  ;
	input \s11_msel_arb0_state_reg[1]/NET0131  ;
	input \s11_msel_arb0_state_reg[2]/NET0131  ;
	input \s11_msel_arb1_state_reg[0]/NET0131  ;
	input \s11_msel_arb1_state_reg[1]/NET0131  ;
	input \s11_msel_arb1_state_reg[2]/NET0131  ;
	input \s11_msel_arb2_state_reg[0]/NET0131  ;
	input \s11_msel_arb2_state_reg[1]/NET0131  ;
	input \s11_msel_arb2_state_reg[2]/NET0131  ;
	input \s11_msel_arb3_state_reg[0]/NET0131  ;
	input \s11_msel_arb3_state_reg[1]/NET0131  ;
	input \s11_msel_arb3_state_reg[2]/NET0131  ;
	input \s11_msel_pri_out_reg[0]/NET0131  ;
	input \s11_msel_pri_out_reg[1]/NET0131  ;
	input \s11_next_reg/P0001  ;
	input \s11_rty_i_pad  ;
	input \s12_ack_i_pad  ;
	input \s12_data_i[0]_pad  ;
	input \s12_data_i[10]_pad  ;
	input \s12_data_i[11]_pad  ;
	input \s12_data_i[12]_pad  ;
	input \s12_data_i[13]_pad  ;
	input \s12_data_i[14]_pad  ;
	input \s12_data_i[15]_pad  ;
	input \s12_data_i[16]_pad  ;
	input \s12_data_i[17]_pad  ;
	input \s12_data_i[18]_pad  ;
	input \s12_data_i[19]_pad  ;
	input \s12_data_i[1]_pad  ;
	input \s12_data_i[20]_pad  ;
	input \s12_data_i[21]_pad  ;
	input \s12_data_i[22]_pad  ;
	input \s12_data_i[23]_pad  ;
	input \s12_data_i[24]_pad  ;
	input \s12_data_i[25]_pad  ;
	input \s12_data_i[26]_pad  ;
	input \s12_data_i[27]_pad  ;
	input \s12_data_i[28]_pad  ;
	input \s12_data_i[29]_pad  ;
	input \s12_data_i[2]_pad  ;
	input \s12_data_i[30]_pad  ;
	input \s12_data_i[31]_pad  ;
	input \s12_data_i[3]_pad  ;
	input \s12_data_i[4]_pad  ;
	input \s12_data_i[5]_pad  ;
	input \s12_data_i[6]_pad  ;
	input \s12_data_i[7]_pad  ;
	input \s12_data_i[8]_pad  ;
	input \s12_data_i[9]_pad  ;
	input \s12_err_i_pad  ;
	input \s12_m0_cyc_r_reg/P0001  ;
	input \s12_m1_cyc_r_reg/P0001  ;
	input \s12_m2_cyc_r_reg/P0001  ;
	input \s12_m3_cyc_r_reg/P0001  ;
	input \s12_m4_cyc_r_reg/P0001  ;
	input \s12_m5_cyc_r_reg/P0001  ;
	input \s12_m6_cyc_r_reg/P0001  ;
	input \s12_m7_cyc_r_reg/P0001  ;
	input \s12_msel_arb0_state_reg[0]/NET0131  ;
	input \s12_msel_arb0_state_reg[1]/NET0131  ;
	input \s12_msel_arb0_state_reg[2]/NET0131  ;
	input \s12_msel_arb1_state_reg[0]/NET0131  ;
	input \s12_msel_arb1_state_reg[1]/NET0131  ;
	input \s12_msel_arb1_state_reg[2]/NET0131  ;
	input \s12_msel_arb2_state_reg[0]/NET0131  ;
	input \s12_msel_arb2_state_reg[1]/NET0131  ;
	input \s12_msel_arb2_state_reg[2]/NET0131  ;
	input \s12_msel_arb3_state_reg[0]/NET0131  ;
	input \s12_msel_arb3_state_reg[1]/NET0131  ;
	input \s12_msel_arb3_state_reg[2]/NET0131  ;
	input \s12_msel_pri_out_reg[0]/NET0131  ;
	input \s12_msel_pri_out_reg[1]/NET0131  ;
	input \s12_next_reg/P0001  ;
	input \s12_rty_i_pad  ;
	input \s13_ack_i_pad  ;
	input \s13_data_i[0]_pad  ;
	input \s13_data_i[10]_pad  ;
	input \s13_data_i[11]_pad  ;
	input \s13_data_i[12]_pad  ;
	input \s13_data_i[13]_pad  ;
	input \s13_data_i[14]_pad  ;
	input \s13_data_i[15]_pad  ;
	input \s13_data_i[16]_pad  ;
	input \s13_data_i[17]_pad  ;
	input \s13_data_i[18]_pad  ;
	input \s13_data_i[19]_pad  ;
	input \s13_data_i[1]_pad  ;
	input \s13_data_i[20]_pad  ;
	input \s13_data_i[21]_pad  ;
	input \s13_data_i[22]_pad  ;
	input \s13_data_i[23]_pad  ;
	input \s13_data_i[24]_pad  ;
	input \s13_data_i[25]_pad  ;
	input \s13_data_i[26]_pad  ;
	input \s13_data_i[27]_pad  ;
	input \s13_data_i[28]_pad  ;
	input \s13_data_i[29]_pad  ;
	input \s13_data_i[2]_pad  ;
	input \s13_data_i[30]_pad  ;
	input \s13_data_i[31]_pad  ;
	input \s13_data_i[3]_pad  ;
	input \s13_data_i[4]_pad  ;
	input \s13_data_i[5]_pad  ;
	input \s13_data_i[6]_pad  ;
	input \s13_data_i[7]_pad  ;
	input \s13_data_i[8]_pad  ;
	input \s13_data_i[9]_pad  ;
	input \s13_err_i_pad  ;
	input \s13_m0_cyc_r_reg/P0001  ;
	input \s13_m1_cyc_r_reg/P0001  ;
	input \s13_m2_cyc_r_reg/P0001  ;
	input \s13_m3_cyc_r_reg/P0001  ;
	input \s13_m4_cyc_r_reg/P0001  ;
	input \s13_m5_cyc_r_reg/P0001  ;
	input \s13_m6_cyc_r_reg/P0001  ;
	input \s13_m7_cyc_r_reg/P0001  ;
	input \s13_msel_arb0_state_reg[0]/NET0131  ;
	input \s13_msel_arb0_state_reg[1]/NET0131  ;
	input \s13_msel_arb0_state_reg[2]/NET0131  ;
	input \s13_msel_arb1_state_reg[0]/NET0131  ;
	input \s13_msel_arb1_state_reg[1]/NET0131  ;
	input \s13_msel_arb1_state_reg[2]/NET0131  ;
	input \s13_msel_arb2_state_reg[0]/NET0131  ;
	input \s13_msel_arb2_state_reg[1]/NET0131  ;
	input \s13_msel_arb2_state_reg[2]/NET0131  ;
	input \s13_msel_arb3_state_reg[0]/NET0131  ;
	input \s13_msel_arb3_state_reg[1]/NET0131  ;
	input \s13_msel_arb3_state_reg[2]/NET0131  ;
	input \s13_msel_pri_out_reg[0]/NET0131  ;
	input \s13_msel_pri_out_reg[1]/NET0131  ;
	input \s13_next_reg/P0001  ;
	input \s13_rty_i_pad  ;
	input \s14_ack_i_pad  ;
	input \s14_data_i[0]_pad  ;
	input \s14_data_i[10]_pad  ;
	input \s14_data_i[11]_pad  ;
	input \s14_data_i[12]_pad  ;
	input \s14_data_i[13]_pad  ;
	input \s14_data_i[14]_pad  ;
	input \s14_data_i[15]_pad  ;
	input \s14_data_i[16]_pad  ;
	input \s14_data_i[17]_pad  ;
	input \s14_data_i[18]_pad  ;
	input \s14_data_i[19]_pad  ;
	input \s14_data_i[1]_pad  ;
	input \s14_data_i[20]_pad  ;
	input \s14_data_i[21]_pad  ;
	input \s14_data_i[22]_pad  ;
	input \s14_data_i[23]_pad  ;
	input \s14_data_i[24]_pad  ;
	input \s14_data_i[25]_pad  ;
	input \s14_data_i[26]_pad  ;
	input \s14_data_i[27]_pad  ;
	input \s14_data_i[28]_pad  ;
	input \s14_data_i[29]_pad  ;
	input \s14_data_i[2]_pad  ;
	input \s14_data_i[30]_pad  ;
	input \s14_data_i[31]_pad  ;
	input \s14_data_i[3]_pad  ;
	input \s14_data_i[4]_pad  ;
	input \s14_data_i[5]_pad  ;
	input \s14_data_i[6]_pad  ;
	input \s14_data_i[7]_pad  ;
	input \s14_data_i[8]_pad  ;
	input \s14_data_i[9]_pad  ;
	input \s14_err_i_pad  ;
	input \s14_m0_cyc_r_reg/P0001  ;
	input \s14_m1_cyc_r_reg/P0001  ;
	input \s14_m2_cyc_r_reg/P0001  ;
	input \s14_m3_cyc_r_reg/P0001  ;
	input \s14_m4_cyc_r_reg/P0001  ;
	input \s14_m5_cyc_r_reg/P0001  ;
	input \s14_m6_cyc_r_reg/P0001  ;
	input \s14_m7_cyc_r_reg/P0001  ;
	input \s14_msel_arb0_state_reg[0]/NET0131  ;
	input \s14_msel_arb0_state_reg[1]/NET0131  ;
	input \s14_msel_arb0_state_reg[2]/NET0131  ;
	input \s14_msel_arb1_state_reg[0]/NET0131  ;
	input \s14_msel_arb1_state_reg[1]/NET0131  ;
	input \s14_msel_arb1_state_reg[2]/NET0131  ;
	input \s14_msel_arb2_state_reg[0]/NET0131  ;
	input \s14_msel_arb2_state_reg[1]/NET0131  ;
	input \s14_msel_arb2_state_reg[2]/NET0131  ;
	input \s14_msel_arb3_state_reg[0]/NET0131  ;
	input \s14_msel_arb3_state_reg[1]/NET0131  ;
	input \s14_msel_arb3_state_reg[2]/NET0131  ;
	input \s14_msel_pri_out_reg[0]/NET0131  ;
	input \s14_msel_pri_out_reg[1]/NET0131  ;
	input \s14_next_reg/P0001  ;
	input \s14_rty_i_pad  ;
	input \s15_ack_i_pad  ;
	input \s15_data_i[0]_pad  ;
	input \s15_data_i[10]_pad  ;
	input \s15_data_i[11]_pad  ;
	input \s15_data_i[12]_pad  ;
	input \s15_data_i[13]_pad  ;
	input \s15_data_i[14]_pad  ;
	input \s15_data_i[15]_pad  ;
	input \s15_data_i[16]_pad  ;
	input \s15_data_i[17]_pad  ;
	input \s15_data_i[18]_pad  ;
	input \s15_data_i[19]_pad  ;
	input \s15_data_i[1]_pad  ;
	input \s15_data_i[20]_pad  ;
	input \s15_data_i[21]_pad  ;
	input \s15_data_i[22]_pad  ;
	input \s15_data_i[23]_pad  ;
	input \s15_data_i[24]_pad  ;
	input \s15_data_i[25]_pad  ;
	input \s15_data_i[26]_pad  ;
	input \s15_data_i[27]_pad  ;
	input \s15_data_i[28]_pad  ;
	input \s15_data_i[29]_pad  ;
	input \s15_data_i[2]_pad  ;
	input \s15_data_i[30]_pad  ;
	input \s15_data_i[31]_pad  ;
	input \s15_data_i[3]_pad  ;
	input \s15_data_i[4]_pad  ;
	input \s15_data_i[5]_pad  ;
	input \s15_data_i[6]_pad  ;
	input \s15_data_i[7]_pad  ;
	input \s15_data_i[8]_pad  ;
	input \s15_data_i[9]_pad  ;
	input \s15_err_i_pad  ;
	input \s15_m0_cyc_r_reg/P0001  ;
	input \s15_m1_cyc_r_reg/P0001  ;
	input \s15_m2_cyc_r_reg/P0001  ;
	input \s15_m3_cyc_r_reg/P0001  ;
	input \s15_m4_cyc_r_reg/P0001  ;
	input \s15_m5_cyc_r_reg/P0001  ;
	input \s15_m6_cyc_r_reg/P0001  ;
	input \s15_m7_cyc_r_reg/P0001  ;
	input \s15_msel_arb0_state_reg[0]/NET0131  ;
	input \s15_msel_arb0_state_reg[1]/NET0131  ;
	input \s15_msel_arb0_state_reg[2]/NET0131  ;
	input \s15_msel_arb1_state_reg[0]/NET0131  ;
	input \s15_msel_arb1_state_reg[1]/NET0131  ;
	input \s15_msel_arb1_state_reg[2]/NET0131  ;
	input \s15_msel_arb2_state_reg[0]/NET0131  ;
	input \s15_msel_arb2_state_reg[1]/NET0131  ;
	input \s15_msel_arb2_state_reg[2]/NET0131  ;
	input \s15_msel_arb3_state_reg[0]/NET0131  ;
	input \s15_msel_arb3_state_reg[1]/NET0131  ;
	input \s15_msel_arb3_state_reg[2]/NET0131  ;
	input \s15_msel_pri_out_reg[0]/NET0131  ;
	input \s15_msel_pri_out_reg[1]/NET0131  ;
	input \s15_next_reg/P0001  ;
	input \s15_rty_i_pad  ;
	input \s1_ack_i_pad  ;
	input \s1_data_i[0]_pad  ;
	input \s1_data_i[10]_pad  ;
	input \s1_data_i[11]_pad  ;
	input \s1_data_i[12]_pad  ;
	input \s1_data_i[13]_pad  ;
	input \s1_data_i[14]_pad  ;
	input \s1_data_i[15]_pad  ;
	input \s1_data_i[16]_pad  ;
	input \s1_data_i[17]_pad  ;
	input \s1_data_i[18]_pad  ;
	input \s1_data_i[19]_pad  ;
	input \s1_data_i[1]_pad  ;
	input \s1_data_i[20]_pad  ;
	input \s1_data_i[21]_pad  ;
	input \s1_data_i[22]_pad  ;
	input \s1_data_i[23]_pad  ;
	input \s1_data_i[24]_pad  ;
	input \s1_data_i[25]_pad  ;
	input \s1_data_i[26]_pad  ;
	input \s1_data_i[27]_pad  ;
	input \s1_data_i[28]_pad  ;
	input \s1_data_i[29]_pad  ;
	input \s1_data_i[2]_pad  ;
	input \s1_data_i[30]_pad  ;
	input \s1_data_i[31]_pad  ;
	input \s1_data_i[3]_pad  ;
	input \s1_data_i[4]_pad  ;
	input \s1_data_i[5]_pad  ;
	input \s1_data_i[6]_pad  ;
	input \s1_data_i[7]_pad  ;
	input \s1_data_i[8]_pad  ;
	input \s1_data_i[9]_pad  ;
	input \s1_err_i_pad  ;
	input \s1_m0_cyc_r_reg/P0001  ;
	input \s1_m1_cyc_r_reg/P0001  ;
	input \s1_m2_cyc_r_reg/P0001  ;
	input \s1_m3_cyc_r_reg/P0001  ;
	input \s1_m4_cyc_r_reg/P0001  ;
	input \s1_m5_cyc_r_reg/P0001  ;
	input \s1_m6_cyc_r_reg/P0001  ;
	input \s1_m7_cyc_r_reg/P0001  ;
	input \s1_msel_arb0_state_reg[0]/NET0131  ;
	input \s1_msel_arb0_state_reg[1]/NET0131  ;
	input \s1_msel_arb0_state_reg[2]/NET0131  ;
	input \s1_msel_arb1_state_reg[0]/NET0131  ;
	input \s1_msel_arb1_state_reg[1]/NET0131  ;
	input \s1_msel_arb1_state_reg[2]/NET0131  ;
	input \s1_msel_arb2_state_reg[0]/NET0131  ;
	input \s1_msel_arb2_state_reg[1]/NET0131  ;
	input \s1_msel_arb2_state_reg[2]/NET0131  ;
	input \s1_msel_arb3_state_reg[0]/NET0131  ;
	input \s1_msel_arb3_state_reg[1]/NET0131  ;
	input \s1_msel_arb3_state_reg[2]/NET0131  ;
	input \s1_msel_pri_out_reg[0]/NET0131  ;
	input \s1_msel_pri_out_reg[1]/NET0131  ;
	input \s1_next_reg/P0001  ;
	input \s1_rty_i_pad  ;
	input \s2_ack_i_pad  ;
	input \s2_data_i[0]_pad  ;
	input \s2_data_i[10]_pad  ;
	input \s2_data_i[11]_pad  ;
	input \s2_data_i[12]_pad  ;
	input \s2_data_i[13]_pad  ;
	input \s2_data_i[14]_pad  ;
	input \s2_data_i[15]_pad  ;
	input \s2_data_i[16]_pad  ;
	input \s2_data_i[17]_pad  ;
	input \s2_data_i[18]_pad  ;
	input \s2_data_i[19]_pad  ;
	input \s2_data_i[1]_pad  ;
	input \s2_data_i[20]_pad  ;
	input \s2_data_i[21]_pad  ;
	input \s2_data_i[22]_pad  ;
	input \s2_data_i[23]_pad  ;
	input \s2_data_i[24]_pad  ;
	input \s2_data_i[25]_pad  ;
	input \s2_data_i[26]_pad  ;
	input \s2_data_i[27]_pad  ;
	input \s2_data_i[28]_pad  ;
	input \s2_data_i[29]_pad  ;
	input \s2_data_i[2]_pad  ;
	input \s2_data_i[30]_pad  ;
	input \s2_data_i[31]_pad  ;
	input \s2_data_i[3]_pad  ;
	input \s2_data_i[4]_pad  ;
	input \s2_data_i[5]_pad  ;
	input \s2_data_i[6]_pad  ;
	input \s2_data_i[7]_pad  ;
	input \s2_data_i[8]_pad  ;
	input \s2_data_i[9]_pad  ;
	input \s2_err_i_pad  ;
	input \s2_m0_cyc_r_reg/P0001  ;
	input \s2_m1_cyc_r_reg/P0001  ;
	input \s2_m2_cyc_r_reg/P0001  ;
	input \s2_m3_cyc_r_reg/P0001  ;
	input \s2_m4_cyc_r_reg/P0001  ;
	input \s2_m5_cyc_r_reg/P0001  ;
	input \s2_m6_cyc_r_reg/P0001  ;
	input \s2_m7_cyc_r_reg/P0001  ;
	input \s2_msel_arb0_state_reg[0]/NET0131  ;
	input \s2_msel_arb0_state_reg[1]/NET0131  ;
	input \s2_msel_arb0_state_reg[2]/NET0131  ;
	input \s2_msel_arb1_state_reg[0]/NET0131  ;
	input \s2_msel_arb1_state_reg[1]/NET0131  ;
	input \s2_msel_arb1_state_reg[2]/NET0131  ;
	input \s2_msel_arb2_state_reg[0]/NET0131  ;
	input \s2_msel_arb2_state_reg[1]/NET0131  ;
	input \s2_msel_arb2_state_reg[2]/NET0131  ;
	input \s2_msel_arb3_state_reg[0]/NET0131  ;
	input \s2_msel_arb3_state_reg[1]/NET0131  ;
	input \s2_msel_arb3_state_reg[2]/NET0131  ;
	input \s2_msel_pri_out_reg[0]/NET0131  ;
	input \s2_msel_pri_out_reg[1]/NET0131  ;
	input \s2_next_reg/P0001  ;
	input \s2_rty_i_pad  ;
	input \s3_ack_i_pad  ;
	input \s3_data_i[0]_pad  ;
	input \s3_data_i[10]_pad  ;
	input \s3_data_i[11]_pad  ;
	input \s3_data_i[12]_pad  ;
	input \s3_data_i[13]_pad  ;
	input \s3_data_i[14]_pad  ;
	input \s3_data_i[15]_pad  ;
	input \s3_data_i[16]_pad  ;
	input \s3_data_i[17]_pad  ;
	input \s3_data_i[18]_pad  ;
	input \s3_data_i[19]_pad  ;
	input \s3_data_i[1]_pad  ;
	input \s3_data_i[20]_pad  ;
	input \s3_data_i[21]_pad  ;
	input \s3_data_i[22]_pad  ;
	input \s3_data_i[23]_pad  ;
	input \s3_data_i[24]_pad  ;
	input \s3_data_i[25]_pad  ;
	input \s3_data_i[26]_pad  ;
	input \s3_data_i[27]_pad  ;
	input \s3_data_i[28]_pad  ;
	input \s3_data_i[29]_pad  ;
	input \s3_data_i[2]_pad  ;
	input \s3_data_i[30]_pad  ;
	input \s3_data_i[31]_pad  ;
	input \s3_data_i[3]_pad  ;
	input \s3_data_i[4]_pad  ;
	input \s3_data_i[5]_pad  ;
	input \s3_data_i[6]_pad  ;
	input \s3_data_i[7]_pad  ;
	input \s3_data_i[8]_pad  ;
	input \s3_data_i[9]_pad  ;
	input \s3_err_i_pad  ;
	input \s3_m0_cyc_r_reg/P0001  ;
	input \s3_m1_cyc_r_reg/P0001  ;
	input \s3_m2_cyc_r_reg/P0001  ;
	input \s3_m3_cyc_r_reg/P0001  ;
	input \s3_m4_cyc_r_reg/P0001  ;
	input \s3_m5_cyc_r_reg/P0001  ;
	input \s3_m6_cyc_r_reg/P0001  ;
	input \s3_m7_cyc_r_reg/P0001  ;
	input \s3_msel_arb0_state_reg[0]/NET0131  ;
	input \s3_msel_arb0_state_reg[1]/NET0131  ;
	input \s3_msel_arb0_state_reg[2]/NET0131  ;
	input \s3_msel_arb1_state_reg[0]/NET0131  ;
	input \s3_msel_arb1_state_reg[1]/NET0131  ;
	input \s3_msel_arb1_state_reg[2]/NET0131  ;
	input \s3_msel_arb2_state_reg[0]/NET0131  ;
	input \s3_msel_arb2_state_reg[1]/NET0131  ;
	input \s3_msel_arb2_state_reg[2]/NET0131  ;
	input \s3_msel_arb3_state_reg[0]/NET0131  ;
	input \s3_msel_arb3_state_reg[1]/NET0131  ;
	input \s3_msel_arb3_state_reg[2]/NET0131  ;
	input \s3_msel_pri_out_reg[0]/NET0131  ;
	input \s3_msel_pri_out_reg[1]/NET0131  ;
	input \s3_next_reg/P0001  ;
	input \s3_rty_i_pad  ;
	input \s4_ack_i_pad  ;
	input \s4_data_i[0]_pad  ;
	input \s4_data_i[10]_pad  ;
	input \s4_data_i[11]_pad  ;
	input \s4_data_i[12]_pad  ;
	input \s4_data_i[13]_pad  ;
	input \s4_data_i[14]_pad  ;
	input \s4_data_i[15]_pad  ;
	input \s4_data_i[16]_pad  ;
	input \s4_data_i[17]_pad  ;
	input \s4_data_i[18]_pad  ;
	input \s4_data_i[19]_pad  ;
	input \s4_data_i[1]_pad  ;
	input \s4_data_i[20]_pad  ;
	input \s4_data_i[21]_pad  ;
	input \s4_data_i[22]_pad  ;
	input \s4_data_i[23]_pad  ;
	input \s4_data_i[24]_pad  ;
	input \s4_data_i[25]_pad  ;
	input \s4_data_i[26]_pad  ;
	input \s4_data_i[27]_pad  ;
	input \s4_data_i[28]_pad  ;
	input \s4_data_i[29]_pad  ;
	input \s4_data_i[2]_pad  ;
	input \s4_data_i[30]_pad  ;
	input \s4_data_i[31]_pad  ;
	input \s4_data_i[3]_pad  ;
	input \s4_data_i[4]_pad  ;
	input \s4_data_i[5]_pad  ;
	input \s4_data_i[6]_pad  ;
	input \s4_data_i[7]_pad  ;
	input \s4_data_i[8]_pad  ;
	input \s4_data_i[9]_pad  ;
	input \s4_err_i_pad  ;
	input \s4_m0_cyc_r_reg/P0001  ;
	input \s4_m1_cyc_r_reg/P0001  ;
	input \s4_m2_cyc_r_reg/P0001  ;
	input \s4_m3_cyc_r_reg/P0001  ;
	input \s4_m4_cyc_r_reg/P0001  ;
	input \s4_m5_cyc_r_reg/P0001  ;
	input \s4_m6_cyc_r_reg/P0001  ;
	input \s4_m7_cyc_r_reg/P0001  ;
	input \s4_msel_arb0_state_reg[0]/NET0131  ;
	input \s4_msel_arb0_state_reg[1]/NET0131  ;
	input \s4_msel_arb0_state_reg[2]/NET0131  ;
	input \s4_msel_arb1_state_reg[0]/NET0131  ;
	input \s4_msel_arb1_state_reg[1]/NET0131  ;
	input \s4_msel_arb1_state_reg[2]/NET0131  ;
	input \s4_msel_arb2_state_reg[0]/NET0131  ;
	input \s4_msel_arb2_state_reg[1]/NET0131  ;
	input \s4_msel_arb2_state_reg[2]/NET0131  ;
	input \s4_msel_arb3_state_reg[0]/NET0131  ;
	input \s4_msel_arb3_state_reg[1]/NET0131  ;
	input \s4_msel_arb3_state_reg[2]/NET0131  ;
	input \s4_msel_pri_out_reg[0]/NET0131  ;
	input \s4_msel_pri_out_reg[1]/NET0131  ;
	input \s4_next_reg/P0001  ;
	input \s4_rty_i_pad  ;
	input \s5_ack_i_pad  ;
	input \s5_data_i[0]_pad  ;
	input \s5_data_i[10]_pad  ;
	input \s5_data_i[11]_pad  ;
	input \s5_data_i[12]_pad  ;
	input \s5_data_i[13]_pad  ;
	input \s5_data_i[14]_pad  ;
	input \s5_data_i[15]_pad  ;
	input \s5_data_i[16]_pad  ;
	input \s5_data_i[17]_pad  ;
	input \s5_data_i[18]_pad  ;
	input \s5_data_i[19]_pad  ;
	input \s5_data_i[1]_pad  ;
	input \s5_data_i[20]_pad  ;
	input \s5_data_i[21]_pad  ;
	input \s5_data_i[22]_pad  ;
	input \s5_data_i[23]_pad  ;
	input \s5_data_i[24]_pad  ;
	input \s5_data_i[25]_pad  ;
	input \s5_data_i[26]_pad  ;
	input \s5_data_i[27]_pad  ;
	input \s5_data_i[28]_pad  ;
	input \s5_data_i[29]_pad  ;
	input \s5_data_i[2]_pad  ;
	input \s5_data_i[30]_pad  ;
	input \s5_data_i[31]_pad  ;
	input \s5_data_i[3]_pad  ;
	input \s5_data_i[4]_pad  ;
	input \s5_data_i[5]_pad  ;
	input \s5_data_i[6]_pad  ;
	input \s5_data_i[7]_pad  ;
	input \s5_data_i[8]_pad  ;
	input \s5_data_i[9]_pad  ;
	input \s5_err_i_pad  ;
	input \s5_m0_cyc_r_reg/P0001  ;
	input \s5_m1_cyc_r_reg/P0001  ;
	input \s5_m2_cyc_r_reg/P0001  ;
	input \s5_m3_cyc_r_reg/P0001  ;
	input \s5_m4_cyc_r_reg/P0001  ;
	input \s5_m5_cyc_r_reg/P0001  ;
	input \s5_m6_cyc_r_reg/P0001  ;
	input \s5_m7_cyc_r_reg/P0001  ;
	input \s5_msel_arb0_state_reg[0]/NET0131  ;
	input \s5_msel_arb0_state_reg[1]/NET0131  ;
	input \s5_msel_arb0_state_reg[2]/NET0131  ;
	input \s5_msel_arb1_state_reg[0]/NET0131  ;
	input \s5_msel_arb1_state_reg[1]/NET0131  ;
	input \s5_msel_arb1_state_reg[2]/NET0131  ;
	input \s5_msel_arb2_state_reg[0]/NET0131  ;
	input \s5_msel_arb2_state_reg[1]/NET0131  ;
	input \s5_msel_arb2_state_reg[2]/NET0131  ;
	input \s5_msel_arb3_state_reg[0]/NET0131  ;
	input \s5_msel_arb3_state_reg[1]/NET0131  ;
	input \s5_msel_arb3_state_reg[2]/NET0131  ;
	input \s5_msel_pri_out_reg[0]/NET0131  ;
	input \s5_msel_pri_out_reg[1]/NET0131  ;
	input \s5_next_reg/P0001  ;
	input \s5_rty_i_pad  ;
	input \s6_ack_i_pad  ;
	input \s6_data_i[0]_pad  ;
	input \s6_data_i[10]_pad  ;
	input \s6_data_i[11]_pad  ;
	input \s6_data_i[12]_pad  ;
	input \s6_data_i[13]_pad  ;
	input \s6_data_i[14]_pad  ;
	input \s6_data_i[15]_pad  ;
	input \s6_data_i[16]_pad  ;
	input \s6_data_i[17]_pad  ;
	input \s6_data_i[18]_pad  ;
	input \s6_data_i[19]_pad  ;
	input \s6_data_i[1]_pad  ;
	input \s6_data_i[20]_pad  ;
	input \s6_data_i[21]_pad  ;
	input \s6_data_i[22]_pad  ;
	input \s6_data_i[23]_pad  ;
	input \s6_data_i[24]_pad  ;
	input \s6_data_i[25]_pad  ;
	input \s6_data_i[26]_pad  ;
	input \s6_data_i[27]_pad  ;
	input \s6_data_i[28]_pad  ;
	input \s6_data_i[29]_pad  ;
	input \s6_data_i[2]_pad  ;
	input \s6_data_i[30]_pad  ;
	input \s6_data_i[31]_pad  ;
	input \s6_data_i[3]_pad  ;
	input \s6_data_i[4]_pad  ;
	input \s6_data_i[5]_pad  ;
	input \s6_data_i[6]_pad  ;
	input \s6_data_i[7]_pad  ;
	input \s6_data_i[8]_pad  ;
	input \s6_data_i[9]_pad  ;
	input \s6_err_i_pad  ;
	input \s6_m0_cyc_r_reg/P0001  ;
	input \s6_m1_cyc_r_reg/P0001  ;
	input \s6_m2_cyc_r_reg/P0001  ;
	input \s6_m3_cyc_r_reg/P0001  ;
	input \s6_m4_cyc_r_reg/P0001  ;
	input \s6_m5_cyc_r_reg/P0001  ;
	input \s6_m6_cyc_r_reg/P0001  ;
	input \s6_m7_cyc_r_reg/P0001  ;
	input \s6_msel_arb0_state_reg[0]/NET0131  ;
	input \s6_msel_arb0_state_reg[1]/NET0131  ;
	input \s6_msel_arb0_state_reg[2]/NET0131  ;
	input \s6_msel_arb1_state_reg[0]/NET0131  ;
	input \s6_msel_arb1_state_reg[1]/NET0131  ;
	input \s6_msel_arb1_state_reg[2]/NET0131  ;
	input \s6_msel_arb2_state_reg[0]/NET0131  ;
	input \s6_msel_arb2_state_reg[1]/NET0131  ;
	input \s6_msel_arb2_state_reg[2]/NET0131  ;
	input \s6_msel_arb3_state_reg[0]/NET0131  ;
	input \s6_msel_arb3_state_reg[1]/NET0131  ;
	input \s6_msel_arb3_state_reg[2]/NET0131  ;
	input \s6_msel_pri_out_reg[0]/NET0131  ;
	input \s6_msel_pri_out_reg[1]/NET0131  ;
	input \s6_next_reg/P0001  ;
	input \s6_rty_i_pad  ;
	input \s7_ack_i_pad  ;
	input \s7_data_i[0]_pad  ;
	input \s7_data_i[10]_pad  ;
	input \s7_data_i[11]_pad  ;
	input \s7_data_i[12]_pad  ;
	input \s7_data_i[13]_pad  ;
	input \s7_data_i[14]_pad  ;
	input \s7_data_i[15]_pad  ;
	input \s7_data_i[16]_pad  ;
	input \s7_data_i[17]_pad  ;
	input \s7_data_i[18]_pad  ;
	input \s7_data_i[19]_pad  ;
	input \s7_data_i[1]_pad  ;
	input \s7_data_i[20]_pad  ;
	input \s7_data_i[21]_pad  ;
	input \s7_data_i[22]_pad  ;
	input \s7_data_i[23]_pad  ;
	input \s7_data_i[24]_pad  ;
	input \s7_data_i[25]_pad  ;
	input \s7_data_i[26]_pad  ;
	input \s7_data_i[27]_pad  ;
	input \s7_data_i[28]_pad  ;
	input \s7_data_i[29]_pad  ;
	input \s7_data_i[2]_pad  ;
	input \s7_data_i[30]_pad  ;
	input \s7_data_i[31]_pad  ;
	input \s7_data_i[3]_pad  ;
	input \s7_data_i[4]_pad  ;
	input \s7_data_i[5]_pad  ;
	input \s7_data_i[6]_pad  ;
	input \s7_data_i[7]_pad  ;
	input \s7_data_i[8]_pad  ;
	input \s7_data_i[9]_pad  ;
	input \s7_err_i_pad  ;
	input \s7_m0_cyc_r_reg/P0001  ;
	input \s7_m1_cyc_r_reg/P0001  ;
	input \s7_m2_cyc_r_reg/P0001  ;
	input \s7_m3_cyc_r_reg/P0001  ;
	input \s7_m4_cyc_r_reg/P0001  ;
	input \s7_m5_cyc_r_reg/P0001  ;
	input \s7_m6_cyc_r_reg/P0001  ;
	input \s7_m7_cyc_r_reg/P0001  ;
	input \s7_msel_arb0_state_reg[0]/NET0131  ;
	input \s7_msel_arb0_state_reg[1]/NET0131  ;
	input \s7_msel_arb0_state_reg[2]/NET0131  ;
	input \s7_msel_arb1_state_reg[0]/NET0131  ;
	input \s7_msel_arb1_state_reg[1]/NET0131  ;
	input \s7_msel_arb1_state_reg[2]/NET0131  ;
	input \s7_msel_arb2_state_reg[0]/NET0131  ;
	input \s7_msel_arb2_state_reg[1]/NET0131  ;
	input \s7_msel_arb2_state_reg[2]/NET0131  ;
	input \s7_msel_arb3_state_reg[0]/NET0131  ;
	input \s7_msel_arb3_state_reg[1]/NET0131  ;
	input \s7_msel_arb3_state_reg[2]/NET0131  ;
	input \s7_msel_pri_out_reg[0]/NET0131  ;
	input \s7_msel_pri_out_reg[1]/NET0131  ;
	input \s7_next_reg/P0001  ;
	input \s7_rty_i_pad  ;
	input \s8_ack_i_pad  ;
	input \s8_data_i[0]_pad  ;
	input \s8_data_i[10]_pad  ;
	input \s8_data_i[11]_pad  ;
	input \s8_data_i[12]_pad  ;
	input \s8_data_i[13]_pad  ;
	input \s8_data_i[14]_pad  ;
	input \s8_data_i[15]_pad  ;
	input \s8_data_i[16]_pad  ;
	input \s8_data_i[17]_pad  ;
	input \s8_data_i[18]_pad  ;
	input \s8_data_i[19]_pad  ;
	input \s8_data_i[1]_pad  ;
	input \s8_data_i[20]_pad  ;
	input \s8_data_i[21]_pad  ;
	input \s8_data_i[22]_pad  ;
	input \s8_data_i[23]_pad  ;
	input \s8_data_i[24]_pad  ;
	input \s8_data_i[25]_pad  ;
	input \s8_data_i[26]_pad  ;
	input \s8_data_i[27]_pad  ;
	input \s8_data_i[28]_pad  ;
	input \s8_data_i[29]_pad  ;
	input \s8_data_i[2]_pad  ;
	input \s8_data_i[30]_pad  ;
	input \s8_data_i[31]_pad  ;
	input \s8_data_i[3]_pad  ;
	input \s8_data_i[4]_pad  ;
	input \s8_data_i[5]_pad  ;
	input \s8_data_i[6]_pad  ;
	input \s8_data_i[7]_pad  ;
	input \s8_data_i[8]_pad  ;
	input \s8_data_i[9]_pad  ;
	input \s8_err_i_pad  ;
	input \s8_m0_cyc_r_reg/P0001  ;
	input \s8_m1_cyc_r_reg/P0001  ;
	input \s8_m2_cyc_r_reg/P0001  ;
	input \s8_m3_cyc_r_reg/P0001  ;
	input \s8_m4_cyc_r_reg/P0001  ;
	input \s8_m5_cyc_r_reg/P0001  ;
	input \s8_m6_cyc_r_reg/P0001  ;
	input \s8_m7_cyc_r_reg/P0001  ;
	input \s8_msel_arb0_state_reg[0]/NET0131  ;
	input \s8_msel_arb0_state_reg[1]/NET0131  ;
	input \s8_msel_arb0_state_reg[2]/NET0131  ;
	input \s8_msel_arb1_state_reg[0]/NET0131  ;
	input \s8_msel_arb1_state_reg[1]/NET0131  ;
	input \s8_msel_arb1_state_reg[2]/NET0131  ;
	input \s8_msel_arb2_state_reg[0]/NET0131  ;
	input \s8_msel_arb2_state_reg[1]/NET0131  ;
	input \s8_msel_arb2_state_reg[2]/NET0131  ;
	input \s8_msel_arb3_state_reg[0]/NET0131  ;
	input \s8_msel_arb3_state_reg[1]/NET0131  ;
	input \s8_msel_arb3_state_reg[2]/NET0131  ;
	input \s8_msel_pri_out_reg[0]/NET0131  ;
	input \s8_msel_pri_out_reg[1]/NET0131  ;
	input \s8_next_reg/P0001  ;
	input \s8_rty_i_pad  ;
	input \s9_ack_i_pad  ;
	input \s9_data_i[0]_pad  ;
	input \s9_data_i[10]_pad  ;
	input \s9_data_i[11]_pad  ;
	input \s9_data_i[12]_pad  ;
	input \s9_data_i[13]_pad  ;
	input \s9_data_i[14]_pad  ;
	input \s9_data_i[15]_pad  ;
	input \s9_data_i[16]_pad  ;
	input \s9_data_i[17]_pad  ;
	input \s9_data_i[18]_pad  ;
	input \s9_data_i[19]_pad  ;
	input \s9_data_i[1]_pad  ;
	input \s9_data_i[20]_pad  ;
	input \s9_data_i[21]_pad  ;
	input \s9_data_i[22]_pad  ;
	input \s9_data_i[23]_pad  ;
	input \s9_data_i[24]_pad  ;
	input \s9_data_i[25]_pad  ;
	input \s9_data_i[26]_pad  ;
	input \s9_data_i[27]_pad  ;
	input \s9_data_i[28]_pad  ;
	input \s9_data_i[29]_pad  ;
	input \s9_data_i[2]_pad  ;
	input \s9_data_i[30]_pad  ;
	input \s9_data_i[31]_pad  ;
	input \s9_data_i[3]_pad  ;
	input \s9_data_i[4]_pad  ;
	input \s9_data_i[5]_pad  ;
	input \s9_data_i[6]_pad  ;
	input \s9_data_i[7]_pad  ;
	input \s9_data_i[8]_pad  ;
	input \s9_data_i[9]_pad  ;
	input \s9_err_i_pad  ;
	input \s9_m0_cyc_r_reg/P0001  ;
	input \s9_m1_cyc_r_reg/P0001  ;
	input \s9_m2_cyc_r_reg/P0001  ;
	input \s9_m3_cyc_r_reg/P0001  ;
	input \s9_m4_cyc_r_reg/P0001  ;
	input \s9_m5_cyc_r_reg/P0001  ;
	input \s9_m6_cyc_r_reg/P0001  ;
	input \s9_m7_cyc_r_reg/P0001  ;
	input \s9_msel_arb0_state_reg[0]/NET0131  ;
	input \s9_msel_arb0_state_reg[1]/NET0131  ;
	input \s9_msel_arb0_state_reg[2]/NET0131  ;
	input \s9_msel_arb1_state_reg[0]/NET0131  ;
	input \s9_msel_arb1_state_reg[1]/NET0131  ;
	input \s9_msel_arb1_state_reg[2]/NET0131  ;
	input \s9_msel_arb2_state_reg[0]/NET0131  ;
	input \s9_msel_arb2_state_reg[1]/NET0131  ;
	input \s9_msel_arb2_state_reg[2]/NET0131  ;
	input \s9_msel_arb3_state_reg[0]/NET0131  ;
	input \s9_msel_arb3_state_reg[1]/NET0131  ;
	input \s9_msel_arb3_state_reg[2]/NET0131  ;
	input \s9_msel_pri_out_reg[0]/NET0131  ;
	input \s9_msel_pri_out_reg[1]/NET0131  ;
	input \s9_next_reg/P0001  ;
	input \s9_rty_i_pad  ;
	output \_al_n0  ;
	output \_al_n1  ;
	output \g106655/_1_  ;
	output \g106703/_1_  ;
	output \g69412/_0_  ;
	output \g69413/_0_  ;
	output \g69417/_1_  ;
	output \g69418/_0_  ;
	output \g69420/_1_  ;
	output \g69421/_0_  ;
	output \g69423/_1_  ;
	output \g69424/_0_  ;
	output \g69426/_1_  ;
	output \g69428/_1_  ;
	output \g69430/_1_  ;
	output \g69432/_1_  ;
	output \g69434/_1_  ;
	output \g69436/_1_  ;
	output \g69438/_1_  ;
	output \g69757/_2_  ;
	output \g69758/_2_  ;
	output \g69759/_2_  ;
	output \g69760/_2_  ;
	output \g69761/_0_  ;
	output \g69762/_2_  ;
	output \g69763/_2_  ;
	output \g69764/_2_  ;
	output \g69765/_2_  ;
	output \g69766/_2_  ;
	output \g69767/_0_  ;
	output \g69768/_0_  ;
	output \g69769/_0_  ;
	output \g69770/_0_  ;
	output \g69771/_0_  ;
	output \g69772/_0_  ;
	output \g70206/_0_  ;
	output \g70392/_0_  ;
	output \g70393/_0_  ;
	output \g70394/_0_  ;
	output \g70395/_0_  ;
	output \g70396/_0_  ;
	output \g70397/_0_  ;
	output \g70398/_0_  ;
	output \g70399/_0_  ;
	output \g70400/_0_  ;
	output \g70401/_0_  ;
	output \g70402/_0_  ;
	output \g70403/_0_  ;
	output \g70404/_0_  ;
	output \g70405/_0_  ;
	output \g70406/_0_  ;
	output \g70407/_0_  ;
	output \g70408/_0_  ;
	output \g70409/_0_  ;
	output \g70410/_0_  ;
	output \g70411/_0_  ;
	output \g70412/_0_  ;
	output \g70413/_0_  ;
	output \g70414/_0_  ;
	output \g70415/_0_  ;
	output \g70416/_0_  ;
	output \g70417/_0_  ;
	output \g70418/_0_  ;
	output \g70419/_0_  ;
	output \g70420/_0_  ;
	output \g70421/_0_  ;
	output \g70422/_0_  ;
	output \g70423/_0_  ;
	output \g70424/_0_  ;
	output \g70425/_0_  ;
	output \g70426/_0_  ;
	output \g70427/_0_  ;
	output \g70428/_0_  ;
	output \g70429/_0_  ;
	output \g70430/_0_  ;
	output \g70431/_0_  ;
	output \g70432/_0_  ;
	output \g70433/_0_  ;
	output \g70434/_0_  ;
	output \g70435/_0_  ;
	output \g70436/_0_  ;
	output \g70437/_0_  ;
	output \g70438/_0_  ;
	output \g70439/_0_  ;
	output \g70440/_0_  ;
	output \g70441/_0_  ;
	output \g70442/_0_  ;
	output \g70443/_0_  ;
	output \g70444/_0_  ;
	output \g70445/_0_  ;
	output \g70446/_0_  ;
	output \g70447/_0_  ;
	output \g70448/_0_  ;
	output \g70449/_0_  ;
	output \g70450/_0_  ;
	output \g70451/_0_  ;
	output \g70452/_0_  ;
	output \g70453/_0_  ;
	output \g70454/_0_  ;
	output \g70455/_0_  ;
	output \g70456/_0_  ;
	output \g70457/_0_  ;
	output \g70458/_0_  ;
	output \g70459/_0_  ;
	output \g70460/_0_  ;
	output \g70461/_0_  ;
	output \g70462/_0_  ;
	output \g70463/_0_  ;
	output \g70464/_0_  ;
	output \g70465/_0_  ;
	output \g70466/_0_  ;
	output \g70467/_0_  ;
	output \g70468/_0_  ;
	output \g70469/_0_  ;
	output \g70470/_0_  ;
	output \g70471/_0_  ;
	output \g70472/_0_  ;
	output \g70473/_0_  ;
	output \g70474/_0_  ;
	output \g70475/_0_  ;
	output \g70476/_0_  ;
	output \g70477/_0_  ;
	output \g70478/_0_  ;
	output \g70479/_0_  ;
	output \g70480/_0_  ;
	output \g70481/_0_  ;
	output \g70482/_0_  ;
	output \g70483/_0_  ;
	output \g70484/_0_  ;
	output \g70485/_0_  ;
	output \g70486/_0_  ;
	output \g70487/_0_  ;
	output \g70488/_0_  ;
	output \g70489/_0_  ;
	output \g70490/_0_  ;
	output \g70491/_0_  ;
	output \g70492/_0_  ;
	output \g70493/_0_  ;
	output \g70494/_0_  ;
	output \g70495/_0_  ;
	output \g70496/_0_  ;
	output \g70497/_0_  ;
	output \g70498/_0_  ;
	output \g70499/_0_  ;
	output \g70500/_0_  ;
	output \g70501/_0_  ;
	output \g70502/_0_  ;
	output \g70503/_0_  ;
	output \g70504/_0_  ;
	output \g70505/_0_  ;
	output \g70506/_0_  ;
	output \g70507/_0_  ;
	output \g70508/_0_  ;
	output \g70509/_0_  ;
	output \g70510/_0_  ;
	output \g70511/_0_  ;
	output \g70513/_0_  ;
	output \g70515/_0_  ;
	output \g70516/_0_  ;
	output \g70517/_0_  ;
	output \g70518/_0_  ;
	output \g70519/_0_  ;
	output \g70521/_0_  ;
	output \g70522/_0_  ;
	output \g70524/_0_  ;
	output \g70557/_0_  ;
	output \g70559/_0_  ;
	output \g70560/_0_  ;
	output \g70561/_0_  ;
	output \g70562/_0_  ;
	output \g70563/_0_  ;
	output \g70564/_0_  ;
	output \g70565/_0_  ;
	output \g70566/_0_  ;
	output \g70567/_0_  ;
	output \g70568/_0_  ;
	output \g70569/_0_  ;
	output \g70570/_0_  ;
	output \g70571/_0_  ;
	output \g70572/_0_  ;
	output \g70573/_0_  ;
	output \g70574/_0_  ;
	output \g70575/_0_  ;
	output \g70576/_0_  ;
	output \g70577/_0_  ;
	output \g70578/_0_  ;
	output \g70579/_0_  ;
	output \g70580/_0_  ;
	output \g70581/_0_  ;
	output \g70582/_0_  ;
	output \g70583/_0_  ;
	output \g70584/_0_  ;
	output \g70585/_0_  ;
	output \g70586/_0_  ;
	output \g70587/_0_  ;
	output \g70588/_0_  ;
	output \g70589/_0_  ;
	output \g70590/_0_  ;
	output \g70591/_0_  ;
	output \g70592/_0_  ;
	output \g70593/_0_  ;
	output \g70594/_0_  ;
	output \g70595/_0_  ;
	output \g70596/_0_  ;
	output \g70597/_0_  ;
	output \g70598/_0_  ;
	output \g70599/_0_  ;
	output \g70600/_0_  ;
	output \g70601/_0_  ;
	output \g70602/_0_  ;
	output \g70603/_0_  ;
	output \g70604/_0_  ;
	output \g70605/_0_  ;
	output \g70606/_0_  ;
	output \g70607/_0_  ;
	output \g70608/_0_  ;
	output \g70609/_0_  ;
	output \g70610/_0_  ;
	output \g70611/_0_  ;
	output \g70612/_0_  ;
	output \g70613/_0_  ;
	output \g70614/_0_  ;
	output \g70615/_0_  ;
	output \g70616/_0_  ;
	output \g70617/_0_  ;
	output \g70618/_0_  ;
	output \g70619/_0_  ;
	output \g70620/_0_  ;
	output \g70621/_0_  ;
	output \g70622/_0_  ;
	output \g70623/_0_  ;
	output \g70624/_0_  ;
	output \g70625/_0_  ;
	output \g70626/_0_  ;
	output \g70627/_0_  ;
	output \g70628/_0_  ;
	output \g70629/_0_  ;
	output \g70630/_0_  ;
	output \g70631/_0_  ;
	output \g70632/_0_  ;
	output \g70633/_0_  ;
	output \g70634/_0_  ;
	output \g70635/_0_  ;
	output \g70636/_0_  ;
	output \g70637/_0_  ;
	output \g70638/_0_  ;
	output \g70639/_0_  ;
	output \g70640/_0_  ;
	output \g70641/_0_  ;
	output \g70642/_0_  ;
	output \g70643/_0_  ;
	output \g70644/_0_  ;
	output \g70645/_0_  ;
	output \g70646/_0_  ;
	output \g70647/_0_  ;
	output \g70648/_0_  ;
	output \g70649/_0_  ;
	output \g70650/_0_  ;
	output \g70651/_0_  ;
	output \g70652/_0_  ;
	output \g70653/_0_  ;
	output \g70654/_0_  ;
	output \g70655/_0_  ;
	output \g70656/_0_  ;
	output \g70657/_0_  ;
	output \g70658/_0_  ;
	output \g70659/_0_  ;
	output \g70660/_0_  ;
	output \g70661/_0_  ;
	output \g70662/_0_  ;
	output \g70663/_0_  ;
	output \g70664/_0_  ;
	output \g70665/_0_  ;
	output \g70666/_0_  ;
	output \g70667/_0_  ;
	output \g70668/_0_  ;
	output \g70669/_0_  ;
	output \g70670/_0_  ;
	output \g70671/_0_  ;
	output \g70672/_0_  ;
	output \g70673/_0_  ;
	output \g70674/_0_  ;
	output \g70675/_0_  ;
	output \g70676/_0_  ;
	output \g70677/_0_  ;
	output \g70678/_0_  ;
	output \g70679/_0_  ;
	output \g70680/_0_  ;
	output \g70681/_0_  ;
	output \g70682/_0_  ;
	output \g70683/_0_  ;
	output \g70684/_0_  ;
	output \g70685/_0_  ;
	output \g70686/_0_  ;
	output \g70687/_0_  ;
	output \g70688/_0_  ;
	output \g70689/_0_  ;
	output \g70690/_0_  ;
	output \g70691/_0_  ;
	output \g70692/_0_  ;
	output \g70693/_0_  ;
	output \g70694/_0_  ;
	output \g70695/_0_  ;
	output \g70696/_0_  ;
	output \g70697/_0_  ;
	output \g70698/_0_  ;
	output \g70699/_0_  ;
	output \g70700/_0_  ;
	output \g70701/_0_  ;
	output \g70702/_0_  ;
	output \g70703/_0_  ;
	output \g70704/_0_  ;
	output \g70705/_0_  ;
	output \g70706/_0_  ;
	output \g70707/_0_  ;
	output \g70708/_0_  ;
	output \g70709/_0_  ;
	output \g70710/_0_  ;
	output \g70711/_0_  ;
	output \g70712/_0_  ;
	output \g70713/_0_  ;
	output \g70714/_0_  ;
	output \g70715/_0_  ;
	output \g70716/_0_  ;
	output \g70717/_0_  ;
	output \g70718/_0_  ;
	output \g70719/_0_  ;
	output \g70720/_0_  ;
	output \g70721/_0_  ;
	output \g70722/_0_  ;
	output \g70723/_0_  ;
	output \g70724/_0_  ;
	output \g70725/_0_  ;
	output \g70726/_0_  ;
	output \g70727/_0_  ;
	output \g70728/_0_  ;
	output \g70729/_0_  ;
	output \g70730/_0_  ;
	output \g70731/_0_  ;
	output \g70732/_0_  ;
	output \g70733/_0_  ;
	output \g70734/_0_  ;
	output \g70735/_0_  ;
	output \g70736/_0_  ;
	output \g70737/_0_  ;
	output \g70738/_0_  ;
	output \g70739/_0_  ;
	output \g70740/_0_  ;
	output \g70741/_0_  ;
	output \g70742/_0_  ;
	output \g70743/_0_  ;
	output \g70744/_0_  ;
	output \g70745/_0_  ;
	output \g70746/_0_  ;
	output \g70747/_0_  ;
	output \g70748/_0_  ;
	output \g70749/_0_  ;
	output \g70750/_0_  ;
	output \g70751/_0_  ;
	output \g70752/_0_  ;
	output \g70753/_0_  ;
	output \g70754/_0_  ;
	output \g70755/_0_  ;
	output \g70756/_0_  ;
	output \g70757/_0_  ;
	output \g70758/_0_  ;
	output \g70759/_0_  ;
	output \g70760/_0_  ;
	output \g70761/_0_  ;
	output \g70762/_0_  ;
	output \g70763/_0_  ;
	output \g70764/_0_  ;
	output \g70765/_0_  ;
	output \g70766/_0_  ;
	output \g70767/_0_  ;
	output \g70768/_0_  ;
	output \g70769/_0_  ;
	output \g70770/_0_  ;
	output \g70771/_0_  ;
	output \g70772/_0_  ;
	output \g70773/_0_  ;
	output \g70774/_0_  ;
	output \g70775/_0_  ;
	output \g70776/_0_  ;
	output \g70777/_0_  ;
	output \g70778/_0_  ;
	output \g70779/_0_  ;
	output \g70780/_0_  ;
	output \g70781/_0_  ;
	output \g70782/_0_  ;
	output \g70783/_0_  ;
	output \g70784/_0_  ;
	output \g70785/_0_  ;
	output \g70786/_0_  ;
	output \g70787/_0_  ;
	output \g70788/_0_  ;
	output \g70789/_0_  ;
	output \g70790/_0_  ;
	output \g70791/_0_  ;
	output \g70792/_0_  ;
	output \g70793/_0_  ;
	output \g70794/_0_  ;
	output \g70795/_0_  ;
	output \g70796/_0_  ;
	output \g70797/_0_  ;
	output \g70798/_0_  ;
	output \g70799/_0_  ;
	output \g70800/_0_  ;
	output \g70801/_0_  ;
	output \g70802/_0_  ;
	output \g70803/_0_  ;
	output \g70804/_0_  ;
	output \g70805/_0_  ;
	output \g70806/_0_  ;
	output \g70807/_0_  ;
	output \g70808/_0_  ;
	output \g70809/_0_  ;
	output \g70810/_0_  ;
	output \g70811/_0_  ;
	output \g70812/_0_  ;
	output \g70813/_0_  ;
	output \g70814/_0_  ;
	output \g70815/_0_  ;
	output \g70816/_0_  ;
	output \g70817/_0_  ;
	output \g70818/_0_  ;
	output \g70819/_0_  ;
	output \g70820/_0_  ;
	output \g70821/_0_  ;
	output \g70822/_0_  ;
	output \g70823/_0_  ;
	output \g70824/_0_  ;
	output \g70825/_0_  ;
	output \g70826/_0_  ;
	output \g70827/_0_  ;
	output \g70828/_0_  ;
	output \g70829/_0_  ;
	output \g70830/_0_  ;
	output \g70831/_0_  ;
	output \g70832/_0_  ;
	output \g70833/_0_  ;
	output \g70834/_0_  ;
	output \g70835/_0_  ;
	output \g70836/_0_  ;
	output \g70837/_0_  ;
	output \g70838/_0_  ;
	output \g70839/_0_  ;
	output \g70840/_0_  ;
	output \g70841/_0_  ;
	output \g70842/_0_  ;
	output \g70843/_0_  ;
	output \g70844/_0_  ;
	output \g70845/_0_  ;
	output \g70846/_0_  ;
	output \g70847/_0_  ;
	output \g70848/_0_  ;
	output \g70849/_0_  ;
	output \g70850/_0_  ;
	output \g70851/_0_  ;
	output \g70852/_0_  ;
	output \g70853/_0_  ;
	output \g70854/_0_  ;
	output \g70855/_0_  ;
	output \g70856/_0_  ;
	output \g70857/_0_  ;
	output \g70858/_0_  ;
	output \g70859/_0_  ;
	output \g70860/_0_  ;
	output \g70861/_0_  ;
	output \g71404/_0_  ;
	output \g71407/_0_  ;
	output \g72631/_0_  ;
	output \g72631/_1_  ;
	output \g72633/_0_  ;
	output \g72642/_0_  ;
	output \g72649/_0_  ;
	output \g72649/_1_  ;
	output \g72652/_0_  ;
	output \g72660/_0_  ;
	output \g72666/_0_  ;
	output \g72666/_1_  ;
	output \g72671/_0_  ;
	output \g72681/_0_  ;
	output \g72681/_1_  ;
	output \g72689/_0_  ;
	output \g72696/_0_  ;
	output \g72696/_1_  ;
	output \g72698/_0_  ;
	output \g72707/_0_  ;
	output \g72715/_0_  ;
	output \g72715/_1_  ;
	output \g72718/_0_  ;
	output \g72726/_0_  ;
	output \g72732/_0_  ;
	output \g72732/_1_  ;
	output \g72736/_0_  ;
	output \g72743/_0_  ;
	output \g72745/_0_  ;
	output \g72745/_1_  ;
	output \g72752/_0_  ;
	output \g72752/_1_  ;
	output \g72756/_0_  ;
	output \g72763/_0_  ;
	output \g72763/_1_  ;
	output \g72765/_0_  ;
	output \g72767/_0_  ;
	output \g72767/_1_  ;
	output \g72769/_0_  ;
	output \g72769/_1_  ;
	output \g72772/_0_  ;
	output \g72772/_1_  ;
	output \g72774/_0_  ;
	output \g72774/_1_  ;
	output \g72790/_0_  ;
	output \g72790/_1_  ;
	output \g72797/_0_  ;
	output \g73807/_0_  ;
	output \g73820/_0_  ;
	output \g73832/_0_  ;
	output \g73844/_0_  ;
	output \g73856/_0_  ;
	output \g73871/_0_  ;
	output \g73883/_0_  ;
	output \g73895/_0_  ;
	output \g73905/_3_  ;
	output \g73910/_0_  ;
	output \g73922/_0_  ;
	output \g73934/_0_  ;
	output \g73946/_0_  ;
	output \g73958/_0_  ;
	output \g73970/_0_  ;
	output \g73982/_0_  ;
	output \g87036/_0_  ;
	output \g87042/_0_  ;
	output \g87043/_0_  ;
	output \g87044/_0_  ;
	output \g87045/_0_  ;
	output \g87046/_0_  ;
	output \g87047/_0_  ;
	output \g87048/_0_  ;
	output \g87049/_0_  ;
	output \g87050/_0_  ;
	output \g87051/_0_  ;
	output \g87052/_0_  ;
	output \g87053/_0_  ;
	output \g87054/_0_  ;
	output \g87055/_0_  ;
	output \g87062/_0_  ;
	output \g88572/_0_  ;
	output \g88681/_0_  ;
	output \g88682/_0_  ;
	output \g88683/_0_  ;
	output \g88684/_0_  ;
	output \g88685/_0_  ;
	output \g88686/_0_  ;
	output \g88687/_0_  ;
	output \g88688/_0_  ;
	output \g88689/_0_  ;
	output \g88690/_0_  ;
	output \g88691/_0_  ;
	output \g88692/_0_  ;
	output \g88693/_0_  ;
	output \g88695/_0_  ;
	output \g88697/_0_  ;
	output \g88698/_0_  ;
	output \g88700/_0_  ;
	output \g88701/_0_  ;
	output \g88703/_0_  ;
	output \g88704/_0_  ;
	output \g88705/_0_  ;
	output \g88706/_0_  ;
	output \g88707/_0_  ;
	output \g88709/_0_  ;
	output \g88710/_0_  ;
	output \g88711/_0_  ;
	output \g88712/_0_  ;
	output \g88713/_0_  ;
	output \g88714/_0_  ;
	output \g88716/_0_  ;
	output \g88717/_0_  ;
	output \g88718/_0_  ;
	output \g88719/_0_  ;
	output \g88720/_0_  ;
	output \g88722/_0_  ;
	output \g88723/_0_  ;
	output \g88724/_0_  ;
	output \g88725/_0_  ;
	output \g88726/_0_  ;
	output \g88727/_0_  ;
	output \g88728/_0_  ;
	output \g88729/_0_  ;
	output \g88731/_0_  ;
	output \g88732/_0_  ;
	output \g88733/_0_  ;
	output \g88734/_0_  ;
	output \g88736/_0_  ;
	output \g88737/_0_  ;
	output \g88738/_0_  ;
	output \g88739/_0_  ;
	output \g88740/_0_  ;
	output \g88741/_0_  ;
	output \g88742/_0_  ;
	output \g88743/_0_  ;
	output \g88744/_0_  ;
	output \g88745/_0_  ;
	output \g88746/_0_  ;
	output \g88748/_0_  ;
	output \g88749/_0_  ;
	output \g88750/_0_  ;
	output \g88752/_0_  ;
	output \g88753/_0_  ;
	output \g88754/_0_  ;
	output \g88755/_0_  ;
	output \g88756/_0_  ;
	output \g88757/_0_  ;
	output \g88759/_0_  ;
	output \g88760/_0_  ;
	output \g88761/_0_  ;
	output \g88762/_0_  ;
	output \g88764/_0_  ;
	output \g88765/_0_  ;
	output \g88766/_0_  ;
	output \g88768/_0_  ;
	output \g88769/_0_  ;
	output \g88770/_0_  ;
	output \g88771/_0_  ;
	output \g88772/_0_  ;
	output \g88773/_0_  ;
	output \g88775/_0_  ;
	output \g88776/_0_  ;
	output \g88777/_0_  ;
	output \g88778/_0_  ;
	output \g88779/_0_  ;
	output \g88780/_0_  ;
	output \g88782/_0_  ;
	output \g88783/_0_  ;
	output \g88784/_0_  ;
	output \g88785/_0_  ;
	output \g88786/_0_  ;
	output \g88787/_0_  ;
	output \g88789/_0_  ;
	output \g88790/_0_  ;
	output \g88791/_0_  ;
	output \g88792/_0_  ;
	output \g88793/_0_  ;
	output \g88795/_0_  ;
	output \g88796/_0_  ;
	output \g88797/_0_  ;
	output \g88799/_0_  ;
	output \g88800/_0_  ;
	output \g88801/_0_  ;
	output \g88802/_0_  ;
	output \g88806/_0_  ;
	output \g88807/_0_  ;
	output \g88808/_0_  ;
	output \g88809/_0_  ;
	output \g88810/_0_  ;
	output \g88813/_0_  ;
	output \g88814/_0_  ;
	output \g88815/_0_  ;
	output \m0_ack_o_pad  ;
	output \m0_data_o[0]_pad  ;
	output \m0_data_o[10]_pad  ;
	output \m0_data_o[11]_pad  ;
	output \m0_data_o[12]_pad  ;
	output \m0_data_o[13]_pad  ;
	output \m0_data_o[14]_pad  ;
	output \m0_data_o[15]_pad  ;
	output \m0_data_o[16]_pad  ;
	output \m0_data_o[17]_pad  ;
	output \m0_data_o[18]_pad  ;
	output \m0_data_o[19]_pad  ;
	output \m0_data_o[1]_pad  ;
	output \m0_data_o[20]_pad  ;
	output \m0_data_o[21]_pad  ;
	output \m0_data_o[22]_pad  ;
	output \m0_data_o[23]_pad  ;
	output \m0_data_o[24]_pad  ;
	output \m0_data_o[25]_pad  ;
	output \m0_data_o[26]_pad  ;
	output \m0_data_o[27]_pad  ;
	output \m0_data_o[28]_pad  ;
	output \m0_data_o[29]_pad  ;
	output \m0_data_o[2]_pad  ;
	output \m0_data_o[30]_pad  ;
	output \m0_data_o[31]_pad  ;
	output \m0_data_o[3]_pad  ;
	output \m0_data_o[4]_pad  ;
	output \m0_data_o[5]_pad  ;
	output \m0_data_o[6]_pad  ;
	output \m0_data_o[7]_pad  ;
	output \m0_data_o[8]_pad  ;
	output \m0_data_o[9]_pad  ;
	output \m0_err_o_pad  ;
	output \m0_rty_o_pad  ;
	output \m1_ack_o_pad  ;
	output \m1_data_o[0]_pad  ;
	output \m1_data_o[10]_pad  ;
	output \m1_data_o[11]_pad  ;
	output \m1_data_o[12]_pad  ;
	output \m1_data_o[13]_pad  ;
	output \m1_data_o[14]_pad  ;
	output \m1_data_o[15]_pad  ;
	output \m1_data_o[16]_pad  ;
	output \m1_data_o[17]_pad  ;
	output \m1_data_o[18]_pad  ;
	output \m1_data_o[19]_pad  ;
	output \m1_data_o[1]_pad  ;
	output \m1_data_o[20]_pad  ;
	output \m1_data_o[21]_pad  ;
	output \m1_data_o[22]_pad  ;
	output \m1_data_o[23]_pad  ;
	output \m1_data_o[24]_pad  ;
	output \m1_data_o[25]_pad  ;
	output \m1_data_o[26]_pad  ;
	output \m1_data_o[27]_pad  ;
	output \m1_data_o[28]_pad  ;
	output \m1_data_o[29]_pad  ;
	output \m1_data_o[2]_pad  ;
	output \m1_data_o[30]_pad  ;
	output \m1_data_o[31]_pad  ;
	output \m1_data_o[3]_pad  ;
	output \m1_data_o[4]_pad  ;
	output \m1_data_o[5]_pad  ;
	output \m1_data_o[6]_pad  ;
	output \m1_data_o[7]_pad  ;
	output \m1_data_o[8]_pad  ;
	output \m1_data_o[9]_pad  ;
	output \m1_err_o_pad  ;
	output \m1_rty_o_pad  ;
	output \m2_ack_o_pad  ;
	output \m2_data_o[0]_pad  ;
	output \m2_data_o[10]_pad  ;
	output \m2_data_o[11]_pad  ;
	output \m2_data_o[12]_pad  ;
	output \m2_data_o[13]_pad  ;
	output \m2_data_o[14]_pad  ;
	output \m2_data_o[15]_pad  ;
	output \m2_data_o[16]_pad  ;
	output \m2_data_o[17]_pad  ;
	output \m2_data_o[18]_pad  ;
	output \m2_data_o[19]_pad  ;
	output \m2_data_o[1]_pad  ;
	output \m2_data_o[20]_pad  ;
	output \m2_data_o[21]_pad  ;
	output \m2_data_o[22]_pad  ;
	output \m2_data_o[23]_pad  ;
	output \m2_data_o[24]_pad  ;
	output \m2_data_o[25]_pad  ;
	output \m2_data_o[26]_pad  ;
	output \m2_data_o[27]_pad  ;
	output \m2_data_o[28]_pad  ;
	output \m2_data_o[29]_pad  ;
	output \m2_data_o[2]_pad  ;
	output \m2_data_o[30]_pad  ;
	output \m2_data_o[31]_pad  ;
	output \m2_data_o[3]_pad  ;
	output \m2_data_o[4]_pad  ;
	output \m2_data_o[5]_pad  ;
	output \m2_data_o[6]_pad  ;
	output \m2_data_o[7]_pad  ;
	output \m2_data_o[8]_pad  ;
	output \m2_data_o[9]_pad  ;
	output \m2_err_o_pad  ;
	output \m2_rty_o_pad  ;
	output \m3_ack_o_pad  ;
	output \m3_data_o[0]_pad  ;
	output \m3_data_o[10]_pad  ;
	output \m3_data_o[11]_pad  ;
	output \m3_data_o[12]_pad  ;
	output \m3_data_o[13]_pad  ;
	output \m3_data_o[14]_pad  ;
	output \m3_data_o[15]_pad  ;
	output \m3_data_o[16]_pad  ;
	output \m3_data_o[17]_pad  ;
	output \m3_data_o[18]_pad  ;
	output \m3_data_o[19]_pad  ;
	output \m3_data_o[1]_pad  ;
	output \m3_data_o[20]_pad  ;
	output \m3_data_o[21]_pad  ;
	output \m3_data_o[22]_pad  ;
	output \m3_data_o[23]_pad  ;
	output \m3_data_o[24]_pad  ;
	output \m3_data_o[25]_pad  ;
	output \m3_data_o[26]_pad  ;
	output \m3_data_o[27]_pad  ;
	output \m3_data_o[28]_pad  ;
	output \m3_data_o[29]_pad  ;
	output \m3_data_o[2]_pad  ;
	output \m3_data_o[30]_pad  ;
	output \m3_data_o[31]_pad  ;
	output \m3_data_o[3]_pad  ;
	output \m3_data_o[4]_pad  ;
	output \m3_data_o[5]_pad  ;
	output \m3_data_o[6]_pad  ;
	output \m3_data_o[7]_pad  ;
	output \m3_data_o[8]_pad  ;
	output \m3_data_o[9]_pad  ;
	output \m3_err_o_pad  ;
	output \m3_rty_o_pad  ;
	output \m4_ack_o_pad  ;
	output \m4_data_o[0]_pad  ;
	output \m4_data_o[10]_pad  ;
	output \m4_data_o[11]_pad  ;
	output \m4_data_o[12]_pad  ;
	output \m4_data_o[13]_pad  ;
	output \m4_data_o[14]_pad  ;
	output \m4_data_o[15]_pad  ;
	output \m4_data_o[16]_pad  ;
	output \m4_data_o[17]_pad  ;
	output \m4_data_o[18]_pad  ;
	output \m4_data_o[19]_pad  ;
	output \m4_data_o[1]_pad  ;
	output \m4_data_o[20]_pad  ;
	output \m4_data_o[21]_pad  ;
	output \m4_data_o[22]_pad  ;
	output \m4_data_o[23]_pad  ;
	output \m4_data_o[24]_pad  ;
	output \m4_data_o[25]_pad  ;
	output \m4_data_o[26]_pad  ;
	output \m4_data_o[27]_pad  ;
	output \m4_data_o[28]_pad  ;
	output \m4_data_o[29]_pad  ;
	output \m4_data_o[2]_pad  ;
	output \m4_data_o[30]_pad  ;
	output \m4_data_o[31]_pad  ;
	output \m4_data_o[3]_pad  ;
	output \m4_data_o[4]_pad  ;
	output \m4_data_o[5]_pad  ;
	output \m4_data_o[6]_pad  ;
	output \m4_data_o[7]_pad  ;
	output \m4_data_o[8]_pad  ;
	output \m4_data_o[9]_pad  ;
	output \m4_err_o_pad  ;
	output \m4_rty_o_pad  ;
	output \m5_ack_o_pad  ;
	output \m5_data_o[0]_pad  ;
	output \m5_data_o[10]_pad  ;
	output \m5_data_o[11]_pad  ;
	output \m5_data_o[12]_pad  ;
	output \m5_data_o[13]_pad  ;
	output \m5_data_o[14]_pad  ;
	output \m5_data_o[15]_pad  ;
	output \m5_data_o[16]_pad  ;
	output \m5_data_o[17]_pad  ;
	output \m5_data_o[18]_pad  ;
	output \m5_data_o[19]_pad  ;
	output \m5_data_o[1]_pad  ;
	output \m5_data_o[20]_pad  ;
	output \m5_data_o[21]_pad  ;
	output \m5_data_o[22]_pad  ;
	output \m5_data_o[23]_pad  ;
	output \m5_data_o[24]_pad  ;
	output \m5_data_o[25]_pad  ;
	output \m5_data_o[26]_pad  ;
	output \m5_data_o[27]_pad  ;
	output \m5_data_o[28]_pad  ;
	output \m5_data_o[29]_pad  ;
	output \m5_data_o[2]_pad  ;
	output \m5_data_o[30]_pad  ;
	output \m5_data_o[31]_pad  ;
	output \m5_data_o[3]_pad  ;
	output \m5_data_o[4]_pad  ;
	output \m5_data_o[5]_pad  ;
	output \m5_data_o[6]_pad  ;
	output \m5_data_o[7]_pad  ;
	output \m5_data_o[8]_pad  ;
	output \m5_data_o[9]_pad  ;
	output \m5_err_o_pad  ;
	output \m5_rty_o_pad  ;
	output \m6_ack_o_pad  ;
	output \m6_data_o[0]_pad  ;
	output \m6_data_o[10]_pad  ;
	output \m6_data_o[11]_pad  ;
	output \m6_data_o[12]_pad  ;
	output \m6_data_o[13]_pad  ;
	output \m6_data_o[14]_pad  ;
	output \m6_data_o[15]_pad  ;
	output \m6_data_o[16]_pad  ;
	output \m6_data_o[17]_pad  ;
	output \m6_data_o[18]_pad  ;
	output \m6_data_o[19]_pad  ;
	output \m6_data_o[1]_pad  ;
	output \m6_data_o[20]_pad  ;
	output \m6_data_o[21]_pad  ;
	output \m6_data_o[22]_pad  ;
	output \m6_data_o[23]_pad  ;
	output \m6_data_o[24]_pad  ;
	output \m6_data_o[25]_pad  ;
	output \m6_data_o[26]_pad  ;
	output \m6_data_o[27]_pad  ;
	output \m6_data_o[28]_pad  ;
	output \m6_data_o[29]_pad  ;
	output \m6_data_o[2]_pad  ;
	output \m6_data_o[30]_pad  ;
	output \m6_data_o[31]_pad  ;
	output \m6_data_o[3]_pad  ;
	output \m6_data_o[4]_pad  ;
	output \m6_data_o[5]_pad  ;
	output \m6_data_o[6]_pad  ;
	output \m6_data_o[7]_pad  ;
	output \m6_data_o[8]_pad  ;
	output \m6_data_o[9]_pad  ;
	output \m6_err_o_pad  ;
	output \m6_rty_o_pad  ;
	output \m7_ack_o_pad  ;
	output \m7_data_o[0]_pad  ;
	output \m7_data_o[10]_pad  ;
	output \m7_data_o[11]_pad  ;
	output \m7_data_o[12]_pad  ;
	output \m7_data_o[13]_pad  ;
	output \m7_data_o[14]_pad  ;
	output \m7_data_o[15]_pad  ;
	output \m7_data_o[16]_pad  ;
	output \m7_data_o[17]_pad  ;
	output \m7_data_o[18]_pad  ;
	output \m7_data_o[19]_pad  ;
	output \m7_data_o[1]_pad  ;
	output \m7_data_o[20]_pad  ;
	output \m7_data_o[21]_pad  ;
	output \m7_data_o[22]_pad  ;
	output \m7_data_o[23]_pad  ;
	output \m7_data_o[24]_pad  ;
	output \m7_data_o[25]_pad  ;
	output \m7_data_o[26]_pad  ;
	output \m7_data_o[27]_pad  ;
	output \m7_data_o[28]_pad  ;
	output \m7_data_o[29]_pad  ;
	output \m7_data_o[2]_pad  ;
	output \m7_data_o[30]_pad  ;
	output \m7_data_o[31]_pad  ;
	output \m7_data_o[3]_pad  ;
	output \m7_data_o[4]_pad  ;
	output \m7_data_o[5]_pad  ;
	output \m7_data_o[6]_pad  ;
	output \m7_data_o[7]_pad  ;
	output \m7_data_o[8]_pad  ;
	output \m7_data_o[9]_pad  ;
	output \m7_err_o_pad  ;
	output \m7_rty_o_pad  ;
	output \s0_addr_o[0]_pad  ;
	output \s0_addr_o[10]_pad  ;
	output \s0_addr_o[11]_pad  ;
	output \s0_addr_o[12]_pad  ;
	output \s0_addr_o[13]_pad  ;
	output \s0_addr_o[14]_pad  ;
	output \s0_addr_o[15]_pad  ;
	output \s0_addr_o[16]_pad  ;
	output \s0_addr_o[17]_pad  ;
	output \s0_addr_o[18]_pad  ;
	output \s0_addr_o[19]_pad  ;
	output \s0_addr_o[1]_pad  ;
	output \s0_addr_o[20]_pad  ;
	output \s0_addr_o[21]_pad  ;
	output \s0_addr_o[22]_pad  ;
	output \s0_addr_o[23]_pad  ;
	output \s0_addr_o[24]_pad  ;
	output \s0_addr_o[25]_pad  ;
	output \s0_addr_o[26]_pad  ;
	output \s0_addr_o[27]_pad  ;
	output \s0_addr_o[28]_pad  ;
	output \s0_addr_o[29]_pad  ;
	output \s0_addr_o[2]_pad  ;
	output \s0_addr_o[30]_pad  ;
	output \s0_addr_o[31]_pad  ;
	output \s0_addr_o[3]_pad  ;
	output \s0_addr_o[4]_pad  ;
	output \s0_addr_o[5]_pad  ;
	output \s0_addr_o[6]_pad  ;
	output \s0_addr_o[7]_pad  ;
	output \s0_addr_o[8]_pad  ;
	output \s0_addr_o[9]_pad  ;
	output \s0_data_o[0]_pad  ;
	output \s0_data_o[10]_pad  ;
	output \s0_data_o[11]_pad  ;
	output \s0_data_o[12]_pad  ;
	output \s0_data_o[13]_pad  ;
	output \s0_data_o[14]_pad  ;
	output \s0_data_o[15]_pad  ;
	output \s0_data_o[16]_pad  ;
	output \s0_data_o[17]_pad  ;
	output \s0_data_o[18]_pad  ;
	output \s0_data_o[19]_pad  ;
	output \s0_data_o[1]_pad  ;
	output \s0_data_o[20]_pad  ;
	output \s0_data_o[21]_pad  ;
	output \s0_data_o[22]_pad  ;
	output \s0_data_o[23]_pad  ;
	output \s0_data_o[24]_pad  ;
	output \s0_data_o[25]_pad  ;
	output \s0_data_o[26]_pad  ;
	output \s0_data_o[27]_pad  ;
	output \s0_data_o[28]_pad  ;
	output \s0_data_o[29]_pad  ;
	output \s0_data_o[2]_pad  ;
	output \s0_data_o[30]_pad  ;
	output \s0_data_o[31]_pad  ;
	output \s0_data_o[3]_pad  ;
	output \s0_data_o[4]_pad  ;
	output \s0_data_o[5]_pad  ;
	output \s0_data_o[6]_pad  ;
	output \s0_data_o[7]_pad  ;
	output \s0_data_o[8]_pad  ;
	output \s0_data_o[9]_pad  ;
	output \s0_sel_o[0]_pad  ;
	output \s0_sel_o[1]_pad  ;
	output \s0_sel_o[2]_pad  ;
	output \s0_sel_o[3]_pad  ;
	output \s0_stb_o_pad  ;
	output \s0_we_o_pad  ;
	output \s10_addr_o[0]_pad  ;
	output \s10_addr_o[10]_pad  ;
	output \s10_addr_o[11]_pad  ;
	output \s10_addr_o[12]_pad  ;
	output \s10_addr_o[13]_pad  ;
	output \s10_addr_o[14]_pad  ;
	output \s10_addr_o[15]_pad  ;
	output \s10_addr_o[16]_pad  ;
	output \s10_addr_o[17]_pad  ;
	output \s10_addr_o[18]_pad  ;
	output \s10_addr_o[19]_pad  ;
	output \s10_addr_o[1]_pad  ;
	output \s10_addr_o[20]_pad  ;
	output \s10_addr_o[21]_pad  ;
	output \s10_addr_o[22]_pad  ;
	output \s10_addr_o[23]_pad  ;
	output \s10_addr_o[24]_pad  ;
	output \s10_addr_o[25]_pad  ;
	output \s10_addr_o[26]_pad  ;
	output \s10_addr_o[27]_pad  ;
	output \s10_addr_o[28]_pad  ;
	output \s10_addr_o[29]_pad  ;
	output \s10_addr_o[2]_pad  ;
	output \s10_addr_o[30]_pad  ;
	output \s10_addr_o[31]_pad  ;
	output \s10_addr_o[3]_pad  ;
	output \s10_addr_o[4]_pad  ;
	output \s10_addr_o[5]_pad  ;
	output \s10_addr_o[6]_pad  ;
	output \s10_addr_o[7]_pad  ;
	output \s10_addr_o[8]_pad  ;
	output \s10_addr_o[9]_pad  ;
	output \s10_data_o[0]_pad  ;
	output \s10_data_o[10]_pad  ;
	output \s10_data_o[11]_pad  ;
	output \s10_data_o[12]_pad  ;
	output \s10_data_o[13]_pad  ;
	output \s10_data_o[14]_pad  ;
	output \s10_data_o[15]_pad  ;
	output \s10_data_o[16]_pad  ;
	output \s10_data_o[17]_pad  ;
	output \s10_data_o[18]_pad  ;
	output \s10_data_o[19]_pad  ;
	output \s10_data_o[1]_pad  ;
	output \s10_data_o[20]_pad  ;
	output \s10_data_o[21]_pad  ;
	output \s10_data_o[22]_pad  ;
	output \s10_data_o[23]_pad  ;
	output \s10_data_o[24]_pad  ;
	output \s10_data_o[25]_pad  ;
	output \s10_data_o[26]_pad  ;
	output \s10_data_o[27]_pad  ;
	output \s10_data_o[28]_pad  ;
	output \s10_data_o[29]_pad  ;
	output \s10_data_o[2]_pad  ;
	output \s10_data_o[30]_pad  ;
	output \s10_data_o[31]_pad  ;
	output \s10_data_o[3]_pad  ;
	output \s10_data_o[4]_pad  ;
	output \s10_data_o[5]_pad  ;
	output \s10_data_o[6]_pad  ;
	output \s10_data_o[7]_pad  ;
	output \s10_data_o[8]_pad  ;
	output \s10_data_o[9]_pad  ;
	output \s10_sel_o[0]_pad  ;
	output \s10_sel_o[1]_pad  ;
	output \s10_sel_o[2]_pad  ;
	output \s10_sel_o[3]_pad  ;
	output \s10_stb_o_pad  ;
	output \s10_we_o_pad  ;
	output \s11_addr_o[0]_pad  ;
	output \s11_addr_o[10]_pad  ;
	output \s11_addr_o[11]_pad  ;
	output \s11_addr_o[12]_pad  ;
	output \s11_addr_o[13]_pad  ;
	output \s11_addr_o[14]_pad  ;
	output \s11_addr_o[15]_pad  ;
	output \s11_addr_o[16]_pad  ;
	output \s11_addr_o[17]_pad  ;
	output \s11_addr_o[18]_pad  ;
	output \s11_addr_o[19]_pad  ;
	output \s11_addr_o[1]_pad  ;
	output \s11_addr_o[20]_pad  ;
	output \s11_addr_o[21]_pad  ;
	output \s11_addr_o[22]_pad  ;
	output \s11_addr_o[23]_pad  ;
	output \s11_addr_o[24]_pad  ;
	output \s11_addr_o[25]_pad  ;
	output \s11_addr_o[26]_pad  ;
	output \s11_addr_o[27]_pad  ;
	output \s11_addr_o[28]_pad  ;
	output \s11_addr_o[29]_pad  ;
	output \s11_addr_o[2]_pad  ;
	output \s11_addr_o[30]_pad  ;
	output \s11_addr_o[31]_pad  ;
	output \s11_addr_o[3]_pad  ;
	output \s11_addr_o[4]_pad  ;
	output \s11_addr_o[5]_pad  ;
	output \s11_addr_o[6]_pad  ;
	output \s11_addr_o[7]_pad  ;
	output \s11_addr_o[8]_pad  ;
	output \s11_addr_o[9]_pad  ;
	output \s11_data_o[0]_pad  ;
	output \s11_data_o[10]_pad  ;
	output \s11_data_o[11]_pad  ;
	output \s11_data_o[12]_pad  ;
	output \s11_data_o[13]_pad  ;
	output \s11_data_o[14]_pad  ;
	output \s11_data_o[15]_pad  ;
	output \s11_data_o[16]_pad  ;
	output \s11_data_o[17]_pad  ;
	output \s11_data_o[18]_pad  ;
	output \s11_data_o[19]_pad  ;
	output \s11_data_o[1]_pad  ;
	output \s11_data_o[20]_pad  ;
	output \s11_data_o[21]_pad  ;
	output \s11_data_o[22]_pad  ;
	output \s11_data_o[23]_pad  ;
	output \s11_data_o[24]_pad  ;
	output \s11_data_o[25]_pad  ;
	output \s11_data_o[26]_pad  ;
	output \s11_data_o[27]_pad  ;
	output \s11_data_o[28]_pad  ;
	output \s11_data_o[29]_pad  ;
	output \s11_data_o[2]_pad  ;
	output \s11_data_o[30]_pad  ;
	output \s11_data_o[31]_pad  ;
	output \s11_data_o[3]_pad  ;
	output \s11_data_o[4]_pad  ;
	output \s11_data_o[5]_pad  ;
	output \s11_data_o[6]_pad  ;
	output \s11_data_o[7]_pad  ;
	output \s11_data_o[8]_pad  ;
	output \s11_data_o[9]_pad  ;
	output \s11_sel_o[0]_pad  ;
	output \s11_sel_o[1]_pad  ;
	output \s11_sel_o[2]_pad  ;
	output \s11_sel_o[3]_pad  ;
	output \s11_stb_o_pad  ;
	output \s11_we_o_pad  ;
	output \s12_addr_o[0]_pad  ;
	output \s12_addr_o[10]_pad  ;
	output \s12_addr_o[11]_pad  ;
	output \s12_addr_o[12]_pad  ;
	output \s12_addr_o[13]_pad  ;
	output \s12_addr_o[14]_pad  ;
	output \s12_addr_o[15]_pad  ;
	output \s12_addr_o[16]_pad  ;
	output \s12_addr_o[17]_pad  ;
	output \s12_addr_o[18]_pad  ;
	output \s12_addr_o[19]_pad  ;
	output \s12_addr_o[1]_pad  ;
	output \s12_addr_o[20]_pad  ;
	output \s12_addr_o[21]_pad  ;
	output \s12_addr_o[22]_pad  ;
	output \s12_addr_o[23]_pad  ;
	output \s12_addr_o[24]_pad  ;
	output \s12_addr_o[25]_pad  ;
	output \s12_addr_o[26]_pad  ;
	output \s12_addr_o[27]_pad  ;
	output \s12_addr_o[28]_pad  ;
	output \s12_addr_o[29]_pad  ;
	output \s12_addr_o[2]_pad  ;
	output \s12_addr_o[30]_pad  ;
	output \s12_addr_o[31]_pad  ;
	output \s12_addr_o[3]_pad  ;
	output \s12_addr_o[4]_pad  ;
	output \s12_addr_o[5]_pad  ;
	output \s12_addr_o[6]_pad  ;
	output \s12_addr_o[7]_pad  ;
	output \s12_addr_o[8]_pad  ;
	output \s12_addr_o[9]_pad  ;
	output \s12_data_o[0]_pad  ;
	output \s12_data_o[10]_pad  ;
	output \s12_data_o[11]_pad  ;
	output \s12_data_o[12]_pad  ;
	output \s12_data_o[13]_pad  ;
	output \s12_data_o[14]_pad  ;
	output \s12_data_o[15]_pad  ;
	output \s12_data_o[16]_pad  ;
	output \s12_data_o[17]_pad  ;
	output \s12_data_o[18]_pad  ;
	output \s12_data_o[19]_pad  ;
	output \s12_data_o[1]_pad  ;
	output \s12_data_o[20]_pad  ;
	output \s12_data_o[21]_pad  ;
	output \s12_data_o[22]_pad  ;
	output \s12_data_o[23]_pad  ;
	output \s12_data_o[24]_pad  ;
	output \s12_data_o[25]_pad  ;
	output \s12_data_o[26]_pad  ;
	output \s12_data_o[27]_pad  ;
	output \s12_data_o[28]_pad  ;
	output \s12_data_o[29]_pad  ;
	output \s12_data_o[2]_pad  ;
	output \s12_data_o[30]_pad  ;
	output \s12_data_o[31]_pad  ;
	output \s12_data_o[3]_pad  ;
	output \s12_data_o[4]_pad  ;
	output \s12_data_o[5]_pad  ;
	output \s12_data_o[6]_pad  ;
	output \s12_data_o[7]_pad  ;
	output \s12_data_o[8]_pad  ;
	output \s12_data_o[9]_pad  ;
	output \s12_sel_o[0]_pad  ;
	output \s12_sel_o[1]_pad  ;
	output \s12_sel_o[2]_pad  ;
	output \s12_sel_o[3]_pad  ;
	output \s12_stb_o_pad  ;
	output \s12_we_o_pad  ;
	output \s13_addr_o[0]_pad  ;
	output \s13_addr_o[10]_pad  ;
	output \s13_addr_o[11]_pad  ;
	output \s13_addr_o[12]_pad  ;
	output \s13_addr_o[13]_pad  ;
	output \s13_addr_o[14]_pad  ;
	output \s13_addr_o[15]_pad  ;
	output \s13_addr_o[16]_pad  ;
	output \s13_addr_o[17]_pad  ;
	output \s13_addr_o[18]_pad  ;
	output \s13_addr_o[19]_pad  ;
	output \s13_addr_o[1]_pad  ;
	output \s13_addr_o[20]_pad  ;
	output \s13_addr_o[21]_pad  ;
	output \s13_addr_o[22]_pad  ;
	output \s13_addr_o[23]_pad  ;
	output \s13_addr_o[24]_pad  ;
	output \s13_addr_o[25]_pad  ;
	output \s13_addr_o[26]_pad  ;
	output \s13_addr_o[27]_pad  ;
	output \s13_addr_o[28]_pad  ;
	output \s13_addr_o[29]_pad  ;
	output \s13_addr_o[2]_pad  ;
	output \s13_addr_o[30]_pad  ;
	output \s13_addr_o[31]_pad  ;
	output \s13_addr_o[3]_pad  ;
	output \s13_addr_o[4]_pad  ;
	output \s13_addr_o[5]_pad  ;
	output \s13_addr_o[6]_pad  ;
	output \s13_addr_o[7]_pad  ;
	output \s13_addr_o[8]_pad  ;
	output \s13_addr_o[9]_pad  ;
	output \s13_data_o[0]_pad  ;
	output \s13_data_o[10]_pad  ;
	output \s13_data_o[11]_pad  ;
	output \s13_data_o[12]_pad  ;
	output \s13_data_o[13]_pad  ;
	output \s13_data_o[14]_pad  ;
	output \s13_data_o[15]_pad  ;
	output \s13_data_o[16]_pad  ;
	output \s13_data_o[17]_pad  ;
	output \s13_data_o[18]_pad  ;
	output \s13_data_o[19]_pad  ;
	output \s13_data_o[1]_pad  ;
	output \s13_data_o[20]_pad  ;
	output \s13_data_o[21]_pad  ;
	output \s13_data_o[22]_pad  ;
	output \s13_data_o[23]_pad  ;
	output \s13_data_o[24]_pad  ;
	output \s13_data_o[25]_pad  ;
	output \s13_data_o[26]_pad  ;
	output \s13_data_o[27]_pad  ;
	output \s13_data_o[28]_pad  ;
	output \s13_data_o[29]_pad  ;
	output \s13_data_o[2]_pad  ;
	output \s13_data_o[30]_pad  ;
	output \s13_data_o[31]_pad  ;
	output \s13_data_o[3]_pad  ;
	output \s13_data_o[4]_pad  ;
	output \s13_data_o[5]_pad  ;
	output \s13_data_o[6]_pad  ;
	output \s13_data_o[7]_pad  ;
	output \s13_data_o[8]_pad  ;
	output \s13_data_o[9]_pad  ;
	output \s13_sel_o[0]_pad  ;
	output \s13_sel_o[1]_pad  ;
	output \s13_sel_o[2]_pad  ;
	output \s13_sel_o[3]_pad  ;
	output \s13_stb_o_pad  ;
	output \s13_we_o_pad  ;
	output \s14_addr_o[0]_pad  ;
	output \s14_addr_o[10]_pad  ;
	output \s14_addr_o[11]_pad  ;
	output \s14_addr_o[12]_pad  ;
	output \s14_addr_o[13]_pad  ;
	output \s14_addr_o[14]_pad  ;
	output \s14_addr_o[15]_pad  ;
	output \s14_addr_o[16]_pad  ;
	output \s14_addr_o[17]_pad  ;
	output \s14_addr_o[18]_pad  ;
	output \s14_addr_o[19]_pad  ;
	output \s14_addr_o[1]_pad  ;
	output \s14_addr_o[20]_pad  ;
	output \s14_addr_o[21]_pad  ;
	output \s14_addr_o[22]_pad  ;
	output \s14_addr_o[23]_pad  ;
	output \s14_addr_o[24]_pad  ;
	output \s14_addr_o[25]_pad  ;
	output \s14_addr_o[26]_pad  ;
	output \s14_addr_o[27]_pad  ;
	output \s14_addr_o[28]_pad  ;
	output \s14_addr_o[29]_pad  ;
	output \s14_addr_o[2]_pad  ;
	output \s14_addr_o[30]_pad  ;
	output \s14_addr_o[31]_pad  ;
	output \s14_addr_o[3]_pad  ;
	output \s14_addr_o[4]_pad  ;
	output \s14_addr_o[5]_pad  ;
	output \s14_addr_o[6]_pad  ;
	output \s14_addr_o[7]_pad  ;
	output \s14_addr_o[8]_pad  ;
	output \s14_addr_o[9]_pad  ;
	output \s14_data_o[0]_pad  ;
	output \s14_data_o[10]_pad  ;
	output \s14_data_o[11]_pad  ;
	output \s14_data_o[12]_pad  ;
	output \s14_data_o[13]_pad  ;
	output \s14_data_o[14]_pad  ;
	output \s14_data_o[15]_pad  ;
	output \s14_data_o[16]_pad  ;
	output \s14_data_o[17]_pad  ;
	output \s14_data_o[18]_pad  ;
	output \s14_data_o[19]_pad  ;
	output \s14_data_o[1]_pad  ;
	output \s14_data_o[20]_pad  ;
	output \s14_data_o[21]_pad  ;
	output \s14_data_o[22]_pad  ;
	output \s14_data_o[23]_pad  ;
	output \s14_data_o[24]_pad  ;
	output \s14_data_o[25]_pad  ;
	output \s14_data_o[26]_pad  ;
	output \s14_data_o[27]_pad  ;
	output \s14_data_o[28]_pad  ;
	output \s14_data_o[29]_pad  ;
	output \s14_data_o[2]_pad  ;
	output \s14_data_o[30]_pad  ;
	output \s14_data_o[31]_pad  ;
	output \s14_data_o[3]_pad  ;
	output \s14_data_o[4]_pad  ;
	output \s14_data_o[5]_pad  ;
	output \s14_data_o[6]_pad  ;
	output \s14_data_o[7]_pad  ;
	output \s14_data_o[8]_pad  ;
	output \s14_data_o[9]_pad  ;
	output \s14_sel_o[0]_pad  ;
	output \s14_sel_o[1]_pad  ;
	output \s14_sel_o[2]_pad  ;
	output \s14_sel_o[3]_pad  ;
	output \s14_stb_o_pad  ;
	output \s14_we_o_pad  ;
	output \s15_addr_o[0]_pad  ;
	output \s15_addr_o[10]_pad  ;
	output \s15_addr_o[11]_pad  ;
	output \s15_addr_o[12]_pad  ;
	output \s15_addr_o[13]_pad  ;
	output \s15_addr_o[14]_pad  ;
	output \s15_addr_o[15]_pad  ;
	output \s15_addr_o[16]_pad  ;
	output \s15_addr_o[17]_pad  ;
	output \s15_addr_o[18]_pad  ;
	output \s15_addr_o[19]_pad  ;
	output \s15_addr_o[1]_pad  ;
	output \s15_addr_o[20]_pad  ;
	output \s15_addr_o[21]_pad  ;
	output \s15_addr_o[22]_pad  ;
	output \s15_addr_o[23]_pad  ;
	output \s15_addr_o[24]_pad  ;
	output \s15_addr_o[25]_pad  ;
	output \s15_addr_o[26]_pad  ;
	output \s15_addr_o[27]_pad  ;
	output \s15_addr_o[28]_pad  ;
	output \s15_addr_o[29]_pad  ;
	output \s15_addr_o[2]_pad  ;
	output \s15_addr_o[30]_pad  ;
	output \s15_addr_o[31]_pad  ;
	output \s15_addr_o[3]_pad  ;
	output \s15_addr_o[4]_pad  ;
	output \s15_addr_o[6]_pad  ;
	output \s15_addr_o[7]_pad  ;
	output \s15_addr_o[8]_pad  ;
	output \s15_addr_o[9]_pad  ;
	output \s15_cyc_o_pad  ;
	output \s15_data_o[0]_pad  ;
	output \s15_data_o[10]_pad  ;
	output \s15_data_o[11]_pad  ;
	output \s15_data_o[12]_pad  ;
	output \s15_data_o[13]_pad  ;
	output \s15_data_o[14]_pad  ;
	output \s15_data_o[15]_pad  ;
	output \s15_data_o[16]_pad  ;
	output \s15_data_o[17]_pad  ;
	output \s15_data_o[18]_pad  ;
	output \s15_data_o[19]_pad  ;
	output \s15_data_o[1]_pad  ;
	output \s15_data_o[20]_pad  ;
	output \s15_data_o[21]_pad  ;
	output \s15_data_o[22]_pad  ;
	output \s15_data_o[23]_pad  ;
	output \s15_data_o[24]_pad  ;
	output \s15_data_o[25]_pad  ;
	output \s15_data_o[26]_pad  ;
	output \s15_data_o[27]_pad  ;
	output \s15_data_o[28]_pad  ;
	output \s15_data_o[29]_pad  ;
	output \s15_data_o[2]_pad  ;
	output \s15_data_o[30]_pad  ;
	output \s15_data_o[31]_pad  ;
	output \s15_data_o[3]_pad  ;
	output \s15_data_o[4]_pad  ;
	output \s15_data_o[5]_pad  ;
	output \s15_data_o[6]_pad  ;
	output \s15_data_o[7]_pad  ;
	output \s15_data_o[8]_pad  ;
	output \s15_data_o[9]_pad  ;
	output \s15_sel_o[0]_pad  ;
	output \s15_sel_o[1]_pad  ;
	output \s15_sel_o[2]_pad  ;
	output \s15_sel_o[3]_pad  ;
	output \s15_stb_o_pad  ;
	output \s15_we_o_pad  ;
	output \s1_addr_o[0]_pad  ;
	output \s1_addr_o[10]_pad  ;
	output \s1_addr_o[11]_pad  ;
	output \s1_addr_o[12]_pad  ;
	output \s1_addr_o[13]_pad  ;
	output \s1_addr_o[14]_pad  ;
	output \s1_addr_o[15]_pad  ;
	output \s1_addr_o[16]_pad  ;
	output \s1_addr_o[17]_pad  ;
	output \s1_addr_o[18]_pad  ;
	output \s1_addr_o[19]_pad  ;
	output \s1_addr_o[1]_pad  ;
	output \s1_addr_o[20]_pad  ;
	output \s1_addr_o[21]_pad  ;
	output \s1_addr_o[22]_pad  ;
	output \s1_addr_o[23]_pad  ;
	output \s1_addr_o[24]_pad  ;
	output \s1_addr_o[25]_pad  ;
	output \s1_addr_o[26]_pad  ;
	output \s1_addr_o[27]_pad  ;
	output \s1_addr_o[28]_pad  ;
	output \s1_addr_o[29]_pad  ;
	output \s1_addr_o[2]_pad  ;
	output \s1_addr_o[30]_pad  ;
	output \s1_addr_o[31]_pad  ;
	output \s1_addr_o[3]_pad  ;
	output \s1_addr_o[4]_pad  ;
	output \s1_addr_o[5]_pad  ;
	output \s1_addr_o[6]_pad  ;
	output \s1_addr_o[7]_pad  ;
	output \s1_addr_o[8]_pad  ;
	output \s1_addr_o[9]_pad  ;
	output \s1_data_o[0]_pad  ;
	output \s1_data_o[10]_pad  ;
	output \s1_data_o[11]_pad  ;
	output \s1_data_o[12]_pad  ;
	output \s1_data_o[13]_pad  ;
	output \s1_data_o[14]_pad  ;
	output \s1_data_o[15]_pad  ;
	output \s1_data_o[16]_pad  ;
	output \s1_data_o[17]_pad  ;
	output \s1_data_o[18]_pad  ;
	output \s1_data_o[19]_pad  ;
	output \s1_data_o[1]_pad  ;
	output \s1_data_o[20]_pad  ;
	output \s1_data_o[21]_pad  ;
	output \s1_data_o[22]_pad  ;
	output \s1_data_o[23]_pad  ;
	output \s1_data_o[24]_pad  ;
	output \s1_data_o[25]_pad  ;
	output \s1_data_o[26]_pad  ;
	output \s1_data_o[27]_pad  ;
	output \s1_data_o[28]_pad  ;
	output \s1_data_o[29]_pad  ;
	output \s1_data_o[2]_pad  ;
	output \s1_data_o[30]_pad  ;
	output \s1_data_o[31]_pad  ;
	output \s1_data_o[3]_pad  ;
	output \s1_data_o[4]_pad  ;
	output \s1_data_o[5]_pad  ;
	output \s1_data_o[6]_pad  ;
	output \s1_data_o[7]_pad  ;
	output \s1_data_o[8]_pad  ;
	output \s1_data_o[9]_pad  ;
	output \s1_sel_o[0]_pad  ;
	output \s1_sel_o[1]_pad  ;
	output \s1_sel_o[2]_pad  ;
	output \s1_sel_o[3]_pad  ;
	output \s1_stb_o_pad  ;
	output \s1_we_o_pad  ;
	output \s2_addr_o[0]_pad  ;
	output \s2_addr_o[10]_pad  ;
	output \s2_addr_o[11]_pad  ;
	output \s2_addr_o[12]_pad  ;
	output \s2_addr_o[13]_pad  ;
	output \s2_addr_o[14]_pad  ;
	output \s2_addr_o[15]_pad  ;
	output \s2_addr_o[16]_pad  ;
	output \s2_addr_o[17]_pad  ;
	output \s2_addr_o[18]_pad  ;
	output \s2_addr_o[19]_pad  ;
	output \s2_addr_o[1]_pad  ;
	output \s2_addr_o[20]_pad  ;
	output \s2_addr_o[21]_pad  ;
	output \s2_addr_o[22]_pad  ;
	output \s2_addr_o[23]_pad  ;
	output \s2_addr_o[24]_pad  ;
	output \s2_addr_o[25]_pad  ;
	output \s2_addr_o[26]_pad  ;
	output \s2_addr_o[27]_pad  ;
	output \s2_addr_o[28]_pad  ;
	output \s2_addr_o[29]_pad  ;
	output \s2_addr_o[2]_pad  ;
	output \s2_addr_o[30]_pad  ;
	output \s2_addr_o[31]_pad  ;
	output \s2_addr_o[3]_pad  ;
	output \s2_addr_o[4]_pad  ;
	output \s2_addr_o[5]_pad  ;
	output \s2_addr_o[6]_pad  ;
	output \s2_addr_o[7]_pad  ;
	output \s2_addr_o[8]_pad  ;
	output \s2_addr_o[9]_pad  ;
	output \s2_data_o[0]_pad  ;
	output \s2_data_o[10]_pad  ;
	output \s2_data_o[11]_pad  ;
	output \s2_data_o[12]_pad  ;
	output \s2_data_o[13]_pad  ;
	output \s2_data_o[14]_pad  ;
	output \s2_data_o[15]_pad  ;
	output \s2_data_o[16]_pad  ;
	output \s2_data_o[17]_pad  ;
	output \s2_data_o[18]_pad  ;
	output \s2_data_o[19]_pad  ;
	output \s2_data_o[1]_pad  ;
	output \s2_data_o[20]_pad  ;
	output \s2_data_o[21]_pad  ;
	output \s2_data_o[22]_pad  ;
	output \s2_data_o[23]_pad  ;
	output \s2_data_o[24]_pad  ;
	output \s2_data_o[25]_pad  ;
	output \s2_data_o[26]_pad  ;
	output \s2_data_o[27]_pad  ;
	output \s2_data_o[28]_pad  ;
	output \s2_data_o[29]_pad  ;
	output \s2_data_o[2]_pad  ;
	output \s2_data_o[30]_pad  ;
	output \s2_data_o[31]_pad  ;
	output \s2_data_o[3]_pad  ;
	output \s2_data_o[4]_pad  ;
	output \s2_data_o[5]_pad  ;
	output \s2_data_o[6]_pad  ;
	output \s2_data_o[7]_pad  ;
	output \s2_data_o[8]_pad  ;
	output \s2_data_o[9]_pad  ;
	output \s2_sel_o[0]_pad  ;
	output \s2_sel_o[1]_pad  ;
	output \s2_sel_o[2]_pad  ;
	output \s2_sel_o[3]_pad  ;
	output \s2_stb_o_pad  ;
	output \s2_we_o_pad  ;
	output \s3_addr_o[0]_pad  ;
	output \s3_addr_o[10]_pad  ;
	output \s3_addr_o[11]_pad  ;
	output \s3_addr_o[12]_pad  ;
	output \s3_addr_o[13]_pad  ;
	output \s3_addr_o[14]_pad  ;
	output \s3_addr_o[15]_pad  ;
	output \s3_addr_o[16]_pad  ;
	output \s3_addr_o[17]_pad  ;
	output \s3_addr_o[18]_pad  ;
	output \s3_addr_o[19]_pad  ;
	output \s3_addr_o[1]_pad  ;
	output \s3_addr_o[20]_pad  ;
	output \s3_addr_o[21]_pad  ;
	output \s3_addr_o[22]_pad  ;
	output \s3_addr_o[23]_pad  ;
	output \s3_addr_o[24]_pad  ;
	output \s3_addr_o[25]_pad  ;
	output \s3_addr_o[26]_pad  ;
	output \s3_addr_o[27]_pad  ;
	output \s3_addr_o[28]_pad  ;
	output \s3_addr_o[29]_pad  ;
	output \s3_addr_o[2]_pad  ;
	output \s3_addr_o[30]_pad  ;
	output \s3_addr_o[31]_pad  ;
	output \s3_addr_o[3]_pad  ;
	output \s3_addr_o[4]_pad  ;
	output \s3_addr_o[5]_pad  ;
	output \s3_addr_o[6]_pad  ;
	output \s3_addr_o[7]_pad  ;
	output \s3_addr_o[8]_pad  ;
	output \s3_addr_o[9]_pad  ;
	output \s3_data_o[0]_pad  ;
	output \s3_data_o[10]_pad  ;
	output \s3_data_o[11]_pad  ;
	output \s3_data_o[12]_pad  ;
	output \s3_data_o[13]_pad  ;
	output \s3_data_o[14]_pad  ;
	output \s3_data_o[15]_pad  ;
	output \s3_data_o[16]_pad  ;
	output \s3_data_o[17]_pad  ;
	output \s3_data_o[18]_pad  ;
	output \s3_data_o[19]_pad  ;
	output \s3_data_o[1]_pad  ;
	output \s3_data_o[20]_pad  ;
	output \s3_data_o[21]_pad  ;
	output \s3_data_o[22]_pad  ;
	output \s3_data_o[23]_pad  ;
	output \s3_data_o[24]_pad  ;
	output \s3_data_o[25]_pad  ;
	output \s3_data_o[26]_pad  ;
	output \s3_data_o[27]_pad  ;
	output \s3_data_o[28]_pad  ;
	output \s3_data_o[29]_pad  ;
	output \s3_data_o[2]_pad  ;
	output \s3_data_o[30]_pad  ;
	output \s3_data_o[31]_pad  ;
	output \s3_data_o[3]_pad  ;
	output \s3_data_o[4]_pad  ;
	output \s3_data_o[5]_pad  ;
	output \s3_data_o[6]_pad  ;
	output \s3_data_o[7]_pad  ;
	output \s3_data_o[8]_pad  ;
	output \s3_data_o[9]_pad  ;
	output \s3_sel_o[0]_pad  ;
	output \s3_sel_o[1]_pad  ;
	output \s3_sel_o[2]_pad  ;
	output \s3_sel_o[3]_pad  ;
	output \s3_stb_o_pad  ;
	output \s3_we_o_pad  ;
	output \s4_addr_o[0]_pad  ;
	output \s4_addr_o[10]_pad  ;
	output \s4_addr_o[11]_pad  ;
	output \s4_addr_o[12]_pad  ;
	output \s4_addr_o[13]_pad  ;
	output \s4_addr_o[14]_pad  ;
	output \s4_addr_o[15]_pad  ;
	output \s4_addr_o[16]_pad  ;
	output \s4_addr_o[17]_pad  ;
	output \s4_addr_o[18]_pad  ;
	output \s4_addr_o[19]_pad  ;
	output \s4_addr_o[1]_pad  ;
	output \s4_addr_o[20]_pad  ;
	output \s4_addr_o[21]_pad  ;
	output \s4_addr_o[22]_pad  ;
	output \s4_addr_o[23]_pad  ;
	output \s4_addr_o[24]_pad  ;
	output \s4_addr_o[25]_pad  ;
	output \s4_addr_o[26]_pad  ;
	output \s4_addr_o[27]_pad  ;
	output \s4_addr_o[28]_pad  ;
	output \s4_addr_o[29]_pad  ;
	output \s4_addr_o[2]_pad  ;
	output \s4_addr_o[30]_pad  ;
	output \s4_addr_o[31]_pad  ;
	output \s4_addr_o[3]_pad  ;
	output \s4_addr_o[4]_pad  ;
	output \s4_addr_o[5]_pad  ;
	output \s4_addr_o[6]_pad  ;
	output \s4_addr_o[7]_pad  ;
	output \s4_addr_o[8]_pad  ;
	output \s4_addr_o[9]_pad  ;
	output \s4_data_o[0]_pad  ;
	output \s4_data_o[10]_pad  ;
	output \s4_data_o[11]_pad  ;
	output \s4_data_o[12]_pad  ;
	output \s4_data_o[13]_pad  ;
	output \s4_data_o[14]_pad  ;
	output \s4_data_o[15]_pad  ;
	output \s4_data_o[16]_pad  ;
	output \s4_data_o[17]_pad  ;
	output \s4_data_o[18]_pad  ;
	output \s4_data_o[19]_pad  ;
	output \s4_data_o[1]_pad  ;
	output \s4_data_o[20]_pad  ;
	output \s4_data_o[21]_pad  ;
	output \s4_data_o[22]_pad  ;
	output \s4_data_o[23]_pad  ;
	output \s4_data_o[24]_pad  ;
	output \s4_data_o[25]_pad  ;
	output \s4_data_o[26]_pad  ;
	output \s4_data_o[27]_pad  ;
	output \s4_data_o[28]_pad  ;
	output \s4_data_o[29]_pad  ;
	output \s4_data_o[2]_pad  ;
	output \s4_data_o[30]_pad  ;
	output \s4_data_o[31]_pad  ;
	output \s4_data_o[3]_pad  ;
	output \s4_data_o[4]_pad  ;
	output \s4_data_o[5]_pad  ;
	output \s4_data_o[6]_pad  ;
	output \s4_data_o[7]_pad  ;
	output \s4_data_o[8]_pad  ;
	output \s4_data_o[9]_pad  ;
	output \s4_sel_o[0]_pad  ;
	output \s4_sel_o[1]_pad  ;
	output \s4_sel_o[2]_pad  ;
	output \s4_sel_o[3]_pad  ;
	output \s4_stb_o_pad  ;
	output \s4_we_o_pad  ;
	output \s5_addr_o[0]_pad  ;
	output \s5_addr_o[10]_pad  ;
	output \s5_addr_o[11]_pad  ;
	output \s5_addr_o[12]_pad  ;
	output \s5_addr_o[13]_pad  ;
	output \s5_addr_o[14]_pad  ;
	output \s5_addr_o[15]_pad  ;
	output \s5_addr_o[16]_pad  ;
	output \s5_addr_o[17]_pad  ;
	output \s5_addr_o[18]_pad  ;
	output \s5_addr_o[19]_pad  ;
	output \s5_addr_o[1]_pad  ;
	output \s5_addr_o[20]_pad  ;
	output \s5_addr_o[21]_pad  ;
	output \s5_addr_o[22]_pad  ;
	output \s5_addr_o[23]_pad  ;
	output \s5_addr_o[24]_pad  ;
	output \s5_addr_o[25]_pad  ;
	output \s5_addr_o[26]_pad  ;
	output \s5_addr_o[27]_pad  ;
	output \s5_addr_o[28]_pad  ;
	output \s5_addr_o[29]_pad  ;
	output \s5_addr_o[2]_pad  ;
	output \s5_addr_o[30]_pad  ;
	output \s5_addr_o[31]_pad  ;
	output \s5_addr_o[3]_pad  ;
	output \s5_addr_o[4]_pad  ;
	output \s5_addr_o[5]_pad  ;
	output \s5_addr_o[6]_pad  ;
	output \s5_addr_o[7]_pad  ;
	output \s5_addr_o[8]_pad  ;
	output \s5_addr_o[9]_pad  ;
	output \s5_data_o[0]_pad  ;
	output \s5_data_o[10]_pad  ;
	output \s5_data_o[11]_pad  ;
	output \s5_data_o[12]_pad  ;
	output \s5_data_o[13]_pad  ;
	output \s5_data_o[14]_pad  ;
	output \s5_data_o[15]_pad  ;
	output \s5_data_o[16]_pad  ;
	output \s5_data_o[17]_pad  ;
	output \s5_data_o[18]_pad  ;
	output \s5_data_o[19]_pad  ;
	output \s5_data_o[1]_pad  ;
	output \s5_data_o[20]_pad  ;
	output \s5_data_o[21]_pad  ;
	output \s5_data_o[22]_pad  ;
	output \s5_data_o[23]_pad  ;
	output \s5_data_o[24]_pad  ;
	output \s5_data_o[25]_pad  ;
	output \s5_data_o[26]_pad  ;
	output \s5_data_o[27]_pad  ;
	output \s5_data_o[28]_pad  ;
	output \s5_data_o[29]_pad  ;
	output \s5_data_o[2]_pad  ;
	output \s5_data_o[30]_pad  ;
	output \s5_data_o[31]_pad  ;
	output \s5_data_o[3]_pad  ;
	output \s5_data_o[4]_pad  ;
	output \s5_data_o[5]_pad  ;
	output \s5_data_o[6]_pad  ;
	output \s5_data_o[7]_pad  ;
	output \s5_data_o[8]_pad  ;
	output \s5_data_o[9]_pad  ;
	output \s5_sel_o[0]_pad  ;
	output \s5_sel_o[1]_pad  ;
	output \s5_sel_o[2]_pad  ;
	output \s5_sel_o[3]_pad  ;
	output \s5_stb_o_pad  ;
	output \s5_we_o_pad  ;
	output \s6_addr_o[0]_pad  ;
	output \s6_addr_o[10]_pad  ;
	output \s6_addr_o[11]_pad  ;
	output \s6_addr_o[12]_pad  ;
	output \s6_addr_o[13]_pad  ;
	output \s6_addr_o[14]_pad  ;
	output \s6_addr_o[15]_pad  ;
	output \s6_addr_o[16]_pad  ;
	output \s6_addr_o[17]_pad  ;
	output \s6_addr_o[18]_pad  ;
	output \s6_addr_o[19]_pad  ;
	output \s6_addr_o[1]_pad  ;
	output \s6_addr_o[20]_pad  ;
	output \s6_addr_o[21]_pad  ;
	output \s6_addr_o[22]_pad  ;
	output \s6_addr_o[23]_pad  ;
	output \s6_addr_o[24]_pad  ;
	output \s6_addr_o[25]_pad  ;
	output \s6_addr_o[26]_pad  ;
	output \s6_addr_o[27]_pad  ;
	output \s6_addr_o[28]_pad  ;
	output \s6_addr_o[29]_pad  ;
	output \s6_addr_o[2]_pad  ;
	output \s6_addr_o[30]_pad  ;
	output \s6_addr_o[31]_pad  ;
	output \s6_addr_o[3]_pad  ;
	output \s6_addr_o[4]_pad  ;
	output \s6_addr_o[5]_pad  ;
	output \s6_addr_o[6]_pad  ;
	output \s6_addr_o[7]_pad  ;
	output \s6_addr_o[8]_pad  ;
	output \s6_addr_o[9]_pad  ;
	output \s6_data_o[0]_pad  ;
	output \s6_data_o[10]_pad  ;
	output \s6_data_o[11]_pad  ;
	output \s6_data_o[12]_pad  ;
	output \s6_data_o[13]_pad  ;
	output \s6_data_o[14]_pad  ;
	output \s6_data_o[15]_pad  ;
	output \s6_data_o[16]_pad  ;
	output \s6_data_o[17]_pad  ;
	output \s6_data_o[18]_pad  ;
	output \s6_data_o[19]_pad  ;
	output \s6_data_o[1]_pad  ;
	output \s6_data_o[20]_pad  ;
	output \s6_data_o[21]_pad  ;
	output \s6_data_o[22]_pad  ;
	output \s6_data_o[23]_pad  ;
	output \s6_data_o[24]_pad  ;
	output \s6_data_o[25]_pad  ;
	output \s6_data_o[26]_pad  ;
	output \s6_data_o[27]_pad  ;
	output \s6_data_o[28]_pad  ;
	output \s6_data_o[29]_pad  ;
	output \s6_data_o[2]_pad  ;
	output \s6_data_o[30]_pad  ;
	output \s6_data_o[31]_pad  ;
	output \s6_data_o[3]_pad  ;
	output \s6_data_o[4]_pad  ;
	output \s6_data_o[5]_pad  ;
	output \s6_data_o[6]_pad  ;
	output \s6_data_o[7]_pad  ;
	output \s6_data_o[8]_pad  ;
	output \s6_data_o[9]_pad  ;
	output \s6_sel_o[0]_pad  ;
	output \s6_sel_o[1]_pad  ;
	output \s6_sel_o[2]_pad  ;
	output \s6_sel_o[3]_pad  ;
	output \s6_stb_o_pad  ;
	output \s6_we_o_pad  ;
	output \s7_addr_o[0]_pad  ;
	output \s7_addr_o[10]_pad  ;
	output \s7_addr_o[11]_pad  ;
	output \s7_addr_o[12]_pad  ;
	output \s7_addr_o[13]_pad  ;
	output \s7_addr_o[14]_pad  ;
	output \s7_addr_o[15]_pad  ;
	output \s7_addr_o[16]_pad  ;
	output \s7_addr_o[17]_pad  ;
	output \s7_addr_o[18]_pad  ;
	output \s7_addr_o[19]_pad  ;
	output \s7_addr_o[1]_pad  ;
	output \s7_addr_o[20]_pad  ;
	output \s7_addr_o[21]_pad  ;
	output \s7_addr_o[22]_pad  ;
	output \s7_addr_o[23]_pad  ;
	output \s7_addr_o[24]_pad  ;
	output \s7_addr_o[25]_pad  ;
	output \s7_addr_o[26]_pad  ;
	output \s7_addr_o[27]_pad  ;
	output \s7_addr_o[28]_pad  ;
	output \s7_addr_o[29]_pad  ;
	output \s7_addr_o[2]_pad  ;
	output \s7_addr_o[30]_pad  ;
	output \s7_addr_o[31]_pad  ;
	output \s7_addr_o[3]_pad  ;
	output \s7_addr_o[4]_pad  ;
	output \s7_addr_o[5]_pad  ;
	output \s7_addr_o[6]_pad  ;
	output \s7_addr_o[7]_pad  ;
	output \s7_addr_o[8]_pad  ;
	output \s7_addr_o[9]_pad  ;
	output \s7_data_o[0]_pad  ;
	output \s7_data_o[10]_pad  ;
	output \s7_data_o[11]_pad  ;
	output \s7_data_o[12]_pad  ;
	output \s7_data_o[13]_pad  ;
	output \s7_data_o[14]_pad  ;
	output \s7_data_o[15]_pad  ;
	output \s7_data_o[16]_pad  ;
	output \s7_data_o[17]_pad  ;
	output \s7_data_o[18]_pad  ;
	output \s7_data_o[19]_pad  ;
	output \s7_data_o[1]_pad  ;
	output \s7_data_o[20]_pad  ;
	output \s7_data_o[21]_pad  ;
	output \s7_data_o[22]_pad  ;
	output \s7_data_o[23]_pad  ;
	output \s7_data_o[24]_pad  ;
	output \s7_data_o[25]_pad  ;
	output \s7_data_o[26]_pad  ;
	output \s7_data_o[27]_pad  ;
	output \s7_data_o[28]_pad  ;
	output \s7_data_o[29]_pad  ;
	output \s7_data_o[2]_pad  ;
	output \s7_data_o[30]_pad  ;
	output \s7_data_o[31]_pad  ;
	output \s7_data_o[3]_pad  ;
	output \s7_data_o[4]_pad  ;
	output \s7_data_o[5]_pad  ;
	output \s7_data_o[6]_pad  ;
	output \s7_data_o[7]_pad  ;
	output \s7_data_o[8]_pad  ;
	output \s7_data_o[9]_pad  ;
	output \s7_sel_o[0]_pad  ;
	output \s7_sel_o[1]_pad  ;
	output \s7_sel_o[2]_pad  ;
	output \s7_sel_o[3]_pad  ;
	output \s7_stb_o_pad  ;
	output \s7_we_o_pad  ;
	output \s8_addr_o[0]_pad  ;
	output \s8_addr_o[10]_pad  ;
	output \s8_addr_o[11]_pad  ;
	output \s8_addr_o[12]_pad  ;
	output \s8_addr_o[13]_pad  ;
	output \s8_addr_o[14]_pad  ;
	output \s8_addr_o[15]_pad  ;
	output \s8_addr_o[16]_pad  ;
	output \s8_addr_o[17]_pad  ;
	output \s8_addr_o[18]_pad  ;
	output \s8_addr_o[19]_pad  ;
	output \s8_addr_o[1]_pad  ;
	output \s8_addr_o[20]_pad  ;
	output \s8_addr_o[21]_pad  ;
	output \s8_addr_o[22]_pad  ;
	output \s8_addr_o[23]_pad  ;
	output \s8_addr_o[24]_pad  ;
	output \s8_addr_o[25]_pad  ;
	output \s8_addr_o[26]_pad  ;
	output \s8_addr_o[27]_pad  ;
	output \s8_addr_o[28]_pad  ;
	output \s8_addr_o[29]_pad  ;
	output \s8_addr_o[2]_pad  ;
	output \s8_addr_o[30]_pad  ;
	output \s8_addr_o[31]_pad  ;
	output \s8_addr_o[3]_pad  ;
	output \s8_addr_o[4]_pad  ;
	output \s8_addr_o[5]_pad  ;
	output \s8_addr_o[6]_pad  ;
	output \s8_addr_o[7]_pad  ;
	output \s8_addr_o[8]_pad  ;
	output \s8_addr_o[9]_pad  ;
	output \s8_data_o[0]_pad  ;
	output \s8_data_o[10]_pad  ;
	output \s8_data_o[11]_pad  ;
	output \s8_data_o[12]_pad  ;
	output \s8_data_o[13]_pad  ;
	output \s8_data_o[14]_pad  ;
	output \s8_data_o[15]_pad  ;
	output \s8_data_o[16]_pad  ;
	output \s8_data_o[17]_pad  ;
	output \s8_data_o[18]_pad  ;
	output \s8_data_o[19]_pad  ;
	output \s8_data_o[1]_pad  ;
	output \s8_data_o[20]_pad  ;
	output \s8_data_o[21]_pad  ;
	output \s8_data_o[22]_pad  ;
	output \s8_data_o[23]_pad  ;
	output \s8_data_o[24]_pad  ;
	output \s8_data_o[25]_pad  ;
	output \s8_data_o[26]_pad  ;
	output \s8_data_o[27]_pad  ;
	output \s8_data_o[28]_pad  ;
	output \s8_data_o[29]_pad  ;
	output \s8_data_o[2]_pad  ;
	output \s8_data_o[30]_pad  ;
	output \s8_data_o[31]_pad  ;
	output \s8_data_o[3]_pad  ;
	output \s8_data_o[4]_pad  ;
	output \s8_data_o[5]_pad  ;
	output \s8_data_o[6]_pad  ;
	output \s8_data_o[7]_pad  ;
	output \s8_data_o[8]_pad  ;
	output \s8_data_o[9]_pad  ;
	output \s8_sel_o[0]_pad  ;
	output \s8_sel_o[1]_pad  ;
	output \s8_sel_o[2]_pad  ;
	output \s8_sel_o[3]_pad  ;
	output \s8_stb_o_pad  ;
	output \s8_we_o_pad  ;
	output \s9_addr_o[0]_pad  ;
	output \s9_addr_o[10]_pad  ;
	output \s9_addr_o[11]_pad  ;
	output \s9_addr_o[12]_pad  ;
	output \s9_addr_o[13]_pad  ;
	output \s9_addr_o[14]_pad  ;
	output \s9_addr_o[15]_pad  ;
	output \s9_addr_o[16]_pad  ;
	output \s9_addr_o[17]_pad  ;
	output \s9_addr_o[18]_pad  ;
	output \s9_addr_o[19]_pad  ;
	output \s9_addr_o[1]_pad  ;
	output \s9_addr_o[20]_pad  ;
	output \s9_addr_o[21]_pad  ;
	output \s9_addr_o[22]_pad  ;
	output \s9_addr_o[23]_pad  ;
	output \s9_addr_o[24]_pad  ;
	output \s9_addr_o[25]_pad  ;
	output \s9_addr_o[26]_pad  ;
	output \s9_addr_o[27]_pad  ;
	output \s9_addr_o[28]_pad  ;
	output \s9_addr_o[29]_pad  ;
	output \s9_addr_o[2]_pad  ;
	output \s9_addr_o[30]_pad  ;
	output \s9_addr_o[31]_pad  ;
	output \s9_addr_o[3]_pad  ;
	output \s9_addr_o[4]_pad  ;
	output \s9_addr_o[5]_pad  ;
	output \s9_addr_o[6]_pad  ;
	output \s9_addr_o[7]_pad  ;
	output \s9_addr_o[8]_pad  ;
	output \s9_addr_o[9]_pad  ;
	output \s9_data_o[0]_pad  ;
	output \s9_data_o[10]_pad  ;
	output \s9_data_o[11]_pad  ;
	output \s9_data_o[12]_pad  ;
	output \s9_data_o[13]_pad  ;
	output \s9_data_o[14]_pad  ;
	output \s9_data_o[15]_pad  ;
	output \s9_data_o[16]_pad  ;
	output \s9_data_o[17]_pad  ;
	output \s9_data_o[18]_pad  ;
	output \s9_data_o[19]_pad  ;
	output \s9_data_o[1]_pad  ;
	output \s9_data_o[20]_pad  ;
	output \s9_data_o[21]_pad  ;
	output \s9_data_o[22]_pad  ;
	output \s9_data_o[23]_pad  ;
	output \s9_data_o[24]_pad  ;
	output \s9_data_o[25]_pad  ;
	output \s9_data_o[26]_pad  ;
	output \s9_data_o[27]_pad  ;
	output \s9_data_o[28]_pad  ;
	output \s9_data_o[29]_pad  ;
	output \s9_data_o[2]_pad  ;
	output \s9_data_o[30]_pad  ;
	output \s9_data_o[31]_pad  ;
	output \s9_data_o[3]_pad  ;
	output \s9_data_o[4]_pad  ;
	output \s9_data_o[5]_pad  ;
	output \s9_data_o[6]_pad  ;
	output \s9_data_o[7]_pad  ;
	output \s9_data_o[8]_pad  ;
	output \s9_data_o[9]_pad  ;
	output \s9_sel_o[0]_pad  ;
	output \s9_sel_o[1]_pad  ;
	output \s9_sel_o[2]_pad  ;
	output \s9_sel_o[3]_pad  ;
	output \s9_stb_o_pad  ;
	output \s9_we_o_pad  ;
	wire _w28163_ ;
	wire _w28162_ ;
	wire _w28161_ ;
	wire _w28160_ ;
	wire _w28159_ ;
	wire _w28158_ ;
	wire _w28157_ ;
	wire _w28156_ ;
	wire _w28155_ ;
	wire _w28154_ ;
	wire _w28153_ ;
	wire _w28152_ ;
	wire _w28151_ ;
	wire _w28150_ ;
	wire _w28149_ ;
	wire _w28148_ ;
	wire _w28147_ ;
	wire _w28146_ ;
	wire _w28145_ ;
	wire _w28144_ ;
	wire _w28143_ ;
	wire _w28142_ ;
	wire _w28141_ ;
	wire _w28140_ ;
	wire _w28139_ ;
	wire _w28138_ ;
	wire _w28137_ ;
	wire _w28136_ ;
	wire _w28135_ ;
	wire _w28134_ ;
	wire _w28133_ ;
	wire _w28132_ ;
	wire _w28131_ ;
	wire _w28130_ ;
	wire _w28129_ ;
	wire _w28128_ ;
	wire _w28127_ ;
	wire _w28126_ ;
	wire _w28125_ ;
	wire _w28124_ ;
	wire _w28123_ ;
	wire _w28122_ ;
	wire _w28121_ ;
	wire _w28120_ ;
	wire _w28119_ ;
	wire _w28118_ ;
	wire _w28117_ ;
	wire _w28116_ ;
	wire _w28115_ ;
	wire _w28114_ ;
	wire _w28113_ ;
	wire _w28112_ ;
	wire _w28111_ ;
	wire _w28110_ ;
	wire _w28109_ ;
	wire _w28108_ ;
	wire _w28107_ ;
	wire _w28106_ ;
	wire _w28105_ ;
	wire _w28104_ ;
	wire _w28103_ ;
	wire _w28102_ ;
	wire _w28101_ ;
	wire _w28100_ ;
	wire _w28099_ ;
	wire _w28098_ ;
	wire _w28097_ ;
	wire _w28096_ ;
	wire _w28095_ ;
	wire _w28094_ ;
	wire _w28093_ ;
	wire _w28092_ ;
	wire _w28091_ ;
	wire _w28090_ ;
	wire _w28089_ ;
	wire _w28088_ ;
	wire _w28087_ ;
	wire _w28086_ ;
	wire _w28085_ ;
	wire _w28084_ ;
	wire _w28083_ ;
	wire _w28082_ ;
	wire _w28081_ ;
	wire _w28080_ ;
	wire _w28079_ ;
	wire _w28078_ ;
	wire _w28077_ ;
	wire _w28076_ ;
	wire _w28075_ ;
	wire _w28074_ ;
	wire _w28073_ ;
	wire _w28072_ ;
	wire _w28071_ ;
	wire _w28070_ ;
	wire _w28069_ ;
	wire _w28068_ ;
	wire _w28067_ ;
	wire _w28066_ ;
	wire _w28065_ ;
	wire _w28064_ ;
	wire _w28063_ ;
	wire _w28062_ ;
	wire _w28061_ ;
	wire _w28060_ ;
	wire _w28059_ ;
	wire _w28058_ ;
	wire _w28057_ ;
	wire _w28056_ ;
	wire _w28055_ ;
	wire _w28054_ ;
	wire _w28053_ ;
	wire _w28052_ ;
	wire _w28051_ ;
	wire _w28050_ ;
	wire _w28049_ ;
	wire _w28048_ ;
	wire _w28047_ ;
	wire _w28046_ ;
	wire _w28045_ ;
	wire _w28044_ ;
	wire _w28043_ ;
	wire _w28042_ ;
	wire _w28041_ ;
	wire _w28040_ ;
	wire _w28039_ ;
	wire _w28038_ ;
	wire _w28037_ ;
	wire _w28036_ ;
	wire _w28035_ ;
	wire _w28034_ ;
	wire _w28033_ ;
	wire _w28032_ ;
	wire _w28031_ ;
	wire _w28030_ ;
	wire _w28029_ ;
	wire _w28028_ ;
	wire _w28027_ ;
	wire _w28026_ ;
	wire _w28025_ ;
	wire _w28024_ ;
	wire _w28023_ ;
	wire _w28022_ ;
	wire _w28021_ ;
	wire _w28020_ ;
	wire _w28019_ ;
	wire _w28018_ ;
	wire _w28017_ ;
	wire _w28016_ ;
	wire _w28015_ ;
	wire _w28014_ ;
	wire _w28013_ ;
	wire _w28012_ ;
	wire _w28011_ ;
	wire _w28010_ ;
	wire _w28009_ ;
	wire _w28008_ ;
	wire _w28007_ ;
	wire _w28006_ ;
	wire _w28005_ ;
	wire _w28004_ ;
	wire _w28003_ ;
	wire _w28002_ ;
	wire _w28001_ ;
	wire _w28000_ ;
	wire _w27999_ ;
	wire _w27998_ ;
	wire _w27997_ ;
	wire _w27996_ ;
	wire _w27995_ ;
	wire _w27994_ ;
	wire _w27993_ ;
	wire _w27992_ ;
	wire _w27991_ ;
	wire _w27990_ ;
	wire _w27989_ ;
	wire _w27988_ ;
	wire _w27987_ ;
	wire _w27986_ ;
	wire _w27985_ ;
	wire _w27984_ ;
	wire _w27983_ ;
	wire _w27982_ ;
	wire _w27981_ ;
	wire _w27980_ ;
	wire _w27979_ ;
	wire _w27978_ ;
	wire _w27977_ ;
	wire _w27976_ ;
	wire _w27975_ ;
	wire _w27974_ ;
	wire _w27973_ ;
	wire _w27972_ ;
	wire _w27971_ ;
	wire _w27970_ ;
	wire _w27969_ ;
	wire _w27968_ ;
	wire _w27967_ ;
	wire _w27966_ ;
	wire _w27965_ ;
	wire _w27964_ ;
	wire _w27963_ ;
	wire _w27962_ ;
	wire _w27961_ ;
	wire _w27960_ ;
	wire _w27959_ ;
	wire _w27958_ ;
	wire _w27957_ ;
	wire _w27956_ ;
	wire _w27955_ ;
	wire _w27954_ ;
	wire _w27953_ ;
	wire _w27952_ ;
	wire _w27951_ ;
	wire _w27950_ ;
	wire _w27949_ ;
	wire _w27948_ ;
	wire _w27947_ ;
	wire _w27946_ ;
	wire _w27945_ ;
	wire _w27944_ ;
	wire _w27943_ ;
	wire _w27942_ ;
	wire _w27941_ ;
	wire _w27940_ ;
	wire _w27939_ ;
	wire _w27938_ ;
	wire _w27937_ ;
	wire _w27936_ ;
	wire _w27935_ ;
	wire _w27934_ ;
	wire _w27933_ ;
	wire _w27932_ ;
	wire _w27931_ ;
	wire _w27930_ ;
	wire _w27929_ ;
	wire _w27928_ ;
	wire _w27927_ ;
	wire _w27926_ ;
	wire _w27925_ ;
	wire _w27924_ ;
	wire _w27923_ ;
	wire _w27922_ ;
	wire _w27921_ ;
	wire _w27920_ ;
	wire _w27919_ ;
	wire _w27918_ ;
	wire _w27917_ ;
	wire _w27916_ ;
	wire _w27915_ ;
	wire _w27914_ ;
	wire _w27913_ ;
	wire _w27912_ ;
	wire _w27911_ ;
	wire _w27910_ ;
	wire _w27909_ ;
	wire _w27908_ ;
	wire _w27907_ ;
	wire _w27906_ ;
	wire _w27905_ ;
	wire _w27904_ ;
	wire _w27903_ ;
	wire _w27902_ ;
	wire _w27901_ ;
	wire _w27900_ ;
	wire _w27899_ ;
	wire _w27898_ ;
	wire _w27897_ ;
	wire _w27896_ ;
	wire _w27895_ ;
	wire _w27894_ ;
	wire _w27893_ ;
	wire _w27892_ ;
	wire _w27891_ ;
	wire _w27890_ ;
	wire _w27889_ ;
	wire _w27888_ ;
	wire _w27887_ ;
	wire _w27886_ ;
	wire _w27885_ ;
	wire _w27884_ ;
	wire _w27883_ ;
	wire _w27882_ ;
	wire _w27881_ ;
	wire _w27880_ ;
	wire _w27879_ ;
	wire _w27878_ ;
	wire _w27877_ ;
	wire _w27876_ ;
	wire _w27875_ ;
	wire _w27874_ ;
	wire _w27873_ ;
	wire _w27872_ ;
	wire _w27871_ ;
	wire _w27870_ ;
	wire _w27869_ ;
	wire _w27868_ ;
	wire _w27867_ ;
	wire _w27866_ ;
	wire _w27865_ ;
	wire _w27864_ ;
	wire _w27863_ ;
	wire _w27862_ ;
	wire _w27861_ ;
	wire _w27860_ ;
	wire _w27859_ ;
	wire _w27858_ ;
	wire _w27857_ ;
	wire _w27856_ ;
	wire _w27855_ ;
	wire _w27854_ ;
	wire _w27853_ ;
	wire _w27852_ ;
	wire _w27851_ ;
	wire _w27850_ ;
	wire _w27849_ ;
	wire _w27848_ ;
	wire _w27847_ ;
	wire _w27846_ ;
	wire _w27845_ ;
	wire _w27844_ ;
	wire _w27843_ ;
	wire _w27842_ ;
	wire _w27841_ ;
	wire _w27840_ ;
	wire _w27839_ ;
	wire _w27838_ ;
	wire _w27837_ ;
	wire _w27836_ ;
	wire _w27835_ ;
	wire _w27834_ ;
	wire _w27833_ ;
	wire _w27832_ ;
	wire _w27831_ ;
	wire _w27830_ ;
	wire _w27829_ ;
	wire _w27828_ ;
	wire _w27827_ ;
	wire _w27826_ ;
	wire _w27825_ ;
	wire _w27824_ ;
	wire _w27823_ ;
	wire _w27822_ ;
	wire _w27821_ ;
	wire _w27820_ ;
	wire _w27819_ ;
	wire _w27818_ ;
	wire _w27817_ ;
	wire _w27816_ ;
	wire _w27815_ ;
	wire _w27814_ ;
	wire _w27813_ ;
	wire _w27812_ ;
	wire _w27811_ ;
	wire _w27810_ ;
	wire _w27809_ ;
	wire _w27808_ ;
	wire _w27807_ ;
	wire _w27806_ ;
	wire _w27805_ ;
	wire _w27804_ ;
	wire _w27803_ ;
	wire _w27802_ ;
	wire _w27801_ ;
	wire _w27800_ ;
	wire _w27799_ ;
	wire _w27798_ ;
	wire _w27797_ ;
	wire _w27796_ ;
	wire _w27795_ ;
	wire _w27794_ ;
	wire _w27793_ ;
	wire _w27792_ ;
	wire _w27791_ ;
	wire _w27790_ ;
	wire _w27789_ ;
	wire _w27788_ ;
	wire _w27787_ ;
	wire _w27786_ ;
	wire _w27785_ ;
	wire _w27784_ ;
	wire _w27783_ ;
	wire _w27782_ ;
	wire _w27781_ ;
	wire _w27780_ ;
	wire _w27779_ ;
	wire _w27778_ ;
	wire _w27777_ ;
	wire _w27776_ ;
	wire _w27775_ ;
	wire _w27774_ ;
	wire _w27773_ ;
	wire _w27772_ ;
	wire _w27771_ ;
	wire _w27770_ ;
	wire _w27769_ ;
	wire _w27768_ ;
	wire _w27767_ ;
	wire _w27766_ ;
	wire _w27765_ ;
	wire _w27764_ ;
	wire _w27763_ ;
	wire _w27762_ ;
	wire _w27761_ ;
	wire _w27760_ ;
	wire _w27759_ ;
	wire _w27758_ ;
	wire _w27757_ ;
	wire _w27756_ ;
	wire _w27755_ ;
	wire _w27754_ ;
	wire _w27753_ ;
	wire _w27752_ ;
	wire _w27751_ ;
	wire _w27750_ ;
	wire _w27749_ ;
	wire _w27748_ ;
	wire _w27747_ ;
	wire _w27746_ ;
	wire _w27745_ ;
	wire _w27744_ ;
	wire _w27743_ ;
	wire _w27742_ ;
	wire _w27741_ ;
	wire _w27740_ ;
	wire _w27739_ ;
	wire _w27738_ ;
	wire _w27737_ ;
	wire _w27736_ ;
	wire _w27735_ ;
	wire _w27734_ ;
	wire _w27733_ ;
	wire _w27732_ ;
	wire _w27731_ ;
	wire _w27730_ ;
	wire _w27729_ ;
	wire _w27728_ ;
	wire _w27727_ ;
	wire _w27726_ ;
	wire _w27725_ ;
	wire _w27724_ ;
	wire _w27723_ ;
	wire _w27722_ ;
	wire _w27721_ ;
	wire _w27720_ ;
	wire _w27719_ ;
	wire _w27718_ ;
	wire _w27717_ ;
	wire _w27716_ ;
	wire _w27715_ ;
	wire _w27714_ ;
	wire _w27713_ ;
	wire _w27712_ ;
	wire _w27711_ ;
	wire _w27710_ ;
	wire _w27709_ ;
	wire _w27708_ ;
	wire _w27707_ ;
	wire _w27706_ ;
	wire _w27705_ ;
	wire _w27704_ ;
	wire _w27703_ ;
	wire _w27702_ ;
	wire _w27701_ ;
	wire _w27700_ ;
	wire _w27699_ ;
	wire _w27698_ ;
	wire _w27697_ ;
	wire _w27696_ ;
	wire _w27695_ ;
	wire _w27694_ ;
	wire _w27693_ ;
	wire _w27692_ ;
	wire _w27691_ ;
	wire _w27690_ ;
	wire _w27689_ ;
	wire _w27688_ ;
	wire _w27687_ ;
	wire _w27686_ ;
	wire _w27685_ ;
	wire _w27684_ ;
	wire _w27683_ ;
	wire _w27682_ ;
	wire _w27681_ ;
	wire _w27680_ ;
	wire _w27679_ ;
	wire _w27678_ ;
	wire _w27677_ ;
	wire _w27676_ ;
	wire _w27675_ ;
	wire _w27674_ ;
	wire _w27673_ ;
	wire _w27672_ ;
	wire _w27671_ ;
	wire _w27670_ ;
	wire _w27669_ ;
	wire _w27668_ ;
	wire _w27667_ ;
	wire _w27666_ ;
	wire _w27665_ ;
	wire _w27664_ ;
	wire _w27663_ ;
	wire _w27662_ ;
	wire _w27661_ ;
	wire _w27660_ ;
	wire _w27659_ ;
	wire _w27658_ ;
	wire _w27657_ ;
	wire _w27656_ ;
	wire _w27655_ ;
	wire _w27654_ ;
	wire _w27653_ ;
	wire _w27652_ ;
	wire _w27651_ ;
	wire _w27650_ ;
	wire _w27649_ ;
	wire _w27648_ ;
	wire _w27647_ ;
	wire _w27646_ ;
	wire _w27645_ ;
	wire _w27644_ ;
	wire _w27643_ ;
	wire _w27642_ ;
	wire _w27641_ ;
	wire _w27640_ ;
	wire _w27639_ ;
	wire _w27638_ ;
	wire _w27637_ ;
	wire _w27636_ ;
	wire _w27635_ ;
	wire _w27634_ ;
	wire _w27633_ ;
	wire _w27632_ ;
	wire _w27631_ ;
	wire _w27630_ ;
	wire _w27629_ ;
	wire _w27628_ ;
	wire _w27627_ ;
	wire _w27626_ ;
	wire _w27625_ ;
	wire _w27624_ ;
	wire _w27623_ ;
	wire _w27622_ ;
	wire _w27621_ ;
	wire _w27620_ ;
	wire _w27619_ ;
	wire _w27618_ ;
	wire _w27617_ ;
	wire _w27616_ ;
	wire _w27615_ ;
	wire _w27614_ ;
	wire _w27613_ ;
	wire _w27612_ ;
	wire _w27611_ ;
	wire _w27610_ ;
	wire _w27609_ ;
	wire _w27608_ ;
	wire _w27607_ ;
	wire _w27606_ ;
	wire _w27605_ ;
	wire _w27604_ ;
	wire _w27603_ ;
	wire _w27602_ ;
	wire _w27601_ ;
	wire _w27600_ ;
	wire _w27599_ ;
	wire _w27598_ ;
	wire _w27597_ ;
	wire _w27596_ ;
	wire _w27595_ ;
	wire _w27594_ ;
	wire _w27593_ ;
	wire _w27592_ ;
	wire _w27591_ ;
	wire _w27590_ ;
	wire _w27589_ ;
	wire _w27588_ ;
	wire _w27587_ ;
	wire _w27586_ ;
	wire _w27585_ ;
	wire _w27584_ ;
	wire _w27583_ ;
	wire _w27582_ ;
	wire _w27581_ ;
	wire _w27580_ ;
	wire _w27579_ ;
	wire _w27578_ ;
	wire _w27577_ ;
	wire _w27576_ ;
	wire _w27575_ ;
	wire _w27574_ ;
	wire _w27573_ ;
	wire _w27572_ ;
	wire _w27571_ ;
	wire _w27570_ ;
	wire _w27569_ ;
	wire _w27568_ ;
	wire _w27567_ ;
	wire _w27566_ ;
	wire _w27565_ ;
	wire _w27564_ ;
	wire _w27563_ ;
	wire _w27562_ ;
	wire _w27561_ ;
	wire _w27560_ ;
	wire _w27559_ ;
	wire _w27558_ ;
	wire _w27557_ ;
	wire _w27556_ ;
	wire _w27555_ ;
	wire _w27554_ ;
	wire _w27553_ ;
	wire _w27552_ ;
	wire _w27551_ ;
	wire _w27550_ ;
	wire _w27549_ ;
	wire _w27548_ ;
	wire _w27547_ ;
	wire _w27546_ ;
	wire _w27545_ ;
	wire _w27544_ ;
	wire _w27543_ ;
	wire _w27542_ ;
	wire _w27541_ ;
	wire _w27540_ ;
	wire _w27539_ ;
	wire _w27538_ ;
	wire _w27537_ ;
	wire _w27536_ ;
	wire _w27535_ ;
	wire _w27534_ ;
	wire _w27533_ ;
	wire _w27532_ ;
	wire _w27531_ ;
	wire _w27530_ ;
	wire _w27529_ ;
	wire _w27528_ ;
	wire _w27527_ ;
	wire _w27526_ ;
	wire _w27525_ ;
	wire _w27524_ ;
	wire _w27523_ ;
	wire _w27522_ ;
	wire _w27521_ ;
	wire _w27520_ ;
	wire _w27519_ ;
	wire _w27518_ ;
	wire _w27517_ ;
	wire _w27516_ ;
	wire _w27515_ ;
	wire _w27514_ ;
	wire _w27513_ ;
	wire _w27512_ ;
	wire _w27511_ ;
	wire _w27510_ ;
	wire _w27509_ ;
	wire _w27508_ ;
	wire _w27507_ ;
	wire _w27506_ ;
	wire _w27505_ ;
	wire _w27504_ ;
	wire _w27503_ ;
	wire _w27502_ ;
	wire _w27501_ ;
	wire _w27500_ ;
	wire _w27499_ ;
	wire _w27498_ ;
	wire _w27497_ ;
	wire _w27496_ ;
	wire _w27495_ ;
	wire _w27494_ ;
	wire _w27493_ ;
	wire _w27492_ ;
	wire _w27491_ ;
	wire _w27490_ ;
	wire _w27489_ ;
	wire _w27488_ ;
	wire _w27487_ ;
	wire _w27486_ ;
	wire _w27485_ ;
	wire _w27484_ ;
	wire _w27483_ ;
	wire _w27482_ ;
	wire _w27481_ ;
	wire _w27480_ ;
	wire _w27479_ ;
	wire _w27478_ ;
	wire _w27477_ ;
	wire _w27476_ ;
	wire _w27475_ ;
	wire _w27474_ ;
	wire _w27473_ ;
	wire _w27472_ ;
	wire _w27471_ ;
	wire _w27470_ ;
	wire _w27469_ ;
	wire _w27468_ ;
	wire _w27467_ ;
	wire _w27466_ ;
	wire _w27465_ ;
	wire _w27464_ ;
	wire _w27463_ ;
	wire _w27462_ ;
	wire _w27461_ ;
	wire _w27460_ ;
	wire _w27459_ ;
	wire _w27458_ ;
	wire _w27457_ ;
	wire _w27456_ ;
	wire _w27455_ ;
	wire _w27454_ ;
	wire _w27453_ ;
	wire _w27452_ ;
	wire _w27451_ ;
	wire _w27450_ ;
	wire _w27449_ ;
	wire _w27448_ ;
	wire _w27447_ ;
	wire _w27446_ ;
	wire _w27445_ ;
	wire _w27444_ ;
	wire _w27443_ ;
	wire _w27442_ ;
	wire _w27441_ ;
	wire _w27440_ ;
	wire _w27439_ ;
	wire _w27438_ ;
	wire _w27437_ ;
	wire _w27436_ ;
	wire _w27435_ ;
	wire _w27434_ ;
	wire _w27433_ ;
	wire _w27432_ ;
	wire _w27431_ ;
	wire _w27430_ ;
	wire _w27429_ ;
	wire _w27428_ ;
	wire _w27427_ ;
	wire _w27426_ ;
	wire _w27425_ ;
	wire _w27424_ ;
	wire _w27423_ ;
	wire _w27422_ ;
	wire _w27421_ ;
	wire _w27420_ ;
	wire _w27419_ ;
	wire _w27418_ ;
	wire _w27417_ ;
	wire _w27416_ ;
	wire _w27415_ ;
	wire _w27414_ ;
	wire _w27413_ ;
	wire _w27412_ ;
	wire _w27411_ ;
	wire _w27410_ ;
	wire _w27409_ ;
	wire _w27408_ ;
	wire _w27407_ ;
	wire _w27406_ ;
	wire _w27405_ ;
	wire _w27404_ ;
	wire _w27403_ ;
	wire _w27402_ ;
	wire _w27401_ ;
	wire _w27400_ ;
	wire _w27399_ ;
	wire _w27398_ ;
	wire _w27397_ ;
	wire _w27396_ ;
	wire _w27395_ ;
	wire _w27394_ ;
	wire _w27393_ ;
	wire _w27392_ ;
	wire _w27391_ ;
	wire _w27390_ ;
	wire _w27389_ ;
	wire _w27388_ ;
	wire _w27387_ ;
	wire _w27386_ ;
	wire _w27385_ ;
	wire _w27384_ ;
	wire _w27383_ ;
	wire _w27382_ ;
	wire _w27381_ ;
	wire _w27380_ ;
	wire _w27379_ ;
	wire _w27378_ ;
	wire _w27377_ ;
	wire _w27376_ ;
	wire _w27375_ ;
	wire _w27374_ ;
	wire _w27373_ ;
	wire _w27372_ ;
	wire _w27371_ ;
	wire _w27370_ ;
	wire _w27369_ ;
	wire _w27368_ ;
	wire _w27367_ ;
	wire _w27366_ ;
	wire _w27365_ ;
	wire _w27364_ ;
	wire _w27363_ ;
	wire _w27362_ ;
	wire _w27361_ ;
	wire _w27360_ ;
	wire _w27359_ ;
	wire _w27358_ ;
	wire _w27357_ ;
	wire _w27356_ ;
	wire _w27355_ ;
	wire _w27354_ ;
	wire _w27353_ ;
	wire _w27352_ ;
	wire _w27351_ ;
	wire _w27350_ ;
	wire _w27349_ ;
	wire _w27348_ ;
	wire _w27347_ ;
	wire _w27346_ ;
	wire _w27345_ ;
	wire _w27344_ ;
	wire _w27343_ ;
	wire _w27342_ ;
	wire _w27341_ ;
	wire _w27340_ ;
	wire _w27339_ ;
	wire _w27338_ ;
	wire _w27337_ ;
	wire _w27336_ ;
	wire _w27335_ ;
	wire _w27334_ ;
	wire _w27333_ ;
	wire _w27332_ ;
	wire _w27331_ ;
	wire _w27330_ ;
	wire _w27329_ ;
	wire _w27328_ ;
	wire _w27327_ ;
	wire _w27326_ ;
	wire _w27325_ ;
	wire _w27324_ ;
	wire _w27323_ ;
	wire _w27322_ ;
	wire _w27321_ ;
	wire _w27320_ ;
	wire _w27319_ ;
	wire _w27318_ ;
	wire _w27317_ ;
	wire _w27316_ ;
	wire _w27315_ ;
	wire _w27314_ ;
	wire _w27313_ ;
	wire _w27312_ ;
	wire _w27311_ ;
	wire _w27310_ ;
	wire _w27309_ ;
	wire _w27308_ ;
	wire _w27307_ ;
	wire _w27306_ ;
	wire _w27305_ ;
	wire _w27304_ ;
	wire _w27303_ ;
	wire _w27302_ ;
	wire _w27301_ ;
	wire _w27300_ ;
	wire _w27299_ ;
	wire _w27298_ ;
	wire _w27297_ ;
	wire _w27296_ ;
	wire _w27295_ ;
	wire _w27294_ ;
	wire _w27293_ ;
	wire _w27292_ ;
	wire _w27291_ ;
	wire _w27290_ ;
	wire _w27289_ ;
	wire _w27288_ ;
	wire _w27287_ ;
	wire _w27286_ ;
	wire _w27285_ ;
	wire _w27284_ ;
	wire _w27283_ ;
	wire _w27282_ ;
	wire _w27281_ ;
	wire _w27280_ ;
	wire _w27279_ ;
	wire _w27278_ ;
	wire _w27277_ ;
	wire _w27276_ ;
	wire _w27275_ ;
	wire _w27274_ ;
	wire _w27273_ ;
	wire _w27272_ ;
	wire _w27271_ ;
	wire _w27270_ ;
	wire _w27269_ ;
	wire _w27268_ ;
	wire _w27267_ ;
	wire _w27266_ ;
	wire _w27265_ ;
	wire _w27264_ ;
	wire _w27263_ ;
	wire _w27262_ ;
	wire _w27261_ ;
	wire _w27260_ ;
	wire _w27259_ ;
	wire _w27258_ ;
	wire _w27257_ ;
	wire _w27256_ ;
	wire _w27255_ ;
	wire _w27254_ ;
	wire _w27253_ ;
	wire _w27252_ ;
	wire _w27251_ ;
	wire _w27250_ ;
	wire _w27249_ ;
	wire _w27248_ ;
	wire _w27247_ ;
	wire _w27246_ ;
	wire _w27245_ ;
	wire _w27244_ ;
	wire _w27243_ ;
	wire _w27242_ ;
	wire _w27241_ ;
	wire _w27240_ ;
	wire _w27239_ ;
	wire _w27238_ ;
	wire _w27237_ ;
	wire _w27236_ ;
	wire _w27235_ ;
	wire _w27234_ ;
	wire _w27233_ ;
	wire _w27232_ ;
	wire _w27231_ ;
	wire _w27230_ ;
	wire _w27229_ ;
	wire _w27228_ ;
	wire _w27227_ ;
	wire _w27226_ ;
	wire _w27225_ ;
	wire _w27224_ ;
	wire _w27223_ ;
	wire _w27222_ ;
	wire _w27221_ ;
	wire _w27220_ ;
	wire _w27219_ ;
	wire _w27218_ ;
	wire _w27217_ ;
	wire _w27216_ ;
	wire _w27215_ ;
	wire _w27214_ ;
	wire _w27213_ ;
	wire _w27212_ ;
	wire _w27211_ ;
	wire _w27210_ ;
	wire _w27209_ ;
	wire _w27208_ ;
	wire _w27207_ ;
	wire _w27206_ ;
	wire _w27205_ ;
	wire _w27204_ ;
	wire _w27203_ ;
	wire _w27202_ ;
	wire _w27201_ ;
	wire _w27200_ ;
	wire _w27199_ ;
	wire _w27198_ ;
	wire _w27197_ ;
	wire _w27196_ ;
	wire _w27195_ ;
	wire _w27194_ ;
	wire _w27193_ ;
	wire _w27192_ ;
	wire _w27191_ ;
	wire _w27190_ ;
	wire _w27189_ ;
	wire _w27188_ ;
	wire _w27187_ ;
	wire _w27186_ ;
	wire _w27185_ ;
	wire _w27184_ ;
	wire _w27183_ ;
	wire _w27182_ ;
	wire _w27181_ ;
	wire _w27180_ ;
	wire _w27179_ ;
	wire _w27178_ ;
	wire _w27177_ ;
	wire _w27176_ ;
	wire _w27175_ ;
	wire _w27174_ ;
	wire _w27173_ ;
	wire _w27172_ ;
	wire _w27171_ ;
	wire _w27170_ ;
	wire _w27169_ ;
	wire _w27168_ ;
	wire _w27167_ ;
	wire _w27166_ ;
	wire _w27165_ ;
	wire _w27164_ ;
	wire _w27163_ ;
	wire _w27162_ ;
	wire _w27161_ ;
	wire _w27160_ ;
	wire _w27159_ ;
	wire _w27158_ ;
	wire _w27157_ ;
	wire _w27156_ ;
	wire _w27155_ ;
	wire _w27154_ ;
	wire _w27153_ ;
	wire _w27152_ ;
	wire _w27151_ ;
	wire _w27150_ ;
	wire _w27149_ ;
	wire _w27148_ ;
	wire _w27147_ ;
	wire _w27146_ ;
	wire _w27145_ ;
	wire _w27144_ ;
	wire _w27143_ ;
	wire _w27142_ ;
	wire _w27141_ ;
	wire _w27140_ ;
	wire _w27139_ ;
	wire _w27138_ ;
	wire _w27137_ ;
	wire _w27136_ ;
	wire _w27135_ ;
	wire _w27134_ ;
	wire _w27133_ ;
	wire _w27132_ ;
	wire _w27131_ ;
	wire _w27130_ ;
	wire _w27129_ ;
	wire _w27128_ ;
	wire _w27127_ ;
	wire _w27126_ ;
	wire _w27125_ ;
	wire _w27124_ ;
	wire _w27123_ ;
	wire _w27122_ ;
	wire _w27121_ ;
	wire _w27120_ ;
	wire _w27119_ ;
	wire _w27118_ ;
	wire _w27117_ ;
	wire _w27116_ ;
	wire _w27115_ ;
	wire _w27114_ ;
	wire _w27113_ ;
	wire _w27112_ ;
	wire _w27111_ ;
	wire _w27110_ ;
	wire _w27109_ ;
	wire _w27108_ ;
	wire _w27107_ ;
	wire _w27106_ ;
	wire _w27105_ ;
	wire _w27104_ ;
	wire _w27103_ ;
	wire _w27102_ ;
	wire _w27101_ ;
	wire _w27100_ ;
	wire _w27099_ ;
	wire _w27098_ ;
	wire _w27097_ ;
	wire _w27096_ ;
	wire _w27095_ ;
	wire _w27094_ ;
	wire _w27093_ ;
	wire _w27092_ ;
	wire _w27091_ ;
	wire _w27090_ ;
	wire _w27089_ ;
	wire _w27088_ ;
	wire _w27087_ ;
	wire _w27086_ ;
	wire _w27085_ ;
	wire _w27084_ ;
	wire _w27083_ ;
	wire _w27082_ ;
	wire _w27081_ ;
	wire _w27080_ ;
	wire _w27079_ ;
	wire _w27078_ ;
	wire _w27077_ ;
	wire _w27076_ ;
	wire _w27075_ ;
	wire _w27074_ ;
	wire _w27073_ ;
	wire _w27072_ ;
	wire _w27071_ ;
	wire _w27070_ ;
	wire _w27069_ ;
	wire _w27068_ ;
	wire _w27067_ ;
	wire _w27066_ ;
	wire _w27065_ ;
	wire _w27064_ ;
	wire _w27063_ ;
	wire _w27062_ ;
	wire _w27061_ ;
	wire _w27060_ ;
	wire _w27059_ ;
	wire _w27058_ ;
	wire _w27057_ ;
	wire _w27056_ ;
	wire _w27055_ ;
	wire _w27054_ ;
	wire _w27053_ ;
	wire _w27052_ ;
	wire _w27051_ ;
	wire _w27050_ ;
	wire _w27049_ ;
	wire _w27048_ ;
	wire _w27047_ ;
	wire _w27046_ ;
	wire _w27045_ ;
	wire _w27044_ ;
	wire _w27043_ ;
	wire _w27042_ ;
	wire _w27041_ ;
	wire _w27040_ ;
	wire _w27039_ ;
	wire _w27038_ ;
	wire _w27037_ ;
	wire _w27036_ ;
	wire _w27035_ ;
	wire _w27034_ ;
	wire _w27033_ ;
	wire _w27032_ ;
	wire _w27031_ ;
	wire _w27030_ ;
	wire _w27029_ ;
	wire _w27028_ ;
	wire _w27027_ ;
	wire _w27026_ ;
	wire _w27025_ ;
	wire _w27024_ ;
	wire _w27023_ ;
	wire _w27022_ ;
	wire _w27021_ ;
	wire _w27020_ ;
	wire _w27019_ ;
	wire _w27018_ ;
	wire _w27017_ ;
	wire _w27016_ ;
	wire _w27015_ ;
	wire _w27014_ ;
	wire _w27013_ ;
	wire _w27012_ ;
	wire _w27011_ ;
	wire _w27010_ ;
	wire _w27009_ ;
	wire _w27008_ ;
	wire _w27007_ ;
	wire _w27006_ ;
	wire _w27005_ ;
	wire _w27004_ ;
	wire _w27003_ ;
	wire _w27002_ ;
	wire _w27001_ ;
	wire _w27000_ ;
	wire _w26999_ ;
	wire _w26998_ ;
	wire _w26997_ ;
	wire _w26996_ ;
	wire _w26995_ ;
	wire _w26994_ ;
	wire _w26993_ ;
	wire _w26992_ ;
	wire _w26991_ ;
	wire _w26990_ ;
	wire _w26989_ ;
	wire _w26988_ ;
	wire _w26987_ ;
	wire _w26986_ ;
	wire _w26985_ ;
	wire _w26984_ ;
	wire _w26983_ ;
	wire _w26982_ ;
	wire _w26981_ ;
	wire _w26980_ ;
	wire _w26979_ ;
	wire _w26978_ ;
	wire _w26977_ ;
	wire _w26976_ ;
	wire _w26975_ ;
	wire _w26974_ ;
	wire _w26973_ ;
	wire _w26972_ ;
	wire _w26971_ ;
	wire _w26970_ ;
	wire _w26969_ ;
	wire _w26968_ ;
	wire _w26967_ ;
	wire _w26966_ ;
	wire _w26965_ ;
	wire _w26964_ ;
	wire _w26963_ ;
	wire _w26962_ ;
	wire _w26961_ ;
	wire _w26960_ ;
	wire _w26959_ ;
	wire _w26958_ ;
	wire _w26957_ ;
	wire _w26956_ ;
	wire _w26955_ ;
	wire _w26954_ ;
	wire _w26953_ ;
	wire _w26952_ ;
	wire _w26951_ ;
	wire _w26950_ ;
	wire _w26949_ ;
	wire _w26948_ ;
	wire _w26947_ ;
	wire _w26946_ ;
	wire _w26945_ ;
	wire _w26944_ ;
	wire _w26943_ ;
	wire _w26942_ ;
	wire _w26941_ ;
	wire _w26940_ ;
	wire _w26939_ ;
	wire _w26938_ ;
	wire _w26937_ ;
	wire _w26936_ ;
	wire _w26935_ ;
	wire _w26934_ ;
	wire _w26933_ ;
	wire _w26932_ ;
	wire _w26931_ ;
	wire _w26930_ ;
	wire _w26929_ ;
	wire _w26928_ ;
	wire _w26927_ ;
	wire _w26926_ ;
	wire _w26925_ ;
	wire _w26924_ ;
	wire _w26923_ ;
	wire _w26922_ ;
	wire _w26921_ ;
	wire _w26920_ ;
	wire _w26919_ ;
	wire _w26918_ ;
	wire _w26917_ ;
	wire _w26916_ ;
	wire _w26915_ ;
	wire _w26914_ ;
	wire _w26913_ ;
	wire _w26912_ ;
	wire _w26911_ ;
	wire _w26910_ ;
	wire _w26909_ ;
	wire _w26908_ ;
	wire _w26907_ ;
	wire _w26906_ ;
	wire _w26905_ ;
	wire _w26904_ ;
	wire _w26903_ ;
	wire _w26902_ ;
	wire _w26901_ ;
	wire _w26900_ ;
	wire _w26899_ ;
	wire _w26898_ ;
	wire _w26897_ ;
	wire _w26896_ ;
	wire _w26895_ ;
	wire _w26894_ ;
	wire _w26893_ ;
	wire _w26892_ ;
	wire _w26891_ ;
	wire _w26890_ ;
	wire _w26889_ ;
	wire _w26888_ ;
	wire _w26887_ ;
	wire _w26886_ ;
	wire _w26885_ ;
	wire _w26884_ ;
	wire _w26883_ ;
	wire _w26882_ ;
	wire _w26881_ ;
	wire _w26880_ ;
	wire _w26879_ ;
	wire _w26878_ ;
	wire _w26877_ ;
	wire _w26876_ ;
	wire _w26875_ ;
	wire _w26874_ ;
	wire _w26873_ ;
	wire _w26872_ ;
	wire _w26871_ ;
	wire _w26870_ ;
	wire _w26869_ ;
	wire _w26868_ ;
	wire _w26867_ ;
	wire _w26866_ ;
	wire _w26865_ ;
	wire _w26864_ ;
	wire _w26863_ ;
	wire _w26862_ ;
	wire _w26861_ ;
	wire _w26860_ ;
	wire _w26859_ ;
	wire _w26858_ ;
	wire _w26857_ ;
	wire _w26856_ ;
	wire _w26855_ ;
	wire _w26854_ ;
	wire _w26853_ ;
	wire _w26852_ ;
	wire _w26851_ ;
	wire _w26850_ ;
	wire _w26849_ ;
	wire _w26848_ ;
	wire _w26847_ ;
	wire _w26846_ ;
	wire _w26845_ ;
	wire _w26844_ ;
	wire _w26843_ ;
	wire _w26842_ ;
	wire _w26841_ ;
	wire _w26840_ ;
	wire _w26839_ ;
	wire _w26838_ ;
	wire _w26837_ ;
	wire _w26836_ ;
	wire _w26835_ ;
	wire _w26834_ ;
	wire _w26833_ ;
	wire _w26832_ ;
	wire _w26831_ ;
	wire _w26830_ ;
	wire _w26829_ ;
	wire _w26828_ ;
	wire _w26827_ ;
	wire _w26826_ ;
	wire _w26825_ ;
	wire _w26824_ ;
	wire _w26823_ ;
	wire _w26822_ ;
	wire _w26821_ ;
	wire _w26820_ ;
	wire _w26819_ ;
	wire _w26818_ ;
	wire _w26817_ ;
	wire _w26816_ ;
	wire _w26815_ ;
	wire _w26814_ ;
	wire _w26813_ ;
	wire _w26812_ ;
	wire _w26811_ ;
	wire _w26810_ ;
	wire _w26809_ ;
	wire _w26808_ ;
	wire _w26807_ ;
	wire _w26806_ ;
	wire _w26805_ ;
	wire _w26804_ ;
	wire _w26803_ ;
	wire _w26802_ ;
	wire _w26801_ ;
	wire _w26800_ ;
	wire _w26799_ ;
	wire _w26798_ ;
	wire _w26797_ ;
	wire _w26796_ ;
	wire _w26795_ ;
	wire _w26794_ ;
	wire _w26793_ ;
	wire _w26792_ ;
	wire _w26791_ ;
	wire _w26790_ ;
	wire _w26789_ ;
	wire _w26788_ ;
	wire _w26787_ ;
	wire _w26786_ ;
	wire _w26785_ ;
	wire _w26784_ ;
	wire _w26783_ ;
	wire _w26782_ ;
	wire _w26781_ ;
	wire _w26780_ ;
	wire _w26779_ ;
	wire _w26778_ ;
	wire _w26777_ ;
	wire _w26776_ ;
	wire _w26775_ ;
	wire _w26774_ ;
	wire _w26773_ ;
	wire _w26772_ ;
	wire _w26771_ ;
	wire _w26770_ ;
	wire _w26769_ ;
	wire _w26768_ ;
	wire _w26767_ ;
	wire _w26766_ ;
	wire _w26765_ ;
	wire _w26764_ ;
	wire _w26763_ ;
	wire _w26762_ ;
	wire _w26761_ ;
	wire _w26760_ ;
	wire _w26759_ ;
	wire _w26758_ ;
	wire _w26757_ ;
	wire _w26756_ ;
	wire _w26755_ ;
	wire _w26754_ ;
	wire _w26753_ ;
	wire _w26752_ ;
	wire _w26751_ ;
	wire _w26750_ ;
	wire _w26749_ ;
	wire _w26748_ ;
	wire _w26747_ ;
	wire _w26746_ ;
	wire _w26745_ ;
	wire _w26744_ ;
	wire _w26743_ ;
	wire _w26742_ ;
	wire _w26741_ ;
	wire _w26740_ ;
	wire _w26739_ ;
	wire _w26738_ ;
	wire _w26737_ ;
	wire _w26736_ ;
	wire _w26735_ ;
	wire _w26734_ ;
	wire _w26733_ ;
	wire _w26732_ ;
	wire _w26731_ ;
	wire _w26730_ ;
	wire _w26729_ ;
	wire _w26728_ ;
	wire _w26727_ ;
	wire _w26726_ ;
	wire _w26725_ ;
	wire _w26724_ ;
	wire _w26723_ ;
	wire _w26722_ ;
	wire _w26721_ ;
	wire _w26720_ ;
	wire _w26719_ ;
	wire _w26718_ ;
	wire _w26717_ ;
	wire _w26716_ ;
	wire _w26715_ ;
	wire _w26714_ ;
	wire _w26713_ ;
	wire _w26712_ ;
	wire _w26711_ ;
	wire _w26710_ ;
	wire _w26709_ ;
	wire _w26708_ ;
	wire _w26707_ ;
	wire _w26706_ ;
	wire _w26705_ ;
	wire _w26704_ ;
	wire _w26703_ ;
	wire _w26702_ ;
	wire _w26701_ ;
	wire _w26700_ ;
	wire _w26699_ ;
	wire _w26698_ ;
	wire _w26697_ ;
	wire _w26696_ ;
	wire _w26695_ ;
	wire _w26694_ ;
	wire _w26693_ ;
	wire _w26692_ ;
	wire _w26691_ ;
	wire _w26690_ ;
	wire _w26689_ ;
	wire _w26688_ ;
	wire _w26687_ ;
	wire _w26686_ ;
	wire _w26685_ ;
	wire _w26684_ ;
	wire _w26683_ ;
	wire _w26682_ ;
	wire _w26681_ ;
	wire _w26680_ ;
	wire _w26679_ ;
	wire _w26678_ ;
	wire _w26677_ ;
	wire _w26676_ ;
	wire _w26675_ ;
	wire _w26674_ ;
	wire _w26673_ ;
	wire _w26672_ ;
	wire _w26671_ ;
	wire _w26670_ ;
	wire _w26669_ ;
	wire _w26668_ ;
	wire _w26667_ ;
	wire _w26666_ ;
	wire _w26665_ ;
	wire _w26664_ ;
	wire _w26663_ ;
	wire _w26662_ ;
	wire _w26661_ ;
	wire _w26660_ ;
	wire _w26659_ ;
	wire _w26658_ ;
	wire _w26657_ ;
	wire _w26656_ ;
	wire _w26655_ ;
	wire _w26654_ ;
	wire _w26653_ ;
	wire _w26652_ ;
	wire _w26651_ ;
	wire _w26650_ ;
	wire _w26649_ ;
	wire _w26648_ ;
	wire _w26647_ ;
	wire _w26646_ ;
	wire _w26645_ ;
	wire _w26644_ ;
	wire _w26643_ ;
	wire _w26642_ ;
	wire _w26641_ ;
	wire _w26640_ ;
	wire _w26639_ ;
	wire _w26638_ ;
	wire _w26637_ ;
	wire _w26636_ ;
	wire _w26635_ ;
	wire _w26634_ ;
	wire _w26633_ ;
	wire _w26632_ ;
	wire _w26631_ ;
	wire _w26630_ ;
	wire _w26629_ ;
	wire _w26628_ ;
	wire _w26627_ ;
	wire _w26626_ ;
	wire _w26625_ ;
	wire _w26624_ ;
	wire _w26623_ ;
	wire _w26622_ ;
	wire _w26621_ ;
	wire _w26620_ ;
	wire _w26619_ ;
	wire _w26618_ ;
	wire _w26617_ ;
	wire _w26616_ ;
	wire _w26615_ ;
	wire _w26614_ ;
	wire _w26613_ ;
	wire _w26612_ ;
	wire _w26611_ ;
	wire _w26610_ ;
	wire _w26609_ ;
	wire _w26608_ ;
	wire _w26607_ ;
	wire _w26606_ ;
	wire _w26605_ ;
	wire _w26604_ ;
	wire _w26603_ ;
	wire _w26602_ ;
	wire _w26601_ ;
	wire _w26600_ ;
	wire _w26599_ ;
	wire _w26598_ ;
	wire _w26597_ ;
	wire _w26596_ ;
	wire _w26595_ ;
	wire _w26594_ ;
	wire _w26593_ ;
	wire _w26592_ ;
	wire _w26591_ ;
	wire _w26590_ ;
	wire _w26589_ ;
	wire _w26588_ ;
	wire _w26587_ ;
	wire _w26586_ ;
	wire _w26585_ ;
	wire _w26584_ ;
	wire _w26583_ ;
	wire _w26582_ ;
	wire _w26581_ ;
	wire _w26580_ ;
	wire _w26579_ ;
	wire _w26578_ ;
	wire _w26577_ ;
	wire _w26576_ ;
	wire _w26575_ ;
	wire _w26574_ ;
	wire _w26573_ ;
	wire _w26572_ ;
	wire _w26571_ ;
	wire _w26570_ ;
	wire _w26569_ ;
	wire _w26568_ ;
	wire _w26567_ ;
	wire _w26566_ ;
	wire _w26565_ ;
	wire _w26564_ ;
	wire _w26563_ ;
	wire _w26562_ ;
	wire _w26561_ ;
	wire _w26560_ ;
	wire _w26559_ ;
	wire _w26558_ ;
	wire _w26557_ ;
	wire _w26556_ ;
	wire _w26555_ ;
	wire _w26554_ ;
	wire _w26553_ ;
	wire _w26552_ ;
	wire _w26551_ ;
	wire _w26550_ ;
	wire _w26549_ ;
	wire _w26548_ ;
	wire _w26547_ ;
	wire _w26546_ ;
	wire _w26545_ ;
	wire _w26544_ ;
	wire _w26543_ ;
	wire _w26542_ ;
	wire _w26541_ ;
	wire _w26540_ ;
	wire _w26539_ ;
	wire _w26538_ ;
	wire _w26537_ ;
	wire _w26536_ ;
	wire _w26535_ ;
	wire _w26534_ ;
	wire _w26533_ ;
	wire _w26532_ ;
	wire _w26531_ ;
	wire _w26530_ ;
	wire _w26529_ ;
	wire _w26528_ ;
	wire _w26527_ ;
	wire _w26526_ ;
	wire _w26525_ ;
	wire _w26524_ ;
	wire _w26523_ ;
	wire _w26522_ ;
	wire _w26521_ ;
	wire _w26520_ ;
	wire _w26519_ ;
	wire _w26518_ ;
	wire _w26517_ ;
	wire _w26516_ ;
	wire _w26515_ ;
	wire _w26514_ ;
	wire _w26513_ ;
	wire _w26512_ ;
	wire _w26511_ ;
	wire _w26510_ ;
	wire _w26509_ ;
	wire _w26508_ ;
	wire _w26507_ ;
	wire _w26506_ ;
	wire _w26505_ ;
	wire _w26504_ ;
	wire _w26503_ ;
	wire _w26502_ ;
	wire _w26501_ ;
	wire _w26500_ ;
	wire _w26499_ ;
	wire _w26498_ ;
	wire _w26497_ ;
	wire _w26496_ ;
	wire _w26495_ ;
	wire _w26494_ ;
	wire _w26493_ ;
	wire _w26492_ ;
	wire _w26491_ ;
	wire _w26490_ ;
	wire _w26489_ ;
	wire _w26488_ ;
	wire _w26487_ ;
	wire _w26486_ ;
	wire _w26485_ ;
	wire _w26484_ ;
	wire _w26483_ ;
	wire _w26482_ ;
	wire _w26481_ ;
	wire _w26480_ ;
	wire _w26479_ ;
	wire _w26478_ ;
	wire _w26477_ ;
	wire _w26476_ ;
	wire _w26475_ ;
	wire _w26474_ ;
	wire _w26473_ ;
	wire _w26472_ ;
	wire _w26471_ ;
	wire _w26470_ ;
	wire _w26469_ ;
	wire _w26468_ ;
	wire _w26467_ ;
	wire _w26466_ ;
	wire _w26465_ ;
	wire _w26464_ ;
	wire _w26463_ ;
	wire _w26462_ ;
	wire _w26461_ ;
	wire _w26460_ ;
	wire _w26459_ ;
	wire _w26458_ ;
	wire _w26457_ ;
	wire _w26456_ ;
	wire _w26455_ ;
	wire _w26454_ ;
	wire _w26453_ ;
	wire _w26452_ ;
	wire _w26451_ ;
	wire _w26450_ ;
	wire _w26449_ ;
	wire _w26448_ ;
	wire _w26447_ ;
	wire _w26446_ ;
	wire _w26445_ ;
	wire _w26444_ ;
	wire _w26443_ ;
	wire _w26442_ ;
	wire _w26441_ ;
	wire _w26440_ ;
	wire _w26439_ ;
	wire _w26438_ ;
	wire _w26437_ ;
	wire _w26436_ ;
	wire _w26435_ ;
	wire _w26434_ ;
	wire _w26433_ ;
	wire _w26432_ ;
	wire _w26431_ ;
	wire _w26430_ ;
	wire _w26429_ ;
	wire _w26428_ ;
	wire _w26427_ ;
	wire _w26426_ ;
	wire _w26425_ ;
	wire _w26424_ ;
	wire _w26423_ ;
	wire _w26422_ ;
	wire _w26421_ ;
	wire _w26420_ ;
	wire _w26419_ ;
	wire _w26418_ ;
	wire _w26417_ ;
	wire _w26416_ ;
	wire _w26415_ ;
	wire _w26414_ ;
	wire _w26413_ ;
	wire _w26412_ ;
	wire _w26411_ ;
	wire _w26410_ ;
	wire _w26409_ ;
	wire _w26408_ ;
	wire _w26407_ ;
	wire _w26406_ ;
	wire _w26405_ ;
	wire _w26404_ ;
	wire _w26403_ ;
	wire _w26402_ ;
	wire _w26401_ ;
	wire _w26400_ ;
	wire _w26399_ ;
	wire _w26398_ ;
	wire _w26397_ ;
	wire _w26396_ ;
	wire _w26395_ ;
	wire _w26394_ ;
	wire _w26393_ ;
	wire _w26392_ ;
	wire _w26391_ ;
	wire _w26390_ ;
	wire _w26389_ ;
	wire _w26388_ ;
	wire _w26387_ ;
	wire _w26386_ ;
	wire _w26385_ ;
	wire _w26384_ ;
	wire _w26383_ ;
	wire _w26382_ ;
	wire _w26381_ ;
	wire _w26380_ ;
	wire _w26379_ ;
	wire _w26378_ ;
	wire _w26377_ ;
	wire _w26376_ ;
	wire _w26375_ ;
	wire _w26374_ ;
	wire _w26373_ ;
	wire _w26372_ ;
	wire _w26371_ ;
	wire _w26370_ ;
	wire _w26369_ ;
	wire _w26368_ ;
	wire _w26367_ ;
	wire _w26366_ ;
	wire _w26365_ ;
	wire _w26364_ ;
	wire _w26363_ ;
	wire _w26362_ ;
	wire _w26361_ ;
	wire _w26360_ ;
	wire _w26359_ ;
	wire _w26358_ ;
	wire _w26357_ ;
	wire _w26356_ ;
	wire _w26355_ ;
	wire _w26354_ ;
	wire _w26353_ ;
	wire _w26352_ ;
	wire _w26351_ ;
	wire _w26350_ ;
	wire _w26349_ ;
	wire _w26348_ ;
	wire _w26347_ ;
	wire _w26346_ ;
	wire _w26345_ ;
	wire _w26344_ ;
	wire _w26343_ ;
	wire _w26342_ ;
	wire _w26341_ ;
	wire _w26340_ ;
	wire _w26339_ ;
	wire _w26338_ ;
	wire _w26337_ ;
	wire _w26336_ ;
	wire _w26335_ ;
	wire _w26334_ ;
	wire _w26333_ ;
	wire _w26332_ ;
	wire _w26331_ ;
	wire _w26330_ ;
	wire _w26329_ ;
	wire _w26328_ ;
	wire _w26327_ ;
	wire _w26326_ ;
	wire _w26325_ ;
	wire _w26324_ ;
	wire _w26323_ ;
	wire _w26322_ ;
	wire _w26321_ ;
	wire _w26320_ ;
	wire _w26319_ ;
	wire _w26318_ ;
	wire _w26317_ ;
	wire _w26316_ ;
	wire _w26315_ ;
	wire _w26314_ ;
	wire _w26313_ ;
	wire _w26312_ ;
	wire _w26311_ ;
	wire _w26310_ ;
	wire _w26309_ ;
	wire _w26308_ ;
	wire _w26307_ ;
	wire _w26306_ ;
	wire _w26305_ ;
	wire _w26304_ ;
	wire _w26303_ ;
	wire _w26302_ ;
	wire _w26301_ ;
	wire _w26300_ ;
	wire _w26299_ ;
	wire _w26298_ ;
	wire _w26297_ ;
	wire _w26296_ ;
	wire _w26295_ ;
	wire _w26294_ ;
	wire _w26293_ ;
	wire _w26292_ ;
	wire _w26291_ ;
	wire _w26290_ ;
	wire _w26289_ ;
	wire _w26288_ ;
	wire _w26287_ ;
	wire _w26286_ ;
	wire _w26285_ ;
	wire _w26284_ ;
	wire _w26283_ ;
	wire _w26282_ ;
	wire _w26281_ ;
	wire _w26280_ ;
	wire _w26279_ ;
	wire _w26278_ ;
	wire _w26277_ ;
	wire _w26276_ ;
	wire _w26275_ ;
	wire _w26274_ ;
	wire _w26273_ ;
	wire _w26272_ ;
	wire _w26271_ ;
	wire _w26270_ ;
	wire _w26269_ ;
	wire _w26268_ ;
	wire _w26267_ ;
	wire _w26266_ ;
	wire _w26265_ ;
	wire _w26264_ ;
	wire _w26263_ ;
	wire _w26262_ ;
	wire _w26261_ ;
	wire _w26260_ ;
	wire _w26259_ ;
	wire _w26258_ ;
	wire _w26257_ ;
	wire _w26256_ ;
	wire _w26255_ ;
	wire _w26254_ ;
	wire _w26253_ ;
	wire _w26252_ ;
	wire _w26251_ ;
	wire _w26250_ ;
	wire _w26249_ ;
	wire _w26248_ ;
	wire _w26247_ ;
	wire _w26246_ ;
	wire _w26245_ ;
	wire _w26244_ ;
	wire _w26243_ ;
	wire _w26242_ ;
	wire _w26241_ ;
	wire _w26240_ ;
	wire _w26239_ ;
	wire _w26238_ ;
	wire _w26237_ ;
	wire _w26236_ ;
	wire _w26235_ ;
	wire _w26234_ ;
	wire _w26233_ ;
	wire _w26232_ ;
	wire _w26231_ ;
	wire _w26230_ ;
	wire _w26229_ ;
	wire _w26228_ ;
	wire _w26227_ ;
	wire _w26226_ ;
	wire _w26225_ ;
	wire _w26224_ ;
	wire _w26223_ ;
	wire _w26222_ ;
	wire _w26221_ ;
	wire _w26220_ ;
	wire _w26219_ ;
	wire _w26218_ ;
	wire _w26217_ ;
	wire _w26216_ ;
	wire _w26215_ ;
	wire _w26214_ ;
	wire _w26213_ ;
	wire _w26212_ ;
	wire _w26211_ ;
	wire _w26210_ ;
	wire _w26209_ ;
	wire _w26208_ ;
	wire _w26207_ ;
	wire _w26206_ ;
	wire _w26205_ ;
	wire _w26204_ ;
	wire _w26203_ ;
	wire _w26202_ ;
	wire _w26201_ ;
	wire _w26200_ ;
	wire _w26199_ ;
	wire _w26198_ ;
	wire _w26197_ ;
	wire _w26196_ ;
	wire _w26195_ ;
	wire _w26194_ ;
	wire _w26193_ ;
	wire _w26192_ ;
	wire _w26191_ ;
	wire _w26190_ ;
	wire _w26189_ ;
	wire _w26188_ ;
	wire _w26187_ ;
	wire _w26186_ ;
	wire _w26185_ ;
	wire _w26184_ ;
	wire _w26183_ ;
	wire _w26182_ ;
	wire _w26181_ ;
	wire _w26180_ ;
	wire _w26179_ ;
	wire _w26178_ ;
	wire _w26177_ ;
	wire _w26176_ ;
	wire _w26175_ ;
	wire _w26174_ ;
	wire _w26173_ ;
	wire _w26172_ ;
	wire _w26171_ ;
	wire _w26170_ ;
	wire _w26169_ ;
	wire _w26168_ ;
	wire _w26167_ ;
	wire _w26166_ ;
	wire _w26165_ ;
	wire _w26164_ ;
	wire _w26163_ ;
	wire _w26162_ ;
	wire _w26161_ ;
	wire _w26160_ ;
	wire _w26159_ ;
	wire _w26158_ ;
	wire _w26157_ ;
	wire _w26156_ ;
	wire _w26155_ ;
	wire _w26154_ ;
	wire _w26153_ ;
	wire _w26152_ ;
	wire _w26151_ ;
	wire _w26150_ ;
	wire _w26149_ ;
	wire _w26148_ ;
	wire _w26147_ ;
	wire _w26146_ ;
	wire _w26145_ ;
	wire _w26144_ ;
	wire _w26143_ ;
	wire _w26142_ ;
	wire _w26141_ ;
	wire _w26140_ ;
	wire _w26139_ ;
	wire _w26138_ ;
	wire _w26137_ ;
	wire _w26136_ ;
	wire _w26135_ ;
	wire _w26134_ ;
	wire _w26133_ ;
	wire _w26132_ ;
	wire _w26131_ ;
	wire _w26130_ ;
	wire _w26129_ ;
	wire _w26128_ ;
	wire _w26127_ ;
	wire _w26126_ ;
	wire _w26125_ ;
	wire _w26124_ ;
	wire _w26123_ ;
	wire _w26122_ ;
	wire _w26121_ ;
	wire _w26120_ ;
	wire _w26119_ ;
	wire _w26118_ ;
	wire _w26117_ ;
	wire _w26116_ ;
	wire _w26115_ ;
	wire _w26114_ ;
	wire _w26113_ ;
	wire _w26112_ ;
	wire _w26111_ ;
	wire _w26110_ ;
	wire _w26109_ ;
	wire _w26108_ ;
	wire _w26107_ ;
	wire _w26106_ ;
	wire _w26105_ ;
	wire _w26104_ ;
	wire _w26103_ ;
	wire _w26102_ ;
	wire _w26101_ ;
	wire _w26100_ ;
	wire _w26099_ ;
	wire _w26098_ ;
	wire _w26097_ ;
	wire _w26096_ ;
	wire _w26095_ ;
	wire _w26094_ ;
	wire _w26093_ ;
	wire _w26092_ ;
	wire _w26091_ ;
	wire _w26090_ ;
	wire _w26089_ ;
	wire _w26088_ ;
	wire _w26087_ ;
	wire _w26086_ ;
	wire _w26085_ ;
	wire _w26084_ ;
	wire _w26083_ ;
	wire _w26082_ ;
	wire _w26081_ ;
	wire _w26080_ ;
	wire _w26079_ ;
	wire _w26078_ ;
	wire _w26077_ ;
	wire _w26076_ ;
	wire _w26075_ ;
	wire _w26074_ ;
	wire _w26073_ ;
	wire _w26072_ ;
	wire _w26071_ ;
	wire _w26070_ ;
	wire _w26069_ ;
	wire _w26068_ ;
	wire _w26067_ ;
	wire _w26066_ ;
	wire _w26065_ ;
	wire _w26064_ ;
	wire _w26063_ ;
	wire _w26062_ ;
	wire _w26061_ ;
	wire _w26060_ ;
	wire _w26059_ ;
	wire _w26058_ ;
	wire _w26057_ ;
	wire _w26056_ ;
	wire _w26055_ ;
	wire _w26054_ ;
	wire _w26053_ ;
	wire _w26052_ ;
	wire _w26051_ ;
	wire _w26050_ ;
	wire _w26049_ ;
	wire _w26048_ ;
	wire _w26047_ ;
	wire _w26046_ ;
	wire _w26045_ ;
	wire _w26044_ ;
	wire _w26043_ ;
	wire _w26042_ ;
	wire _w26041_ ;
	wire _w26040_ ;
	wire _w26039_ ;
	wire _w26038_ ;
	wire _w26037_ ;
	wire _w26036_ ;
	wire _w26035_ ;
	wire _w26034_ ;
	wire _w26033_ ;
	wire _w26032_ ;
	wire _w26031_ ;
	wire _w26030_ ;
	wire _w26029_ ;
	wire _w26028_ ;
	wire _w26027_ ;
	wire _w26026_ ;
	wire _w26025_ ;
	wire _w26024_ ;
	wire _w26023_ ;
	wire _w26022_ ;
	wire _w26021_ ;
	wire _w26020_ ;
	wire _w26019_ ;
	wire _w26018_ ;
	wire _w26017_ ;
	wire _w26016_ ;
	wire _w26015_ ;
	wire _w26014_ ;
	wire _w26013_ ;
	wire _w26012_ ;
	wire _w26011_ ;
	wire _w26010_ ;
	wire _w26009_ ;
	wire _w26008_ ;
	wire _w26007_ ;
	wire _w26006_ ;
	wire _w26005_ ;
	wire _w26004_ ;
	wire _w26003_ ;
	wire _w26002_ ;
	wire _w26001_ ;
	wire _w26000_ ;
	wire _w25999_ ;
	wire _w25998_ ;
	wire _w25997_ ;
	wire _w25996_ ;
	wire _w25995_ ;
	wire _w25994_ ;
	wire _w25993_ ;
	wire _w25992_ ;
	wire _w25991_ ;
	wire _w25990_ ;
	wire _w25989_ ;
	wire _w25988_ ;
	wire _w25987_ ;
	wire _w25986_ ;
	wire _w25985_ ;
	wire _w25984_ ;
	wire _w25983_ ;
	wire _w25982_ ;
	wire _w25981_ ;
	wire _w25980_ ;
	wire _w25979_ ;
	wire _w25978_ ;
	wire _w25977_ ;
	wire _w25976_ ;
	wire _w25975_ ;
	wire _w25974_ ;
	wire _w25973_ ;
	wire _w25972_ ;
	wire _w25971_ ;
	wire _w25970_ ;
	wire _w25969_ ;
	wire _w25968_ ;
	wire _w25967_ ;
	wire _w25966_ ;
	wire _w25965_ ;
	wire _w25964_ ;
	wire _w25963_ ;
	wire _w25962_ ;
	wire _w25961_ ;
	wire _w25960_ ;
	wire _w25959_ ;
	wire _w25958_ ;
	wire _w25957_ ;
	wire _w25956_ ;
	wire _w25955_ ;
	wire _w25954_ ;
	wire _w25953_ ;
	wire _w25952_ ;
	wire _w25951_ ;
	wire _w25950_ ;
	wire _w25949_ ;
	wire _w25948_ ;
	wire _w25947_ ;
	wire _w25946_ ;
	wire _w25945_ ;
	wire _w25944_ ;
	wire _w25943_ ;
	wire _w25942_ ;
	wire _w25941_ ;
	wire _w25940_ ;
	wire _w25939_ ;
	wire _w25938_ ;
	wire _w25937_ ;
	wire _w25936_ ;
	wire _w25935_ ;
	wire _w25934_ ;
	wire _w25933_ ;
	wire _w25932_ ;
	wire _w25931_ ;
	wire _w25930_ ;
	wire _w25929_ ;
	wire _w25928_ ;
	wire _w25927_ ;
	wire _w25926_ ;
	wire _w25925_ ;
	wire _w25924_ ;
	wire _w25923_ ;
	wire _w25922_ ;
	wire _w25921_ ;
	wire _w25920_ ;
	wire _w25919_ ;
	wire _w25918_ ;
	wire _w25917_ ;
	wire _w25916_ ;
	wire _w25915_ ;
	wire _w25914_ ;
	wire _w25913_ ;
	wire _w25912_ ;
	wire _w25911_ ;
	wire _w25910_ ;
	wire _w25909_ ;
	wire _w25908_ ;
	wire _w25907_ ;
	wire _w25906_ ;
	wire _w25905_ ;
	wire _w25904_ ;
	wire _w25903_ ;
	wire _w25902_ ;
	wire _w25901_ ;
	wire _w25900_ ;
	wire _w25899_ ;
	wire _w25898_ ;
	wire _w25897_ ;
	wire _w25896_ ;
	wire _w25895_ ;
	wire _w25894_ ;
	wire _w25893_ ;
	wire _w25892_ ;
	wire _w25891_ ;
	wire _w25890_ ;
	wire _w25889_ ;
	wire _w25888_ ;
	wire _w25887_ ;
	wire _w25886_ ;
	wire _w25885_ ;
	wire _w25884_ ;
	wire _w25883_ ;
	wire _w25882_ ;
	wire _w25881_ ;
	wire _w25880_ ;
	wire _w25879_ ;
	wire _w25878_ ;
	wire _w25877_ ;
	wire _w25876_ ;
	wire _w25875_ ;
	wire _w25874_ ;
	wire _w25873_ ;
	wire _w25872_ ;
	wire _w25871_ ;
	wire _w25870_ ;
	wire _w25869_ ;
	wire _w25868_ ;
	wire _w25867_ ;
	wire _w25866_ ;
	wire _w25865_ ;
	wire _w25864_ ;
	wire _w25863_ ;
	wire _w25862_ ;
	wire _w25861_ ;
	wire _w25860_ ;
	wire _w25859_ ;
	wire _w25858_ ;
	wire _w25857_ ;
	wire _w25856_ ;
	wire _w25855_ ;
	wire _w25854_ ;
	wire _w25853_ ;
	wire _w25852_ ;
	wire _w25851_ ;
	wire _w25850_ ;
	wire _w25849_ ;
	wire _w25848_ ;
	wire _w25847_ ;
	wire _w25846_ ;
	wire _w25845_ ;
	wire _w25844_ ;
	wire _w25843_ ;
	wire _w25842_ ;
	wire _w25841_ ;
	wire _w25840_ ;
	wire _w25839_ ;
	wire _w25838_ ;
	wire _w25837_ ;
	wire _w25836_ ;
	wire _w25835_ ;
	wire _w25834_ ;
	wire _w25833_ ;
	wire _w25832_ ;
	wire _w25831_ ;
	wire _w25830_ ;
	wire _w25829_ ;
	wire _w25828_ ;
	wire _w25827_ ;
	wire _w25826_ ;
	wire _w25825_ ;
	wire _w25824_ ;
	wire _w25823_ ;
	wire _w25822_ ;
	wire _w25821_ ;
	wire _w25820_ ;
	wire _w25819_ ;
	wire _w25818_ ;
	wire _w25817_ ;
	wire _w25816_ ;
	wire _w25815_ ;
	wire _w25814_ ;
	wire _w25813_ ;
	wire _w25812_ ;
	wire _w25811_ ;
	wire _w25810_ ;
	wire _w25809_ ;
	wire _w25808_ ;
	wire _w25807_ ;
	wire _w25806_ ;
	wire _w25805_ ;
	wire _w25804_ ;
	wire _w25803_ ;
	wire _w25802_ ;
	wire _w25801_ ;
	wire _w25800_ ;
	wire _w25799_ ;
	wire _w25798_ ;
	wire _w25797_ ;
	wire _w25796_ ;
	wire _w25795_ ;
	wire _w25794_ ;
	wire _w25793_ ;
	wire _w25792_ ;
	wire _w25791_ ;
	wire _w25790_ ;
	wire _w25789_ ;
	wire _w25788_ ;
	wire _w25787_ ;
	wire _w25786_ ;
	wire _w25785_ ;
	wire _w25784_ ;
	wire _w25783_ ;
	wire _w25782_ ;
	wire _w25781_ ;
	wire _w25780_ ;
	wire _w25779_ ;
	wire _w25778_ ;
	wire _w25777_ ;
	wire _w25776_ ;
	wire _w25775_ ;
	wire _w25774_ ;
	wire _w25773_ ;
	wire _w25772_ ;
	wire _w25771_ ;
	wire _w25770_ ;
	wire _w25769_ ;
	wire _w25768_ ;
	wire _w25767_ ;
	wire _w25766_ ;
	wire _w25765_ ;
	wire _w25764_ ;
	wire _w25763_ ;
	wire _w25762_ ;
	wire _w25761_ ;
	wire _w25760_ ;
	wire _w25759_ ;
	wire _w25758_ ;
	wire _w25757_ ;
	wire _w25756_ ;
	wire _w25755_ ;
	wire _w25754_ ;
	wire _w25753_ ;
	wire _w25752_ ;
	wire _w25751_ ;
	wire _w25750_ ;
	wire _w25749_ ;
	wire _w25748_ ;
	wire _w25747_ ;
	wire _w25746_ ;
	wire _w25745_ ;
	wire _w25744_ ;
	wire _w25743_ ;
	wire _w25742_ ;
	wire _w25741_ ;
	wire _w25740_ ;
	wire _w25739_ ;
	wire _w25738_ ;
	wire _w25737_ ;
	wire _w25736_ ;
	wire _w25735_ ;
	wire _w25734_ ;
	wire _w25733_ ;
	wire _w25732_ ;
	wire _w25731_ ;
	wire _w25730_ ;
	wire _w25729_ ;
	wire _w25728_ ;
	wire _w25727_ ;
	wire _w25726_ ;
	wire _w25725_ ;
	wire _w25724_ ;
	wire _w25723_ ;
	wire _w25722_ ;
	wire _w25721_ ;
	wire _w25720_ ;
	wire _w25719_ ;
	wire _w25718_ ;
	wire _w25717_ ;
	wire _w25716_ ;
	wire _w25715_ ;
	wire _w25714_ ;
	wire _w25713_ ;
	wire _w25712_ ;
	wire _w25711_ ;
	wire _w25710_ ;
	wire _w25709_ ;
	wire _w25708_ ;
	wire _w25707_ ;
	wire _w25706_ ;
	wire _w25705_ ;
	wire _w25704_ ;
	wire _w25703_ ;
	wire _w25702_ ;
	wire _w25701_ ;
	wire _w25700_ ;
	wire _w25699_ ;
	wire _w25698_ ;
	wire _w25697_ ;
	wire _w25696_ ;
	wire _w25695_ ;
	wire _w25694_ ;
	wire _w25693_ ;
	wire _w25692_ ;
	wire _w25691_ ;
	wire _w25690_ ;
	wire _w25689_ ;
	wire _w25688_ ;
	wire _w25687_ ;
	wire _w25686_ ;
	wire _w25685_ ;
	wire _w25684_ ;
	wire _w25683_ ;
	wire _w25682_ ;
	wire _w25681_ ;
	wire _w25680_ ;
	wire _w25679_ ;
	wire _w25678_ ;
	wire _w25677_ ;
	wire _w25676_ ;
	wire _w25675_ ;
	wire _w25674_ ;
	wire _w25673_ ;
	wire _w25672_ ;
	wire _w25671_ ;
	wire _w25670_ ;
	wire _w25669_ ;
	wire _w25668_ ;
	wire _w25667_ ;
	wire _w25666_ ;
	wire _w25665_ ;
	wire _w25664_ ;
	wire _w25663_ ;
	wire _w25662_ ;
	wire _w25661_ ;
	wire _w25660_ ;
	wire _w25659_ ;
	wire _w25658_ ;
	wire _w25657_ ;
	wire _w25656_ ;
	wire _w25655_ ;
	wire _w25654_ ;
	wire _w25653_ ;
	wire _w25652_ ;
	wire _w25651_ ;
	wire _w25650_ ;
	wire _w25649_ ;
	wire _w25648_ ;
	wire _w25647_ ;
	wire _w25646_ ;
	wire _w25645_ ;
	wire _w25644_ ;
	wire _w25643_ ;
	wire _w25642_ ;
	wire _w25641_ ;
	wire _w25640_ ;
	wire _w25639_ ;
	wire _w25638_ ;
	wire _w25637_ ;
	wire _w25636_ ;
	wire _w25635_ ;
	wire _w25634_ ;
	wire _w25633_ ;
	wire _w25632_ ;
	wire _w25631_ ;
	wire _w25630_ ;
	wire _w25629_ ;
	wire _w25628_ ;
	wire _w25627_ ;
	wire _w25626_ ;
	wire _w25625_ ;
	wire _w25624_ ;
	wire _w25623_ ;
	wire _w25622_ ;
	wire _w25621_ ;
	wire _w25620_ ;
	wire _w25619_ ;
	wire _w25618_ ;
	wire _w25617_ ;
	wire _w25616_ ;
	wire _w25615_ ;
	wire _w25614_ ;
	wire _w25613_ ;
	wire _w25612_ ;
	wire _w25611_ ;
	wire _w25610_ ;
	wire _w25609_ ;
	wire _w25608_ ;
	wire _w25607_ ;
	wire _w25606_ ;
	wire _w25605_ ;
	wire _w25604_ ;
	wire _w25603_ ;
	wire _w25602_ ;
	wire _w25601_ ;
	wire _w25600_ ;
	wire _w25599_ ;
	wire _w25598_ ;
	wire _w25597_ ;
	wire _w25596_ ;
	wire _w25595_ ;
	wire _w25594_ ;
	wire _w25593_ ;
	wire _w25592_ ;
	wire _w25591_ ;
	wire _w25590_ ;
	wire _w25589_ ;
	wire _w25588_ ;
	wire _w25587_ ;
	wire _w25586_ ;
	wire _w25585_ ;
	wire _w25584_ ;
	wire _w25583_ ;
	wire _w25582_ ;
	wire _w25581_ ;
	wire _w25580_ ;
	wire _w25579_ ;
	wire _w25578_ ;
	wire _w25577_ ;
	wire _w25576_ ;
	wire _w25575_ ;
	wire _w25574_ ;
	wire _w25573_ ;
	wire _w25572_ ;
	wire _w25571_ ;
	wire _w25570_ ;
	wire _w25569_ ;
	wire _w25568_ ;
	wire _w25567_ ;
	wire _w25566_ ;
	wire _w25565_ ;
	wire _w25564_ ;
	wire _w25563_ ;
	wire _w25562_ ;
	wire _w25561_ ;
	wire _w25560_ ;
	wire _w25559_ ;
	wire _w25558_ ;
	wire _w25557_ ;
	wire _w25556_ ;
	wire _w25555_ ;
	wire _w25554_ ;
	wire _w25553_ ;
	wire _w25552_ ;
	wire _w25551_ ;
	wire _w25550_ ;
	wire _w25549_ ;
	wire _w25548_ ;
	wire _w25547_ ;
	wire _w25546_ ;
	wire _w25545_ ;
	wire _w25544_ ;
	wire _w25543_ ;
	wire _w25542_ ;
	wire _w25541_ ;
	wire _w25540_ ;
	wire _w25539_ ;
	wire _w25538_ ;
	wire _w25537_ ;
	wire _w25536_ ;
	wire _w25535_ ;
	wire _w25534_ ;
	wire _w25533_ ;
	wire _w25532_ ;
	wire _w25531_ ;
	wire _w25530_ ;
	wire _w25529_ ;
	wire _w25528_ ;
	wire _w25527_ ;
	wire _w25526_ ;
	wire _w25525_ ;
	wire _w25524_ ;
	wire _w25523_ ;
	wire _w25522_ ;
	wire _w25521_ ;
	wire _w25520_ ;
	wire _w25519_ ;
	wire _w25518_ ;
	wire _w25517_ ;
	wire _w25516_ ;
	wire _w25515_ ;
	wire _w25514_ ;
	wire _w25513_ ;
	wire _w25512_ ;
	wire _w25511_ ;
	wire _w25510_ ;
	wire _w25509_ ;
	wire _w25508_ ;
	wire _w25507_ ;
	wire _w25506_ ;
	wire _w25505_ ;
	wire _w25504_ ;
	wire _w25503_ ;
	wire _w25502_ ;
	wire _w25501_ ;
	wire _w25500_ ;
	wire _w25499_ ;
	wire _w25498_ ;
	wire _w25497_ ;
	wire _w25496_ ;
	wire _w25495_ ;
	wire _w25494_ ;
	wire _w25493_ ;
	wire _w25492_ ;
	wire _w25491_ ;
	wire _w25490_ ;
	wire _w25489_ ;
	wire _w25488_ ;
	wire _w25487_ ;
	wire _w25486_ ;
	wire _w25485_ ;
	wire _w25484_ ;
	wire _w25483_ ;
	wire _w25482_ ;
	wire _w25481_ ;
	wire _w25480_ ;
	wire _w25479_ ;
	wire _w25478_ ;
	wire _w25477_ ;
	wire _w25476_ ;
	wire _w25475_ ;
	wire _w25474_ ;
	wire _w25473_ ;
	wire _w25472_ ;
	wire _w25471_ ;
	wire _w25470_ ;
	wire _w25469_ ;
	wire _w25468_ ;
	wire _w25467_ ;
	wire _w25466_ ;
	wire _w25465_ ;
	wire _w25464_ ;
	wire _w25463_ ;
	wire _w25462_ ;
	wire _w25461_ ;
	wire _w25460_ ;
	wire _w25459_ ;
	wire _w25458_ ;
	wire _w25457_ ;
	wire _w25456_ ;
	wire _w25455_ ;
	wire _w25454_ ;
	wire _w25453_ ;
	wire _w25452_ ;
	wire _w25451_ ;
	wire _w25450_ ;
	wire _w25449_ ;
	wire _w25448_ ;
	wire _w25447_ ;
	wire _w25446_ ;
	wire _w25445_ ;
	wire _w25444_ ;
	wire _w25443_ ;
	wire _w25442_ ;
	wire _w25441_ ;
	wire _w25440_ ;
	wire _w25439_ ;
	wire _w25438_ ;
	wire _w25437_ ;
	wire _w25436_ ;
	wire _w25435_ ;
	wire _w25434_ ;
	wire _w25433_ ;
	wire _w25432_ ;
	wire _w25431_ ;
	wire _w25430_ ;
	wire _w25429_ ;
	wire _w25428_ ;
	wire _w25427_ ;
	wire _w25426_ ;
	wire _w25425_ ;
	wire _w25424_ ;
	wire _w25423_ ;
	wire _w25422_ ;
	wire _w25421_ ;
	wire _w25420_ ;
	wire _w25419_ ;
	wire _w25418_ ;
	wire _w25417_ ;
	wire _w25416_ ;
	wire _w25415_ ;
	wire _w25414_ ;
	wire _w25413_ ;
	wire _w25412_ ;
	wire _w25411_ ;
	wire _w25410_ ;
	wire _w25409_ ;
	wire _w25408_ ;
	wire _w25407_ ;
	wire _w25406_ ;
	wire _w25405_ ;
	wire _w25404_ ;
	wire _w25403_ ;
	wire _w25402_ ;
	wire _w25401_ ;
	wire _w25400_ ;
	wire _w25399_ ;
	wire _w25398_ ;
	wire _w25397_ ;
	wire _w25396_ ;
	wire _w25395_ ;
	wire _w25394_ ;
	wire _w25393_ ;
	wire _w25392_ ;
	wire _w25391_ ;
	wire _w25390_ ;
	wire _w25389_ ;
	wire _w25388_ ;
	wire _w25387_ ;
	wire _w25386_ ;
	wire _w25385_ ;
	wire _w25384_ ;
	wire _w25383_ ;
	wire _w25382_ ;
	wire _w25381_ ;
	wire _w25380_ ;
	wire _w25379_ ;
	wire _w25378_ ;
	wire _w25377_ ;
	wire _w25376_ ;
	wire _w25375_ ;
	wire _w25374_ ;
	wire _w25373_ ;
	wire _w25372_ ;
	wire _w25371_ ;
	wire _w25370_ ;
	wire _w25369_ ;
	wire _w25368_ ;
	wire _w25367_ ;
	wire _w25366_ ;
	wire _w25365_ ;
	wire _w25364_ ;
	wire _w25363_ ;
	wire _w25362_ ;
	wire _w25361_ ;
	wire _w25360_ ;
	wire _w25359_ ;
	wire _w25358_ ;
	wire _w25357_ ;
	wire _w25356_ ;
	wire _w25355_ ;
	wire _w25354_ ;
	wire _w25353_ ;
	wire _w25352_ ;
	wire _w25351_ ;
	wire _w25350_ ;
	wire _w25349_ ;
	wire _w25348_ ;
	wire _w25347_ ;
	wire _w25346_ ;
	wire _w25345_ ;
	wire _w25344_ ;
	wire _w25343_ ;
	wire _w25342_ ;
	wire _w25341_ ;
	wire _w25340_ ;
	wire _w25339_ ;
	wire _w25338_ ;
	wire _w25337_ ;
	wire _w25336_ ;
	wire _w25335_ ;
	wire _w25334_ ;
	wire _w25333_ ;
	wire _w25332_ ;
	wire _w25331_ ;
	wire _w25330_ ;
	wire _w25329_ ;
	wire _w25328_ ;
	wire _w25327_ ;
	wire _w25326_ ;
	wire _w25325_ ;
	wire _w25324_ ;
	wire _w25323_ ;
	wire _w25322_ ;
	wire _w25321_ ;
	wire _w25320_ ;
	wire _w25319_ ;
	wire _w25318_ ;
	wire _w25317_ ;
	wire _w25316_ ;
	wire _w25315_ ;
	wire _w25314_ ;
	wire _w25313_ ;
	wire _w25312_ ;
	wire _w25311_ ;
	wire _w25310_ ;
	wire _w25309_ ;
	wire _w25308_ ;
	wire _w25307_ ;
	wire _w25306_ ;
	wire _w25305_ ;
	wire _w25304_ ;
	wire _w25303_ ;
	wire _w25302_ ;
	wire _w25301_ ;
	wire _w25300_ ;
	wire _w25299_ ;
	wire _w25298_ ;
	wire _w25297_ ;
	wire _w25296_ ;
	wire _w25295_ ;
	wire _w25294_ ;
	wire _w25293_ ;
	wire _w25292_ ;
	wire _w25291_ ;
	wire _w25290_ ;
	wire _w25289_ ;
	wire _w25288_ ;
	wire _w25287_ ;
	wire _w25286_ ;
	wire _w25285_ ;
	wire _w25284_ ;
	wire _w25283_ ;
	wire _w25282_ ;
	wire _w25281_ ;
	wire _w25280_ ;
	wire _w25279_ ;
	wire _w25278_ ;
	wire _w25277_ ;
	wire _w25276_ ;
	wire _w25275_ ;
	wire _w25274_ ;
	wire _w25273_ ;
	wire _w25272_ ;
	wire _w25271_ ;
	wire _w25270_ ;
	wire _w25269_ ;
	wire _w25268_ ;
	wire _w25267_ ;
	wire _w25266_ ;
	wire _w25265_ ;
	wire _w25264_ ;
	wire _w25263_ ;
	wire _w25262_ ;
	wire _w25261_ ;
	wire _w25260_ ;
	wire _w25259_ ;
	wire _w25258_ ;
	wire _w25257_ ;
	wire _w25256_ ;
	wire _w25255_ ;
	wire _w25254_ ;
	wire _w25253_ ;
	wire _w25252_ ;
	wire _w25251_ ;
	wire _w25250_ ;
	wire _w25249_ ;
	wire _w25248_ ;
	wire _w25247_ ;
	wire _w25246_ ;
	wire _w25245_ ;
	wire _w25244_ ;
	wire _w25243_ ;
	wire _w25242_ ;
	wire _w25241_ ;
	wire _w25240_ ;
	wire _w25239_ ;
	wire _w25238_ ;
	wire _w25237_ ;
	wire _w25236_ ;
	wire _w25235_ ;
	wire _w25234_ ;
	wire _w25233_ ;
	wire _w25232_ ;
	wire _w25231_ ;
	wire _w25230_ ;
	wire _w25229_ ;
	wire _w25228_ ;
	wire _w25227_ ;
	wire _w25226_ ;
	wire _w25225_ ;
	wire _w25224_ ;
	wire _w25223_ ;
	wire _w25222_ ;
	wire _w25221_ ;
	wire _w25220_ ;
	wire _w25219_ ;
	wire _w25218_ ;
	wire _w25217_ ;
	wire _w25216_ ;
	wire _w25215_ ;
	wire _w25214_ ;
	wire _w25213_ ;
	wire _w25212_ ;
	wire _w25211_ ;
	wire _w25210_ ;
	wire _w25209_ ;
	wire _w25208_ ;
	wire _w25207_ ;
	wire _w25206_ ;
	wire _w25205_ ;
	wire _w25204_ ;
	wire _w25203_ ;
	wire _w25202_ ;
	wire _w25201_ ;
	wire _w25200_ ;
	wire _w25199_ ;
	wire _w25198_ ;
	wire _w25197_ ;
	wire _w25196_ ;
	wire _w25195_ ;
	wire _w25194_ ;
	wire _w25193_ ;
	wire _w25192_ ;
	wire _w25191_ ;
	wire _w25190_ ;
	wire _w25189_ ;
	wire _w25188_ ;
	wire _w25187_ ;
	wire _w25186_ ;
	wire _w25185_ ;
	wire _w25184_ ;
	wire _w25183_ ;
	wire _w25182_ ;
	wire _w25181_ ;
	wire _w25180_ ;
	wire _w25179_ ;
	wire _w25178_ ;
	wire _w25177_ ;
	wire _w25176_ ;
	wire _w25175_ ;
	wire _w25174_ ;
	wire _w25173_ ;
	wire _w25172_ ;
	wire _w25171_ ;
	wire _w25170_ ;
	wire _w25169_ ;
	wire _w25168_ ;
	wire _w25167_ ;
	wire _w25166_ ;
	wire _w25165_ ;
	wire _w25164_ ;
	wire _w25163_ ;
	wire _w25162_ ;
	wire _w25161_ ;
	wire _w25160_ ;
	wire _w25159_ ;
	wire _w25158_ ;
	wire _w25157_ ;
	wire _w25156_ ;
	wire _w25155_ ;
	wire _w25154_ ;
	wire _w25153_ ;
	wire _w25152_ ;
	wire _w25151_ ;
	wire _w25150_ ;
	wire _w25149_ ;
	wire _w25148_ ;
	wire _w25147_ ;
	wire _w25146_ ;
	wire _w25145_ ;
	wire _w25144_ ;
	wire _w25143_ ;
	wire _w25142_ ;
	wire _w25141_ ;
	wire _w25140_ ;
	wire _w25139_ ;
	wire _w25138_ ;
	wire _w25137_ ;
	wire _w25136_ ;
	wire _w25135_ ;
	wire _w25134_ ;
	wire _w25133_ ;
	wire _w25132_ ;
	wire _w25131_ ;
	wire _w25130_ ;
	wire _w25129_ ;
	wire _w25128_ ;
	wire _w25127_ ;
	wire _w25126_ ;
	wire _w25125_ ;
	wire _w25124_ ;
	wire _w25123_ ;
	wire _w25122_ ;
	wire _w25121_ ;
	wire _w25120_ ;
	wire _w25119_ ;
	wire _w25118_ ;
	wire _w25117_ ;
	wire _w25116_ ;
	wire _w25115_ ;
	wire _w25114_ ;
	wire _w25113_ ;
	wire _w25112_ ;
	wire _w25111_ ;
	wire _w25110_ ;
	wire _w25109_ ;
	wire _w25108_ ;
	wire _w25107_ ;
	wire _w25106_ ;
	wire _w25105_ ;
	wire _w25104_ ;
	wire _w25103_ ;
	wire _w25102_ ;
	wire _w25101_ ;
	wire _w25100_ ;
	wire _w25099_ ;
	wire _w25098_ ;
	wire _w25097_ ;
	wire _w25096_ ;
	wire _w25095_ ;
	wire _w25094_ ;
	wire _w25093_ ;
	wire _w25092_ ;
	wire _w25091_ ;
	wire _w25090_ ;
	wire _w25089_ ;
	wire _w25088_ ;
	wire _w25087_ ;
	wire _w25086_ ;
	wire _w25085_ ;
	wire _w25084_ ;
	wire _w25083_ ;
	wire _w25082_ ;
	wire _w25081_ ;
	wire _w25080_ ;
	wire _w25079_ ;
	wire _w25078_ ;
	wire _w25077_ ;
	wire _w25076_ ;
	wire _w25075_ ;
	wire _w25074_ ;
	wire _w25073_ ;
	wire _w25072_ ;
	wire _w25071_ ;
	wire _w25070_ ;
	wire _w25069_ ;
	wire _w25068_ ;
	wire _w25067_ ;
	wire _w25066_ ;
	wire _w25065_ ;
	wire _w25064_ ;
	wire _w25063_ ;
	wire _w25062_ ;
	wire _w25061_ ;
	wire _w25060_ ;
	wire _w25059_ ;
	wire _w25058_ ;
	wire _w25057_ ;
	wire _w25056_ ;
	wire _w25055_ ;
	wire _w25054_ ;
	wire _w25053_ ;
	wire _w25052_ ;
	wire _w25051_ ;
	wire _w25050_ ;
	wire _w25049_ ;
	wire _w25048_ ;
	wire _w25047_ ;
	wire _w25046_ ;
	wire _w25045_ ;
	wire _w25044_ ;
	wire _w25043_ ;
	wire _w25042_ ;
	wire _w25041_ ;
	wire _w25040_ ;
	wire _w25039_ ;
	wire _w25038_ ;
	wire _w25037_ ;
	wire _w25036_ ;
	wire _w25035_ ;
	wire _w25034_ ;
	wire _w25033_ ;
	wire _w25032_ ;
	wire _w25031_ ;
	wire _w25030_ ;
	wire _w25029_ ;
	wire _w25028_ ;
	wire _w25027_ ;
	wire _w25026_ ;
	wire _w25025_ ;
	wire _w25024_ ;
	wire _w25023_ ;
	wire _w25022_ ;
	wire _w25021_ ;
	wire _w25020_ ;
	wire _w25019_ ;
	wire _w25018_ ;
	wire _w25017_ ;
	wire _w25016_ ;
	wire _w25015_ ;
	wire _w25014_ ;
	wire _w25013_ ;
	wire _w25012_ ;
	wire _w25011_ ;
	wire _w25010_ ;
	wire _w25009_ ;
	wire _w25008_ ;
	wire _w25007_ ;
	wire _w25006_ ;
	wire _w25005_ ;
	wire _w25004_ ;
	wire _w25003_ ;
	wire _w25002_ ;
	wire _w25001_ ;
	wire _w25000_ ;
	wire _w24999_ ;
	wire _w24998_ ;
	wire _w24997_ ;
	wire _w24996_ ;
	wire _w24995_ ;
	wire _w24994_ ;
	wire _w24993_ ;
	wire _w24992_ ;
	wire _w24991_ ;
	wire _w24990_ ;
	wire _w24989_ ;
	wire _w24988_ ;
	wire _w24987_ ;
	wire _w24986_ ;
	wire _w24985_ ;
	wire _w24984_ ;
	wire _w24983_ ;
	wire _w24982_ ;
	wire _w24981_ ;
	wire _w24980_ ;
	wire _w24979_ ;
	wire _w24978_ ;
	wire _w24977_ ;
	wire _w24976_ ;
	wire _w24975_ ;
	wire _w24974_ ;
	wire _w24973_ ;
	wire _w24972_ ;
	wire _w24971_ ;
	wire _w24970_ ;
	wire _w24969_ ;
	wire _w24968_ ;
	wire _w24967_ ;
	wire _w24966_ ;
	wire _w24965_ ;
	wire _w24964_ ;
	wire _w24963_ ;
	wire _w24962_ ;
	wire _w24961_ ;
	wire _w24960_ ;
	wire _w24959_ ;
	wire _w24958_ ;
	wire _w24957_ ;
	wire _w24956_ ;
	wire _w24955_ ;
	wire _w24954_ ;
	wire _w24953_ ;
	wire _w24952_ ;
	wire _w24951_ ;
	wire _w24950_ ;
	wire _w24949_ ;
	wire _w24948_ ;
	wire _w24947_ ;
	wire _w24946_ ;
	wire _w24945_ ;
	wire _w24944_ ;
	wire _w24943_ ;
	wire _w24942_ ;
	wire _w24941_ ;
	wire _w24940_ ;
	wire _w24939_ ;
	wire _w24938_ ;
	wire _w24937_ ;
	wire _w24936_ ;
	wire _w24935_ ;
	wire _w24934_ ;
	wire _w24933_ ;
	wire _w24932_ ;
	wire _w24931_ ;
	wire _w24930_ ;
	wire _w24929_ ;
	wire _w24928_ ;
	wire _w24927_ ;
	wire _w24926_ ;
	wire _w24925_ ;
	wire _w24924_ ;
	wire _w24923_ ;
	wire _w24922_ ;
	wire _w24921_ ;
	wire _w24920_ ;
	wire _w24919_ ;
	wire _w24918_ ;
	wire _w24917_ ;
	wire _w24916_ ;
	wire _w24915_ ;
	wire _w24914_ ;
	wire _w24913_ ;
	wire _w24912_ ;
	wire _w24911_ ;
	wire _w24910_ ;
	wire _w24909_ ;
	wire _w24908_ ;
	wire _w24907_ ;
	wire _w24906_ ;
	wire _w24905_ ;
	wire _w24904_ ;
	wire _w24903_ ;
	wire _w24902_ ;
	wire _w24901_ ;
	wire _w24900_ ;
	wire _w24899_ ;
	wire _w24898_ ;
	wire _w24897_ ;
	wire _w24896_ ;
	wire _w24895_ ;
	wire _w24894_ ;
	wire _w24893_ ;
	wire _w24892_ ;
	wire _w24891_ ;
	wire _w24890_ ;
	wire _w24889_ ;
	wire _w24888_ ;
	wire _w24887_ ;
	wire _w24886_ ;
	wire _w24885_ ;
	wire _w24884_ ;
	wire _w24883_ ;
	wire _w24882_ ;
	wire _w24881_ ;
	wire _w24880_ ;
	wire _w24879_ ;
	wire _w24878_ ;
	wire _w24877_ ;
	wire _w24876_ ;
	wire _w24875_ ;
	wire _w24874_ ;
	wire _w24873_ ;
	wire _w24872_ ;
	wire _w24871_ ;
	wire _w24870_ ;
	wire _w24869_ ;
	wire _w24868_ ;
	wire _w24867_ ;
	wire _w24866_ ;
	wire _w24865_ ;
	wire _w24864_ ;
	wire _w24863_ ;
	wire _w24862_ ;
	wire _w24861_ ;
	wire _w24860_ ;
	wire _w24859_ ;
	wire _w24858_ ;
	wire _w24857_ ;
	wire _w24856_ ;
	wire _w24855_ ;
	wire _w24854_ ;
	wire _w24853_ ;
	wire _w24852_ ;
	wire _w24851_ ;
	wire _w24850_ ;
	wire _w24849_ ;
	wire _w24848_ ;
	wire _w24847_ ;
	wire _w24846_ ;
	wire _w24845_ ;
	wire _w24844_ ;
	wire _w24843_ ;
	wire _w24842_ ;
	wire _w24841_ ;
	wire _w24840_ ;
	wire _w24839_ ;
	wire _w24838_ ;
	wire _w24837_ ;
	wire _w24836_ ;
	wire _w24835_ ;
	wire _w24834_ ;
	wire _w24833_ ;
	wire _w24832_ ;
	wire _w24831_ ;
	wire _w24830_ ;
	wire _w24829_ ;
	wire _w24828_ ;
	wire _w24827_ ;
	wire _w24826_ ;
	wire _w24825_ ;
	wire _w24824_ ;
	wire _w24823_ ;
	wire _w24822_ ;
	wire _w24821_ ;
	wire _w24820_ ;
	wire _w24819_ ;
	wire _w24818_ ;
	wire _w24817_ ;
	wire _w24816_ ;
	wire _w24815_ ;
	wire _w24814_ ;
	wire _w24813_ ;
	wire _w24812_ ;
	wire _w24811_ ;
	wire _w24810_ ;
	wire _w24809_ ;
	wire _w24808_ ;
	wire _w24807_ ;
	wire _w24806_ ;
	wire _w24805_ ;
	wire _w24804_ ;
	wire _w24803_ ;
	wire _w24802_ ;
	wire _w24801_ ;
	wire _w24800_ ;
	wire _w24799_ ;
	wire _w24798_ ;
	wire _w24797_ ;
	wire _w24796_ ;
	wire _w24795_ ;
	wire _w24794_ ;
	wire _w24793_ ;
	wire _w24792_ ;
	wire _w24791_ ;
	wire _w24790_ ;
	wire _w24789_ ;
	wire _w24788_ ;
	wire _w24787_ ;
	wire _w24786_ ;
	wire _w24785_ ;
	wire _w24784_ ;
	wire _w24783_ ;
	wire _w24782_ ;
	wire _w24781_ ;
	wire _w24780_ ;
	wire _w24779_ ;
	wire _w24778_ ;
	wire _w24777_ ;
	wire _w24776_ ;
	wire _w24775_ ;
	wire _w24774_ ;
	wire _w24773_ ;
	wire _w24772_ ;
	wire _w24771_ ;
	wire _w24770_ ;
	wire _w24769_ ;
	wire _w24768_ ;
	wire _w24767_ ;
	wire _w24766_ ;
	wire _w24765_ ;
	wire _w24764_ ;
	wire _w24763_ ;
	wire _w24762_ ;
	wire _w24761_ ;
	wire _w24760_ ;
	wire _w24759_ ;
	wire _w24758_ ;
	wire _w24757_ ;
	wire _w24756_ ;
	wire _w24755_ ;
	wire _w24754_ ;
	wire _w24753_ ;
	wire _w24752_ ;
	wire _w24751_ ;
	wire _w24750_ ;
	wire _w24749_ ;
	wire _w24748_ ;
	wire _w24747_ ;
	wire _w24746_ ;
	wire _w24745_ ;
	wire _w24744_ ;
	wire _w24743_ ;
	wire _w24742_ ;
	wire _w24741_ ;
	wire _w24740_ ;
	wire _w24739_ ;
	wire _w24738_ ;
	wire _w24737_ ;
	wire _w24736_ ;
	wire _w24735_ ;
	wire _w24734_ ;
	wire _w24733_ ;
	wire _w24732_ ;
	wire _w24731_ ;
	wire _w24730_ ;
	wire _w24729_ ;
	wire _w24728_ ;
	wire _w24727_ ;
	wire _w24726_ ;
	wire _w24725_ ;
	wire _w24724_ ;
	wire _w24723_ ;
	wire _w24722_ ;
	wire _w24721_ ;
	wire _w24720_ ;
	wire _w24719_ ;
	wire _w24718_ ;
	wire _w24717_ ;
	wire _w24716_ ;
	wire _w24715_ ;
	wire _w24714_ ;
	wire _w24713_ ;
	wire _w24712_ ;
	wire _w24711_ ;
	wire _w24710_ ;
	wire _w24709_ ;
	wire _w24708_ ;
	wire _w24707_ ;
	wire _w24706_ ;
	wire _w24705_ ;
	wire _w24704_ ;
	wire _w24703_ ;
	wire _w24702_ ;
	wire _w24701_ ;
	wire _w24700_ ;
	wire _w24699_ ;
	wire _w24698_ ;
	wire _w24697_ ;
	wire _w24696_ ;
	wire _w24695_ ;
	wire _w24694_ ;
	wire _w24693_ ;
	wire _w24692_ ;
	wire _w24691_ ;
	wire _w24690_ ;
	wire _w24689_ ;
	wire _w24688_ ;
	wire _w24687_ ;
	wire _w24686_ ;
	wire _w24685_ ;
	wire _w24684_ ;
	wire _w24683_ ;
	wire _w24682_ ;
	wire _w24681_ ;
	wire _w24680_ ;
	wire _w24679_ ;
	wire _w24678_ ;
	wire _w24677_ ;
	wire _w24676_ ;
	wire _w24675_ ;
	wire _w24674_ ;
	wire _w24673_ ;
	wire _w24672_ ;
	wire _w24671_ ;
	wire _w24670_ ;
	wire _w24669_ ;
	wire _w24668_ ;
	wire _w24667_ ;
	wire _w24666_ ;
	wire _w24665_ ;
	wire _w24664_ ;
	wire _w24663_ ;
	wire _w24662_ ;
	wire _w24661_ ;
	wire _w24660_ ;
	wire _w24659_ ;
	wire _w24658_ ;
	wire _w24657_ ;
	wire _w24656_ ;
	wire _w24655_ ;
	wire _w24654_ ;
	wire _w24653_ ;
	wire _w24652_ ;
	wire _w24651_ ;
	wire _w24650_ ;
	wire _w24649_ ;
	wire _w24648_ ;
	wire _w24647_ ;
	wire _w24646_ ;
	wire _w24645_ ;
	wire _w24644_ ;
	wire _w24643_ ;
	wire _w24642_ ;
	wire _w24641_ ;
	wire _w24640_ ;
	wire _w24639_ ;
	wire _w24638_ ;
	wire _w24637_ ;
	wire _w24636_ ;
	wire _w24635_ ;
	wire _w24634_ ;
	wire _w24633_ ;
	wire _w24632_ ;
	wire _w24631_ ;
	wire _w24630_ ;
	wire _w24629_ ;
	wire _w24628_ ;
	wire _w24627_ ;
	wire _w24626_ ;
	wire _w24625_ ;
	wire _w24624_ ;
	wire _w24623_ ;
	wire _w24622_ ;
	wire _w24621_ ;
	wire _w24620_ ;
	wire _w24619_ ;
	wire _w24618_ ;
	wire _w24617_ ;
	wire _w24616_ ;
	wire _w24615_ ;
	wire _w24614_ ;
	wire _w24613_ ;
	wire _w24612_ ;
	wire _w24611_ ;
	wire _w24610_ ;
	wire _w24609_ ;
	wire _w24608_ ;
	wire _w24607_ ;
	wire _w24606_ ;
	wire _w24605_ ;
	wire _w24604_ ;
	wire _w24603_ ;
	wire _w24602_ ;
	wire _w24601_ ;
	wire _w24600_ ;
	wire _w24599_ ;
	wire _w24598_ ;
	wire _w24597_ ;
	wire _w24596_ ;
	wire _w24595_ ;
	wire _w24594_ ;
	wire _w24593_ ;
	wire _w24592_ ;
	wire _w24591_ ;
	wire _w24590_ ;
	wire _w24589_ ;
	wire _w24588_ ;
	wire _w24587_ ;
	wire _w24586_ ;
	wire _w24585_ ;
	wire _w24584_ ;
	wire _w24583_ ;
	wire _w24582_ ;
	wire _w24581_ ;
	wire _w24580_ ;
	wire _w24579_ ;
	wire _w24578_ ;
	wire _w24577_ ;
	wire _w24576_ ;
	wire _w24575_ ;
	wire _w24574_ ;
	wire _w24573_ ;
	wire _w24572_ ;
	wire _w24571_ ;
	wire _w24570_ ;
	wire _w24569_ ;
	wire _w24568_ ;
	wire _w24567_ ;
	wire _w24566_ ;
	wire _w24565_ ;
	wire _w24564_ ;
	wire _w24563_ ;
	wire _w24562_ ;
	wire _w24561_ ;
	wire _w24560_ ;
	wire _w24559_ ;
	wire _w24558_ ;
	wire _w24557_ ;
	wire _w24556_ ;
	wire _w24555_ ;
	wire _w24554_ ;
	wire _w24553_ ;
	wire _w24552_ ;
	wire _w24551_ ;
	wire _w24550_ ;
	wire _w24549_ ;
	wire _w24548_ ;
	wire _w24547_ ;
	wire _w24546_ ;
	wire _w24545_ ;
	wire _w24544_ ;
	wire _w24543_ ;
	wire _w24542_ ;
	wire _w24541_ ;
	wire _w24540_ ;
	wire _w24539_ ;
	wire _w24538_ ;
	wire _w24537_ ;
	wire _w24536_ ;
	wire _w24535_ ;
	wire _w24534_ ;
	wire _w24533_ ;
	wire _w24532_ ;
	wire _w24531_ ;
	wire _w24530_ ;
	wire _w24529_ ;
	wire _w24528_ ;
	wire _w24527_ ;
	wire _w24526_ ;
	wire _w24525_ ;
	wire _w24524_ ;
	wire _w24523_ ;
	wire _w24522_ ;
	wire _w24521_ ;
	wire _w24520_ ;
	wire _w24519_ ;
	wire _w24518_ ;
	wire _w24517_ ;
	wire _w24516_ ;
	wire _w24515_ ;
	wire _w24514_ ;
	wire _w24513_ ;
	wire _w24512_ ;
	wire _w24511_ ;
	wire _w24510_ ;
	wire _w24509_ ;
	wire _w24508_ ;
	wire _w24507_ ;
	wire _w24506_ ;
	wire _w24505_ ;
	wire _w24504_ ;
	wire _w24503_ ;
	wire _w24502_ ;
	wire _w24501_ ;
	wire _w24500_ ;
	wire _w24499_ ;
	wire _w24498_ ;
	wire _w24497_ ;
	wire _w24496_ ;
	wire _w24495_ ;
	wire _w24494_ ;
	wire _w24493_ ;
	wire _w24492_ ;
	wire _w24491_ ;
	wire _w24490_ ;
	wire _w24489_ ;
	wire _w24488_ ;
	wire _w24487_ ;
	wire _w24486_ ;
	wire _w24485_ ;
	wire _w24484_ ;
	wire _w24483_ ;
	wire _w24482_ ;
	wire _w24481_ ;
	wire _w24480_ ;
	wire _w24479_ ;
	wire _w24478_ ;
	wire _w24477_ ;
	wire _w24476_ ;
	wire _w24475_ ;
	wire _w24474_ ;
	wire _w24473_ ;
	wire _w24472_ ;
	wire _w24471_ ;
	wire _w24470_ ;
	wire _w24469_ ;
	wire _w24468_ ;
	wire _w24467_ ;
	wire _w24466_ ;
	wire _w24465_ ;
	wire _w24464_ ;
	wire _w24463_ ;
	wire _w24462_ ;
	wire _w24461_ ;
	wire _w24460_ ;
	wire _w24459_ ;
	wire _w24458_ ;
	wire _w24457_ ;
	wire _w24456_ ;
	wire _w24455_ ;
	wire _w24454_ ;
	wire _w24453_ ;
	wire _w24452_ ;
	wire _w24451_ ;
	wire _w24450_ ;
	wire _w24449_ ;
	wire _w24448_ ;
	wire _w24447_ ;
	wire _w24446_ ;
	wire _w24445_ ;
	wire _w24444_ ;
	wire _w24443_ ;
	wire _w24442_ ;
	wire _w24441_ ;
	wire _w24440_ ;
	wire _w24439_ ;
	wire _w24438_ ;
	wire _w24437_ ;
	wire _w24436_ ;
	wire _w24435_ ;
	wire _w24434_ ;
	wire _w24433_ ;
	wire _w24432_ ;
	wire _w24431_ ;
	wire _w24430_ ;
	wire _w24429_ ;
	wire _w24428_ ;
	wire _w24427_ ;
	wire _w24426_ ;
	wire _w24425_ ;
	wire _w24424_ ;
	wire _w24423_ ;
	wire _w24422_ ;
	wire _w24421_ ;
	wire _w24420_ ;
	wire _w24419_ ;
	wire _w24418_ ;
	wire _w24417_ ;
	wire _w24416_ ;
	wire _w24415_ ;
	wire _w24414_ ;
	wire _w24413_ ;
	wire _w24412_ ;
	wire _w24411_ ;
	wire _w24410_ ;
	wire _w24409_ ;
	wire _w24408_ ;
	wire _w24407_ ;
	wire _w24406_ ;
	wire _w24405_ ;
	wire _w24404_ ;
	wire _w24403_ ;
	wire _w24402_ ;
	wire _w24401_ ;
	wire _w24400_ ;
	wire _w24399_ ;
	wire _w24398_ ;
	wire _w24397_ ;
	wire _w24396_ ;
	wire _w24395_ ;
	wire _w24394_ ;
	wire _w24393_ ;
	wire _w24392_ ;
	wire _w24391_ ;
	wire _w24390_ ;
	wire _w24389_ ;
	wire _w24388_ ;
	wire _w24387_ ;
	wire _w24386_ ;
	wire _w24385_ ;
	wire _w24384_ ;
	wire _w24383_ ;
	wire _w24382_ ;
	wire _w24381_ ;
	wire _w24380_ ;
	wire _w24379_ ;
	wire _w24378_ ;
	wire _w24377_ ;
	wire _w24376_ ;
	wire _w24375_ ;
	wire _w24374_ ;
	wire _w24373_ ;
	wire _w24372_ ;
	wire _w24371_ ;
	wire _w24370_ ;
	wire _w24369_ ;
	wire _w24368_ ;
	wire _w24367_ ;
	wire _w24366_ ;
	wire _w24365_ ;
	wire _w24364_ ;
	wire _w24363_ ;
	wire _w24362_ ;
	wire _w24361_ ;
	wire _w24360_ ;
	wire _w24359_ ;
	wire _w24358_ ;
	wire _w24357_ ;
	wire _w24356_ ;
	wire _w24355_ ;
	wire _w24354_ ;
	wire _w24353_ ;
	wire _w24352_ ;
	wire _w24351_ ;
	wire _w24350_ ;
	wire _w24349_ ;
	wire _w24348_ ;
	wire _w24347_ ;
	wire _w24346_ ;
	wire _w24345_ ;
	wire _w24344_ ;
	wire _w24343_ ;
	wire _w24342_ ;
	wire _w24341_ ;
	wire _w24340_ ;
	wire _w24339_ ;
	wire _w24338_ ;
	wire _w24337_ ;
	wire _w24336_ ;
	wire _w24335_ ;
	wire _w24334_ ;
	wire _w24333_ ;
	wire _w24332_ ;
	wire _w24331_ ;
	wire _w24330_ ;
	wire _w24329_ ;
	wire _w24328_ ;
	wire _w24327_ ;
	wire _w24326_ ;
	wire _w24325_ ;
	wire _w24324_ ;
	wire _w24323_ ;
	wire _w24322_ ;
	wire _w24321_ ;
	wire _w24320_ ;
	wire _w24319_ ;
	wire _w24318_ ;
	wire _w24317_ ;
	wire _w24316_ ;
	wire _w24315_ ;
	wire _w24314_ ;
	wire _w24313_ ;
	wire _w24312_ ;
	wire _w24311_ ;
	wire _w24310_ ;
	wire _w24309_ ;
	wire _w24308_ ;
	wire _w24307_ ;
	wire _w24306_ ;
	wire _w24305_ ;
	wire _w24304_ ;
	wire _w24303_ ;
	wire _w24302_ ;
	wire _w24301_ ;
	wire _w24300_ ;
	wire _w24299_ ;
	wire _w24298_ ;
	wire _w24297_ ;
	wire _w24296_ ;
	wire _w24295_ ;
	wire _w24294_ ;
	wire _w24293_ ;
	wire _w24292_ ;
	wire _w24291_ ;
	wire _w24290_ ;
	wire _w24289_ ;
	wire _w24288_ ;
	wire _w24287_ ;
	wire _w24286_ ;
	wire _w24285_ ;
	wire _w24284_ ;
	wire _w24283_ ;
	wire _w24282_ ;
	wire _w24281_ ;
	wire _w24280_ ;
	wire _w24279_ ;
	wire _w24278_ ;
	wire _w24277_ ;
	wire _w24276_ ;
	wire _w24275_ ;
	wire _w24274_ ;
	wire _w24273_ ;
	wire _w24272_ ;
	wire _w24271_ ;
	wire _w24270_ ;
	wire _w24269_ ;
	wire _w24268_ ;
	wire _w24267_ ;
	wire _w24266_ ;
	wire _w24265_ ;
	wire _w24264_ ;
	wire _w24263_ ;
	wire _w24262_ ;
	wire _w24261_ ;
	wire _w24260_ ;
	wire _w24259_ ;
	wire _w24258_ ;
	wire _w24257_ ;
	wire _w24256_ ;
	wire _w24255_ ;
	wire _w24254_ ;
	wire _w24253_ ;
	wire _w24252_ ;
	wire _w24251_ ;
	wire _w24250_ ;
	wire _w24249_ ;
	wire _w24248_ ;
	wire _w24247_ ;
	wire _w24246_ ;
	wire _w24245_ ;
	wire _w24244_ ;
	wire _w24243_ ;
	wire _w24242_ ;
	wire _w24241_ ;
	wire _w24240_ ;
	wire _w24239_ ;
	wire _w24238_ ;
	wire _w24237_ ;
	wire _w24236_ ;
	wire _w24235_ ;
	wire _w24234_ ;
	wire _w24233_ ;
	wire _w24232_ ;
	wire _w24231_ ;
	wire _w24230_ ;
	wire _w24229_ ;
	wire _w24228_ ;
	wire _w24227_ ;
	wire _w24226_ ;
	wire _w24225_ ;
	wire _w24224_ ;
	wire _w24223_ ;
	wire _w24222_ ;
	wire _w24221_ ;
	wire _w24220_ ;
	wire _w24219_ ;
	wire _w24218_ ;
	wire _w24217_ ;
	wire _w24216_ ;
	wire _w24215_ ;
	wire _w24214_ ;
	wire _w24213_ ;
	wire _w24212_ ;
	wire _w24211_ ;
	wire _w24210_ ;
	wire _w24209_ ;
	wire _w24208_ ;
	wire _w24207_ ;
	wire _w24206_ ;
	wire _w24205_ ;
	wire _w24204_ ;
	wire _w24203_ ;
	wire _w24202_ ;
	wire _w24201_ ;
	wire _w24200_ ;
	wire _w24199_ ;
	wire _w24198_ ;
	wire _w24197_ ;
	wire _w24196_ ;
	wire _w24195_ ;
	wire _w24194_ ;
	wire _w24193_ ;
	wire _w24192_ ;
	wire _w24191_ ;
	wire _w24190_ ;
	wire _w24189_ ;
	wire _w24188_ ;
	wire _w24187_ ;
	wire _w24186_ ;
	wire _w24185_ ;
	wire _w24184_ ;
	wire _w24183_ ;
	wire _w24182_ ;
	wire _w24181_ ;
	wire _w24180_ ;
	wire _w24179_ ;
	wire _w24178_ ;
	wire _w24177_ ;
	wire _w24176_ ;
	wire _w24175_ ;
	wire _w24174_ ;
	wire _w24173_ ;
	wire _w24172_ ;
	wire _w24171_ ;
	wire _w24170_ ;
	wire _w24169_ ;
	wire _w24168_ ;
	wire _w24167_ ;
	wire _w24166_ ;
	wire _w24165_ ;
	wire _w24164_ ;
	wire _w24163_ ;
	wire _w24162_ ;
	wire _w24161_ ;
	wire _w24160_ ;
	wire _w24159_ ;
	wire _w24158_ ;
	wire _w24157_ ;
	wire _w24156_ ;
	wire _w24155_ ;
	wire _w24154_ ;
	wire _w24153_ ;
	wire _w24152_ ;
	wire _w24151_ ;
	wire _w24150_ ;
	wire _w24149_ ;
	wire _w24148_ ;
	wire _w24147_ ;
	wire _w24146_ ;
	wire _w24145_ ;
	wire _w24144_ ;
	wire _w24143_ ;
	wire _w24142_ ;
	wire _w24141_ ;
	wire _w24140_ ;
	wire _w24139_ ;
	wire _w24138_ ;
	wire _w24137_ ;
	wire _w24136_ ;
	wire _w24135_ ;
	wire _w24134_ ;
	wire _w24133_ ;
	wire _w24132_ ;
	wire _w24131_ ;
	wire _w24130_ ;
	wire _w24129_ ;
	wire _w24128_ ;
	wire _w24127_ ;
	wire _w24126_ ;
	wire _w24125_ ;
	wire _w24124_ ;
	wire _w24123_ ;
	wire _w24122_ ;
	wire _w24121_ ;
	wire _w24120_ ;
	wire _w24119_ ;
	wire _w24118_ ;
	wire _w24117_ ;
	wire _w24116_ ;
	wire _w24115_ ;
	wire _w24114_ ;
	wire _w24113_ ;
	wire _w24112_ ;
	wire _w24111_ ;
	wire _w24110_ ;
	wire _w24109_ ;
	wire _w24108_ ;
	wire _w24107_ ;
	wire _w24106_ ;
	wire _w24105_ ;
	wire _w24104_ ;
	wire _w24103_ ;
	wire _w24102_ ;
	wire _w24101_ ;
	wire _w24100_ ;
	wire _w24099_ ;
	wire _w24098_ ;
	wire _w24097_ ;
	wire _w24096_ ;
	wire _w24095_ ;
	wire _w24094_ ;
	wire _w24093_ ;
	wire _w24092_ ;
	wire _w24091_ ;
	wire _w24090_ ;
	wire _w24089_ ;
	wire _w24088_ ;
	wire _w24087_ ;
	wire _w24086_ ;
	wire _w24085_ ;
	wire _w24084_ ;
	wire _w24083_ ;
	wire _w24082_ ;
	wire _w24081_ ;
	wire _w24080_ ;
	wire _w24079_ ;
	wire _w24078_ ;
	wire _w24077_ ;
	wire _w24076_ ;
	wire _w24075_ ;
	wire _w24074_ ;
	wire _w24073_ ;
	wire _w24072_ ;
	wire _w24071_ ;
	wire _w24070_ ;
	wire _w24069_ ;
	wire _w24068_ ;
	wire _w24067_ ;
	wire _w24066_ ;
	wire _w24065_ ;
	wire _w24064_ ;
	wire _w24063_ ;
	wire _w24062_ ;
	wire _w24061_ ;
	wire _w24060_ ;
	wire _w24059_ ;
	wire _w24058_ ;
	wire _w24057_ ;
	wire _w24056_ ;
	wire _w24055_ ;
	wire _w24054_ ;
	wire _w24053_ ;
	wire _w24052_ ;
	wire _w24051_ ;
	wire _w24050_ ;
	wire _w24049_ ;
	wire _w24048_ ;
	wire _w24047_ ;
	wire _w24046_ ;
	wire _w24045_ ;
	wire _w24044_ ;
	wire _w24043_ ;
	wire _w24042_ ;
	wire _w24041_ ;
	wire _w24040_ ;
	wire _w24039_ ;
	wire _w24038_ ;
	wire _w24037_ ;
	wire _w24036_ ;
	wire _w24035_ ;
	wire _w24034_ ;
	wire _w24033_ ;
	wire _w24032_ ;
	wire _w24031_ ;
	wire _w24030_ ;
	wire _w24029_ ;
	wire _w24028_ ;
	wire _w24027_ ;
	wire _w24026_ ;
	wire _w24025_ ;
	wire _w24024_ ;
	wire _w24023_ ;
	wire _w24022_ ;
	wire _w24021_ ;
	wire _w24020_ ;
	wire _w24019_ ;
	wire _w24018_ ;
	wire _w24017_ ;
	wire _w24016_ ;
	wire _w24015_ ;
	wire _w24014_ ;
	wire _w24013_ ;
	wire _w24012_ ;
	wire _w24011_ ;
	wire _w24010_ ;
	wire _w24009_ ;
	wire _w24008_ ;
	wire _w24007_ ;
	wire _w24006_ ;
	wire _w24005_ ;
	wire _w24004_ ;
	wire _w24003_ ;
	wire _w24002_ ;
	wire _w24001_ ;
	wire _w24000_ ;
	wire _w23999_ ;
	wire _w23998_ ;
	wire _w23997_ ;
	wire _w23996_ ;
	wire _w23995_ ;
	wire _w23994_ ;
	wire _w23993_ ;
	wire _w23992_ ;
	wire _w23991_ ;
	wire _w23990_ ;
	wire _w23989_ ;
	wire _w23988_ ;
	wire _w23987_ ;
	wire _w23986_ ;
	wire _w23985_ ;
	wire _w23984_ ;
	wire _w23983_ ;
	wire _w23982_ ;
	wire _w23981_ ;
	wire _w23980_ ;
	wire _w23979_ ;
	wire _w23978_ ;
	wire _w23977_ ;
	wire _w23976_ ;
	wire _w23975_ ;
	wire _w23974_ ;
	wire _w23973_ ;
	wire _w23972_ ;
	wire _w23971_ ;
	wire _w23970_ ;
	wire _w23969_ ;
	wire _w23968_ ;
	wire _w23967_ ;
	wire _w23966_ ;
	wire _w23965_ ;
	wire _w23964_ ;
	wire _w23963_ ;
	wire _w23962_ ;
	wire _w23961_ ;
	wire _w23960_ ;
	wire _w23959_ ;
	wire _w23958_ ;
	wire _w23957_ ;
	wire _w23956_ ;
	wire _w23955_ ;
	wire _w23954_ ;
	wire _w23953_ ;
	wire _w23952_ ;
	wire _w23951_ ;
	wire _w23950_ ;
	wire _w23949_ ;
	wire _w23948_ ;
	wire _w23947_ ;
	wire _w23946_ ;
	wire _w23945_ ;
	wire _w23944_ ;
	wire _w23943_ ;
	wire _w23942_ ;
	wire _w23941_ ;
	wire _w23940_ ;
	wire _w23939_ ;
	wire _w23938_ ;
	wire _w23937_ ;
	wire _w23936_ ;
	wire _w23935_ ;
	wire _w23934_ ;
	wire _w23933_ ;
	wire _w23932_ ;
	wire _w23931_ ;
	wire _w23930_ ;
	wire _w23929_ ;
	wire _w23928_ ;
	wire _w23927_ ;
	wire _w23926_ ;
	wire _w23925_ ;
	wire _w23924_ ;
	wire _w23923_ ;
	wire _w23922_ ;
	wire _w23921_ ;
	wire _w23920_ ;
	wire _w23919_ ;
	wire _w23918_ ;
	wire _w23917_ ;
	wire _w23916_ ;
	wire _w23915_ ;
	wire _w23914_ ;
	wire _w23913_ ;
	wire _w23912_ ;
	wire _w23911_ ;
	wire _w23910_ ;
	wire _w23909_ ;
	wire _w23908_ ;
	wire _w23907_ ;
	wire _w23906_ ;
	wire _w23905_ ;
	wire _w23904_ ;
	wire _w23903_ ;
	wire _w23902_ ;
	wire _w23901_ ;
	wire _w23900_ ;
	wire _w23899_ ;
	wire _w23898_ ;
	wire _w23897_ ;
	wire _w23896_ ;
	wire _w23895_ ;
	wire _w23894_ ;
	wire _w23893_ ;
	wire _w23892_ ;
	wire _w23891_ ;
	wire _w23890_ ;
	wire _w23889_ ;
	wire _w23888_ ;
	wire _w23887_ ;
	wire _w23886_ ;
	wire _w23885_ ;
	wire _w23884_ ;
	wire _w23883_ ;
	wire _w23882_ ;
	wire _w23881_ ;
	wire _w23880_ ;
	wire _w23879_ ;
	wire _w23878_ ;
	wire _w23877_ ;
	wire _w23876_ ;
	wire _w23875_ ;
	wire _w23874_ ;
	wire _w23873_ ;
	wire _w23872_ ;
	wire _w23871_ ;
	wire _w23870_ ;
	wire _w23869_ ;
	wire _w23868_ ;
	wire _w23867_ ;
	wire _w23866_ ;
	wire _w23865_ ;
	wire _w23864_ ;
	wire _w23863_ ;
	wire _w23862_ ;
	wire _w23861_ ;
	wire _w23860_ ;
	wire _w23859_ ;
	wire _w23858_ ;
	wire _w23857_ ;
	wire _w23856_ ;
	wire _w23855_ ;
	wire _w23854_ ;
	wire _w23853_ ;
	wire _w23852_ ;
	wire _w23851_ ;
	wire _w23850_ ;
	wire _w23849_ ;
	wire _w23848_ ;
	wire _w23847_ ;
	wire _w23846_ ;
	wire _w23845_ ;
	wire _w23844_ ;
	wire _w23843_ ;
	wire _w23842_ ;
	wire _w23841_ ;
	wire _w23840_ ;
	wire _w23839_ ;
	wire _w23838_ ;
	wire _w23837_ ;
	wire _w23836_ ;
	wire _w23835_ ;
	wire _w23834_ ;
	wire _w23833_ ;
	wire _w23832_ ;
	wire _w23831_ ;
	wire _w23830_ ;
	wire _w23829_ ;
	wire _w23828_ ;
	wire _w23827_ ;
	wire _w23826_ ;
	wire _w23825_ ;
	wire _w23824_ ;
	wire _w23823_ ;
	wire _w23822_ ;
	wire _w23821_ ;
	wire _w23820_ ;
	wire _w23819_ ;
	wire _w23818_ ;
	wire _w23817_ ;
	wire _w23816_ ;
	wire _w23815_ ;
	wire _w23814_ ;
	wire _w23813_ ;
	wire _w23812_ ;
	wire _w23811_ ;
	wire _w23810_ ;
	wire _w23809_ ;
	wire _w23808_ ;
	wire _w23807_ ;
	wire _w23806_ ;
	wire _w23805_ ;
	wire _w23804_ ;
	wire _w23803_ ;
	wire _w23802_ ;
	wire _w23801_ ;
	wire _w23800_ ;
	wire _w23799_ ;
	wire _w23798_ ;
	wire _w23797_ ;
	wire _w23796_ ;
	wire _w23795_ ;
	wire _w23794_ ;
	wire _w23793_ ;
	wire _w23792_ ;
	wire _w23791_ ;
	wire _w23790_ ;
	wire _w23789_ ;
	wire _w23788_ ;
	wire _w23787_ ;
	wire _w23786_ ;
	wire _w23785_ ;
	wire _w23784_ ;
	wire _w23783_ ;
	wire _w23782_ ;
	wire _w23781_ ;
	wire _w23780_ ;
	wire _w23779_ ;
	wire _w23778_ ;
	wire _w23777_ ;
	wire _w23776_ ;
	wire _w23775_ ;
	wire _w23774_ ;
	wire _w23773_ ;
	wire _w23772_ ;
	wire _w23771_ ;
	wire _w23770_ ;
	wire _w23769_ ;
	wire _w23768_ ;
	wire _w23767_ ;
	wire _w23766_ ;
	wire _w23765_ ;
	wire _w23764_ ;
	wire _w23763_ ;
	wire _w23762_ ;
	wire _w23761_ ;
	wire _w23760_ ;
	wire _w23759_ ;
	wire _w23758_ ;
	wire _w23757_ ;
	wire _w23756_ ;
	wire _w23755_ ;
	wire _w23754_ ;
	wire _w23753_ ;
	wire _w23752_ ;
	wire _w23751_ ;
	wire _w23750_ ;
	wire _w23749_ ;
	wire _w23748_ ;
	wire _w23747_ ;
	wire _w23746_ ;
	wire _w23745_ ;
	wire _w23744_ ;
	wire _w23743_ ;
	wire _w23742_ ;
	wire _w23741_ ;
	wire _w23740_ ;
	wire _w23739_ ;
	wire _w23738_ ;
	wire _w23737_ ;
	wire _w23736_ ;
	wire _w23735_ ;
	wire _w23734_ ;
	wire _w23733_ ;
	wire _w23732_ ;
	wire _w23731_ ;
	wire _w23730_ ;
	wire _w23729_ ;
	wire _w23728_ ;
	wire _w23727_ ;
	wire _w23726_ ;
	wire _w23725_ ;
	wire _w23724_ ;
	wire _w23723_ ;
	wire _w23722_ ;
	wire _w23721_ ;
	wire _w23720_ ;
	wire _w23719_ ;
	wire _w23718_ ;
	wire _w23717_ ;
	wire _w23716_ ;
	wire _w23715_ ;
	wire _w23714_ ;
	wire _w23713_ ;
	wire _w23712_ ;
	wire _w23711_ ;
	wire _w23710_ ;
	wire _w23709_ ;
	wire _w23708_ ;
	wire _w23707_ ;
	wire _w23706_ ;
	wire _w23705_ ;
	wire _w23704_ ;
	wire _w23703_ ;
	wire _w23702_ ;
	wire _w23701_ ;
	wire _w23700_ ;
	wire _w23699_ ;
	wire _w23698_ ;
	wire _w23697_ ;
	wire _w23696_ ;
	wire _w23695_ ;
	wire _w23694_ ;
	wire _w23693_ ;
	wire _w23692_ ;
	wire _w23691_ ;
	wire _w23690_ ;
	wire _w23689_ ;
	wire _w23688_ ;
	wire _w23687_ ;
	wire _w23686_ ;
	wire _w23685_ ;
	wire _w23684_ ;
	wire _w23683_ ;
	wire _w23682_ ;
	wire _w23681_ ;
	wire _w23680_ ;
	wire _w23679_ ;
	wire _w23678_ ;
	wire _w23677_ ;
	wire _w23676_ ;
	wire _w23675_ ;
	wire _w23674_ ;
	wire _w23673_ ;
	wire _w23672_ ;
	wire _w23671_ ;
	wire _w23670_ ;
	wire _w23669_ ;
	wire _w23668_ ;
	wire _w23667_ ;
	wire _w23666_ ;
	wire _w23665_ ;
	wire _w23664_ ;
	wire _w23663_ ;
	wire _w23662_ ;
	wire _w23661_ ;
	wire _w23660_ ;
	wire _w23659_ ;
	wire _w23658_ ;
	wire _w23657_ ;
	wire _w23656_ ;
	wire _w23655_ ;
	wire _w23654_ ;
	wire _w23653_ ;
	wire _w23652_ ;
	wire _w23651_ ;
	wire _w23650_ ;
	wire _w23649_ ;
	wire _w23648_ ;
	wire _w23647_ ;
	wire _w23646_ ;
	wire _w23645_ ;
	wire _w23644_ ;
	wire _w23643_ ;
	wire _w23642_ ;
	wire _w23641_ ;
	wire _w23640_ ;
	wire _w23639_ ;
	wire _w23638_ ;
	wire _w23637_ ;
	wire _w23636_ ;
	wire _w23635_ ;
	wire _w23634_ ;
	wire _w23633_ ;
	wire _w23632_ ;
	wire _w23631_ ;
	wire _w23630_ ;
	wire _w23629_ ;
	wire _w23628_ ;
	wire _w23627_ ;
	wire _w23626_ ;
	wire _w23625_ ;
	wire _w23624_ ;
	wire _w23623_ ;
	wire _w23622_ ;
	wire _w23621_ ;
	wire _w23620_ ;
	wire _w23619_ ;
	wire _w23618_ ;
	wire _w23617_ ;
	wire _w23616_ ;
	wire _w23615_ ;
	wire _w23614_ ;
	wire _w23613_ ;
	wire _w23612_ ;
	wire _w23611_ ;
	wire _w23610_ ;
	wire _w23609_ ;
	wire _w23608_ ;
	wire _w23607_ ;
	wire _w23606_ ;
	wire _w23605_ ;
	wire _w23604_ ;
	wire _w23603_ ;
	wire _w23602_ ;
	wire _w23601_ ;
	wire _w23600_ ;
	wire _w23599_ ;
	wire _w23598_ ;
	wire _w23597_ ;
	wire _w23596_ ;
	wire _w23595_ ;
	wire _w23594_ ;
	wire _w23593_ ;
	wire _w23592_ ;
	wire _w23591_ ;
	wire _w23590_ ;
	wire _w23589_ ;
	wire _w23588_ ;
	wire _w23587_ ;
	wire _w23586_ ;
	wire _w23585_ ;
	wire _w23584_ ;
	wire _w23583_ ;
	wire _w23582_ ;
	wire _w23581_ ;
	wire _w23580_ ;
	wire _w23579_ ;
	wire _w23578_ ;
	wire _w23577_ ;
	wire _w23576_ ;
	wire _w23575_ ;
	wire _w23574_ ;
	wire _w23573_ ;
	wire _w23572_ ;
	wire _w23571_ ;
	wire _w23570_ ;
	wire _w23569_ ;
	wire _w23568_ ;
	wire _w23567_ ;
	wire _w23566_ ;
	wire _w23565_ ;
	wire _w23564_ ;
	wire _w23563_ ;
	wire _w23562_ ;
	wire _w23561_ ;
	wire _w23560_ ;
	wire _w23559_ ;
	wire _w23558_ ;
	wire _w23557_ ;
	wire _w23556_ ;
	wire _w23555_ ;
	wire _w23554_ ;
	wire _w23553_ ;
	wire _w23552_ ;
	wire _w23551_ ;
	wire _w23550_ ;
	wire _w23549_ ;
	wire _w23548_ ;
	wire _w23547_ ;
	wire _w23546_ ;
	wire _w23545_ ;
	wire _w23544_ ;
	wire _w23543_ ;
	wire _w23542_ ;
	wire _w23541_ ;
	wire _w23540_ ;
	wire _w23539_ ;
	wire _w23538_ ;
	wire _w23537_ ;
	wire _w23536_ ;
	wire _w23535_ ;
	wire _w23534_ ;
	wire _w23533_ ;
	wire _w23532_ ;
	wire _w23531_ ;
	wire _w23530_ ;
	wire _w23529_ ;
	wire _w23528_ ;
	wire _w23527_ ;
	wire _w23526_ ;
	wire _w23525_ ;
	wire _w23524_ ;
	wire _w23523_ ;
	wire _w23522_ ;
	wire _w23521_ ;
	wire _w23520_ ;
	wire _w23519_ ;
	wire _w23518_ ;
	wire _w23517_ ;
	wire _w23516_ ;
	wire _w23515_ ;
	wire _w23514_ ;
	wire _w23513_ ;
	wire _w23512_ ;
	wire _w23511_ ;
	wire _w23510_ ;
	wire _w23509_ ;
	wire _w23508_ ;
	wire _w23507_ ;
	wire _w23506_ ;
	wire _w23505_ ;
	wire _w23504_ ;
	wire _w23503_ ;
	wire _w23502_ ;
	wire _w23501_ ;
	wire _w23500_ ;
	wire _w23499_ ;
	wire _w23498_ ;
	wire _w23497_ ;
	wire _w23496_ ;
	wire _w23495_ ;
	wire _w23494_ ;
	wire _w23493_ ;
	wire _w23492_ ;
	wire _w23491_ ;
	wire _w23490_ ;
	wire _w23489_ ;
	wire _w23488_ ;
	wire _w23487_ ;
	wire _w23486_ ;
	wire _w23485_ ;
	wire _w23484_ ;
	wire _w23483_ ;
	wire _w23482_ ;
	wire _w23481_ ;
	wire _w23480_ ;
	wire _w23479_ ;
	wire _w23478_ ;
	wire _w23477_ ;
	wire _w23476_ ;
	wire _w23475_ ;
	wire _w23474_ ;
	wire _w23473_ ;
	wire _w23472_ ;
	wire _w23471_ ;
	wire _w23470_ ;
	wire _w23469_ ;
	wire _w23468_ ;
	wire _w23467_ ;
	wire _w23466_ ;
	wire _w23465_ ;
	wire _w23464_ ;
	wire _w23463_ ;
	wire _w23462_ ;
	wire _w23461_ ;
	wire _w23460_ ;
	wire _w23459_ ;
	wire _w23458_ ;
	wire _w23457_ ;
	wire _w23456_ ;
	wire _w23455_ ;
	wire _w23454_ ;
	wire _w23453_ ;
	wire _w23452_ ;
	wire _w23451_ ;
	wire _w23450_ ;
	wire _w23449_ ;
	wire _w23448_ ;
	wire _w23447_ ;
	wire _w23446_ ;
	wire _w23445_ ;
	wire _w23444_ ;
	wire _w23443_ ;
	wire _w23442_ ;
	wire _w23441_ ;
	wire _w23440_ ;
	wire _w23439_ ;
	wire _w23438_ ;
	wire _w23437_ ;
	wire _w23436_ ;
	wire _w23435_ ;
	wire _w23434_ ;
	wire _w23433_ ;
	wire _w23432_ ;
	wire _w23431_ ;
	wire _w23430_ ;
	wire _w23429_ ;
	wire _w23428_ ;
	wire _w23427_ ;
	wire _w23426_ ;
	wire _w23425_ ;
	wire _w23424_ ;
	wire _w23423_ ;
	wire _w23422_ ;
	wire _w23421_ ;
	wire _w23420_ ;
	wire _w23419_ ;
	wire _w23418_ ;
	wire _w23417_ ;
	wire _w23416_ ;
	wire _w23415_ ;
	wire _w23414_ ;
	wire _w23413_ ;
	wire _w23412_ ;
	wire _w23411_ ;
	wire _w23410_ ;
	wire _w23409_ ;
	wire _w23408_ ;
	wire _w23407_ ;
	wire _w23406_ ;
	wire _w23405_ ;
	wire _w23404_ ;
	wire _w23403_ ;
	wire _w23402_ ;
	wire _w23401_ ;
	wire _w23400_ ;
	wire _w23399_ ;
	wire _w23398_ ;
	wire _w23397_ ;
	wire _w23396_ ;
	wire _w23395_ ;
	wire _w23394_ ;
	wire _w23393_ ;
	wire _w23392_ ;
	wire _w23391_ ;
	wire _w23390_ ;
	wire _w23389_ ;
	wire _w23388_ ;
	wire _w23387_ ;
	wire _w23386_ ;
	wire _w23385_ ;
	wire _w23384_ ;
	wire _w23383_ ;
	wire _w23382_ ;
	wire _w23381_ ;
	wire _w23380_ ;
	wire _w23379_ ;
	wire _w23378_ ;
	wire _w23377_ ;
	wire _w23376_ ;
	wire _w23375_ ;
	wire _w23374_ ;
	wire _w23373_ ;
	wire _w23372_ ;
	wire _w23371_ ;
	wire _w23370_ ;
	wire _w23369_ ;
	wire _w23368_ ;
	wire _w23367_ ;
	wire _w23366_ ;
	wire _w23365_ ;
	wire _w23364_ ;
	wire _w23363_ ;
	wire _w23362_ ;
	wire _w23361_ ;
	wire _w23360_ ;
	wire _w23359_ ;
	wire _w23358_ ;
	wire _w23357_ ;
	wire _w23356_ ;
	wire _w23355_ ;
	wire _w23354_ ;
	wire _w23353_ ;
	wire _w23352_ ;
	wire _w23351_ ;
	wire _w23350_ ;
	wire _w23349_ ;
	wire _w23348_ ;
	wire _w23347_ ;
	wire _w23346_ ;
	wire _w23345_ ;
	wire _w23344_ ;
	wire _w23343_ ;
	wire _w23342_ ;
	wire _w23341_ ;
	wire _w23340_ ;
	wire _w23339_ ;
	wire _w23338_ ;
	wire _w23337_ ;
	wire _w23336_ ;
	wire _w23335_ ;
	wire _w23334_ ;
	wire _w23333_ ;
	wire _w23332_ ;
	wire _w23331_ ;
	wire _w23330_ ;
	wire _w23329_ ;
	wire _w23328_ ;
	wire _w23327_ ;
	wire _w23326_ ;
	wire _w23325_ ;
	wire _w23324_ ;
	wire _w23323_ ;
	wire _w23322_ ;
	wire _w23321_ ;
	wire _w23320_ ;
	wire _w23319_ ;
	wire _w23318_ ;
	wire _w23317_ ;
	wire _w23316_ ;
	wire _w23315_ ;
	wire _w23314_ ;
	wire _w23313_ ;
	wire _w23312_ ;
	wire _w23311_ ;
	wire _w23310_ ;
	wire _w23309_ ;
	wire _w23308_ ;
	wire _w23307_ ;
	wire _w23306_ ;
	wire _w23305_ ;
	wire _w23304_ ;
	wire _w23303_ ;
	wire _w23302_ ;
	wire _w23301_ ;
	wire _w23300_ ;
	wire _w23299_ ;
	wire _w23298_ ;
	wire _w23297_ ;
	wire _w23296_ ;
	wire _w23295_ ;
	wire _w23294_ ;
	wire _w23293_ ;
	wire _w23292_ ;
	wire _w23291_ ;
	wire _w23290_ ;
	wire _w23289_ ;
	wire _w23288_ ;
	wire _w23287_ ;
	wire _w23286_ ;
	wire _w23285_ ;
	wire _w23284_ ;
	wire _w23283_ ;
	wire _w23282_ ;
	wire _w23281_ ;
	wire _w23280_ ;
	wire _w23279_ ;
	wire _w23278_ ;
	wire _w23277_ ;
	wire _w23276_ ;
	wire _w23275_ ;
	wire _w23274_ ;
	wire _w23273_ ;
	wire _w23272_ ;
	wire _w23271_ ;
	wire _w23270_ ;
	wire _w23269_ ;
	wire _w23268_ ;
	wire _w23267_ ;
	wire _w23266_ ;
	wire _w23265_ ;
	wire _w23264_ ;
	wire _w23263_ ;
	wire _w23262_ ;
	wire _w23261_ ;
	wire _w23260_ ;
	wire _w23259_ ;
	wire _w23258_ ;
	wire _w23257_ ;
	wire _w23256_ ;
	wire _w23255_ ;
	wire _w23254_ ;
	wire _w23253_ ;
	wire _w23252_ ;
	wire _w23251_ ;
	wire _w23250_ ;
	wire _w23249_ ;
	wire _w23248_ ;
	wire _w23247_ ;
	wire _w23246_ ;
	wire _w23245_ ;
	wire _w23244_ ;
	wire _w23243_ ;
	wire _w23242_ ;
	wire _w23241_ ;
	wire _w23240_ ;
	wire _w23239_ ;
	wire _w23238_ ;
	wire _w23237_ ;
	wire _w23236_ ;
	wire _w23235_ ;
	wire _w23234_ ;
	wire _w23233_ ;
	wire _w23232_ ;
	wire _w23231_ ;
	wire _w23230_ ;
	wire _w23229_ ;
	wire _w23228_ ;
	wire _w23227_ ;
	wire _w23226_ ;
	wire _w23225_ ;
	wire _w23224_ ;
	wire _w23223_ ;
	wire _w23222_ ;
	wire _w23221_ ;
	wire _w23220_ ;
	wire _w23219_ ;
	wire _w23218_ ;
	wire _w23217_ ;
	wire _w23216_ ;
	wire _w23215_ ;
	wire _w23214_ ;
	wire _w23213_ ;
	wire _w23212_ ;
	wire _w23211_ ;
	wire _w23210_ ;
	wire _w23209_ ;
	wire _w23208_ ;
	wire _w23207_ ;
	wire _w23206_ ;
	wire _w23205_ ;
	wire _w23204_ ;
	wire _w23203_ ;
	wire _w23202_ ;
	wire _w23201_ ;
	wire _w23200_ ;
	wire _w23199_ ;
	wire _w23198_ ;
	wire _w23197_ ;
	wire _w23196_ ;
	wire _w23195_ ;
	wire _w23194_ ;
	wire _w23193_ ;
	wire _w23192_ ;
	wire _w23191_ ;
	wire _w23190_ ;
	wire _w23189_ ;
	wire _w23188_ ;
	wire _w23187_ ;
	wire _w23186_ ;
	wire _w23185_ ;
	wire _w23184_ ;
	wire _w23183_ ;
	wire _w23182_ ;
	wire _w23181_ ;
	wire _w23180_ ;
	wire _w23179_ ;
	wire _w23178_ ;
	wire _w23177_ ;
	wire _w23176_ ;
	wire _w23175_ ;
	wire _w23174_ ;
	wire _w23173_ ;
	wire _w23172_ ;
	wire _w23171_ ;
	wire _w23170_ ;
	wire _w23169_ ;
	wire _w23168_ ;
	wire _w23167_ ;
	wire _w23166_ ;
	wire _w23165_ ;
	wire _w23164_ ;
	wire _w23163_ ;
	wire _w23162_ ;
	wire _w23161_ ;
	wire _w23160_ ;
	wire _w23159_ ;
	wire _w23158_ ;
	wire _w23157_ ;
	wire _w23156_ ;
	wire _w23155_ ;
	wire _w23154_ ;
	wire _w23153_ ;
	wire _w23152_ ;
	wire _w23151_ ;
	wire _w23150_ ;
	wire _w23149_ ;
	wire _w23148_ ;
	wire _w23147_ ;
	wire _w23146_ ;
	wire _w23145_ ;
	wire _w23144_ ;
	wire _w23143_ ;
	wire _w23142_ ;
	wire _w23141_ ;
	wire _w23140_ ;
	wire _w23139_ ;
	wire _w23138_ ;
	wire _w23137_ ;
	wire _w23136_ ;
	wire _w23135_ ;
	wire _w23134_ ;
	wire _w23133_ ;
	wire _w23132_ ;
	wire _w23131_ ;
	wire _w23130_ ;
	wire _w23129_ ;
	wire _w23128_ ;
	wire _w23127_ ;
	wire _w23126_ ;
	wire _w23125_ ;
	wire _w23124_ ;
	wire _w23123_ ;
	wire _w23122_ ;
	wire _w23121_ ;
	wire _w23120_ ;
	wire _w23119_ ;
	wire _w23118_ ;
	wire _w23117_ ;
	wire _w23116_ ;
	wire _w23115_ ;
	wire _w23114_ ;
	wire _w23113_ ;
	wire _w23112_ ;
	wire _w23111_ ;
	wire _w23110_ ;
	wire _w23109_ ;
	wire _w23108_ ;
	wire _w23107_ ;
	wire _w23106_ ;
	wire _w23105_ ;
	wire _w23104_ ;
	wire _w23103_ ;
	wire _w23102_ ;
	wire _w23101_ ;
	wire _w23100_ ;
	wire _w23099_ ;
	wire _w23098_ ;
	wire _w23097_ ;
	wire _w23096_ ;
	wire _w23095_ ;
	wire _w23094_ ;
	wire _w23093_ ;
	wire _w23092_ ;
	wire _w23091_ ;
	wire _w23090_ ;
	wire _w23089_ ;
	wire _w23088_ ;
	wire _w23087_ ;
	wire _w23086_ ;
	wire _w23085_ ;
	wire _w23084_ ;
	wire _w23083_ ;
	wire _w23082_ ;
	wire _w23081_ ;
	wire _w23080_ ;
	wire _w23079_ ;
	wire _w23078_ ;
	wire _w23077_ ;
	wire _w23076_ ;
	wire _w23075_ ;
	wire _w23074_ ;
	wire _w23073_ ;
	wire _w23072_ ;
	wire _w23071_ ;
	wire _w23070_ ;
	wire _w23069_ ;
	wire _w23068_ ;
	wire _w23067_ ;
	wire _w23066_ ;
	wire _w23065_ ;
	wire _w23064_ ;
	wire _w23063_ ;
	wire _w23062_ ;
	wire _w23061_ ;
	wire _w23060_ ;
	wire _w23059_ ;
	wire _w23058_ ;
	wire _w23057_ ;
	wire _w23056_ ;
	wire _w23055_ ;
	wire _w23054_ ;
	wire _w23053_ ;
	wire _w23052_ ;
	wire _w23051_ ;
	wire _w23050_ ;
	wire _w23049_ ;
	wire _w23048_ ;
	wire _w23047_ ;
	wire _w23046_ ;
	wire _w23045_ ;
	wire _w23044_ ;
	wire _w23043_ ;
	wire _w23042_ ;
	wire _w23041_ ;
	wire _w23040_ ;
	wire _w23039_ ;
	wire _w23038_ ;
	wire _w23037_ ;
	wire _w23036_ ;
	wire _w23035_ ;
	wire _w23034_ ;
	wire _w23033_ ;
	wire _w23032_ ;
	wire _w23031_ ;
	wire _w23030_ ;
	wire _w23029_ ;
	wire _w23028_ ;
	wire _w23027_ ;
	wire _w23026_ ;
	wire _w23025_ ;
	wire _w23024_ ;
	wire _w23023_ ;
	wire _w23022_ ;
	wire _w23021_ ;
	wire _w23020_ ;
	wire _w23019_ ;
	wire _w23018_ ;
	wire _w23017_ ;
	wire _w23016_ ;
	wire _w23015_ ;
	wire _w23014_ ;
	wire _w23013_ ;
	wire _w23012_ ;
	wire _w23011_ ;
	wire _w23010_ ;
	wire _w23009_ ;
	wire _w23008_ ;
	wire _w23007_ ;
	wire _w23006_ ;
	wire _w23005_ ;
	wire _w23004_ ;
	wire _w23003_ ;
	wire _w23002_ ;
	wire _w23001_ ;
	wire _w23000_ ;
	wire _w22999_ ;
	wire _w22998_ ;
	wire _w22997_ ;
	wire _w22996_ ;
	wire _w22995_ ;
	wire _w22994_ ;
	wire _w22993_ ;
	wire _w22992_ ;
	wire _w22991_ ;
	wire _w22990_ ;
	wire _w22989_ ;
	wire _w22988_ ;
	wire _w22987_ ;
	wire _w22986_ ;
	wire _w22985_ ;
	wire _w22984_ ;
	wire _w22983_ ;
	wire _w22982_ ;
	wire _w22981_ ;
	wire _w22980_ ;
	wire _w22979_ ;
	wire _w22978_ ;
	wire _w22977_ ;
	wire _w22976_ ;
	wire _w22975_ ;
	wire _w22974_ ;
	wire _w22973_ ;
	wire _w22972_ ;
	wire _w22971_ ;
	wire _w22970_ ;
	wire _w22969_ ;
	wire _w22968_ ;
	wire _w22967_ ;
	wire _w22966_ ;
	wire _w22965_ ;
	wire _w22964_ ;
	wire _w22963_ ;
	wire _w22962_ ;
	wire _w22961_ ;
	wire _w22960_ ;
	wire _w22959_ ;
	wire _w22958_ ;
	wire _w22957_ ;
	wire _w22956_ ;
	wire _w22955_ ;
	wire _w22954_ ;
	wire _w22953_ ;
	wire _w22952_ ;
	wire _w22951_ ;
	wire _w22950_ ;
	wire _w22949_ ;
	wire _w22948_ ;
	wire _w22947_ ;
	wire _w22946_ ;
	wire _w22945_ ;
	wire _w22944_ ;
	wire _w22943_ ;
	wire _w22942_ ;
	wire _w22941_ ;
	wire _w22940_ ;
	wire _w22939_ ;
	wire _w22938_ ;
	wire _w22937_ ;
	wire _w22936_ ;
	wire _w22935_ ;
	wire _w22934_ ;
	wire _w22933_ ;
	wire _w22932_ ;
	wire _w22931_ ;
	wire _w22930_ ;
	wire _w22929_ ;
	wire _w22928_ ;
	wire _w22927_ ;
	wire _w22926_ ;
	wire _w22925_ ;
	wire _w22924_ ;
	wire _w22923_ ;
	wire _w22922_ ;
	wire _w22921_ ;
	wire _w22920_ ;
	wire _w22919_ ;
	wire _w22918_ ;
	wire _w22917_ ;
	wire _w22916_ ;
	wire _w22915_ ;
	wire _w22914_ ;
	wire _w22913_ ;
	wire _w22912_ ;
	wire _w22911_ ;
	wire _w22910_ ;
	wire _w22909_ ;
	wire _w22908_ ;
	wire _w22907_ ;
	wire _w22906_ ;
	wire _w22905_ ;
	wire _w22904_ ;
	wire _w22903_ ;
	wire _w22902_ ;
	wire _w22901_ ;
	wire _w22900_ ;
	wire _w22899_ ;
	wire _w22898_ ;
	wire _w22897_ ;
	wire _w22896_ ;
	wire _w22895_ ;
	wire _w22894_ ;
	wire _w22893_ ;
	wire _w22892_ ;
	wire _w22891_ ;
	wire _w22890_ ;
	wire _w22889_ ;
	wire _w22888_ ;
	wire _w22887_ ;
	wire _w22886_ ;
	wire _w22885_ ;
	wire _w22884_ ;
	wire _w22883_ ;
	wire _w22882_ ;
	wire _w22881_ ;
	wire _w22880_ ;
	wire _w22879_ ;
	wire _w22878_ ;
	wire _w22877_ ;
	wire _w22876_ ;
	wire _w22875_ ;
	wire _w22874_ ;
	wire _w22873_ ;
	wire _w22872_ ;
	wire _w22871_ ;
	wire _w22870_ ;
	wire _w22869_ ;
	wire _w22868_ ;
	wire _w22867_ ;
	wire _w22866_ ;
	wire _w22865_ ;
	wire _w22864_ ;
	wire _w22863_ ;
	wire _w22862_ ;
	wire _w22861_ ;
	wire _w22860_ ;
	wire _w22859_ ;
	wire _w22858_ ;
	wire _w22857_ ;
	wire _w22856_ ;
	wire _w22855_ ;
	wire _w22854_ ;
	wire _w22853_ ;
	wire _w22852_ ;
	wire _w22851_ ;
	wire _w22850_ ;
	wire _w22849_ ;
	wire _w22848_ ;
	wire _w22847_ ;
	wire _w22846_ ;
	wire _w22845_ ;
	wire _w22844_ ;
	wire _w22843_ ;
	wire _w22842_ ;
	wire _w22841_ ;
	wire _w22840_ ;
	wire _w22839_ ;
	wire _w22838_ ;
	wire _w22837_ ;
	wire _w22836_ ;
	wire _w22835_ ;
	wire _w22834_ ;
	wire _w22833_ ;
	wire _w22832_ ;
	wire _w22831_ ;
	wire _w22830_ ;
	wire _w22829_ ;
	wire _w22828_ ;
	wire _w22827_ ;
	wire _w22826_ ;
	wire _w22825_ ;
	wire _w22824_ ;
	wire _w22823_ ;
	wire _w22822_ ;
	wire _w22821_ ;
	wire _w22820_ ;
	wire _w22819_ ;
	wire _w22818_ ;
	wire _w22817_ ;
	wire _w22816_ ;
	wire _w22815_ ;
	wire _w22814_ ;
	wire _w22813_ ;
	wire _w22812_ ;
	wire _w22811_ ;
	wire _w22810_ ;
	wire _w22809_ ;
	wire _w22808_ ;
	wire _w22807_ ;
	wire _w22806_ ;
	wire _w22805_ ;
	wire _w22804_ ;
	wire _w22803_ ;
	wire _w22802_ ;
	wire _w22801_ ;
	wire _w22800_ ;
	wire _w22799_ ;
	wire _w22798_ ;
	wire _w22797_ ;
	wire _w22796_ ;
	wire _w22795_ ;
	wire _w22794_ ;
	wire _w22793_ ;
	wire _w22792_ ;
	wire _w22791_ ;
	wire _w22790_ ;
	wire _w22789_ ;
	wire _w22788_ ;
	wire _w22787_ ;
	wire _w22786_ ;
	wire _w22785_ ;
	wire _w22784_ ;
	wire _w22783_ ;
	wire _w22782_ ;
	wire _w22781_ ;
	wire _w22780_ ;
	wire _w22779_ ;
	wire _w22778_ ;
	wire _w22777_ ;
	wire _w22776_ ;
	wire _w22775_ ;
	wire _w22774_ ;
	wire _w22773_ ;
	wire _w22772_ ;
	wire _w22771_ ;
	wire _w22770_ ;
	wire _w22769_ ;
	wire _w22768_ ;
	wire _w22767_ ;
	wire _w22766_ ;
	wire _w22765_ ;
	wire _w22764_ ;
	wire _w22763_ ;
	wire _w22762_ ;
	wire _w22761_ ;
	wire _w22760_ ;
	wire _w22759_ ;
	wire _w22758_ ;
	wire _w22757_ ;
	wire _w22756_ ;
	wire _w22755_ ;
	wire _w22754_ ;
	wire _w22753_ ;
	wire _w22752_ ;
	wire _w22751_ ;
	wire _w22750_ ;
	wire _w22749_ ;
	wire _w22748_ ;
	wire _w22747_ ;
	wire _w22746_ ;
	wire _w22745_ ;
	wire _w22744_ ;
	wire _w22743_ ;
	wire _w22742_ ;
	wire _w22741_ ;
	wire _w22740_ ;
	wire _w22739_ ;
	wire _w22738_ ;
	wire _w22737_ ;
	wire _w22736_ ;
	wire _w22735_ ;
	wire _w22734_ ;
	wire _w22733_ ;
	wire _w22732_ ;
	wire _w22731_ ;
	wire _w22730_ ;
	wire _w22729_ ;
	wire _w22728_ ;
	wire _w22727_ ;
	wire _w22726_ ;
	wire _w22725_ ;
	wire _w22724_ ;
	wire _w22723_ ;
	wire _w22722_ ;
	wire _w22721_ ;
	wire _w22720_ ;
	wire _w22719_ ;
	wire _w22718_ ;
	wire _w22717_ ;
	wire _w22716_ ;
	wire _w22715_ ;
	wire _w22714_ ;
	wire _w22713_ ;
	wire _w22712_ ;
	wire _w22711_ ;
	wire _w22710_ ;
	wire _w22709_ ;
	wire _w22708_ ;
	wire _w22707_ ;
	wire _w22706_ ;
	wire _w22705_ ;
	wire _w22704_ ;
	wire _w22703_ ;
	wire _w22702_ ;
	wire _w22701_ ;
	wire _w22700_ ;
	wire _w22699_ ;
	wire _w22698_ ;
	wire _w22697_ ;
	wire _w22696_ ;
	wire _w22695_ ;
	wire _w22694_ ;
	wire _w22693_ ;
	wire _w22692_ ;
	wire _w22691_ ;
	wire _w22690_ ;
	wire _w22689_ ;
	wire _w22688_ ;
	wire _w22687_ ;
	wire _w22686_ ;
	wire _w22685_ ;
	wire _w22684_ ;
	wire _w22683_ ;
	wire _w22682_ ;
	wire _w22681_ ;
	wire _w22680_ ;
	wire _w22679_ ;
	wire _w22678_ ;
	wire _w22677_ ;
	wire _w22676_ ;
	wire _w22675_ ;
	wire _w22674_ ;
	wire _w22673_ ;
	wire _w22672_ ;
	wire _w22671_ ;
	wire _w22670_ ;
	wire _w22669_ ;
	wire _w22668_ ;
	wire _w22667_ ;
	wire _w22666_ ;
	wire _w22665_ ;
	wire _w22664_ ;
	wire _w22663_ ;
	wire _w22662_ ;
	wire _w22661_ ;
	wire _w22660_ ;
	wire _w22659_ ;
	wire _w22658_ ;
	wire _w22657_ ;
	wire _w22656_ ;
	wire _w22655_ ;
	wire _w22654_ ;
	wire _w12173_ ;
	wire _w12172_ ;
	wire _w12171_ ;
	wire _w12170_ ;
	wire _w12169_ ;
	wire _w12168_ ;
	wire _w12167_ ;
	wire _w12166_ ;
	wire _w12165_ ;
	wire _w12164_ ;
	wire _w12163_ ;
	wire _w12162_ ;
	wire _w12161_ ;
	wire _w12160_ ;
	wire _w12159_ ;
	wire _w12158_ ;
	wire _w12157_ ;
	wire _w12156_ ;
	wire _w12155_ ;
	wire _w12154_ ;
	wire _w12153_ ;
	wire _w12152_ ;
	wire _w12151_ ;
	wire _w12150_ ;
	wire _w12149_ ;
	wire _w12148_ ;
	wire _w12147_ ;
	wire _w12146_ ;
	wire _w12145_ ;
	wire _w12144_ ;
	wire _w12143_ ;
	wire _w12142_ ;
	wire _w12141_ ;
	wire _w12140_ ;
	wire _w12139_ ;
	wire _w12138_ ;
	wire _w12137_ ;
	wire _w12136_ ;
	wire _w12135_ ;
	wire _w12134_ ;
	wire _w12133_ ;
	wire _w12132_ ;
	wire _w12131_ ;
	wire _w12130_ ;
	wire _w12129_ ;
	wire _w12128_ ;
	wire _w12127_ ;
	wire _w12126_ ;
	wire _w12125_ ;
	wire _w12124_ ;
	wire _w12123_ ;
	wire _w12122_ ;
	wire _w12121_ ;
	wire _w12120_ ;
	wire _w12119_ ;
	wire _w12118_ ;
	wire _w12117_ ;
	wire _w12116_ ;
	wire _w12115_ ;
	wire _w12114_ ;
	wire _w12113_ ;
	wire _w12112_ ;
	wire _w12111_ ;
	wire _w12110_ ;
	wire _w12109_ ;
	wire _w12108_ ;
	wire _w12107_ ;
	wire _w12106_ ;
	wire _w12105_ ;
	wire _w12104_ ;
	wire _w12103_ ;
	wire _w12102_ ;
	wire _w12101_ ;
	wire _w12100_ ;
	wire _w12099_ ;
	wire _w12098_ ;
	wire _w12097_ ;
	wire _w12096_ ;
	wire _w12095_ ;
	wire _w12094_ ;
	wire _w12093_ ;
	wire _w12092_ ;
	wire _w12091_ ;
	wire _w12090_ ;
	wire _w12089_ ;
	wire _w12088_ ;
	wire _w12087_ ;
	wire _w12086_ ;
	wire _w12085_ ;
	wire _w12084_ ;
	wire _w12083_ ;
	wire _w12082_ ;
	wire _w12081_ ;
	wire _w12080_ ;
	wire _w12079_ ;
	wire _w12078_ ;
	wire _w12077_ ;
	wire _w12076_ ;
	wire _w12075_ ;
	wire _w12074_ ;
	wire _w12073_ ;
	wire _w12072_ ;
	wire _w12071_ ;
	wire _w12070_ ;
	wire _w12069_ ;
	wire _w12068_ ;
	wire _w12067_ ;
	wire _w12066_ ;
	wire _w12065_ ;
	wire _w12064_ ;
	wire _w12063_ ;
	wire _w12062_ ;
	wire _w12061_ ;
	wire _w12060_ ;
	wire _w12059_ ;
	wire _w12058_ ;
	wire _w12057_ ;
	wire _w12056_ ;
	wire _w12055_ ;
	wire _w12054_ ;
	wire _w12053_ ;
	wire _w12052_ ;
	wire _w12051_ ;
	wire _w12050_ ;
	wire _w12049_ ;
	wire _w12048_ ;
	wire _w12047_ ;
	wire _w12046_ ;
	wire _w12045_ ;
	wire _w12044_ ;
	wire _w12043_ ;
	wire _w12042_ ;
	wire _w12041_ ;
	wire _w12040_ ;
	wire _w12039_ ;
	wire _w12038_ ;
	wire _w12037_ ;
	wire _w12036_ ;
	wire _w12035_ ;
	wire _w12034_ ;
	wire _w12033_ ;
	wire _w12032_ ;
	wire _w12031_ ;
	wire _w12030_ ;
	wire _w12029_ ;
	wire _w12028_ ;
	wire _w12027_ ;
	wire _w12026_ ;
	wire _w12025_ ;
	wire _w12024_ ;
	wire _w12023_ ;
	wire _w12022_ ;
	wire _w12021_ ;
	wire _w12020_ ;
	wire _w12019_ ;
	wire _w12018_ ;
	wire _w12017_ ;
	wire _w12016_ ;
	wire _w12015_ ;
	wire _w12014_ ;
	wire _w12013_ ;
	wire _w12012_ ;
	wire _w12011_ ;
	wire _w12010_ ;
	wire _w12009_ ;
	wire _w12008_ ;
	wire _w12007_ ;
	wire _w12006_ ;
	wire _w12005_ ;
	wire _w12004_ ;
	wire _w12003_ ;
	wire _w12002_ ;
	wire _w12001_ ;
	wire _w12000_ ;
	wire _w11999_ ;
	wire _w11998_ ;
	wire _w11997_ ;
	wire _w11996_ ;
	wire _w11995_ ;
	wire _w11994_ ;
	wire _w11993_ ;
	wire _w11992_ ;
	wire _w11991_ ;
	wire _w11990_ ;
	wire _w11989_ ;
	wire _w11988_ ;
	wire _w11987_ ;
	wire _w11986_ ;
	wire _w11985_ ;
	wire _w11984_ ;
	wire _w11983_ ;
	wire _w11982_ ;
	wire _w11981_ ;
	wire _w11980_ ;
	wire _w11979_ ;
	wire _w11978_ ;
	wire _w11977_ ;
	wire _w11976_ ;
	wire _w11975_ ;
	wire _w11974_ ;
	wire _w11973_ ;
	wire _w11972_ ;
	wire _w11971_ ;
	wire _w11970_ ;
	wire _w11969_ ;
	wire _w11968_ ;
	wire _w11967_ ;
	wire _w11966_ ;
	wire _w11965_ ;
	wire _w11964_ ;
	wire _w11963_ ;
	wire _w11962_ ;
	wire _w11961_ ;
	wire _w11960_ ;
	wire _w11959_ ;
	wire _w11958_ ;
	wire _w11957_ ;
	wire _w11956_ ;
	wire _w11955_ ;
	wire _w11954_ ;
	wire _w11953_ ;
	wire _w11952_ ;
	wire _w11951_ ;
	wire _w11950_ ;
	wire _w11949_ ;
	wire _w11948_ ;
	wire _w11947_ ;
	wire _w11946_ ;
	wire _w11945_ ;
	wire _w11944_ ;
	wire _w11943_ ;
	wire _w11942_ ;
	wire _w11941_ ;
	wire _w11940_ ;
	wire _w11939_ ;
	wire _w11938_ ;
	wire _w11937_ ;
	wire _w11936_ ;
	wire _w11935_ ;
	wire _w11934_ ;
	wire _w11933_ ;
	wire _w11932_ ;
	wire _w11931_ ;
	wire _w11930_ ;
	wire _w11929_ ;
	wire _w11928_ ;
	wire _w11927_ ;
	wire _w11926_ ;
	wire _w11925_ ;
	wire _w11924_ ;
	wire _w11923_ ;
	wire _w11922_ ;
	wire _w11921_ ;
	wire _w11920_ ;
	wire _w11919_ ;
	wire _w11918_ ;
	wire _w11917_ ;
	wire _w11916_ ;
	wire _w11915_ ;
	wire _w11914_ ;
	wire _w11913_ ;
	wire _w11912_ ;
	wire _w11911_ ;
	wire _w11910_ ;
	wire _w11909_ ;
	wire _w11908_ ;
	wire _w11907_ ;
	wire _w11906_ ;
	wire _w11905_ ;
	wire _w11904_ ;
	wire _w11903_ ;
	wire _w11902_ ;
	wire _w11901_ ;
	wire _w11900_ ;
	wire _w11899_ ;
	wire _w11898_ ;
	wire _w11897_ ;
	wire _w11896_ ;
	wire _w11895_ ;
	wire _w11894_ ;
	wire _w11893_ ;
	wire _w11892_ ;
	wire _w11891_ ;
	wire _w11890_ ;
	wire _w11889_ ;
	wire _w11888_ ;
	wire _w11887_ ;
	wire _w11886_ ;
	wire _w11885_ ;
	wire _w11884_ ;
	wire _w11883_ ;
	wire _w11882_ ;
	wire _w11881_ ;
	wire _w11880_ ;
	wire _w11879_ ;
	wire _w11878_ ;
	wire _w11877_ ;
	wire _w11876_ ;
	wire _w11875_ ;
	wire _w11874_ ;
	wire _w11873_ ;
	wire _w11872_ ;
	wire _w11871_ ;
	wire _w11870_ ;
	wire _w11869_ ;
	wire _w11868_ ;
	wire _w11867_ ;
	wire _w11866_ ;
	wire _w11865_ ;
	wire _w11864_ ;
	wire _w11863_ ;
	wire _w11862_ ;
	wire _w11861_ ;
	wire _w11860_ ;
	wire _w11859_ ;
	wire _w11858_ ;
	wire _w11857_ ;
	wire _w11856_ ;
	wire _w11855_ ;
	wire _w11854_ ;
	wire _w11853_ ;
	wire _w11852_ ;
	wire _w11851_ ;
	wire _w11850_ ;
	wire _w11849_ ;
	wire _w11848_ ;
	wire _w11847_ ;
	wire _w11846_ ;
	wire _w11845_ ;
	wire _w11844_ ;
	wire _w11843_ ;
	wire _w11842_ ;
	wire _w11841_ ;
	wire _w11840_ ;
	wire _w11839_ ;
	wire _w11838_ ;
	wire _w11837_ ;
	wire _w11836_ ;
	wire _w11835_ ;
	wire _w11834_ ;
	wire _w11833_ ;
	wire _w11832_ ;
	wire _w11831_ ;
	wire _w11830_ ;
	wire _w11829_ ;
	wire _w11828_ ;
	wire _w11827_ ;
	wire _w11826_ ;
	wire _w11825_ ;
	wire _w11824_ ;
	wire _w11823_ ;
	wire _w11822_ ;
	wire _w11821_ ;
	wire _w11820_ ;
	wire _w11819_ ;
	wire _w11818_ ;
	wire _w11817_ ;
	wire _w11816_ ;
	wire _w11815_ ;
	wire _w11814_ ;
	wire _w11813_ ;
	wire _w11812_ ;
	wire _w11811_ ;
	wire _w11810_ ;
	wire _w11809_ ;
	wire _w11808_ ;
	wire _w11807_ ;
	wire _w11806_ ;
	wire _w11805_ ;
	wire _w11804_ ;
	wire _w11803_ ;
	wire _w11802_ ;
	wire _w11801_ ;
	wire _w11800_ ;
	wire _w11799_ ;
	wire _w11798_ ;
	wire _w11797_ ;
	wire _w11796_ ;
	wire _w11795_ ;
	wire _w11794_ ;
	wire _w11793_ ;
	wire _w11792_ ;
	wire _w11791_ ;
	wire _w11790_ ;
	wire _w11789_ ;
	wire _w11788_ ;
	wire _w11787_ ;
	wire _w11786_ ;
	wire _w11785_ ;
	wire _w11784_ ;
	wire _w11783_ ;
	wire _w11782_ ;
	wire _w11781_ ;
	wire _w11780_ ;
	wire _w11779_ ;
	wire _w11778_ ;
	wire _w11777_ ;
	wire _w11776_ ;
	wire _w11775_ ;
	wire _w11774_ ;
	wire _w11773_ ;
	wire _w11772_ ;
	wire _w11771_ ;
	wire _w11770_ ;
	wire _w11769_ ;
	wire _w11768_ ;
	wire _w11767_ ;
	wire _w11766_ ;
	wire _w11765_ ;
	wire _w11764_ ;
	wire _w11763_ ;
	wire _w11762_ ;
	wire _w11761_ ;
	wire _w11760_ ;
	wire _w11759_ ;
	wire _w11758_ ;
	wire _w11757_ ;
	wire _w11756_ ;
	wire _w11755_ ;
	wire _w11754_ ;
	wire _w11753_ ;
	wire _w11752_ ;
	wire _w11751_ ;
	wire _w11750_ ;
	wire _w11749_ ;
	wire _w11748_ ;
	wire _w11747_ ;
	wire _w11746_ ;
	wire _w11745_ ;
	wire _w11744_ ;
	wire _w11743_ ;
	wire _w11742_ ;
	wire _w11741_ ;
	wire _w11740_ ;
	wire _w11739_ ;
	wire _w11738_ ;
	wire _w11737_ ;
	wire _w11736_ ;
	wire _w11735_ ;
	wire _w11734_ ;
	wire _w11733_ ;
	wire _w11732_ ;
	wire _w11731_ ;
	wire _w11730_ ;
	wire _w11729_ ;
	wire _w11728_ ;
	wire _w11727_ ;
	wire _w11726_ ;
	wire _w11725_ ;
	wire _w11724_ ;
	wire _w11723_ ;
	wire _w11722_ ;
	wire _w11721_ ;
	wire _w11720_ ;
	wire _w11719_ ;
	wire _w11718_ ;
	wire _w11717_ ;
	wire _w11716_ ;
	wire _w11715_ ;
	wire _w11714_ ;
	wire _w11713_ ;
	wire _w11712_ ;
	wire _w11711_ ;
	wire _w11710_ ;
	wire _w11709_ ;
	wire _w11708_ ;
	wire _w11707_ ;
	wire _w11706_ ;
	wire _w11705_ ;
	wire _w11704_ ;
	wire _w11703_ ;
	wire _w11702_ ;
	wire _w11701_ ;
	wire _w11700_ ;
	wire _w11699_ ;
	wire _w11698_ ;
	wire _w11697_ ;
	wire _w11696_ ;
	wire _w11695_ ;
	wire _w11694_ ;
	wire _w11693_ ;
	wire _w11692_ ;
	wire _w11691_ ;
	wire _w11690_ ;
	wire _w11689_ ;
	wire _w11688_ ;
	wire _w11687_ ;
	wire _w11686_ ;
	wire _w11685_ ;
	wire _w11684_ ;
	wire _w11683_ ;
	wire _w11682_ ;
	wire _w11681_ ;
	wire _w11680_ ;
	wire _w11679_ ;
	wire _w11678_ ;
	wire _w11677_ ;
	wire _w11676_ ;
	wire _w11675_ ;
	wire _w11674_ ;
	wire _w11673_ ;
	wire _w11672_ ;
	wire _w11671_ ;
	wire _w11670_ ;
	wire _w11669_ ;
	wire _w11668_ ;
	wire _w11667_ ;
	wire _w11666_ ;
	wire _w11665_ ;
	wire _w11664_ ;
	wire _w11663_ ;
	wire _w11662_ ;
	wire _w11661_ ;
	wire _w11660_ ;
	wire _w11659_ ;
	wire _w11658_ ;
	wire _w11657_ ;
	wire _w11656_ ;
	wire _w11655_ ;
	wire _w11654_ ;
	wire _w11653_ ;
	wire _w11652_ ;
	wire _w11651_ ;
	wire _w11650_ ;
	wire _w11649_ ;
	wire _w11648_ ;
	wire _w11647_ ;
	wire _w11646_ ;
	wire _w11645_ ;
	wire _w11644_ ;
	wire _w11643_ ;
	wire _w11642_ ;
	wire _w11641_ ;
	wire _w11640_ ;
	wire _w11639_ ;
	wire _w11638_ ;
	wire _w11637_ ;
	wire _w11636_ ;
	wire _w11635_ ;
	wire _w11634_ ;
	wire _w11633_ ;
	wire _w11632_ ;
	wire _w11631_ ;
	wire _w11630_ ;
	wire _w11629_ ;
	wire _w11628_ ;
	wire _w11627_ ;
	wire _w11626_ ;
	wire _w11625_ ;
	wire _w11624_ ;
	wire _w11623_ ;
	wire _w11622_ ;
	wire _w11621_ ;
	wire _w11620_ ;
	wire _w11619_ ;
	wire _w11618_ ;
	wire _w11617_ ;
	wire _w11616_ ;
	wire _w11615_ ;
	wire _w11614_ ;
	wire _w11613_ ;
	wire _w11612_ ;
	wire _w11611_ ;
	wire _w11610_ ;
	wire _w11609_ ;
	wire _w11608_ ;
	wire _w11607_ ;
	wire _w11606_ ;
	wire _w11605_ ;
	wire _w11604_ ;
	wire _w11603_ ;
	wire _w11602_ ;
	wire _w11601_ ;
	wire _w11600_ ;
	wire _w11599_ ;
	wire _w11598_ ;
	wire _w11597_ ;
	wire _w11596_ ;
	wire _w11595_ ;
	wire _w11594_ ;
	wire _w11593_ ;
	wire _w11592_ ;
	wire _w11591_ ;
	wire _w11590_ ;
	wire _w11589_ ;
	wire _w11588_ ;
	wire _w11587_ ;
	wire _w11586_ ;
	wire _w11585_ ;
	wire _w11584_ ;
	wire _w11583_ ;
	wire _w11582_ ;
	wire _w11581_ ;
	wire _w11580_ ;
	wire _w11579_ ;
	wire _w11578_ ;
	wire _w11577_ ;
	wire _w11576_ ;
	wire _w11575_ ;
	wire _w11574_ ;
	wire _w11573_ ;
	wire _w11572_ ;
	wire _w11571_ ;
	wire _w11570_ ;
	wire _w11569_ ;
	wire _w11568_ ;
	wire _w11567_ ;
	wire _w11566_ ;
	wire _w11565_ ;
	wire _w11564_ ;
	wire _w11563_ ;
	wire _w11562_ ;
	wire _w11561_ ;
	wire _w11560_ ;
	wire _w11559_ ;
	wire _w11558_ ;
	wire _w11557_ ;
	wire _w11556_ ;
	wire _w11555_ ;
	wire _w11554_ ;
	wire _w11553_ ;
	wire _w11552_ ;
	wire _w11551_ ;
	wire _w11550_ ;
	wire _w11549_ ;
	wire _w11548_ ;
	wire _w11547_ ;
	wire _w11546_ ;
	wire _w11545_ ;
	wire _w11544_ ;
	wire _w11543_ ;
	wire _w11542_ ;
	wire _w11541_ ;
	wire _w11540_ ;
	wire _w11539_ ;
	wire _w11538_ ;
	wire _w11537_ ;
	wire _w11536_ ;
	wire _w11535_ ;
	wire _w11534_ ;
	wire _w11533_ ;
	wire _w11532_ ;
	wire _w11531_ ;
	wire _w11530_ ;
	wire _w11529_ ;
	wire _w11528_ ;
	wire _w11527_ ;
	wire _w11526_ ;
	wire _w11525_ ;
	wire _w11524_ ;
	wire _w11523_ ;
	wire _w11522_ ;
	wire _w11521_ ;
	wire _w11520_ ;
	wire _w11519_ ;
	wire _w11518_ ;
	wire _w11517_ ;
	wire _w11516_ ;
	wire _w11515_ ;
	wire _w11514_ ;
	wire _w11513_ ;
	wire _w11512_ ;
	wire _w11511_ ;
	wire _w11510_ ;
	wire _w11509_ ;
	wire _w11508_ ;
	wire _w11507_ ;
	wire _w11506_ ;
	wire _w11505_ ;
	wire _w11504_ ;
	wire _w11503_ ;
	wire _w11502_ ;
	wire _w11501_ ;
	wire _w11500_ ;
	wire _w11499_ ;
	wire _w11498_ ;
	wire _w11497_ ;
	wire _w11496_ ;
	wire _w11495_ ;
	wire _w11494_ ;
	wire _w11493_ ;
	wire _w11492_ ;
	wire _w11491_ ;
	wire _w11490_ ;
	wire _w11489_ ;
	wire _w11488_ ;
	wire _w11487_ ;
	wire _w11486_ ;
	wire _w11485_ ;
	wire _w11484_ ;
	wire _w11483_ ;
	wire _w11482_ ;
	wire _w11481_ ;
	wire _w11480_ ;
	wire _w11479_ ;
	wire _w11478_ ;
	wire _w11477_ ;
	wire _w11476_ ;
	wire _w11475_ ;
	wire _w11474_ ;
	wire _w11473_ ;
	wire _w11472_ ;
	wire _w11471_ ;
	wire _w11470_ ;
	wire _w11469_ ;
	wire _w11468_ ;
	wire _w11467_ ;
	wire _w11466_ ;
	wire _w11465_ ;
	wire _w11464_ ;
	wire _w11463_ ;
	wire _w11462_ ;
	wire _w11461_ ;
	wire _w11460_ ;
	wire _w11459_ ;
	wire _w11458_ ;
	wire _w11457_ ;
	wire _w11456_ ;
	wire _w11455_ ;
	wire _w11454_ ;
	wire _w11453_ ;
	wire _w11452_ ;
	wire _w11451_ ;
	wire _w11450_ ;
	wire _w11449_ ;
	wire _w11448_ ;
	wire _w11447_ ;
	wire _w11446_ ;
	wire _w11445_ ;
	wire _w11444_ ;
	wire _w11443_ ;
	wire _w11442_ ;
	wire _w11441_ ;
	wire _w11440_ ;
	wire _w11439_ ;
	wire _w11438_ ;
	wire _w11437_ ;
	wire _w11436_ ;
	wire _w11435_ ;
	wire _w11434_ ;
	wire _w11433_ ;
	wire _w11432_ ;
	wire _w11431_ ;
	wire _w11430_ ;
	wire _w11429_ ;
	wire _w11428_ ;
	wire _w11427_ ;
	wire _w11426_ ;
	wire _w11425_ ;
	wire _w11424_ ;
	wire _w11423_ ;
	wire _w11422_ ;
	wire _w11421_ ;
	wire _w11420_ ;
	wire _w11419_ ;
	wire _w11418_ ;
	wire _w11417_ ;
	wire _w11416_ ;
	wire _w11415_ ;
	wire _w11414_ ;
	wire _w11413_ ;
	wire _w11412_ ;
	wire _w11411_ ;
	wire _w11410_ ;
	wire _w11409_ ;
	wire _w11408_ ;
	wire _w11407_ ;
	wire _w11406_ ;
	wire _w11405_ ;
	wire _w11404_ ;
	wire _w11403_ ;
	wire _w11402_ ;
	wire _w11401_ ;
	wire _w11400_ ;
	wire _w11399_ ;
	wire _w11398_ ;
	wire _w11397_ ;
	wire _w11396_ ;
	wire _w11395_ ;
	wire _w11394_ ;
	wire _w11393_ ;
	wire _w11392_ ;
	wire _w11391_ ;
	wire _w11390_ ;
	wire _w11389_ ;
	wire _w11388_ ;
	wire _w11387_ ;
	wire _w11386_ ;
	wire _w11385_ ;
	wire _w11384_ ;
	wire _w11383_ ;
	wire _w11382_ ;
	wire _w11381_ ;
	wire _w11380_ ;
	wire _w11379_ ;
	wire _w11378_ ;
	wire _w11377_ ;
	wire _w11376_ ;
	wire _w11375_ ;
	wire _w11374_ ;
	wire _w11373_ ;
	wire _w11372_ ;
	wire _w11371_ ;
	wire _w11370_ ;
	wire _w11369_ ;
	wire _w11368_ ;
	wire _w11367_ ;
	wire _w11366_ ;
	wire _w11365_ ;
	wire _w11364_ ;
	wire _w11363_ ;
	wire _w11362_ ;
	wire _w11361_ ;
	wire _w11360_ ;
	wire _w11359_ ;
	wire _w11358_ ;
	wire _w11357_ ;
	wire _w11356_ ;
	wire _w11355_ ;
	wire _w11354_ ;
	wire _w11353_ ;
	wire _w11352_ ;
	wire _w11351_ ;
	wire _w11350_ ;
	wire _w11349_ ;
	wire _w11348_ ;
	wire _w11347_ ;
	wire _w11346_ ;
	wire _w11345_ ;
	wire _w11344_ ;
	wire _w11343_ ;
	wire _w11342_ ;
	wire _w11341_ ;
	wire _w11340_ ;
	wire _w11339_ ;
	wire _w11338_ ;
	wire _w11337_ ;
	wire _w11336_ ;
	wire _w11335_ ;
	wire _w11334_ ;
	wire _w11333_ ;
	wire _w11332_ ;
	wire _w11331_ ;
	wire _w11330_ ;
	wire _w11329_ ;
	wire _w11328_ ;
	wire _w11327_ ;
	wire _w11326_ ;
	wire _w11325_ ;
	wire _w11324_ ;
	wire _w11323_ ;
	wire _w11322_ ;
	wire _w11321_ ;
	wire _w11320_ ;
	wire _w11319_ ;
	wire _w11318_ ;
	wire _w11317_ ;
	wire _w11316_ ;
	wire _w11315_ ;
	wire _w11314_ ;
	wire _w11313_ ;
	wire _w11312_ ;
	wire _w11311_ ;
	wire _w11310_ ;
	wire _w11309_ ;
	wire _w11308_ ;
	wire _w11307_ ;
	wire _w11306_ ;
	wire _w11305_ ;
	wire _w11304_ ;
	wire _w11303_ ;
	wire _w11302_ ;
	wire _w11301_ ;
	wire _w11300_ ;
	wire _w11299_ ;
	wire _w11298_ ;
	wire _w11297_ ;
	wire _w11296_ ;
	wire _w11295_ ;
	wire _w11294_ ;
	wire _w11293_ ;
	wire _w11292_ ;
	wire _w11291_ ;
	wire _w11290_ ;
	wire _w11289_ ;
	wire _w11288_ ;
	wire _w11287_ ;
	wire _w11286_ ;
	wire _w11285_ ;
	wire _w11284_ ;
	wire _w11283_ ;
	wire _w11282_ ;
	wire _w11281_ ;
	wire _w11280_ ;
	wire _w11279_ ;
	wire _w11278_ ;
	wire _w11277_ ;
	wire _w11276_ ;
	wire _w11275_ ;
	wire _w11274_ ;
	wire _w11273_ ;
	wire _w11272_ ;
	wire _w11271_ ;
	wire _w11270_ ;
	wire _w11269_ ;
	wire _w11268_ ;
	wire _w11267_ ;
	wire _w11266_ ;
	wire _w11265_ ;
	wire _w11264_ ;
	wire _w11263_ ;
	wire _w11262_ ;
	wire _w11261_ ;
	wire _w11260_ ;
	wire _w11259_ ;
	wire _w11258_ ;
	wire _w11257_ ;
	wire _w11256_ ;
	wire _w11255_ ;
	wire _w11254_ ;
	wire _w11253_ ;
	wire _w11252_ ;
	wire _w11251_ ;
	wire _w11250_ ;
	wire _w11249_ ;
	wire _w11248_ ;
	wire _w11247_ ;
	wire _w11246_ ;
	wire _w11245_ ;
	wire _w11244_ ;
	wire _w11243_ ;
	wire _w11242_ ;
	wire _w11241_ ;
	wire _w11240_ ;
	wire _w11239_ ;
	wire _w11238_ ;
	wire _w11237_ ;
	wire _w11236_ ;
	wire _w11235_ ;
	wire _w11234_ ;
	wire _w11233_ ;
	wire _w11232_ ;
	wire _w11231_ ;
	wire _w11230_ ;
	wire _w11229_ ;
	wire _w11228_ ;
	wire _w11227_ ;
	wire _w11226_ ;
	wire _w11225_ ;
	wire _w11224_ ;
	wire _w11223_ ;
	wire _w11222_ ;
	wire _w11221_ ;
	wire _w11220_ ;
	wire _w11219_ ;
	wire _w11218_ ;
	wire _w11217_ ;
	wire _w11216_ ;
	wire _w11215_ ;
	wire _w11214_ ;
	wire _w11213_ ;
	wire _w11212_ ;
	wire _w11211_ ;
	wire _w11210_ ;
	wire _w11209_ ;
	wire _w11208_ ;
	wire _w11207_ ;
	wire _w11206_ ;
	wire _w11205_ ;
	wire _w11204_ ;
	wire _w11203_ ;
	wire _w11202_ ;
	wire _w11201_ ;
	wire _w11200_ ;
	wire _w11199_ ;
	wire _w11198_ ;
	wire _w11197_ ;
	wire _w11196_ ;
	wire _w11195_ ;
	wire _w11194_ ;
	wire _w11193_ ;
	wire _w11192_ ;
	wire _w11191_ ;
	wire _w11190_ ;
	wire _w11189_ ;
	wire _w11188_ ;
	wire _w11187_ ;
	wire _w11186_ ;
	wire _w11185_ ;
	wire _w11184_ ;
	wire _w11183_ ;
	wire _w11182_ ;
	wire _w11181_ ;
	wire _w11180_ ;
	wire _w11179_ ;
	wire _w11178_ ;
	wire _w11177_ ;
	wire _w11176_ ;
	wire _w11175_ ;
	wire _w11174_ ;
	wire _w11173_ ;
	wire _w11172_ ;
	wire _w11171_ ;
	wire _w11170_ ;
	wire _w11169_ ;
	wire _w11168_ ;
	wire _w11167_ ;
	wire _w11166_ ;
	wire _w11165_ ;
	wire _w11164_ ;
	wire _w11163_ ;
	wire _w11162_ ;
	wire _w11161_ ;
	wire _w11160_ ;
	wire _w11159_ ;
	wire _w11158_ ;
	wire _w11157_ ;
	wire _w11156_ ;
	wire _w11155_ ;
	wire _w11154_ ;
	wire _w11153_ ;
	wire _w11152_ ;
	wire _w11151_ ;
	wire _w11150_ ;
	wire _w11149_ ;
	wire _w11148_ ;
	wire _w11147_ ;
	wire _w11146_ ;
	wire _w11145_ ;
	wire _w11144_ ;
	wire _w11143_ ;
	wire _w11142_ ;
	wire _w11141_ ;
	wire _w11140_ ;
	wire _w11139_ ;
	wire _w11138_ ;
	wire _w11137_ ;
	wire _w11136_ ;
	wire _w11135_ ;
	wire _w11134_ ;
	wire _w11133_ ;
	wire _w11132_ ;
	wire _w11131_ ;
	wire _w11130_ ;
	wire _w11129_ ;
	wire _w11128_ ;
	wire _w11127_ ;
	wire _w11126_ ;
	wire _w11125_ ;
	wire _w11124_ ;
	wire _w11123_ ;
	wire _w11122_ ;
	wire _w11121_ ;
	wire _w11120_ ;
	wire _w11119_ ;
	wire _w11118_ ;
	wire _w11117_ ;
	wire _w11116_ ;
	wire _w11115_ ;
	wire _w11114_ ;
	wire _w11113_ ;
	wire _w11112_ ;
	wire _w11111_ ;
	wire _w11110_ ;
	wire _w11109_ ;
	wire _w11108_ ;
	wire _w11107_ ;
	wire _w11106_ ;
	wire _w11105_ ;
	wire _w11104_ ;
	wire _w11103_ ;
	wire _w11102_ ;
	wire _w11101_ ;
	wire _w11100_ ;
	wire _w11099_ ;
	wire _w11098_ ;
	wire _w11097_ ;
	wire _w11096_ ;
	wire _w11095_ ;
	wire _w11094_ ;
	wire _w11093_ ;
	wire _w11092_ ;
	wire _w11091_ ;
	wire _w11090_ ;
	wire _w11089_ ;
	wire _w11088_ ;
	wire _w11087_ ;
	wire _w11086_ ;
	wire _w11085_ ;
	wire _w11084_ ;
	wire _w11083_ ;
	wire _w11082_ ;
	wire _w11081_ ;
	wire _w11080_ ;
	wire _w11079_ ;
	wire _w11078_ ;
	wire _w11077_ ;
	wire _w11076_ ;
	wire _w11075_ ;
	wire _w11074_ ;
	wire _w11073_ ;
	wire _w11072_ ;
	wire _w11071_ ;
	wire _w11070_ ;
	wire _w11069_ ;
	wire _w11068_ ;
	wire _w11067_ ;
	wire _w11066_ ;
	wire _w11065_ ;
	wire _w11064_ ;
	wire _w11063_ ;
	wire _w11062_ ;
	wire _w11061_ ;
	wire _w11060_ ;
	wire _w11059_ ;
	wire _w11058_ ;
	wire _w11057_ ;
	wire _w11056_ ;
	wire _w11055_ ;
	wire _w11054_ ;
	wire _w11053_ ;
	wire _w11052_ ;
	wire _w11051_ ;
	wire _w11050_ ;
	wire _w11049_ ;
	wire _w11048_ ;
	wire _w11047_ ;
	wire _w11046_ ;
	wire _w11045_ ;
	wire _w11044_ ;
	wire _w11043_ ;
	wire _w11042_ ;
	wire _w11041_ ;
	wire _w11040_ ;
	wire _w11039_ ;
	wire _w11038_ ;
	wire _w11037_ ;
	wire _w11036_ ;
	wire _w11035_ ;
	wire _w11034_ ;
	wire _w11033_ ;
	wire _w11032_ ;
	wire _w11031_ ;
	wire _w11030_ ;
	wire _w11029_ ;
	wire _w11028_ ;
	wire _w11027_ ;
	wire _w11026_ ;
	wire _w11025_ ;
	wire _w11024_ ;
	wire _w11023_ ;
	wire _w11022_ ;
	wire _w11021_ ;
	wire _w11020_ ;
	wire _w11019_ ;
	wire _w11018_ ;
	wire _w11017_ ;
	wire _w11016_ ;
	wire _w11015_ ;
	wire _w11014_ ;
	wire _w11013_ ;
	wire _w11012_ ;
	wire _w11011_ ;
	wire _w11010_ ;
	wire _w11009_ ;
	wire _w11008_ ;
	wire _w11007_ ;
	wire _w11006_ ;
	wire _w11005_ ;
	wire _w11004_ ;
	wire _w11003_ ;
	wire _w11002_ ;
	wire _w11001_ ;
	wire _w11000_ ;
	wire _w10999_ ;
	wire _w10998_ ;
	wire _w10997_ ;
	wire _w10996_ ;
	wire _w10995_ ;
	wire _w10994_ ;
	wire _w10993_ ;
	wire _w10992_ ;
	wire _w10991_ ;
	wire _w10990_ ;
	wire _w10989_ ;
	wire _w10988_ ;
	wire _w10987_ ;
	wire _w10986_ ;
	wire _w10985_ ;
	wire _w10984_ ;
	wire _w10983_ ;
	wire _w10982_ ;
	wire _w10981_ ;
	wire _w10980_ ;
	wire _w10979_ ;
	wire _w10978_ ;
	wire _w10977_ ;
	wire _w10976_ ;
	wire _w10975_ ;
	wire _w10974_ ;
	wire _w10973_ ;
	wire _w10972_ ;
	wire _w10971_ ;
	wire _w10970_ ;
	wire _w10969_ ;
	wire _w10968_ ;
	wire _w10967_ ;
	wire _w10966_ ;
	wire _w10965_ ;
	wire _w10964_ ;
	wire _w10963_ ;
	wire _w10962_ ;
	wire _w10961_ ;
	wire _w10960_ ;
	wire _w10959_ ;
	wire _w10958_ ;
	wire _w10957_ ;
	wire _w10956_ ;
	wire _w10955_ ;
	wire _w10954_ ;
	wire _w10953_ ;
	wire _w10952_ ;
	wire _w10951_ ;
	wire _w10950_ ;
	wire _w10949_ ;
	wire _w10948_ ;
	wire _w10947_ ;
	wire _w10946_ ;
	wire _w10945_ ;
	wire _w10944_ ;
	wire _w10943_ ;
	wire _w10942_ ;
	wire _w10941_ ;
	wire _w10940_ ;
	wire _w10939_ ;
	wire _w10938_ ;
	wire _w10937_ ;
	wire _w10936_ ;
	wire _w10935_ ;
	wire _w10934_ ;
	wire _w10933_ ;
	wire _w10932_ ;
	wire _w10931_ ;
	wire _w10930_ ;
	wire _w10929_ ;
	wire _w10928_ ;
	wire _w10927_ ;
	wire _w10926_ ;
	wire _w10925_ ;
	wire _w10924_ ;
	wire _w10923_ ;
	wire _w10922_ ;
	wire _w10921_ ;
	wire _w10920_ ;
	wire _w10919_ ;
	wire _w10918_ ;
	wire _w10917_ ;
	wire _w10916_ ;
	wire _w10915_ ;
	wire _w10914_ ;
	wire _w10913_ ;
	wire _w10912_ ;
	wire _w10911_ ;
	wire _w10910_ ;
	wire _w10909_ ;
	wire _w10908_ ;
	wire _w10907_ ;
	wire _w10906_ ;
	wire _w10905_ ;
	wire _w10904_ ;
	wire _w10903_ ;
	wire _w10902_ ;
	wire _w10901_ ;
	wire _w10900_ ;
	wire _w10899_ ;
	wire _w10898_ ;
	wire _w10897_ ;
	wire _w10896_ ;
	wire _w10895_ ;
	wire _w10894_ ;
	wire _w10893_ ;
	wire _w10892_ ;
	wire _w10891_ ;
	wire _w10890_ ;
	wire _w10889_ ;
	wire _w10888_ ;
	wire _w10887_ ;
	wire _w10886_ ;
	wire _w10885_ ;
	wire _w10884_ ;
	wire _w10883_ ;
	wire _w10882_ ;
	wire _w10881_ ;
	wire _w10880_ ;
	wire _w10879_ ;
	wire _w10878_ ;
	wire _w10877_ ;
	wire _w10876_ ;
	wire _w10875_ ;
	wire _w10874_ ;
	wire _w10873_ ;
	wire _w10872_ ;
	wire _w10871_ ;
	wire _w10870_ ;
	wire _w10869_ ;
	wire _w10868_ ;
	wire _w10867_ ;
	wire _w10866_ ;
	wire _w10865_ ;
	wire _w10864_ ;
	wire _w10863_ ;
	wire _w10862_ ;
	wire _w10861_ ;
	wire _w10860_ ;
	wire _w10859_ ;
	wire _w10858_ ;
	wire _w10857_ ;
	wire _w10856_ ;
	wire _w10855_ ;
	wire _w10854_ ;
	wire _w10853_ ;
	wire _w10852_ ;
	wire _w10851_ ;
	wire _w10850_ ;
	wire _w10849_ ;
	wire _w10848_ ;
	wire _w10847_ ;
	wire _w10846_ ;
	wire _w10845_ ;
	wire _w10844_ ;
	wire _w10843_ ;
	wire _w10842_ ;
	wire _w10841_ ;
	wire _w10840_ ;
	wire _w10839_ ;
	wire _w10838_ ;
	wire _w10837_ ;
	wire _w10836_ ;
	wire _w10835_ ;
	wire _w10834_ ;
	wire _w10833_ ;
	wire _w10832_ ;
	wire _w10831_ ;
	wire _w10830_ ;
	wire _w10829_ ;
	wire _w10828_ ;
	wire _w10827_ ;
	wire _w10826_ ;
	wire _w10825_ ;
	wire _w10824_ ;
	wire _w10823_ ;
	wire _w10822_ ;
	wire _w10821_ ;
	wire _w10820_ ;
	wire _w10819_ ;
	wire _w10818_ ;
	wire _w10817_ ;
	wire _w10816_ ;
	wire _w10815_ ;
	wire _w10814_ ;
	wire _w10813_ ;
	wire _w10812_ ;
	wire _w10811_ ;
	wire _w10810_ ;
	wire _w10809_ ;
	wire _w10808_ ;
	wire _w10807_ ;
	wire _w10806_ ;
	wire _w10805_ ;
	wire _w10804_ ;
	wire _w10803_ ;
	wire _w10802_ ;
	wire _w10801_ ;
	wire _w10800_ ;
	wire _w10799_ ;
	wire _w10798_ ;
	wire _w10797_ ;
	wire _w10796_ ;
	wire _w10795_ ;
	wire _w10794_ ;
	wire _w10793_ ;
	wire _w10792_ ;
	wire _w10791_ ;
	wire _w10790_ ;
	wire _w10789_ ;
	wire _w10788_ ;
	wire _w10787_ ;
	wire _w10786_ ;
	wire _w10785_ ;
	wire _w10784_ ;
	wire _w10783_ ;
	wire _w10782_ ;
	wire _w10781_ ;
	wire _w10780_ ;
	wire _w10779_ ;
	wire _w10778_ ;
	wire _w10777_ ;
	wire _w10776_ ;
	wire _w10775_ ;
	wire _w10774_ ;
	wire _w10773_ ;
	wire _w10772_ ;
	wire _w10771_ ;
	wire _w10770_ ;
	wire _w10769_ ;
	wire _w10768_ ;
	wire _w10767_ ;
	wire _w10766_ ;
	wire _w10765_ ;
	wire _w10764_ ;
	wire _w10763_ ;
	wire _w10762_ ;
	wire _w10761_ ;
	wire _w10760_ ;
	wire _w10759_ ;
	wire _w10758_ ;
	wire _w10757_ ;
	wire _w10756_ ;
	wire _w10755_ ;
	wire _w10754_ ;
	wire _w10753_ ;
	wire _w10752_ ;
	wire _w10751_ ;
	wire _w10750_ ;
	wire _w10749_ ;
	wire _w10748_ ;
	wire _w10747_ ;
	wire _w10746_ ;
	wire _w10745_ ;
	wire _w10744_ ;
	wire _w10743_ ;
	wire _w10742_ ;
	wire _w10741_ ;
	wire _w10740_ ;
	wire _w10739_ ;
	wire _w10738_ ;
	wire _w10737_ ;
	wire _w10736_ ;
	wire _w10735_ ;
	wire _w10734_ ;
	wire _w10733_ ;
	wire _w10732_ ;
	wire _w10731_ ;
	wire _w10730_ ;
	wire _w10729_ ;
	wire _w10728_ ;
	wire _w10727_ ;
	wire _w10726_ ;
	wire _w10725_ ;
	wire _w10724_ ;
	wire _w10723_ ;
	wire _w10722_ ;
	wire _w10721_ ;
	wire _w10720_ ;
	wire _w10719_ ;
	wire _w10718_ ;
	wire _w10717_ ;
	wire _w10716_ ;
	wire _w10715_ ;
	wire _w10714_ ;
	wire _w10713_ ;
	wire _w10712_ ;
	wire _w10711_ ;
	wire _w10710_ ;
	wire _w10709_ ;
	wire _w10708_ ;
	wire _w10707_ ;
	wire _w10706_ ;
	wire _w10705_ ;
	wire _w10704_ ;
	wire _w10703_ ;
	wire _w10702_ ;
	wire _w10701_ ;
	wire _w10700_ ;
	wire _w10699_ ;
	wire _w10698_ ;
	wire _w10697_ ;
	wire _w10696_ ;
	wire _w10695_ ;
	wire _w10694_ ;
	wire _w10693_ ;
	wire _w10692_ ;
	wire _w10691_ ;
	wire _w10690_ ;
	wire _w10689_ ;
	wire _w10688_ ;
	wire _w10687_ ;
	wire _w10686_ ;
	wire _w10685_ ;
	wire _w10684_ ;
	wire _w10683_ ;
	wire _w10682_ ;
	wire _w10681_ ;
	wire _w10680_ ;
	wire _w10679_ ;
	wire _w10678_ ;
	wire _w10677_ ;
	wire _w10676_ ;
	wire _w10675_ ;
	wire _w10674_ ;
	wire _w10673_ ;
	wire _w10672_ ;
	wire _w10671_ ;
	wire _w10670_ ;
	wire _w10669_ ;
	wire _w10668_ ;
	wire _w10667_ ;
	wire _w10666_ ;
	wire _w10665_ ;
	wire _w10664_ ;
	wire _w10663_ ;
	wire _w10662_ ;
	wire _w10661_ ;
	wire _w10660_ ;
	wire _w10659_ ;
	wire _w10658_ ;
	wire _w10657_ ;
	wire _w10656_ ;
	wire _w10655_ ;
	wire _w10654_ ;
	wire _w10653_ ;
	wire _w10652_ ;
	wire _w10651_ ;
	wire _w10650_ ;
	wire _w10649_ ;
	wire _w10648_ ;
	wire _w10647_ ;
	wire _w10646_ ;
	wire _w10645_ ;
	wire _w10644_ ;
	wire _w10643_ ;
	wire _w10642_ ;
	wire _w10641_ ;
	wire _w10640_ ;
	wire _w10639_ ;
	wire _w10638_ ;
	wire _w10637_ ;
	wire _w10636_ ;
	wire _w10635_ ;
	wire _w10634_ ;
	wire _w10633_ ;
	wire _w10632_ ;
	wire _w10631_ ;
	wire _w10630_ ;
	wire _w10629_ ;
	wire _w10628_ ;
	wire _w10627_ ;
	wire _w10626_ ;
	wire _w10625_ ;
	wire _w10624_ ;
	wire _w10623_ ;
	wire _w10622_ ;
	wire _w10621_ ;
	wire _w10620_ ;
	wire _w10619_ ;
	wire _w10618_ ;
	wire _w10617_ ;
	wire _w10616_ ;
	wire _w10615_ ;
	wire _w10614_ ;
	wire _w10613_ ;
	wire _w10612_ ;
	wire _w10611_ ;
	wire _w10610_ ;
	wire _w10609_ ;
	wire _w10608_ ;
	wire _w10607_ ;
	wire _w10606_ ;
	wire _w10605_ ;
	wire _w10604_ ;
	wire _w10603_ ;
	wire _w10602_ ;
	wire _w10601_ ;
	wire _w10600_ ;
	wire _w10599_ ;
	wire _w10598_ ;
	wire _w10597_ ;
	wire _w10596_ ;
	wire _w10595_ ;
	wire _w10594_ ;
	wire _w10593_ ;
	wire _w10592_ ;
	wire _w10591_ ;
	wire _w10590_ ;
	wire _w10589_ ;
	wire _w10588_ ;
	wire _w10587_ ;
	wire _w10586_ ;
	wire _w10585_ ;
	wire _w10584_ ;
	wire _w10583_ ;
	wire _w10582_ ;
	wire _w10581_ ;
	wire _w10580_ ;
	wire _w10579_ ;
	wire _w10578_ ;
	wire _w10577_ ;
	wire _w10576_ ;
	wire _w10575_ ;
	wire _w10574_ ;
	wire _w10573_ ;
	wire _w10572_ ;
	wire _w10571_ ;
	wire _w10570_ ;
	wire _w10569_ ;
	wire _w10568_ ;
	wire _w10567_ ;
	wire _w10566_ ;
	wire _w10565_ ;
	wire _w10564_ ;
	wire _w10563_ ;
	wire _w10562_ ;
	wire _w10561_ ;
	wire _w10560_ ;
	wire _w10559_ ;
	wire _w10558_ ;
	wire _w10557_ ;
	wire _w10556_ ;
	wire _w10555_ ;
	wire _w10554_ ;
	wire _w10553_ ;
	wire _w10552_ ;
	wire _w10551_ ;
	wire _w10550_ ;
	wire _w10549_ ;
	wire _w10548_ ;
	wire _w10547_ ;
	wire _w10546_ ;
	wire _w10545_ ;
	wire _w10544_ ;
	wire _w10543_ ;
	wire _w10542_ ;
	wire _w10541_ ;
	wire _w10540_ ;
	wire _w10539_ ;
	wire _w10538_ ;
	wire _w10537_ ;
	wire _w10536_ ;
	wire _w10535_ ;
	wire _w10534_ ;
	wire _w10533_ ;
	wire _w10532_ ;
	wire _w10531_ ;
	wire _w10530_ ;
	wire _w10529_ ;
	wire _w10528_ ;
	wire _w10527_ ;
	wire _w10526_ ;
	wire _w10525_ ;
	wire _w10524_ ;
	wire _w10523_ ;
	wire _w10522_ ;
	wire _w10521_ ;
	wire _w10520_ ;
	wire _w10519_ ;
	wire _w10518_ ;
	wire _w10517_ ;
	wire _w10516_ ;
	wire _w10515_ ;
	wire _w10514_ ;
	wire _w10513_ ;
	wire _w10512_ ;
	wire _w10511_ ;
	wire _w10510_ ;
	wire _w10509_ ;
	wire _w10508_ ;
	wire _w10507_ ;
	wire _w10506_ ;
	wire _w10505_ ;
	wire _w10504_ ;
	wire _w10503_ ;
	wire _w10502_ ;
	wire _w10501_ ;
	wire _w10500_ ;
	wire _w10499_ ;
	wire _w10498_ ;
	wire _w10497_ ;
	wire _w10496_ ;
	wire _w10495_ ;
	wire _w10494_ ;
	wire _w10493_ ;
	wire _w10492_ ;
	wire _w10491_ ;
	wire _w10490_ ;
	wire _w10489_ ;
	wire _w10488_ ;
	wire _w10487_ ;
	wire _w10486_ ;
	wire _w10485_ ;
	wire _w10484_ ;
	wire _w10483_ ;
	wire _w10482_ ;
	wire _w10481_ ;
	wire _w10480_ ;
	wire _w10479_ ;
	wire _w10478_ ;
	wire _w10477_ ;
	wire _w10476_ ;
	wire _w10475_ ;
	wire _w10474_ ;
	wire _w10473_ ;
	wire _w10472_ ;
	wire _w10471_ ;
	wire _w10470_ ;
	wire _w10469_ ;
	wire _w10468_ ;
	wire _w10467_ ;
	wire _w10466_ ;
	wire _w10465_ ;
	wire _w10464_ ;
	wire _w10463_ ;
	wire _w10462_ ;
	wire _w10461_ ;
	wire _w10460_ ;
	wire _w10459_ ;
	wire _w10458_ ;
	wire _w10457_ ;
	wire _w10456_ ;
	wire _w10455_ ;
	wire _w10454_ ;
	wire _w10453_ ;
	wire _w10452_ ;
	wire _w10451_ ;
	wire _w10450_ ;
	wire _w10449_ ;
	wire _w10448_ ;
	wire _w10447_ ;
	wire _w10446_ ;
	wire _w10445_ ;
	wire _w10444_ ;
	wire _w10443_ ;
	wire _w10442_ ;
	wire _w10441_ ;
	wire _w10440_ ;
	wire _w10439_ ;
	wire _w10438_ ;
	wire _w10437_ ;
	wire _w10436_ ;
	wire _w10435_ ;
	wire _w10434_ ;
	wire _w10433_ ;
	wire _w10432_ ;
	wire _w10431_ ;
	wire _w10430_ ;
	wire _w10429_ ;
	wire _w10428_ ;
	wire _w10427_ ;
	wire _w10426_ ;
	wire _w10425_ ;
	wire _w10424_ ;
	wire _w10423_ ;
	wire _w10422_ ;
	wire _w10421_ ;
	wire _w10420_ ;
	wire _w10419_ ;
	wire _w10418_ ;
	wire _w10417_ ;
	wire _w10416_ ;
	wire _w10415_ ;
	wire _w10414_ ;
	wire _w10413_ ;
	wire _w10412_ ;
	wire _w10411_ ;
	wire _w10410_ ;
	wire _w10409_ ;
	wire _w10408_ ;
	wire _w10407_ ;
	wire _w10406_ ;
	wire _w10405_ ;
	wire _w10404_ ;
	wire _w10403_ ;
	wire _w10402_ ;
	wire _w10401_ ;
	wire _w10400_ ;
	wire _w10399_ ;
	wire _w10398_ ;
	wire _w10397_ ;
	wire _w10396_ ;
	wire _w10395_ ;
	wire _w10394_ ;
	wire _w10393_ ;
	wire _w10392_ ;
	wire _w10391_ ;
	wire _w10390_ ;
	wire _w10389_ ;
	wire _w10388_ ;
	wire _w10387_ ;
	wire _w10386_ ;
	wire _w10385_ ;
	wire _w10384_ ;
	wire _w10383_ ;
	wire _w10382_ ;
	wire _w10381_ ;
	wire _w10380_ ;
	wire _w10379_ ;
	wire _w10378_ ;
	wire _w10377_ ;
	wire _w10376_ ;
	wire _w10375_ ;
	wire _w10374_ ;
	wire _w10373_ ;
	wire _w10372_ ;
	wire _w10371_ ;
	wire _w10370_ ;
	wire _w10369_ ;
	wire _w10368_ ;
	wire _w10367_ ;
	wire _w10366_ ;
	wire _w10365_ ;
	wire _w10364_ ;
	wire _w10363_ ;
	wire _w10362_ ;
	wire _w10361_ ;
	wire _w10360_ ;
	wire _w10359_ ;
	wire _w10358_ ;
	wire _w10357_ ;
	wire _w10356_ ;
	wire _w10355_ ;
	wire _w10354_ ;
	wire _w10353_ ;
	wire _w10352_ ;
	wire _w10351_ ;
	wire _w10350_ ;
	wire _w10349_ ;
	wire _w10348_ ;
	wire _w10347_ ;
	wire _w10346_ ;
	wire _w10345_ ;
	wire _w10344_ ;
	wire _w10343_ ;
	wire _w10342_ ;
	wire _w10341_ ;
	wire _w10340_ ;
	wire _w10339_ ;
	wire _w10338_ ;
	wire _w10337_ ;
	wire _w10336_ ;
	wire _w10335_ ;
	wire _w10334_ ;
	wire _w10333_ ;
	wire _w10332_ ;
	wire _w10331_ ;
	wire _w10330_ ;
	wire _w10329_ ;
	wire _w10328_ ;
	wire _w10327_ ;
	wire _w10326_ ;
	wire _w10325_ ;
	wire _w10324_ ;
	wire _w10323_ ;
	wire _w10322_ ;
	wire _w10321_ ;
	wire _w10320_ ;
	wire _w10319_ ;
	wire _w10318_ ;
	wire _w10317_ ;
	wire _w10316_ ;
	wire _w10315_ ;
	wire _w10314_ ;
	wire _w10313_ ;
	wire _w10312_ ;
	wire _w10311_ ;
	wire _w10310_ ;
	wire _w10309_ ;
	wire _w10308_ ;
	wire _w10307_ ;
	wire _w10306_ ;
	wire _w10305_ ;
	wire _w10304_ ;
	wire _w10303_ ;
	wire _w10302_ ;
	wire _w10301_ ;
	wire _w10300_ ;
	wire _w10299_ ;
	wire _w10298_ ;
	wire _w10297_ ;
	wire _w10296_ ;
	wire _w10295_ ;
	wire _w10294_ ;
	wire _w10293_ ;
	wire _w10292_ ;
	wire _w10291_ ;
	wire _w10290_ ;
	wire _w10289_ ;
	wire _w10288_ ;
	wire _w10287_ ;
	wire _w10286_ ;
	wire _w10285_ ;
	wire _w10284_ ;
	wire _w10283_ ;
	wire _w10282_ ;
	wire _w10281_ ;
	wire _w10280_ ;
	wire _w10279_ ;
	wire _w10278_ ;
	wire _w10277_ ;
	wire _w10276_ ;
	wire _w10275_ ;
	wire _w10274_ ;
	wire _w10273_ ;
	wire _w10272_ ;
	wire _w10271_ ;
	wire _w10270_ ;
	wire _w10269_ ;
	wire _w10268_ ;
	wire _w10267_ ;
	wire _w10266_ ;
	wire _w10265_ ;
	wire _w10264_ ;
	wire _w10263_ ;
	wire _w10262_ ;
	wire _w10261_ ;
	wire _w10260_ ;
	wire _w10259_ ;
	wire _w10258_ ;
	wire _w10257_ ;
	wire _w10256_ ;
	wire _w10255_ ;
	wire _w10254_ ;
	wire _w10253_ ;
	wire _w10252_ ;
	wire _w10251_ ;
	wire _w10250_ ;
	wire _w10249_ ;
	wire _w10248_ ;
	wire _w10247_ ;
	wire _w10246_ ;
	wire _w10245_ ;
	wire _w10244_ ;
	wire _w10243_ ;
	wire _w10242_ ;
	wire _w10241_ ;
	wire _w10240_ ;
	wire _w10239_ ;
	wire _w10238_ ;
	wire _w10237_ ;
	wire _w10236_ ;
	wire _w10235_ ;
	wire _w10234_ ;
	wire _w10233_ ;
	wire _w10232_ ;
	wire _w10231_ ;
	wire _w10230_ ;
	wire _w10229_ ;
	wire _w10228_ ;
	wire _w10227_ ;
	wire _w10226_ ;
	wire _w10225_ ;
	wire _w10224_ ;
	wire _w10223_ ;
	wire _w10222_ ;
	wire _w10221_ ;
	wire _w10220_ ;
	wire _w10219_ ;
	wire _w10218_ ;
	wire _w10217_ ;
	wire _w10216_ ;
	wire _w10215_ ;
	wire _w10214_ ;
	wire _w10213_ ;
	wire _w10212_ ;
	wire _w10211_ ;
	wire _w10210_ ;
	wire _w10209_ ;
	wire _w10208_ ;
	wire _w10207_ ;
	wire _w10206_ ;
	wire _w10205_ ;
	wire _w10204_ ;
	wire _w10203_ ;
	wire _w10202_ ;
	wire _w10201_ ;
	wire _w10200_ ;
	wire _w10199_ ;
	wire _w10198_ ;
	wire _w10197_ ;
	wire _w10196_ ;
	wire _w10195_ ;
	wire _w10194_ ;
	wire _w10193_ ;
	wire _w10192_ ;
	wire _w10191_ ;
	wire _w10190_ ;
	wire _w10189_ ;
	wire _w10188_ ;
	wire _w10187_ ;
	wire _w10186_ ;
	wire _w10185_ ;
	wire _w10184_ ;
	wire _w10183_ ;
	wire _w10182_ ;
	wire _w10181_ ;
	wire _w10180_ ;
	wire _w10179_ ;
	wire _w10178_ ;
	wire _w10177_ ;
	wire _w10176_ ;
	wire _w10175_ ;
	wire _w10174_ ;
	wire _w10173_ ;
	wire _w10172_ ;
	wire _w10171_ ;
	wire _w10170_ ;
	wire _w10169_ ;
	wire _w10168_ ;
	wire _w10167_ ;
	wire _w10166_ ;
	wire _w10165_ ;
	wire _w10164_ ;
	wire _w10163_ ;
	wire _w10162_ ;
	wire _w10161_ ;
	wire _w10160_ ;
	wire _w10159_ ;
	wire _w10158_ ;
	wire _w10157_ ;
	wire _w10156_ ;
	wire _w10155_ ;
	wire _w10154_ ;
	wire _w10153_ ;
	wire _w10152_ ;
	wire _w10151_ ;
	wire _w10150_ ;
	wire _w10149_ ;
	wire _w10148_ ;
	wire _w10147_ ;
	wire _w10146_ ;
	wire _w10145_ ;
	wire _w10144_ ;
	wire _w10143_ ;
	wire _w10142_ ;
	wire _w10141_ ;
	wire _w10140_ ;
	wire _w10139_ ;
	wire _w10138_ ;
	wire _w10137_ ;
	wire _w10136_ ;
	wire _w10135_ ;
	wire _w10134_ ;
	wire _w10133_ ;
	wire _w10132_ ;
	wire _w10131_ ;
	wire _w10130_ ;
	wire _w10129_ ;
	wire _w10128_ ;
	wire _w10127_ ;
	wire _w10126_ ;
	wire _w10125_ ;
	wire _w10124_ ;
	wire _w10123_ ;
	wire _w10122_ ;
	wire _w10121_ ;
	wire _w10120_ ;
	wire _w10119_ ;
	wire _w10118_ ;
	wire _w10117_ ;
	wire _w10116_ ;
	wire _w10115_ ;
	wire _w10114_ ;
	wire _w10113_ ;
	wire _w10112_ ;
	wire _w10111_ ;
	wire _w10110_ ;
	wire _w10109_ ;
	wire _w10108_ ;
	wire _w10107_ ;
	wire _w10106_ ;
	wire _w10105_ ;
	wire _w10104_ ;
	wire _w10103_ ;
	wire _w10102_ ;
	wire _w10101_ ;
	wire _w10100_ ;
	wire _w10099_ ;
	wire _w10098_ ;
	wire _w10097_ ;
	wire _w10096_ ;
	wire _w10095_ ;
	wire _w10094_ ;
	wire _w10093_ ;
	wire _w10092_ ;
	wire _w10091_ ;
	wire _w10090_ ;
	wire _w10089_ ;
	wire _w10088_ ;
	wire _w10087_ ;
	wire _w10086_ ;
	wire _w10085_ ;
	wire _w10084_ ;
	wire _w10083_ ;
	wire _w10082_ ;
	wire _w10081_ ;
	wire _w10080_ ;
	wire _w10079_ ;
	wire _w10078_ ;
	wire _w10077_ ;
	wire _w10076_ ;
	wire _w10075_ ;
	wire _w10074_ ;
	wire _w10073_ ;
	wire _w10072_ ;
	wire _w10071_ ;
	wire _w10070_ ;
	wire _w10069_ ;
	wire _w10068_ ;
	wire _w10067_ ;
	wire _w10066_ ;
	wire _w10065_ ;
	wire _w10064_ ;
	wire _w10063_ ;
	wire _w10062_ ;
	wire _w10061_ ;
	wire _w10060_ ;
	wire _w10059_ ;
	wire _w10058_ ;
	wire _w10057_ ;
	wire _w10056_ ;
	wire _w10055_ ;
	wire _w10054_ ;
	wire _w10053_ ;
	wire _w10052_ ;
	wire _w10051_ ;
	wire _w10050_ ;
	wire _w10049_ ;
	wire _w10048_ ;
	wire _w10047_ ;
	wire _w10046_ ;
	wire _w10045_ ;
	wire _w10044_ ;
	wire _w10043_ ;
	wire _w10042_ ;
	wire _w10041_ ;
	wire _w10040_ ;
	wire _w10039_ ;
	wire _w10038_ ;
	wire _w10037_ ;
	wire _w10036_ ;
	wire _w10035_ ;
	wire _w10034_ ;
	wire _w10033_ ;
	wire _w10032_ ;
	wire _w10031_ ;
	wire _w10030_ ;
	wire _w10029_ ;
	wire _w10028_ ;
	wire _w10027_ ;
	wire _w10026_ ;
	wire _w10025_ ;
	wire _w10024_ ;
	wire _w10023_ ;
	wire _w10022_ ;
	wire _w10021_ ;
	wire _w10020_ ;
	wire _w10019_ ;
	wire _w10018_ ;
	wire _w10017_ ;
	wire _w10016_ ;
	wire _w10015_ ;
	wire _w10014_ ;
	wire _w10013_ ;
	wire _w10012_ ;
	wire _w10011_ ;
	wire _w10010_ ;
	wire _w10009_ ;
	wire _w10008_ ;
	wire _w10007_ ;
	wire _w10006_ ;
	wire _w10005_ ;
	wire _w10004_ ;
	wire _w10003_ ;
	wire _w10002_ ;
	wire _w10001_ ;
	wire _w10000_ ;
	wire _w9999_ ;
	wire _w9998_ ;
	wire _w9997_ ;
	wire _w9996_ ;
	wire _w9995_ ;
	wire _w9994_ ;
	wire _w9993_ ;
	wire _w9992_ ;
	wire _w9991_ ;
	wire _w9990_ ;
	wire _w9989_ ;
	wire _w9988_ ;
	wire _w9987_ ;
	wire _w9986_ ;
	wire _w9985_ ;
	wire _w9984_ ;
	wire _w9983_ ;
	wire _w9982_ ;
	wire _w9981_ ;
	wire _w9980_ ;
	wire _w9979_ ;
	wire _w9978_ ;
	wire _w9977_ ;
	wire _w9976_ ;
	wire _w9975_ ;
	wire _w9974_ ;
	wire _w9973_ ;
	wire _w9972_ ;
	wire _w9971_ ;
	wire _w9970_ ;
	wire _w9969_ ;
	wire _w9968_ ;
	wire _w9967_ ;
	wire _w9966_ ;
	wire _w9965_ ;
	wire _w9964_ ;
	wire _w9963_ ;
	wire _w9962_ ;
	wire _w9961_ ;
	wire _w9960_ ;
	wire _w9959_ ;
	wire _w9958_ ;
	wire _w9957_ ;
	wire _w9956_ ;
	wire _w9955_ ;
	wire _w9954_ ;
	wire _w9953_ ;
	wire _w9952_ ;
	wire _w9951_ ;
	wire _w9950_ ;
	wire _w9949_ ;
	wire _w9948_ ;
	wire _w9947_ ;
	wire _w9946_ ;
	wire _w9945_ ;
	wire _w9944_ ;
	wire _w9943_ ;
	wire _w9942_ ;
	wire _w9941_ ;
	wire _w9940_ ;
	wire _w9939_ ;
	wire _w9938_ ;
	wire _w9937_ ;
	wire _w9936_ ;
	wire _w9935_ ;
	wire _w9934_ ;
	wire _w9933_ ;
	wire _w9932_ ;
	wire _w9931_ ;
	wire _w9930_ ;
	wire _w9929_ ;
	wire _w9928_ ;
	wire _w9927_ ;
	wire _w9926_ ;
	wire _w9925_ ;
	wire _w9924_ ;
	wire _w9923_ ;
	wire _w9922_ ;
	wire _w9921_ ;
	wire _w9920_ ;
	wire _w9919_ ;
	wire _w9918_ ;
	wire _w9917_ ;
	wire _w9916_ ;
	wire _w9915_ ;
	wire _w9914_ ;
	wire _w9913_ ;
	wire _w9912_ ;
	wire _w9911_ ;
	wire _w9910_ ;
	wire _w9909_ ;
	wire _w9908_ ;
	wire _w9907_ ;
	wire _w9906_ ;
	wire _w9905_ ;
	wire _w9904_ ;
	wire _w9903_ ;
	wire _w9902_ ;
	wire _w9901_ ;
	wire _w9900_ ;
	wire _w9899_ ;
	wire _w9898_ ;
	wire _w9897_ ;
	wire _w9896_ ;
	wire _w9895_ ;
	wire _w9894_ ;
	wire _w9893_ ;
	wire _w9892_ ;
	wire _w9891_ ;
	wire _w9890_ ;
	wire _w9889_ ;
	wire _w9888_ ;
	wire _w9887_ ;
	wire _w9886_ ;
	wire _w9885_ ;
	wire _w9884_ ;
	wire _w9883_ ;
	wire _w9882_ ;
	wire _w9881_ ;
	wire _w9880_ ;
	wire _w9879_ ;
	wire _w9878_ ;
	wire _w9877_ ;
	wire _w9876_ ;
	wire _w9875_ ;
	wire _w9874_ ;
	wire _w9873_ ;
	wire _w9872_ ;
	wire _w9871_ ;
	wire _w9870_ ;
	wire _w9869_ ;
	wire _w9868_ ;
	wire _w9867_ ;
	wire _w9866_ ;
	wire _w9865_ ;
	wire _w9864_ ;
	wire _w9863_ ;
	wire _w9862_ ;
	wire _w9861_ ;
	wire _w9860_ ;
	wire _w9859_ ;
	wire _w9858_ ;
	wire _w9857_ ;
	wire _w9856_ ;
	wire _w9855_ ;
	wire _w9854_ ;
	wire _w9853_ ;
	wire _w9852_ ;
	wire _w9851_ ;
	wire _w9850_ ;
	wire _w9849_ ;
	wire _w9848_ ;
	wire _w9847_ ;
	wire _w9846_ ;
	wire _w9845_ ;
	wire _w9844_ ;
	wire _w9843_ ;
	wire _w9842_ ;
	wire _w9841_ ;
	wire _w9840_ ;
	wire _w9839_ ;
	wire _w9838_ ;
	wire _w9837_ ;
	wire _w9836_ ;
	wire _w9835_ ;
	wire _w9834_ ;
	wire _w9833_ ;
	wire _w9832_ ;
	wire _w9831_ ;
	wire _w9830_ ;
	wire _w9829_ ;
	wire _w9828_ ;
	wire _w9827_ ;
	wire _w9826_ ;
	wire _w9825_ ;
	wire _w9824_ ;
	wire _w9823_ ;
	wire _w9822_ ;
	wire _w9821_ ;
	wire _w9820_ ;
	wire _w9819_ ;
	wire _w9818_ ;
	wire _w9817_ ;
	wire _w9816_ ;
	wire _w9815_ ;
	wire _w9814_ ;
	wire _w9813_ ;
	wire _w9812_ ;
	wire _w9811_ ;
	wire _w9810_ ;
	wire _w9809_ ;
	wire _w9808_ ;
	wire _w9807_ ;
	wire _w9806_ ;
	wire _w9805_ ;
	wire _w9804_ ;
	wire _w9803_ ;
	wire _w9802_ ;
	wire _w9801_ ;
	wire _w9800_ ;
	wire _w9799_ ;
	wire _w9798_ ;
	wire _w9797_ ;
	wire _w9796_ ;
	wire _w9795_ ;
	wire _w9794_ ;
	wire _w9793_ ;
	wire _w9792_ ;
	wire _w9791_ ;
	wire _w9790_ ;
	wire _w9789_ ;
	wire _w9788_ ;
	wire _w9787_ ;
	wire _w9786_ ;
	wire _w9785_ ;
	wire _w9784_ ;
	wire _w9783_ ;
	wire _w9782_ ;
	wire _w9781_ ;
	wire _w9780_ ;
	wire _w9779_ ;
	wire _w9778_ ;
	wire _w9777_ ;
	wire _w9776_ ;
	wire _w9775_ ;
	wire _w9774_ ;
	wire _w9773_ ;
	wire _w9772_ ;
	wire _w9771_ ;
	wire _w9770_ ;
	wire _w9769_ ;
	wire _w9768_ ;
	wire _w9767_ ;
	wire _w9766_ ;
	wire _w9765_ ;
	wire _w9764_ ;
	wire _w9763_ ;
	wire _w9762_ ;
	wire _w9761_ ;
	wire _w9760_ ;
	wire _w9759_ ;
	wire _w9758_ ;
	wire _w9757_ ;
	wire _w9756_ ;
	wire _w9755_ ;
	wire _w9754_ ;
	wire _w9753_ ;
	wire _w9752_ ;
	wire _w9751_ ;
	wire _w9750_ ;
	wire _w9749_ ;
	wire _w9748_ ;
	wire _w9747_ ;
	wire _w9746_ ;
	wire _w9745_ ;
	wire _w9744_ ;
	wire _w9743_ ;
	wire _w9742_ ;
	wire _w9741_ ;
	wire _w9740_ ;
	wire _w9739_ ;
	wire _w9738_ ;
	wire _w9737_ ;
	wire _w9736_ ;
	wire _w9735_ ;
	wire _w9734_ ;
	wire _w9733_ ;
	wire _w9732_ ;
	wire _w9731_ ;
	wire _w9730_ ;
	wire _w9729_ ;
	wire _w9728_ ;
	wire _w9727_ ;
	wire _w9726_ ;
	wire _w9725_ ;
	wire _w9724_ ;
	wire _w9723_ ;
	wire _w9722_ ;
	wire _w9721_ ;
	wire _w9720_ ;
	wire _w9719_ ;
	wire _w9718_ ;
	wire _w9717_ ;
	wire _w9716_ ;
	wire _w9715_ ;
	wire _w9714_ ;
	wire _w9713_ ;
	wire _w9712_ ;
	wire _w9711_ ;
	wire _w9710_ ;
	wire _w9709_ ;
	wire _w9708_ ;
	wire _w9707_ ;
	wire _w9706_ ;
	wire _w9705_ ;
	wire _w9704_ ;
	wire _w9703_ ;
	wire _w9702_ ;
	wire _w9701_ ;
	wire _w9700_ ;
	wire _w9699_ ;
	wire _w9698_ ;
	wire _w9697_ ;
	wire _w9696_ ;
	wire _w9695_ ;
	wire _w9694_ ;
	wire _w9693_ ;
	wire _w9692_ ;
	wire _w9691_ ;
	wire _w9690_ ;
	wire _w9689_ ;
	wire _w9688_ ;
	wire _w9687_ ;
	wire _w9686_ ;
	wire _w9685_ ;
	wire _w9684_ ;
	wire _w9683_ ;
	wire _w9682_ ;
	wire _w9681_ ;
	wire _w9680_ ;
	wire _w9679_ ;
	wire _w9678_ ;
	wire _w9677_ ;
	wire _w9676_ ;
	wire _w9675_ ;
	wire _w9674_ ;
	wire _w9673_ ;
	wire _w9672_ ;
	wire _w9671_ ;
	wire _w9670_ ;
	wire _w9669_ ;
	wire _w9668_ ;
	wire _w9667_ ;
	wire _w9666_ ;
	wire _w9665_ ;
	wire _w9664_ ;
	wire _w9663_ ;
	wire _w9662_ ;
	wire _w9661_ ;
	wire _w9660_ ;
	wire _w9659_ ;
	wire _w9658_ ;
	wire _w9657_ ;
	wire _w9656_ ;
	wire _w9655_ ;
	wire _w9654_ ;
	wire _w9653_ ;
	wire _w9652_ ;
	wire _w9651_ ;
	wire _w9650_ ;
	wire _w9649_ ;
	wire _w9648_ ;
	wire _w9647_ ;
	wire _w9646_ ;
	wire _w9645_ ;
	wire _w9644_ ;
	wire _w9643_ ;
	wire _w9642_ ;
	wire _w9641_ ;
	wire _w9640_ ;
	wire _w9639_ ;
	wire _w9638_ ;
	wire _w9637_ ;
	wire _w9636_ ;
	wire _w9635_ ;
	wire _w9634_ ;
	wire _w9633_ ;
	wire _w9632_ ;
	wire _w9631_ ;
	wire _w9630_ ;
	wire _w9629_ ;
	wire _w9628_ ;
	wire _w9627_ ;
	wire _w9626_ ;
	wire _w9625_ ;
	wire _w9624_ ;
	wire _w9623_ ;
	wire _w9622_ ;
	wire _w9621_ ;
	wire _w9620_ ;
	wire _w9619_ ;
	wire _w9618_ ;
	wire _w9617_ ;
	wire _w9616_ ;
	wire _w9615_ ;
	wire _w9614_ ;
	wire _w9613_ ;
	wire _w9612_ ;
	wire _w9611_ ;
	wire _w9610_ ;
	wire _w9609_ ;
	wire _w9608_ ;
	wire _w9607_ ;
	wire _w9606_ ;
	wire _w9605_ ;
	wire _w9604_ ;
	wire _w9603_ ;
	wire _w9602_ ;
	wire _w9601_ ;
	wire _w9600_ ;
	wire _w9599_ ;
	wire _w9598_ ;
	wire _w9597_ ;
	wire _w9596_ ;
	wire _w9595_ ;
	wire _w9594_ ;
	wire _w9593_ ;
	wire _w9592_ ;
	wire _w9591_ ;
	wire _w9590_ ;
	wire _w9589_ ;
	wire _w9588_ ;
	wire _w9587_ ;
	wire _w9586_ ;
	wire _w9585_ ;
	wire _w9584_ ;
	wire _w9583_ ;
	wire _w9582_ ;
	wire _w9581_ ;
	wire _w9580_ ;
	wire _w9579_ ;
	wire _w9578_ ;
	wire _w9577_ ;
	wire _w9576_ ;
	wire _w9575_ ;
	wire _w9574_ ;
	wire _w9573_ ;
	wire _w9572_ ;
	wire _w9571_ ;
	wire _w9570_ ;
	wire _w9569_ ;
	wire _w9568_ ;
	wire _w9567_ ;
	wire _w9566_ ;
	wire _w9565_ ;
	wire _w9564_ ;
	wire _w9563_ ;
	wire _w9562_ ;
	wire _w9561_ ;
	wire _w9560_ ;
	wire _w9559_ ;
	wire _w9558_ ;
	wire _w9557_ ;
	wire _w9556_ ;
	wire _w9555_ ;
	wire _w9554_ ;
	wire _w9553_ ;
	wire _w9552_ ;
	wire _w9551_ ;
	wire _w9550_ ;
	wire _w9549_ ;
	wire _w9548_ ;
	wire _w9547_ ;
	wire _w9546_ ;
	wire _w9545_ ;
	wire _w9544_ ;
	wire _w9543_ ;
	wire _w9542_ ;
	wire _w9541_ ;
	wire _w9540_ ;
	wire _w9539_ ;
	wire _w9538_ ;
	wire _w9537_ ;
	wire _w9536_ ;
	wire _w9535_ ;
	wire _w9534_ ;
	wire _w9533_ ;
	wire _w9532_ ;
	wire _w9531_ ;
	wire _w9530_ ;
	wire _w9529_ ;
	wire _w9528_ ;
	wire _w9527_ ;
	wire _w9526_ ;
	wire _w9525_ ;
	wire _w9524_ ;
	wire _w9523_ ;
	wire _w9522_ ;
	wire _w9521_ ;
	wire _w9520_ ;
	wire _w9519_ ;
	wire _w9518_ ;
	wire _w9517_ ;
	wire _w9516_ ;
	wire _w9515_ ;
	wire _w9514_ ;
	wire _w9513_ ;
	wire _w9512_ ;
	wire _w9511_ ;
	wire _w9510_ ;
	wire _w9509_ ;
	wire _w9508_ ;
	wire _w9507_ ;
	wire _w9506_ ;
	wire _w9505_ ;
	wire _w9504_ ;
	wire _w9503_ ;
	wire _w9502_ ;
	wire _w9501_ ;
	wire _w9500_ ;
	wire _w9499_ ;
	wire _w9498_ ;
	wire _w9497_ ;
	wire _w9496_ ;
	wire _w9495_ ;
	wire _w9494_ ;
	wire _w9493_ ;
	wire _w9492_ ;
	wire _w9491_ ;
	wire _w9490_ ;
	wire _w9489_ ;
	wire _w9488_ ;
	wire _w9487_ ;
	wire _w9486_ ;
	wire _w9485_ ;
	wire _w9484_ ;
	wire _w9483_ ;
	wire _w9482_ ;
	wire _w9481_ ;
	wire _w9480_ ;
	wire _w9479_ ;
	wire _w9478_ ;
	wire _w9477_ ;
	wire _w9476_ ;
	wire _w9475_ ;
	wire _w9474_ ;
	wire _w9473_ ;
	wire _w9472_ ;
	wire _w9471_ ;
	wire _w9470_ ;
	wire _w9469_ ;
	wire _w9468_ ;
	wire _w9467_ ;
	wire _w9466_ ;
	wire _w9465_ ;
	wire _w9464_ ;
	wire _w9463_ ;
	wire _w9462_ ;
	wire _w9461_ ;
	wire _w9460_ ;
	wire _w9459_ ;
	wire _w9458_ ;
	wire _w9457_ ;
	wire _w9456_ ;
	wire _w9455_ ;
	wire _w9454_ ;
	wire _w9453_ ;
	wire _w9452_ ;
	wire _w9451_ ;
	wire _w9450_ ;
	wire _w9449_ ;
	wire _w9448_ ;
	wire _w9447_ ;
	wire _w9446_ ;
	wire _w9445_ ;
	wire _w9444_ ;
	wire _w9443_ ;
	wire _w9442_ ;
	wire _w9441_ ;
	wire _w9440_ ;
	wire _w9439_ ;
	wire _w9438_ ;
	wire _w9437_ ;
	wire _w9436_ ;
	wire _w9435_ ;
	wire _w9434_ ;
	wire _w9433_ ;
	wire _w9432_ ;
	wire _w9431_ ;
	wire _w9430_ ;
	wire _w9429_ ;
	wire _w9428_ ;
	wire _w9427_ ;
	wire _w9426_ ;
	wire _w9425_ ;
	wire _w9424_ ;
	wire _w9423_ ;
	wire _w9422_ ;
	wire _w9421_ ;
	wire _w9420_ ;
	wire _w9419_ ;
	wire _w9418_ ;
	wire _w9417_ ;
	wire _w9416_ ;
	wire _w9415_ ;
	wire _w9414_ ;
	wire _w9413_ ;
	wire _w9412_ ;
	wire _w9411_ ;
	wire _w9410_ ;
	wire _w9409_ ;
	wire _w9408_ ;
	wire _w9407_ ;
	wire _w9406_ ;
	wire _w9405_ ;
	wire _w9404_ ;
	wire _w9403_ ;
	wire _w9402_ ;
	wire _w9401_ ;
	wire _w9400_ ;
	wire _w9399_ ;
	wire _w9398_ ;
	wire _w9397_ ;
	wire _w9396_ ;
	wire _w9395_ ;
	wire _w9394_ ;
	wire _w9393_ ;
	wire _w9392_ ;
	wire _w9391_ ;
	wire _w9390_ ;
	wire _w9389_ ;
	wire _w9388_ ;
	wire _w9387_ ;
	wire _w9386_ ;
	wire _w9385_ ;
	wire _w9384_ ;
	wire _w9383_ ;
	wire _w9382_ ;
	wire _w9381_ ;
	wire _w9380_ ;
	wire _w9379_ ;
	wire _w9378_ ;
	wire _w9377_ ;
	wire _w9376_ ;
	wire _w9375_ ;
	wire _w9374_ ;
	wire _w9373_ ;
	wire _w9372_ ;
	wire _w9371_ ;
	wire _w9370_ ;
	wire _w9369_ ;
	wire _w9368_ ;
	wire _w9367_ ;
	wire _w9366_ ;
	wire _w9365_ ;
	wire _w9364_ ;
	wire _w9363_ ;
	wire _w9362_ ;
	wire _w9361_ ;
	wire _w9360_ ;
	wire _w9359_ ;
	wire _w9358_ ;
	wire _w9357_ ;
	wire _w9356_ ;
	wire _w9355_ ;
	wire _w9354_ ;
	wire _w9353_ ;
	wire _w9352_ ;
	wire _w9351_ ;
	wire _w9350_ ;
	wire _w9349_ ;
	wire _w9348_ ;
	wire _w9347_ ;
	wire _w9346_ ;
	wire _w9345_ ;
	wire _w9344_ ;
	wire _w9343_ ;
	wire _w9342_ ;
	wire _w9341_ ;
	wire _w9340_ ;
	wire _w9339_ ;
	wire _w9338_ ;
	wire _w9337_ ;
	wire _w9336_ ;
	wire _w9335_ ;
	wire _w9334_ ;
	wire _w9333_ ;
	wire _w9332_ ;
	wire _w9331_ ;
	wire _w9330_ ;
	wire _w9329_ ;
	wire _w9328_ ;
	wire _w9327_ ;
	wire _w9326_ ;
	wire _w9325_ ;
	wire _w9324_ ;
	wire _w9323_ ;
	wire _w9322_ ;
	wire _w9321_ ;
	wire _w9320_ ;
	wire _w9319_ ;
	wire _w9318_ ;
	wire _w9317_ ;
	wire _w9316_ ;
	wire _w9315_ ;
	wire _w9314_ ;
	wire _w9313_ ;
	wire _w9312_ ;
	wire _w9311_ ;
	wire _w9310_ ;
	wire _w9309_ ;
	wire _w9308_ ;
	wire _w9307_ ;
	wire _w9306_ ;
	wire _w9305_ ;
	wire _w9304_ ;
	wire _w9303_ ;
	wire _w9302_ ;
	wire _w9301_ ;
	wire _w9300_ ;
	wire _w9299_ ;
	wire _w9298_ ;
	wire _w9297_ ;
	wire _w9296_ ;
	wire _w9295_ ;
	wire _w9294_ ;
	wire _w9293_ ;
	wire _w9292_ ;
	wire _w9291_ ;
	wire _w9290_ ;
	wire _w9289_ ;
	wire _w9288_ ;
	wire _w9287_ ;
	wire _w9286_ ;
	wire _w9285_ ;
	wire _w9284_ ;
	wire _w9283_ ;
	wire _w9282_ ;
	wire _w9281_ ;
	wire _w9280_ ;
	wire _w9279_ ;
	wire _w9278_ ;
	wire _w9277_ ;
	wire _w9276_ ;
	wire _w9275_ ;
	wire _w9274_ ;
	wire _w9273_ ;
	wire _w9272_ ;
	wire _w9271_ ;
	wire _w9270_ ;
	wire _w9269_ ;
	wire _w9268_ ;
	wire _w9267_ ;
	wire _w9266_ ;
	wire _w9265_ ;
	wire _w9264_ ;
	wire _w9263_ ;
	wire _w9262_ ;
	wire _w9261_ ;
	wire _w9260_ ;
	wire _w9259_ ;
	wire _w9258_ ;
	wire _w9257_ ;
	wire _w9256_ ;
	wire _w9255_ ;
	wire _w9254_ ;
	wire _w9253_ ;
	wire _w9252_ ;
	wire _w9251_ ;
	wire _w9250_ ;
	wire _w9249_ ;
	wire _w9248_ ;
	wire _w9247_ ;
	wire _w9246_ ;
	wire _w9245_ ;
	wire _w9244_ ;
	wire _w9243_ ;
	wire _w9242_ ;
	wire _w9241_ ;
	wire _w9240_ ;
	wire _w9239_ ;
	wire _w9238_ ;
	wire _w9237_ ;
	wire _w9236_ ;
	wire _w9235_ ;
	wire _w9234_ ;
	wire _w9233_ ;
	wire _w9232_ ;
	wire _w9231_ ;
	wire _w9230_ ;
	wire _w9229_ ;
	wire _w9228_ ;
	wire _w9227_ ;
	wire _w9226_ ;
	wire _w9225_ ;
	wire _w9224_ ;
	wire _w9223_ ;
	wire _w9222_ ;
	wire _w9221_ ;
	wire _w9220_ ;
	wire _w9219_ ;
	wire _w9218_ ;
	wire _w9217_ ;
	wire _w9216_ ;
	wire _w9215_ ;
	wire _w9214_ ;
	wire _w9213_ ;
	wire _w9212_ ;
	wire _w9211_ ;
	wire _w9210_ ;
	wire _w9209_ ;
	wire _w9208_ ;
	wire _w9207_ ;
	wire _w9206_ ;
	wire _w9205_ ;
	wire _w9204_ ;
	wire _w9203_ ;
	wire _w9202_ ;
	wire _w9201_ ;
	wire _w9200_ ;
	wire _w9199_ ;
	wire _w9198_ ;
	wire _w9197_ ;
	wire _w9196_ ;
	wire _w9195_ ;
	wire _w9194_ ;
	wire _w9193_ ;
	wire _w9192_ ;
	wire _w9191_ ;
	wire _w9190_ ;
	wire _w9189_ ;
	wire _w9188_ ;
	wire _w9187_ ;
	wire _w9186_ ;
	wire _w9185_ ;
	wire _w9184_ ;
	wire _w9183_ ;
	wire _w9182_ ;
	wire _w9181_ ;
	wire _w9180_ ;
	wire _w9179_ ;
	wire _w9178_ ;
	wire _w9177_ ;
	wire _w9176_ ;
	wire _w9175_ ;
	wire _w9174_ ;
	wire _w9173_ ;
	wire _w9172_ ;
	wire _w9171_ ;
	wire _w9170_ ;
	wire _w9169_ ;
	wire _w9168_ ;
	wire _w9167_ ;
	wire _w9166_ ;
	wire _w9165_ ;
	wire _w9164_ ;
	wire _w9163_ ;
	wire _w9162_ ;
	wire _w9161_ ;
	wire _w9160_ ;
	wire _w9159_ ;
	wire _w9158_ ;
	wire _w9157_ ;
	wire _w9156_ ;
	wire _w9155_ ;
	wire _w9154_ ;
	wire _w9153_ ;
	wire _w9152_ ;
	wire _w9151_ ;
	wire _w9150_ ;
	wire _w9149_ ;
	wire _w9148_ ;
	wire _w9147_ ;
	wire _w9146_ ;
	wire _w9145_ ;
	wire _w9144_ ;
	wire _w9143_ ;
	wire _w9142_ ;
	wire _w9141_ ;
	wire _w9140_ ;
	wire _w9139_ ;
	wire _w9138_ ;
	wire _w9137_ ;
	wire _w9136_ ;
	wire _w9135_ ;
	wire _w9134_ ;
	wire _w9133_ ;
	wire _w9132_ ;
	wire _w9131_ ;
	wire _w9130_ ;
	wire _w9129_ ;
	wire _w9128_ ;
	wire _w9127_ ;
	wire _w9126_ ;
	wire _w9125_ ;
	wire _w9124_ ;
	wire _w9123_ ;
	wire _w9122_ ;
	wire _w9121_ ;
	wire _w9120_ ;
	wire _w9119_ ;
	wire _w9118_ ;
	wire _w9117_ ;
	wire _w9116_ ;
	wire _w9115_ ;
	wire _w9114_ ;
	wire _w9113_ ;
	wire _w9112_ ;
	wire _w9111_ ;
	wire _w9110_ ;
	wire _w9109_ ;
	wire _w9108_ ;
	wire _w9107_ ;
	wire _w9106_ ;
	wire _w9105_ ;
	wire _w9104_ ;
	wire _w9103_ ;
	wire _w9102_ ;
	wire _w9101_ ;
	wire _w9100_ ;
	wire _w9099_ ;
	wire _w9098_ ;
	wire _w9097_ ;
	wire _w9096_ ;
	wire _w9095_ ;
	wire _w9094_ ;
	wire _w9093_ ;
	wire _w9092_ ;
	wire _w9091_ ;
	wire _w9090_ ;
	wire _w9089_ ;
	wire _w9088_ ;
	wire _w9087_ ;
	wire _w9086_ ;
	wire _w9085_ ;
	wire _w9084_ ;
	wire _w9083_ ;
	wire _w9082_ ;
	wire _w9081_ ;
	wire _w9080_ ;
	wire _w9079_ ;
	wire _w9078_ ;
	wire _w9077_ ;
	wire _w9076_ ;
	wire _w9075_ ;
	wire _w9074_ ;
	wire _w9073_ ;
	wire _w9072_ ;
	wire _w9071_ ;
	wire _w9070_ ;
	wire _w9069_ ;
	wire _w9068_ ;
	wire _w9067_ ;
	wire _w9066_ ;
	wire _w9065_ ;
	wire _w9064_ ;
	wire _w9063_ ;
	wire _w9062_ ;
	wire _w9061_ ;
	wire _w9060_ ;
	wire _w9059_ ;
	wire _w9058_ ;
	wire _w9057_ ;
	wire _w9056_ ;
	wire _w9055_ ;
	wire _w9054_ ;
	wire _w9053_ ;
	wire _w9052_ ;
	wire _w9051_ ;
	wire _w9050_ ;
	wire _w9049_ ;
	wire _w9048_ ;
	wire _w9047_ ;
	wire _w9046_ ;
	wire _w9045_ ;
	wire _w9044_ ;
	wire _w9043_ ;
	wire _w9042_ ;
	wire _w9041_ ;
	wire _w9040_ ;
	wire _w9039_ ;
	wire _w9038_ ;
	wire _w9037_ ;
	wire _w9036_ ;
	wire _w9035_ ;
	wire _w9034_ ;
	wire _w9033_ ;
	wire _w9032_ ;
	wire _w9031_ ;
	wire _w9030_ ;
	wire _w9029_ ;
	wire _w9028_ ;
	wire _w9027_ ;
	wire _w9026_ ;
	wire _w9025_ ;
	wire _w9024_ ;
	wire _w9023_ ;
	wire _w9022_ ;
	wire _w9021_ ;
	wire _w9020_ ;
	wire _w9019_ ;
	wire _w9018_ ;
	wire _w9017_ ;
	wire _w9016_ ;
	wire _w9015_ ;
	wire _w9014_ ;
	wire _w9013_ ;
	wire _w9012_ ;
	wire _w9011_ ;
	wire _w9010_ ;
	wire _w9009_ ;
	wire _w9008_ ;
	wire _w9007_ ;
	wire _w9006_ ;
	wire _w9005_ ;
	wire _w9004_ ;
	wire _w9003_ ;
	wire _w9002_ ;
	wire _w9001_ ;
	wire _w9000_ ;
	wire _w8999_ ;
	wire _w8998_ ;
	wire _w8997_ ;
	wire _w8996_ ;
	wire _w8995_ ;
	wire _w8994_ ;
	wire _w8993_ ;
	wire _w8992_ ;
	wire _w8991_ ;
	wire _w8990_ ;
	wire _w8989_ ;
	wire _w8988_ ;
	wire _w8987_ ;
	wire _w8986_ ;
	wire _w8985_ ;
	wire _w8984_ ;
	wire _w8983_ ;
	wire _w8982_ ;
	wire _w8981_ ;
	wire _w8980_ ;
	wire _w8979_ ;
	wire _w8978_ ;
	wire _w8977_ ;
	wire _w8976_ ;
	wire _w8975_ ;
	wire _w8974_ ;
	wire _w8973_ ;
	wire _w8972_ ;
	wire _w8971_ ;
	wire _w8970_ ;
	wire _w8969_ ;
	wire _w8968_ ;
	wire _w8967_ ;
	wire _w8966_ ;
	wire _w8965_ ;
	wire _w8964_ ;
	wire _w8963_ ;
	wire _w8962_ ;
	wire _w8961_ ;
	wire _w8960_ ;
	wire _w8959_ ;
	wire _w8958_ ;
	wire _w8957_ ;
	wire _w8956_ ;
	wire _w8955_ ;
	wire _w8954_ ;
	wire _w8953_ ;
	wire _w8952_ ;
	wire _w8951_ ;
	wire _w8950_ ;
	wire _w8949_ ;
	wire _w8948_ ;
	wire _w8947_ ;
	wire _w8946_ ;
	wire _w8945_ ;
	wire _w8944_ ;
	wire _w8943_ ;
	wire _w8942_ ;
	wire _w8941_ ;
	wire _w8940_ ;
	wire _w8939_ ;
	wire _w8938_ ;
	wire _w8937_ ;
	wire _w8936_ ;
	wire _w8935_ ;
	wire _w8934_ ;
	wire _w8933_ ;
	wire _w8932_ ;
	wire _w8931_ ;
	wire _w8930_ ;
	wire _w8929_ ;
	wire _w8928_ ;
	wire _w8927_ ;
	wire _w8926_ ;
	wire _w8925_ ;
	wire _w8924_ ;
	wire _w8923_ ;
	wire _w8922_ ;
	wire _w8921_ ;
	wire _w8920_ ;
	wire _w8919_ ;
	wire _w8918_ ;
	wire _w8917_ ;
	wire _w8916_ ;
	wire _w8915_ ;
	wire _w8914_ ;
	wire _w8913_ ;
	wire _w8912_ ;
	wire _w8911_ ;
	wire _w8910_ ;
	wire _w8909_ ;
	wire _w8908_ ;
	wire _w8907_ ;
	wire _w8906_ ;
	wire _w8905_ ;
	wire _w8904_ ;
	wire _w8903_ ;
	wire _w8902_ ;
	wire _w8901_ ;
	wire _w8900_ ;
	wire _w8899_ ;
	wire _w8898_ ;
	wire _w8897_ ;
	wire _w8896_ ;
	wire _w8895_ ;
	wire _w8894_ ;
	wire _w8893_ ;
	wire _w8892_ ;
	wire _w8891_ ;
	wire _w8890_ ;
	wire _w8889_ ;
	wire _w8888_ ;
	wire _w8887_ ;
	wire _w8886_ ;
	wire _w8885_ ;
	wire _w8884_ ;
	wire _w8883_ ;
	wire _w8882_ ;
	wire _w8881_ ;
	wire _w8880_ ;
	wire _w8879_ ;
	wire _w8878_ ;
	wire _w8877_ ;
	wire _w8876_ ;
	wire _w8875_ ;
	wire _w8874_ ;
	wire _w8873_ ;
	wire _w8872_ ;
	wire _w8871_ ;
	wire _w8870_ ;
	wire _w8869_ ;
	wire _w8868_ ;
	wire _w8867_ ;
	wire _w8866_ ;
	wire _w8865_ ;
	wire _w8864_ ;
	wire _w8863_ ;
	wire _w8862_ ;
	wire _w8861_ ;
	wire _w8860_ ;
	wire _w8859_ ;
	wire _w8858_ ;
	wire _w8857_ ;
	wire _w8856_ ;
	wire _w8855_ ;
	wire _w8854_ ;
	wire _w8853_ ;
	wire _w8852_ ;
	wire _w8851_ ;
	wire _w8850_ ;
	wire _w8849_ ;
	wire _w8848_ ;
	wire _w8847_ ;
	wire _w8846_ ;
	wire _w8845_ ;
	wire _w8844_ ;
	wire _w8843_ ;
	wire _w8842_ ;
	wire _w8841_ ;
	wire _w8840_ ;
	wire _w8839_ ;
	wire _w8838_ ;
	wire _w8837_ ;
	wire _w8836_ ;
	wire _w8835_ ;
	wire _w8834_ ;
	wire _w8833_ ;
	wire _w8832_ ;
	wire _w8831_ ;
	wire _w8830_ ;
	wire _w8829_ ;
	wire _w8828_ ;
	wire _w8827_ ;
	wire _w8826_ ;
	wire _w8825_ ;
	wire _w8824_ ;
	wire _w8823_ ;
	wire _w8822_ ;
	wire _w8821_ ;
	wire _w8820_ ;
	wire _w8819_ ;
	wire _w8818_ ;
	wire _w8817_ ;
	wire _w8816_ ;
	wire _w8815_ ;
	wire _w8814_ ;
	wire _w8813_ ;
	wire _w8812_ ;
	wire _w8811_ ;
	wire _w8810_ ;
	wire _w8809_ ;
	wire _w8808_ ;
	wire _w8807_ ;
	wire _w8806_ ;
	wire _w8805_ ;
	wire _w8804_ ;
	wire _w8803_ ;
	wire _w8802_ ;
	wire _w8801_ ;
	wire _w8800_ ;
	wire _w8799_ ;
	wire _w8798_ ;
	wire _w8797_ ;
	wire _w8796_ ;
	wire _w8795_ ;
	wire _w8794_ ;
	wire _w8793_ ;
	wire _w8792_ ;
	wire _w8791_ ;
	wire _w8790_ ;
	wire _w8789_ ;
	wire _w8788_ ;
	wire _w8787_ ;
	wire _w8786_ ;
	wire _w8785_ ;
	wire _w8784_ ;
	wire _w8783_ ;
	wire _w8782_ ;
	wire _w8781_ ;
	wire _w8780_ ;
	wire _w8779_ ;
	wire _w8778_ ;
	wire _w8777_ ;
	wire _w8776_ ;
	wire _w8775_ ;
	wire _w8774_ ;
	wire _w8773_ ;
	wire _w8772_ ;
	wire _w8771_ ;
	wire _w8770_ ;
	wire _w8769_ ;
	wire _w8768_ ;
	wire _w8767_ ;
	wire _w8766_ ;
	wire _w8765_ ;
	wire _w8764_ ;
	wire _w8763_ ;
	wire _w8762_ ;
	wire _w8761_ ;
	wire _w8760_ ;
	wire _w8759_ ;
	wire _w8758_ ;
	wire _w8757_ ;
	wire _w8756_ ;
	wire _w8755_ ;
	wire _w8754_ ;
	wire _w8753_ ;
	wire _w8752_ ;
	wire _w8751_ ;
	wire _w8750_ ;
	wire _w8749_ ;
	wire _w8748_ ;
	wire _w8747_ ;
	wire _w8746_ ;
	wire _w8745_ ;
	wire _w8744_ ;
	wire _w8743_ ;
	wire _w8742_ ;
	wire _w8741_ ;
	wire _w8740_ ;
	wire _w8739_ ;
	wire _w8738_ ;
	wire _w8737_ ;
	wire _w8736_ ;
	wire _w8735_ ;
	wire _w8734_ ;
	wire _w8733_ ;
	wire _w8732_ ;
	wire _w8731_ ;
	wire _w8730_ ;
	wire _w8729_ ;
	wire _w8728_ ;
	wire _w8727_ ;
	wire _w8726_ ;
	wire _w8725_ ;
	wire _w8724_ ;
	wire _w8723_ ;
	wire _w8722_ ;
	wire _w8721_ ;
	wire _w8720_ ;
	wire _w8719_ ;
	wire _w8718_ ;
	wire _w8717_ ;
	wire _w8716_ ;
	wire _w8715_ ;
	wire _w8714_ ;
	wire _w8713_ ;
	wire _w8712_ ;
	wire _w8711_ ;
	wire _w8710_ ;
	wire _w8709_ ;
	wire _w8708_ ;
	wire _w8707_ ;
	wire _w8706_ ;
	wire _w8705_ ;
	wire _w8704_ ;
	wire _w8703_ ;
	wire _w8702_ ;
	wire _w8701_ ;
	wire _w8700_ ;
	wire _w8699_ ;
	wire _w8698_ ;
	wire _w8697_ ;
	wire _w8696_ ;
	wire _w8695_ ;
	wire _w8694_ ;
	wire _w8693_ ;
	wire _w8692_ ;
	wire _w8691_ ;
	wire _w8690_ ;
	wire _w8689_ ;
	wire _w8688_ ;
	wire _w8687_ ;
	wire _w8686_ ;
	wire _w8685_ ;
	wire _w8684_ ;
	wire _w8683_ ;
	wire _w8682_ ;
	wire _w8681_ ;
	wire _w8680_ ;
	wire _w8679_ ;
	wire _w8678_ ;
	wire _w8677_ ;
	wire _w8676_ ;
	wire _w8675_ ;
	wire _w8674_ ;
	wire _w8673_ ;
	wire _w8672_ ;
	wire _w8671_ ;
	wire _w8670_ ;
	wire _w8669_ ;
	wire _w8668_ ;
	wire _w8667_ ;
	wire _w8666_ ;
	wire _w8665_ ;
	wire _w8664_ ;
	wire _w8663_ ;
	wire _w8662_ ;
	wire _w8661_ ;
	wire _w8660_ ;
	wire _w8659_ ;
	wire _w8658_ ;
	wire _w8657_ ;
	wire _w8656_ ;
	wire _w8655_ ;
	wire _w8654_ ;
	wire _w8653_ ;
	wire _w8652_ ;
	wire _w8651_ ;
	wire _w8650_ ;
	wire _w8649_ ;
	wire _w8648_ ;
	wire _w8647_ ;
	wire _w8646_ ;
	wire _w8645_ ;
	wire _w8644_ ;
	wire _w8643_ ;
	wire _w8642_ ;
	wire _w8641_ ;
	wire _w8640_ ;
	wire _w8639_ ;
	wire _w8638_ ;
	wire _w8637_ ;
	wire _w8636_ ;
	wire _w8635_ ;
	wire _w8634_ ;
	wire _w8633_ ;
	wire _w8632_ ;
	wire _w8631_ ;
	wire _w8630_ ;
	wire _w8629_ ;
	wire _w8628_ ;
	wire _w8627_ ;
	wire _w8626_ ;
	wire _w8625_ ;
	wire _w8624_ ;
	wire _w8623_ ;
	wire _w8622_ ;
	wire _w8621_ ;
	wire _w8620_ ;
	wire _w8619_ ;
	wire _w8618_ ;
	wire _w8617_ ;
	wire _w8616_ ;
	wire _w8615_ ;
	wire _w8614_ ;
	wire _w8613_ ;
	wire _w8612_ ;
	wire _w8611_ ;
	wire _w8610_ ;
	wire _w8609_ ;
	wire _w8608_ ;
	wire _w8607_ ;
	wire _w8606_ ;
	wire _w8605_ ;
	wire _w8604_ ;
	wire _w8603_ ;
	wire _w8602_ ;
	wire _w8601_ ;
	wire _w8600_ ;
	wire _w8599_ ;
	wire _w8598_ ;
	wire _w8597_ ;
	wire _w8596_ ;
	wire _w8595_ ;
	wire _w8594_ ;
	wire _w8593_ ;
	wire _w8592_ ;
	wire _w8591_ ;
	wire _w8590_ ;
	wire _w8589_ ;
	wire _w8588_ ;
	wire _w8587_ ;
	wire _w8586_ ;
	wire _w8585_ ;
	wire _w8584_ ;
	wire _w8583_ ;
	wire _w8582_ ;
	wire _w8581_ ;
	wire _w8580_ ;
	wire _w8579_ ;
	wire _w8578_ ;
	wire _w8577_ ;
	wire _w8576_ ;
	wire _w8575_ ;
	wire _w8574_ ;
	wire _w8573_ ;
	wire _w8572_ ;
	wire _w8571_ ;
	wire _w8570_ ;
	wire _w8569_ ;
	wire _w8568_ ;
	wire _w8567_ ;
	wire _w8566_ ;
	wire _w8565_ ;
	wire _w8564_ ;
	wire _w8563_ ;
	wire _w8562_ ;
	wire _w8561_ ;
	wire _w8560_ ;
	wire _w8559_ ;
	wire _w8558_ ;
	wire _w8557_ ;
	wire _w8556_ ;
	wire _w8555_ ;
	wire _w8554_ ;
	wire _w8553_ ;
	wire _w8552_ ;
	wire _w8551_ ;
	wire _w8550_ ;
	wire _w8549_ ;
	wire _w8548_ ;
	wire _w8547_ ;
	wire _w8546_ ;
	wire _w8545_ ;
	wire _w8544_ ;
	wire _w8543_ ;
	wire _w8542_ ;
	wire _w8541_ ;
	wire _w8540_ ;
	wire _w8539_ ;
	wire _w8538_ ;
	wire _w8537_ ;
	wire _w8536_ ;
	wire _w8535_ ;
	wire _w8534_ ;
	wire _w8533_ ;
	wire _w8532_ ;
	wire _w8531_ ;
	wire _w8530_ ;
	wire _w8529_ ;
	wire _w8528_ ;
	wire _w8527_ ;
	wire _w8526_ ;
	wire _w8525_ ;
	wire _w8524_ ;
	wire _w8523_ ;
	wire _w8522_ ;
	wire _w8521_ ;
	wire _w8520_ ;
	wire _w8519_ ;
	wire _w8518_ ;
	wire _w8517_ ;
	wire _w8516_ ;
	wire _w8515_ ;
	wire _w8514_ ;
	wire _w8513_ ;
	wire _w8512_ ;
	wire _w8511_ ;
	wire _w8510_ ;
	wire _w8509_ ;
	wire _w8508_ ;
	wire _w8507_ ;
	wire _w8506_ ;
	wire _w8505_ ;
	wire _w8504_ ;
	wire _w8503_ ;
	wire _w8502_ ;
	wire _w8501_ ;
	wire _w8500_ ;
	wire _w8499_ ;
	wire _w8498_ ;
	wire _w8497_ ;
	wire _w8496_ ;
	wire _w8495_ ;
	wire _w8494_ ;
	wire _w8493_ ;
	wire _w8492_ ;
	wire _w8491_ ;
	wire _w8490_ ;
	wire _w8489_ ;
	wire _w8488_ ;
	wire _w8487_ ;
	wire _w8486_ ;
	wire _w8485_ ;
	wire _w8484_ ;
	wire _w8483_ ;
	wire _w8482_ ;
	wire _w8481_ ;
	wire _w8480_ ;
	wire _w8479_ ;
	wire _w8478_ ;
	wire _w8477_ ;
	wire _w8476_ ;
	wire _w8475_ ;
	wire _w8474_ ;
	wire _w8473_ ;
	wire _w8472_ ;
	wire _w8471_ ;
	wire _w8470_ ;
	wire _w8469_ ;
	wire _w8468_ ;
	wire _w8467_ ;
	wire _w8466_ ;
	wire _w8465_ ;
	wire _w8464_ ;
	wire _w8463_ ;
	wire _w8462_ ;
	wire _w8461_ ;
	wire _w8460_ ;
	wire _w8459_ ;
	wire _w8458_ ;
	wire _w8457_ ;
	wire _w8456_ ;
	wire _w8455_ ;
	wire _w8454_ ;
	wire _w8453_ ;
	wire _w8452_ ;
	wire _w8451_ ;
	wire _w8450_ ;
	wire _w8449_ ;
	wire _w8448_ ;
	wire _w8447_ ;
	wire _w8446_ ;
	wire _w8445_ ;
	wire _w8444_ ;
	wire _w8443_ ;
	wire _w8442_ ;
	wire _w8441_ ;
	wire _w8440_ ;
	wire _w8439_ ;
	wire _w8438_ ;
	wire _w8437_ ;
	wire _w8436_ ;
	wire _w8435_ ;
	wire _w8434_ ;
	wire _w8433_ ;
	wire _w8432_ ;
	wire _w8431_ ;
	wire _w8430_ ;
	wire _w8429_ ;
	wire _w8428_ ;
	wire _w8427_ ;
	wire _w8426_ ;
	wire _w8425_ ;
	wire _w8424_ ;
	wire _w8423_ ;
	wire _w8422_ ;
	wire _w8421_ ;
	wire _w8420_ ;
	wire _w8419_ ;
	wire _w8418_ ;
	wire _w8417_ ;
	wire _w8416_ ;
	wire _w8415_ ;
	wire _w8414_ ;
	wire _w8413_ ;
	wire _w8412_ ;
	wire _w8411_ ;
	wire _w8410_ ;
	wire _w8409_ ;
	wire _w8408_ ;
	wire _w8407_ ;
	wire _w8406_ ;
	wire _w8405_ ;
	wire _w8404_ ;
	wire _w8403_ ;
	wire _w8402_ ;
	wire _w8401_ ;
	wire _w8400_ ;
	wire _w8399_ ;
	wire _w8398_ ;
	wire _w8397_ ;
	wire _w8396_ ;
	wire _w8395_ ;
	wire _w8394_ ;
	wire _w8393_ ;
	wire _w8392_ ;
	wire _w8391_ ;
	wire _w8390_ ;
	wire _w8389_ ;
	wire _w8388_ ;
	wire _w8387_ ;
	wire _w8386_ ;
	wire _w8385_ ;
	wire _w8384_ ;
	wire _w8383_ ;
	wire _w8382_ ;
	wire _w8381_ ;
	wire _w8380_ ;
	wire _w8379_ ;
	wire _w8378_ ;
	wire _w8377_ ;
	wire _w8376_ ;
	wire _w8375_ ;
	wire _w8374_ ;
	wire _w8373_ ;
	wire _w8372_ ;
	wire _w8371_ ;
	wire _w8370_ ;
	wire _w8369_ ;
	wire _w8368_ ;
	wire _w8367_ ;
	wire _w8366_ ;
	wire _w8365_ ;
	wire _w8364_ ;
	wire _w8363_ ;
	wire _w8362_ ;
	wire _w8361_ ;
	wire _w8360_ ;
	wire _w8359_ ;
	wire _w8358_ ;
	wire _w8357_ ;
	wire _w8356_ ;
	wire _w8355_ ;
	wire _w8354_ ;
	wire _w8353_ ;
	wire _w8352_ ;
	wire _w8351_ ;
	wire _w8350_ ;
	wire _w8349_ ;
	wire _w8348_ ;
	wire _w8347_ ;
	wire _w8346_ ;
	wire _w8345_ ;
	wire _w8344_ ;
	wire _w8343_ ;
	wire _w8342_ ;
	wire _w8341_ ;
	wire _w8340_ ;
	wire _w8339_ ;
	wire _w8338_ ;
	wire _w8337_ ;
	wire _w8336_ ;
	wire _w8335_ ;
	wire _w8334_ ;
	wire _w8333_ ;
	wire _w8332_ ;
	wire _w8331_ ;
	wire _w8330_ ;
	wire _w8329_ ;
	wire _w8328_ ;
	wire _w8327_ ;
	wire _w8326_ ;
	wire _w8325_ ;
	wire _w8324_ ;
	wire _w8323_ ;
	wire _w8322_ ;
	wire _w8321_ ;
	wire _w8320_ ;
	wire _w8319_ ;
	wire _w8318_ ;
	wire _w8317_ ;
	wire _w8316_ ;
	wire _w8315_ ;
	wire _w8314_ ;
	wire _w8313_ ;
	wire _w8312_ ;
	wire _w8311_ ;
	wire _w8310_ ;
	wire _w8309_ ;
	wire _w8308_ ;
	wire _w8307_ ;
	wire _w8306_ ;
	wire _w8305_ ;
	wire _w8304_ ;
	wire _w8303_ ;
	wire _w8302_ ;
	wire _w8301_ ;
	wire _w8300_ ;
	wire _w8299_ ;
	wire _w8298_ ;
	wire _w8297_ ;
	wire _w8296_ ;
	wire _w8295_ ;
	wire _w8294_ ;
	wire _w8293_ ;
	wire _w8292_ ;
	wire _w8291_ ;
	wire _w8290_ ;
	wire _w8289_ ;
	wire _w8288_ ;
	wire _w8287_ ;
	wire _w8286_ ;
	wire _w8285_ ;
	wire _w8284_ ;
	wire _w8283_ ;
	wire _w8282_ ;
	wire _w8281_ ;
	wire _w8280_ ;
	wire _w8279_ ;
	wire _w8278_ ;
	wire _w8277_ ;
	wire _w8276_ ;
	wire _w8275_ ;
	wire _w8274_ ;
	wire _w8273_ ;
	wire _w8272_ ;
	wire _w8271_ ;
	wire _w8270_ ;
	wire _w8269_ ;
	wire _w8268_ ;
	wire _w8267_ ;
	wire _w8266_ ;
	wire _w8265_ ;
	wire _w8264_ ;
	wire _w8263_ ;
	wire _w8262_ ;
	wire _w8261_ ;
	wire _w8260_ ;
	wire _w8259_ ;
	wire _w8258_ ;
	wire _w8257_ ;
	wire _w8256_ ;
	wire _w8255_ ;
	wire _w8254_ ;
	wire _w8253_ ;
	wire _w8252_ ;
	wire _w8251_ ;
	wire _w8250_ ;
	wire _w8249_ ;
	wire _w8248_ ;
	wire _w8247_ ;
	wire _w8246_ ;
	wire _w8245_ ;
	wire _w8244_ ;
	wire _w8243_ ;
	wire _w8242_ ;
	wire _w8241_ ;
	wire _w8240_ ;
	wire _w8239_ ;
	wire _w8238_ ;
	wire _w8237_ ;
	wire _w8236_ ;
	wire _w8235_ ;
	wire _w8234_ ;
	wire _w8233_ ;
	wire _w8232_ ;
	wire _w8231_ ;
	wire _w8230_ ;
	wire _w8229_ ;
	wire _w8228_ ;
	wire _w8227_ ;
	wire _w8226_ ;
	wire _w8225_ ;
	wire _w8224_ ;
	wire _w8223_ ;
	wire _w8222_ ;
	wire _w8221_ ;
	wire _w8220_ ;
	wire _w8219_ ;
	wire _w8218_ ;
	wire _w8217_ ;
	wire _w8216_ ;
	wire _w8215_ ;
	wire _w8214_ ;
	wire _w8213_ ;
	wire _w8212_ ;
	wire _w8211_ ;
	wire _w8210_ ;
	wire _w8209_ ;
	wire _w8208_ ;
	wire _w8207_ ;
	wire _w8206_ ;
	wire _w8205_ ;
	wire _w8204_ ;
	wire _w8203_ ;
	wire _w8202_ ;
	wire _w8201_ ;
	wire _w8200_ ;
	wire _w8199_ ;
	wire _w8198_ ;
	wire _w8197_ ;
	wire _w8196_ ;
	wire _w8195_ ;
	wire _w8194_ ;
	wire _w8193_ ;
	wire _w8192_ ;
	wire _w8191_ ;
	wire _w8190_ ;
	wire _w8189_ ;
	wire _w8188_ ;
	wire _w8187_ ;
	wire _w8186_ ;
	wire _w8185_ ;
	wire _w8184_ ;
	wire _w8183_ ;
	wire _w8182_ ;
	wire _w8181_ ;
	wire _w8180_ ;
	wire _w8179_ ;
	wire _w8178_ ;
	wire _w8177_ ;
	wire _w8176_ ;
	wire _w8175_ ;
	wire _w8174_ ;
	wire _w8173_ ;
	wire _w8172_ ;
	wire _w8171_ ;
	wire _w8170_ ;
	wire _w8169_ ;
	wire _w8168_ ;
	wire _w8167_ ;
	wire _w8166_ ;
	wire _w8165_ ;
	wire _w8164_ ;
	wire _w8163_ ;
	wire _w8162_ ;
	wire _w8161_ ;
	wire _w8160_ ;
	wire _w8159_ ;
	wire _w8158_ ;
	wire _w8157_ ;
	wire _w8156_ ;
	wire _w8155_ ;
	wire _w8154_ ;
	wire _w8153_ ;
	wire _w8152_ ;
	wire _w8151_ ;
	wire _w8150_ ;
	wire _w8149_ ;
	wire _w8148_ ;
	wire _w8147_ ;
	wire _w8146_ ;
	wire _w8145_ ;
	wire _w8144_ ;
	wire _w8143_ ;
	wire _w8142_ ;
	wire _w8141_ ;
	wire _w8140_ ;
	wire _w8139_ ;
	wire _w8138_ ;
	wire _w8137_ ;
	wire _w8136_ ;
	wire _w8135_ ;
	wire _w8134_ ;
	wire _w8133_ ;
	wire _w8132_ ;
	wire _w8131_ ;
	wire _w8130_ ;
	wire _w8129_ ;
	wire _w8128_ ;
	wire _w8127_ ;
	wire _w8126_ ;
	wire _w8125_ ;
	wire _w8124_ ;
	wire _w8123_ ;
	wire _w8122_ ;
	wire _w8121_ ;
	wire _w8120_ ;
	wire _w8119_ ;
	wire _w8118_ ;
	wire _w8117_ ;
	wire _w8116_ ;
	wire _w8115_ ;
	wire _w8114_ ;
	wire _w8113_ ;
	wire _w8112_ ;
	wire _w8111_ ;
	wire _w8110_ ;
	wire _w8109_ ;
	wire _w8108_ ;
	wire _w8107_ ;
	wire _w8106_ ;
	wire _w8105_ ;
	wire _w8104_ ;
	wire _w8103_ ;
	wire _w8102_ ;
	wire _w8101_ ;
	wire _w8100_ ;
	wire _w8099_ ;
	wire _w8098_ ;
	wire _w8097_ ;
	wire _w8096_ ;
	wire _w8095_ ;
	wire _w8094_ ;
	wire _w8093_ ;
	wire _w8092_ ;
	wire _w8091_ ;
	wire _w8090_ ;
	wire _w8089_ ;
	wire _w8088_ ;
	wire _w8087_ ;
	wire _w8086_ ;
	wire _w8085_ ;
	wire _w8084_ ;
	wire _w8083_ ;
	wire _w8082_ ;
	wire _w8081_ ;
	wire _w8080_ ;
	wire _w8079_ ;
	wire _w8078_ ;
	wire _w8077_ ;
	wire _w8076_ ;
	wire _w8075_ ;
	wire _w8074_ ;
	wire _w8073_ ;
	wire _w8072_ ;
	wire _w8071_ ;
	wire _w8070_ ;
	wire _w8069_ ;
	wire _w8068_ ;
	wire _w8067_ ;
	wire _w8066_ ;
	wire _w8065_ ;
	wire _w8064_ ;
	wire _w8063_ ;
	wire _w8062_ ;
	wire _w8061_ ;
	wire _w8060_ ;
	wire _w8059_ ;
	wire _w8058_ ;
	wire _w8057_ ;
	wire _w8056_ ;
	wire _w8055_ ;
	wire _w8054_ ;
	wire _w8053_ ;
	wire _w8052_ ;
	wire _w8051_ ;
	wire _w8050_ ;
	wire _w8049_ ;
	wire _w8048_ ;
	wire _w8047_ ;
	wire _w8046_ ;
	wire _w8045_ ;
	wire _w8044_ ;
	wire _w8043_ ;
	wire _w8042_ ;
	wire _w8041_ ;
	wire _w8040_ ;
	wire _w8039_ ;
	wire _w8038_ ;
	wire _w8037_ ;
	wire _w8036_ ;
	wire _w8035_ ;
	wire _w8034_ ;
	wire _w8033_ ;
	wire _w8032_ ;
	wire _w8031_ ;
	wire _w8030_ ;
	wire _w8029_ ;
	wire _w8028_ ;
	wire _w8027_ ;
	wire _w8026_ ;
	wire _w8025_ ;
	wire _w8024_ ;
	wire _w8023_ ;
	wire _w8022_ ;
	wire _w8021_ ;
	wire _w8020_ ;
	wire _w8019_ ;
	wire _w8018_ ;
	wire _w8017_ ;
	wire _w8016_ ;
	wire _w8015_ ;
	wire _w8014_ ;
	wire _w8013_ ;
	wire _w8012_ ;
	wire _w8011_ ;
	wire _w8010_ ;
	wire _w8009_ ;
	wire _w8008_ ;
	wire _w8007_ ;
	wire _w8006_ ;
	wire _w8005_ ;
	wire _w8004_ ;
	wire _w8003_ ;
	wire _w8002_ ;
	wire _w8001_ ;
	wire _w8000_ ;
	wire _w7999_ ;
	wire _w7998_ ;
	wire _w7997_ ;
	wire _w7996_ ;
	wire _w7995_ ;
	wire _w7994_ ;
	wire _w7993_ ;
	wire _w7992_ ;
	wire _w7991_ ;
	wire _w7990_ ;
	wire _w7989_ ;
	wire _w7988_ ;
	wire _w7987_ ;
	wire _w7986_ ;
	wire _w7985_ ;
	wire _w7984_ ;
	wire _w7983_ ;
	wire _w7982_ ;
	wire _w7981_ ;
	wire _w7980_ ;
	wire _w7979_ ;
	wire _w7978_ ;
	wire _w7977_ ;
	wire _w7976_ ;
	wire _w7975_ ;
	wire _w7974_ ;
	wire _w7973_ ;
	wire _w7972_ ;
	wire _w7971_ ;
	wire _w7970_ ;
	wire _w7969_ ;
	wire _w7968_ ;
	wire _w7967_ ;
	wire _w7966_ ;
	wire _w7965_ ;
	wire _w7964_ ;
	wire _w7963_ ;
	wire _w7962_ ;
	wire _w7961_ ;
	wire _w7960_ ;
	wire _w7959_ ;
	wire _w7958_ ;
	wire _w7957_ ;
	wire _w7956_ ;
	wire _w7955_ ;
	wire _w7954_ ;
	wire _w7953_ ;
	wire _w7952_ ;
	wire _w7951_ ;
	wire _w7950_ ;
	wire _w7949_ ;
	wire _w7948_ ;
	wire _w7947_ ;
	wire _w7946_ ;
	wire _w7945_ ;
	wire _w7944_ ;
	wire _w7943_ ;
	wire _w7942_ ;
	wire _w7941_ ;
	wire _w7940_ ;
	wire _w7939_ ;
	wire _w7938_ ;
	wire _w7937_ ;
	wire _w7936_ ;
	wire _w7935_ ;
	wire _w7934_ ;
	wire _w7933_ ;
	wire _w7932_ ;
	wire _w7931_ ;
	wire _w7930_ ;
	wire _w7929_ ;
	wire _w7928_ ;
	wire _w7927_ ;
	wire _w7926_ ;
	wire _w7925_ ;
	wire _w7924_ ;
	wire _w7923_ ;
	wire _w7922_ ;
	wire _w7921_ ;
	wire _w7920_ ;
	wire _w7919_ ;
	wire _w7918_ ;
	wire _w7917_ ;
	wire _w7916_ ;
	wire _w7915_ ;
	wire _w7914_ ;
	wire _w7913_ ;
	wire _w7912_ ;
	wire _w7911_ ;
	wire _w7910_ ;
	wire _w7909_ ;
	wire _w7908_ ;
	wire _w7907_ ;
	wire _w7906_ ;
	wire _w7905_ ;
	wire _w7904_ ;
	wire _w7903_ ;
	wire _w7902_ ;
	wire _w7901_ ;
	wire _w7900_ ;
	wire _w7899_ ;
	wire _w7898_ ;
	wire _w7897_ ;
	wire _w7896_ ;
	wire _w7895_ ;
	wire _w7894_ ;
	wire _w7893_ ;
	wire _w7892_ ;
	wire _w7891_ ;
	wire _w7890_ ;
	wire _w7889_ ;
	wire _w7888_ ;
	wire _w7887_ ;
	wire _w7886_ ;
	wire _w7885_ ;
	wire _w7884_ ;
	wire _w7883_ ;
	wire _w7882_ ;
	wire _w7881_ ;
	wire _w7880_ ;
	wire _w7879_ ;
	wire _w7878_ ;
	wire _w7877_ ;
	wire _w7876_ ;
	wire _w7875_ ;
	wire _w7874_ ;
	wire _w7873_ ;
	wire _w7872_ ;
	wire _w7871_ ;
	wire _w7870_ ;
	wire _w7869_ ;
	wire _w7868_ ;
	wire _w7867_ ;
	wire _w7866_ ;
	wire _w7865_ ;
	wire _w7864_ ;
	wire _w7863_ ;
	wire _w7862_ ;
	wire _w7861_ ;
	wire _w7860_ ;
	wire _w7859_ ;
	wire _w7858_ ;
	wire _w7857_ ;
	wire _w7856_ ;
	wire _w7855_ ;
	wire _w7854_ ;
	wire _w7853_ ;
	wire _w7852_ ;
	wire _w7851_ ;
	wire _w7850_ ;
	wire _w7849_ ;
	wire _w7848_ ;
	wire _w7847_ ;
	wire _w7846_ ;
	wire _w7845_ ;
	wire _w7844_ ;
	wire _w7843_ ;
	wire _w7842_ ;
	wire _w7841_ ;
	wire _w7840_ ;
	wire _w7839_ ;
	wire _w7838_ ;
	wire _w7837_ ;
	wire _w7836_ ;
	wire _w7835_ ;
	wire _w7834_ ;
	wire _w7833_ ;
	wire _w7832_ ;
	wire _w7831_ ;
	wire _w7830_ ;
	wire _w7829_ ;
	wire _w7828_ ;
	wire _w7827_ ;
	wire _w7826_ ;
	wire _w7825_ ;
	wire _w7824_ ;
	wire _w7823_ ;
	wire _w7822_ ;
	wire _w7821_ ;
	wire _w7820_ ;
	wire _w7819_ ;
	wire _w7818_ ;
	wire _w7817_ ;
	wire _w7816_ ;
	wire _w7815_ ;
	wire _w7814_ ;
	wire _w7813_ ;
	wire _w7812_ ;
	wire _w7811_ ;
	wire _w7810_ ;
	wire _w7809_ ;
	wire _w7808_ ;
	wire _w7807_ ;
	wire _w7806_ ;
	wire _w7805_ ;
	wire _w7804_ ;
	wire _w7803_ ;
	wire _w7802_ ;
	wire _w7801_ ;
	wire _w7800_ ;
	wire _w7799_ ;
	wire _w7798_ ;
	wire _w7797_ ;
	wire _w7796_ ;
	wire _w7795_ ;
	wire _w7794_ ;
	wire _w7793_ ;
	wire _w7792_ ;
	wire _w7791_ ;
	wire _w7790_ ;
	wire _w7789_ ;
	wire _w7788_ ;
	wire _w7787_ ;
	wire _w7786_ ;
	wire _w7785_ ;
	wire _w7784_ ;
	wire _w7783_ ;
	wire _w7782_ ;
	wire _w7781_ ;
	wire _w7780_ ;
	wire _w7779_ ;
	wire _w7778_ ;
	wire _w7777_ ;
	wire _w7776_ ;
	wire _w7775_ ;
	wire _w7774_ ;
	wire _w7773_ ;
	wire _w7772_ ;
	wire _w7771_ ;
	wire _w7770_ ;
	wire _w7769_ ;
	wire _w7768_ ;
	wire _w7767_ ;
	wire _w7766_ ;
	wire _w7765_ ;
	wire _w7764_ ;
	wire _w7763_ ;
	wire _w7762_ ;
	wire _w7761_ ;
	wire _w7760_ ;
	wire _w7759_ ;
	wire _w7758_ ;
	wire _w7757_ ;
	wire _w7756_ ;
	wire _w7755_ ;
	wire _w7754_ ;
	wire _w7753_ ;
	wire _w7752_ ;
	wire _w7751_ ;
	wire _w7750_ ;
	wire _w7749_ ;
	wire _w7748_ ;
	wire _w7747_ ;
	wire _w7746_ ;
	wire _w7745_ ;
	wire _w7744_ ;
	wire _w7743_ ;
	wire _w7742_ ;
	wire _w7741_ ;
	wire _w7740_ ;
	wire _w7739_ ;
	wire _w7738_ ;
	wire _w7737_ ;
	wire _w7736_ ;
	wire _w7735_ ;
	wire _w7734_ ;
	wire _w7733_ ;
	wire _w7732_ ;
	wire _w7731_ ;
	wire _w7730_ ;
	wire _w7729_ ;
	wire _w7728_ ;
	wire _w7727_ ;
	wire _w7726_ ;
	wire _w7725_ ;
	wire _w7724_ ;
	wire _w7723_ ;
	wire _w7722_ ;
	wire _w7721_ ;
	wire _w7720_ ;
	wire _w7719_ ;
	wire _w7718_ ;
	wire _w7717_ ;
	wire _w7716_ ;
	wire _w7715_ ;
	wire _w7714_ ;
	wire _w7713_ ;
	wire _w7712_ ;
	wire _w7711_ ;
	wire _w7710_ ;
	wire _w7709_ ;
	wire _w7708_ ;
	wire _w7707_ ;
	wire _w7706_ ;
	wire _w7705_ ;
	wire _w7704_ ;
	wire _w7703_ ;
	wire _w7702_ ;
	wire _w7701_ ;
	wire _w7700_ ;
	wire _w7699_ ;
	wire _w7698_ ;
	wire _w7697_ ;
	wire _w7696_ ;
	wire _w7695_ ;
	wire _w7694_ ;
	wire _w7693_ ;
	wire _w7692_ ;
	wire _w7691_ ;
	wire _w7690_ ;
	wire _w7689_ ;
	wire _w7688_ ;
	wire _w7687_ ;
	wire _w7686_ ;
	wire _w7685_ ;
	wire _w7684_ ;
	wire _w7683_ ;
	wire _w7682_ ;
	wire _w7681_ ;
	wire _w7680_ ;
	wire _w7679_ ;
	wire _w7678_ ;
	wire _w7677_ ;
	wire _w7676_ ;
	wire _w7675_ ;
	wire _w7674_ ;
	wire _w7673_ ;
	wire _w7672_ ;
	wire _w7671_ ;
	wire _w7670_ ;
	wire _w7669_ ;
	wire _w7668_ ;
	wire _w7667_ ;
	wire _w7666_ ;
	wire _w7665_ ;
	wire _w7664_ ;
	wire _w7663_ ;
	wire _w7662_ ;
	wire _w7661_ ;
	wire _w7660_ ;
	wire _w7659_ ;
	wire _w7658_ ;
	wire _w7657_ ;
	wire _w7656_ ;
	wire _w7655_ ;
	wire _w7654_ ;
	wire _w7653_ ;
	wire _w7652_ ;
	wire _w7651_ ;
	wire _w7650_ ;
	wire _w7649_ ;
	wire _w7648_ ;
	wire _w7647_ ;
	wire _w7646_ ;
	wire _w7645_ ;
	wire _w7644_ ;
	wire _w7643_ ;
	wire _w7642_ ;
	wire _w7641_ ;
	wire _w7640_ ;
	wire _w7639_ ;
	wire _w7638_ ;
	wire _w7637_ ;
	wire _w7636_ ;
	wire _w7635_ ;
	wire _w7634_ ;
	wire _w7633_ ;
	wire _w7632_ ;
	wire _w7631_ ;
	wire _w7630_ ;
	wire _w7629_ ;
	wire _w7628_ ;
	wire _w7627_ ;
	wire _w7626_ ;
	wire _w7625_ ;
	wire _w7624_ ;
	wire _w7623_ ;
	wire _w7622_ ;
	wire _w7621_ ;
	wire _w7620_ ;
	wire _w7619_ ;
	wire _w7618_ ;
	wire _w7617_ ;
	wire _w7616_ ;
	wire _w7615_ ;
	wire _w7614_ ;
	wire _w7613_ ;
	wire _w7612_ ;
	wire _w7611_ ;
	wire _w7610_ ;
	wire _w7609_ ;
	wire _w7608_ ;
	wire _w7607_ ;
	wire _w7606_ ;
	wire _w7605_ ;
	wire _w7604_ ;
	wire _w7603_ ;
	wire _w7602_ ;
	wire _w7601_ ;
	wire _w7600_ ;
	wire _w7599_ ;
	wire _w7598_ ;
	wire _w7597_ ;
	wire _w7596_ ;
	wire _w7595_ ;
	wire _w7594_ ;
	wire _w7593_ ;
	wire _w7592_ ;
	wire _w7591_ ;
	wire _w7590_ ;
	wire _w7589_ ;
	wire _w7588_ ;
	wire _w7587_ ;
	wire _w7586_ ;
	wire _w7585_ ;
	wire _w7584_ ;
	wire _w7583_ ;
	wire _w7582_ ;
	wire _w7581_ ;
	wire _w7580_ ;
	wire _w7579_ ;
	wire _w7578_ ;
	wire _w7577_ ;
	wire _w7576_ ;
	wire _w7575_ ;
	wire _w7574_ ;
	wire _w7573_ ;
	wire _w7572_ ;
	wire _w7571_ ;
	wire _w7570_ ;
	wire _w7569_ ;
	wire _w7568_ ;
	wire _w7567_ ;
	wire _w7566_ ;
	wire _w7565_ ;
	wire _w7564_ ;
	wire _w7563_ ;
	wire _w7562_ ;
	wire _w7561_ ;
	wire _w7560_ ;
	wire _w7559_ ;
	wire _w7558_ ;
	wire _w7557_ ;
	wire _w7556_ ;
	wire _w7555_ ;
	wire _w7554_ ;
	wire _w7553_ ;
	wire _w7552_ ;
	wire _w7551_ ;
	wire _w7550_ ;
	wire _w7549_ ;
	wire _w7548_ ;
	wire _w7547_ ;
	wire _w7546_ ;
	wire _w7545_ ;
	wire _w7544_ ;
	wire _w7543_ ;
	wire _w7542_ ;
	wire _w7541_ ;
	wire _w7540_ ;
	wire _w7539_ ;
	wire _w7538_ ;
	wire _w7537_ ;
	wire _w7536_ ;
	wire _w7535_ ;
	wire _w7534_ ;
	wire _w7533_ ;
	wire _w7532_ ;
	wire _w7531_ ;
	wire _w7530_ ;
	wire _w7529_ ;
	wire _w7528_ ;
	wire _w7527_ ;
	wire _w7526_ ;
	wire _w7525_ ;
	wire _w7524_ ;
	wire _w7523_ ;
	wire _w7522_ ;
	wire _w7521_ ;
	wire _w7520_ ;
	wire _w7519_ ;
	wire _w7518_ ;
	wire _w7517_ ;
	wire _w7516_ ;
	wire _w7515_ ;
	wire _w7514_ ;
	wire _w7513_ ;
	wire _w7512_ ;
	wire _w7511_ ;
	wire _w7510_ ;
	wire _w7509_ ;
	wire _w7508_ ;
	wire _w7507_ ;
	wire _w7506_ ;
	wire _w7505_ ;
	wire _w7504_ ;
	wire _w7503_ ;
	wire _w7502_ ;
	wire _w7501_ ;
	wire _w7500_ ;
	wire _w7499_ ;
	wire _w7498_ ;
	wire _w7497_ ;
	wire _w7496_ ;
	wire _w7495_ ;
	wire _w7494_ ;
	wire _w7493_ ;
	wire _w7492_ ;
	wire _w7491_ ;
	wire _w7490_ ;
	wire _w7489_ ;
	wire _w7488_ ;
	wire _w7487_ ;
	wire _w7486_ ;
	wire _w7485_ ;
	wire _w7484_ ;
	wire _w7483_ ;
	wire _w7482_ ;
	wire _w7481_ ;
	wire _w7480_ ;
	wire _w7479_ ;
	wire _w7478_ ;
	wire _w7477_ ;
	wire _w7476_ ;
	wire _w7475_ ;
	wire _w7474_ ;
	wire _w7473_ ;
	wire _w7472_ ;
	wire _w7471_ ;
	wire _w7470_ ;
	wire _w7469_ ;
	wire _w7468_ ;
	wire _w7467_ ;
	wire _w7466_ ;
	wire _w7465_ ;
	wire _w7464_ ;
	wire _w7463_ ;
	wire _w7462_ ;
	wire _w7461_ ;
	wire _w7460_ ;
	wire _w7459_ ;
	wire _w7458_ ;
	wire _w7457_ ;
	wire _w7456_ ;
	wire _w7455_ ;
	wire _w7454_ ;
	wire _w7453_ ;
	wire _w7452_ ;
	wire _w7451_ ;
	wire _w7450_ ;
	wire _w7449_ ;
	wire _w7448_ ;
	wire _w7447_ ;
	wire _w7446_ ;
	wire _w7445_ ;
	wire _w7444_ ;
	wire _w7443_ ;
	wire _w7442_ ;
	wire _w7441_ ;
	wire _w7440_ ;
	wire _w7439_ ;
	wire _w7438_ ;
	wire _w7437_ ;
	wire _w7436_ ;
	wire _w7435_ ;
	wire _w7434_ ;
	wire _w7433_ ;
	wire _w7432_ ;
	wire _w7431_ ;
	wire _w7430_ ;
	wire _w7429_ ;
	wire _w7428_ ;
	wire _w7427_ ;
	wire _w7426_ ;
	wire _w7425_ ;
	wire _w7424_ ;
	wire _w7423_ ;
	wire _w7422_ ;
	wire _w7421_ ;
	wire _w7420_ ;
	wire _w7419_ ;
	wire _w7418_ ;
	wire _w7417_ ;
	wire _w7416_ ;
	wire _w7415_ ;
	wire _w7414_ ;
	wire _w7413_ ;
	wire _w7412_ ;
	wire _w7411_ ;
	wire _w7410_ ;
	wire _w7409_ ;
	wire _w7408_ ;
	wire _w7407_ ;
	wire _w7406_ ;
	wire _w7405_ ;
	wire _w7404_ ;
	wire _w7403_ ;
	wire _w7402_ ;
	wire _w7401_ ;
	wire _w7400_ ;
	wire _w7399_ ;
	wire _w7398_ ;
	wire _w7397_ ;
	wire _w7396_ ;
	wire _w7395_ ;
	wire _w7394_ ;
	wire _w7393_ ;
	wire _w7392_ ;
	wire _w7391_ ;
	wire _w7390_ ;
	wire _w7389_ ;
	wire _w7388_ ;
	wire _w7387_ ;
	wire _w7386_ ;
	wire _w7385_ ;
	wire _w7384_ ;
	wire _w7383_ ;
	wire _w7382_ ;
	wire _w7381_ ;
	wire _w7380_ ;
	wire _w7379_ ;
	wire _w7378_ ;
	wire _w7377_ ;
	wire _w7376_ ;
	wire _w7375_ ;
	wire _w7374_ ;
	wire _w7373_ ;
	wire _w7372_ ;
	wire _w7371_ ;
	wire _w7370_ ;
	wire _w7369_ ;
	wire _w7368_ ;
	wire _w7367_ ;
	wire _w7366_ ;
	wire _w7365_ ;
	wire _w7364_ ;
	wire _w7363_ ;
	wire _w7362_ ;
	wire _w7361_ ;
	wire _w7360_ ;
	wire _w7359_ ;
	wire _w7358_ ;
	wire _w7357_ ;
	wire _w7356_ ;
	wire _w7355_ ;
	wire _w7354_ ;
	wire _w7353_ ;
	wire _w7352_ ;
	wire _w7351_ ;
	wire _w7350_ ;
	wire _w7349_ ;
	wire _w7348_ ;
	wire _w7347_ ;
	wire _w7346_ ;
	wire _w7345_ ;
	wire _w7344_ ;
	wire _w7343_ ;
	wire _w7342_ ;
	wire _w7341_ ;
	wire _w7340_ ;
	wire _w7339_ ;
	wire _w7338_ ;
	wire _w7337_ ;
	wire _w7336_ ;
	wire _w7335_ ;
	wire _w7334_ ;
	wire _w7333_ ;
	wire _w7332_ ;
	wire _w7331_ ;
	wire _w7330_ ;
	wire _w7329_ ;
	wire _w7328_ ;
	wire _w7327_ ;
	wire _w7326_ ;
	wire _w7325_ ;
	wire _w7324_ ;
	wire _w7323_ ;
	wire _w7322_ ;
	wire _w7321_ ;
	wire _w7320_ ;
	wire _w7319_ ;
	wire _w7318_ ;
	wire _w7317_ ;
	wire _w7316_ ;
	wire _w7315_ ;
	wire _w7314_ ;
	wire _w7313_ ;
	wire _w7312_ ;
	wire _w7311_ ;
	wire _w7310_ ;
	wire _w7309_ ;
	wire _w7308_ ;
	wire _w7307_ ;
	wire _w7306_ ;
	wire _w7305_ ;
	wire _w7304_ ;
	wire _w7303_ ;
	wire _w7302_ ;
	wire _w7301_ ;
	wire _w7300_ ;
	wire _w7299_ ;
	wire _w7298_ ;
	wire _w7297_ ;
	wire _w7296_ ;
	wire _w7295_ ;
	wire _w7294_ ;
	wire _w7293_ ;
	wire _w7292_ ;
	wire _w7291_ ;
	wire _w7290_ ;
	wire _w7289_ ;
	wire _w7288_ ;
	wire _w7287_ ;
	wire _w7286_ ;
	wire _w7285_ ;
	wire _w7284_ ;
	wire _w7283_ ;
	wire _w7282_ ;
	wire _w7281_ ;
	wire _w7280_ ;
	wire _w7279_ ;
	wire _w7278_ ;
	wire _w7277_ ;
	wire _w7276_ ;
	wire _w7275_ ;
	wire _w7274_ ;
	wire _w7273_ ;
	wire _w7272_ ;
	wire _w7271_ ;
	wire _w7270_ ;
	wire _w7269_ ;
	wire _w7268_ ;
	wire _w7267_ ;
	wire _w7266_ ;
	wire _w7265_ ;
	wire _w7264_ ;
	wire _w7263_ ;
	wire _w7262_ ;
	wire _w7261_ ;
	wire _w7260_ ;
	wire _w7259_ ;
	wire _w7258_ ;
	wire _w7257_ ;
	wire _w7256_ ;
	wire _w7255_ ;
	wire _w7254_ ;
	wire _w7253_ ;
	wire _w7252_ ;
	wire _w7251_ ;
	wire _w7250_ ;
	wire _w7249_ ;
	wire _w7248_ ;
	wire _w7247_ ;
	wire _w7246_ ;
	wire _w7245_ ;
	wire _w7244_ ;
	wire _w7243_ ;
	wire _w7242_ ;
	wire _w7241_ ;
	wire _w7240_ ;
	wire _w7239_ ;
	wire _w7238_ ;
	wire _w7237_ ;
	wire _w7236_ ;
	wire _w7235_ ;
	wire _w7234_ ;
	wire _w7233_ ;
	wire _w7232_ ;
	wire _w7231_ ;
	wire _w7230_ ;
	wire _w7229_ ;
	wire _w7228_ ;
	wire _w7227_ ;
	wire _w7226_ ;
	wire _w7225_ ;
	wire _w7224_ ;
	wire _w7223_ ;
	wire _w7222_ ;
	wire _w7221_ ;
	wire _w7220_ ;
	wire _w7219_ ;
	wire _w7218_ ;
	wire _w7217_ ;
	wire _w7216_ ;
	wire _w7215_ ;
	wire _w7214_ ;
	wire _w7213_ ;
	wire _w7212_ ;
	wire _w7211_ ;
	wire _w7210_ ;
	wire _w7209_ ;
	wire _w7208_ ;
	wire _w7207_ ;
	wire _w7206_ ;
	wire _w7205_ ;
	wire _w7204_ ;
	wire _w7203_ ;
	wire _w7202_ ;
	wire _w7201_ ;
	wire _w7200_ ;
	wire _w7199_ ;
	wire _w7198_ ;
	wire _w7197_ ;
	wire _w7196_ ;
	wire _w7195_ ;
	wire _w7194_ ;
	wire _w7193_ ;
	wire _w7192_ ;
	wire _w7191_ ;
	wire _w7190_ ;
	wire _w7189_ ;
	wire _w7188_ ;
	wire _w7187_ ;
	wire _w7186_ ;
	wire _w7185_ ;
	wire _w7184_ ;
	wire _w7183_ ;
	wire _w7182_ ;
	wire _w7181_ ;
	wire _w7180_ ;
	wire _w7179_ ;
	wire _w7178_ ;
	wire _w7177_ ;
	wire _w7176_ ;
	wire _w7175_ ;
	wire _w7174_ ;
	wire _w7173_ ;
	wire _w7172_ ;
	wire _w7171_ ;
	wire _w7170_ ;
	wire _w7169_ ;
	wire _w7168_ ;
	wire _w7167_ ;
	wire _w7166_ ;
	wire _w7165_ ;
	wire _w7164_ ;
	wire _w7163_ ;
	wire _w7162_ ;
	wire _w7161_ ;
	wire _w7160_ ;
	wire _w7159_ ;
	wire _w7158_ ;
	wire _w7157_ ;
	wire _w7156_ ;
	wire _w7155_ ;
	wire _w7154_ ;
	wire _w7153_ ;
	wire _w7152_ ;
	wire _w7151_ ;
	wire _w7150_ ;
	wire _w7149_ ;
	wire _w7148_ ;
	wire _w7147_ ;
	wire _w7146_ ;
	wire _w7145_ ;
	wire _w7144_ ;
	wire _w7143_ ;
	wire _w7142_ ;
	wire _w7141_ ;
	wire _w7140_ ;
	wire _w7139_ ;
	wire _w7138_ ;
	wire _w7137_ ;
	wire _w7136_ ;
	wire _w7135_ ;
	wire _w7134_ ;
	wire _w7133_ ;
	wire _w7132_ ;
	wire _w7131_ ;
	wire _w7130_ ;
	wire _w7129_ ;
	wire _w7128_ ;
	wire _w7127_ ;
	wire _w7126_ ;
	wire _w7125_ ;
	wire _w7124_ ;
	wire _w7123_ ;
	wire _w7122_ ;
	wire _w7121_ ;
	wire _w7120_ ;
	wire _w7119_ ;
	wire _w7118_ ;
	wire _w7117_ ;
	wire _w7116_ ;
	wire _w7115_ ;
	wire _w7114_ ;
	wire _w7113_ ;
	wire _w7112_ ;
	wire _w7111_ ;
	wire _w7110_ ;
	wire _w7109_ ;
	wire _w7108_ ;
	wire _w7107_ ;
	wire _w7106_ ;
	wire _w7105_ ;
	wire _w7104_ ;
	wire _w7103_ ;
	wire _w7102_ ;
	wire _w7101_ ;
	wire _w7100_ ;
	wire _w7099_ ;
	wire _w7098_ ;
	wire _w7097_ ;
	wire _w7096_ ;
	wire _w7095_ ;
	wire _w7094_ ;
	wire _w7093_ ;
	wire _w7092_ ;
	wire _w7091_ ;
	wire _w7090_ ;
	wire _w7089_ ;
	wire _w7088_ ;
	wire _w7087_ ;
	wire _w7086_ ;
	wire _w7085_ ;
	wire _w7084_ ;
	wire _w7083_ ;
	wire _w7082_ ;
	wire _w7081_ ;
	wire _w7080_ ;
	wire _w7079_ ;
	wire _w7078_ ;
	wire _w7077_ ;
	wire _w7076_ ;
	wire _w7075_ ;
	wire _w7074_ ;
	wire _w7073_ ;
	wire _w7072_ ;
	wire _w7071_ ;
	wire _w7070_ ;
	wire _w7069_ ;
	wire _w7068_ ;
	wire _w7067_ ;
	wire _w7066_ ;
	wire _w7065_ ;
	wire _w7064_ ;
	wire _w7063_ ;
	wire _w7062_ ;
	wire _w7061_ ;
	wire _w7060_ ;
	wire _w7059_ ;
	wire _w7058_ ;
	wire _w7057_ ;
	wire _w7056_ ;
	wire _w7055_ ;
	wire _w7054_ ;
	wire _w7053_ ;
	wire _w7052_ ;
	wire _w7051_ ;
	wire _w7050_ ;
	wire _w7049_ ;
	wire _w7048_ ;
	wire _w7047_ ;
	wire _w7046_ ;
	wire _w7045_ ;
	wire _w7044_ ;
	wire _w7043_ ;
	wire _w7042_ ;
	wire _w7041_ ;
	wire _w7040_ ;
	wire _w7039_ ;
	wire _w7038_ ;
	wire _w7037_ ;
	wire _w7036_ ;
	wire _w7035_ ;
	wire _w7034_ ;
	wire _w7033_ ;
	wire _w7032_ ;
	wire _w7031_ ;
	wire _w7030_ ;
	wire _w7029_ ;
	wire _w7028_ ;
	wire _w7027_ ;
	wire _w7026_ ;
	wire _w7025_ ;
	wire _w7024_ ;
	wire _w7023_ ;
	wire _w7022_ ;
	wire _w7021_ ;
	wire _w7020_ ;
	wire _w7019_ ;
	wire _w7018_ ;
	wire _w7017_ ;
	wire _w7016_ ;
	wire _w7015_ ;
	wire _w7014_ ;
	wire _w7013_ ;
	wire _w7012_ ;
	wire _w7011_ ;
	wire _w7010_ ;
	wire _w7009_ ;
	wire _w7008_ ;
	wire _w7007_ ;
	wire _w7006_ ;
	wire _w7005_ ;
	wire _w7004_ ;
	wire _w7003_ ;
	wire _w7002_ ;
	wire _w7001_ ;
	wire _w7000_ ;
	wire _w6999_ ;
	wire _w6998_ ;
	wire _w6997_ ;
	wire _w6996_ ;
	wire _w6995_ ;
	wire _w6994_ ;
	wire _w6993_ ;
	wire _w6992_ ;
	wire _w6991_ ;
	wire _w6990_ ;
	wire _w6989_ ;
	wire _w6988_ ;
	wire _w4257_ ;
	wire _w4256_ ;
	wire _w4255_ ;
	wire _w4254_ ;
	wire _w4253_ ;
	wire _w4252_ ;
	wire _w4251_ ;
	wire _w4250_ ;
	wire _w4249_ ;
	wire _w4248_ ;
	wire _w4247_ ;
	wire _w4246_ ;
	wire _w4245_ ;
	wire _w4244_ ;
	wire _w4243_ ;
	wire _w4242_ ;
	wire _w4241_ ;
	wire _w4240_ ;
	wire _w4239_ ;
	wire _w4238_ ;
	wire _w4237_ ;
	wire _w4236_ ;
	wire _w4235_ ;
	wire _w4234_ ;
	wire _w4233_ ;
	wire _w4232_ ;
	wire _w4231_ ;
	wire _w4230_ ;
	wire _w4229_ ;
	wire _w4228_ ;
	wire _w4227_ ;
	wire _w4226_ ;
	wire _w4225_ ;
	wire _w4224_ ;
	wire _w4223_ ;
	wire _w4222_ ;
	wire _w4221_ ;
	wire _w4220_ ;
	wire _w4219_ ;
	wire _w4218_ ;
	wire _w4217_ ;
	wire _w4216_ ;
	wire _w4215_ ;
	wire _w4214_ ;
	wire _w4213_ ;
	wire _w4212_ ;
	wire _w4211_ ;
	wire _w4210_ ;
	wire _w4209_ ;
	wire _w4208_ ;
	wire _w4207_ ;
	wire _w4206_ ;
	wire _w4205_ ;
	wire _w4204_ ;
	wire _w4203_ ;
	wire _w4202_ ;
	wire _w4201_ ;
	wire _w4200_ ;
	wire _w4199_ ;
	wire _w4198_ ;
	wire _w4197_ ;
	wire _w4196_ ;
	wire _w4195_ ;
	wire _w4194_ ;
	wire _w4193_ ;
	wire _w4192_ ;
	wire _w4191_ ;
	wire _w4190_ ;
	wire _w4189_ ;
	wire _w4188_ ;
	wire _w4187_ ;
	wire _w4186_ ;
	wire _w4185_ ;
	wire _w4184_ ;
	wire _w4183_ ;
	wire _w4182_ ;
	wire _w4181_ ;
	wire _w4180_ ;
	wire _w4179_ ;
	wire _w4178_ ;
	wire _w4177_ ;
	wire _w4176_ ;
	wire _w4175_ ;
	wire _w4174_ ;
	wire _w4173_ ;
	wire _w4172_ ;
	wire _w4171_ ;
	wire _w4170_ ;
	wire _w4169_ ;
	wire _w4168_ ;
	wire _w4167_ ;
	wire _w4166_ ;
	wire _w4165_ ;
	wire _w4164_ ;
	wire _w4163_ ;
	wire _w4162_ ;
	wire _w4161_ ;
	wire _w4160_ ;
	wire _w4159_ ;
	wire _w4158_ ;
	wire _w4157_ ;
	wire _w4156_ ;
	wire _w4155_ ;
	wire _w4154_ ;
	wire _w4153_ ;
	wire _w4152_ ;
	wire _w4151_ ;
	wire _w4150_ ;
	wire _w4149_ ;
	wire _w4148_ ;
	wire _w4147_ ;
	wire _w4146_ ;
	wire _w4145_ ;
	wire _w4144_ ;
	wire _w4143_ ;
	wire _w4142_ ;
	wire _w4141_ ;
	wire _w4140_ ;
	wire _w4139_ ;
	wire _w4138_ ;
	wire _w4137_ ;
	wire _w4136_ ;
	wire _w4135_ ;
	wire _w4134_ ;
	wire _w4133_ ;
	wire _w4132_ ;
	wire _w4131_ ;
	wire _w4130_ ;
	wire _w4129_ ;
	wire _w4128_ ;
	wire _w4127_ ;
	wire _w4126_ ;
	wire _w4125_ ;
	wire _w4124_ ;
	wire _w4123_ ;
	wire _w4122_ ;
	wire _w4121_ ;
	wire _w4120_ ;
	wire _w4119_ ;
	wire _w4118_ ;
	wire _w4117_ ;
	wire _w4116_ ;
	wire _w4115_ ;
	wire _w4114_ ;
	wire _w4113_ ;
	wire _w4112_ ;
	wire _w4111_ ;
	wire _w4110_ ;
	wire _w4109_ ;
	wire _w4108_ ;
	wire _w4107_ ;
	wire _w4106_ ;
	wire _w4105_ ;
	wire _w4104_ ;
	wire _w4103_ ;
	wire _w4102_ ;
	wire _w4101_ ;
	wire _w4100_ ;
	wire _w4099_ ;
	wire _w4098_ ;
	wire _w4097_ ;
	wire _w4096_ ;
	wire _w4095_ ;
	wire _w4094_ ;
	wire _w4093_ ;
	wire _w4092_ ;
	wire _w4091_ ;
	wire _w4090_ ;
	wire _w4089_ ;
	wire _w4088_ ;
	wire _w4087_ ;
	wire _w4086_ ;
	wire _w4085_ ;
	wire _w4084_ ;
	wire _w4083_ ;
	wire _w4082_ ;
	wire _w4081_ ;
	wire _w4080_ ;
	wire _w4079_ ;
	wire _w4078_ ;
	wire _w4077_ ;
	wire _w4076_ ;
	wire _w4075_ ;
	wire _w4074_ ;
	wire _w4073_ ;
	wire _w4072_ ;
	wire _w4071_ ;
	wire _w4070_ ;
	wire _w4069_ ;
	wire _w4068_ ;
	wire _w4067_ ;
	wire _w4066_ ;
	wire _w4065_ ;
	wire _w4064_ ;
	wire _w4063_ ;
	wire _w4062_ ;
	wire _w4061_ ;
	wire _w4060_ ;
	wire _w4059_ ;
	wire _w4058_ ;
	wire _w4057_ ;
	wire _w4056_ ;
	wire _w4055_ ;
	wire _w4054_ ;
	wire _w4053_ ;
	wire _w4052_ ;
	wire _w4051_ ;
	wire _w4050_ ;
	wire _w4049_ ;
	wire _w4048_ ;
	wire _w4047_ ;
	wire _w4046_ ;
	wire _w4045_ ;
	wire _w4044_ ;
	wire _w4043_ ;
	wire _w4042_ ;
	wire _w4041_ ;
	wire _w4040_ ;
	wire _w4039_ ;
	wire _w4038_ ;
	wire _w4037_ ;
	wire _w4036_ ;
	wire _w4035_ ;
	wire _w4034_ ;
	wire _w4033_ ;
	wire _w4032_ ;
	wire _w4031_ ;
	wire _w4030_ ;
	wire _w4029_ ;
	wire _w4028_ ;
	wire _w4027_ ;
	wire _w4026_ ;
	wire _w4025_ ;
	wire _w4024_ ;
	wire _w4023_ ;
	wire _w4022_ ;
	wire _w4021_ ;
	wire _w4020_ ;
	wire _w4019_ ;
	wire _w4018_ ;
	wire _w4017_ ;
	wire _w4016_ ;
	wire _w4015_ ;
	wire _w4014_ ;
	wire _w4013_ ;
	wire _w4012_ ;
	wire _w4011_ ;
	wire _w4010_ ;
	wire _w4009_ ;
	wire _w4008_ ;
	wire _w4007_ ;
	wire _w4006_ ;
	wire _w4005_ ;
	wire _w4004_ ;
	wire _w4003_ ;
	wire _w4002_ ;
	wire _w4001_ ;
	wire _w4000_ ;
	wire _w3999_ ;
	wire _w3998_ ;
	wire _w3997_ ;
	wire _w3996_ ;
	wire _w3995_ ;
	wire _w3994_ ;
	wire _w3993_ ;
	wire _w3992_ ;
	wire _w3991_ ;
	wire _w3990_ ;
	wire _w3989_ ;
	wire _w3988_ ;
	wire _w3987_ ;
	wire _w3986_ ;
	wire _w3985_ ;
	wire _w3984_ ;
	wire _w3983_ ;
	wire _w3982_ ;
	wire _w3981_ ;
	wire _w3980_ ;
	wire _w3979_ ;
	wire _w3978_ ;
	wire _w3977_ ;
	wire _w3976_ ;
	wire _w3975_ ;
	wire _w3974_ ;
	wire _w3973_ ;
	wire _w3972_ ;
	wire _w3971_ ;
	wire _w3970_ ;
	wire _w3969_ ;
	wire _w3968_ ;
	wire _w3967_ ;
	wire _w3966_ ;
	wire _w3965_ ;
	wire _w3964_ ;
	wire _w3963_ ;
	wire _w3962_ ;
	wire _w3961_ ;
	wire _w3960_ ;
	wire _w3959_ ;
	wire _w3958_ ;
	wire _w3957_ ;
	wire _w3956_ ;
	wire _w3955_ ;
	wire _w3954_ ;
	wire _w3953_ ;
	wire _w3952_ ;
	wire _w3951_ ;
	wire _w3950_ ;
	wire _w3949_ ;
	wire _w3948_ ;
	wire _w3947_ ;
	wire _w3946_ ;
	wire _w3945_ ;
	wire _w3944_ ;
	wire _w3943_ ;
	wire _w3942_ ;
	wire _w3941_ ;
	wire _w3940_ ;
	wire _w3939_ ;
	wire _w3938_ ;
	wire _w3937_ ;
	wire _w3936_ ;
	wire _w3935_ ;
	wire _w3934_ ;
	wire _w3933_ ;
	wire _w3932_ ;
	wire _w3931_ ;
	wire _w3930_ ;
	wire _w3929_ ;
	wire _w3928_ ;
	wire _w3927_ ;
	wire _w3926_ ;
	wire _w3925_ ;
	wire _w3924_ ;
	wire _w3923_ ;
	wire _w3922_ ;
	wire _w3921_ ;
	wire _w3920_ ;
	wire _w3919_ ;
	wire _w3918_ ;
	wire _w3917_ ;
	wire _w3916_ ;
	wire _w3915_ ;
	wire _w3914_ ;
	wire _w3913_ ;
	wire _w3912_ ;
	wire _w3911_ ;
	wire _w3910_ ;
	wire _w3909_ ;
	wire _w3908_ ;
	wire _w3907_ ;
	wire _w3906_ ;
	wire _w3905_ ;
	wire _w3904_ ;
	wire _w3903_ ;
	wire _w3902_ ;
	wire _w3901_ ;
	wire _w3900_ ;
	wire _w3899_ ;
	wire _w3898_ ;
	wire _w3897_ ;
	wire _w3896_ ;
	wire _w3895_ ;
	wire _w3894_ ;
	wire _w3893_ ;
	wire _w3892_ ;
	wire _w3891_ ;
	wire _w3890_ ;
	wire _w3889_ ;
	wire _w3888_ ;
	wire _w3887_ ;
	wire _w3886_ ;
	wire _w3885_ ;
	wire _w3884_ ;
	wire _w3883_ ;
	wire _w3882_ ;
	wire _w3881_ ;
	wire _w3880_ ;
	wire _w3879_ ;
	wire _w3878_ ;
	wire _w3877_ ;
	wire _w3876_ ;
	wire _w3875_ ;
	wire _w3874_ ;
	wire _w3873_ ;
	wire _w3872_ ;
	wire _w3871_ ;
	wire _w3870_ ;
	wire _w3869_ ;
	wire _w3868_ ;
	wire _w3867_ ;
	wire _w3866_ ;
	wire _w3865_ ;
	wire _w3864_ ;
	wire _w3863_ ;
	wire _w3862_ ;
	wire _w3861_ ;
	wire _w3860_ ;
	wire _w3859_ ;
	wire _w3858_ ;
	wire _w3857_ ;
	wire _w3856_ ;
	wire _w3855_ ;
	wire _w3854_ ;
	wire _w3853_ ;
	wire _w3852_ ;
	wire _w3851_ ;
	wire _w3850_ ;
	wire _w3849_ ;
	wire _w3848_ ;
	wire _w3847_ ;
	wire _w3846_ ;
	wire _w3845_ ;
	wire _w3844_ ;
	wire _w3843_ ;
	wire _w3842_ ;
	wire _w3841_ ;
	wire _w3840_ ;
	wire _w3839_ ;
	wire _w3838_ ;
	wire _w3837_ ;
	wire _w3836_ ;
	wire _w3835_ ;
	wire _w3834_ ;
	wire _w3833_ ;
	wire _w3832_ ;
	wire _w3831_ ;
	wire _w3830_ ;
	wire _w3829_ ;
	wire _w3828_ ;
	wire _w3827_ ;
	wire _w3826_ ;
	wire _w3825_ ;
	wire _w3824_ ;
	wire _w3823_ ;
	wire _w3822_ ;
	wire _w3821_ ;
	wire _w3820_ ;
	wire _w3819_ ;
	wire _w3818_ ;
	wire _w3817_ ;
	wire _w3816_ ;
	wire _w3815_ ;
	wire _w3814_ ;
	wire _w3813_ ;
	wire _w3812_ ;
	wire _w3811_ ;
	wire _w3810_ ;
	wire _w3809_ ;
	wire _w3808_ ;
	wire _w3807_ ;
	wire _w3806_ ;
	wire _w3805_ ;
	wire _w3804_ ;
	wire _w3803_ ;
	wire _w3802_ ;
	wire _w3801_ ;
	wire _w3800_ ;
	wire _w3799_ ;
	wire _w3798_ ;
	wire _w3797_ ;
	wire _w3796_ ;
	wire _w3795_ ;
	wire _w3794_ ;
	wire _w3793_ ;
	wire _w3792_ ;
	wire _w3791_ ;
	wire _w3790_ ;
	wire _w3789_ ;
	wire _w3788_ ;
	wire _w3787_ ;
	wire _w3786_ ;
	wire _w3785_ ;
	wire _w3784_ ;
	wire _w3783_ ;
	wire _w3782_ ;
	wire _w3781_ ;
	wire _w3780_ ;
	wire _w3779_ ;
	wire _w3778_ ;
	wire _w3777_ ;
	wire _w3776_ ;
	wire _w3775_ ;
	wire _w3774_ ;
	wire _w3773_ ;
	wire _w3772_ ;
	wire _w3771_ ;
	wire _w3770_ ;
	wire _w3769_ ;
	wire _w3768_ ;
	wire _w3767_ ;
	wire _w3766_ ;
	wire _w3765_ ;
	wire _w3764_ ;
	wire _w3763_ ;
	wire _w3762_ ;
	wire _w3761_ ;
	wire _w3760_ ;
	wire _w3759_ ;
	wire _w3758_ ;
	wire _w3757_ ;
	wire _w3756_ ;
	wire _w3755_ ;
	wire _w3754_ ;
	wire _w3753_ ;
	wire _w3752_ ;
	wire _w3751_ ;
	wire _w3750_ ;
	wire _w3749_ ;
	wire _w3748_ ;
	wire _w3747_ ;
	wire _w3746_ ;
	wire _w3745_ ;
	wire _w3744_ ;
	wire _w3743_ ;
	wire _w3742_ ;
	wire _w3741_ ;
	wire _w3740_ ;
	wire _w3739_ ;
	wire _w3738_ ;
	wire _w3737_ ;
	wire _w3736_ ;
	wire _w3735_ ;
	wire _w3734_ ;
	wire _w3733_ ;
	wire _w3732_ ;
	wire _w3731_ ;
	wire _w3730_ ;
	wire _w3729_ ;
	wire _w3728_ ;
	wire _w3727_ ;
	wire _w3726_ ;
	wire _w3725_ ;
	wire _w3724_ ;
	wire _w3723_ ;
	wire _w3722_ ;
	wire _w3721_ ;
	wire _w3720_ ;
	wire _w3719_ ;
	wire _w3718_ ;
	wire _w3717_ ;
	wire _w3716_ ;
	wire _w3715_ ;
	wire _w3714_ ;
	wire _w3713_ ;
	wire _w3712_ ;
	wire _w3711_ ;
	wire _w3710_ ;
	wire _w3709_ ;
	wire _w3708_ ;
	wire _w3707_ ;
	wire _w3706_ ;
	wire _w3705_ ;
	wire _w3704_ ;
	wire _w3703_ ;
	wire _w3702_ ;
	wire _w3701_ ;
	wire _w3700_ ;
	wire _w3699_ ;
	wire _w3698_ ;
	wire _w3697_ ;
	wire _w3696_ ;
	wire _w3695_ ;
	wire _w3694_ ;
	wire _w3693_ ;
	wire _w3692_ ;
	wire _w3691_ ;
	wire _w3690_ ;
	wire _w3689_ ;
	wire _w3688_ ;
	wire _w3687_ ;
	wire _w3686_ ;
	wire _w3685_ ;
	wire _w3684_ ;
	wire _w3683_ ;
	wire _w3682_ ;
	wire _w3681_ ;
	wire _w3680_ ;
	wire _w3679_ ;
	wire _w3678_ ;
	wire _w3677_ ;
	wire _w3676_ ;
	wire _w3675_ ;
	wire _w3674_ ;
	wire _w3673_ ;
	wire _w3672_ ;
	wire _w3671_ ;
	wire _w3670_ ;
	wire _w3669_ ;
	wire _w3668_ ;
	wire _w3667_ ;
	wire _w3666_ ;
	wire _w3665_ ;
	wire _w3664_ ;
	wire _w3663_ ;
	wire _w3662_ ;
	wire _w3661_ ;
	wire _w3660_ ;
	wire _w3659_ ;
	wire _w3658_ ;
	wire _w3657_ ;
	wire _w3656_ ;
	wire _w3655_ ;
	wire _w3654_ ;
	wire _w3653_ ;
	wire _w3652_ ;
	wire _w3651_ ;
	wire _w3650_ ;
	wire _w3649_ ;
	wire _w3648_ ;
	wire _w3647_ ;
	wire _w3646_ ;
	wire _w3645_ ;
	wire _w3644_ ;
	wire _w3643_ ;
	wire _w3642_ ;
	wire _w3641_ ;
	wire _w3640_ ;
	wire _w3639_ ;
	wire _w3638_ ;
	wire _w3637_ ;
	wire _w3636_ ;
	wire _w3635_ ;
	wire _w3634_ ;
	wire _w3633_ ;
	wire _w3632_ ;
	wire _w3631_ ;
	wire _w3630_ ;
	wire _w3629_ ;
	wire _w3628_ ;
	wire _w3627_ ;
	wire _w3626_ ;
	wire _w3625_ ;
	wire _w3624_ ;
	wire _w3623_ ;
	wire _w3622_ ;
	wire _w3621_ ;
	wire _w3620_ ;
	wire _w3619_ ;
	wire _w3618_ ;
	wire _w3617_ ;
	wire _w3616_ ;
	wire _w3615_ ;
	wire _w3614_ ;
	wire _w3613_ ;
	wire _w3612_ ;
	wire _w3611_ ;
	wire _w3610_ ;
	wire _w3609_ ;
	wire _w3608_ ;
	wire _w3607_ ;
	wire _w3606_ ;
	wire _w3605_ ;
	wire _w3604_ ;
	wire _w3603_ ;
	wire _w3602_ ;
	wire _w3601_ ;
	wire _w3600_ ;
	wire _w3599_ ;
	wire _w3598_ ;
	wire _w3597_ ;
	wire _w3596_ ;
	wire _w3595_ ;
	wire _w3594_ ;
	wire _w3593_ ;
	wire _w3592_ ;
	wire _w3591_ ;
	wire _w3590_ ;
	wire _w3589_ ;
	wire _w3588_ ;
	wire _w3587_ ;
	wire _w3586_ ;
	wire _w3585_ ;
	wire _w3584_ ;
	wire _w3583_ ;
	wire _w3582_ ;
	wire _w3581_ ;
	wire _w3580_ ;
	wire _w3579_ ;
	wire _w3578_ ;
	wire _w3577_ ;
	wire _w3576_ ;
	wire _w3575_ ;
	wire _w3574_ ;
	wire _w3573_ ;
	wire _w3572_ ;
	wire _w3571_ ;
	wire _w3570_ ;
	wire _w3569_ ;
	wire _w3568_ ;
	wire _w3567_ ;
	wire _w3566_ ;
	wire _w3565_ ;
	wire _w3564_ ;
	wire _w3563_ ;
	wire _w3562_ ;
	wire _w3561_ ;
	wire _w3560_ ;
	wire _w3559_ ;
	wire _w3558_ ;
	wire _w3557_ ;
	wire _w3556_ ;
	wire _w3555_ ;
	wire _w3554_ ;
	wire _w3553_ ;
	wire _w3552_ ;
	wire _w3551_ ;
	wire _w3550_ ;
	wire _w3549_ ;
	wire _w3548_ ;
	wire _w3547_ ;
	wire _w3546_ ;
	wire _w3545_ ;
	wire _w3544_ ;
	wire _w3543_ ;
	wire _w3542_ ;
	wire _w3541_ ;
	wire _w3540_ ;
	wire _w3539_ ;
	wire _w3538_ ;
	wire _w3537_ ;
	wire _w3536_ ;
	wire _w3535_ ;
	wire _w3534_ ;
	wire _w3533_ ;
	wire _w3532_ ;
	wire _w3531_ ;
	wire _w3530_ ;
	wire _w3529_ ;
	wire _w3528_ ;
	wire _w3527_ ;
	wire _w3526_ ;
	wire _w3525_ ;
	wire _w3524_ ;
	wire _w3523_ ;
	wire _w3522_ ;
	wire _w3521_ ;
	wire _w3520_ ;
	wire _w3519_ ;
	wire _w3518_ ;
	wire _w3517_ ;
	wire _w3516_ ;
	wire _w3515_ ;
	wire _w3514_ ;
	wire _w3513_ ;
	wire _w3512_ ;
	wire _w3511_ ;
	wire _w3510_ ;
	wire _w3509_ ;
	wire _w3508_ ;
	wire _w3507_ ;
	wire _w3506_ ;
	wire _w3505_ ;
	wire _w3504_ ;
	wire _w3503_ ;
	wire _w3502_ ;
	wire _w3501_ ;
	wire _w3500_ ;
	wire _w3499_ ;
	wire _w3498_ ;
	wire _w3497_ ;
	wire _w3496_ ;
	wire _w3495_ ;
	wire _w3494_ ;
	wire _w3493_ ;
	wire _w3492_ ;
	wire _w3491_ ;
	wire _w3490_ ;
	wire _w3489_ ;
	wire _w3488_ ;
	wire _w3487_ ;
	wire _w3486_ ;
	wire _w3485_ ;
	wire _w3484_ ;
	wire _w3483_ ;
	wire _w3482_ ;
	wire _w3481_ ;
	wire _w3480_ ;
	wire _w3479_ ;
	wire _w3478_ ;
	wire _w3477_ ;
	wire _w3476_ ;
	wire _w3475_ ;
	wire _w3474_ ;
	wire _w3473_ ;
	wire _w3472_ ;
	wire _w3471_ ;
	wire _w3470_ ;
	wire _w3469_ ;
	wire _w3468_ ;
	wire _w3467_ ;
	wire _w3466_ ;
	wire _w3465_ ;
	wire _w3464_ ;
	wire _w3463_ ;
	wire _w3462_ ;
	wire _w3461_ ;
	wire _w3460_ ;
	wire _w3459_ ;
	wire _w3458_ ;
	wire _w3457_ ;
	wire _w3456_ ;
	wire _w3455_ ;
	wire _w3454_ ;
	wire _w3453_ ;
	wire _w3452_ ;
	wire _w3451_ ;
	wire _w3450_ ;
	wire _w3449_ ;
	wire _w3448_ ;
	wire _w3447_ ;
	wire _w3446_ ;
	wire _w3445_ ;
	wire _w3444_ ;
	wire _w3443_ ;
	wire _w3442_ ;
	wire _w3441_ ;
	wire _w3440_ ;
	wire _w3439_ ;
	wire _w3438_ ;
	wire _w3437_ ;
	wire _w3436_ ;
	wire _w3435_ ;
	wire _w3434_ ;
	wire _w3433_ ;
	wire _w3432_ ;
	wire _w3431_ ;
	wire _w3430_ ;
	wire _w3429_ ;
	wire _w3428_ ;
	wire _w3427_ ;
	wire _w3426_ ;
	wire _w3425_ ;
	wire _w3424_ ;
	wire _w3423_ ;
	wire _w3422_ ;
	wire _w3421_ ;
	wire _w3420_ ;
	wire _w3419_ ;
	wire _w3418_ ;
	wire _w3417_ ;
	wire _w3416_ ;
	wire _w3415_ ;
	wire _w3414_ ;
	wire _w3413_ ;
	wire _w3412_ ;
	wire _w3411_ ;
	wire _w3410_ ;
	wire _w3409_ ;
	wire _w3408_ ;
	wire _w3407_ ;
	wire _w3406_ ;
	wire _w3405_ ;
	wire _w3404_ ;
	wire _w3403_ ;
	wire _w3402_ ;
	wire _w3401_ ;
	wire _w3400_ ;
	wire _w3399_ ;
	wire _w3398_ ;
	wire _w3397_ ;
	wire _w3396_ ;
	wire _w3395_ ;
	wire _w3394_ ;
	wire _w3393_ ;
	wire _w3392_ ;
	wire _w3391_ ;
	wire _w3390_ ;
	wire _w3389_ ;
	wire _w3388_ ;
	wire _w3387_ ;
	wire _w3386_ ;
	wire _w3385_ ;
	wire _w3384_ ;
	wire _w3383_ ;
	wire _w3382_ ;
	wire _w3381_ ;
	wire _w3380_ ;
	wire _w3379_ ;
	wire _w3378_ ;
	wire _w3377_ ;
	wire _w3376_ ;
	wire _w3375_ ;
	wire _w3374_ ;
	wire _w3373_ ;
	wire _w3372_ ;
	wire _w3371_ ;
	wire _w3370_ ;
	wire _w3369_ ;
	wire _w3368_ ;
	wire _w3367_ ;
	wire _w3366_ ;
	wire _w3365_ ;
	wire _w3364_ ;
	wire _w3363_ ;
	wire _w3362_ ;
	wire _w3361_ ;
	wire _w3360_ ;
	wire _w3359_ ;
	wire _w3358_ ;
	wire _w3357_ ;
	wire _w3356_ ;
	wire _w3355_ ;
	wire _w3354_ ;
	wire _w3353_ ;
	wire _w3352_ ;
	wire _w3351_ ;
	wire _w3350_ ;
	wire _w3349_ ;
	wire _w3348_ ;
	wire _w3347_ ;
	wire _w3346_ ;
	wire _w3345_ ;
	wire _w3344_ ;
	wire _w3343_ ;
	wire _w3342_ ;
	wire _w3341_ ;
	wire _w3340_ ;
	wire _w3339_ ;
	wire _w3338_ ;
	wire _w3337_ ;
	wire _w3336_ ;
	wire _w3335_ ;
	wire _w3334_ ;
	wire _w3333_ ;
	wire _w3332_ ;
	wire _w3331_ ;
	wire _w3330_ ;
	wire _w3329_ ;
	wire _w3328_ ;
	wire _w3327_ ;
	wire _w3326_ ;
	wire _w3325_ ;
	wire _w3324_ ;
	wire _w3323_ ;
	wire _w3322_ ;
	wire _w3321_ ;
	wire _w3320_ ;
	wire _w3319_ ;
	wire _w3318_ ;
	wire _w3317_ ;
	wire _w3316_ ;
	wire _w3315_ ;
	wire _w3314_ ;
	wire _w3313_ ;
	wire _w3312_ ;
	wire _w3311_ ;
	wire _w3310_ ;
	wire _w3309_ ;
	wire _w3308_ ;
	wire _w3307_ ;
	wire _w3306_ ;
	wire _w3305_ ;
	wire _w3304_ ;
	wire _w3303_ ;
	wire _w3302_ ;
	wire _w3301_ ;
	wire _w3300_ ;
	wire _w3299_ ;
	wire _w3298_ ;
	wire _w3297_ ;
	wire _w3296_ ;
	wire _w3295_ ;
	wire _w3294_ ;
	wire _w3293_ ;
	wire _w3292_ ;
	wire _w3291_ ;
	wire _w3290_ ;
	wire _w3289_ ;
	wire _w3288_ ;
	wire _w3287_ ;
	wire _w3286_ ;
	wire _w3285_ ;
	wire _w3284_ ;
	wire _w3283_ ;
	wire _w3282_ ;
	wire _w3281_ ;
	wire _w3280_ ;
	wire _w3279_ ;
	wire _w3278_ ;
	wire _w3277_ ;
	wire _w3276_ ;
	wire _w3275_ ;
	wire _w3274_ ;
	wire _w3273_ ;
	wire _w3272_ ;
	wire _w3271_ ;
	wire _w3270_ ;
	wire _w3269_ ;
	wire _w3268_ ;
	wire _w3267_ ;
	wire _w3266_ ;
	wire _w3265_ ;
	wire _w3264_ ;
	wire _w3263_ ;
	wire _w3262_ ;
	wire _w3261_ ;
	wire _w3260_ ;
	wire _w3259_ ;
	wire _w3258_ ;
	wire _w3257_ ;
	wire _w3256_ ;
	wire _w3255_ ;
	wire _w3254_ ;
	wire _w3253_ ;
	wire _w3252_ ;
	wire _w3251_ ;
	wire _w3250_ ;
	wire _w3249_ ;
	wire _w3248_ ;
	wire _w3247_ ;
	wire _w3246_ ;
	wire _w3245_ ;
	wire _w3244_ ;
	wire _w3243_ ;
	wire _w3242_ ;
	wire _w3241_ ;
	wire _w3240_ ;
	wire _w3239_ ;
	wire _w3238_ ;
	wire _w3237_ ;
	wire _w3236_ ;
	wire _w3235_ ;
	wire _w3234_ ;
	wire _w3233_ ;
	wire _w3232_ ;
	wire _w3231_ ;
	wire _w3230_ ;
	wire _w3229_ ;
	wire _w3228_ ;
	wire _w3227_ ;
	wire _w3226_ ;
	wire _w3225_ ;
	wire _w3224_ ;
	wire _w3223_ ;
	wire _w3222_ ;
	wire _w3221_ ;
	wire _w3220_ ;
	wire _w3219_ ;
	wire _w3218_ ;
	wire _w3217_ ;
	wire _w3216_ ;
	wire _w3215_ ;
	wire _w3214_ ;
	wire _w3213_ ;
	wire _w3212_ ;
	wire _w3211_ ;
	wire _w3210_ ;
	wire _w3209_ ;
	wire _w3208_ ;
	wire _w3207_ ;
	wire _w3206_ ;
	wire _w3205_ ;
	wire _w3204_ ;
	wire _w3203_ ;
	wire _w3202_ ;
	wire _w3201_ ;
	wire _w3200_ ;
	wire _w3199_ ;
	wire _w3198_ ;
	wire _w3197_ ;
	wire _w3196_ ;
	wire _w3195_ ;
	wire _w3194_ ;
	wire _w3193_ ;
	wire _w3192_ ;
	wire _w3191_ ;
	wire _w3190_ ;
	wire _w3189_ ;
	wire _w3188_ ;
	wire _w3187_ ;
	wire _w3186_ ;
	wire _w3185_ ;
	wire _w3184_ ;
	wire _w3183_ ;
	wire _w3182_ ;
	wire _w3181_ ;
	wire _w3180_ ;
	wire _w3179_ ;
	wire _w3178_ ;
	wire _w3177_ ;
	wire _w3176_ ;
	wire _w3175_ ;
	wire _w3174_ ;
	wire _w3173_ ;
	wire _w3172_ ;
	wire _w3171_ ;
	wire _w3170_ ;
	wire _w3169_ ;
	wire _w3168_ ;
	wire _w3167_ ;
	wire _w3166_ ;
	wire _w3165_ ;
	wire _w3164_ ;
	wire _w3163_ ;
	wire _w3162_ ;
	wire _w3161_ ;
	wire _w3160_ ;
	wire _w3159_ ;
	wire _w3158_ ;
	wire _w3157_ ;
	wire _w3156_ ;
	wire _w3155_ ;
	wire _w3154_ ;
	wire _w3153_ ;
	wire _w3152_ ;
	wire _w3151_ ;
	wire _w3150_ ;
	wire _w3149_ ;
	wire _w3148_ ;
	wire _w3147_ ;
	wire _w3146_ ;
	wire _w3145_ ;
	wire _w3144_ ;
	wire _w3143_ ;
	wire _w3142_ ;
	wire _w3141_ ;
	wire _w3140_ ;
	wire _w3139_ ;
	wire _w3138_ ;
	wire _w3137_ ;
	wire _w3136_ ;
	wire _w3135_ ;
	wire _w3134_ ;
	wire _w3133_ ;
	wire _w3132_ ;
	wire _w3131_ ;
	wire _w3130_ ;
	wire _w3129_ ;
	wire _w3128_ ;
	wire _w3127_ ;
	wire _w3126_ ;
	wire _w3125_ ;
	wire _w3124_ ;
	wire _w3123_ ;
	wire _w3122_ ;
	wire _w3121_ ;
	wire _w3120_ ;
	wire _w3119_ ;
	wire _w3118_ ;
	wire _w3117_ ;
	wire _w3116_ ;
	wire _w3115_ ;
	wire _w3114_ ;
	wire _w3113_ ;
	wire _w3112_ ;
	wire _w3111_ ;
	wire _w3110_ ;
	wire _w3109_ ;
	wire _w3108_ ;
	wire _w3107_ ;
	wire _w3106_ ;
	wire _w3105_ ;
	wire _w3104_ ;
	wire _w3103_ ;
	wire _w3102_ ;
	wire _w3101_ ;
	wire _w3100_ ;
	wire _w3099_ ;
	wire _w3098_ ;
	wire _w3097_ ;
	wire _w3096_ ;
	wire _w3095_ ;
	wire _w3094_ ;
	wire _w3093_ ;
	wire _w3092_ ;
	wire _w3091_ ;
	wire _w3090_ ;
	wire _w3089_ ;
	wire _w3088_ ;
	wire _w3087_ ;
	wire _w3086_ ;
	wire _w3085_ ;
	wire _w3084_ ;
	wire _w3083_ ;
	wire _w3082_ ;
	wire _w3081_ ;
	wire _w3080_ ;
	wire _w3079_ ;
	wire _w3078_ ;
	wire _w3077_ ;
	wire _w3076_ ;
	wire _w3075_ ;
	wire _w3074_ ;
	wire _w3073_ ;
	wire _w3072_ ;
	wire _w3071_ ;
	wire _w3070_ ;
	wire _w3069_ ;
	wire _w3068_ ;
	wire _w3067_ ;
	wire _w3066_ ;
	wire _w3065_ ;
	wire _w3064_ ;
	wire _w3063_ ;
	wire _w3062_ ;
	wire _w3061_ ;
	wire _w3060_ ;
	wire _w3059_ ;
	wire _w3058_ ;
	wire _w3057_ ;
	wire _w3056_ ;
	wire _w3055_ ;
	wire _w3054_ ;
	wire _w3053_ ;
	wire _w3052_ ;
	wire _w3051_ ;
	wire _w3050_ ;
	wire _w3049_ ;
	wire _w3048_ ;
	wire _w3047_ ;
	wire _w3046_ ;
	wire _w3045_ ;
	wire _w3044_ ;
	wire _w3043_ ;
	wire _w3042_ ;
	wire _w3041_ ;
	wire _w3040_ ;
	wire _w3039_ ;
	wire _w3038_ ;
	wire _w3037_ ;
	wire _w3036_ ;
	wire _w3035_ ;
	wire _w3034_ ;
	wire _w3033_ ;
	wire _w3032_ ;
	wire _w3031_ ;
	wire _w3030_ ;
	wire _w3029_ ;
	wire _w3028_ ;
	wire _w3027_ ;
	wire _w3026_ ;
	wire _w3025_ ;
	wire _w3024_ ;
	wire _w3023_ ;
	wire _w3022_ ;
	wire _w3021_ ;
	wire _w3020_ ;
	wire _w3019_ ;
	wire _w3018_ ;
	wire _w3017_ ;
	wire _w3016_ ;
	wire _w3015_ ;
	wire _w3014_ ;
	wire _w3013_ ;
	wire _w3012_ ;
	wire _w3011_ ;
	wire _w3010_ ;
	wire _w2441_ ;
	wire _w2440_ ;
	wire _w2439_ ;
	wire _w2438_ ;
	wire _w2437_ ;
	wire _w2436_ ;
	wire _w2435_ ;
	wire _w2434_ ;
	wire _w2433_ ;
	wire _w2432_ ;
	wire _w2431_ ;
	wire _w2430_ ;
	wire _w2429_ ;
	wire _w2428_ ;
	wire _w2427_ ;
	wire _w2426_ ;
	wire _w2425_ ;
	wire _w2424_ ;
	wire _w2423_ ;
	wire _w2422_ ;
	wire _w2421_ ;
	wire _w2420_ ;
	wire _w2419_ ;
	wire _w2418_ ;
	wire _w2417_ ;
	wire _w2416_ ;
	wire _w2415_ ;
	wire _w2414_ ;
	wire _w2413_ ;
	wire _w2412_ ;
	wire _w2411_ ;
	wire _w2410_ ;
	wire _w2409_ ;
	wire _w2408_ ;
	wire _w2407_ ;
	wire _w2406_ ;
	wire _w2405_ ;
	wire _w2404_ ;
	wire _w2403_ ;
	wire _w2402_ ;
	wire _w2401_ ;
	wire _w2400_ ;
	wire _w2399_ ;
	wire _w2398_ ;
	wire _w2397_ ;
	wire _w2396_ ;
	wire _w2395_ ;
	wire _w2394_ ;
	wire _w2393_ ;
	wire _w2392_ ;
	wire _w2391_ ;
	wire _w2390_ ;
	wire _w2389_ ;
	wire _w2388_ ;
	wire _w2387_ ;
	wire _w2386_ ;
	wire _w2385_ ;
	wire _w2384_ ;
	wire _w2383_ ;
	wire _w2382_ ;
	wire _w2381_ ;
	wire _w2380_ ;
	wire _w2379_ ;
	wire _w2378_ ;
	wire _w2377_ ;
	wire _w2376_ ;
	wire _w2375_ ;
	wire _w2374_ ;
	wire _w2373_ ;
	wire _w2372_ ;
	wire _w2371_ ;
	wire _w2370_ ;
	wire _w2369_ ;
	wire _w2368_ ;
	wire _w2367_ ;
	wire _w2366_ ;
	wire _w2365_ ;
	wire _w2364_ ;
	wire _w2363_ ;
	wire _w2362_ ;
	wire _w2361_ ;
	wire _w2360_ ;
	wire _w2359_ ;
	wire _w2358_ ;
	wire _w2357_ ;
	wire _w2356_ ;
	wire _w2355_ ;
	wire _w2354_ ;
	wire _w2353_ ;
	wire _w2352_ ;
	wire _w2351_ ;
	wire _w2350_ ;
	wire _w2349_ ;
	wire _w2348_ ;
	wire _w2347_ ;
	wire _w2346_ ;
	wire _w2345_ ;
	wire _w2344_ ;
	wire _w2343_ ;
	wire _w2342_ ;
	wire _w2341_ ;
	wire _w2340_ ;
	wire _w2339_ ;
	wire _w2338_ ;
	wire _w2337_ ;
	wire _w2336_ ;
	wire _w2335_ ;
	wire _w2334_ ;
	wire _w2333_ ;
	wire _w2332_ ;
	wire _w2331_ ;
	wire _w2330_ ;
	wire _w2329_ ;
	wire _w2328_ ;
	wire _w2327_ ;
	wire _w2326_ ;
	wire _w2325_ ;
	wire _w2324_ ;
	wire _w2323_ ;
	wire _w2322_ ;
	wire _w2321_ ;
	wire _w2320_ ;
	wire _w2319_ ;
	wire _w2318_ ;
	wire _w2317_ ;
	wire _w2316_ ;
	wire _w2315_ ;
	wire _w2314_ ;
	wire _w2313_ ;
	wire _w2312_ ;
	wire _w2311_ ;
	wire _w2310_ ;
	wire _w2309_ ;
	wire _w2308_ ;
	wire _w2307_ ;
	wire _w2306_ ;
	wire _w2305_ ;
	wire _w2304_ ;
	wire _w2303_ ;
	wire _w2302_ ;
	wire _w2301_ ;
	wire _w2300_ ;
	wire _w2299_ ;
	wire _w2298_ ;
	wire _w2297_ ;
	wire _w2296_ ;
	wire _w2295_ ;
	wire _w2294_ ;
	wire _w2293_ ;
	wire _w2292_ ;
	wire _w2291_ ;
	wire _w2290_ ;
	wire _w2289_ ;
	wire _w2288_ ;
	wire _w2287_ ;
	wire _w2286_ ;
	wire _w2285_ ;
	wire _w2284_ ;
	wire _w2283_ ;
	wire _w2282_ ;
	wire _w2281_ ;
	wire _w2280_ ;
	wire _w2279_ ;
	wire _w2278_ ;
	wire _w2277_ ;
	wire _w2276_ ;
	wire _w2275_ ;
	wire _w2274_ ;
	wire _w2273_ ;
	wire _w2272_ ;
	wire _w2271_ ;
	wire _w2270_ ;
	wire _w2269_ ;
	wire _w2268_ ;
	wire _w2267_ ;
	wire _w2266_ ;
	wire _w2265_ ;
	wire _w2264_ ;
	wire _w2263_ ;
	wire _w2262_ ;
	wire _w2261_ ;
	wire _w2260_ ;
	wire _w2259_ ;
	wire _w2258_ ;
	wire _w2257_ ;
	wire _w2256_ ;
	wire _w2255_ ;
	wire _w2254_ ;
	wire _w2253_ ;
	wire _w2252_ ;
	wire _w2251_ ;
	wire _w2250_ ;
	wire _w2249_ ;
	wire _w2248_ ;
	wire _w2247_ ;
	wire _w2246_ ;
	wire _w2245_ ;
	wire _w2244_ ;
	wire _w2243_ ;
	wire _w2242_ ;
	wire _w2241_ ;
	wire _w2240_ ;
	wire _w2239_ ;
	wire _w2238_ ;
	wire _w2237_ ;
	wire _w2236_ ;
	wire _w2235_ ;
	wire _w2234_ ;
	wire _w2233_ ;
	wire _w2232_ ;
	wire _w2231_ ;
	wire _w2230_ ;
	wire _w2229_ ;
	wire _w2228_ ;
	wire _w2227_ ;
	wire _w2226_ ;
	wire _w2225_ ;
	wire _w2224_ ;
	wire _w2223_ ;
	wire _w2222_ ;
	wire _w2221_ ;
	wire _w2220_ ;
	wire _w2219_ ;
	wire _w2218_ ;
	wire _w2217_ ;
	wire _w2216_ ;
	wire _w2215_ ;
	wire _w2214_ ;
	wire _w2213_ ;
	wire _w2212_ ;
	wire _w2211_ ;
	wire _w2210_ ;
	wire _w2209_ ;
	wire _w2208_ ;
	wire _w2207_ ;
	wire _w2206_ ;
	wire _w2205_ ;
	wire _w2204_ ;
	wire _w2203_ ;
	wire _w2202_ ;
	wire _w2201_ ;
	wire _w2200_ ;
	wire _w2199_ ;
	wire _w2198_ ;
	wire _w2197_ ;
	wire _w2196_ ;
	wire _w2195_ ;
	wire _w2194_ ;
	wire _w2193_ ;
	wire _w2192_ ;
	wire _w2191_ ;
	wire _w2190_ ;
	wire _w2189_ ;
	wire _w2188_ ;
	wire _w2187_ ;
	wire _w2186_ ;
	wire _w2185_ ;
	wire _w2184_ ;
	wire _w2183_ ;
	wire _w2182_ ;
	wire _w2181_ ;
	wire _w2180_ ;
	wire _w2179_ ;
	wire _w2178_ ;
	wire _w2177_ ;
	wire _w2176_ ;
	wire _w2175_ ;
	wire _w2174_ ;
	wire _w2173_ ;
	wire _w2172_ ;
	wire _w2171_ ;
	wire _w2170_ ;
	wire _w2169_ ;
	wire _w2168_ ;
	wire _w2167_ ;
	wire _w2166_ ;
	wire _w2165_ ;
	wire _w2164_ ;
	wire _w2163_ ;
	wire _w2162_ ;
	wire _w2161_ ;
	wire _w2160_ ;
	wire _w2159_ ;
	wire _w2158_ ;
	wire _w2027_ ;
	wire _w2026_ ;
	wire _w2025_ ;
	wire _w2024_ ;
	wire _w2023_ ;
	wire _w2022_ ;
	wire _w2021_ ;
	wire _w2020_ ;
	wire _w2019_ ;
	wire _w2018_ ;
	wire _w2017_ ;
	wire _w2016_ ;
	wire _w2015_ ;
	wire _w2014_ ;
	wire _w2013_ ;
	wire _w2012_ ;
	wire _w2011_ ;
	wire _w2010_ ;
	wire _w2009_ ;
	wire _w2008_ ;
	wire _w2007_ ;
	wire _w2006_ ;
	wire _w2005_ ;
	wire _w2004_ ;
	wire _w2003_ ;
	wire _w2002_ ;
	wire _w2001_ ;
	wire _w2000_ ;
	wire _w1999_ ;
	wire _w1998_ ;
	wire _w1997_ ;
	wire _w1996_ ;
	wire _w1995_ ;
	wire _w1994_ ;
	wire _w1993_ ;
	wire _w1992_ ;
	wire _w1991_ ;
	wire _w1990_ ;
	wire _w1989_ ;
	wire _w1988_ ;
	wire _w1987_ ;
	wire _w1986_ ;
	wire _w1985_ ;
	wire _w1984_ ;
	wire _w1983_ ;
	wire _w1982_ ;
	wire _w1981_ ;
	wire _w1980_ ;
	wire _w1979_ ;
	wire _w1978_ ;
	wire _w1977_ ;
	wire _w1976_ ;
	wire _w1975_ ;
	wire _w1974_ ;
	wire _w1973_ ;
	wire _w1972_ ;
	wire _w1971_ ;
	wire _w1970_ ;
	wire _w1969_ ;
	wire _w1968_ ;
	wire _w1967_ ;
	wire _w1966_ ;
	wire _w1965_ ;
	wire _w1964_ ;
	wire _w1963_ ;
	wire _w1962_ ;
	wire _w1961_ ;
	wire _w1960_ ;
	wire _w1929_ ;
	wire _w1928_ ;
	wire _w1927_ ;
	wire _w1926_ ;
	wire _w1925_ ;
	wire _w1924_ ;
	wire _w1923_ ;
	wire _w1922_ ;
	wire _w1921_ ;
	wire _w1920_ ;
	wire _w1919_ ;
	wire _w1918_ ;
	wire _w1917_ ;
	wire _w1916_ ;
	wire _w1915_ ;
	wire _w1914_ ;
	wire _w1901_ ;
	wire _w1902_ ;
	wire _w1903_ ;
	wire _w1904_ ;
	wire _w1905_ ;
	wire _w1906_ ;
	wire _w1907_ ;
	wire _w1908_ ;
	wire _w1909_ ;
	wire _w1910_ ;
	wire _w1911_ ;
	wire _w1912_ ;
	wire _w1913_ ;
	wire _w1930_ ;
	wire _w1931_ ;
	wire _w1932_ ;
	wire _w1933_ ;
	wire _w1934_ ;
	wire _w1935_ ;
	wire _w1936_ ;
	wire _w1937_ ;
	wire _w1938_ ;
	wire _w1939_ ;
	wire _w1940_ ;
	wire _w1941_ ;
	wire _w1942_ ;
	wire _w1943_ ;
	wire _w1944_ ;
	wire _w1945_ ;
	wire _w1946_ ;
	wire _w1947_ ;
	wire _w1948_ ;
	wire _w1949_ ;
	wire _w1950_ ;
	wire _w1951_ ;
	wire _w1952_ ;
	wire _w1953_ ;
	wire _w1954_ ;
	wire _w1955_ ;
	wire _w1956_ ;
	wire _w1957_ ;
	wire _w1958_ ;
	wire _w1959_ ;
	wire _w2028_ ;
	wire _w2029_ ;
	wire _w2030_ ;
	wire _w2031_ ;
	wire _w2032_ ;
	wire _w2033_ ;
	wire _w2034_ ;
	wire _w2035_ ;
	wire _w2036_ ;
	wire _w2037_ ;
	wire _w2038_ ;
	wire _w2039_ ;
	wire _w2040_ ;
	wire _w2041_ ;
	wire _w2042_ ;
	wire _w2043_ ;
	wire _w2044_ ;
	wire _w2045_ ;
	wire _w2046_ ;
	wire _w2047_ ;
	wire _w2048_ ;
	wire _w2049_ ;
	wire _w2050_ ;
	wire _w2051_ ;
	wire _w2052_ ;
	wire _w2053_ ;
	wire _w2054_ ;
	wire _w2055_ ;
	wire _w2056_ ;
	wire _w2057_ ;
	wire _w2058_ ;
	wire _w2059_ ;
	wire _w2060_ ;
	wire _w2061_ ;
	wire _w2062_ ;
	wire _w2063_ ;
	wire _w2064_ ;
	wire _w2065_ ;
	wire _w2066_ ;
	wire _w2067_ ;
	wire _w2068_ ;
	wire _w2069_ ;
	wire _w2070_ ;
	wire _w2071_ ;
	wire _w2072_ ;
	wire _w2073_ ;
	wire _w2074_ ;
	wire _w2075_ ;
	wire _w2076_ ;
	wire _w2077_ ;
	wire _w2078_ ;
	wire _w2079_ ;
	wire _w2080_ ;
	wire _w2081_ ;
	wire _w2082_ ;
	wire _w2083_ ;
	wire _w2084_ ;
	wire _w2085_ ;
	wire _w2086_ ;
	wire _w2087_ ;
	wire _w2088_ ;
	wire _w2089_ ;
	wire _w2090_ ;
	wire _w2091_ ;
	wire _w2092_ ;
	wire _w2093_ ;
	wire _w2094_ ;
	wire _w2095_ ;
	wire _w2096_ ;
	wire _w2097_ ;
	wire _w2098_ ;
	wire _w2099_ ;
	wire _w2100_ ;
	wire _w2101_ ;
	wire _w2102_ ;
	wire _w2103_ ;
	wire _w2104_ ;
	wire _w2105_ ;
	wire _w2106_ ;
	wire _w2107_ ;
	wire _w2108_ ;
	wire _w2109_ ;
	wire _w2110_ ;
	wire _w2111_ ;
	wire _w2112_ ;
	wire _w2113_ ;
	wire _w2114_ ;
	wire _w2115_ ;
	wire _w2116_ ;
	wire _w2117_ ;
	wire _w2118_ ;
	wire _w2119_ ;
	wire _w2120_ ;
	wire _w2121_ ;
	wire _w2122_ ;
	wire _w2123_ ;
	wire _w2124_ ;
	wire _w2125_ ;
	wire _w2126_ ;
	wire _w2127_ ;
	wire _w2128_ ;
	wire _w2129_ ;
	wire _w2130_ ;
	wire _w2131_ ;
	wire _w2132_ ;
	wire _w2133_ ;
	wire _w2134_ ;
	wire _w2135_ ;
	wire _w2136_ ;
	wire _w2137_ ;
	wire _w2138_ ;
	wire _w2139_ ;
	wire _w2140_ ;
	wire _w2141_ ;
	wire _w2142_ ;
	wire _w2143_ ;
	wire _w2144_ ;
	wire _w2145_ ;
	wire _w2146_ ;
	wire _w2147_ ;
	wire _w2148_ ;
	wire _w2149_ ;
	wire _w2150_ ;
	wire _w2151_ ;
	wire _w2152_ ;
	wire _w2153_ ;
	wire _w2154_ ;
	wire _w2155_ ;
	wire _w2156_ ;
	wire _w2157_ ;
	wire _w2442_ ;
	wire _w2443_ ;
	wire _w2444_ ;
	wire _w2445_ ;
	wire _w2446_ ;
	wire _w2447_ ;
	wire _w2448_ ;
	wire _w2449_ ;
	wire _w2450_ ;
	wire _w2451_ ;
	wire _w2452_ ;
	wire _w2453_ ;
	wire _w2454_ ;
	wire _w2455_ ;
	wire _w2456_ ;
	wire _w2457_ ;
	wire _w2458_ ;
	wire _w2459_ ;
	wire _w2460_ ;
	wire _w2461_ ;
	wire _w2462_ ;
	wire _w2463_ ;
	wire _w2464_ ;
	wire _w2465_ ;
	wire _w2466_ ;
	wire _w2467_ ;
	wire _w2468_ ;
	wire _w2469_ ;
	wire _w2470_ ;
	wire _w2471_ ;
	wire _w2472_ ;
	wire _w2473_ ;
	wire _w2474_ ;
	wire _w2475_ ;
	wire _w2476_ ;
	wire _w2477_ ;
	wire _w2478_ ;
	wire _w2479_ ;
	wire _w2480_ ;
	wire _w2481_ ;
	wire _w2482_ ;
	wire _w2483_ ;
	wire _w2484_ ;
	wire _w2485_ ;
	wire _w2486_ ;
	wire _w2487_ ;
	wire _w2488_ ;
	wire _w2489_ ;
	wire _w2490_ ;
	wire _w2491_ ;
	wire _w2492_ ;
	wire _w2493_ ;
	wire _w2494_ ;
	wire _w2495_ ;
	wire _w2496_ ;
	wire _w2497_ ;
	wire _w2498_ ;
	wire _w2499_ ;
	wire _w2500_ ;
	wire _w2501_ ;
	wire _w2502_ ;
	wire _w2503_ ;
	wire _w2504_ ;
	wire _w2505_ ;
	wire _w2506_ ;
	wire _w2507_ ;
	wire _w2508_ ;
	wire _w2509_ ;
	wire _w2510_ ;
	wire _w2511_ ;
	wire _w2512_ ;
	wire _w2513_ ;
	wire _w2514_ ;
	wire _w2515_ ;
	wire _w2516_ ;
	wire _w2517_ ;
	wire _w2518_ ;
	wire _w2519_ ;
	wire _w2520_ ;
	wire _w2521_ ;
	wire _w2522_ ;
	wire _w2523_ ;
	wire _w2524_ ;
	wire _w2525_ ;
	wire _w2526_ ;
	wire _w2527_ ;
	wire _w2528_ ;
	wire _w2529_ ;
	wire _w2530_ ;
	wire _w2531_ ;
	wire _w2532_ ;
	wire _w2533_ ;
	wire _w2534_ ;
	wire _w2535_ ;
	wire _w2536_ ;
	wire _w2537_ ;
	wire _w2538_ ;
	wire _w2539_ ;
	wire _w2540_ ;
	wire _w2541_ ;
	wire _w2542_ ;
	wire _w2543_ ;
	wire _w2544_ ;
	wire _w2545_ ;
	wire _w2546_ ;
	wire _w2547_ ;
	wire _w2548_ ;
	wire _w2549_ ;
	wire _w2550_ ;
	wire _w2551_ ;
	wire _w2552_ ;
	wire _w2553_ ;
	wire _w2554_ ;
	wire _w2555_ ;
	wire _w2556_ ;
	wire _w2557_ ;
	wire _w2558_ ;
	wire _w2559_ ;
	wire _w2560_ ;
	wire _w2561_ ;
	wire _w2562_ ;
	wire _w2563_ ;
	wire _w2564_ ;
	wire _w2565_ ;
	wire _w2566_ ;
	wire _w2567_ ;
	wire _w2568_ ;
	wire _w2569_ ;
	wire _w2570_ ;
	wire _w2571_ ;
	wire _w2572_ ;
	wire _w2573_ ;
	wire _w2574_ ;
	wire _w2575_ ;
	wire _w2576_ ;
	wire _w2577_ ;
	wire _w2578_ ;
	wire _w2579_ ;
	wire _w2580_ ;
	wire _w2581_ ;
	wire _w2582_ ;
	wire _w2583_ ;
	wire _w2584_ ;
	wire _w2585_ ;
	wire _w2586_ ;
	wire _w2587_ ;
	wire _w2588_ ;
	wire _w2589_ ;
	wire _w2590_ ;
	wire _w2591_ ;
	wire _w2592_ ;
	wire _w2593_ ;
	wire _w2594_ ;
	wire _w2595_ ;
	wire _w2596_ ;
	wire _w2597_ ;
	wire _w2598_ ;
	wire _w2599_ ;
	wire _w2600_ ;
	wire _w2601_ ;
	wire _w2602_ ;
	wire _w2603_ ;
	wire _w2604_ ;
	wire _w2605_ ;
	wire _w2606_ ;
	wire _w2607_ ;
	wire _w2608_ ;
	wire _w2609_ ;
	wire _w2610_ ;
	wire _w2611_ ;
	wire _w2612_ ;
	wire _w2613_ ;
	wire _w2614_ ;
	wire _w2615_ ;
	wire _w2616_ ;
	wire _w2617_ ;
	wire _w2618_ ;
	wire _w2619_ ;
	wire _w2620_ ;
	wire _w2621_ ;
	wire _w2622_ ;
	wire _w2623_ ;
	wire _w2624_ ;
	wire _w2625_ ;
	wire _w2626_ ;
	wire _w2627_ ;
	wire _w2628_ ;
	wire _w2629_ ;
	wire _w2630_ ;
	wire _w2631_ ;
	wire _w2632_ ;
	wire _w2633_ ;
	wire _w2634_ ;
	wire _w2635_ ;
	wire _w2636_ ;
	wire _w2637_ ;
	wire _w2638_ ;
	wire _w2639_ ;
	wire _w2640_ ;
	wire _w2641_ ;
	wire _w2642_ ;
	wire _w2643_ ;
	wire _w2644_ ;
	wire _w2645_ ;
	wire _w2646_ ;
	wire _w2647_ ;
	wire _w2648_ ;
	wire _w2649_ ;
	wire _w2650_ ;
	wire _w2651_ ;
	wire _w2652_ ;
	wire _w2653_ ;
	wire _w2654_ ;
	wire _w2655_ ;
	wire _w2656_ ;
	wire _w2657_ ;
	wire _w2658_ ;
	wire _w2659_ ;
	wire _w2660_ ;
	wire _w2661_ ;
	wire _w2662_ ;
	wire _w2663_ ;
	wire _w2664_ ;
	wire _w2665_ ;
	wire _w2666_ ;
	wire _w2667_ ;
	wire _w2668_ ;
	wire _w2669_ ;
	wire _w2670_ ;
	wire _w2671_ ;
	wire _w2672_ ;
	wire _w2673_ ;
	wire _w2674_ ;
	wire _w2675_ ;
	wire _w2676_ ;
	wire _w2677_ ;
	wire _w2678_ ;
	wire _w2679_ ;
	wire _w2680_ ;
	wire _w2681_ ;
	wire _w2682_ ;
	wire _w2683_ ;
	wire _w2684_ ;
	wire _w2685_ ;
	wire _w2686_ ;
	wire _w2687_ ;
	wire _w2688_ ;
	wire _w2689_ ;
	wire _w2690_ ;
	wire _w2691_ ;
	wire _w2692_ ;
	wire _w2693_ ;
	wire _w2694_ ;
	wire _w2695_ ;
	wire _w2696_ ;
	wire _w2697_ ;
	wire _w2698_ ;
	wire _w2699_ ;
	wire _w2700_ ;
	wire _w2701_ ;
	wire _w2702_ ;
	wire _w2703_ ;
	wire _w2704_ ;
	wire _w2705_ ;
	wire _w2706_ ;
	wire _w2707_ ;
	wire _w2708_ ;
	wire _w2709_ ;
	wire _w2710_ ;
	wire _w2711_ ;
	wire _w2712_ ;
	wire _w2713_ ;
	wire _w2714_ ;
	wire _w2715_ ;
	wire _w2716_ ;
	wire _w2717_ ;
	wire _w2718_ ;
	wire _w2719_ ;
	wire _w2720_ ;
	wire _w2721_ ;
	wire _w2722_ ;
	wire _w2723_ ;
	wire _w2724_ ;
	wire _w2725_ ;
	wire _w2726_ ;
	wire _w2727_ ;
	wire _w2728_ ;
	wire _w2729_ ;
	wire _w2730_ ;
	wire _w2731_ ;
	wire _w2732_ ;
	wire _w2733_ ;
	wire _w2734_ ;
	wire _w2735_ ;
	wire _w2736_ ;
	wire _w2737_ ;
	wire _w2738_ ;
	wire _w2739_ ;
	wire _w2740_ ;
	wire _w2741_ ;
	wire _w2742_ ;
	wire _w2743_ ;
	wire _w2744_ ;
	wire _w2745_ ;
	wire _w2746_ ;
	wire _w2747_ ;
	wire _w2748_ ;
	wire _w2749_ ;
	wire _w2750_ ;
	wire _w2751_ ;
	wire _w2752_ ;
	wire _w2753_ ;
	wire _w2754_ ;
	wire _w2755_ ;
	wire _w2756_ ;
	wire _w2757_ ;
	wire _w2758_ ;
	wire _w2759_ ;
	wire _w2760_ ;
	wire _w2761_ ;
	wire _w2762_ ;
	wire _w2763_ ;
	wire _w2764_ ;
	wire _w2765_ ;
	wire _w2766_ ;
	wire _w2767_ ;
	wire _w2768_ ;
	wire _w2769_ ;
	wire _w2770_ ;
	wire _w2771_ ;
	wire _w2772_ ;
	wire _w2773_ ;
	wire _w2774_ ;
	wire _w2775_ ;
	wire _w2776_ ;
	wire _w2777_ ;
	wire _w2778_ ;
	wire _w2779_ ;
	wire _w2780_ ;
	wire _w2781_ ;
	wire _w2782_ ;
	wire _w2783_ ;
	wire _w2784_ ;
	wire _w2785_ ;
	wire _w2786_ ;
	wire _w2787_ ;
	wire _w2788_ ;
	wire _w2789_ ;
	wire _w2790_ ;
	wire _w2791_ ;
	wire _w2792_ ;
	wire _w2793_ ;
	wire _w2794_ ;
	wire _w2795_ ;
	wire _w2796_ ;
	wire _w2797_ ;
	wire _w2798_ ;
	wire _w2799_ ;
	wire _w2800_ ;
	wire _w2801_ ;
	wire _w2802_ ;
	wire _w2803_ ;
	wire _w2804_ ;
	wire _w2805_ ;
	wire _w2806_ ;
	wire _w2807_ ;
	wire _w2808_ ;
	wire _w2809_ ;
	wire _w2810_ ;
	wire _w2811_ ;
	wire _w2812_ ;
	wire _w2813_ ;
	wire _w2814_ ;
	wire _w2815_ ;
	wire _w2816_ ;
	wire _w2817_ ;
	wire _w2818_ ;
	wire _w2819_ ;
	wire _w2820_ ;
	wire _w2821_ ;
	wire _w2822_ ;
	wire _w2823_ ;
	wire _w2824_ ;
	wire _w2825_ ;
	wire _w2826_ ;
	wire _w2827_ ;
	wire _w2828_ ;
	wire _w2829_ ;
	wire _w2830_ ;
	wire _w2831_ ;
	wire _w2832_ ;
	wire _w2833_ ;
	wire _w2834_ ;
	wire _w2835_ ;
	wire _w2836_ ;
	wire _w2837_ ;
	wire _w2838_ ;
	wire _w2839_ ;
	wire _w2840_ ;
	wire _w2841_ ;
	wire _w2842_ ;
	wire _w2843_ ;
	wire _w2844_ ;
	wire _w2845_ ;
	wire _w2846_ ;
	wire _w2847_ ;
	wire _w2848_ ;
	wire _w2849_ ;
	wire _w2850_ ;
	wire _w2851_ ;
	wire _w2852_ ;
	wire _w2853_ ;
	wire _w2854_ ;
	wire _w2855_ ;
	wire _w2856_ ;
	wire _w2857_ ;
	wire _w2858_ ;
	wire _w2859_ ;
	wire _w2860_ ;
	wire _w2861_ ;
	wire _w2862_ ;
	wire _w2863_ ;
	wire _w2864_ ;
	wire _w2865_ ;
	wire _w2866_ ;
	wire _w2867_ ;
	wire _w2868_ ;
	wire _w2869_ ;
	wire _w2870_ ;
	wire _w2871_ ;
	wire _w2872_ ;
	wire _w2873_ ;
	wire _w2874_ ;
	wire _w2875_ ;
	wire _w2876_ ;
	wire _w2877_ ;
	wire _w2878_ ;
	wire _w2879_ ;
	wire _w2880_ ;
	wire _w2881_ ;
	wire _w2882_ ;
	wire _w2883_ ;
	wire _w2884_ ;
	wire _w2885_ ;
	wire _w2886_ ;
	wire _w2887_ ;
	wire _w2888_ ;
	wire _w2889_ ;
	wire _w2890_ ;
	wire _w2891_ ;
	wire _w2892_ ;
	wire _w2893_ ;
	wire _w2894_ ;
	wire _w2895_ ;
	wire _w2896_ ;
	wire _w2897_ ;
	wire _w2898_ ;
	wire _w2899_ ;
	wire _w2900_ ;
	wire _w2901_ ;
	wire _w2902_ ;
	wire _w2903_ ;
	wire _w2904_ ;
	wire _w2905_ ;
	wire _w2906_ ;
	wire _w2907_ ;
	wire _w2908_ ;
	wire _w2909_ ;
	wire _w2910_ ;
	wire _w2911_ ;
	wire _w2912_ ;
	wire _w2913_ ;
	wire _w2914_ ;
	wire _w2915_ ;
	wire _w2916_ ;
	wire _w2917_ ;
	wire _w2918_ ;
	wire _w2919_ ;
	wire _w2920_ ;
	wire _w2921_ ;
	wire _w2922_ ;
	wire _w2923_ ;
	wire _w2924_ ;
	wire _w2925_ ;
	wire _w2926_ ;
	wire _w2927_ ;
	wire _w2928_ ;
	wire _w2929_ ;
	wire _w2930_ ;
	wire _w2931_ ;
	wire _w2932_ ;
	wire _w2933_ ;
	wire _w2934_ ;
	wire _w2935_ ;
	wire _w2936_ ;
	wire _w2937_ ;
	wire _w2938_ ;
	wire _w2939_ ;
	wire _w2940_ ;
	wire _w2941_ ;
	wire _w2942_ ;
	wire _w2943_ ;
	wire _w2944_ ;
	wire _w2945_ ;
	wire _w2946_ ;
	wire _w2947_ ;
	wire _w2948_ ;
	wire _w2949_ ;
	wire _w2950_ ;
	wire _w2951_ ;
	wire _w2952_ ;
	wire _w2953_ ;
	wire _w2954_ ;
	wire _w2955_ ;
	wire _w2956_ ;
	wire _w2957_ ;
	wire _w2958_ ;
	wire _w2959_ ;
	wire _w2960_ ;
	wire _w2961_ ;
	wire _w2962_ ;
	wire _w2963_ ;
	wire _w2964_ ;
	wire _w2965_ ;
	wire _w2966_ ;
	wire _w2967_ ;
	wire _w2968_ ;
	wire _w2969_ ;
	wire _w2970_ ;
	wire _w2971_ ;
	wire _w2972_ ;
	wire _w2973_ ;
	wire _w2974_ ;
	wire _w2975_ ;
	wire _w2976_ ;
	wire _w2977_ ;
	wire _w2978_ ;
	wire _w2979_ ;
	wire _w2980_ ;
	wire _w2981_ ;
	wire _w2982_ ;
	wire _w2983_ ;
	wire _w2984_ ;
	wire _w2985_ ;
	wire _w2986_ ;
	wire _w2987_ ;
	wire _w2988_ ;
	wire _w2989_ ;
	wire _w2990_ ;
	wire _w2991_ ;
	wire _w2992_ ;
	wire _w2993_ ;
	wire _w2994_ ;
	wire _w2995_ ;
	wire _w2996_ ;
	wire _w2997_ ;
	wire _w2998_ ;
	wire _w2999_ ;
	wire _w3000_ ;
	wire _w3001_ ;
	wire _w3002_ ;
	wire _w3003_ ;
	wire _w3004_ ;
	wire _w3005_ ;
	wire _w3006_ ;
	wire _w3007_ ;
	wire _w3008_ ;
	wire _w3009_ ;
	wire _w4258_ ;
	wire _w4259_ ;
	wire _w4260_ ;
	wire _w4261_ ;
	wire _w4262_ ;
	wire _w4263_ ;
	wire _w4264_ ;
	wire _w4265_ ;
	wire _w4266_ ;
	wire _w4267_ ;
	wire _w4268_ ;
	wire _w4269_ ;
	wire _w4270_ ;
	wire _w4271_ ;
	wire _w4272_ ;
	wire _w4273_ ;
	wire _w4274_ ;
	wire _w4275_ ;
	wire _w4276_ ;
	wire _w4277_ ;
	wire _w4278_ ;
	wire _w4279_ ;
	wire _w4280_ ;
	wire _w4281_ ;
	wire _w4282_ ;
	wire _w4283_ ;
	wire _w4284_ ;
	wire _w4285_ ;
	wire _w4286_ ;
	wire _w4287_ ;
	wire _w4288_ ;
	wire _w4289_ ;
	wire _w4290_ ;
	wire _w4291_ ;
	wire _w4292_ ;
	wire _w4293_ ;
	wire _w4294_ ;
	wire _w4295_ ;
	wire _w4296_ ;
	wire _w4297_ ;
	wire _w4298_ ;
	wire _w4299_ ;
	wire _w4300_ ;
	wire _w4301_ ;
	wire _w4302_ ;
	wire _w4303_ ;
	wire _w4304_ ;
	wire _w4305_ ;
	wire _w4306_ ;
	wire _w4307_ ;
	wire _w4308_ ;
	wire _w4309_ ;
	wire _w4310_ ;
	wire _w4311_ ;
	wire _w4312_ ;
	wire _w4313_ ;
	wire _w4314_ ;
	wire _w4315_ ;
	wire _w4316_ ;
	wire _w4317_ ;
	wire _w4318_ ;
	wire _w4319_ ;
	wire _w4320_ ;
	wire _w4321_ ;
	wire _w4322_ ;
	wire _w4323_ ;
	wire _w4324_ ;
	wire _w4325_ ;
	wire _w4326_ ;
	wire _w4327_ ;
	wire _w4328_ ;
	wire _w4329_ ;
	wire _w4330_ ;
	wire _w4331_ ;
	wire _w4332_ ;
	wire _w4333_ ;
	wire _w4334_ ;
	wire _w4335_ ;
	wire _w4336_ ;
	wire _w4337_ ;
	wire _w4338_ ;
	wire _w4339_ ;
	wire _w4340_ ;
	wire _w4341_ ;
	wire _w4342_ ;
	wire _w4343_ ;
	wire _w4344_ ;
	wire _w4345_ ;
	wire _w4346_ ;
	wire _w4347_ ;
	wire _w4348_ ;
	wire _w4349_ ;
	wire _w4350_ ;
	wire _w4351_ ;
	wire _w4352_ ;
	wire _w4353_ ;
	wire _w4354_ ;
	wire _w4355_ ;
	wire _w4356_ ;
	wire _w4357_ ;
	wire _w4358_ ;
	wire _w4359_ ;
	wire _w4360_ ;
	wire _w4361_ ;
	wire _w4362_ ;
	wire _w4363_ ;
	wire _w4364_ ;
	wire _w4365_ ;
	wire _w4366_ ;
	wire _w4367_ ;
	wire _w4368_ ;
	wire _w4369_ ;
	wire _w4370_ ;
	wire _w4371_ ;
	wire _w4372_ ;
	wire _w4373_ ;
	wire _w4374_ ;
	wire _w4375_ ;
	wire _w4376_ ;
	wire _w4377_ ;
	wire _w4378_ ;
	wire _w4379_ ;
	wire _w4380_ ;
	wire _w4381_ ;
	wire _w4382_ ;
	wire _w4383_ ;
	wire _w4384_ ;
	wire _w4385_ ;
	wire _w4386_ ;
	wire _w4387_ ;
	wire _w4388_ ;
	wire _w4389_ ;
	wire _w4390_ ;
	wire _w4391_ ;
	wire _w4392_ ;
	wire _w4393_ ;
	wire _w4394_ ;
	wire _w4395_ ;
	wire _w4396_ ;
	wire _w4397_ ;
	wire _w4398_ ;
	wire _w4399_ ;
	wire _w4400_ ;
	wire _w4401_ ;
	wire _w4402_ ;
	wire _w4403_ ;
	wire _w4404_ ;
	wire _w4405_ ;
	wire _w4406_ ;
	wire _w4407_ ;
	wire _w4408_ ;
	wire _w4409_ ;
	wire _w4410_ ;
	wire _w4411_ ;
	wire _w4412_ ;
	wire _w4413_ ;
	wire _w4414_ ;
	wire _w4415_ ;
	wire _w4416_ ;
	wire _w4417_ ;
	wire _w4418_ ;
	wire _w4419_ ;
	wire _w4420_ ;
	wire _w4421_ ;
	wire _w4422_ ;
	wire _w4423_ ;
	wire _w4424_ ;
	wire _w4425_ ;
	wire _w4426_ ;
	wire _w4427_ ;
	wire _w4428_ ;
	wire _w4429_ ;
	wire _w4430_ ;
	wire _w4431_ ;
	wire _w4432_ ;
	wire _w4433_ ;
	wire _w4434_ ;
	wire _w4435_ ;
	wire _w4436_ ;
	wire _w4437_ ;
	wire _w4438_ ;
	wire _w4439_ ;
	wire _w4440_ ;
	wire _w4441_ ;
	wire _w4442_ ;
	wire _w4443_ ;
	wire _w4444_ ;
	wire _w4445_ ;
	wire _w4446_ ;
	wire _w4447_ ;
	wire _w4448_ ;
	wire _w4449_ ;
	wire _w4450_ ;
	wire _w4451_ ;
	wire _w4452_ ;
	wire _w4453_ ;
	wire _w4454_ ;
	wire _w4455_ ;
	wire _w4456_ ;
	wire _w4457_ ;
	wire _w4458_ ;
	wire _w4459_ ;
	wire _w4460_ ;
	wire _w4461_ ;
	wire _w4462_ ;
	wire _w4463_ ;
	wire _w4464_ ;
	wire _w4465_ ;
	wire _w4466_ ;
	wire _w4467_ ;
	wire _w4468_ ;
	wire _w4469_ ;
	wire _w4470_ ;
	wire _w4471_ ;
	wire _w4472_ ;
	wire _w4473_ ;
	wire _w4474_ ;
	wire _w4475_ ;
	wire _w4476_ ;
	wire _w4477_ ;
	wire _w4478_ ;
	wire _w4479_ ;
	wire _w4480_ ;
	wire _w4481_ ;
	wire _w4482_ ;
	wire _w4483_ ;
	wire _w4484_ ;
	wire _w4485_ ;
	wire _w4486_ ;
	wire _w4487_ ;
	wire _w4488_ ;
	wire _w4489_ ;
	wire _w4490_ ;
	wire _w4491_ ;
	wire _w4492_ ;
	wire _w4493_ ;
	wire _w4494_ ;
	wire _w4495_ ;
	wire _w4496_ ;
	wire _w4497_ ;
	wire _w4498_ ;
	wire _w4499_ ;
	wire _w4500_ ;
	wire _w4501_ ;
	wire _w4502_ ;
	wire _w4503_ ;
	wire _w4504_ ;
	wire _w4505_ ;
	wire _w4506_ ;
	wire _w4507_ ;
	wire _w4508_ ;
	wire _w4509_ ;
	wire _w4510_ ;
	wire _w4511_ ;
	wire _w4512_ ;
	wire _w4513_ ;
	wire _w4514_ ;
	wire _w4515_ ;
	wire _w4516_ ;
	wire _w4517_ ;
	wire _w4518_ ;
	wire _w4519_ ;
	wire _w4520_ ;
	wire _w4521_ ;
	wire _w4522_ ;
	wire _w4523_ ;
	wire _w4524_ ;
	wire _w4525_ ;
	wire _w4526_ ;
	wire _w4527_ ;
	wire _w4528_ ;
	wire _w4529_ ;
	wire _w4530_ ;
	wire _w4531_ ;
	wire _w4532_ ;
	wire _w4533_ ;
	wire _w4534_ ;
	wire _w4535_ ;
	wire _w4536_ ;
	wire _w4537_ ;
	wire _w4538_ ;
	wire _w4539_ ;
	wire _w4540_ ;
	wire _w4541_ ;
	wire _w4542_ ;
	wire _w4543_ ;
	wire _w4544_ ;
	wire _w4545_ ;
	wire _w4546_ ;
	wire _w4547_ ;
	wire _w4548_ ;
	wire _w4549_ ;
	wire _w4550_ ;
	wire _w4551_ ;
	wire _w4552_ ;
	wire _w4553_ ;
	wire _w4554_ ;
	wire _w4555_ ;
	wire _w4556_ ;
	wire _w4557_ ;
	wire _w4558_ ;
	wire _w4559_ ;
	wire _w4560_ ;
	wire _w4561_ ;
	wire _w4562_ ;
	wire _w4563_ ;
	wire _w4564_ ;
	wire _w4565_ ;
	wire _w4566_ ;
	wire _w4567_ ;
	wire _w4568_ ;
	wire _w4569_ ;
	wire _w4570_ ;
	wire _w4571_ ;
	wire _w4572_ ;
	wire _w4573_ ;
	wire _w4574_ ;
	wire _w4575_ ;
	wire _w4576_ ;
	wire _w4577_ ;
	wire _w4578_ ;
	wire _w4579_ ;
	wire _w4580_ ;
	wire _w4581_ ;
	wire _w4582_ ;
	wire _w4583_ ;
	wire _w4584_ ;
	wire _w4585_ ;
	wire _w4586_ ;
	wire _w4587_ ;
	wire _w4588_ ;
	wire _w4589_ ;
	wire _w4590_ ;
	wire _w4591_ ;
	wire _w4592_ ;
	wire _w4593_ ;
	wire _w4594_ ;
	wire _w4595_ ;
	wire _w4596_ ;
	wire _w4597_ ;
	wire _w4598_ ;
	wire _w4599_ ;
	wire _w4600_ ;
	wire _w4601_ ;
	wire _w4602_ ;
	wire _w4603_ ;
	wire _w4604_ ;
	wire _w4605_ ;
	wire _w4606_ ;
	wire _w4607_ ;
	wire _w4608_ ;
	wire _w4609_ ;
	wire _w4610_ ;
	wire _w4611_ ;
	wire _w4612_ ;
	wire _w4613_ ;
	wire _w4614_ ;
	wire _w4615_ ;
	wire _w4616_ ;
	wire _w4617_ ;
	wire _w4618_ ;
	wire _w4619_ ;
	wire _w4620_ ;
	wire _w4621_ ;
	wire _w4622_ ;
	wire _w4623_ ;
	wire _w4624_ ;
	wire _w4625_ ;
	wire _w4626_ ;
	wire _w4627_ ;
	wire _w4628_ ;
	wire _w4629_ ;
	wire _w4630_ ;
	wire _w4631_ ;
	wire _w4632_ ;
	wire _w4633_ ;
	wire _w4634_ ;
	wire _w4635_ ;
	wire _w4636_ ;
	wire _w4637_ ;
	wire _w4638_ ;
	wire _w4639_ ;
	wire _w4640_ ;
	wire _w4641_ ;
	wire _w4642_ ;
	wire _w4643_ ;
	wire _w4644_ ;
	wire _w4645_ ;
	wire _w4646_ ;
	wire _w4647_ ;
	wire _w4648_ ;
	wire _w4649_ ;
	wire _w4650_ ;
	wire _w4651_ ;
	wire _w4652_ ;
	wire _w4653_ ;
	wire _w4654_ ;
	wire _w4655_ ;
	wire _w4656_ ;
	wire _w4657_ ;
	wire _w4658_ ;
	wire _w4659_ ;
	wire _w4660_ ;
	wire _w4661_ ;
	wire _w4662_ ;
	wire _w4663_ ;
	wire _w4664_ ;
	wire _w4665_ ;
	wire _w4666_ ;
	wire _w4667_ ;
	wire _w4668_ ;
	wire _w4669_ ;
	wire _w4670_ ;
	wire _w4671_ ;
	wire _w4672_ ;
	wire _w4673_ ;
	wire _w4674_ ;
	wire _w4675_ ;
	wire _w4676_ ;
	wire _w4677_ ;
	wire _w4678_ ;
	wire _w4679_ ;
	wire _w4680_ ;
	wire _w4681_ ;
	wire _w4682_ ;
	wire _w4683_ ;
	wire _w4684_ ;
	wire _w4685_ ;
	wire _w4686_ ;
	wire _w4687_ ;
	wire _w4688_ ;
	wire _w4689_ ;
	wire _w4690_ ;
	wire _w4691_ ;
	wire _w4692_ ;
	wire _w4693_ ;
	wire _w4694_ ;
	wire _w4695_ ;
	wire _w4696_ ;
	wire _w4697_ ;
	wire _w4698_ ;
	wire _w4699_ ;
	wire _w4700_ ;
	wire _w4701_ ;
	wire _w4702_ ;
	wire _w4703_ ;
	wire _w4704_ ;
	wire _w4705_ ;
	wire _w4706_ ;
	wire _w4707_ ;
	wire _w4708_ ;
	wire _w4709_ ;
	wire _w4710_ ;
	wire _w4711_ ;
	wire _w4712_ ;
	wire _w4713_ ;
	wire _w4714_ ;
	wire _w4715_ ;
	wire _w4716_ ;
	wire _w4717_ ;
	wire _w4718_ ;
	wire _w4719_ ;
	wire _w4720_ ;
	wire _w4721_ ;
	wire _w4722_ ;
	wire _w4723_ ;
	wire _w4724_ ;
	wire _w4725_ ;
	wire _w4726_ ;
	wire _w4727_ ;
	wire _w4728_ ;
	wire _w4729_ ;
	wire _w4730_ ;
	wire _w4731_ ;
	wire _w4732_ ;
	wire _w4733_ ;
	wire _w4734_ ;
	wire _w4735_ ;
	wire _w4736_ ;
	wire _w4737_ ;
	wire _w4738_ ;
	wire _w4739_ ;
	wire _w4740_ ;
	wire _w4741_ ;
	wire _w4742_ ;
	wire _w4743_ ;
	wire _w4744_ ;
	wire _w4745_ ;
	wire _w4746_ ;
	wire _w4747_ ;
	wire _w4748_ ;
	wire _w4749_ ;
	wire _w4750_ ;
	wire _w4751_ ;
	wire _w4752_ ;
	wire _w4753_ ;
	wire _w4754_ ;
	wire _w4755_ ;
	wire _w4756_ ;
	wire _w4757_ ;
	wire _w4758_ ;
	wire _w4759_ ;
	wire _w4760_ ;
	wire _w4761_ ;
	wire _w4762_ ;
	wire _w4763_ ;
	wire _w4764_ ;
	wire _w4765_ ;
	wire _w4766_ ;
	wire _w4767_ ;
	wire _w4768_ ;
	wire _w4769_ ;
	wire _w4770_ ;
	wire _w4771_ ;
	wire _w4772_ ;
	wire _w4773_ ;
	wire _w4774_ ;
	wire _w4775_ ;
	wire _w4776_ ;
	wire _w4777_ ;
	wire _w4778_ ;
	wire _w4779_ ;
	wire _w4780_ ;
	wire _w4781_ ;
	wire _w4782_ ;
	wire _w4783_ ;
	wire _w4784_ ;
	wire _w4785_ ;
	wire _w4786_ ;
	wire _w4787_ ;
	wire _w4788_ ;
	wire _w4789_ ;
	wire _w4790_ ;
	wire _w4791_ ;
	wire _w4792_ ;
	wire _w4793_ ;
	wire _w4794_ ;
	wire _w4795_ ;
	wire _w4796_ ;
	wire _w4797_ ;
	wire _w4798_ ;
	wire _w4799_ ;
	wire _w4800_ ;
	wire _w4801_ ;
	wire _w4802_ ;
	wire _w4803_ ;
	wire _w4804_ ;
	wire _w4805_ ;
	wire _w4806_ ;
	wire _w4807_ ;
	wire _w4808_ ;
	wire _w4809_ ;
	wire _w4810_ ;
	wire _w4811_ ;
	wire _w4812_ ;
	wire _w4813_ ;
	wire _w4814_ ;
	wire _w4815_ ;
	wire _w4816_ ;
	wire _w4817_ ;
	wire _w4818_ ;
	wire _w4819_ ;
	wire _w4820_ ;
	wire _w4821_ ;
	wire _w4822_ ;
	wire _w4823_ ;
	wire _w4824_ ;
	wire _w4825_ ;
	wire _w4826_ ;
	wire _w4827_ ;
	wire _w4828_ ;
	wire _w4829_ ;
	wire _w4830_ ;
	wire _w4831_ ;
	wire _w4832_ ;
	wire _w4833_ ;
	wire _w4834_ ;
	wire _w4835_ ;
	wire _w4836_ ;
	wire _w4837_ ;
	wire _w4838_ ;
	wire _w4839_ ;
	wire _w4840_ ;
	wire _w4841_ ;
	wire _w4842_ ;
	wire _w4843_ ;
	wire _w4844_ ;
	wire _w4845_ ;
	wire _w4846_ ;
	wire _w4847_ ;
	wire _w4848_ ;
	wire _w4849_ ;
	wire _w4850_ ;
	wire _w4851_ ;
	wire _w4852_ ;
	wire _w4853_ ;
	wire _w4854_ ;
	wire _w4855_ ;
	wire _w4856_ ;
	wire _w4857_ ;
	wire _w4858_ ;
	wire _w4859_ ;
	wire _w4860_ ;
	wire _w4861_ ;
	wire _w4862_ ;
	wire _w4863_ ;
	wire _w4864_ ;
	wire _w4865_ ;
	wire _w4866_ ;
	wire _w4867_ ;
	wire _w4868_ ;
	wire _w4869_ ;
	wire _w4870_ ;
	wire _w4871_ ;
	wire _w4872_ ;
	wire _w4873_ ;
	wire _w4874_ ;
	wire _w4875_ ;
	wire _w4876_ ;
	wire _w4877_ ;
	wire _w4878_ ;
	wire _w4879_ ;
	wire _w4880_ ;
	wire _w4881_ ;
	wire _w4882_ ;
	wire _w4883_ ;
	wire _w4884_ ;
	wire _w4885_ ;
	wire _w4886_ ;
	wire _w4887_ ;
	wire _w4888_ ;
	wire _w4889_ ;
	wire _w4890_ ;
	wire _w4891_ ;
	wire _w4892_ ;
	wire _w4893_ ;
	wire _w4894_ ;
	wire _w4895_ ;
	wire _w4896_ ;
	wire _w4897_ ;
	wire _w4898_ ;
	wire _w4899_ ;
	wire _w4900_ ;
	wire _w4901_ ;
	wire _w4902_ ;
	wire _w4903_ ;
	wire _w4904_ ;
	wire _w4905_ ;
	wire _w4906_ ;
	wire _w4907_ ;
	wire _w4908_ ;
	wire _w4909_ ;
	wire _w4910_ ;
	wire _w4911_ ;
	wire _w4912_ ;
	wire _w4913_ ;
	wire _w4914_ ;
	wire _w4915_ ;
	wire _w4916_ ;
	wire _w4917_ ;
	wire _w4918_ ;
	wire _w4919_ ;
	wire _w4920_ ;
	wire _w4921_ ;
	wire _w4922_ ;
	wire _w4923_ ;
	wire _w4924_ ;
	wire _w4925_ ;
	wire _w4926_ ;
	wire _w4927_ ;
	wire _w4928_ ;
	wire _w4929_ ;
	wire _w4930_ ;
	wire _w4931_ ;
	wire _w4932_ ;
	wire _w4933_ ;
	wire _w4934_ ;
	wire _w4935_ ;
	wire _w4936_ ;
	wire _w4937_ ;
	wire _w4938_ ;
	wire _w4939_ ;
	wire _w4940_ ;
	wire _w4941_ ;
	wire _w4942_ ;
	wire _w4943_ ;
	wire _w4944_ ;
	wire _w4945_ ;
	wire _w4946_ ;
	wire _w4947_ ;
	wire _w4948_ ;
	wire _w4949_ ;
	wire _w4950_ ;
	wire _w4951_ ;
	wire _w4952_ ;
	wire _w4953_ ;
	wire _w4954_ ;
	wire _w4955_ ;
	wire _w4956_ ;
	wire _w4957_ ;
	wire _w4958_ ;
	wire _w4959_ ;
	wire _w4960_ ;
	wire _w4961_ ;
	wire _w4962_ ;
	wire _w4963_ ;
	wire _w4964_ ;
	wire _w4965_ ;
	wire _w4966_ ;
	wire _w4967_ ;
	wire _w4968_ ;
	wire _w4969_ ;
	wire _w4970_ ;
	wire _w4971_ ;
	wire _w4972_ ;
	wire _w4973_ ;
	wire _w4974_ ;
	wire _w4975_ ;
	wire _w4976_ ;
	wire _w4977_ ;
	wire _w4978_ ;
	wire _w4979_ ;
	wire _w4980_ ;
	wire _w4981_ ;
	wire _w4982_ ;
	wire _w4983_ ;
	wire _w4984_ ;
	wire _w4985_ ;
	wire _w4986_ ;
	wire _w4987_ ;
	wire _w4988_ ;
	wire _w4989_ ;
	wire _w4990_ ;
	wire _w4991_ ;
	wire _w4992_ ;
	wire _w4993_ ;
	wire _w4994_ ;
	wire _w4995_ ;
	wire _w4996_ ;
	wire _w4997_ ;
	wire _w4998_ ;
	wire _w4999_ ;
	wire _w5000_ ;
	wire _w5001_ ;
	wire _w5002_ ;
	wire _w5003_ ;
	wire _w5004_ ;
	wire _w5005_ ;
	wire _w5006_ ;
	wire _w5007_ ;
	wire _w5008_ ;
	wire _w5009_ ;
	wire _w5010_ ;
	wire _w5011_ ;
	wire _w5012_ ;
	wire _w5013_ ;
	wire _w5014_ ;
	wire _w5015_ ;
	wire _w5016_ ;
	wire _w5017_ ;
	wire _w5018_ ;
	wire _w5019_ ;
	wire _w5020_ ;
	wire _w5021_ ;
	wire _w5022_ ;
	wire _w5023_ ;
	wire _w5024_ ;
	wire _w5025_ ;
	wire _w5026_ ;
	wire _w5027_ ;
	wire _w5028_ ;
	wire _w5029_ ;
	wire _w5030_ ;
	wire _w5031_ ;
	wire _w5032_ ;
	wire _w5033_ ;
	wire _w5034_ ;
	wire _w5035_ ;
	wire _w5036_ ;
	wire _w5037_ ;
	wire _w5038_ ;
	wire _w5039_ ;
	wire _w5040_ ;
	wire _w5041_ ;
	wire _w5042_ ;
	wire _w5043_ ;
	wire _w5044_ ;
	wire _w5045_ ;
	wire _w5046_ ;
	wire _w5047_ ;
	wire _w5048_ ;
	wire _w5049_ ;
	wire _w5050_ ;
	wire _w5051_ ;
	wire _w5052_ ;
	wire _w5053_ ;
	wire _w5054_ ;
	wire _w5055_ ;
	wire _w5056_ ;
	wire _w5057_ ;
	wire _w5058_ ;
	wire _w5059_ ;
	wire _w5060_ ;
	wire _w5061_ ;
	wire _w5062_ ;
	wire _w5063_ ;
	wire _w5064_ ;
	wire _w5065_ ;
	wire _w5066_ ;
	wire _w5067_ ;
	wire _w5068_ ;
	wire _w5069_ ;
	wire _w5070_ ;
	wire _w5071_ ;
	wire _w5072_ ;
	wire _w5073_ ;
	wire _w5074_ ;
	wire _w5075_ ;
	wire _w5076_ ;
	wire _w5077_ ;
	wire _w5078_ ;
	wire _w5079_ ;
	wire _w5080_ ;
	wire _w5081_ ;
	wire _w5082_ ;
	wire _w5083_ ;
	wire _w5084_ ;
	wire _w5085_ ;
	wire _w5086_ ;
	wire _w5087_ ;
	wire _w5088_ ;
	wire _w5089_ ;
	wire _w5090_ ;
	wire _w5091_ ;
	wire _w5092_ ;
	wire _w5093_ ;
	wire _w5094_ ;
	wire _w5095_ ;
	wire _w5096_ ;
	wire _w5097_ ;
	wire _w5098_ ;
	wire _w5099_ ;
	wire _w5100_ ;
	wire _w5101_ ;
	wire _w5102_ ;
	wire _w5103_ ;
	wire _w5104_ ;
	wire _w5105_ ;
	wire _w5106_ ;
	wire _w5107_ ;
	wire _w5108_ ;
	wire _w5109_ ;
	wire _w5110_ ;
	wire _w5111_ ;
	wire _w5112_ ;
	wire _w5113_ ;
	wire _w5114_ ;
	wire _w5115_ ;
	wire _w5116_ ;
	wire _w5117_ ;
	wire _w5118_ ;
	wire _w5119_ ;
	wire _w5120_ ;
	wire _w5121_ ;
	wire _w5122_ ;
	wire _w5123_ ;
	wire _w5124_ ;
	wire _w5125_ ;
	wire _w5126_ ;
	wire _w5127_ ;
	wire _w5128_ ;
	wire _w5129_ ;
	wire _w5130_ ;
	wire _w5131_ ;
	wire _w5132_ ;
	wire _w5133_ ;
	wire _w5134_ ;
	wire _w5135_ ;
	wire _w5136_ ;
	wire _w5137_ ;
	wire _w5138_ ;
	wire _w5139_ ;
	wire _w5140_ ;
	wire _w5141_ ;
	wire _w5142_ ;
	wire _w5143_ ;
	wire _w5144_ ;
	wire _w5145_ ;
	wire _w5146_ ;
	wire _w5147_ ;
	wire _w5148_ ;
	wire _w5149_ ;
	wire _w5150_ ;
	wire _w5151_ ;
	wire _w5152_ ;
	wire _w5153_ ;
	wire _w5154_ ;
	wire _w5155_ ;
	wire _w5156_ ;
	wire _w5157_ ;
	wire _w5158_ ;
	wire _w5159_ ;
	wire _w5160_ ;
	wire _w5161_ ;
	wire _w5162_ ;
	wire _w5163_ ;
	wire _w5164_ ;
	wire _w5165_ ;
	wire _w5166_ ;
	wire _w5167_ ;
	wire _w5168_ ;
	wire _w5169_ ;
	wire _w5170_ ;
	wire _w5171_ ;
	wire _w5172_ ;
	wire _w5173_ ;
	wire _w5174_ ;
	wire _w5175_ ;
	wire _w5176_ ;
	wire _w5177_ ;
	wire _w5178_ ;
	wire _w5179_ ;
	wire _w5180_ ;
	wire _w5181_ ;
	wire _w5182_ ;
	wire _w5183_ ;
	wire _w5184_ ;
	wire _w5185_ ;
	wire _w5186_ ;
	wire _w5187_ ;
	wire _w5188_ ;
	wire _w5189_ ;
	wire _w5190_ ;
	wire _w5191_ ;
	wire _w5192_ ;
	wire _w5193_ ;
	wire _w5194_ ;
	wire _w5195_ ;
	wire _w5196_ ;
	wire _w5197_ ;
	wire _w5198_ ;
	wire _w5199_ ;
	wire _w5200_ ;
	wire _w5201_ ;
	wire _w5202_ ;
	wire _w5203_ ;
	wire _w5204_ ;
	wire _w5205_ ;
	wire _w5206_ ;
	wire _w5207_ ;
	wire _w5208_ ;
	wire _w5209_ ;
	wire _w5210_ ;
	wire _w5211_ ;
	wire _w5212_ ;
	wire _w5213_ ;
	wire _w5214_ ;
	wire _w5215_ ;
	wire _w5216_ ;
	wire _w5217_ ;
	wire _w5218_ ;
	wire _w5219_ ;
	wire _w5220_ ;
	wire _w5221_ ;
	wire _w5222_ ;
	wire _w5223_ ;
	wire _w5224_ ;
	wire _w5225_ ;
	wire _w5226_ ;
	wire _w5227_ ;
	wire _w5228_ ;
	wire _w5229_ ;
	wire _w5230_ ;
	wire _w5231_ ;
	wire _w5232_ ;
	wire _w5233_ ;
	wire _w5234_ ;
	wire _w5235_ ;
	wire _w5236_ ;
	wire _w5237_ ;
	wire _w5238_ ;
	wire _w5239_ ;
	wire _w5240_ ;
	wire _w5241_ ;
	wire _w5242_ ;
	wire _w5243_ ;
	wire _w5244_ ;
	wire _w5245_ ;
	wire _w5246_ ;
	wire _w5247_ ;
	wire _w5248_ ;
	wire _w5249_ ;
	wire _w5250_ ;
	wire _w5251_ ;
	wire _w5252_ ;
	wire _w5253_ ;
	wire _w5254_ ;
	wire _w5255_ ;
	wire _w5256_ ;
	wire _w5257_ ;
	wire _w5258_ ;
	wire _w5259_ ;
	wire _w5260_ ;
	wire _w5261_ ;
	wire _w5262_ ;
	wire _w5263_ ;
	wire _w5264_ ;
	wire _w5265_ ;
	wire _w5266_ ;
	wire _w5267_ ;
	wire _w5268_ ;
	wire _w5269_ ;
	wire _w5270_ ;
	wire _w5271_ ;
	wire _w5272_ ;
	wire _w5273_ ;
	wire _w5274_ ;
	wire _w5275_ ;
	wire _w5276_ ;
	wire _w5277_ ;
	wire _w5278_ ;
	wire _w5279_ ;
	wire _w5280_ ;
	wire _w5281_ ;
	wire _w5282_ ;
	wire _w5283_ ;
	wire _w5284_ ;
	wire _w5285_ ;
	wire _w5286_ ;
	wire _w5287_ ;
	wire _w5288_ ;
	wire _w5289_ ;
	wire _w5290_ ;
	wire _w5291_ ;
	wire _w5292_ ;
	wire _w5293_ ;
	wire _w5294_ ;
	wire _w5295_ ;
	wire _w5296_ ;
	wire _w5297_ ;
	wire _w5298_ ;
	wire _w5299_ ;
	wire _w5300_ ;
	wire _w5301_ ;
	wire _w5302_ ;
	wire _w5303_ ;
	wire _w5304_ ;
	wire _w5305_ ;
	wire _w5306_ ;
	wire _w5307_ ;
	wire _w5308_ ;
	wire _w5309_ ;
	wire _w5310_ ;
	wire _w5311_ ;
	wire _w5312_ ;
	wire _w5313_ ;
	wire _w5314_ ;
	wire _w5315_ ;
	wire _w5316_ ;
	wire _w5317_ ;
	wire _w5318_ ;
	wire _w5319_ ;
	wire _w5320_ ;
	wire _w5321_ ;
	wire _w5322_ ;
	wire _w5323_ ;
	wire _w5324_ ;
	wire _w5325_ ;
	wire _w5326_ ;
	wire _w5327_ ;
	wire _w5328_ ;
	wire _w5329_ ;
	wire _w5330_ ;
	wire _w5331_ ;
	wire _w5332_ ;
	wire _w5333_ ;
	wire _w5334_ ;
	wire _w5335_ ;
	wire _w5336_ ;
	wire _w5337_ ;
	wire _w5338_ ;
	wire _w5339_ ;
	wire _w5340_ ;
	wire _w5341_ ;
	wire _w5342_ ;
	wire _w5343_ ;
	wire _w5344_ ;
	wire _w5345_ ;
	wire _w5346_ ;
	wire _w5347_ ;
	wire _w5348_ ;
	wire _w5349_ ;
	wire _w5350_ ;
	wire _w5351_ ;
	wire _w5352_ ;
	wire _w5353_ ;
	wire _w5354_ ;
	wire _w5355_ ;
	wire _w5356_ ;
	wire _w5357_ ;
	wire _w5358_ ;
	wire _w5359_ ;
	wire _w5360_ ;
	wire _w5361_ ;
	wire _w5362_ ;
	wire _w5363_ ;
	wire _w5364_ ;
	wire _w5365_ ;
	wire _w5366_ ;
	wire _w5367_ ;
	wire _w5368_ ;
	wire _w5369_ ;
	wire _w5370_ ;
	wire _w5371_ ;
	wire _w5372_ ;
	wire _w5373_ ;
	wire _w5374_ ;
	wire _w5375_ ;
	wire _w5376_ ;
	wire _w5377_ ;
	wire _w5378_ ;
	wire _w5379_ ;
	wire _w5380_ ;
	wire _w5381_ ;
	wire _w5382_ ;
	wire _w5383_ ;
	wire _w5384_ ;
	wire _w5385_ ;
	wire _w5386_ ;
	wire _w5387_ ;
	wire _w5388_ ;
	wire _w5389_ ;
	wire _w5390_ ;
	wire _w5391_ ;
	wire _w5392_ ;
	wire _w5393_ ;
	wire _w5394_ ;
	wire _w5395_ ;
	wire _w5396_ ;
	wire _w5397_ ;
	wire _w5398_ ;
	wire _w5399_ ;
	wire _w5400_ ;
	wire _w5401_ ;
	wire _w5402_ ;
	wire _w5403_ ;
	wire _w5404_ ;
	wire _w5405_ ;
	wire _w5406_ ;
	wire _w5407_ ;
	wire _w5408_ ;
	wire _w5409_ ;
	wire _w5410_ ;
	wire _w5411_ ;
	wire _w5412_ ;
	wire _w5413_ ;
	wire _w5414_ ;
	wire _w5415_ ;
	wire _w5416_ ;
	wire _w5417_ ;
	wire _w5418_ ;
	wire _w5419_ ;
	wire _w5420_ ;
	wire _w5421_ ;
	wire _w5422_ ;
	wire _w5423_ ;
	wire _w5424_ ;
	wire _w5425_ ;
	wire _w5426_ ;
	wire _w5427_ ;
	wire _w5428_ ;
	wire _w5429_ ;
	wire _w5430_ ;
	wire _w5431_ ;
	wire _w5432_ ;
	wire _w5433_ ;
	wire _w5434_ ;
	wire _w5435_ ;
	wire _w5436_ ;
	wire _w5437_ ;
	wire _w5438_ ;
	wire _w5439_ ;
	wire _w5440_ ;
	wire _w5441_ ;
	wire _w5442_ ;
	wire _w5443_ ;
	wire _w5444_ ;
	wire _w5445_ ;
	wire _w5446_ ;
	wire _w5447_ ;
	wire _w5448_ ;
	wire _w5449_ ;
	wire _w5450_ ;
	wire _w5451_ ;
	wire _w5452_ ;
	wire _w5453_ ;
	wire _w5454_ ;
	wire _w5455_ ;
	wire _w5456_ ;
	wire _w5457_ ;
	wire _w5458_ ;
	wire _w5459_ ;
	wire _w5460_ ;
	wire _w5461_ ;
	wire _w5462_ ;
	wire _w5463_ ;
	wire _w5464_ ;
	wire _w5465_ ;
	wire _w5466_ ;
	wire _w5467_ ;
	wire _w5468_ ;
	wire _w5469_ ;
	wire _w5470_ ;
	wire _w5471_ ;
	wire _w5472_ ;
	wire _w5473_ ;
	wire _w5474_ ;
	wire _w5475_ ;
	wire _w5476_ ;
	wire _w5477_ ;
	wire _w5478_ ;
	wire _w5479_ ;
	wire _w5480_ ;
	wire _w5481_ ;
	wire _w5482_ ;
	wire _w5483_ ;
	wire _w5484_ ;
	wire _w5485_ ;
	wire _w5486_ ;
	wire _w5487_ ;
	wire _w5488_ ;
	wire _w5489_ ;
	wire _w5490_ ;
	wire _w5491_ ;
	wire _w5492_ ;
	wire _w5493_ ;
	wire _w5494_ ;
	wire _w5495_ ;
	wire _w5496_ ;
	wire _w5497_ ;
	wire _w5498_ ;
	wire _w5499_ ;
	wire _w5500_ ;
	wire _w5501_ ;
	wire _w5502_ ;
	wire _w5503_ ;
	wire _w5504_ ;
	wire _w5505_ ;
	wire _w5506_ ;
	wire _w5507_ ;
	wire _w5508_ ;
	wire _w5509_ ;
	wire _w5510_ ;
	wire _w5511_ ;
	wire _w5512_ ;
	wire _w5513_ ;
	wire _w5514_ ;
	wire _w5515_ ;
	wire _w5516_ ;
	wire _w5517_ ;
	wire _w5518_ ;
	wire _w5519_ ;
	wire _w5520_ ;
	wire _w5521_ ;
	wire _w5522_ ;
	wire _w5523_ ;
	wire _w5524_ ;
	wire _w5525_ ;
	wire _w5526_ ;
	wire _w5527_ ;
	wire _w5528_ ;
	wire _w5529_ ;
	wire _w5530_ ;
	wire _w5531_ ;
	wire _w5532_ ;
	wire _w5533_ ;
	wire _w5534_ ;
	wire _w5535_ ;
	wire _w5536_ ;
	wire _w5537_ ;
	wire _w5538_ ;
	wire _w5539_ ;
	wire _w5540_ ;
	wire _w5541_ ;
	wire _w5542_ ;
	wire _w5543_ ;
	wire _w5544_ ;
	wire _w5545_ ;
	wire _w5546_ ;
	wire _w5547_ ;
	wire _w5548_ ;
	wire _w5549_ ;
	wire _w5550_ ;
	wire _w5551_ ;
	wire _w5552_ ;
	wire _w5553_ ;
	wire _w5554_ ;
	wire _w5555_ ;
	wire _w5556_ ;
	wire _w5557_ ;
	wire _w5558_ ;
	wire _w5559_ ;
	wire _w5560_ ;
	wire _w5561_ ;
	wire _w5562_ ;
	wire _w5563_ ;
	wire _w5564_ ;
	wire _w5565_ ;
	wire _w5566_ ;
	wire _w5567_ ;
	wire _w5568_ ;
	wire _w5569_ ;
	wire _w5570_ ;
	wire _w5571_ ;
	wire _w5572_ ;
	wire _w5573_ ;
	wire _w5574_ ;
	wire _w5575_ ;
	wire _w5576_ ;
	wire _w5577_ ;
	wire _w5578_ ;
	wire _w5579_ ;
	wire _w5580_ ;
	wire _w5581_ ;
	wire _w5582_ ;
	wire _w5583_ ;
	wire _w5584_ ;
	wire _w5585_ ;
	wire _w5586_ ;
	wire _w5587_ ;
	wire _w5588_ ;
	wire _w5589_ ;
	wire _w5590_ ;
	wire _w5591_ ;
	wire _w5592_ ;
	wire _w5593_ ;
	wire _w5594_ ;
	wire _w5595_ ;
	wire _w5596_ ;
	wire _w5597_ ;
	wire _w5598_ ;
	wire _w5599_ ;
	wire _w5600_ ;
	wire _w5601_ ;
	wire _w5602_ ;
	wire _w5603_ ;
	wire _w5604_ ;
	wire _w5605_ ;
	wire _w5606_ ;
	wire _w5607_ ;
	wire _w5608_ ;
	wire _w5609_ ;
	wire _w5610_ ;
	wire _w5611_ ;
	wire _w5612_ ;
	wire _w5613_ ;
	wire _w5614_ ;
	wire _w5615_ ;
	wire _w5616_ ;
	wire _w5617_ ;
	wire _w5618_ ;
	wire _w5619_ ;
	wire _w5620_ ;
	wire _w5621_ ;
	wire _w5622_ ;
	wire _w5623_ ;
	wire _w5624_ ;
	wire _w5625_ ;
	wire _w5626_ ;
	wire _w5627_ ;
	wire _w5628_ ;
	wire _w5629_ ;
	wire _w5630_ ;
	wire _w5631_ ;
	wire _w5632_ ;
	wire _w5633_ ;
	wire _w5634_ ;
	wire _w5635_ ;
	wire _w5636_ ;
	wire _w5637_ ;
	wire _w5638_ ;
	wire _w5639_ ;
	wire _w5640_ ;
	wire _w5641_ ;
	wire _w5642_ ;
	wire _w5643_ ;
	wire _w5644_ ;
	wire _w5645_ ;
	wire _w5646_ ;
	wire _w5647_ ;
	wire _w5648_ ;
	wire _w5649_ ;
	wire _w5650_ ;
	wire _w5651_ ;
	wire _w5652_ ;
	wire _w5653_ ;
	wire _w5654_ ;
	wire _w5655_ ;
	wire _w5656_ ;
	wire _w5657_ ;
	wire _w5658_ ;
	wire _w5659_ ;
	wire _w5660_ ;
	wire _w5661_ ;
	wire _w5662_ ;
	wire _w5663_ ;
	wire _w5664_ ;
	wire _w5665_ ;
	wire _w5666_ ;
	wire _w5667_ ;
	wire _w5668_ ;
	wire _w5669_ ;
	wire _w5670_ ;
	wire _w5671_ ;
	wire _w5672_ ;
	wire _w5673_ ;
	wire _w5674_ ;
	wire _w5675_ ;
	wire _w5676_ ;
	wire _w5677_ ;
	wire _w5678_ ;
	wire _w5679_ ;
	wire _w5680_ ;
	wire _w5681_ ;
	wire _w5682_ ;
	wire _w5683_ ;
	wire _w5684_ ;
	wire _w5685_ ;
	wire _w5686_ ;
	wire _w5687_ ;
	wire _w5688_ ;
	wire _w5689_ ;
	wire _w5690_ ;
	wire _w5691_ ;
	wire _w5692_ ;
	wire _w5693_ ;
	wire _w5694_ ;
	wire _w5695_ ;
	wire _w5696_ ;
	wire _w5697_ ;
	wire _w5698_ ;
	wire _w5699_ ;
	wire _w5700_ ;
	wire _w5701_ ;
	wire _w5702_ ;
	wire _w5703_ ;
	wire _w5704_ ;
	wire _w5705_ ;
	wire _w5706_ ;
	wire _w5707_ ;
	wire _w5708_ ;
	wire _w5709_ ;
	wire _w5710_ ;
	wire _w5711_ ;
	wire _w5712_ ;
	wire _w5713_ ;
	wire _w5714_ ;
	wire _w5715_ ;
	wire _w5716_ ;
	wire _w5717_ ;
	wire _w5718_ ;
	wire _w5719_ ;
	wire _w5720_ ;
	wire _w5721_ ;
	wire _w5722_ ;
	wire _w5723_ ;
	wire _w5724_ ;
	wire _w5725_ ;
	wire _w5726_ ;
	wire _w5727_ ;
	wire _w5728_ ;
	wire _w5729_ ;
	wire _w5730_ ;
	wire _w5731_ ;
	wire _w5732_ ;
	wire _w5733_ ;
	wire _w5734_ ;
	wire _w5735_ ;
	wire _w5736_ ;
	wire _w5737_ ;
	wire _w5738_ ;
	wire _w5739_ ;
	wire _w5740_ ;
	wire _w5741_ ;
	wire _w5742_ ;
	wire _w5743_ ;
	wire _w5744_ ;
	wire _w5745_ ;
	wire _w5746_ ;
	wire _w5747_ ;
	wire _w5748_ ;
	wire _w5749_ ;
	wire _w5750_ ;
	wire _w5751_ ;
	wire _w5752_ ;
	wire _w5753_ ;
	wire _w5754_ ;
	wire _w5755_ ;
	wire _w5756_ ;
	wire _w5757_ ;
	wire _w5758_ ;
	wire _w5759_ ;
	wire _w5760_ ;
	wire _w5761_ ;
	wire _w5762_ ;
	wire _w5763_ ;
	wire _w5764_ ;
	wire _w5765_ ;
	wire _w5766_ ;
	wire _w5767_ ;
	wire _w5768_ ;
	wire _w5769_ ;
	wire _w5770_ ;
	wire _w5771_ ;
	wire _w5772_ ;
	wire _w5773_ ;
	wire _w5774_ ;
	wire _w5775_ ;
	wire _w5776_ ;
	wire _w5777_ ;
	wire _w5778_ ;
	wire _w5779_ ;
	wire _w5780_ ;
	wire _w5781_ ;
	wire _w5782_ ;
	wire _w5783_ ;
	wire _w5784_ ;
	wire _w5785_ ;
	wire _w5786_ ;
	wire _w5787_ ;
	wire _w5788_ ;
	wire _w5789_ ;
	wire _w5790_ ;
	wire _w5791_ ;
	wire _w5792_ ;
	wire _w5793_ ;
	wire _w5794_ ;
	wire _w5795_ ;
	wire _w5796_ ;
	wire _w5797_ ;
	wire _w5798_ ;
	wire _w5799_ ;
	wire _w5800_ ;
	wire _w5801_ ;
	wire _w5802_ ;
	wire _w5803_ ;
	wire _w5804_ ;
	wire _w5805_ ;
	wire _w5806_ ;
	wire _w5807_ ;
	wire _w5808_ ;
	wire _w5809_ ;
	wire _w5810_ ;
	wire _w5811_ ;
	wire _w5812_ ;
	wire _w5813_ ;
	wire _w5814_ ;
	wire _w5815_ ;
	wire _w5816_ ;
	wire _w5817_ ;
	wire _w5818_ ;
	wire _w5819_ ;
	wire _w5820_ ;
	wire _w5821_ ;
	wire _w5822_ ;
	wire _w5823_ ;
	wire _w5824_ ;
	wire _w5825_ ;
	wire _w5826_ ;
	wire _w5827_ ;
	wire _w5828_ ;
	wire _w5829_ ;
	wire _w5830_ ;
	wire _w5831_ ;
	wire _w5832_ ;
	wire _w5833_ ;
	wire _w5834_ ;
	wire _w5835_ ;
	wire _w5836_ ;
	wire _w5837_ ;
	wire _w5838_ ;
	wire _w5839_ ;
	wire _w5840_ ;
	wire _w5841_ ;
	wire _w5842_ ;
	wire _w5843_ ;
	wire _w5844_ ;
	wire _w5845_ ;
	wire _w5846_ ;
	wire _w5847_ ;
	wire _w5848_ ;
	wire _w5849_ ;
	wire _w5850_ ;
	wire _w5851_ ;
	wire _w5852_ ;
	wire _w5853_ ;
	wire _w5854_ ;
	wire _w5855_ ;
	wire _w5856_ ;
	wire _w5857_ ;
	wire _w5858_ ;
	wire _w5859_ ;
	wire _w5860_ ;
	wire _w5861_ ;
	wire _w5862_ ;
	wire _w5863_ ;
	wire _w5864_ ;
	wire _w5865_ ;
	wire _w5866_ ;
	wire _w5867_ ;
	wire _w5868_ ;
	wire _w5869_ ;
	wire _w5870_ ;
	wire _w5871_ ;
	wire _w5872_ ;
	wire _w5873_ ;
	wire _w5874_ ;
	wire _w5875_ ;
	wire _w5876_ ;
	wire _w5877_ ;
	wire _w5878_ ;
	wire _w5879_ ;
	wire _w5880_ ;
	wire _w5881_ ;
	wire _w5882_ ;
	wire _w5883_ ;
	wire _w5884_ ;
	wire _w5885_ ;
	wire _w5886_ ;
	wire _w5887_ ;
	wire _w5888_ ;
	wire _w5889_ ;
	wire _w5890_ ;
	wire _w5891_ ;
	wire _w5892_ ;
	wire _w5893_ ;
	wire _w5894_ ;
	wire _w5895_ ;
	wire _w5896_ ;
	wire _w5897_ ;
	wire _w5898_ ;
	wire _w5899_ ;
	wire _w5900_ ;
	wire _w5901_ ;
	wire _w5902_ ;
	wire _w5903_ ;
	wire _w5904_ ;
	wire _w5905_ ;
	wire _w5906_ ;
	wire _w5907_ ;
	wire _w5908_ ;
	wire _w5909_ ;
	wire _w5910_ ;
	wire _w5911_ ;
	wire _w5912_ ;
	wire _w5913_ ;
	wire _w5914_ ;
	wire _w5915_ ;
	wire _w5916_ ;
	wire _w5917_ ;
	wire _w5918_ ;
	wire _w5919_ ;
	wire _w5920_ ;
	wire _w5921_ ;
	wire _w5922_ ;
	wire _w5923_ ;
	wire _w5924_ ;
	wire _w5925_ ;
	wire _w5926_ ;
	wire _w5927_ ;
	wire _w5928_ ;
	wire _w5929_ ;
	wire _w5930_ ;
	wire _w5931_ ;
	wire _w5932_ ;
	wire _w5933_ ;
	wire _w5934_ ;
	wire _w5935_ ;
	wire _w5936_ ;
	wire _w5937_ ;
	wire _w5938_ ;
	wire _w5939_ ;
	wire _w5940_ ;
	wire _w5941_ ;
	wire _w5942_ ;
	wire _w5943_ ;
	wire _w5944_ ;
	wire _w5945_ ;
	wire _w5946_ ;
	wire _w5947_ ;
	wire _w5948_ ;
	wire _w5949_ ;
	wire _w5950_ ;
	wire _w5951_ ;
	wire _w5952_ ;
	wire _w5953_ ;
	wire _w5954_ ;
	wire _w5955_ ;
	wire _w5956_ ;
	wire _w5957_ ;
	wire _w5958_ ;
	wire _w5959_ ;
	wire _w5960_ ;
	wire _w5961_ ;
	wire _w5962_ ;
	wire _w5963_ ;
	wire _w5964_ ;
	wire _w5965_ ;
	wire _w5966_ ;
	wire _w5967_ ;
	wire _w5968_ ;
	wire _w5969_ ;
	wire _w5970_ ;
	wire _w5971_ ;
	wire _w5972_ ;
	wire _w5973_ ;
	wire _w5974_ ;
	wire _w5975_ ;
	wire _w5976_ ;
	wire _w5977_ ;
	wire _w5978_ ;
	wire _w5979_ ;
	wire _w5980_ ;
	wire _w5981_ ;
	wire _w5982_ ;
	wire _w5983_ ;
	wire _w5984_ ;
	wire _w5985_ ;
	wire _w5986_ ;
	wire _w5987_ ;
	wire _w5988_ ;
	wire _w5989_ ;
	wire _w5990_ ;
	wire _w5991_ ;
	wire _w5992_ ;
	wire _w5993_ ;
	wire _w5994_ ;
	wire _w5995_ ;
	wire _w5996_ ;
	wire _w5997_ ;
	wire _w5998_ ;
	wire _w5999_ ;
	wire _w6000_ ;
	wire _w6001_ ;
	wire _w6002_ ;
	wire _w6003_ ;
	wire _w6004_ ;
	wire _w6005_ ;
	wire _w6006_ ;
	wire _w6007_ ;
	wire _w6008_ ;
	wire _w6009_ ;
	wire _w6010_ ;
	wire _w6011_ ;
	wire _w6012_ ;
	wire _w6013_ ;
	wire _w6014_ ;
	wire _w6015_ ;
	wire _w6016_ ;
	wire _w6017_ ;
	wire _w6018_ ;
	wire _w6019_ ;
	wire _w6020_ ;
	wire _w6021_ ;
	wire _w6022_ ;
	wire _w6023_ ;
	wire _w6024_ ;
	wire _w6025_ ;
	wire _w6026_ ;
	wire _w6027_ ;
	wire _w6028_ ;
	wire _w6029_ ;
	wire _w6030_ ;
	wire _w6031_ ;
	wire _w6032_ ;
	wire _w6033_ ;
	wire _w6034_ ;
	wire _w6035_ ;
	wire _w6036_ ;
	wire _w6037_ ;
	wire _w6038_ ;
	wire _w6039_ ;
	wire _w6040_ ;
	wire _w6041_ ;
	wire _w6042_ ;
	wire _w6043_ ;
	wire _w6044_ ;
	wire _w6045_ ;
	wire _w6046_ ;
	wire _w6047_ ;
	wire _w6048_ ;
	wire _w6049_ ;
	wire _w6050_ ;
	wire _w6051_ ;
	wire _w6052_ ;
	wire _w6053_ ;
	wire _w6054_ ;
	wire _w6055_ ;
	wire _w6056_ ;
	wire _w6057_ ;
	wire _w6058_ ;
	wire _w6059_ ;
	wire _w6060_ ;
	wire _w6061_ ;
	wire _w6062_ ;
	wire _w6063_ ;
	wire _w6064_ ;
	wire _w6065_ ;
	wire _w6066_ ;
	wire _w6067_ ;
	wire _w6068_ ;
	wire _w6069_ ;
	wire _w6070_ ;
	wire _w6071_ ;
	wire _w6072_ ;
	wire _w6073_ ;
	wire _w6074_ ;
	wire _w6075_ ;
	wire _w6076_ ;
	wire _w6077_ ;
	wire _w6078_ ;
	wire _w6079_ ;
	wire _w6080_ ;
	wire _w6081_ ;
	wire _w6082_ ;
	wire _w6083_ ;
	wire _w6084_ ;
	wire _w6085_ ;
	wire _w6086_ ;
	wire _w6087_ ;
	wire _w6088_ ;
	wire _w6089_ ;
	wire _w6090_ ;
	wire _w6091_ ;
	wire _w6092_ ;
	wire _w6093_ ;
	wire _w6094_ ;
	wire _w6095_ ;
	wire _w6096_ ;
	wire _w6097_ ;
	wire _w6098_ ;
	wire _w6099_ ;
	wire _w6100_ ;
	wire _w6101_ ;
	wire _w6102_ ;
	wire _w6103_ ;
	wire _w6104_ ;
	wire _w6105_ ;
	wire _w6106_ ;
	wire _w6107_ ;
	wire _w6108_ ;
	wire _w6109_ ;
	wire _w6110_ ;
	wire _w6111_ ;
	wire _w6112_ ;
	wire _w6113_ ;
	wire _w6114_ ;
	wire _w6115_ ;
	wire _w6116_ ;
	wire _w6117_ ;
	wire _w6118_ ;
	wire _w6119_ ;
	wire _w6120_ ;
	wire _w6121_ ;
	wire _w6122_ ;
	wire _w6123_ ;
	wire _w6124_ ;
	wire _w6125_ ;
	wire _w6126_ ;
	wire _w6127_ ;
	wire _w6128_ ;
	wire _w6129_ ;
	wire _w6130_ ;
	wire _w6131_ ;
	wire _w6132_ ;
	wire _w6133_ ;
	wire _w6134_ ;
	wire _w6135_ ;
	wire _w6136_ ;
	wire _w6137_ ;
	wire _w6138_ ;
	wire _w6139_ ;
	wire _w6140_ ;
	wire _w6141_ ;
	wire _w6142_ ;
	wire _w6143_ ;
	wire _w6144_ ;
	wire _w6145_ ;
	wire _w6146_ ;
	wire _w6147_ ;
	wire _w6148_ ;
	wire _w6149_ ;
	wire _w6150_ ;
	wire _w6151_ ;
	wire _w6152_ ;
	wire _w6153_ ;
	wire _w6154_ ;
	wire _w6155_ ;
	wire _w6156_ ;
	wire _w6157_ ;
	wire _w6158_ ;
	wire _w6159_ ;
	wire _w6160_ ;
	wire _w6161_ ;
	wire _w6162_ ;
	wire _w6163_ ;
	wire _w6164_ ;
	wire _w6165_ ;
	wire _w6166_ ;
	wire _w6167_ ;
	wire _w6168_ ;
	wire _w6169_ ;
	wire _w6170_ ;
	wire _w6171_ ;
	wire _w6172_ ;
	wire _w6173_ ;
	wire _w6174_ ;
	wire _w6175_ ;
	wire _w6176_ ;
	wire _w6177_ ;
	wire _w6178_ ;
	wire _w6179_ ;
	wire _w6180_ ;
	wire _w6181_ ;
	wire _w6182_ ;
	wire _w6183_ ;
	wire _w6184_ ;
	wire _w6185_ ;
	wire _w6186_ ;
	wire _w6187_ ;
	wire _w6188_ ;
	wire _w6189_ ;
	wire _w6190_ ;
	wire _w6191_ ;
	wire _w6192_ ;
	wire _w6193_ ;
	wire _w6194_ ;
	wire _w6195_ ;
	wire _w6196_ ;
	wire _w6197_ ;
	wire _w6198_ ;
	wire _w6199_ ;
	wire _w6200_ ;
	wire _w6201_ ;
	wire _w6202_ ;
	wire _w6203_ ;
	wire _w6204_ ;
	wire _w6205_ ;
	wire _w6206_ ;
	wire _w6207_ ;
	wire _w6208_ ;
	wire _w6209_ ;
	wire _w6210_ ;
	wire _w6211_ ;
	wire _w6212_ ;
	wire _w6213_ ;
	wire _w6214_ ;
	wire _w6215_ ;
	wire _w6216_ ;
	wire _w6217_ ;
	wire _w6218_ ;
	wire _w6219_ ;
	wire _w6220_ ;
	wire _w6221_ ;
	wire _w6222_ ;
	wire _w6223_ ;
	wire _w6224_ ;
	wire _w6225_ ;
	wire _w6226_ ;
	wire _w6227_ ;
	wire _w6228_ ;
	wire _w6229_ ;
	wire _w6230_ ;
	wire _w6231_ ;
	wire _w6232_ ;
	wire _w6233_ ;
	wire _w6234_ ;
	wire _w6235_ ;
	wire _w6236_ ;
	wire _w6237_ ;
	wire _w6238_ ;
	wire _w6239_ ;
	wire _w6240_ ;
	wire _w6241_ ;
	wire _w6242_ ;
	wire _w6243_ ;
	wire _w6244_ ;
	wire _w6245_ ;
	wire _w6246_ ;
	wire _w6247_ ;
	wire _w6248_ ;
	wire _w6249_ ;
	wire _w6250_ ;
	wire _w6251_ ;
	wire _w6252_ ;
	wire _w6253_ ;
	wire _w6254_ ;
	wire _w6255_ ;
	wire _w6256_ ;
	wire _w6257_ ;
	wire _w6258_ ;
	wire _w6259_ ;
	wire _w6260_ ;
	wire _w6261_ ;
	wire _w6262_ ;
	wire _w6263_ ;
	wire _w6264_ ;
	wire _w6265_ ;
	wire _w6266_ ;
	wire _w6267_ ;
	wire _w6268_ ;
	wire _w6269_ ;
	wire _w6270_ ;
	wire _w6271_ ;
	wire _w6272_ ;
	wire _w6273_ ;
	wire _w6274_ ;
	wire _w6275_ ;
	wire _w6276_ ;
	wire _w6277_ ;
	wire _w6278_ ;
	wire _w6279_ ;
	wire _w6280_ ;
	wire _w6281_ ;
	wire _w6282_ ;
	wire _w6283_ ;
	wire _w6284_ ;
	wire _w6285_ ;
	wire _w6286_ ;
	wire _w6287_ ;
	wire _w6288_ ;
	wire _w6289_ ;
	wire _w6290_ ;
	wire _w6291_ ;
	wire _w6292_ ;
	wire _w6293_ ;
	wire _w6294_ ;
	wire _w6295_ ;
	wire _w6296_ ;
	wire _w6297_ ;
	wire _w6298_ ;
	wire _w6299_ ;
	wire _w6300_ ;
	wire _w6301_ ;
	wire _w6302_ ;
	wire _w6303_ ;
	wire _w6304_ ;
	wire _w6305_ ;
	wire _w6306_ ;
	wire _w6307_ ;
	wire _w6308_ ;
	wire _w6309_ ;
	wire _w6310_ ;
	wire _w6311_ ;
	wire _w6312_ ;
	wire _w6313_ ;
	wire _w6314_ ;
	wire _w6315_ ;
	wire _w6316_ ;
	wire _w6317_ ;
	wire _w6318_ ;
	wire _w6319_ ;
	wire _w6320_ ;
	wire _w6321_ ;
	wire _w6322_ ;
	wire _w6323_ ;
	wire _w6324_ ;
	wire _w6325_ ;
	wire _w6326_ ;
	wire _w6327_ ;
	wire _w6328_ ;
	wire _w6329_ ;
	wire _w6330_ ;
	wire _w6331_ ;
	wire _w6332_ ;
	wire _w6333_ ;
	wire _w6334_ ;
	wire _w6335_ ;
	wire _w6336_ ;
	wire _w6337_ ;
	wire _w6338_ ;
	wire _w6339_ ;
	wire _w6340_ ;
	wire _w6341_ ;
	wire _w6342_ ;
	wire _w6343_ ;
	wire _w6344_ ;
	wire _w6345_ ;
	wire _w6346_ ;
	wire _w6347_ ;
	wire _w6348_ ;
	wire _w6349_ ;
	wire _w6350_ ;
	wire _w6351_ ;
	wire _w6352_ ;
	wire _w6353_ ;
	wire _w6354_ ;
	wire _w6355_ ;
	wire _w6356_ ;
	wire _w6357_ ;
	wire _w6358_ ;
	wire _w6359_ ;
	wire _w6360_ ;
	wire _w6361_ ;
	wire _w6362_ ;
	wire _w6363_ ;
	wire _w6364_ ;
	wire _w6365_ ;
	wire _w6366_ ;
	wire _w6367_ ;
	wire _w6368_ ;
	wire _w6369_ ;
	wire _w6370_ ;
	wire _w6371_ ;
	wire _w6372_ ;
	wire _w6373_ ;
	wire _w6374_ ;
	wire _w6375_ ;
	wire _w6376_ ;
	wire _w6377_ ;
	wire _w6378_ ;
	wire _w6379_ ;
	wire _w6380_ ;
	wire _w6381_ ;
	wire _w6382_ ;
	wire _w6383_ ;
	wire _w6384_ ;
	wire _w6385_ ;
	wire _w6386_ ;
	wire _w6387_ ;
	wire _w6388_ ;
	wire _w6389_ ;
	wire _w6390_ ;
	wire _w6391_ ;
	wire _w6392_ ;
	wire _w6393_ ;
	wire _w6394_ ;
	wire _w6395_ ;
	wire _w6396_ ;
	wire _w6397_ ;
	wire _w6398_ ;
	wire _w6399_ ;
	wire _w6400_ ;
	wire _w6401_ ;
	wire _w6402_ ;
	wire _w6403_ ;
	wire _w6404_ ;
	wire _w6405_ ;
	wire _w6406_ ;
	wire _w6407_ ;
	wire _w6408_ ;
	wire _w6409_ ;
	wire _w6410_ ;
	wire _w6411_ ;
	wire _w6412_ ;
	wire _w6413_ ;
	wire _w6414_ ;
	wire _w6415_ ;
	wire _w6416_ ;
	wire _w6417_ ;
	wire _w6418_ ;
	wire _w6419_ ;
	wire _w6420_ ;
	wire _w6421_ ;
	wire _w6422_ ;
	wire _w6423_ ;
	wire _w6424_ ;
	wire _w6425_ ;
	wire _w6426_ ;
	wire _w6427_ ;
	wire _w6428_ ;
	wire _w6429_ ;
	wire _w6430_ ;
	wire _w6431_ ;
	wire _w6432_ ;
	wire _w6433_ ;
	wire _w6434_ ;
	wire _w6435_ ;
	wire _w6436_ ;
	wire _w6437_ ;
	wire _w6438_ ;
	wire _w6439_ ;
	wire _w6440_ ;
	wire _w6441_ ;
	wire _w6442_ ;
	wire _w6443_ ;
	wire _w6444_ ;
	wire _w6445_ ;
	wire _w6446_ ;
	wire _w6447_ ;
	wire _w6448_ ;
	wire _w6449_ ;
	wire _w6450_ ;
	wire _w6451_ ;
	wire _w6452_ ;
	wire _w6453_ ;
	wire _w6454_ ;
	wire _w6455_ ;
	wire _w6456_ ;
	wire _w6457_ ;
	wire _w6458_ ;
	wire _w6459_ ;
	wire _w6460_ ;
	wire _w6461_ ;
	wire _w6462_ ;
	wire _w6463_ ;
	wire _w6464_ ;
	wire _w6465_ ;
	wire _w6466_ ;
	wire _w6467_ ;
	wire _w6468_ ;
	wire _w6469_ ;
	wire _w6470_ ;
	wire _w6471_ ;
	wire _w6472_ ;
	wire _w6473_ ;
	wire _w6474_ ;
	wire _w6475_ ;
	wire _w6476_ ;
	wire _w6477_ ;
	wire _w6478_ ;
	wire _w6479_ ;
	wire _w6480_ ;
	wire _w6481_ ;
	wire _w6482_ ;
	wire _w6483_ ;
	wire _w6484_ ;
	wire _w6485_ ;
	wire _w6486_ ;
	wire _w6487_ ;
	wire _w6488_ ;
	wire _w6489_ ;
	wire _w6490_ ;
	wire _w6491_ ;
	wire _w6492_ ;
	wire _w6493_ ;
	wire _w6494_ ;
	wire _w6495_ ;
	wire _w6496_ ;
	wire _w6497_ ;
	wire _w6498_ ;
	wire _w6499_ ;
	wire _w6500_ ;
	wire _w6501_ ;
	wire _w6502_ ;
	wire _w6503_ ;
	wire _w6504_ ;
	wire _w6505_ ;
	wire _w6506_ ;
	wire _w6507_ ;
	wire _w6508_ ;
	wire _w6509_ ;
	wire _w6510_ ;
	wire _w6511_ ;
	wire _w6512_ ;
	wire _w6513_ ;
	wire _w6514_ ;
	wire _w6515_ ;
	wire _w6516_ ;
	wire _w6517_ ;
	wire _w6518_ ;
	wire _w6519_ ;
	wire _w6520_ ;
	wire _w6521_ ;
	wire _w6522_ ;
	wire _w6523_ ;
	wire _w6524_ ;
	wire _w6525_ ;
	wire _w6526_ ;
	wire _w6527_ ;
	wire _w6528_ ;
	wire _w6529_ ;
	wire _w6530_ ;
	wire _w6531_ ;
	wire _w6532_ ;
	wire _w6533_ ;
	wire _w6534_ ;
	wire _w6535_ ;
	wire _w6536_ ;
	wire _w6537_ ;
	wire _w6538_ ;
	wire _w6539_ ;
	wire _w6540_ ;
	wire _w6541_ ;
	wire _w6542_ ;
	wire _w6543_ ;
	wire _w6544_ ;
	wire _w6545_ ;
	wire _w6546_ ;
	wire _w6547_ ;
	wire _w6548_ ;
	wire _w6549_ ;
	wire _w6550_ ;
	wire _w6551_ ;
	wire _w6552_ ;
	wire _w6553_ ;
	wire _w6554_ ;
	wire _w6555_ ;
	wire _w6556_ ;
	wire _w6557_ ;
	wire _w6558_ ;
	wire _w6559_ ;
	wire _w6560_ ;
	wire _w6561_ ;
	wire _w6562_ ;
	wire _w6563_ ;
	wire _w6564_ ;
	wire _w6565_ ;
	wire _w6566_ ;
	wire _w6567_ ;
	wire _w6568_ ;
	wire _w6569_ ;
	wire _w6570_ ;
	wire _w6571_ ;
	wire _w6572_ ;
	wire _w6573_ ;
	wire _w6574_ ;
	wire _w6575_ ;
	wire _w6576_ ;
	wire _w6577_ ;
	wire _w6578_ ;
	wire _w6579_ ;
	wire _w6580_ ;
	wire _w6581_ ;
	wire _w6582_ ;
	wire _w6583_ ;
	wire _w6584_ ;
	wire _w6585_ ;
	wire _w6586_ ;
	wire _w6587_ ;
	wire _w6588_ ;
	wire _w6589_ ;
	wire _w6590_ ;
	wire _w6591_ ;
	wire _w6592_ ;
	wire _w6593_ ;
	wire _w6594_ ;
	wire _w6595_ ;
	wire _w6596_ ;
	wire _w6597_ ;
	wire _w6598_ ;
	wire _w6599_ ;
	wire _w6600_ ;
	wire _w6601_ ;
	wire _w6602_ ;
	wire _w6603_ ;
	wire _w6604_ ;
	wire _w6605_ ;
	wire _w6606_ ;
	wire _w6607_ ;
	wire _w6608_ ;
	wire _w6609_ ;
	wire _w6610_ ;
	wire _w6611_ ;
	wire _w6612_ ;
	wire _w6613_ ;
	wire _w6614_ ;
	wire _w6615_ ;
	wire _w6616_ ;
	wire _w6617_ ;
	wire _w6618_ ;
	wire _w6619_ ;
	wire _w6620_ ;
	wire _w6621_ ;
	wire _w6622_ ;
	wire _w6623_ ;
	wire _w6624_ ;
	wire _w6625_ ;
	wire _w6626_ ;
	wire _w6627_ ;
	wire _w6628_ ;
	wire _w6629_ ;
	wire _w6630_ ;
	wire _w6631_ ;
	wire _w6632_ ;
	wire _w6633_ ;
	wire _w6634_ ;
	wire _w6635_ ;
	wire _w6636_ ;
	wire _w6637_ ;
	wire _w6638_ ;
	wire _w6639_ ;
	wire _w6640_ ;
	wire _w6641_ ;
	wire _w6642_ ;
	wire _w6643_ ;
	wire _w6644_ ;
	wire _w6645_ ;
	wire _w6646_ ;
	wire _w6647_ ;
	wire _w6648_ ;
	wire _w6649_ ;
	wire _w6650_ ;
	wire _w6651_ ;
	wire _w6652_ ;
	wire _w6653_ ;
	wire _w6654_ ;
	wire _w6655_ ;
	wire _w6656_ ;
	wire _w6657_ ;
	wire _w6658_ ;
	wire _w6659_ ;
	wire _w6660_ ;
	wire _w6661_ ;
	wire _w6662_ ;
	wire _w6663_ ;
	wire _w6664_ ;
	wire _w6665_ ;
	wire _w6666_ ;
	wire _w6667_ ;
	wire _w6668_ ;
	wire _w6669_ ;
	wire _w6670_ ;
	wire _w6671_ ;
	wire _w6672_ ;
	wire _w6673_ ;
	wire _w6674_ ;
	wire _w6675_ ;
	wire _w6676_ ;
	wire _w6677_ ;
	wire _w6678_ ;
	wire _w6679_ ;
	wire _w6680_ ;
	wire _w6681_ ;
	wire _w6682_ ;
	wire _w6683_ ;
	wire _w6684_ ;
	wire _w6685_ ;
	wire _w6686_ ;
	wire _w6687_ ;
	wire _w6688_ ;
	wire _w6689_ ;
	wire _w6690_ ;
	wire _w6691_ ;
	wire _w6692_ ;
	wire _w6693_ ;
	wire _w6694_ ;
	wire _w6695_ ;
	wire _w6696_ ;
	wire _w6697_ ;
	wire _w6698_ ;
	wire _w6699_ ;
	wire _w6700_ ;
	wire _w6701_ ;
	wire _w6702_ ;
	wire _w6703_ ;
	wire _w6704_ ;
	wire _w6705_ ;
	wire _w6706_ ;
	wire _w6707_ ;
	wire _w6708_ ;
	wire _w6709_ ;
	wire _w6710_ ;
	wire _w6711_ ;
	wire _w6712_ ;
	wire _w6713_ ;
	wire _w6714_ ;
	wire _w6715_ ;
	wire _w6716_ ;
	wire _w6717_ ;
	wire _w6718_ ;
	wire _w6719_ ;
	wire _w6720_ ;
	wire _w6721_ ;
	wire _w6722_ ;
	wire _w6723_ ;
	wire _w6724_ ;
	wire _w6725_ ;
	wire _w6726_ ;
	wire _w6727_ ;
	wire _w6728_ ;
	wire _w6729_ ;
	wire _w6730_ ;
	wire _w6731_ ;
	wire _w6732_ ;
	wire _w6733_ ;
	wire _w6734_ ;
	wire _w6735_ ;
	wire _w6736_ ;
	wire _w6737_ ;
	wire _w6738_ ;
	wire _w6739_ ;
	wire _w6740_ ;
	wire _w6741_ ;
	wire _w6742_ ;
	wire _w6743_ ;
	wire _w6744_ ;
	wire _w6745_ ;
	wire _w6746_ ;
	wire _w6747_ ;
	wire _w6748_ ;
	wire _w6749_ ;
	wire _w6750_ ;
	wire _w6751_ ;
	wire _w6752_ ;
	wire _w6753_ ;
	wire _w6754_ ;
	wire _w6755_ ;
	wire _w6756_ ;
	wire _w6757_ ;
	wire _w6758_ ;
	wire _w6759_ ;
	wire _w6760_ ;
	wire _w6761_ ;
	wire _w6762_ ;
	wire _w6763_ ;
	wire _w6764_ ;
	wire _w6765_ ;
	wire _w6766_ ;
	wire _w6767_ ;
	wire _w6768_ ;
	wire _w6769_ ;
	wire _w6770_ ;
	wire _w6771_ ;
	wire _w6772_ ;
	wire _w6773_ ;
	wire _w6774_ ;
	wire _w6775_ ;
	wire _w6776_ ;
	wire _w6777_ ;
	wire _w6778_ ;
	wire _w6779_ ;
	wire _w6780_ ;
	wire _w6781_ ;
	wire _w6782_ ;
	wire _w6783_ ;
	wire _w6784_ ;
	wire _w6785_ ;
	wire _w6786_ ;
	wire _w6787_ ;
	wire _w6788_ ;
	wire _w6789_ ;
	wire _w6790_ ;
	wire _w6791_ ;
	wire _w6792_ ;
	wire _w6793_ ;
	wire _w6794_ ;
	wire _w6795_ ;
	wire _w6796_ ;
	wire _w6797_ ;
	wire _w6798_ ;
	wire _w6799_ ;
	wire _w6800_ ;
	wire _w6801_ ;
	wire _w6802_ ;
	wire _w6803_ ;
	wire _w6804_ ;
	wire _w6805_ ;
	wire _w6806_ ;
	wire _w6807_ ;
	wire _w6808_ ;
	wire _w6809_ ;
	wire _w6810_ ;
	wire _w6811_ ;
	wire _w6812_ ;
	wire _w6813_ ;
	wire _w6814_ ;
	wire _w6815_ ;
	wire _w6816_ ;
	wire _w6817_ ;
	wire _w6818_ ;
	wire _w6819_ ;
	wire _w6820_ ;
	wire _w6821_ ;
	wire _w6822_ ;
	wire _w6823_ ;
	wire _w6824_ ;
	wire _w6825_ ;
	wire _w6826_ ;
	wire _w6827_ ;
	wire _w6828_ ;
	wire _w6829_ ;
	wire _w6830_ ;
	wire _w6831_ ;
	wire _w6832_ ;
	wire _w6833_ ;
	wire _w6834_ ;
	wire _w6835_ ;
	wire _w6836_ ;
	wire _w6837_ ;
	wire _w6838_ ;
	wire _w6839_ ;
	wire _w6840_ ;
	wire _w6841_ ;
	wire _w6842_ ;
	wire _w6843_ ;
	wire _w6844_ ;
	wire _w6845_ ;
	wire _w6846_ ;
	wire _w6847_ ;
	wire _w6848_ ;
	wire _w6849_ ;
	wire _w6850_ ;
	wire _w6851_ ;
	wire _w6852_ ;
	wire _w6853_ ;
	wire _w6854_ ;
	wire _w6855_ ;
	wire _w6856_ ;
	wire _w6857_ ;
	wire _w6858_ ;
	wire _w6859_ ;
	wire _w6860_ ;
	wire _w6861_ ;
	wire _w6862_ ;
	wire _w6863_ ;
	wire _w6864_ ;
	wire _w6865_ ;
	wire _w6866_ ;
	wire _w6867_ ;
	wire _w6868_ ;
	wire _w6869_ ;
	wire _w6870_ ;
	wire _w6871_ ;
	wire _w6872_ ;
	wire _w6873_ ;
	wire _w6874_ ;
	wire _w6875_ ;
	wire _w6876_ ;
	wire _w6877_ ;
	wire _w6878_ ;
	wire _w6879_ ;
	wire _w6880_ ;
	wire _w6881_ ;
	wire _w6882_ ;
	wire _w6883_ ;
	wire _w6884_ ;
	wire _w6885_ ;
	wire _w6886_ ;
	wire _w6887_ ;
	wire _w6888_ ;
	wire _w6889_ ;
	wire _w6890_ ;
	wire _w6891_ ;
	wire _w6892_ ;
	wire _w6893_ ;
	wire _w6894_ ;
	wire _w6895_ ;
	wire _w6896_ ;
	wire _w6897_ ;
	wire _w6898_ ;
	wire _w6899_ ;
	wire _w6900_ ;
	wire _w6901_ ;
	wire _w6902_ ;
	wire _w6903_ ;
	wire _w6904_ ;
	wire _w6905_ ;
	wire _w6906_ ;
	wire _w6907_ ;
	wire _w6908_ ;
	wire _w6909_ ;
	wire _w6910_ ;
	wire _w6911_ ;
	wire _w6912_ ;
	wire _w6913_ ;
	wire _w6914_ ;
	wire _w6915_ ;
	wire _w6916_ ;
	wire _w6917_ ;
	wire _w6918_ ;
	wire _w6919_ ;
	wire _w6920_ ;
	wire _w6921_ ;
	wire _w6922_ ;
	wire _w6923_ ;
	wire _w6924_ ;
	wire _w6925_ ;
	wire _w6926_ ;
	wire _w6927_ ;
	wire _w6928_ ;
	wire _w6929_ ;
	wire _w6930_ ;
	wire _w6931_ ;
	wire _w6932_ ;
	wire _w6933_ ;
	wire _w6934_ ;
	wire _w6935_ ;
	wire _w6936_ ;
	wire _w6937_ ;
	wire _w6938_ ;
	wire _w6939_ ;
	wire _w6940_ ;
	wire _w6941_ ;
	wire _w6942_ ;
	wire _w6943_ ;
	wire _w6944_ ;
	wire _w6945_ ;
	wire _w6946_ ;
	wire _w6947_ ;
	wire _w6948_ ;
	wire _w6949_ ;
	wire _w6950_ ;
	wire _w6951_ ;
	wire _w6952_ ;
	wire _w6953_ ;
	wire _w6954_ ;
	wire _w6955_ ;
	wire _w6956_ ;
	wire _w6957_ ;
	wire _w6958_ ;
	wire _w6959_ ;
	wire _w6960_ ;
	wire _w6961_ ;
	wire _w6962_ ;
	wire _w6963_ ;
	wire _w6964_ ;
	wire _w6965_ ;
	wire _w6966_ ;
	wire _w6967_ ;
	wire _w6968_ ;
	wire _w6969_ ;
	wire _w6970_ ;
	wire _w6971_ ;
	wire _w6972_ ;
	wire _w6973_ ;
	wire _w6974_ ;
	wire _w6975_ ;
	wire _w6976_ ;
	wire _w6977_ ;
	wire _w6978_ ;
	wire _w6979_ ;
	wire _w6980_ ;
	wire _w6981_ ;
	wire _w6982_ ;
	wire _w6983_ ;
	wire _w6984_ ;
	wire _w6985_ ;
	wire _w6986_ ;
	wire _w6987_ ;
	wire _w12174_ ;
	wire _w12175_ ;
	wire _w12176_ ;
	wire _w12177_ ;
	wire _w12178_ ;
	wire _w12179_ ;
	wire _w12180_ ;
	wire _w12181_ ;
	wire _w12182_ ;
	wire _w12183_ ;
	wire _w12184_ ;
	wire _w12185_ ;
	wire _w12186_ ;
	wire _w12187_ ;
	wire _w12188_ ;
	wire _w12189_ ;
	wire _w12190_ ;
	wire _w12191_ ;
	wire _w12192_ ;
	wire _w12193_ ;
	wire _w12194_ ;
	wire _w12195_ ;
	wire _w12196_ ;
	wire _w12197_ ;
	wire _w12198_ ;
	wire _w12199_ ;
	wire _w12200_ ;
	wire _w12201_ ;
	wire _w12202_ ;
	wire _w12203_ ;
	wire _w12204_ ;
	wire _w12205_ ;
	wire _w12206_ ;
	wire _w12207_ ;
	wire _w12208_ ;
	wire _w12209_ ;
	wire _w12210_ ;
	wire _w12211_ ;
	wire _w12212_ ;
	wire _w12213_ ;
	wire _w12214_ ;
	wire _w12215_ ;
	wire _w12216_ ;
	wire _w12217_ ;
	wire _w12218_ ;
	wire _w12219_ ;
	wire _w12220_ ;
	wire _w12221_ ;
	wire _w12222_ ;
	wire _w12223_ ;
	wire _w12224_ ;
	wire _w12225_ ;
	wire _w12226_ ;
	wire _w12227_ ;
	wire _w12228_ ;
	wire _w12229_ ;
	wire _w12230_ ;
	wire _w12231_ ;
	wire _w12232_ ;
	wire _w12233_ ;
	wire _w12234_ ;
	wire _w12235_ ;
	wire _w12236_ ;
	wire _w12237_ ;
	wire _w12238_ ;
	wire _w12239_ ;
	wire _w12240_ ;
	wire _w12241_ ;
	wire _w12242_ ;
	wire _w12243_ ;
	wire _w12244_ ;
	wire _w12245_ ;
	wire _w12246_ ;
	wire _w12247_ ;
	wire _w12248_ ;
	wire _w12249_ ;
	wire _w12250_ ;
	wire _w12251_ ;
	wire _w12252_ ;
	wire _w12253_ ;
	wire _w12254_ ;
	wire _w12255_ ;
	wire _w12256_ ;
	wire _w12257_ ;
	wire _w12258_ ;
	wire _w12259_ ;
	wire _w12260_ ;
	wire _w12261_ ;
	wire _w12262_ ;
	wire _w12263_ ;
	wire _w12264_ ;
	wire _w12265_ ;
	wire _w12266_ ;
	wire _w12267_ ;
	wire _w12268_ ;
	wire _w12269_ ;
	wire _w12270_ ;
	wire _w12271_ ;
	wire _w12272_ ;
	wire _w12273_ ;
	wire _w12274_ ;
	wire _w12275_ ;
	wire _w12276_ ;
	wire _w12277_ ;
	wire _w12278_ ;
	wire _w12279_ ;
	wire _w12280_ ;
	wire _w12281_ ;
	wire _w12282_ ;
	wire _w12283_ ;
	wire _w12284_ ;
	wire _w12285_ ;
	wire _w12286_ ;
	wire _w12287_ ;
	wire _w12288_ ;
	wire _w12289_ ;
	wire _w12290_ ;
	wire _w12291_ ;
	wire _w12292_ ;
	wire _w12293_ ;
	wire _w12294_ ;
	wire _w12295_ ;
	wire _w12296_ ;
	wire _w12297_ ;
	wire _w12298_ ;
	wire _w12299_ ;
	wire _w12300_ ;
	wire _w12301_ ;
	wire _w12302_ ;
	wire _w12303_ ;
	wire _w12304_ ;
	wire _w12305_ ;
	wire _w12306_ ;
	wire _w12307_ ;
	wire _w12308_ ;
	wire _w12309_ ;
	wire _w12310_ ;
	wire _w12311_ ;
	wire _w12312_ ;
	wire _w12313_ ;
	wire _w12314_ ;
	wire _w12315_ ;
	wire _w12316_ ;
	wire _w12317_ ;
	wire _w12318_ ;
	wire _w12319_ ;
	wire _w12320_ ;
	wire _w12321_ ;
	wire _w12322_ ;
	wire _w12323_ ;
	wire _w12324_ ;
	wire _w12325_ ;
	wire _w12326_ ;
	wire _w12327_ ;
	wire _w12328_ ;
	wire _w12329_ ;
	wire _w12330_ ;
	wire _w12331_ ;
	wire _w12332_ ;
	wire _w12333_ ;
	wire _w12334_ ;
	wire _w12335_ ;
	wire _w12336_ ;
	wire _w12337_ ;
	wire _w12338_ ;
	wire _w12339_ ;
	wire _w12340_ ;
	wire _w12341_ ;
	wire _w12342_ ;
	wire _w12343_ ;
	wire _w12344_ ;
	wire _w12345_ ;
	wire _w12346_ ;
	wire _w12347_ ;
	wire _w12348_ ;
	wire _w12349_ ;
	wire _w12350_ ;
	wire _w12351_ ;
	wire _w12352_ ;
	wire _w12353_ ;
	wire _w12354_ ;
	wire _w12355_ ;
	wire _w12356_ ;
	wire _w12357_ ;
	wire _w12358_ ;
	wire _w12359_ ;
	wire _w12360_ ;
	wire _w12361_ ;
	wire _w12362_ ;
	wire _w12363_ ;
	wire _w12364_ ;
	wire _w12365_ ;
	wire _w12366_ ;
	wire _w12367_ ;
	wire _w12368_ ;
	wire _w12369_ ;
	wire _w12370_ ;
	wire _w12371_ ;
	wire _w12372_ ;
	wire _w12373_ ;
	wire _w12374_ ;
	wire _w12375_ ;
	wire _w12376_ ;
	wire _w12377_ ;
	wire _w12378_ ;
	wire _w12379_ ;
	wire _w12380_ ;
	wire _w12381_ ;
	wire _w12382_ ;
	wire _w12383_ ;
	wire _w12384_ ;
	wire _w12385_ ;
	wire _w12386_ ;
	wire _w12387_ ;
	wire _w12388_ ;
	wire _w12389_ ;
	wire _w12390_ ;
	wire _w12391_ ;
	wire _w12392_ ;
	wire _w12393_ ;
	wire _w12394_ ;
	wire _w12395_ ;
	wire _w12396_ ;
	wire _w12397_ ;
	wire _w12398_ ;
	wire _w12399_ ;
	wire _w12400_ ;
	wire _w12401_ ;
	wire _w12402_ ;
	wire _w12403_ ;
	wire _w12404_ ;
	wire _w12405_ ;
	wire _w12406_ ;
	wire _w12407_ ;
	wire _w12408_ ;
	wire _w12409_ ;
	wire _w12410_ ;
	wire _w12411_ ;
	wire _w12412_ ;
	wire _w12413_ ;
	wire _w12414_ ;
	wire _w12415_ ;
	wire _w12416_ ;
	wire _w12417_ ;
	wire _w12418_ ;
	wire _w12419_ ;
	wire _w12420_ ;
	wire _w12421_ ;
	wire _w12422_ ;
	wire _w12423_ ;
	wire _w12424_ ;
	wire _w12425_ ;
	wire _w12426_ ;
	wire _w12427_ ;
	wire _w12428_ ;
	wire _w12429_ ;
	wire _w12430_ ;
	wire _w12431_ ;
	wire _w12432_ ;
	wire _w12433_ ;
	wire _w12434_ ;
	wire _w12435_ ;
	wire _w12436_ ;
	wire _w12437_ ;
	wire _w12438_ ;
	wire _w12439_ ;
	wire _w12440_ ;
	wire _w12441_ ;
	wire _w12442_ ;
	wire _w12443_ ;
	wire _w12444_ ;
	wire _w12445_ ;
	wire _w12446_ ;
	wire _w12447_ ;
	wire _w12448_ ;
	wire _w12449_ ;
	wire _w12450_ ;
	wire _w12451_ ;
	wire _w12452_ ;
	wire _w12453_ ;
	wire _w12454_ ;
	wire _w12455_ ;
	wire _w12456_ ;
	wire _w12457_ ;
	wire _w12458_ ;
	wire _w12459_ ;
	wire _w12460_ ;
	wire _w12461_ ;
	wire _w12462_ ;
	wire _w12463_ ;
	wire _w12464_ ;
	wire _w12465_ ;
	wire _w12466_ ;
	wire _w12467_ ;
	wire _w12468_ ;
	wire _w12469_ ;
	wire _w12470_ ;
	wire _w12471_ ;
	wire _w12472_ ;
	wire _w12473_ ;
	wire _w12474_ ;
	wire _w12475_ ;
	wire _w12476_ ;
	wire _w12477_ ;
	wire _w12478_ ;
	wire _w12479_ ;
	wire _w12480_ ;
	wire _w12481_ ;
	wire _w12482_ ;
	wire _w12483_ ;
	wire _w12484_ ;
	wire _w12485_ ;
	wire _w12486_ ;
	wire _w12487_ ;
	wire _w12488_ ;
	wire _w12489_ ;
	wire _w12490_ ;
	wire _w12491_ ;
	wire _w12492_ ;
	wire _w12493_ ;
	wire _w12494_ ;
	wire _w12495_ ;
	wire _w12496_ ;
	wire _w12497_ ;
	wire _w12498_ ;
	wire _w12499_ ;
	wire _w12500_ ;
	wire _w12501_ ;
	wire _w12502_ ;
	wire _w12503_ ;
	wire _w12504_ ;
	wire _w12505_ ;
	wire _w12506_ ;
	wire _w12507_ ;
	wire _w12508_ ;
	wire _w12509_ ;
	wire _w12510_ ;
	wire _w12511_ ;
	wire _w12512_ ;
	wire _w12513_ ;
	wire _w12514_ ;
	wire _w12515_ ;
	wire _w12516_ ;
	wire _w12517_ ;
	wire _w12518_ ;
	wire _w12519_ ;
	wire _w12520_ ;
	wire _w12521_ ;
	wire _w12522_ ;
	wire _w12523_ ;
	wire _w12524_ ;
	wire _w12525_ ;
	wire _w12526_ ;
	wire _w12527_ ;
	wire _w12528_ ;
	wire _w12529_ ;
	wire _w12530_ ;
	wire _w12531_ ;
	wire _w12532_ ;
	wire _w12533_ ;
	wire _w12534_ ;
	wire _w12535_ ;
	wire _w12536_ ;
	wire _w12537_ ;
	wire _w12538_ ;
	wire _w12539_ ;
	wire _w12540_ ;
	wire _w12541_ ;
	wire _w12542_ ;
	wire _w12543_ ;
	wire _w12544_ ;
	wire _w12545_ ;
	wire _w12546_ ;
	wire _w12547_ ;
	wire _w12548_ ;
	wire _w12549_ ;
	wire _w12550_ ;
	wire _w12551_ ;
	wire _w12552_ ;
	wire _w12553_ ;
	wire _w12554_ ;
	wire _w12555_ ;
	wire _w12556_ ;
	wire _w12557_ ;
	wire _w12558_ ;
	wire _w12559_ ;
	wire _w12560_ ;
	wire _w12561_ ;
	wire _w12562_ ;
	wire _w12563_ ;
	wire _w12564_ ;
	wire _w12565_ ;
	wire _w12566_ ;
	wire _w12567_ ;
	wire _w12568_ ;
	wire _w12569_ ;
	wire _w12570_ ;
	wire _w12571_ ;
	wire _w12572_ ;
	wire _w12573_ ;
	wire _w12574_ ;
	wire _w12575_ ;
	wire _w12576_ ;
	wire _w12577_ ;
	wire _w12578_ ;
	wire _w12579_ ;
	wire _w12580_ ;
	wire _w12581_ ;
	wire _w12582_ ;
	wire _w12583_ ;
	wire _w12584_ ;
	wire _w12585_ ;
	wire _w12586_ ;
	wire _w12587_ ;
	wire _w12588_ ;
	wire _w12589_ ;
	wire _w12590_ ;
	wire _w12591_ ;
	wire _w12592_ ;
	wire _w12593_ ;
	wire _w12594_ ;
	wire _w12595_ ;
	wire _w12596_ ;
	wire _w12597_ ;
	wire _w12598_ ;
	wire _w12599_ ;
	wire _w12600_ ;
	wire _w12601_ ;
	wire _w12602_ ;
	wire _w12603_ ;
	wire _w12604_ ;
	wire _w12605_ ;
	wire _w12606_ ;
	wire _w12607_ ;
	wire _w12608_ ;
	wire _w12609_ ;
	wire _w12610_ ;
	wire _w12611_ ;
	wire _w12612_ ;
	wire _w12613_ ;
	wire _w12614_ ;
	wire _w12615_ ;
	wire _w12616_ ;
	wire _w12617_ ;
	wire _w12618_ ;
	wire _w12619_ ;
	wire _w12620_ ;
	wire _w12621_ ;
	wire _w12622_ ;
	wire _w12623_ ;
	wire _w12624_ ;
	wire _w12625_ ;
	wire _w12626_ ;
	wire _w12627_ ;
	wire _w12628_ ;
	wire _w12629_ ;
	wire _w12630_ ;
	wire _w12631_ ;
	wire _w12632_ ;
	wire _w12633_ ;
	wire _w12634_ ;
	wire _w12635_ ;
	wire _w12636_ ;
	wire _w12637_ ;
	wire _w12638_ ;
	wire _w12639_ ;
	wire _w12640_ ;
	wire _w12641_ ;
	wire _w12642_ ;
	wire _w12643_ ;
	wire _w12644_ ;
	wire _w12645_ ;
	wire _w12646_ ;
	wire _w12647_ ;
	wire _w12648_ ;
	wire _w12649_ ;
	wire _w12650_ ;
	wire _w12651_ ;
	wire _w12652_ ;
	wire _w12653_ ;
	wire _w12654_ ;
	wire _w12655_ ;
	wire _w12656_ ;
	wire _w12657_ ;
	wire _w12658_ ;
	wire _w12659_ ;
	wire _w12660_ ;
	wire _w12661_ ;
	wire _w12662_ ;
	wire _w12663_ ;
	wire _w12664_ ;
	wire _w12665_ ;
	wire _w12666_ ;
	wire _w12667_ ;
	wire _w12668_ ;
	wire _w12669_ ;
	wire _w12670_ ;
	wire _w12671_ ;
	wire _w12672_ ;
	wire _w12673_ ;
	wire _w12674_ ;
	wire _w12675_ ;
	wire _w12676_ ;
	wire _w12677_ ;
	wire _w12678_ ;
	wire _w12679_ ;
	wire _w12680_ ;
	wire _w12681_ ;
	wire _w12682_ ;
	wire _w12683_ ;
	wire _w12684_ ;
	wire _w12685_ ;
	wire _w12686_ ;
	wire _w12687_ ;
	wire _w12688_ ;
	wire _w12689_ ;
	wire _w12690_ ;
	wire _w12691_ ;
	wire _w12692_ ;
	wire _w12693_ ;
	wire _w12694_ ;
	wire _w12695_ ;
	wire _w12696_ ;
	wire _w12697_ ;
	wire _w12698_ ;
	wire _w12699_ ;
	wire _w12700_ ;
	wire _w12701_ ;
	wire _w12702_ ;
	wire _w12703_ ;
	wire _w12704_ ;
	wire _w12705_ ;
	wire _w12706_ ;
	wire _w12707_ ;
	wire _w12708_ ;
	wire _w12709_ ;
	wire _w12710_ ;
	wire _w12711_ ;
	wire _w12712_ ;
	wire _w12713_ ;
	wire _w12714_ ;
	wire _w12715_ ;
	wire _w12716_ ;
	wire _w12717_ ;
	wire _w12718_ ;
	wire _w12719_ ;
	wire _w12720_ ;
	wire _w12721_ ;
	wire _w12722_ ;
	wire _w12723_ ;
	wire _w12724_ ;
	wire _w12725_ ;
	wire _w12726_ ;
	wire _w12727_ ;
	wire _w12728_ ;
	wire _w12729_ ;
	wire _w12730_ ;
	wire _w12731_ ;
	wire _w12732_ ;
	wire _w12733_ ;
	wire _w12734_ ;
	wire _w12735_ ;
	wire _w12736_ ;
	wire _w12737_ ;
	wire _w12738_ ;
	wire _w12739_ ;
	wire _w12740_ ;
	wire _w12741_ ;
	wire _w12742_ ;
	wire _w12743_ ;
	wire _w12744_ ;
	wire _w12745_ ;
	wire _w12746_ ;
	wire _w12747_ ;
	wire _w12748_ ;
	wire _w12749_ ;
	wire _w12750_ ;
	wire _w12751_ ;
	wire _w12752_ ;
	wire _w12753_ ;
	wire _w12754_ ;
	wire _w12755_ ;
	wire _w12756_ ;
	wire _w12757_ ;
	wire _w12758_ ;
	wire _w12759_ ;
	wire _w12760_ ;
	wire _w12761_ ;
	wire _w12762_ ;
	wire _w12763_ ;
	wire _w12764_ ;
	wire _w12765_ ;
	wire _w12766_ ;
	wire _w12767_ ;
	wire _w12768_ ;
	wire _w12769_ ;
	wire _w12770_ ;
	wire _w12771_ ;
	wire _w12772_ ;
	wire _w12773_ ;
	wire _w12774_ ;
	wire _w12775_ ;
	wire _w12776_ ;
	wire _w12777_ ;
	wire _w12778_ ;
	wire _w12779_ ;
	wire _w12780_ ;
	wire _w12781_ ;
	wire _w12782_ ;
	wire _w12783_ ;
	wire _w12784_ ;
	wire _w12785_ ;
	wire _w12786_ ;
	wire _w12787_ ;
	wire _w12788_ ;
	wire _w12789_ ;
	wire _w12790_ ;
	wire _w12791_ ;
	wire _w12792_ ;
	wire _w12793_ ;
	wire _w12794_ ;
	wire _w12795_ ;
	wire _w12796_ ;
	wire _w12797_ ;
	wire _w12798_ ;
	wire _w12799_ ;
	wire _w12800_ ;
	wire _w12801_ ;
	wire _w12802_ ;
	wire _w12803_ ;
	wire _w12804_ ;
	wire _w12805_ ;
	wire _w12806_ ;
	wire _w12807_ ;
	wire _w12808_ ;
	wire _w12809_ ;
	wire _w12810_ ;
	wire _w12811_ ;
	wire _w12812_ ;
	wire _w12813_ ;
	wire _w12814_ ;
	wire _w12815_ ;
	wire _w12816_ ;
	wire _w12817_ ;
	wire _w12818_ ;
	wire _w12819_ ;
	wire _w12820_ ;
	wire _w12821_ ;
	wire _w12822_ ;
	wire _w12823_ ;
	wire _w12824_ ;
	wire _w12825_ ;
	wire _w12826_ ;
	wire _w12827_ ;
	wire _w12828_ ;
	wire _w12829_ ;
	wire _w12830_ ;
	wire _w12831_ ;
	wire _w12832_ ;
	wire _w12833_ ;
	wire _w12834_ ;
	wire _w12835_ ;
	wire _w12836_ ;
	wire _w12837_ ;
	wire _w12838_ ;
	wire _w12839_ ;
	wire _w12840_ ;
	wire _w12841_ ;
	wire _w12842_ ;
	wire _w12843_ ;
	wire _w12844_ ;
	wire _w12845_ ;
	wire _w12846_ ;
	wire _w12847_ ;
	wire _w12848_ ;
	wire _w12849_ ;
	wire _w12850_ ;
	wire _w12851_ ;
	wire _w12852_ ;
	wire _w12853_ ;
	wire _w12854_ ;
	wire _w12855_ ;
	wire _w12856_ ;
	wire _w12857_ ;
	wire _w12858_ ;
	wire _w12859_ ;
	wire _w12860_ ;
	wire _w12861_ ;
	wire _w12862_ ;
	wire _w12863_ ;
	wire _w12864_ ;
	wire _w12865_ ;
	wire _w12866_ ;
	wire _w12867_ ;
	wire _w12868_ ;
	wire _w12869_ ;
	wire _w12870_ ;
	wire _w12871_ ;
	wire _w12872_ ;
	wire _w12873_ ;
	wire _w12874_ ;
	wire _w12875_ ;
	wire _w12876_ ;
	wire _w12877_ ;
	wire _w12878_ ;
	wire _w12879_ ;
	wire _w12880_ ;
	wire _w12881_ ;
	wire _w12882_ ;
	wire _w12883_ ;
	wire _w12884_ ;
	wire _w12885_ ;
	wire _w12886_ ;
	wire _w12887_ ;
	wire _w12888_ ;
	wire _w12889_ ;
	wire _w12890_ ;
	wire _w12891_ ;
	wire _w12892_ ;
	wire _w12893_ ;
	wire _w12894_ ;
	wire _w12895_ ;
	wire _w12896_ ;
	wire _w12897_ ;
	wire _w12898_ ;
	wire _w12899_ ;
	wire _w12900_ ;
	wire _w12901_ ;
	wire _w12902_ ;
	wire _w12903_ ;
	wire _w12904_ ;
	wire _w12905_ ;
	wire _w12906_ ;
	wire _w12907_ ;
	wire _w12908_ ;
	wire _w12909_ ;
	wire _w12910_ ;
	wire _w12911_ ;
	wire _w12912_ ;
	wire _w12913_ ;
	wire _w12914_ ;
	wire _w12915_ ;
	wire _w12916_ ;
	wire _w12917_ ;
	wire _w12918_ ;
	wire _w12919_ ;
	wire _w12920_ ;
	wire _w12921_ ;
	wire _w12922_ ;
	wire _w12923_ ;
	wire _w12924_ ;
	wire _w12925_ ;
	wire _w12926_ ;
	wire _w12927_ ;
	wire _w12928_ ;
	wire _w12929_ ;
	wire _w12930_ ;
	wire _w12931_ ;
	wire _w12932_ ;
	wire _w12933_ ;
	wire _w12934_ ;
	wire _w12935_ ;
	wire _w12936_ ;
	wire _w12937_ ;
	wire _w12938_ ;
	wire _w12939_ ;
	wire _w12940_ ;
	wire _w12941_ ;
	wire _w12942_ ;
	wire _w12943_ ;
	wire _w12944_ ;
	wire _w12945_ ;
	wire _w12946_ ;
	wire _w12947_ ;
	wire _w12948_ ;
	wire _w12949_ ;
	wire _w12950_ ;
	wire _w12951_ ;
	wire _w12952_ ;
	wire _w12953_ ;
	wire _w12954_ ;
	wire _w12955_ ;
	wire _w12956_ ;
	wire _w12957_ ;
	wire _w12958_ ;
	wire _w12959_ ;
	wire _w12960_ ;
	wire _w12961_ ;
	wire _w12962_ ;
	wire _w12963_ ;
	wire _w12964_ ;
	wire _w12965_ ;
	wire _w12966_ ;
	wire _w12967_ ;
	wire _w12968_ ;
	wire _w12969_ ;
	wire _w12970_ ;
	wire _w12971_ ;
	wire _w12972_ ;
	wire _w12973_ ;
	wire _w12974_ ;
	wire _w12975_ ;
	wire _w12976_ ;
	wire _w12977_ ;
	wire _w12978_ ;
	wire _w12979_ ;
	wire _w12980_ ;
	wire _w12981_ ;
	wire _w12982_ ;
	wire _w12983_ ;
	wire _w12984_ ;
	wire _w12985_ ;
	wire _w12986_ ;
	wire _w12987_ ;
	wire _w12988_ ;
	wire _w12989_ ;
	wire _w12990_ ;
	wire _w12991_ ;
	wire _w12992_ ;
	wire _w12993_ ;
	wire _w12994_ ;
	wire _w12995_ ;
	wire _w12996_ ;
	wire _w12997_ ;
	wire _w12998_ ;
	wire _w12999_ ;
	wire _w13000_ ;
	wire _w13001_ ;
	wire _w13002_ ;
	wire _w13003_ ;
	wire _w13004_ ;
	wire _w13005_ ;
	wire _w13006_ ;
	wire _w13007_ ;
	wire _w13008_ ;
	wire _w13009_ ;
	wire _w13010_ ;
	wire _w13011_ ;
	wire _w13012_ ;
	wire _w13013_ ;
	wire _w13014_ ;
	wire _w13015_ ;
	wire _w13016_ ;
	wire _w13017_ ;
	wire _w13018_ ;
	wire _w13019_ ;
	wire _w13020_ ;
	wire _w13021_ ;
	wire _w13022_ ;
	wire _w13023_ ;
	wire _w13024_ ;
	wire _w13025_ ;
	wire _w13026_ ;
	wire _w13027_ ;
	wire _w13028_ ;
	wire _w13029_ ;
	wire _w13030_ ;
	wire _w13031_ ;
	wire _w13032_ ;
	wire _w13033_ ;
	wire _w13034_ ;
	wire _w13035_ ;
	wire _w13036_ ;
	wire _w13037_ ;
	wire _w13038_ ;
	wire _w13039_ ;
	wire _w13040_ ;
	wire _w13041_ ;
	wire _w13042_ ;
	wire _w13043_ ;
	wire _w13044_ ;
	wire _w13045_ ;
	wire _w13046_ ;
	wire _w13047_ ;
	wire _w13048_ ;
	wire _w13049_ ;
	wire _w13050_ ;
	wire _w13051_ ;
	wire _w13052_ ;
	wire _w13053_ ;
	wire _w13054_ ;
	wire _w13055_ ;
	wire _w13056_ ;
	wire _w13057_ ;
	wire _w13058_ ;
	wire _w13059_ ;
	wire _w13060_ ;
	wire _w13061_ ;
	wire _w13062_ ;
	wire _w13063_ ;
	wire _w13064_ ;
	wire _w13065_ ;
	wire _w13066_ ;
	wire _w13067_ ;
	wire _w13068_ ;
	wire _w13069_ ;
	wire _w13070_ ;
	wire _w13071_ ;
	wire _w13072_ ;
	wire _w13073_ ;
	wire _w13074_ ;
	wire _w13075_ ;
	wire _w13076_ ;
	wire _w13077_ ;
	wire _w13078_ ;
	wire _w13079_ ;
	wire _w13080_ ;
	wire _w13081_ ;
	wire _w13082_ ;
	wire _w13083_ ;
	wire _w13084_ ;
	wire _w13085_ ;
	wire _w13086_ ;
	wire _w13087_ ;
	wire _w13088_ ;
	wire _w13089_ ;
	wire _w13090_ ;
	wire _w13091_ ;
	wire _w13092_ ;
	wire _w13093_ ;
	wire _w13094_ ;
	wire _w13095_ ;
	wire _w13096_ ;
	wire _w13097_ ;
	wire _w13098_ ;
	wire _w13099_ ;
	wire _w13100_ ;
	wire _w13101_ ;
	wire _w13102_ ;
	wire _w13103_ ;
	wire _w13104_ ;
	wire _w13105_ ;
	wire _w13106_ ;
	wire _w13107_ ;
	wire _w13108_ ;
	wire _w13109_ ;
	wire _w13110_ ;
	wire _w13111_ ;
	wire _w13112_ ;
	wire _w13113_ ;
	wire _w13114_ ;
	wire _w13115_ ;
	wire _w13116_ ;
	wire _w13117_ ;
	wire _w13118_ ;
	wire _w13119_ ;
	wire _w13120_ ;
	wire _w13121_ ;
	wire _w13122_ ;
	wire _w13123_ ;
	wire _w13124_ ;
	wire _w13125_ ;
	wire _w13126_ ;
	wire _w13127_ ;
	wire _w13128_ ;
	wire _w13129_ ;
	wire _w13130_ ;
	wire _w13131_ ;
	wire _w13132_ ;
	wire _w13133_ ;
	wire _w13134_ ;
	wire _w13135_ ;
	wire _w13136_ ;
	wire _w13137_ ;
	wire _w13138_ ;
	wire _w13139_ ;
	wire _w13140_ ;
	wire _w13141_ ;
	wire _w13142_ ;
	wire _w13143_ ;
	wire _w13144_ ;
	wire _w13145_ ;
	wire _w13146_ ;
	wire _w13147_ ;
	wire _w13148_ ;
	wire _w13149_ ;
	wire _w13150_ ;
	wire _w13151_ ;
	wire _w13152_ ;
	wire _w13153_ ;
	wire _w13154_ ;
	wire _w13155_ ;
	wire _w13156_ ;
	wire _w13157_ ;
	wire _w13158_ ;
	wire _w13159_ ;
	wire _w13160_ ;
	wire _w13161_ ;
	wire _w13162_ ;
	wire _w13163_ ;
	wire _w13164_ ;
	wire _w13165_ ;
	wire _w13166_ ;
	wire _w13167_ ;
	wire _w13168_ ;
	wire _w13169_ ;
	wire _w13170_ ;
	wire _w13171_ ;
	wire _w13172_ ;
	wire _w13173_ ;
	wire _w13174_ ;
	wire _w13175_ ;
	wire _w13176_ ;
	wire _w13177_ ;
	wire _w13178_ ;
	wire _w13179_ ;
	wire _w13180_ ;
	wire _w13181_ ;
	wire _w13182_ ;
	wire _w13183_ ;
	wire _w13184_ ;
	wire _w13185_ ;
	wire _w13186_ ;
	wire _w13187_ ;
	wire _w13188_ ;
	wire _w13189_ ;
	wire _w13190_ ;
	wire _w13191_ ;
	wire _w13192_ ;
	wire _w13193_ ;
	wire _w13194_ ;
	wire _w13195_ ;
	wire _w13196_ ;
	wire _w13197_ ;
	wire _w13198_ ;
	wire _w13199_ ;
	wire _w13200_ ;
	wire _w13201_ ;
	wire _w13202_ ;
	wire _w13203_ ;
	wire _w13204_ ;
	wire _w13205_ ;
	wire _w13206_ ;
	wire _w13207_ ;
	wire _w13208_ ;
	wire _w13209_ ;
	wire _w13210_ ;
	wire _w13211_ ;
	wire _w13212_ ;
	wire _w13213_ ;
	wire _w13214_ ;
	wire _w13215_ ;
	wire _w13216_ ;
	wire _w13217_ ;
	wire _w13218_ ;
	wire _w13219_ ;
	wire _w13220_ ;
	wire _w13221_ ;
	wire _w13222_ ;
	wire _w13223_ ;
	wire _w13224_ ;
	wire _w13225_ ;
	wire _w13226_ ;
	wire _w13227_ ;
	wire _w13228_ ;
	wire _w13229_ ;
	wire _w13230_ ;
	wire _w13231_ ;
	wire _w13232_ ;
	wire _w13233_ ;
	wire _w13234_ ;
	wire _w13235_ ;
	wire _w13236_ ;
	wire _w13237_ ;
	wire _w13238_ ;
	wire _w13239_ ;
	wire _w13240_ ;
	wire _w13241_ ;
	wire _w13242_ ;
	wire _w13243_ ;
	wire _w13244_ ;
	wire _w13245_ ;
	wire _w13246_ ;
	wire _w13247_ ;
	wire _w13248_ ;
	wire _w13249_ ;
	wire _w13250_ ;
	wire _w13251_ ;
	wire _w13252_ ;
	wire _w13253_ ;
	wire _w13254_ ;
	wire _w13255_ ;
	wire _w13256_ ;
	wire _w13257_ ;
	wire _w13258_ ;
	wire _w13259_ ;
	wire _w13260_ ;
	wire _w13261_ ;
	wire _w13262_ ;
	wire _w13263_ ;
	wire _w13264_ ;
	wire _w13265_ ;
	wire _w13266_ ;
	wire _w13267_ ;
	wire _w13268_ ;
	wire _w13269_ ;
	wire _w13270_ ;
	wire _w13271_ ;
	wire _w13272_ ;
	wire _w13273_ ;
	wire _w13274_ ;
	wire _w13275_ ;
	wire _w13276_ ;
	wire _w13277_ ;
	wire _w13278_ ;
	wire _w13279_ ;
	wire _w13280_ ;
	wire _w13281_ ;
	wire _w13282_ ;
	wire _w13283_ ;
	wire _w13284_ ;
	wire _w13285_ ;
	wire _w13286_ ;
	wire _w13287_ ;
	wire _w13288_ ;
	wire _w13289_ ;
	wire _w13290_ ;
	wire _w13291_ ;
	wire _w13292_ ;
	wire _w13293_ ;
	wire _w13294_ ;
	wire _w13295_ ;
	wire _w13296_ ;
	wire _w13297_ ;
	wire _w13298_ ;
	wire _w13299_ ;
	wire _w13300_ ;
	wire _w13301_ ;
	wire _w13302_ ;
	wire _w13303_ ;
	wire _w13304_ ;
	wire _w13305_ ;
	wire _w13306_ ;
	wire _w13307_ ;
	wire _w13308_ ;
	wire _w13309_ ;
	wire _w13310_ ;
	wire _w13311_ ;
	wire _w13312_ ;
	wire _w13313_ ;
	wire _w13314_ ;
	wire _w13315_ ;
	wire _w13316_ ;
	wire _w13317_ ;
	wire _w13318_ ;
	wire _w13319_ ;
	wire _w13320_ ;
	wire _w13321_ ;
	wire _w13322_ ;
	wire _w13323_ ;
	wire _w13324_ ;
	wire _w13325_ ;
	wire _w13326_ ;
	wire _w13327_ ;
	wire _w13328_ ;
	wire _w13329_ ;
	wire _w13330_ ;
	wire _w13331_ ;
	wire _w13332_ ;
	wire _w13333_ ;
	wire _w13334_ ;
	wire _w13335_ ;
	wire _w13336_ ;
	wire _w13337_ ;
	wire _w13338_ ;
	wire _w13339_ ;
	wire _w13340_ ;
	wire _w13341_ ;
	wire _w13342_ ;
	wire _w13343_ ;
	wire _w13344_ ;
	wire _w13345_ ;
	wire _w13346_ ;
	wire _w13347_ ;
	wire _w13348_ ;
	wire _w13349_ ;
	wire _w13350_ ;
	wire _w13351_ ;
	wire _w13352_ ;
	wire _w13353_ ;
	wire _w13354_ ;
	wire _w13355_ ;
	wire _w13356_ ;
	wire _w13357_ ;
	wire _w13358_ ;
	wire _w13359_ ;
	wire _w13360_ ;
	wire _w13361_ ;
	wire _w13362_ ;
	wire _w13363_ ;
	wire _w13364_ ;
	wire _w13365_ ;
	wire _w13366_ ;
	wire _w13367_ ;
	wire _w13368_ ;
	wire _w13369_ ;
	wire _w13370_ ;
	wire _w13371_ ;
	wire _w13372_ ;
	wire _w13373_ ;
	wire _w13374_ ;
	wire _w13375_ ;
	wire _w13376_ ;
	wire _w13377_ ;
	wire _w13378_ ;
	wire _w13379_ ;
	wire _w13380_ ;
	wire _w13381_ ;
	wire _w13382_ ;
	wire _w13383_ ;
	wire _w13384_ ;
	wire _w13385_ ;
	wire _w13386_ ;
	wire _w13387_ ;
	wire _w13388_ ;
	wire _w13389_ ;
	wire _w13390_ ;
	wire _w13391_ ;
	wire _w13392_ ;
	wire _w13393_ ;
	wire _w13394_ ;
	wire _w13395_ ;
	wire _w13396_ ;
	wire _w13397_ ;
	wire _w13398_ ;
	wire _w13399_ ;
	wire _w13400_ ;
	wire _w13401_ ;
	wire _w13402_ ;
	wire _w13403_ ;
	wire _w13404_ ;
	wire _w13405_ ;
	wire _w13406_ ;
	wire _w13407_ ;
	wire _w13408_ ;
	wire _w13409_ ;
	wire _w13410_ ;
	wire _w13411_ ;
	wire _w13412_ ;
	wire _w13413_ ;
	wire _w13414_ ;
	wire _w13415_ ;
	wire _w13416_ ;
	wire _w13417_ ;
	wire _w13418_ ;
	wire _w13419_ ;
	wire _w13420_ ;
	wire _w13421_ ;
	wire _w13422_ ;
	wire _w13423_ ;
	wire _w13424_ ;
	wire _w13425_ ;
	wire _w13426_ ;
	wire _w13427_ ;
	wire _w13428_ ;
	wire _w13429_ ;
	wire _w13430_ ;
	wire _w13431_ ;
	wire _w13432_ ;
	wire _w13433_ ;
	wire _w13434_ ;
	wire _w13435_ ;
	wire _w13436_ ;
	wire _w13437_ ;
	wire _w13438_ ;
	wire _w13439_ ;
	wire _w13440_ ;
	wire _w13441_ ;
	wire _w13442_ ;
	wire _w13443_ ;
	wire _w13444_ ;
	wire _w13445_ ;
	wire _w13446_ ;
	wire _w13447_ ;
	wire _w13448_ ;
	wire _w13449_ ;
	wire _w13450_ ;
	wire _w13451_ ;
	wire _w13452_ ;
	wire _w13453_ ;
	wire _w13454_ ;
	wire _w13455_ ;
	wire _w13456_ ;
	wire _w13457_ ;
	wire _w13458_ ;
	wire _w13459_ ;
	wire _w13460_ ;
	wire _w13461_ ;
	wire _w13462_ ;
	wire _w13463_ ;
	wire _w13464_ ;
	wire _w13465_ ;
	wire _w13466_ ;
	wire _w13467_ ;
	wire _w13468_ ;
	wire _w13469_ ;
	wire _w13470_ ;
	wire _w13471_ ;
	wire _w13472_ ;
	wire _w13473_ ;
	wire _w13474_ ;
	wire _w13475_ ;
	wire _w13476_ ;
	wire _w13477_ ;
	wire _w13478_ ;
	wire _w13479_ ;
	wire _w13480_ ;
	wire _w13481_ ;
	wire _w13482_ ;
	wire _w13483_ ;
	wire _w13484_ ;
	wire _w13485_ ;
	wire _w13486_ ;
	wire _w13487_ ;
	wire _w13488_ ;
	wire _w13489_ ;
	wire _w13490_ ;
	wire _w13491_ ;
	wire _w13492_ ;
	wire _w13493_ ;
	wire _w13494_ ;
	wire _w13495_ ;
	wire _w13496_ ;
	wire _w13497_ ;
	wire _w13498_ ;
	wire _w13499_ ;
	wire _w13500_ ;
	wire _w13501_ ;
	wire _w13502_ ;
	wire _w13503_ ;
	wire _w13504_ ;
	wire _w13505_ ;
	wire _w13506_ ;
	wire _w13507_ ;
	wire _w13508_ ;
	wire _w13509_ ;
	wire _w13510_ ;
	wire _w13511_ ;
	wire _w13512_ ;
	wire _w13513_ ;
	wire _w13514_ ;
	wire _w13515_ ;
	wire _w13516_ ;
	wire _w13517_ ;
	wire _w13518_ ;
	wire _w13519_ ;
	wire _w13520_ ;
	wire _w13521_ ;
	wire _w13522_ ;
	wire _w13523_ ;
	wire _w13524_ ;
	wire _w13525_ ;
	wire _w13526_ ;
	wire _w13527_ ;
	wire _w13528_ ;
	wire _w13529_ ;
	wire _w13530_ ;
	wire _w13531_ ;
	wire _w13532_ ;
	wire _w13533_ ;
	wire _w13534_ ;
	wire _w13535_ ;
	wire _w13536_ ;
	wire _w13537_ ;
	wire _w13538_ ;
	wire _w13539_ ;
	wire _w13540_ ;
	wire _w13541_ ;
	wire _w13542_ ;
	wire _w13543_ ;
	wire _w13544_ ;
	wire _w13545_ ;
	wire _w13546_ ;
	wire _w13547_ ;
	wire _w13548_ ;
	wire _w13549_ ;
	wire _w13550_ ;
	wire _w13551_ ;
	wire _w13552_ ;
	wire _w13553_ ;
	wire _w13554_ ;
	wire _w13555_ ;
	wire _w13556_ ;
	wire _w13557_ ;
	wire _w13558_ ;
	wire _w13559_ ;
	wire _w13560_ ;
	wire _w13561_ ;
	wire _w13562_ ;
	wire _w13563_ ;
	wire _w13564_ ;
	wire _w13565_ ;
	wire _w13566_ ;
	wire _w13567_ ;
	wire _w13568_ ;
	wire _w13569_ ;
	wire _w13570_ ;
	wire _w13571_ ;
	wire _w13572_ ;
	wire _w13573_ ;
	wire _w13574_ ;
	wire _w13575_ ;
	wire _w13576_ ;
	wire _w13577_ ;
	wire _w13578_ ;
	wire _w13579_ ;
	wire _w13580_ ;
	wire _w13581_ ;
	wire _w13582_ ;
	wire _w13583_ ;
	wire _w13584_ ;
	wire _w13585_ ;
	wire _w13586_ ;
	wire _w13587_ ;
	wire _w13588_ ;
	wire _w13589_ ;
	wire _w13590_ ;
	wire _w13591_ ;
	wire _w13592_ ;
	wire _w13593_ ;
	wire _w13594_ ;
	wire _w13595_ ;
	wire _w13596_ ;
	wire _w13597_ ;
	wire _w13598_ ;
	wire _w13599_ ;
	wire _w13600_ ;
	wire _w13601_ ;
	wire _w13602_ ;
	wire _w13603_ ;
	wire _w13604_ ;
	wire _w13605_ ;
	wire _w13606_ ;
	wire _w13607_ ;
	wire _w13608_ ;
	wire _w13609_ ;
	wire _w13610_ ;
	wire _w13611_ ;
	wire _w13612_ ;
	wire _w13613_ ;
	wire _w13614_ ;
	wire _w13615_ ;
	wire _w13616_ ;
	wire _w13617_ ;
	wire _w13618_ ;
	wire _w13619_ ;
	wire _w13620_ ;
	wire _w13621_ ;
	wire _w13622_ ;
	wire _w13623_ ;
	wire _w13624_ ;
	wire _w13625_ ;
	wire _w13626_ ;
	wire _w13627_ ;
	wire _w13628_ ;
	wire _w13629_ ;
	wire _w13630_ ;
	wire _w13631_ ;
	wire _w13632_ ;
	wire _w13633_ ;
	wire _w13634_ ;
	wire _w13635_ ;
	wire _w13636_ ;
	wire _w13637_ ;
	wire _w13638_ ;
	wire _w13639_ ;
	wire _w13640_ ;
	wire _w13641_ ;
	wire _w13642_ ;
	wire _w13643_ ;
	wire _w13644_ ;
	wire _w13645_ ;
	wire _w13646_ ;
	wire _w13647_ ;
	wire _w13648_ ;
	wire _w13649_ ;
	wire _w13650_ ;
	wire _w13651_ ;
	wire _w13652_ ;
	wire _w13653_ ;
	wire _w13654_ ;
	wire _w13655_ ;
	wire _w13656_ ;
	wire _w13657_ ;
	wire _w13658_ ;
	wire _w13659_ ;
	wire _w13660_ ;
	wire _w13661_ ;
	wire _w13662_ ;
	wire _w13663_ ;
	wire _w13664_ ;
	wire _w13665_ ;
	wire _w13666_ ;
	wire _w13667_ ;
	wire _w13668_ ;
	wire _w13669_ ;
	wire _w13670_ ;
	wire _w13671_ ;
	wire _w13672_ ;
	wire _w13673_ ;
	wire _w13674_ ;
	wire _w13675_ ;
	wire _w13676_ ;
	wire _w13677_ ;
	wire _w13678_ ;
	wire _w13679_ ;
	wire _w13680_ ;
	wire _w13681_ ;
	wire _w13682_ ;
	wire _w13683_ ;
	wire _w13684_ ;
	wire _w13685_ ;
	wire _w13686_ ;
	wire _w13687_ ;
	wire _w13688_ ;
	wire _w13689_ ;
	wire _w13690_ ;
	wire _w13691_ ;
	wire _w13692_ ;
	wire _w13693_ ;
	wire _w13694_ ;
	wire _w13695_ ;
	wire _w13696_ ;
	wire _w13697_ ;
	wire _w13698_ ;
	wire _w13699_ ;
	wire _w13700_ ;
	wire _w13701_ ;
	wire _w13702_ ;
	wire _w13703_ ;
	wire _w13704_ ;
	wire _w13705_ ;
	wire _w13706_ ;
	wire _w13707_ ;
	wire _w13708_ ;
	wire _w13709_ ;
	wire _w13710_ ;
	wire _w13711_ ;
	wire _w13712_ ;
	wire _w13713_ ;
	wire _w13714_ ;
	wire _w13715_ ;
	wire _w13716_ ;
	wire _w13717_ ;
	wire _w13718_ ;
	wire _w13719_ ;
	wire _w13720_ ;
	wire _w13721_ ;
	wire _w13722_ ;
	wire _w13723_ ;
	wire _w13724_ ;
	wire _w13725_ ;
	wire _w13726_ ;
	wire _w13727_ ;
	wire _w13728_ ;
	wire _w13729_ ;
	wire _w13730_ ;
	wire _w13731_ ;
	wire _w13732_ ;
	wire _w13733_ ;
	wire _w13734_ ;
	wire _w13735_ ;
	wire _w13736_ ;
	wire _w13737_ ;
	wire _w13738_ ;
	wire _w13739_ ;
	wire _w13740_ ;
	wire _w13741_ ;
	wire _w13742_ ;
	wire _w13743_ ;
	wire _w13744_ ;
	wire _w13745_ ;
	wire _w13746_ ;
	wire _w13747_ ;
	wire _w13748_ ;
	wire _w13749_ ;
	wire _w13750_ ;
	wire _w13751_ ;
	wire _w13752_ ;
	wire _w13753_ ;
	wire _w13754_ ;
	wire _w13755_ ;
	wire _w13756_ ;
	wire _w13757_ ;
	wire _w13758_ ;
	wire _w13759_ ;
	wire _w13760_ ;
	wire _w13761_ ;
	wire _w13762_ ;
	wire _w13763_ ;
	wire _w13764_ ;
	wire _w13765_ ;
	wire _w13766_ ;
	wire _w13767_ ;
	wire _w13768_ ;
	wire _w13769_ ;
	wire _w13770_ ;
	wire _w13771_ ;
	wire _w13772_ ;
	wire _w13773_ ;
	wire _w13774_ ;
	wire _w13775_ ;
	wire _w13776_ ;
	wire _w13777_ ;
	wire _w13778_ ;
	wire _w13779_ ;
	wire _w13780_ ;
	wire _w13781_ ;
	wire _w13782_ ;
	wire _w13783_ ;
	wire _w13784_ ;
	wire _w13785_ ;
	wire _w13786_ ;
	wire _w13787_ ;
	wire _w13788_ ;
	wire _w13789_ ;
	wire _w13790_ ;
	wire _w13791_ ;
	wire _w13792_ ;
	wire _w13793_ ;
	wire _w13794_ ;
	wire _w13795_ ;
	wire _w13796_ ;
	wire _w13797_ ;
	wire _w13798_ ;
	wire _w13799_ ;
	wire _w13800_ ;
	wire _w13801_ ;
	wire _w13802_ ;
	wire _w13803_ ;
	wire _w13804_ ;
	wire _w13805_ ;
	wire _w13806_ ;
	wire _w13807_ ;
	wire _w13808_ ;
	wire _w13809_ ;
	wire _w13810_ ;
	wire _w13811_ ;
	wire _w13812_ ;
	wire _w13813_ ;
	wire _w13814_ ;
	wire _w13815_ ;
	wire _w13816_ ;
	wire _w13817_ ;
	wire _w13818_ ;
	wire _w13819_ ;
	wire _w13820_ ;
	wire _w13821_ ;
	wire _w13822_ ;
	wire _w13823_ ;
	wire _w13824_ ;
	wire _w13825_ ;
	wire _w13826_ ;
	wire _w13827_ ;
	wire _w13828_ ;
	wire _w13829_ ;
	wire _w13830_ ;
	wire _w13831_ ;
	wire _w13832_ ;
	wire _w13833_ ;
	wire _w13834_ ;
	wire _w13835_ ;
	wire _w13836_ ;
	wire _w13837_ ;
	wire _w13838_ ;
	wire _w13839_ ;
	wire _w13840_ ;
	wire _w13841_ ;
	wire _w13842_ ;
	wire _w13843_ ;
	wire _w13844_ ;
	wire _w13845_ ;
	wire _w13846_ ;
	wire _w13847_ ;
	wire _w13848_ ;
	wire _w13849_ ;
	wire _w13850_ ;
	wire _w13851_ ;
	wire _w13852_ ;
	wire _w13853_ ;
	wire _w13854_ ;
	wire _w13855_ ;
	wire _w13856_ ;
	wire _w13857_ ;
	wire _w13858_ ;
	wire _w13859_ ;
	wire _w13860_ ;
	wire _w13861_ ;
	wire _w13862_ ;
	wire _w13863_ ;
	wire _w13864_ ;
	wire _w13865_ ;
	wire _w13866_ ;
	wire _w13867_ ;
	wire _w13868_ ;
	wire _w13869_ ;
	wire _w13870_ ;
	wire _w13871_ ;
	wire _w13872_ ;
	wire _w13873_ ;
	wire _w13874_ ;
	wire _w13875_ ;
	wire _w13876_ ;
	wire _w13877_ ;
	wire _w13878_ ;
	wire _w13879_ ;
	wire _w13880_ ;
	wire _w13881_ ;
	wire _w13882_ ;
	wire _w13883_ ;
	wire _w13884_ ;
	wire _w13885_ ;
	wire _w13886_ ;
	wire _w13887_ ;
	wire _w13888_ ;
	wire _w13889_ ;
	wire _w13890_ ;
	wire _w13891_ ;
	wire _w13892_ ;
	wire _w13893_ ;
	wire _w13894_ ;
	wire _w13895_ ;
	wire _w13896_ ;
	wire _w13897_ ;
	wire _w13898_ ;
	wire _w13899_ ;
	wire _w13900_ ;
	wire _w13901_ ;
	wire _w13902_ ;
	wire _w13903_ ;
	wire _w13904_ ;
	wire _w13905_ ;
	wire _w13906_ ;
	wire _w13907_ ;
	wire _w13908_ ;
	wire _w13909_ ;
	wire _w13910_ ;
	wire _w13911_ ;
	wire _w13912_ ;
	wire _w13913_ ;
	wire _w13914_ ;
	wire _w13915_ ;
	wire _w13916_ ;
	wire _w13917_ ;
	wire _w13918_ ;
	wire _w13919_ ;
	wire _w13920_ ;
	wire _w13921_ ;
	wire _w13922_ ;
	wire _w13923_ ;
	wire _w13924_ ;
	wire _w13925_ ;
	wire _w13926_ ;
	wire _w13927_ ;
	wire _w13928_ ;
	wire _w13929_ ;
	wire _w13930_ ;
	wire _w13931_ ;
	wire _w13932_ ;
	wire _w13933_ ;
	wire _w13934_ ;
	wire _w13935_ ;
	wire _w13936_ ;
	wire _w13937_ ;
	wire _w13938_ ;
	wire _w13939_ ;
	wire _w13940_ ;
	wire _w13941_ ;
	wire _w13942_ ;
	wire _w13943_ ;
	wire _w13944_ ;
	wire _w13945_ ;
	wire _w13946_ ;
	wire _w13947_ ;
	wire _w13948_ ;
	wire _w13949_ ;
	wire _w13950_ ;
	wire _w13951_ ;
	wire _w13952_ ;
	wire _w13953_ ;
	wire _w13954_ ;
	wire _w13955_ ;
	wire _w13956_ ;
	wire _w13957_ ;
	wire _w13958_ ;
	wire _w13959_ ;
	wire _w13960_ ;
	wire _w13961_ ;
	wire _w13962_ ;
	wire _w13963_ ;
	wire _w13964_ ;
	wire _w13965_ ;
	wire _w13966_ ;
	wire _w13967_ ;
	wire _w13968_ ;
	wire _w13969_ ;
	wire _w13970_ ;
	wire _w13971_ ;
	wire _w13972_ ;
	wire _w13973_ ;
	wire _w13974_ ;
	wire _w13975_ ;
	wire _w13976_ ;
	wire _w13977_ ;
	wire _w13978_ ;
	wire _w13979_ ;
	wire _w13980_ ;
	wire _w13981_ ;
	wire _w13982_ ;
	wire _w13983_ ;
	wire _w13984_ ;
	wire _w13985_ ;
	wire _w13986_ ;
	wire _w13987_ ;
	wire _w13988_ ;
	wire _w13989_ ;
	wire _w13990_ ;
	wire _w13991_ ;
	wire _w13992_ ;
	wire _w13993_ ;
	wire _w13994_ ;
	wire _w13995_ ;
	wire _w13996_ ;
	wire _w13997_ ;
	wire _w13998_ ;
	wire _w13999_ ;
	wire _w14000_ ;
	wire _w14001_ ;
	wire _w14002_ ;
	wire _w14003_ ;
	wire _w14004_ ;
	wire _w14005_ ;
	wire _w14006_ ;
	wire _w14007_ ;
	wire _w14008_ ;
	wire _w14009_ ;
	wire _w14010_ ;
	wire _w14011_ ;
	wire _w14012_ ;
	wire _w14013_ ;
	wire _w14014_ ;
	wire _w14015_ ;
	wire _w14016_ ;
	wire _w14017_ ;
	wire _w14018_ ;
	wire _w14019_ ;
	wire _w14020_ ;
	wire _w14021_ ;
	wire _w14022_ ;
	wire _w14023_ ;
	wire _w14024_ ;
	wire _w14025_ ;
	wire _w14026_ ;
	wire _w14027_ ;
	wire _w14028_ ;
	wire _w14029_ ;
	wire _w14030_ ;
	wire _w14031_ ;
	wire _w14032_ ;
	wire _w14033_ ;
	wire _w14034_ ;
	wire _w14035_ ;
	wire _w14036_ ;
	wire _w14037_ ;
	wire _w14038_ ;
	wire _w14039_ ;
	wire _w14040_ ;
	wire _w14041_ ;
	wire _w14042_ ;
	wire _w14043_ ;
	wire _w14044_ ;
	wire _w14045_ ;
	wire _w14046_ ;
	wire _w14047_ ;
	wire _w14048_ ;
	wire _w14049_ ;
	wire _w14050_ ;
	wire _w14051_ ;
	wire _w14052_ ;
	wire _w14053_ ;
	wire _w14054_ ;
	wire _w14055_ ;
	wire _w14056_ ;
	wire _w14057_ ;
	wire _w14058_ ;
	wire _w14059_ ;
	wire _w14060_ ;
	wire _w14061_ ;
	wire _w14062_ ;
	wire _w14063_ ;
	wire _w14064_ ;
	wire _w14065_ ;
	wire _w14066_ ;
	wire _w14067_ ;
	wire _w14068_ ;
	wire _w14069_ ;
	wire _w14070_ ;
	wire _w14071_ ;
	wire _w14072_ ;
	wire _w14073_ ;
	wire _w14074_ ;
	wire _w14075_ ;
	wire _w14076_ ;
	wire _w14077_ ;
	wire _w14078_ ;
	wire _w14079_ ;
	wire _w14080_ ;
	wire _w14081_ ;
	wire _w14082_ ;
	wire _w14083_ ;
	wire _w14084_ ;
	wire _w14085_ ;
	wire _w14086_ ;
	wire _w14087_ ;
	wire _w14088_ ;
	wire _w14089_ ;
	wire _w14090_ ;
	wire _w14091_ ;
	wire _w14092_ ;
	wire _w14093_ ;
	wire _w14094_ ;
	wire _w14095_ ;
	wire _w14096_ ;
	wire _w14097_ ;
	wire _w14098_ ;
	wire _w14099_ ;
	wire _w14100_ ;
	wire _w14101_ ;
	wire _w14102_ ;
	wire _w14103_ ;
	wire _w14104_ ;
	wire _w14105_ ;
	wire _w14106_ ;
	wire _w14107_ ;
	wire _w14108_ ;
	wire _w14109_ ;
	wire _w14110_ ;
	wire _w14111_ ;
	wire _w14112_ ;
	wire _w14113_ ;
	wire _w14114_ ;
	wire _w14115_ ;
	wire _w14116_ ;
	wire _w14117_ ;
	wire _w14118_ ;
	wire _w14119_ ;
	wire _w14120_ ;
	wire _w14121_ ;
	wire _w14122_ ;
	wire _w14123_ ;
	wire _w14124_ ;
	wire _w14125_ ;
	wire _w14126_ ;
	wire _w14127_ ;
	wire _w14128_ ;
	wire _w14129_ ;
	wire _w14130_ ;
	wire _w14131_ ;
	wire _w14132_ ;
	wire _w14133_ ;
	wire _w14134_ ;
	wire _w14135_ ;
	wire _w14136_ ;
	wire _w14137_ ;
	wire _w14138_ ;
	wire _w14139_ ;
	wire _w14140_ ;
	wire _w14141_ ;
	wire _w14142_ ;
	wire _w14143_ ;
	wire _w14144_ ;
	wire _w14145_ ;
	wire _w14146_ ;
	wire _w14147_ ;
	wire _w14148_ ;
	wire _w14149_ ;
	wire _w14150_ ;
	wire _w14151_ ;
	wire _w14152_ ;
	wire _w14153_ ;
	wire _w14154_ ;
	wire _w14155_ ;
	wire _w14156_ ;
	wire _w14157_ ;
	wire _w14158_ ;
	wire _w14159_ ;
	wire _w14160_ ;
	wire _w14161_ ;
	wire _w14162_ ;
	wire _w14163_ ;
	wire _w14164_ ;
	wire _w14165_ ;
	wire _w14166_ ;
	wire _w14167_ ;
	wire _w14168_ ;
	wire _w14169_ ;
	wire _w14170_ ;
	wire _w14171_ ;
	wire _w14172_ ;
	wire _w14173_ ;
	wire _w14174_ ;
	wire _w14175_ ;
	wire _w14176_ ;
	wire _w14177_ ;
	wire _w14178_ ;
	wire _w14179_ ;
	wire _w14180_ ;
	wire _w14181_ ;
	wire _w14182_ ;
	wire _w14183_ ;
	wire _w14184_ ;
	wire _w14185_ ;
	wire _w14186_ ;
	wire _w14187_ ;
	wire _w14188_ ;
	wire _w14189_ ;
	wire _w14190_ ;
	wire _w14191_ ;
	wire _w14192_ ;
	wire _w14193_ ;
	wire _w14194_ ;
	wire _w14195_ ;
	wire _w14196_ ;
	wire _w14197_ ;
	wire _w14198_ ;
	wire _w14199_ ;
	wire _w14200_ ;
	wire _w14201_ ;
	wire _w14202_ ;
	wire _w14203_ ;
	wire _w14204_ ;
	wire _w14205_ ;
	wire _w14206_ ;
	wire _w14207_ ;
	wire _w14208_ ;
	wire _w14209_ ;
	wire _w14210_ ;
	wire _w14211_ ;
	wire _w14212_ ;
	wire _w14213_ ;
	wire _w14214_ ;
	wire _w14215_ ;
	wire _w14216_ ;
	wire _w14217_ ;
	wire _w14218_ ;
	wire _w14219_ ;
	wire _w14220_ ;
	wire _w14221_ ;
	wire _w14222_ ;
	wire _w14223_ ;
	wire _w14224_ ;
	wire _w14225_ ;
	wire _w14226_ ;
	wire _w14227_ ;
	wire _w14228_ ;
	wire _w14229_ ;
	wire _w14230_ ;
	wire _w14231_ ;
	wire _w14232_ ;
	wire _w14233_ ;
	wire _w14234_ ;
	wire _w14235_ ;
	wire _w14236_ ;
	wire _w14237_ ;
	wire _w14238_ ;
	wire _w14239_ ;
	wire _w14240_ ;
	wire _w14241_ ;
	wire _w14242_ ;
	wire _w14243_ ;
	wire _w14244_ ;
	wire _w14245_ ;
	wire _w14246_ ;
	wire _w14247_ ;
	wire _w14248_ ;
	wire _w14249_ ;
	wire _w14250_ ;
	wire _w14251_ ;
	wire _w14252_ ;
	wire _w14253_ ;
	wire _w14254_ ;
	wire _w14255_ ;
	wire _w14256_ ;
	wire _w14257_ ;
	wire _w14258_ ;
	wire _w14259_ ;
	wire _w14260_ ;
	wire _w14261_ ;
	wire _w14262_ ;
	wire _w14263_ ;
	wire _w14264_ ;
	wire _w14265_ ;
	wire _w14266_ ;
	wire _w14267_ ;
	wire _w14268_ ;
	wire _w14269_ ;
	wire _w14270_ ;
	wire _w14271_ ;
	wire _w14272_ ;
	wire _w14273_ ;
	wire _w14274_ ;
	wire _w14275_ ;
	wire _w14276_ ;
	wire _w14277_ ;
	wire _w14278_ ;
	wire _w14279_ ;
	wire _w14280_ ;
	wire _w14281_ ;
	wire _w14282_ ;
	wire _w14283_ ;
	wire _w14284_ ;
	wire _w14285_ ;
	wire _w14286_ ;
	wire _w14287_ ;
	wire _w14288_ ;
	wire _w14289_ ;
	wire _w14290_ ;
	wire _w14291_ ;
	wire _w14292_ ;
	wire _w14293_ ;
	wire _w14294_ ;
	wire _w14295_ ;
	wire _w14296_ ;
	wire _w14297_ ;
	wire _w14298_ ;
	wire _w14299_ ;
	wire _w14300_ ;
	wire _w14301_ ;
	wire _w14302_ ;
	wire _w14303_ ;
	wire _w14304_ ;
	wire _w14305_ ;
	wire _w14306_ ;
	wire _w14307_ ;
	wire _w14308_ ;
	wire _w14309_ ;
	wire _w14310_ ;
	wire _w14311_ ;
	wire _w14312_ ;
	wire _w14313_ ;
	wire _w14314_ ;
	wire _w14315_ ;
	wire _w14316_ ;
	wire _w14317_ ;
	wire _w14318_ ;
	wire _w14319_ ;
	wire _w14320_ ;
	wire _w14321_ ;
	wire _w14322_ ;
	wire _w14323_ ;
	wire _w14324_ ;
	wire _w14325_ ;
	wire _w14326_ ;
	wire _w14327_ ;
	wire _w14328_ ;
	wire _w14329_ ;
	wire _w14330_ ;
	wire _w14331_ ;
	wire _w14332_ ;
	wire _w14333_ ;
	wire _w14334_ ;
	wire _w14335_ ;
	wire _w14336_ ;
	wire _w14337_ ;
	wire _w14338_ ;
	wire _w14339_ ;
	wire _w14340_ ;
	wire _w14341_ ;
	wire _w14342_ ;
	wire _w14343_ ;
	wire _w14344_ ;
	wire _w14345_ ;
	wire _w14346_ ;
	wire _w14347_ ;
	wire _w14348_ ;
	wire _w14349_ ;
	wire _w14350_ ;
	wire _w14351_ ;
	wire _w14352_ ;
	wire _w14353_ ;
	wire _w14354_ ;
	wire _w14355_ ;
	wire _w14356_ ;
	wire _w14357_ ;
	wire _w14358_ ;
	wire _w14359_ ;
	wire _w14360_ ;
	wire _w14361_ ;
	wire _w14362_ ;
	wire _w14363_ ;
	wire _w14364_ ;
	wire _w14365_ ;
	wire _w14366_ ;
	wire _w14367_ ;
	wire _w14368_ ;
	wire _w14369_ ;
	wire _w14370_ ;
	wire _w14371_ ;
	wire _w14372_ ;
	wire _w14373_ ;
	wire _w14374_ ;
	wire _w14375_ ;
	wire _w14376_ ;
	wire _w14377_ ;
	wire _w14378_ ;
	wire _w14379_ ;
	wire _w14380_ ;
	wire _w14381_ ;
	wire _w14382_ ;
	wire _w14383_ ;
	wire _w14384_ ;
	wire _w14385_ ;
	wire _w14386_ ;
	wire _w14387_ ;
	wire _w14388_ ;
	wire _w14389_ ;
	wire _w14390_ ;
	wire _w14391_ ;
	wire _w14392_ ;
	wire _w14393_ ;
	wire _w14394_ ;
	wire _w14395_ ;
	wire _w14396_ ;
	wire _w14397_ ;
	wire _w14398_ ;
	wire _w14399_ ;
	wire _w14400_ ;
	wire _w14401_ ;
	wire _w14402_ ;
	wire _w14403_ ;
	wire _w14404_ ;
	wire _w14405_ ;
	wire _w14406_ ;
	wire _w14407_ ;
	wire _w14408_ ;
	wire _w14409_ ;
	wire _w14410_ ;
	wire _w14411_ ;
	wire _w14412_ ;
	wire _w14413_ ;
	wire _w14414_ ;
	wire _w14415_ ;
	wire _w14416_ ;
	wire _w14417_ ;
	wire _w14418_ ;
	wire _w14419_ ;
	wire _w14420_ ;
	wire _w14421_ ;
	wire _w14422_ ;
	wire _w14423_ ;
	wire _w14424_ ;
	wire _w14425_ ;
	wire _w14426_ ;
	wire _w14427_ ;
	wire _w14428_ ;
	wire _w14429_ ;
	wire _w14430_ ;
	wire _w14431_ ;
	wire _w14432_ ;
	wire _w14433_ ;
	wire _w14434_ ;
	wire _w14435_ ;
	wire _w14436_ ;
	wire _w14437_ ;
	wire _w14438_ ;
	wire _w14439_ ;
	wire _w14440_ ;
	wire _w14441_ ;
	wire _w14442_ ;
	wire _w14443_ ;
	wire _w14444_ ;
	wire _w14445_ ;
	wire _w14446_ ;
	wire _w14447_ ;
	wire _w14448_ ;
	wire _w14449_ ;
	wire _w14450_ ;
	wire _w14451_ ;
	wire _w14452_ ;
	wire _w14453_ ;
	wire _w14454_ ;
	wire _w14455_ ;
	wire _w14456_ ;
	wire _w14457_ ;
	wire _w14458_ ;
	wire _w14459_ ;
	wire _w14460_ ;
	wire _w14461_ ;
	wire _w14462_ ;
	wire _w14463_ ;
	wire _w14464_ ;
	wire _w14465_ ;
	wire _w14466_ ;
	wire _w14467_ ;
	wire _w14468_ ;
	wire _w14469_ ;
	wire _w14470_ ;
	wire _w14471_ ;
	wire _w14472_ ;
	wire _w14473_ ;
	wire _w14474_ ;
	wire _w14475_ ;
	wire _w14476_ ;
	wire _w14477_ ;
	wire _w14478_ ;
	wire _w14479_ ;
	wire _w14480_ ;
	wire _w14481_ ;
	wire _w14482_ ;
	wire _w14483_ ;
	wire _w14484_ ;
	wire _w14485_ ;
	wire _w14486_ ;
	wire _w14487_ ;
	wire _w14488_ ;
	wire _w14489_ ;
	wire _w14490_ ;
	wire _w14491_ ;
	wire _w14492_ ;
	wire _w14493_ ;
	wire _w14494_ ;
	wire _w14495_ ;
	wire _w14496_ ;
	wire _w14497_ ;
	wire _w14498_ ;
	wire _w14499_ ;
	wire _w14500_ ;
	wire _w14501_ ;
	wire _w14502_ ;
	wire _w14503_ ;
	wire _w14504_ ;
	wire _w14505_ ;
	wire _w14506_ ;
	wire _w14507_ ;
	wire _w14508_ ;
	wire _w14509_ ;
	wire _w14510_ ;
	wire _w14511_ ;
	wire _w14512_ ;
	wire _w14513_ ;
	wire _w14514_ ;
	wire _w14515_ ;
	wire _w14516_ ;
	wire _w14517_ ;
	wire _w14518_ ;
	wire _w14519_ ;
	wire _w14520_ ;
	wire _w14521_ ;
	wire _w14522_ ;
	wire _w14523_ ;
	wire _w14524_ ;
	wire _w14525_ ;
	wire _w14526_ ;
	wire _w14527_ ;
	wire _w14528_ ;
	wire _w14529_ ;
	wire _w14530_ ;
	wire _w14531_ ;
	wire _w14532_ ;
	wire _w14533_ ;
	wire _w14534_ ;
	wire _w14535_ ;
	wire _w14536_ ;
	wire _w14537_ ;
	wire _w14538_ ;
	wire _w14539_ ;
	wire _w14540_ ;
	wire _w14541_ ;
	wire _w14542_ ;
	wire _w14543_ ;
	wire _w14544_ ;
	wire _w14545_ ;
	wire _w14546_ ;
	wire _w14547_ ;
	wire _w14548_ ;
	wire _w14549_ ;
	wire _w14550_ ;
	wire _w14551_ ;
	wire _w14552_ ;
	wire _w14553_ ;
	wire _w14554_ ;
	wire _w14555_ ;
	wire _w14556_ ;
	wire _w14557_ ;
	wire _w14558_ ;
	wire _w14559_ ;
	wire _w14560_ ;
	wire _w14561_ ;
	wire _w14562_ ;
	wire _w14563_ ;
	wire _w14564_ ;
	wire _w14565_ ;
	wire _w14566_ ;
	wire _w14567_ ;
	wire _w14568_ ;
	wire _w14569_ ;
	wire _w14570_ ;
	wire _w14571_ ;
	wire _w14572_ ;
	wire _w14573_ ;
	wire _w14574_ ;
	wire _w14575_ ;
	wire _w14576_ ;
	wire _w14577_ ;
	wire _w14578_ ;
	wire _w14579_ ;
	wire _w14580_ ;
	wire _w14581_ ;
	wire _w14582_ ;
	wire _w14583_ ;
	wire _w14584_ ;
	wire _w14585_ ;
	wire _w14586_ ;
	wire _w14587_ ;
	wire _w14588_ ;
	wire _w14589_ ;
	wire _w14590_ ;
	wire _w14591_ ;
	wire _w14592_ ;
	wire _w14593_ ;
	wire _w14594_ ;
	wire _w14595_ ;
	wire _w14596_ ;
	wire _w14597_ ;
	wire _w14598_ ;
	wire _w14599_ ;
	wire _w14600_ ;
	wire _w14601_ ;
	wire _w14602_ ;
	wire _w14603_ ;
	wire _w14604_ ;
	wire _w14605_ ;
	wire _w14606_ ;
	wire _w14607_ ;
	wire _w14608_ ;
	wire _w14609_ ;
	wire _w14610_ ;
	wire _w14611_ ;
	wire _w14612_ ;
	wire _w14613_ ;
	wire _w14614_ ;
	wire _w14615_ ;
	wire _w14616_ ;
	wire _w14617_ ;
	wire _w14618_ ;
	wire _w14619_ ;
	wire _w14620_ ;
	wire _w14621_ ;
	wire _w14622_ ;
	wire _w14623_ ;
	wire _w14624_ ;
	wire _w14625_ ;
	wire _w14626_ ;
	wire _w14627_ ;
	wire _w14628_ ;
	wire _w14629_ ;
	wire _w14630_ ;
	wire _w14631_ ;
	wire _w14632_ ;
	wire _w14633_ ;
	wire _w14634_ ;
	wire _w14635_ ;
	wire _w14636_ ;
	wire _w14637_ ;
	wire _w14638_ ;
	wire _w14639_ ;
	wire _w14640_ ;
	wire _w14641_ ;
	wire _w14642_ ;
	wire _w14643_ ;
	wire _w14644_ ;
	wire _w14645_ ;
	wire _w14646_ ;
	wire _w14647_ ;
	wire _w14648_ ;
	wire _w14649_ ;
	wire _w14650_ ;
	wire _w14651_ ;
	wire _w14652_ ;
	wire _w14653_ ;
	wire _w14654_ ;
	wire _w14655_ ;
	wire _w14656_ ;
	wire _w14657_ ;
	wire _w14658_ ;
	wire _w14659_ ;
	wire _w14660_ ;
	wire _w14661_ ;
	wire _w14662_ ;
	wire _w14663_ ;
	wire _w14664_ ;
	wire _w14665_ ;
	wire _w14666_ ;
	wire _w14667_ ;
	wire _w14668_ ;
	wire _w14669_ ;
	wire _w14670_ ;
	wire _w14671_ ;
	wire _w14672_ ;
	wire _w14673_ ;
	wire _w14674_ ;
	wire _w14675_ ;
	wire _w14676_ ;
	wire _w14677_ ;
	wire _w14678_ ;
	wire _w14679_ ;
	wire _w14680_ ;
	wire _w14681_ ;
	wire _w14682_ ;
	wire _w14683_ ;
	wire _w14684_ ;
	wire _w14685_ ;
	wire _w14686_ ;
	wire _w14687_ ;
	wire _w14688_ ;
	wire _w14689_ ;
	wire _w14690_ ;
	wire _w14691_ ;
	wire _w14692_ ;
	wire _w14693_ ;
	wire _w14694_ ;
	wire _w14695_ ;
	wire _w14696_ ;
	wire _w14697_ ;
	wire _w14698_ ;
	wire _w14699_ ;
	wire _w14700_ ;
	wire _w14701_ ;
	wire _w14702_ ;
	wire _w14703_ ;
	wire _w14704_ ;
	wire _w14705_ ;
	wire _w14706_ ;
	wire _w14707_ ;
	wire _w14708_ ;
	wire _w14709_ ;
	wire _w14710_ ;
	wire _w14711_ ;
	wire _w14712_ ;
	wire _w14713_ ;
	wire _w14714_ ;
	wire _w14715_ ;
	wire _w14716_ ;
	wire _w14717_ ;
	wire _w14718_ ;
	wire _w14719_ ;
	wire _w14720_ ;
	wire _w14721_ ;
	wire _w14722_ ;
	wire _w14723_ ;
	wire _w14724_ ;
	wire _w14725_ ;
	wire _w14726_ ;
	wire _w14727_ ;
	wire _w14728_ ;
	wire _w14729_ ;
	wire _w14730_ ;
	wire _w14731_ ;
	wire _w14732_ ;
	wire _w14733_ ;
	wire _w14734_ ;
	wire _w14735_ ;
	wire _w14736_ ;
	wire _w14737_ ;
	wire _w14738_ ;
	wire _w14739_ ;
	wire _w14740_ ;
	wire _w14741_ ;
	wire _w14742_ ;
	wire _w14743_ ;
	wire _w14744_ ;
	wire _w14745_ ;
	wire _w14746_ ;
	wire _w14747_ ;
	wire _w14748_ ;
	wire _w14749_ ;
	wire _w14750_ ;
	wire _w14751_ ;
	wire _w14752_ ;
	wire _w14753_ ;
	wire _w14754_ ;
	wire _w14755_ ;
	wire _w14756_ ;
	wire _w14757_ ;
	wire _w14758_ ;
	wire _w14759_ ;
	wire _w14760_ ;
	wire _w14761_ ;
	wire _w14762_ ;
	wire _w14763_ ;
	wire _w14764_ ;
	wire _w14765_ ;
	wire _w14766_ ;
	wire _w14767_ ;
	wire _w14768_ ;
	wire _w14769_ ;
	wire _w14770_ ;
	wire _w14771_ ;
	wire _w14772_ ;
	wire _w14773_ ;
	wire _w14774_ ;
	wire _w14775_ ;
	wire _w14776_ ;
	wire _w14777_ ;
	wire _w14778_ ;
	wire _w14779_ ;
	wire _w14780_ ;
	wire _w14781_ ;
	wire _w14782_ ;
	wire _w14783_ ;
	wire _w14784_ ;
	wire _w14785_ ;
	wire _w14786_ ;
	wire _w14787_ ;
	wire _w14788_ ;
	wire _w14789_ ;
	wire _w14790_ ;
	wire _w14791_ ;
	wire _w14792_ ;
	wire _w14793_ ;
	wire _w14794_ ;
	wire _w14795_ ;
	wire _w14796_ ;
	wire _w14797_ ;
	wire _w14798_ ;
	wire _w14799_ ;
	wire _w14800_ ;
	wire _w14801_ ;
	wire _w14802_ ;
	wire _w14803_ ;
	wire _w14804_ ;
	wire _w14805_ ;
	wire _w14806_ ;
	wire _w14807_ ;
	wire _w14808_ ;
	wire _w14809_ ;
	wire _w14810_ ;
	wire _w14811_ ;
	wire _w14812_ ;
	wire _w14813_ ;
	wire _w14814_ ;
	wire _w14815_ ;
	wire _w14816_ ;
	wire _w14817_ ;
	wire _w14818_ ;
	wire _w14819_ ;
	wire _w14820_ ;
	wire _w14821_ ;
	wire _w14822_ ;
	wire _w14823_ ;
	wire _w14824_ ;
	wire _w14825_ ;
	wire _w14826_ ;
	wire _w14827_ ;
	wire _w14828_ ;
	wire _w14829_ ;
	wire _w14830_ ;
	wire _w14831_ ;
	wire _w14832_ ;
	wire _w14833_ ;
	wire _w14834_ ;
	wire _w14835_ ;
	wire _w14836_ ;
	wire _w14837_ ;
	wire _w14838_ ;
	wire _w14839_ ;
	wire _w14840_ ;
	wire _w14841_ ;
	wire _w14842_ ;
	wire _w14843_ ;
	wire _w14844_ ;
	wire _w14845_ ;
	wire _w14846_ ;
	wire _w14847_ ;
	wire _w14848_ ;
	wire _w14849_ ;
	wire _w14850_ ;
	wire _w14851_ ;
	wire _w14852_ ;
	wire _w14853_ ;
	wire _w14854_ ;
	wire _w14855_ ;
	wire _w14856_ ;
	wire _w14857_ ;
	wire _w14858_ ;
	wire _w14859_ ;
	wire _w14860_ ;
	wire _w14861_ ;
	wire _w14862_ ;
	wire _w14863_ ;
	wire _w14864_ ;
	wire _w14865_ ;
	wire _w14866_ ;
	wire _w14867_ ;
	wire _w14868_ ;
	wire _w14869_ ;
	wire _w14870_ ;
	wire _w14871_ ;
	wire _w14872_ ;
	wire _w14873_ ;
	wire _w14874_ ;
	wire _w14875_ ;
	wire _w14876_ ;
	wire _w14877_ ;
	wire _w14878_ ;
	wire _w14879_ ;
	wire _w14880_ ;
	wire _w14881_ ;
	wire _w14882_ ;
	wire _w14883_ ;
	wire _w14884_ ;
	wire _w14885_ ;
	wire _w14886_ ;
	wire _w14887_ ;
	wire _w14888_ ;
	wire _w14889_ ;
	wire _w14890_ ;
	wire _w14891_ ;
	wire _w14892_ ;
	wire _w14893_ ;
	wire _w14894_ ;
	wire _w14895_ ;
	wire _w14896_ ;
	wire _w14897_ ;
	wire _w14898_ ;
	wire _w14899_ ;
	wire _w14900_ ;
	wire _w14901_ ;
	wire _w14902_ ;
	wire _w14903_ ;
	wire _w14904_ ;
	wire _w14905_ ;
	wire _w14906_ ;
	wire _w14907_ ;
	wire _w14908_ ;
	wire _w14909_ ;
	wire _w14910_ ;
	wire _w14911_ ;
	wire _w14912_ ;
	wire _w14913_ ;
	wire _w14914_ ;
	wire _w14915_ ;
	wire _w14916_ ;
	wire _w14917_ ;
	wire _w14918_ ;
	wire _w14919_ ;
	wire _w14920_ ;
	wire _w14921_ ;
	wire _w14922_ ;
	wire _w14923_ ;
	wire _w14924_ ;
	wire _w14925_ ;
	wire _w14926_ ;
	wire _w14927_ ;
	wire _w14928_ ;
	wire _w14929_ ;
	wire _w14930_ ;
	wire _w14931_ ;
	wire _w14932_ ;
	wire _w14933_ ;
	wire _w14934_ ;
	wire _w14935_ ;
	wire _w14936_ ;
	wire _w14937_ ;
	wire _w14938_ ;
	wire _w14939_ ;
	wire _w14940_ ;
	wire _w14941_ ;
	wire _w14942_ ;
	wire _w14943_ ;
	wire _w14944_ ;
	wire _w14945_ ;
	wire _w14946_ ;
	wire _w14947_ ;
	wire _w14948_ ;
	wire _w14949_ ;
	wire _w14950_ ;
	wire _w14951_ ;
	wire _w14952_ ;
	wire _w14953_ ;
	wire _w14954_ ;
	wire _w14955_ ;
	wire _w14956_ ;
	wire _w14957_ ;
	wire _w14958_ ;
	wire _w14959_ ;
	wire _w14960_ ;
	wire _w14961_ ;
	wire _w14962_ ;
	wire _w14963_ ;
	wire _w14964_ ;
	wire _w14965_ ;
	wire _w14966_ ;
	wire _w14967_ ;
	wire _w14968_ ;
	wire _w14969_ ;
	wire _w14970_ ;
	wire _w14971_ ;
	wire _w14972_ ;
	wire _w14973_ ;
	wire _w14974_ ;
	wire _w14975_ ;
	wire _w14976_ ;
	wire _w14977_ ;
	wire _w14978_ ;
	wire _w14979_ ;
	wire _w14980_ ;
	wire _w14981_ ;
	wire _w14982_ ;
	wire _w14983_ ;
	wire _w14984_ ;
	wire _w14985_ ;
	wire _w14986_ ;
	wire _w14987_ ;
	wire _w14988_ ;
	wire _w14989_ ;
	wire _w14990_ ;
	wire _w14991_ ;
	wire _w14992_ ;
	wire _w14993_ ;
	wire _w14994_ ;
	wire _w14995_ ;
	wire _w14996_ ;
	wire _w14997_ ;
	wire _w14998_ ;
	wire _w14999_ ;
	wire _w15000_ ;
	wire _w15001_ ;
	wire _w15002_ ;
	wire _w15003_ ;
	wire _w15004_ ;
	wire _w15005_ ;
	wire _w15006_ ;
	wire _w15007_ ;
	wire _w15008_ ;
	wire _w15009_ ;
	wire _w15010_ ;
	wire _w15011_ ;
	wire _w15012_ ;
	wire _w15013_ ;
	wire _w15014_ ;
	wire _w15015_ ;
	wire _w15016_ ;
	wire _w15017_ ;
	wire _w15018_ ;
	wire _w15019_ ;
	wire _w15020_ ;
	wire _w15021_ ;
	wire _w15022_ ;
	wire _w15023_ ;
	wire _w15024_ ;
	wire _w15025_ ;
	wire _w15026_ ;
	wire _w15027_ ;
	wire _w15028_ ;
	wire _w15029_ ;
	wire _w15030_ ;
	wire _w15031_ ;
	wire _w15032_ ;
	wire _w15033_ ;
	wire _w15034_ ;
	wire _w15035_ ;
	wire _w15036_ ;
	wire _w15037_ ;
	wire _w15038_ ;
	wire _w15039_ ;
	wire _w15040_ ;
	wire _w15041_ ;
	wire _w15042_ ;
	wire _w15043_ ;
	wire _w15044_ ;
	wire _w15045_ ;
	wire _w15046_ ;
	wire _w15047_ ;
	wire _w15048_ ;
	wire _w15049_ ;
	wire _w15050_ ;
	wire _w15051_ ;
	wire _w15052_ ;
	wire _w15053_ ;
	wire _w15054_ ;
	wire _w15055_ ;
	wire _w15056_ ;
	wire _w15057_ ;
	wire _w15058_ ;
	wire _w15059_ ;
	wire _w15060_ ;
	wire _w15061_ ;
	wire _w15062_ ;
	wire _w15063_ ;
	wire _w15064_ ;
	wire _w15065_ ;
	wire _w15066_ ;
	wire _w15067_ ;
	wire _w15068_ ;
	wire _w15069_ ;
	wire _w15070_ ;
	wire _w15071_ ;
	wire _w15072_ ;
	wire _w15073_ ;
	wire _w15074_ ;
	wire _w15075_ ;
	wire _w15076_ ;
	wire _w15077_ ;
	wire _w15078_ ;
	wire _w15079_ ;
	wire _w15080_ ;
	wire _w15081_ ;
	wire _w15082_ ;
	wire _w15083_ ;
	wire _w15084_ ;
	wire _w15085_ ;
	wire _w15086_ ;
	wire _w15087_ ;
	wire _w15088_ ;
	wire _w15089_ ;
	wire _w15090_ ;
	wire _w15091_ ;
	wire _w15092_ ;
	wire _w15093_ ;
	wire _w15094_ ;
	wire _w15095_ ;
	wire _w15096_ ;
	wire _w15097_ ;
	wire _w15098_ ;
	wire _w15099_ ;
	wire _w15100_ ;
	wire _w15101_ ;
	wire _w15102_ ;
	wire _w15103_ ;
	wire _w15104_ ;
	wire _w15105_ ;
	wire _w15106_ ;
	wire _w15107_ ;
	wire _w15108_ ;
	wire _w15109_ ;
	wire _w15110_ ;
	wire _w15111_ ;
	wire _w15112_ ;
	wire _w15113_ ;
	wire _w15114_ ;
	wire _w15115_ ;
	wire _w15116_ ;
	wire _w15117_ ;
	wire _w15118_ ;
	wire _w15119_ ;
	wire _w15120_ ;
	wire _w15121_ ;
	wire _w15122_ ;
	wire _w15123_ ;
	wire _w15124_ ;
	wire _w15125_ ;
	wire _w15126_ ;
	wire _w15127_ ;
	wire _w15128_ ;
	wire _w15129_ ;
	wire _w15130_ ;
	wire _w15131_ ;
	wire _w15132_ ;
	wire _w15133_ ;
	wire _w15134_ ;
	wire _w15135_ ;
	wire _w15136_ ;
	wire _w15137_ ;
	wire _w15138_ ;
	wire _w15139_ ;
	wire _w15140_ ;
	wire _w15141_ ;
	wire _w15142_ ;
	wire _w15143_ ;
	wire _w15144_ ;
	wire _w15145_ ;
	wire _w15146_ ;
	wire _w15147_ ;
	wire _w15148_ ;
	wire _w15149_ ;
	wire _w15150_ ;
	wire _w15151_ ;
	wire _w15152_ ;
	wire _w15153_ ;
	wire _w15154_ ;
	wire _w15155_ ;
	wire _w15156_ ;
	wire _w15157_ ;
	wire _w15158_ ;
	wire _w15159_ ;
	wire _w15160_ ;
	wire _w15161_ ;
	wire _w15162_ ;
	wire _w15163_ ;
	wire _w15164_ ;
	wire _w15165_ ;
	wire _w15166_ ;
	wire _w15167_ ;
	wire _w15168_ ;
	wire _w15169_ ;
	wire _w15170_ ;
	wire _w15171_ ;
	wire _w15172_ ;
	wire _w15173_ ;
	wire _w15174_ ;
	wire _w15175_ ;
	wire _w15176_ ;
	wire _w15177_ ;
	wire _w15178_ ;
	wire _w15179_ ;
	wire _w15180_ ;
	wire _w15181_ ;
	wire _w15182_ ;
	wire _w15183_ ;
	wire _w15184_ ;
	wire _w15185_ ;
	wire _w15186_ ;
	wire _w15187_ ;
	wire _w15188_ ;
	wire _w15189_ ;
	wire _w15190_ ;
	wire _w15191_ ;
	wire _w15192_ ;
	wire _w15193_ ;
	wire _w15194_ ;
	wire _w15195_ ;
	wire _w15196_ ;
	wire _w15197_ ;
	wire _w15198_ ;
	wire _w15199_ ;
	wire _w15200_ ;
	wire _w15201_ ;
	wire _w15202_ ;
	wire _w15203_ ;
	wire _w15204_ ;
	wire _w15205_ ;
	wire _w15206_ ;
	wire _w15207_ ;
	wire _w15208_ ;
	wire _w15209_ ;
	wire _w15210_ ;
	wire _w15211_ ;
	wire _w15212_ ;
	wire _w15213_ ;
	wire _w15214_ ;
	wire _w15215_ ;
	wire _w15216_ ;
	wire _w15217_ ;
	wire _w15218_ ;
	wire _w15219_ ;
	wire _w15220_ ;
	wire _w15221_ ;
	wire _w15222_ ;
	wire _w15223_ ;
	wire _w15224_ ;
	wire _w15225_ ;
	wire _w15226_ ;
	wire _w15227_ ;
	wire _w15228_ ;
	wire _w15229_ ;
	wire _w15230_ ;
	wire _w15231_ ;
	wire _w15232_ ;
	wire _w15233_ ;
	wire _w15234_ ;
	wire _w15235_ ;
	wire _w15236_ ;
	wire _w15237_ ;
	wire _w15238_ ;
	wire _w15239_ ;
	wire _w15240_ ;
	wire _w15241_ ;
	wire _w15242_ ;
	wire _w15243_ ;
	wire _w15244_ ;
	wire _w15245_ ;
	wire _w15246_ ;
	wire _w15247_ ;
	wire _w15248_ ;
	wire _w15249_ ;
	wire _w15250_ ;
	wire _w15251_ ;
	wire _w15252_ ;
	wire _w15253_ ;
	wire _w15254_ ;
	wire _w15255_ ;
	wire _w15256_ ;
	wire _w15257_ ;
	wire _w15258_ ;
	wire _w15259_ ;
	wire _w15260_ ;
	wire _w15261_ ;
	wire _w15262_ ;
	wire _w15263_ ;
	wire _w15264_ ;
	wire _w15265_ ;
	wire _w15266_ ;
	wire _w15267_ ;
	wire _w15268_ ;
	wire _w15269_ ;
	wire _w15270_ ;
	wire _w15271_ ;
	wire _w15272_ ;
	wire _w15273_ ;
	wire _w15274_ ;
	wire _w15275_ ;
	wire _w15276_ ;
	wire _w15277_ ;
	wire _w15278_ ;
	wire _w15279_ ;
	wire _w15280_ ;
	wire _w15281_ ;
	wire _w15282_ ;
	wire _w15283_ ;
	wire _w15284_ ;
	wire _w15285_ ;
	wire _w15286_ ;
	wire _w15287_ ;
	wire _w15288_ ;
	wire _w15289_ ;
	wire _w15290_ ;
	wire _w15291_ ;
	wire _w15292_ ;
	wire _w15293_ ;
	wire _w15294_ ;
	wire _w15295_ ;
	wire _w15296_ ;
	wire _w15297_ ;
	wire _w15298_ ;
	wire _w15299_ ;
	wire _w15300_ ;
	wire _w15301_ ;
	wire _w15302_ ;
	wire _w15303_ ;
	wire _w15304_ ;
	wire _w15305_ ;
	wire _w15306_ ;
	wire _w15307_ ;
	wire _w15308_ ;
	wire _w15309_ ;
	wire _w15310_ ;
	wire _w15311_ ;
	wire _w15312_ ;
	wire _w15313_ ;
	wire _w15314_ ;
	wire _w15315_ ;
	wire _w15316_ ;
	wire _w15317_ ;
	wire _w15318_ ;
	wire _w15319_ ;
	wire _w15320_ ;
	wire _w15321_ ;
	wire _w15322_ ;
	wire _w15323_ ;
	wire _w15324_ ;
	wire _w15325_ ;
	wire _w15326_ ;
	wire _w15327_ ;
	wire _w15328_ ;
	wire _w15329_ ;
	wire _w15330_ ;
	wire _w15331_ ;
	wire _w15332_ ;
	wire _w15333_ ;
	wire _w15334_ ;
	wire _w15335_ ;
	wire _w15336_ ;
	wire _w15337_ ;
	wire _w15338_ ;
	wire _w15339_ ;
	wire _w15340_ ;
	wire _w15341_ ;
	wire _w15342_ ;
	wire _w15343_ ;
	wire _w15344_ ;
	wire _w15345_ ;
	wire _w15346_ ;
	wire _w15347_ ;
	wire _w15348_ ;
	wire _w15349_ ;
	wire _w15350_ ;
	wire _w15351_ ;
	wire _w15352_ ;
	wire _w15353_ ;
	wire _w15354_ ;
	wire _w15355_ ;
	wire _w15356_ ;
	wire _w15357_ ;
	wire _w15358_ ;
	wire _w15359_ ;
	wire _w15360_ ;
	wire _w15361_ ;
	wire _w15362_ ;
	wire _w15363_ ;
	wire _w15364_ ;
	wire _w15365_ ;
	wire _w15366_ ;
	wire _w15367_ ;
	wire _w15368_ ;
	wire _w15369_ ;
	wire _w15370_ ;
	wire _w15371_ ;
	wire _w15372_ ;
	wire _w15373_ ;
	wire _w15374_ ;
	wire _w15375_ ;
	wire _w15376_ ;
	wire _w15377_ ;
	wire _w15378_ ;
	wire _w15379_ ;
	wire _w15380_ ;
	wire _w15381_ ;
	wire _w15382_ ;
	wire _w15383_ ;
	wire _w15384_ ;
	wire _w15385_ ;
	wire _w15386_ ;
	wire _w15387_ ;
	wire _w15388_ ;
	wire _w15389_ ;
	wire _w15390_ ;
	wire _w15391_ ;
	wire _w15392_ ;
	wire _w15393_ ;
	wire _w15394_ ;
	wire _w15395_ ;
	wire _w15396_ ;
	wire _w15397_ ;
	wire _w15398_ ;
	wire _w15399_ ;
	wire _w15400_ ;
	wire _w15401_ ;
	wire _w15402_ ;
	wire _w15403_ ;
	wire _w15404_ ;
	wire _w15405_ ;
	wire _w15406_ ;
	wire _w15407_ ;
	wire _w15408_ ;
	wire _w15409_ ;
	wire _w15410_ ;
	wire _w15411_ ;
	wire _w15412_ ;
	wire _w15413_ ;
	wire _w15414_ ;
	wire _w15415_ ;
	wire _w15416_ ;
	wire _w15417_ ;
	wire _w15418_ ;
	wire _w15419_ ;
	wire _w15420_ ;
	wire _w15421_ ;
	wire _w15422_ ;
	wire _w15423_ ;
	wire _w15424_ ;
	wire _w15425_ ;
	wire _w15426_ ;
	wire _w15427_ ;
	wire _w15428_ ;
	wire _w15429_ ;
	wire _w15430_ ;
	wire _w15431_ ;
	wire _w15432_ ;
	wire _w15433_ ;
	wire _w15434_ ;
	wire _w15435_ ;
	wire _w15436_ ;
	wire _w15437_ ;
	wire _w15438_ ;
	wire _w15439_ ;
	wire _w15440_ ;
	wire _w15441_ ;
	wire _w15442_ ;
	wire _w15443_ ;
	wire _w15444_ ;
	wire _w15445_ ;
	wire _w15446_ ;
	wire _w15447_ ;
	wire _w15448_ ;
	wire _w15449_ ;
	wire _w15450_ ;
	wire _w15451_ ;
	wire _w15452_ ;
	wire _w15453_ ;
	wire _w15454_ ;
	wire _w15455_ ;
	wire _w15456_ ;
	wire _w15457_ ;
	wire _w15458_ ;
	wire _w15459_ ;
	wire _w15460_ ;
	wire _w15461_ ;
	wire _w15462_ ;
	wire _w15463_ ;
	wire _w15464_ ;
	wire _w15465_ ;
	wire _w15466_ ;
	wire _w15467_ ;
	wire _w15468_ ;
	wire _w15469_ ;
	wire _w15470_ ;
	wire _w15471_ ;
	wire _w15472_ ;
	wire _w15473_ ;
	wire _w15474_ ;
	wire _w15475_ ;
	wire _w15476_ ;
	wire _w15477_ ;
	wire _w15478_ ;
	wire _w15479_ ;
	wire _w15480_ ;
	wire _w15481_ ;
	wire _w15482_ ;
	wire _w15483_ ;
	wire _w15484_ ;
	wire _w15485_ ;
	wire _w15486_ ;
	wire _w15487_ ;
	wire _w15488_ ;
	wire _w15489_ ;
	wire _w15490_ ;
	wire _w15491_ ;
	wire _w15492_ ;
	wire _w15493_ ;
	wire _w15494_ ;
	wire _w15495_ ;
	wire _w15496_ ;
	wire _w15497_ ;
	wire _w15498_ ;
	wire _w15499_ ;
	wire _w15500_ ;
	wire _w15501_ ;
	wire _w15502_ ;
	wire _w15503_ ;
	wire _w15504_ ;
	wire _w15505_ ;
	wire _w15506_ ;
	wire _w15507_ ;
	wire _w15508_ ;
	wire _w15509_ ;
	wire _w15510_ ;
	wire _w15511_ ;
	wire _w15512_ ;
	wire _w15513_ ;
	wire _w15514_ ;
	wire _w15515_ ;
	wire _w15516_ ;
	wire _w15517_ ;
	wire _w15518_ ;
	wire _w15519_ ;
	wire _w15520_ ;
	wire _w15521_ ;
	wire _w15522_ ;
	wire _w15523_ ;
	wire _w15524_ ;
	wire _w15525_ ;
	wire _w15526_ ;
	wire _w15527_ ;
	wire _w15528_ ;
	wire _w15529_ ;
	wire _w15530_ ;
	wire _w15531_ ;
	wire _w15532_ ;
	wire _w15533_ ;
	wire _w15534_ ;
	wire _w15535_ ;
	wire _w15536_ ;
	wire _w15537_ ;
	wire _w15538_ ;
	wire _w15539_ ;
	wire _w15540_ ;
	wire _w15541_ ;
	wire _w15542_ ;
	wire _w15543_ ;
	wire _w15544_ ;
	wire _w15545_ ;
	wire _w15546_ ;
	wire _w15547_ ;
	wire _w15548_ ;
	wire _w15549_ ;
	wire _w15550_ ;
	wire _w15551_ ;
	wire _w15552_ ;
	wire _w15553_ ;
	wire _w15554_ ;
	wire _w15555_ ;
	wire _w15556_ ;
	wire _w15557_ ;
	wire _w15558_ ;
	wire _w15559_ ;
	wire _w15560_ ;
	wire _w15561_ ;
	wire _w15562_ ;
	wire _w15563_ ;
	wire _w15564_ ;
	wire _w15565_ ;
	wire _w15566_ ;
	wire _w15567_ ;
	wire _w15568_ ;
	wire _w15569_ ;
	wire _w15570_ ;
	wire _w15571_ ;
	wire _w15572_ ;
	wire _w15573_ ;
	wire _w15574_ ;
	wire _w15575_ ;
	wire _w15576_ ;
	wire _w15577_ ;
	wire _w15578_ ;
	wire _w15579_ ;
	wire _w15580_ ;
	wire _w15581_ ;
	wire _w15582_ ;
	wire _w15583_ ;
	wire _w15584_ ;
	wire _w15585_ ;
	wire _w15586_ ;
	wire _w15587_ ;
	wire _w15588_ ;
	wire _w15589_ ;
	wire _w15590_ ;
	wire _w15591_ ;
	wire _w15592_ ;
	wire _w15593_ ;
	wire _w15594_ ;
	wire _w15595_ ;
	wire _w15596_ ;
	wire _w15597_ ;
	wire _w15598_ ;
	wire _w15599_ ;
	wire _w15600_ ;
	wire _w15601_ ;
	wire _w15602_ ;
	wire _w15603_ ;
	wire _w15604_ ;
	wire _w15605_ ;
	wire _w15606_ ;
	wire _w15607_ ;
	wire _w15608_ ;
	wire _w15609_ ;
	wire _w15610_ ;
	wire _w15611_ ;
	wire _w15612_ ;
	wire _w15613_ ;
	wire _w15614_ ;
	wire _w15615_ ;
	wire _w15616_ ;
	wire _w15617_ ;
	wire _w15618_ ;
	wire _w15619_ ;
	wire _w15620_ ;
	wire _w15621_ ;
	wire _w15622_ ;
	wire _w15623_ ;
	wire _w15624_ ;
	wire _w15625_ ;
	wire _w15626_ ;
	wire _w15627_ ;
	wire _w15628_ ;
	wire _w15629_ ;
	wire _w15630_ ;
	wire _w15631_ ;
	wire _w15632_ ;
	wire _w15633_ ;
	wire _w15634_ ;
	wire _w15635_ ;
	wire _w15636_ ;
	wire _w15637_ ;
	wire _w15638_ ;
	wire _w15639_ ;
	wire _w15640_ ;
	wire _w15641_ ;
	wire _w15642_ ;
	wire _w15643_ ;
	wire _w15644_ ;
	wire _w15645_ ;
	wire _w15646_ ;
	wire _w15647_ ;
	wire _w15648_ ;
	wire _w15649_ ;
	wire _w15650_ ;
	wire _w15651_ ;
	wire _w15652_ ;
	wire _w15653_ ;
	wire _w15654_ ;
	wire _w15655_ ;
	wire _w15656_ ;
	wire _w15657_ ;
	wire _w15658_ ;
	wire _w15659_ ;
	wire _w15660_ ;
	wire _w15661_ ;
	wire _w15662_ ;
	wire _w15663_ ;
	wire _w15664_ ;
	wire _w15665_ ;
	wire _w15666_ ;
	wire _w15667_ ;
	wire _w15668_ ;
	wire _w15669_ ;
	wire _w15670_ ;
	wire _w15671_ ;
	wire _w15672_ ;
	wire _w15673_ ;
	wire _w15674_ ;
	wire _w15675_ ;
	wire _w15676_ ;
	wire _w15677_ ;
	wire _w15678_ ;
	wire _w15679_ ;
	wire _w15680_ ;
	wire _w15681_ ;
	wire _w15682_ ;
	wire _w15683_ ;
	wire _w15684_ ;
	wire _w15685_ ;
	wire _w15686_ ;
	wire _w15687_ ;
	wire _w15688_ ;
	wire _w15689_ ;
	wire _w15690_ ;
	wire _w15691_ ;
	wire _w15692_ ;
	wire _w15693_ ;
	wire _w15694_ ;
	wire _w15695_ ;
	wire _w15696_ ;
	wire _w15697_ ;
	wire _w15698_ ;
	wire _w15699_ ;
	wire _w15700_ ;
	wire _w15701_ ;
	wire _w15702_ ;
	wire _w15703_ ;
	wire _w15704_ ;
	wire _w15705_ ;
	wire _w15706_ ;
	wire _w15707_ ;
	wire _w15708_ ;
	wire _w15709_ ;
	wire _w15710_ ;
	wire _w15711_ ;
	wire _w15712_ ;
	wire _w15713_ ;
	wire _w15714_ ;
	wire _w15715_ ;
	wire _w15716_ ;
	wire _w15717_ ;
	wire _w15718_ ;
	wire _w15719_ ;
	wire _w15720_ ;
	wire _w15721_ ;
	wire _w15722_ ;
	wire _w15723_ ;
	wire _w15724_ ;
	wire _w15725_ ;
	wire _w15726_ ;
	wire _w15727_ ;
	wire _w15728_ ;
	wire _w15729_ ;
	wire _w15730_ ;
	wire _w15731_ ;
	wire _w15732_ ;
	wire _w15733_ ;
	wire _w15734_ ;
	wire _w15735_ ;
	wire _w15736_ ;
	wire _w15737_ ;
	wire _w15738_ ;
	wire _w15739_ ;
	wire _w15740_ ;
	wire _w15741_ ;
	wire _w15742_ ;
	wire _w15743_ ;
	wire _w15744_ ;
	wire _w15745_ ;
	wire _w15746_ ;
	wire _w15747_ ;
	wire _w15748_ ;
	wire _w15749_ ;
	wire _w15750_ ;
	wire _w15751_ ;
	wire _w15752_ ;
	wire _w15753_ ;
	wire _w15754_ ;
	wire _w15755_ ;
	wire _w15756_ ;
	wire _w15757_ ;
	wire _w15758_ ;
	wire _w15759_ ;
	wire _w15760_ ;
	wire _w15761_ ;
	wire _w15762_ ;
	wire _w15763_ ;
	wire _w15764_ ;
	wire _w15765_ ;
	wire _w15766_ ;
	wire _w15767_ ;
	wire _w15768_ ;
	wire _w15769_ ;
	wire _w15770_ ;
	wire _w15771_ ;
	wire _w15772_ ;
	wire _w15773_ ;
	wire _w15774_ ;
	wire _w15775_ ;
	wire _w15776_ ;
	wire _w15777_ ;
	wire _w15778_ ;
	wire _w15779_ ;
	wire _w15780_ ;
	wire _w15781_ ;
	wire _w15782_ ;
	wire _w15783_ ;
	wire _w15784_ ;
	wire _w15785_ ;
	wire _w15786_ ;
	wire _w15787_ ;
	wire _w15788_ ;
	wire _w15789_ ;
	wire _w15790_ ;
	wire _w15791_ ;
	wire _w15792_ ;
	wire _w15793_ ;
	wire _w15794_ ;
	wire _w15795_ ;
	wire _w15796_ ;
	wire _w15797_ ;
	wire _w15798_ ;
	wire _w15799_ ;
	wire _w15800_ ;
	wire _w15801_ ;
	wire _w15802_ ;
	wire _w15803_ ;
	wire _w15804_ ;
	wire _w15805_ ;
	wire _w15806_ ;
	wire _w15807_ ;
	wire _w15808_ ;
	wire _w15809_ ;
	wire _w15810_ ;
	wire _w15811_ ;
	wire _w15812_ ;
	wire _w15813_ ;
	wire _w15814_ ;
	wire _w15815_ ;
	wire _w15816_ ;
	wire _w15817_ ;
	wire _w15818_ ;
	wire _w15819_ ;
	wire _w15820_ ;
	wire _w15821_ ;
	wire _w15822_ ;
	wire _w15823_ ;
	wire _w15824_ ;
	wire _w15825_ ;
	wire _w15826_ ;
	wire _w15827_ ;
	wire _w15828_ ;
	wire _w15829_ ;
	wire _w15830_ ;
	wire _w15831_ ;
	wire _w15832_ ;
	wire _w15833_ ;
	wire _w15834_ ;
	wire _w15835_ ;
	wire _w15836_ ;
	wire _w15837_ ;
	wire _w15838_ ;
	wire _w15839_ ;
	wire _w15840_ ;
	wire _w15841_ ;
	wire _w15842_ ;
	wire _w15843_ ;
	wire _w15844_ ;
	wire _w15845_ ;
	wire _w15846_ ;
	wire _w15847_ ;
	wire _w15848_ ;
	wire _w15849_ ;
	wire _w15850_ ;
	wire _w15851_ ;
	wire _w15852_ ;
	wire _w15853_ ;
	wire _w15854_ ;
	wire _w15855_ ;
	wire _w15856_ ;
	wire _w15857_ ;
	wire _w15858_ ;
	wire _w15859_ ;
	wire _w15860_ ;
	wire _w15861_ ;
	wire _w15862_ ;
	wire _w15863_ ;
	wire _w15864_ ;
	wire _w15865_ ;
	wire _w15866_ ;
	wire _w15867_ ;
	wire _w15868_ ;
	wire _w15869_ ;
	wire _w15870_ ;
	wire _w15871_ ;
	wire _w15872_ ;
	wire _w15873_ ;
	wire _w15874_ ;
	wire _w15875_ ;
	wire _w15876_ ;
	wire _w15877_ ;
	wire _w15878_ ;
	wire _w15879_ ;
	wire _w15880_ ;
	wire _w15881_ ;
	wire _w15882_ ;
	wire _w15883_ ;
	wire _w15884_ ;
	wire _w15885_ ;
	wire _w15886_ ;
	wire _w15887_ ;
	wire _w15888_ ;
	wire _w15889_ ;
	wire _w15890_ ;
	wire _w15891_ ;
	wire _w15892_ ;
	wire _w15893_ ;
	wire _w15894_ ;
	wire _w15895_ ;
	wire _w15896_ ;
	wire _w15897_ ;
	wire _w15898_ ;
	wire _w15899_ ;
	wire _w15900_ ;
	wire _w15901_ ;
	wire _w15902_ ;
	wire _w15903_ ;
	wire _w15904_ ;
	wire _w15905_ ;
	wire _w15906_ ;
	wire _w15907_ ;
	wire _w15908_ ;
	wire _w15909_ ;
	wire _w15910_ ;
	wire _w15911_ ;
	wire _w15912_ ;
	wire _w15913_ ;
	wire _w15914_ ;
	wire _w15915_ ;
	wire _w15916_ ;
	wire _w15917_ ;
	wire _w15918_ ;
	wire _w15919_ ;
	wire _w15920_ ;
	wire _w15921_ ;
	wire _w15922_ ;
	wire _w15923_ ;
	wire _w15924_ ;
	wire _w15925_ ;
	wire _w15926_ ;
	wire _w15927_ ;
	wire _w15928_ ;
	wire _w15929_ ;
	wire _w15930_ ;
	wire _w15931_ ;
	wire _w15932_ ;
	wire _w15933_ ;
	wire _w15934_ ;
	wire _w15935_ ;
	wire _w15936_ ;
	wire _w15937_ ;
	wire _w15938_ ;
	wire _w15939_ ;
	wire _w15940_ ;
	wire _w15941_ ;
	wire _w15942_ ;
	wire _w15943_ ;
	wire _w15944_ ;
	wire _w15945_ ;
	wire _w15946_ ;
	wire _w15947_ ;
	wire _w15948_ ;
	wire _w15949_ ;
	wire _w15950_ ;
	wire _w15951_ ;
	wire _w15952_ ;
	wire _w15953_ ;
	wire _w15954_ ;
	wire _w15955_ ;
	wire _w15956_ ;
	wire _w15957_ ;
	wire _w15958_ ;
	wire _w15959_ ;
	wire _w15960_ ;
	wire _w15961_ ;
	wire _w15962_ ;
	wire _w15963_ ;
	wire _w15964_ ;
	wire _w15965_ ;
	wire _w15966_ ;
	wire _w15967_ ;
	wire _w15968_ ;
	wire _w15969_ ;
	wire _w15970_ ;
	wire _w15971_ ;
	wire _w15972_ ;
	wire _w15973_ ;
	wire _w15974_ ;
	wire _w15975_ ;
	wire _w15976_ ;
	wire _w15977_ ;
	wire _w15978_ ;
	wire _w15979_ ;
	wire _w15980_ ;
	wire _w15981_ ;
	wire _w15982_ ;
	wire _w15983_ ;
	wire _w15984_ ;
	wire _w15985_ ;
	wire _w15986_ ;
	wire _w15987_ ;
	wire _w15988_ ;
	wire _w15989_ ;
	wire _w15990_ ;
	wire _w15991_ ;
	wire _w15992_ ;
	wire _w15993_ ;
	wire _w15994_ ;
	wire _w15995_ ;
	wire _w15996_ ;
	wire _w15997_ ;
	wire _w15998_ ;
	wire _w15999_ ;
	wire _w16000_ ;
	wire _w16001_ ;
	wire _w16002_ ;
	wire _w16003_ ;
	wire _w16004_ ;
	wire _w16005_ ;
	wire _w16006_ ;
	wire _w16007_ ;
	wire _w16008_ ;
	wire _w16009_ ;
	wire _w16010_ ;
	wire _w16011_ ;
	wire _w16012_ ;
	wire _w16013_ ;
	wire _w16014_ ;
	wire _w16015_ ;
	wire _w16016_ ;
	wire _w16017_ ;
	wire _w16018_ ;
	wire _w16019_ ;
	wire _w16020_ ;
	wire _w16021_ ;
	wire _w16022_ ;
	wire _w16023_ ;
	wire _w16024_ ;
	wire _w16025_ ;
	wire _w16026_ ;
	wire _w16027_ ;
	wire _w16028_ ;
	wire _w16029_ ;
	wire _w16030_ ;
	wire _w16031_ ;
	wire _w16032_ ;
	wire _w16033_ ;
	wire _w16034_ ;
	wire _w16035_ ;
	wire _w16036_ ;
	wire _w16037_ ;
	wire _w16038_ ;
	wire _w16039_ ;
	wire _w16040_ ;
	wire _w16041_ ;
	wire _w16042_ ;
	wire _w16043_ ;
	wire _w16044_ ;
	wire _w16045_ ;
	wire _w16046_ ;
	wire _w16047_ ;
	wire _w16048_ ;
	wire _w16049_ ;
	wire _w16050_ ;
	wire _w16051_ ;
	wire _w16052_ ;
	wire _w16053_ ;
	wire _w16054_ ;
	wire _w16055_ ;
	wire _w16056_ ;
	wire _w16057_ ;
	wire _w16058_ ;
	wire _w16059_ ;
	wire _w16060_ ;
	wire _w16061_ ;
	wire _w16062_ ;
	wire _w16063_ ;
	wire _w16064_ ;
	wire _w16065_ ;
	wire _w16066_ ;
	wire _w16067_ ;
	wire _w16068_ ;
	wire _w16069_ ;
	wire _w16070_ ;
	wire _w16071_ ;
	wire _w16072_ ;
	wire _w16073_ ;
	wire _w16074_ ;
	wire _w16075_ ;
	wire _w16076_ ;
	wire _w16077_ ;
	wire _w16078_ ;
	wire _w16079_ ;
	wire _w16080_ ;
	wire _w16081_ ;
	wire _w16082_ ;
	wire _w16083_ ;
	wire _w16084_ ;
	wire _w16085_ ;
	wire _w16086_ ;
	wire _w16087_ ;
	wire _w16088_ ;
	wire _w16089_ ;
	wire _w16090_ ;
	wire _w16091_ ;
	wire _w16092_ ;
	wire _w16093_ ;
	wire _w16094_ ;
	wire _w16095_ ;
	wire _w16096_ ;
	wire _w16097_ ;
	wire _w16098_ ;
	wire _w16099_ ;
	wire _w16100_ ;
	wire _w16101_ ;
	wire _w16102_ ;
	wire _w16103_ ;
	wire _w16104_ ;
	wire _w16105_ ;
	wire _w16106_ ;
	wire _w16107_ ;
	wire _w16108_ ;
	wire _w16109_ ;
	wire _w16110_ ;
	wire _w16111_ ;
	wire _w16112_ ;
	wire _w16113_ ;
	wire _w16114_ ;
	wire _w16115_ ;
	wire _w16116_ ;
	wire _w16117_ ;
	wire _w16118_ ;
	wire _w16119_ ;
	wire _w16120_ ;
	wire _w16121_ ;
	wire _w16122_ ;
	wire _w16123_ ;
	wire _w16124_ ;
	wire _w16125_ ;
	wire _w16126_ ;
	wire _w16127_ ;
	wire _w16128_ ;
	wire _w16129_ ;
	wire _w16130_ ;
	wire _w16131_ ;
	wire _w16132_ ;
	wire _w16133_ ;
	wire _w16134_ ;
	wire _w16135_ ;
	wire _w16136_ ;
	wire _w16137_ ;
	wire _w16138_ ;
	wire _w16139_ ;
	wire _w16140_ ;
	wire _w16141_ ;
	wire _w16142_ ;
	wire _w16143_ ;
	wire _w16144_ ;
	wire _w16145_ ;
	wire _w16146_ ;
	wire _w16147_ ;
	wire _w16148_ ;
	wire _w16149_ ;
	wire _w16150_ ;
	wire _w16151_ ;
	wire _w16152_ ;
	wire _w16153_ ;
	wire _w16154_ ;
	wire _w16155_ ;
	wire _w16156_ ;
	wire _w16157_ ;
	wire _w16158_ ;
	wire _w16159_ ;
	wire _w16160_ ;
	wire _w16161_ ;
	wire _w16162_ ;
	wire _w16163_ ;
	wire _w16164_ ;
	wire _w16165_ ;
	wire _w16166_ ;
	wire _w16167_ ;
	wire _w16168_ ;
	wire _w16169_ ;
	wire _w16170_ ;
	wire _w16171_ ;
	wire _w16172_ ;
	wire _w16173_ ;
	wire _w16174_ ;
	wire _w16175_ ;
	wire _w16176_ ;
	wire _w16177_ ;
	wire _w16178_ ;
	wire _w16179_ ;
	wire _w16180_ ;
	wire _w16181_ ;
	wire _w16182_ ;
	wire _w16183_ ;
	wire _w16184_ ;
	wire _w16185_ ;
	wire _w16186_ ;
	wire _w16187_ ;
	wire _w16188_ ;
	wire _w16189_ ;
	wire _w16190_ ;
	wire _w16191_ ;
	wire _w16192_ ;
	wire _w16193_ ;
	wire _w16194_ ;
	wire _w16195_ ;
	wire _w16196_ ;
	wire _w16197_ ;
	wire _w16198_ ;
	wire _w16199_ ;
	wire _w16200_ ;
	wire _w16201_ ;
	wire _w16202_ ;
	wire _w16203_ ;
	wire _w16204_ ;
	wire _w16205_ ;
	wire _w16206_ ;
	wire _w16207_ ;
	wire _w16208_ ;
	wire _w16209_ ;
	wire _w16210_ ;
	wire _w16211_ ;
	wire _w16212_ ;
	wire _w16213_ ;
	wire _w16214_ ;
	wire _w16215_ ;
	wire _w16216_ ;
	wire _w16217_ ;
	wire _w16218_ ;
	wire _w16219_ ;
	wire _w16220_ ;
	wire _w16221_ ;
	wire _w16222_ ;
	wire _w16223_ ;
	wire _w16224_ ;
	wire _w16225_ ;
	wire _w16226_ ;
	wire _w16227_ ;
	wire _w16228_ ;
	wire _w16229_ ;
	wire _w16230_ ;
	wire _w16231_ ;
	wire _w16232_ ;
	wire _w16233_ ;
	wire _w16234_ ;
	wire _w16235_ ;
	wire _w16236_ ;
	wire _w16237_ ;
	wire _w16238_ ;
	wire _w16239_ ;
	wire _w16240_ ;
	wire _w16241_ ;
	wire _w16242_ ;
	wire _w16243_ ;
	wire _w16244_ ;
	wire _w16245_ ;
	wire _w16246_ ;
	wire _w16247_ ;
	wire _w16248_ ;
	wire _w16249_ ;
	wire _w16250_ ;
	wire _w16251_ ;
	wire _w16252_ ;
	wire _w16253_ ;
	wire _w16254_ ;
	wire _w16255_ ;
	wire _w16256_ ;
	wire _w16257_ ;
	wire _w16258_ ;
	wire _w16259_ ;
	wire _w16260_ ;
	wire _w16261_ ;
	wire _w16262_ ;
	wire _w16263_ ;
	wire _w16264_ ;
	wire _w16265_ ;
	wire _w16266_ ;
	wire _w16267_ ;
	wire _w16268_ ;
	wire _w16269_ ;
	wire _w16270_ ;
	wire _w16271_ ;
	wire _w16272_ ;
	wire _w16273_ ;
	wire _w16274_ ;
	wire _w16275_ ;
	wire _w16276_ ;
	wire _w16277_ ;
	wire _w16278_ ;
	wire _w16279_ ;
	wire _w16280_ ;
	wire _w16281_ ;
	wire _w16282_ ;
	wire _w16283_ ;
	wire _w16284_ ;
	wire _w16285_ ;
	wire _w16286_ ;
	wire _w16287_ ;
	wire _w16288_ ;
	wire _w16289_ ;
	wire _w16290_ ;
	wire _w16291_ ;
	wire _w16292_ ;
	wire _w16293_ ;
	wire _w16294_ ;
	wire _w16295_ ;
	wire _w16296_ ;
	wire _w16297_ ;
	wire _w16298_ ;
	wire _w16299_ ;
	wire _w16300_ ;
	wire _w16301_ ;
	wire _w16302_ ;
	wire _w16303_ ;
	wire _w16304_ ;
	wire _w16305_ ;
	wire _w16306_ ;
	wire _w16307_ ;
	wire _w16308_ ;
	wire _w16309_ ;
	wire _w16310_ ;
	wire _w16311_ ;
	wire _w16312_ ;
	wire _w16313_ ;
	wire _w16314_ ;
	wire _w16315_ ;
	wire _w16316_ ;
	wire _w16317_ ;
	wire _w16318_ ;
	wire _w16319_ ;
	wire _w16320_ ;
	wire _w16321_ ;
	wire _w16322_ ;
	wire _w16323_ ;
	wire _w16324_ ;
	wire _w16325_ ;
	wire _w16326_ ;
	wire _w16327_ ;
	wire _w16328_ ;
	wire _w16329_ ;
	wire _w16330_ ;
	wire _w16331_ ;
	wire _w16332_ ;
	wire _w16333_ ;
	wire _w16334_ ;
	wire _w16335_ ;
	wire _w16336_ ;
	wire _w16337_ ;
	wire _w16338_ ;
	wire _w16339_ ;
	wire _w16340_ ;
	wire _w16341_ ;
	wire _w16342_ ;
	wire _w16343_ ;
	wire _w16344_ ;
	wire _w16345_ ;
	wire _w16346_ ;
	wire _w16347_ ;
	wire _w16348_ ;
	wire _w16349_ ;
	wire _w16350_ ;
	wire _w16351_ ;
	wire _w16352_ ;
	wire _w16353_ ;
	wire _w16354_ ;
	wire _w16355_ ;
	wire _w16356_ ;
	wire _w16357_ ;
	wire _w16358_ ;
	wire _w16359_ ;
	wire _w16360_ ;
	wire _w16361_ ;
	wire _w16362_ ;
	wire _w16363_ ;
	wire _w16364_ ;
	wire _w16365_ ;
	wire _w16366_ ;
	wire _w16367_ ;
	wire _w16368_ ;
	wire _w16369_ ;
	wire _w16370_ ;
	wire _w16371_ ;
	wire _w16372_ ;
	wire _w16373_ ;
	wire _w16374_ ;
	wire _w16375_ ;
	wire _w16376_ ;
	wire _w16377_ ;
	wire _w16378_ ;
	wire _w16379_ ;
	wire _w16380_ ;
	wire _w16381_ ;
	wire _w16382_ ;
	wire _w16383_ ;
	wire _w16384_ ;
	wire _w16385_ ;
	wire _w16386_ ;
	wire _w16387_ ;
	wire _w16388_ ;
	wire _w16389_ ;
	wire _w16390_ ;
	wire _w16391_ ;
	wire _w16392_ ;
	wire _w16393_ ;
	wire _w16394_ ;
	wire _w16395_ ;
	wire _w16396_ ;
	wire _w16397_ ;
	wire _w16398_ ;
	wire _w16399_ ;
	wire _w16400_ ;
	wire _w16401_ ;
	wire _w16402_ ;
	wire _w16403_ ;
	wire _w16404_ ;
	wire _w16405_ ;
	wire _w16406_ ;
	wire _w16407_ ;
	wire _w16408_ ;
	wire _w16409_ ;
	wire _w16410_ ;
	wire _w16411_ ;
	wire _w16412_ ;
	wire _w16413_ ;
	wire _w16414_ ;
	wire _w16415_ ;
	wire _w16416_ ;
	wire _w16417_ ;
	wire _w16418_ ;
	wire _w16419_ ;
	wire _w16420_ ;
	wire _w16421_ ;
	wire _w16422_ ;
	wire _w16423_ ;
	wire _w16424_ ;
	wire _w16425_ ;
	wire _w16426_ ;
	wire _w16427_ ;
	wire _w16428_ ;
	wire _w16429_ ;
	wire _w16430_ ;
	wire _w16431_ ;
	wire _w16432_ ;
	wire _w16433_ ;
	wire _w16434_ ;
	wire _w16435_ ;
	wire _w16436_ ;
	wire _w16437_ ;
	wire _w16438_ ;
	wire _w16439_ ;
	wire _w16440_ ;
	wire _w16441_ ;
	wire _w16442_ ;
	wire _w16443_ ;
	wire _w16444_ ;
	wire _w16445_ ;
	wire _w16446_ ;
	wire _w16447_ ;
	wire _w16448_ ;
	wire _w16449_ ;
	wire _w16450_ ;
	wire _w16451_ ;
	wire _w16452_ ;
	wire _w16453_ ;
	wire _w16454_ ;
	wire _w16455_ ;
	wire _w16456_ ;
	wire _w16457_ ;
	wire _w16458_ ;
	wire _w16459_ ;
	wire _w16460_ ;
	wire _w16461_ ;
	wire _w16462_ ;
	wire _w16463_ ;
	wire _w16464_ ;
	wire _w16465_ ;
	wire _w16466_ ;
	wire _w16467_ ;
	wire _w16468_ ;
	wire _w16469_ ;
	wire _w16470_ ;
	wire _w16471_ ;
	wire _w16472_ ;
	wire _w16473_ ;
	wire _w16474_ ;
	wire _w16475_ ;
	wire _w16476_ ;
	wire _w16477_ ;
	wire _w16478_ ;
	wire _w16479_ ;
	wire _w16480_ ;
	wire _w16481_ ;
	wire _w16482_ ;
	wire _w16483_ ;
	wire _w16484_ ;
	wire _w16485_ ;
	wire _w16486_ ;
	wire _w16487_ ;
	wire _w16488_ ;
	wire _w16489_ ;
	wire _w16490_ ;
	wire _w16491_ ;
	wire _w16492_ ;
	wire _w16493_ ;
	wire _w16494_ ;
	wire _w16495_ ;
	wire _w16496_ ;
	wire _w16497_ ;
	wire _w16498_ ;
	wire _w16499_ ;
	wire _w16500_ ;
	wire _w16501_ ;
	wire _w16502_ ;
	wire _w16503_ ;
	wire _w16504_ ;
	wire _w16505_ ;
	wire _w16506_ ;
	wire _w16507_ ;
	wire _w16508_ ;
	wire _w16509_ ;
	wire _w16510_ ;
	wire _w16511_ ;
	wire _w16512_ ;
	wire _w16513_ ;
	wire _w16514_ ;
	wire _w16515_ ;
	wire _w16516_ ;
	wire _w16517_ ;
	wire _w16518_ ;
	wire _w16519_ ;
	wire _w16520_ ;
	wire _w16521_ ;
	wire _w16522_ ;
	wire _w16523_ ;
	wire _w16524_ ;
	wire _w16525_ ;
	wire _w16526_ ;
	wire _w16527_ ;
	wire _w16528_ ;
	wire _w16529_ ;
	wire _w16530_ ;
	wire _w16531_ ;
	wire _w16532_ ;
	wire _w16533_ ;
	wire _w16534_ ;
	wire _w16535_ ;
	wire _w16536_ ;
	wire _w16537_ ;
	wire _w16538_ ;
	wire _w16539_ ;
	wire _w16540_ ;
	wire _w16541_ ;
	wire _w16542_ ;
	wire _w16543_ ;
	wire _w16544_ ;
	wire _w16545_ ;
	wire _w16546_ ;
	wire _w16547_ ;
	wire _w16548_ ;
	wire _w16549_ ;
	wire _w16550_ ;
	wire _w16551_ ;
	wire _w16552_ ;
	wire _w16553_ ;
	wire _w16554_ ;
	wire _w16555_ ;
	wire _w16556_ ;
	wire _w16557_ ;
	wire _w16558_ ;
	wire _w16559_ ;
	wire _w16560_ ;
	wire _w16561_ ;
	wire _w16562_ ;
	wire _w16563_ ;
	wire _w16564_ ;
	wire _w16565_ ;
	wire _w16566_ ;
	wire _w16567_ ;
	wire _w16568_ ;
	wire _w16569_ ;
	wire _w16570_ ;
	wire _w16571_ ;
	wire _w16572_ ;
	wire _w16573_ ;
	wire _w16574_ ;
	wire _w16575_ ;
	wire _w16576_ ;
	wire _w16577_ ;
	wire _w16578_ ;
	wire _w16579_ ;
	wire _w16580_ ;
	wire _w16581_ ;
	wire _w16582_ ;
	wire _w16583_ ;
	wire _w16584_ ;
	wire _w16585_ ;
	wire _w16586_ ;
	wire _w16587_ ;
	wire _w16588_ ;
	wire _w16589_ ;
	wire _w16590_ ;
	wire _w16591_ ;
	wire _w16592_ ;
	wire _w16593_ ;
	wire _w16594_ ;
	wire _w16595_ ;
	wire _w16596_ ;
	wire _w16597_ ;
	wire _w16598_ ;
	wire _w16599_ ;
	wire _w16600_ ;
	wire _w16601_ ;
	wire _w16602_ ;
	wire _w16603_ ;
	wire _w16604_ ;
	wire _w16605_ ;
	wire _w16606_ ;
	wire _w16607_ ;
	wire _w16608_ ;
	wire _w16609_ ;
	wire _w16610_ ;
	wire _w16611_ ;
	wire _w16612_ ;
	wire _w16613_ ;
	wire _w16614_ ;
	wire _w16615_ ;
	wire _w16616_ ;
	wire _w16617_ ;
	wire _w16618_ ;
	wire _w16619_ ;
	wire _w16620_ ;
	wire _w16621_ ;
	wire _w16622_ ;
	wire _w16623_ ;
	wire _w16624_ ;
	wire _w16625_ ;
	wire _w16626_ ;
	wire _w16627_ ;
	wire _w16628_ ;
	wire _w16629_ ;
	wire _w16630_ ;
	wire _w16631_ ;
	wire _w16632_ ;
	wire _w16633_ ;
	wire _w16634_ ;
	wire _w16635_ ;
	wire _w16636_ ;
	wire _w16637_ ;
	wire _w16638_ ;
	wire _w16639_ ;
	wire _w16640_ ;
	wire _w16641_ ;
	wire _w16642_ ;
	wire _w16643_ ;
	wire _w16644_ ;
	wire _w16645_ ;
	wire _w16646_ ;
	wire _w16647_ ;
	wire _w16648_ ;
	wire _w16649_ ;
	wire _w16650_ ;
	wire _w16651_ ;
	wire _w16652_ ;
	wire _w16653_ ;
	wire _w16654_ ;
	wire _w16655_ ;
	wire _w16656_ ;
	wire _w16657_ ;
	wire _w16658_ ;
	wire _w16659_ ;
	wire _w16660_ ;
	wire _w16661_ ;
	wire _w16662_ ;
	wire _w16663_ ;
	wire _w16664_ ;
	wire _w16665_ ;
	wire _w16666_ ;
	wire _w16667_ ;
	wire _w16668_ ;
	wire _w16669_ ;
	wire _w16670_ ;
	wire _w16671_ ;
	wire _w16672_ ;
	wire _w16673_ ;
	wire _w16674_ ;
	wire _w16675_ ;
	wire _w16676_ ;
	wire _w16677_ ;
	wire _w16678_ ;
	wire _w16679_ ;
	wire _w16680_ ;
	wire _w16681_ ;
	wire _w16682_ ;
	wire _w16683_ ;
	wire _w16684_ ;
	wire _w16685_ ;
	wire _w16686_ ;
	wire _w16687_ ;
	wire _w16688_ ;
	wire _w16689_ ;
	wire _w16690_ ;
	wire _w16691_ ;
	wire _w16692_ ;
	wire _w16693_ ;
	wire _w16694_ ;
	wire _w16695_ ;
	wire _w16696_ ;
	wire _w16697_ ;
	wire _w16698_ ;
	wire _w16699_ ;
	wire _w16700_ ;
	wire _w16701_ ;
	wire _w16702_ ;
	wire _w16703_ ;
	wire _w16704_ ;
	wire _w16705_ ;
	wire _w16706_ ;
	wire _w16707_ ;
	wire _w16708_ ;
	wire _w16709_ ;
	wire _w16710_ ;
	wire _w16711_ ;
	wire _w16712_ ;
	wire _w16713_ ;
	wire _w16714_ ;
	wire _w16715_ ;
	wire _w16716_ ;
	wire _w16717_ ;
	wire _w16718_ ;
	wire _w16719_ ;
	wire _w16720_ ;
	wire _w16721_ ;
	wire _w16722_ ;
	wire _w16723_ ;
	wire _w16724_ ;
	wire _w16725_ ;
	wire _w16726_ ;
	wire _w16727_ ;
	wire _w16728_ ;
	wire _w16729_ ;
	wire _w16730_ ;
	wire _w16731_ ;
	wire _w16732_ ;
	wire _w16733_ ;
	wire _w16734_ ;
	wire _w16735_ ;
	wire _w16736_ ;
	wire _w16737_ ;
	wire _w16738_ ;
	wire _w16739_ ;
	wire _w16740_ ;
	wire _w16741_ ;
	wire _w16742_ ;
	wire _w16743_ ;
	wire _w16744_ ;
	wire _w16745_ ;
	wire _w16746_ ;
	wire _w16747_ ;
	wire _w16748_ ;
	wire _w16749_ ;
	wire _w16750_ ;
	wire _w16751_ ;
	wire _w16752_ ;
	wire _w16753_ ;
	wire _w16754_ ;
	wire _w16755_ ;
	wire _w16756_ ;
	wire _w16757_ ;
	wire _w16758_ ;
	wire _w16759_ ;
	wire _w16760_ ;
	wire _w16761_ ;
	wire _w16762_ ;
	wire _w16763_ ;
	wire _w16764_ ;
	wire _w16765_ ;
	wire _w16766_ ;
	wire _w16767_ ;
	wire _w16768_ ;
	wire _w16769_ ;
	wire _w16770_ ;
	wire _w16771_ ;
	wire _w16772_ ;
	wire _w16773_ ;
	wire _w16774_ ;
	wire _w16775_ ;
	wire _w16776_ ;
	wire _w16777_ ;
	wire _w16778_ ;
	wire _w16779_ ;
	wire _w16780_ ;
	wire _w16781_ ;
	wire _w16782_ ;
	wire _w16783_ ;
	wire _w16784_ ;
	wire _w16785_ ;
	wire _w16786_ ;
	wire _w16787_ ;
	wire _w16788_ ;
	wire _w16789_ ;
	wire _w16790_ ;
	wire _w16791_ ;
	wire _w16792_ ;
	wire _w16793_ ;
	wire _w16794_ ;
	wire _w16795_ ;
	wire _w16796_ ;
	wire _w16797_ ;
	wire _w16798_ ;
	wire _w16799_ ;
	wire _w16800_ ;
	wire _w16801_ ;
	wire _w16802_ ;
	wire _w16803_ ;
	wire _w16804_ ;
	wire _w16805_ ;
	wire _w16806_ ;
	wire _w16807_ ;
	wire _w16808_ ;
	wire _w16809_ ;
	wire _w16810_ ;
	wire _w16811_ ;
	wire _w16812_ ;
	wire _w16813_ ;
	wire _w16814_ ;
	wire _w16815_ ;
	wire _w16816_ ;
	wire _w16817_ ;
	wire _w16818_ ;
	wire _w16819_ ;
	wire _w16820_ ;
	wire _w16821_ ;
	wire _w16822_ ;
	wire _w16823_ ;
	wire _w16824_ ;
	wire _w16825_ ;
	wire _w16826_ ;
	wire _w16827_ ;
	wire _w16828_ ;
	wire _w16829_ ;
	wire _w16830_ ;
	wire _w16831_ ;
	wire _w16832_ ;
	wire _w16833_ ;
	wire _w16834_ ;
	wire _w16835_ ;
	wire _w16836_ ;
	wire _w16837_ ;
	wire _w16838_ ;
	wire _w16839_ ;
	wire _w16840_ ;
	wire _w16841_ ;
	wire _w16842_ ;
	wire _w16843_ ;
	wire _w16844_ ;
	wire _w16845_ ;
	wire _w16846_ ;
	wire _w16847_ ;
	wire _w16848_ ;
	wire _w16849_ ;
	wire _w16850_ ;
	wire _w16851_ ;
	wire _w16852_ ;
	wire _w16853_ ;
	wire _w16854_ ;
	wire _w16855_ ;
	wire _w16856_ ;
	wire _w16857_ ;
	wire _w16858_ ;
	wire _w16859_ ;
	wire _w16860_ ;
	wire _w16861_ ;
	wire _w16862_ ;
	wire _w16863_ ;
	wire _w16864_ ;
	wire _w16865_ ;
	wire _w16866_ ;
	wire _w16867_ ;
	wire _w16868_ ;
	wire _w16869_ ;
	wire _w16870_ ;
	wire _w16871_ ;
	wire _w16872_ ;
	wire _w16873_ ;
	wire _w16874_ ;
	wire _w16875_ ;
	wire _w16876_ ;
	wire _w16877_ ;
	wire _w16878_ ;
	wire _w16879_ ;
	wire _w16880_ ;
	wire _w16881_ ;
	wire _w16882_ ;
	wire _w16883_ ;
	wire _w16884_ ;
	wire _w16885_ ;
	wire _w16886_ ;
	wire _w16887_ ;
	wire _w16888_ ;
	wire _w16889_ ;
	wire _w16890_ ;
	wire _w16891_ ;
	wire _w16892_ ;
	wire _w16893_ ;
	wire _w16894_ ;
	wire _w16895_ ;
	wire _w16896_ ;
	wire _w16897_ ;
	wire _w16898_ ;
	wire _w16899_ ;
	wire _w16900_ ;
	wire _w16901_ ;
	wire _w16902_ ;
	wire _w16903_ ;
	wire _w16904_ ;
	wire _w16905_ ;
	wire _w16906_ ;
	wire _w16907_ ;
	wire _w16908_ ;
	wire _w16909_ ;
	wire _w16910_ ;
	wire _w16911_ ;
	wire _w16912_ ;
	wire _w16913_ ;
	wire _w16914_ ;
	wire _w16915_ ;
	wire _w16916_ ;
	wire _w16917_ ;
	wire _w16918_ ;
	wire _w16919_ ;
	wire _w16920_ ;
	wire _w16921_ ;
	wire _w16922_ ;
	wire _w16923_ ;
	wire _w16924_ ;
	wire _w16925_ ;
	wire _w16926_ ;
	wire _w16927_ ;
	wire _w16928_ ;
	wire _w16929_ ;
	wire _w16930_ ;
	wire _w16931_ ;
	wire _w16932_ ;
	wire _w16933_ ;
	wire _w16934_ ;
	wire _w16935_ ;
	wire _w16936_ ;
	wire _w16937_ ;
	wire _w16938_ ;
	wire _w16939_ ;
	wire _w16940_ ;
	wire _w16941_ ;
	wire _w16942_ ;
	wire _w16943_ ;
	wire _w16944_ ;
	wire _w16945_ ;
	wire _w16946_ ;
	wire _w16947_ ;
	wire _w16948_ ;
	wire _w16949_ ;
	wire _w16950_ ;
	wire _w16951_ ;
	wire _w16952_ ;
	wire _w16953_ ;
	wire _w16954_ ;
	wire _w16955_ ;
	wire _w16956_ ;
	wire _w16957_ ;
	wire _w16958_ ;
	wire _w16959_ ;
	wire _w16960_ ;
	wire _w16961_ ;
	wire _w16962_ ;
	wire _w16963_ ;
	wire _w16964_ ;
	wire _w16965_ ;
	wire _w16966_ ;
	wire _w16967_ ;
	wire _w16968_ ;
	wire _w16969_ ;
	wire _w16970_ ;
	wire _w16971_ ;
	wire _w16972_ ;
	wire _w16973_ ;
	wire _w16974_ ;
	wire _w16975_ ;
	wire _w16976_ ;
	wire _w16977_ ;
	wire _w16978_ ;
	wire _w16979_ ;
	wire _w16980_ ;
	wire _w16981_ ;
	wire _w16982_ ;
	wire _w16983_ ;
	wire _w16984_ ;
	wire _w16985_ ;
	wire _w16986_ ;
	wire _w16987_ ;
	wire _w16988_ ;
	wire _w16989_ ;
	wire _w16990_ ;
	wire _w16991_ ;
	wire _w16992_ ;
	wire _w16993_ ;
	wire _w16994_ ;
	wire _w16995_ ;
	wire _w16996_ ;
	wire _w16997_ ;
	wire _w16998_ ;
	wire _w16999_ ;
	wire _w17000_ ;
	wire _w17001_ ;
	wire _w17002_ ;
	wire _w17003_ ;
	wire _w17004_ ;
	wire _w17005_ ;
	wire _w17006_ ;
	wire _w17007_ ;
	wire _w17008_ ;
	wire _w17009_ ;
	wire _w17010_ ;
	wire _w17011_ ;
	wire _w17012_ ;
	wire _w17013_ ;
	wire _w17014_ ;
	wire _w17015_ ;
	wire _w17016_ ;
	wire _w17017_ ;
	wire _w17018_ ;
	wire _w17019_ ;
	wire _w17020_ ;
	wire _w17021_ ;
	wire _w17022_ ;
	wire _w17023_ ;
	wire _w17024_ ;
	wire _w17025_ ;
	wire _w17026_ ;
	wire _w17027_ ;
	wire _w17028_ ;
	wire _w17029_ ;
	wire _w17030_ ;
	wire _w17031_ ;
	wire _w17032_ ;
	wire _w17033_ ;
	wire _w17034_ ;
	wire _w17035_ ;
	wire _w17036_ ;
	wire _w17037_ ;
	wire _w17038_ ;
	wire _w17039_ ;
	wire _w17040_ ;
	wire _w17041_ ;
	wire _w17042_ ;
	wire _w17043_ ;
	wire _w17044_ ;
	wire _w17045_ ;
	wire _w17046_ ;
	wire _w17047_ ;
	wire _w17048_ ;
	wire _w17049_ ;
	wire _w17050_ ;
	wire _w17051_ ;
	wire _w17052_ ;
	wire _w17053_ ;
	wire _w17054_ ;
	wire _w17055_ ;
	wire _w17056_ ;
	wire _w17057_ ;
	wire _w17058_ ;
	wire _w17059_ ;
	wire _w17060_ ;
	wire _w17061_ ;
	wire _w17062_ ;
	wire _w17063_ ;
	wire _w17064_ ;
	wire _w17065_ ;
	wire _w17066_ ;
	wire _w17067_ ;
	wire _w17068_ ;
	wire _w17069_ ;
	wire _w17070_ ;
	wire _w17071_ ;
	wire _w17072_ ;
	wire _w17073_ ;
	wire _w17074_ ;
	wire _w17075_ ;
	wire _w17076_ ;
	wire _w17077_ ;
	wire _w17078_ ;
	wire _w17079_ ;
	wire _w17080_ ;
	wire _w17081_ ;
	wire _w17082_ ;
	wire _w17083_ ;
	wire _w17084_ ;
	wire _w17085_ ;
	wire _w17086_ ;
	wire _w17087_ ;
	wire _w17088_ ;
	wire _w17089_ ;
	wire _w17090_ ;
	wire _w17091_ ;
	wire _w17092_ ;
	wire _w17093_ ;
	wire _w17094_ ;
	wire _w17095_ ;
	wire _w17096_ ;
	wire _w17097_ ;
	wire _w17098_ ;
	wire _w17099_ ;
	wire _w17100_ ;
	wire _w17101_ ;
	wire _w17102_ ;
	wire _w17103_ ;
	wire _w17104_ ;
	wire _w17105_ ;
	wire _w17106_ ;
	wire _w17107_ ;
	wire _w17108_ ;
	wire _w17109_ ;
	wire _w17110_ ;
	wire _w17111_ ;
	wire _w17112_ ;
	wire _w17113_ ;
	wire _w17114_ ;
	wire _w17115_ ;
	wire _w17116_ ;
	wire _w17117_ ;
	wire _w17118_ ;
	wire _w17119_ ;
	wire _w17120_ ;
	wire _w17121_ ;
	wire _w17122_ ;
	wire _w17123_ ;
	wire _w17124_ ;
	wire _w17125_ ;
	wire _w17126_ ;
	wire _w17127_ ;
	wire _w17128_ ;
	wire _w17129_ ;
	wire _w17130_ ;
	wire _w17131_ ;
	wire _w17132_ ;
	wire _w17133_ ;
	wire _w17134_ ;
	wire _w17135_ ;
	wire _w17136_ ;
	wire _w17137_ ;
	wire _w17138_ ;
	wire _w17139_ ;
	wire _w17140_ ;
	wire _w17141_ ;
	wire _w17142_ ;
	wire _w17143_ ;
	wire _w17144_ ;
	wire _w17145_ ;
	wire _w17146_ ;
	wire _w17147_ ;
	wire _w17148_ ;
	wire _w17149_ ;
	wire _w17150_ ;
	wire _w17151_ ;
	wire _w17152_ ;
	wire _w17153_ ;
	wire _w17154_ ;
	wire _w17155_ ;
	wire _w17156_ ;
	wire _w17157_ ;
	wire _w17158_ ;
	wire _w17159_ ;
	wire _w17160_ ;
	wire _w17161_ ;
	wire _w17162_ ;
	wire _w17163_ ;
	wire _w17164_ ;
	wire _w17165_ ;
	wire _w17166_ ;
	wire _w17167_ ;
	wire _w17168_ ;
	wire _w17169_ ;
	wire _w17170_ ;
	wire _w17171_ ;
	wire _w17172_ ;
	wire _w17173_ ;
	wire _w17174_ ;
	wire _w17175_ ;
	wire _w17176_ ;
	wire _w17177_ ;
	wire _w17178_ ;
	wire _w17179_ ;
	wire _w17180_ ;
	wire _w17181_ ;
	wire _w17182_ ;
	wire _w17183_ ;
	wire _w17184_ ;
	wire _w17185_ ;
	wire _w17186_ ;
	wire _w17187_ ;
	wire _w17188_ ;
	wire _w17189_ ;
	wire _w17190_ ;
	wire _w17191_ ;
	wire _w17192_ ;
	wire _w17193_ ;
	wire _w17194_ ;
	wire _w17195_ ;
	wire _w17196_ ;
	wire _w17197_ ;
	wire _w17198_ ;
	wire _w17199_ ;
	wire _w17200_ ;
	wire _w17201_ ;
	wire _w17202_ ;
	wire _w17203_ ;
	wire _w17204_ ;
	wire _w17205_ ;
	wire _w17206_ ;
	wire _w17207_ ;
	wire _w17208_ ;
	wire _w17209_ ;
	wire _w17210_ ;
	wire _w17211_ ;
	wire _w17212_ ;
	wire _w17213_ ;
	wire _w17214_ ;
	wire _w17215_ ;
	wire _w17216_ ;
	wire _w17217_ ;
	wire _w17218_ ;
	wire _w17219_ ;
	wire _w17220_ ;
	wire _w17221_ ;
	wire _w17222_ ;
	wire _w17223_ ;
	wire _w17224_ ;
	wire _w17225_ ;
	wire _w17226_ ;
	wire _w17227_ ;
	wire _w17228_ ;
	wire _w17229_ ;
	wire _w17230_ ;
	wire _w17231_ ;
	wire _w17232_ ;
	wire _w17233_ ;
	wire _w17234_ ;
	wire _w17235_ ;
	wire _w17236_ ;
	wire _w17237_ ;
	wire _w17238_ ;
	wire _w17239_ ;
	wire _w17240_ ;
	wire _w17241_ ;
	wire _w17242_ ;
	wire _w17243_ ;
	wire _w17244_ ;
	wire _w17245_ ;
	wire _w17246_ ;
	wire _w17247_ ;
	wire _w17248_ ;
	wire _w17249_ ;
	wire _w17250_ ;
	wire _w17251_ ;
	wire _w17252_ ;
	wire _w17253_ ;
	wire _w17254_ ;
	wire _w17255_ ;
	wire _w17256_ ;
	wire _w17257_ ;
	wire _w17258_ ;
	wire _w17259_ ;
	wire _w17260_ ;
	wire _w17261_ ;
	wire _w17262_ ;
	wire _w17263_ ;
	wire _w17264_ ;
	wire _w17265_ ;
	wire _w17266_ ;
	wire _w17267_ ;
	wire _w17268_ ;
	wire _w17269_ ;
	wire _w17270_ ;
	wire _w17271_ ;
	wire _w17272_ ;
	wire _w17273_ ;
	wire _w17274_ ;
	wire _w17275_ ;
	wire _w17276_ ;
	wire _w17277_ ;
	wire _w17278_ ;
	wire _w17279_ ;
	wire _w17280_ ;
	wire _w17281_ ;
	wire _w17282_ ;
	wire _w17283_ ;
	wire _w17284_ ;
	wire _w17285_ ;
	wire _w17286_ ;
	wire _w17287_ ;
	wire _w17288_ ;
	wire _w17289_ ;
	wire _w17290_ ;
	wire _w17291_ ;
	wire _w17292_ ;
	wire _w17293_ ;
	wire _w17294_ ;
	wire _w17295_ ;
	wire _w17296_ ;
	wire _w17297_ ;
	wire _w17298_ ;
	wire _w17299_ ;
	wire _w17300_ ;
	wire _w17301_ ;
	wire _w17302_ ;
	wire _w17303_ ;
	wire _w17304_ ;
	wire _w17305_ ;
	wire _w17306_ ;
	wire _w17307_ ;
	wire _w17308_ ;
	wire _w17309_ ;
	wire _w17310_ ;
	wire _w17311_ ;
	wire _w17312_ ;
	wire _w17313_ ;
	wire _w17314_ ;
	wire _w17315_ ;
	wire _w17316_ ;
	wire _w17317_ ;
	wire _w17318_ ;
	wire _w17319_ ;
	wire _w17320_ ;
	wire _w17321_ ;
	wire _w17322_ ;
	wire _w17323_ ;
	wire _w17324_ ;
	wire _w17325_ ;
	wire _w17326_ ;
	wire _w17327_ ;
	wire _w17328_ ;
	wire _w17329_ ;
	wire _w17330_ ;
	wire _w17331_ ;
	wire _w17332_ ;
	wire _w17333_ ;
	wire _w17334_ ;
	wire _w17335_ ;
	wire _w17336_ ;
	wire _w17337_ ;
	wire _w17338_ ;
	wire _w17339_ ;
	wire _w17340_ ;
	wire _w17341_ ;
	wire _w17342_ ;
	wire _w17343_ ;
	wire _w17344_ ;
	wire _w17345_ ;
	wire _w17346_ ;
	wire _w17347_ ;
	wire _w17348_ ;
	wire _w17349_ ;
	wire _w17350_ ;
	wire _w17351_ ;
	wire _w17352_ ;
	wire _w17353_ ;
	wire _w17354_ ;
	wire _w17355_ ;
	wire _w17356_ ;
	wire _w17357_ ;
	wire _w17358_ ;
	wire _w17359_ ;
	wire _w17360_ ;
	wire _w17361_ ;
	wire _w17362_ ;
	wire _w17363_ ;
	wire _w17364_ ;
	wire _w17365_ ;
	wire _w17366_ ;
	wire _w17367_ ;
	wire _w17368_ ;
	wire _w17369_ ;
	wire _w17370_ ;
	wire _w17371_ ;
	wire _w17372_ ;
	wire _w17373_ ;
	wire _w17374_ ;
	wire _w17375_ ;
	wire _w17376_ ;
	wire _w17377_ ;
	wire _w17378_ ;
	wire _w17379_ ;
	wire _w17380_ ;
	wire _w17381_ ;
	wire _w17382_ ;
	wire _w17383_ ;
	wire _w17384_ ;
	wire _w17385_ ;
	wire _w17386_ ;
	wire _w17387_ ;
	wire _w17388_ ;
	wire _w17389_ ;
	wire _w17390_ ;
	wire _w17391_ ;
	wire _w17392_ ;
	wire _w17393_ ;
	wire _w17394_ ;
	wire _w17395_ ;
	wire _w17396_ ;
	wire _w17397_ ;
	wire _w17398_ ;
	wire _w17399_ ;
	wire _w17400_ ;
	wire _w17401_ ;
	wire _w17402_ ;
	wire _w17403_ ;
	wire _w17404_ ;
	wire _w17405_ ;
	wire _w17406_ ;
	wire _w17407_ ;
	wire _w17408_ ;
	wire _w17409_ ;
	wire _w17410_ ;
	wire _w17411_ ;
	wire _w17412_ ;
	wire _w17413_ ;
	wire _w17414_ ;
	wire _w17415_ ;
	wire _w17416_ ;
	wire _w17417_ ;
	wire _w17418_ ;
	wire _w17419_ ;
	wire _w17420_ ;
	wire _w17421_ ;
	wire _w17422_ ;
	wire _w17423_ ;
	wire _w17424_ ;
	wire _w17425_ ;
	wire _w17426_ ;
	wire _w17427_ ;
	wire _w17428_ ;
	wire _w17429_ ;
	wire _w17430_ ;
	wire _w17431_ ;
	wire _w17432_ ;
	wire _w17433_ ;
	wire _w17434_ ;
	wire _w17435_ ;
	wire _w17436_ ;
	wire _w17437_ ;
	wire _w17438_ ;
	wire _w17439_ ;
	wire _w17440_ ;
	wire _w17441_ ;
	wire _w17442_ ;
	wire _w17443_ ;
	wire _w17444_ ;
	wire _w17445_ ;
	wire _w17446_ ;
	wire _w17447_ ;
	wire _w17448_ ;
	wire _w17449_ ;
	wire _w17450_ ;
	wire _w17451_ ;
	wire _w17452_ ;
	wire _w17453_ ;
	wire _w17454_ ;
	wire _w17455_ ;
	wire _w17456_ ;
	wire _w17457_ ;
	wire _w17458_ ;
	wire _w17459_ ;
	wire _w17460_ ;
	wire _w17461_ ;
	wire _w17462_ ;
	wire _w17463_ ;
	wire _w17464_ ;
	wire _w17465_ ;
	wire _w17466_ ;
	wire _w17467_ ;
	wire _w17468_ ;
	wire _w17469_ ;
	wire _w17470_ ;
	wire _w17471_ ;
	wire _w17472_ ;
	wire _w17473_ ;
	wire _w17474_ ;
	wire _w17475_ ;
	wire _w17476_ ;
	wire _w17477_ ;
	wire _w17478_ ;
	wire _w17479_ ;
	wire _w17480_ ;
	wire _w17481_ ;
	wire _w17482_ ;
	wire _w17483_ ;
	wire _w17484_ ;
	wire _w17485_ ;
	wire _w17486_ ;
	wire _w17487_ ;
	wire _w17488_ ;
	wire _w17489_ ;
	wire _w17490_ ;
	wire _w17491_ ;
	wire _w17492_ ;
	wire _w17493_ ;
	wire _w17494_ ;
	wire _w17495_ ;
	wire _w17496_ ;
	wire _w17497_ ;
	wire _w17498_ ;
	wire _w17499_ ;
	wire _w17500_ ;
	wire _w17501_ ;
	wire _w17502_ ;
	wire _w17503_ ;
	wire _w17504_ ;
	wire _w17505_ ;
	wire _w17506_ ;
	wire _w17507_ ;
	wire _w17508_ ;
	wire _w17509_ ;
	wire _w17510_ ;
	wire _w17511_ ;
	wire _w17512_ ;
	wire _w17513_ ;
	wire _w17514_ ;
	wire _w17515_ ;
	wire _w17516_ ;
	wire _w17517_ ;
	wire _w17518_ ;
	wire _w17519_ ;
	wire _w17520_ ;
	wire _w17521_ ;
	wire _w17522_ ;
	wire _w17523_ ;
	wire _w17524_ ;
	wire _w17525_ ;
	wire _w17526_ ;
	wire _w17527_ ;
	wire _w17528_ ;
	wire _w17529_ ;
	wire _w17530_ ;
	wire _w17531_ ;
	wire _w17532_ ;
	wire _w17533_ ;
	wire _w17534_ ;
	wire _w17535_ ;
	wire _w17536_ ;
	wire _w17537_ ;
	wire _w17538_ ;
	wire _w17539_ ;
	wire _w17540_ ;
	wire _w17541_ ;
	wire _w17542_ ;
	wire _w17543_ ;
	wire _w17544_ ;
	wire _w17545_ ;
	wire _w17546_ ;
	wire _w17547_ ;
	wire _w17548_ ;
	wire _w17549_ ;
	wire _w17550_ ;
	wire _w17551_ ;
	wire _w17552_ ;
	wire _w17553_ ;
	wire _w17554_ ;
	wire _w17555_ ;
	wire _w17556_ ;
	wire _w17557_ ;
	wire _w17558_ ;
	wire _w17559_ ;
	wire _w17560_ ;
	wire _w17561_ ;
	wire _w17562_ ;
	wire _w17563_ ;
	wire _w17564_ ;
	wire _w17565_ ;
	wire _w17566_ ;
	wire _w17567_ ;
	wire _w17568_ ;
	wire _w17569_ ;
	wire _w17570_ ;
	wire _w17571_ ;
	wire _w17572_ ;
	wire _w17573_ ;
	wire _w17574_ ;
	wire _w17575_ ;
	wire _w17576_ ;
	wire _w17577_ ;
	wire _w17578_ ;
	wire _w17579_ ;
	wire _w17580_ ;
	wire _w17581_ ;
	wire _w17582_ ;
	wire _w17583_ ;
	wire _w17584_ ;
	wire _w17585_ ;
	wire _w17586_ ;
	wire _w17587_ ;
	wire _w17588_ ;
	wire _w17589_ ;
	wire _w17590_ ;
	wire _w17591_ ;
	wire _w17592_ ;
	wire _w17593_ ;
	wire _w17594_ ;
	wire _w17595_ ;
	wire _w17596_ ;
	wire _w17597_ ;
	wire _w17598_ ;
	wire _w17599_ ;
	wire _w17600_ ;
	wire _w17601_ ;
	wire _w17602_ ;
	wire _w17603_ ;
	wire _w17604_ ;
	wire _w17605_ ;
	wire _w17606_ ;
	wire _w17607_ ;
	wire _w17608_ ;
	wire _w17609_ ;
	wire _w17610_ ;
	wire _w17611_ ;
	wire _w17612_ ;
	wire _w17613_ ;
	wire _w17614_ ;
	wire _w17615_ ;
	wire _w17616_ ;
	wire _w17617_ ;
	wire _w17618_ ;
	wire _w17619_ ;
	wire _w17620_ ;
	wire _w17621_ ;
	wire _w17622_ ;
	wire _w17623_ ;
	wire _w17624_ ;
	wire _w17625_ ;
	wire _w17626_ ;
	wire _w17627_ ;
	wire _w17628_ ;
	wire _w17629_ ;
	wire _w17630_ ;
	wire _w17631_ ;
	wire _w17632_ ;
	wire _w17633_ ;
	wire _w17634_ ;
	wire _w17635_ ;
	wire _w17636_ ;
	wire _w17637_ ;
	wire _w17638_ ;
	wire _w17639_ ;
	wire _w17640_ ;
	wire _w17641_ ;
	wire _w17642_ ;
	wire _w17643_ ;
	wire _w17644_ ;
	wire _w17645_ ;
	wire _w17646_ ;
	wire _w17647_ ;
	wire _w17648_ ;
	wire _w17649_ ;
	wire _w17650_ ;
	wire _w17651_ ;
	wire _w17652_ ;
	wire _w17653_ ;
	wire _w17654_ ;
	wire _w17655_ ;
	wire _w17656_ ;
	wire _w17657_ ;
	wire _w17658_ ;
	wire _w17659_ ;
	wire _w17660_ ;
	wire _w17661_ ;
	wire _w17662_ ;
	wire _w17663_ ;
	wire _w17664_ ;
	wire _w17665_ ;
	wire _w17666_ ;
	wire _w17667_ ;
	wire _w17668_ ;
	wire _w17669_ ;
	wire _w17670_ ;
	wire _w17671_ ;
	wire _w17672_ ;
	wire _w17673_ ;
	wire _w17674_ ;
	wire _w17675_ ;
	wire _w17676_ ;
	wire _w17677_ ;
	wire _w17678_ ;
	wire _w17679_ ;
	wire _w17680_ ;
	wire _w17681_ ;
	wire _w17682_ ;
	wire _w17683_ ;
	wire _w17684_ ;
	wire _w17685_ ;
	wire _w17686_ ;
	wire _w17687_ ;
	wire _w17688_ ;
	wire _w17689_ ;
	wire _w17690_ ;
	wire _w17691_ ;
	wire _w17692_ ;
	wire _w17693_ ;
	wire _w17694_ ;
	wire _w17695_ ;
	wire _w17696_ ;
	wire _w17697_ ;
	wire _w17698_ ;
	wire _w17699_ ;
	wire _w17700_ ;
	wire _w17701_ ;
	wire _w17702_ ;
	wire _w17703_ ;
	wire _w17704_ ;
	wire _w17705_ ;
	wire _w17706_ ;
	wire _w17707_ ;
	wire _w17708_ ;
	wire _w17709_ ;
	wire _w17710_ ;
	wire _w17711_ ;
	wire _w17712_ ;
	wire _w17713_ ;
	wire _w17714_ ;
	wire _w17715_ ;
	wire _w17716_ ;
	wire _w17717_ ;
	wire _w17718_ ;
	wire _w17719_ ;
	wire _w17720_ ;
	wire _w17721_ ;
	wire _w17722_ ;
	wire _w17723_ ;
	wire _w17724_ ;
	wire _w17725_ ;
	wire _w17726_ ;
	wire _w17727_ ;
	wire _w17728_ ;
	wire _w17729_ ;
	wire _w17730_ ;
	wire _w17731_ ;
	wire _w17732_ ;
	wire _w17733_ ;
	wire _w17734_ ;
	wire _w17735_ ;
	wire _w17736_ ;
	wire _w17737_ ;
	wire _w17738_ ;
	wire _w17739_ ;
	wire _w17740_ ;
	wire _w17741_ ;
	wire _w17742_ ;
	wire _w17743_ ;
	wire _w17744_ ;
	wire _w17745_ ;
	wire _w17746_ ;
	wire _w17747_ ;
	wire _w17748_ ;
	wire _w17749_ ;
	wire _w17750_ ;
	wire _w17751_ ;
	wire _w17752_ ;
	wire _w17753_ ;
	wire _w17754_ ;
	wire _w17755_ ;
	wire _w17756_ ;
	wire _w17757_ ;
	wire _w17758_ ;
	wire _w17759_ ;
	wire _w17760_ ;
	wire _w17761_ ;
	wire _w17762_ ;
	wire _w17763_ ;
	wire _w17764_ ;
	wire _w17765_ ;
	wire _w17766_ ;
	wire _w17767_ ;
	wire _w17768_ ;
	wire _w17769_ ;
	wire _w17770_ ;
	wire _w17771_ ;
	wire _w17772_ ;
	wire _w17773_ ;
	wire _w17774_ ;
	wire _w17775_ ;
	wire _w17776_ ;
	wire _w17777_ ;
	wire _w17778_ ;
	wire _w17779_ ;
	wire _w17780_ ;
	wire _w17781_ ;
	wire _w17782_ ;
	wire _w17783_ ;
	wire _w17784_ ;
	wire _w17785_ ;
	wire _w17786_ ;
	wire _w17787_ ;
	wire _w17788_ ;
	wire _w17789_ ;
	wire _w17790_ ;
	wire _w17791_ ;
	wire _w17792_ ;
	wire _w17793_ ;
	wire _w17794_ ;
	wire _w17795_ ;
	wire _w17796_ ;
	wire _w17797_ ;
	wire _w17798_ ;
	wire _w17799_ ;
	wire _w17800_ ;
	wire _w17801_ ;
	wire _w17802_ ;
	wire _w17803_ ;
	wire _w17804_ ;
	wire _w17805_ ;
	wire _w17806_ ;
	wire _w17807_ ;
	wire _w17808_ ;
	wire _w17809_ ;
	wire _w17810_ ;
	wire _w17811_ ;
	wire _w17812_ ;
	wire _w17813_ ;
	wire _w17814_ ;
	wire _w17815_ ;
	wire _w17816_ ;
	wire _w17817_ ;
	wire _w17818_ ;
	wire _w17819_ ;
	wire _w17820_ ;
	wire _w17821_ ;
	wire _w17822_ ;
	wire _w17823_ ;
	wire _w17824_ ;
	wire _w17825_ ;
	wire _w17826_ ;
	wire _w17827_ ;
	wire _w17828_ ;
	wire _w17829_ ;
	wire _w17830_ ;
	wire _w17831_ ;
	wire _w17832_ ;
	wire _w17833_ ;
	wire _w17834_ ;
	wire _w17835_ ;
	wire _w17836_ ;
	wire _w17837_ ;
	wire _w17838_ ;
	wire _w17839_ ;
	wire _w17840_ ;
	wire _w17841_ ;
	wire _w17842_ ;
	wire _w17843_ ;
	wire _w17844_ ;
	wire _w17845_ ;
	wire _w17846_ ;
	wire _w17847_ ;
	wire _w17848_ ;
	wire _w17849_ ;
	wire _w17850_ ;
	wire _w17851_ ;
	wire _w17852_ ;
	wire _w17853_ ;
	wire _w17854_ ;
	wire _w17855_ ;
	wire _w17856_ ;
	wire _w17857_ ;
	wire _w17858_ ;
	wire _w17859_ ;
	wire _w17860_ ;
	wire _w17861_ ;
	wire _w17862_ ;
	wire _w17863_ ;
	wire _w17864_ ;
	wire _w17865_ ;
	wire _w17866_ ;
	wire _w17867_ ;
	wire _w17868_ ;
	wire _w17869_ ;
	wire _w17870_ ;
	wire _w17871_ ;
	wire _w17872_ ;
	wire _w17873_ ;
	wire _w17874_ ;
	wire _w17875_ ;
	wire _w17876_ ;
	wire _w17877_ ;
	wire _w17878_ ;
	wire _w17879_ ;
	wire _w17880_ ;
	wire _w17881_ ;
	wire _w17882_ ;
	wire _w17883_ ;
	wire _w17884_ ;
	wire _w17885_ ;
	wire _w17886_ ;
	wire _w17887_ ;
	wire _w17888_ ;
	wire _w17889_ ;
	wire _w17890_ ;
	wire _w17891_ ;
	wire _w17892_ ;
	wire _w17893_ ;
	wire _w17894_ ;
	wire _w17895_ ;
	wire _w17896_ ;
	wire _w17897_ ;
	wire _w17898_ ;
	wire _w17899_ ;
	wire _w17900_ ;
	wire _w17901_ ;
	wire _w17902_ ;
	wire _w17903_ ;
	wire _w17904_ ;
	wire _w17905_ ;
	wire _w17906_ ;
	wire _w17907_ ;
	wire _w17908_ ;
	wire _w17909_ ;
	wire _w17910_ ;
	wire _w17911_ ;
	wire _w17912_ ;
	wire _w17913_ ;
	wire _w17914_ ;
	wire _w17915_ ;
	wire _w17916_ ;
	wire _w17917_ ;
	wire _w17918_ ;
	wire _w17919_ ;
	wire _w17920_ ;
	wire _w17921_ ;
	wire _w17922_ ;
	wire _w17923_ ;
	wire _w17924_ ;
	wire _w17925_ ;
	wire _w17926_ ;
	wire _w17927_ ;
	wire _w17928_ ;
	wire _w17929_ ;
	wire _w17930_ ;
	wire _w17931_ ;
	wire _w17932_ ;
	wire _w17933_ ;
	wire _w17934_ ;
	wire _w17935_ ;
	wire _w17936_ ;
	wire _w17937_ ;
	wire _w17938_ ;
	wire _w17939_ ;
	wire _w17940_ ;
	wire _w17941_ ;
	wire _w17942_ ;
	wire _w17943_ ;
	wire _w17944_ ;
	wire _w17945_ ;
	wire _w17946_ ;
	wire _w17947_ ;
	wire _w17948_ ;
	wire _w17949_ ;
	wire _w17950_ ;
	wire _w17951_ ;
	wire _w17952_ ;
	wire _w17953_ ;
	wire _w17954_ ;
	wire _w17955_ ;
	wire _w17956_ ;
	wire _w17957_ ;
	wire _w17958_ ;
	wire _w17959_ ;
	wire _w17960_ ;
	wire _w17961_ ;
	wire _w17962_ ;
	wire _w17963_ ;
	wire _w17964_ ;
	wire _w17965_ ;
	wire _w17966_ ;
	wire _w17967_ ;
	wire _w17968_ ;
	wire _w17969_ ;
	wire _w17970_ ;
	wire _w17971_ ;
	wire _w17972_ ;
	wire _w17973_ ;
	wire _w17974_ ;
	wire _w17975_ ;
	wire _w17976_ ;
	wire _w17977_ ;
	wire _w17978_ ;
	wire _w17979_ ;
	wire _w17980_ ;
	wire _w17981_ ;
	wire _w17982_ ;
	wire _w17983_ ;
	wire _w17984_ ;
	wire _w17985_ ;
	wire _w17986_ ;
	wire _w17987_ ;
	wire _w17988_ ;
	wire _w17989_ ;
	wire _w17990_ ;
	wire _w17991_ ;
	wire _w17992_ ;
	wire _w17993_ ;
	wire _w17994_ ;
	wire _w17995_ ;
	wire _w17996_ ;
	wire _w17997_ ;
	wire _w17998_ ;
	wire _w17999_ ;
	wire _w18000_ ;
	wire _w18001_ ;
	wire _w18002_ ;
	wire _w18003_ ;
	wire _w18004_ ;
	wire _w18005_ ;
	wire _w18006_ ;
	wire _w18007_ ;
	wire _w18008_ ;
	wire _w18009_ ;
	wire _w18010_ ;
	wire _w18011_ ;
	wire _w18012_ ;
	wire _w18013_ ;
	wire _w18014_ ;
	wire _w18015_ ;
	wire _w18016_ ;
	wire _w18017_ ;
	wire _w18018_ ;
	wire _w18019_ ;
	wire _w18020_ ;
	wire _w18021_ ;
	wire _w18022_ ;
	wire _w18023_ ;
	wire _w18024_ ;
	wire _w18025_ ;
	wire _w18026_ ;
	wire _w18027_ ;
	wire _w18028_ ;
	wire _w18029_ ;
	wire _w18030_ ;
	wire _w18031_ ;
	wire _w18032_ ;
	wire _w18033_ ;
	wire _w18034_ ;
	wire _w18035_ ;
	wire _w18036_ ;
	wire _w18037_ ;
	wire _w18038_ ;
	wire _w18039_ ;
	wire _w18040_ ;
	wire _w18041_ ;
	wire _w18042_ ;
	wire _w18043_ ;
	wire _w18044_ ;
	wire _w18045_ ;
	wire _w18046_ ;
	wire _w18047_ ;
	wire _w18048_ ;
	wire _w18049_ ;
	wire _w18050_ ;
	wire _w18051_ ;
	wire _w18052_ ;
	wire _w18053_ ;
	wire _w18054_ ;
	wire _w18055_ ;
	wire _w18056_ ;
	wire _w18057_ ;
	wire _w18058_ ;
	wire _w18059_ ;
	wire _w18060_ ;
	wire _w18061_ ;
	wire _w18062_ ;
	wire _w18063_ ;
	wire _w18064_ ;
	wire _w18065_ ;
	wire _w18066_ ;
	wire _w18067_ ;
	wire _w18068_ ;
	wire _w18069_ ;
	wire _w18070_ ;
	wire _w18071_ ;
	wire _w18072_ ;
	wire _w18073_ ;
	wire _w18074_ ;
	wire _w18075_ ;
	wire _w18076_ ;
	wire _w18077_ ;
	wire _w18078_ ;
	wire _w18079_ ;
	wire _w18080_ ;
	wire _w18081_ ;
	wire _w18082_ ;
	wire _w18083_ ;
	wire _w18084_ ;
	wire _w18085_ ;
	wire _w18086_ ;
	wire _w18087_ ;
	wire _w18088_ ;
	wire _w18089_ ;
	wire _w18090_ ;
	wire _w18091_ ;
	wire _w18092_ ;
	wire _w18093_ ;
	wire _w18094_ ;
	wire _w18095_ ;
	wire _w18096_ ;
	wire _w18097_ ;
	wire _w18098_ ;
	wire _w18099_ ;
	wire _w18100_ ;
	wire _w18101_ ;
	wire _w18102_ ;
	wire _w18103_ ;
	wire _w18104_ ;
	wire _w18105_ ;
	wire _w18106_ ;
	wire _w18107_ ;
	wire _w18108_ ;
	wire _w18109_ ;
	wire _w18110_ ;
	wire _w18111_ ;
	wire _w18112_ ;
	wire _w18113_ ;
	wire _w18114_ ;
	wire _w18115_ ;
	wire _w18116_ ;
	wire _w18117_ ;
	wire _w18118_ ;
	wire _w18119_ ;
	wire _w18120_ ;
	wire _w18121_ ;
	wire _w18122_ ;
	wire _w18123_ ;
	wire _w18124_ ;
	wire _w18125_ ;
	wire _w18126_ ;
	wire _w18127_ ;
	wire _w18128_ ;
	wire _w18129_ ;
	wire _w18130_ ;
	wire _w18131_ ;
	wire _w18132_ ;
	wire _w18133_ ;
	wire _w18134_ ;
	wire _w18135_ ;
	wire _w18136_ ;
	wire _w18137_ ;
	wire _w18138_ ;
	wire _w18139_ ;
	wire _w18140_ ;
	wire _w18141_ ;
	wire _w18142_ ;
	wire _w18143_ ;
	wire _w18144_ ;
	wire _w18145_ ;
	wire _w18146_ ;
	wire _w18147_ ;
	wire _w18148_ ;
	wire _w18149_ ;
	wire _w18150_ ;
	wire _w18151_ ;
	wire _w18152_ ;
	wire _w18153_ ;
	wire _w18154_ ;
	wire _w18155_ ;
	wire _w18156_ ;
	wire _w18157_ ;
	wire _w18158_ ;
	wire _w18159_ ;
	wire _w18160_ ;
	wire _w18161_ ;
	wire _w18162_ ;
	wire _w18163_ ;
	wire _w18164_ ;
	wire _w18165_ ;
	wire _w18166_ ;
	wire _w18167_ ;
	wire _w18168_ ;
	wire _w18169_ ;
	wire _w18170_ ;
	wire _w18171_ ;
	wire _w18172_ ;
	wire _w18173_ ;
	wire _w18174_ ;
	wire _w18175_ ;
	wire _w18176_ ;
	wire _w18177_ ;
	wire _w18178_ ;
	wire _w18179_ ;
	wire _w18180_ ;
	wire _w18181_ ;
	wire _w18182_ ;
	wire _w18183_ ;
	wire _w18184_ ;
	wire _w18185_ ;
	wire _w18186_ ;
	wire _w18187_ ;
	wire _w18188_ ;
	wire _w18189_ ;
	wire _w18190_ ;
	wire _w18191_ ;
	wire _w18192_ ;
	wire _w18193_ ;
	wire _w18194_ ;
	wire _w18195_ ;
	wire _w18196_ ;
	wire _w18197_ ;
	wire _w18198_ ;
	wire _w18199_ ;
	wire _w18200_ ;
	wire _w18201_ ;
	wire _w18202_ ;
	wire _w18203_ ;
	wire _w18204_ ;
	wire _w18205_ ;
	wire _w18206_ ;
	wire _w18207_ ;
	wire _w18208_ ;
	wire _w18209_ ;
	wire _w18210_ ;
	wire _w18211_ ;
	wire _w18212_ ;
	wire _w18213_ ;
	wire _w18214_ ;
	wire _w18215_ ;
	wire _w18216_ ;
	wire _w18217_ ;
	wire _w18218_ ;
	wire _w18219_ ;
	wire _w18220_ ;
	wire _w18221_ ;
	wire _w18222_ ;
	wire _w18223_ ;
	wire _w18224_ ;
	wire _w18225_ ;
	wire _w18226_ ;
	wire _w18227_ ;
	wire _w18228_ ;
	wire _w18229_ ;
	wire _w18230_ ;
	wire _w18231_ ;
	wire _w18232_ ;
	wire _w18233_ ;
	wire _w18234_ ;
	wire _w18235_ ;
	wire _w18236_ ;
	wire _w18237_ ;
	wire _w18238_ ;
	wire _w18239_ ;
	wire _w18240_ ;
	wire _w18241_ ;
	wire _w18242_ ;
	wire _w18243_ ;
	wire _w18244_ ;
	wire _w18245_ ;
	wire _w18246_ ;
	wire _w18247_ ;
	wire _w18248_ ;
	wire _w18249_ ;
	wire _w18250_ ;
	wire _w18251_ ;
	wire _w18252_ ;
	wire _w18253_ ;
	wire _w18254_ ;
	wire _w18255_ ;
	wire _w18256_ ;
	wire _w18257_ ;
	wire _w18258_ ;
	wire _w18259_ ;
	wire _w18260_ ;
	wire _w18261_ ;
	wire _w18262_ ;
	wire _w18263_ ;
	wire _w18264_ ;
	wire _w18265_ ;
	wire _w18266_ ;
	wire _w18267_ ;
	wire _w18268_ ;
	wire _w18269_ ;
	wire _w18270_ ;
	wire _w18271_ ;
	wire _w18272_ ;
	wire _w18273_ ;
	wire _w18274_ ;
	wire _w18275_ ;
	wire _w18276_ ;
	wire _w18277_ ;
	wire _w18278_ ;
	wire _w18279_ ;
	wire _w18280_ ;
	wire _w18281_ ;
	wire _w18282_ ;
	wire _w18283_ ;
	wire _w18284_ ;
	wire _w18285_ ;
	wire _w18286_ ;
	wire _w18287_ ;
	wire _w18288_ ;
	wire _w18289_ ;
	wire _w18290_ ;
	wire _w18291_ ;
	wire _w18292_ ;
	wire _w18293_ ;
	wire _w18294_ ;
	wire _w18295_ ;
	wire _w18296_ ;
	wire _w18297_ ;
	wire _w18298_ ;
	wire _w18299_ ;
	wire _w18300_ ;
	wire _w18301_ ;
	wire _w18302_ ;
	wire _w18303_ ;
	wire _w18304_ ;
	wire _w18305_ ;
	wire _w18306_ ;
	wire _w18307_ ;
	wire _w18308_ ;
	wire _w18309_ ;
	wire _w18310_ ;
	wire _w18311_ ;
	wire _w18312_ ;
	wire _w18313_ ;
	wire _w18314_ ;
	wire _w18315_ ;
	wire _w18316_ ;
	wire _w18317_ ;
	wire _w18318_ ;
	wire _w18319_ ;
	wire _w18320_ ;
	wire _w18321_ ;
	wire _w18322_ ;
	wire _w18323_ ;
	wire _w18324_ ;
	wire _w18325_ ;
	wire _w18326_ ;
	wire _w18327_ ;
	wire _w18328_ ;
	wire _w18329_ ;
	wire _w18330_ ;
	wire _w18331_ ;
	wire _w18332_ ;
	wire _w18333_ ;
	wire _w18334_ ;
	wire _w18335_ ;
	wire _w18336_ ;
	wire _w18337_ ;
	wire _w18338_ ;
	wire _w18339_ ;
	wire _w18340_ ;
	wire _w18341_ ;
	wire _w18342_ ;
	wire _w18343_ ;
	wire _w18344_ ;
	wire _w18345_ ;
	wire _w18346_ ;
	wire _w18347_ ;
	wire _w18348_ ;
	wire _w18349_ ;
	wire _w18350_ ;
	wire _w18351_ ;
	wire _w18352_ ;
	wire _w18353_ ;
	wire _w18354_ ;
	wire _w18355_ ;
	wire _w18356_ ;
	wire _w18357_ ;
	wire _w18358_ ;
	wire _w18359_ ;
	wire _w18360_ ;
	wire _w18361_ ;
	wire _w18362_ ;
	wire _w18363_ ;
	wire _w18364_ ;
	wire _w18365_ ;
	wire _w18366_ ;
	wire _w18367_ ;
	wire _w18368_ ;
	wire _w18369_ ;
	wire _w18370_ ;
	wire _w18371_ ;
	wire _w18372_ ;
	wire _w18373_ ;
	wire _w18374_ ;
	wire _w18375_ ;
	wire _w18376_ ;
	wire _w18377_ ;
	wire _w18378_ ;
	wire _w18379_ ;
	wire _w18380_ ;
	wire _w18381_ ;
	wire _w18382_ ;
	wire _w18383_ ;
	wire _w18384_ ;
	wire _w18385_ ;
	wire _w18386_ ;
	wire _w18387_ ;
	wire _w18388_ ;
	wire _w18389_ ;
	wire _w18390_ ;
	wire _w18391_ ;
	wire _w18392_ ;
	wire _w18393_ ;
	wire _w18394_ ;
	wire _w18395_ ;
	wire _w18396_ ;
	wire _w18397_ ;
	wire _w18398_ ;
	wire _w18399_ ;
	wire _w18400_ ;
	wire _w18401_ ;
	wire _w18402_ ;
	wire _w18403_ ;
	wire _w18404_ ;
	wire _w18405_ ;
	wire _w18406_ ;
	wire _w18407_ ;
	wire _w18408_ ;
	wire _w18409_ ;
	wire _w18410_ ;
	wire _w18411_ ;
	wire _w18412_ ;
	wire _w18413_ ;
	wire _w18414_ ;
	wire _w18415_ ;
	wire _w18416_ ;
	wire _w18417_ ;
	wire _w18418_ ;
	wire _w18419_ ;
	wire _w18420_ ;
	wire _w18421_ ;
	wire _w18422_ ;
	wire _w18423_ ;
	wire _w18424_ ;
	wire _w18425_ ;
	wire _w18426_ ;
	wire _w18427_ ;
	wire _w18428_ ;
	wire _w18429_ ;
	wire _w18430_ ;
	wire _w18431_ ;
	wire _w18432_ ;
	wire _w18433_ ;
	wire _w18434_ ;
	wire _w18435_ ;
	wire _w18436_ ;
	wire _w18437_ ;
	wire _w18438_ ;
	wire _w18439_ ;
	wire _w18440_ ;
	wire _w18441_ ;
	wire _w18442_ ;
	wire _w18443_ ;
	wire _w18444_ ;
	wire _w18445_ ;
	wire _w18446_ ;
	wire _w18447_ ;
	wire _w18448_ ;
	wire _w18449_ ;
	wire _w18450_ ;
	wire _w18451_ ;
	wire _w18452_ ;
	wire _w18453_ ;
	wire _w18454_ ;
	wire _w18455_ ;
	wire _w18456_ ;
	wire _w18457_ ;
	wire _w18458_ ;
	wire _w18459_ ;
	wire _w18460_ ;
	wire _w18461_ ;
	wire _w18462_ ;
	wire _w18463_ ;
	wire _w18464_ ;
	wire _w18465_ ;
	wire _w18466_ ;
	wire _w18467_ ;
	wire _w18468_ ;
	wire _w18469_ ;
	wire _w18470_ ;
	wire _w18471_ ;
	wire _w18472_ ;
	wire _w18473_ ;
	wire _w18474_ ;
	wire _w18475_ ;
	wire _w18476_ ;
	wire _w18477_ ;
	wire _w18478_ ;
	wire _w18479_ ;
	wire _w18480_ ;
	wire _w18481_ ;
	wire _w18482_ ;
	wire _w18483_ ;
	wire _w18484_ ;
	wire _w18485_ ;
	wire _w18486_ ;
	wire _w18487_ ;
	wire _w18488_ ;
	wire _w18489_ ;
	wire _w18490_ ;
	wire _w18491_ ;
	wire _w18492_ ;
	wire _w18493_ ;
	wire _w18494_ ;
	wire _w18495_ ;
	wire _w18496_ ;
	wire _w18497_ ;
	wire _w18498_ ;
	wire _w18499_ ;
	wire _w18500_ ;
	wire _w18501_ ;
	wire _w18502_ ;
	wire _w18503_ ;
	wire _w18504_ ;
	wire _w18505_ ;
	wire _w18506_ ;
	wire _w18507_ ;
	wire _w18508_ ;
	wire _w18509_ ;
	wire _w18510_ ;
	wire _w18511_ ;
	wire _w18512_ ;
	wire _w18513_ ;
	wire _w18514_ ;
	wire _w18515_ ;
	wire _w18516_ ;
	wire _w18517_ ;
	wire _w18518_ ;
	wire _w18519_ ;
	wire _w18520_ ;
	wire _w18521_ ;
	wire _w18522_ ;
	wire _w18523_ ;
	wire _w18524_ ;
	wire _w18525_ ;
	wire _w18526_ ;
	wire _w18527_ ;
	wire _w18528_ ;
	wire _w18529_ ;
	wire _w18530_ ;
	wire _w18531_ ;
	wire _w18532_ ;
	wire _w18533_ ;
	wire _w18534_ ;
	wire _w18535_ ;
	wire _w18536_ ;
	wire _w18537_ ;
	wire _w18538_ ;
	wire _w18539_ ;
	wire _w18540_ ;
	wire _w18541_ ;
	wire _w18542_ ;
	wire _w18543_ ;
	wire _w18544_ ;
	wire _w18545_ ;
	wire _w18546_ ;
	wire _w18547_ ;
	wire _w18548_ ;
	wire _w18549_ ;
	wire _w18550_ ;
	wire _w18551_ ;
	wire _w18552_ ;
	wire _w18553_ ;
	wire _w18554_ ;
	wire _w18555_ ;
	wire _w18556_ ;
	wire _w18557_ ;
	wire _w18558_ ;
	wire _w18559_ ;
	wire _w18560_ ;
	wire _w18561_ ;
	wire _w18562_ ;
	wire _w18563_ ;
	wire _w18564_ ;
	wire _w18565_ ;
	wire _w18566_ ;
	wire _w18567_ ;
	wire _w18568_ ;
	wire _w18569_ ;
	wire _w18570_ ;
	wire _w18571_ ;
	wire _w18572_ ;
	wire _w18573_ ;
	wire _w18574_ ;
	wire _w18575_ ;
	wire _w18576_ ;
	wire _w18577_ ;
	wire _w18578_ ;
	wire _w18579_ ;
	wire _w18580_ ;
	wire _w18581_ ;
	wire _w18582_ ;
	wire _w18583_ ;
	wire _w18584_ ;
	wire _w18585_ ;
	wire _w18586_ ;
	wire _w18587_ ;
	wire _w18588_ ;
	wire _w18589_ ;
	wire _w18590_ ;
	wire _w18591_ ;
	wire _w18592_ ;
	wire _w18593_ ;
	wire _w18594_ ;
	wire _w18595_ ;
	wire _w18596_ ;
	wire _w18597_ ;
	wire _w18598_ ;
	wire _w18599_ ;
	wire _w18600_ ;
	wire _w18601_ ;
	wire _w18602_ ;
	wire _w18603_ ;
	wire _w18604_ ;
	wire _w18605_ ;
	wire _w18606_ ;
	wire _w18607_ ;
	wire _w18608_ ;
	wire _w18609_ ;
	wire _w18610_ ;
	wire _w18611_ ;
	wire _w18612_ ;
	wire _w18613_ ;
	wire _w18614_ ;
	wire _w18615_ ;
	wire _w18616_ ;
	wire _w18617_ ;
	wire _w18618_ ;
	wire _w18619_ ;
	wire _w18620_ ;
	wire _w18621_ ;
	wire _w18622_ ;
	wire _w18623_ ;
	wire _w18624_ ;
	wire _w18625_ ;
	wire _w18626_ ;
	wire _w18627_ ;
	wire _w18628_ ;
	wire _w18629_ ;
	wire _w18630_ ;
	wire _w18631_ ;
	wire _w18632_ ;
	wire _w18633_ ;
	wire _w18634_ ;
	wire _w18635_ ;
	wire _w18636_ ;
	wire _w18637_ ;
	wire _w18638_ ;
	wire _w18639_ ;
	wire _w18640_ ;
	wire _w18641_ ;
	wire _w18642_ ;
	wire _w18643_ ;
	wire _w18644_ ;
	wire _w18645_ ;
	wire _w18646_ ;
	wire _w18647_ ;
	wire _w18648_ ;
	wire _w18649_ ;
	wire _w18650_ ;
	wire _w18651_ ;
	wire _w18652_ ;
	wire _w18653_ ;
	wire _w18654_ ;
	wire _w18655_ ;
	wire _w18656_ ;
	wire _w18657_ ;
	wire _w18658_ ;
	wire _w18659_ ;
	wire _w18660_ ;
	wire _w18661_ ;
	wire _w18662_ ;
	wire _w18663_ ;
	wire _w18664_ ;
	wire _w18665_ ;
	wire _w18666_ ;
	wire _w18667_ ;
	wire _w18668_ ;
	wire _w18669_ ;
	wire _w18670_ ;
	wire _w18671_ ;
	wire _w18672_ ;
	wire _w18673_ ;
	wire _w18674_ ;
	wire _w18675_ ;
	wire _w18676_ ;
	wire _w18677_ ;
	wire _w18678_ ;
	wire _w18679_ ;
	wire _w18680_ ;
	wire _w18681_ ;
	wire _w18682_ ;
	wire _w18683_ ;
	wire _w18684_ ;
	wire _w18685_ ;
	wire _w18686_ ;
	wire _w18687_ ;
	wire _w18688_ ;
	wire _w18689_ ;
	wire _w18690_ ;
	wire _w18691_ ;
	wire _w18692_ ;
	wire _w18693_ ;
	wire _w18694_ ;
	wire _w18695_ ;
	wire _w18696_ ;
	wire _w18697_ ;
	wire _w18698_ ;
	wire _w18699_ ;
	wire _w18700_ ;
	wire _w18701_ ;
	wire _w18702_ ;
	wire _w18703_ ;
	wire _w18704_ ;
	wire _w18705_ ;
	wire _w18706_ ;
	wire _w18707_ ;
	wire _w18708_ ;
	wire _w18709_ ;
	wire _w18710_ ;
	wire _w18711_ ;
	wire _w18712_ ;
	wire _w18713_ ;
	wire _w18714_ ;
	wire _w18715_ ;
	wire _w18716_ ;
	wire _w18717_ ;
	wire _w18718_ ;
	wire _w18719_ ;
	wire _w18720_ ;
	wire _w18721_ ;
	wire _w18722_ ;
	wire _w18723_ ;
	wire _w18724_ ;
	wire _w18725_ ;
	wire _w18726_ ;
	wire _w18727_ ;
	wire _w18728_ ;
	wire _w18729_ ;
	wire _w18730_ ;
	wire _w18731_ ;
	wire _w18732_ ;
	wire _w18733_ ;
	wire _w18734_ ;
	wire _w18735_ ;
	wire _w18736_ ;
	wire _w18737_ ;
	wire _w18738_ ;
	wire _w18739_ ;
	wire _w18740_ ;
	wire _w18741_ ;
	wire _w18742_ ;
	wire _w18743_ ;
	wire _w18744_ ;
	wire _w18745_ ;
	wire _w18746_ ;
	wire _w18747_ ;
	wire _w18748_ ;
	wire _w18749_ ;
	wire _w18750_ ;
	wire _w18751_ ;
	wire _w18752_ ;
	wire _w18753_ ;
	wire _w18754_ ;
	wire _w18755_ ;
	wire _w18756_ ;
	wire _w18757_ ;
	wire _w18758_ ;
	wire _w18759_ ;
	wire _w18760_ ;
	wire _w18761_ ;
	wire _w18762_ ;
	wire _w18763_ ;
	wire _w18764_ ;
	wire _w18765_ ;
	wire _w18766_ ;
	wire _w18767_ ;
	wire _w18768_ ;
	wire _w18769_ ;
	wire _w18770_ ;
	wire _w18771_ ;
	wire _w18772_ ;
	wire _w18773_ ;
	wire _w18774_ ;
	wire _w18775_ ;
	wire _w18776_ ;
	wire _w18777_ ;
	wire _w18778_ ;
	wire _w18779_ ;
	wire _w18780_ ;
	wire _w18781_ ;
	wire _w18782_ ;
	wire _w18783_ ;
	wire _w18784_ ;
	wire _w18785_ ;
	wire _w18786_ ;
	wire _w18787_ ;
	wire _w18788_ ;
	wire _w18789_ ;
	wire _w18790_ ;
	wire _w18791_ ;
	wire _w18792_ ;
	wire _w18793_ ;
	wire _w18794_ ;
	wire _w18795_ ;
	wire _w18796_ ;
	wire _w18797_ ;
	wire _w18798_ ;
	wire _w18799_ ;
	wire _w18800_ ;
	wire _w18801_ ;
	wire _w18802_ ;
	wire _w18803_ ;
	wire _w18804_ ;
	wire _w18805_ ;
	wire _w18806_ ;
	wire _w18807_ ;
	wire _w18808_ ;
	wire _w18809_ ;
	wire _w18810_ ;
	wire _w18811_ ;
	wire _w18812_ ;
	wire _w18813_ ;
	wire _w18814_ ;
	wire _w18815_ ;
	wire _w18816_ ;
	wire _w18817_ ;
	wire _w18818_ ;
	wire _w18819_ ;
	wire _w18820_ ;
	wire _w18821_ ;
	wire _w18822_ ;
	wire _w18823_ ;
	wire _w18824_ ;
	wire _w18825_ ;
	wire _w18826_ ;
	wire _w18827_ ;
	wire _w18828_ ;
	wire _w18829_ ;
	wire _w18830_ ;
	wire _w18831_ ;
	wire _w18832_ ;
	wire _w18833_ ;
	wire _w18834_ ;
	wire _w18835_ ;
	wire _w18836_ ;
	wire _w18837_ ;
	wire _w18838_ ;
	wire _w18839_ ;
	wire _w18840_ ;
	wire _w18841_ ;
	wire _w18842_ ;
	wire _w18843_ ;
	wire _w18844_ ;
	wire _w18845_ ;
	wire _w18846_ ;
	wire _w18847_ ;
	wire _w18848_ ;
	wire _w18849_ ;
	wire _w18850_ ;
	wire _w18851_ ;
	wire _w18852_ ;
	wire _w18853_ ;
	wire _w18854_ ;
	wire _w18855_ ;
	wire _w18856_ ;
	wire _w18857_ ;
	wire _w18858_ ;
	wire _w18859_ ;
	wire _w18860_ ;
	wire _w18861_ ;
	wire _w18862_ ;
	wire _w18863_ ;
	wire _w18864_ ;
	wire _w18865_ ;
	wire _w18866_ ;
	wire _w18867_ ;
	wire _w18868_ ;
	wire _w18869_ ;
	wire _w18870_ ;
	wire _w18871_ ;
	wire _w18872_ ;
	wire _w18873_ ;
	wire _w18874_ ;
	wire _w18875_ ;
	wire _w18876_ ;
	wire _w18877_ ;
	wire _w18878_ ;
	wire _w18879_ ;
	wire _w18880_ ;
	wire _w18881_ ;
	wire _w18882_ ;
	wire _w18883_ ;
	wire _w18884_ ;
	wire _w18885_ ;
	wire _w18886_ ;
	wire _w18887_ ;
	wire _w18888_ ;
	wire _w18889_ ;
	wire _w18890_ ;
	wire _w18891_ ;
	wire _w18892_ ;
	wire _w18893_ ;
	wire _w18894_ ;
	wire _w18895_ ;
	wire _w18896_ ;
	wire _w18897_ ;
	wire _w18898_ ;
	wire _w18899_ ;
	wire _w18900_ ;
	wire _w18901_ ;
	wire _w18902_ ;
	wire _w18903_ ;
	wire _w18904_ ;
	wire _w18905_ ;
	wire _w18906_ ;
	wire _w18907_ ;
	wire _w18908_ ;
	wire _w18909_ ;
	wire _w18910_ ;
	wire _w18911_ ;
	wire _w18912_ ;
	wire _w18913_ ;
	wire _w18914_ ;
	wire _w18915_ ;
	wire _w18916_ ;
	wire _w18917_ ;
	wire _w18918_ ;
	wire _w18919_ ;
	wire _w18920_ ;
	wire _w18921_ ;
	wire _w18922_ ;
	wire _w18923_ ;
	wire _w18924_ ;
	wire _w18925_ ;
	wire _w18926_ ;
	wire _w18927_ ;
	wire _w18928_ ;
	wire _w18929_ ;
	wire _w18930_ ;
	wire _w18931_ ;
	wire _w18932_ ;
	wire _w18933_ ;
	wire _w18934_ ;
	wire _w18935_ ;
	wire _w18936_ ;
	wire _w18937_ ;
	wire _w18938_ ;
	wire _w18939_ ;
	wire _w18940_ ;
	wire _w18941_ ;
	wire _w18942_ ;
	wire _w18943_ ;
	wire _w18944_ ;
	wire _w18945_ ;
	wire _w18946_ ;
	wire _w18947_ ;
	wire _w18948_ ;
	wire _w18949_ ;
	wire _w18950_ ;
	wire _w18951_ ;
	wire _w18952_ ;
	wire _w18953_ ;
	wire _w18954_ ;
	wire _w18955_ ;
	wire _w18956_ ;
	wire _w18957_ ;
	wire _w18958_ ;
	wire _w18959_ ;
	wire _w18960_ ;
	wire _w18961_ ;
	wire _w18962_ ;
	wire _w18963_ ;
	wire _w18964_ ;
	wire _w18965_ ;
	wire _w18966_ ;
	wire _w18967_ ;
	wire _w18968_ ;
	wire _w18969_ ;
	wire _w18970_ ;
	wire _w18971_ ;
	wire _w18972_ ;
	wire _w18973_ ;
	wire _w18974_ ;
	wire _w18975_ ;
	wire _w18976_ ;
	wire _w18977_ ;
	wire _w18978_ ;
	wire _w18979_ ;
	wire _w18980_ ;
	wire _w18981_ ;
	wire _w18982_ ;
	wire _w18983_ ;
	wire _w18984_ ;
	wire _w18985_ ;
	wire _w18986_ ;
	wire _w18987_ ;
	wire _w18988_ ;
	wire _w18989_ ;
	wire _w18990_ ;
	wire _w18991_ ;
	wire _w18992_ ;
	wire _w18993_ ;
	wire _w18994_ ;
	wire _w18995_ ;
	wire _w18996_ ;
	wire _w18997_ ;
	wire _w18998_ ;
	wire _w18999_ ;
	wire _w19000_ ;
	wire _w19001_ ;
	wire _w19002_ ;
	wire _w19003_ ;
	wire _w19004_ ;
	wire _w19005_ ;
	wire _w19006_ ;
	wire _w19007_ ;
	wire _w19008_ ;
	wire _w19009_ ;
	wire _w19010_ ;
	wire _w19011_ ;
	wire _w19012_ ;
	wire _w19013_ ;
	wire _w19014_ ;
	wire _w19015_ ;
	wire _w19016_ ;
	wire _w19017_ ;
	wire _w19018_ ;
	wire _w19019_ ;
	wire _w19020_ ;
	wire _w19021_ ;
	wire _w19022_ ;
	wire _w19023_ ;
	wire _w19024_ ;
	wire _w19025_ ;
	wire _w19026_ ;
	wire _w19027_ ;
	wire _w19028_ ;
	wire _w19029_ ;
	wire _w19030_ ;
	wire _w19031_ ;
	wire _w19032_ ;
	wire _w19033_ ;
	wire _w19034_ ;
	wire _w19035_ ;
	wire _w19036_ ;
	wire _w19037_ ;
	wire _w19038_ ;
	wire _w19039_ ;
	wire _w19040_ ;
	wire _w19041_ ;
	wire _w19042_ ;
	wire _w19043_ ;
	wire _w19044_ ;
	wire _w19045_ ;
	wire _w19046_ ;
	wire _w19047_ ;
	wire _w19048_ ;
	wire _w19049_ ;
	wire _w19050_ ;
	wire _w19051_ ;
	wire _w19052_ ;
	wire _w19053_ ;
	wire _w19054_ ;
	wire _w19055_ ;
	wire _w19056_ ;
	wire _w19057_ ;
	wire _w19058_ ;
	wire _w19059_ ;
	wire _w19060_ ;
	wire _w19061_ ;
	wire _w19062_ ;
	wire _w19063_ ;
	wire _w19064_ ;
	wire _w19065_ ;
	wire _w19066_ ;
	wire _w19067_ ;
	wire _w19068_ ;
	wire _w19069_ ;
	wire _w19070_ ;
	wire _w19071_ ;
	wire _w19072_ ;
	wire _w19073_ ;
	wire _w19074_ ;
	wire _w19075_ ;
	wire _w19076_ ;
	wire _w19077_ ;
	wire _w19078_ ;
	wire _w19079_ ;
	wire _w19080_ ;
	wire _w19081_ ;
	wire _w19082_ ;
	wire _w19083_ ;
	wire _w19084_ ;
	wire _w19085_ ;
	wire _w19086_ ;
	wire _w19087_ ;
	wire _w19088_ ;
	wire _w19089_ ;
	wire _w19090_ ;
	wire _w19091_ ;
	wire _w19092_ ;
	wire _w19093_ ;
	wire _w19094_ ;
	wire _w19095_ ;
	wire _w19096_ ;
	wire _w19097_ ;
	wire _w19098_ ;
	wire _w19099_ ;
	wire _w19100_ ;
	wire _w19101_ ;
	wire _w19102_ ;
	wire _w19103_ ;
	wire _w19104_ ;
	wire _w19105_ ;
	wire _w19106_ ;
	wire _w19107_ ;
	wire _w19108_ ;
	wire _w19109_ ;
	wire _w19110_ ;
	wire _w19111_ ;
	wire _w19112_ ;
	wire _w19113_ ;
	wire _w19114_ ;
	wire _w19115_ ;
	wire _w19116_ ;
	wire _w19117_ ;
	wire _w19118_ ;
	wire _w19119_ ;
	wire _w19120_ ;
	wire _w19121_ ;
	wire _w19122_ ;
	wire _w19123_ ;
	wire _w19124_ ;
	wire _w19125_ ;
	wire _w19126_ ;
	wire _w19127_ ;
	wire _w19128_ ;
	wire _w19129_ ;
	wire _w19130_ ;
	wire _w19131_ ;
	wire _w19132_ ;
	wire _w19133_ ;
	wire _w19134_ ;
	wire _w19135_ ;
	wire _w19136_ ;
	wire _w19137_ ;
	wire _w19138_ ;
	wire _w19139_ ;
	wire _w19140_ ;
	wire _w19141_ ;
	wire _w19142_ ;
	wire _w19143_ ;
	wire _w19144_ ;
	wire _w19145_ ;
	wire _w19146_ ;
	wire _w19147_ ;
	wire _w19148_ ;
	wire _w19149_ ;
	wire _w19150_ ;
	wire _w19151_ ;
	wire _w19152_ ;
	wire _w19153_ ;
	wire _w19154_ ;
	wire _w19155_ ;
	wire _w19156_ ;
	wire _w19157_ ;
	wire _w19158_ ;
	wire _w19159_ ;
	wire _w19160_ ;
	wire _w19161_ ;
	wire _w19162_ ;
	wire _w19163_ ;
	wire _w19164_ ;
	wire _w19165_ ;
	wire _w19166_ ;
	wire _w19167_ ;
	wire _w19168_ ;
	wire _w19169_ ;
	wire _w19170_ ;
	wire _w19171_ ;
	wire _w19172_ ;
	wire _w19173_ ;
	wire _w19174_ ;
	wire _w19175_ ;
	wire _w19176_ ;
	wire _w19177_ ;
	wire _w19178_ ;
	wire _w19179_ ;
	wire _w19180_ ;
	wire _w19181_ ;
	wire _w19182_ ;
	wire _w19183_ ;
	wire _w19184_ ;
	wire _w19185_ ;
	wire _w19186_ ;
	wire _w19187_ ;
	wire _w19188_ ;
	wire _w19189_ ;
	wire _w19190_ ;
	wire _w19191_ ;
	wire _w19192_ ;
	wire _w19193_ ;
	wire _w19194_ ;
	wire _w19195_ ;
	wire _w19196_ ;
	wire _w19197_ ;
	wire _w19198_ ;
	wire _w19199_ ;
	wire _w19200_ ;
	wire _w19201_ ;
	wire _w19202_ ;
	wire _w19203_ ;
	wire _w19204_ ;
	wire _w19205_ ;
	wire _w19206_ ;
	wire _w19207_ ;
	wire _w19208_ ;
	wire _w19209_ ;
	wire _w19210_ ;
	wire _w19211_ ;
	wire _w19212_ ;
	wire _w19213_ ;
	wire _w19214_ ;
	wire _w19215_ ;
	wire _w19216_ ;
	wire _w19217_ ;
	wire _w19218_ ;
	wire _w19219_ ;
	wire _w19220_ ;
	wire _w19221_ ;
	wire _w19222_ ;
	wire _w19223_ ;
	wire _w19224_ ;
	wire _w19225_ ;
	wire _w19226_ ;
	wire _w19227_ ;
	wire _w19228_ ;
	wire _w19229_ ;
	wire _w19230_ ;
	wire _w19231_ ;
	wire _w19232_ ;
	wire _w19233_ ;
	wire _w19234_ ;
	wire _w19235_ ;
	wire _w19236_ ;
	wire _w19237_ ;
	wire _w19238_ ;
	wire _w19239_ ;
	wire _w19240_ ;
	wire _w19241_ ;
	wire _w19242_ ;
	wire _w19243_ ;
	wire _w19244_ ;
	wire _w19245_ ;
	wire _w19246_ ;
	wire _w19247_ ;
	wire _w19248_ ;
	wire _w19249_ ;
	wire _w19250_ ;
	wire _w19251_ ;
	wire _w19252_ ;
	wire _w19253_ ;
	wire _w19254_ ;
	wire _w19255_ ;
	wire _w19256_ ;
	wire _w19257_ ;
	wire _w19258_ ;
	wire _w19259_ ;
	wire _w19260_ ;
	wire _w19261_ ;
	wire _w19262_ ;
	wire _w19263_ ;
	wire _w19264_ ;
	wire _w19265_ ;
	wire _w19266_ ;
	wire _w19267_ ;
	wire _w19268_ ;
	wire _w19269_ ;
	wire _w19270_ ;
	wire _w19271_ ;
	wire _w19272_ ;
	wire _w19273_ ;
	wire _w19274_ ;
	wire _w19275_ ;
	wire _w19276_ ;
	wire _w19277_ ;
	wire _w19278_ ;
	wire _w19279_ ;
	wire _w19280_ ;
	wire _w19281_ ;
	wire _w19282_ ;
	wire _w19283_ ;
	wire _w19284_ ;
	wire _w19285_ ;
	wire _w19286_ ;
	wire _w19287_ ;
	wire _w19288_ ;
	wire _w19289_ ;
	wire _w19290_ ;
	wire _w19291_ ;
	wire _w19292_ ;
	wire _w19293_ ;
	wire _w19294_ ;
	wire _w19295_ ;
	wire _w19296_ ;
	wire _w19297_ ;
	wire _w19298_ ;
	wire _w19299_ ;
	wire _w19300_ ;
	wire _w19301_ ;
	wire _w19302_ ;
	wire _w19303_ ;
	wire _w19304_ ;
	wire _w19305_ ;
	wire _w19306_ ;
	wire _w19307_ ;
	wire _w19308_ ;
	wire _w19309_ ;
	wire _w19310_ ;
	wire _w19311_ ;
	wire _w19312_ ;
	wire _w19313_ ;
	wire _w19314_ ;
	wire _w19315_ ;
	wire _w19316_ ;
	wire _w19317_ ;
	wire _w19318_ ;
	wire _w19319_ ;
	wire _w19320_ ;
	wire _w19321_ ;
	wire _w19322_ ;
	wire _w19323_ ;
	wire _w19324_ ;
	wire _w19325_ ;
	wire _w19326_ ;
	wire _w19327_ ;
	wire _w19328_ ;
	wire _w19329_ ;
	wire _w19330_ ;
	wire _w19331_ ;
	wire _w19332_ ;
	wire _w19333_ ;
	wire _w19334_ ;
	wire _w19335_ ;
	wire _w19336_ ;
	wire _w19337_ ;
	wire _w19338_ ;
	wire _w19339_ ;
	wire _w19340_ ;
	wire _w19341_ ;
	wire _w19342_ ;
	wire _w19343_ ;
	wire _w19344_ ;
	wire _w19345_ ;
	wire _w19346_ ;
	wire _w19347_ ;
	wire _w19348_ ;
	wire _w19349_ ;
	wire _w19350_ ;
	wire _w19351_ ;
	wire _w19352_ ;
	wire _w19353_ ;
	wire _w19354_ ;
	wire _w19355_ ;
	wire _w19356_ ;
	wire _w19357_ ;
	wire _w19358_ ;
	wire _w19359_ ;
	wire _w19360_ ;
	wire _w19361_ ;
	wire _w19362_ ;
	wire _w19363_ ;
	wire _w19364_ ;
	wire _w19365_ ;
	wire _w19366_ ;
	wire _w19367_ ;
	wire _w19368_ ;
	wire _w19369_ ;
	wire _w19370_ ;
	wire _w19371_ ;
	wire _w19372_ ;
	wire _w19373_ ;
	wire _w19374_ ;
	wire _w19375_ ;
	wire _w19376_ ;
	wire _w19377_ ;
	wire _w19378_ ;
	wire _w19379_ ;
	wire _w19380_ ;
	wire _w19381_ ;
	wire _w19382_ ;
	wire _w19383_ ;
	wire _w19384_ ;
	wire _w19385_ ;
	wire _w19386_ ;
	wire _w19387_ ;
	wire _w19388_ ;
	wire _w19389_ ;
	wire _w19390_ ;
	wire _w19391_ ;
	wire _w19392_ ;
	wire _w19393_ ;
	wire _w19394_ ;
	wire _w19395_ ;
	wire _w19396_ ;
	wire _w19397_ ;
	wire _w19398_ ;
	wire _w19399_ ;
	wire _w19400_ ;
	wire _w19401_ ;
	wire _w19402_ ;
	wire _w19403_ ;
	wire _w19404_ ;
	wire _w19405_ ;
	wire _w19406_ ;
	wire _w19407_ ;
	wire _w19408_ ;
	wire _w19409_ ;
	wire _w19410_ ;
	wire _w19411_ ;
	wire _w19412_ ;
	wire _w19413_ ;
	wire _w19414_ ;
	wire _w19415_ ;
	wire _w19416_ ;
	wire _w19417_ ;
	wire _w19418_ ;
	wire _w19419_ ;
	wire _w19420_ ;
	wire _w19421_ ;
	wire _w19422_ ;
	wire _w19423_ ;
	wire _w19424_ ;
	wire _w19425_ ;
	wire _w19426_ ;
	wire _w19427_ ;
	wire _w19428_ ;
	wire _w19429_ ;
	wire _w19430_ ;
	wire _w19431_ ;
	wire _w19432_ ;
	wire _w19433_ ;
	wire _w19434_ ;
	wire _w19435_ ;
	wire _w19436_ ;
	wire _w19437_ ;
	wire _w19438_ ;
	wire _w19439_ ;
	wire _w19440_ ;
	wire _w19441_ ;
	wire _w19442_ ;
	wire _w19443_ ;
	wire _w19444_ ;
	wire _w19445_ ;
	wire _w19446_ ;
	wire _w19447_ ;
	wire _w19448_ ;
	wire _w19449_ ;
	wire _w19450_ ;
	wire _w19451_ ;
	wire _w19452_ ;
	wire _w19453_ ;
	wire _w19454_ ;
	wire _w19455_ ;
	wire _w19456_ ;
	wire _w19457_ ;
	wire _w19458_ ;
	wire _w19459_ ;
	wire _w19460_ ;
	wire _w19461_ ;
	wire _w19462_ ;
	wire _w19463_ ;
	wire _w19464_ ;
	wire _w19465_ ;
	wire _w19466_ ;
	wire _w19467_ ;
	wire _w19468_ ;
	wire _w19469_ ;
	wire _w19470_ ;
	wire _w19471_ ;
	wire _w19472_ ;
	wire _w19473_ ;
	wire _w19474_ ;
	wire _w19475_ ;
	wire _w19476_ ;
	wire _w19477_ ;
	wire _w19478_ ;
	wire _w19479_ ;
	wire _w19480_ ;
	wire _w19481_ ;
	wire _w19482_ ;
	wire _w19483_ ;
	wire _w19484_ ;
	wire _w19485_ ;
	wire _w19486_ ;
	wire _w19487_ ;
	wire _w19488_ ;
	wire _w19489_ ;
	wire _w19490_ ;
	wire _w19491_ ;
	wire _w19492_ ;
	wire _w19493_ ;
	wire _w19494_ ;
	wire _w19495_ ;
	wire _w19496_ ;
	wire _w19497_ ;
	wire _w19498_ ;
	wire _w19499_ ;
	wire _w19500_ ;
	wire _w19501_ ;
	wire _w19502_ ;
	wire _w19503_ ;
	wire _w19504_ ;
	wire _w19505_ ;
	wire _w19506_ ;
	wire _w19507_ ;
	wire _w19508_ ;
	wire _w19509_ ;
	wire _w19510_ ;
	wire _w19511_ ;
	wire _w19512_ ;
	wire _w19513_ ;
	wire _w19514_ ;
	wire _w19515_ ;
	wire _w19516_ ;
	wire _w19517_ ;
	wire _w19518_ ;
	wire _w19519_ ;
	wire _w19520_ ;
	wire _w19521_ ;
	wire _w19522_ ;
	wire _w19523_ ;
	wire _w19524_ ;
	wire _w19525_ ;
	wire _w19526_ ;
	wire _w19527_ ;
	wire _w19528_ ;
	wire _w19529_ ;
	wire _w19530_ ;
	wire _w19531_ ;
	wire _w19532_ ;
	wire _w19533_ ;
	wire _w19534_ ;
	wire _w19535_ ;
	wire _w19536_ ;
	wire _w19537_ ;
	wire _w19538_ ;
	wire _w19539_ ;
	wire _w19540_ ;
	wire _w19541_ ;
	wire _w19542_ ;
	wire _w19543_ ;
	wire _w19544_ ;
	wire _w19545_ ;
	wire _w19546_ ;
	wire _w19547_ ;
	wire _w19548_ ;
	wire _w19549_ ;
	wire _w19550_ ;
	wire _w19551_ ;
	wire _w19552_ ;
	wire _w19553_ ;
	wire _w19554_ ;
	wire _w19555_ ;
	wire _w19556_ ;
	wire _w19557_ ;
	wire _w19558_ ;
	wire _w19559_ ;
	wire _w19560_ ;
	wire _w19561_ ;
	wire _w19562_ ;
	wire _w19563_ ;
	wire _w19564_ ;
	wire _w19565_ ;
	wire _w19566_ ;
	wire _w19567_ ;
	wire _w19568_ ;
	wire _w19569_ ;
	wire _w19570_ ;
	wire _w19571_ ;
	wire _w19572_ ;
	wire _w19573_ ;
	wire _w19574_ ;
	wire _w19575_ ;
	wire _w19576_ ;
	wire _w19577_ ;
	wire _w19578_ ;
	wire _w19579_ ;
	wire _w19580_ ;
	wire _w19581_ ;
	wire _w19582_ ;
	wire _w19583_ ;
	wire _w19584_ ;
	wire _w19585_ ;
	wire _w19586_ ;
	wire _w19587_ ;
	wire _w19588_ ;
	wire _w19589_ ;
	wire _w19590_ ;
	wire _w19591_ ;
	wire _w19592_ ;
	wire _w19593_ ;
	wire _w19594_ ;
	wire _w19595_ ;
	wire _w19596_ ;
	wire _w19597_ ;
	wire _w19598_ ;
	wire _w19599_ ;
	wire _w19600_ ;
	wire _w19601_ ;
	wire _w19602_ ;
	wire _w19603_ ;
	wire _w19604_ ;
	wire _w19605_ ;
	wire _w19606_ ;
	wire _w19607_ ;
	wire _w19608_ ;
	wire _w19609_ ;
	wire _w19610_ ;
	wire _w19611_ ;
	wire _w19612_ ;
	wire _w19613_ ;
	wire _w19614_ ;
	wire _w19615_ ;
	wire _w19616_ ;
	wire _w19617_ ;
	wire _w19618_ ;
	wire _w19619_ ;
	wire _w19620_ ;
	wire _w19621_ ;
	wire _w19622_ ;
	wire _w19623_ ;
	wire _w19624_ ;
	wire _w19625_ ;
	wire _w19626_ ;
	wire _w19627_ ;
	wire _w19628_ ;
	wire _w19629_ ;
	wire _w19630_ ;
	wire _w19631_ ;
	wire _w19632_ ;
	wire _w19633_ ;
	wire _w19634_ ;
	wire _w19635_ ;
	wire _w19636_ ;
	wire _w19637_ ;
	wire _w19638_ ;
	wire _w19639_ ;
	wire _w19640_ ;
	wire _w19641_ ;
	wire _w19642_ ;
	wire _w19643_ ;
	wire _w19644_ ;
	wire _w19645_ ;
	wire _w19646_ ;
	wire _w19647_ ;
	wire _w19648_ ;
	wire _w19649_ ;
	wire _w19650_ ;
	wire _w19651_ ;
	wire _w19652_ ;
	wire _w19653_ ;
	wire _w19654_ ;
	wire _w19655_ ;
	wire _w19656_ ;
	wire _w19657_ ;
	wire _w19658_ ;
	wire _w19659_ ;
	wire _w19660_ ;
	wire _w19661_ ;
	wire _w19662_ ;
	wire _w19663_ ;
	wire _w19664_ ;
	wire _w19665_ ;
	wire _w19666_ ;
	wire _w19667_ ;
	wire _w19668_ ;
	wire _w19669_ ;
	wire _w19670_ ;
	wire _w19671_ ;
	wire _w19672_ ;
	wire _w19673_ ;
	wire _w19674_ ;
	wire _w19675_ ;
	wire _w19676_ ;
	wire _w19677_ ;
	wire _w19678_ ;
	wire _w19679_ ;
	wire _w19680_ ;
	wire _w19681_ ;
	wire _w19682_ ;
	wire _w19683_ ;
	wire _w19684_ ;
	wire _w19685_ ;
	wire _w19686_ ;
	wire _w19687_ ;
	wire _w19688_ ;
	wire _w19689_ ;
	wire _w19690_ ;
	wire _w19691_ ;
	wire _w19692_ ;
	wire _w19693_ ;
	wire _w19694_ ;
	wire _w19695_ ;
	wire _w19696_ ;
	wire _w19697_ ;
	wire _w19698_ ;
	wire _w19699_ ;
	wire _w19700_ ;
	wire _w19701_ ;
	wire _w19702_ ;
	wire _w19703_ ;
	wire _w19704_ ;
	wire _w19705_ ;
	wire _w19706_ ;
	wire _w19707_ ;
	wire _w19708_ ;
	wire _w19709_ ;
	wire _w19710_ ;
	wire _w19711_ ;
	wire _w19712_ ;
	wire _w19713_ ;
	wire _w19714_ ;
	wire _w19715_ ;
	wire _w19716_ ;
	wire _w19717_ ;
	wire _w19718_ ;
	wire _w19719_ ;
	wire _w19720_ ;
	wire _w19721_ ;
	wire _w19722_ ;
	wire _w19723_ ;
	wire _w19724_ ;
	wire _w19725_ ;
	wire _w19726_ ;
	wire _w19727_ ;
	wire _w19728_ ;
	wire _w19729_ ;
	wire _w19730_ ;
	wire _w19731_ ;
	wire _w19732_ ;
	wire _w19733_ ;
	wire _w19734_ ;
	wire _w19735_ ;
	wire _w19736_ ;
	wire _w19737_ ;
	wire _w19738_ ;
	wire _w19739_ ;
	wire _w19740_ ;
	wire _w19741_ ;
	wire _w19742_ ;
	wire _w19743_ ;
	wire _w19744_ ;
	wire _w19745_ ;
	wire _w19746_ ;
	wire _w19747_ ;
	wire _w19748_ ;
	wire _w19749_ ;
	wire _w19750_ ;
	wire _w19751_ ;
	wire _w19752_ ;
	wire _w19753_ ;
	wire _w19754_ ;
	wire _w19755_ ;
	wire _w19756_ ;
	wire _w19757_ ;
	wire _w19758_ ;
	wire _w19759_ ;
	wire _w19760_ ;
	wire _w19761_ ;
	wire _w19762_ ;
	wire _w19763_ ;
	wire _w19764_ ;
	wire _w19765_ ;
	wire _w19766_ ;
	wire _w19767_ ;
	wire _w19768_ ;
	wire _w19769_ ;
	wire _w19770_ ;
	wire _w19771_ ;
	wire _w19772_ ;
	wire _w19773_ ;
	wire _w19774_ ;
	wire _w19775_ ;
	wire _w19776_ ;
	wire _w19777_ ;
	wire _w19778_ ;
	wire _w19779_ ;
	wire _w19780_ ;
	wire _w19781_ ;
	wire _w19782_ ;
	wire _w19783_ ;
	wire _w19784_ ;
	wire _w19785_ ;
	wire _w19786_ ;
	wire _w19787_ ;
	wire _w19788_ ;
	wire _w19789_ ;
	wire _w19790_ ;
	wire _w19791_ ;
	wire _w19792_ ;
	wire _w19793_ ;
	wire _w19794_ ;
	wire _w19795_ ;
	wire _w19796_ ;
	wire _w19797_ ;
	wire _w19798_ ;
	wire _w19799_ ;
	wire _w19800_ ;
	wire _w19801_ ;
	wire _w19802_ ;
	wire _w19803_ ;
	wire _w19804_ ;
	wire _w19805_ ;
	wire _w19806_ ;
	wire _w19807_ ;
	wire _w19808_ ;
	wire _w19809_ ;
	wire _w19810_ ;
	wire _w19811_ ;
	wire _w19812_ ;
	wire _w19813_ ;
	wire _w19814_ ;
	wire _w19815_ ;
	wire _w19816_ ;
	wire _w19817_ ;
	wire _w19818_ ;
	wire _w19819_ ;
	wire _w19820_ ;
	wire _w19821_ ;
	wire _w19822_ ;
	wire _w19823_ ;
	wire _w19824_ ;
	wire _w19825_ ;
	wire _w19826_ ;
	wire _w19827_ ;
	wire _w19828_ ;
	wire _w19829_ ;
	wire _w19830_ ;
	wire _w19831_ ;
	wire _w19832_ ;
	wire _w19833_ ;
	wire _w19834_ ;
	wire _w19835_ ;
	wire _w19836_ ;
	wire _w19837_ ;
	wire _w19838_ ;
	wire _w19839_ ;
	wire _w19840_ ;
	wire _w19841_ ;
	wire _w19842_ ;
	wire _w19843_ ;
	wire _w19844_ ;
	wire _w19845_ ;
	wire _w19846_ ;
	wire _w19847_ ;
	wire _w19848_ ;
	wire _w19849_ ;
	wire _w19850_ ;
	wire _w19851_ ;
	wire _w19852_ ;
	wire _w19853_ ;
	wire _w19854_ ;
	wire _w19855_ ;
	wire _w19856_ ;
	wire _w19857_ ;
	wire _w19858_ ;
	wire _w19859_ ;
	wire _w19860_ ;
	wire _w19861_ ;
	wire _w19862_ ;
	wire _w19863_ ;
	wire _w19864_ ;
	wire _w19865_ ;
	wire _w19866_ ;
	wire _w19867_ ;
	wire _w19868_ ;
	wire _w19869_ ;
	wire _w19870_ ;
	wire _w19871_ ;
	wire _w19872_ ;
	wire _w19873_ ;
	wire _w19874_ ;
	wire _w19875_ ;
	wire _w19876_ ;
	wire _w19877_ ;
	wire _w19878_ ;
	wire _w19879_ ;
	wire _w19880_ ;
	wire _w19881_ ;
	wire _w19882_ ;
	wire _w19883_ ;
	wire _w19884_ ;
	wire _w19885_ ;
	wire _w19886_ ;
	wire _w19887_ ;
	wire _w19888_ ;
	wire _w19889_ ;
	wire _w19890_ ;
	wire _w19891_ ;
	wire _w19892_ ;
	wire _w19893_ ;
	wire _w19894_ ;
	wire _w19895_ ;
	wire _w19896_ ;
	wire _w19897_ ;
	wire _w19898_ ;
	wire _w19899_ ;
	wire _w19900_ ;
	wire _w19901_ ;
	wire _w19902_ ;
	wire _w19903_ ;
	wire _w19904_ ;
	wire _w19905_ ;
	wire _w19906_ ;
	wire _w19907_ ;
	wire _w19908_ ;
	wire _w19909_ ;
	wire _w19910_ ;
	wire _w19911_ ;
	wire _w19912_ ;
	wire _w19913_ ;
	wire _w19914_ ;
	wire _w19915_ ;
	wire _w19916_ ;
	wire _w19917_ ;
	wire _w19918_ ;
	wire _w19919_ ;
	wire _w19920_ ;
	wire _w19921_ ;
	wire _w19922_ ;
	wire _w19923_ ;
	wire _w19924_ ;
	wire _w19925_ ;
	wire _w19926_ ;
	wire _w19927_ ;
	wire _w19928_ ;
	wire _w19929_ ;
	wire _w19930_ ;
	wire _w19931_ ;
	wire _w19932_ ;
	wire _w19933_ ;
	wire _w19934_ ;
	wire _w19935_ ;
	wire _w19936_ ;
	wire _w19937_ ;
	wire _w19938_ ;
	wire _w19939_ ;
	wire _w19940_ ;
	wire _w19941_ ;
	wire _w19942_ ;
	wire _w19943_ ;
	wire _w19944_ ;
	wire _w19945_ ;
	wire _w19946_ ;
	wire _w19947_ ;
	wire _w19948_ ;
	wire _w19949_ ;
	wire _w19950_ ;
	wire _w19951_ ;
	wire _w19952_ ;
	wire _w19953_ ;
	wire _w19954_ ;
	wire _w19955_ ;
	wire _w19956_ ;
	wire _w19957_ ;
	wire _w19958_ ;
	wire _w19959_ ;
	wire _w19960_ ;
	wire _w19961_ ;
	wire _w19962_ ;
	wire _w19963_ ;
	wire _w19964_ ;
	wire _w19965_ ;
	wire _w19966_ ;
	wire _w19967_ ;
	wire _w19968_ ;
	wire _w19969_ ;
	wire _w19970_ ;
	wire _w19971_ ;
	wire _w19972_ ;
	wire _w19973_ ;
	wire _w19974_ ;
	wire _w19975_ ;
	wire _w19976_ ;
	wire _w19977_ ;
	wire _w19978_ ;
	wire _w19979_ ;
	wire _w19980_ ;
	wire _w19981_ ;
	wire _w19982_ ;
	wire _w19983_ ;
	wire _w19984_ ;
	wire _w19985_ ;
	wire _w19986_ ;
	wire _w19987_ ;
	wire _w19988_ ;
	wire _w19989_ ;
	wire _w19990_ ;
	wire _w19991_ ;
	wire _w19992_ ;
	wire _w19993_ ;
	wire _w19994_ ;
	wire _w19995_ ;
	wire _w19996_ ;
	wire _w19997_ ;
	wire _w19998_ ;
	wire _w19999_ ;
	wire _w20000_ ;
	wire _w20001_ ;
	wire _w20002_ ;
	wire _w20003_ ;
	wire _w20004_ ;
	wire _w20005_ ;
	wire _w20006_ ;
	wire _w20007_ ;
	wire _w20008_ ;
	wire _w20009_ ;
	wire _w20010_ ;
	wire _w20011_ ;
	wire _w20012_ ;
	wire _w20013_ ;
	wire _w20014_ ;
	wire _w20015_ ;
	wire _w20016_ ;
	wire _w20017_ ;
	wire _w20018_ ;
	wire _w20019_ ;
	wire _w20020_ ;
	wire _w20021_ ;
	wire _w20022_ ;
	wire _w20023_ ;
	wire _w20024_ ;
	wire _w20025_ ;
	wire _w20026_ ;
	wire _w20027_ ;
	wire _w20028_ ;
	wire _w20029_ ;
	wire _w20030_ ;
	wire _w20031_ ;
	wire _w20032_ ;
	wire _w20033_ ;
	wire _w20034_ ;
	wire _w20035_ ;
	wire _w20036_ ;
	wire _w20037_ ;
	wire _w20038_ ;
	wire _w20039_ ;
	wire _w20040_ ;
	wire _w20041_ ;
	wire _w20042_ ;
	wire _w20043_ ;
	wire _w20044_ ;
	wire _w20045_ ;
	wire _w20046_ ;
	wire _w20047_ ;
	wire _w20048_ ;
	wire _w20049_ ;
	wire _w20050_ ;
	wire _w20051_ ;
	wire _w20052_ ;
	wire _w20053_ ;
	wire _w20054_ ;
	wire _w20055_ ;
	wire _w20056_ ;
	wire _w20057_ ;
	wire _w20058_ ;
	wire _w20059_ ;
	wire _w20060_ ;
	wire _w20061_ ;
	wire _w20062_ ;
	wire _w20063_ ;
	wire _w20064_ ;
	wire _w20065_ ;
	wire _w20066_ ;
	wire _w20067_ ;
	wire _w20068_ ;
	wire _w20069_ ;
	wire _w20070_ ;
	wire _w20071_ ;
	wire _w20072_ ;
	wire _w20073_ ;
	wire _w20074_ ;
	wire _w20075_ ;
	wire _w20076_ ;
	wire _w20077_ ;
	wire _w20078_ ;
	wire _w20079_ ;
	wire _w20080_ ;
	wire _w20081_ ;
	wire _w20082_ ;
	wire _w20083_ ;
	wire _w20084_ ;
	wire _w20085_ ;
	wire _w20086_ ;
	wire _w20087_ ;
	wire _w20088_ ;
	wire _w20089_ ;
	wire _w20090_ ;
	wire _w20091_ ;
	wire _w20092_ ;
	wire _w20093_ ;
	wire _w20094_ ;
	wire _w20095_ ;
	wire _w20096_ ;
	wire _w20097_ ;
	wire _w20098_ ;
	wire _w20099_ ;
	wire _w20100_ ;
	wire _w20101_ ;
	wire _w20102_ ;
	wire _w20103_ ;
	wire _w20104_ ;
	wire _w20105_ ;
	wire _w20106_ ;
	wire _w20107_ ;
	wire _w20108_ ;
	wire _w20109_ ;
	wire _w20110_ ;
	wire _w20111_ ;
	wire _w20112_ ;
	wire _w20113_ ;
	wire _w20114_ ;
	wire _w20115_ ;
	wire _w20116_ ;
	wire _w20117_ ;
	wire _w20118_ ;
	wire _w20119_ ;
	wire _w20120_ ;
	wire _w20121_ ;
	wire _w20122_ ;
	wire _w20123_ ;
	wire _w20124_ ;
	wire _w20125_ ;
	wire _w20126_ ;
	wire _w20127_ ;
	wire _w20128_ ;
	wire _w20129_ ;
	wire _w20130_ ;
	wire _w20131_ ;
	wire _w20132_ ;
	wire _w20133_ ;
	wire _w20134_ ;
	wire _w20135_ ;
	wire _w20136_ ;
	wire _w20137_ ;
	wire _w20138_ ;
	wire _w20139_ ;
	wire _w20140_ ;
	wire _w20141_ ;
	wire _w20142_ ;
	wire _w20143_ ;
	wire _w20144_ ;
	wire _w20145_ ;
	wire _w20146_ ;
	wire _w20147_ ;
	wire _w20148_ ;
	wire _w20149_ ;
	wire _w20150_ ;
	wire _w20151_ ;
	wire _w20152_ ;
	wire _w20153_ ;
	wire _w20154_ ;
	wire _w20155_ ;
	wire _w20156_ ;
	wire _w20157_ ;
	wire _w20158_ ;
	wire _w20159_ ;
	wire _w20160_ ;
	wire _w20161_ ;
	wire _w20162_ ;
	wire _w20163_ ;
	wire _w20164_ ;
	wire _w20165_ ;
	wire _w20166_ ;
	wire _w20167_ ;
	wire _w20168_ ;
	wire _w20169_ ;
	wire _w20170_ ;
	wire _w20171_ ;
	wire _w20172_ ;
	wire _w20173_ ;
	wire _w20174_ ;
	wire _w20175_ ;
	wire _w20176_ ;
	wire _w20177_ ;
	wire _w20178_ ;
	wire _w20179_ ;
	wire _w20180_ ;
	wire _w20181_ ;
	wire _w20182_ ;
	wire _w20183_ ;
	wire _w20184_ ;
	wire _w20185_ ;
	wire _w20186_ ;
	wire _w20187_ ;
	wire _w20188_ ;
	wire _w20189_ ;
	wire _w20190_ ;
	wire _w20191_ ;
	wire _w20192_ ;
	wire _w20193_ ;
	wire _w20194_ ;
	wire _w20195_ ;
	wire _w20196_ ;
	wire _w20197_ ;
	wire _w20198_ ;
	wire _w20199_ ;
	wire _w20200_ ;
	wire _w20201_ ;
	wire _w20202_ ;
	wire _w20203_ ;
	wire _w20204_ ;
	wire _w20205_ ;
	wire _w20206_ ;
	wire _w20207_ ;
	wire _w20208_ ;
	wire _w20209_ ;
	wire _w20210_ ;
	wire _w20211_ ;
	wire _w20212_ ;
	wire _w20213_ ;
	wire _w20214_ ;
	wire _w20215_ ;
	wire _w20216_ ;
	wire _w20217_ ;
	wire _w20218_ ;
	wire _w20219_ ;
	wire _w20220_ ;
	wire _w20221_ ;
	wire _w20222_ ;
	wire _w20223_ ;
	wire _w20224_ ;
	wire _w20225_ ;
	wire _w20226_ ;
	wire _w20227_ ;
	wire _w20228_ ;
	wire _w20229_ ;
	wire _w20230_ ;
	wire _w20231_ ;
	wire _w20232_ ;
	wire _w20233_ ;
	wire _w20234_ ;
	wire _w20235_ ;
	wire _w20236_ ;
	wire _w20237_ ;
	wire _w20238_ ;
	wire _w20239_ ;
	wire _w20240_ ;
	wire _w20241_ ;
	wire _w20242_ ;
	wire _w20243_ ;
	wire _w20244_ ;
	wire _w20245_ ;
	wire _w20246_ ;
	wire _w20247_ ;
	wire _w20248_ ;
	wire _w20249_ ;
	wire _w20250_ ;
	wire _w20251_ ;
	wire _w20252_ ;
	wire _w20253_ ;
	wire _w20254_ ;
	wire _w20255_ ;
	wire _w20256_ ;
	wire _w20257_ ;
	wire _w20258_ ;
	wire _w20259_ ;
	wire _w20260_ ;
	wire _w20261_ ;
	wire _w20262_ ;
	wire _w20263_ ;
	wire _w20264_ ;
	wire _w20265_ ;
	wire _w20266_ ;
	wire _w20267_ ;
	wire _w20268_ ;
	wire _w20269_ ;
	wire _w20270_ ;
	wire _w20271_ ;
	wire _w20272_ ;
	wire _w20273_ ;
	wire _w20274_ ;
	wire _w20275_ ;
	wire _w20276_ ;
	wire _w20277_ ;
	wire _w20278_ ;
	wire _w20279_ ;
	wire _w20280_ ;
	wire _w20281_ ;
	wire _w20282_ ;
	wire _w20283_ ;
	wire _w20284_ ;
	wire _w20285_ ;
	wire _w20286_ ;
	wire _w20287_ ;
	wire _w20288_ ;
	wire _w20289_ ;
	wire _w20290_ ;
	wire _w20291_ ;
	wire _w20292_ ;
	wire _w20293_ ;
	wire _w20294_ ;
	wire _w20295_ ;
	wire _w20296_ ;
	wire _w20297_ ;
	wire _w20298_ ;
	wire _w20299_ ;
	wire _w20300_ ;
	wire _w20301_ ;
	wire _w20302_ ;
	wire _w20303_ ;
	wire _w20304_ ;
	wire _w20305_ ;
	wire _w20306_ ;
	wire _w20307_ ;
	wire _w20308_ ;
	wire _w20309_ ;
	wire _w20310_ ;
	wire _w20311_ ;
	wire _w20312_ ;
	wire _w20313_ ;
	wire _w20314_ ;
	wire _w20315_ ;
	wire _w20316_ ;
	wire _w20317_ ;
	wire _w20318_ ;
	wire _w20319_ ;
	wire _w20320_ ;
	wire _w20321_ ;
	wire _w20322_ ;
	wire _w20323_ ;
	wire _w20324_ ;
	wire _w20325_ ;
	wire _w20326_ ;
	wire _w20327_ ;
	wire _w20328_ ;
	wire _w20329_ ;
	wire _w20330_ ;
	wire _w20331_ ;
	wire _w20332_ ;
	wire _w20333_ ;
	wire _w20334_ ;
	wire _w20335_ ;
	wire _w20336_ ;
	wire _w20337_ ;
	wire _w20338_ ;
	wire _w20339_ ;
	wire _w20340_ ;
	wire _w20341_ ;
	wire _w20342_ ;
	wire _w20343_ ;
	wire _w20344_ ;
	wire _w20345_ ;
	wire _w20346_ ;
	wire _w20347_ ;
	wire _w20348_ ;
	wire _w20349_ ;
	wire _w20350_ ;
	wire _w20351_ ;
	wire _w20352_ ;
	wire _w20353_ ;
	wire _w20354_ ;
	wire _w20355_ ;
	wire _w20356_ ;
	wire _w20357_ ;
	wire _w20358_ ;
	wire _w20359_ ;
	wire _w20360_ ;
	wire _w20361_ ;
	wire _w20362_ ;
	wire _w20363_ ;
	wire _w20364_ ;
	wire _w20365_ ;
	wire _w20366_ ;
	wire _w20367_ ;
	wire _w20368_ ;
	wire _w20369_ ;
	wire _w20370_ ;
	wire _w20371_ ;
	wire _w20372_ ;
	wire _w20373_ ;
	wire _w20374_ ;
	wire _w20375_ ;
	wire _w20376_ ;
	wire _w20377_ ;
	wire _w20378_ ;
	wire _w20379_ ;
	wire _w20380_ ;
	wire _w20381_ ;
	wire _w20382_ ;
	wire _w20383_ ;
	wire _w20384_ ;
	wire _w20385_ ;
	wire _w20386_ ;
	wire _w20387_ ;
	wire _w20388_ ;
	wire _w20389_ ;
	wire _w20390_ ;
	wire _w20391_ ;
	wire _w20392_ ;
	wire _w20393_ ;
	wire _w20394_ ;
	wire _w20395_ ;
	wire _w20396_ ;
	wire _w20397_ ;
	wire _w20398_ ;
	wire _w20399_ ;
	wire _w20400_ ;
	wire _w20401_ ;
	wire _w20402_ ;
	wire _w20403_ ;
	wire _w20404_ ;
	wire _w20405_ ;
	wire _w20406_ ;
	wire _w20407_ ;
	wire _w20408_ ;
	wire _w20409_ ;
	wire _w20410_ ;
	wire _w20411_ ;
	wire _w20412_ ;
	wire _w20413_ ;
	wire _w20414_ ;
	wire _w20415_ ;
	wire _w20416_ ;
	wire _w20417_ ;
	wire _w20418_ ;
	wire _w20419_ ;
	wire _w20420_ ;
	wire _w20421_ ;
	wire _w20422_ ;
	wire _w20423_ ;
	wire _w20424_ ;
	wire _w20425_ ;
	wire _w20426_ ;
	wire _w20427_ ;
	wire _w20428_ ;
	wire _w20429_ ;
	wire _w20430_ ;
	wire _w20431_ ;
	wire _w20432_ ;
	wire _w20433_ ;
	wire _w20434_ ;
	wire _w20435_ ;
	wire _w20436_ ;
	wire _w20437_ ;
	wire _w20438_ ;
	wire _w20439_ ;
	wire _w20440_ ;
	wire _w20441_ ;
	wire _w20442_ ;
	wire _w20443_ ;
	wire _w20444_ ;
	wire _w20445_ ;
	wire _w20446_ ;
	wire _w20447_ ;
	wire _w20448_ ;
	wire _w20449_ ;
	wire _w20450_ ;
	wire _w20451_ ;
	wire _w20452_ ;
	wire _w20453_ ;
	wire _w20454_ ;
	wire _w20455_ ;
	wire _w20456_ ;
	wire _w20457_ ;
	wire _w20458_ ;
	wire _w20459_ ;
	wire _w20460_ ;
	wire _w20461_ ;
	wire _w20462_ ;
	wire _w20463_ ;
	wire _w20464_ ;
	wire _w20465_ ;
	wire _w20466_ ;
	wire _w20467_ ;
	wire _w20468_ ;
	wire _w20469_ ;
	wire _w20470_ ;
	wire _w20471_ ;
	wire _w20472_ ;
	wire _w20473_ ;
	wire _w20474_ ;
	wire _w20475_ ;
	wire _w20476_ ;
	wire _w20477_ ;
	wire _w20478_ ;
	wire _w20479_ ;
	wire _w20480_ ;
	wire _w20481_ ;
	wire _w20482_ ;
	wire _w20483_ ;
	wire _w20484_ ;
	wire _w20485_ ;
	wire _w20486_ ;
	wire _w20487_ ;
	wire _w20488_ ;
	wire _w20489_ ;
	wire _w20490_ ;
	wire _w20491_ ;
	wire _w20492_ ;
	wire _w20493_ ;
	wire _w20494_ ;
	wire _w20495_ ;
	wire _w20496_ ;
	wire _w20497_ ;
	wire _w20498_ ;
	wire _w20499_ ;
	wire _w20500_ ;
	wire _w20501_ ;
	wire _w20502_ ;
	wire _w20503_ ;
	wire _w20504_ ;
	wire _w20505_ ;
	wire _w20506_ ;
	wire _w20507_ ;
	wire _w20508_ ;
	wire _w20509_ ;
	wire _w20510_ ;
	wire _w20511_ ;
	wire _w20512_ ;
	wire _w20513_ ;
	wire _w20514_ ;
	wire _w20515_ ;
	wire _w20516_ ;
	wire _w20517_ ;
	wire _w20518_ ;
	wire _w20519_ ;
	wire _w20520_ ;
	wire _w20521_ ;
	wire _w20522_ ;
	wire _w20523_ ;
	wire _w20524_ ;
	wire _w20525_ ;
	wire _w20526_ ;
	wire _w20527_ ;
	wire _w20528_ ;
	wire _w20529_ ;
	wire _w20530_ ;
	wire _w20531_ ;
	wire _w20532_ ;
	wire _w20533_ ;
	wire _w20534_ ;
	wire _w20535_ ;
	wire _w20536_ ;
	wire _w20537_ ;
	wire _w20538_ ;
	wire _w20539_ ;
	wire _w20540_ ;
	wire _w20541_ ;
	wire _w20542_ ;
	wire _w20543_ ;
	wire _w20544_ ;
	wire _w20545_ ;
	wire _w20546_ ;
	wire _w20547_ ;
	wire _w20548_ ;
	wire _w20549_ ;
	wire _w20550_ ;
	wire _w20551_ ;
	wire _w20552_ ;
	wire _w20553_ ;
	wire _w20554_ ;
	wire _w20555_ ;
	wire _w20556_ ;
	wire _w20557_ ;
	wire _w20558_ ;
	wire _w20559_ ;
	wire _w20560_ ;
	wire _w20561_ ;
	wire _w20562_ ;
	wire _w20563_ ;
	wire _w20564_ ;
	wire _w20565_ ;
	wire _w20566_ ;
	wire _w20567_ ;
	wire _w20568_ ;
	wire _w20569_ ;
	wire _w20570_ ;
	wire _w20571_ ;
	wire _w20572_ ;
	wire _w20573_ ;
	wire _w20574_ ;
	wire _w20575_ ;
	wire _w20576_ ;
	wire _w20577_ ;
	wire _w20578_ ;
	wire _w20579_ ;
	wire _w20580_ ;
	wire _w20581_ ;
	wire _w20582_ ;
	wire _w20583_ ;
	wire _w20584_ ;
	wire _w20585_ ;
	wire _w20586_ ;
	wire _w20587_ ;
	wire _w20588_ ;
	wire _w20589_ ;
	wire _w20590_ ;
	wire _w20591_ ;
	wire _w20592_ ;
	wire _w20593_ ;
	wire _w20594_ ;
	wire _w20595_ ;
	wire _w20596_ ;
	wire _w20597_ ;
	wire _w20598_ ;
	wire _w20599_ ;
	wire _w20600_ ;
	wire _w20601_ ;
	wire _w20602_ ;
	wire _w20603_ ;
	wire _w20604_ ;
	wire _w20605_ ;
	wire _w20606_ ;
	wire _w20607_ ;
	wire _w20608_ ;
	wire _w20609_ ;
	wire _w20610_ ;
	wire _w20611_ ;
	wire _w20612_ ;
	wire _w20613_ ;
	wire _w20614_ ;
	wire _w20615_ ;
	wire _w20616_ ;
	wire _w20617_ ;
	wire _w20618_ ;
	wire _w20619_ ;
	wire _w20620_ ;
	wire _w20621_ ;
	wire _w20622_ ;
	wire _w20623_ ;
	wire _w20624_ ;
	wire _w20625_ ;
	wire _w20626_ ;
	wire _w20627_ ;
	wire _w20628_ ;
	wire _w20629_ ;
	wire _w20630_ ;
	wire _w20631_ ;
	wire _w20632_ ;
	wire _w20633_ ;
	wire _w20634_ ;
	wire _w20635_ ;
	wire _w20636_ ;
	wire _w20637_ ;
	wire _w20638_ ;
	wire _w20639_ ;
	wire _w20640_ ;
	wire _w20641_ ;
	wire _w20642_ ;
	wire _w20643_ ;
	wire _w20644_ ;
	wire _w20645_ ;
	wire _w20646_ ;
	wire _w20647_ ;
	wire _w20648_ ;
	wire _w20649_ ;
	wire _w20650_ ;
	wire _w20651_ ;
	wire _w20652_ ;
	wire _w20653_ ;
	wire _w20654_ ;
	wire _w20655_ ;
	wire _w20656_ ;
	wire _w20657_ ;
	wire _w20658_ ;
	wire _w20659_ ;
	wire _w20660_ ;
	wire _w20661_ ;
	wire _w20662_ ;
	wire _w20663_ ;
	wire _w20664_ ;
	wire _w20665_ ;
	wire _w20666_ ;
	wire _w20667_ ;
	wire _w20668_ ;
	wire _w20669_ ;
	wire _w20670_ ;
	wire _w20671_ ;
	wire _w20672_ ;
	wire _w20673_ ;
	wire _w20674_ ;
	wire _w20675_ ;
	wire _w20676_ ;
	wire _w20677_ ;
	wire _w20678_ ;
	wire _w20679_ ;
	wire _w20680_ ;
	wire _w20681_ ;
	wire _w20682_ ;
	wire _w20683_ ;
	wire _w20684_ ;
	wire _w20685_ ;
	wire _w20686_ ;
	wire _w20687_ ;
	wire _w20688_ ;
	wire _w20689_ ;
	wire _w20690_ ;
	wire _w20691_ ;
	wire _w20692_ ;
	wire _w20693_ ;
	wire _w20694_ ;
	wire _w20695_ ;
	wire _w20696_ ;
	wire _w20697_ ;
	wire _w20698_ ;
	wire _w20699_ ;
	wire _w20700_ ;
	wire _w20701_ ;
	wire _w20702_ ;
	wire _w20703_ ;
	wire _w20704_ ;
	wire _w20705_ ;
	wire _w20706_ ;
	wire _w20707_ ;
	wire _w20708_ ;
	wire _w20709_ ;
	wire _w20710_ ;
	wire _w20711_ ;
	wire _w20712_ ;
	wire _w20713_ ;
	wire _w20714_ ;
	wire _w20715_ ;
	wire _w20716_ ;
	wire _w20717_ ;
	wire _w20718_ ;
	wire _w20719_ ;
	wire _w20720_ ;
	wire _w20721_ ;
	wire _w20722_ ;
	wire _w20723_ ;
	wire _w20724_ ;
	wire _w20725_ ;
	wire _w20726_ ;
	wire _w20727_ ;
	wire _w20728_ ;
	wire _w20729_ ;
	wire _w20730_ ;
	wire _w20731_ ;
	wire _w20732_ ;
	wire _w20733_ ;
	wire _w20734_ ;
	wire _w20735_ ;
	wire _w20736_ ;
	wire _w20737_ ;
	wire _w20738_ ;
	wire _w20739_ ;
	wire _w20740_ ;
	wire _w20741_ ;
	wire _w20742_ ;
	wire _w20743_ ;
	wire _w20744_ ;
	wire _w20745_ ;
	wire _w20746_ ;
	wire _w20747_ ;
	wire _w20748_ ;
	wire _w20749_ ;
	wire _w20750_ ;
	wire _w20751_ ;
	wire _w20752_ ;
	wire _w20753_ ;
	wire _w20754_ ;
	wire _w20755_ ;
	wire _w20756_ ;
	wire _w20757_ ;
	wire _w20758_ ;
	wire _w20759_ ;
	wire _w20760_ ;
	wire _w20761_ ;
	wire _w20762_ ;
	wire _w20763_ ;
	wire _w20764_ ;
	wire _w20765_ ;
	wire _w20766_ ;
	wire _w20767_ ;
	wire _w20768_ ;
	wire _w20769_ ;
	wire _w20770_ ;
	wire _w20771_ ;
	wire _w20772_ ;
	wire _w20773_ ;
	wire _w20774_ ;
	wire _w20775_ ;
	wire _w20776_ ;
	wire _w20777_ ;
	wire _w20778_ ;
	wire _w20779_ ;
	wire _w20780_ ;
	wire _w20781_ ;
	wire _w20782_ ;
	wire _w20783_ ;
	wire _w20784_ ;
	wire _w20785_ ;
	wire _w20786_ ;
	wire _w20787_ ;
	wire _w20788_ ;
	wire _w20789_ ;
	wire _w20790_ ;
	wire _w20791_ ;
	wire _w20792_ ;
	wire _w20793_ ;
	wire _w20794_ ;
	wire _w20795_ ;
	wire _w20796_ ;
	wire _w20797_ ;
	wire _w20798_ ;
	wire _w20799_ ;
	wire _w20800_ ;
	wire _w20801_ ;
	wire _w20802_ ;
	wire _w20803_ ;
	wire _w20804_ ;
	wire _w20805_ ;
	wire _w20806_ ;
	wire _w20807_ ;
	wire _w20808_ ;
	wire _w20809_ ;
	wire _w20810_ ;
	wire _w20811_ ;
	wire _w20812_ ;
	wire _w20813_ ;
	wire _w20814_ ;
	wire _w20815_ ;
	wire _w20816_ ;
	wire _w20817_ ;
	wire _w20818_ ;
	wire _w20819_ ;
	wire _w20820_ ;
	wire _w20821_ ;
	wire _w20822_ ;
	wire _w20823_ ;
	wire _w20824_ ;
	wire _w20825_ ;
	wire _w20826_ ;
	wire _w20827_ ;
	wire _w20828_ ;
	wire _w20829_ ;
	wire _w20830_ ;
	wire _w20831_ ;
	wire _w20832_ ;
	wire _w20833_ ;
	wire _w20834_ ;
	wire _w20835_ ;
	wire _w20836_ ;
	wire _w20837_ ;
	wire _w20838_ ;
	wire _w20839_ ;
	wire _w20840_ ;
	wire _w20841_ ;
	wire _w20842_ ;
	wire _w20843_ ;
	wire _w20844_ ;
	wire _w20845_ ;
	wire _w20846_ ;
	wire _w20847_ ;
	wire _w20848_ ;
	wire _w20849_ ;
	wire _w20850_ ;
	wire _w20851_ ;
	wire _w20852_ ;
	wire _w20853_ ;
	wire _w20854_ ;
	wire _w20855_ ;
	wire _w20856_ ;
	wire _w20857_ ;
	wire _w20858_ ;
	wire _w20859_ ;
	wire _w20860_ ;
	wire _w20861_ ;
	wire _w20862_ ;
	wire _w20863_ ;
	wire _w20864_ ;
	wire _w20865_ ;
	wire _w20866_ ;
	wire _w20867_ ;
	wire _w20868_ ;
	wire _w20869_ ;
	wire _w20870_ ;
	wire _w20871_ ;
	wire _w20872_ ;
	wire _w20873_ ;
	wire _w20874_ ;
	wire _w20875_ ;
	wire _w20876_ ;
	wire _w20877_ ;
	wire _w20878_ ;
	wire _w20879_ ;
	wire _w20880_ ;
	wire _w20881_ ;
	wire _w20882_ ;
	wire _w20883_ ;
	wire _w20884_ ;
	wire _w20885_ ;
	wire _w20886_ ;
	wire _w20887_ ;
	wire _w20888_ ;
	wire _w20889_ ;
	wire _w20890_ ;
	wire _w20891_ ;
	wire _w20892_ ;
	wire _w20893_ ;
	wire _w20894_ ;
	wire _w20895_ ;
	wire _w20896_ ;
	wire _w20897_ ;
	wire _w20898_ ;
	wire _w20899_ ;
	wire _w20900_ ;
	wire _w20901_ ;
	wire _w20902_ ;
	wire _w20903_ ;
	wire _w20904_ ;
	wire _w20905_ ;
	wire _w20906_ ;
	wire _w20907_ ;
	wire _w20908_ ;
	wire _w20909_ ;
	wire _w20910_ ;
	wire _w20911_ ;
	wire _w20912_ ;
	wire _w20913_ ;
	wire _w20914_ ;
	wire _w20915_ ;
	wire _w20916_ ;
	wire _w20917_ ;
	wire _w20918_ ;
	wire _w20919_ ;
	wire _w20920_ ;
	wire _w20921_ ;
	wire _w20922_ ;
	wire _w20923_ ;
	wire _w20924_ ;
	wire _w20925_ ;
	wire _w20926_ ;
	wire _w20927_ ;
	wire _w20928_ ;
	wire _w20929_ ;
	wire _w20930_ ;
	wire _w20931_ ;
	wire _w20932_ ;
	wire _w20933_ ;
	wire _w20934_ ;
	wire _w20935_ ;
	wire _w20936_ ;
	wire _w20937_ ;
	wire _w20938_ ;
	wire _w20939_ ;
	wire _w20940_ ;
	wire _w20941_ ;
	wire _w20942_ ;
	wire _w20943_ ;
	wire _w20944_ ;
	wire _w20945_ ;
	wire _w20946_ ;
	wire _w20947_ ;
	wire _w20948_ ;
	wire _w20949_ ;
	wire _w20950_ ;
	wire _w20951_ ;
	wire _w20952_ ;
	wire _w20953_ ;
	wire _w20954_ ;
	wire _w20955_ ;
	wire _w20956_ ;
	wire _w20957_ ;
	wire _w20958_ ;
	wire _w20959_ ;
	wire _w20960_ ;
	wire _w20961_ ;
	wire _w20962_ ;
	wire _w20963_ ;
	wire _w20964_ ;
	wire _w20965_ ;
	wire _w20966_ ;
	wire _w20967_ ;
	wire _w20968_ ;
	wire _w20969_ ;
	wire _w20970_ ;
	wire _w20971_ ;
	wire _w20972_ ;
	wire _w20973_ ;
	wire _w20974_ ;
	wire _w20975_ ;
	wire _w20976_ ;
	wire _w20977_ ;
	wire _w20978_ ;
	wire _w20979_ ;
	wire _w20980_ ;
	wire _w20981_ ;
	wire _w20982_ ;
	wire _w20983_ ;
	wire _w20984_ ;
	wire _w20985_ ;
	wire _w20986_ ;
	wire _w20987_ ;
	wire _w20988_ ;
	wire _w20989_ ;
	wire _w20990_ ;
	wire _w20991_ ;
	wire _w20992_ ;
	wire _w20993_ ;
	wire _w20994_ ;
	wire _w20995_ ;
	wire _w20996_ ;
	wire _w20997_ ;
	wire _w20998_ ;
	wire _w20999_ ;
	wire _w21000_ ;
	wire _w21001_ ;
	wire _w21002_ ;
	wire _w21003_ ;
	wire _w21004_ ;
	wire _w21005_ ;
	wire _w21006_ ;
	wire _w21007_ ;
	wire _w21008_ ;
	wire _w21009_ ;
	wire _w21010_ ;
	wire _w21011_ ;
	wire _w21012_ ;
	wire _w21013_ ;
	wire _w21014_ ;
	wire _w21015_ ;
	wire _w21016_ ;
	wire _w21017_ ;
	wire _w21018_ ;
	wire _w21019_ ;
	wire _w21020_ ;
	wire _w21021_ ;
	wire _w21022_ ;
	wire _w21023_ ;
	wire _w21024_ ;
	wire _w21025_ ;
	wire _w21026_ ;
	wire _w21027_ ;
	wire _w21028_ ;
	wire _w21029_ ;
	wire _w21030_ ;
	wire _w21031_ ;
	wire _w21032_ ;
	wire _w21033_ ;
	wire _w21034_ ;
	wire _w21035_ ;
	wire _w21036_ ;
	wire _w21037_ ;
	wire _w21038_ ;
	wire _w21039_ ;
	wire _w21040_ ;
	wire _w21041_ ;
	wire _w21042_ ;
	wire _w21043_ ;
	wire _w21044_ ;
	wire _w21045_ ;
	wire _w21046_ ;
	wire _w21047_ ;
	wire _w21048_ ;
	wire _w21049_ ;
	wire _w21050_ ;
	wire _w21051_ ;
	wire _w21052_ ;
	wire _w21053_ ;
	wire _w21054_ ;
	wire _w21055_ ;
	wire _w21056_ ;
	wire _w21057_ ;
	wire _w21058_ ;
	wire _w21059_ ;
	wire _w21060_ ;
	wire _w21061_ ;
	wire _w21062_ ;
	wire _w21063_ ;
	wire _w21064_ ;
	wire _w21065_ ;
	wire _w21066_ ;
	wire _w21067_ ;
	wire _w21068_ ;
	wire _w21069_ ;
	wire _w21070_ ;
	wire _w21071_ ;
	wire _w21072_ ;
	wire _w21073_ ;
	wire _w21074_ ;
	wire _w21075_ ;
	wire _w21076_ ;
	wire _w21077_ ;
	wire _w21078_ ;
	wire _w21079_ ;
	wire _w21080_ ;
	wire _w21081_ ;
	wire _w21082_ ;
	wire _w21083_ ;
	wire _w21084_ ;
	wire _w21085_ ;
	wire _w21086_ ;
	wire _w21087_ ;
	wire _w21088_ ;
	wire _w21089_ ;
	wire _w21090_ ;
	wire _w21091_ ;
	wire _w21092_ ;
	wire _w21093_ ;
	wire _w21094_ ;
	wire _w21095_ ;
	wire _w21096_ ;
	wire _w21097_ ;
	wire _w21098_ ;
	wire _w21099_ ;
	wire _w21100_ ;
	wire _w21101_ ;
	wire _w21102_ ;
	wire _w21103_ ;
	wire _w21104_ ;
	wire _w21105_ ;
	wire _w21106_ ;
	wire _w21107_ ;
	wire _w21108_ ;
	wire _w21109_ ;
	wire _w21110_ ;
	wire _w21111_ ;
	wire _w21112_ ;
	wire _w21113_ ;
	wire _w21114_ ;
	wire _w21115_ ;
	wire _w21116_ ;
	wire _w21117_ ;
	wire _w21118_ ;
	wire _w21119_ ;
	wire _w21120_ ;
	wire _w21121_ ;
	wire _w21122_ ;
	wire _w21123_ ;
	wire _w21124_ ;
	wire _w21125_ ;
	wire _w21126_ ;
	wire _w21127_ ;
	wire _w21128_ ;
	wire _w21129_ ;
	wire _w21130_ ;
	wire _w21131_ ;
	wire _w21132_ ;
	wire _w21133_ ;
	wire _w21134_ ;
	wire _w21135_ ;
	wire _w21136_ ;
	wire _w21137_ ;
	wire _w21138_ ;
	wire _w21139_ ;
	wire _w21140_ ;
	wire _w21141_ ;
	wire _w21142_ ;
	wire _w21143_ ;
	wire _w21144_ ;
	wire _w21145_ ;
	wire _w21146_ ;
	wire _w21147_ ;
	wire _w21148_ ;
	wire _w21149_ ;
	wire _w21150_ ;
	wire _w21151_ ;
	wire _w21152_ ;
	wire _w21153_ ;
	wire _w21154_ ;
	wire _w21155_ ;
	wire _w21156_ ;
	wire _w21157_ ;
	wire _w21158_ ;
	wire _w21159_ ;
	wire _w21160_ ;
	wire _w21161_ ;
	wire _w21162_ ;
	wire _w21163_ ;
	wire _w21164_ ;
	wire _w21165_ ;
	wire _w21166_ ;
	wire _w21167_ ;
	wire _w21168_ ;
	wire _w21169_ ;
	wire _w21170_ ;
	wire _w21171_ ;
	wire _w21172_ ;
	wire _w21173_ ;
	wire _w21174_ ;
	wire _w21175_ ;
	wire _w21176_ ;
	wire _w21177_ ;
	wire _w21178_ ;
	wire _w21179_ ;
	wire _w21180_ ;
	wire _w21181_ ;
	wire _w21182_ ;
	wire _w21183_ ;
	wire _w21184_ ;
	wire _w21185_ ;
	wire _w21186_ ;
	wire _w21187_ ;
	wire _w21188_ ;
	wire _w21189_ ;
	wire _w21190_ ;
	wire _w21191_ ;
	wire _w21192_ ;
	wire _w21193_ ;
	wire _w21194_ ;
	wire _w21195_ ;
	wire _w21196_ ;
	wire _w21197_ ;
	wire _w21198_ ;
	wire _w21199_ ;
	wire _w21200_ ;
	wire _w21201_ ;
	wire _w21202_ ;
	wire _w21203_ ;
	wire _w21204_ ;
	wire _w21205_ ;
	wire _w21206_ ;
	wire _w21207_ ;
	wire _w21208_ ;
	wire _w21209_ ;
	wire _w21210_ ;
	wire _w21211_ ;
	wire _w21212_ ;
	wire _w21213_ ;
	wire _w21214_ ;
	wire _w21215_ ;
	wire _w21216_ ;
	wire _w21217_ ;
	wire _w21218_ ;
	wire _w21219_ ;
	wire _w21220_ ;
	wire _w21221_ ;
	wire _w21222_ ;
	wire _w21223_ ;
	wire _w21224_ ;
	wire _w21225_ ;
	wire _w21226_ ;
	wire _w21227_ ;
	wire _w21228_ ;
	wire _w21229_ ;
	wire _w21230_ ;
	wire _w21231_ ;
	wire _w21232_ ;
	wire _w21233_ ;
	wire _w21234_ ;
	wire _w21235_ ;
	wire _w21236_ ;
	wire _w21237_ ;
	wire _w21238_ ;
	wire _w21239_ ;
	wire _w21240_ ;
	wire _w21241_ ;
	wire _w21242_ ;
	wire _w21243_ ;
	wire _w21244_ ;
	wire _w21245_ ;
	wire _w21246_ ;
	wire _w21247_ ;
	wire _w21248_ ;
	wire _w21249_ ;
	wire _w21250_ ;
	wire _w21251_ ;
	wire _w21252_ ;
	wire _w21253_ ;
	wire _w21254_ ;
	wire _w21255_ ;
	wire _w21256_ ;
	wire _w21257_ ;
	wire _w21258_ ;
	wire _w21259_ ;
	wire _w21260_ ;
	wire _w21261_ ;
	wire _w21262_ ;
	wire _w21263_ ;
	wire _w21264_ ;
	wire _w21265_ ;
	wire _w21266_ ;
	wire _w21267_ ;
	wire _w21268_ ;
	wire _w21269_ ;
	wire _w21270_ ;
	wire _w21271_ ;
	wire _w21272_ ;
	wire _w21273_ ;
	wire _w21274_ ;
	wire _w21275_ ;
	wire _w21276_ ;
	wire _w21277_ ;
	wire _w21278_ ;
	wire _w21279_ ;
	wire _w21280_ ;
	wire _w21281_ ;
	wire _w21282_ ;
	wire _w21283_ ;
	wire _w21284_ ;
	wire _w21285_ ;
	wire _w21286_ ;
	wire _w21287_ ;
	wire _w21288_ ;
	wire _w21289_ ;
	wire _w21290_ ;
	wire _w21291_ ;
	wire _w21292_ ;
	wire _w21293_ ;
	wire _w21294_ ;
	wire _w21295_ ;
	wire _w21296_ ;
	wire _w21297_ ;
	wire _w21298_ ;
	wire _w21299_ ;
	wire _w21300_ ;
	wire _w21301_ ;
	wire _w21302_ ;
	wire _w21303_ ;
	wire _w21304_ ;
	wire _w21305_ ;
	wire _w21306_ ;
	wire _w21307_ ;
	wire _w21308_ ;
	wire _w21309_ ;
	wire _w21310_ ;
	wire _w21311_ ;
	wire _w21312_ ;
	wire _w21313_ ;
	wire _w21314_ ;
	wire _w21315_ ;
	wire _w21316_ ;
	wire _w21317_ ;
	wire _w21318_ ;
	wire _w21319_ ;
	wire _w21320_ ;
	wire _w21321_ ;
	wire _w21322_ ;
	wire _w21323_ ;
	wire _w21324_ ;
	wire _w21325_ ;
	wire _w21326_ ;
	wire _w21327_ ;
	wire _w21328_ ;
	wire _w21329_ ;
	wire _w21330_ ;
	wire _w21331_ ;
	wire _w21332_ ;
	wire _w21333_ ;
	wire _w21334_ ;
	wire _w21335_ ;
	wire _w21336_ ;
	wire _w21337_ ;
	wire _w21338_ ;
	wire _w21339_ ;
	wire _w21340_ ;
	wire _w21341_ ;
	wire _w21342_ ;
	wire _w21343_ ;
	wire _w21344_ ;
	wire _w21345_ ;
	wire _w21346_ ;
	wire _w21347_ ;
	wire _w21348_ ;
	wire _w21349_ ;
	wire _w21350_ ;
	wire _w21351_ ;
	wire _w21352_ ;
	wire _w21353_ ;
	wire _w21354_ ;
	wire _w21355_ ;
	wire _w21356_ ;
	wire _w21357_ ;
	wire _w21358_ ;
	wire _w21359_ ;
	wire _w21360_ ;
	wire _w21361_ ;
	wire _w21362_ ;
	wire _w21363_ ;
	wire _w21364_ ;
	wire _w21365_ ;
	wire _w21366_ ;
	wire _w21367_ ;
	wire _w21368_ ;
	wire _w21369_ ;
	wire _w21370_ ;
	wire _w21371_ ;
	wire _w21372_ ;
	wire _w21373_ ;
	wire _w21374_ ;
	wire _w21375_ ;
	wire _w21376_ ;
	wire _w21377_ ;
	wire _w21378_ ;
	wire _w21379_ ;
	wire _w21380_ ;
	wire _w21381_ ;
	wire _w21382_ ;
	wire _w21383_ ;
	wire _w21384_ ;
	wire _w21385_ ;
	wire _w21386_ ;
	wire _w21387_ ;
	wire _w21388_ ;
	wire _w21389_ ;
	wire _w21390_ ;
	wire _w21391_ ;
	wire _w21392_ ;
	wire _w21393_ ;
	wire _w21394_ ;
	wire _w21395_ ;
	wire _w21396_ ;
	wire _w21397_ ;
	wire _w21398_ ;
	wire _w21399_ ;
	wire _w21400_ ;
	wire _w21401_ ;
	wire _w21402_ ;
	wire _w21403_ ;
	wire _w21404_ ;
	wire _w21405_ ;
	wire _w21406_ ;
	wire _w21407_ ;
	wire _w21408_ ;
	wire _w21409_ ;
	wire _w21410_ ;
	wire _w21411_ ;
	wire _w21412_ ;
	wire _w21413_ ;
	wire _w21414_ ;
	wire _w21415_ ;
	wire _w21416_ ;
	wire _w21417_ ;
	wire _w21418_ ;
	wire _w21419_ ;
	wire _w21420_ ;
	wire _w21421_ ;
	wire _w21422_ ;
	wire _w21423_ ;
	wire _w21424_ ;
	wire _w21425_ ;
	wire _w21426_ ;
	wire _w21427_ ;
	wire _w21428_ ;
	wire _w21429_ ;
	wire _w21430_ ;
	wire _w21431_ ;
	wire _w21432_ ;
	wire _w21433_ ;
	wire _w21434_ ;
	wire _w21435_ ;
	wire _w21436_ ;
	wire _w21437_ ;
	wire _w21438_ ;
	wire _w21439_ ;
	wire _w21440_ ;
	wire _w21441_ ;
	wire _w21442_ ;
	wire _w21443_ ;
	wire _w21444_ ;
	wire _w21445_ ;
	wire _w21446_ ;
	wire _w21447_ ;
	wire _w21448_ ;
	wire _w21449_ ;
	wire _w21450_ ;
	wire _w21451_ ;
	wire _w21452_ ;
	wire _w21453_ ;
	wire _w21454_ ;
	wire _w21455_ ;
	wire _w21456_ ;
	wire _w21457_ ;
	wire _w21458_ ;
	wire _w21459_ ;
	wire _w21460_ ;
	wire _w21461_ ;
	wire _w21462_ ;
	wire _w21463_ ;
	wire _w21464_ ;
	wire _w21465_ ;
	wire _w21466_ ;
	wire _w21467_ ;
	wire _w21468_ ;
	wire _w21469_ ;
	wire _w21470_ ;
	wire _w21471_ ;
	wire _w21472_ ;
	wire _w21473_ ;
	wire _w21474_ ;
	wire _w21475_ ;
	wire _w21476_ ;
	wire _w21477_ ;
	wire _w21478_ ;
	wire _w21479_ ;
	wire _w21480_ ;
	wire _w21481_ ;
	wire _w21482_ ;
	wire _w21483_ ;
	wire _w21484_ ;
	wire _w21485_ ;
	wire _w21486_ ;
	wire _w21487_ ;
	wire _w21488_ ;
	wire _w21489_ ;
	wire _w21490_ ;
	wire _w21491_ ;
	wire _w21492_ ;
	wire _w21493_ ;
	wire _w21494_ ;
	wire _w21495_ ;
	wire _w21496_ ;
	wire _w21497_ ;
	wire _w21498_ ;
	wire _w21499_ ;
	wire _w21500_ ;
	wire _w21501_ ;
	wire _w21502_ ;
	wire _w21503_ ;
	wire _w21504_ ;
	wire _w21505_ ;
	wire _w21506_ ;
	wire _w21507_ ;
	wire _w21508_ ;
	wire _w21509_ ;
	wire _w21510_ ;
	wire _w21511_ ;
	wire _w21512_ ;
	wire _w21513_ ;
	wire _w21514_ ;
	wire _w21515_ ;
	wire _w21516_ ;
	wire _w21517_ ;
	wire _w21518_ ;
	wire _w21519_ ;
	wire _w21520_ ;
	wire _w21521_ ;
	wire _w21522_ ;
	wire _w21523_ ;
	wire _w21524_ ;
	wire _w21525_ ;
	wire _w21526_ ;
	wire _w21527_ ;
	wire _w21528_ ;
	wire _w21529_ ;
	wire _w21530_ ;
	wire _w21531_ ;
	wire _w21532_ ;
	wire _w21533_ ;
	wire _w21534_ ;
	wire _w21535_ ;
	wire _w21536_ ;
	wire _w21537_ ;
	wire _w21538_ ;
	wire _w21539_ ;
	wire _w21540_ ;
	wire _w21541_ ;
	wire _w21542_ ;
	wire _w21543_ ;
	wire _w21544_ ;
	wire _w21545_ ;
	wire _w21546_ ;
	wire _w21547_ ;
	wire _w21548_ ;
	wire _w21549_ ;
	wire _w21550_ ;
	wire _w21551_ ;
	wire _w21552_ ;
	wire _w21553_ ;
	wire _w21554_ ;
	wire _w21555_ ;
	wire _w21556_ ;
	wire _w21557_ ;
	wire _w21558_ ;
	wire _w21559_ ;
	wire _w21560_ ;
	wire _w21561_ ;
	wire _w21562_ ;
	wire _w21563_ ;
	wire _w21564_ ;
	wire _w21565_ ;
	wire _w21566_ ;
	wire _w21567_ ;
	wire _w21568_ ;
	wire _w21569_ ;
	wire _w21570_ ;
	wire _w21571_ ;
	wire _w21572_ ;
	wire _w21573_ ;
	wire _w21574_ ;
	wire _w21575_ ;
	wire _w21576_ ;
	wire _w21577_ ;
	wire _w21578_ ;
	wire _w21579_ ;
	wire _w21580_ ;
	wire _w21581_ ;
	wire _w21582_ ;
	wire _w21583_ ;
	wire _w21584_ ;
	wire _w21585_ ;
	wire _w21586_ ;
	wire _w21587_ ;
	wire _w21588_ ;
	wire _w21589_ ;
	wire _w21590_ ;
	wire _w21591_ ;
	wire _w21592_ ;
	wire _w21593_ ;
	wire _w21594_ ;
	wire _w21595_ ;
	wire _w21596_ ;
	wire _w21597_ ;
	wire _w21598_ ;
	wire _w21599_ ;
	wire _w21600_ ;
	wire _w21601_ ;
	wire _w21602_ ;
	wire _w21603_ ;
	wire _w21604_ ;
	wire _w21605_ ;
	wire _w21606_ ;
	wire _w21607_ ;
	wire _w21608_ ;
	wire _w21609_ ;
	wire _w21610_ ;
	wire _w21611_ ;
	wire _w21612_ ;
	wire _w21613_ ;
	wire _w21614_ ;
	wire _w21615_ ;
	wire _w21616_ ;
	wire _w21617_ ;
	wire _w21618_ ;
	wire _w21619_ ;
	wire _w21620_ ;
	wire _w21621_ ;
	wire _w21622_ ;
	wire _w21623_ ;
	wire _w21624_ ;
	wire _w21625_ ;
	wire _w21626_ ;
	wire _w21627_ ;
	wire _w21628_ ;
	wire _w21629_ ;
	wire _w21630_ ;
	wire _w21631_ ;
	wire _w21632_ ;
	wire _w21633_ ;
	wire _w21634_ ;
	wire _w21635_ ;
	wire _w21636_ ;
	wire _w21637_ ;
	wire _w21638_ ;
	wire _w21639_ ;
	wire _w21640_ ;
	wire _w21641_ ;
	wire _w21642_ ;
	wire _w21643_ ;
	wire _w21644_ ;
	wire _w21645_ ;
	wire _w21646_ ;
	wire _w21647_ ;
	wire _w21648_ ;
	wire _w21649_ ;
	wire _w21650_ ;
	wire _w21651_ ;
	wire _w21652_ ;
	wire _w21653_ ;
	wire _w21654_ ;
	wire _w21655_ ;
	wire _w21656_ ;
	wire _w21657_ ;
	wire _w21658_ ;
	wire _w21659_ ;
	wire _w21660_ ;
	wire _w21661_ ;
	wire _w21662_ ;
	wire _w21663_ ;
	wire _w21664_ ;
	wire _w21665_ ;
	wire _w21666_ ;
	wire _w21667_ ;
	wire _w21668_ ;
	wire _w21669_ ;
	wire _w21670_ ;
	wire _w21671_ ;
	wire _w21672_ ;
	wire _w21673_ ;
	wire _w21674_ ;
	wire _w21675_ ;
	wire _w21676_ ;
	wire _w21677_ ;
	wire _w21678_ ;
	wire _w21679_ ;
	wire _w21680_ ;
	wire _w21681_ ;
	wire _w21682_ ;
	wire _w21683_ ;
	wire _w21684_ ;
	wire _w21685_ ;
	wire _w21686_ ;
	wire _w21687_ ;
	wire _w21688_ ;
	wire _w21689_ ;
	wire _w21690_ ;
	wire _w21691_ ;
	wire _w21692_ ;
	wire _w21693_ ;
	wire _w21694_ ;
	wire _w21695_ ;
	wire _w21696_ ;
	wire _w21697_ ;
	wire _w21698_ ;
	wire _w21699_ ;
	wire _w21700_ ;
	wire _w21701_ ;
	wire _w21702_ ;
	wire _w21703_ ;
	wire _w21704_ ;
	wire _w21705_ ;
	wire _w21706_ ;
	wire _w21707_ ;
	wire _w21708_ ;
	wire _w21709_ ;
	wire _w21710_ ;
	wire _w21711_ ;
	wire _w21712_ ;
	wire _w21713_ ;
	wire _w21714_ ;
	wire _w21715_ ;
	wire _w21716_ ;
	wire _w21717_ ;
	wire _w21718_ ;
	wire _w21719_ ;
	wire _w21720_ ;
	wire _w21721_ ;
	wire _w21722_ ;
	wire _w21723_ ;
	wire _w21724_ ;
	wire _w21725_ ;
	wire _w21726_ ;
	wire _w21727_ ;
	wire _w21728_ ;
	wire _w21729_ ;
	wire _w21730_ ;
	wire _w21731_ ;
	wire _w21732_ ;
	wire _w21733_ ;
	wire _w21734_ ;
	wire _w21735_ ;
	wire _w21736_ ;
	wire _w21737_ ;
	wire _w21738_ ;
	wire _w21739_ ;
	wire _w21740_ ;
	wire _w21741_ ;
	wire _w21742_ ;
	wire _w21743_ ;
	wire _w21744_ ;
	wire _w21745_ ;
	wire _w21746_ ;
	wire _w21747_ ;
	wire _w21748_ ;
	wire _w21749_ ;
	wire _w21750_ ;
	wire _w21751_ ;
	wire _w21752_ ;
	wire _w21753_ ;
	wire _w21754_ ;
	wire _w21755_ ;
	wire _w21756_ ;
	wire _w21757_ ;
	wire _w21758_ ;
	wire _w21759_ ;
	wire _w21760_ ;
	wire _w21761_ ;
	wire _w21762_ ;
	wire _w21763_ ;
	wire _w21764_ ;
	wire _w21765_ ;
	wire _w21766_ ;
	wire _w21767_ ;
	wire _w21768_ ;
	wire _w21769_ ;
	wire _w21770_ ;
	wire _w21771_ ;
	wire _w21772_ ;
	wire _w21773_ ;
	wire _w21774_ ;
	wire _w21775_ ;
	wire _w21776_ ;
	wire _w21777_ ;
	wire _w21778_ ;
	wire _w21779_ ;
	wire _w21780_ ;
	wire _w21781_ ;
	wire _w21782_ ;
	wire _w21783_ ;
	wire _w21784_ ;
	wire _w21785_ ;
	wire _w21786_ ;
	wire _w21787_ ;
	wire _w21788_ ;
	wire _w21789_ ;
	wire _w21790_ ;
	wire _w21791_ ;
	wire _w21792_ ;
	wire _w21793_ ;
	wire _w21794_ ;
	wire _w21795_ ;
	wire _w21796_ ;
	wire _w21797_ ;
	wire _w21798_ ;
	wire _w21799_ ;
	wire _w21800_ ;
	wire _w21801_ ;
	wire _w21802_ ;
	wire _w21803_ ;
	wire _w21804_ ;
	wire _w21805_ ;
	wire _w21806_ ;
	wire _w21807_ ;
	wire _w21808_ ;
	wire _w21809_ ;
	wire _w21810_ ;
	wire _w21811_ ;
	wire _w21812_ ;
	wire _w21813_ ;
	wire _w21814_ ;
	wire _w21815_ ;
	wire _w21816_ ;
	wire _w21817_ ;
	wire _w21818_ ;
	wire _w21819_ ;
	wire _w21820_ ;
	wire _w21821_ ;
	wire _w21822_ ;
	wire _w21823_ ;
	wire _w21824_ ;
	wire _w21825_ ;
	wire _w21826_ ;
	wire _w21827_ ;
	wire _w21828_ ;
	wire _w21829_ ;
	wire _w21830_ ;
	wire _w21831_ ;
	wire _w21832_ ;
	wire _w21833_ ;
	wire _w21834_ ;
	wire _w21835_ ;
	wire _w21836_ ;
	wire _w21837_ ;
	wire _w21838_ ;
	wire _w21839_ ;
	wire _w21840_ ;
	wire _w21841_ ;
	wire _w21842_ ;
	wire _w21843_ ;
	wire _w21844_ ;
	wire _w21845_ ;
	wire _w21846_ ;
	wire _w21847_ ;
	wire _w21848_ ;
	wire _w21849_ ;
	wire _w21850_ ;
	wire _w21851_ ;
	wire _w21852_ ;
	wire _w21853_ ;
	wire _w21854_ ;
	wire _w21855_ ;
	wire _w21856_ ;
	wire _w21857_ ;
	wire _w21858_ ;
	wire _w21859_ ;
	wire _w21860_ ;
	wire _w21861_ ;
	wire _w21862_ ;
	wire _w21863_ ;
	wire _w21864_ ;
	wire _w21865_ ;
	wire _w21866_ ;
	wire _w21867_ ;
	wire _w21868_ ;
	wire _w21869_ ;
	wire _w21870_ ;
	wire _w21871_ ;
	wire _w21872_ ;
	wire _w21873_ ;
	wire _w21874_ ;
	wire _w21875_ ;
	wire _w21876_ ;
	wire _w21877_ ;
	wire _w21878_ ;
	wire _w21879_ ;
	wire _w21880_ ;
	wire _w21881_ ;
	wire _w21882_ ;
	wire _w21883_ ;
	wire _w21884_ ;
	wire _w21885_ ;
	wire _w21886_ ;
	wire _w21887_ ;
	wire _w21888_ ;
	wire _w21889_ ;
	wire _w21890_ ;
	wire _w21891_ ;
	wire _w21892_ ;
	wire _w21893_ ;
	wire _w21894_ ;
	wire _w21895_ ;
	wire _w21896_ ;
	wire _w21897_ ;
	wire _w21898_ ;
	wire _w21899_ ;
	wire _w21900_ ;
	wire _w21901_ ;
	wire _w21902_ ;
	wire _w21903_ ;
	wire _w21904_ ;
	wire _w21905_ ;
	wire _w21906_ ;
	wire _w21907_ ;
	wire _w21908_ ;
	wire _w21909_ ;
	wire _w21910_ ;
	wire _w21911_ ;
	wire _w21912_ ;
	wire _w21913_ ;
	wire _w21914_ ;
	wire _w21915_ ;
	wire _w21916_ ;
	wire _w21917_ ;
	wire _w21918_ ;
	wire _w21919_ ;
	wire _w21920_ ;
	wire _w21921_ ;
	wire _w21922_ ;
	wire _w21923_ ;
	wire _w21924_ ;
	wire _w21925_ ;
	wire _w21926_ ;
	wire _w21927_ ;
	wire _w21928_ ;
	wire _w21929_ ;
	wire _w21930_ ;
	wire _w21931_ ;
	wire _w21932_ ;
	wire _w21933_ ;
	wire _w21934_ ;
	wire _w21935_ ;
	wire _w21936_ ;
	wire _w21937_ ;
	wire _w21938_ ;
	wire _w21939_ ;
	wire _w21940_ ;
	wire _w21941_ ;
	wire _w21942_ ;
	wire _w21943_ ;
	wire _w21944_ ;
	wire _w21945_ ;
	wire _w21946_ ;
	wire _w21947_ ;
	wire _w21948_ ;
	wire _w21949_ ;
	wire _w21950_ ;
	wire _w21951_ ;
	wire _w21952_ ;
	wire _w21953_ ;
	wire _w21954_ ;
	wire _w21955_ ;
	wire _w21956_ ;
	wire _w21957_ ;
	wire _w21958_ ;
	wire _w21959_ ;
	wire _w21960_ ;
	wire _w21961_ ;
	wire _w21962_ ;
	wire _w21963_ ;
	wire _w21964_ ;
	wire _w21965_ ;
	wire _w21966_ ;
	wire _w21967_ ;
	wire _w21968_ ;
	wire _w21969_ ;
	wire _w21970_ ;
	wire _w21971_ ;
	wire _w21972_ ;
	wire _w21973_ ;
	wire _w21974_ ;
	wire _w21975_ ;
	wire _w21976_ ;
	wire _w21977_ ;
	wire _w21978_ ;
	wire _w21979_ ;
	wire _w21980_ ;
	wire _w21981_ ;
	wire _w21982_ ;
	wire _w21983_ ;
	wire _w21984_ ;
	wire _w21985_ ;
	wire _w21986_ ;
	wire _w21987_ ;
	wire _w21988_ ;
	wire _w21989_ ;
	wire _w21990_ ;
	wire _w21991_ ;
	wire _w21992_ ;
	wire _w21993_ ;
	wire _w21994_ ;
	wire _w21995_ ;
	wire _w21996_ ;
	wire _w21997_ ;
	wire _w21998_ ;
	wire _w21999_ ;
	wire _w22000_ ;
	wire _w22001_ ;
	wire _w22002_ ;
	wire _w22003_ ;
	wire _w22004_ ;
	wire _w22005_ ;
	wire _w22006_ ;
	wire _w22007_ ;
	wire _w22008_ ;
	wire _w22009_ ;
	wire _w22010_ ;
	wire _w22011_ ;
	wire _w22012_ ;
	wire _w22013_ ;
	wire _w22014_ ;
	wire _w22015_ ;
	wire _w22016_ ;
	wire _w22017_ ;
	wire _w22018_ ;
	wire _w22019_ ;
	wire _w22020_ ;
	wire _w22021_ ;
	wire _w22022_ ;
	wire _w22023_ ;
	wire _w22024_ ;
	wire _w22025_ ;
	wire _w22026_ ;
	wire _w22027_ ;
	wire _w22028_ ;
	wire _w22029_ ;
	wire _w22030_ ;
	wire _w22031_ ;
	wire _w22032_ ;
	wire _w22033_ ;
	wire _w22034_ ;
	wire _w22035_ ;
	wire _w22036_ ;
	wire _w22037_ ;
	wire _w22038_ ;
	wire _w22039_ ;
	wire _w22040_ ;
	wire _w22041_ ;
	wire _w22042_ ;
	wire _w22043_ ;
	wire _w22044_ ;
	wire _w22045_ ;
	wire _w22046_ ;
	wire _w22047_ ;
	wire _w22048_ ;
	wire _w22049_ ;
	wire _w22050_ ;
	wire _w22051_ ;
	wire _w22052_ ;
	wire _w22053_ ;
	wire _w22054_ ;
	wire _w22055_ ;
	wire _w22056_ ;
	wire _w22057_ ;
	wire _w22058_ ;
	wire _w22059_ ;
	wire _w22060_ ;
	wire _w22061_ ;
	wire _w22062_ ;
	wire _w22063_ ;
	wire _w22064_ ;
	wire _w22065_ ;
	wire _w22066_ ;
	wire _w22067_ ;
	wire _w22068_ ;
	wire _w22069_ ;
	wire _w22070_ ;
	wire _w22071_ ;
	wire _w22072_ ;
	wire _w22073_ ;
	wire _w22074_ ;
	wire _w22075_ ;
	wire _w22076_ ;
	wire _w22077_ ;
	wire _w22078_ ;
	wire _w22079_ ;
	wire _w22080_ ;
	wire _w22081_ ;
	wire _w22082_ ;
	wire _w22083_ ;
	wire _w22084_ ;
	wire _w22085_ ;
	wire _w22086_ ;
	wire _w22087_ ;
	wire _w22088_ ;
	wire _w22089_ ;
	wire _w22090_ ;
	wire _w22091_ ;
	wire _w22092_ ;
	wire _w22093_ ;
	wire _w22094_ ;
	wire _w22095_ ;
	wire _w22096_ ;
	wire _w22097_ ;
	wire _w22098_ ;
	wire _w22099_ ;
	wire _w22100_ ;
	wire _w22101_ ;
	wire _w22102_ ;
	wire _w22103_ ;
	wire _w22104_ ;
	wire _w22105_ ;
	wire _w22106_ ;
	wire _w22107_ ;
	wire _w22108_ ;
	wire _w22109_ ;
	wire _w22110_ ;
	wire _w22111_ ;
	wire _w22112_ ;
	wire _w22113_ ;
	wire _w22114_ ;
	wire _w22115_ ;
	wire _w22116_ ;
	wire _w22117_ ;
	wire _w22118_ ;
	wire _w22119_ ;
	wire _w22120_ ;
	wire _w22121_ ;
	wire _w22122_ ;
	wire _w22123_ ;
	wire _w22124_ ;
	wire _w22125_ ;
	wire _w22126_ ;
	wire _w22127_ ;
	wire _w22128_ ;
	wire _w22129_ ;
	wire _w22130_ ;
	wire _w22131_ ;
	wire _w22132_ ;
	wire _w22133_ ;
	wire _w22134_ ;
	wire _w22135_ ;
	wire _w22136_ ;
	wire _w22137_ ;
	wire _w22138_ ;
	wire _w22139_ ;
	wire _w22140_ ;
	wire _w22141_ ;
	wire _w22142_ ;
	wire _w22143_ ;
	wire _w22144_ ;
	wire _w22145_ ;
	wire _w22146_ ;
	wire _w22147_ ;
	wire _w22148_ ;
	wire _w22149_ ;
	wire _w22150_ ;
	wire _w22151_ ;
	wire _w22152_ ;
	wire _w22153_ ;
	wire _w22154_ ;
	wire _w22155_ ;
	wire _w22156_ ;
	wire _w22157_ ;
	wire _w22158_ ;
	wire _w22159_ ;
	wire _w22160_ ;
	wire _w22161_ ;
	wire _w22162_ ;
	wire _w22163_ ;
	wire _w22164_ ;
	wire _w22165_ ;
	wire _w22166_ ;
	wire _w22167_ ;
	wire _w22168_ ;
	wire _w22169_ ;
	wire _w22170_ ;
	wire _w22171_ ;
	wire _w22172_ ;
	wire _w22173_ ;
	wire _w22174_ ;
	wire _w22175_ ;
	wire _w22176_ ;
	wire _w22177_ ;
	wire _w22178_ ;
	wire _w22179_ ;
	wire _w22180_ ;
	wire _w22181_ ;
	wire _w22182_ ;
	wire _w22183_ ;
	wire _w22184_ ;
	wire _w22185_ ;
	wire _w22186_ ;
	wire _w22187_ ;
	wire _w22188_ ;
	wire _w22189_ ;
	wire _w22190_ ;
	wire _w22191_ ;
	wire _w22192_ ;
	wire _w22193_ ;
	wire _w22194_ ;
	wire _w22195_ ;
	wire _w22196_ ;
	wire _w22197_ ;
	wire _w22198_ ;
	wire _w22199_ ;
	wire _w22200_ ;
	wire _w22201_ ;
	wire _w22202_ ;
	wire _w22203_ ;
	wire _w22204_ ;
	wire _w22205_ ;
	wire _w22206_ ;
	wire _w22207_ ;
	wire _w22208_ ;
	wire _w22209_ ;
	wire _w22210_ ;
	wire _w22211_ ;
	wire _w22212_ ;
	wire _w22213_ ;
	wire _w22214_ ;
	wire _w22215_ ;
	wire _w22216_ ;
	wire _w22217_ ;
	wire _w22218_ ;
	wire _w22219_ ;
	wire _w22220_ ;
	wire _w22221_ ;
	wire _w22222_ ;
	wire _w22223_ ;
	wire _w22224_ ;
	wire _w22225_ ;
	wire _w22226_ ;
	wire _w22227_ ;
	wire _w22228_ ;
	wire _w22229_ ;
	wire _w22230_ ;
	wire _w22231_ ;
	wire _w22232_ ;
	wire _w22233_ ;
	wire _w22234_ ;
	wire _w22235_ ;
	wire _w22236_ ;
	wire _w22237_ ;
	wire _w22238_ ;
	wire _w22239_ ;
	wire _w22240_ ;
	wire _w22241_ ;
	wire _w22242_ ;
	wire _w22243_ ;
	wire _w22244_ ;
	wire _w22245_ ;
	wire _w22246_ ;
	wire _w22247_ ;
	wire _w22248_ ;
	wire _w22249_ ;
	wire _w22250_ ;
	wire _w22251_ ;
	wire _w22252_ ;
	wire _w22253_ ;
	wire _w22254_ ;
	wire _w22255_ ;
	wire _w22256_ ;
	wire _w22257_ ;
	wire _w22258_ ;
	wire _w22259_ ;
	wire _w22260_ ;
	wire _w22261_ ;
	wire _w22262_ ;
	wire _w22263_ ;
	wire _w22264_ ;
	wire _w22265_ ;
	wire _w22266_ ;
	wire _w22267_ ;
	wire _w22268_ ;
	wire _w22269_ ;
	wire _w22270_ ;
	wire _w22271_ ;
	wire _w22272_ ;
	wire _w22273_ ;
	wire _w22274_ ;
	wire _w22275_ ;
	wire _w22276_ ;
	wire _w22277_ ;
	wire _w22278_ ;
	wire _w22279_ ;
	wire _w22280_ ;
	wire _w22281_ ;
	wire _w22282_ ;
	wire _w22283_ ;
	wire _w22284_ ;
	wire _w22285_ ;
	wire _w22286_ ;
	wire _w22287_ ;
	wire _w22288_ ;
	wire _w22289_ ;
	wire _w22290_ ;
	wire _w22291_ ;
	wire _w22292_ ;
	wire _w22293_ ;
	wire _w22294_ ;
	wire _w22295_ ;
	wire _w22296_ ;
	wire _w22297_ ;
	wire _w22298_ ;
	wire _w22299_ ;
	wire _w22300_ ;
	wire _w22301_ ;
	wire _w22302_ ;
	wire _w22303_ ;
	wire _w22304_ ;
	wire _w22305_ ;
	wire _w22306_ ;
	wire _w22307_ ;
	wire _w22308_ ;
	wire _w22309_ ;
	wire _w22310_ ;
	wire _w22311_ ;
	wire _w22312_ ;
	wire _w22313_ ;
	wire _w22314_ ;
	wire _w22315_ ;
	wire _w22316_ ;
	wire _w22317_ ;
	wire _w22318_ ;
	wire _w22319_ ;
	wire _w22320_ ;
	wire _w22321_ ;
	wire _w22322_ ;
	wire _w22323_ ;
	wire _w22324_ ;
	wire _w22325_ ;
	wire _w22326_ ;
	wire _w22327_ ;
	wire _w22328_ ;
	wire _w22329_ ;
	wire _w22330_ ;
	wire _w22331_ ;
	wire _w22332_ ;
	wire _w22333_ ;
	wire _w22334_ ;
	wire _w22335_ ;
	wire _w22336_ ;
	wire _w22337_ ;
	wire _w22338_ ;
	wire _w22339_ ;
	wire _w22340_ ;
	wire _w22341_ ;
	wire _w22342_ ;
	wire _w22343_ ;
	wire _w22344_ ;
	wire _w22345_ ;
	wire _w22346_ ;
	wire _w22347_ ;
	wire _w22348_ ;
	wire _w22349_ ;
	wire _w22350_ ;
	wire _w22351_ ;
	wire _w22352_ ;
	wire _w22353_ ;
	wire _w22354_ ;
	wire _w22355_ ;
	wire _w22356_ ;
	wire _w22357_ ;
	wire _w22358_ ;
	wire _w22359_ ;
	wire _w22360_ ;
	wire _w22361_ ;
	wire _w22362_ ;
	wire _w22363_ ;
	wire _w22364_ ;
	wire _w22365_ ;
	wire _w22366_ ;
	wire _w22367_ ;
	wire _w22368_ ;
	wire _w22369_ ;
	wire _w22370_ ;
	wire _w22371_ ;
	wire _w22372_ ;
	wire _w22373_ ;
	wire _w22374_ ;
	wire _w22375_ ;
	wire _w22376_ ;
	wire _w22377_ ;
	wire _w22378_ ;
	wire _w22379_ ;
	wire _w22380_ ;
	wire _w22381_ ;
	wire _w22382_ ;
	wire _w22383_ ;
	wire _w22384_ ;
	wire _w22385_ ;
	wire _w22386_ ;
	wire _w22387_ ;
	wire _w22388_ ;
	wire _w22389_ ;
	wire _w22390_ ;
	wire _w22391_ ;
	wire _w22392_ ;
	wire _w22393_ ;
	wire _w22394_ ;
	wire _w22395_ ;
	wire _w22396_ ;
	wire _w22397_ ;
	wire _w22398_ ;
	wire _w22399_ ;
	wire _w22400_ ;
	wire _w22401_ ;
	wire _w22402_ ;
	wire _w22403_ ;
	wire _w22404_ ;
	wire _w22405_ ;
	wire _w22406_ ;
	wire _w22407_ ;
	wire _w22408_ ;
	wire _w22409_ ;
	wire _w22410_ ;
	wire _w22411_ ;
	wire _w22412_ ;
	wire _w22413_ ;
	wire _w22414_ ;
	wire _w22415_ ;
	wire _w22416_ ;
	wire _w22417_ ;
	wire _w22418_ ;
	wire _w22419_ ;
	wire _w22420_ ;
	wire _w22421_ ;
	wire _w22422_ ;
	wire _w22423_ ;
	wire _w22424_ ;
	wire _w22425_ ;
	wire _w22426_ ;
	wire _w22427_ ;
	wire _w22428_ ;
	wire _w22429_ ;
	wire _w22430_ ;
	wire _w22431_ ;
	wire _w22432_ ;
	wire _w22433_ ;
	wire _w22434_ ;
	wire _w22435_ ;
	wire _w22436_ ;
	wire _w22437_ ;
	wire _w22438_ ;
	wire _w22439_ ;
	wire _w22440_ ;
	wire _w22441_ ;
	wire _w22442_ ;
	wire _w22443_ ;
	wire _w22444_ ;
	wire _w22445_ ;
	wire _w22446_ ;
	wire _w22447_ ;
	wire _w22448_ ;
	wire _w22449_ ;
	wire _w22450_ ;
	wire _w22451_ ;
	wire _w22452_ ;
	wire _w22453_ ;
	wire _w22454_ ;
	wire _w22455_ ;
	wire _w22456_ ;
	wire _w22457_ ;
	wire _w22458_ ;
	wire _w22459_ ;
	wire _w22460_ ;
	wire _w22461_ ;
	wire _w22462_ ;
	wire _w22463_ ;
	wire _w22464_ ;
	wire _w22465_ ;
	wire _w22466_ ;
	wire _w22467_ ;
	wire _w22468_ ;
	wire _w22469_ ;
	wire _w22470_ ;
	wire _w22471_ ;
	wire _w22472_ ;
	wire _w22473_ ;
	wire _w22474_ ;
	wire _w22475_ ;
	wire _w22476_ ;
	wire _w22477_ ;
	wire _w22478_ ;
	wire _w22479_ ;
	wire _w22480_ ;
	wire _w22481_ ;
	wire _w22482_ ;
	wire _w22483_ ;
	wire _w22484_ ;
	wire _w22485_ ;
	wire _w22486_ ;
	wire _w22487_ ;
	wire _w22488_ ;
	wire _w22489_ ;
	wire _w22490_ ;
	wire _w22491_ ;
	wire _w22492_ ;
	wire _w22493_ ;
	wire _w22494_ ;
	wire _w22495_ ;
	wire _w22496_ ;
	wire _w22497_ ;
	wire _w22498_ ;
	wire _w22499_ ;
	wire _w22500_ ;
	wire _w22501_ ;
	wire _w22502_ ;
	wire _w22503_ ;
	wire _w22504_ ;
	wire _w22505_ ;
	wire _w22506_ ;
	wire _w22507_ ;
	wire _w22508_ ;
	wire _w22509_ ;
	wire _w22510_ ;
	wire _w22511_ ;
	wire _w22512_ ;
	wire _w22513_ ;
	wire _w22514_ ;
	wire _w22515_ ;
	wire _w22516_ ;
	wire _w22517_ ;
	wire _w22518_ ;
	wire _w22519_ ;
	wire _w22520_ ;
	wire _w22521_ ;
	wire _w22522_ ;
	wire _w22523_ ;
	wire _w22524_ ;
	wire _w22525_ ;
	wire _w22526_ ;
	wire _w22527_ ;
	wire _w22528_ ;
	wire _w22529_ ;
	wire _w22530_ ;
	wire _w22531_ ;
	wire _w22532_ ;
	wire _w22533_ ;
	wire _w22534_ ;
	wire _w22535_ ;
	wire _w22536_ ;
	wire _w22537_ ;
	wire _w22538_ ;
	wire _w22539_ ;
	wire _w22540_ ;
	wire _w22541_ ;
	wire _w22542_ ;
	wire _w22543_ ;
	wire _w22544_ ;
	wire _w22545_ ;
	wire _w22546_ ;
	wire _w22547_ ;
	wire _w22548_ ;
	wire _w22549_ ;
	wire _w22550_ ;
	wire _w22551_ ;
	wire _w22552_ ;
	wire _w22553_ ;
	wire _w22554_ ;
	wire _w22555_ ;
	wire _w22556_ ;
	wire _w22557_ ;
	wire _w22558_ ;
	wire _w22559_ ;
	wire _w22560_ ;
	wire _w22561_ ;
	wire _w22562_ ;
	wire _w22563_ ;
	wire _w22564_ ;
	wire _w22565_ ;
	wire _w22566_ ;
	wire _w22567_ ;
	wire _w22568_ ;
	wire _w22569_ ;
	wire _w22570_ ;
	wire _w22571_ ;
	wire _w22572_ ;
	wire _w22573_ ;
	wire _w22574_ ;
	wire _w22575_ ;
	wire _w22576_ ;
	wire _w22577_ ;
	wire _w22578_ ;
	wire _w22579_ ;
	wire _w22580_ ;
	wire _w22581_ ;
	wire _w22582_ ;
	wire _w22583_ ;
	wire _w22584_ ;
	wire _w22585_ ;
	wire _w22586_ ;
	wire _w22587_ ;
	wire _w22588_ ;
	wire _w22589_ ;
	wire _w22590_ ;
	wire _w22591_ ;
	wire _w22592_ ;
	wire _w22593_ ;
	wire _w22594_ ;
	wire _w22595_ ;
	wire _w22596_ ;
	wire _w22597_ ;
	wire _w22598_ ;
	wire _w22599_ ;
	wire _w22600_ ;
	wire _w22601_ ;
	wire _w22602_ ;
	wire _w22603_ ;
	wire _w22604_ ;
	wire _w22605_ ;
	wire _w22606_ ;
	wire _w22607_ ;
	wire _w22608_ ;
	wire _w22609_ ;
	wire _w22610_ ;
	wire _w22611_ ;
	wire _w22612_ ;
	wire _w22613_ ;
	wire _w22614_ ;
	wire _w22615_ ;
	wire _w22616_ ;
	wire _w22617_ ;
	wire _w22618_ ;
	wire _w22619_ ;
	wire _w22620_ ;
	wire _w22621_ ;
	wire _w22622_ ;
	wire _w22623_ ;
	wire _w22624_ ;
	wire _w22625_ ;
	wire _w22626_ ;
	wire _w22627_ ;
	wire _w22628_ ;
	wire _w22629_ ;
	wire _w22630_ ;
	wire _w22631_ ;
	wire _w22632_ ;
	wire _w22633_ ;
	wire _w22634_ ;
	wire _w22635_ ;
	wire _w22636_ ;
	wire _w22637_ ;
	wire _w22638_ ;
	wire _w22639_ ;
	wire _w22640_ ;
	wire _w22641_ ;
	wire _w22642_ ;
	wire _w22643_ ;
	wire _w22644_ ;
	wire _w22645_ ;
	wire _w22646_ ;
	wire _w22647_ ;
	wire _w22648_ ;
	wire _w22649_ ;
	wire _w22650_ ;
	wire _w22651_ ;
	wire _w22652_ ;
	wire _w22653_ ;
	LUT4 #(
		.INIT('hf35f)
	) name0 (
		\s15_msel_arb1_state_reg[2]/NET0131 ,
		\s15_msel_arb2_state_reg[2]/NET0131 ,
		\s15_msel_pri_out_reg[0]/NET0131 ,
		\s15_msel_pri_out_reg[1]/NET0131 ,
		_w1901_
	);
	LUT4 #(
		.INIT('h3ff5)
	) name1 (
		\s15_msel_arb0_state_reg[2]/NET0131 ,
		\s15_msel_arb3_state_reg[2]/NET0131 ,
		\s15_msel_pri_out_reg[0]/NET0131 ,
		\s15_msel_pri_out_reg[1]/NET0131 ,
		_w1902_
	);
	LUT2 #(
		.INIT('h8)
	) name2 (
		_w1901_,
		_w1902_,
		_w1903_
	);
	LUT4 #(
		.INIT('hff35)
	) name3 (
		\s15_msel_arb0_state_reg[0]/NET0131 ,
		\s15_msel_arb1_state_reg[0]/NET0131 ,
		\s15_msel_pri_out_reg[0]/NET0131 ,
		\s15_msel_pri_out_reg[1]/NET0131 ,
		_w1904_
	);
	LUT4 #(
		.INIT('h35ff)
	) name4 (
		\s15_msel_arb2_state_reg[0]/NET0131 ,
		\s15_msel_arb3_state_reg[0]/NET0131 ,
		\s15_msel_pri_out_reg[0]/NET0131 ,
		\s15_msel_pri_out_reg[1]/NET0131 ,
		_w1905_
	);
	LUT2 #(
		.INIT('h8)
	) name5 (
		_w1904_,
		_w1905_,
		_w1906_
	);
	LUT4 #(
		.INIT('h7000)
	) name6 (
		_w1901_,
		_w1902_,
		_w1904_,
		_w1905_,
		_w1907_
	);
	LUT4 #(
		.INIT('hff35)
	) name7 (
		\s15_msel_arb0_state_reg[1]/NET0131 ,
		\s15_msel_arb1_state_reg[1]/NET0131 ,
		\s15_msel_pri_out_reg[0]/NET0131 ,
		\s15_msel_pri_out_reg[1]/NET0131 ,
		_w1908_
	);
	LUT4 #(
		.INIT('h35ff)
	) name8 (
		\s15_msel_arb2_state_reg[1]/NET0131 ,
		\s15_msel_arb3_state_reg[1]/NET0131 ,
		\s15_msel_pri_out_reg[0]/NET0131 ,
		\s15_msel_pri_out_reg[1]/NET0131 ,
		_w1909_
	);
	LUT2 #(
		.INIT('h8)
	) name9 (
		_w1908_,
		_w1909_,
		_w1910_
	);
	LUT3 #(
		.INIT('h80)
	) name10 (
		\m4_addr_i[2]_pad ,
		_w1908_,
		_w1909_,
		_w1911_
	);
	LUT3 #(
		.INIT('h2a)
	) name11 (
		\m6_addr_i[2]_pad ,
		_w1908_,
		_w1909_,
		_w1912_
	);
	LUT3 #(
		.INIT('h57)
	) name12 (
		_w1907_,
		_w1911_,
		_w1912_,
		_w1913_
	);
	LUT4 #(
		.INIT('h8000)
	) name13 (
		_w1901_,
		_w1902_,
		_w1904_,
		_w1905_,
		_w1914_
	);
	LUT3 #(
		.INIT('h2a)
	) name14 (
		\m2_addr_i[2]_pad ,
		_w1908_,
		_w1909_,
		_w1915_
	);
	LUT3 #(
		.INIT('h80)
	) name15 (
		\m0_addr_i[2]_pad ,
		_w1908_,
		_w1909_,
		_w1916_
	);
	LUT3 #(
		.INIT('h57)
	) name16 (
		_w1914_,
		_w1915_,
		_w1916_,
		_w1917_
	);
	LUT4 #(
		.INIT('h0777)
	) name17 (
		_w1904_,
		_w1905_,
		_w1908_,
		_w1909_,
		_w1918_
	);
	LUT3 #(
		.INIT('h2a)
	) name18 (
		\m7_addr_i[2]_pad ,
		_w1901_,
		_w1902_,
		_w1919_
	);
	LUT4 #(
		.INIT('h7000)
	) name19 (
		_w1904_,
		_w1905_,
		_w1908_,
		_w1909_,
		_w1920_
	);
	LUT3 #(
		.INIT('h2a)
	) name20 (
		\m5_addr_i[2]_pad ,
		_w1901_,
		_w1902_,
		_w1921_
	);
	LUT4 #(
		.INIT('habef)
	) name21 (
		_w1906_,
		_w1910_,
		_w1919_,
		_w1921_,
		_w1922_
	);
	LUT3 #(
		.INIT('h80)
	) name22 (
		\m1_addr_i[2]_pad ,
		_w1901_,
		_w1902_,
		_w1923_
	);
	LUT3 #(
		.INIT('h80)
	) name23 (
		\m3_addr_i[2]_pad ,
		_w1901_,
		_w1902_,
		_w1924_
	);
	LUT4 #(
		.INIT('haebf)
	) name24 (
		_w1906_,
		_w1910_,
		_w1923_,
		_w1924_,
		_w1925_
	);
	LUT4 #(
		.INIT('h8000)
	) name25 (
		_w1913_,
		_w1917_,
		_w1922_,
		_w1925_,
		_w1926_
	);
	LUT4 #(
		.INIT('h7fff)
	) name26 (
		_w1913_,
		_w1917_,
		_w1922_,
		_w1925_,
		_w1927_
	);
	LUT3 #(
		.INIT('h2a)
	) name27 (
		\m7_addr_i[3]_pad ,
		_w1901_,
		_w1902_,
		_w1928_
	);
	LUT3 #(
		.INIT('h80)
	) name28 (
		\m3_addr_i[3]_pad ,
		_w1901_,
		_w1902_,
		_w1929_
	);
	LUT3 #(
		.INIT('h57)
	) name29 (
		_w1918_,
		_w1928_,
		_w1929_,
		_w1930_
	);
	LUT3 #(
		.INIT('h2a)
	) name30 (
		\m6_addr_i[3]_pad ,
		_w1908_,
		_w1909_,
		_w1931_
	);
	LUT3 #(
		.INIT('h2a)
	) name31 (
		\m5_addr_i[3]_pad ,
		_w1901_,
		_w1902_,
		_w1932_
	);
	LUT4 #(
		.INIT('h135f)
	) name32 (
		_w1907_,
		_w1920_,
		_w1931_,
		_w1932_,
		_w1933_
	);
	LUT3 #(
		.INIT('h80)
	) name33 (
		\m4_addr_i[3]_pad ,
		_w1908_,
		_w1909_,
		_w1934_
	);
	LUT3 #(
		.INIT('h80)
	) name34 (
		\m0_addr_i[3]_pad ,
		_w1908_,
		_w1909_,
		_w1935_
	);
	LUT4 #(
		.INIT('h37bf)
	) name35 (
		_w1903_,
		_w1906_,
		_w1934_,
		_w1935_,
		_w1936_
	);
	LUT3 #(
		.INIT('h80)
	) name36 (
		\m1_addr_i[3]_pad ,
		_w1901_,
		_w1902_,
		_w1937_
	);
	LUT3 #(
		.INIT('h2a)
	) name37 (
		\m2_addr_i[3]_pad ,
		_w1908_,
		_w1909_,
		_w1938_
	);
	LUT4 #(
		.INIT('h153f)
	) name38 (
		_w1914_,
		_w1920_,
		_w1937_,
		_w1938_,
		_w1939_
	);
	LUT4 #(
		.INIT('h8000)
	) name39 (
		_w1930_,
		_w1933_,
		_w1936_,
		_w1939_,
		_w1940_
	);
	LUT4 #(
		.INIT('h7fff)
	) name40 (
		_w1930_,
		_w1933_,
		_w1936_,
		_w1939_,
		_w1941_
	);
	LUT3 #(
		.INIT('h2a)
	) name41 (
		\m6_addr_i[5]_pad ,
		_w1908_,
		_w1909_,
		_w1942_
	);
	LUT3 #(
		.INIT('h2a)
	) name42 (
		\m7_addr_i[5]_pad ,
		_w1901_,
		_w1902_,
		_w1943_
	);
	LUT4 #(
		.INIT('h135f)
	) name43 (
		_w1907_,
		_w1918_,
		_w1942_,
		_w1943_,
		_w1944_
	);
	LUT3 #(
		.INIT('h80)
	) name44 (
		\m4_addr_i[5]_pad ,
		_w1908_,
		_w1909_,
		_w1945_
	);
	LUT3 #(
		.INIT('h2a)
	) name45 (
		\m5_addr_i[5]_pad ,
		_w1901_,
		_w1902_,
		_w1946_
	);
	LUT4 #(
		.INIT('h135f)
	) name46 (
		_w1907_,
		_w1920_,
		_w1945_,
		_w1946_,
		_w1947_
	);
	LUT3 #(
		.INIT('h80)
	) name47 (
		\m0_addr_i[5]_pad ,
		_w1908_,
		_w1909_,
		_w1948_
	);
	LUT3 #(
		.INIT('h80)
	) name48 (
		\m1_addr_i[5]_pad ,
		_w1901_,
		_w1902_,
		_w1949_
	);
	LUT4 #(
		.INIT('h135f)
	) name49 (
		_w1914_,
		_w1920_,
		_w1948_,
		_w1949_,
		_w1950_
	);
	LUT3 #(
		.INIT('h2a)
	) name50 (
		\m2_addr_i[5]_pad ,
		_w1908_,
		_w1909_,
		_w1951_
	);
	LUT3 #(
		.INIT('h80)
	) name51 (
		\m3_addr_i[5]_pad ,
		_w1901_,
		_w1902_,
		_w1952_
	);
	LUT4 #(
		.INIT('h135f)
	) name52 (
		_w1914_,
		_w1918_,
		_w1951_,
		_w1952_,
		_w1953_
	);
	LUT4 #(
		.INIT('h8000)
	) name53 (
		_w1944_,
		_w1947_,
		_w1950_,
		_w1953_,
		_w1954_
	);
	LUT4 #(
		.INIT('h7fff)
	) name54 (
		_w1944_,
		_w1947_,
		_w1950_,
		_w1953_,
		_w1955_
	);
	LUT3 #(
		.INIT('h80)
	) name55 (
		\m1_addr_i[4]_pad ,
		_w1901_,
		_w1902_,
		_w1956_
	);
	LUT3 #(
		.INIT('h80)
	) name56 (
		\m0_addr_i[4]_pad ,
		_w1908_,
		_w1909_,
		_w1957_
	);
	LUT4 #(
		.INIT('h153f)
	) name57 (
		_w1914_,
		_w1920_,
		_w1956_,
		_w1957_,
		_w1958_
	);
	LUT3 #(
		.INIT('h80)
	) name58 (
		\m4_addr_i[4]_pad ,
		_w1908_,
		_w1909_,
		_w1959_
	);
	LUT3 #(
		.INIT('h2a)
	) name59 (
		\m5_addr_i[4]_pad ,
		_w1901_,
		_w1902_,
		_w1960_
	);
	LUT4 #(
		.INIT('h135f)
	) name60 (
		_w1907_,
		_w1920_,
		_w1959_,
		_w1960_,
		_w1961_
	);
	LUT3 #(
		.INIT('h2a)
	) name61 (
		\m6_addr_i[4]_pad ,
		_w1908_,
		_w1909_,
		_w1962_
	);
	LUT3 #(
		.INIT('h2a)
	) name62 (
		\m7_addr_i[4]_pad ,
		_w1901_,
		_w1902_,
		_w1963_
	);
	LUT4 #(
		.INIT('h135f)
	) name63 (
		_w1907_,
		_w1918_,
		_w1962_,
		_w1963_,
		_w1964_
	);
	LUT3 #(
		.INIT('h80)
	) name64 (
		\m3_addr_i[4]_pad ,
		_w1901_,
		_w1902_,
		_w1965_
	);
	LUT3 #(
		.INIT('h2a)
	) name65 (
		\m2_addr_i[4]_pad ,
		_w1908_,
		_w1909_,
		_w1966_
	);
	LUT4 #(
		.INIT('h153f)
	) name66 (
		_w1914_,
		_w1918_,
		_w1965_,
		_w1966_,
		_w1967_
	);
	LUT4 #(
		.INIT('h8000)
	) name67 (
		_w1958_,
		_w1961_,
		_w1964_,
		_w1967_,
		_w1968_
	);
	LUT4 #(
		.INIT('h7fff)
	) name68 (
		_w1958_,
		_w1961_,
		_w1964_,
		_w1967_,
		_w1969_
	);
	LUT4 #(
		.INIT('h0040)
	) name69 (
		_w1926_,
		_w1940_,
		_w1954_,
		_w1968_,
		_w1970_
	);
	LUT4 #(
		.INIT('h1000)
	) name70 (
		_w1926_,
		_w1940_,
		_w1954_,
		_w1968_,
		_w1971_
	);
	LUT4 #(
		.INIT('h153f)
	) name71 (
		\rf_conf3_reg[11]/NET0131 ,
		\rf_conf5_reg[11]/NET0131 ,
		_w1970_,
		_w1971_,
		_w1972_
	);
	LUT4 #(
		.INIT('h0008)
	) name72 (
		_w1926_,
		_w1940_,
		_w1954_,
		_w1968_,
		_w1973_
	);
	LUT4 #(
		.INIT('h0002)
	) name73 (
		_w1926_,
		_w1940_,
		_w1954_,
		_w1968_,
		_w1974_
	);
	LUT4 #(
		.INIT('h135f)
	) name74 (
		\rf_conf12_reg[11]/NET0131 ,
		\rf_conf14_reg[11]/NET0131 ,
		_w1973_,
		_w1974_,
		_w1975_
	);
	LUT4 #(
		.INIT('h2000)
	) name75 (
		_w1926_,
		_w1940_,
		_w1954_,
		_w1968_,
		_w1976_
	);
	LUT4 #(
		.INIT('h4000)
	) name76 (
		_w1926_,
		_w1940_,
		_w1954_,
		_w1968_,
		_w1977_
	);
	LUT4 #(
		.INIT('h153f)
	) name77 (
		\rf_conf1_reg[11]/NET0131 ,
		\rf_conf2_reg[11]/NET0131 ,
		_w1976_,
		_w1977_,
		_w1978_
	);
	LUT4 #(
		.INIT('h8000)
	) name78 (
		_w1926_,
		_w1940_,
		_w1954_,
		_w1968_,
		_w1979_
	);
	LUT4 #(
		.INIT('h0080)
	) name79 (
		_w1926_,
		_w1940_,
		_w1954_,
		_w1968_,
		_w1980_
	);
	LUT4 #(
		.INIT('h135f)
	) name80 (
		\rf_conf0_reg[11]/NET0131 ,
		\rf_conf4_reg[11]/NET0131 ,
		_w1979_,
		_w1980_,
		_w1981_
	);
	LUT4 #(
		.INIT('h8000)
	) name81 (
		_w1972_,
		_w1975_,
		_w1978_,
		_w1981_,
		_w1982_
	);
	LUT4 #(
		.INIT('h0020)
	) name82 (
		_w1926_,
		_w1940_,
		_w1954_,
		_w1968_,
		_w1983_
	);
	LUT4 #(
		.INIT('h0010)
	) name83 (
		_w1926_,
		_w1940_,
		_w1954_,
		_w1968_,
		_w1984_
	);
	LUT4 #(
		.INIT('h135f)
	) name84 (
		\rf_conf6_reg[11]/NET0131 ,
		\rf_conf7_reg[11]/NET0131 ,
		_w1983_,
		_w1984_,
		_w1985_
	);
	LUT4 #(
		.INIT('h0800)
	) name85 (
		_w1926_,
		_w1940_,
		_w1954_,
		_w1968_,
		_w1986_
	);
	LUT4 #(
		.INIT('h0100)
	) name86 (
		_w1926_,
		_w1940_,
		_w1954_,
		_w1968_,
		_w1987_
	);
	LUT4 #(
		.INIT('h153f)
	) name87 (
		\rf_conf11_reg[11]/NET0131 ,
		\rf_conf8_reg[11]/NET0131 ,
		_w1986_,
		_w1987_,
		_w1988_
	);
	LUT4 #(
		.INIT('h0400)
	) name88 (
		_w1926_,
		_w1940_,
		_w1954_,
		_w1968_,
		_w1989_
	);
	LUT4 #(
		.INIT('h0200)
	) name89 (
		_w1926_,
		_w1940_,
		_w1954_,
		_w1968_,
		_w1990_
	);
	LUT4 #(
		.INIT('h153f)
	) name90 (
		\rf_conf10_reg[11]/NET0131 ,
		\rf_conf9_reg[11]/NET0131 ,
		_w1989_,
		_w1990_,
		_w1991_
	);
	LUT4 #(
		.INIT('h0004)
	) name91 (
		_w1926_,
		_w1940_,
		_w1954_,
		_w1968_,
		_w1992_
	);
	LUT4 #(
		.INIT('h0001)
	) name92 (
		_w1926_,
		_w1940_,
		_w1954_,
		_w1968_,
		_w1993_
	);
	LUT4 #(
		.INIT('h135f)
	) name93 (
		\rf_conf13_reg[11]/NET0131 ,
		\rf_conf15_reg[11]/NET0131 ,
		_w1992_,
		_w1993_,
		_w1994_
	);
	LUT4 #(
		.INIT('h8000)
	) name94 (
		_w1985_,
		_w1988_,
		_w1991_,
		_w1994_,
		_w1995_
	);
	LUT2 #(
		.INIT('h8)
	) name95 (
		\m5_s15_cyc_o_reg/NET0131 ,
		\s15_m5_cyc_r_reg/P0001 ,
		_w1996_
	);
	LUT3 #(
		.INIT('h70)
	) name96 (
		_w1901_,
		_w1902_,
		_w1996_,
		_w1997_
	);
	LUT2 #(
		.INIT('h8)
	) name97 (
		\m4_s15_cyc_o_reg/NET0131 ,
		\s15_m4_cyc_r_reg/P0001 ,
		_w1998_
	);
	LUT3 #(
		.INIT('h80)
	) name98 (
		_w1908_,
		_w1909_,
		_w1998_,
		_w1999_
	);
	LUT4 #(
		.INIT('h153f)
	) name99 (
		_w1907_,
		_w1920_,
		_w1997_,
		_w1999_,
		_w2000_
	);
	LUT2 #(
		.INIT('h8)
	) name100 (
		\m2_s15_cyc_o_reg/NET0131 ,
		\s15_m2_cyc_r_reg/P0001 ,
		_w2001_
	);
	LUT3 #(
		.INIT('h70)
	) name101 (
		_w1908_,
		_w1909_,
		_w2001_,
		_w2002_
	);
	LUT2 #(
		.INIT('h8)
	) name102 (
		\m3_s15_cyc_o_reg/NET0131 ,
		\s15_m3_cyc_r_reg/P0001 ,
		_w2003_
	);
	LUT3 #(
		.INIT('h80)
	) name103 (
		_w1901_,
		_w1902_,
		_w2003_,
		_w2004_
	);
	LUT4 #(
		.INIT('h135f)
	) name104 (
		_w1914_,
		_w1918_,
		_w2002_,
		_w2004_,
		_w2005_
	);
	LUT2 #(
		.INIT('h8)
	) name105 (
		\m0_s15_cyc_o_reg/NET0131 ,
		\s15_m0_cyc_r_reg/P0001 ,
		_w2006_
	);
	LUT3 #(
		.INIT('h80)
	) name106 (
		_w1908_,
		_w1909_,
		_w2006_,
		_w2007_
	);
	LUT2 #(
		.INIT('h8)
	) name107 (
		\m1_s15_cyc_o_reg/NET0131 ,
		\s15_m1_cyc_r_reg/P0001 ,
		_w2008_
	);
	LUT3 #(
		.INIT('h80)
	) name108 (
		_w1901_,
		_w1902_,
		_w2008_,
		_w2009_
	);
	LUT4 #(
		.INIT('h135f)
	) name109 (
		_w1914_,
		_w1920_,
		_w2007_,
		_w2009_,
		_w2010_
	);
	LUT2 #(
		.INIT('h8)
	) name110 (
		\m6_s15_cyc_o_reg/NET0131 ,
		\s15_m6_cyc_r_reg/P0001 ,
		_w2011_
	);
	LUT3 #(
		.INIT('h70)
	) name111 (
		_w1908_,
		_w1909_,
		_w2011_,
		_w2012_
	);
	LUT2 #(
		.INIT('h8)
	) name112 (
		\m7_s15_cyc_o_reg/NET0131 ,
		\s15_m7_cyc_r_reg/P0001 ,
		_w2013_
	);
	LUT3 #(
		.INIT('h70)
	) name113 (
		_w1901_,
		_w1902_,
		_w2013_,
		_w2014_
	);
	LUT4 #(
		.INIT('h135f)
	) name114 (
		_w1907_,
		_w1918_,
		_w2012_,
		_w2014_,
		_w2015_
	);
	LUT4 #(
		.INIT('h8000)
	) name115 (
		_w2000_,
		_w2005_,
		_w2010_,
		_w2015_,
		_w2016_
	);
	LUT3 #(
		.INIT('h80)
	) name116 (
		\m3_addr_i[27]_pad ,
		_w1901_,
		_w1902_,
		_w2017_
	);
	LUT3 #(
		.INIT('h2a)
	) name117 (
		\m7_addr_i[27]_pad ,
		_w1901_,
		_w1902_,
		_w2018_
	);
	LUT3 #(
		.INIT('h57)
	) name118 (
		_w1918_,
		_w2017_,
		_w2018_,
		_w2019_
	);
	LUT3 #(
		.INIT('h80)
	) name119 (
		\m4_addr_i[27]_pad ,
		_w1908_,
		_w1909_,
		_w2020_
	);
	LUT3 #(
		.INIT('h80)
	) name120 (
		\m1_addr_i[27]_pad ,
		_w1901_,
		_w1902_,
		_w2021_
	);
	LUT4 #(
		.INIT('h135f)
	) name121 (
		_w1907_,
		_w1920_,
		_w2020_,
		_w2021_,
		_w2022_
	);
	LUT3 #(
		.INIT('h80)
	) name122 (
		\m0_addr_i[27]_pad ,
		_w1908_,
		_w1909_,
		_w2023_
	);
	LUT3 #(
		.INIT('h2a)
	) name123 (
		\m5_addr_i[27]_pad ,
		_w1901_,
		_w1902_,
		_w2024_
	);
	LUT4 #(
		.INIT('h135f)
	) name124 (
		_w1914_,
		_w1920_,
		_w2023_,
		_w2024_,
		_w2025_
	);
	LUT3 #(
		.INIT('h2a)
	) name125 (
		\m2_addr_i[27]_pad ,
		_w1908_,
		_w1909_,
		_w2026_
	);
	LUT3 #(
		.INIT('h2a)
	) name126 (
		\m6_addr_i[27]_pad ,
		_w1908_,
		_w1909_,
		_w2027_
	);
	LUT4 #(
		.INIT('h3b7f)
	) name127 (
		_w1903_,
		_w1906_,
		_w2026_,
		_w2027_,
		_w2028_
	);
	LUT4 #(
		.INIT('h8000)
	) name128 (
		_w2019_,
		_w2022_,
		_w2025_,
		_w2028_,
		_w2029_
	);
	LUT4 #(
		.INIT('h7fff)
	) name129 (
		_w2019_,
		_w2022_,
		_w2025_,
		_w2028_,
		_w2030_
	);
	LUT3 #(
		.INIT('h2a)
	) name130 (
		\m2_addr_i[24]_pad ,
		_w1908_,
		_w1909_,
		_w2031_
	);
	LUT3 #(
		.INIT('h2a)
	) name131 (
		\m7_addr_i[24]_pad ,
		_w1901_,
		_w1902_,
		_w2032_
	);
	LUT4 #(
		.INIT('h135f)
	) name132 (
		_w1914_,
		_w1918_,
		_w2031_,
		_w2032_,
		_w2033_
	);
	LUT3 #(
		.INIT('h80)
	) name133 (
		\m0_addr_i[24]_pad ,
		_w1908_,
		_w1909_,
		_w2034_
	);
	LUT3 #(
		.INIT('h2a)
	) name134 (
		\m6_addr_i[24]_pad ,
		_w1908_,
		_w1909_,
		_w2035_
	);
	LUT4 #(
		.INIT('h3b7f)
	) name135 (
		_w1903_,
		_w1906_,
		_w2034_,
		_w2035_,
		_w2036_
	);
	LUT3 #(
		.INIT('h80)
	) name136 (
		\m1_addr_i[24]_pad ,
		_w1901_,
		_w1902_,
		_w2037_
	);
	LUT3 #(
		.INIT('h80)
	) name137 (
		\m4_addr_i[24]_pad ,
		_w1908_,
		_w1909_,
		_w2038_
	);
	LUT4 #(
		.INIT('h153f)
	) name138 (
		_w1907_,
		_w1920_,
		_w2037_,
		_w2038_,
		_w2039_
	);
	LUT3 #(
		.INIT('h2a)
	) name139 (
		\m5_addr_i[24]_pad ,
		_w1901_,
		_w1902_,
		_w2040_
	);
	LUT3 #(
		.INIT('h80)
	) name140 (
		\m3_addr_i[24]_pad ,
		_w1901_,
		_w1902_,
		_w2041_
	);
	LUT4 #(
		.INIT('haebf)
	) name141 (
		_w1906_,
		_w1910_,
		_w2040_,
		_w2041_,
		_w2042_
	);
	LUT4 #(
		.INIT('h8000)
	) name142 (
		_w2033_,
		_w2036_,
		_w2039_,
		_w2042_,
		_w2043_
	);
	LUT4 #(
		.INIT('h7fff)
	) name143 (
		_w2033_,
		_w2036_,
		_w2039_,
		_w2042_,
		_w2044_
	);
	LUT2 #(
		.INIT('h1)
	) name144 (
		_w2029_,
		_w2043_,
		_w2045_
	);
	LUT3 #(
		.INIT('h01)
	) name145 (
		_w2016_,
		_w2029_,
		_w2043_,
		_w2046_
	);
	LUT4 #(
		.INIT('h8000)
	) name146 (
		\m1_addr_i[28]_pad ,
		\m1_addr_i[29]_pad ,
		\m1_addr_i[30]_pad ,
		\m1_addr_i[31]_pad ,
		_w2047_
	);
	LUT4 #(
		.INIT('h8000)
	) name147 (
		\m1_stb_i_pad ,
		_w1901_,
		_w1902_,
		_w2047_,
		_w2048_
	);
	LUT4 #(
		.INIT('h8000)
	) name148 (
		\m0_addr_i[28]_pad ,
		\m0_addr_i[29]_pad ,
		\m0_addr_i[30]_pad ,
		\m0_addr_i[31]_pad ,
		_w2049_
	);
	LUT4 #(
		.INIT('h8000)
	) name149 (
		\m0_stb_i_pad ,
		_w1908_,
		_w1909_,
		_w2049_,
		_w2050_
	);
	LUT4 #(
		.INIT('h153f)
	) name150 (
		_w1914_,
		_w1920_,
		_w2048_,
		_w2050_,
		_w2051_
	);
	LUT4 #(
		.INIT('h8000)
	) name151 (
		\m7_addr_i[28]_pad ,
		\m7_addr_i[29]_pad ,
		\m7_addr_i[30]_pad ,
		\m7_addr_i[31]_pad ,
		_w2052_
	);
	LUT4 #(
		.INIT('h2a00)
	) name152 (
		\m7_stb_i_pad ,
		_w1901_,
		_w1902_,
		_w2052_,
		_w2053_
	);
	LUT4 #(
		.INIT('h8000)
	) name153 (
		\m6_addr_i[28]_pad ,
		\m6_addr_i[29]_pad ,
		\m6_addr_i[30]_pad ,
		\m6_addr_i[31]_pad ,
		_w2054_
	);
	LUT4 #(
		.INIT('h2a00)
	) name154 (
		\m6_stb_i_pad ,
		_w1908_,
		_w1909_,
		_w2054_,
		_w2055_
	);
	LUT4 #(
		.INIT('h153f)
	) name155 (
		_w1907_,
		_w1918_,
		_w2053_,
		_w2055_,
		_w2056_
	);
	LUT4 #(
		.INIT('h8000)
	) name156 (
		\m2_addr_i[28]_pad ,
		\m2_addr_i[29]_pad ,
		\m2_addr_i[30]_pad ,
		\m2_addr_i[31]_pad ,
		_w2057_
	);
	LUT4 #(
		.INIT('h2a00)
	) name157 (
		\m2_stb_i_pad ,
		_w1908_,
		_w1909_,
		_w2057_,
		_w2058_
	);
	LUT4 #(
		.INIT('h8000)
	) name158 (
		\m3_addr_i[28]_pad ,
		\m3_addr_i[29]_pad ,
		\m3_addr_i[30]_pad ,
		\m3_addr_i[31]_pad ,
		_w2059_
	);
	LUT4 #(
		.INIT('h8000)
	) name159 (
		\m3_stb_i_pad ,
		_w1901_,
		_w1902_,
		_w2059_,
		_w2060_
	);
	LUT4 #(
		.INIT('h135f)
	) name160 (
		_w1914_,
		_w1918_,
		_w2058_,
		_w2060_,
		_w2061_
	);
	LUT4 #(
		.INIT('h8000)
	) name161 (
		\m4_addr_i[28]_pad ,
		\m4_addr_i[29]_pad ,
		\m4_addr_i[30]_pad ,
		\m4_addr_i[31]_pad ,
		_w2062_
	);
	LUT4 #(
		.INIT('h8000)
	) name162 (
		\m4_stb_i_pad ,
		_w1908_,
		_w1909_,
		_w2062_,
		_w2063_
	);
	LUT4 #(
		.INIT('h8000)
	) name163 (
		\m5_addr_i[28]_pad ,
		\m5_addr_i[29]_pad ,
		\m5_addr_i[30]_pad ,
		\m5_addr_i[31]_pad ,
		_w2064_
	);
	LUT4 #(
		.INIT('h2a00)
	) name164 (
		\m5_stb_i_pad ,
		_w1901_,
		_w1902_,
		_w2064_,
		_w2065_
	);
	LUT4 #(
		.INIT('h135f)
	) name165 (
		_w1907_,
		_w1920_,
		_w2063_,
		_w2065_,
		_w2066_
	);
	LUT4 #(
		.INIT('h8000)
	) name166 (
		_w2051_,
		_w2056_,
		_w2061_,
		_w2066_,
		_w2067_
	);
	LUT4 #(
		.INIT('h7fff)
	) name167 (
		_w2051_,
		_w2056_,
		_w2061_,
		_w2066_,
		_w2068_
	);
	LUT3 #(
		.INIT('h2a)
	) name168 (
		\m7_addr_i[25]_pad ,
		_w1901_,
		_w1902_,
		_w2069_
	);
	LUT3 #(
		.INIT('h2a)
	) name169 (
		\m5_addr_i[25]_pad ,
		_w1901_,
		_w1902_,
		_w2070_
	);
	LUT4 #(
		.INIT('habef)
	) name170 (
		_w1906_,
		_w1910_,
		_w2069_,
		_w2070_,
		_w2071_
	);
	LUT3 #(
		.INIT('h2a)
	) name171 (
		\m6_addr_i[25]_pad ,
		_w1908_,
		_w1909_,
		_w2072_
	);
	LUT3 #(
		.INIT('h80)
	) name172 (
		\m1_addr_i[25]_pad ,
		_w1901_,
		_w1902_,
		_w2073_
	);
	LUT4 #(
		.INIT('h135f)
	) name173 (
		_w1907_,
		_w1920_,
		_w2072_,
		_w2073_,
		_w2074_
	);
	LUT3 #(
		.INIT('h80)
	) name174 (
		\m3_addr_i[25]_pad ,
		_w1901_,
		_w1902_,
		_w2075_
	);
	LUT3 #(
		.INIT('h80)
	) name175 (
		\m4_addr_i[25]_pad ,
		_w1908_,
		_w1909_,
		_w2076_
	);
	LUT4 #(
		.INIT('h153f)
	) name176 (
		_w1907_,
		_w1918_,
		_w2075_,
		_w2076_,
		_w2077_
	);
	LUT3 #(
		.INIT('h80)
	) name177 (
		\m0_addr_i[25]_pad ,
		_w1908_,
		_w1909_,
		_w2078_
	);
	LUT3 #(
		.INIT('h2a)
	) name178 (
		\m2_addr_i[25]_pad ,
		_w1908_,
		_w1909_,
		_w2079_
	);
	LUT3 #(
		.INIT('h57)
	) name179 (
		_w1914_,
		_w2078_,
		_w2079_,
		_w2080_
	);
	LUT4 #(
		.INIT('h8000)
	) name180 (
		_w2071_,
		_w2074_,
		_w2077_,
		_w2080_,
		_w2081_
	);
	LUT4 #(
		.INIT('h7fff)
	) name181 (
		_w2071_,
		_w2074_,
		_w2077_,
		_w2080_,
		_w2082_
	);
	LUT3 #(
		.INIT('h80)
	) name182 (
		\m1_addr_i[26]_pad ,
		_w1901_,
		_w1902_,
		_w2083_
	);
	LUT3 #(
		.INIT('h2a)
	) name183 (
		\m2_addr_i[26]_pad ,
		_w1908_,
		_w1909_,
		_w2084_
	);
	LUT4 #(
		.INIT('h153f)
	) name184 (
		_w1914_,
		_w1920_,
		_w2083_,
		_w2084_,
		_w2085_
	);
	LUT3 #(
		.INIT('h2a)
	) name185 (
		\m7_addr_i[26]_pad ,
		_w1901_,
		_w1902_,
		_w2086_
	);
	LUT3 #(
		.INIT('h80)
	) name186 (
		\m3_addr_i[26]_pad ,
		_w1901_,
		_w1902_,
		_w2087_
	);
	LUT3 #(
		.INIT('h57)
	) name187 (
		_w1918_,
		_w2086_,
		_w2087_,
		_w2088_
	);
	LUT3 #(
		.INIT('h2a)
	) name188 (
		\m6_addr_i[26]_pad ,
		_w1908_,
		_w1909_,
		_w2089_
	);
	LUT3 #(
		.INIT('h2a)
	) name189 (
		\m5_addr_i[26]_pad ,
		_w1901_,
		_w1902_,
		_w2090_
	);
	LUT4 #(
		.INIT('h135f)
	) name190 (
		_w1907_,
		_w1920_,
		_w2089_,
		_w2090_,
		_w2091_
	);
	LUT3 #(
		.INIT('h80)
	) name191 (
		\m4_addr_i[26]_pad ,
		_w1908_,
		_w1909_,
		_w2092_
	);
	LUT3 #(
		.INIT('h80)
	) name192 (
		\m0_addr_i[26]_pad ,
		_w1908_,
		_w1909_,
		_w2093_
	);
	LUT4 #(
		.INIT('h37bf)
	) name193 (
		_w1903_,
		_w1906_,
		_w2092_,
		_w2093_,
		_w2094_
	);
	LUT4 #(
		.INIT('h8000)
	) name194 (
		_w2085_,
		_w2088_,
		_w2091_,
		_w2094_,
		_w2095_
	);
	LUT4 #(
		.INIT('h7fff)
	) name195 (
		_w2085_,
		_w2088_,
		_w2091_,
		_w2094_,
		_w2096_
	);
	LUT3 #(
		.INIT('h01)
	) name196 (
		_w2067_,
		_w2081_,
		_w2095_,
		_w2097_
	);
	LUT2 #(
		.INIT('h8)
	) name197 (
		_w2046_,
		_w2097_,
		_w2098_
	);
	LUT3 #(
		.INIT('h70)
	) name198 (
		_w1982_,
		_w1995_,
		_w2098_,
		_w2099_
	);
	LUT4 #(
		.INIT('h153f)
	) name199 (
		\rf_conf11_reg[0]/NET0131 ,
		\rf_conf8_reg[0]/NET0131 ,
		_w1986_,
		_w1987_,
		_w2100_
	);
	LUT4 #(
		.INIT('h135f)
	) name200 (
		\rf_conf6_reg[0]/NET0131 ,
		\rf_conf7_reg[0]/NET0131 ,
		_w1983_,
		_w1984_,
		_w2101_
	);
	LUT4 #(
		.INIT('h135f)
	) name201 (
		\rf_conf12_reg[0]/NET0131 ,
		\rf_conf14_reg[0]/NET0131 ,
		_w1973_,
		_w1974_,
		_w2102_
	);
	LUT4 #(
		.INIT('h153f)
	) name202 (
		\rf_conf3_reg[0]/NET0131 ,
		\rf_conf5_reg[0]/NET0131 ,
		_w1970_,
		_w1971_,
		_w2103_
	);
	LUT4 #(
		.INIT('h8000)
	) name203 (
		_w2100_,
		_w2101_,
		_w2102_,
		_w2103_,
		_w2104_
	);
	LUT4 #(
		.INIT('h153f)
	) name204 (
		\rf_conf1_reg[0]/NET0131 ,
		\rf_conf2_reg[0]/NET0131 ,
		_w1976_,
		_w1977_,
		_w2105_
	);
	LUT4 #(
		.INIT('h135f)
	) name205 (
		\rf_conf13_reg[0]/NET0131 ,
		\rf_conf15_reg[0]/NET0131 ,
		_w1992_,
		_w1993_,
		_w2106_
	);
	LUT4 #(
		.INIT('h153f)
	) name206 (
		\rf_conf10_reg[0]/NET0131 ,
		\rf_conf9_reg[0]/NET0131 ,
		_w1989_,
		_w1990_,
		_w2107_
	);
	LUT4 #(
		.INIT('h135f)
	) name207 (
		\rf_conf0_reg[0]/NET0131 ,
		\rf_conf4_reg[0]/NET0131 ,
		_w1979_,
		_w1980_,
		_w2108_
	);
	LUT4 #(
		.INIT('h8000)
	) name208 (
		_w2105_,
		_w2106_,
		_w2107_,
		_w2108_,
		_w2109_
	);
	LUT3 #(
		.INIT('h2a)
	) name209 (
		_w2098_,
		_w2104_,
		_w2109_,
		_w2110_
	);
	LUT4 #(
		.INIT('h135f)
	) name210 (
		\rf_conf12_reg[10]/NET0131 ,
		\rf_conf14_reg[10]/NET0131 ,
		_w1973_,
		_w1974_,
		_w2111_
	);
	LUT4 #(
		.INIT('h135f)
	) name211 (
		\rf_conf6_reg[10]/NET0131 ,
		\rf_conf7_reg[10]/NET0131 ,
		_w1983_,
		_w1984_,
		_w2112_
	);
	LUT4 #(
		.INIT('h153f)
	) name212 (
		\rf_conf11_reg[10]/NET0131 ,
		\rf_conf8_reg[10]/NET0131 ,
		_w1986_,
		_w1987_,
		_w2113_
	);
	LUT4 #(
		.INIT('h153f)
	) name213 (
		\rf_conf1_reg[10]/NET0131 ,
		\rf_conf2_reg[10]/NET0131 ,
		_w1976_,
		_w1977_,
		_w2114_
	);
	LUT4 #(
		.INIT('h8000)
	) name214 (
		_w2111_,
		_w2112_,
		_w2113_,
		_w2114_,
		_w2115_
	);
	LUT4 #(
		.INIT('h153f)
	) name215 (
		\rf_conf3_reg[10]/NET0131 ,
		\rf_conf5_reg[10]/NET0131 ,
		_w1970_,
		_w1971_,
		_w2116_
	);
	LUT4 #(
		.INIT('h135f)
	) name216 (
		\rf_conf13_reg[10]/NET0131 ,
		\rf_conf15_reg[10]/NET0131 ,
		_w1992_,
		_w1993_,
		_w2117_
	);
	LUT4 #(
		.INIT('h135f)
	) name217 (
		\rf_conf0_reg[10]/NET0131 ,
		\rf_conf4_reg[10]/NET0131 ,
		_w1979_,
		_w1980_,
		_w2118_
	);
	LUT4 #(
		.INIT('h153f)
	) name218 (
		\rf_conf10_reg[10]/NET0131 ,
		\rf_conf9_reg[10]/NET0131 ,
		_w1989_,
		_w1990_,
		_w2119_
	);
	LUT4 #(
		.INIT('h8000)
	) name219 (
		_w2116_,
		_w2117_,
		_w2118_,
		_w2119_,
		_w2120_
	);
	LUT3 #(
		.INIT('h2a)
	) name220 (
		_w2098_,
		_w2115_,
		_w2120_,
		_w2121_
	);
	LUT4 #(
		.INIT('h153f)
	) name221 (
		\rf_conf10_reg[12]/NET0131 ,
		\rf_conf9_reg[12]/NET0131 ,
		_w1989_,
		_w1990_,
		_w2122_
	);
	LUT4 #(
		.INIT('h135f)
	) name222 (
		\rf_conf12_reg[12]/NET0131 ,
		\rf_conf14_reg[12]/NET0131 ,
		_w1973_,
		_w1974_,
		_w2123_
	);
	LUT4 #(
		.INIT('h135f)
	) name223 (
		\rf_conf0_reg[12]/NET0131 ,
		\rf_conf4_reg[12]/NET0131 ,
		_w1979_,
		_w1980_,
		_w2124_
	);
	LUT4 #(
		.INIT('h135f)
	) name224 (
		\rf_conf13_reg[12]/NET0131 ,
		\rf_conf15_reg[12]/NET0131 ,
		_w1992_,
		_w1993_,
		_w2125_
	);
	LUT4 #(
		.INIT('h8000)
	) name225 (
		_w2122_,
		_w2123_,
		_w2124_,
		_w2125_,
		_w2126_
	);
	LUT4 #(
		.INIT('h135f)
	) name226 (
		\rf_conf6_reg[12]/NET0131 ,
		\rf_conf7_reg[12]/NET0131 ,
		_w1983_,
		_w1984_,
		_w2127_
	);
	LUT4 #(
		.INIT('h153f)
	) name227 (
		\rf_conf11_reg[12]/NET0131 ,
		\rf_conf8_reg[12]/NET0131 ,
		_w1986_,
		_w1987_,
		_w2128_
	);
	LUT4 #(
		.INIT('h153f)
	) name228 (
		\rf_conf3_reg[12]/NET0131 ,
		\rf_conf5_reg[12]/NET0131 ,
		_w1970_,
		_w1971_,
		_w2129_
	);
	LUT4 #(
		.INIT('h153f)
	) name229 (
		\rf_conf1_reg[12]/NET0131 ,
		\rf_conf2_reg[12]/NET0131 ,
		_w1976_,
		_w1977_,
		_w2130_
	);
	LUT4 #(
		.INIT('h8000)
	) name230 (
		_w2127_,
		_w2128_,
		_w2129_,
		_w2130_,
		_w2131_
	);
	LUT3 #(
		.INIT('h2a)
	) name231 (
		_w2098_,
		_w2126_,
		_w2131_,
		_w2132_
	);
	LUT4 #(
		.INIT('h135f)
	) name232 (
		\rf_conf12_reg[13]/NET0131 ,
		\rf_conf14_reg[13]/NET0131 ,
		_w1973_,
		_w1974_,
		_w2133_
	);
	LUT4 #(
		.INIT('h153f)
	) name233 (
		\rf_conf10_reg[13]/NET0131 ,
		\rf_conf9_reg[13]/NET0131 ,
		_w1989_,
		_w1990_,
		_w2134_
	);
	LUT4 #(
		.INIT('h153f)
	) name234 (
		\rf_conf11_reg[13]/NET0131 ,
		\rf_conf8_reg[13]/NET0131 ,
		_w1986_,
		_w1987_,
		_w2135_
	);
	LUT4 #(
		.INIT('h153f)
	) name235 (
		\rf_conf1_reg[13]/NET0131 ,
		\rf_conf2_reg[13]/NET0131 ,
		_w1976_,
		_w1977_,
		_w2136_
	);
	LUT4 #(
		.INIT('h8000)
	) name236 (
		_w2133_,
		_w2134_,
		_w2135_,
		_w2136_,
		_w2137_
	);
	LUT4 #(
		.INIT('h153f)
	) name237 (
		\rf_conf3_reg[13]/NET0131 ,
		\rf_conf5_reg[13]/NET0131 ,
		_w1970_,
		_w1971_,
		_w2138_
	);
	LUT4 #(
		.INIT('h135f)
	) name238 (
		\rf_conf6_reg[13]/NET0131 ,
		\rf_conf7_reg[13]/NET0131 ,
		_w1983_,
		_w1984_,
		_w2139_
	);
	LUT4 #(
		.INIT('h135f)
	) name239 (
		\rf_conf13_reg[13]/NET0131 ,
		\rf_conf15_reg[13]/NET0131 ,
		_w1992_,
		_w1993_,
		_w2140_
	);
	LUT4 #(
		.INIT('h135f)
	) name240 (
		\rf_conf0_reg[13]/NET0131 ,
		\rf_conf4_reg[13]/NET0131 ,
		_w1979_,
		_w1980_,
		_w2141_
	);
	LUT4 #(
		.INIT('h8000)
	) name241 (
		_w2138_,
		_w2139_,
		_w2140_,
		_w2141_,
		_w2142_
	);
	LUT3 #(
		.INIT('h2a)
	) name242 (
		_w2098_,
		_w2137_,
		_w2142_,
		_w2143_
	);
	LUT4 #(
		.INIT('h135f)
	) name243 (
		\rf_conf6_reg[14]/NET0131 ,
		\rf_conf7_reg[14]/NET0131 ,
		_w1983_,
		_w1984_,
		_w2144_
	);
	LUT4 #(
		.INIT('h153f)
	) name244 (
		\rf_conf11_reg[14]/NET0131 ,
		\rf_conf8_reg[14]/NET0131 ,
		_w1986_,
		_w1987_,
		_w2145_
	);
	LUT4 #(
		.INIT('h135f)
	) name245 (
		\rf_conf13_reg[14]/NET0131 ,
		\rf_conf15_reg[14]/NET0131 ,
		_w1992_,
		_w1993_,
		_w2146_
	);
	LUT4 #(
		.INIT('h135f)
	) name246 (
		\rf_conf0_reg[14]/NET0131 ,
		\rf_conf4_reg[14]/NET0131 ,
		_w1979_,
		_w1980_,
		_w2147_
	);
	LUT4 #(
		.INIT('h8000)
	) name247 (
		_w2144_,
		_w2145_,
		_w2146_,
		_w2147_,
		_w2148_
	);
	LUT4 #(
		.INIT('h153f)
	) name248 (
		\rf_conf10_reg[14]/NET0131 ,
		\rf_conf9_reg[14]/NET0131 ,
		_w1989_,
		_w1990_,
		_w2149_
	);
	LUT4 #(
		.INIT('h153f)
	) name249 (
		\rf_conf2_reg[14]/NET0131 ,
		\rf_conf3_reg[14]/NET0131 ,
		_w1971_,
		_w1976_,
		_w2150_
	);
	LUT4 #(
		.INIT('h135f)
	) name250 (
		\rf_conf14_reg[14]/NET0131 ,
		\rf_conf1_reg[14]/NET0131 ,
		_w1974_,
		_w1977_,
		_w2151_
	);
	LUT4 #(
		.INIT('h153f)
	) name251 (
		\rf_conf12_reg[14]/NET0131 ,
		\rf_conf5_reg[14]/NET0131 ,
		_w1970_,
		_w1973_,
		_w2152_
	);
	LUT4 #(
		.INIT('h8000)
	) name252 (
		_w2149_,
		_w2150_,
		_w2151_,
		_w2152_,
		_w2153_
	);
	LUT3 #(
		.INIT('h2a)
	) name253 (
		_w2098_,
		_w2148_,
		_w2153_,
		_w2154_
	);
	LUT4 #(
		.INIT('h135f)
	) name254 (
		\rf_conf12_reg[15]/NET0131 ,
		\rf_conf14_reg[15]/NET0131 ,
		_w1973_,
		_w1974_,
		_w2155_
	);
	LUT4 #(
		.INIT('h135f)
	) name255 (
		\rf_conf6_reg[15]/NET0131 ,
		\rf_conf7_reg[15]/NET0131 ,
		_w1983_,
		_w1984_,
		_w2156_
	);
	LUT4 #(
		.INIT('h153f)
	) name256 (
		\rf_conf11_reg[15]/NET0131 ,
		\rf_conf8_reg[15]/NET0131 ,
		_w1986_,
		_w1987_,
		_w2157_
	);
	LUT4 #(
		.INIT('h153f)
	) name257 (
		\rf_conf1_reg[15]/NET0131 ,
		\rf_conf2_reg[15]/NET0131 ,
		_w1976_,
		_w1977_,
		_w2158_
	);
	LUT4 #(
		.INIT('h8000)
	) name258 (
		_w2155_,
		_w2156_,
		_w2157_,
		_w2158_,
		_w2159_
	);
	LUT4 #(
		.INIT('h153f)
	) name259 (
		\rf_conf3_reg[15]/NET0131 ,
		\rf_conf5_reg[15]/NET0131 ,
		_w1970_,
		_w1971_,
		_w2160_
	);
	LUT4 #(
		.INIT('h153f)
	) name260 (
		\rf_conf10_reg[15]/NET0131 ,
		\rf_conf9_reg[15]/NET0131 ,
		_w1989_,
		_w1990_,
		_w2161_
	);
	LUT4 #(
		.INIT('h135f)
	) name261 (
		\rf_conf0_reg[15]/NET0131 ,
		\rf_conf4_reg[15]/NET0131 ,
		_w1979_,
		_w1980_,
		_w2162_
	);
	LUT4 #(
		.INIT('h135f)
	) name262 (
		\rf_conf13_reg[15]/NET0131 ,
		\rf_conf15_reg[15]/NET0131 ,
		_w1992_,
		_w1993_,
		_w2163_
	);
	LUT4 #(
		.INIT('h8000)
	) name263 (
		_w2160_,
		_w2161_,
		_w2162_,
		_w2163_,
		_w2164_
	);
	LUT3 #(
		.INIT('h2a)
	) name264 (
		_w2098_,
		_w2159_,
		_w2164_,
		_w2165_
	);
	LUT4 #(
		.INIT('h135f)
	) name265 (
		\rf_conf0_reg[1]/NET0131 ,
		\rf_conf4_reg[1]/NET0131 ,
		_w1979_,
		_w1980_,
		_w2166_
	);
	LUT4 #(
		.INIT('h153f)
	) name266 (
		\rf_conf11_reg[1]/NET0131 ,
		\rf_conf8_reg[1]/NET0131 ,
		_w1986_,
		_w1987_,
		_w2167_
	);
	LUT4 #(
		.INIT('h135f)
	) name267 (
		\rf_conf6_reg[1]/NET0131 ,
		\rf_conf7_reg[1]/NET0131 ,
		_w1983_,
		_w1984_,
		_w2168_
	);
	LUT4 #(
		.INIT('h135f)
	) name268 (
		\rf_conf13_reg[1]/NET0131 ,
		\rf_conf15_reg[1]/NET0131 ,
		_w1992_,
		_w1993_,
		_w2169_
	);
	LUT4 #(
		.INIT('h8000)
	) name269 (
		_w2166_,
		_w2167_,
		_w2168_,
		_w2169_,
		_w2170_
	);
	LUT4 #(
		.INIT('h153f)
	) name270 (
		\rf_conf10_reg[1]/NET0131 ,
		\rf_conf9_reg[1]/NET0131 ,
		_w1989_,
		_w1990_,
		_w2171_
	);
	LUT4 #(
		.INIT('h135f)
	) name271 (
		\rf_conf12_reg[1]/NET0131 ,
		\rf_conf14_reg[1]/NET0131 ,
		_w1973_,
		_w1974_,
		_w2172_
	);
	LUT4 #(
		.INIT('h153f)
	) name272 (
		\rf_conf3_reg[1]/NET0131 ,
		\rf_conf5_reg[1]/NET0131 ,
		_w1970_,
		_w1971_,
		_w2173_
	);
	LUT4 #(
		.INIT('h153f)
	) name273 (
		\rf_conf1_reg[1]/NET0131 ,
		\rf_conf2_reg[1]/NET0131 ,
		_w1976_,
		_w1977_,
		_w2174_
	);
	LUT4 #(
		.INIT('h8000)
	) name274 (
		_w2171_,
		_w2172_,
		_w2173_,
		_w2174_,
		_w2175_
	);
	LUT3 #(
		.INIT('h2a)
	) name275 (
		_w2098_,
		_w2170_,
		_w2175_,
		_w2176_
	);
	LUT4 #(
		.INIT('h135f)
	) name276 (
		\rf_conf0_reg[2]/NET0131 ,
		\rf_conf4_reg[2]/NET0131 ,
		_w1979_,
		_w1980_,
		_w2177_
	);
	LUT4 #(
		.INIT('h153f)
	) name277 (
		\rf_conf3_reg[2]/NET0131 ,
		\rf_conf5_reg[2]/NET0131 ,
		_w1970_,
		_w1971_,
		_w2178_
	);
	LUT4 #(
		.INIT('h135f)
	) name278 (
		\rf_conf13_reg[2]/NET0131 ,
		\rf_conf15_reg[2]/NET0131 ,
		_w1992_,
		_w1993_,
		_w2179_
	);
	LUT4 #(
		.INIT('h153f)
	) name279 (
		\rf_conf10_reg[2]/NET0131 ,
		\rf_conf9_reg[2]/NET0131 ,
		_w1989_,
		_w1990_,
		_w2180_
	);
	LUT4 #(
		.INIT('h8000)
	) name280 (
		_w2177_,
		_w2178_,
		_w2179_,
		_w2180_,
		_w2181_
	);
	LUT4 #(
		.INIT('h135f)
	) name281 (
		\rf_conf6_reg[2]/NET0131 ,
		\rf_conf7_reg[2]/NET0131 ,
		_w1983_,
		_w1984_,
		_w2182_
	);
	LUT4 #(
		.INIT('h153f)
	) name282 (
		\rf_conf11_reg[2]/NET0131 ,
		\rf_conf8_reg[2]/NET0131 ,
		_w1986_,
		_w1987_,
		_w2183_
	);
	LUT4 #(
		.INIT('h153f)
	) name283 (
		\rf_conf1_reg[2]/NET0131 ,
		\rf_conf2_reg[2]/NET0131 ,
		_w1976_,
		_w1977_,
		_w2184_
	);
	LUT4 #(
		.INIT('h135f)
	) name284 (
		\rf_conf12_reg[2]/NET0131 ,
		\rf_conf14_reg[2]/NET0131 ,
		_w1973_,
		_w1974_,
		_w2185_
	);
	LUT4 #(
		.INIT('h8000)
	) name285 (
		_w2182_,
		_w2183_,
		_w2184_,
		_w2185_,
		_w2186_
	);
	LUT3 #(
		.INIT('h2a)
	) name286 (
		_w2098_,
		_w2181_,
		_w2186_,
		_w2187_
	);
	LUT4 #(
		.INIT('h153f)
	) name287 (
		\rf_conf3_reg[3]/NET0131 ,
		\rf_conf5_reg[3]/NET0131 ,
		_w1970_,
		_w1971_,
		_w2188_
	);
	LUT4 #(
		.INIT('h135f)
	) name288 (
		\rf_conf13_reg[3]/NET0131 ,
		\rf_conf15_reg[3]/NET0131 ,
		_w1992_,
		_w1993_,
		_w2189_
	);
	LUT4 #(
		.INIT('h153f)
	) name289 (
		\rf_conf11_reg[3]/NET0131 ,
		\rf_conf8_reg[3]/NET0131 ,
		_w1986_,
		_w1987_,
		_w2190_
	);
	LUT4 #(
		.INIT('h153f)
	) name290 (
		\rf_conf1_reg[3]/NET0131 ,
		\rf_conf2_reg[3]/NET0131 ,
		_w1976_,
		_w1977_,
		_w2191_
	);
	LUT4 #(
		.INIT('h8000)
	) name291 (
		_w2188_,
		_w2189_,
		_w2190_,
		_w2191_,
		_w2192_
	);
	LUT4 #(
		.INIT('h135f)
	) name292 (
		\rf_conf12_reg[3]/NET0131 ,
		\rf_conf14_reg[3]/NET0131 ,
		_w1973_,
		_w1974_,
		_w2193_
	);
	LUT4 #(
		.INIT('h153f)
	) name293 (
		\rf_conf10_reg[3]/NET0131 ,
		\rf_conf9_reg[3]/NET0131 ,
		_w1989_,
		_w1990_,
		_w2194_
	);
	LUT4 #(
		.INIT('h135f)
	) name294 (
		\rf_conf6_reg[3]/NET0131 ,
		\rf_conf7_reg[3]/NET0131 ,
		_w1983_,
		_w1984_,
		_w2195_
	);
	LUT4 #(
		.INIT('h135f)
	) name295 (
		\rf_conf0_reg[3]/NET0131 ,
		\rf_conf4_reg[3]/NET0131 ,
		_w1979_,
		_w1980_,
		_w2196_
	);
	LUT4 #(
		.INIT('h8000)
	) name296 (
		_w2193_,
		_w2194_,
		_w2195_,
		_w2196_,
		_w2197_
	);
	LUT3 #(
		.INIT('h2a)
	) name297 (
		_w2098_,
		_w2192_,
		_w2197_,
		_w2198_
	);
	LUT4 #(
		.INIT('h135f)
	) name298 (
		\rf_conf6_reg[4]/NET0131 ,
		\rf_conf7_reg[4]/NET0131 ,
		_w1983_,
		_w1984_,
		_w2199_
	);
	LUT4 #(
		.INIT('h153f)
	) name299 (
		\rf_conf11_reg[4]/NET0131 ,
		\rf_conf8_reg[4]/NET0131 ,
		_w1986_,
		_w1987_,
		_w2200_
	);
	LUT4 #(
		.INIT('h135f)
	) name300 (
		\rf_conf13_reg[4]/NET0131 ,
		\rf_conf15_reg[4]/NET0131 ,
		_w1992_,
		_w1993_,
		_w2201_
	);
	LUT4 #(
		.INIT('h153f)
	) name301 (
		\rf_conf10_reg[4]/NET0131 ,
		\rf_conf9_reg[4]/NET0131 ,
		_w1989_,
		_w1990_,
		_w2202_
	);
	LUT4 #(
		.INIT('h8000)
	) name302 (
		_w2199_,
		_w2200_,
		_w2201_,
		_w2202_,
		_w2203_
	);
	LUT4 #(
		.INIT('h135f)
	) name303 (
		\rf_conf0_reg[4]/NET0131 ,
		\rf_conf4_reg[4]/NET0131 ,
		_w1979_,
		_w1980_,
		_w2204_
	);
	LUT4 #(
		.INIT('h135f)
	) name304 (
		\rf_conf12_reg[4]/NET0131 ,
		\rf_conf14_reg[4]/NET0131 ,
		_w1973_,
		_w1974_,
		_w2205_
	);
	LUT4 #(
		.INIT('h153f)
	) name305 (
		\rf_conf3_reg[4]/NET0131 ,
		\rf_conf5_reg[4]/NET0131 ,
		_w1970_,
		_w1971_,
		_w2206_
	);
	LUT4 #(
		.INIT('h153f)
	) name306 (
		\rf_conf1_reg[4]/NET0131 ,
		\rf_conf2_reg[4]/NET0131 ,
		_w1976_,
		_w1977_,
		_w2207_
	);
	LUT4 #(
		.INIT('h8000)
	) name307 (
		_w2204_,
		_w2205_,
		_w2206_,
		_w2207_,
		_w2208_
	);
	LUT3 #(
		.INIT('h2a)
	) name308 (
		_w2098_,
		_w2203_,
		_w2208_,
		_w2209_
	);
	LUT4 #(
		.INIT('h135f)
	) name309 (
		\rf_conf6_reg[5]/NET0131 ,
		\rf_conf7_reg[5]/NET0131 ,
		_w1983_,
		_w1984_,
		_w2210_
	);
	LUT4 #(
		.INIT('h153f)
	) name310 (
		\rf_conf11_reg[5]/NET0131 ,
		\rf_conf8_reg[5]/NET0131 ,
		_w1986_,
		_w1987_,
		_w2211_
	);
	LUT4 #(
		.INIT('h135f)
	) name311 (
		\rf_conf13_reg[5]/NET0131 ,
		\rf_conf15_reg[5]/NET0131 ,
		_w1992_,
		_w1993_,
		_w2212_
	);
	LUT4 #(
		.INIT('h153f)
	) name312 (
		\rf_conf10_reg[5]/NET0131 ,
		\rf_conf9_reg[5]/NET0131 ,
		_w1989_,
		_w1990_,
		_w2213_
	);
	LUT4 #(
		.INIT('h8000)
	) name313 (
		_w2210_,
		_w2211_,
		_w2212_,
		_w2213_,
		_w2214_
	);
	LUT4 #(
		.INIT('h135f)
	) name314 (
		\rf_conf0_reg[5]/NET0131 ,
		\rf_conf4_reg[5]/NET0131 ,
		_w1979_,
		_w1980_,
		_w2215_
	);
	LUT4 #(
		.INIT('h135f)
	) name315 (
		\rf_conf12_reg[5]/NET0131 ,
		\rf_conf14_reg[5]/NET0131 ,
		_w1973_,
		_w1974_,
		_w2216_
	);
	LUT4 #(
		.INIT('h153f)
	) name316 (
		\rf_conf3_reg[5]/NET0131 ,
		\rf_conf5_reg[5]/NET0131 ,
		_w1970_,
		_w1971_,
		_w2217_
	);
	LUT4 #(
		.INIT('h153f)
	) name317 (
		\rf_conf1_reg[5]/NET0131 ,
		\rf_conf2_reg[5]/NET0131 ,
		_w1976_,
		_w1977_,
		_w2218_
	);
	LUT4 #(
		.INIT('h8000)
	) name318 (
		_w2215_,
		_w2216_,
		_w2217_,
		_w2218_,
		_w2219_
	);
	LUT3 #(
		.INIT('h2a)
	) name319 (
		_w2098_,
		_w2214_,
		_w2219_,
		_w2220_
	);
	LUT4 #(
		.INIT('h135f)
	) name320 (
		\rf_conf11_reg[6]/NET0131 ,
		\rf_conf15_reg[6]/NET0131 ,
		_w1987_,
		_w1993_,
		_w2221_
	);
	LUT4 #(
		.INIT('h135f)
	) name321 (
		\rf_conf0_reg[6]/NET0131 ,
		\rf_conf4_reg[6]/NET0131 ,
		_w1979_,
		_w1980_,
		_w2222_
	);
	LUT4 #(
		.INIT('h135f)
	) name322 (
		\rf_conf6_reg[6]/NET0131 ,
		\rf_conf9_reg[6]/NET0131 ,
		_w1983_,
		_w1989_,
		_w2223_
	);
	LUT4 #(
		.INIT('h153f)
	) name323 (
		\rf_conf13_reg[6]/NET0131 ,
		\rf_conf8_reg[6]/NET0131 ,
		_w1986_,
		_w1992_,
		_w2224_
	);
	LUT4 #(
		.INIT('h8000)
	) name324 (
		_w2221_,
		_w2222_,
		_w2223_,
		_w2224_,
		_w2225_
	);
	LUT4 #(
		.INIT('h153f)
	) name325 (
		\rf_conf10_reg[6]/NET0131 ,
		\rf_conf7_reg[6]/NET0131 ,
		_w1984_,
		_w1990_,
		_w2226_
	);
	LUT4 #(
		.INIT('h153f)
	) name326 (
		\rf_conf1_reg[6]/NET0131 ,
		\rf_conf2_reg[6]/NET0131 ,
		_w1976_,
		_w1977_,
		_w2227_
	);
	LUT4 #(
		.INIT('h135f)
	) name327 (
		\rf_conf12_reg[6]/NET0131 ,
		\rf_conf14_reg[6]/NET0131 ,
		_w1973_,
		_w1974_,
		_w2228_
	);
	LUT4 #(
		.INIT('h153f)
	) name328 (
		\rf_conf3_reg[6]/NET0131 ,
		\rf_conf5_reg[6]/NET0131 ,
		_w1970_,
		_w1971_,
		_w2229_
	);
	LUT4 #(
		.INIT('h8000)
	) name329 (
		_w2226_,
		_w2227_,
		_w2228_,
		_w2229_,
		_w2230_
	);
	LUT3 #(
		.INIT('h2a)
	) name330 (
		_w2098_,
		_w2225_,
		_w2230_,
		_w2231_
	);
	LUT4 #(
		.INIT('h153f)
	) name331 (
		\rf_conf11_reg[7]/NET0131 ,
		\rf_conf8_reg[7]/NET0131 ,
		_w1986_,
		_w1987_,
		_w2232_
	);
	LUT4 #(
		.INIT('h135f)
	) name332 (
		\rf_conf13_reg[7]/NET0131 ,
		\rf_conf15_reg[7]/NET0131 ,
		_w1992_,
		_w1993_,
		_w2233_
	);
	LUT4 #(
		.INIT('h135f)
	) name333 (
		\rf_conf12_reg[7]/NET0131 ,
		\rf_conf14_reg[7]/NET0131 ,
		_w1973_,
		_w1974_,
		_w2234_
	);
	LUT4 #(
		.INIT('h153f)
	) name334 (
		\rf_conf3_reg[7]/NET0131 ,
		\rf_conf5_reg[7]/NET0131 ,
		_w1970_,
		_w1971_,
		_w2235_
	);
	LUT4 #(
		.INIT('h8000)
	) name335 (
		_w2232_,
		_w2233_,
		_w2234_,
		_w2235_,
		_w2236_
	);
	LUT4 #(
		.INIT('h153f)
	) name336 (
		\rf_conf1_reg[7]/NET0131 ,
		\rf_conf2_reg[7]/NET0131 ,
		_w1976_,
		_w1977_,
		_w2237_
	);
	LUT4 #(
		.INIT('h135f)
	) name337 (
		\rf_conf6_reg[7]/NET0131 ,
		\rf_conf7_reg[7]/NET0131 ,
		_w1983_,
		_w1984_,
		_w2238_
	);
	LUT4 #(
		.INIT('h153f)
	) name338 (
		\rf_conf10_reg[7]/NET0131 ,
		\rf_conf9_reg[7]/NET0131 ,
		_w1989_,
		_w1990_,
		_w2239_
	);
	LUT4 #(
		.INIT('h135f)
	) name339 (
		\rf_conf0_reg[7]/NET0131 ,
		\rf_conf4_reg[7]/NET0131 ,
		_w1979_,
		_w1980_,
		_w2240_
	);
	LUT4 #(
		.INIT('h8000)
	) name340 (
		_w2237_,
		_w2238_,
		_w2239_,
		_w2240_,
		_w2241_
	);
	LUT3 #(
		.INIT('h2a)
	) name341 (
		_w2098_,
		_w2236_,
		_w2241_,
		_w2242_
	);
	LUT4 #(
		.INIT('h135f)
	) name342 (
		\rf_conf12_reg[8]/NET0131 ,
		\rf_conf14_reg[8]/NET0131 ,
		_w1973_,
		_w1974_,
		_w2243_
	);
	LUT4 #(
		.INIT('h135f)
	) name343 (
		\rf_conf13_reg[8]/NET0131 ,
		\rf_conf15_reg[8]/NET0131 ,
		_w1992_,
		_w1993_,
		_w2244_
	);
	LUT4 #(
		.INIT('h153f)
	) name344 (
		\rf_conf11_reg[8]/NET0131 ,
		\rf_conf8_reg[8]/NET0131 ,
		_w1986_,
		_w1987_,
		_w2245_
	);
	LUT4 #(
		.INIT('h153f)
	) name345 (
		\rf_conf1_reg[8]/NET0131 ,
		\rf_conf2_reg[8]/NET0131 ,
		_w1976_,
		_w1977_,
		_w2246_
	);
	LUT4 #(
		.INIT('h8000)
	) name346 (
		_w2243_,
		_w2244_,
		_w2245_,
		_w2246_,
		_w2247_
	);
	LUT4 #(
		.INIT('h153f)
	) name347 (
		\rf_conf3_reg[8]/NET0131 ,
		\rf_conf5_reg[8]/NET0131 ,
		_w1970_,
		_w1971_,
		_w2248_
	);
	LUT4 #(
		.INIT('h153f)
	) name348 (
		\rf_conf10_reg[8]/NET0131 ,
		\rf_conf9_reg[8]/NET0131 ,
		_w1989_,
		_w1990_,
		_w2249_
	);
	LUT4 #(
		.INIT('h135f)
	) name349 (
		\rf_conf6_reg[8]/NET0131 ,
		\rf_conf7_reg[8]/NET0131 ,
		_w1983_,
		_w1984_,
		_w2250_
	);
	LUT4 #(
		.INIT('h135f)
	) name350 (
		\rf_conf0_reg[8]/NET0131 ,
		\rf_conf4_reg[8]/NET0131 ,
		_w1979_,
		_w1980_,
		_w2251_
	);
	LUT4 #(
		.INIT('h8000)
	) name351 (
		_w2248_,
		_w2249_,
		_w2250_,
		_w2251_,
		_w2252_
	);
	LUT3 #(
		.INIT('h2a)
	) name352 (
		_w2098_,
		_w2247_,
		_w2252_,
		_w2253_
	);
	LUT4 #(
		.INIT('h135f)
	) name353 (
		\rf_conf6_reg[9]/NET0131 ,
		\rf_conf7_reg[9]/NET0131 ,
		_w1983_,
		_w1984_,
		_w2254_
	);
	LUT4 #(
		.INIT('h135f)
	) name354 (
		\rf_conf12_reg[9]/NET0131 ,
		\rf_conf14_reg[9]/NET0131 ,
		_w1973_,
		_w1974_,
		_w2255_
	);
	LUT4 #(
		.INIT('h135f)
	) name355 (
		\rf_conf13_reg[9]/NET0131 ,
		\rf_conf15_reg[9]/NET0131 ,
		_w1992_,
		_w1993_,
		_w2256_
	);
	LUT4 #(
		.INIT('h153f)
	) name356 (
		\rf_conf10_reg[9]/NET0131 ,
		\rf_conf9_reg[9]/NET0131 ,
		_w1989_,
		_w1990_,
		_w2257_
	);
	LUT4 #(
		.INIT('h8000)
	) name357 (
		_w2254_,
		_w2255_,
		_w2256_,
		_w2257_,
		_w2258_
	);
	LUT4 #(
		.INIT('h135f)
	) name358 (
		\rf_conf0_reg[9]/NET0131 ,
		\rf_conf4_reg[9]/NET0131 ,
		_w1979_,
		_w1980_,
		_w2259_
	);
	LUT4 #(
		.INIT('h153f)
	) name359 (
		\rf_conf11_reg[9]/NET0131 ,
		\rf_conf8_reg[9]/NET0131 ,
		_w1986_,
		_w1987_,
		_w2260_
	);
	LUT4 #(
		.INIT('h153f)
	) name360 (
		\rf_conf3_reg[9]/NET0131 ,
		\rf_conf5_reg[9]/NET0131 ,
		_w1970_,
		_w1971_,
		_w2261_
	);
	LUT4 #(
		.INIT('h153f)
	) name361 (
		\rf_conf1_reg[9]/NET0131 ,
		\rf_conf2_reg[9]/NET0131 ,
		_w1976_,
		_w1977_,
		_w2262_
	);
	LUT4 #(
		.INIT('h8000)
	) name362 (
		_w2259_,
		_w2260_,
		_w2261_,
		_w2262_,
		_w2263_
	);
	LUT3 #(
		.INIT('h2a)
	) name363 (
		_w2098_,
		_w2258_,
		_w2263_,
		_w2264_
	);
	LUT3 #(
		.INIT('h02)
	) name364 (
		\m5_s11_cyc_o_reg/NET0131 ,
		\rf_conf11_reg[10]/NET0131 ,
		\rf_conf11_reg[11]/NET0131 ,
		_w2265_
	);
	LUT3 #(
		.INIT('h02)
	) name365 (
		\m4_s11_cyc_o_reg/NET0131 ,
		\rf_conf11_reg[8]/NET0131 ,
		\rf_conf11_reg[9]/NET0131 ,
		_w2266_
	);
	LUT2 #(
		.INIT('h1)
	) name366 (
		_w2265_,
		_w2266_,
		_w2267_
	);
	LUT3 #(
		.INIT('h02)
	) name367 (
		\m7_s11_cyc_o_reg/NET0131 ,
		\rf_conf11_reg[14]/NET0131 ,
		\rf_conf11_reg[15]/NET0131 ,
		_w2268_
	);
	LUT3 #(
		.INIT('h02)
	) name368 (
		\m6_s11_cyc_o_reg/NET0131 ,
		\rf_conf11_reg[12]/NET0131 ,
		\rf_conf11_reg[13]/NET0131 ,
		_w2269_
	);
	LUT3 #(
		.INIT('h02)
	) name369 (
		\m1_s11_cyc_o_reg/NET0131 ,
		\rf_conf11_reg[2]/NET0131 ,
		\rf_conf11_reg[3]/NET0131 ,
		_w2270_
	);
	LUT3 #(
		.INIT('h02)
	) name370 (
		\m0_s11_cyc_o_reg/NET0131 ,
		\rf_conf11_reg[0]/NET0131 ,
		\rf_conf11_reg[1]/NET0131 ,
		_w2271_
	);
	LUT4 #(
		.INIT('h1110)
	) name371 (
		_w2268_,
		_w2269_,
		_w2270_,
		_w2271_,
		_w2272_
	);
	LUT3 #(
		.INIT('h02)
	) name372 (
		\m3_s11_cyc_o_reg/NET0131 ,
		\rf_conf11_reg[6]/NET0131 ,
		\rf_conf11_reg[7]/NET0131 ,
		_w2273_
	);
	LUT4 #(
		.INIT('h00fd)
	) name373 (
		\m3_s11_cyc_o_reg/NET0131 ,
		\rf_conf11_reg[6]/NET0131 ,
		\rf_conf11_reg[7]/NET0131 ,
		\s11_msel_arb0_state_reg[2]/NET0131 ,
		_w2274_
	);
	LUT3 #(
		.INIT('hd0)
	) name374 (
		_w2267_,
		_w2272_,
		_w2274_,
		_w2275_
	);
	LUT4 #(
		.INIT('hfd00)
	) name375 (
		\m7_s11_cyc_o_reg/NET0131 ,
		\rf_conf11_reg[14]/NET0131 ,
		\rf_conf11_reg[15]/NET0131 ,
		\s11_msel_arb0_state_reg[2]/NET0131 ,
		_w2276_
	);
	LUT2 #(
		.INIT('h2)
	) name376 (
		\s11_msel_arb0_state_reg[1]/NET0131 ,
		_w2276_,
		_w2277_
	);
	LUT3 #(
		.INIT('h02)
	) name377 (
		\m2_s11_cyc_o_reg/NET0131 ,
		\rf_conf11_reg[4]/NET0131 ,
		\rf_conf11_reg[5]/NET0131 ,
		_w2278_
	);
	LUT4 #(
		.INIT('h000e)
	) name378 (
		_w2265_,
		_w2266_,
		_w2273_,
		_w2278_,
		_w2279_
	);
	LUT3 #(
		.INIT('h02)
	) name379 (
		\s11_msel_arb0_state_reg[1]/NET0131 ,
		_w2270_,
		_w2271_,
		_w2280_
	);
	LUT3 #(
		.INIT('h45)
	) name380 (
		_w2277_,
		_w2279_,
		_w2280_,
		_w2281_
	);
	LUT3 #(
		.INIT('h02)
	) name381 (
		\s11_msel_arb0_state_reg[0]/NET0131 ,
		_w2275_,
		_w2281_,
		_w2282_
	);
	LUT4 #(
		.INIT('h2220)
	) name382 (
		\s11_msel_arb0_state_reg[2]/NET0131 ,
		_w2265_,
		_w2268_,
		_w2269_,
		_w2283_
	);
	LUT3 #(
		.INIT('h54)
	) name383 (
		_w2266_,
		_w2268_,
		_w2269_,
		_w2284_
	);
	LUT3 #(
		.INIT('h54)
	) name384 (
		_w2271_,
		_w2273_,
		_w2278_,
		_w2285_
	);
	LUT2 #(
		.INIT('h1)
	) name385 (
		_w2265_,
		_w2270_,
		_w2286_
	);
	LUT4 #(
		.INIT('h0155)
	) name386 (
		_w2283_,
		_w2284_,
		_w2285_,
		_w2286_,
		_w2287_
	);
	LUT4 #(
		.INIT('h00fd)
	) name387 (
		\m1_s11_cyc_o_reg/NET0131 ,
		\rf_conf11_reg[2]/NET0131 ,
		\rf_conf11_reg[3]/NET0131 ,
		\s11_msel_arb0_state_reg[2]/NET0131 ,
		_w2288_
	);
	LUT3 #(
		.INIT('he0)
	) name388 (
		_w2273_,
		_w2278_,
		_w2288_,
		_w2289_
	);
	LUT2 #(
		.INIT('h2)
	) name389 (
		\s11_msel_arb0_state_reg[0]/NET0131 ,
		\s11_msel_arb0_state_reg[1]/NET0131 ,
		_w2290_
	);
	LUT3 #(
		.INIT('hd0)
	) name390 (
		_w2287_,
		_w2289_,
		_w2290_,
		_w2291_
	);
	LUT2 #(
		.INIT('h1)
	) name391 (
		\s11_msel_arb0_state_reg[1]/NET0131 ,
		\s11_msel_arb0_state_reg[2]/NET0131 ,
		_w2292_
	);
	LUT3 #(
		.INIT('he0)
	) name392 (
		_w2270_,
		_w2271_,
		_w2292_,
		_w2293_
	);
	LUT3 #(
		.INIT('h0b)
	) name393 (
		\s11_msel_arb0_state_reg[2]/NET0131 ,
		_w2279_,
		_w2293_,
		_w2294_
	);
	LUT2 #(
		.INIT('h4)
	) name394 (
		\s11_msel_arb0_state_reg[1]/NET0131 ,
		\s11_msel_arb0_state_reg[2]/NET0131 ,
		_w2295_
	);
	LUT3 #(
		.INIT('he0)
	) name395 (
		_w2265_,
		_w2266_,
		_w2295_,
		_w2296_
	);
	LUT3 #(
		.INIT('h07)
	) name396 (
		\s11_msel_arb0_state_reg[2]/NET0131 ,
		_w2272_,
		_w2296_,
		_w2297_
	);
	LUT4 #(
		.INIT('h0001)
	) name397 (
		_w2268_,
		_w2269_,
		_w2273_,
		_w2278_,
		_w2298_
	);
	LUT4 #(
		.INIT('hbfaa)
	) name398 (
		\s11_msel_arb0_state_reg[0]/NET0131 ,
		_w2267_,
		_w2280_,
		_w2298_,
		_w2299_
	);
	LUT3 #(
		.INIT('h08)
	) name399 (
		_w2294_,
		_w2297_,
		_w2299_,
		_w2300_
	);
	LUT3 #(
		.INIT('hfe)
	) name400 (
		_w2282_,
		_w2291_,
		_w2300_,
		_w2301_
	);
	LUT3 #(
		.INIT('h02)
	) name401 (
		\m5_s12_cyc_o_reg/NET0131 ,
		\rf_conf12_reg[10]/NET0131 ,
		\rf_conf12_reg[11]/NET0131 ,
		_w2302_
	);
	LUT3 #(
		.INIT('h02)
	) name402 (
		\m4_s12_cyc_o_reg/NET0131 ,
		\rf_conf12_reg[8]/NET0131 ,
		\rf_conf12_reg[9]/NET0131 ,
		_w2303_
	);
	LUT2 #(
		.INIT('h1)
	) name403 (
		_w2302_,
		_w2303_,
		_w2304_
	);
	LUT3 #(
		.INIT('h02)
	) name404 (
		\m7_s12_cyc_o_reg/NET0131 ,
		\rf_conf12_reg[14]/NET0131 ,
		\rf_conf12_reg[15]/NET0131 ,
		_w2305_
	);
	LUT3 #(
		.INIT('h02)
	) name405 (
		\m6_s12_cyc_o_reg/NET0131 ,
		\rf_conf12_reg[12]/NET0131 ,
		\rf_conf12_reg[13]/NET0131 ,
		_w2306_
	);
	LUT3 #(
		.INIT('h02)
	) name406 (
		\m1_s12_cyc_o_reg/NET0131 ,
		\rf_conf12_reg[2]/NET0131 ,
		\rf_conf12_reg[3]/NET0131 ,
		_w2307_
	);
	LUT3 #(
		.INIT('h02)
	) name407 (
		\m0_s12_cyc_o_reg/NET0131 ,
		\rf_conf12_reg[0]/NET0131 ,
		\rf_conf12_reg[1]/NET0131 ,
		_w2308_
	);
	LUT4 #(
		.INIT('h1110)
	) name408 (
		_w2305_,
		_w2306_,
		_w2307_,
		_w2308_,
		_w2309_
	);
	LUT3 #(
		.INIT('h02)
	) name409 (
		\m3_s12_cyc_o_reg/NET0131 ,
		\rf_conf12_reg[6]/NET0131 ,
		\rf_conf12_reg[7]/NET0131 ,
		_w2310_
	);
	LUT4 #(
		.INIT('h00fd)
	) name410 (
		\m3_s12_cyc_o_reg/NET0131 ,
		\rf_conf12_reg[6]/NET0131 ,
		\rf_conf12_reg[7]/NET0131 ,
		\s12_msel_arb0_state_reg[2]/NET0131 ,
		_w2311_
	);
	LUT3 #(
		.INIT('hd0)
	) name411 (
		_w2304_,
		_w2309_,
		_w2311_,
		_w2312_
	);
	LUT4 #(
		.INIT('hfd00)
	) name412 (
		\m7_s12_cyc_o_reg/NET0131 ,
		\rf_conf12_reg[14]/NET0131 ,
		\rf_conf12_reg[15]/NET0131 ,
		\s12_msel_arb0_state_reg[2]/NET0131 ,
		_w2313_
	);
	LUT2 #(
		.INIT('h2)
	) name413 (
		\s12_msel_arb0_state_reg[1]/NET0131 ,
		_w2313_,
		_w2314_
	);
	LUT3 #(
		.INIT('h02)
	) name414 (
		\m2_s12_cyc_o_reg/NET0131 ,
		\rf_conf12_reg[4]/NET0131 ,
		\rf_conf12_reg[5]/NET0131 ,
		_w2315_
	);
	LUT4 #(
		.INIT('h000e)
	) name415 (
		_w2302_,
		_w2303_,
		_w2310_,
		_w2315_,
		_w2316_
	);
	LUT3 #(
		.INIT('h02)
	) name416 (
		\s12_msel_arb0_state_reg[1]/NET0131 ,
		_w2307_,
		_w2308_,
		_w2317_
	);
	LUT3 #(
		.INIT('h45)
	) name417 (
		_w2314_,
		_w2316_,
		_w2317_,
		_w2318_
	);
	LUT3 #(
		.INIT('h02)
	) name418 (
		\s12_msel_arb0_state_reg[0]/NET0131 ,
		_w2312_,
		_w2318_,
		_w2319_
	);
	LUT4 #(
		.INIT('h2220)
	) name419 (
		\s12_msel_arb0_state_reg[2]/NET0131 ,
		_w2302_,
		_w2305_,
		_w2306_,
		_w2320_
	);
	LUT3 #(
		.INIT('h54)
	) name420 (
		_w2303_,
		_w2305_,
		_w2306_,
		_w2321_
	);
	LUT3 #(
		.INIT('h54)
	) name421 (
		_w2308_,
		_w2310_,
		_w2315_,
		_w2322_
	);
	LUT2 #(
		.INIT('h1)
	) name422 (
		_w2302_,
		_w2307_,
		_w2323_
	);
	LUT4 #(
		.INIT('h0155)
	) name423 (
		_w2320_,
		_w2321_,
		_w2322_,
		_w2323_,
		_w2324_
	);
	LUT4 #(
		.INIT('h00fd)
	) name424 (
		\m1_s12_cyc_o_reg/NET0131 ,
		\rf_conf12_reg[2]/NET0131 ,
		\rf_conf12_reg[3]/NET0131 ,
		\s12_msel_arb0_state_reg[2]/NET0131 ,
		_w2325_
	);
	LUT3 #(
		.INIT('he0)
	) name425 (
		_w2310_,
		_w2315_,
		_w2325_,
		_w2326_
	);
	LUT2 #(
		.INIT('h2)
	) name426 (
		\s12_msel_arb0_state_reg[0]/NET0131 ,
		\s12_msel_arb0_state_reg[1]/NET0131 ,
		_w2327_
	);
	LUT3 #(
		.INIT('hd0)
	) name427 (
		_w2324_,
		_w2326_,
		_w2327_,
		_w2328_
	);
	LUT2 #(
		.INIT('h1)
	) name428 (
		\s12_msel_arb0_state_reg[1]/NET0131 ,
		\s12_msel_arb0_state_reg[2]/NET0131 ,
		_w2329_
	);
	LUT3 #(
		.INIT('he0)
	) name429 (
		_w2307_,
		_w2308_,
		_w2329_,
		_w2330_
	);
	LUT3 #(
		.INIT('h0b)
	) name430 (
		\s12_msel_arb0_state_reg[2]/NET0131 ,
		_w2316_,
		_w2330_,
		_w2331_
	);
	LUT2 #(
		.INIT('h4)
	) name431 (
		\s12_msel_arb0_state_reg[1]/NET0131 ,
		\s12_msel_arb0_state_reg[2]/NET0131 ,
		_w2332_
	);
	LUT3 #(
		.INIT('he0)
	) name432 (
		_w2302_,
		_w2303_,
		_w2332_,
		_w2333_
	);
	LUT3 #(
		.INIT('h07)
	) name433 (
		\s12_msel_arb0_state_reg[2]/NET0131 ,
		_w2309_,
		_w2333_,
		_w2334_
	);
	LUT4 #(
		.INIT('h0001)
	) name434 (
		_w2305_,
		_w2306_,
		_w2310_,
		_w2315_,
		_w2335_
	);
	LUT4 #(
		.INIT('hbfaa)
	) name435 (
		\s12_msel_arb0_state_reg[0]/NET0131 ,
		_w2304_,
		_w2317_,
		_w2335_,
		_w2336_
	);
	LUT3 #(
		.INIT('h08)
	) name436 (
		_w2331_,
		_w2334_,
		_w2336_,
		_w2337_
	);
	LUT3 #(
		.INIT('hfe)
	) name437 (
		_w2319_,
		_w2328_,
		_w2337_,
		_w2338_
	);
	LUT3 #(
		.INIT('h02)
	) name438 (
		\m5_s13_cyc_o_reg/NET0131 ,
		\rf_conf13_reg[10]/NET0131 ,
		\rf_conf13_reg[11]/NET0131 ,
		_w2339_
	);
	LUT3 #(
		.INIT('h02)
	) name439 (
		\m4_s13_cyc_o_reg/NET0131 ,
		\rf_conf13_reg[8]/NET0131 ,
		\rf_conf13_reg[9]/NET0131 ,
		_w2340_
	);
	LUT2 #(
		.INIT('h1)
	) name440 (
		_w2339_,
		_w2340_,
		_w2341_
	);
	LUT3 #(
		.INIT('h02)
	) name441 (
		\m7_s13_cyc_o_reg/NET0131 ,
		\rf_conf13_reg[14]/NET0131 ,
		\rf_conf13_reg[15]/NET0131 ,
		_w2342_
	);
	LUT3 #(
		.INIT('h02)
	) name442 (
		\m6_s13_cyc_o_reg/NET0131 ,
		\rf_conf13_reg[12]/NET0131 ,
		\rf_conf13_reg[13]/NET0131 ,
		_w2343_
	);
	LUT3 #(
		.INIT('h02)
	) name443 (
		\m1_s13_cyc_o_reg/NET0131 ,
		\rf_conf13_reg[2]/NET0131 ,
		\rf_conf13_reg[3]/NET0131 ,
		_w2344_
	);
	LUT3 #(
		.INIT('h02)
	) name444 (
		\m0_s13_cyc_o_reg/NET0131 ,
		\rf_conf13_reg[0]/NET0131 ,
		\rf_conf13_reg[1]/NET0131 ,
		_w2345_
	);
	LUT4 #(
		.INIT('h1110)
	) name445 (
		_w2342_,
		_w2343_,
		_w2344_,
		_w2345_,
		_w2346_
	);
	LUT3 #(
		.INIT('h02)
	) name446 (
		\m3_s13_cyc_o_reg/NET0131 ,
		\rf_conf13_reg[6]/NET0131 ,
		\rf_conf13_reg[7]/NET0131 ,
		_w2347_
	);
	LUT4 #(
		.INIT('h00fd)
	) name447 (
		\m3_s13_cyc_o_reg/NET0131 ,
		\rf_conf13_reg[6]/NET0131 ,
		\rf_conf13_reg[7]/NET0131 ,
		\s13_msel_arb0_state_reg[2]/NET0131 ,
		_w2348_
	);
	LUT3 #(
		.INIT('hd0)
	) name448 (
		_w2341_,
		_w2346_,
		_w2348_,
		_w2349_
	);
	LUT4 #(
		.INIT('hfd00)
	) name449 (
		\m7_s13_cyc_o_reg/NET0131 ,
		\rf_conf13_reg[14]/NET0131 ,
		\rf_conf13_reg[15]/NET0131 ,
		\s13_msel_arb0_state_reg[2]/NET0131 ,
		_w2350_
	);
	LUT2 #(
		.INIT('h2)
	) name450 (
		\s13_msel_arb0_state_reg[1]/NET0131 ,
		_w2350_,
		_w2351_
	);
	LUT3 #(
		.INIT('h02)
	) name451 (
		\m2_s13_cyc_o_reg/NET0131 ,
		\rf_conf13_reg[4]/NET0131 ,
		\rf_conf13_reg[5]/NET0131 ,
		_w2352_
	);
	LUT4 #(
		.INIT('h000e)
	) name452 (
		_w2339_,
		_w2340_,
		_w2347_,
		_w2352_,
		_w2353_
	);
	LUT3 #(
		.INIT('h02)
	) name453 (
		\s13_msel_arb0_state_reg[1]/NET0131 ,
		_w2344_,
		_w2345_,
		_w2354_
	);
	LUT3 #(
		.INIT('h45)
	) name454 (
		_w2351_,
		_w2353_,
		_w2354_,
		_w2355_
	);
	LUT3 #(
		.INIT('h02)
	) name455 (
		\s13_msel_arb0_state_reg[0]/NET0131 ,
		_w2349_,
		_w2355_,
		_w2356_
	);
	LUT4 #(
		.INIT('h2220)
	) name456 (
		\s13_msel_arb0_state_reg[2]/NET0131 ,
		_w2339_,
		_w2342_,
		_w2343_,
		_w2357_
	);
	LUT3 #(
		.INIT('h54)
	) name457 (
		_w2340_,
		_w2342_,
		_w2343_,
		_w2358_
	);
	LUT3 #(
		.INIT('h54)
	) name458 (
		_w2345_,
		_w2347_,
		_w2352_,
		_w2359_
	);
	LUT2 #(
		.INIT('h1)
	) name459 (
		_w2339_,
		_w2344_,
		_w2360_
	);
	LUT4 #(
		.INIT('h0155)
	) name460 (
		_w2357_,
		_w2358_,
		_w2359_,
		_w2360_,
		_w2361_
	);
	LUT4 #(
		.INIT('h00fd)
	) name461 (
		\m1_s13_cyc_o_reg/NET0131 ,
		\rf_conf13_reg[2]/NET0131 ,
		\rf_conf13_reg[3]/NET0131 ,
		\s13_msel_arb0_state_reg[2]/NET0131 ,
		_w2362_
	);
	LUT3 #(
		.INIT('he0)
	) name462 (
		_w2347_,
		_w2352_,
		_w2362_,
		_w2363_
	);
	LUT2 #(
		.INIT('h2)
	) name463 (
		\s13_msel_arb0_state_reg[0]/NET0131 ,
		\s13_msel_arb0_state_reg[1]/NET0131 ,
		_w2364_
	);
	LUT3 #(
		.INIT('hd0)
	) name464 (
		_w2361_,
		_w2363_,
		_w2364_,
		_w2365_
	);
	LUT2 #(
		.INIT('h1)
	) name465 (
		\s13_msel_arb0_state_reg[1]/NET0131 ,
		\s13_msel_arb0_state_reg[2]/NET0131 ,
		_w2366_
	);
	LUT3 #(
		.INIT('he0)
	) name466 (
		_w2344_,
		_w2345_,
		_w2366_,
		_w2367_
	);
	LUT3 #(
		.INIT('h0b)
	) name467 (
		\s13_msel_arb0_state_reg[2]/NET0131 ,
		_w2353_,
		_w2367_,
		_w2368_
	);
	LUT2 #(
		.INIT('h4)
	) name468 (
		\s13_msel_arb0_state_reg[1]/NET0131 ,
		\s13_msel_arb0_state_reg[2]/NET0131 ,
		_w2369_
	);
	LUT3 #(
		.INIT('he0)
	) name469 (
		_w2339_,
		_w2340_,
		_w2369_,
		_w2370_
	);
	LUT3 #(
		.INIT('h07)
	) name470 (
		\s13_msel_arb0_state_reg[2]/NET0131 ,
		_w2346_,
		_w2370_,
		_w2371_
	);
	LUT4 #(
		.INIT('h0001)
	) name471 (
		_w2342_,
		_w2343_,
		_w2347_,
		_w2352_,
		_w2372_
	);
	LUT4 #(
		.INIT('hbfaa)
	) name472 (
		\s13_msel_arb0_state_reg[0]/NET0131 ,
		_w2341_,
		_w2354_,
		_w2372_,
		_w2373_
	);
	LUT3 #(
		.INIT('h08)
	) name473 (
		_w2368_,
		_w2371_,
		_w2373_,
		_w2374_
	);
	LUT3 #(
		.INIT('hfe)
	) name474 (
		_w2356_,
		_w2365_,
		_w2374_,
		_w2375_
	);
	LUT3 #(
		.INIT('h02)
	) name475 (
		\m5_s14_cyc_o_reg/NET0131 ,
		\rf_conf14_reg[10]/NET0131 ,
		\rf_conf14_reg[11]/NET0131 ,
		_w2376_
	);
	LUT3 #(
		.INIT('h02)
	) name476 (
		\m4_s14_cyc_o_reg/NET0131 ,
		\rf_conf14_reg[8]/NET0131 ,
		\rf_conf14_reg[9]/NET0131 ,
		_w2377_
	);
	LUT2 #(
		.INIT('h1)
	) name477 (
		_w2376_,
		_w2377_,
		_w2378_
	);
	LUT3 #(
		.INIT('h02)
	) name478 (
		\m7_s14_cyc_o_reg/NET0131 ,
		\rf_conf14_reg[14]/NET0131 ,
		\rf_conf14_reg[15]/NET0131 ,
		_w2379_
	);
	LUT3 #(
		.INIT('h02)
	) name479 (
		\m6_s14_cyc_o_reg/NET0131 ,
		\rf_conf14_reg[12]/NET0131 ,
		\rf_conf14_reg[13]/NET0131 ,
		_w2380_
	);
	LUT3 #(
		.INIT('h02)
	) name480 (
		\m1_s14_cyc_o_reg/NET0131 ,
		\rf_conf14_reg[2]/NET0131 ,
		\rf_conf14_reg[3]/NET0131 ,
		_w2381_
	);
	LUT3 #(
		.INIT('h02)
	) name481 (
		\m0_s14_cyc_o_reg/NET0131 ,
		\rf_conf14_reg[0]/NET0131 ,
		\rf_conf14_reg[1]/NET0131 ,
		_w2382_
	);
	LUT4 #(
		.INIT('h1110)
	) name482 (
		_w2379_,
		_w2380_,
		_w2381_,
		_w2382_,
		_w2383_
	);
	LUT3 #(
		.INIT('h02)
	) name483 (
		\m3_s14_cyc_o_reg/NET0131 ,
		\rf_conf14_reg[6]/NET0131 ,
		\rf_conf14_reg[7]/NET0131 ,
		_w2384_
	);
	LUT4 #(
		.INIT('h00fd)
	) name484 (
		\m3_s14_cyc_o_reg/NET0131 ,
		\rf_conf14_reg[6]/NET0131 ,
		\rf_conf14_reg[7]/NET0131 ,
		\s14_msel_arb0_state_reg[2]/NET0131 ,
		_w2385_
	);
	LUT3 #(
		.INIT('hd0)
	) name485 (
		_w2378_,
		_w2383_,
		_w2385_,
		_w2386_
	);
	LUT4 #(
		.INIT('hfd00)
	) name486 (
		\m7_s14_cyc_o_reg/NET0131 ,
		\rf_conf14_reg[14]/NET0131 ,
		\rf_conf14_reg[15]/NET0131 ,
		\s14_msel_arb0_state_reg[2]/NET0131 ,
		_w2387_
	);
	LUT2 #(
		.INIT('h2)
	) name487 (
		\s14_msel_arb0_state_reg[1]/NET0131 ,
		_w2387_,
		_w2388_
	);
	LUT3 #(
		.INIT('h02)
	) name488 (
		\m2_s14_cyc_o_reg/NET0131 ,
		\rf_conf14_reg[4]/NET0131 ,
		\rf_conf14_reg[5]/NET0131 ,
		_w2389_
	);
	LUT4 #(
		.INIT('h000e)
	) name489 (
		_w2376_,
		_w2377_,
		_w2384_,
		_w2389_,
		_w2390_
	);
	LUT3 #(
		.INIT('h02)
	) name490 (
		\s14_msel_arb0_state_reg[1]/NET0131 ,
		_w2381_,
		_w2382_,
		_w2391_
	);
	LUT3 #(
		.INIT('h45)
	) name491 (
		_w2388_,
		_w2390_,
		_w2391_,
		_w2392_
	);
	LUT3 #(
		.INIT('h02)
	) name492 (
		\s14_msel_arb0_state_reg[0]/NET0131 ,
		_w2386_,
		_w2392_,
		_w2393_
	);
	LUT4 #(
		.INIT('h2220)
	) name493 (
		\s14_msel_arb0_state_reg[2]/NET0131 ,
		_w2376_,
		_w2379_,
		_w2380_,
		_w2394_
	);
	LUT3 #(
		.INIT('h54)
	) name494 (
		_w2377_,
		_w2379_,
		_w2380_,
		_w2395_
	);
	LUT3 #(
		.INIT('h54)
	) name495 (
		_w2382_,
		_w2384_,
		_w2389_,
		_w2396_
	);
	LUT2 #(
		.INIT('h1)
	) name496 (
		_w2376_,
		_w2381_,
		_w2397_
	);
	LUT4 #(
		.INIT('h0155)
	) name497 (
		_w2394_,
		_w2395_,
		_w2396_,
		_w2397_,
		_w2398_
	);
	LUT4 #(
		.INIT('h00fd)
	) name498 (
		\m1_s14_cyc_o_reg/NET0131 ,
		\rf_conf14_reg[2]/NET0131 ,
		\rf_conf14_reg[3]/NET0131 ,
		\s14_msel_arb0_state_reg[2]/NET0131 ,
		_w2399_
	);
	LUT3 #(
		.INIT('he0)
	) name499 (
		_w2384_,
		_w2389_,
		_w2399_,
		_w2400_
	);
	LUT2 #(
		.INIT('h2)
	) name500 (
		\s14_msel_arb0_state_reg[0]/NET0131 ,
		\s14_msel_arb0_state_reg[1]/NET0131 ,
		_w2401_
	);
	LUT3 #(
		.INIT('hd0)
	) name501 (
		_w2398_,
		_w2400_,
		_w2401_,
		_w2402_
	);
	LUT2 #(
		.INIT('h1)
	) name502 (
		\s14_msel_arb0_state_reg[1]/NET0131 ,
		\s14_msel_arb0_state_reg[2]/NET0131 ,
		_w2403_
	);
	LUT3 #(
		.INIT('he0)
	) name503 (
		_w2381_,
		_w2382_,
		_w2403_,
		_w2404_
	);
	LUT3 #(
		.INIT('h0b)
	) name504 (
		\s14_msel_arb0_state_reg[2]/NET0131 ,
		_w2390_,
		_w2404_,
		_w2405_
	);
	LUT2 #(
		.INIT('h4)
	) name505 (
		\s14_msel_arb0_state_reg[1]/NET0131 ,
		\s14_msel_arb0_state_reg[2]/NET0131 ,
		_w2406_
	);
	LUT3 #(
		.INIT('he0)
	) name506 (
		_w2376_,
		_w2377_,
		_w2406_,
		_w2407_
	);
	LUT3 #(
		.INIT('h07)
	) name507 (
		\s14_msel_arb0_state_reg[2]/NET0131 ,
		_w2383_,
		_w2407_,
		_w2408_
	);
	LUT4 #(
		.INIT('h0001)
	) name508 (
		_w2379_,
		_w2380_,
		_w2384_,
		_w2389_,
		_w2409_
	);
	LUT4 #(
		.INIT('hbfaa)
	) name509 (
		\s14_msel_arb0_state_reg[0]/NET0131 ,
		_w2378_,
		_w2391_,
		_w2409_,
		_w2410_
	);
	LUT3 #(
		.INIT('h08)
	) name510 (
		_w2405_,
		_w2408_,
		_w2410_,
		_w2411_
	);
	LUT3 #(
		.INIT('hfe)
	) name511 (
		_w2393_,
		_w2402_,
		_w2411_,
		_w2412_
	);
	LUT3 #(
		.INIT('h02)
	) name512 (
		\m5_s15_cyc_o_reg/NET0131 ,
		\rf_conf15_reg[10]/NET0131 ,
		\rf_conf15_reg[11]/NET0131 ,
		_w2413_
	);
	LUT3 #(
		.INIT('h02)
	) name513 (
		\m4_s15_cyc_o_reg/NET0131 ,
		\rf_conf15_reg[8]/NET0131 ,
		\rf_conf15_reg[9]/NET0131 ,
		_w2414_
	);
	LUT2 #(
		.INIT('h1)
	) name514 (
		_w2413_,
		_w2414_,
		_w2415_
	);
	LUT3 #(
		.INIT('h02)
	) name515 (
		\m6_s15_cyc_o_reg/NET0131 ,
		\rf_conf15_reg[12]/NET0131 ,
		\rf_conf15_reg[13]/NET0131 ,
		_w2416_
	);
	LUT3 #(
		.INIT('h02)
	) name516 (
		\m7_s15_cyc_o_reg/NET0131 ,
		\rf_conf15_reg[14]/NET0131 ,
		\rf_conf15_reg[15]/NET0131 ,
		_w2417_
	);
	LUT3 #(
		.INIT('h10)
	) name517 (
		\s15_msel_arb0_state_reg[0]/NET0131 ,
		\s15_msel_arb0_state_reg[1]/NET0131 ,
		\s15_msel_arb0_state_reg[2]/NET0131 ,
		_w2418_
	);
	LUT3 #(
		.INIT('he0)
	) name518 (
		_w2416_,
		_w2417_,
		_w2418_,
		_w2419_
	);
	LUT3 #(
		.INIT('h02)
	) name519 (
		\m3_s15_cyc_o_reg/NET0131 ,
		\rf_conf15_reg[6]/NET0131 ,
		\rf_conf15_reg[7]/NET0131 ,
		_w2420_
	);
	LUT3 #(
		.INIT('h02)
	) name520 (
		\m2_s15_cyc_o_reg/NET0131 ,
		\rf_conf15_reg[4]/NET0131 ,
		\rf_conf15_reg[5]/NET0131 ,
		_w2421_
	);
	LUT2 #(
		.INIT('h1)
	) name521 (
		_w2420_,
		_w2421_,
		_w2422_
	);
	LUT3 #(
		.INIT('h01)
	) name522 (
		\s15_msel_arb0_state_reg[1]/NET0131 ,
		_w2420_,
		_w2421_,
		_w2423_
	);
	LUT3 #(
		.INIT('h02)
	) name523 (
		\m1_s15_cyc_o_reg/NET0131 ,
		\rf_conf15_reg[2]/NET0131 ,
		\rf_conf15_reg[3]/NET0131 ,
		_w2424_
	);
	LUT3 #(
		.INIT('h02)
	) name524 (
		\m0_s15_cyc_o_reg/NET0131 ,
		\rf_conf15_reg[0]/NET0131 ,
		\rf_conf15_reg[1]/NET0131 ,
		_w2425_
	);
	LUT3 #(
		.INIT('h02)
	) name525 (
		_w2418_,
		_w2424_,
		_w2425_,
		_w2426_
	);
	LUT3 #(
		.INIT('h45)
	) name526 (
		_w2419_,
		_w2423_,
		_w2426_,
		_w2427_
	);
	LUT4 #(
		.INIT('h1110)
	) name527 (
		_w2416_,
		_w2417_,
		_w2424_,
		_w2425_,
		_w2428_
	);
	LUT2 #(
		.INIT('h8)
	) name528 (
		\s15_msel_arb0_state_reg[0]/NET0131 ,
		\s15_msel_arb0_state_reg[1]/NET0131 ,
		_w2429_
	);
	LUT3 #(
		.INIT('h08)
	) name529 (
		\s15_msel_arb0_state_reg[0]/NET0131 ,
		\s15_msel_arb0_state_reg[1]/NET0131 ,
		\s15_msel_arb0_state_reg[2]/NET0131 ,
		_w2430_
	);
	LUT2 #(
		.INIT('h4)
	) name530 (
		_w2420_,
		_w2430_,
		_w2431_
	);
	LUT2 #(
		.INIT('h4)
	) name531 (
		_w2428_,
		_w2431_,
		_w2432_
	);
	LUT3 #(
		.INIT('ha2)
	) name532 (
		_w2415_,
		_w2427_,
		_w2432_,
		_w2433_
	);
	LUT4 #(
		.INIT('h000e)
	) name533 (
		_w2413_,
		_w2414_,
		_w2420_,
		_w2421_,
		_w2434_
	);
	LUT4 #(
		.INIT('hfd00)
	) name534 (
		\m7_s15_cyc_o_reg/NET0131 ,
		\rf_conf15_reg[14]/NET0131 ,
		\rf_conf15_reg[15]/NET0131 ,
		\s15_msel_arb0_state_reg[1]/NET0131 ,
		_w2435_
	);
	LUT4 #(
		.INIT('h00fd)
	) name535 (
		\m5_s15_cyc_o_reg/NET0131 ,
		\rf_conf15_reg[10]/NET0131 ,
		\rf_conf15_reg[11]/NET0131 ,
		\s15_msel_arb0_state_reg[1]/NET0131 ,
		_w2436_
	);
	LUT3 #(
		.INIT('he0)
	) name536 (
		_w2420_,
		_w2421_,
		_w2436_,
		_w2437_
	);
	LUT2 #(
		.INIT('h8)
	) name537 (
		\s15_msel_arb0_state_reg[0]/NET0131 ,
		\s15_msel_arb0_state_reg[2]/NET0131 ,
		_w2438_
	);
	LUT3 #(
		.INIT('h10)
	) name538 (
		_w2424_,
		_w2425_,
		_w2438_,
		_w2439_
	);
	LUT4 #(
		.INIT('hf400)
	) name539 (
		_w2434_,
		_w2435_,
		_w2437_,
		_w2439_,
		_w2440_
	);
	LUT3 #(
		.INIT('h54)
	) name540 (
		\s15_msel_arb0_state_reg[2]/NET0131 ,
		_w2420_,
		_w2421_,
		_w2441_
	);
	LUT2 #(
		.INIT('h2)
	) name541 (
		_w2428_,
		_w2441_,
		_w2442_
	);
	LUT3 #(
		.INIT('ha8)
	) name542 (
		\s15_msel_arb0_state_reg[2]/NET0131 ,
		_w2416_,
		_w2417_,
		_w2443_
	);
	LUT2 #(
		.INIT('h4)
	) name543 (
		\s15_msel_arb0_state_reg[0]/NET0131 ,
		\s15_msel_arb0_state_reg[1]/NET0131 ,
		_w2444_
	);
	LUT3 #(
		.INIT('hd0)
	) name544 (
		_w2434_,
		_w2443_,
		_w2444_,
		_w2445_
	);
	LUT4 #(
		.INIT('h1110)
	) name545 (
		_w2413_,
		_w2414_,
		_w2416_,
		_w2417_,
		_w2446_
	);
	LUT2 #(
		.INIT('h2)
	) name546 (
		\s15_msel_arb0_state_reg[0]/NET0131 ,
		\s15_msel_arb0_state_reg[1]/NET0131 ,
		_w2447_
	);
	LUT3 #(
		.INIT('h02)
	) name547 (
		\s15_msel_arb0_state_reg[0]/NET0131 ,
		\s15_msel_arb0_state_reg[1]/NET0131 ,
		\s15_msel_arb0_state_reg[2]/NET0131 ,
		_w2448_
	);
	LUT3 #(
		.INIT('h01)
	) name548 (
		\s15_msel_arb0_state_reg[0]/NET0131 ,
		\s15_msel_arb0_state_reg[1]/NET0131 ,
		\s15_msel_arb0_state_reg[2]/NET0131 ,
		_w2449_
	);
	LUT4 #(
		.INIT('haeaf)
	) name549 (
		_w2424_,
		_w2425_,
		_w2448_,
		_w2449_,
		_w2450_
	);
	LUT3 #(
		.INIT('h0d)
	) name550 (
		_w2422_,
		_w2446_,
		_w2450_,
		_w2451_
	);
	LUT3 #(
		.INIT('h20)
	) name551 (
		\s15_msel_arb0_state_reg[0]/NET0131 ,
		\s15_msel_arb0_state_reg[1]/NET0131 ,
		\s15_msel_arb0_state_reg[2]/NET0131 ,
		_w2452_
	);
	LUT4 #(
		.INIT('h5400)
	) name552 (
		_w2413_,
		_w2416_,
		_w2417_,
		_w2452_,
		_w2453_
	);
	LUT3 #(
		.INIT('h80)
	) name553 (
		\s15_msel_arb0_state_reg[0]/NET0131 ,
		\s15_msel_arb0_state_reg[1]/NET0131 ,
		\s15_msel_arb0_state_reg[2]/NET0131 ,
		_w2454_
	);
	LUT4 #(
		.INIT('h27ff)
	) name554 (
		\s15_msel_arb0_state_reg[2]/NET0131 ,
		_w2417_,
		_w2420_,
		_w2429_,
		_w2455_
	);
	LUT2 #(
		.INIT('h4)
	) name555 (
		_w2453_,
		_w2455_,
		_w2456_
	);
	LUT4 #(
		.INIT('h0b00)
	) name556 (
		_w2442_,
		_w2445_,
		_w2451_,
		_w2456_,
		_w2457_
	);
	LUT3 #(
		.INIT('hef)
	) name557 (
		_w2433_,
		_w2440_,
		_w2457_,
		_w2458_
	);
	LUT3 #(
		.INIT('h02)
	) name558 (
		\m5_s3_cyc_o_reg/NET0131 ,
		\rf_conf3_reg[10]/NET0131 ,
		\rf_conf3_reg[11]/NET0131 ,
		_w2459_
	);
	LUT3 #(
		.INIT('h02)
	) name559 (
		\m4_s3_cyc_o_reg/NET0131 ,
		\rf_conf3_reg[8]/NET0131 ,
		\rf_conf3_reg[9]/NET0131 ,
		_w2460_
	);
	LUT2 #(
		.INIT('h1)
	) name560 (
		_w2459_,
		_w2460_,
		_w2461_
	);
	LUT3 #(
		.INIT('h02)
	) name561 (
		\m7_s3_cyc_o_reg/NET0131 ,
		\rf_conf3_reg[14]/NET0131 ,
		\rf_conf3_reg[15]/NET0131 ,
		_w2462_
	);
	LUT3 #(
		.INIT('h02)
	) name562 (
		\m6_s3_cyc_o_reg/NET0131 ,
		\rf_conf3_reg[12]/NET0131 ,
		\rf_conf3_reg[13]/NET0131 ,
		_w2463_
	);
	LUT3 #(
		.INIT('h02)
	) name563 (
		\m1_s3_cyc_o_reg/NET0131 ,
		\rf_conf3_reg[2]/NET0131 ,
		\rf_conf3_reg[3]/NET0131 ,
		_w2464_
	);
	LUT3 #(
		.INIT('h02)
	) name564 (
		\m0_s3_cyc_o_reg/NET0131 ,
		\rf_conf3_reg[0]/NET0131 ,
		\rf_conf3_reg[1]/NET0131 ,
		_w2465_
	);
	LUT4 #(
		.INIT('h1110)
	) name565 (
		_w2462_,
		_w2463_,
		_w2464_,
		_w2465_,
		_w2466_
	);
	LUT3 #(
		.INIT('h02)
	) name566 (
		\m3_s3_cyc_o_reg/NET0131 ,
		\rf_conf3_reg[6]/NET0131 ,
		\rf_conf3_reg[7]/NET0131 ,
		_w2467_
	);
	LUT4 #(
		.INIT('h00fd)
	) name567 (
		\m3_s3_cyc_o_reg/NET0131 ,
		\rf_conf3_reg[6]/NET0131 ,
		\rf_conf3_reg[7]/NET0131 ,
		\s3_msel_arb0_state_reg[2]/NET0131 ,
		_w2468_
	);
	LUT3 #(
		.INIT('hd0)
	) name568 (
		_w2461_,
		_w2466_,
		_w2468_,
		_w2469_
	);
	LUT4 #(
		.INIT('hfd00)
	) name569 (
		\m7_s3_cyc_o_reg/NET0131 ,
		\rf_conf3_reg[14]/NET0131 ,
		\rf_conf3_reg[15]/NET0131 ,
		\s3_msel_arb0_state_reg[2]/NET0131 ,
		_w2470_
	);
	LUT2 #(
		.INIT('h2)
	) name570 (
		\s3_msel_arb0_state_reg[1]/NET0131 ,
		_w2470_,
		_w2471_
	);
	LUT3 #(
		.INIT('h02)
	) name571 (
		\m2_s3_cyc_o_reg/NET0131 ,
		\rf_conf3_reg[4]/NET0131 ,
		\rf_conf3_reg[5]/NET0131 ,
		_w2472_
	);
	LUT4 #(
		.INIT('h000e)
	) name572 (
		_w2459_,
		_w2460_,
		_w2467_,
		_w2472_,
		_w2473_
	);
	LUT3 #(
		.INIT('h02)
	) name573 (
		\s3_msel_arb0_state_reg[1]/NET0131 ,
		_w2464_,
		_w2465_,
		_w2474_
	);
	LUT3 #(
		.INIT('h45)
	) name574 (
		_w2471_,
		_w2473_,
		_w2474_,
		_w2475_
	);
	LUT3 #(
		.INIT('h02)
	) name575 (
		\s3_msel_arb0_state_reg[0]/NET0131 ,
		_w2469_,
		_w2475_,
		_w2476_
	);
	LUT4 #(
		.INIT('h2220)
	) name576 (
		\s3_msel_arb0_state_reg[2]/NET0131 ,
		_w2459_,
		_w2462_,
		_w2463_,
		_w2477_
	);
	LUT3 #(
		.INIT('h54)
	) name577 (
		_w2460_,
		_w2462_,
		_w2463_,
		_w2478_
	);
	LUT3 #(
		.INIT('h54)
	) name578 (
		_w2465_,
		_w2467_,
		_w2472_,
		_w2479_
	);
	LUT2 #(
		.INIT('h1)
	) name579 (
		_w2459_,
		_w2464_,
		_w2480_
	);
	LUT4 #(
		.INIT('h0155)
	) name580 (
		_w2477_,
		_w2478_,
		_w2479_,
		_w2480_,
		_w2481_
	);
	LUT4 #(
		.INIT('h00fd)
	) name581 (
		\m1_s3_cyc_o_reg/NET0131 ,
		\rf_conf3_reg[2]/NET0131 ,
		\rf_conf3_reg[3]/NET0131 ,
		\s3_msel_arb0_state_reg[2]/NET0131 ,
		_w2482_
	);
	LUT3 #(
		.INIT('he0)
	) name582 (
		_w2467_,
		_w2472_,
		_w2482_,
		_w2483_
	);
	LUT2 #(
		.INIT('h2)
	) name583 (
		\s3_msel_arb0_state_reg[0]/NET0131 ,
		\s3_msel_arb0_state_reg[1]/NET0131 ,
		_w2484_
	);
	LUT3 #(
		.INIT('hd0)
	) name584 (
		_w2481_,
		_w2483_,
		_w2484_,
		_w2485_
	);
	LUT2 #(
		.INIT('h1)
	) name585 (
		\s3_msel_arb0_state_reg[1]/NET0131 ,
		\s3_msel_arb0_state_reg[2]/NET0131 ,
		_w2486_
	);
	LUT3 #(
		.INIT('he0)
	) name586 (
		_w2464_,
		_w2465_,
		_w2486_,
		_w2487_
	);
	LUT3 #(
		.INIT('h0b)
	) name587 (
		\s3_msel_arb0_state_reg[2]/NET0131 ,
		_w2473_,
		_w2487_,
		_w2488_
	);
	LUT2 #(
		.INIT('h4)
	) name588 (
		\s3_msel_arb0_state_reg[1]/NET0131 ,
		\s3_msel_arb0_state_reg[2]/NET0131 ,
		_w2489_
	);
	LUT3 #(
		.INIT('he0)
	) name589 (
		_w2459_,
		_w2460_,
		_w2489_,
		_w2490_
	);
	LUT3 #(
		.INIT('h07)
	) name590 (
		\s3_msel_arb0_state_reg[2]/NET0131 ,
		_w2466_,
		_w2490_,
		_w2491_
	);
	LUT4 #(
		.INIT('h0001)
	) name591 (
		_w2462_,
		_w2463_,
		_w2467_,
		_w2472_,
		_w2492_
	);
	LUT4 #(
		.INIT('hbfaa)
	) name592 (
		\s3_msel_arb0_state_reg[0]/NET0131 ,
		_w2461_,
		_w2474_,
		_w2492_,
		_w2493_
	);
	LUT3 #(
		.INIT('h08)
	) name593 (
		_w2488_,
		_w2491_,
		_w2493_,
		_w2494_
	);
	LUT3 #(
		.INIT('hfe)
	) name594 (
		_w2476_,
		_w2485_,
		_w2494_,
		_w2495_
	);
	LUT3 #(
		.INIT('h02)
	) name595 (
		\m5_s4_cyc_o_reg/NET0131 ,
		\rf_conf4_reg[10]/NET0131 ,
		\rf_conf4_reg[11]/NET0131 ,
		_w2496_
	);
	LUT3 #(
		.INIT('h02)
	) name596 (
		\m4_s4_cyc_o_reg/NET0131 ,
		\rf_conf4_reg[8]/NET0131 ,
		\rf_conf4_reg[9]/NET0131 ,
		_w2497_
	);
	LUT2 #(
		.INIT('h1)
	) name597 (
		_w2496_,
		_w2497_,
		_w2498_
	);
	LUT3 #(
		.INIT('h02)
	) name598 (
		\m7_s4_cyc_o_reg/NET0131 ,
		\rf_conf4_reg[14]/NET0131 ,
		\rf_conf4_reg[15]/NET0131 ,
		_w2499_
	);
	LUT3 #(
		.INIT('h02)
	) name599 (
		\m6_s4_cyc_o_reg/NET0131 ,
		\rf_conf4_reg[12]/NET0131 ,
		\rf_conf4_reg[13]/NET0131 ,
		_w2500_
	);
	LUT3 #(
		.INIT('h02)
	) name600 (
		\m1_s4_cyc_o_reg/NET0131 ,
		\rf_conf4_reg[2]/NET0131 ,
		\rf_conf4_reg[3]/NET0131 ,
		_w2501_
	);
	LUT3 #(
		.INIT('h02)
	) name601 (
		\m0_s4_cyc_o_reg/NET0131 ,
		\rf_conf4_reg[0]/NET0131 ,
		\rf_conf4_reg[1]/NET0131 ,
		_w2502_
	);
	LUT4 #(
		.INIT('h1110)
	) name602 (
		_w2499_,
		_w2500_,
		_w2501_,
		_w2502_,
		_w2503_
	);
	LUT3 #(
		.INIT('h02)
	) name603 (
		\m3_s4_cyc_o_reg/NET0131 ,
		\rf_conf4_reg[6]/NET0131 ,
		\rf_conf4_reg[7]/NET0131 ,
		_w2504_
	);
	LUT4 #(
		.INIT('h00fd)
	) name604 (
		\m3_s4_cyc_o_reg/NET0131 ,
		\rf_conf4_reg[6]/NET0131 ,
		\rf_conf4_reg[7]/NET0131 ,
		\s4_msel_arb0_state_reg[2]/NET0131 ,
		_w2505_
	);
	LUT3 #(
		.INIT('hd0)
	) name605 (
		_w2498_,
		_w2503_,
		_w2505_,
		_w2506_
	);
	LUT4 #(
		.INIT('hfd00)
	) name606 (
		\m7_s4_cyc_o_reg/NET0131 ,
		\rf_conf4_reg[14]/NET0131 ,
		\rf_conf4_reg[15]/NET0131 ,
		\s4_msel_arb0_state_reg[2]/NET0131 ,
		_w2507_
	);
	LUT2 #(
		.INIT('h2)
	) name607 (
		\s4_msel_arb0_state_reg[1]/NET0131 ,
		_w2507_,
		_w2508_
	);
	LUT3 #(
		.INIT('h02)
	) name608 (
		\m2_s4_cyc_o_reg/NET0131 ,
		\rf_conf4_reg[4]/NET0131 ,
		\rf_conf4_reg[5]/NET0131 ,
		_w2509_
	);
	LUT4 #(
		.INIT('h000e)
	) name609 (
		_w2496_,
		_w2497_,
		_w2504_,
		_w2509_,
		_w2510_
	);
	LUT3 #(
		.INIT('h02)
	) name610 (
		\s4_msel_arb0_state_reg[1]/NET0131 ,
		_w2501_,
		_w2502_,
		_w2511_
	);
	LUT3 #(
		.INIT('h45)
	) name611 (
		_w2508_,
		_w2510_,
		_w2511_,
		_w2512_
	);
	LUT3 #(
		.INIT('h02)
	) name612 (
		\s4_msel_arb0_state_reg[0]/NET0131 ,
		_w2506_,
		_w2512_,
		_w2513_
	);
	LUT4 #(
		.INIT('h2220)
	) name613 (
		\s4_msel_arb0_state_reg[2]/NET0131 ,
		_w2496_,
		_w2499_,
		_w2500_,
		_w2514_
	);
	LUT3 #(
		.INIT('h54)
	) name614 (
		_w2497_,
		_w2499_,
		_w2500_,
		_w2515_
	);
	LUT3 #(
		.INIT('h54)
	) name615 (
		_w2502_,
		_w2504_,
		_w2509_,
		_w2516_
	);
	LUT2 #(
		.INIT('h1)
	) name616 (
		_w2496_,
		_w2501_,
		_w2517_
	);
	LUT4 #(
		.INIT('h0155)
	) name617 (
		_w2514_,
		_w2515_,
		_w2516_,
		_w2517_,
		_w2518_
	);
	LUT4 #(
		.INIT('h00fd)
	) name618 (
		\m1_s4_cyc_o_reg/NET0131 ,
		\rf_conf4_reg[2]/NET0131 ,
		\rf_conf4_reg[3]/NET0131 ,
		\s4_msel_arb0_state_reg[2]/NET0131 ,
		_w2519_
	);
	LUT3 #(
		.INIT('he0)
	) name619 (
		_w2504_,
		_w2509_,
		_w2519_,
		_w2520_
	);
	LUT2 #(
		.INIT('h2)
	) name620 (
		\s4_msel_arb0_state_reg[0]/NET0131 ,
		\s4_msel_arb0_state_reg[1]/NET0131 ,
		_w2521_
	);
	LUT3 #(
		.INIT('hd0)
	) name621 (
		_w2518_,
		_w2520_,
		_w2521_,
		_w2522_
	);
	LUT2 #(
		.INIT('h1)
	) name622 (
		\s4_msel_arb0_state_reg[1]/NET0131 ,
		\s4_msel_arb0_state_reg[2]/NET0131 ,
		_w2523_
	);
	LUT3 #(
		.INIT('he0)
	) name623 (
		_w2501_,
		_w2502_,
		_w2523_,
		_w2524_
	);
	LUT3 #(
		.INIT('h0b)
	) name624 (
		\s4_msel_arb0_state_reg[2]/NET0131 ,
		_w2510_,
		_w2524_,
		_w2525_
	);
	LUT2 #(
		.INIT('h4)
	) name625 (
		\s4_msel_arb0_state_reg[1]/NET0131 ,
		\s4_msel_arb0_state_reg[2]/NET0131 ,
		_w2526_
	);
	LUT3 #(
		.INIT('he0)
	) name626 (
		_w2496_,
		_w2497_,
		_w2526_,
		_w2527_
	);
	LUT3 #(
		.INIT('h07)
	) name627 (
		\s4_msel_arb0_state_reg[2]/NET0131 ,
		_w2503_,
		_w2527_,
		_w2528_
	);
	LUT4 #(
		.INIT('h0001)
	) name628 (
		_w2499_,
		_w2500_,
		_w2504_,
		_w2509_,
		_w2529_
	);
	LUT4 #(
		.INIT('hbfaa)
	) name629 (
		\s4_msel_arb0_state_reg[0]/NET0131 ,
		_w2498_,
		_w2511_,
		_w2529_,
		_w2530_
	);
	LUT3 #(
		.INIT('h08)
	) name630 (
		_w2525_,
		_w2528_,
		_w2530_,
		_w2531_
	);
	LUT3 #(
		.INIT('hfe)
	) name631 (
		_w2513_,
		_w2522_,
		_w2531_,
		_w2532_
	);
	LUT3 #(
		.INIT('h02)
	) name632 (
		\m5_s5_cyc_o_reg/NET0131 ,
		\rf_conf5_reg[10]/NET0131 ,
		\rf_conf5_reg[11]/NET0131 ,
		_w2533_
	);
	LUT3 #(
		.INIT('h02)
	) name633 (
		\m4_s5_cyc_o_reg/NET0131 ,
		\rf_conf5_reg[8]/NET0131 ,
		\rf_conf5_reg[9]/NET0131 ,
		_w2534_
	);
	LUT2 #(
		.INIT('h1)
	) name634 (
		_w2533_,
		_w2534_,
		_w2535_
	);
	LUT3 #(
		.INIT('h02)
	) name635 (
		\m7_s5_cyc_o_reg/NET0131 ,
		\rf_conf5_reg[14]/NET0131 ,
		\rf_conf5_reg[15]/NET0131 ,
		_w2536_
	);
	LUT3 #(
		.INIT('h02)
	) name636 (
		\m6_s5_cyc_o_reg/NET0131 ,
		\rf_conf5_reg[12]/NET0131 ,
		\rf_conf5_reg[13]/NET0131 ,
		_w2537_
	);
	LUT3 #(
		.INIT('h02)
	) name637 (
		\m1_s5_cyc_o_reg/NET0131 ,
		\rf_conf5_reg[2]/NET0131 ,
		\rf_conf5_reg[3]/NET0131 ,
		_w2538_
	);
	LUT3 #(
		.INIT('h02)
	) name638 (
		\m0_s5_cyc_o_reg/NET0131 ,
		\rf_conf5_reg[0]/NET0131 ,
		\rf_conf5_reg[1]/NET0131 ,
		_w2539_
	);
	LUT4 #(
		.INIT('h1110)
	) name639 (
		_w2536_,
		_w2537_,
		_w2538_,
		_w2539_,
		_w2540_
	);
	LUT3 #(
		.INIT('h02)
	) name640 (
		\m3_s5_cyc_o_reg/NET0131 ,
		\rf_conf5_reg[6]/NET0131 ,
		\rf_conf5_reg[7]/NET0131 ,
		_w2541_
	);
	LUT4 #(
		.INIT('h00fd)
	) name641 (
		\m3_s5_cyc_o_reg/NET0131 ,
		\rf_conf5_reg[6]/NET0131 ,
		\rf_conf5_reg[7]/NET0131 ,
		\s5_msel_arb0_state_reg[2]/NET0131 ,
		_w2542_
	);
	LUT3 #(
		.INIT('hd0)
	) name642 (
		_w2535_,
		_w2540_,
		_w2542_,
		_w2543_
	);
	LUT4 #(
		.INIT('hfd00)
	) name643 (
		\m7_s5_cyc_o_reg/NET0131 ,
		\rf_conf5_reg[14]/NET0131 ,
		\rf_conf5_reg[15]/NET0131 ,
		\s5_msel_arb0_state_reg[2]/NET0131 ,
		_w2544_
	);
	LUT2 #(
		.INIT('h2)
	) name644 (
		\s5_msel_arb0_state_reg[1]/NET0131 ,
		_w2544_,
		_w2545_
	);
	LUT3 #(
		.INIT('h02)
	) name645 (
		\m2_s5_cyc_o_reg/NET0131 ,
		\rf_conf5_reg[4]/NET0131 ,
		\rf_conf5_reg[5]/NET0131 ,
		_w2546_
	);
	LUT4 #(
		.INIT('h000e)
	) name646 (
		_w2533_,
		_w2534_,
		_w2541_,
		_w2546_,
		_w2547_
	);
	LUT3 #(
		.INIT('h02)
	) name647 (
		\s5_msel_arb0_state_reg[1]/NET0131 ,
		_w2538_,
		_w2539_,
		_w2548_
	);
	LUT3 #(
		.INIT('h45)
	) name648 (
		_w2545_,
		_w2547_,
		_w2548_,
		_w2549_
	);
	LUT3 #(
		.INIT('h02)
	) name649 (
		\s5_msel_arb0_state_reg[0]/NET0131 ,
		_w2543_,
		_w2549_,
		_w2550_
	);
	LUT4 #(
		.INIT('h2220)
	) name650 (
		\s5_msel_arb0_state_reg[2]/NET0131 ,
		_w2533_,
		_w2536_,
		_w2537_,
		_w2551_
	);
	LUT3 #(
		.INIT('h54)
	) name651 (
		_w2534_,
		_w2536_,
		_w2537_,
		_w2552_
	);
	LUT3 #(
		.INIT('h54)
	) name652 (
		_w2539_,
		_w2541_,
		_w2546_,
		_w2553_
	);
	LUT2 #(
		.INIT('h1)
	) name653 (
		_w2533_,
		_w2538_,
		_w2554_
	);
	LUT4 #(
		.INIT('h0155)
	) name654 (
		_w2551_,
		_w2552_,
		_w2553_,
		_w2554_,
		_w2555_
	);
	LUT4 #(
		.INIT('h00fd)
	) name655 (
		\m1_s5_cyc_o_reg/NET0131 ,
		\rf_conf5_reg[2]/NET0131 ,
		\rf_conf5_reg[3]/NET0131 ,
		\s5_msel_arb0_state_reg[2]/NET0131 ,
		_w2556_
	);
	LUT3 #(
		.INIT('he0)
	) name656 (
		_w2541_,
		_w2546_,
		_w2556_,
		_w2557_
	);
	LUT2 #(
		.INIT('h2)
	) name657 (
		\s5_msel_arb0_state_reg[0]/NET0131 ,
		\s5_msel_arb0_state_reg[1]/NET0131 ,
		_w2558_
	);
	LUT3 #(
		.INIT('hd0)
	) name658 (
		_w2555_,
		_w2557_,
		_w2558_,
		_w2559_
	);
	LUT2 #(
		.INIT('h1)
	) name659 (
		\s5_msel_arb0_state_reg[1]/NET0131 ,
		\s5_msel_arb0_state_reg[2]/NET0131 ,
		_w2560_
	);
	LUT3 #(
		.INIT('he0)
	) name660 (
		_w2538_,
		_w2539_,
		_w2560_,
		_w2561_
	);
	LUT3 #(
		.INIT('h0b)
	) name661 (
		\s5_msel_arb0_state_reg[2]/NET0131 ,
		_w2547_,
		_w2561_,
		_w2562_
	);
	LUT2 #(
		.INIT('h4)
	) name662 (
		\s5_msel_arb0_state_reg[1]/NET0131 ,
		\s5_msel_arb0_state_reg[2]/NET0131 ,
		_w2563_
	);
	LUT3 #(
		.INIT('he0)
	) name663 (
		_w2533_,
		_w2534_,
		_w2563_,
		_w2564_
	);
	LUT3 #(
		.INIT('h07)
	) name664 (
		\s5_msel_arb0_state_reg[2]/NET0131 ,
		_w2540_,
		_w2564_,
		_w2565_
	);
	LUT4 #(
		.INIT('h0001)
	) name665 (
		_w2536_,
		_w2537_,
		_w2541_,
		_w2546_,
		_w2566_
	);
	LUT4 #(
		.INIT('hbfaa)
	) name666 (
		\s5_msel_arb0_state_reg[0]/NET0131 ,
		_w2535_,
		_w2548_,
		_w2566_,
		_w2567_
	);
	LUT3 #(
		.INIT('h08)
	) name667 (
		_w2562_,
		_w2565_,
		_w2567_,
		_w2568_
	);
	LUT3 #(
		.INIT('hfe)
	) name668 (
		_w2550_,
		_w2559_,
		_w2568_,
		_w2569_
	);
	LUT3 #(
		.INIT('h02)
	) name669 (
		\m5_s6_cyc_o_reg/NET0131 ,
		\rf_conf6_reg[10]/NET0131 ,
		\rf_conf6_reg[11]/NET0131 ,
		_w2570_
	);
	LUT3 #(
		.INIT('h02)
	) name670 (
		\m4_s6_cyc_o_reg/NET0131 ,
		\rf_conf6_reg[8]/NET0131 ,
		\rf_conf6_reg[9]/NET0131 ,
		_w2571_
	);
	LUT2 #(
		.INIT('h1)
	) name671 (
		_w2570_,
		_w2571_,
		_w2572_
	);
	LUT3 #(
		.INIT('h02)
	) name672 (
		\m7_s6_cyc_o_reg/NET0131 ,
		\rf_conf6_reg[14]/NET0131 ,
		\rf_conf6_reg[15]/NET0131 ,
		_w2573_
	);
	LUT3 #(
		.INIT('h02)
	) name673 (
		\m6_s6_cyc_o_reg/NET0131 ,
		\rf_conf6_reg[12]/NET0131 ,
		\rf_conf6_reg[13]/NET0131 ,
		_w2574_
	);
	LUT3 #(
		.INIT('h02)
	) name674 (
		\m1_s6_cyc_o_reg/NET0131 ,
		\rf_conf6_reg[2]/NET0131 ,
		\rf_conf6_reg[3]/NET0131 ,
		_w2575_
	);
	LUT3 #(
		.INIT('h02)
	) name675 (
		\m0_s6_cyc_o_reg/NET0131 ,
		\rf_conf6_reg[0]/NET0131 ,
		\rf_conf6_reg[1]/NET0131 ,
		_w2576_
	);
	LUT4 #(
		.INIT('h1110)
	) name676 (
		_w2573_,
		_w2574_,
		_w2575_,
		_w2576_,
		_w2577_
	);
	LUT3 #(
		.INIT('h02)
	) name677 (
		\m3_s6_cyc_o_reg/NET0131 ,
		\rf_conf6_reg[6]/NET0131 ,
		\rf_conf6_reg[7]/NET0131 ,
		_w2578_
	);
	LUT4 #(
		.INIT('h00fd)
	) name678 (
		\m3_s6_cyc_o_reg/NET0131 ,
		\rf_conf6_reg[6]/NET0131 ,
		\rf_conf6_reg[7]/NET0131 ,
		\s6_msel_arb0_state_reg[2]/NET0131 ,
		_w2579_
	);
	LUT3 #(
		.INIT('hd0)
	) name679 (
		_w2572_,
		_w2577_,
		_w2579_,
		_w2580_
	);
	LUT4 #(
		.INIT('hfd00)
	) name680 (
		\m7_s6_cyc_o_reg/NET0131 ,
		\rf_conf6_reg[14]/NET0131 ,
		\rf_conf6_reg[15]/NET0131 ,
		\s6_msel_arb0_state_reg[2]/NET0131 ,
		_w2581_
	);
	LUT2 #(
		.INIT('h2)
	) name681 (
		\s6_msel_arb0_state_reg[1]/NET0131 ,
		_w2581_,
		_w2582_
	);
	LUT3 #(
		.INIT('h02)
	) name682 (
		\m2_s6_cyc_o_reg/NET0131 ,
		\rf_conf6_reg[4]/NET0131 ,
		\rf_conf6_reg[5]/NET0131 ,
		_w2583_
	);
	LUT4 #(
		.INIT('h000e)
	) name683 (
		_w2570_,
		_w2571_,
		_w2578_,
		_w2583_,
		_w2584_
	);
	LUT3 #(
		.INIT('h02)
	) name684 (
		\s6_msel_arb0_state_reg[1]/NET0131 ,
		_w2575_,
		_w2576_,
		_w2585_
	);
	LUT3 #(
		.INIT('h45)
	) name685 (
		_w2582_,
		_w2584_,
		_w2585_,
		_w2586_
	);
	LUT3 #(
		.INIT('h02)
	) name686 (
		\s6_msel_arb0_state_reg[0]/NET0131 ,
		_w2580_,
		_w2586_,
		_w2587_
	);
	LUT4 #(
		.INIT('h2220)
	) name687 (
		\s6_msel_arb0_state_reg[2]/NET0131 ,
		_w2570_,
		_w2573_,
		_w2574_,
		_w2588_
	);
	LUT3 #(
		.INIT('h54)
	) name688 (
		_w2571_,
		_w2573_,
		_w2574_,
		_w2589_
	);
	LUT3 #(
		.INIT('h54)
	) name689 (
		_w2576_,
		_w2578_,
		_w2583_,
		_w2590_
	);
	LUT2 #(
		.INIT('h1)
	) name690 (
		_w2570_,
		_w2575_,
		_w2591_
	);
	LUT4 #(
		.INIT('h0155)
	) name691 (
		_w2588_,
		_w2589_,
		_w2590_,
		_w2591_,
		_w2592_
	);
	LUT4 #(
		.INIT('h00fd)
	) name692 (
		\m1_s6_cyc_o_reg/NET0131 ,
		\rf_conf6_reg[2]/NET0131 ,
		\rf_conf6_reg[3]/NET0131 ,
		\s6_msel_arb0_state_reg[2]/NET0131 ,
		_w2593_
	);
	LUT3 #(
		.INIT('he0)
	) name693 (
		_w2578_,
		_w2583_,
		_w2593_,
		_w2594_
	);
	LUT2 #(
		.INIT('h2)
	) name694 (
		\s6_msel_arb0_state_reg[0]/NET0131 ,
		\s6_msel_arb0_state_reg[1]/NET0131 ,
		_w2595_
	);
	LUT3 #(
		.INIT('hd0)
	) name695 (
		_w2592_,
		_w2594_,
		_w2595_,
		_w2596_
	);
	LUT2 #(
		.INIT('h1)
	) name696 (
		\s6_msel_arb0_state_reg[1]/NET0131 ,
		\s6_msel_arb0_state_reg[2]/NET0131 ,
		_w2597_
	);
	LUT3 #(
		.INIT('he0)
	) name697 (
		_w2575_,
		_w2576_,
		_w2597_,
		_w2598_
	);
	LUT3 #(
		.INIT('h0b)
	) name698 (
		\s6_msel_arb0_state_reg[2]/NET0131 ,
		_w2584_,
		_w2598_,
		_w2599_
	);
	LUT2 #(
		.INIT('h4)
	) name699 (
		\s6_msel_arb0_state_reg[1]/NET0131 ,
		\s6_msel_arb0_state_reg[2]/NET0131 ,
		_w2600_
	);
	LUT3 #(
		.INIT('he0)
	) name700 (
		_w2570_,
		_w2571_,
		_w2600_,
		_w2601_
	);
	LUT3 #(
		.INIT('h07)
	) name701 (
		\s6_msel_arb0_state_reg[2]/NET0131 ,
		_w2577_,
		_w2601_,
		_w2602_
	);
	LUT4 #(
		.INIT('h0001)
	) name702 (
		_w2573_,
		_w2574_,
		_w2578_,
		_w2583_,
		_w2603_
	);
	LUT4 #(
		.INIT('hbfaa)
	) name703 (
		\s6_msel_arb0_state_reg[0]/NET0131 ,
		_w2572_,
		_w2585_,
		_w2603_,
		_w2604_
	);
	LUT3 #(
		.INIT('h08)
	) name704 (
		_w2599_,
		_w2602_,
		_w2604_,
		_w2605_
	);
	LUT3 #(
		.INIT('hfe)
	) name705 (
		_w2587_,
		_w2596_,
		_w2605_,
		_w2606_
	);
	LUT3 #(
		.INIT('h02)
	) name706 (
		\m5_s8_cyc_o_reg/NET0131 ,
		\rf_conf8_reg[10]/NET0131 ,
		\rf_conf8_reg[11]/NET0131 ,
		_w2607_
	);
	LUT3 #(
		.INIT('h02)
	) name707 (
		\m4_s8_cyc_o_reg/NET0131 ,
		\rf_conf8_reg[8]/NET0131 ,
		\rf_conf8_reg[9]/NET0131 ,
		_w2608_
	);
	LUT2 #(
		.INIT('h1)
	) name708 (
		_w2607_,
		_w2608_,
		_w2609_
	);
	LUT3 #(
		.INIT('h02)
	) name709 (
		\m7_s8_cyc_o_reg/NET0131 ,
		\rf_conf8_reg[14]/NET0131 ,
		\rf_conf8_reg[15]/NET0131 ,
		_w2610_
	);
	LUT3 #(
		.INIT('h02)
	) name710 (
		\m6_s8_cyc_o_reg/NET0131 ,
		\rf_conf8_reg[12]/NET0131 ,
		\rf_conf8_reg[13]/NET0131 ,
		_w2611_
	);
	LUT3 #(
		.INIT('h02)
	) name711 (
		\m1_s8_cyc_o_reg/NET0131 ,
		\rf_conf8_reg[2]/NET0131 ,
		\rf_conf8_reg[3]/NET0131 ,
		_w2612_
	);
	LUT3 #(
		.INIT('h02)
	) name712 (
		\m0_s8_cyc_o_reg/NET0131 ,
		\rf_conf8_reg[0]/NET0131 ,
		\rf_conf8_reg[1]/NET0131 ,
		_w2613_
	);
	LUT4 #(
		.INIT('h1110)
	) name713 (
		_w2610_,
		_w2611_,
		_w2612_,
		_w2613_,
		_w2614_
	);
	LUT3 #(
		.INIT('h02)
	) name714 (
		\m3_s8_cyc_o_reg/NET0131 ,
		\rf_conf8_reg[6]/NET0131 ,
		\rf_conf8_reg[7]/NET0131 ,
		_w2615_
	);
	LUT4 #(
		.INIT('h00fd)
	) name715 (
		\m3_s8_cyc_o_reg/NET0131 ,
		\rf_conf8_reg[6]/NET0131 ,
		\rf_conf8_reg[7]/NET0131 ,
		\s8_msel_arb0_state_reg[2]/NET0131 ,
		_w2616_
	);
	LUT3 #(
		.INIT('hd0)
	) name716 (
		_w2609_,
		_w2614_,
		_w2616_,
		_w2617_
	);
	LUT4 #(
		.INIT('hfd00)
	) name717 (
		\m7_s8_cyc_o_reg/NET0131 ,
		\rf_conf8_reg[14]/NET0131 ,
		\rf_conf8_reg[15]/NET0131 ,
		\s8_msel_arb0_state_reg[2]/NET0131 ,
		_w2618_
	);
	LUT2 #(
		.INIT('h2)
	) name718 (
		\s8_msel_arb0_state_reg[1]/NET0131 ,
		_w2618_,
		_w2619_
	);
	LUT3 #(
		.INIT('h02)
	) name719 (
		\m2_s8_cyc_o_reg/NET0131 ,
		\rf_conf8_reg[4]/NET0131 ,
		\rf_conf8_reg[5]/NET0131 ,
		_w2620_
	);
	LUT4 #(
		.INIT('h000e)
	) name720 (
		_w2607_,
		_w2608_,
		_w2615_,
		_w2620_,
		_w2621_
	);
	LUT3 #(
		.INIT('h02)
	) name721 (
		\s8_msel_arb0_state_reg[1]/NET0131 ,
		_w2612_,
		_w2613_,
		_w2622_
	);
	LUT3 #(
		.INIT('h45)
	) name722 (
		_w2619_,
		_w2621_,
		_w2622_,
		_w2623_
	);
	LUT3 #(
		.INIT('h02)
	) name723 (
		\s8_msel_arb0_state_reg[0]/NET0131 ,
		_w2617_,
		_w2623_,
		_w2624_
	);
	LUT4 #(
		.INIT('h2220)
	) name724 (
		\s8_msel_arb0_state_reg[2]/NET0131 ,
		_w2607_,
		_w2610_,
		_w2611_,
		_w2625_
	);
	LUT3 #(
		.INIT('h54)
	) name725 (
		_w2608_,
		_w2610_,
		_w2611_,
		_w2626_
	);
	LUT3 #(
		.INIT('h54)
	) name726 (
		_w2613_,
		_w2615_,
		_w2620_,
		_w2627_
	);
	LUT2 #(
		.INIT('h1)
	) name727 (
		_w2607_,
		_w2612_,
		_w2628_
	);
	LUT4 #(
		.INIT('h0155)
	) name728 (
		_w2625_,
		_w2626_,
		_w2627_,
		_w2628_,
		_w2629_
	);
	LUT4 #(
		.INIT('h00fd)
	) name729 (
		\m1_s8_cyc_o_reg/NET0131 ,
		\rf_conf8_reg[2]/NET0131 ,
		\rf_conf8_reg[3]/NET0131 ,
		\s8_msel_arb0_state_reg[2]/NET0131 ,
		_w2630_
	);
	LUT3 #(
		.INIT('he0)
	) name730 (
		_w2615_,
		_w2620_,
		_w2630_,
		_w2631_
	);
	LUT2 #(
		.INIT('h2)
	) name731 (
		\s8_msel_arb0_state_reg[0]/NET0131 ,
		\s8_msel_arb0_state_reg[1]/NET0131 ,
		_w2632_
	);
	LUT3 #(
		.INIT('hd0)
	) name732 (
		_w2629_,
		_w2631_,
		_w2632_,
		_w2633_
	);
	LUT2 #(
		.INIT('h1)
	) name733 (
		\s8_msel_arb0_state_reg[1]/NET0131 ,
		\s8_msel_arb0_state_reg[2]/NET0131 ,
		_w2634_
	);
	LUT3 #(
		.INIT('he0)
	) name734 (
		_w2612_,
		_w2613_,
		_w2634_,
		_w2635_
	);
	LUT3 #(
		.INIT('h0b)
	) name735 (
		\s8_msel_arb0_state_reg[2]/NET0131 ,
		_w2621_,
		_w2635_,
		_w2636_
	);
	LUT2 #(
		.INIT('h4)
	) name736 (
		\s8_msel_arb0_state_reg[1]/NET0131 ,
		\s8_msel_arb0_state_reg[2]/NET0131 ,
		_w2637_
	);
	LUT3 #(
		.INIT('he0)
	) name737 (
		_w2607_,
		_w2608_,
		_w2637_,
		_w2638_
	);
	LUT3 #(
		.INIT('h07)
	) name738 (
		\s8_msel_arb0_state_reg[2]/NET0131 ,
		_w2614_,
		_w2638_,
		_w2639_
	);
	LUT4 #(
		.INIT('h0001)
	) name739 (
		_w2610_,
		_w2611_,
		_w2615_,
		_w2620_,
		_w2640_
	);
	LUT4 #(
		.INIT('hbfaa)
	) name740 (
		\s8_msel_arb0_state_reg[0]/NET0131 ,
		_w2609_,
		_w2622_,
		_w2640_,
		_w2641_
	);
	LUT3 #(
		.INIT('h08)
	) name741 (
		_w2636_,
		_w2639_,
		_w2641_,
		_w2642_
	);
	LUT3 #(
		.INIT('hfe)
	) name742 (
		_w2624_,
		_w2633_,
		_w2642_,
		_w2643_
	);
	LUT3 #(
		.INIT('h02)
	) name743 (
		\m3_s1_cyc_o_reg/NET0131 ,
		\rf_conf1_reg[6]/NET0131 ,
		\rf_conf1_reg[7]/NET0131 ,
		_w2644_
	);
	LUT3 #(
		.INIT('h02)
	) name744 (
		\m2_s1_cyc_o_reg/NET0131 ,
		\rf_conf1_reg[4]/NET0131 ,
		\rf_conf1_reg[5]/NET0131 ,
		_w2645_
	);
	LUT2 #(
		.INIT('h1)
	) name745 (
		_w2644_,
		_w2645_,
		_w2646_
	);
	LUT3 #(
		.INIT('h02)
	) name746 (
		\m4_s1_cyc_o_reg/NET0131 ,
		\rf_conf1_reg[8]/NET0131 ,
		\rf_conf1_reg[9]/NET0131 ,
		_w2647_
	);
	LUT3 #(
		.INIT('h02)
	) name747 (
		\m5_s1_cyc_o_reg/NET0131 ,
		\rf_conf1_reg[10]/NET0131 ,
		\rf_conf1_reg[11]/NET0131 ,
		_w2648_
	);
	LUT3 #(
		.INIT('h02)
	) name748 (
		\m7_s1_cyc_o_reg/NET0131 ,
		\rf_conf1_reg[14]/NET0131 ,
		\rf_conf1_reg[15]/NET0131 ,
		_w2649_
	);
	LUT3 #(
		.INIT('h02)
	) name749 (
		\m6_s1_cyc_o_reg/NET0131 ,
		\rf_conf1_reg[12]/NET0131 ,
		\rf_conf1_reg[13]/NET0131 ,
		_w2650_
	);
	LUT2 #(
		.INIT('h1)
	) name750 (
		_w2649_,
		_w2650_,
		_w2651_
	);
	LUT4 #(
		.INIT('h1110)
	) name751 (
		_w2647_,
		_w2648_,
		_w2649_,
		_w2650_,
		_w2652_
	);
	LUT3 #(
		.INIT('h02)
	) name752 (
		\m1_s1_cyc_o_reg/NET0131 ,
		\rf_conf1_reg[2]/NET0131 ,
		\rf_conf1_reg[3]/NET0131 ,
		_w2653_
	);
	LUT3 #(
		.INIT('h02)
	) name753 (
		\m0_s1_cyc_o_reg/NET0131 ,
		\rf_conf1_reg[0]/NET0131 ,
		\rf_conf1_reg[1]/NET0131 ,
		_w2654_
	);
	LUT2 #(
		.INIT('h1)
	) name754 (
		_w2653_,
		_w2654_,
		_w2655_
	);
	LUT4 #(
		.INIT('h2223)
	) name755 (
		\s1_msel_arb0_state_reg[1]/NET0131 ,
		\s1_msel_arb0_state_reg[2]/NET0131 ,
		_w2653_,
		_w2654_,
		_w2656_
	);
	LUT3 #(
		.INIT('hd0)
	) name756 (
		_w2646_,
		_w2652_,
		_w2656_,
		_w2657_
	);
	LUT4 #(
		.INIT('h8880)
	) name757 (
		\s1_msel_arb0_state_reg[1]/NET0131 ,
		\s1_msel_arb0_state_reg[2]/NET0131 ,
		_w2649_,
		_w2650_,
		_w2658_
	);
	LUT4 #(
		.INIT('h1110)
	) name758 (
		_w2644_,
		_w2645_,
		_w2647_,
		_w2648_,
		_w2659_
	);
	LUT3 #(
		.INIT('h02)
	) name759 (
		\s1_msel_arb0_state_reg[1]/NET0131 ,
		_w2653_,
		_w2654_,
		_w2660_
	);
	LUT3 #(
		.INIT('h45)
	) name760 (
		_w2658_,
		_w2659_,
		_w2660_,
		_w2661_
	);
	LUT3 #(
		.INIT('h45)
	) name761 (
		\s1_msel_arb0_state_reg[0]/NET0131 ,
		_w2657_,
		_w2661_,
		_w2662_
	);
	LUT4 #(
		.INIT('hfd00)
	) name762 (
		\m1_s1_cyc_o_reg/NET0131 ,
		\rf_conf1_reg[2]/NET0131 ,
		\rf_conf1_reg[3]/NET0131 ,
		\s1_msel_arb0_state_reg[0]/NET0131 ,
		_w2663_
	);
	LUT2 #(
		.INIT('h4)
	) name763 (
		\s1_msel_arb0_state_reg[2]/NET0131 ,
		_w2663_,
		_w2664_
	);
	LUT4 #(
		.INIT('h5100)
	) name764 (
		\s1_msel_arb0_state_reg[1]/NET0131 ,
		_w2646_,
		_w2652_,
		_w2664_,
		_w2665_
	);
	LUT2 #(
		.INIT('h4)
	) name765 (
		\s1_msel_arb0_state_reg[0]/NET0131 ,
		\s1_msel_arb0_state_reg[1]/NET0131 ,
		_w2666_
	);
	LUT3 #(
		.INIT('h01)
	) name766 (
		_w2644_,
		_w2645_,
		_w2666_,
		_w2667_
	);
	LUT4 #(
		.INIT('h0002)
	) name767 (
		\m4_s1_cyc_o_reg/NET0131 ,
		\rf_conf1_reg[8]/NET0131 ,
		\rf_conf1_reg[9]/NET0131 ,
		\s1_msel_arb0_state_reg[0]/NET0131 ,
		_w2668_
	);
	LUT4 #(
		.INIT('h0004)
	) name768 (
		\s1_msel_arb0_state_reg[1]/NET0131 ,
		\s1_msel_arb0_state_reg[2]/NET0131 ,
		_w2648_,
		_w2668_,
		_w2669_
	);
	LUT4 #(
		.INIT('h5d00)
	) name769 (
		_w2651_,
		_w2655_,
		_w2667_,
		_w2669_,
		_w2670_
	);
	LUT2 #(
		.INIT('h1)
	) name770 (
		_w2665_,
		_w2670_,
		_w2671_
	);
	LUT2 #(
		.INIT('h2)
	) name771 (
		\s1_msel_arb0_state_reg[1]/NET0131 ,
		\s1_msel_arb0_state_reg[2]/NET0131 ,
		_w2672_
	);
	LUT2 #(
		.INIT('h8)
	) name772 (
		_w2644_,
		_w2672_,
		_w2673_
	);
	LUT4 #(
		.INIT('h1110)
	) name773 (
		_w2649_,
		_w2650_,
		_w2653_,
		_w2654_,
		_w2674_
	);
	LUT3 #(
		.INIT('h10)
	) name774 (
		_w2647_,
		_w2648_,
		_w2672_,
		_w2675_
	);
	LUT3 #(
		.INIT('h45)
	) name775 (
		_w2673_,
		_w2674_,
		_w2675_,
		_w2676_
	);
	LUT2 #(
		.INIT('h8)
	) name776 (
		\s1_msel_arb0_state_reg[1]/NET0131 ,
		\s1_msel_arb0_state_reg[2]/NET0131 ,
		_w2677_
	);
	LUT2 #(
		.INIT('h8)
	) name777 (
		_w2649_,
		_w2677_,
		_w2678_
	);
	LUT3 #(
		.INIT('h10)
	) name778 (
		_w2653_,
		_w2654_,
		_w2677_,
		_w2679_
	);
	LUT3 #(
		.INIT('h23)
	) name779 (
		_w2659_,
		_w2678_,
		_w2679_,
		_w2680_
	);
	LUT3 #(
		.INIT('h2a)
	) name780 (
		\s1_msel_arb0_state_reg[0]/NET0131 ,
		_w2676_,
		_w2680_,
		_w2681_
	);
	LUT3 #(
		.INIT('hfb)
	) name781 (
		_w2662_,
		_w2671_,
		_w2681_,
		_w2682_
	);
	LUT3 #(
		.INIT('h02)
	) name782 (
		\m3_s2_cyc_o_reg/NET0131 ,
		\rf_conf2_reg[6]/NET0131 ,
		\rf_conf2_reg[7]/NET0131 ,
		_w2683_
	);
	LUT3 #(
		.INIT('h02)
	) name783 (
		\m2_s2_cyc_o_reg/NET0131 ,
		\rf_conf2_reg[4]/NET0131 ,
		\rf_conf2_reg[5]/NET0131 ,
		_w2684_
	);
	LUT2 #(
		.INIT('h1)
	) name784 (
		_w2683_,
		_w2684_,
		_w2685_
	);
	LUT3 #(
		.INIT('h02)
	) name785 (
		\m4_s2_cyc_o_reg/NET0131 ,
		\rf_conf2_reg[8]/NET0131 ,
		\rf_conf2_reg[9]/NET0131 ,
		_w2686_
	);
	LUT3 #(
		.INIT('h02)
	) name786 (
		\m5_s2_cyc_o_reg/NET0131 ,
		\rf_conf2_reg[10]/NET0131 ,
		\rf_conf2_reg[11]/NET0131 ,
		_w2687_
	);
	LUT3 #(
		.INIT('h02)
	) name787 (
		\m7_s2_cyc_o_reg/NET0131 ,
		\rf_conf2_reg[14]/NET0131 ,
		\rf_conf2_reg[15]/NET0131 ,
		_w2688_
	);
	LUT3 #(
		.INIT('h02)
	) name788 (
		\m6_s2_cyc_o_reg/NET0131 ,
		\rf_conf2_reg[12]/NET0131 ,
		\rf_conf2_reg[13]/NET0131 ,
		_w2689_
	);
	LUT2 #(
		.INIT('h1)
	) name789 (
		_w2688_,
		_w2689_,
		_w2690_
	);
	LUT4 #(
		.INIT('h1110)
	) name790 (
		_w2686_,
		_w2687_,
		_w2688_,
		_w2689_,
		_w2691_
	);
	LUT3 #(
		.INIT('h02)
	) name791 (
		\m1_s2_cyc_o_reg/NET0131 ,
		\rf_conf2_reg[2]/NET0131 ,
		\rf_conf2_reg[3]/NET0131 ,
		_w2692_
	);
	LUT3 #(
		.INIT('h02)
	) name792 (
		\m0_s2_cyc_o_reg/NET0131 ,
		\rf_conf2_reg[0]/NET0131 ,
		\rf_conf2_reg[1]/NET0131 ,
		_w2693_
	);
	LUT2 #(
		.INIT('h1)
	) name793 (
		_w2692_,
		_w2693_,
		_w2694_
	);
	LUT4 #(
		.INIT('h2223)
	) name794 (
		\s2_msel_arb0_state_reg[1]/NET0131 ,
		\s2_msel_arb0_state_reg[2]/NET0131 ,
		_w2692_,
		_w2693_,
		_w2695_
	);
	LUT3 #(
		.INIT('hd0)
	) name795 (
		_w2685_,
		_w2691_,
		_w2695_,
		_w2696_
	);
	LUT4 #(
		.INIT('h8880)
	) name796 (
		\s2_msel_arb0_state_reg[1]/NET0131 ,
		\s2_msel_arb0_state_reg[2]/NET0131 ,
		_w2688_,
		_w2689_,
		_w2697_
	);
	LUT4 #(
		.INIT('h1110)
	) name797 (
		_w2683_,
		_w2684_,
		_w2686_,
		_w2687_,
		_w2698_
	);
	LUT3 #(
		.INIT('h02)
	) name798 (
		\s2_msel_arb0_state_reg[1]/NET0131 ,
		_w2692_,
		_w2693_,
		_w2699_
	);
	LUT3 #(
		.INIT('h45)
	) name799 (
		_w2697_,
		_w2698_,
		_w2699_,
		_w2700_
	);
	LUT3 #(
		.INIT('h45)
	) name800 (
		\s2_msel_arb0_state_reg[0]/NET0131 ,
		_w2696_,
		_w2700_,
		_w2701_
	);
	LUT4 #(
		.INIT('hfd00)
	) name801 (
		\m1_s2_cyc_o_reg/NET0131 ,
		\rf_conf2_reg[2]/NET0131 ,
		\rf_conf2_reg[3]/NET0131 ,
		\s2_msel_arb0_state_reg[0]/NET0131 ,
		_w2702_
	);
	LUT2 #(
		.INIT('h4)
	) name802 (
		\s2_msel_arb0_state_reg[2]/NET0131 ,
		_w2702_,
		_w2703_
	);
	LUT4 #(
		.INIT('h5100)
	) name803 (
		\s2_msel_arb0_state_reg[1]/NET0131 ,
		_w2685_,
		_w2691_,
		_w2703_,
		_w2704_
	);
	LUT2 #(
		.INIT('h4)
	) name804 (
		\s2_msel_arb0_state_reg[0]/NET0131 ,
		\s2_msel_arb0_state_reg[1]/NET0131 ,
		_w2705_
	);
	LUT3 #(
		.INIT('h01)
	) name805 (
		_w2683_,
		_w2684_,
		_w2705_,
		_w2706_
	);
	LUT4 #(
		.INIT('h0002)
	) name806 (
		\m4_s2_cyc_o_reg/NET0131 ,
		\rf_conf2_reg[8]/NET0131 ,
		\rf_conf2_reg[9]/NET0131 ,
		\s2_msel_arb0_state_reg[0]/NET0131 ,
		_w2707_
	);
	LUT4 #(
		.INIT('h0004)
	) name807 (
		\s2_msel_arb0_state_reg[1]/NET0131 ,
		\s2_msel_arb0_state_reg[2]/NET0131 ,
		_w2687_,
		_w2707_,
		_w2708_
	);
	LUT4 #(
		.INIT('h5d00)
	) name808 (
		_w2690_,
		_w2694_,
		_w2706_,
		_w2708_,
		_w2709_
	);
	LUT2 #(
		.INIT('h1)
	) name809 (
		_w2704_,
		_w2709_,
		_w2710_
	);
	LUT2 #(
		.INIT('h2)
	) name810 (
		\s2_msel_arb0_state_reg[1]/NET0131 ,
		\s2_msel_arb0_state_reg[2]/NET0131 ,
		_w2711_
	);
	LUT2 #(
		.INIT('h8)
	) name811 (
		_w2683_,
		_w2711_,
		_w2712_
	);
	LUT4 #(
		.INIT('h1110)
	) name812 (
		_w2688_,
		_w2689_,
		_w2692_,
		_w2693_,
		_w2713_
	);
	LUT3 #(
		.INIT('h10)
	) name813 (
		_w2686_,
		_w2687_,
		_w2711_,
		_w2714_
	);
	LUT3 #(
		.INIT('h45)
	) name814 (
		_w2712_,
		_w2713_,
		_w2714_,
		_w2715_
	);
	LUT2 #(
		.INIT('h8)
	) name815 (
		\s2_msel_arb0_state_reg[1]/NET0131 ,
		\s2_msel_arb0_state_reg[2]/NET0131 ,
		_w2716_
	);
	LUT2 #(
		.INIT('h8)
	) name816 (
		_w2688_,
		_w2716_,
		_w2717_
	);
	LUT3 #(
		.INIT('h10)
	) name817 (
		_w2692_,
		_w2693_,
		_w2716_,
		_w2718_
	);
	LUT3 #(
		.INIT('h23)
	) name818 (
		_w2698_,
		_w2717_,
		_w2718_,
		_w2719_
	);
	LUT3 #(
		.INIT('h2a)
	) name819 (
		\s2_msel_arb0_state_reg[0]/NET0131 ,
		_w2715_,
		_w2719_,
		_w2720_
	);
	LUT3 #(
		.INIT('hfb)
	) name820 (
		_w2701_,
		_w2710_,
		_w2720_,
		_w2721_
	);
	LUT3 #(
		.INIT('h02)
	) name821 (
		\m3_s7_cyc_o_reg/NET0131 ,
		\rf_conf7_reg[6]/NET0131 ,
		\rf_conf7_reg[7]/NET0131 ,
		_w2722_
	);
	LUT3 #(
		.INIT('h02)
	) name822 (
		\m2_s7_cyc_o_reg/NET0131 ,
		\rf_conf7_reg[4]/NET0131 ,
		\rf_conf7_reg[5]/NET0131 ,
		_w2723_
	);
	LUT2 #(
		.INIT('h1)
	) name823 (
		_w2722_,
		_w2723_,
		_w2724_
	);
	LUT3 #(
		.INIT('h02)
	) name824 (
		\m4_s7_cyc_o_reg/NET0131 ,
		\rf_conf7_reg[8]/NET0131 ,
		\rf_conf7_reg[9]/NET0131 ,
		_w2725_
	);
	LUT3 #(
		.INIT('h02)
	) name825 (
		\m5_s7_cyc_o_reg/NET0131 ,
		\rf_conf7_reg[10]/NET0131 ,
		\rf_conf7_reg[11]/NET0131 ,
		_w2726_
	);
	LUT3 #(
		.INIT('h02)
	) name826 (
		\m7_s7_cyc_o_reg/NET0131 ,
		\rf_conf7_reg[14]/NET0131 ,
		\rf_conf7_reg[15]/NET0131 ,
		_w2727_
	);
	LUT3 #(
		.INIT('h02)
	) name827 (
		\m6_s7_cyc_o_reg/NET0131 ,
		\rf_conf7_reg[12]/NET0131 ,
		\rf_conf7_reg[13]/NET0131 ,
		_w2728_
	);
	LUT2 #(
		.INIT('h1)
	) name828 (
		_w2727_,
		_w2728_,
		_w2729_
	);
	LUT4 #(
		.INIT('h1110)
	) name829 (
		_w2725_,
		_w2726_,
		_w2727_,
		_w2728_,
		_w2730_
	);
	LUT3 #(
		.INIT('h02)
	) name830 (
		\m1_s7_cyc_o_reg/NET0131 ,
		\rf_conf7_reg[2]/NET0131 ,
		\rf_conf7_reg[3]/NET0131 ,
		_w2731_
	);
	LUT3 #(
		.INIT('h02)
	) name831 (
		\m0_s7_cyc_o_reg/NET0131 ,
		\rf_conf7_reg[0]/NET0131 ,
		\rf_conf7_reg[1]/NET0131 ,
		_w2732_
	);
	LUT2 #(
		.INIT('h1)
	) name832 (
		_w2731_,
		_w2732_,
		_w2733_
	);
	LUT4 #(
		.INIT('h2223)
	) name833 (
		\s7_msel_arb0_state_reg[1]/NET0131 ,
		\s7_msel_arb0_state_reg[2]/NET0131 ,
		_w2731_,
		_w2732_,
		_w2734_
	);
	LUT3 #(
		.INIT('hd0)
	) name834 (
		_w2724_,
		_w2730_,
		_w2734_,
		_w2735_
	);
	LUT4 #(
		.INIT('h8880)
	) name835 (
		\s7_msel_arb0_state_reg[1]/NET0131 ,
		\s7_msel_arb0_state_reg[2]/NET0131 ,
		_w2727_,
		_w2728_,
		_w2736_
	);
	LUT4 #(
		.INIT('h1110)
	) name836 (
		_w2722_,
		_w2723_,
		_w2725_,
		_w2726_,
		_w2737_
	);
	LUT3 #(
		.INIT('h02)
	) name837 (
		\s7_msel_arb0_state_reg[1]/NET0131 ,
		_w2731_,
		_w2732_,
		_w2738_
	);
	LUT3 #(
		.INIT('h45)
	) name838 (
		_w2736_,
		_w2737_,
		_w2738_,
		_w2739_
	);
	LUT3 #(
		.INIT('h45)
	) name839 (
		\s7_msel_arb0_state_reg[0]/NET0131 ,
		_w2735_,
		_w2739_,
		_w2740_
	);
	LUT4 #(
		.INIT('hfd00)
	) name840 (
		\m1_s7_cyc_o_reg/NET0131 ,
		\rf_conf7_reg[2]/NET0131 ,
		\rf_conf7_reg[3]/NET0131 ,
		\s7_msel_arb0_state_reg[0]/NET0131 ,
		_w2741_
	);
	LUT2 #(
		.INIT('h4)
	) name841 (
		\s7_msel_arb0_state_reg[2]/NET0131 ,
		_w2741_,
		_w2742_
	);
	LUT4 #(
		.INIT('h5100)
	) name842 (
		\s7_msel_arb0_state_reg[1]/NET0131 ,
		_w2724_,
		_w2730_,
		_w2742_,
		_w2743_
	);
	LUT2 #(
		.INIT('h4)
	) name843 (
		\s7_msel_arb0_state_reg[0]/NET0131 ,
		\s7_msel_arb0_state_reg[1]/NET0131 ,
		_w2744_
	);
	LUT3 #(
		.INIT('h01)
	) name844 (
		_w2722_,
		_w2723_,
		_w2744_,
		_w2745_
	);
	LUT4 #(
		.INIT('h0002)
	) name845 (
		\m4_s7_cyc_o_reg/NET0131 ,
		\rf_conf7_reg[8]/NET0131 ,
		\rf_conf7_reg[9]/NET0131 ,
		\s7_msel_arb0_state_reg[0]/NET0131 ,
		_w2746_
	);
	LUT4 #(
		.INIT('h0004)
	) name846 (
		\s7_msel_arb0_state_reg[1]/NET0131 ,
		\s7_msel_arb0_state_reg[2]/NET0131 ,
		_w2726_,
		_w2746_,
		_w2747_
	);
	LUT4 #(
		.INIT('h5d00)
	) name847 (
		_w2729_,
		_w2733_,
		_w2745_,
		_w2747_,
		_w2748_
	);
	LUT2 #(
		.INIT('h1)
	) name848 (
		_w2743_,
		_w2748_,
		_w2749_
	);
	LUT2 #(
		.INIT('h2)
	) name849 (
		\s7_msel_arb0_state_reg[1]/NET0131 ,
		\s7_msel_arb0_state_reg[2]/NET0131 ,
		_w2750_
	);
	LUT2 #(
		.INIT('h8)
	) name850 (
		_w2722_,
		_w2750_,
		_w2751_
	);
	LUT4 #(
		.INIT('h1110)
	) name851 (
		_w2727_,
		_w2728_,
		_w2731_,
		_w2732_,
		_w2752_
	);
	LUT3 #(
		.INIT('h10)
	) name852 (
		_w2725_,
		_w2726_,
		_w2750_,
		_w2753_
	);
	LUT3 #(
		.INIT('h45)
	) name853 (
		_w2751_,
		_w2752_,
		_w2753_,
		_w2754_
	);
	LUT2 #(
		.INIT('h8)
	) name854 (
		\s7_msel_arb0_state_reg[1]/NET0131 ,
		\s7_msel_arb0_state_reg[2]/NET0131 ,
		_w2755_
	);
	LUT2 #(
		.INIT('h8)
	) name855 (
		_w2727_,
		_w2755_,
		_w2756_
	);
	LUT3 #(
		.INIT('h10)
	) name856 (
		_w2731_,
		_w2732_,
		_w2755_,
		_w2757_
	);
	LUT3 #(
		.INIT('h23)
	) name857 (
		_w2737_,
		_w2756_,
		_w2757_,
		_w2758_
	);
	LUT3 #(
		.INIT('h2a)
	) name858 (
		\s7_msel_arb0_state_reg[0]/NET0131 ,
		_w2754_,
		_w2758_,
		_w2759_
	);
	LUT3 #(
		.INIT('hfb)
	) name859 (
		_w2740_,
		_w2749_,
		_w2759_,
		_w2760_
	);
	LUT3 #(
		.INIT('h02)
	) name860 (
		\m3_s9_cyc_o_reg/NET0131 ,
		\rf_conf9_reg[6]/NET0131 ,
		\rf_conf9_reg[7]/NET0131 ,
		_w2761_
	);
	LUT3 #(
		.INIT('h02)
	) name861 (
		\m2_s9_cyc_o_reg/NET0131 ,
		\rf_conf9_reg[4]/NET0131 ,
		\rf_conf9_reg[5]/NET0131 ,
		_w2762_
	);
	LUT2 #(
		.INIT('h1)
	) name862 (
		_w2761_,
		_w2762_,
		_w2763_
	);
	LUT3 #(
		.INIT('h02)
	) name863 (
		\m4_s9_cyc_o_reg/NET0131 ,
		\rf_conf9_reg[8]/NET0131 ,
		\rf_conf9_reg[9]/NET0131 ,
		_w2764_
	);
	LUT3 #(
		.INIT('h02)
	) name864 (
		\m5_s9_cyc_o_reg/NET0131 ,
		\rf_conf9_reg[10]/NET0131 ,
		\rf_conf9_reg[11]/NET0131 ,
		_w2765_
	);
	LUT3 #(
		.INIT('h02)
	) name865 (
		\m7_s9_cyc_o_reg/NET0131 ,
		\rf_conf9_reg[14]/NET0131 ,
		\rf_conf9_reg[15]/NET0131 ,
		_w2766_
	);
	LUT3 #(
		.INIT('h02)
	) name866 (
		\m6_s9_cyc_o_reg/NET0131 ,
		\rf_conf9_reg[12]/NET0131 ,
		\rf_conf9_reg[13]/NET0131 ,
		_w2767_
	);
	LUT2 #(
		.INIT('h1)
	) name867 (
		_w2766_,
		_w2767_,
		_w2768_
	);
	LUT4 #(
		.INIT('h1110)
	) name868 (
		_w2764_,
		_w2765_,
		_w2766_,
		_w2767_,
		_w2769_
	);
	LUT3 #(
		.INIT('h02)
	) name869 (
		\m1_s9_cyc_o_reg/NET0131 ,
		\rf_conf9_reg[2]/NET0131 ,
		\rf_conf9_reg[3]/NET0131 ,
		_w2770_
	);
	LUT3 #(
		.INIT('h02)
	) name870 (
		\m0_s9_cyc_o_reg/NET0131 ,
		\rf_conf9_reg[0]/NET0131 ,
		\rf_conf9_reg[1]/NET0131 ,
		_w2771_
	);
	LUT2 #(
		.INIT('h1)
	) name871 (
		_w2770_,
		_w2771_,
		_w2772_
	);
	LUT4 #(
		.INIT('h2223)
	) name872 (
		\s9_msel_arb0_state_reg[1]/NET0131 ,
		\s9_msel_arb0_state_reg[2]/NET0131 ,
		_w2770_,
		_w2771_,
		_w2773_
	);
	LUT3 #(
		.INIT('hd0)
	) name873 (
		_w2763_,
		_w2769_,
		_w2773_,
		_w2774_
	);
	LUT4 #(
		.INIT('h8880)
	) name874 (
		\s9_msel_arb0_state_reg[1]/NET0131 ,
		\s9_msel_arb0_state_reg[2]/NET0131 ,
		_w2766_,
		_w2767_,
		_w2775_
	);
	LUT4 #(
		.INIT('h1110)
	) name875 (
		_w2761_,
		_w2762_,
		_w2764_,
		_w2765_,
		_w2776_
	);
	LUT3 #(
		.INIT('h02)
	) name876 (
		\s9_msel_arb0_state_reg[1]/NET0131 ,
		_w2770_,
		_w2771_,
		_w2777_
	);
	LUT3 #(
		.INIT('h45)
	) name877 (
		_w2775_,
		_w2776_,
		_w2777_,
		_w2778_
	);
	LUT3 #(
		.INIT('h45)
	) name878 (
		\s9_msel_arb0_state_reg[0]/NET0131 ,
		_w2774_,
		_w2778_,
		_w2779_
	);
	LUT4 #(
		.INIT('hfd00)
	) name879 (
		\m1_s9_cyc_o_reg/NET0131 ,
		\rf_conf9_reg[2]/NET0131 ,
		\rf_conf9_reg[3]/NET0131 ,
		\s9_msel_arb0_state_reg[0]/NET0131 ,
		_w2780_
	);
	LUT2 #(
		.INIT('h4)
	) name880 (
		\s9_msel_arb0_state_reg[2]/NET0131 ,
		_w2780_,
		_w2781_
	);
	LUT4 #(
		.INIT('h5100)
	) name881 (
		\s9_msel_arb0_state_reg[1]/NET0131 ,
		_w2763_,
		_w2769_,
		_w2781_,
		_w2782_
	);
	LUT2 #(
		.INIT('h4)
	) name882 (
		\s9_msel_arb0_state_reg[0]/NET0131 ,
		\s9_msel_arb0_state_reg[1]/NET0131 ,
		_w2783_
	);
	LUT3 #(
		.INIT('h01)
	) name883 (
		_w2761_,
		_w2762_,
		_w2783_,
		_w2784_
	);
	LUT4 #(
		.INIT('h0002)
	) name884 (
		\m4_s9_cyc_o_reg/NET0131 ,
		\rf_conf9_reg[8]/NET0131 ,
		\rf_conf9_reg[9]/NET0131 ,
		\s9_msel_arb0_state_reg[0]/NET0131 ,
		_w2785_
	);
	LUT4 #(
		.INIT('h0004)
	) name885 (
		\s9_msel_arb0_state_reg[1]/NET0131 ,
		\s9_msel_arb0_state_reg[2]/NET0131 ,
		_w2765_,
		_w2785_,
		_w2786_
	);
	LUT4 #(
		.INIT('h5d00)
	) name886 (
		_w2768_,
		_w2772_,
		_w2784_,
		_w2786_,
		_w2787_
	);
	LUT2 #(
		.INIT('h1)
	) name887 (
		_w2782_,
		_w2787_,
		_w2788_
	);
	LUT2 #(
		.INIT('h2)
	) name888 (
		\s9_msel_arb0_state_reg[1]/NET0131 ,
		\s9_msel_arb0_state_reg[2]/NET0131 ,
		_w2789_
	);
	LUT2 #(
		.INIT('h8)
	) name889 (
		_w2761_,
		_w2789_,
		_w2790_
	);
	LUT4 #(
		.INIT('h1110)
	) name890 (
		_w2766_,
		_w2767_,
		_w2770_,
		_w2771_,
		_w2791_
	);
	LUT3 #(
		.INIT('h10)
	) name891 (
		_w2764_,
		_w2765_,
		_w2789_,
		_w2792_
	);
	LUT3 #(
		.INIT('h45)
	) name892 (
		_w2790_,
		_w2791_,
		_w2792_,
		_w2793_
	);
	LUT2 #(
		.INIT('h8)
	) name893 (
		\s9_msel_arb0_state_reg[1]/NET0131 ,
		\s9_msel_arb0_state_reg[2]/NET0131 ,
		_w2794_
	);
	LUT2 #(
		.INIT('h8)
	) name894 (
		_w2766_,
		_w2794_,
		_w2795_
	);
	LUT3 #(
		.INIT('h10)
	) name895 (
		_w2770_,
		_w2771_,
		_w2794_,
		_w2796_
	);
	LUT3 #(
		.INIT('h23)
	) name896 (
		_w2776_,
		_w2795_,
		_w2796_,
		_w2797_
	);
	LUT3 #(
		.INIT('h2a)
	) name897 (
		\s9_msel_arb0_state_reg[0]/NET0131 ,
		_w2793_,
		_w2797_,
		_w2798_
	);
	LUT3 #(
		.INIT('hfb)
	) name898 (
		_w2779_,
		_w2788_,
		_w2798_,
		_w2799_
	);
	LUT3 #(
		.INIT('h02)
	) name899 (
		\m3_s0_cyc_o_reg/NET0131 ,
		\rf_conf0_reg[6]/NET0131 ,
		\rf_conf0_reg[7]/NET0131 ,
		_w2800_
	);
	LUT3 #(
		.INIT('h02)
	) name900 (
		\m2_s0_cyc_o_reg/NET0131 ,
		\rf_conf0_reg[4]/NET0131 ,
		\rf_conf0_reg[5]/NET0131 ,
		_w2801_
	);
	LUT2 #(
		.INIT('h1)
	) name901 (
		_w2800_,
		_w2801_,
		_w2802_
	);
	LUT3 #(
		.INIT('h02)
	) name902 (
		\m4_s0_cyc_o_reg/NET0131 ,
		\rf_conf0_reg[8]/NET0131 ,
		\rf_conf0_reg[9]/NET0131 ,
		_w2803_
	);
	LUT3 #(
		.INIT('h02)
	) name903 (
		\m5_s0_cyc_o_reg/NET0131 ,
		\rf_conf0_reg[10]/NET0131 ,
		\rf_conf0_reg[11]/NET0131 ,
		_w2804_
	);
	LUT3 #(
		.INIT('h02)
	) name904 (
		\m7_s0_cyc_o_reg/NET0131 ,
		\rf_conf0_reg[14]/NET0131 ,
		\rf_conf0_reg[15]/NET0131 ,
		_w2805_
	);
	LUT3 #(
		.INIT('h02)
	) name905 (
		\m6_s0_cyc_o_reg/NET0131 ,
		\rf_conf0_reg[12]/NET0131 ,
		\rf_conf0_reg[13]/NET0131 ,
		_w2806_
	);
	LUT2 #(
		.INIT('h1)
	) name906 (
		_w2805_,
		_w2806_,
		_w2807_
	);
	LUT4 #(
		.INIT('h1110)
	) name907 (
		_w2803_,
		_w2804_,
		_w2805_,
		_w2806_,
		_w2808_
	);
	LUT3 #(
		.INIT('h02)
	) name908 (
		\m1_s0_cyc_o_reg/NET0131 ,
		\rf_conf0_reg[2]/NET0131 ,
		\rf_conf0_reg[3]/NET0131 ,
		_w2809_
	);
	LUT3 #(
		.INIT('h02)
	) name909 (
		\m0_s0_cyc_o_reg/NET0131 ,
		\rf_conf0_reg[0]/NET0131 ,
		\rf_conf0_reg[1]/NET0131 ,
		_w2810_
	);
	LUT2 #(
		.INIT('h1)
	) name910 (
		_w2809_,
		_w2810_,
		_w2811_
	);
	LUT4 #(
		.INIT('h2223)
	) name911 (
		\s0_msel_arb0_state_reg[1]/NET0131 ,
		\s0_msel_arb0_state_reg[2]/NET0131 ,
		_w2809_,
		_w2810_,
		_w2812_
	);
	LUT3 #(
		.INIT('hd0)
	) name912 (
		_w2802_,
		_w2808_,
		_w2812_,
		_w2813_
	);
	LUT4 #(
		.INIT('h8880)
	) name913 (
		\s0_msel_arb0_state_reg[1]/NET0131 ,
		\s0_msel_arb0_state_reg[2]/NET0131 ,
		_w2805_,
		_w2806_,
		_w2814_
	);
	LUT4 #(
		.INIT('h1110)
	) name914 (
		_w2800_,
		_w2801_,
		_w2803_,
		_w2804_,
		_w2815_
	);
	LUT3 #(
		.INIT('h02)
	) name915 (
		\s0_msel_arb0_state_reg[1]/NET0131 ,
		_w2809_,
		_w2810_,
		_w2816_
	);
	LUT3 #(
		.INIT('h45)
	) name916 (
		_w2814_,
		_w2815_,
		_w2816_,
		_w2817_
	);
	LUT3 #(
		.INIT('h45)
	) name917 (
		\s0_msel_arb0_state_reg[0]/NET0131 ,
		_w2813_,
		_w2817_,
		_w2818_
	);
	LUT4 #(
		.INIT('hfd00)
	) name918 (
		\m1_s0_cyc_o_reg/NET0131 ,
		\rf_conf0_reg[2]/NET0131 ,
		\rf_conf0_reg[3]/NET0131 ,
		\s0_msel_arb0_state_reg[0]/NET0131 ,
		_w2819_
	);
	LUT2 #(
		.INIT('h4)
	) name919 (
		\s0_msel_arb0_state_reg[2]/NET0131 ,
		_w2819_,
		_w2820_
	);
	LUT4 #(
		.INIT('h5100)
	) name920 (
		\s0_msel_arb0_state_reg[1]/NET0131 ,
		_w2802_,
		_w2808_,
		_w2820_,
		_w2821_
	);
	LUT2 #(
		.INIT('h4)
	) name921 (
		\s0_msel_arb0_state_reg[0]/NET0131 ,
		\s0_msel_arb0_state_reg[1]/NET0131 ,
		_w2822_
	);
	LUT3 #(
		.INIT('h01)
	) name922 (
		_w2800_,
		_w2801_,
		_w2822_,
		_w2823_
	);
	LUT4 #(
		.INIT('h0002)
	) name923 (
		\m4_s0_cyc_o_reg/NET0131 ,
		\rf_conf0_reg[8]/NET0131 ,
		\rf_conf0_reg[9]/NET0131 ,
		\s0_msel_arb0_state_reg[0]/NET0131 ,
		_w2824_
	);
	LUT4 #(
		.INIT('h0004)
	) name924 (
		\s0_msel_arb0_state_reg[1]/NET0131 ,
		\s0_msel_arb0_state_reg[2]/NET0131 ,
		_w2804_,
		_w2824_,
		_w2825_
	);
	LUT4 #(
		.INIT('h5d00)
	) name925 (
		_w2807_,
		_w2811_,
		_w2823_,
		_w2825_,
		_w2826_
	);
	LUT2 #(
		.INIT('h1)
	) name926 (
		_w2821_,
		_w2826_,
		_w2827_
	);
	LUT2 #(
		.INIT('h2)
	) name927 (
		\s0_msel_arb0_state_reg[1]/NET0131 ,
		\s0_msel_arb0_state_reg[2]/NET0131 ,
		_w2828_
	);
	LUT2 #(
		.INIT('h8)
	) name928 (
		_w2800_,
		_w2828_,
		_w2829_
	);
	LUT4 #(
		.INIT('h1110)
	) name929 (
		_w2805_,
		_w2806_,
		_w2809_,
		_w2810_,
		_w2830_
	);
	LUT3 #(
		.INIT('h10)
	) name930 (
		_w2803_,
		_w2804_,
		_w2828_,
		_w2831_
	);
	LUT3 #(
		.INIT('h45)
	) name931 (
		_w2829_,
		_w2830_,
		_w2831_,
		_w2832_
	);
	LUT2 #(
		.INIT('h8)
	) name932 (
		\s0_msel_arb0_state_reg[1]/NET0131 ,
		\s0_msel_arb0_state_reg[2]/NET0131 ,
		_w2833_
	);
	LUT2 #(
		.INIT('h8)
	) name933 (
		_w2805_,
		_w2833_,
		_w2834_
	);
	LUT3 #(
		.INIT('h10)
	) name934 (
		_w2809_,
		_w2810_,
		_w2833_,
		_w2835_
	);
	LUT3 #(
		.INIT('h23)
	) name935 (
		_w2815_,
		_w2834_,
		_w2835_,
		_w2836_
	);
	LUT3 #(
		.INIT('h2a)
	) name936 (
		\s0_msel_arb0_state_reg[0]/NET0131 ,
		_w2832_,
		_w2836_,
		_w2837_
	);
	LUT3 #(
		.INIT('hfb)
	) name937 (
		_w2818_,
		_w2827_,
		_w2837_,
		_w2838_
	);
	LUT3 #(
		.INIT('h02)
	) name938 (
		\m3_s10_cyc_o_reg/NET0131 ,
		\rf_conf10_reg[6]/NET0131 ,
		\rf_conf10_reg[7]/NET0131 ,
		_w2839_
	);
	LUT3 #(
		.INIT('h02)
	) name939 (
		\m2_s10_cyc_o_reg/NET0131 ,
		\rf_conf10_reg[4]/NET0131 ,
		\rf_conf10_reg[5]/NET0131 ,
		_w2840_
	);
	LUT2 #(
		.INIT('h1)
	) name940 (
		_w2839_,
		_w2840_,
		_w2841_
	);
	LUT3 #(
		.INIT('h02)
	) name941 (
		\m4_s10_cyc_o_reg/NET0131 ,
		\rf_conf10_reg[8]/NET0131 ,
		\rf_conf10_reg[9]/NET0131 ,
		_w2842_
	);
	LUT3 #(
		.INIT('h02)
	) name942 (
		\m5_s10_cyc_o_reg/NET0131 ,
		\rf_conf10_reg[10]/NET0131 ,
		\rf_conf10_reg[11]/NET0131 ,
		_w2843_
	);
	LUT3 #(
		.INIT('h02)
	) name943 (
		\m7_s10_cyc_o_reg/NET0131 ,
		\rf_conf10_reg[14]/NET0131 ,
		\rf_conf10_reg[15]/NET0131 ,
		_w2844_
	);
	LUT3 #(
		.INIT('h02)
	) name944 (
		\m6_s10_cyc_o_reg/NET0131 ,
		\rf_conf10_reg[12]/NET0131 ,
		\rf_conf10_reg[13]/NET0131 ,
		_w2845_
	);
	LUT2 #(
		.INIT('h1)
	) name945 (
		_w2844_,
		_w2845_,
		_w2846_
	);
	LUT4 #(
		.INIT('h1110)
	) name946 (
		_w2842_,
		_w2843_,
		_w2844_,
		_w2845_,
		_w2847_
	);
	LUT3 #(
		.INIT('h02)
	) name947 (
		\m1_s10_cyc_o_reg/NET0131 ,
		\rf_conf10_reg[2]/NET0131 ,
		\rf_conf10_reg[3]/NET0131 ,
		_w2848_
	);
	LUT3 #(
		.INIT('h02)
	) name948 (
		\m0_s10_cyc_o_reg/NET0131 ,
		\rf_conf10_reg[0]/NET0131 ,
		\rf_conf10_reg[1]/NET0131 ,
		_w2849_
	);
	LUT2 #(
		.INIT('h1)
	) name949 (
		_w2848_,
		_w2849_,
		_w2850_
	);
	LUT4 #(
		.INIT('h2223)
	) name950 (
		\s10_msel_arb0_state_reg[1]/NET0131 ,
		\s10_msel_arb0_state_reg[2]/NET0131 ,
		_w2848_,
		_w2849_,
		_w2851_
	);
	LUT3 #(
		.INIT('hd0)
	) name951 (
		_w2841_,
		_w2847_,
		_w2851_,
		_w2852_
	);
	LUT4 #(
		.INIT('h8880)
	) name952 (
		\s10_msel_arb0_state_reg[1]/NET0131 ,
		\s10_msel_arb0_state_reg[2]/NET0131 ,
		_w2844_,
		_w2845_,
		_w2853_
	);
	LUT4 #(
		.INIT('h1110)
	) name953 (
		_w2839_,
		_w2840_,
		_w2842_,
		_w2843_,
		_w2854_
	);
	LUT3 #(
		.INIT('h02)
	) name954 (
		\s10_msel_arb0_state_reg[1]/NET0131 ,
		_w2848_,
		_w2849_,
		_w2855_
	);
	LUT3 #(
		.INIT('h45)
	) name955 (
		_w2853_,
		_w2854_,
		_w2855_,
		_w2856_
	);
	LUT3 #(
		.INIT('h45)
	) name956 (
		\s10_msel_arb0_state_reg[0]/NET0131 ,
		_w2852_,
		_w2856_,
		_w2857_
	);
	LUT4 #(
		.INIT('hfd00)
	) name957 (
		\m1_s10_cyc_o_reg/NET0131 ,
		\rf_conf10_reg[2]/NET0131 ,
		\rf_conf10_reg[3]/NET0131 ,
		\s10_msel_arb0_state_reg[0]/NET0131 ,
		_w2858_
	);
	LUT2 #(
		.INIT('h4)
	) name958 (
		\s10_msel_arb0_state_reg[2]/NET0131 ,
		_w2858_,
		_w2859_
	);
	LUT4 #(
		.INIT('h5100)
	) name959 (
		\s10_msel_arb0_state_reg[1]/NET0131 ,
		_w2841_,
		_w2847_,
		_w2859_,
		_w2860_
	);
	LUT2 #(
		.INIT('h4)
	) name960 (
		\s10_msel_arb0_state_reg[0]/NET0131 ,
		\s10_msel_arb0_state_reg[1]/NET0131 ,
		_w2861_
	);
	LUT3 #(
		.INIT('h01)
	) name961 (
		_w2839_,
		_w2840_,
		_w2861_,
		_w2862_
	);
	LUT4 #(
		.INIT('h0002)
	) name962 (
		\m4_s10_cyc_o_reg/NET0131 ,
		\rf_conf10_reg[8]/NET0131 ,
		\rf_conf10_reg[9]/NET0131 ,
		\s10_msel_arb0_state_reg[0]/NET0131 ,
		_w2863_
	);
	LUT4 #(
		.INIT('h0004)
	) name963 (
		\s10_msel_arb0_state_reg[1]/NET0131 ,
		\s10_msel_arb0_state_reg[2]/NET0131 ,
		_w2843_,
		_w2863_,
		_w2864_
	);
	LUT4 #(
		.INIT('h5d00)
	) name964 (
		_w2846_,
		_w2850_,
		_w2862_,
		_w2864_,
		_w2865_
	);
	LUT2 #(
		.INIT('h1)
	) name965 (
		_w2860_,
		_w2865_,
		_w2866_
	);
	LUT2 #(
		.INIT('h2)
	) name966 (
		\s10_msel_arb0_state_reg[1]/NET0131 ,
		\s10_msel_arb0_state_reg[2]/NET0131 ,
		_w2867_
	);
	LUT2 #(
		.INIT('h8)
	) name967 (
		_w2839_,
		_w2867_,
		_w2868_
	);
	LUT4 #(
		.INIT('h1110)
	) name968 (
		_w2844_,
		_w2845_,
		_w2848_,
		_w2849_,
		_w2869_
	);
	LUT3 #(
		.INIT('h10)
	) name969 (
		_w2842_,
		_w2843_,
		_w2867_,
		_w2870_
	);
	LUT3 #(
		.INIT('h45)
	) name970 (
		_w2868_,
		_w2869_,
		_w2870_,
		_w2871_
	);
	LUT2 #(
		.INIT('h8)
	) name971 (
		\s10_msel_arb0_state_reg[1]/NET0131 ,
		\s10_msel_arb0_state_reg[2]/NET0131 ,
		_w2872_
	);
	LUT2 #(
		.INIT('h8)
	) name972 (
		_w2844_,
		_w2872_,
		_w2873_
	);
	LUT3 #(
		.INIT('h10)
	) name973 (
		_w2848_,
		_w2849_,
		_w2872_,
		_w2874_
	);
	LUT3 #(
		.INIT('h23)
	) name974 (
		_w2854_,
		_w2873_,
		_w2874_,
		_w2875_
	);
	LUT3 #(
		.INIT('h2a)
	) name975 (
		\s10_msel_arb0_state_reg[0]/NET0131 ,
		_w2871_,
		_w2875_,
		_w2876_
	);
	LUT3 #(
		.INIT('hfb)
	) name976 (
		_w2857_,
		_w2866_,
		_w2876_,
		_w2877_
	);
	LUT3 #(
		.INIT('h08)
	) name977 (
		\m3_s15_cyc_o_reg/NET0131 ,
		\rf_conf15_reg[6]/NET0131 ,
		\rf_conf15_reg[7]/NET0131 ,
		_w2878_
	);
	LUT3 #(
		.INIT('h08)
	) name978 (
		\m2_s15_cyc_o_reg/NET0131 ,
		\rf_conf15_reg[4]/NET0131 ,
		\rf_conf15_reg[5]/NET0131 ,
		_w2879_
	);
	LUT3 #(
		.INIT('h08)
	) name979 (
		\m0_s15_cyc_o_reg/NET0131 ,
		\rf_conf15_reg[0]/NET0131 ,
		\rf_conf15_reg[1]/NET0131 ,
		_w2880_
	);
	LUT3 #(
		.INIT('h08)
	) name980 (
		\m1_s15_cyc_o_reg/NET0131 ,
		\rf_conf15_reg[2]/NET0131 ,
		\rf_conf15_reg[3]/NET0131 ,
		_w2881_
	);
	LUT2 #(
		.INIT('h1)
	) name981 (
		_w2880_,
		_w2881_,
		_w2882_
	);
	LUT4 #(
		.INIT('h0001)
	) name982 (
		_w2878_,
		_w2879_,
		_w2880_,
		_w2881_,
		_w2883_
	);
	LUT3 #(
		.INIT('h08)
	) name983 (
		\m6_s15_cyc_o_reg/NET0131 ,
		\rf_conf15_reg[12]/NET0131 ,
		\rf_conf15_reg[13]/NET0131 ,
		_w2884_
	);
	LUT3 #(
		.INIT('h08)
	) name984 (
		\m7_s15_cyc_o_reg/NET0131 ,
		\rf_conf15_reg[14]/NET0131 ,
		\rf_conf15_reg[15]/NET0131 ,
		_w2885_
	);
	LUT3 #(
		.INIT('h08)
	) name985 (
		\m5_s15_cyc_o_reg/NET0131 ,
		\rf_conf15_reg[10]/NET0131 ,
		\rf_conf15_reg[11]/NET0131 ,
		_w2886_
	);
	LUT3 #(
		.INIT('h08)
	) name986 (
		\m4_s15_cyc_o_reg/NET0131 ,
		\rf_conf15_reg[8]/NET0131 ,
		\rf_conf15_reg[9]/NET0131 ,
		_w2887_
	);
	LUT2 #(
		.INIT('h1)
	) name987 (
		_w2886_,
		_w2887_,
		_w2888_
	);
	LUT4 #(
		.INIT('h0001)
	) name988 (
		_w2884_,
		_w2885_,
		_w2886_,
		_w2887_,
		_w2889_
	);
	LUT2 #(
		.INIT('h8)
	) name989 (
		_w2883_,
		_w2889_,
		_w2890_
	);
	LUT3 #(
		.INIT('h20)
	) name990 (
		\m3_s15_cyc_o_reg/NET0131 ,
		\rf_conf15_reg[6]/NET0131 ,
		\rf_conf15_reg[7]/NET0131 ,
		_w2891_
	);
	LUT3 #(
		.INIT('h20)
	) name991 (
		\m2_s15_cyc_o_reg/NET0131 ,
		\rf_conf15_reg[4]/NET0131 ,
		\rf_conf15_reg[5]/NET0131 ,
		_w2892_
	);
	LUT2 #(
		.INIT('h1)
	) name992 (
		_w2891_,
		_w2892_,
		_w2893_
	);
	LUT3 #(
		.INIT('h20)
	) name993 (
		\m0_s15_cyc_o_reg/NET0131 ,
		\rf_conf15_reg[0]/NET0131 ,
		\rf_conf15_reg[1]/NET0131 ,
		_w2894_
	);
	LUT3 #(
		.INIT('h20)
	) name994 (
		\m1_s15_cyc_o_reg/NET0131 ,
		\rf_conf15_reg[2]/NET0131 ,
		\rf_conf15_reg[3]/NET0131 ,
		_w2895_
	);
	LUT2 #(
		.INIT('h1)
	) name995 (
		_w2894_,
		_w2895_,
		_w2896_
	);
	LUT4 #(
		.INIT('h0001)
	) name996 (
		_w2891_,
		_w2892_,
		_w2894_,
		_w2895_,
		_w2897_
	);
	LUT3 #(
		.INIT('h20)
	) name997 (
		\m4_s15_cyc_o_reg/NET0131 ,
		\rf_conf15_reg[8]/NET0131 ,
		\rf_conf15_reg[9]/NET0131 ,
		_w2898_
	);
	LUT3 #(
		.INIT('h20)
	) name998 (
		\m5_s15_cyc_o_reg/NET0131 ,
		\rf_conf15_reg[10]/NET0131 ,
		\rf_conf15_reg[11]/NET0131 ,
		_w2899_
	);
	LUT3 #(
		.INIT('h20)
	) name999 (
		\m7_s15_cyc_o_reg/NET0131 ,
		\rf_conf15_reg[14]/NET0131 ,
		\rf_conf15_reg[15]/NET0131 ,
		_w2900_
	);
	LUT3 #(
		.INIT('h20)
	) name1000 (
		\m6_s15_cyc_o_reg/NET0131 ,
		\rf_conf15_reg[12]/NET0131 ,
		\rf_conf15_reg[13]/NET0131 ,
		_w2901_
	);
	LUT2 #(
		.INIT('h1)
	) name1001 (
		_w2900_,
		_w2901_,
		_w2902_
	);
	LUT4 #(
		.INIT('h0001)
	) name1002 (
		_w2898_,
		_w2899_,
		_w2900_,
		_w2901_,
		_w2903_
	);
	LUT3 #(
		.INIT('h80)
	) name1003 (
		\s15_next_reg/P0001 ,
		_w2897_,
		_w2903_,
		_w2904_
	);
	LUT3 #(
		.INIT('h80)
	) name1004 (
		\m3_s15_cyc_o_reg/NET0131 ,
		\rf_conf15_reg[6]/NET0131 ,
		\rf_conf15_reg[7]/NET0131 ,
		_w2905_
	);
	LUT3 #(
		.INIT('h80)
	) name1005 (
		\m2_s15_cyc_o_reg/NET0131 ,
		\rf_conf15_reg[4]/NET0131 ,
		\rf_conf15_reg[5]/NET0131 ,
		_w2906_
	);
	LUT2 #(
		.INIT('h1)
	) name1006 (
		_w2905_,
		_w2906_,
		_w2907_
	);
	LUT3 #(
		.INIT('h80)
	) name1007 (
		\m0_s15_cyc_o_reg/NET0131 ,
		\rf_conf15_reg[0]/NET0131 ,
		\rf_conf15_reg[1]/NET0131 ,
		_w2908_
	);
	LUT3 #(
		.INIT('h80)
	) name1008 (
		\m1_s15_cyc_o_reg/NET0131 ,
		\rf_conf15_reg[2]/NET0131 ,
		\rf_conf15_reg[3]/NET0131 ,
		_w2909_
	);
	LUT2 #(
		.INIT('h1)
	) name1009 (
		_w2908_,
		_w2909_,
		_w2910_
	);
	LUT4 #(
		.INIT('h0001)
	) name1010 (
		_w2905_,
		_w2906_,
		_w2908_,
		_w2909_,
		_w2911_
	);
	LUT3 #(
		.INIT('h80)
	) name1011 (
		\m7_s15_cyc_o_reg/NET0131 ,
		\rf_conf15_reg[14]/NET0131 ,
		\rf_conf15_reg[15]/NET0131 ,
		_w2912_
	);
	LUT3 #(
		.INIT('h80)
	) name1012 (
		\m6_s15_cyc_o_reg/NET0131 ,
		\rf_conf15_reg[12]/NET0131 ,
		\rf_conf15_reg[13]/NET0131 ,
		_w2913_
	);
	LUT3 #(
		.INIT('h80)
	) name1013 (
		\m4_s15_cyc_o_reg/NET0131 ,
		\rf_conf15_reg[8]/NET0131 ,
		\rf_conf15_reg[9]/NET0131 ,
		_w2914_
	);
	LUT3 #(
		.INIT('h80)
	) name1014 (
		\m5_s15_cyc_o_reg/NET0131 ,
		\rf_conf15_reg[10]/NET0131 ,
		\rf_conf15_reg[11]/NET0131 ,
		_w2915_
	);
	LUT4 #(
		.INIT('h0001)
	) name1015 (
		_w2912_,
		_w2913_,
		_w2914_,
		_w2915_,
		_w2916_
	);
	LUT2 #(
		.INIT('h8)
	) name1016 (
		_w2911_,
		_w2916_,
		_w2917_
	);
	LUT4 #(
		.INIT('hd111)
	) name1017 (
		\s15_msel_pri_out_reg[0]/NET0131 ,
		\s15_next_reg/P0001 ,
		_w2911_,
		_w2916_,
		_w2918_
	);
	LUT4 #(
		.INIT('h1055)
	) name1018 (
		rst_i_pad,
		_w2890_,
		_w2904_,
		_w2918_,
		_w2919_
	);
	LUT2 #(
		.INIT('h1)
	) name1019 (
		\s15_msel_arb3_state_reg[0]/NET0131 ,
		\s15_msel_arb3_state_reg[1]/NET0131 ,
		_w2920_
	);
	LUT4 #(
		.INIT('h0080)
	) name1020 (
		\m1_s15_cyc_o_reg/NET0131 ,
		\rf_conf15_reg[2]/NET0131 ,
		\rf_conf15_reg[3]/NET0131 ,
		\s15_msel_arb3_state_reg[1]/NET0131 ,
		_w2921_
	);
	LUT2 #(
		.INIT('h8)
	) name1021 (
		\s15_msel_arb3_state_reg[0]/NET0131 ,
		\s15_msel_arb3_state_reg[1]/NET0131 ,
		_w2922_
	);
	LUT4 #(
		.INIT('h007f)
	) name1022 (
		\m3_s15_cyc_o_reg/NET0131 ,
		\rf_conf15_reg[6]/NET0131 ,
		\rf_conf15_reg[7]/NET0131 ,
		\s15_msel_arb3_state_reg[2]/NET0131 ,
		_w2923_
	);
	LUT3 #(
		.INIT('hd0)
	) name1023 (
		_w2906_,
		_w2922_,
		_w2923_,
		_w2924_
	);
	LUT4 #(
		.INIT('h7477)
	) name1024 (
		_w2911_,
		_w2920_,
		_w2921_,
		_w2924_,
		_w2925_
	);
	LUT4 #(
		.INIT('h0080)
	) name1025 (
		\m5_s15_cyc_o_reg/NET0131 ,
		\rf_conf15_reg[10]/NET0131 ,
		\rf_conf15_reg[11]/NET0131 ,
		\s15_msel_arb3_state_reg[1]/NET0131 ,
		_w2926_
	);
	LUT3 #(
		.INIT('h07)
	) name1026 (
		_w2914_,
		_w2920_,
		_w2926_,
		_w2927_
	);
	LUT3 #(
		.INIT('h51)
	) name1027 (
		_w2912_,
		_w2913_,
		_w2922_,
		_w2928_
	);
	LUT4 #(
		.INIT('h8aaa)
	) name1028 (
		\s15_msel_arb3_state_reg[2]/NET0131 ,
		_w2911_,
		_w2927_,
		_w2928_,
		_w2929_
	);
	LUT3 #(
		.INIT('hf1)
	) name1029 (
		_w2916_,
		_w2925_,
		_w2929_,
		_w2930_
	);
	LUT4 #(
		.INIT('h0008)
	) name1030 (
		\m1_s15_cyc_o_reg/NET0131 ,
		\rf_conf15_reg[2]/NET0131 ,
		\rf_conf15_reg[3]/NET0131 ,
		\s15_msel_arb1_state_reg[1]/NET0131 ,
		_w2931_
	);
	LUT2 #(
		.INIT('h1)
	) name1031 (
		\s15_msel_arb1_state_reg[0]/NET0131 ,
		\s15_msel_arb1_state_reg[1]/NET0131 ,
		_w2932_
	);
	LUT3 #(
		.INIT('h13)
	) name1032 (
		_w2880_,
		_w2931_,
		_w2932_,
		_w2933_
	);
	LUT2 #(
		.INIT('h8)
	) name1033 (
		\s15_msel_arb1_state_reg[0]/NET0131 ,
		\s15_msel_arb1_state_reg[1]/NET0131 ,
		_w2934_
	);
	LUT3 #(
		.INIT('h51)
	) name1034 (
		_w2878_,
		_w2879_,
		_w2934_,
		_w2935_
	);
	LUT4 #(
		.INIT('h4555)
	) name1035 (
		\s15_msel_arb1_state_reg[2]/NET0131 ,
		_w2889_,
		_w2933_,
		_w2935_,
		_w2936_
	);
	LUT4 #(
		.INIT('h0008)
	) name1036 (
		\m4_s15_cyc_o_reg/NET0131 ,
		\rf_conf15_reg[8]/NET0131 ,
		\rf_conf15_reg[9]/NET0131 ,
		\s15_msel_arb1_state_reg[0]/NET0131 ,
		_w2937_
	);
	LUT3 #(
		.INIT('h54)
	) name1037 (
		\s15_msel_arb1_state_reg[1]/NET0131 ,
		_w2886_,
		_w2937_,
		_w2938_
	);
	LUT4 #(
		.INIT('hf700)
	) name1038 (
		\m7_s15_cyc_o_reg/NET0131 ,
		\rf_conf15_reg[14]/NET0131 ,
		\rf_conf15_reg[15]/NET0131 ,
		\s15_msel_arb1_state_reg[2]/NET0131 ,
		_w2939_
	);
	LUT3 #(
		.INIT('hd0)
	) name1039 (
		_w2884_,
		_w2934_,
		_w2939_,
		_w2940_
	);
	LUT3 #(
		.INIT('h10)
	) name1040 (
		_w2883_,
		_w2938_,
		_w2940_,
		_w2941_
	);
	LUT2 #(
		.INIT('h1)
	) name1041 (
		_w2936_,
		_w2941_,
		_w2942_
	);
	LUT3 #(
		.INIT('h80)
	) name1042 (
		\m5_s13_cyc_o_reg/NET0131 ,
		\rf_conf13_reg[10]/NET0131 ,
		\rf_conf13_reg[11]/NET0131 ,
		_w2943_
	);
	LUT3 #(
		.INIT('h80)
	) name1043 (
		\m4_s13_cyc_o_reg/NET0131 ,
		\rf_conf13_reg[8]/NET0131 ,
		\rf_conf13_reg[9]/NET0131 ,
		_w2944_
	);
	LUT3 #(
		.INIT('h01)
	) name1044 (
		\s13_msel_arb3_state_reg[0]/NET0131 ,
		_w2943_,
		_w2944_,
		_w2945_
	);
	LUT2 #(
		.INIT('h8)
	) name1045 (
		\s13_msel_arb3_state_reg[0]/NET0131 ,
		\s13_msel_arb3_state_reg[2]/NET0131 ,
		_w2946_
	);
	LUT3 #(
		.INIT('h13)
	) name1046 (
		\s13_msel_arb3_state_reg[0]/NET0131 ,
		\s13_msel_arb3_state_reg[1]/NET0131 ,
		\s13_msel_arb3_state_reg[2]/NET0131 ,
		_w2947_
	);
	LUT4 #(
		.INIT('h0080)
	) name1047 (
		\m5_s13_cyc_o_reg/NET0131 ,
		\rf_conf13_reg[10]/NET0131 ,
		\rf_conf13_reg[11]/NET0131 ,
		\s13_msel_arb3_state_reg[1]/NET0131 ,
		_w2948_
	);
	LUT2 #(
		.INIT('h1)
	) name1048 (
		_w2947_,
		_w2948_,
		_w2949_
	);
	LUT3 #(
		.INIT('h80)
	) name1049 (
		\m7_s13_cyc_o_reg/NET0131 ,
		\rf_conf13_reg[14]/NET0131 ,
		\rf_conf13_reg[15]/NET0131 ,
		_w2950_
	);
	LUT3 #(
		.INIT('h80)
	) name1050 (
		\m6_s13_cyc_o_reg/NET0131 ,
		\rf_conf13_reg[12]/NET0131 ,
		\rf_conf13_reg[13]/NET0131 ,
		_w2951_
	);
	LUT2 #(
		.INIT('h1)
	) name1051 (
		_w2950_,
		_w2951_,
		_w2952_
	);
	LUT3 #(
		.INIT('h80)
	) name1052 (
		\m3_s13_cyc_o_reg/NET0131 ,
		\rf_conf13_reg[6]/NET0131 ,
		\rf_conf13_reg[7]/NET0131 ,
		_w2953_
	);
	LUT3 #(
		.INIT('h80)
	) name1053 (
		\m2_s13_cyc_o_reg/NET0131 ,
		\rf_conf13_reg[4]/NET0131 ,
		\rf_conf13_reg[5]/NET0131 ,
		_w2954_
	);
	LUT3 #(
		.INIT('h80)
	) name1054 (
		\m1_s13_cyc_o_reg/NET0131 ,
		\rf_conf13_reg[2]/NET0131 ,
		\rf_conf13_reg[3]/NET0131 ,
		_w2955_
	);
	LUT3 #(
		.INIT('h80)
	) name1055 (
		\m0_s13_cyc_o_reg/NET0131 ,
		\rf_conf13_reg[0]/NET0131 ,
		\rf_conf13_reg[1]/NET0131 ,
		_w2956_
	);
	LUT4 #(
		.INIT('h0001)
	) name1056 (
		_w2953_,
		_w2954_,
		_w2955_,
		_w2956_,
		_w2957_
	);
	LUT4 #(
		.INIT('h00e0)
	) name1057 (
		_w2945_,
		_w2949_,
		_w2952_,
		_w2957_,
		_w2958_
	);
	LUT4 #(
		.INIT('h3332)
	) name1058 (
		\s13_msel_arb3_state_reg[0]/NET0131 ,
		\s13_msel_arb3_state_reg[1]/NET0131 ,
		_w2955_,
		_w2956_,
		_w2959_
	);
	LUT4 #(
		.INIT('h0001)
	) name1059 (
		_w2943_,
		_w2944_,
		_w2950_,
		_w2951_,
		_w2960_
	);
	LUT4 #(
		.INIT('h0080)
	) name1060 (
		\m2_s13_cyc_o_reg/NET0131 ,
		\rf_conf13_reg[4]/NET0131 ,
		\rf_conf13_reg[5]/NET0131 ,
		\s13_msel_arb3_state_reg[0]/NET0131 ,
		_w2961_
	);
	LUT2 #(
		.INIT('h1)
	) name1061 (
		\s13_msel_arb3_state_reg[2]/NET0131 ,
		_w2961_,
		_w2962_
	);
	LUT3 #(
		.INIT('h01)
	) name1062 (
		\s13_msel_arb3_state_reg[2]/NET0131 ,
		_w2953_,
		_w2961_,
		_w2963_
	);
	LUT3 #(
		.INIT('h10)
	) name1063 (
		_w2959_,
		_w2960_,
		_w2963_,
		_w2964_
	);
	LUT2 #(
		.INIT('h8)
	) name1064 (
		\s13_msel_arb3_state_reg[0]/NET0131 ,
		\s13_msel_arb3_state_reg[1]/NET0131 ,
		_w2965_
	);
	LUT4 #(
		.INIT('h7f00)
	) name1065 (
		\m2_s13_cyc_o_reg/NET0131 ,
		\rf_conf13_reg[4]/NET0131 ,
		\rf_conf13_reg[5]/NET0131 ,
		\s13_msel_arb3_state_reg[0]/NET0131 ,
		_w2966_
	);
	LUT3 #(
		.INIT('h10)
	) name1066 (
		_w2953_,
		_w2955_,
		_w2966_,
		_w2967_
	);
	LUT4 #(
		.INIT('h0b0a)
	) name1067 (
		\s13_msel_arb3_state_reg[2]/NET0131 ,
		_w2960_,
		_w2965_,
		_w2967_,
		_w2968_
	);
	LUT2 #(
		.INIT('h8)
	) name1068 (
		\s13_msel_arb3_state_reg[1]/NET0131 ,
		\s13_msel_arb3_state_reg[2]/NET0131 ,
		_w2969_
	);
	LUT3 #(
		.INIT('h80)
	) name1069 (
		\s13_msel_arb3_state_reg[0]/NET0131 ,
		\s13_msel_arb3_state_reg[1]/NET0131 ,
		\s13_msel_arb3_state_reg[2]/NET0131 ,
		_w2970_
	);
	LUT3 #(
		.INIT('he0)
	) name1070 (
		_w2950_,
		_w2957_,
		_w2970_,
		_w2971_
	);
	LUT4 #(
		.INIT('hdddc)
	) name1071 (
		_w2958_,
		_w2964_,
		_w2968_,
		_w2971_,
		_w2972_
	);
	LUT3 #(
		.INIT('h20)
	) name1072 (
		\m5_s14_cyc_o_reg/NET0131 ,
		\rf_conf14_reg[10]/NET0131 ,
		\rf_conf14_reg[11]/NET0131 ,
		_w2973_
	);
	LUT3 #(
		.INIT('h20)
	) name1073 (
		\m4_s14_cyc_o_reg/NET0131 ,
		\rf_conf14_reg[8]/NET0131 ,
		\rf_conf14_reg[9]/NET0131 ,
		_w2974_
	);
	LUT3 #(
		.INIT('h01)
	) name1074 (
		\s14_msel_arb2_state_reg[0]/NET0131 ,
		_w2973_,
		_w2974_,
		_w2975_
	);
	LUT2 #(
		.INIT('h8)
	) name1075 (
		\s14_msel_arb2_state_reg[0]/NET0131 ,
		\s14_msel_arb2_state_reg[2]/NET0131 ,
		_w2976_
	);
	LUT3 #(
		.INIT('h13)
	) name1076 (
		\s14_msel_arb2_state_reg[0]/NET0131 ,
		\s14_msel_arb2_state_reg[1]/NET0131 ,
		\s14_msel_arb2_state_reg[2]/NET0131 ,
		_w2977_
	);
	LUT4 #(
		.INIT('h0020)
	) name1077 (
		\m5_s14_cyc_o_reg/NET0131 ,
		\rf_conf14_reg[10]/NET0131 ,
		\rf_conf14_reg[11]/NET0131 ,
		\s14_msel_arb2_state_reg[1]/NET0131 ,
		_w2978_
	);
	LUT2 #(
		.INIT('h1)
	) name1078 (
		_w2977_,
		_w2978_,
		_w2979_
	);
	LUT3 #(
		.INIT('h20)
	) name1079 (
		\m7_s14_cyc_o_reg/NET0131 ,
		\rf_conf14_reg[14]/NET0131 ,
		\rf_conf14_reg[15]/NET0131 ,
		_w2980_
	);
	LUT3 #(
		.INIT('h20)
	) name1080 (
		\m6_s14_cyc_o_reg/NET0131 ,
		\rf_conf14_reg[12]/NET0131 ,
		\rf_conf14_reg[13]/NET0131 ,
		_w2981_
	);
	LUT2 #(
		.INIT('h1)
	) name1081 (
		_w2980_,
		_w2981_,
		_w2982_
	);
	LUT3 #(
		.INIT('h20)
	) name1082 (
		\m3_s14_cyc_o_reg/NET0131 ,
		\rf_conf14_reg[6]/NET0131 ,
		\rf_conf14_reg[7]/NET0131 ,
		_w2983_
	);
	LUT3 #(
		.INIT('h20)
	) name1083 (
		\m2_s14_cyc_o_reg/NET0131 ,
		\rf_conf14_reg[4]/NET0131 ,
		\rf_conf14_reg[5]/NET0131 ,
		_w2984_
	);
	LUT3 #(
		.INIT('h20)
	) name1084 (
		\m1_s14_cyc_o_reg/NET0131 ,
		\rf_conf14_reg[2]/NET0131 ,
		\rf_conf14_reg[3]/NET0131 ,
		_w2985_
	);
	LUT3 #(
		.INIT('h20)
	) name1085 (
		\m0_s14_cyc_o_reg/NET0131 ,
		\rf_conf14_reg[0]/NET0131 ,
		\rf_conf14_reg[1]/NET0131 ,
		_w2986_
	);
	LUT4 #(
		.INIT('h0001)
	) name1086 (
		_w2983_,
		_w2984_,
		_w2985_,
		_w2986_,
		_w2987_
	);
	LUT4 #(
		.INIT('h00e0)
	) name1087 (
		_w2975_,
		_w2979_,
		_w2982_,
		_w2987_,
		_w2988_
	);
	LUT4 #(
		.INIT('h3332)
	) name1088 (
		\s14_msel_arb2_state_reg[0]/NET0131 ,
		\s14_msel_arb2_state_reg[1]/NET0131 ,
		_w2985_,
		_w2986_,
		_w2989_
	);
	LUT4 #(
		.INIT('h0001)
	) name1089 (
		_w2973_,
		_w2974_,
		_w2980_,
		_w2981_,
		_w2990_
	);
	LUT4 #(
		.INIT('h0020)
	) name1090 (
		\m2_s14_cyc_o_reg/NET0131 ,
		\rf_conf14_reg[4]/NET0131 ,
		\rf_conf14_reg[5]/NET0131 ,
		\s14_msel_arb2_state_reg[0]/NET0131 ,
		_w2991_
	);
	LUT2 #(
		.INIT('h1)
	) name1091 (
		\s14_msel_arb2_state_reg[2]/NET0131 ,
		_w2991_,
		_w2992_
	);
	LUT3 #(
		.INIT('h01)
	) name1092 (
		\s14_msel_arb2_state_reg[2]/NET0131 ,
		_w2983_,
		_w2991_,
		_w2993_
	);
	LUT3 #(
		.INIT('h10)
	) name1093 (
		_w2989_,
		_w2990_,
		_w2993_,
		_w2994_
	);
	LUT2 #(
		.INIT('h8)
	) name1094 (
		\s14_msel_arb2_state_reg[0]/NET0131 ,
		\s14_msel_arb2_state_reg[1]/NET0131 ,
		_w2995_
	);
	LUT4 #(
		.INIT('hdf00)
	) name1095 (
		\m2_s14_cyc_o_reg/NET0131 ,
		\rf_conf14_reg[4]/NET0131 ,
		\rf_conf14_reg[5]/NET0131 ,
		\s14_msel_arb2_state_reg[0]/NET0131 ,
		_w2996_
	);
	LUT3 #(
		.INIT('h10)
	) name1096 (
		_w2983_,
		_w2985_,
		_w2996_,
		_w2997_
	);
	LUT4 #(
		.INIT('h0b0a)
	) name1097 (
		\s14_msel_arb2_state_reg[2]/NET0131 ,
		_w2990_,
		_w2995_,
		_w2997_,
		_w2998_
	);
	LUT2 #(
		.INIT('h8)
	) name1098 (
		\s14_msel_arb2_state_reg[1]/NET0131 ,
		\s14_msel_arb2_state_reg[2]/NET0131 ,
		_w2999_
	);
	LUT3 #(
		.INIT('h80)
	) name1099 (
		\s14_msel_arb2_state_reg[0]/NET0131 ,
		\s14_msel_arb2_state_reg[1]/NET0131 ,
		\s14_msel_arb2_state_reg[2]/NET0131 ,
		_w3000_
	);
	LUT3 #(
		.INIT('he0)
	) name1100 (
		_w2980_,
		_w2987_,
		_w3000_,
		_w3001_
	);
	LUT4 #(
		.INIT('hdddc)
	) name1101 (
		_w2988_,
		_w2994_,
		_w2998_,
		_w3001_,
		_w3002_
	);
	LUT3 #(
		.INIT('h80)
	) name1102 (
		\m5_s2_cyc_o_reg/NET0131 ,
		\rf_conf2_reg[10]/NET0131 ,
		\rf_conf2_reg[11]/NET0131 ,
		_w3003_
	);
	LUT3 #(
		.INIT('h80)
	) name1103 (
		\m4_s2_cyc_o_reg/NET0131 ,
		\rf_conf2_reg[8]/NET0131 ,
		\rf_conf2_reg[9]/NET0131 ,
		_w3004_
	);
	LUT3 #(
		.INIT('h01)
	) name1104 (
		\s2_msel_arb3_state_reg[0]/NET0131 ,
		_w3003_,
		_w3004_,
		_w3005_
	);
	LUT2 #(
		.INIT('h8)
	) name1105 (
		\s2_msel_arb3_state_reg[0]/NET0131 ,
		\s2_msel_arb3_state_reg[2]/NET0131 ,
		_w3006_
	);
	LUT3 #(
		.INIT('h13)
	) name1106 (
		\s2_msel_arb3_state_reg[0]/NET0131 ,
		\s2_msel_arb3_state_reg[1]/NET0131 ,
		\s2_msel_arb3_state_reg[2]/NET0131 ,
		_w3007_
	);
	LUT4 #(
		.INIT('h0080)
	) name1107 (
		\m5_s2_cyc_o_reg/NET0131 ,
		\rf_conf2_reg[10]/NET0131 ,
		\rf_conf2_reg[11]/NET0131 ,
		\s2_msel_arb3_state_reg[1]/NET0131 ,
		_w3008_
	);
	LUT2 #(
		.INIT('h1)
	) name1108 (
		_w3007_,
		_w3008_,
		_w3009_
	);
	LUT3 #(
		.INIT('h80)
	) name1109 (
		\m7_s2_cyc_o_reg/NET0131 ,
		\rf_conf2_reg[14]/NET0131 ,
		\rf_conf2_reg[15]/NET0131 ,
		_w3010_
	);
	LUT3 #(
		.INIT('h80)
	) name1110 (
		\m6_s2_cyc_o_reg/NET0131 ,
		\rf_conf2_reg[12]/NET0131 ,
		\rf_conf2_reg[13]/NET0131 ,
		_w3011_
	);
	LUT2 #(
		.INIT('h1)
	) name1111 (
		_w3010_,
		_w3011_,
		_w3012_
	);
	LUT3 #(
		.INIT('h80)
	) name1112 (
		\m3_s2_cyc_o_reg/NET0131 ,
		\rf_conf2_reg[6]/NET0131 ,
		\rf_conf2_reg[7]/NET0131 ,
		_w3013_
	);
	LUT3 #(
		.INIT('h80)
	) name1113 (
		\m2_s2_cyc_o_reg/NET0131 ,
		\rf_conf2_reg[4]/NET0131 ,
		\rf_conf2_reg[5]/NET0131 ,
		_w3014_
	);
	LUT3 #(
		.INIT('h80)
	) name1114 (
		\m1_s2_cyc_o_reg/NET0131 ,
		\rf_conf2_reg[2]/NET0131 ,
		\rf_conf2_reg[3]/NET0131 ,
		_w3015_
	);
	LUT3 #(
		.INIT('h80)
	) name1115 (
		\m0_s2_cyc_o_reg/NET0131 ,
		\rf_conf2_reg[0]/NET0131 ,
		\rf_conf2_reg[1]/NET0131 ,
		_w3016_
	);
	LUT4 #(
		.INIT('h0001)
	) name1116 (
		_w3013_,
		_w3014_,
		_w3015_,
		_w3016_,
		_w3017_
	);
	LUT4 #(
		.INIT('h00e0)
	) name1117 (
		_w3005_,
		_w3009_,
		_w3012_,
		_w3017_,
		_w3018_
	);
	LUT4 #(
		.INIT('h3332)
	) name1118 (
		\s2_msel_arb3_state_reg[0]/NET0131 ,
		\s2_msel_arb3_state_reg[1]/NET0131 ,
		_w3015_,
		_w3016_,
		_w3019_
	);
	LUT4 #(
		.INIT('h0001)
	) name1119 (
		_w3003_,
		_w3004_,
		_w3010_,
		_w3011_,
		_w3020_
	);
	LUT4 #(
		.INIT('h0080)
	) name1120 (
		\m2_s2_cyc_o_reg/NET0131 ,
		\rf_conf2_reg[4]/NET0131 ,
		\rf_conf2_reg[5]/NET0131 ,
		\s2_msel_arb3_state_reg[0]/NET0131 ,
		_w3021_
	);
	LUT2 #(
		.INIT('h1)
	) name1121 (
		\s2_msel_arb3_state_reg[2]/NET0131 ,
		_w3021_,
		_w3022_
	);
	LUT3 #(
		.INIT('h01)
	) name1122 (
		\s2_msel_arb3_state_reg[2]/NET0131 ,
		_w3013_,
		_w3021_,
		_w3023_
	);
	LUT3 #(
		.INIT('h10)
	) name1123 (
		_w3019_,
		_w3020_,
		_w3023_,
		_w3024_
	);
	LUT2 #(
		.INIT('h8)
	) name1124 (
		\s2_msel_arb3_state_reg[0]/NET0131 ,
		\s2_msel_arb3_state_reg[1]/NET0131 ,
		_w3025_
	);
	LUT4 #(
		.INIT('h7f00)
	) name1125 (
		\m2_s2_cyc_o_reg/NET0131 ,
		\rf_conf2_reg[4]/NET0131 ,
		\rf_conf2_reg[5]/NET0131 ,
		\s2_msel_arb3_state_reg[0]/NET0131 ,
		_w3026_
	);
	LUT3 #(
		.INIT('h10)
	) name1126 (
		_w3013_,
		_w3015_,
		_w3026_,
		_w3027_
	);
	LUT4 #(
		.INIT('h0b0a)
	) name1127 (
		\s2_msel_arb3_state_reg[2]/NET0131 ,
		_w3020_,
		_w3025_,
		_w3027_,
		_w3028_
	);
	LUT2 #(
		.INIT('h8)
	) name1128 (
		\s2_msel_arb3_state_reg[1]/NET0131 ,
		\s2_msel_arb3_state_reg[2]/NET0131 ,
		_w3029_
	);
	LUT3 #(
		.INIT('h80)
	) name1129 (
		\s2_msel_arb3_state_reg[0]/NET0131 ,
		\s2_msel_arb3_state_reg[1]/NET0131 ,
		\s2_msel_arb3_state_reg[2]/NET0131 ,
		_w3030_
	);
	LUT3 #(
		.INIT('he0)
	) name1130 (
		_w3010_,
		_w3017_,
		_w3030_,
		_w3031_
	);
	LUT4 #(
		.INIT('hdddc)
	) name1131 (
		_w3018_,
		_w3024_,
		_w3028_,
		_w3031_,
		_w3032_
	);
	LUT3 #(
		.INIT('h20)
	) name1132 (
		\m5_s3_cyc_o_reg/NET0131 ,
		\rf_conf3_reg[10]/NET0131 ,
		\rf_conf3_reg[11]/NET0131 ,
		_w3033_
	);
	LUT3 #(
		.INIT('h20)
	) name1133 (
		\m4_s3_cyc_o_reg/NET0131 ,
		\rf_conf3_reg[8]/NET0131 ,
		\rf_conf3_reg[9]/NET0131 ,
		_w3034_
	);
	LUT3 #(
		.INIT('h20)
	) name1134 (
		\m6_s3_cyc_o_reg/NET0131 ,
		\rf_conf3_reg[12]/NET0131 ,
		\rf_conf3_reg[13]/NET0131 ,
		_w3035_
	);
	LUT3 #(
		.INIT('h20)
	) name1135 (
		\m7_s3_cyc_o_reg/NET0131 ,
		\rf_conf3_reg[14]/NET0131 ,
		\rf_conf3_reg[15]/NET0131 ,
		_w3036_
	);
	LUT2 #(
		.INIT('h1)
	) name1136 (
		_w3035_,
		_w3036_,
		_w3037_
	);
	LUT4 #(
		.INIT('h0001)
	) name1137 (
		_w3033_,
		_w3034_,
		_w3035_,
		_w3036_,
		_w3038_
	);
	LUT3 #(
		.INIT('h20)
	) name1138 (
		\m3_s3_cyc_o_reg/NET0131 ,
		\rf_conf3_reg[6]/NET0131 ,
		\rf_conf3_reg[7]/NET0131 ,
		_w3039_
	);
	LUT4 #(
		.INIT('h00df)
	) name1139 (
		\m3_s3_cyc_o_reg/NET0131 ,
		\rf_conf3_reg[6]/NET0131 ,
		\rf_conf3_reg[7]/NET0131 ,
		\s3_msel_arb2_state_reg[2]/NET0131 ,
		_w3040_
	);
	LUT3 #(
		.INIT('h20)
	) name1140 (
		\m2_s3_cyc_o_reg/NET0131 ,
		\rf_conf3_reg[4]/NET0131 ,
		\rf_conf3_reg[5]/NET0131 ,
		_w3041_
	);
	LUT4 #(
		.INIT('h0020)
	) name1141 (
		\m0_s3_cyc_o_reg/NET0131 ,
		\rf_conf3_reg[0]/NET0131 ,
		\rf_conf3_reg[1]/NET0131 ,
		\s3_msel_arb2_state_reg[1]/NET0131 ,
		_w3042_
	);
	LUT3 #(
		.INIT('h54)
	) name1142 (
		\s3_msel_arb2_state_reg[0]/NET0131 ,
		_w3041_,
		_w3042_,
		_w3043_
	);
	LUT3 #(
		.INIT('h20)
	) name1143 (
		\m1_s3_cyc_o_reg/NET0131 ,
		\rf_conf3_reg[2]/NET0131 ,
		\rf_conf3_reg[3]/NET0131 ,
		_w3044_
	);
	LUT3 #(
		.INIT('h54)
	) name1144 (
		\s3_msel_arb2_state_reg[1]/NET0131 ,
		_w3041_,
		_w3044_,
		_w3045_
	);
	LUT4 #(
		.INIT('h0004)
	) name1145 (
		_w3038_,
		_w3040_,
		_w3043_,
		_w3045_,
		_w3046_
	);
	LUT2 #(
		.INIT('h1)
	) name1146 (
		_w3039_,
		_w3041_,
		_w3047_
	);
	LUT3 #(
		.INIT('h20)
	) name1147 (
		\m0_s3_cyc_o_reg/NET0131 ,
		\rf_conf3_reg[0]/NET0131 ,
		\rf_conf3_reg[1]/NET0131 ,
		_w3048_
	);
	LUT4 #(
		.INIT('h0001)
	) name1148 (
		_w3039_,
		_w3041_,
		_w3044_,
		_w3048_,
		_w3049_
	);
	LUT4 #(
		.INIT('h0020)
	) name1149 (
		\m4_s3_cyc_o_reg/NET0131 ,
		\rf_conf3_reg[8]/NET0131 ,
		\rf_conf3_reg[9]/NET0131 ,
		\s3_msel_arb2_state_reg[1]/NET0131 ,
		_w3050_
	);
	LUT3 #(
		.INIT('h54)
	) name1150 (
		\s3_msel_arb2_state_reg[0]/NET0131 ,
		_w3035_,
		_w3050_,
		_w3051_
	);
	LUT3 #(
		.INIT('h54)
	) name1151 (
		\s3_msel_arb2_state_reg[1]/NET0131 ,
		_w3033_,
		_w3035_,
		_w3052_
	);
	LUT4 #(
		.INIT('h0001)
	) name1152 (
		_w3036_,
		_w3049_,
		_w3051_,
		_w3052_,
		_w3053_
	);
	LUT3 #(
		.INIT('hce)
	) name1153 (
		\s3_msel_arb2_state_reg[2]/NET0131 ,
		_w3046_,
		_w3053_,
		_w3054_
	);
	LUT2 #(
		.INIT('h4)
	) name1154 (
		\s4_msel_arb3_state_reg[1]/NET0131 ,
		\s4_msel_arb3_state_reg[2]/NET0131 ,
		_w3055_
	);
	LUT3 #(
		.INIT('h80)
	) name1155 (
		\m1_s4_cyc_o_reg/NET0131 ,
		\rf_conf4_reg[2]/NET0131 ,
		\rf_conf4_reg[3]/NET0131 ,
		_w3056_
	);
	LUT3 #(
		.INIT('h80)
	) name1156 (
		\m0_s4_cyc_o_reg/NET0131 ,
		\rf_conf4_reg[0]/NET0131 ,
		\rf_conf4_reg[1]/NET0131 ,
		_w3057_
	);
	LUT3 #(
		.INIT('h80)
	) name1157 (
		\m3_s4_cyc_o_reg/NET0131 ,
		\rf_conf4_reg[6]/NET0131 ,
		\rf_conf4_reg[7]/NET0131 ,
		_w3058_
	);
	LUT3 #(
		.INIT('h80)
	) name1158 (
		\m2_s4_cyc_o_reg/NET0131 ,
		\rf_conf4_reg[4]/NET0131 ,
		\rf_conf4_reg[5]/NET0131 ,
		_w3059_
	);
	LUT4 #(
		.INIT('h0001)
	) name1159 (
		_w3056_,
		_w3057_,
		_w3058_,
		_w3059_,
		_w3060_
	);
	LUT3 #(
		.INIT('h80)
	) name1160 (
		\m5_s4_cyc_o_reg/NET0131 ,
		\rf_conf4_reg[10]/NET0131 ,
		\rf_conf4_reg[11]/NET0131 ,
		_w3061_
	);
	LUT3 #(
		.INIT('h80)
	) name1161 (
		\m7_s4_cyc_o_reg/NET0131 ,
		\rf_conf4_reg[14]/NET0131 ,
		\rf_conf4_reg[15]/NET0131 ,
		_w3062_
	);
	LUT3 #(
		.INIT('h80)
	) name1162 (
		\m6_s4_cyc_o_reg/NET0131 ,
		\rf_conf4_reg[12]/NET0131 ,
		\rf_conf4_reg[13]/NET0131 ,
		_w3063_
	);
	LUT2 #(
		.INIT('h1)
	) name1163 (
		_w3062_,
		_w3063_,
		_w3064_
	);
	LUT3 #(
		.INIT('h01)
	) name1164 (
		_w3061_,
		_w3062_,
		_w3063_,
		_w3065_
	);
	LUT3 #(
		.INIT('h8a)
	) name1165 (
		_w3055_,
		_w3060_,
		_w3065_,
		_w3066_
	);
	LUT2 #(
		.INIT('h8)
	) name1166 (
		\s4_msel_arb3_state_reg[1]/NET0131 ,
		\s4_msel_arb3_state_reg[2]/NET0131 ,
		_w3067_
	);
	LUT3 #(
		.INIT('he0)
	) name1167 (
		_w3060_,
		_w3062_,
		_w3067_,
		_w3068_
	);
	LUT3 #(
		.INIT('h80)
	) name1168 (
		\m4_s4_cyc_o_reg/NET0131 ,
		\rf_conf4_reg[8]/NET0131 ,
		\rf_conf4_reg[9]/NET0131 ,
		_w3069_
	);
	LUT2 #(
		.INIT('h1)
	) name1169 (
		_w3061_,
		_w3069_,
		_w3070_
	);
	LUT4 #(
		.INIT('h0001)
	) name1170 (
		_w3061_,
		_w3062_,
		_w3063_,
		_w3069_,
		_w3071_
	);
	LUT4 #(
		.INIT('h007f)
	) name1171 (
		\m1_s4_cyc_o_reg/NET0131 ,
		\rf_conf4_reg[2]/NET0131 ,
		\rf_conf4_reg[3]/NET0131 ,
		\s4_msel_arb3_state_reg[2]/NET0131 ,
		_w3072_
	);
	LUT4 #(
		.INIT('h007f)
	) name1172 (
		\m2_s4_cyc_o_reg/NET0131 ,
		\rf_conf4_reg[4]/NET0131 ,
		\rf_conf4_reg[5]/NET0131 ,
		\s4_msel_arb3_state_reg[1]/NET0131 ,
		_w3073_
	);
	LUT2 #(
		.INIT('h8)
	) name1173 (
		_w3072_,
		_w3073_,
		_w3074_
	);
	LUT3 #(
		.INIT('h10)
	) name1174 (
		_w3058_,
		_w3071_,
		_w3074_,
		_w3075_
	);
	LUT4 #(
		.INIT('haaa8)
	) name1175 (
		\s4_msel_arb3_state_reg[0]/NET0131 ,
		_w3066_,
		_w3068_,
		_w3075_,
		_w3076_
	);
	LUT4 #(
		.INIT('h0080)
	) name1176 (
		\m2_s4_cyc_o_reg/NET0131 ,
		\rf_conf4_reg[4]/NET0131 ,
		\rf_conf4_reg[5]/NET0131 ,
		\s4_msel_arb3_state_reg[0]/NET0131 ,
		_w3077_
	);
	LUT3 #(
		.INIT('h54)
	) name1177 (
		\s4_msel_arb3_state_reg[1]/NET0131 ,
		_w3056_,
		_w3057_,
		_w3078_
	);
	LUT4 #(
		.INIT('h00ab)
	) name1178 (
		\s4_msel_arb3_state_reg[1]/NET0131 ,
		_w3056_,
		_w3057_,
		_w3077_,
		_w3079_
	);
	LUT4 #(
		.INIT('h5455)
	) name1179 (
		\s4_msel_arb3_state_reg[2]/NET0131 ,
		_w3058_,
		_w3071_,
		_w3079_,
		_w3080_
	);
	LUT2 #(
		.INIT('h2)
	) name1180 (
		\s4_msel_arb3_state_reg[1]/NET0131 ,
		\s4_msel_arb3_state_reg[2]/NET0131 ,
		_w3081_
	);
	LUT3 #(
		.INIT('ha2)
	) name1181 (
		\s4_msel_arb3_state_reg[0]/NET0131 ,
		\s4_msel_arb3_state_reg[1]/NET0131 ,
		\s4_msel_arb3_state_reg[2]/NET0131 ,
		_w3082_
	);
	LUT3 #(
		.INIT('h32)
	) name1182 (
		_w3061_,
		_w3067_,
		_w3069_,
		_w3083_
	);
	LUT4 #(
		.INIT('h0f0b)
	) name1183 (
		_w3060_,
		_w3064_,
		_w3082_,
		_w3083_,
		_w3084_
	);
	LUT2 #(
		.INIT('h4)
	) name1184 (
		_w3080_,
		_w3084_,
		_w3085_
	);
	LUT2 #(
		.INIT('he)
	) name1185 (
		_w3076_,
		_w3085_,
		_w3086_
	);
	LUT3 #(
		.INIT('h20)
	) name1186 (
		\m5_s6_cyc_o_reg/NET0131 ,
		\rf_conf6_reg[10]/NET0131 ,
		\rf_conf6_reg[11]/NET0131 ,
		_w3087_
	);
	LUT3 #(
		.INIT('h20)
	) name1187 (
		\m4_s6_cyc_o_reg/NET0131 ,
		\rf_conf6_reg[8]/NET0131 ,
		\rf_conf6_reg[9]/NET0131 ,
		_w3088_
	);
	LUT3 #(
		.INIT('h20)
	) name1188 (
		\m6_s6_cyc_o_reg/NET0131 ,
		\rf_conf6_reg[12]/NET0131 ,
		\rf_conf6_reg[13]/NET0131 ,
		_w3089_
	);
	LUT3 #(
		.INIT('h20)
	) name1189 (
		\m7_s6_cyc_o_reg/NET0131 ,
		\rf_conf6_reg[14]/NET0131 ,
		\rf_conf6_reg[15]/NET0131 ,
		_w3090_
	);
	LUT2 #(
		.INIT('h1)
	) name1190 (
		_w3089_,
		_w3090_,
		_w3091_
	);
	LUT4 #(
		.INIT('h0001)
	) name1191 (
		_w3087_,
		_w3088_,
		_w3089_,
		_w3090_,
		_w3092_
	);
	LUT3 #(
		.INIT('h20)
	) name1192 (
		\m3_s6_cyc_o_reg/NET0131 ,
		\rf_conf6_reg[6]/NET0131 ,
		\rf_conf6_reg[7]/NET0131 ,
		_w3093_
	);
	LUT4 #(
		.INIT('h00df)
	) name1193 (
		\m3_s6_cyc_o_reg/NET0131 ,
		\rf_conf6_reg[6]/NET0131 ,
		\rf_conf6_reg[7]/NET0131 ,
		\s6_msel_arb2_state_reg[2]/NET0131 ,
		_w3094_
	);
	LUT3 #(
		.INIT('h20)
	) name1194 (
		\m2_s6_cyc_o_reg/NET0131 ,
		\rf_conf6_reg[4]/NET0131 ,
		\rf_conf6_reg[5]/NET0131 ,
		_w3095_
	);
	LUT4 #(
		.INIT('h0020)
	) name1195 (
		\m0_s6_cyc_o_reg/NET0131 ,
		\rf_conf6_reg[0]/NET0131 ,
		\rf_conf6_reg[1]/NET0131 ,
		\s6_msel_arb2_state_reg[1]/NET0131 ,
		_w3096_
	);
	LUT3 #(
		.INIT('h54)
	) name1196 (
		\s6_msel_arb2_state_reg[0]/NET0131 ,
		_w3095_,
		_w3096_,
		_w3097_
	);
	LUT3 #(
		.INIT('h20)
	) name1197 (
		\m1_s6_cyc_o_reg/NET0131 ,
		\rf_conf6_reg[2]/NET0131 ,
		\rf_conf6_reg[3]/NET0131 ,
		_w3098_
	);
	LUT3 #(
		.INIT('h54)
	) name1198 (
		\s6_msel_arb2_state_reg[1]/NET0131 ,
		_w3095_,
		_w3098_,
		_w3099_
	);
	LUT4 #(
		.INIT('h0004)
	) name1199 (
		_w3092_,
		_w3094_,
		_w3097_,
		_w3099_,
		_w3100_
	);
	LUT2 #(
		.INIT('h1)
	) name1200 (
		_w3093_,
		_w3095_,
		_w3101_
	);
	LUT3 #(
		.INIT('h20)
	) name1201 (
		\m0_s6_cyc_o_reg/NET0131 ,
		\rf_conf6_reg[0]/NET0131 ,
		\rf_conf6_reg[1]/NET0131 ,
		_w3102_
	);
	LUT4 #(
		.INIT('h0001)
	) name1202 (
		_w3093_,
		_w3095_,
		_w3098_,
		_w3102_,
		_w3103_
	);
	LUT4 #(
		.INIT('h0020)
	) name1203 (
		\m4_s6_cyc_o_reg/NET0131 ,
		\rf_conf6_reg[8]/NET0131 ,
		\rf_conf6_reg[9]/NET0131 ,
		\s6_msel_arb2_state_reg[1]/NET0131 ,
		_w3104_
	);
	LUT3 #(
		.INIT('h54)
	) name1204 (
		\s6_msel_arb2_state_reg[0]/NET0131 ,
		_w3089_,
		_w3104_,
		_w3105_
	);
	LUT3 #(
		.INIT('h54)
	) name1205 (
		\s6_msel_arb2_state_reg[1]/NET0131 ,
		_w3087_,
		_w3089_,
		_w3106_
	);
	LUT4 #(
		.INIT('h0001)
	) name1206 (
		_w3090_,
		_w3103_,
		_w3105_,
		_w3106_,
		_w3107_
	);
	LUT3 #(
		.INIT('hce)
	) name1207 (
		\s6_msel_arb2_state_reg[2]/NET0131 ,
		_w3100_,
		_w3107_,
		_w3108_
	);
	LUT3 #(
		.INIT('h20)
	) name1208 (
		\m5_s8_cyc_o_reg/NET0131 ,
		\rf_conf8_reg[10]/NET0131 ,
		\rf_conf8_reg[11]/NET0131 ,
		_w3109_
	);
	LUT3 #(
		.INIT('h20)
	) name1209 (
		\m4_s8_cyc_o_reg/NET0131 ,
		\rf_conf8_reg[8]/NET0131 ,
		\rf_conf8_reg[9]/NET0131 ,
		_w3110_
	);
	LUT3 #(
		.INIT('h20)
	) name1210 (
		\m6_s8_cyc_o_reg/NET0131 ,
		\rf_conf8_reg[12]/NET0131 ,
		\rf_conf8_reg[13]/NET0131 ,
		_w3111_
	);
	LUT3 #(
		.INIT('h20)
	) name1211 (
		\m7_s8_cyc_o_reg/NET0131 ,
		\rf_conf8_reg[14]/NET0131 ,
		\rf_conf8_reg[15]/NET0131 ,
		_w3112_
	);
	LUT2 #(
		.INIT('h1)
	) name1212 (
		_w3111_,
		_w3112_,
		_w3113_
	);
	LUT4 #(
		.INIT('h0001)
	) name1213 (
		_w3109_,
		_w3110_,
		_w3111_,
		_w3112_,
		_w3114_
	);
	LUT3 #(
		.INIT('h20)
	) name1214 (
		\m3_s8_cyc_o_reg/NET0131 ,
		\rf_conf8_reg[6]/NET0131 ,
		\rf_conf8_reg[7]/NET0131 ,
		_w3115_
	);
	LUT4 #(
		.INIT('h00df)
	) name1215 (
		\m3_s8_cyc_o_reg/NET0131 ,
		\rf_conf8_reg[6]/NET0131 ,
		\rf_conf8_reg[7]/NET0131 ,
		\s8_msel_arb2_state_reg[2]/NET0131 ,
		_w3116_
	);
	LUT3 #(
		.INIT('h20)
	) name1216 (
		\m2_s8_cyc_o_reg/NET0131 ,
		\rf_conf8_reg[4]/NET0131 ,
		\rf_conf8_reg[5]/NET0131 ,
		_w3117_
	);
	LUT4 #(
		.INIT('h0020)
	) name1217 (
		\m0_s8_cyc_o_reg/NET0131 ,
		\rf_conf8_reg[0]/NET0131 ,
		\rf_conf8_reg[1]/NET0131 ,
		\s8_msel_arb2_state_reg[1]/NET0131 ,
		_w3118_
	);
	LUT3 #(
		.INIT('h54)
	) name1218 (
		\s8_msel_arb2_state_reg[0]/NET0131 ,
		_w3117_,
		_w3118_,
		_w3119_
	);
	LUT3 #(
		.INIT('h20)
	) name1219 (
		\m1_s8_cyc_o_reg/NET0131 ,
		\rf_conf8_reg[2]/NET0131 ,
		\rf_conf8_reg[3]/NET0131 ,
		_w3120_
	);
	LUT3 #(
		.INIT('h54)
	) name1220 (
		\s8_msel_arb2_state_reg[1]/NET0131 ,
		_w3117_,
		_w3120_,
		_w3121_
	);
	LUT4 #(
		.INIT('h0004)
	) name1221 (
		_w3114_,
		_w3116_,
		_w3119_,
		_w3121_,
		_w3122_
	);
	LUT2 #(
		.INIT('h1)
	) name1222 (
		_w3115_,
		_w3117_,
		_w3123_
	);
	LUT3 #(
		.INIT('h20)
	) name1223 (
		\m0_s8_cyc_o_reg/NET0131 ,
		\rf_conf8_reg[0]/NET0131 ,
		\rf_conf8_reg[1]/NET0131 ,
		_w3124_
	);
	LUT4 #(
		.INIT('h0001)
	) name1224 (
		_w3115_,
		_w3117_,
		_w3120_,
		_w3124_,
		_w3125_
	);
	LUT4 #(
		.INIT('h0020)
	) name1225 (
		\m4_s8_cyc_o_reg/NET0131 ,
		\rf_conf8_reg[8]/NET0131 ,
		\rf_conf8_reg[9]/NET0131 ,
		\s8_msel_arb2_state_reg[1]/NET0131 ,
		_w3126_
	);
	LUT3 #(
		.INIT('h54)
	) name1226 (
		\s8_msel_arb2_state_reg[0]/NET0131 ,
		_w3111_,
		_w3126_,
		_w3127_
	);
	LUT3 #(
		.INIT('h54)
	) name1227 (
		\s8_msel_arb2_state_reg[1]/NET0131 ,
		_w3109_,
		_w3111_,
		_w3128_
	);
	LUT4 #(
		.INIT('h0001)
	) name1228 (
		_w3112_,
		_w3125_,
		_w3127_,
		_w3128_,
		_w3129_
	);
	LUT3 #(
		.INIT('hce)
	) name1229 (
		\s8_msel_arb2_state_reg[2]/NET0131 ,
		_w3122_,
		_w3129_,
		_w3130_
	);
	LUT3 #(
		.INIT('h20)
	) name1230 (
		\m5_s0_cyc_o_reg/NET0131 ,
		\rf_conf0_reg[10]/NET0131 ,
		\rf_conf0_reg[11]/NET0131 ,
		_w3131_
	);
	LUT3 #(
		.INIT('h20)
	) name1231 (
		\m4_s0_cyc_o_reg/NET0131 ,
		\rf_conf0_reg[8]/NET0131 ,
		\rf_conf0_reg[9]/NET0131 ,
		_w3132_
	);
	LUT3 #(
		.INIT('h20)
	) name1232 (
		\m6_s0_cyc_o_reg/NET0131 ,
		\rf_conf0_reg[12]/NET0131 ,
		\rf_conf0_reg[13]/NET0131 ,
		_w3133_
	);
	LUT3 #(
		.INIT('h20)
	) name1233 (
		\m7_s0_cyc_o_reg/NET0131 ,
		\rf_conf0_reg[14]/NET0131 ,
		\rf_conf0_reg[15]/NET0131 ,
		_w3134_
	);
	LUT2 #(
		.INIT('h1)
	) name1234 (
		_w3133_,
		_w3134_,
		_w3135_
	);
	LUT4 #(
		.INIT('h0001)
	) name1235 (
		_w3131_,
		_w3132_,
		_w3133_,
		_w3134_,
		_w3136_
	);
	LUT3 #(
		.INIT('h20)
	) name1236 (
		\m3_s0_cyc_o_reg/NET0131 ,
		\rf_conf0_reg[6]/NET0131 ,
		\rf_conf0_reg[7]/NET0131 ,
		_w3137_
	);
	LUT4 #(
		.INIT('h00df)
	) name1237 (
		\m3_s0_cyc_o_reg/NET0131 ,
		\rf_conf0_reg[6]/NET0131 ,
		\rf_conf0_reg[7]/NET0131 ,
		\s0_msel_arb2_state_reg[2]/NET0131 ,
		_w3138_
	);
	LUT3 #(
		.INIT('h20)
	) name1238 (
		\m2_s0_cyc_o_reg/NET0131 ,
		\rf_conf0_reg[4]/NET0131 ,
		\rf_conf0_reg[5]/NET0131 ,
		_w3139_
	);
	LUT4 #(
		.INIT('h0020)
	) name1239 (
		\m0_s0_cyc_o_reg/NET0131 ,
		\rf_conf0_reg[0]/NET0131 ,
		\rf_conf0_reg[1]/NET0131 ,
		\s0_msel_arb2_state_reg[1]/NET0131 ,
		_w3140_
	);
	LUT3 #(
		.INIT('h54)
	) name1240 (
		\s0_msel_arb2_state_reg[0]/NET0131 ,
		_w3139_,
		_w3140_,
		_w3141_
	);
	LUT3 #(
		.INIT('h20)
	) name1241 (
		\m1_s0_cyc_o_reg/NET0131 ,
		\rf_conf0_reg[2]/NET0131 ,
		\rf_conf0_reg[3]/NET0131 ,
		_w3142_
	);
	LUT3 #(
		.INIT('h54)
	) name1242 (
		\s0_msel_arb2_state_reg[1]/NET0131 ,
		_w3139_,
		_w3142_,
		_w3143_
	);
	LUT4 #(
		.INIT('h0004)
	) name1243 (
		_w3136_,
		_w3138_,
		_w3141_,
		_w3143_,
		_w3144_
	);
	LUT2 #(
		.INIT('h1)
	) name1244 (
		_w3137_,
		_w3139_,
		_w3145_
	);
	LUT3 #(
		.INIT('h20)
	) name1245 (
		\m0_s0_cyc_o_reg/NET0131 ,
		\rf_conf0_reg[0]/NET0131 ,
		\rf_conf0_reg[1]/NET0131 ,
		_w3146_
	);
	LUT4 #(
		.INIT('h0001)
	) name1246 (
		_w3137_,
		_w3139_,
		_w3142_,
		_w3146_,
		_w3147_
	);
	LUT4 #(
		.INIT('h0020)
	) name1247 (
		\m4_s0_cyc_o_reg/NET0131 ,
		\rf_conf0_reg[8]/NET0131 ,
		\rf_conf0_reg[9]/NET0131 ,
		\s0_msel_arb2_state_reg[1]/NET0131 ,
		_w3148_
	);
	LUT3 #(
		.INIT('h54)
	) name1248 (
		\s0_msel_arb2_state_reg[0]/NET0131 ,
		_w3133_,
		_w3148_,
		_w3149_
	);
	LUT3 #(
		.INIT('h54)
	) name1249 (
		\s0_msel_arb2_state_reg[1]/NET0131 ,
		_w3131_,
		_w3133_,
		_w3150_
	);
	LUT4 #(
		.INIT('h0001)
	) name1250 (
		_w3134_,
		_w3147_,
		_w3149_,
		_w3150_,
		_w3151_
	);
	LUT3 #(
		.INIT('hce)
	) name1251 (
		\s0_msel_arb2_state_reg[2]/NET0131 ,
		_w3144_,
		_w3151_,
		_w3152_
	);
	LUT3 #(
		.INIT('h80)
	) name1252 (
		\m5_s10_cyc_o_reg/NET0131 ,
		\rf_conf10_reg[10]/NET0131 ,
		\rf_conf10_reg[11]/NET0131 ,
		_w3153_
	);
	LUT3 #(
		.INIT('h80)
	) name1253 (
		\m4_s10_cyc_o_reg/NET0131 ,
		\rf_conf10_reg[8]/NET0131 ,
		\rf_conf10_reg[9]/NET0131 ,
		_w3154_
	);
	LUT3 #(
		.INIT('h01)
	) name1254 (
		\s10_msel_arb3_state_reg[0]/NET0131 ,
		_w3153_,
		_w3154_,
		_w3155_
	);
	LUT2 #(
		.INIT('h8)
	) name1255 (
		\s10_msel_arb3_state_reg[0]/NET0131 ,
		\s10_msel_arb3_state_reg[2]/NET0131 ,
		_w3156_
	);
	LUT3 #(
		.INIT('h13)
	) name1256 (
		\s10_msel_arb3_state_reg[0]/NET0131 ,
		\s10_msel_arb3_state_reg[1]/NET0131 ,
		\s10_msel_arb3_state_reg[2]/NET0131 ,
		_w3157_
	);
	LUT4 #(
		.INIT('h0080)
	) name1257 (
		\m5_s10_cyc_o_reg/NET0131 ,
		\rf_conf10_reg[10]/NET0131 ,
		\rf_conf10_reg[11]/NET0131 ,
		\s10_msel_arb3_state_reg[1]/NET0131 ,
		_w3158_
	);
	LUT2 #(
		.INIT('h1)
	) name1258 (
		_w3157_,
		_w3158_,
		_w3159_
	);
	LUT3 #(
		.INIT('h80)
	) name1259 (
		\m7_s10_cyc_o_reg/NET0131 ,
		\rf_conf10_reg[14]/NET0131 ,
		\rf_conf10_reg[15]/NET0131 ,
		_w3160_
	);
	LUT3 #(
		.INIT('h80)
	) name1260 (
		\m6_s10_cyc_o_reg/NET0131 ,
		\rf_conf10_reg[12]/NET0131 ,
		\rf_conf10_reg[13]/NET0131 ,
		_w3161_
	);
	LUT2 #(
		.INIT('h1)
	) name1261 (
		_w3160_,
		_w3161_,
		_w3162_
	);
	LUT3 #(
		.INIT('h80)
	) name1262 (
		\m3_s10_cyc_o_reg/NET0131 ,
		\rf_conf10_reg[6]/NET0131 ,
		\rf_conf10_reg[7]/NET0131 ,
		_w3163_
	);
	LUT3 #(
		.INIT('h80)
	) name1263 (
		\m2_s10_cyc_o_reg/NET0131 ,
		\rf_conf10_reg[4]/NET0131 ,
		\rf_conf10_reg[5]/NET0131 ,
		_w3164_
	);
	LUT3 #(
		.INIT('h80)
	) name1264 (
		\m1_s10_cyc_o_reg/NET0131 ,
		\rf_conf10_reg[2]/NET0131 ,
		\rf_conf10_reg[3]/NET0131 ,
		_w3165_
	);
	LUT3 #(
		.INIT('h80)
	) name1265 (
		\m0_s10_cyc_o_reg/NET0131 ,
		\rf_conf10_reg[0]/NET0131 ,
		\rf_conf10_reg[1]/NET0131 ,
		_w3166_
	);
	LUT4 #(
		.INIT('h0001)
	) name1266 (
		_w3163_,
		_w3164_,
		_w3165_,
		_w3166_,
		_w3167_
	);
	LUT4 #(
		.INIT('h00e0)
	) name1267 (
		_w3155_,
		_w3159_,
		_w3162_,
		_w3167_,
		_w3168_
	);
	LUT4 #(
		.INIT('h3332)
	) name1268 (
		\s10_msel_arb3_state_reg[0]/NET0131 ,
		\s10_msel_arb3_state_reg[1]/NET0131 ,
		_w3165_,
		_w3166_,
		_w3169_
	);
	LUT4 #(
		.INIT('h0001)
	) name1269 (
		_w3153_,
		_w3154_,
		_w3160_,
		_w3161_,
		_w3170_
	);
	LUT4 #(
		.INIT('h0080)
	) name1270 (
		\m2_s10_cyc_o_reg/NET0131 ,
		\rf_conf10_reg[4]/NET0131 ,
		\rf_conf10_reg[5]/NET0131 ,
		\s10_msel_arb3_state_reg[0]/NET0131 ,
		_w3171_
	);
	LUT2 #(
		.INIT('h1)
	) name1271 (
		\s10_msel_arb3_state_reg[2]/NET0131 ,
		_w3171_,
		_w3172_
	);
	LUT3 #(
		.INIT('h01)
	) name1272 (
		\s10_msel_arb3_state_reg[2]/NET0131 ,
		_w3163_,
		_w3171_,
		_w3173_
	);
	LUT3 #(
		.INIT('h10)
	) name1273 (
		_w3169_,
		_w3170_,
		_w3173_,
		_w3174_
	);
	LUT2 #(
		.INIT('h8)
	) name1274 (
		\s10_msel_arb3_state_reg[0]/NET0131 ,
		\s10_msel_arb3_state_reg[1]/NET0131 ,
		_w3175_
	);
	LUT4 #(
		.INIT('h7f00)
	) name1275 (
		\m2_s10_cyc_o_reg/NET0131 ,
		\rf_conf10_reg[4]/NET0131 ,
		\rf_conf10_reg[5]/NET0131 ,
		\s10_msel_arb3_state_reg[0]/NET0131 ,
		_w3176_
	);
	LUT3 #(
		.INIT('h10)
	) name1276 (
		_w3163_,
		_w3165_,
		_w3176_,
		_w3177_
	);
	LUT4 #(
		.INIT('h0b0a)
	) name1277 (
		\s10_msel_arb3_state_reg[2]/NET0131 ,
		_w3170_,
		_w3175_,
		_w3177_,
		_w3178_
	);
	LUT2 #(
		.INIT('h8)
	) name1278 (
		\s10_msel_arb3_state_reg[1]/NET0131 ,
		\s10_msel_arb3_state_reg[2]/NET0131 ,
		_w3179_
	);
	LUT3 #(
		.INIT('h80)
	) name1279 (
		\s10_msel_arb3_state_reg[0]/NET0131 ,
		\s10_msel_arb3_state_reg[1]/NET0131 ,
		\s10_msel_arb3_state_reg[2]/NET0131 ,
		_w3180_
	);
	LUT3 #(
		.INIT('he0)
	) name1280 (
		_w3160_,
		_w3167_,
		_w3180_,
		_w3181_
	);
	LUT4 #(
		.INIT('hdddc)
	) name1281 (
		_w3168_,
		_w3174_,
		_w3178_,
		_w3181_,
		_w3182_
	);
	LUT3 #(
		.INIT('h20)
	) name1282 (
		\m5_s11_cyc_o_reg/NET0131 ,
		\rf_conf11_reg[10]/NET0131 ,
		\rf_conf11_reg[11]/NET0131 ,
		_w3183_
	);
	LUT3 #(
		.INIT('h20)
	) name1283 (
		\m4_s11_cyc_o_reg/NET0131 ,
		\rf_conf11_reg[8]/NET0131 ,
		\rf_conf11_reg[9]/NET0131 ,
		_w3184_
	);
	LUT3 #(
		.INIT('h20)
	) name1284 (
		\m6_s11_cyc_o_reg/NET0131 ,
		\rf_conf11_reg[12]/NET0131 ,
		\rf_conf11_reg[13]/NET0131 ,
		_w3185_
	);
	LUT3 #(
		.INIT('h20)
	) name1285 (
		\m7_s11_cyc_o_reg/NET0131 ,
		\rf_conf11_reg[14]/NET0131 ,
		\rf_conf11_reg[15]/NET0131 ,
		_w3186_
	);
	LUT2 #(
		.INIT('h1)
	) name1286 (
		_w3185_,
		_w3186_,
		_w3187_
	);
	LUT4 #(
		.INIT('h0001)
	) name1287 (
		_w3183_,
		_w3184_,
		_w3185_,
		_w3186_,
		_w3188_
	);
	LUT3 #(
		.INIT('h20)
	) name1288 (
		\m3_s11_cyc_o_reg/NET0131 ,
		\rf_conf11_reg[6]/NET0131 ,
		\rf_conf11_reg[7]/NET0131 ,
		_w3189_
	);
	LUT4 #(
		.INIT('h00df)
	) name1289 (
		\m3_s11_cyc_o_reg/NET0131 ,
		\rf_conf11_reg[6]/NET0131 ,
		\rf_conf11_reg[7]/NET0131 ,
		\s11_msel_arb2_state_reg[2]/NET0131 ,
		_w3190_
	);
	LUT3 #(
		.INIT('h20)
	) name1290 (
		\m2_s11_cyc_o_reg/NET0131 ,
		\rf_conf11_reg[4]/NET0131 ,
		\rf_conf11_reg[5]/NET0131 ,
		_w3191_
	);
	LUT4 #(
		.INIT('h0020)
	) name1291 (
		\m0_s11_cyc_o_reg/NET0131 ,
		\rf_conf11_reg[0]/NET0131 ,
		\rf_conf11_reg[1]/NET0131 ,
		\s11_msel_arb2_state_reg[1]/NET0131 ,
		_w3192_
	);
	LUT3 #(
		.INIT('h54)
	) name1292 (
		\s11_msel_arb2_state_reg[0]/NET0131 ,
		_w3191_,
		_w3192_,
		_w3193_
	);
	LUT3 #(
		.INIT('h20)
	) name1293 (
		\m1_s11_cyc_o_reg/NET0131 ,
		\rf_conf11_reg[2]/NET0131 ,
		\rf_conf11_reg[3]/NET0131 ,
		_w3194_
	);
	LUT3 #(
		.INIT('h54)
	) name1294 (
		\s11_msel_arb2_state_reg[1]/NET0131 ,
		_w3191_,
		_w3194_,
		_w3195_
	);
	LUT4 #(
		.INIT('h0004)
	) name1295 (
		_w3188_,
		_w3190_,
		_w3193_,
		_w3195_,
		_w3196_
	);
	LUT2 #(
		.INIT('h1)
	) name1296 (
		_w3189_,
		_w3191_,
		_w3197_
	);
	LUT3 #(
		.INIT('h20)
	) name1297 (
		\m0_s11_cyc_o_reg/NET0131 ,
		\rf_conf11_reg[0]/NET0131 ,
		\rf_conf11_reg[1]/NET0131 ,
		_w3198_
	);
	LUT4 #(
		.INIT('h0001)
	) name1298 (
		_w3189_,
		_w3191_,
		_w3194_,
		_w3198_,
		_w3199_
	);
	LUT4 #(
		.INIT('h0020)
	) name1299 (
		\m4_s11_cyc_o_reg/NET0131 ,
		\rf_conf11_reg[8]/NET0131 ,
		\rf_conf11_reg[9]/NET0131 ,
		\s11_msel_arb2_state_reg[1]/NET0131 ,
		_w3200_
	);
	LUT3 #(
		.INIT('h54)
	) name1300 (
		\s11_msel_arb2_state_reg[0]/NET0131 ,
		_w3185_,
		_w3200_,
		_w3201_
	);
	LUT3 #(
		.INIT('h54)
	) name1301 (
		\s11_msel_arb2_state_reg[1]/NET0131 ,
		_w3183_,
		_w3185_,
		_w3202_
	);
	LUT4 #(
		.INIT('h0001)
	) name1302 (
		_w3186_,
		_w3199_,
		_w3201_,
		_w3202_,
		_w3203_
	);
	LUT3 #(
		.INIT('hce)
	) name1303 (
		\s11_msel_arb2_state_reg[2]/NET0131 ,
		_w3196_,
		_w3203_,
		_w3204_
	);
	LUT2 #(
		.INIT('h4)
	) name1304 (
		\s11_msel_arb3_state_reg[1]/NET0131 ,
		\s11_msel_arb3_state_reg[2]/NET0131 ,
		_w3205_
	);
	LUT3 #(
		.INIT('h80)
	) name1305 (
		\m1_s11_cyc_o_reg/NET0131 ,
		\rf_conf11_reg[2]/NET0131 ,
		\rf_conf11_reg[3]/NET0131 ,
		_w3206_
	);
	LUT3 #(
		.INIT('h80)
	) name1306 (
		\m0_s11_cyc_o_reg/NET0131 ,
		\rf_conf11_reg[0]/NET0131 ,
		\rf_conf11_reg[1]/NET0131 ,
		_w3207_
	);
	LUT3 #(
		.INIT('h80)
	) name1307 (
		\m3_s11_cyc_o_reg/NET0131 ,
		\rf_conf11_reg[6]/NET0131 ,
		\rf_conf11_reg[7]/NET0131 ,
		_w3208_
	);
	LUT3 #(
		.INIT('h80)
	) name1308 (
		\m2_s11_cyc_o_reg/NET0131 ,
		\rf_conf11_reg[4]/NET0131 ,
		\rf_conf11_reg[5]/NET0131 ,
		_w3209_
	);
	LUT4 #(
		.INIT('h0001)
	) name1309 (
		_w3206_,
		_w3207_,
		_w3208_,
		_w3209_,
		_w3210_
	);
	LUT3 #(
		.INIT('h80)
	) name1310 (
		\m5_s11_cyc_o_reg/NET0131 ,
		\rf_conf11_reg[10]/NET0131 ,
		\rf_conf11_reg[11]/NET0131 ,
		_w3211_
	);
	LUT3 #(
		.INIT('h80)
	) name1311 (
		\m7_s11_cyc_o_reg/NET0131 ,
		\rf_conf11_reg[14]/NET0131 ,
		\rf_conf11_reg[15]/NET0131 ,
		_w3212_
	);
	LUT3 #(
		.INIT('h80)
	) name1312 (
		\m6_s11_cyc_o_reg/NET0131 ,
		\rf_conf11_reg[12]/NET0131 ,
		\rf_conf11_reg[13]/NET0131 ,
		_w3213_
	);
	LUT2 #(
		.INIT('h1)
	) name1313 (
		_w3212_,
		_w3213_,
		_w3214_
	);
	LUT3 #(
		.INIT('h01)
	) name1314 (
		_w3211_,
		_w3212_,
		_w3213_,
		_w3215_
	);
	LUT3 #(
		.INIT('h8a)
	) name1315 (
		_w3205_,
		_w3210_,
		_w3215_,
		_w3216_
	);
	LUT2 #(
		.INIT('h8)
	) name1316 (
		\s11_msel_arb3_state_reg[1]/NET0131 ,
		\s11_msel_arb3_state_reg[2]/NET0131 ,
		_w3217_
	);
	LUT3 #(
		.INIT('he0)
	) name1317 (
		_w3210_,
		_w3212_,
		_w3217_,
		_w3218_
	);
	LUT3 #(
		.INIT('h80)
	) name1318 (
		\m4_s11_cyc_o_reg/NET0131 ,
		\rf_conf11_reg[8]/NET0131 ,
		\rf_conf11_reg[9]/NET0131 ,
		_w3219_
	);
	LUT2 #(
		.INIT('h1)
	) name1319 (
		_w3211_,
		_w3219_,
		_w3220_
	);
	LUT4 #(
		.INIT('h0001)
	) name1320 (
		_w3211_,
		_w3212_,
		_w3213_,
		_w3219_,
		_w3221_
	);
	LUT4 #(
		.INIT('h007f)
	) name1321 (
		\m1_s11_cyc_o_reg/NET0131 ,
		\rf_conf11_reg[2]/NET0131 ,
		\rf_conf11_reg[3]/NET0131 ,
		\s11_msel_arb3_state_reg[2]/NET0131 ,
		_w3222_
	);
	LUT4 #(
		.INIT('h007f)
	) name1322 (
		\m2_s11_cyc_o_reg/NET0131 ,
		\rf_conf11_reg[4]/NET0131 ,
		\rf_conf11_reg[5]/NET0131 ,
		\s11_msel_arb3_state_reg[1]/NET0131 ,
		_w3223_
	);
	LUT2 #(
		.INIT('h8)
	) name1323 (
		_w3222_,
		_w3223_,
		_w3224_
	);
	LUT3 #(
		.INIT('h10)
	) name1324 (
		_w3208_,
		_w3221_,
		_w3224_,
		_w3225_
	);
	LUT4 #(
		.INIT('haaa8)
	) name1325 (
		\s11_msel_arb3_state_reg[0]/NET0131 ,
		_w3216_,
		_w3218_,
		_w3225_,
		_w3226_
	);
	LUT4 #(
		.INIT('h0080)
	) name1326 (
		\m2_s11_cyc_o_reg/NET0131 ,
		\rf_conf11_reg[4]/NET0131 ,
		\rf_conf11_reg[5]/NET0131 ,
		\s11_msel_arb3_state_reg[0]/NET0131 ,
		_w3227_
	);
	LUT3 #(
		.INIT('h54)
	) name1327 (
		\s11_msel_arb3_state_reg[1]/NET0131 ,
		_w3206_,
		_w3207_,
		_w3228_
	);
	LUT4 #(
		.INIT('h00ab)
	) name1328 (
		\s11_msel_arb3_state_reg[1]/NET0131 ,
		_w3206_,
		_w3207_,
		_w3227_,
		_w3229_
	);
	LUT4 #(
		.INIT('h5455)
	) name1329 (
		\s11_msel_arb3_state_reg[2]/NET0131 ,
		_w3208_,
		_w3221_,
		_w3229_,
		_w3230_
	);
	LUT2 #(
		.INIT('h2)
	) name1330 (
		\s11_msel_arb3_state_reg[1]/NET0131 ,
		\s11_msel_arb3_state_reg[2]/NET0131 ,
		_w3231_
	);
	LUT3 #(
		.INIT('ha2)
	) name1331 (
		\s11_msel_arb3_state_reg[0]/NET0131 ,
		\s11_msel_arb3_state_reg[1]/NET0131 ,
		\s11_msel_arb3_state_reg[2]/NET0131 ,
		_w3232_
	);
	LUT3 #(
		.INIT('h32)
	) name1332 (
		_w3211_,
		_w3217_,
		_w3219_,
		_w3233_
	);
	LUT4 #(
		.INIT('h0f0b)
	) name1333 (
		_w3210_,
		_w3214_,
		_w3232_,
		_w3233_,
		_w3234_
	);
	LUT2 #(
		.INIT('h4)
	) name1334 (
		_w3230_,
		_w3234_,
		_w3235_
	);
	LUT2 #(
		.INIT('he)
	) name1335 (
		_w3226_,
		_w3235_,
		_w3236_
	);
	LUT3 #(
		.INIT('h80)
	) name1336 (
		\m5_s12_cyc_o_reg/NET0131 ,
		\rf_conf12_reg[10]/NET0131 ,
		\rf_conf12_reg[11]/NET0131 ,
		_w3237_
	);
	LUT3 #(
		.INIT('h80)
	) name1337 (
		\m4_s12_cyc_o_reg/NET0131 ,
		\rf_conf12_reg[8]/NET0131 ,
		\rf_conf12_reg[9]/NET0131 ,
		_w3238_
	);
	LUT3 #(
		.INIT('h01)
	) name1338 (
		\s12_msel_arb3_state_reg[0]/NET0131 ,
		_w3237_,
		_w3238_,
		_w3239_
	);
	LUT2 #(
		.INIT('h8)
	) name1339 (
		\s12_msel_arb3_state_reg[0]/NET0131 ,
		\s12_msel_arb3_state_reg[2]/NET0131 ,
		_w3240_
	);
	LUT3 #(
		.INIT('h13)
	) name1340 (
		\s12_msel_arb3_state_reg[0]/NET0131 ,
		\s12_msel_arb3_state_reg[1]/NET0131 ,
		\s12_msel_arb3_state_reg[2]/NET0131 ,
		_w3241_
	);
	LUT4 #(
		.INIT('h0080)
	) name1341 (
		\m5_s12_cyc_o_reg/NET0131 ,
		\rf_conf12_reg[10]/NET0131 ,
		\rf_conf12_reg[11]/NET0131 ,
		\s12_msel_arb3_state_reg[1]/NET0131 ,
		_w3242_
	);
	LUT2 #(
		.INIT('h1)
	) name1342 (
		_w3241_,
		_w3242_,
		_w3243_
	);
	LUT3 #(
		.INIT('h80)
	) name1343 (
		\m7_s12_cyc_o_reg/NET0131 ,
		\rf_conf12_reg[14]/NET0131 ,
		\rf_conf12_reg[15]/NET0131 ,
		_w3244_
	);
	LUT3 #(
		.INIT('h80)
	) name1344 (
		\m6_s12_cyc_o_reg/NET0131 ,
		\rf_conf12_reg[12]/NET0131 ,
		\rf_conf12_reg[13]/NET0131 ,
		_w3245_
	);
	LUT2 #(
		.INIT('h1)
	) name1345 (
		_w3244_,
		_w3245_,
		_w3246_
	);
	LUT3 #(
		.INIT('h80)
	) name1346 (
		\m3_s12_cyc_o_reg/NET0131 ,
		\rf_conf12_reg[6]/NET0131 ,
		\rf_conf12_reg[7]/NET0131 ,
		_w3247_
	);
	LUT3 #(
		.INIT('h80)
	) name1347 (
		\m2_s12_cyc_o_reg/NET0131 ,
		\rf_conf12_reg[4]/NET0131 ,
		\rf_conf12_reg[5]/NET0131 ,
		_w3248_
	);
	LUT3 #(
		.INIT('h80)
	) name1348 (
		\m1_s12_cyc_o_reg/NET0131 ,
		\rf_conf12_reg[2]/NET0131 ,
		\rf_conf12_reg[3]/NET0131 ,
		_w3249_
	);
	LUT3 #(
		.INIT('h80)
	) name1349 (
		\m0_s12_cyc_o_reg/NET0131 ,
		\rf_conf12_reg[0]/NET0131 ,
		\rf_conf12_reg[1]/NET0131 ,
		_w3250_
	);
	LUT4 #(
		.INIT('h0001)
	) name1350 (
		_w3247_,
		_w3248_,
		_w3249_,
		_w3250_,
		_w3251_
	);
	LUT4 #(
		.INIT('h00e0)
	) name1351 (
		_w3239_,
		_w3243_,
		_w3246_,
		_w3251_,
		_w3252_
	);
	LUT4 #(
		.INIT('h3332)
	) name1352 (
		\s12_msel_arb3_state_reg[0]/NET0131 ,
		\s12_msel_arb3_state_reg[1]/NET0131 ,
		_w3249_,
		_w3250_,
		_w3253_
	);
	LUT4 #(
		.INIT('h0001)
	) name1353 (
		_w3237_,
		_w3238_,
		_w3244_,
		_w3245_,
		_w3254_
	);
	LUT4 #(
		.INIT('h0080)
	) name1354 (
		\m2_s12_cyc_o_reg/NET0131 ,
		\rf_conf12_reg[4]/NET0131 ,
		\rf_conf12_reg[5]/NET0131 ,
		\s12_msel_arb3_state_reg[0]/NET0131 ,
		_w3255_
	);
	LUT2 #(
		.INIT('h1)
	) name1355 (
		\s12_msel_arb3_state_reg[2]/NET0131 ,
		_w3255_,
		_w3256_
	);
	LUT3 #(
		.INIT('h01)
	) name1356 (
		\s12_msel_arb3_state_reg[2]/NET0131 ,
		_w3247_,
		_w3255_,
		_w3257_
	);
	LUT3 #(
		.INIT('h10)
	) name1357 (
		_w3253_,
		_w3254_,
		_w3257_,
		_w3258_
	);
	LUT2 #(
		.INIT('h8)
	) name1358 (
		\s12_msel_arb3_state_reg[0]/NET0131 ,
		\s12_msel_arb3_state_reg[1]/NET0131 ,
		_w3259_
	);
	LUT4 #(
		.INIT('h7f00)
	) name1359 (
		\m2_s12_cyc_o_reg/NET0131 ,
		\rf_conf12_reg[4]/NET0131 ,
		\rf_conf12_reg[5]/NET0131 ,
		\s12_msel_arb3_state_reg[0]/NET0131 ,
		_w3260_
	);
	LUT3 #(
		.INIT('h10)
	) name1360 (
		_w3247_,
		_w3249_,
		_w3260_,
		_w3261_
	);
	LUT4 #(
		.INIT('h0b0a)
	) name1361 (
		\s12_msel_arb3_state_reg[2]/NET0131 ,
		_w3254_,
		_w3259_,
		_w3261_,
		_w3262_
	);
	LUT2 #(
		.INIT('h8)
	) name1362 (
		\s12_msel_arb3_state_reg[1]/NET0131 ,
		\s12_msel_arb3_state_reg[2]/NET0131 ,
		_w3263_
	);
	LUT3 #(
		.INIT('h80)
	) name1363 (
		\s12_msel_arb3_state_reg[0]/NET0131 ,
		\s12_msel_arb3_state_reg[1]/NET0131 ,
		\s12_msel_arb3_state_reg[2]/NET0131 ,
		_w3264_
	);
	LUT3 #(
		.INIT('he0)
	) name1364 (
		_w3244_,
		_w3251_,
		_w3264_,
		_w3265_
	);
	LUT4 #(
		.INIT('hdddc)
	) name1365 (
		_w3252_,
		_w3258_,
		_w3262_,
		_w3265_,
		_w3266_
	);
	LUT2 #(
		.INIT('h4)
	) name1366 (
		\s14_msel_arb3_state_reg[1]/NET0131 ,
		\s14_msel_arb3_state_reg[2]/NET0131 ,
		_w3267_
	);
	LUT3 #(
		.INIT('h80)
	) name1367 (
		\m1_s14_cyc_o_reg/NET0131 ,
		\rf_conf14_reg[2]/NET0131 ,
		\rf_conf14_reg[3]/NET0131 ,
		_w3268_
	);
	LUT3 #(
		.INIT('h80)
	) name1368 (
		\m0_s14_cyc_o_reg/NET0131 ,
		\rf_conf14_reg[0]/NET0131 ,
		\rf_conf14_reg[1]/NET0131 ,
		_w3269_
	);
	LUT3 #(
		.INIT('h80)
	) name1369 (
		\m3_s14_cyc_o_reg/NET0131 ,
		\rf_conf14_reg[6]/NET0131 ,
		\rf_conf14_reg[7]/NET0131 ,
		_w3270_
	);
	LUT3 #(
		.INIT('h80)
	) name1370 (
		\m2_s14_cyc_o_reg/NET0131 ,
		\rf_conf14_reg[4]/NET0131 ,
		\rf_conf14_reg[5]/NET0131 ,
		_w3271_
	);
	LUT4 #(
		.INIT('h0001)
	) name1371 (
		_w3268_,
		_w3269_,
		_w3270_,
		_w3271_,
		_w3272_
	);
	LUT3 #(
		.INIT('h80)
	) name1372 (
		\m5_s14_cyc_o_reg/NET0131 ,
		\rf_conf14_reg[10]/NET0131 ,
		\rf_conf14_reg[11]/NET0131 ,
		_w3273_
	);
	LUT3 #(
		.INIT('h80)
	) name1373 (
		\m7_s14_cyc_o_reg/NET0131 ,
		\rf_conf14_reg[14]/NET0131 ,
		\rf_conf14_reg[15]/NET0131 ,
		_w3274_
	);
	LUT3 #(
		.INIT('h80)
	) name1374 (
		\m6_s14_cyc_o_reg/NET0131 ,
		\rf_conf14_reg[12]/NET0131 ,
		\rf_conf14_reg[13]/NET0131 ,
		_w3275_
	);
	LUT2 #(
		.INIT('h1)
	) name1375 (
		_w3274_,
		_w3275_,
		_w3276_
	);
	LUT3 #(
		.INIT('h01)
	) name1376 (
		_w3273_,
		_w3274_,
		_w3275_,
		_w3277_
	);
	LUT3 #(
		.INIT('h8a)
	) name1377 (
		_w3267_,
		_w3272_,
		_w3277_,
		_w3278_
	);
	LUT2 #(
		.INIT('h8)
	) name1378 (
		\s14_msel_arb3_state_reg[1]/NET0131 ,
		\s14_msel_arb3_state_reg[2]/NET0131 ,
		_w3279_
	);
	LUT3 #(
		.INIT('he0)
	) name1379 (
		_w3272_,
		_w3274_,
		_w3279_,
		_w3280_
	);
	LUT3 #(
		.INIT('h80)
	) name1380 (
		\m4_s14_cyc_o_reg/NET0131 ,
		\rf_conf14_reg[8]/NET0131 ,
		\rf_conf14_reg[9]/NET0131 ,
		_w3281_
	);
	LUT2 #(
		.INIT('h1)
	) name1381 (
		_w3273_,
		_w3281_,
		_w3282_
	);
	LUT4 #(
		.INIT('h0001)
	) name1382 (
		_w3273_,
		_w3274_,
		_w3275_,
		_w3281_,
		_w3283_
	);
	LUT4 #(
		.INIT('h007f)
	) name1383 (
		\m1_s14_cyc_o_reg/NET0131 ,
		\rf_conf14_reg[2]/NET0131 ,
		\rf_conf14_reg[3]/NET0131 ,
		\s14_msel_arb3_state_reg[2]/NET0131 ,
		_w3284_
	);
	LUT4 #(
		.INIT('h007f)
	) name1384 (
		\m2_s14_cyc_o_reg/NET0131 ,
		\rf_conf14_reg[4]/NET0131 ,
		\rf_conf14_reg[5]/NET0131 ,
		\s14_msel_arb3_state_reg[1]/NET0131 ,
		_w3285_
	);
	LUT2 #(
		.INIT('h8)
	) name1385 (
		_w3284_,
		_w3285_,
		_w3286_
	);
	LUT3 #(
		.INIT('h10)
	) name1386 (
		_w3270_,
		_w3283_,
		_w3286_,
		_w3287_
	);
	LUT4 #(
		.INIT('haaa8)
	) name1387 (
		\s14_msel_arb3_state_reg[0]/NET0131 ,
		_w3278_,
		_w3280_,
		_w3287_,
		_w3288_
	);
	LUT4 #(
		.INIT('h0080)
	) name1388 (
		\m2_s14_cyc_o_reg/NET0131 ,
		\rf_conf14_reg[4]/NET0131 ,
		\rf_conf14_reg[5]/NET0131 ,
		\s14_msel_arb3_state_reg[0]/NET0131 ,
		_w3289_
	);
	LUT3 #(
		.INIT('h54)
	) name1389 (
		\s14_msel_arb3_state_reg[1]/NET0131 ,
		_w3268_,
		_w3269_,
		_w3290_
	);
	LUT4 #(
		.INIT('h00ab)
	) name1390 (
		\s14_msel_arb3_state_reg[1]/NET0131 ,
		_w3268_,
		_w3269_,
		_w3289_,
		_w3291_
	);
	LUT4 #(
		.INIT('h5455)
	) name1391 (
		\s14_msel_arb3_state_reg[2]/NET0131 ,
		_w3270_,
		_w3283_,
		_w3291_,
		_w3292_
	);
	LUT2 #(
		.INIT('h2)
	) name1392 (
		\s14_msel_arb3_state_reg[1]/NET0131 ,
		\s14_msel_arb3_state_reg[2]/NET0131 ,
		_w3293_
	);
	LUT3 #(
		.INIT('ha2)
	) name1393 (
		\s14_msel_arb3_state_reg[0]/NET0131 ,
		\s14_msel_arb3_state_reg[1]/NET0131 ,
		\s14_msel_arb3_state_reg[2]/NET0131 ,
		_w3294_
	);
	LUT3 #(
		.INIT('h32)
	) name1394 (
		_w3273_,
		_w3279_,
		_w3281_,
		_w3295_
	);
	LUT4 #(
		.INIT('h0f0b)
	) name1395 (
		_w3272_,
		_w3276_,
		_w3294_,
		_w3295_,
		_w3296_
	);
	LUT2 #(
		.INIT('h4)
	) name1396 (
		_w3292_,
		_w3296_,
		_w3297_
	);
	LUT2 #(
		.INIT('he)
	) name1397 (
		_w3288_,
		_w3297_,
		_w3298_
	);
	LUT3 #(
		.INIT('h20)
	) name1398 (
		\m5_s1_cyc_o_reg/NET0131 ,
		\rf_conf1_reg[10]/NET0131 ,
		\rf_conf1_reg[11]/NET0131 ,
		_w3299_
	);
	LUT3 #(
		.INIT('h20)
	) name1399 (
		\m4_s1_cyc_o_reg/NET0131 ,
		\rf_conf1_reg[8]/NET0131 ,
		\rf_conf1_reg[9]/NET0131 ,
		_w3300_
	);
	LUT3 #(
		.INIT('h20)
	) name1400 (
		\m6_s1_cyc_o_reg/NET0131 ,
		\rf_conf1_reg[12]/NET0131 ,
		\rf_conf1_reg[13]/NET0131 ,
		_w3301_
	);
	LUT3 #(
		.INIT('h20)
	) name1401 (
		\m7_s1_cyc_o_reg/NET0131 ,
		\rf_conf1_reg[14]/NET0131 ,
		\rf_conf1_reg[15]/NET0131 ,
		_w3302_
	);
	LUT2 #(
		.INIT('h1)
	) name1402 (
		_w3301_,
		_w3302_,
		_w3303_
	);
	LUT4 #(
		.INIT('h0001)
	) name1403 (
		_w3299_,
		_w3300_,
		_w3301_,
		_w3302_,
		_w3304_
	);
	LUT3 #(
		.INIT('h20)
	) name1404 (
		\m3_s1_cyc_o_reg/NET0131 ,
		\rf_conf1_reg[6]/NET0131 ,
		\rf_conf1_reg[7]/NET0131 ,
		_w3305_
	);
	LUT4 #(
		.INIT('h00df)
	) name1405 (
		\m3_s1_cyc_o_reg/NET0131 ,
		\rf_conf1_reg[6]/NET0131 ,
		\rf_conf1_reg[7]/NET0131 ,
		\s1_msel_arb2_state_reg[2]/NET0131 ,
		_w3306_
	);
	LUT3 #(
		.INIT('h20)
	) name1406 (
		\m2_s1_cyc_o_reg/NET0131 ,
		\rf_conf1_reg[4]/NET0131 ,
		\rf_conf1_reg[5]/NET0131 ,
		_w3307_
	);
	LUT4 #(
		.INIT('h0020)
	) name1407 (
		\m0_s1_cyc_o_reg/NET0131 ,
		\rf_conf1_reg[0]/NET0131 ,
		\rf_conf1_reg[1]/NET0131 ,
		\s1_msel_arb2_state_reg[1]/NET0131 ,
		_w3308_
	);
	LUT3 #(
		.INIT('h54)
	) name1408 (
		\s1_msel_arb2_state_reg[0]/NET0131 ,
		_w3307_,
		_w3308_,
		_w3309_
	);
	LUT3 #(
		.INIT('h20)
	) name1409 (
		\m1_s1_cyc_o_reg/NET0131 ,
		\rf_conf1_reg[2]/NET0131 ,
		\rf_conf1_reg[3]/NET0131 ,
		_w3310_
	);
	LUT3 #(
		.INIT('h54)
	) name1410 (
		\s1_msel_arb2_state_reg[1]/NET0131 ,
		_w3307_,
		_w3310_,
		_w3311_
	);
	LUT4 #(
		.INIT('h0004)
	) name1411 (
		_w3304_,
		_w3306_,
		_w3309_,
		_w3311_,
		_w3312_
	);
	LUT2 #(
		.INIT('h1)
	) name1412 (
		_w3305_,
		_w3307_,
		_w3313_
	);
	LUT3 #(
		.INIT('h20)
	) name1413 (
		\m0_s1_cyc_o_reg/NET0131 ,
		\rf_conf1_reg[0]/NET0131 ,
		\rf_conf1_reg[1]/NET0131 ,
		_w3314_
	);
	LUT4 #(
		.INIT('h0001)
	) name1414 (
		_w3305_,
		_w3307_,
		_w3310_,
		_w3314_,
		_w3315_
	);
	LUT4 #(
		.INIT('h0020)
	) name1415 (
		\m4_s1_cyc_o_reg/NET0131 ,
		\rf_conf1_reg[8]/NET0131 ,
		\rf_conf1_reg[9]/NET0131 ,
		\s1_msel_arb2_state_reg[1]/NET0131 ,
		_w3316_
	);
	LUT3 #(
		.INIT('h54)
	) name1416 (
		\s1_msel_arb2_state_reg[0]/NET0131 ,
		_w3301_,
		_w3316_,
		_w3317_
	);
	LUT3 #(
		.INIT('h54)
	) name1417 (
		\s1_msel_arb2_state_reg[1]/NET0131 ,
		_w3299_,
		_w3301_,
		_w3318_
	);
	LUT4 #(
		.INIT('h0001)
	) name1418 (
		_w3302_,
		_w3315_,
		_w3317_,
		_w3318_,
		_w3319_
	);
	LUT3 #(
		.INIT('hce)
	) name1419 (
		\s1_msel_arb2_state_reg[2]/NET0131 ,
		_w3312_,
		_w3319_,
		_w3320_
	);
	LUT2 #(
		.INIT('h4)
	) name1420 (
		\s1_msel_arb3_state_reg[1]/NET0131 ,
		\s1_msel_arb3_state_reg[2]/NET0131 ,
		_w3321_
	);
	LUT3 #(
		.INIT('h80)
	) name1421 (
		\m1_s1_cyc_o_reg/NET0131 ,
		\rf_conf1_reg[2]/NET0131 ,
		\rf_conf1_reg[3]/NET0131 ,
		_w3322_
	);
	LUT3 #(
		.INIT('h80)
	) name1422 (
		\m0_s1_cyc_o_reg/NET0131 ,
		\rf_conf1_reg[0]/NET0131 ,
		\rf_conf1_reg[1]/NET0131 ,
		_w3323_
	);
	LUT3 #(
		.INIT('h80)
	) name1423 (
		\m3_s1_cyc_o_reg/NET0131 ,
		\rf_conf1_reg[6]/NET0131 ,
		\rf_conf1_reg[7]/NET0131 ,
		_w3324_
	);
	LUT3 #(
		.INIT('h80)
	) name1424 (
		\m2_s1_cyc_o_reg/NET0131 ,
		\rf_conf1_reg[4]/NET0131 ,
		\rf_conf1_reg[5]/NET0131 ,
		_w3325_
	);
	LUT4 #(
		.INIT('h0001)
	) name1425 (
		_w3322_,
		_w3323_,
		_w3324_,
		_w3325_,
		_w3326_
	);
	LUT3 #(
		.INIT('h80)
	) name1426 (
		\m5_s1_cyc_o_reg/NET0131 ,
		\rf_conf1_reg[10]/NET0131 ,
		\rf_conf1_reg[11]/NET0131 ,
		_w3327_
	);
	LUT3 #(
		.INIT('h80)
	) name1427 (
		\m7_s1_cyc_o_reg/NET0131 ,
		\rf_conf1_reg[14]/NET0131 ,
		\rf_conf1_reg[15]/NET0131 ,
		_w3328_
	);
	LUT3 #(
		.INIT('h80)
	) name1428 (
		\m6_s1_cyc_o_reg/NET0131 ,
		\rf_conf1_reg[12]/NET0131 ,
		\rf_conf1_reg[13]/NET0131 ,
		_w3329_
	);
	LUT2 #(
		.INIT('h1)
	) name1429 (
		_w3328_,
		_w3329_,
		_w3330_
	);
	LUT3 #(
		.INIT('h01)
	) name1430 (
		_w3327_,
		_w3328_,
		_w3329_,
		_w3331_
	);
	LUT3 #(
		.INIT('h8a)
	) name1431 (
		_w3321_,
		_w3326_,
		_w3331_,
		_w3332_
	);
	LUT2 #(
		.INIT('h8)
	) name1432 (
		\s1_msel_arb3_state_reg[1]/NET0131 ,
		\s1_msel_arb3_state_reg[2]/NET0131 ,
		_w3333_
	);
	LUT3 #(
		.INIT('he0)
	) name1433 (
		_w3326_,
		_w3328_,
		_w3333_,
		_w3334_
	);
	LUT3 #(
		.INIT('h80)
	) name1434 (
		\m4_s1_cyc_o_reg/NET0131 ,
		\rf_conf1_reg[8]/NET0131 ,
		\rf_conf1_reg[9]/NET0131 ,
		_w3335_
	);
	LUT2 #(
		.INIT('h1)
	) name1435 (
		_w3327_,
		_w3335_,
		_w3336_
	);
	LUT4 #(
		.INIT('h0001)
	) name1436 (
		_w3327_,
		_w3328_,
		_w3329_,
		_w3335_,
		_w3337_
	);
	LUT4 #(
		.INIT('h007f)
	) name1437 (
		\m1_s1_cyc_o_reg/NET0131 ,
		\rf_conf1_reg[2]/NET0131 ,
		\rf_conf1_reg[3]/NET0131 ,
		\s1_msel_arb3_state_reg[2]/NET0131 ,
		_w3338_
	);
	LUT4 #(
		.INIT('h007f)
	) name1438 (
		\m2_s1_cyc_o_reg/NET0131 ,
		\rf_conf1_reg[4]/NET0131 ,
		\rf_conf1_reg[5]/NET0131 ,
		\s1_msel_arb3_state_reg[1]/NET0131 ,
		_w3339_
	);
	LUT2 #(
		.INIT('h8)
	) name1439 (
		_w3338_,
		_w3339_,
		_w3340_
	);
	LUT3 #(
		.INIT('h10)
	) name1440 (
		_w3324_,
		_w3337_,
		_w3340_,
		_w3341_
	);
	LUT4 #(
		.INIT('haaa8)
	) name1441 (
		\s1_msel_arb3_state_reg[0]/NET0131 ,
		_w3332_,
		_w3334_,
		_w3341_,
		_w3342_
	);
	LUT4 #(
		.INIT('h0080)
	) name1442 (
		\m2_s1_cyc_o_reg/NET0131 ,
		\rf_conf1_reg[4]/NET0131 ,
		\rf_conf1_reg[5]/NET0131 ,
		\s1_msel_arb3_state_reg[0]/NET0131 ,
		_w3343_
	);
	LUT3 #(
		.INIT('h54)
	) name1443 (
		\s1_msel_arb3_state_reg[1]/NET0131 ,
		_w3322_,
		_w3323_,
		_w3344_
	);
	LUT4 #(
		.INIT('h00ab)
	) name1444 (
		\s1_msel_arb3_state_reg[1]/NET0131 ,
		_w3322_,
		_w3323_,
		_w3343_,
		_w3345_
	);
	LUT4 #(
		.INIT('h5455)
	) name1445 (
		\s1_msel_arb3_state_reg[2]/NET0131 ,
		_w3324_,
		_w3337_,
		_w3345_,
		_w3346_
	);
	LUT2 #(
		.INIT('h2)
	) name1446 (
		\s1_msel_arb3_state_reg[1]/NET0131 ,
		\s1_msel_arb3_state_reg[2]/NET0131 ,
		_w3347_
	);
	LUT3 #(
		.INIT('ha2)
	) name1447 (
		\s1_msel_arb3_state_reg[0]/NET0131 ,
		\s1_msel_arb3_state_reg[1]/NET0131 ,
		\s1_msel_arb3_state_reg[2]/NET0131 ,
		_w3348_
	);
	LUT3 #(
		.INIT('h32)
	) name1448 (
		_w3327_,
		_w3333_,
		_w3335_,
		_w3349_
	);
	LUT4 #(
		.INIT('h0f0b)
	) name1449 (
		_w3326_,
		_w3330_,
		_w3348_,
		_w3349_,
		_w3350_
	);
	LUT2 #(
		.INIT('h4)
	) name1450 (
		_w3346_,
		_w3350_,
		_w3351_
	);
	LUT2 #(
		.INIT('he)
	) name1451 (
		_w3342_,
		_w3351_,
		_w3352_
	);
	LUT2 #(
		.INIT('h4)
	) name1452 (
		\s3_msel_arb3_state_reg[1]/NET0131 ,
		\s3_msel_arb3_state_reg[2]/NET0131 ,
		_w3353_
	);
	LUT3 #(
		.INIT('h80)
	) name1453 (
		\m1_s3_cyc_o_reg/NET0131 ,
		\rf_conf3_reg[2]/NET0131 ,
		\rf_conf3_reg[3]/NET0131 ,
		_w3354_
	);
	LUT3 #(
		.INIT('h80)
	) name1454 (
		\m0_s3_cyc_o_reg/NET0131 ,
		\rf_conf3_reg[0]/NET0131 ,
		\rf_conf3_reg[1]/NET0131 ,
		_w3355_
	);
	LUT3 #(
		.INIT('h80)
	) name1455 (
		\m3_s3_cyc_o_reg/NET0131 ,
		\rf_conf3_reg[6]/NET0131 ,
		\rf_conf3_reg[7]/NET0131 ,
		_w3356_
	);
	LUT3 #(
		.INIT('h80)
	) name1456 (
		\m2_s3_cyc_o_reg/NET0131 ,
		\rf_conf3_reg[4]/NET0131 ,
		\rf_conf3_reg[5]/NET0131 ,
		_w3357_
	);
	LUT4 #(
		.INIT('h0001)
	) name1457 (
		_w3354_,
		_w3355_,
		_w3356_,
		_w3357_,
		_w3358_
	);
	LUT3 #(
		.INIT('h80)
	) name1458 (
		\m5_s3_cyc_o_reg/NET0131 ,
		\rf_conf3_reg[10]/NET0131 ,
		\rf_conf3_reg[11]/NET0131 ,
		_w3359_
	);
	LUT3 #(
		.INIT('h80)
	) name1459 (
		\m7_s3_cyc_o_reg/NET0131 ,
		\rf_conf3_reg[14]/NET0131 ,
		\rf_conf3_reg[15]/NET0131 ,
		_w3360_
	);
	LUT3 #(
		.INIT('h80)
	) name1460 (
		\m6_s3_cyc_o_reg/NET0131 ,
		\rf_conf3_reg[12]/NET0131 ,
		\rf_conf3_reg[13]/NET0131 ,
		_w3361_
	);
	LUT2 #(
		.INIT('h1)
	) name1461 (
		_w3360_,
		_w3361_,
		_w3362_
	);
	LUT3 #(
		.INIT('h01)
	) name1462 (
		_w3359_,
		_w3360_,
		_w3361_,
		_w3363_
	);
	LUT3 #(
		.INIT('h8a)
	) name1463 (
		_w3353_,
		_w3358_,
		_w3363_,
		_w3364_
	);
	LUT2 #(
		.INIT('h8)
	) name1464 (
		\s3_msel_arb3_state_reg[1]/NET0131 ,
		\s3_msel_arb3_state_reg[2]/NET0131 ,
		_w3365_
	);
	LUT3 #(
		.INIT('he0)
	) name1465 (
		_w3358_,
		_w3360_,
		_w3365_,
		_w3366_
	);
	LUT3 #(
		.INIT('h80)
	) name1466 (
		\m4_s3_cyc_o_reg/NET0131 ,
		\rf_conf3_reg[8]/NET0131 ,
		\rf_conf3_reg[9]/NET0131 ,
		_w3367_
	);
	LUT2 #(
		.INIT('h1)
	) name1467 (
		_w3359_,
		_w3367_,
		_w3368_
	);
	LUT4 #(
		.INIT('h0001)
	) name1468 (
		_w3359_,
		_w3360_,
		_w3361_,
		_w3367_,
		_w3369_
	);
	LUT4 #(
		.INIT('h007f)
	) name1469 (
		\m1_s3_cyc_o_reg/NET0131 ,
		\rf_conf3_reg[2]/NET0131 ,
		\rf_conf3_reg[3]/NET0131 ,
		\s3_msel_arb3_state_reg[2]/NET0131 ,
		_w3370_
	);
	LUT4 #(
		.INIT('h007f)
	) name1470 (
		\m2_s3_cyc_o_reg/NET0131 ,
		\rf_conf3_reg[4]/NET0131 ,
		\rf_conf3_reg[5]/NET0131 ,
		\s3_msel_arb3_state_reg[1]/NET0131 ,
		_w3371_
	);
	LUT2 #(
		.INIT('h8)
	) name1471 (
		_w3370_,
		_w3371_,
		_w3372_
	);
	LUT3 #(
		.INIT('h10)
	) name1472 (
		_w3356_,
		_w3369_,
		_w3372_,
		_w3373_
	);
	LUT4 #(
		.INIT('haaa8)
	) name1473 (
		\s3_msel_arb3_state_reg[0]/NET0131 ,
		_w3364_,
		_w3366_,
		_w3373_,
		_w3374_
	);
	LUT4 #(
		.INIT('h0080)
	) name1474 (
		\m2_s3_cyc_o_reg/NET0131 ,
		\rf_conf3_reg[4]/NET0131 ,
		\rf_conf3_reg[5]/NET0131 ,
		\s3_msel_arb3_state_reg[0]/NET0131 ,
		_w3375_
	);
	LUT3 #(
		.INIT('h54)
	) name1475 (
		\s3_msel_arb3_state_reg[1]/NET0131 ,
		_w3354_,
		_w3355_,
		_w3376_
	);
	LUT4 #(
		.INIT('h00ab)
	) name1476 (
		\s3_msel_arb3_state_reg[1]/NET0131 ,
		_w3354_,
		_w3355_,
		_w3375_,
		_w3377_
	);
	LUT4 #(
		.INIT('h5455)
	) name1477 (
		\s3_msel_arb3_state_reg[2]/NET0131 ,
		_w3356_,
		_w3369_,
		_w3377_,
		_w3378_
	);
	LUT2 #(
		.INIT('h2)
	) name1478 (
		\s3_msel_arb3_state_reg[1]/NET0131 ,
		\s3_msel_arb3_state_reg[2]/NET0131 ,
		_w3379_
	);
	LUT3 #(
		.INIT('ha2)
	) name1479 (
		\s3_msel_arb3_state_reg[0]/NET0131 ,
		\s3_msel_arb3_state_reg[1]/NET0131 ,
		\s3_msel_arb3_state_reg[2]/NET0131 ,
		_w3380_
	);
	LUT3 #(
		.INIT('h32)
	) name1480 (
		_w3359_,
		_w3365_,
		_w3367_,
		_w3381_
	);
	LUT4 #(
		.INIT('h0f0b)
	) name1481 (
		_w3358_,
		_w3362_,
		_w3380_,
		_w3381_,
		_w3382_
	);
	LUT2 #(
		.INIT('h4)
	) name1482 (
		_w3378_,
		_w3382_,
		_w3383_
	);
	LUT2 #(
		.INIT('he)
	) name1483 (
		_w3374_,
		_w3383_,
		_w3384_
	);
	LUT3 #(
		.INIT('h20)
	) name1484 (
		\m5_s5_cyc_o_reg/NET0131 ,
		\rf_conf5_reg[10]/NET0131 ,
		\rf_conf5_reg[11]/NET0131 ,
		_w3385_
	);
	LUT3 #(
		.INIT('h20)
	) name1485 (
		\m4_s5_cyc_o_reg/NET0131 ,
		\rf_conf5_reg[8]/NET0131 ,
		\rf_conf5_reg[9]/NET0131 ,
		_w3386_
	);
	LUT3 #(
		.INIT('h20)
	) name1486 (
		\m6_s5_cyc_o_reg/NET0131 ,
		\rf_conf5_reg[12]/NET0131 ,
		\rf_conf5_reg[13]/NET0131 ,
		_w3387_
	);
	LUT3 #(
		.INIT('h20)
	) name1487 (
		\m7_s5_cyc_o_reg/NET0131 ,
		\rf_conf5_reg[14]/NET0131 ,
		\rf_conf5_reg[15]/NET0131 ,
		_w3388_
	);
	LUT2 #(
		.INIT('h1)
	) name1488 (
		_w3387_,
		_w3388_,
		_w3389_
	);
	LUT4 #(
		.INIT('h0001)
	) name1489 (
		_w3385_,
		_w3386_,
		_w3387_,
		_w3388_,
		_w3390_
	);
	LUT3 #(
		.INIT('h20)
	) name1490 (
		\m3_s5_cyc_o_reg/NET0131 ,
		\rf_conf5_reg[6]/NET0131 ,
		\rf_conf5_reg[7]/NET0131 ,
		_w3391_
	);
	LUT4 #(
		.INIT('h00df)
	) name1491 (
		\m3_s5_cyc_o_reg/NET0131 ,
		\rf_conf5_reg[6]/NET0131 ,
		\rf_conf5_reg[7]/NET0131 ,
		\s5_msel_arb2_state_reg[2]/NET0131 ,
		_w3392_
	);
	LUT3 #(
		.INIT('h20)
	) name1492 (
		\m2_s5_cyc_o_reg/NET0131 ,
		\rf_conf5_reg[4]/NET0131 ,
		\rf_conf5_reg[5]/NET0131 ,
		_w3393_
	);
	LUT4 #(
		.INIT('h0020)
	) name1493 (
		\m0_s5_cyc_o_reg/NET0131 ,
		\rf_conf5_reg[0]/NET0131 ,
		\rf_conf5_reg[1]/NET0131 ,
		\s5_msel_arb2_state_reg[1]/NET0131 ,
		_w3394_
	);
	LUT3 #(
		.INIT('h54)
	) name1494 (
		\s5_msel_arb2_state_reg[0]/NET0131 ,
		_w3393_,
		_w3394_,
		_w3395_
	);
	LUT3 #(
		.INIT('h20)
	) name1495 (
		\m1_s5_cyc_o_reg/NET0131 ,
		\rf_conf5_reg[2]/NET0131 ,
		\rf_conf5_reg[3]/NET0131 ,
		_w3396_
	);
	LUT3 #(
		.INIT('h54)
	) name1496 (
		\s5_msel_arb2_state_reg[1]/NET0131 ,
		_w3393_,
		_w3396_,
		_w3397_
	);
	LUT4 #(
		.INIT('h0004)
	) name1497 (
		_w3390_,
		_w3392_,
		_w3395_,
		_w3397_,
		_w3398_
	);
	LUT2 #(
		.INIT('h1)
	) name1498 (
		_w3391_,
		_w3393_,
		_w3399_
	);
	LUT3 #(
		.INIT('h20)
	) name1499 (
		\m0_s5_cyc_o_reg/NET0131 ,
		\rf_conf5_reg[0]/NET0131 ,
		\rf_conf5_reg[1]/NET0131 ,
		_w3400_
	);
	LUT4 #(
		.INIT('h0001)
	) name1500 (
		_w3391_,
		_w3393_,
		_w3396_,
		_w3400_,
		_w3401_
	);
	LUT4 #(
		.INIT('h0020)
	) name1501 (
		\m4_s5_cyc_o_reg/NET0131 ,
		\rf_conf5_reg[8]/NET0131 ,
		\rf_conf5_reg[9]/NET0131 ,
		\s5_msel_arb2_state_reg[1]/NET0131 ,
		_w3402_
	);
	LUT3 #(
		.INIT('h54)
	) name1502 (
		\s5_msel_arb2_state_reg[0]/NET0131 ,
		_w3387_,
		_w3402_,
		_w3403_
	);
	LUT3 #(
		.INIT('h54)
	) name1503 (
		\s5_msel_arb2_state_reg[1]/NET0131 ,
		_w3385_,
		_w3387_,
		_w3404_
	);
	LUT4 #(
		.INIT('h0001)
	) name1504 (
		_w3388_,
		_w3401_,
		_w3403_,
		_w3404_,
		_w3405_
	);
	LUT3 #(
		.INIT('hce)
	) name1505 (
		\s5_msel_arb2_state_reg[2]/NET0131 ,
		_w3398_,
		_w3405_,
		_w3406_
	);
	LUT3 #(
		.INIT('h80)
	) name1506 (
		\m5_s5_cyc_o_reg/NET0131 ,
		\rf_conf5_reg[10]/NET0131 ,
		\rf_conf5_reg[11]/NET0131 ,
		_w3407_
	);
	LUT3 #(
		.INIT('h80)
	) name1507 (
		\m4_s5_cyc_o_reg/NET0131 ,
		\rf_conf5_reg[8]/NET0131 ,
		\rf_conf5_reg[9]/NET0131 ,
		_w3408_
	);
	LUT3 #(
		.INIT('h01)
	) name1508 (
		\s5_msel_arb3_state_reg[0]/NET0131 ,
		_w3407_,
		_w3408_,
		_w3409_
	);
	LUT2 #(
		.INIT('h8)
	) name1509 (
		\s5_msel_arb3_state_reg[0]/NET0131 ,
		\s5_msel_arb3_state_reg[2]/NET0131 ,
		_w3410_
	);
	LUT3 #(
		.INIT('h13)
	) name1510 (
		\s5_msel_arb3_state_reg[0]/NET0131 ,
		\s5_msel_arb3_state_reg[1]/NET0131 ,
		\s5_msel_arb3_state_reg[2]/NET0131 ,
		_w3411_
	);
	LUT4 #(
		.INIT('h0080)
	) name1511 (
		\m5_s5_cyc_o_reg/NET0131 ,
		\rf_conf5_reg[10]/NET0131 ,
		\rf_conf5_reg[11]/NET0131 ,
		\s5_msel_arb3_state_reg[1]/NET0131 ,
		_w3412_
	);
	LUT2 #(
		.INIT('h1)
	) name1512 (
		_w3411_,
		_w3412_,
		_w3413_
	);
	LUT3 #(
		.INIT('h80)
	) name1513 (
		\m7_s5_cyc_o_reg/NET0131 ,
		\rf_conf5_reg[14]/NET0131 ,
		\rf_conf5_reg[15]/NET0131 ,
		_w3414_
	);
	LUT3 #(
		.INIT('h80)
	) name1514 (
		\m6_s5_cyc_o_reg/NET0131 ,
		\rf_conf5_reg[12]/NET0131 ,
		\rf_conf5_reg[13]/NET0131 ,
		_w3415_
	);
	LUT2 #(
		.INIT('h1)
	) name1515 (
		_w3414_,
		_w3415_,
		_w3416_
	);
	LUT3 #(
		.INIT('h80)
	) name1516 (
		\m3_s5_cyc_o_reg/NET0131 ,
		\rf_conf5_reg[6]/NET0131 ,
		\rf_conf5_reg[7]/NET0131 ,
		_w3417_
	);
	LUT3 #(
		.INIT('h80)
	) name1517 (
		\m2_s5_cyc_o_reg/NET0131 ,
		\rf_conf5_reg[4]/NET0131 ,
		\rf_conf5_reg[5]/NET0131 ,
		_w3418_
	);
	LUT3 #(
		.INIT('h80)
	) name1518 (
		\m1_s5_cyc_o_reg/NET0131 ,
		\rf_conf5_reg[2]/NET0131 ,
		\rf_conf5_reg[3]/NET0131 ,
		_w3419_
	);
	LUT3 #(
		.INIT('h80)
	) name1519 (
		\m0_s5_cyc_o_reg/NET0131 ,
		\rf_conf5_reg[0]/NET0131 ,
		\rf_conf5_reg[1]/NET0131 ,
		_w3420_
	);
	LUT4 #(
		.INIT('h0001)
	) name1520 (
		_w3417_,
		_w3418_,
		_w3419_,
		_w3420_,
		_w3421_
	);
	LUT4 #(
		.INIT('h00e0)
	) name1521 (
		_w3409_,
		_w3413_,
		_w3416_,
		_w3421_,
		_w3422_
	);
	LUT4 #(
		.INIT('h3332)
	) name1522 (
		\s5_msel_arb3_state_reg[0]/NET0131 ,
		\s5_msel_arb3_state_reg[1]/NET0131 ,
		_w3419_,
		_w3420_,
		_w3423_
	);
	LUT4 #(
		.INIT('h0001)
	) name1523 (
		_w3407_,
		_w3408_,
		_w3414_,
		_w3415_,
		_w3424_
	);
	LUT4 #(
		.INIT('h0080)
	) name1524 (
		\m2_s5_cyc_o_reg/NET0131 ,
		\rf_conf5_reg[4]/NET0131 ,
		\rf_conf5_reg[5]/NET0131 ,
		\s5_msel_arb3_state_reg[0]/NET0131 ,
		_w3425_
	);
	LUT2 #(
		.INIT('h1)
	) name1525 (
		\s5_msel_arb3_state_reg[2]/NET0131 ,
		_w3425_,
		_w3426_
	);
	LUT3 #(
		.INIT('h01)
	) name1526 (
		\s5_msel_arb3_state_reg[2]/NET0131 ,
		_w3417_,
		_w3425_,
		_w3427_
	);
	LUT3 #(
		.INIT('h10)
	) name1527 (
		_w3423_,
		_w3424_,
		_w3427_,
		_w3428_
	);
	LUT2 #(
		.INIT('h8)
	) name1528 (
		\s5_msel_arb3_state_reg[0]/NET0131 ,
		\s5_msel_arb3_state_reg[1]/NET0131 ,
		_w3429_
	);
	LUT4 #(
		.INIT('h7f00)
	) name1529 (
		\m2_s5_cyc_o_reg/NET0131 ,
		\rf_conf5_reg[4]/NET0131 ,
		\rf_conf5_reg[5]/NET0131 ,
		\s5_msel_arb3_state_reg[0]/NET0131 ,
		_w3430_
	);
	LUT3 #(
		.INIT('h10)
	) name1530 (
		_w3417_,
		_w3419_,
		_w3430_,
		_w3431_
	);
	LUT4 #(
		.INIT('h0b0a)
	) name1531 (
		\s5_msel_arb3_state_reg[2]/NET0131 ,
		_w3424_,
		_w3429_,
		_w3431_,
		_w3432_
	);
	LUT2 #(
		.INIT('h8)
	) name1532 (
		\s5_msel_arb3_state_reg[1]/NET0131 ,
		\s5_msel_arb3_state_reg[2]/NET0131 ,
		_w3433_
	);
	LUT3 #(
		.INIT('h80)
	) name1533 (
		\s5_msel_arb3_state_reg[0]/NET0131 ,
		\s5_msel_arb3_state_reg[1]/NET0131 ,
		\s5_msel_arb3_state_reg[2]/NET0131 ,
		_w3434_
	);
	LUT3 #(
		.INIT('he0)
	) name1534 (
		_w3414_,
		_w3421_,
		_w3434_,
		_w3435_
	);
	LUT4 #(
		.INIT('hdddc)
	) name1535 (
		_w3422_,
		_w3428_,
		_w3432_,
		_w3435_,
		_w3436_
	);
	LUT3 #(
		.INIT('h80)
	) name1536 (
		\m5_s6_cyc_o_reg/NET0131 ,
		\rf_conf6_reg[10]/NET0131 ,
		\rf_conf6_reg[11]/NET0131 ,
		_w3437_
	);
	LUT3 #(
		.INIT('h80)
	) name1537 (
		\m4_s6_cyc_o_reg/NET0131 ,
		\rf_conf6_reg[8]/NET0131 ,
		\rf_conf6_reg[9]/NET0131 ,
		_w3438_
	);
	LUT3 #(
		.INIT('h01)
	) name1538 (
		\s6_msel_arb3_state_reg[0]/NET0131 ,
		_w3437_,
		_w3438_,
		_w3439_
	);
	LUT2 #(
		.INIT('h8)
	) name1539 (
		\s6_msel_arb3_state_reg[0]/NET0131 ,
		\s6_msel_arb3_state_reg[2]/NET0131 ,
		_w3440_
	);
	LUT3 #(
		.INIT('h13)
	) name1540 (
		\s6_msel_arb3_state_reg[0]/NET0131 ,
		\s6_msel_arb3_state_reg[1]/NET0131 ,
		\s6_msel_arb3_state_reg[2]/NET0131 ,
		_w3441_
	);
	LUT4 #(
		.INIT('h0080)
	) name1541 (
		\m5_s6_cyc_o_reg/NET0131 ,
		\rf_conf6_reg[10]/NET0131 ,
		\rf_conf6_reg[11]/NET0131 ,
		\s6_msel_arb3_state_reg[1]/NET0131 ,
		_w3442_
	);
	LUT2 #(
		.INIT('h1)
	) name1542 (
		_w3441_,
		_w3442_,
		_w3443_
	);
	LUT3 #(
		.INIT('h80)
	) name1543 (
		\m7_s6_cyc_o_reg/NET0131 ,
		\rf_conf6_reg[14]/NET0131 ,
		\rf_conf6_reg[15]/NET0131 ,
		_w3444_
	);
	LUT3 #(
		.INIT('h80)
	) name1544 (
		\m6_s6_cyc_o_reg/NET0131 ,
		\rf_conf6_reg[12]/NET0131 ,
		\rf_conf6_reg[13]/NET0131 ,
		_w3445_
	);
	LUT2 #(
		.INIT('h1)
	) name1545 (
		_w3444_,
		_w3445_,
		_w3446_
	);
	LUT3 #(
		.INIT('h80)
	) name1546 (
		\m3_s6_cyc_o_reg/NET0131 ,
		\rf_conf6_reg[6]/NET0131 ,
		\rf_conf6_reg[7]/NET0131 ,
		_w3447_
	);
	LUT3 #(
		.INIT('h80)
	) name1547 (
		\m2_s6_cyc_o_reg/NET0131 ,
		\rf_conf6_reg[4]/NET0131 ,
		\rf_conf6_reg[5]/NET0131 ,
		_w3448_
	);
	LUT3 #(
		.INIT('h80)
	) name1548 (
		\m1_s6_cyc_o_reg/NET0131 ,
		\rf_conf6_reg[2]/NET0131 ,
		\rf_conf6_reg[3]/NET0131 ,
		_w3449_
	);
	LUT3 #(
		.INIT('h80)
	) name1549 (
		\m0_s6_cyc_o_reg/NET0131 ,
		\rf_conf6_reg[0]/NET0131 ,
		\rf_conf6_reg[1]/NET0131 ,
		_w3450_
	);
	LUT4 #(
		.INIT('h0001)
	) name1550 (
		_w3447_,
		_w3448_,
		_w3449_,
		_w3450_,
		_w3451_
	);
	LUT4 #(
		.INIT('h00e0)
	) name1551 (
		_w3439_,
		_w3443_,
		_w3446_,
		_w3451_,
		_w3452_
	);
	LUT4 #(
		.INIT('h3332)
	) name1552 (
		\s6_msel_arb3_state_reg[0]/NET0131 ,
		\s6_msel_arb3_state_reg[1]/NET0131 ,
		_w3449_,
		_w3450_,
		_w3453_
	);
	LUT4 #(
		.INIT('h0001)
	) name1553 (
		_w3437_,
		_w3438_,
		_w3444_,
		_w3445_,
		_w3454_
	);
	LUT4 #(
		.INIT('h0080)
	) name1554 (
		\m2_s6_cyc_o_reg/NET0131 ,
		\rf_conf6_reg[4]/NET0131 ,
		\rf_conf6_reg[5]/NET0131 ,
		\s6_msel_arb3_state_reg[0]/NET0131 ,
		_w3455_
	);
	LUT2 #(
		.INIT('h1)
	) name1555 (
		\s6_msel_arb3_state_reg[2]/NET0131 ,
		_w3455_,
		_w3456_
	);
	LUT3 #(
		.INIT('h01)
	) name1556 (
		\s6_msel_arb3_state_reg[2]/NET0131 ,
		_w3447_,
		_w3455_,
		_w3457_
	);
	LUT3 #(
		.INIT('h10)
	) name1557 (
		_w3453_,
		_w3454_,
		_w3457_,
		_w3458_
	);
	LUT2 #(
		.INIT('h8)
	) name1558 (
		\s6_msel_arb3_state_reg[0]/NET0131 ,
		\s6_msel_arb3_state_reg[1]/NET0131 ,
		_w3459_
	);
	LUT4 #(
		.INIT('h7f00)
	) name1559 (
		\m2_s6_cyc_o_reg/NET0131 ,
		\rf_conf6_reg[4]/NET0131 ,
		\rf_conf6_reg[5]/NET0131 ,
		\s6_msel_arb3_state_reg[0]/NET0131 ,
		_w3460_
	);
	LUT3 #(
		.INIT('h10)
	) name1560 (
		_w3447_,
		_w3449_,
		_w3460_,
		_w3461_
	);
	LUT4 #(
		.INIT('h0b0a)
	) name1561 (
		\s6_msel_arb3_state_reg[2]/NET0131 ,
		_w3454_,
		_w3459_,
		_w3461_,
		_w3462_
	);
	LUT2 #(
		.INIT('h8)
	) name1562 (
		\s6_msel_arb3_state_reg[1]/NET0131 ,
		\s6_msel_arb3_state_reg[2]/NET0131 ,
		_w3463_
	);
	LUT3 #(
		.INIT('h80)
	) name1563 (
		\s6_msel_arb3_state_reg[0]/NET0131 ,
		\s6_msel_arb3_state_reg[1]/NET0131 ,
		\s6_msel_arb3_state_reg[2]/NET0131 ,
		_w3464_
	);
	LUT3 #(
		.INIT('he0)
	) name1564 (
		_w3444_,
		_w3451_,
		_w3464_,
		_w3465_
	);
	LUT4 #(
		.INIT('hdddc)
	) name1565 (
		_w3452_,
		_w3458_,
		_w3462_,
		_w3465_,
		_w3466_
	);
	LUT3 #(
		.INIT('h80)
	) name1566 (
		\m5_s7_cyc_o_reg/NET0131 ,
		\rf_conf7_reg[10]/NET0131 ,
		\rf_conf7_reg[11]/NET0131 ,
		_w3467_
	);
	LUT3 #(
		.INIT('h80)
	) name1567 (
		\m4_s7_cyc_o_reg/NET0131 ,
		\rf_conf7_reg[8]/NET0131 ,
		\rf_conf7_reg[9]/NET0131 ,
		_w3468_
	);
	LUT3 #(
		.INIT('h01)
	) name1568 (
		\s7_msel_arb3_state_reg[0]/NET0131 ,
		_w3467_,
		_w3468_,
		_w3469_
	);
	LUT2 #(
		.INIT('h8)
	) name1569 (
		\s7_msel_arb3_state_reg[0]/NET0131 ,
		\s7_msel_arb3_state_reg[2]/NET0131 ,
		_w3470_
	);
	LUT3 #(
		.INIT('h13)
	) name1570 (
		\s7_msel_arb3_state_reg[0]/NET0131 ,
		\s7_msel_arb3_state_reg[1]/NET0131 ,
		\s7_msel_arb3_state_reg[2]/NET0131 ,
		_w3471_
	);
	LUT4 #(
		.INIT('h0080)
	) name1571 (
		\m5_s7_cyc_o_reg/NET0131 ,
		\rf_conf7_reg[10]/NET0131 ,
		\rf_conf7_reg[11]/NET0131 ,
		\s7_msel_arb3_state_reg[1]/NET0131 ,
		_w3472_
	);
	LUT2 #(
		.INIT('h1)
	) name1572 (
		_w3471_,
		_w3472_,
		_w3473_
	);
	LUT3 #(
		.INIT('h80)
	) name1573 (
		\m7_s7_cyc_o_reg/NET0131 ,
		\rf_conf7_reg[14]/NET0131 ,
		\rf_conf7_reg[15]/NET0131 ,
		_w3474_
	);
	LUT3 #(
		.INIT('h80)
	) name1574 (
		\m6_s7_cyc_o_reg/NET0131 ,
		\rf_conf7_reg[12]/NET0131 ,
		\rf_conf7_reg[13]/NET0131 ,
		_w3475_
	);
	LUT2 #(
		.INIT('h1)
	) name1575 (
		_w3474_,
		_w3475_,
		_w3476_
	);
	LUT3 #(
		.INIT('h80)
	) name1576 (
		\m3_s7_cyc_o_reg/NET0131 ,
		\rf_conf7_reg[6]/NET0131 ,
		\rf_conf7_reg[7]/NET0131 ,
		_w3477_
	);
	LUT3 #(
		.INIT('h80)
	) name1577 (
		\m2_s7_cyc_o_reg/NET0131 ,
		\rf_conf7_reg[4]/NET0131 ,
		\rf_conf7_reg[5]/NET0131 ,
		_w3478_
	);
	LUT3 #(
		.INIT('h80)
	) name1578 (
		\m1_s7_cyc_o_reg/NET0131 ,
		\rf_conf7_reg[2]/NET0131 ,
		\rf_conf7_reg[3]/NET0131 ,
		_w3479_
	);
	LUT3 #(
		.INIT('h80)
	) name1579 (
		\m0_s7_cyc_o_reg/NET0131 ,
		\rf_conf7_reg[0]/NET0131 ,
		\rf_conf7_reg[1]/NET0131 ,
		_w3480_
	);
	LUT4 #(
		.INIT('h0001)
	) name1580 (
		_w3477_,
		_w3478_,
		_w3479_,
		_w3480_,
		_w3481_
	);
	LUT4 #(
		.INIT('h00e0)
	) name1581 (
		_w3469_,
		_w3473_,
		_w3476_,
		_w3481_,
		_w3482_
	);
	LUT4 #(
		.INIT('h3332)
	) name1582 (
		\s7_msel_arb3_state_reg[0]/NET0131 ,
		\s7_msel_arb3_state_reg[1]/NET0131 ,
		_w3479_,
		_w3480_,
		_w3483_
	);
	LUT4 #(
		.INIT('h0001)
	) name1583 (
		_w3467_,
		_w3468_,
		_w3474_,
		_w3475_,
		_w3484_
	);
	LUT4 #(
		.INIT('h0080)
	) name1584 (
		\m2_s7_cyc_o_reg/NET0131 ,
		\rf_conf7_reg[4]/NET0131 ,
		\rf_conf7_reg[5]/NET0131 ,
		\s7_msel_arb3_state_reg[0]/NET0131 ,
		_w3485_
	);
	LUT2 #(
		.INIT('h1)
	) name1585 (
		\s7_msel_arb3_state_reg[2]/NET0131 ,
		_w3485_,
		_w3486_
	);
	LUT3 #(
		.INIT('h01)
	) name1586 (
		\s7_msel_arb3_state_reg[2]/NET0131 ,
		_w3477_,
		_w3485_,
		_w3487_
	);
	LUT3 #(
		.INIT('h10)
	) name1587 (
		_w3483_,
		_w3484_,
		_w3487_,
		_w3488_
	);
	LUT2 #(
		.INIT('h8)
	) name1588 (
		\s7_msel_arb3_state_reg[0]/NET0131 ,
		\s7_msel_arb3_state_reg[1]/NET0131 ,
		_w3489_
	);
	LUT4 #(
		.INIT('h7f00)
	) name1589 (
		\m2_s7_cyc_o_reg/NET0131 ,
		\rf_conf7_reg[4]/NET0131 ,
		\rf_conf7_reg[5]/NET0131 ,
		\s7_msel_arb3_state_reg[0]/NET0131 ,
		_w3490_
	);
	LUT3 #(
		.INIT('h10)
	) name1590 (
		_w3477_,
		_w3479_,
		_w3490_,
		_w3491_
	);
	LUT4 #(
		.INIT('h0b0a)
	) name1591 (
		\s7_msel_arb3_state_reg[2]/NET0131 ,
		_w3484_,
		_w3489_,
		_w3491_,
		_w3492_
	);
	LUT2 #(
		.INIT('h8)
	) name1592 (
		\s7_msel_arb3_state_reg[1]/NET0131 ,
		\s7_msel_arb3_state_reg[2]/NET0131 ,
		_w3493_
	);
	LUT3 #(
		.INIT('h80)
	) name1593 (
		\s7_msel_arb3_state_reg[0]/NET0131 ,
		\s7_msel_arb3_state_reg[1]/NET0131 ,
		\s7_msel_arb3_state_reg[2]/NET0131 ,
		_w3494_
	);
	LUT3 #(
		.INIT('he0)
	) name1594 (
		_w3474_,
		_w3481_,
		_w3494_,
		_w3495_
	);
	LUT4 #(
		.INIT('hdddc)
	) name1595 (
		_w3482_,
		_w3488_,
		_w3492_,
		_w3495_,
		_w3496_
	);
	LUT2 #(
		.INIT('h4)
	) name1596 (
		\s8_msel_arb3_state_reg[1]/NET0131 ,
		\s8_msel_arb3_state_reg[2]/NET0131 ,
		_w3497_
	);
	LUT3 #(
		.INIT('h80)
	) name1597 (
		\m1_s8_cyc_o_reg/NET0131 ,
		\rf_conf8_reg[2]/NET0131 ,
		\rf_conf8_reg[3]/NET0131 ,
		_w3498_
	);
	LUT3 #(
		.INIT('h80)
	) name1598 (
		\m0_s8_cyc_o_reg/NET0131 ,
		\rf_conf8_reg[0]/NET0131 ,
		\rf_conf8_reg[1]/NET0131 ,
		_w3499_
	);
	LUT3 #(
		.INIT('h80)
	) name1599 (
		\m3_s8_cyc_o_reg/NET0131 ,
		\rf_conf8_reg[6]/NET0131 ,
		\rf_conf8_reg[7]/NET0131 ,
		_w3500_
	);
	LUT3 #(
		.INIT('h80)
	) name1600 (
		\m2_s8_cyc_o_reg/NET0131 ,
		\rf_conf8_reg[4]/NET0131 ,
		\rf_conf8_reg[5]/NET0131 ,
		_w3501_
	);
	LUT4 #(
		.INIT('h0001)
	) name1601 (
		_w3498_,
		_w3499_,
		_w3500_,
		_w3501_,
		_w3502_
	);
	LUT3 #(
		.INIT('h80)
	) name1602 (
		\m5_s8_cyc_o_reg/NET0131 ,
		\rf_conf8_reg[10]/NET0131 ,
		\rf_conf8_reg[11]/NET0131 ,
		_w3503_
	);
	LUT3 #(
		.INIT('h80)
	) name1603 (
		\m7_s8_cyc_o_reg/NET0131 ,
		\rf_conf8_reg[14]/NET0131 ,
		\rf_conf8_reg[15]/NET0131 ,
		_w3504_
	);
	LUT3 #(
		.INIT('h80)
	) name1604 (
		\m6_s8_cyc_o_reg/NET0131 ,
		\rf_conf8_reg[12]/NET0131 ,
		\rf_conf8_reg[13]/NET0131 ,
		_w3505_
	);
	LUT2 #(
		.INIT('h1)
	) name1605 (
		_w3504_,
		_w3505_,
		_w3506_
	);
	LUT3 #(
		.INIT('h01)
	) name1606 (
		_w3503_,
		_w3504_,
		_w3505_,
		_w3507_
	);
	LUT3 #(
		.INIT('h8a)
	) name1607 (
		_w3497_,
		_w3502_,
		_w3507_,
		_w3508_
	);
	LUT2 #(
		.INIT('h8)
	) name1608 (
		\s8_msel_arb3_state_reg[1]/NET0131 ,
		\s8_msel_arb3_state_reg[2]/NET0131 ,
		_w3509_
	);
	LUT3 #(
		.INIT('he0)
	) name1609 (
		_w3502_,
		_w3504_,
		_w3509_,
		_w3510_
	);
	LUT3 #(
		.INIT('h80)
	) name1610 (
		\m4_s8_cyc_o_reg/NET0131 ,
		\rf_conf8_reg[8]/NET0131 ,
		\rf_conf8_reg[9]/NET0131 ,
		_w3511_
	);
	LUT2 #(
		.INIT('h1)
	) name1611 (
		_w3503_,
		_w3511_,
		_w3512_
	);
	LUT4 #(
		.INIT('h0001)
	) name1612 (
		_w3503_,
		_w3504_,
		_w3505_,
		_w3511_,
		_w3513_
	);
	LUT4 #(
		.INIT('h007f)
	) name1613 (
		\m1_s8_cyc_o_reg/NET0131 ,
		\rf_conf8_reg[2]/NET0131 ,
		\rf_conf8_reg[3]/NET0131 ,
		\s8_msel_arb3_state_reg[2]/NET0131 ,
		_w3514_
	);
	LUT4 #(
		.INIT('h007f)
	) name1614 (
		\m2_s8_cyc_o_reg/NET0131 ,
		\rf_conf8_reg[4]/NET0131 ,
		\rf_conf8_reg[5]/NET0131 ,
		\s8_msel_arb3_state_reg[1]/NET0131 ,
		_w3515_
	);
	LUT2 #(
		.INIT('h8)
	) name1615 (
		_w3514_,
		_w3515_,
		_w3516_
	);
	LUT3 #(
		.INIT('h10)
	) name1616 (
		_w3500_,
		_w3513_,
		_w3516_,
		_w3517_
	);
	LUT4 #(
		.INIT('haaa8)
	) name1617 (
		\s8_msel_arb3_state_reg[0]/NET0131 ,
		_w3508_,
		_w3510_,
		_w3517_,
		_w3518_
	);
	LUT4 #(
		.INIT('h0080)
	) name1618 (
		\m2_s8_cyc_o_reg/NET0131 ,
		\rf_conf8_reg[4]/NET0131 ,
		\rf_conf8_reg[5]/NET0131 ,
		\s8_msel_arb3_state_reg[0]/NET0131 ,
		_w3519_
	);
	LUT3 #(
		.INIT('h54)
	) name1619 (
		\s8_msel_arb3_state_reg[1]/NET0131 ,
		_w3498_,
		_w3499_,
		_w3520_
	);
	LUT4 #(
		.INIT('h00ab)
	) name1620 (
		\s8_msel_arb3_state_reg[1]/NET0131 ,
		_w3498_,
		_w3499_,
		_w3519_,
		_w3521_
	);
	LUT4 #(
		.INIT('h5455)
	) name1621 (
		\s8_msel_arb3_state_reg[2]/NET0131 ,
		_w3500_,
		_w3513_,
		_w3521_,
		_w3522_
	);
	LUT2 #(
		.INIT('h2)
	) name1622 (
		\s8_msel_arb3_state_reg[1]/NET0131 ,
		\s8_msel_arb3_state_reg[2]/NET0131 ,
		_w3523_
	);
	LUT3 #(
		.INIT('ha2)
	) name1623 (
		\s8_msel_arb3_state_reg[0]/NET0131 ,
		\s8_msel_arb3_state_reg[1]/NET0131 ,
		\s8_msel_arb3_state_reg[2]/NET0131 ,
		_w3524_
	);
	LUT3 #(
		.INIT('h32)
	) name1624 (
		_w3503_,
		_w3509_,
		_w3511_,
		_w3525_
	);
	LUT4 #(
		.INIT('h0f0b)
	) name1625 (
		_w3502_,
		_w3506_,
		_w3524_,
		_w3525_,
		_w3526_
	);
	LUT2 #(
		.INIT('h4)
	) name1626 (
		_w3522_,
		_w3526_,
		_w3527_
	);
	LUT2 #(
		.INIT('he)
	) name1627 (
		_w3518_,
		_w3527_,
		_w3528_
	);
	LUT3 #(
		.INIT('h80)
	) name1628 (
		\m5_s0_cyc_o_reg/NET0131 ,
		\rf_conf0_reg[10]/NET0131 ,
		\rf_conf0_reg[11]/NET0131 ,
		_w3529_
	);
	LUT3 #(
		.INIT('h80)
	) name1629 (
		\m4_s0_cyc_o_reg/NET0131 ,
		\rf_conf0_reg[8]/NET0131 ,
		\rf_conf0_reg[9]/NET0131 ,
		_w3530_
	);
	LUT3 #(
		.INIT('h01)
	) name1630 (
		\s0_msel_arb3_state_reg[0]/NET0131 ,
		_w3529_,
		_w3530_,
		_w3531_
	);
	LUT2 #(
		.INIT('h8)
	) name1631 (
		\s0_msel_arb3_state_reg[0]/NET0131 ,
		\s0_msel_arb3_state_reg[2]/NET0131 ,
		_w3532_
	);
	LUT3 #(
		.INIT('h13)
	) name1632 (
		\s0_msel_arb3_state_reg[0]/NET0131 ,
		\s0_msel_arb3_state_reg[1]/NET0131 ,
		\s0_msel_arb3_state_reg[2]/NET0131 ,
		_w3533_
	);
	LUT4 #(
		.INIT('h0080)
	) name1633 (
		\m5_s0_cyc_o_reg/NET0131 ,
		\rf_conf0_reg[10]/NET0131 ,
		\rf_conf0_reg[11]/NET0131 ,
		\s0_msel_arb3_state_reg[1]/NET0131 ,
		_w3534_
	);
	LUT2 #(
		.INIT('h1)
	) name1634 (
		_w3533_,
		_w3534_,
		_w3535_
	);
	LUT3 #(
		.INIT('h80)
	) name1635 (
		\m7_s0_cyc_o_reg/NET0131 ,
		\rf_conf0_reg[14]/NET0131 ,
		\rf_conf0_reg[15]/NET0131 ,
		_w3536_
	);
	LUT3 #(
		.INIT('h80)
	) name1636 (
		\m6_s0_cyc_o_reg/NET0131 ,
		\rf_conf0_reg[12]/NET0131 ,
		\rf_conf0_reg[13]/NET0131 ,
		_w3537_
	);
	LUT2 #(
		.INIT('h1)
	) name1637 (
		_w3536_,
		_w3537_,
		_w3538_
	);
	LUT3 #(
		.INIT('h80)
	) name1638 (
		\m3_s0_cyc_o_reg/NET0131 ,
		\rf_conf0_reg[6]/NET0131 ,
		\rf_conf0_reg[7]/NET0131 ,
		_w3539_
	);
	LUT3 #(
		.INIT('h80)
	) name1639 (
		\m2_s0_cyc_o_reg/NET0131 ,
		\rf_conf0_reg[4]/NET0131 ,
		\rf_conf0_reg[5]/NET0131 ,
		_w3540_
	);
	LUT3 #(
		.INIT('h80)
	) name1640 (
		\m1_s0_cyc_o_reg/NET0131 ,
		\rf_conf0_reg[2]/NET0131 ,
		\rf_conf0_reg[3]/NET0131 ,
		_w3541_
	);
	LUT3 #(
		.INIT('h80)
	) name1641 (
		\m0_s0_cyc_o_reg/NET0131 ,
		\rf_conf0_reg[0]/NET0131 ,
		\rf_conf0_reg[1]/NET0131 ,
		_w3542_
	);
	LUT4 #(
		.INIT('h0001)
	) name1642 (
		_w3539_,
		_w3540_,
		_w3541_,
		_w3542_,
		_w3543_
	);
	LUT4 #(
		.INIT('h00e0)
	) name1643 (
		_w3531_,
		_w3535_,
		_w3538_,
		_w3543_,
		_w3544_
	);
	LUT4 #(
		.INIT('h3332)
	) name1644 (
		\s0_msel_arb3_state_reg[0]/NET0131 ,
		\s0_msel_arb3_state_reg[1]/NET0131 ,
		_w3541_,
		_w3542_,
		_w3545_
	);
	LUT4 #(
		.INIT('h0001)
	) name1645 (
		_w3529_,
		_w3530_,
		_w3536_,
		_w3537_,
		_w3546_
	);
	LUT4 #(
		.INIT('h0080)
	) name1646 (
		\m2_s0_cyc_o_reg/NET0131 ,
		\rf_conf0_reg[4]/NET0131 ,
		\rf_conf0_reg[5]/NET0131 ,
		\s0_msel_arb3_state_reg[0]/NET0131 ,
		_w3547_
	);
	LUT2 #(
		.INIT('h1)
	) name1647 (
		\s0_msel_arb3_state_reg[2]/NET0131 ,
		_w3547_,
		_w3548_
	);
	LUT3 #(
		.INIT('h01)
	) name1648 (
		\s0_msel_arb3_state_reg[2]/NET0131 ,
		_w3539_,
		_w3547_,
		_w3549_
	);
	LUT3 #(
		.INIT('h10)
	) name1649 (
		_w3545_,
		_w3546_,
		_w3549_,
		_w3550_
	);
	LUT2 #(
		.INIT('h8)
	) name1650 (
		\s0_msel_arb3_state_reg[0]/NET0131 ,
		\s0_msel_arb3_state_reg[1]/NET0131 ,
		_w3551_
	);
	LUT4 #(
		.INIT('h7f00)
	) name1651 (
		\m2_s0_cyc_o_reg/NET0131 ,
		\rf_conf0_reg[4]/NET0131 ,
		\rf_conf0_reg[5]/NET0131 ,
		\s0_msel_arb3_state_reg[0]/NET0131 ,
		_w3552_
	);
	LUT3 #(
		.INIT('h10)
	) name1652 (
		_w3539_,
		_w3541_,
		_w3552_,
		_w3553_
	);
	LUT4 #(
		.INIT('h0b0a)
	) name1653 (
		\s0_msel_arb3_state_reg[2]/NET0131 ,
		_w3546_,
		_w3551_,
		_w3553_,
		_w3554_
	);
	LUT2 #(
		.INIT('h8)
	) name1654 (
		\s0_msel_arb3_state_reg[1]/NET0131 ,
		\s0_msel_arb3_state_reg[2]/NET0131 ,
		_w3555_
	);
	LUT3 #(
		.INIT('h80)
	) name1655 (
		\s0_msel_arb3_state_reg[0]/NET0131 ,
		\s0_msel_arb3_state_reg[1]/NET0131 ,
		\s0_msel_arb3_state_reg[2]/NET0131 ,
		_w3556_
	);
	LUT3 #(
		.INIT('he0)
	) name1656 (
		_w3536_,
		_w3543_,
		_w3556_,
		_w3557_
	);
	LUT4 #(
		.INIT('hdddc)
	) name1657 (
		_w3544_,
		_w3550_,
		_w3554_,
		_w3557_,
		_w3558_
	);
	LUT3 #(
		.INIT('h08)
	) name1658 (
		\m5_s10_cyc_o_reg/NET0131 ,
		\rf_conf10_reg[10]/NET0131 ,
		\rf_conf10_reg[11]/NET0131 ,
		_w3559_
	);
	LUT4 #(
		.INIT('h0008)
	) name1659 (
		\m5_s10_cyc_o_reg/NET0131 ,
		\rf_conf10_reg[10]/NET0131 ,
		\rf_conf10_reg[11]/NET0131 ,
		\s10_msel_arb1_state_reg[1]/NET0131 ,
		_w3560_
	);
	LUT3 #(
		.INIT('h08)
	) name1660 (
		\m4_s10_cyc_o_reg/NET0131 ,
		\rf_conf10_reg[8]/NET0131 ,
		\rf_conf10_reg[9]/NET0131 ,
		_w3561_
	);
	LUT2 #(
		.INIT('h1)
	) name1661 (
		\s10_msel_arb1_state_reg[0]/NET0131 ,
		\s10_msel_arb1_state_reg[1]/NET0131 ,
		_w3562_
	);
	LUT3 #(
		.INIT('h15)
	) name1662 (
		_w3560_,
		_w3561_,
		_w3562_,
		_w3563_
	);
	LUT3 #(
		.INIT('h08)
	) name1663 (
		\m2_s10_cyc_o_reg/NET0131 ,
		\rf_conf10_reg[4]/NET0131 ,
		\rf_conf10_reg[5]/NET0131 ,
		_w3564_
	);
	LUT3 #(
		.INIT('h08)
	) name1664 (
		\m3_s10_cyc_o_reg/NET0131 ,
		\rf_conf10_reg[6]/NET0131 ,
		\rf_conf10_reg[7]/NET0131 ,
		_w3565_
	);
	LUT2 #(
		.INIT('h1)
	) name1665 (
		_w3564_,
		_w3565_,
		_w3566_
	);
	LUT3 #(
		.INIT('h08)
	) name1666 (
		\m1_s10_cyc_o_reg/NET0131 ,
		\rf_conf10_reg[2]/NET0131 ,
		\rf_conf10_reg[3]/NET0131 ,
		_w3567_
	);
	LUT3 #(
		.INIT('h08)
	) name1667 (
		\m0_s10_cyc_o_reg/NET0131 ,
		\rf_conf10_reg[0]/NET0131 ,
		\rf_conf10_reg[1]/NET0131 ,
		_w3568_
	);
	LUT4 #(
		.INIT('h0001)
	) name1668 (
		_w3564_,
		_w3565_,
		_w3567_,
		_w3568_,
		_w3569_
	);
	LUT3 #(
		.INIT('h08)
	) name1669 (
		\m7_s10_cyc_o_reg/NET0131 ,
		\rf_conf10_reg[14]/NET0131 ,
		\rf_conf10_reg[15]/NET0131 ,
		_w3570_
	);
	LUT3 #(
		.INIT('h08)
	) name1670 (
		\m6_s10_cyc_o_reg/NET0131 ,
		\rf_conf10_reg[12]/NET0131 ,
		\rf_conf10_reg[13]/NET0131 ,
		_w3571_
	);
	LUT2 #(
		.INIT('h8)
	) name1671 (
		\s10_msel_arb1_state_reg[0]/NET0131 ,
		\s10_msel_arb1_state_reg[1]/NET0131 ,
		_w3572_
	);
	LUT3 #(
		.INIT('h51)
	) name1672 (
		_w3570_,
		_w3571_,
		_w3572_,
		_w3573_
	);
	LUT4 #(
		.INIT('ha2aa)
	) name1673 (
		\s10_msel_arb1_state_reg[2]/NET0131 ,
		_w3563_,
		_w3569_,
		_w3573_,
		_w3574_
	);
	LUT4 #(
		.INIT('h0008)
	) name1674 (
		\m0_s10_cyc_o_reg/NET0131 ,
		\rf_conf10_reg[0]/NET0131 ,
		\rf_conf10_reg[1]/NET0131 ,
		\s10_msel_arb1_state_reg[0]/NET0131 ,
		_w3575_
	);
	LUT3 #(
		.INIT('h54)
	) name1675 (
		\s10_msel_arb1_state_reg[1]/NET0131 ,
		_w3567_,
		_w3575_,
		_w3576_
	);
	LUT2 #(
		.INIT('h1)
	) name1676 (
		_w3559_,
		_w3561_,
		_w3577_
	);
	LUT2 #(
		.INIT('h1)
	) name1677 (
		_w3570_,
		_w3571_,
		_w3578_
	);
	LUT4 #(
		.INIT('h0001)
	) name1678 (
		_w3559_,
		_w3561_,
		_w3570_,
		_w3571_,
		_w3579_
	);
	LUT4 #(
		.INIT('h00f7)
	) name1679 (
		\m3_s10_cyc_o_reg/NET0131 ,
		\rf_conf10_reg[6]/NET0131 ,
		\rf_conf10_reg[7]/NET0131 ,
		\s10_msel_arb1_state_reg[2]/NET0131 ,
		_w3580_
	);
	LUT3 #(
		.INIT('hd0)
	) name1680 (
		_w3564_,
		_w3572_,
		_w3580_,
		_w3581_
	);
	LUT3 #(
		.INIT('h10)
	) name1681 (
		_w3576_,
		_w3579_,
		_w3581_,
		_w3582_
	);
	LUT2 #(
		.INIT('he)
	) name1682 (
		_w3574_,
		_w3582_,
		_w3583_
	);
	LUT3 #(
		.INIT('h08)
	) name1683 (
		\m3_s11_cyc_o_reg/NET0131 ,
		\rf_conf11_reg[6]/NET0131 ,
		\rf_conf11_reg[7]/NET0131 ,
		_w3584_
	);
	LUT2 #(
		.INIT('h2)
	) name1684 (
		\s11_msel_arb1_state_reg[1]/NET0131 ,
		\s11_msel_arb1_state_reg[2]/NET0131 ,
		_w3585_
	);
	LUT3 #(
		.INIT('h08)
	) name1685 (
		\s11_msel_arb1_state_reg[0]/NET0131 ,
		\s11_msel_arb1_state_reg[1]/NET0131 ,
		\s11_msel_arb1_state_reg[2]/NET0131 ,
		_w3586_
	);
	LUT3 #(
		.INIT('h08)
	) name1686 (
		\m7_s11_cyc_o_reg/NET0131 ,
		\rf_conf11_reg[14]/NET0131 ,
		\rf_conf11_reg[15]/NET0131 ,
		_w3587_
	);
	LUT3 #(
		.INIT('h08)
	) name1687 (
		\m6_s11_cyc_o_reg/NET0131 ,
		\rf_conf11_reg[12]/NET0131 ,
		\rf_conf11_reg[13]/NET0131 ,
		_w3588_
	);
	LUT2 #(
		.INIT('h1)
	) name1688 (
		_w3587_,
		_w3588_,
		_w3589_
	);
	LUT3 #(
		.INIT('h08)
	) name1689 (
		\m4_s11_cyc_o_reg/NET0131 ,
		\rf_conf11_reg[8]/NET0131 ,
		\rf_conf11_reg[9]/NET0131 ,
		_w3590_
	);
	LUT3 #(
		.INIT('h08)
	) name1690 (
		\m5_s11_cyc_o_reg/NET0131 ,
		\rf_conf11_reg[10]/NET0131 ,
		\rf_conf11_reg[11]/NET0131 ,
		_w3591_
	);
	LUT4 #(
		.INIT('h0001)
	) name1691 (
		_w3587_,
		_w3588_,
		_w3590_,
		_w3591_,
		_w3592_
	);
	LUT3 #(
		.INIT('h04)
	) name1692 (
		_w3584_,
		_w3586_,
		_w3592_,
		_w3593_
	);
	LUT3 #(
		.INIT('h08)
	) name1693 (
		\m0_s11_cyc_o_reg/NET0131 ,
		\rf_conf11_reg[0]/NET0131 ,
		\rf_conf11_reg[1]/NET0131 ,
		_w3594_
	);
	LUT2 #(
		.INIT('h8)
	) name1694 (
		\s11_msel_arb1_state_reg[1]/NET0131 ,
		\s11_msel_arb1_state_reg[2]/NET0131 ,
		_w3595_
	);
	LUT2 #(
		.INIT('h4)
	) name1695 (
		_w3594_,
		_w3595_,
		_w3596_
	);
	LUT2 #(
		.INIT('h4)
	) name1696 (
		\s11_msel_arb1_state_reg[0]/NET0131 ,
		\s11_msel_arb1_state_reg[1]/NET0131 ,
		_w3597_
	);
	LUT4 #(
		.INIT('h0008)
	) name1697 (
		\m0_s11_cyc_o_reg/NET0131 ,
		\rf_conf11_reg[0]/NET0131 ,
		\rf_conf11_reg[1]/NET0131 ,
		\s11_msel_arb1_state_reg[0]/NET0131 ,
		_w3598_
	);
	LUT3 #(
		.INIT('h01)
	) name1698 (
		\s11_msel_arb1_state_reg[2]/NET0131 ,
		_w3597_,
		_w3598_,
		_w3599_
	);
	LUT3 #(
		.INIT('h08)
	) name1699 (
		\m2_s11_cyc_o_reg/NET0131 ,
		\rf_conf11_reg[4]/NET0131 ,
		\rf_conf11_reg[5]/NET0131 ,
		_w3600_
	);
	LUT3 #(
		.INIT('h08)
	) name1700 (
		\m1_s11_cyc_o_reg/NET0131 ,
		\rf_conf11_reg[2]/NET0131 ,
		\rf_conf11_reg[3]/NET0131 ,
		_w3601_
	);
	LUT3 #(
		.INIT('h01)
	) name1701 (
		_w3584_,
		_w3600_,
		_w3601_,
		_w3602_
	);
	LUT4 #(
		.INIT('hdc00)
	) name1702 (
		_w3592_,
		_w3596_,
		_w3599_,
		_w3602_,
		_w3603_
	);
	LUT2 #(
		.INIT('h1)
	) name1703 (
		_w3593_,
		_w3603_,
		_w3604_
	);
	LUT2 #(
		.INIT('h1)
	) name1704 (
		_w3584_,
		_w3600_,
		_w3605_
	);
	LUT3 #(
		.INIT('h04)
	) name1705 (
		_w3584_,
		_w3585_,
		_w3600_,
		_w3606_
	);
	LUT3 #(
		.INIT('h10)
	) name1706 (
		\s11_msel_arb1_state_reg[0]/NET0131 ,
		_w3592_,
		_w3606_,
		_w3607_
	);
	LUT4 #(
		.INIT('h0001)
	) name1707 (
		_w3584_,
		_w3594_,
		_w3600_,
		_w3601_,
		_w3608_
	);
	LUT2 #(
		.INIT('h4)
	) name1708 (
		\s11_msel_arb1_state_reg[1]/NET0131 ,
		\s11_msel_arb1_state_reg[2]/NET0131 ,
		_w3609_
	);
	LUT3 #(
		.INIT('h10)
	) name1709 (
		\s11_msel_arb1_state_reg[0]/NET0131 ,
		\s11_msel_arb1_state_reg[1]/NET0131 ,
		\s11_msel_arb1_state_reg[2]/NET0131 ,
		_w3610_
	);
	LUT3 #(
		.INIT('hd0)
	) name1710 (
		_w3592_,
		_w3608_,
		_w3610_,
		_w3611_
	);
	LUT4 #(
		.INIT('h0008)
	) name1711 (
		\m6_s11_cyc_o_reg/NET0131 ,
		\rf_conf11_reg[12]/NET0131 ,
		\rf_conf11_reg[13]/NET0131 ,
		\s11_msel_arb1_state_reg[0]/NET0131 ,
		_w3612_
	);
	LUT4 #(
		.INIT('h8880)
	) name1712 (
		\s11_msel_arb1_state_reg[1]/NET0131 ,
		\s11_msel_arb1_state_reg[2]/NET0131 ,
		_w3587_,
		_w3612_,
		_w3613_
	);
	LUT3 #(
		.INIT('h01)
	) name1713 (
		_w3587_,
		_w3588_,
		_w3591_,
		_w3614_
	);
	LUT3 #(
		.INIT('h20)
	) name1714 (
		\s11_msel_arb1_state_reg[0]/NET0131 ,
		\s11_msel_arb1_state_reg[1]/NET0131 ,
		\s11_msel_arb1_state_reg[2]/NET0131 ,
		_w3615_
	);
	LUT4 #(
		.INIT('h1033)
	) name1715 (
		_w3608_,
		_w3613_,
		_w3614_,
		_w3615_,
		_w3616_
	);
	LUT3 #(
		.INIT('h10)
	) name1716 (
		_w3607_,
		_w3611_,
		_w3616_,
		_w3617_
	);
	LUT2 #(
		.INIT('h7)
	) name1717 (
		_w3604_,
		_w3617_,
		_w3618_
	);
	LUT3 #(
		.INIT('h08)
	) name1718 (
		\m1_s12_cyc_o_reg/NET0131 ,
		\rf_conf12_reg[2]/NET0131 ,
		\rf_conf12_reg[3]/NET0131 ,
		_w3619_
	);
	LUT4 #(
		.INIT('h0008)
	) name1719 (
		\m0_s12_cyc_o_reg/NET0131 ,
		\rf_conf12_reg[0]/NET0131 ,
		\rf_conf12_reg[1]/NET0131 ,
		\s12_msel_arb1_state_reg[0]/NET0131 ,
		_w3620_
	);
	LUT3 #(
		.INIT('h54)
	) name1720 (
		\s12_msel_arb1_state_reg[1]/NET0131 ,
		_w3619_,
		_w3620_,
		_w3621_
	);
	LUT3 #(
		.INIT('h08)
	) name1721 (
		\m7_s12_cyc_o_reg/NET0131 ,
		\rf_conf12_reg[14]/NET0131 ,
		\rf_conf12_reg[15]/NET0131 ,
		_w3622_
	);
	LUT3 #(
		.INIT('h08)
	) name1722 (
		\m6_s12_cyc_o_reg/NET0131 ,
		\rf_conf12_reg[12]/NET0131 ,
		\rf_conf12_reg[13]/NET0131 ,
		_w3623_
	);
	LUT2 #(
		.INIT('h1)
	) name1723 (
		_w3622_,
		_w3623_,
		_w3624_
	);
	LUT3 #(
		.INIT('h08)
	) name1724 (
		\m4_s12_cyc_o_reg/NET0131 ,
		\rf_conf12_reg[8]/NET0131 ,
		\rf_conf12_reg[9]/NET0131 ,
		_w3625_
	);
	LUT3 #(
		.INIT('h08)
	) name1725 (
		\m5_s12_cyc_o_reg/NET0131 ,
		\rf_conf12_reg[10]/NET0131 ,
		\rf_conf12_reg[11]/NET0131 ,
		_w3626_
	);
	LUT2 #(
		.INIT('h1)
	) name1726 (
		_w3625_,
		_w3626_,
		_w3627_
	);
	LUT4 #(
		.INIT('h0001)
	) name1727 (
		_w3622_,
		_w3623_,
		_w3625_,
		_w3626_,
		_w3628_
	);
	LUT2 #(
		.INIT('h8)
	) name1728 (
		\s12_msel_arb1_state_reg[0]/NET0131 ,
		\s12_msel_arb1_state_reg[1]/NET0131 ,
		_w3629_
	);
	LUT3 #(
		.INIT('h08)
	) name1729 (
		\m2_s12_cyc_o_reg/NET0131 ,
		\rf_conf12_reg[4]/NET0131 ,
		\rf_conf12_reg[5]/NET0131 ,
		_w3630_
	);
	LUT3 #(
		.INIT('h08)
	) name1730 (
		\m3_s12_cyc_o_reg/NET0131 ,
		\rf_conf12_reg[6]/NET0131 ,
		\rf_conf12_reg[7]/NET0131 ,
		_w3631_
	);
	LUT3 #(
		.INIT('h0b)
	) name1731 (
		_w3629_,
		_w3630_,
		_w3631_,
		_w3632_
	);
	LUT4 #(
		.INIT('h5455)
	) name1732 (
		\s12_msel_arb1_state_reg[2]/NET0131 ,
		_w3621_,
		_w3628_,
		_w3632_,
		_w3633_
	);
	LUT4 #(
		.INIT('h0008)
	) name1733 (
		\m6_s12_cyc_o_reg/NET0131 ,
		\rf_conf12_reg[12]/NET0131 ,
		\rf_conf12_reg[13]/NET0131 ,
		\s12_msel_arb1_state_reg[0]/NET0131 ,
		_w3634_
	);
	LUT2 #(
		.INIT('h2)
	) name1734 (
		\s12_msel_arb1_state_reg[1]/NET0131 ,
		_w3634_,
		_w3635_
	);
	LUT4 #(
		.INIT('h0008)
	) name1735 (
		\m4_s12_cyc_o_reg/NET0131 ,
		\rf_conf12_reg[8]/NET0131 ,
		\rf_conf12_reg[9]/NET0131 ,
		\s12_msel_arb1_state_reg[0]/NET0131 ,
		_w3636_
	);
	LUT3 #(
		.INIT('h01)
	) name1736 (
		_w3623_,
		_w3626_,
		_w3636_,
		_w3637_
	);
	LUT4 #(
		.INIT('hf700)
	) name1737 (
		\m7_s12_cyc_o_reg/NET0131 ,
		\rf_conf12_reg[14]/NET0131 ,
		\rf_conf12_reg[15]/NET0131 ,
		\s12_msel_arb1_state_reg[2]/NET0131 ,
		_w3638_
	);
	LUT3 #(
		.INIT('h08)
	) name1738 (
		\m0_s12_cyc_o_reg/NET0131 ,
		\rf_conf12_reg[0]/NET0131 ,
		\rf_conf12_reg[1]/NET0131 ,
		_w3639_
	);
	LUT2 #(
		.INIT('h1)
	) name1739 (
		_w3619_,
		_w3639_,
		_w3640_
	);
	LUT2 #(
		.INIT('h1)
	) name1740 (
		_w3630_,
		_w3631_,
		_w3641_
	);
	LUT4 #(
		.INIT('h0001)
	) name1741 (
		_w3619_,
		_w3630_,
		_w3631_,
		_w3639_,
		_w3642_
	);
	LUT4 #(
		.INIT('h00e0)
	) name1742 (
		_w3635_,
		_w3637_,
		_w3638_,
		_w3642_,
		_w3643_
	);
	LUT2 #(
		.INIT('h1)
	) name1743 (
		_w3633_,
		_w3643_,
		_w3644_
	);
	LUT3 #(
		.INIT('h08)
	) name1744 (
		\m5_s13_cyc_o_reg/NET0131 ,
		\rf_conf13_reg[10]/NET0131 ,
		\rf_conf13_reg[11]/NET0131 ,
		_w3645_
	);
	LUT4 #(
		.INIT('h0008)
	) name1745 (
		\m5_s13_cyc_o_reg/NET0131 ,
		\rf_conf13_reg[10]/NET0131 ,
		\rf_conf13_reg[11]/NET0131 ,
		\s13_msel_arb1_state_reg[1]/NET0131 ,
		_w3646_
	);
	LUT3 #(
		.INIT('h08)
	) name1746 (
		\m4_s13_cyc_o_reg/NET0131 ,
		\rf_conf13_reg[8]/NET0131 ,
		\rf_conf13_reg[9]/NET0131 ,
		_w3647_
	);
	LUT2 #(
		.INIT('h1)
	) name1747 (
		\s13_msel_arb1_state_reg[0]/NET0131 ,
		\s13_msel_arb1_state_reg[1]/NET0131 ,
		_w3648_
	);
	LUT3 #(
		.INIT('h15)
	) name1748 (
		_w3646_,
		_w3647_,
		_w3648_,
		_w3649_
	);
	LUT3 #(
		.INIT('h08)
	) name1749 (
		\m2_s13_cyc_o_reg/NET0131 ,
		\rf_conf13_reg[4]/NET0131 ,
		\rf_conf13_reg[5]/NET0131 ,
		_w3650_
	);
	LUT3 #(
		.INIT('h08)
	) name1750 (
		\m3_s13_cyc_o_reg/NET0131 ,
		\rf_conf13_reg[6]/NET0131 ,
		\rf_conf13_reg[7]/NET0131 ,
		_w3651_
	);
	LUT2 #(
		.INIT('h1)
	) name1751 (
		_w3650_,
		_w3651_,
		_w3652_
	);
	LUT3 #(
		.INIT('h08)
	) name1752 (
		\m1_s13_cyc_o_reg/NET0131 ,
		\rf_conf13_reg[2]/NET0131 ,
		\rf_conf13_reg[3]/NET0131 ,
		_w3653_
	);
	LUT3 #(
		.INIT('h08)
	) name1753 (
		\m0_s13_cyc_o_reg/NET0131 ,
		\rf_conf13_reg[0]/NET0131 ,
		\rf_conf13_reg[1]/NET0131 ,
		_w3654_
	);
	LUT4 #(
		.INIT('h0001)
	) name1754 (
		_w3650_,
		_w3651_,
		_w3653_,
		_w3654_,
		_w3655_
	);
	LUT3 #(
		.INIT('h08)
	) name1755 (
		\m7_s13_cyc_o_reg/NET0131 ,
		\rf_conf13_reg[14]/NET0131 ,
		\rf_conf13_reg[15]/NET0131 ,
		_w3656_
	);
	LUT3 #(
		.INIT('h08)
	) name1756 (
		\m6_s13_cyc_o_reg/NET0131 ,
		\rf_conf13_reg[12]/NET0131 ,
		\rf_conf13_reg[13]/NET0131 ,
		_w3657_
	);
	LUT2 #(
		.INIT('h8)
	) name1757 (
		\s13_msel_arb1_state_reg[0]/NET0131 ,
		\s13_msel_arb1_state_reg[1]/NET0131 ,
		_w3658_
	);
	LUT3 #(
		.INIT('h51)
	) name1758 (
		_w3656_,
		_w3657_,
		_w3658_,
		_w3659_
	);
	LUT4 #(
		.INIT('ha2aa)
	) name1759 (
		\s13_msel_arb1_state_reg[2]/NET0131 ,
		_w3649_,
		_w3655_,
		_w3659_,
		_w3660_
	);
	LUT4 #(
		.INIT('h0008)
	) name1760 (
		\m0_s13_cyc_o_reg/NET0131 ,
		\rf_conf13_reg[0]/NET0131 ,
		\rf_conf13_reg[1]/NET0131 ,
		\s13_msel_arb1_state_reg[0]/NET0131 ,
		_w3661_
	);
	LUT3 #(
		.INIT('h54)
	) name1761 (
		\s13_msel_arb1_state_reg[1]/NET0131 ,
		_w3653_,
		_w3661_,
		_w3662_
	);
	LUT2 #(
		.INIT('h1)
	) name1762 (
		_w3645_,
		_w3647_,
		_w3663_
	);
	LUT2 #(
		.INIT('h1)
	) name1763 (
		_w3656_,
		_w3657_,
		_w3664_
	);
	LUT4 #(
		.INIT('h0001)
	) name1764 (
		_w3645_,
		_w3647_,
		_w3656_,
		_w3657_,
		_w3665_
	);
	LUT4 #(
		.INIT('h00f7)
	) name1765 (
		\m3_s13_cyc_o_reg/NET0131 ,
		\rf_conf13_reg[6]/NET0131 ,
		\rf_conf13_reg[7]/NET0131 ,
		\s13_msel_arb1_state_reg[2]/NET0131 ,
		_w3666_
	);
	LUT3 #(
		.INIT('hd0)
	) name1766 (
		_w3650_,
		_w3658_,
		_w3666_,
		_w3667_
	);
	LUT3 #(
		.INIT('h10)
	) name1767 (
		_w3662_,
		_w3665_,
		_w3667_,
		_w3668_
	);
	LUT2 #(
		.INIT('he)
	) name1768 (
		_w3660_,
		_w3668_,
		_w3669_
	);
	LUT3 #(
		.INIT('h08)
	) name1769 (
		\m6_s14_cyc_o_reg/NET0131 ,
		\rf_conf14_reg[12]/NET0131 ,
		\rf_conf14_reg[13]/NET0131 ,
		_w3670_
	);
	LUT3 #(
		.INIT('h08)
	) name1770 (
		\m7_s14_cyc_o_reg/NET0131 ,
		\rf_conf14_reg[14]/NET0131 ,
		\rf_conf14_reg[15]/NET0131 ,
		_w3671_
	);
	LUT2 #(
		.INIT('h1)
	) name1771 (
		_w3670_,
		_w3671_,
		_w3672_
	);
	LUT3 #(
		.INIT('h08)
	) name1772 (
		\m4_s14_cyc_o_reg/NET0131 ,
		\rf_conf14_reg[8]/NET0131 ,
		\rf_conf14_reg[9]/NET0131 ,
		_w3673_
	);
	LUT3 #(
		.INIT('h08)
	) name1773 (
		\m5_s14_cyc_o_reg/NET0131 ,
		\rf_conf14_reg[10]/NET0131 ,
		\rf_conf14_reg[11]/NET0131 ,
		_w3674_
	);
	LUT4 #(
		.INIT('h0001)
	) name1774 (
		_w3670_,
		_w3671_,
		_w3673_,
		_w3674_,
		_w3675_
	);
	LUT2 #(
		.INIT('h4)
	) name1775 (
		\s14_msel_arb1_state_reg[1]/NET0131 ,
		\s14_msel_arb1_state_reg[2]/NET0131 ,
		_w3676_
	);
	LUT3 #(
		.INIT('h10)
	) name1776 (
		\s14_msel_arb1_state_reg[0]/NET0131 ,
		\s14_msel_arb1_state_reg[1]/NET0131 ,
		\s14_msel_arb1_state_reg[2]/NET0131 ,
		_w3677_
	);
	LUT3 #(
		.INIT('h08)
	) name1777 (
		\m3_s14_cyc_o_reg/NET0131 ,
		\rf_conf14_reg[6]/NET0131 ,
		\rf_conf14_reg[7]/NET0131 ,
		_w3678_
	);
	LUT4 #(
		.INIT('h00f7)
	) name1778 (
		\m3_s14_cyc_o_reg/NET0131 ,
		\rf_conf14_reg[6]/NET0131 ,
		\rf_conf14_reg[7]/NET0131 ,
		\s14_msel_arb1_state_reg[2]/NET0131 ,
		_w3679_
	);
	LUT2 #(
		.INIT('h1)
	) name1779 (
		_w3677_,
		_w3679_,
		_w3680_
	);
	LUT4 #(
		.INIT('h0008)
	) name1780 (
		\m0_s14_cyc_o_reg/NET0131 ,
		\rf_conf14_reg[0]/NET0131 ,
		\rf_conf14_reg[1]/NET0131 ,
		\s14_msel_arb1_state_reg[0]/NET0131 ,
		_w3681_
	);
	LUT3 #(
		.INIT('h08)
	) name1781 (
		\m2_s14_cyc_o_reg/NET0131 ,
		\rf_conf14_reg[4]/NET0131 ,
		\rf_conf14_reg[5]/NET0131 ,
		_w3682_
	);
	LUT3 #(
		.INIT('h08)
	) name1782 (
		\m1_s14_cyc_o_reg/NET0131 ,
		\rf_conf14_reg[2]/NET0131 ,
		\rf_conf14_reg[3]/NET0131 ,
		_w3683_
	);
	LUT3 #(
		.INIT('h01)
	) name1783 (
		_w3681_,
		_w3682_,
		_w3683_,
		_w3684_
	);
	LUT4 #(
		.INIT('h0008)
	) name1784 (
		\m2_s14_cyc_o_reg/NET0131 ,
		\rf_conf14_reg[4]/NET0131 ,
		\rf_conf14_reg[5]/NET0131 ,
		\s14_msel_arb1_state_reg[0]/NET0131 ,
		_w3685_
	);
	LUT3 #(
		.INIT('h31)
	) name1785 (
		\s14_msel_arb1_state_reg[1]/NET0131 ,
		_w3677_,
		_w3685_,
		_w3686_
	);
	LUT4 #(
		.INIT('h1011)
	) name1786 (
		_w3675_,
		_w3680_,
		_w3684_,
		_w3686_,
		_w3687_
	);
	LUT3 #(
		.INIT('h08)
	) name1787 (
		\m0_s14_cyc_o_reg/NET0131 ,
		\rf_conf14_reg[0]/NET0131 ,
		\rf_conf14_reg[1]/NET0131 ,
		_w3688_
	);
	LUT2 #(
		.INIT('h1)
	) name1788 (
		_w3678_,
		_w3682_,
		_w3689_
	);
	LUT4 #(
		.INIT('h0001)
	) name1789 (
		_w3678_,
		_w3682_,
		_w3683_,
		_w3688_,
		_w3690_
	);
	LUT4 #(
		.INIT('h1115)
	) name1790 (
		\s14_msel_arb1_state_reg[0]/NET0131 ,
		\s14_msel_arb1_state_reg[1]/NET0131 ,
		_w3670_,
		_w3671_,
		_w3691_
	);
	LUT2 #(
		.INIT('h8)
	) name1791 (
		\s14_msel_arb1_state_reg[0]/NET0131 ,
		\s14_msel_arb1_state_reg[1]/NET0131 ,
		_w3692_
	);
	LUT4 #(
		.INIT('h3301)
	) name1792 (
		_w3670_,
		_w3671_,
		_w3674_,
		_w3692_,
		_w3693_
	);
	LUT4 #(
		.INIT('h888a)
	) name1793 (
		\s14_msel_arb1_state_reg[2]/NET0131 ,
		_w3690_,
		_w3691_,
		_w3693_,
		_w3694_
	);
	LUT2 #(
		.INIT('he)
	) name1794 (
		_w3687_,
		_w3694_,
		_w3695_
	);
	LUT3 #(
		.INIT('h08)
	) name1795 (
		\m6_s1_cyc_o_reg/NET0131 ,
		\rf_conf1_reg[12]/NET0131 ,
		\rf_conf1_reg[13]/NET0131 ,
		_w3696_
	);
	LUT3 #(
		.INIT('h08)
	) name1796 (
		\m7_s1_cyc_o_reg/NET0131 ,
		\rf_conf1_reg[14]/NET0131 ,
		\rf_conf1_reg[15]/NET0131 ,
		_w3697_
	);
	LUT2 #(
		.INIT('h1)
	) name1797 (
		_w3696_,
		_w3697_,
		_w3698_
	);
	LUT3 #(
		.INIT('h08)
	) name1798 (
		\m4_s1_cyc_o_reg/NET0131 ,
		\rf_conf1_reg[8]/NET0131 ,
		\rf_conf1_reg[9]/NET0131 ,
		_w3699_
	);
	LUT3 #(
		.INIT('h08)
	) name1799 (
		\m5_s1_cyc_o_reg/NET0131 ,
		\rf_conf1_reg[10]/NET0131 ,
		\rf_conf1_reg[11]/NET0131 ,
		_w3700_
	);
	LUT4 #(
		.INIT('h0001)
	) name1800 (
		_w3696_,
		_w3697_,
		_w3699_,
		_w3700_,
		_w3701_
	);
	LUT2 #(
		.INIT('h4)
	) name1801 (
		\s1_msel_arb1_state_reg[1]/NET0131 ,
		\s1_msel_arb1_state_reg[2]/NET0131 ,
		_w3702_
	);
	LUT3 #(
		.INIT('h10)
	) name1802 (
		\s1_msel_arb1_state_reg[0]/NET0131 ,
		\s1_msel_arb1_state_reg[1]/NET0131 ,
		\s1_msel_arb1_state_reg[2]/NET0131 ,
		_w3703_
	);
	LUT3 #(
		.INIT('h08)
	) name1803 (
		\m3_s1_cyc_o_reg/NET0131 ,
		\rf_conf1_reg[6]/NET0131 ,
		\rf_conf1_reg[7]/NET0131 ,
		_w3704_
	);
	LUT4 #(
		.INIT('h00f7)
	) name1804 (
		\m3_s1_cyc_o_reg/NET0131 ,
		\rf_conf1_reg[6]/NET0131 ,
		\rf_conf1_reg[7]/NET0131 ,
		\s1_msel_arb1_state_reg[2]/NET0131 ,
		_w3705_
	);
	LUT2 #(
		.INIT('h1)
	) name1805 (
		_w3703_,
		_w3705_,
		_w3706_
	);
	LUT4 #(
		.INIT('h0008)
	) name1806 (
		\m0_s1_cyc_o_reg/NET0131 ,
		\rf_conf1_reg[0]/NET0131 ,
		\rf_conf1_reg[1]/NET0131 ,
		\s1_msel_arb1_state_reg[0]/NET0131 ,
		_w3707_
	);
	LUT3 #(
		.INIT('h08)
	) name1807 (
		\m2_s1_cyc_o_reg/NET0131 ,
		\rf_conf1_reg[4]/NET0131 ,
		\rf_conf1_reg[5]/NET0131 ,
		_w3708_
	);
	LUT3 #(
		.INIT('h08)
	) name1808 (
		\m1_s1_cyc_o_reg/NET0131 ,
		\rf_conf1_reg[2]/NET0131 ,
		\rf_conf1_reg[3]/NET0131 ,
		_w3709_
	);
	LUT3 #(
		.INIT('h01)
	) name1809 (
		_w3707_,
		_w3708_,
		_w3709_,
		_w3710_
	);
	LUT4 #(
		.INIT('h0008)
	) name1810 (
		\m2_s1_cyc_o_reg/NET0131 ,
		\rf_conf1_reg[4]/NET0131 ,
		\rf_conf1_reg[5]/NET0131 ,
		\s1_msel_arb1_state_reg[0]/NET0131 ,
		_w3711_
	);
	LUT3 #(
		.INIT('h31)
	) name1811 (
		\s1_msel_arb1_state_reg[1]/NET0131 ,
		_w3703_,
		_w3711_,
		_w3712_
	);
	LUT4 #(
		.INIT('h1011)
	) name1812 (
		_w3701_,
		_w3706_,
		_w3710_,
		_w3712_,
		_w3713_
	);
	LUT3 #(
		.INIT('h08)
	) name1813 (
		\m0_s1_cyc_o_reg/NET0131 ,
		\rf_conf1_reg[0]/NET0131 ,
		\rf_conf1_reg[1]/NET0131 ,
		_w3714_
	);
	LUT2 #(
		.INIT('h1)
	) name1814 (
		_w3704_,
		_w3708_,
		_w3715_
	);
	LUT4 #(
		.INIT('h0001)
	) name1815 (
		_w3704_,
		_w3708_,
		_w3709_,
		_w3714_,
		_w3716_
	);
	LUT4 #(
		.INIT('h1115)
	) name1816 (
		\s1_msel_arb1_state_reg[0]/NET0131 ,
		\s1_msel_arb1_state_reg[1]/NET0131 ,
		_w3696_,
		_w3697_,
		_w3717_
	);
	LUT2 #(
		.INIT('h8)
	) name1817 (
		\s1_msel_arb1_state_reg[0]/NET0131 ,
		\s1_msel_arb1_state_reg[1]/NET0131 ,
		_w3718_
	);
	LUT4 #(
		.INIT('h3301)
	) name1818 (
		_w3696_,
		_w3697_,
		_w3700_,
		_w3718_,
		_w3719_
	);
	LUT4 #(
		.INIT('h888a)
	) name1819 (
		\s1_msel_arb1_state_reg[2]/NET0131 ,
		_w3716_,
		_w3717_,
		_w3719_,
		_w3720_
	);
	LUT2 #(
		.INIT('he)
	) name1820 (
		_w3713_,
		_w3720_,
		_w3721_
	);
	LUT3 #(
		.INIT('h08)
	) name1821 (
		\m5_s2_cyc_o_reg/NET0131 ,
		\rf_conf2_reg[10]/NET0131 ,
		\rf_conf2_reg[11]/NET0131 ,
		_w3722_
	);
	LUT4 #(
		.INIT('h0008)
	) name1822 (
		\m5_s2_cyc_o_reg/NET0131 ,
		\rf_conf2_reg[10]/NET0131 ,
		\rf_conf2_reg[11]/NET0131 ,
		\s2_msel_arb1_state_reg[1]/NET0131 ,
		_w3723_
	);
	LUT3 #(
		.INIT('h08)
	) name1823 (
		\m4_s2_cyc_o_reg/NET0131 ,
		\rf_conf2_reg[8]/NET0131 ,
		\rf_conf2_reg[9]/NET0131 ,
		_w3724_
	);
	LUT2 #(
		.INIT('h1)
	) name1824 (
		\s2_msel_arb1_state_reg[0]/NET0131 ,
		\s2_msel_arb1_state_reg[1]/NET0131 ,
		_w3725_
	);
	LUT3 #(
		.INIT('h15)
	) name1825 (
		_w3723_,
		_w3724_,
		_w3725_,
		_w3726_
	);
	LUT3 #(
		.INIT('h08)
	) name1826 (
		\m2_s2_cyc_o_reg/NET0131 ,
		\rf_conf2_reg[4]/NET0131 ,
		\rf_conf2_reg[5]/NET0131 ,
		_w3727_
	);
	LUT3 #(
		.INIT('h08)
	) name1827 (
		\m3_s2_cyc_o_reg/NET0131 ,
		\rf_conf2_reg[6]/NET0131 ,
		\rf_conf2_reg[7]/NET0131 ,
		_w3728_
	);
	LUT2 #(
		.INIT('h1)
	) name1828 (
		_w3727_,
		_w3728_,
		_w3729_
	);
	LUT3 #(
		.INIT('h08)
	) name1829 (
		\m1_s2_cyc_o_reg/NET0131 ,
		\rf_conf2_reg[2]/NET0131 ,
		\rf_conf2_reg[3]/NET0131 ,
		_w3730_
	);
	LUT3 #(
		.INIT('h08)
	) name1830 (
		\m0_s2_cyc_o_reg/NET0131 ,
		\rf_conf2_reg[0]/NET0131 ,
		\rf_conf2_reg[1]/NET0131 ,
		_w3731_
	);
	LUT4 #(
		.INIT('h0001)
	) name1831 (
		_w3727_,
		_w3728_,
		_w3730_,
		_w3731_,
		_w3732_
	);
	LUT3 #(
		.INIT('h08)
	) name1832 (
		\m7_s2_cyc_o_reg/NET0131 ,
		\rf_conf2_reg[14]/NET0131 ,
		\rf_conf2_reg[15]/NET0131 ,
		_w3733_
	);
	LUT3 #(
		.INIT('h08)
	) name1833 (
		\m6_s2_cyc_o_reg/NET0131 ,
		\rf_conf2_reg[12]/NET0131 ,
		\rf_conf2_reg[13]/NET0131 ,
		_w3734_
	);
	LUT2 #(
		.INIT('h8)
	) name1834 (
		\s2_msel_arb1_state_reg[0]/NET0131 ,
		\s2_msel_arb1_state_reg[1]/NET0131 ,
		_w3735_
	);
	LUT3 #(
		.INIT('h51)
	) name1835 (
		_w3733_,
		_w3734_,
		_w3735_,
		_w3736_
	);
	LUT4 #(
		.INIT('ha2aa)
	) name1836 (
		\s2_msel_arb1_state_reg[2]/NET0131 ,
		_w3726_,
		_w3732_,
		_w3736_,
		_w3737_
	);
	LUT4 #(
		.INIT('h0008)
	) name1837 (
		\m0_s2_cyc_o_reg/NET0131 ,
		\rf_conf2_reg[0]/NET0131 ,
		\rf_conf2_reg[1]/NET0131 ,
		\s2_msel_arb1_state_reg[0]/NET0131 ,
		_w3738_
	);
	LUT3 #(
		.INIT('h54)
	) name1838 (
		\s2_msel_arb1_state_reg[1]/NET0131 ,
		_w3730_,
		_w3738_,
		_w3739_
	);
	LUT2 #(
		.INIT('h1)
	) name1839 (
		_w3722_,
		_w3724_,
		_w3740_
	);
	LUT2 #(
		.INIT('h1)
	) name1840 (
		_w3733_,
		_w3734_,
		_w3741_
	);
	LUT4 #(
		.INIT('h0001)
	) name1841 (
		_w3722_,
		_w3724_,
		_w3733_,
		_w3734_,
		_w3742_
	);
	LUT4 #(
		.INIT('h00f7)
	) name1842 (
		\m3_s2_cyc_o_reg/NET0131 ,
		\rf_conf2_reg[6]/NET0131 ,
		\rf_conf2_reg[7]/NET0131 ,
		\s2_msel_arb1_state_reg[2]/NET0131 ,
		_w3743_
	);
	LUT3 #(
		.INIT('hd0)
	) name1843 (
		_w3727_,
		_w3735_,
		_w3743_,
		_w3744_
	);
	LUT3 #(
		.INIT('h10)
	) name1844 (
		_w3739_,
		_w3742_,
		_w3744_,
		_w3745_
	);
	LUT2 #(
		.INIT('he)
	) name1845 (
		_w3737_,
		_w3745_,
		_w3746_
	);
	LUT2 #(
		.INIT('h4)
	) name1846 (
		\s3_msel_arb1_state_reg[0]/NET0131 ,
		\s3_msel_arb1_state_reg[1]/NET0131 ,
		_w3747_
	);
	LUT3 #(
		.INIT('h08)
	) name1847 (
		\m7_s3_cyc_o_reg/NET0131 ,
		\rf_conf3_reg[14]/NET0131 ,
		\rf_conf3_reg[15]/NET0131 ,
		_w3748_
	);
	LUT3 #(
		.INIT('h08)
	) name1848 (
		\m6_s3_cyc_o_reg/NET0131 ,
		\rf_conf3_reg[12]/NET0131 ,
		\rf_conf3_reg[13]/NET0131 ,
		_w3749_
	);
	LUT2 #(
		.INIT('h1)
	) name1849 (
		_w3748_,
		_w3749_,
		_w3750_
	);
	LUT3 #(
		.INIT('ha8)
	) name1850 (
		\s3_msel_arb1_state_reg[2]/NET0131 ,
		_w3748_,
		_w3749_,
		_w3751_
	);
	LUT3 #(
		.INIT('h08)
	) name1851 (
		\m4_s3_cyc_o_reg/NET0131 ,
		\rf_conf3_reg[8]/NET0131 ,
		\rf_conf3_reg[9]/NET0131 ,
		_w3752_
	);
	LUT3 #(
		.INIT('h08)
	) name1852 (
		\m5_s3_cyc_o_reg/NET0131 ,
		\rf_conf3_reg[10]/NET0131 ,
		\rf_conf3_reg[11]/NET0131 ,
		_w3753_
	);
	LUT2 #(
		.INIT('h1)
	) name1853 (
		_w3752_,
		_w3753_,
		_w3754_
	);
	LUT4 #(
		.INIT('h0001)
	) name1854 (
		_w3748_,
		_w3749_,
		_w3752_,
		_w3753_,
		_w3755_
	);
	LUT3 #(
		.INIT('h08)
	) name1855 (
		\m2_s3_cyc_o_reg/NET0131 ,
		\rf_conf3_reg[4]/NET0131 ,
		\rf_conf3_reg[5]/NET0131 ,
		_w3756_
	);
	LUT3 #(
		.INIT('h08)
	) name1856 (
		\m3_s3_cyc_o_reg/NET0131 ,
		\rf_conf3_reg[6]/NET0131 ,
		\rf_conf3_reg[7]/NET0131 ,
		_w3757_
	);
	LUT2 #(
		.INIT('h1)
	) name1857 (
		_w3756_,
		_w3757_,
		_w3758_
	);
	LUT3 #(
		.INIT('h08)
	) name1858 (
		\m1_s3_cyc_o_reg/NET0131 ,
		\rf_conf3_reg[2]/NET0131 ,
		\rf_conf3_reg[3]/NET0131 ,
		_w3759_
	);
	LUT3 #(
		.INIT('h08)
	) name1859 (
		\m0_s3_cyc_o_reg/NET0131 ,
		\rf_conf3_reg[0]/NET0131 ,
		\rf_conf3_reg[1]/NET0131 ,
		_w3760_
	);
	LUT2 #(
		.INIT('h1)
	) name1860 (
		_w3759_,
		_w3760_,
		_w3761_
	);
	LUT4 #(
		.INIT('hb010)
	) name1861 (
		\s3_msel_arb1_state_reg[2]/NET0131 ,
		_w3755_,
		_w3758_,
		_w3761_,
		_w3762_
	);
	LUT3 #(
		.INIT('ha8)
	) name1862 (
		_w3747_,
		_w3751_,
		_w3762_,
		_w3763_
	);
	LUT4 #(
		.INIT('h00f7)
	) name1863 (
		\m3_s3_cyc_o_reg/NET0131 ,
		\rf_conf3_reg[6]/NET0131 ,
		\rf_conf3_reg[7]/NET0131 ,
		\s3_msel_arb1_state_reg[2]/NET0131 ,
		_w3764_
	);
	LUT4 #(
		.INIT('h0008)
	) name1864 (
		\m0_s3_cyc_o_reg/NET0131 ,
		\rf_conf3_reg[0]/NET0131 ,
		\rf_conf3_reg[1]/NET0131 ,
		\s3_msel_arb1_state_reg[0]/NET0131 ,
		_w3765_
	);
	LUT2 #(
		.INIT('h1)
	) name1865 (
		_w3747_,
		_w3765_,
		_w3766_
	);
	LUT3 #(
		.INIT('h54)
	) name1866 (
		\s3_msel_arb1_state_reg[1]/NET0131 ,
		_w3756_,
		_w3759_,
		_w3767_
	);
	LUT4 #(
		.INIT('h0040)
	) name1867 (
		_w3755_,
		_w3764_,
		_w3766_,
		_w3767_,
		_w3768_
	);
	LUT4 #(
		.INIT('h0008)
	) name1868 (
		\m4_s3_cyc_o_reg/NET0131 ,
		\rf_conf3_reg[8]/NET0131 ,
		\rf_conf3_reg[9]/NET0131 ,
		\s3_msel_arb1_state_reg[0]/NET0131 ,
		_w3769_
	);
	LUT4 #(
		.INIT('h5554)
	) name1869 (
		\s3_msel_arb1_state_reg[1]/NET0131 ,
		_w3749_,
		_w3753_,
		_w3769_,
		_w3770_
	);
	LUT4 #(
		.INIT('h0001)
	) name1870 (
		_w3756_,
		_w3757_,
		_w3759_,
		_w3760_,
		_w3771_
	);
	LUT3 #(
		.INIT('hb0)
	) name1871 (
		\s3_msel_arb1_state_reg[0]/NET0131 ,
		\s3_msel_arb1_state_reg[1]/NET0131 ,
		\s3_msel_arb1_state_reg[2]/NET0131 ,
		_w3772_
	);
	LUT4 #(
		.INIT('hfe00)
	) name1872 (
		_w3748_,
		_w3770_,
		_w3771_,
		_w3772_,
		_w3773_
	);
	LUT2 #(
		.INIT('h1)
	) name1873 (
		_w3768_,
		_w3773_,
		_w3774_
	);
	LUT2 #(
		.INIT('hb)
	) name1874 (
		_w3763_,
		_w3774_,
		_w3775_
	);
	LUT3 #(
		.INIT('h08)
	) name1875 (
		\m6_s4_cyc_o_reg/NET0131 ,
		\rf_conf4_reg[12]/NET0131 ,
		\rf_conf4_reg[13]/NET0131 ,
		_w3776_
	);
	LUT3 #(
		.INIT('h08)
	) name1876 (
		\m7_s4_cyc_o_reg/NET0131 ,
		\rf_conf4_reg[14]/NET0131 ,
		\rf_conf4_reg[15]/NET0131 ,
		_w3777_
	);
	LUT2 #(
		.INIT('h1)
	) name1877 (
		_w3776_,
		_w3777_,
		_w3778_
	);
	LUT3 #(
		.INIT('h08)
	) name1878 (
		\m4_s4_cyc_o_reg/NET0131 ,
		\rf_conf4_reg[8]/NET0131 ,
		\rf_conf4_reg[9]/NET0131 ,
		_w3779_
	);
	LUT3 #(
		.INIT('h08)
	) name1879 (
		\m5_s4_cyc_o_reg/NET0131 ,
		\rf_conf4_reg[10]/NET0131 ,
		\rf_conf4_reg[11]/NET0131 ,
		_w3780_
	);
	LUT4 #(
		.INIT('h0001)
	) name1880 (
		_w3776_,
		_w3777_,
		_w3779_,
		_w3780_,
		_w3781_
	);
	LUT2 #(
		.INIT('h4)
	) name1881 (
		\s4_msel_arb1_state_reg[1]/NET0131 ,
		\s4_msel_arb1_state_reg[2]/NET0131 ,
		_w3782_
	);
	LUT3 #(
		.INIT('h10)
	) name1882 (
		\s4_msel_arb1_state_reg[0]/NET0131 ,
		\s4_msel_arb1_state_reg[1]/NET0131 ,
		\s4_msel_arb1_state_reg[2]/NET0131 ,
		_w3783_
	);
	LUT3 #(
		.INIT('h08)
	) name1883 (
		\m3_s4_cyc_o_reg/NET0131 ,
		\rf_conf4_reg[6]/NET0131 ,
		\rf_conf4_reg[7]/NET0131 ,
		_w3784_
	);
	LUT4 #(
		.INIT('h00f7)
	) name1884 (
		\m3_s4_cyc_o_reg/NET0131 ,
		\rf_conf4_reg[6]/NET0131 ,
		\rf_conf4_reg[7]/NET0131 ,
		\s4_msel_arb1_state_reg[2]/NET0131 ,
		_w3785_
	);
	LUT2 #(
		.INIT('h1)
	) name1885 (
		_w3783_,
		_w3785_,
		_w3786_
	);
	LUT4 #(
		.INIT('h0008)
	) name1886 (
		\m0_s4_cyc_o_reg/NET0131 ,
		\rf_conf4_reg[0]/NET0131 ,
		\rf_conf4_reg[1]/NET0131 ,
		\s4_msel_arb1_state_reg[0]/NET0131 ,
		_w3787_
	);
	LUT3 #(
		.INIT('h08)
	) name1887 (
		\m2_s4_cyc_o_reg/NET0131 ,
		\rf_conf4_reg[4]/NET0131 ,
		\rf_conf4_reg[5]/NET0131 ,
		_w3788_
	);
	LUT3 #(
		.INIT('h08)
	) name1888 (
		\m1_s4_cyc_o_reg/NET0131 ,
		\rf_conf4_reg[2]/NET0131 ,
		\rf_conf4_reg[3]/NET0131 ,
		_w3789_
	);
	LUT3 #(
		.INIT('h01)
	) name1889 (
		_w3787_,
		_w3788_,
		_w3789_,
		_w3790_
	);
	LUT4 #(
		.INIT('h0008)
	) name1890 (
		\m2_s4_cyc_o_reg/NET0131 ,
		\rf_conf4_reg[4]/NET0131 ,
		\rf_conf4_reg[5]/NET0131 ,
		\s4_msel_arb1_state_reg[0]/NET0131 ,
		_w3791_
	);
	LUT3 #(
		.INIT('h31)
	) name1891 (
		\s4_msel_arb1_state_reg[1]/NET0131 ,
		_w3783_,
		_w3791_,
		_w3792_
	);
	LUT4 #(
		.INIT('h1011)
	) name1892 (
		_w3781_,
		_w3786_,
		_w3790_,
		_w3792_,
		_w3793_
	);
	LUT3 #(
		.INIT('h08)
	) name1893 (
		\m0_s4_cyc_o_reg/NET0131 ,
		\rf_conf4_reg[0]/NET0131 ,
		\rf_conf4_reg[1]/NET0131 ,
		_w3794_
	);
	LUT2 #(
		.INIT('h1)
	) name1894 (
		_w3784_,
		_w3788_,
		_w3795_
	);
	LUT4 #(
		.INIT('h0001)
	) name1895 (
		_w3784_,
		_w3788_,
		_w3789_,
		_w3794_,
		_w3796_
	);
	LUT4 #(
		.INIT('h1115)
	) name1896 (
		\s4_msel_arb1_state_reg[0]/NET0131 ,
		\s4_msel_arb1_state_reg[1]/NET0131 ,
		_w3776_,
		_w3777_,
		_w3797_
	);
	LUT2 #(
		.INIT('h8)
	) name1897 (
		\s4_msel_arb1_state_reg[0]/NET0131 ,
		\s4_msel_arb1_state_reg[1]/NET0131 ,
		_w3798_
	);
	LUT4 #(
		.INIT('h3301)
	) name1898 (
		_w3776_,
		_w3777_,
		_w3780_,
		_w3798_,
		_w3799_
	);
	LUT4 #(
		.INIT('h888a)
	) name1899 (
		\s4_msel_arb1_state_reg[2]/NET0131 ,
		_w3796_,
		_w3797_,
		_w3799_,
		_w3800_
	);
	LUT2 #(
		.INIT('he)
	) name1900 (
		_w3793_,
		_w3800_,
		_w3801_
	);
	LUT3 #(
		.INIT('h08)
	) name1901 (
		\m3_s5_cyc_o_reg/NET0131 ,
		\rf_conf5_reg[6]/NET0131 ,
		\rf_conf5_reg[7]/NET0131 ,
		_w3802_
	);
	LUT3 #(
		.INIT('h08)
	) name1902 (
		\m2_s5_cyc_o_reg/NET0131 ,
		\rf_conf5_reg[4]/NET0131 ,
		\rf_conf5_reg[5]/NET0131 ,
		_w3803_
	);
	LUT2 #(
		.INIT('h1)
	) name1903 (
		_w3802_,
		_w3803_,
		_w3804_
	);
	LUT3 #(
		.INIT('h08)
	) name1904 (
		\m0_s5_cyc_o_reg/NET0131 ,
		\rf_conf5_reg[0]/NET0131 ,
		\rf_conf5_reg[1]/NET0131 ,
		_w3805_
	);
	LUT3 #(
		.INIT('h08)
	) name1905 (
		\m1_s5_cyc_o_reg/NET0131 ,
		\rf_conf5_reg[2]/NET0131 ,
		\rf_conf5_reg[3]/NET0131 ,
		_w3806_
	);
	LUT3 #(
		.INIT('h02)
	) name1906 (
		\s5_msel_arb1_state_reg[2]/NET0131 ,
		_w3805_,
		_w3806_,
		_w3807_
	);
	LUT3 #(
		.INIT('h08)
	) name1907 (
		\m7_s5_cyc_o_reg/NET0131 ,
		\rf_conf5_reg[14]/NET0131 ,
		\rf_conf5_reg[15]/NET0131 ,
		_w3808_
	);
	LUT3 #(
		.INIT('h08)
	) name1908 (
		\m6_s5_cyc_o_reg/NET0131 ,
		\rf_conf5_reg[12]/NET0131 ,
		\rf_conf5_reg[13]/NET0131 ,
		_w3809_
	);
	LUT2 #(
		.INIT('h1)
	) name1909 (
		_w3808_,
		_w3809_,
		_w3810_
	);
	LUT3 #(
		.INIT('h08)
	) name1910 (
		\m4_s5_cyc_o_reg/NET0131 ,
		\rf_conf5_reg[8]/NET0131 ,
		\rf_conf5_reg[9]/NET0131 ,
		_w3811_
	);
	LUT3 #(
		.INIT('h08)
	) name1911 (
		\m5_s5_cyc_o_reg/NET0131 ,
		\rf_conf5_reg[10]/NET0131 ,
		\rf_conf5_reg[11]/NET0131 ,
		_w3812_
	);
	LUT4 #(
		.INIT('h0001)
	) name1912 (
		_w3808_,
		_w3809_,
		_w3811_,
		_w3812_,
		_w3813_
	);
	LUT2 #(
		.INIT('h1)
	) name1913 (
		\s5_msel_arb1_state_reg[1]/NET0131 ,
		\s5_msel_arb1_state_reg[2]/NET0131 ,
		_w3814_
	);
	LUT2 #(
		.INIT('h4)
	) name1914 (
		_w3806_,
		_w3814_,
		_w3815_
	);
	LUT4 #(
		.INIT('h7577)
	) name1915 (
		_w3804_,
		_w3807_,
		_w3813_,
		_w3815_,
		_w3816_
	);
	LUT4 #(
		.INIT('h0800)
	) name1916 (
		\m7_s5_cyc_o_reg/NET0131 ,
		\rf_conf5_reg[14]/NET0131 ,
		\rf_conf5_reg[15]/NET0131 ,
		\s5_msel_arb1_state_reg[2]/NET0131 ,
		_w3817_
	);
	LUT2 #(
		.INIT('h4)
	) name1917 (
		\s5_msel_arb1_state_reg[1]/NET0131 ,
		\s5_msel_arb1_state_reg[2]/NET0131 ,
		_w3818_
	);
	LUT4 #(
		.INIT('h010f)
	) name1918 (
		_w3809_,
		_w3812_,
		_w3817_,
		_w3818_,
		_w3819_
	);
	LUT3 #(
		.INIT('h2a)
	) name1919 (
		\s5_msel_arb1_state_reg[0]/NET0131 ,
		_w3816_,
		_w3819_,
		_w3820_
	);
	LUT2 #(
		.INIT('h2)
	) name1920 (
		\s5_msel_arb1_state_reg[1]/NET0131 ,
		\s5_msel_arb1_state_reg[2]/NET0131 ,
		_w3821_
	);
	LUT4 #(
		.INIT('h00fe)
	) name1921 (
		\s5_msel_arb1_state_reg[0]/NET0131 ,
		_w3805_,
		_w3806_,
		_w3821_,
		_w3822_
	);
	LUT4 #(
		.INIT('h0008)
	) name1922 (
		\m2_s5_cyc_o_reg/NET0131 ,
		\rf_conf5_reg[4]/NET0131 ,
		\rf_conf5_reg[5]/NET0131 ,
		\s5_msel_arb1_state_reg[0]/NET0131 ,
		_w3823_
	);
	LUT2 #(
		.INIT('h1)
	) name1923 (
		_w3802_,
		_w3823_,
		_w3824_
	);
	LUT4 #(
		.INIT('h0b00)
	) name1924 (
		\s5_msel_arb1_state_reg[2]/NET0131 ,
		_w3813_,
		_w3822_,
		_w3824_,
		_w3825_
	);
	LUT2 #(
		.INIT('h4)
	) name1925 (
		\s5_msel_arb1_state_reg[0]/NET0131 ,
		\s5_msel_arb1_state_reg[2]/NET0131 ,
		_w3826_
	);
	LUT3 #(
		.INIT('he0)
	) name1926 (
		_w3808_,
		_w3809_,
		_w3826_,
		_w3827_
	);
	LUT3 #(
		.INIT('h10)
	) name1927 (
		\s5_msel_arb1_state_reg[0]/NET0131 ,
		\s5_msel_arb1_state_reg[1]/NET0131 ,
		\s5_msel_arb1_state_reg[2]/NET0131 ,
		_w3828_
	);
	LUT3 #(
		.INIT('he0)
	) name1928 (
		_w3811_,
		_w3812_,
		_w3828_,
		_w3829_
	);
	LUT2 #(
		.INIT('h1)
	) name1929 (
		_w3827_,
		_w3829_,
		_w3830_
	);
	LUT2 #(
		.INIT('h4)
	) name1930 (
		_w3825_,
		_w3830_,
		_w3831_
	);
	LUT2 #(
		.INIT('hb)
	) name1931 (
		_w3820_,
		_w3831_,
		_w3832_
	);
	LUT3 #(
		.INIT('h08)
	) name1932 (
		\m3_s6_cyc_o_reg/NET0131 ,
		\rf_conf6_reg[6]/NET0131 ,
		\rf_conf6_reg[7]/NET0131 ,
		_w3833_
	);
	LUT3 #(
		.INIT('h08)
	) name1933 (
		\m2_s6_cyc_o_reg/NET0131 ,
		\rf_conf6_reg[4]/NET0131 ,
		\rf_conf6_reg[5]/NET0131 ,
		_w3834_
	);
	LUT2 #(
		.INIT('h1)
	) name1934 (
		_w3833_,
		_w3834_,
		_w3835_
	);
	LUT3 #(
		.INIT('h08)
	) name1935 (
		\m0_s6_cyc_o_reg/NET0131 ,
		\rf_conf6_reg[0]/NET0131 ,
		\rf_conf6_reg[1]/NET0131 ,
		_w3836_
	);
	LUT3 #(
		.INIT('h08)
	) name1936 (
		\m1_s6_cyc_o_reg/NET0131 ,
		\rf_conf6_reg[2]/NET0131 ,
		\rf_conf6_reg[3]/NET0131 ,
		_w3837_
	);
	LUT3 #(
		.INIT('h02)
	) name1937 (
		\s6_msel_arb1_state_reg[2]/NET0131 ,
		_w3836_,
		_w3837_,
		_w3838_
	);
	LUT3 #(
		.INIT('h08)
	) name1938 (
		\m7_s6_cyc_o_reg/NET0131 ,
		\rf_conf6_reg[14]/NET0131 ,
		\rf_conf6_reg[15]/NET0131 ,
		_w3839_
	);
	LUT3 #(
		.INIT('h08)
	) name1939 (
		\m6_s6_cyc_o_reg/NET0131 ,
		\rf_conf6_reg[12]/NET0131 ,
		\rf_conf6_reg[13]/NET0131 ,
		_w3840_
	);
	LUT2 #(
		.INIT('h1)
	) name1940 (
		_w3839_,
		_w3840_,
		_w3841_
	);
	LUT3 #(
		.INIT('h08)
	) name1941 (
		\m4_s6_cyc_o_reg/NET0131 ,
		\rf_conf6_reg[8]/NET0131 ,
		\rf_conf6_reg[9]/NET0131 ,
		_w3842_
	);
	LUT3 #(
		.INIT('h08)
	) name1942 (
		\m5_s6_cyc_o_reg/NET0131 ,
		\rf_conf6_reg[10]/NET0131 ,
		\rf_conf6_reg[11]/NET0131 ,
		_w3843_
	);
	LUT4 #(
		.INIT('h0001)
	) name1943 (
		_w3839_,
		_w3840_,
		_w3842_,
		_w3843_,
		_w3844_
	);
	LUT2 #(
		.INIT('h1)
	) name1944 (
		\s6_msel_arb1_state_reg[1]/NET0131 ,
		\s6_msel_arb1_state_reg[2]/NET0131 ,
		_w3845_
	);
	LUT2 #(
		.INIT('h4)
	) name1945 (
		_w3837_,
		_w3845_,
		_w3846_
	);
	LUT4 #(
		.INIT('h7577)
	) name1946 (
		_w3835_,
		_w3838_,
		_w3844_,
		_w3846_,
		_w3847_
	);
	LUT4 #(
		.INIT('h0800)
	) name1947 (
		\m7_s6_cyc_o_reg/NET0131 ,
		\rf_conf6_reg[14]/NET0131 ,
		\rf_conf6_reg[15]/NET0131 ,
		\s6_msel_arb1_state_reg[2]/NET0131 ,
		_w3848_
	);
	LUT2 #(
		.INIT('h4)
	) name1948 (
		\s6_msel_arb1_state_reg[1]/NET0131 ,
		\s6_msel_arb1_state_reg[2]/NET0131 ,
		_w3849_
	);
	LUT4 #(
		.INIT('h010f)
	) name1949 (
		_w3840_,
		_w3843_,
		_w3848_,
		_w3849_,
		_w3850_
	);
	LUT3 #(
		.INIT('h2a)
	) name1950 (
		\s6_msel_arb1_state_reg[0]/NET0131 ,
		_w3847_,
		_w3850_,
		_w3851_
	);
	LUT2 #(
		.INIT('h2)
	) name1951 (
		\s6_msel_arb1_state_reg[1]/NET0131 ,
		\s6_msel_arb1_state_reg[2]/NET0131 ,
		_w3852_
	);
	LUT4 #(
		.INIT('h00fe)
	) name1952 (
		\s6_msel_arb1_state_reg[0]/NET0131 ,
		_w3836_,
		_w3837_,
		_w3852_,
		_w3853_
	);
	LUT4 #(
		.INIT('h0008)
	) name1953 (
		\m2_s6_cyc_o_reg/NET0131 ,
		\rf_conf6_reg[4]/NET0131 ,
		\rf_conf6_reg[5]/NET0131 ,
		\s6_msel_arb1_state_reg[0]/NET0131 ,
		_w3854_
	);
	LUT2 #(
		.INIT('h1)
	) name1954 (
		_w3833_,
		_w3854_,
		_w3855_
	);
	LUT4 #(
		.INIT('h0b00)
	) name1955 (
		\s6_msel_arb1_state_reg[2]/NET0131 ,
		_w3844_,
		_w3853_,
		_w3855_,
		_w3856_
	);
	LUT2 #(
		.INIT('h4)
	) name1956 (
		\s6_msel_arb1_state_reg[0]/NET0131 ,
		\s6_msel_arb1_state_reg[2]/NET0131 ,
		_w3857_
	);
	LUT3 #(
		.INIT('he0)
	) name1957 (
		_w3839_,
		_w3840_,
		_w3857_,
		_w3858_
	);
	LUT3 #(
		.INIT('h10)
	) name1958 (
		\s6_msel_arb1_state_reg[0]/NET0131 ,
		\s6_msel_arb1_state_reg[1]/NET0131 ,
		\s6_msel_arb1_state_reg[2]/NET0131 ,
		_w3859_
	);
	LUT3 #(
		.INIT('he0)
	) name1959 (
		_w3842_,
		_w3843_,
		_w3859_,
		_w3860_
	);
	LUT2 #(
		.INIT('h1)
	) name1960 (
		_w3858_,
		_w3860_,
		_w3861_
	);
	LUT2 #(
		.INIT('h4)
	) name1961 (
		_w3856_,
		_w3861_,
		_w3862_
	);
	LUT2 #(
		.INIT('hb)
	) name1962 (
		_w3851_,
		_w3862_,
		_w3863_
	);
	LUT3 #(
		.INIT('h08)
	) name1963 (
		\m1_s7_cyc_o_reg/NET0131 ,
		\rf_conf7_reg[2]/NET0131 ,
		\rf_conf7_reg[3]/NET0131 ,
		_w3864_
	);
	LUT3 #(
		.INIT('h08)
	) name1964 (
		\m0_s7_cyc_o_reg/NET0131 ,
		\rf_conf7_reg[0]/NET0131 ,
		\rf_conf7_reg[1]/NET0131 ,
		_w3865_
	);
	LUT2 #(
		.INIT('h1)
	) name1965 (
		_w3864_,
		_w3865_,
		_w3866_
	);
	LUT3 #(
		.INIT('h08)
	) name1966 (
		\m3_s7_cyc_o_reg/NET0131 ,
		\rf_conf7_reg[6]/NET0131 ,
		\rf_conf7_reg[7]/NET0131 ,
		_w3867_
	);
	LUT3 #(
		.INIT('h08)
	) name1967 (
		\m2_s7_cyc_o_reg/NET0131 ,
		\rf_conf7_reg[4]/NET0131 ,
		\rf_conf7_reg[5]/NET0131 ,
		_w3868_
	);
	LUT2 #(
		.INIT('h1)
	) name1968 (
		_w3867_,
		_w3868_,
		_w3869_
	);
	LUT4 #(
		.INIT('h0001)
	) name1969 (
		_w3864_,
		_w3865_,
		_w3867_,
		_w3868_,
		_w3870_
	);
	LUT3 #(
		.INIT('h08)
	) name1970 (
		\m5_s7_cyc_o_reg/NET0131 ,
		\rf_conf7_reg[10]/NET0131 ,
		\rf_conf7_reg[11]/NET0131 ,
		_w3871_
	);
	LUT3 #(
		.INIT('h08)
	) name1971 (
		\m4_s7_cyc_o_reg/NET0131 ,
		\rf_conf7_reg[8]/NET0131 ,
		\rf_conf7_reg[9]/NET0131 ,
		_w3872_
	);
	LUT2 #(
		.INIT('h1)
	) name1972 (
		_w3871_,
		_w3872_,
		_w3873_
	);
	LUT3 #(
		.INIT('h08)
	) name1973 (
		\m7_s7_cyc_o_reg/NET0131 ,
		\rf_conf7_reg[14]/NET0131 ,
		\rf_conf7_reg[15]/NET0131 ,
		_w3874_
	);
	LUT3 #(
		.INIT('h08)
	) name1974 (
		\m6_s7_cyc_o_reg/NET0131 ,
		\rf_conf7_reg[12]/NET0131 ,
		\rf_conf7_reg[13]/NET0131 ,
		_w3875_
	);
	LUT4 #(
		.INIT('h0001)
	) name1975 (
		_w3871_,
		_w3872_,
		_w3874_,
		_w3875_,
		_w3876_
	);
	LUT2 #(
		.INIT('h1)
	) name1976 (
		\s7_msel_arb1_state_reg[0]/NET0131 ,
		\s7_msel_arb1_state_reg[1]/NET0131 ,
		_w3877_
	);
	LUT3 #(
		.INIT('h40)
	) name1977 (
		_w3870_,
		_w3876_,
		_w3877_,
		_w3878_
	);
	LUT4 #(
		.INIT('h0008)
	) name1978 (
		\m6_s7_cyc_o_reg/NET0131 ,
		\rf_conf7_reg[12]/NET0131 ,
		\rf_conf7_reg[13]/NET0131 ,
		\s7_msel_arb1_state_reg[0]/NET0131 ,
		_w3879_
	);
	LUT4 #(
		.INIT('hf700)
	) name1979 (
		\m6_s7_cyc_o_reg/NET0131 ,
		\rf_conf7_reg[12]/NET0131 ,
		\rf_conf7_reg[13]/NET0131 ,
		\s7_msel_arb1_state_reg[0]/NET0131 ,
		_w3880_
	);
	LUT4 #(
		.INIT('hc4f5)
	) name1980 (
		\s7_msel_arb1_state_reg[1]/NET0131 ,
		_w3871_,
		_w3879_,
		_w3880_,
		_w3881_
	);
	LUT4 #(
		.INIT('hf700)
	) name1981 (
		\m7_s7_cyc_o_reg/NET0131 ,
		\rf_conf7_reg[14]/NET0131 ,
		\rf_conf7_reg[15]/NET0131 ,
		\s7_msel_arb1_state_reg[2]/NET0131 ,
		_w3882_
	);
	LUT3 #(
		.INIT('h10)
	) name1982 (
		_w3870_,
		_w3881_,
		_w3882_,
		_w3883_
	);
	LUT4 #(
		.INIT('h0008)
	) name1983 (
		\m0_s7_cyc_o_reg/NET0131 ,
		\rf_conf7_reg[0]/NET0131 ,
		\rf_conf7_reg[1]/NET0131 ,
		\s7_msel_arb1_state_reg[0]/NET0131 ,
		_w3884_
	);
	LUT3 #(
		.INIT('h54)
	) name1984 (
		\s7_msel_arb1_state_reg[1]/NET0131 ,
		_w3864_,
		_w3884_,
		_w3885_
	);
	LUT2 #(
		.INIT('h8)
	) name1985 (
		\s7_msel_arb1_state_reg[0]/NET0131 ,
		\s7_msel_arb1_state_reg[1]/NET0131 ,
		_w3886_
	);
	LUT3 #(
		.INIT('h51)
	) name1986 (
		_w3867_,
		_w3868_,
		_w3886_,
		_w3887_
	);
	LUT4 #(
		.INIT('h5455)
	) name1987 (
		\s7_msel_arb1_state_reg[2]/NET0131 ,
		_w3876_,
		_w3885_,
		_w3887_,
		_w3888_
	);
	LUT3 #(
		.INIT('h01)
	) name1988 (
		_w3878_,
		_w3883_,
		_w3888_,
		_w3889_
	);
	LUT3 #(
		.INIT('h08)
	) name1989 (
		\m3_s8_cyc_o_reg/NET0131 ,
		\rf_conf8_reg[6]/NET0131 ,
		\rf_conf8_reg[7]/NET0131 ,
		_w3890_
	);
	LUT3 #(
		.INIT('h08)
	) name1990 (
		\m2_s8_cyc_o_reg/NET0131 ,
		\rf_conf8_reg[4]/NET0131 ,
		\rf_conf8_reg[5]/NET0131 ,
		_w3891_
	);
	LUT2 #(
		.INIT('h1)
	) name1991 (
		_w3890_,
		_w3891_,
		_w3892_
	);
	LUT3 #(
		.INIT('h08)
	) name1992 (
		\m0_s8_cyc_o_reg/NET0131 ,
		\rf_conf8_reg[0]/NET0131 ,
		\rf_conf8_reg[1]/NET0131 ,
		_w3893_
	);
	LUT3 #(
		.INIT('h08)
	) name1993 (
		\m1_s8_cyc_o_reg/NET0131 ,
		\rf_conf8_reg[2]/NET0131 ,
		\rf_conf8_reg[3]/NET0131 ,
		_w3894_
	);
	LUT3 #(
		.INIT('h02)
	) name1994 (
		\s8_msel_arb1_state_reg[2]/NET0131 ,
		_w3893_,
		_w3894_,
		_w3895_
	);
	LUT3 #(
		.INIT('h08)
	) name1995 (
		\m7_s8_cyc_o_reg/NET0131 ,
		\rf_conf8_reg[14]/NET0131 ,
		\rf_conf8_reg[15]/NET0131 ,
		_w3896_
	);
	LUT3 #(
		.INIT('h08)
	) name1996 (
		\m6_s8_cyc_o_reg/NET0131 ,
		\rf_conf8_reg[12]/NET0131 ,
		\rf_conf8_reg[13]/NET0131 ,
		_w3897_
	);
	LUT2 #(
		.INIT('h1)
	) name1997 (
		_w3896_,
		_w3897_,
		_w3898_
	);
	LUT3 #(
		.INIT('h08)
	) name1998 (
		\m4_s8_cyc_o_reg/NET0131 ,
		\rf_conf8_reg[8]/NET0131 ,
		\rf_conf8_reg[9]/NET0131 ,
		_w3899_
	);
	LUT3 #(
		.INIT('h08)
	) name1999 (
		\m5_s8_cyc_o_reg/NET0131 ,
		\rf_conf8_reg[10]/NET0131 ,
		\rf_conf8_reg[11]/NET0131 ,
		_w3900_
	);
	LUT4 #(
		.INIT('h0001)
	) name2000 (
		_w3896_,
		_w3897_,
		_w3899_,
		_w3900_,
		_w3901_
	);
	LUT2 #(
		.INIT('h1)
	) name2001 (
		\s8_msel_arb1_state_reg[1]/NET0131 ,
		\s8_msel_arb1_state_reg[2]/NET0131 ,
		_w3902_
	);
	LUT2 #(
		.INIT('h4)
	) name2002 (
		_w3894_,
		_w3902_,
		_w3903_
	);
	LUT4 #(
		.INIT('h7577)
	) name2003 (
		_w3892_,
		_w3895_,
		_w3901_,
		_w3903_,
		_w3904_
	);
	LUT4 #(
		.INIT('h0800)
	) name2004 (
		\m7_s8_cyc_o_reg/NET0131 ,
		\rf_conf8_reg[14]/NET0131 ,
		\rf_conf8_reg[15]/NET0131 ,
		\s8_msel_arb1_state_reg[2]/NET0131 ,
		_w3905_
	);
	LUT2 #(
		.INIT('h4)
	) name2005 (
		\s8_msel_arb1_state_reg[1]/NET0131 ,
		\s8_msel_arb1_state_reg[2]/NET0131 ,
		_w3906_
	);
	LUT4 #(
		.INIT('h010f)
	) name2006 (
		_w3897_,
		_w3900_,
		_w3905_,
		_w3906_,
		_w3907_
	);
	LUT3 #(
		.INIT('h2a)
	) name2007 (
		\s8_msel_arb1_state_reg[0]/NET0131 ,
		_w3904_,
		_w3907_,
		_w3908_
	);
	LUT2 #(
		.INIT('h2)
	) name2008 (
		\s8_msel_arb1_state_reg[1]/NET0131 ,
		\s8_msel_arb1_state_reg[2]/NET0131 ,
		_w3909_
	);
	LUT4 #(
		.INIT('h00fe)
	) name2009 (
		\s8_msel_arb1_state_reg[0]/NET0131 ,
		_w3893_,
		_w3894_,
		_w3909_,
		_w3910_
	);
	LUT4 #(
		.INIT('h0008)
	) name2010 (
		\m2_s8_cyc_o_reg/NET0131 ,
		\rf_conf8_reg[4]/NET0131 ,
		\rf_conf8_reg[5]/NET0131 ,
		\s8_msel_arb1_state_reg[0]/NET0131 ,
		_w3911_
	);
	LUT2 #(
		.INIT('h1)
	) name2011 (
		_w3890_,
		_w3911_,
		_w3912_
	);
	LUT4 #(
		.INIT('h0b00)
	) name2012 (
		\s8_msel_arb1_state_reg[2]/NET0131 ,
		_w3901_,
		_w3910_,
		_w3912_,
		_w3913_
	);
	LUT2 #(
		.INIT('h4)
	) name2013 (
		\s8_msel_arb1_state_reg[0]/NET0131 ,
		\s8_msel_arb1_state_reg[2]/NET0131 ,
		_w3914_
	);
	LUT3 #(
		.INIT('he0)
	) name2014 (
		_w3896_,
		_w3897_,
		_w3914_,
		_w3915_
	);
	LUT3 #(
		.INIT('h10)
	) name2015 (
		\s8_msel_arb1_state_reg[0]/NET0131 ,
		\s8_msel_arb1_state_reg[1]/NET0131 ,
		\s8_msel_arb1_state_reg[2]/NET0131 ,
		_w3916_
	);
	LUT3 #(
		.INIT('he0)
	) name2016 (
		_w3899_,
		_w3900_,
		_w3916_,
		_w3917_
	);
	LUT2 #(
		.INIT('h1)
	) name2017 (
		_w3915_,
		_w3917_,
		_w3918_
	);
	LUT2 #(
		.INIT('h4)
	) name2018 (
		_w3913_,
		_w3918_,
		_w3919_
	);
	LUT2 #(
		.INIT('hb)
	) name2019 (
		_w3908_,
		_w3919_,
		_w3920_
	);
	LUT3 #(
		.INIT('h08)
	) name2020 (
		\m3_s9_cyc_o_reg/NET0131 ,
		\rf_conf9_reg[6]/NET0131 ,
		\rf_conf9_reg[7]/NET0131 ,
		_w3921_
	);
	LUT3 #(
		.INIT('h08)
	) name2021 (
		\m2_s9_cyc_o_reg/NET0131 ,
		\rf_conf9_reg[4]/NET0131 ,
		\rf_conf9_reg[5]/NET0131 ,
		_w3922_
	);
	LUT2 #(
		.INIT('h1)
	) name2022 (
		_w3921_,
		_w3922_,
		_w3923_
	);
	LUT3 #(
		.INIT('h08)
	) name2023 (
		\m0_s9_cyc_o_reg/NET0131 ,
		\rf_conf9_reg[0]/NET0131 ,
		\rf_conf9_reg[1]/NET0131 ,
		_w3924_
	);
	LUT3 #(
		.INIT('h08)
	) name2024 (
		\m1_s9_cyc_o_reg/NET0131 ,
		\rf_conf9_reg[2]/NET0131 ,
		\rf_conf9_reg[3]/NET0131 ,
		_w3925_
	);
	LUT3 #(
		.INIT('h02)
	) name2025 (
		\s9_msel_arb1_state_reg[2]/NET0131 ,
		_w3924_,
		_w3925_,
		_w3926_
	);
	LUT3 #(
		.INIT('h08)
	) name2026 (
		\m7_s9_cyc_o_reg/NET0131 ,
		\rf_conf9_reg[14]/NET0131 ,
		\rf_conf9_reg[15]/NET0131 ,
		_w3927_
	);
	LUT3 #(
		.INIT('h08)
	) name2027 (
		\m6_s9_cyc_o_reg/NET0131 ,
		\rf_conf9_reg[12]/NET0131 ,
		\rf_conf9_reg[13]/NET0131 ,
		_w3928_
	);
	LUT2 #(
		.INIT('h1)
	) name2028 (
		_w3927_,
		_w3928_,
		_w3929_
	);
	LUT3 #(
		.INIT('h08)
	) name2029 (
		\m4_s9_cyc_o_reg/NET0131 ,
		\rf_conf9_reg[8]/NET0131 ,
		\rf_conf9_reg[9]/NET0131 ,
		_w3930_
	);
	LUT3 #(
		.INIT('h08)
	) name2030 (
		\m5_s9_cyc_o_reg/NET0131 ,
		\rf_conf9_reg[10]/NET0131 ,
		\rf_conf9_reg[11]/NET0131 ,
		_w3931_
	);
	LUT4 #(
		.INIT('h0001)
	) name2031 (
		_w3927_,
		_w3928_,
		_w3930_,
		_w3931_,
		_w3932_
	);
	LUT2 #(
		.INIT('h1)
	) name2032 (
		\s9_msel_arb1_state_reg[1]/NET0131 ,
		\s9_msel_arb1_state_reg[2]/NET0131 ,
		_w3933_
	);
	LUT2 #(
		.INIT('h4)
	) name2033 (
		_w3925_,
		_w3933_,
		_w3934_
	);
	LUT4 #(
		.INIT('h7577)
	) name2034 (
		_w3923_,
		_w3926_,
		_w3932_,
		_w3934_,
		_w3935_
	);
	LUT4 #(
		.INIT('h0800)
	) name2035 (
		\m7_s9_cyc_o_reg/NET0131 ,
		\rf_conf9_reg[14]/NET0131 ,
		\rf_conf9_reg[15]/NET0131 ,
		\s9_msel_arb1_state_reg[2]/NET0131 ,
		_w3936_
	);
	LUT2 #(
		.INIT('h4)
	) name2036 (
		\s9_msel_arb1_state_reg[1]/NET0131 ,
		\s9_msel_arb1_state_reg[2]/NET0131 ,
		_w3937_
	);
	LUT4 #(
		.INIT('h010f)
	) name2037 (
		_w3928_,
		_w3931_,
		_w3936_,
		_w3937_,
		_w3938_
	);
	LUT3 #(
		.INIT('h2a)
	) name2038 (
		\s9_msel_arb1_state_reg[0]/NET0131 ,
		_w3935_,
		_w3938_,
		_w3939_
	);
	LUT2 #(
		.INIT('h2)
	) name2039 (
		\s9_msel_arb1_state_reg[1]/NET0131 ,
		\s9_msel_arb1_state_reg[2]/NET0131 ,
		_w3940_
	);
	LUT4 #(
		.INIT('h00fe)
	) name2040 (
		\s9_msel_arb1_state_reg[0]/NET0131 ,
		_w3924_,
		_w3925_,
		_w3940_,
		_w3941_
	);
	LUT4 #(
		.INIT('h0008)
	) name2041 (
		\m2_s9_cyc_o_reg/NET0131 ,
		\rf_conf9_reg[4]/NET0131 ,
		\rf_conf9_reg[5]/NET0131 ,
		\s9_msel_arb1_state_reg[0]/NET0131 ,
		_w3942_
	);
	LUT2 #(
		.INIT('h1)
	) name2042 (
		_w3921_,
		_w3942_,
		_w3943_
	);
	LUT4 #(
		.INIT('h0b00)
	) name2043 (
		\s9_msel_arb1_state_reg[2]/NET0131 ,
		_w3932_,
		_w3941_,
		_w3943_,
		_w3944_
	);
	LUT2 #(
		.INIT('h4)
	) name2044 (
		\s9_msel_arb1_state_reg[0]/NET0131 ,
		\s9_msel_arb1_state_reg[2]/NET0131 ,
		_w3945_
	);
	LUT3 #(
		.INIT('he0)
	) name2045 (
		_w3927_,
		_w3928_,
		_w3945_,
		_w3946_
	);
	LUT3 #(
		.INIT('h10)
	) name2046 (
		\s9_msel_arb1_state_reg[0]/NET0131 ,
		\s9_msel_arb1_state_reg[1]/NET0131 ,
		\s9_msel_arb1_state_reg[2]/NET0131 ,
		_w3947_
	);
	LUT3 #(
		.INIT('he0)
	) name2047 (
		_w3930_,
		_w3931_,
		_w3947_,
		_w3948_
	);
	LUT2 #(
		.INIT('h1)
	) name2048 (
		_w3946_,
		_w3948_,
		_w3949_
	);
	LUT2 #(
		.INIT('h4)
	) name2049 (
		_w3944_,
		_w3949_,
		_w3950_
	);
	LUT2 #(
		.INIT('hb)
	) name2050 (
		_w3939_,
		_w3950_,
		_w3951_
	);
	LUT3 #(
		.INIT('h08)
	) name2051 (
		\m3_s0_cyc_o_reg/NET0131 ,
		\rf_conf0_reg[6]/NET0131 ,
		\rf_conf0_reg[7]/NET0131 ,
		_w3952_
	);
	LUT3 #(
		.INIT('h08)
	) name2052 (
		\m2_s0_cyc_o_reg/NET0131 ,
		\rf_conf0_reg[4]/NET0131 ,
		\rf_conf0_reg[5]/NET0131 ,
		_w3953_
	);
	LUT2 #(
		.INIT('h1)
	) name2053 (
		_w3952_,
		_w3953_,
		_w3954_
	);
	LUT3 #(
		.INIT('h08)
	) name2054 (
		\m0_s0_cyc_o_reg/NET0131 ,
		\rf_conf0_reg[0]/NET0131 ,
		\rf_conf0_reg[1]/NET0131 ,
		_w3955_
	);
	LUT3 #(
		.INIT('h08)
	) name2055 (
		\m1_s0_cyc_o_reg/NET0131 ,
		\rf_conf0_reg[2]/NET0131 ,
		\rf_conf0_reg[3]/NET0131 ,
		_w3956_
	);
	LUT3 #(
		.INIT('h02)
	) name2056 (
		\s0_msel_arb1_state_reg[2]/NET0131 ,
		_w3955_,
		_w3956_,
		_w3957_
	);
	LUT3 #(
		.INIT('h08)
	) name2057 (
		\m7_s0_cyc_o_reg/NET0131 ,
		\rf_conf0_reg[14]/NET0131 ,
		\rf_conf0_reg[15]/NET0131 ,
		_w3958_
	);
	LUT3 #(
		.INIT('h08)
	) name2058 (
		\m6_s0_cyc_o_reg/NET0131 ,
		\rf_conf0_reg[12]/NET0131 ,
		\rf_conf0_reg[13]/NET0131 ,
		_w3959_
	);
	LUT2 #(
		.INIT('h1)
	) name2059 (
		_w3958_,
		_w3959_,
		_w3960_
	);
	LUT3 #(
		.INIT('h08)
	) name2060 (
		\m4_s0_cyc_o_reg/NET0131 ,
		\rf_conf0_reg[8]/NET0131 ,
		\rf_conf0_reg[9]/NET0131 ,
		_w3961_
	);
	LUT3 #(
		.INIT('h08)
	) name2061 (
		\m5_s0_cyc_o_reg/NET0131 ,
		\rf_conf0_reg[10]/NET0131 ,
		\rf_conf0_reg[11]/NET0131 ,
		_w3962_
	);
	LUT4 #(
		.INIT('h0001)
	) name2062 (
		_w3958_,
		_w3959_,
		_w3961_,
		_w3962_,
		_w3963_
	);
	LUT2 #(
		.INIT('h1)
	) name2063 (
		\s0_msel_arb1_state_reg[1]/NET0131 ,
		\s0_msel_arb1_state_reg[2]/NET0131 ,
		_w3964_
	);
	LUT2 #(
		.INIT('h4)
	) name2064 (
		_w3956_,
		_w3964_,
		_w3965_
	);
	LUT4 #(
		.INIT('h7577)
	) name2065 (
		_w3954_,
		_w3957_,
		_w3963_,
		_w3965_,
		_w3966_
	);
	LUT4 #(
		.INIT('h0800)
	) name2066 (
		\m7_s0_cyc_o_reg/NET0131 ,
		\rf_conf0_reg[14]/NET0131 ,
		\rf_conf0_reg[15]/NET0131 ,
		\s0_msel_arb1_state_reg[2]/NET0131 ,
		_w3967_
	);
	LUT2 #(
		.INIT('h4)
	) name2067 (
		\s0_msel_arb1_state_reg[1]/NET0131 ,
		\s0_msel_arb1_state_reg[2]/NET0131 ,
		_w3968_
	);
	LUT4 #(
		.INIT('h010f)
	) name2068 (
		_w3959_,
		_w3962_,
		_w3967_,
		_w3968_,
		_w3969_
	);
	LUT3 #(
		.INIT('h2a)
	) name2069 (
		\s0_msel_arb1_state_reg[0]/NET0131 ,
		_w3966_,
		_w3969_,
		_w3970_
	);
	LUT2 #(
		.INIT('h2)
	) name2070 (
		\s0_msel_arb1_state_reg[1]/NET0131 ,
		\s0_msel_arb1_state_reg[2]/NET0131 ,
		_w3971_
	);
	LUT4 #(
		.INIT('h00fe)
	) name2071 (
		\s0_msel_arb1_state_reg[0]/NET0131 ,
		_w3955_,
		_w3956_,
		_w3971_,
		_w3972_
	);
	LUT4 #(
		.INIT('h0008)
	) name2072 (
		\m2_s0_cyc_o_reg/NET0131 ,
		\rf_conf0_reg[4]/NET0131 ,
		\rf_conf0_reg[5]/NET0131 ,
		\s0_msel_arb1_state_reg[0]/NET0131 ,
		_w3973_
	);
	LUT2 #(
		.INIT('h1)
	) name2073 (
		_w3952_,
		_w3973_,
		_w3974_
	);
	LUT4 #(
		.INIT('h0b00)
	) name2074 (
		\s0_msel_arb1_state_reg[2]/NET0131 ,
		_w3963_,
		_w3972_,
		_w3974_,
		_w3975_
	);
	LUT2 #(
		.INIT('h4)
	) name2075 (
		\s0_msel_arb1_state_reg[0]/NET0131 ,
		\s0_msel_arb1_state_reg[2]/NET0131 ,
		_w3976_
	);
	LUT3 #(
		.INIT('he0)
	) name2076 (
		_w3958_,
		_w3959_,
		_w3976_,
		_w3977_
	);
	LUT3 #(
		.INIT('h10)
	) name2077 (
		\s0_msel_arb1_state_reg[0]/NET0131 ,
		\s0_msel_arb1_state_reg[1]/NET0131 ,
		\s0_msel_arb1_state_reg[2]/NET0131 ,
		_w3978_
	);
	LUT3 #(
		.INIT('he0)
	) name2078 (
		_w3961_,
		_w3962_,
		_w3978_,
		_w3979_
	);
	LUT2 #(
		.INIT('h1)
	) name2079 (
		_w3977_,
		_w3979_,
		_w3980_
	);
	LUT2 #(
		.INIT('h4)
	) name2080 (
		_w3975_,
		_w3980_,
		_w3981_
	);
	LUT2 #(
		.INIT('hb)
	) name2081 (
		_w3970_,
		_w3981_,
		_w3982_
	);
	LUT3 #(
		.INIT('h23)
	) name2082 (
		_w3559_,
		_w3561_,
		_w3571_,
		_w3983_
	);
	LUT4 #(
		.INIT('h2232)
	) name2083 (
		_w3559_,
		_w3561_,
		_w3570_,
		_w3571_,
		_w3984_
	);
	LUT2 #(
		.INIT('h1)
	) name2084 (
		_w3561_,
		_w3571_,
		_w3985_
	);
	LUT4 #(
		.INIT('h0004)
	) name2085 (
		_w3561_,
		_w3567_,
		_w3568_,
		_w3571_,
		_w3986_
	);
	LUT2 #(
		.INIT('h2)
	) name2086 (
		\s10_msel_arb1_state_reg[1]/NET0131 ,
		\s10_msel_arb1_state_reg[2]/NET0131 ,
		_w3987_
	);
	LUT2 #(
		.INIT('h4)
	) name2087 (
		_w3564_,
		_w3987_,
		_w3988_
	);
	LUT4 #(
		.INIT('hfe00)
	) name2088 (
		_w3565_,
		_w3984_,
		_w3986_,
		_w3988_,
		_w3989_
	);
	LUT3 #(
		.INIT('hdc)
	) name2089 (
		_w3559_,
		_w3561_,
		_w3571_,
		_w3990_
	);
	LUT2 #(
		.INIT('h2)
	) name2090 (
		_w3568_,
		_w3570_,
		_w3991_
	);
	LUT2 #(
		.INIT('h4)
	) name2091 (
		_w3564_,
		_w3565_,
		_w3992_
	);
	LUT4 #(
		.INIT('h000b)
	) name2092 (
		_w3564_,
		_w3565_,
		_w3567_,
		_w3570_,
		_w3993_
	);
	LUT4 #(
		.INIT('hf700)
	) name2093 (
		\m0_s10_cyc_o_reg/NET0131 ,
		\rf_conf10_reg[0]/NET0131 ,
		\rf_conf10_reg[1]/NET0131 ,
		\s10_msel_arb1_state_reg[0]/NET0131 ,
		_w3994_
	);
	LUT4 #(
		.INIT('hd0dd)
	) name2094 (
		_w3559_,
		_w3561_,
		_w3564_,
		_w3994_,
		_w3995_
	);
	LUT4 #(
		.INIT('h0155)
	) name2095 (
		_w3990_,
		_w3991_,
		_w3993_,
		_w3995_,
		_w3996_
	);
	LUT2 #(
		.INIT('h4)
	) name2096 (
		\s10_msel_arb1_state_reg[1]/NET0131 ,
		\s10_msel_arb1_state_reg[2]/NET0131 ,
		_w3997_
	);
	LUT4 #(
		.INIT('habbb)
	) name2097 (
		\s10_msel_arb1_state_reg[0]/NET0131 ,
		_w3989_,
		_w3996_,
		_w3997_,
		_w3998_
	);
	LUT4 #(
		.INIT('hff0d)
	) name2098 (
		\s10_msel_arb1_state_reg[0]/NET0131 ,
		_w3564_,
		_w3567_,
		_w3568_,
		_w3999_
	);
	LUT4 #(
		.INIT('h1101)
	) name2099 (
		_w3565_,
		_w3984_,
		_w3985_,
		_w3999_,
		_w4000_
	);
	LUT2 #(
		.INIT('h2)
	) name2100 (
		_w3987_,
		_w4000_,
		_w4001_
	);
	LUT2 #(
		.INIT('h1)
	) name2101 (
		\s10_msel_arb1_state_reg[1]/NET0131 ,
		\s10_msel_arb1_state_reg[2]/NET0131 ,
		_w4002_
	);
	LUT3 #(
		.INIT('h0b)
	) name2102 (
		_w3564_,
		_w3565_,
		_w3567_,
		_w4003_
	);
	LUT3 #(
		.INIT('h02)
	) name2103 (
		_w3559_,
		_w3561_,
		_w3564_,
		_w4004_
	);
	LUT3 #(
		.INIT('h01)
	) name2104 (
		_w3561_,
		_w3564_,
		_w3571_,
		_w4005_
	);
	LUT2 #(
		.INIT('h1)
	) name2105 (
		_w3570_,
		_w3994_,
		_w4006_
	);
	LUT4 #(
		.INIT('h2202)
	) name2106 (
		_w4003_,
		_w4004_,
		_w4005_,
		_w4006_,
		_w4007_
	);
	LUT4 #(
		.INIT('h5455)
	) name2107 (
		_w3559_,
		_w3561_,
		_w3564_,
		_w3994_,
		_w4008_
	);
	LUT3 #(
		.INIT('hb0)
	) name2108 (
		_w3559_,
		_w3571_,
		_w3997_,
		_w4009_
	);
	LUT4 #(
		.INIT('h1f00)
	) name2109 (
		_w3991_,
		_w3993_,
		_w4008_,
		_w4009_,
		_w4010_
	);
	LUT3 #(
		.INIT('h0d)
	) name2110 (
		_w4002_,
		_w4007_,
		_w4010_,
		_w4011_
	);
	LUT3 #(
		.INIT('h8a)
	) name2111 (
		\s10_msel_arb1_state_reg[0]/NET0131 ,
		_w4001_,
		_w4011_,
		_w4012_
	);
	LUT4 #(
		.INIT('h0008)
	) name2112 (
		\m6_s10_cyc_o_reg/NET0131 ,
		\rf_conf10_reg[12]/NET0131 ,
		\rf_conf10_reg[13]/NET0131 ,
		\s10_msel_arb1_state_reg[0]/NET0131 ,
		_w4013_
	);
	LUT2 #(
		.INIT('h8)
	) name2113 (
		\s10_msel_arb1_state_reg[1]/NET0131 ,
		\s10_msel_arb1_state_reg[2]/NET0131 ,
		_w4014_
	);
	LUT2 #(
		.INIT('h4)
	) name2114 (
		_w4013_,
		_w4014_,
		_w4015_
	);
	LUT3 #(
		.INIT('h20)
	) name2115 (
		_w3570_,
		_w4013_,
		_w4014_,
		_w4016_
	);
	LUT4 #(
		.INIT('hf700)
	) name2116 (
		\m2_s10_cyc_o_reg/NET0131 ,
		\rf_conf10_reg[4]/NET0131 ,
		\rf_conf10_reg[5]/NET0131 ,
		\s10_msel_arb1_state_reg[0]/NET0131 ,
		_w4017_
	);
	LUT3 #(
		.INIT('h10)
	) name2117 (
		_w3561_,
		_w3571_,
		_w4017_,
		_w4018_
	);
	LUT4 #(
		.INIT('hf0d0)
	) name2118 (
		_w4003_,
		_w4004_,
		_w4015_,
		_w4018_,
		_w4019_
	);
	LUT3 #(
		.INIT('h32)
	) name2119 (
		_w3559_,
		_w3564_,
		_w3570_,
		_w4020_
	);
	LUT4 #(
		.INIT('h0105)
	) name2120 (
		_w3567_,
		_w3983_,
		_w3992_,
		_w4020_,
		_w4021_
	);
	LUT3 #(
		.INIT('h01)
	) name2121 (
		\s10_msel_arb1_state_reg[0]/NET0131 ,
		\s10_msel_arb1_state_reg[1]/NET0131 ,
		\s10_msel_arb1_state_reg[2]/NET0131 ,
		_w4022_
	);
	LUT4 #(
		.INIT('hbabb)
	) name2122 (
		_w3568_,
		_w4019_,
		_w4021_,
		_w4022_,
		_w4023_
	);
	LUT2 #(
		.INIT('h4)
	) name2123 (
		_w4016_,
		_w4023_,
		_w4024_
	);
	LUT3 #(
		.INIT('hdf)
	) name2124 (
		_w3998_,
		_w4012_,
		_w4024_,
		_w4025_
	);
	LUT3 #(
		.INIT('h20)
	) name2125 (
		\m2_s10_cyc_o_reg/NET0131 ,
		\rf_conf10_reg[4]/NET0131 ,
		\rf_conf10_reg[5]/NET0131 ,
		_w4026_
	);
	LUT3 #(
		.INIT('h20)
	) name2126 (
		\m3_s10_cyc_o_reg/NET0131 ,
		\rf_conf10_reg[6]/NET0131 ,
		\rf_conf10_reg[7]/NET0131 ,
		_w4027_
	);
	LUT2 #(
		.INIT('h2)
	) name2127 (
		\s10_msel_arb2_state_reg[1]/NET0131 ,
		\s10_msel_arb2_state_reg[2]/NET0131 ,
		_w4028_
	);
	LUT3 #(
		.INIT('h40)
	) name2128 (
		_w4026_,
		_w4027_,
		_w4028_,
		_w4029_
	);
	LUT3 #(
		.INIT('h20)
	) name2129 (
		\m5_s10_cyc_o_reg/NET0131 ,
		\rf_conf10_reg[10]/NET0131 ,
		\rf_conf10_reg[11]/NET0131 ,
		_w4030_
	);
	LUT3 #(
		.INIT('h20)
	) name2130 (
		\m7_s10_cyc_o_reg/NET0131 ,
		\rf_conf10_reg[14]/NET0131 ,
		\rf_conf10_reg[15]/NET0131 ,
		_w4031_
	);
	LUT3 #(
		.INIT('h20)
	) name2131 (
		\m6_s10_cyc_o_reg/NET0131 ,
		\rf_conf10_reg[12]/NET0131 ,
		\rf_conf10_reg[13]/NET0131 ,
		_w4032_
	);
	LUT3 #(
		.INIT('h51)
	) name2132 (
		_w4030_,
		_w4031_,
		_w4032_,
		_w4033_
	);
	LUT3 #(
		.INIT('h20)
	) name2133 (
		\m1_s10_cyc_o_reg/NET0131 ,
		\rf_conf10_reg[2]/NET0131 ,
		\rf_conf10_reg[3]/NET0131 ,
		_w4034_
	);
	LUT3 #(
		.INIT('h20)
	) name2134 (
		\m0_s10_cyc_o_reg/NET0131 ,
		\rf_conf10_reg[0]/NET0131 ,
		\rf_conf10_reg[1]/NET0131 ,
		_w4035_
	);
	LUT2 #(
		.INIT('h1)
	) name2135 (
		_w4032_,
		_w4035_,
		_w4036_
	);
	LUT3 #(
		.INIT('h04)
	) name2136 (
		_w4032_,
		_w4034_,
		_w4035_,
		_w4037_
	);
	LUT3 #(
		.INIT('h20)
	) name2137 (
		\m4_s10_cyc_o_reg/NET0131 ,
		\rf_conf10_reg[8]/NET0131 ,
		\rf_conf10_reg[9]/NET0131 ,
		_w4038_
	);
	LUT2 #(
		.INIT('h1)
	) name2138 (
		_w4026_,
		_w4038_,
		_w4039_
	);
	LUT3 #(
		.INIT('h04)
	) name2139 (
		_w4026_,
		_w4028_,
		_w4038_,
		_w4040_
	);
	LUT4 #(
		.INIT('h0455)
	) name2140 (
		_w4029_,
		_w4033_,
		_w4037_,
		_w4040_,
		_w4041_
	);
	LUT3 #(
		.INIT('h0b)
	) name2141 (
		_w4026_,
		_w4027_,
		_w4034_,
		_w4042_
	);
	LUT2 #(
		.INIT('h1)
	) name2142 (
		\s10_msel_arb2_state_reg[1]/NET0131 ,
		\s10_msel_arb2_state_reg[2]/NET0131 ,
		_w4043_
	);
	LUT2 #(
		.INIT('h4)
	) name2143 (
		_w4035_,
		_w4043_,
		_w4044_
	);
	LUT4 #(
		.INIT('hb0ff)
	) name2144 (
		_w4033_,
		_w4039_,
		_w4042_,
		_w4044_,
		_w4045_
	);
	LUT3 #(
		.INIT('h40)
	) name2145 (
		\s10_msel_arb2_state_reg[0]/NET0131 ,
		_w4041_,
		_w4045_,
		_w4046_
	);
	LUT2 #(
		.INIT('h8)
	) name2146 (
		\s10_msel_arb2_state_reg[1]/NET0131 ,
		\s10_msel_arb2_state_reg[2]/NET0131 ,
		_w4047_
	);
	LUT3 #(
		.INIT('h20)
	) name2147 (
		_w4031_,
		_w4032_,
		_w4047_,
		_w4048_
	);
	LUT3 #(
		.INIT('h04)
	) name2148 (
		_w4026_,
		_w4030_,
		_w4038_,
		_w4049_
	);
	LUT3 #(
		.INIT('h10)
	) name2149 (
		_w4032_,
		_w4035_,
		_w4047_,
		_w4050_
	);
	LUT4 #(
		.INIT('h0233)
	) name2150 (
		_w4042_,
		_w4048_,
		_w4049_,
		_w4050_,
		_w4051_
	);
	LUT2 #(
		.INIT('h4)
	) name2151 (
		\s10_msel_arb2_state_reg[1]/NET0131 ,
		\s10_msel_arb2_state_reg[2]/NET0131 ,
		_w4052_
	);
	LUT3 #(
		.INIT('h20)
	) name2152 (
		_w4030_,
		_w4038_,
		_w4052_,
		_w4053_
	);
	LUT2 #(
		.INIT('h4)
	) name2153 (
		_w4031_,
		_w4035_,
		_w4054_
	);
	LUT4 #(
		.INIT('h000b)
	) name2154 (
		_w4026_,
		_w4027_,
		_w4031_,
		_w4034_,
		_w4055_
	);
	LUT3 #(
		.INIT('h10)
	) name2155 (
		_w4032_,
		_w4038_,
		_w4052_,
		_w4056_
	);
	LUT4 #(
		.INIT('h5455)
	) name2156 (
		_w4053_,
		_w4054_,
		_w4055_,
		_w4056_,
		_w4057_
	);
	LUT2 #(
		.INIT('h8)
	) name2157 (
		_w4051_,
		_w4057_,
		_w4058_
	);
	LUT4 #(
		.INIT('hdf00)
	) name2158 (
		\m0_s10_cyc_o_reg/NET0131 ,
		\rf_conf10_reg[0]/NET0131 ,
		\rf_conf10_reg[1]/NET0131 ,
		\s10_msel_arb2_state_reg[0]/NET0131 ,
		_w4059_
	);
	LUT3 #(
		.INIT('h10)
	) name2159 (
		_w4026_,
		_w4038_,
		_w4059_,
		_w4060_
	);
	LUT3 #(
		.INIT('h20)
	) name2160 (
		\s10_msel_arb2_state_reg[0]/NET0131 ,
		\s10_msel_arb2_state_reg[1]/NET0131 ,
		\s10_msel_arb2_state_reg[2]/NET0131 ,
		_w4061_
	);
	LUT3 #(
		.INIT('h10)
	) name2161 (
		_w4030_,
		_w4032_,
		_w4061_,
		_w4062_
	);
	LUT4 #(
		.INIT('hf100)
	) name2162 (
		_w4054_,
		_w4055_,
		_w4060_,
		_w4062_,
		_w4063_
	);
	LUT3 #(
		.INIT('h08)
	) name2163 (
		_w4046_,
		_w4058_,
		_w4063_,
		_w4064_
	);
	LUT3 #(
		.INIT('hb0)
	) name2164 (
		_w4033_,
		_w4039_,
		_w4042_,
		_w4065_
	);
	LUT3 #(
		.INIT('h02)
	) name2165 (
		\s10_msel_arb2_state_reg[0]/NET0131 ,
		_w4026_,
		_w4038_,
		_w4066_
	);
	LUT2 #(
		.INIT('h8)
	) name2166 (
		_w4036_,
		_w4066_,
		_w4067_
	);
	LUT3 #(
		.INIT('ha2)
	) name2167 (
		_w4043_,
		_w4065_,
		_w4067_,
		_w4068_
	);
	LUT2 #(
		.INIT('h8)
	) name2168 (
		_w4027_,
		_w4028_,
		_w4069_
	);
	LUT4 #(
		.INIT('h0031)
	) name2169 (
		_w4026_,
		_w4032_,
		_w4034_,
		_w4035_,
		_w4070_
	);
	LUT2 #(
		.INIT('h2)
	) name2170 (
		_w4028_,
		_w4038_,
		_w4071_
	);
	LUT4 #(
		.INIT('h0233)
	) name2171 (
		_w4033_,
		_w4069_,
		_w4070_,
		_w4071_,
		_w4072_
	);
	LUT3 #(
		.INIT('h2a)
	) name2172 (
		\s10_msel_arb2_state_reg[0]/NET0131 ,
		_w4030_,
		_w4052_,
		_w4073_
	);
	LUT2 #(
		.INIT('h8)
	) name2173 (
		_w4072_,
		_w4073_,
		_w4074_
	);
	LUT4 #(
		.INIT('hdf00)
	) name2174 (
		\m6_s10_cyc_o_reg/NET0131 ,
		\rf_conf10_reg[12]/NET0131 ,
		\rf_conf10_reg[13]/NET0131 ,
		\s10_msel_arb2_state_reg[0]/NET0131 ,
		_w4075_
	);
	LUT4 #(
		.INIT('h3233)
	) name2175 (
		_w4026_,
		_w4031_,
		_w4038_,
		_w4075_,
		_w4076_
	);
	LUT4 #(
		.INIT('h0d0f)
	) name2176 (
		_w4042_,
		_w4049_,
		_w4054_,
		_w4076_,
		_w4077_
	);
	LUT3 #(
		.INIT('h13)
	) name2177 (
		_w4047_,
		_w4063_,
		_w4077_,
		_w4078_
	);
	LUT3 #(
		.INIT('h40)
	) name2178 (
		_w4068_,
		_w4074_,
		_w4078_,
		_w4079_
	);
	LUT2 #(
		.INIT('h1)
	) name2179 (
		_w4064_,
		_w4079_,
		_w4080_
	);
	LUT2 #(
		.INIT('h2)
	) name2180 (
		\s10_msel_arb3_state_reg[1]/NET0131 ,
		\s10_msel_arb3_state_reg[2]/NET0131 ,
		_w4081_
	);
	LUT2 #(
		.INIT('h4)
	) name2181 (
		_w3171_,
		_w4081_,
		_w4082_
	);
	LUT2 #(
		.INIT('h1)
	) name2182 (
		_w3153_,
		_w3160_,
		_w4083_
	);
	LUT3 #(
		.INIT('hae)
	) name2183 (
		_w3153_,
		_w3160_,
		_w3161_,
		_w4084_
	);
	LUT2 #(
		.INIT('h1)
	) name2184 (
		_w3165_,
		_w3176_,
		_w4085_
	);
	LUT2 #(
		.INIT('h1)
	) name2185 (
		_w3161_,
		_w3166_,
		_w4086_
	);
	LUT4 #(
		.INIT('h7577)
	) name2186 (
		_w4082_,
		_w4084_,
		_w4085_,
		_w4086_,
		_w4087_
	);
	LUT3 #(
		.INIT('h0d)
	) name2187 (
		_w3163_,
		_w3164_,
		_w3165_,
		_w4088_
	);
	LUT4 #(
		.INIT('h00f2)
	) name2188 (
		_w3163_,
		_w3164_,
		_w3165_,
		_w3166_,
		_w4089_
	);
	LUT3 #(
		.INIT('h10)
	) name2189 (
		\s10_msel_arb3_state_reg[0]/NET0131 ,
		\s10_msel_arb3_state_reg[1]/NET0131 ,
		\s10_msel_arb3_state_reg[2]/NET0131 ,
		_w4090_
	);
	LUT4 #(
		.INIT('h2300)
	) name2190 (
		_w3153_,
		_w3154_,
		_w3161_,
		_w4090_,
		_w4091_
	);
	LUT3 #(
		.INIT('hd0)
	) name2191 (
		_w4083_,
		_w4089_,
		_w4091_,
		_w4092_
	);
	LUT3 #(
		.INIT('h0e)
	) name2192 (
		_w3154_,
		_w4087_,
		_w4092_,
		_w4093_
	);
	LUT2 #(
		.INIT('h1)
	) name2193 (
		\s10_msel_arb3_state_reg[1]/NET0131 ,
		\s10_msel_arb3_state_reg[2]/NET0131 ,
		_w4094_
	);
	LUT4 #(
		.INIT('h0080)
	) name2194 (
		\m0_s10_cyc_o_reg/NET0131 ,
		\rf_conf10_reg[0]/NET0131 ,
		\rf_conf10_reg[1]/NET0131 ,
		\s10_msel_arb3_state_reg[0]/NET0131 ,
		_w4095_
	);
	LUT2 #(
		.INIT('h2)
	) name2195 (
		_w4094_,
		_w4095_,
		_w4096_
	);
	LUT2 #(
		.INIT('h1)
	) name2196 (
		_w3154_,
		_w3164_,
		_w4097_
	);
	LUT4 #(
		.INIT('h4fcf)
	) name2197 (
		_w4084_,
		_w4088_,
		_w4096_,
		_w4097_,
		_w4098_
	);
	LUT3 #(
		.INIT('h20)
	) name2198 (
		_w3163_,
		_w3171_,
		_w4081_,
		_w4099_
	);
	LUT3 #(
		.INIT('h20)
	) name2199 (
		\s10_msel_arb3_state_reg[0]/NET0131 ,
		\s10_msel_arb3_state_reg[1]/NET0131 ,
		\s10_msel_arb3_state_reg[2]/NET0131 ,
		_w4100_
	);
	LUT2 #(
		.INIT('h8)
	) name2200 (
		_w3153_,
		_w4100_,
		_w4101_
	);
	LUT2 #(
		.INIT('h1)
	) name2201 (
		_w4099_,
		_w4101_,
		_w4102_
	);
	LUT2 #(
		.INIT('h8)
	) name2202 (
		_w4098_,
		_w4102_,
		_w4103_
	);
	LUT3 #(
		.INIT('h02)
	) name2203 (
		\s10_msel_arb3_state_reg[0]/NET0131 ,
		\s10_msel_arb3_state_reg[1]/NET0131 ,
		\s10_msel_arb3_state_reg[2]/NET0131 ,
		_w4104_
	);
	LUT4 #(
		.INIT('h0100)
	) name2204 (
		_w3154_,
		_w3164_,
		_w3166_,
		_w4104_,
		_w4105_
	);
	LUT2 #(
		.INIT('h4)
	) name2205 (
		_w3153_,
		_w4100_,
		_w4106_
	);
	LUT2 #(
		.INIT('h1)
	) name2206 (
		_w4105_,
		_w4106_,
		_w4107_
	);
	LUT2 #(
		.INIT('h4)
	) name2207 (
		_w3160_,
		_w3166_,
		_w4108_
	);
	LUT4 #(
		.INIT('h0051)
	) name2208 (
		_w3160_,
		_w3163_,
		_w3164_,
		_w3165_,
		_w4109_
	);
	LUT4 #(
		.INIT('h7f00)
	) name2209 (
		\m0_s10_cyc_o_reg/NET0131 ,
		\rf_conf10_reg[0]/NET0131 ,
		\rf_conf10_reg[1]/NET0131 ,
		\s10_msel_arb3_state_reg[0]/NET0131 ,
		_w4110_
	);
	LUT3 #(
		.INIT('h10)
	) name2210 (
		_w3154_,
		_w3164_,
		_w4110_,
		_w4111_
	);
	LUT4 #(
		.INIT('h0054)
	) name2211 (
		_w4105_,
		_w4108_,
		_w4109_,
		_w4111_,
		_w4112_
	);
	LUT3 #(
		.INIT('h01)
	) name2212 (
		_w3161_,
		_w4107_,
		_w4112_,
		_w4113_
	);
	LUT4 #(
		.INIT('h007f)
	) name2213 (
		\m5_s10_cyc_o_reg/NET0131 ,
		\rf_conf10_reg[10]/NET0131 ,
		\rf_conf10_reg[11]/NET0131 ,
		\s10_msel_arb3_state_reg[0]/NET0131 ,
		_w4114_
	);
	LUT4 #(
		.INIT('h0001)
	) name2214 (
		_w3154_,
		_w3164_,
		_w3166_,
		_w4114_,
		_w4115_
	);
	LUT3 #(
		.INIT('h0e)
	) name2215 (
		_w4108_,
		_w4109_,
		_w4115_,
		_w4116_
	);
	LUT4 #(
		.INIT('h0080)
	) name2216 (
		\m6_s10_cyc_o_reg/NET0131 ,
		\rf_conf10_reg[12]/NET0131 ,
		\rf_conf10_reg[13]/NET0131 ,
		\s10_msel_arb3_state_reg[0]/NET0131 ,
		_w4117_
	);
	LUT3 #(
		.INIT('h10)
	) name2217 (
		_w3153_,
		_w3160_,
		_w3161_,
		_w4118_
	);
	LUT4 #(
		.INIT('h020a)
	) name2218 (
		_w3179_,
		_w4088_,
		_w4117_,
		_w4118_,
		_w4119_
	);
	LUT2 #(
		.INIT('h4)
	) name2219 (
		_w4116_,
		_w4119_,
		_w4120_
	);
	LUT4 #(
		.INIT('hfff7)
	) name2220 (
		_w4093_,
		_w4103_,
		_w4113_,
		_w4120_,
		_w4121_
	);
	LUT2 #(
		.INIT('h4)
	) name2221 (
		_w2270_,
		_w2278_,
		_w4122_
	);
	LUT3 #(
		.INIT('h04)
	) name2222 (
		_w2266_,
		_w2268_,
		_w2269_,
		_w4123_
	);
	LUT4 #(
		.INIT('hfd00)
	) name2223 (
		\m4_s11_cyc_o_reg/NET0131 ,
		\rf_conf11_reg[8]/NET0131 ,
		\rf_conf11_reg[9]/NET0131 ,
		\s11_msel_arb0_state_reg[0]/NET0131 ,
		_w4124_
	);
	LUT3 #(
		.INIT('h10)
	) name2224 (
		_w2269_,
		_w2271_,
		_w4124_,
		_w4125_
	);
	LUT3 #(
		.INIT('hf2)
	) name2225 (
		_w2265_,
		_w2266_,
		_w2273_,
		_w4126_
	);
	LUT4 #(
		.INIT('h000d)
	) name2226 (
		_w2265_,
		_w2266_,
		_w2270_,
		_w2273_,
		_w4127_
	);
	LUT4 #(
		.INIT('h5455)
	) name2227 (
		_w4122_,
		_w4123_,
		_w4125_,
		_w4127_,
		_w4128_
	);
	LUT2 #(
		.INIT('h8)
	) name2228 (
		_w2292_,
		_w4128_,
		_w4129_
	);
	LUT2 #(
		.INIT('h8)
	) name2229 (
		\s11_msel_arb0_state_reg[1]/NET0131 ,
		\s11_msel_arb0_state_reg[2]/NET0131 ,
		_w4130_
	);
	LUT2 #(
		.INIT('h2)
	) name2230 (
		_w2273_,
		_w2278_,
		_w4131_
	);
	LUT3 #(
		.INIT('h51)
	) name2231 (
		_w2270_,
		_w2273_,
		_w2278_,
		_w4132_
	);
	LUT4 #(
		.INIT('h2232)
	) name2232 (
		_w2270_,
		_w2271_,
		_w2273_,
		_w2278_,
		_w4133_
	);
	LUT2 #(
		.INIT('h1)
	) name2233 (
		_w2266_,
		_w2278_,
		_w4134_
	);
	LUT4 #(
		.INIT('h00fd)
	) name2234 (
		\m5_s11_cyc_o_reg/NET0131 ,
		\rf_conf11_reg[10]/NET0131 ,
		\rf_conf11_reg[11]/NET0131 ,
		\s11_msel_arb0_state_reg[0]/NET0131 ,
		_w4135_
	);
	LUT3 #(
		.INIT('h01)
	) name2235 (
		_w2266_,
		_w2278_,
		_w4135_,
		_w4136_
	);
	LUT2 #(
		.INIT('h4)
	) name2236 (
		_w2265_,
		_w2269_,
		_w4137_
	);
	LUT3 #(
		.INIT('h0b)
	) name2237 (
		_w2265_,
		_w2269_,
		_w2271_,
		_w4138_
	);
	LUT4 #(
		.INIT('h0111)
	) name2238 (
		_w2268_,
		_w4133_,
		_w4136_,
		_w4138_,
		_w4139_
	);
	LUT4 #(
		.INIT('h1101)
	) name2239 (
		_w2265_,
		_w2268_,
		_w2270_,
		_w2271_,
		_w4140_
	);
	LUT4 #(
		.INIT('hfd00)
	) name2240 (
		\m2_s11_cyc_o_reg/NET0131 ,
		\rf_conf11_reg[4]/NET0131 ,
		\rf_conf11_reg[5]/NET0131 ,
		\s11_msel_arb0_state_reg[0]/NET0131 ,
		_w4141_
	);
	LUT4 #(
		.INIT('h0e0f)
	) name2241 (
		_w2269_,
		_w2271_,
		_w2273_,
		_w4141_,
		_w4142_
	);
	LUT2 #(
		.INIT('h2)
	) name2242 (
		\s11_msel_arb0_state_reg[1]/NET0131 ,
		\s11_msel_arb0_state_reg[2]/NET0131 ,
		_w4143_
	);
	LUT3 #(
		.INIT('hd0)
	) name2243 (
		_w2266_,
		_w2273_,
		_w4143_,
		_w4144_
	);
	LUT4 #(
		.INIT('h1f00)
	) name2244 (
		_w4137_,
		_w4140_,
		_w4142_,
		_w4144_,
		_w4145_
	);
	LUT3 #(
		.INIT('h0d)
	) name2245 (
		_w4130_,
		_w4139_,
		_w4145_,
		_w4146_
	);
	LUT3 #(
		.INIT('h8a)
	) name2246 (
		\s11_msel_arb0_state_reg[0]/NET0131 ,
		_w4129_,
		_w4146_,
		_w4147_
	);
	LUT3 #(
		.INIT('h02)
	) name2247 (
		\s11_msel_arb0_state_reg[0]/NET0131 ,
		_w2269_,
		_w2271_,
		_w4148_
	);
	LUT4 #(
		.INIT('h55fd)
	) name2248 (
		_w4134_,
		_w4137_,
		_w4140_,
		_w4148_,
		_w4149_
	);
	LUT3 #(
		.INIT('h8c)
	) name2249 (
		_w4131_,
		_w4143_,
		_w4149_,
		_w4150_
	);
	LUT3 #(
		.INIT('h20)
	) name2250 (
		_w2268_,
		_w2269_,
		_w4130_,
		_w4151_
	);
	LUT3 #(
		.INIT('h10)
	) name2251 (
		_w2269_,
		_w2271_,
		_w4130_,
		_w4152_
	);
	LUT4 #(
		.INIT('h020f)
	) name2252 (
		_w4132_,
		_w4136_,
		_w4151_,
		_w4152_,
		_w4153_
	);
	LUT3 #(
		.INIT('h20)
	) name2253 (
		_w2270_,
		_w2271_,
		_w2292_,
		_w4154_
	);
	LUT2 #(
		.INIT('h1)
	) name2254 (
		_w2266_,
		_w2269_,
		_w4155_
	);
	LUT4 #(
		.INIT('h00fd)
	) name2255 (
		\m7_s11_cyc_o_reg/NET0131 ,
		\rf_conf11_reg[14]/NET0131 ,
		\rf_conf11_reg[15]/NET0131 ,
		\s11_msel_arb0_state_reg[0]/NET0131 ,
		_w4156_
	);
	LUT3 #(
		.INIT('h01)
	) name2256 (
		_w2266_,
		_w2269_,
		_w4156_,
		_w4157_
	);
	LUT3 #(
		.INIT('h10)
	) name2257 (
		_w2271_,
		_w2278_,
		_w2292_,
		_w4158_
	);
	LUT4 #(
		.INIT('h0133)
	) name2258 (
		_w4126_,
		_w4154_,
		_w4157_,
		_w4158_,
		_w4159_
	);
	LUT2 #(
		.INIT('h8)
	) name2259 (
		_w4153_,
		_w4159_,
		_w4160_
	);
	LUT3 #(
		.INIT('h02)
	) name2260 (
		\s11_msel_arb0_state_reg[0]/NET0131 ,
		_w2271_,
		_w2278_,
		_w4161_
	);
	LUT3 #(
		.INIT('h80)
	) name2261 (
		_w2295_,
		_w4155_,
		_w4161_,
		_w4162_
	);
	LUT3 #(
		.INIT('h04)
	) name2262 (
		_w2271_,
		_w2273_,
		_w2278_,
		_w4163_
	);
	LUT4 #(
		.INIT('h0002)
	) name2263 (
		\m4_s11_cyc_o_reg/NET0131 ,
		\rf_conf11_reg[8]/NET0131 ,
		\rf_conf11_reg[9]/NET0131 ,
		\s11_msel_arb0_state_reg[0]/NET0131 ,
		_w4164_
	);
	LUT4 #(
		.INIT('h00b0)
	) name2264 (
		_w2265_,
		_w2269_,
		_w2295_,
		_w4164_,
		_w4165_
	);
	LUT3 #(
		.INIT('hd0)
	) name2265 (
		_w4140_,
		_w4163_,
		_w4165_,
		_w4166_
	);
	LUT2 #(
		.INIT('h1)
	) name2266 (
		_w4162_,
		_w4166_,
		_w4167_
	);
	LUT4 #(
		.INIT('hba00)
	) name2267 (
		\s11_msel_arb0_state_reg[0]/NET0131 ,
		_w4150_,
		_w4160_,
		_w4167_,
		_w4168_
	);
	LUT2 #(
		.INIT('hb)
	) name2268 (
		_w4147_,
		_w4168_,
		_w4169_
	);
	LUT4 #(
		.INIT('h0008)
	) name2269 (
		\m4_s11_cyc_o_reg/NET0131 ,
		\rf_conf11_reg[8]/NET0131 ,
		\rf_conf11_reg[9]/NET0131 ,
		\s11_msel_arb1_state_reg[0]/NET0131 ,
		_w4170_
	);
	LUT2 #(
		.INIT('h2)
	) name2270 (
		_w3609_,
		_w4170_,
		_w4171_
	);
	LUT2 #(
		.INIT('h4)
	) name2271 (
		_w3587_,
		_w3594_,
		_w4172_
	);
	LUT4 #(
		.INIT('h0031)
	) name2272 (
		_w3584_,
		_w3587_,
		_w3600_,
		_w3601_,
		_w4173_
	);
	LUT2 #(
		.INIT('h1)
	) name2273 (
		_w4172_,
		_w4173_,
		_w4174_
	);
	LUT3 #(
		.INIT('h01)
	) name2274 (
		_w3588_,
		_w4172_,
		_w4173_,
		_w4175_
	);
	LUT2 #(
		.INIT('h1)
	) name2275 (
		_w3588_,
		_w3594_,
		_w4176_
	);
	LUT3 #(
		.INIT('h02)
	) name2276 (
		\s11_msel_arb1_state_reg[0]/NET0131 ,
		_w3590_,
		_w3600_,
		_w4177_
	);
	LUT2 #(
		.INIT('h8)
	) name2277 (
		_w4176_,
		_w4177_,
		_w4178_
	);
	LUT3 #(
		.INIT('h15)
	) name2278 (
		_w3591_,
		_w4176_,
		_w4177_,
		_w4179_
	);
	LUT3 #(
		.INIT('h8a)
	) name2279 (
		_w4171_,
		_w4175_,
		_w4179_,
		_w4180_
	);
	LUT3 #(
		.INIT('h04)
	) name2280 (
		\s11_msel_arb1_state_reg[0]/NET0131 ,
		\s11_msel_arb1_state_reg[1]/NET0131 ,
		\s11_msel_arb1_state_reg[2]/NET0131 ,
		_w4181_
	);
	LUT3 #(
		.INIT('h20)
	) name2281 (
		_w3584_,
		_w3600_,
		_w4181_,
		_w4182_
	);
	LUT3 #(
		.INIT('h0d)
	) name2282 (
		_w3587_,
		_w3588_,
		_w3591_,
		_w4183_
	);
	LUT4 #(
		.INIT('h00f7)
	) name2283 (
		\m1_s11_cyc_o_reg/NET0131 ,
		\rf_conf11_reg[2]/NET0131 ,
		\rf_conf11_reg[3]/NET0131 ,
		\s11_msel_arb1_state_reg[0]/NET0131 ,
		_w4184_
	);
	LUT3 #(
		.INIT('h01)
	) name2284 (
		_w3588_,
		_w3594_,
		_w4184_,
		_w4185_
	);
	LUT3 #(
		.INIT('h10)
	) name2285 (
		_w3590_,
		_w3600_,
		_w4181_,
		_w4186_
	);
	LUT4 #(
		.INIT('h0455)
	) name2286 (
		_w4182_,
		_w4183_,
		_w4185_,
		_w4186_,
		_w4187_
	);
	LUT4 #(
		.INIT('h0004)
	) name2287 (
		_w3590_,
		_w3591_,
		_w3594_,
		_w3600_,
		_w4188_
	);
	LUT3 #(
		.INIT('h07)
	) name2288 (
		_w4176_,
		_w4177_,
		_w4188_,
		_w4189_
	);
	LUT2 #(
		.INIT('h2)
	) name2289 (
		_w3595_,
		_w3612_,
		_w4190_
	);
	LUT4 #(
		.INIT('h40cc)
	) name2290 (
		_w4174_,
		_w4187_,
		_w4189_,
		_w4190_,
		_w4191_
	);
	LUT4 #(
		.INIT('h0f02)
	) name2291 (
		_w3587_,
		_w3588_,
		_w3590_,
		_w3591_,
		_w4192_
	);
	LUT3 #(
		.INIT('h51)
	) name2292 (
		_w3590_,
		_w3600_,
		_w3601_,
		_w4193_
	);
	LUT4 #(
		.INIT('h0105)
	) name2293 (
		_w3584_,
		_w4185_,
		_w4192_,
		_w4193_,
		_w4194_
	);
	LUT2 #(
		.INIT('h2)
	) name2294 (
		_w3586_,
		_w4194_,
		_w4195_
	);
	LUT4 #(
		.INIT('h3302)
	) name2295 (
		_w3584_,
		_w3598_,
		_w3600_,
		_w3601_,
		_w4196_
	);
	LUT3 #(
		.INIT('h01)
	) name2296 (
		_w3590_,
		_w3598_,
		_w3600_,
		_w4197_
	);
	LUT3 #(
		.INIT('h23)
	) name2297 (
		_w4183_,
		_w4196_,
		_w4197_,
		_w4198_
	);
	LUT2 #(
		.INIT('h1)
	) name2298 (
		\s11_msel_arb1_state_reg[1]/NET0131 ,
		\s11_msel_arb1_state_reg[2]/NET0131 ,
		_w4199_
	);
	LUT3 #(
		.INIT('hb0)
	) name2299 (
		_w4178_,
		_w4198_,
		_w4199_,
		_w4200_
	);
	LUT4 #(
		.INIT('hfffb)
	) name2300 (
		_w4180_,
		_w4191_,
		_w4195_,
		_w4200_,
		_w4201_
	);
	LUT2 #(
		.INIT('h4)
	) name2301 (
		\s11_msel_arb2_state_reg[1]/NET0131 ,
		\s11_msel_arb2_state_reg[2]/NET0131 ,
		_w4202_
	);
	LUT3 #(
		.INIT('h20)
	) name2302 (
		_w3183_,
		_w3184_,
		_w4202_,
		_w4203_
	);
	LUT2 #(
		.INIT('h4)
	) name2303 (
		_w3186_,
		_w3198_,
		_w4204_
	);
	LUT2 #(
		.INIT('h2)
	) name2304 (
		_w3189_,
		_w3191_,
		_w4205_
	);
	LUT4 #(
		.INIT('h0051)
	) name2305 (
		_w3186_,
		_w3189_,
		_w3191_,
		_w3194_,
		_w4206_
	);
	LUT3 #(
		.INIT('h10)
	) name2306 (
		_w3184_,
		_w3185_,
		_w4202_,
		_w4207_
	);
	LUT4 #(
		.INIT('h5455)
	) name2307 (
		_w4203_,
		_w4204_,
		_w4206_,
		_w4207_,
		_w4208_
	);
	LUT2 #(
		.INIT('h1)
	) name2308 (
		\s11_msel_arb2_state_reg[0]/NET0131 ,
		_w4208_,
		_w4209_
	);
	LUT2 #(
		.INIT('h1)
	) name2309 (
		_w3184_,
		_w3191_,
		_w4210_
	);
	LUT3 #(
		.INIT('hf2)
	) name2310 (
		_w3184_,
		_w3189_,
		_w3191_,
		_w4211_
	);
	LUT3 #(
		.INIT('h45)
	) name2311 (
		_w3183_,
		_w3185_,
		_w3186_,
		_w4212_
	);
	LUT3 #(
		.INIT('h04)
	) name2312 (
		_w3185_,
		_w3194_,
		_w3198_,
		_w4213_
	);
	LUT3 #(
		.INIT('h02)
	) name2313 (
		\s11_msel_arb2_state_reg[0]/NET0131 ,
		_w3185_,
		_w3198_,
		_w4214_
	);
	LUT4 #(
		.INIT('h0004)
	) name2314 (
		_w4205_,
		_w4212_,
		_w4213_,
		_w4214_,
		_w4215_
	);
	LUT3 #(
		.INIT('h04)
	) name2315 (
		\s11_msel_arb2_state_reg[0]/NET0131 ,
		\s11_msel_arb2_state_reg[1]/NET0131 ,
		\s11_msel_arb2_state_reg[2]/NET0131 ,
		_w4216_
	);
	LUT3 #(
		.INIT('h10)
	) name2316 (
		_w4211_,
		_w4215_,
		_w4216_,
		_w4217_
	);
	LUT2 #(
		.INIT('h1)
	) name2317 (
		_w4209_,
		_w4217_,
		_w4218_
	);
	LUT4 #(
		.INIT('hdf00)
	) name2318 (
		\m6_s11_cyc_o_reg/NET0131 ,
		\rf_conf11_reg[12]/NET0131 ,
		\rf_conf11_reg[13]/NET0131 ,
		\s11_msel_arb2_state_reg[0]/NET0131 ,
		_w4219_
	);
	LUT2 #(
		.INIT('h1)
	) name2319 (
		_w3183_,
		_w4219_,
		_w4220_
	);
	LUT3 #(
		.INIT('h01)
	) name2320 (
		_w3184_,
		_w3191_,
		_w3198_,
		_w4221_
	);
	LUT4 #(
		.INIT('he0ee)
	) name2321 (
		_w4204_,
		_w4206_,
		_w4220_,
		_w4221_,
		_w4222_
	);
	LUT4 #(
		.INIT('h0020)
	) name2322 (
		\m6_s11_cyc_o_reg/NET0131 ,
		\rf_conf11_reg[12]/NET0131 ,
		\rf_conf11_reg[13]/NET0131 ,
		\s11_msel_arb2_state_reg[0]/NET0131 ,
		_w4223_
	);
	LUT2 #(
		.INIT('h8)
	) name2323 (
		\s11_msel_arb2_state_reg[1]/NET0131 ,
		\s11_msel_arb2_state_reg[2]/NET0131 ,
		_w4224_
	);
	LUT2 #(
		.INIT('h4)
	) name2324 (
		_w4223_,
		_w4224_,
		_w4225_
	);
	LUT2 #(
		.INIT('h4)
	) name2325 (
		_w4222_,
		_w4225_,
		_w4226_
	);
	LUT3 #(
		.INIT('h51)
	) name2326 (
		_w3184_,
		_w4212_,
		_w4213_,
		_w4227_
	);
	LUT2 #(
		.INIT('h8)
	) name2327 (
		_w4210_,
		_w4214_,
		_w4228_
	);
	LUT3 #(
		.INIT('h15)
	) name2328 (
		_w3189_,
		_w4210_,
		_w4214_,
		_w4229_
	);
	LUT3 #(
		.INIT('h08)
	) name2329 (
		\s11_msel_arb2_state_reg[0]/NET0131 ,
		\s11_msel_arb2_state_reg[1]/NET0131 ,
		\s11_msel_arb2_state_reg[2]/NET0131 ,
		_w4230_
	);
	LUT3 #(
		.INIT('hb0)
	) name2330 (
		_w4227_,
		_w4229_,
		_w4230_,
		_w4231_
	);
	LUT2 #(
		.INIT('h2)
	) name2331 (
		\s11_msel_arb2_state_reg[0]/NET0131 ,
		\s11_msel_arb2_state_reg[1]/NET0131 ,
		_w4232_
	);
	LUT3 #(
		.INIT('h20)
	) name2332 (
		\s11_msel_arb2_state_reg[0]/NET0131 ,
		\s11_msel_arb2_state_reg[1]/NET0131 ,
		\s11_msel_arb2_state_reg[2]/NET0131 ,
		_w4233_
	);
	LUT3 #(
		.INIT('h01)
	) name2333 (
		_w3185_,
		_w4204_,
		_w4206_,
		_w4234_
	);
	LUT3 #(
		.INIT('h15)
	) name2334 (
		_w3183_,
		_w4210_,
		_w4214_,
		_w4235_
	);
	LUT3 #(
		.INIT('h8a)
	) name2335 (
		_w4233_,
		_w4234_,
		_w4235_,
		_w4236_
	);
	LUT4 #(
		.INIT('h0020)
	) name2336 (
		\m0_s11_cyc_o_reg/NET0131 ,
		\rf_conf11_reg[0]/NET0131 ,
		\rf_conf11_reg[1]/NET0131 ,
		\s11_msel_arb2_state_reg[0]/NET0131 ,
		_w4237_
	);
	LUT4 #(
		.INIT('h00f2)
	) name2337 (
		_w3189_,
		_w3191_,
		_w3194_,
		_w4237_,
		_w4238_
	);
	LUT3 #(
		.INIT('h01)
	) name2338 (
		_w3184_,
		_w3191_,
		_w4237_,
		_w4239_
	);
	LUT3 #(
		.INIT('h23)
	) name2339 (
		_w4212_,
		_w4238_,
		_w4239_,
		_w4240_
	);
	LUT2 #(
		.INIT('h1)
	) name2340 (
		\s11_msel_arb2_state_reg[1]/NET0131 ,
		\s11_msel_arb2_state_reg[2]/NET0131 ,
		_w4241_
	);
	LUT3 #(
		.INIT('hb0)
	) name2341 (
		_w4228_,
		_w4240_,
		_w4241_,
		_w4242_
	);
	LUT4 #(
		.INIT('h0001)
	) name2342 (
		_w4226_,
		_w4231_,
		_w4236_,
		_w4242_,
		_w4243_
	);
	LUT2 #(
		.INIT('h7)
	) name2343 (
		_w4218_,
		_w4243_,
		_w4244_
	);
	LUT3 #(
		.INIT('hdc)
	) name2344 (
		_w3208_,
		_w3209_,
		_w3219_,
		_w4245_
	);
	LUT2 #(
		.INIT('h4)
	) name2345 (
		_w3211_,
		_w3213_,
		_w4246_
	);
	LUT4 #(
		.INIT('h000d)
	) name2346 (
		_w3206_,
		_w3207_,
		_w3211_,
		_w3212_,
		_w4247_
	);
	LUT4 #(
		.INIT('h7f00)
	) name2347 (
		\m6_s11_cyc_o_reg/NET0131 ,
		\rf_conf11_reg[12]/NET0131 ,
		\rf_conf11_reg[13]/NET0131 ,
		\s11_msel_arb3_state_reg[0]/NET0131 ,
		_w4248_
	);
	LUT4 #(
		.INIT('ha2f3)
	) name2348 (
		_w3207_,
		_w3208_,
		_w3209_,
		_w4248_,
		_w4249_
	);
	LUT4 #(
		.INIT('h0155)
	) name2349 (
		_w4245_,
		_w4246_,
		_w4247_,
		_w4249_,
		_w4250_
	);
	LUT2 #(
		.INIT('h8)
	) name2350 (
		_w3231_,
		_w4250_,
		_w4251_
	);
	LUT2 #(
		.INIT('h1)
	) name2351 (
		\s11_msel_arb3_state_reg[1]/NET0131 ,
		\s11_msel_arb3_state_reg[2]/NET0131 ,
		_w4252_
	);
	LUT3 #(
		.INIT('h20)
	) name2352 (
		_w3206_,
		_w3207_,
		_w4252_,
		_w4253_
	);
	LUT2 #(
		.INIT('h4)
	) name2353 (
		_w3208_,
		_w3219_,
		_w4254_
	);
	LUT4 #(
		.INIT('h1101)
	) name2354 (
		_w3208_,
		_w3211_,
		_w3212_,
		_w3213_,
		_w4255_
	);
	LUT3 #(
		.INIT('h10)
	) name2355 (
		_w3207_,
		_w3209_,
		_w4252_,
		_w4256_
	);
	LUT4 #(
		.INIT('h5455)
	) name2356 (
		_w4253_,
		_w4254_,
		_w4255_,
		_w4256_,
		_w4257_
	);
	LUT3 #(
		.INIT('h08)
	) name2357 (
		_w3205_,
		_w3211_,
		_w3219_,
		_w4258_
	);
	LUT3 #(
		.INIT('h0d)
	) name2358 (
		_w3206_,
		_w3207_,
		_w3212_,
		_w4259_
	);
	LUT3 #(
		.INIT('h04)
	) name2359 (
		_w3207_,
		_w3208_,
		_w3209_,
		_w4260_
	);
	LUT3 #(
		.INIT('h02)
	) name2360 (
		_w3205_,
		_w3213_,
		_w3219_,
		_w4261_
	);
	LUT4 #(
		.INIT('h0455)
	) name2361 (
		_w4258_,
		_w4259_,
		_w4260_,
		_w4261_,
		_w4262_
	);
	LUT3 #(
		.INIT('h40)
	) name2362 (
		\s11_msel_arb3_state_reg[0]/NET0131 ,
		_w4257_,
		_w4262_,
		_w4263_
	);
	LUT3 #(
		.INIT('h51)
	) name2363 (
		_w3213_,
		_w4259_,
		_w4260_,
		_w4264_
	);
	LUT4 #(
		.INIT('h0001)
	) name2364 (
		_w3207_,
		_w3209_,
		_w3213_,
		_w3219_,
		_w4265_
	);
	LUT2 #(
		.INIT('h1)
	) name2365 (
		_w3211_,
		_w4265_,
		_w4266_
	);
	LUT3 #(
		.INIT('h2a)
	) name2366 (
		\s11_msel_arb3_state_reg[0]/NET0131 ,
		_w3208_,
		_w3231_,
		_w4267_
	);
	LUT4 #(
		.INIT('h7500)
	) name2367 (
		_w3205_,
		_w4264_,
		_w4266_,
		_w4267_,
		_w4268_
	);
	LUT3 #(
		.INIT('h0b)
	) name2368 (
		_w4251_,
		_w4263_,
		_w4268_,
		_w4269_
	);
	LUT2 #(
		.INIT('h4)
	) name2369 (
		_w3206_,
		_w3209_,
		_w4270_
	);
	LUT4 #(
		.INIT('h5455)
	) name2370 (
		_w3206_,
		_w3207_,
		_w3219_,
		_w4248_,
		_w4271_
	);
	LUT4 #(
		.INIT('h010f)
	) name2371 (
		_w4254_,
		_w4255_,
		_w4270_,
		_w4271_,
		_w4272_
	);
	LUT3 #(
		.INIT('h02)
	) name2372 (
		\s11_msel_arb3_state_reg[0]/NET0131 ,
		\s11_msel_arb3_state_reg[1]/NET0131 ,
		\s11_msel_arb3_state_reg[2]/NET0131 ,
		_w4273_
	);
	LUT2 #(
		.INIT('h8)
	) name2373 (
		_w4272_,
		_w4273_,
		_w4274_
	);
	LUT2 #(
		.INIT('h1)
	) name2374 (
		_w3211_,
		_w4248_,
		_w4275_
	);
	LUT3 #(
		.INIT('h01)
	) name2375 (
		_w3207_,
		_w3209_,
		_w3219_,
		_w4276_
	);
	LUT4 #(
		.INIT('h2022)
	) name2376 (
		_w4259_,
		_w4260_,
		_w4275_,
		_w4276_,
		_w4277_
	);
	LUT4 #(
		.INIT('h0080)
	) name2377 (
		\m6_s11_cyc_o_reg/NET0131 ,
		\rf_conf11_reg[12]/NET0131 ,
		\rf_conf11_reg[13]/NET0131 ,
		\s11_msel_arb3_state_reg[0]/NET0131 ,
		_w4278_
	);
	LUT2 #(
		.INIT('h2)
	) name2378 (
		_w3217_,
		_w4278_,
		_w4279_
	);
	LUT3 #(
		.INIT('h10)
	) name2379 (
		_w3207_,
		_w3209_,
		_w4248_,
		_w4280_
	);
	LUT3 #(
		.INIT('h08)
	) name2380 (
		\s11_msel_arb3_state_reg[0]/NET0131 ,
		\s11_msel_arb3_state_reg[1]/NET0131 ,
		\s11_msel_arb3_state_reg[2]/NET0131 ,
		_w4281_
	);
	LUT3 #(
		.INIT('h10)
	) name2381 (
		_w3208_,
		_w3219_,
		_w4281_,
		_w4282_
	);
	LUT4 #(
		.INIT('hf100)
	) name2382 (
		_w4246_,
		_w4247_,
		_w4280_,
		_w4282_,
		_w4283_
	);
	LUT3 #(
		.INIT('h0b)
	) name2383 (
		_w4277_,
		_w4279_,
		_w4283_,
		_w4284_
	);
	LUT2 #(
		.INIT('h4)
	) name2384 (
		_w4274_,
		_w4284_,
		_w4285_
	);
	LUT2 #(
		.INIT('hb)
	) name2385 (
		_w4269_,
		_w4285_,
		_w4286_
	);
	LUT2 #(
		.INIT('h4)
	) name2386 (
		_w2307_,
		_w2315_,
		_w4287_
	);
	LUT3 #(
		.INIT('h04)
	) name2387 (
		_w2303_,
		_w2305_,
		_w2306_,
		_w4288_
	);
	LUT4 #(
		.INIT('hfd00)
	) name2388 (
		\m4_s12_cyc_o_reg/NET0131 ,
		\rf_conf12_reg[8]/NET0131 ,
		\rf_conf12_reg[9]/NET0131 ,
		\s12_msel_arb0_state_reg[0]/NET0131 ,
		_w4289_
	);
	LUT3 #(
		.INIT('h10)
	) name2389 (
		_w2306_,
		_w2308_,
		_w4289_,
		_w4290_
	);
	LUT3 #(
		.INIT('hf2)
	) name2390 (
		_w2302_,
		_w2303_,
		_w2310_,
		_w4291_
	);
	LUT4 #(
		.INIT('h000d)
	) name2391 (
		_w2302_,
		_w2303_,
		_w2307_,
		_w2310_,
		_w4292_
	);
	LUT4 #(
		.INIT('h5455)
	) name2392 (
		_w4287_,
		_w4288_,
		_w4290_,
		_w4292_,
		_w4293_
	);
	LUT2 #(
		.INIT('h8)
	) name2393 (
		_w2329_,
		_w4293_,
		_w4294_
	);
	LUT2 #(
		.INIT('h8)
	) name2394 (
		\s12_msel_arb0_state_reg[1]/NET0131 ,
		\s12_msel_arb0_state_reg[2]/NET0131 ,
		_w4295_
	);
	LUT2 #(
		.INIT('h2)
	) name2395 (
		_w2310_,
		_w2315_,
		_w4296_
	);
	LUT3 #(
		.INIT('h51)
	) name2396 (
		_w2307_,
		_w2310_,
		_w2315_,
		_w4297_
	);
	LUT4 #(
		.INIT('h2232)
	) name2397 (
		_w2307_,
		_w2308_,
		_w2310_,
		_w2315_,
		_w4298_
	);
	LUT2 #(
		.INIT('h1)
	) name2398 (
		_w2303_,
		_w2315_,
		_w4299_
	);
	LUT4 #(
		.INIT('h00fd)
	) name2399 (
		\m5_s12_cyc_o_reg/NET0131 ,
		\rf_conf12_reg[10]/NET0131 ,
		\rf_conf12_reg[11]/NET0131 ,
		\s12_msel_arb0_state_reg[0]/NET0131 ,
		_w4300_
	);
	LUT3 #(
		.INIT('h01)
	) name2400 (
		_w2303_,
		_w2315_,
		_w4300_,
		_w4301_
	);
	LUT2 #(
		.INIT('h4)
	) name2401 (
		_w2302_,
		_w2306_,
		_w4302_
	);
	LUT3 #(
		.INIT('h0b)
	) name2402 (
		_w2302_,
		_w2306_,
		_w2308_,
		_w4303_
	);
	LUT4 #(
		.INIT('h0111)
	) name2403 (
		_w2305_,
		_w4298_,
		_w4301_,
		_w4303_,
		_w4304_
	);
	LUT4 #(
		.INIT('h1101)
	) name2404 (
		_w2302_,
		_w2305_,
		_w2307_,
		_w2308_,
		_w4305_
	);
	LUT4 #(
		.INIT('hfd00)
	) name2405 (
		\m2_s12_cyc_o_reg/NET0131 ,
		\rf_conf12_reg[4]/NET0131 ,
		\rf_conf12_reg[5]/NET0131 ,
		\s12_msel_arb0_state_reg[0]/NET0131 ,
		_w4306_
	);
	LUT4 #(
		.INIT('h0e0f)
	) name2406 (
		_w2306_,
		_w2308_,
		_w2310_,
		_w4306_,
		_w4307_
	);
	LUT2 #(
		.INIT('h2)
	) name2407 (
		\s12_msel_arb0_state_reg[1]/NET0131 ,
		\s12_msel_arb0_state_reg[2]/NET0131 ,
		_w4308_
	);
	LUT3 #(
		.INIT('hd0)
	) name2408 (
		_w2303_,
		_w2310_,
		_w4308_,
		_w4309_
	);
	LUT4 #(
		.INIT('h1f00)
	) name2409 (
		_w4302_,
		_w4305_,
		_w4307_,
		_w4309_,
		_w4310_
	);
	LUT3 #(
		.INIT('h0d)
	) name2410 (
		_w4295_,
		_w4304_,
		_w4310_,
		_w4311_
	);
	LUT3 #(
		.INIT('h8a)
	) name2411 (
		\s12_msel_arb0_state_reg[0]/NET0131 ,
		_w4294_,
		_w4311_,
		_w4312_
	);
	LUT3 #(
		.INIT('h02)
	) name2412 (
		\s12_msel_arb0_state_reg[0]/NET0131 ,
		_w2306_,
		_w2308_,
		_w4313_
	);
	LUT4 #(
		.INIT('h55fd)
	) name2413 (
		_w4299_,
		_w4302_,
		_w4305_,
		_w4313_,
		_w4314_
	);
	LUT3 #(
		.INIT('h8c)
	) name2414 (
		_w4296_,
		_w4308_,
		_w4314_,
		_w4315_
	);
	LUT3 #(
		.INIT('h20)
	) name2415 (
		_w2305_,
		_w2306_,
		_w4295_,
		_w4316_
	);
	LUT3 #(
		.INIT('h10)
	) name2416 (
		_w2306_,
		_w2308_,
		_w4295_,
		_w4317_
	);
	LUT4 #(
		.INIT('h020f)
	) name2417 (
		_w4297_,
		_w4301_,
		_w4316_,
		_w4317_,
		_w4318_
	);
	LUT3 #(
		.INIT('h20)
	) name2418 (
		_w2307_,
		_w2308_,
		_w2329_,
		_w4319_
	);
	LUT2 #(
		.INIT('h1)
	) name2419 (
		_w2303_,
		_w2306_,
		_w4320_
	);
	LUT4 #(
		.INIT('h00fd)
	) name2420 (
		\m7_s12_cyc_o_reg/NET0131 ,
		\rf_conf12_reg[14]/NET0131 ,
		\rf_conf12_reg[15]/NET0131 ,
		\s12_msel_arb0_state_reg[0]/NET0131 ,
		_w4321_
	);
	LUT3 #(
		.INIT('h01)
	) name2421 (
		_w2303_,
		_w2306_,
		_w4321_,
		_w4322_
	);
	LUT3 #(
		.INIT('h10)
	) name2422 (
		_w2308_,
		_w2315_,
		_w2329_,
		_w4323_
	);
	LUT4 #(
		.INIT('h0133)
	) name2423 (
		_w4291_,
		_w4319_,
		_w4322_,
		_w4323_,
		_w4324_
	);
	LUT2 #(
		.INIT('h8)
	) name2424 (
		_w4318_,
		_w4324_,
		_w4325_
	);
	LUT3 #(
		.INIT('h02)
	) name2425 (
		\s12_msel_arb0_state_reg[0]/NET0131 ,
		_w2308_,
		_w2315_,
		_w4326_
	);
	LUT3 #(
		.INIT('h80)
	) name2426 (
		_w2332_,
		_w4320_,
		_w4326_,
		_w4327_
	);
	LUT3 #(
		.INIT('h04)
	) name2427 (
		_w2308_,
		_w2310_,
		_w2315_,
		_w4328_
	);
	LUT4 #(
		.INIT('h0002)
	) name2428 (
		\m4_s12_cyc_o_reg/NET0131 ,
		\rf_conf12_reg[8]/NET0131 ,
		\rf_conf12_reg[9]/NET0131 ,
		\s12_msel_arb0_state_reg[0]/NET0131 ,
		_w4329_
	);
	LUT4 #(
		.INIT('h00b0)
	) name2429 (
		_w2302_,
		_w2306_,
		_w2332_,
		_w4329_,
		_w4330_
	);
	LUT3 #(
		.INIT('hd0)
	) name2430 (
		_w4305_,
		_w4328_,
		_w4330_,
		_w4331_
	);
	LUT2 #(
		.INIT('h1)
	) name2431 (
		_w4327_,
		_w4331_,
		_w4332_
	);
	LUT4 #(
		.INIT('hba00)
	) name2432 (
		\s12_msel_arb0_state_reg[0]/NET0131 ,
		_w4315_,
		_w4325_,
		_w4332_,
		_w4333_
	);
	LUT2 #(
		.INIT('hb)
	) name2433 (
		_w4312_,
		_w4333_,
		_w4334_
	);
	LUT3 #(
		.INIT('h0b)
	) name2434 (
		_w3625_,
		_w3626_,
		_w3631_,
		_w4335_
	);
	LUT4 #(
		.INIT('h0f04)
	) name2435 (
		_w3625_,
		_w3626_,
		_w3630_,
		_w3631_,
		_w4336_
	);
	LUT2 #(
		.INIT('h1)
	) name2436 (
		_w3623_,
		_w3625_,
		_w4337_
	);
	LUT4 #(
		.INIT('h0002)
	) name2437 (
		_w3622_,
		_w3623_,
		_w3625_,
		_w3630_,
		_w4338_
	);
	LUT4 #(
		.INIT('h3332)
	) name2438 (
		_w3619_,
		_w3620_,
		_w4336_,
		_w4338_,
		_w4339_
	);
	LUT4 #(
		.INIT('hf700)
	) name2439 (
		\m2_s12_cyc_o_reg/NET0131 ,
		\rf_conf12_reg[4]/NET0131 ,
		\rf_conf12_reg[5]/NET0131 ,
		\s12_msel_arb1_state_reg[0]/NET0131 ,
		_w4340_
	);
	LUT4 #(
		.INIT('h0100)
	) name2440 (
		_w3623_,
		_w3625_,
		_w3639_,
		_w4340_,
		_w4341_
	);
	LUT2 #(
		.INIT('h1)
	) name2441 (
		\s12_msel_arb1_state_reg[1]/NET0131 ,
		_w4341_,
		_w4342_
	);
	LUT3 #(
		.INIT('h10)
	) name2442 (
		\s12_msel_arb1_state_reg[2]/NET0131 ,
		_w4339_,
		_w4342_,
		_w4343_
	);
	LUT3 #(
		.INIT('h31)
	) name2443 (
		_w3619_,
		_w3622_,
		_w3639_,
		_w4344_
	);
	LUT4 #(
		.INIT('h3031)
	) name2444 (
		_w3619_,
		_w3622_,
		_w3639_,
		_w4340_,
		_w4345_
	);
	LUT4 #(
		.INIT('hf700)
	) name2445 (
		\m3_s12_cyc_o_reg/NET0131 ,
		\rf_conf12_reg[6]/NET0131 ,
		\rf_conf12_reg[7]/NET0131 ,
		\s12_msel_arb1_state_reg[0]/NET0131 ,
		_w4346_
	);
	LUT3 #(
		.INIT('hb0)
	) name2446 (
		_w3625_,
		_w3626_,
		_w4346_,
		_w4347_
	);
	LUT3 #(
		.INIT('hd0)
	) name2447 (
		_w4337_,
		_w4345_,
		_w4347_,
		_w4348_
	);
	LUT2 #(
		.INIT('h2)
	) name2448 (
		_w3623_,
		_w3626_,
		_w4349_
	);
	LUT4 #(
		.INIT('h0301)
	) name2449 (
		_w3619_,
		_w3622_,
		_w3626_,
		_w3639_,
		_w4350_
	);
	LUT2 #(
		.INIT('h1)
	) name2450 (
		_w3625_,
		_w3630_,
		_w4351_
	);
	LUT3 #(
		.INIT('h45)
	) name2451 (
		\s12_msel_arb1_state_reg[0]/NET0131 ,
		_w3630_,
		_w3631_,
		_w4352_
	);
	LUT4 #(
		.INIT('hef00)
	) name2452 (
		_w4349_,
		_w4350_,
		_w4351_,
		_w4352_,
		_w4353_
	);
	LUT2 #(
		.INIT('h2)
	) name2453 (
		\s12_msel_arb1_state_reg[1]/NET0131 ,
		\s12_msel_arb1_state_reg[2]/NET0131 ,
		_w4354_
	);
	LUT3 #(
		.INIT('he0)
	) name2454 (
		_w4348_,
		_w4353_,
		_w4354_,
		_w4355_
	);
	LUT4 #(
		.INIT('h0010)
	) name2455 (
		_w3623_,
		_w3630_,
		_w3631_,
		_w3639_,
		_w4356_
	);
	LUT2 #(
		.INIT('h1)
	) name2456 (
		\s12_msel_arb1_state_reg[1]/NET0131 ,
		_w3636_,
		_w4357_
	);
	LUT4 #(
		.INIT('hf100)
	) name2457 (
		_w4349_,
		_w4350_,
		_w4356_,
		_w4357_,
		_w4358_
	);
	LUT2 #(
		.INIT('h1)
	) name2458 (
		_w3630_,
		_w3639_,
		_w4359_
	);
	LUT4 #(
		.INIT('h2a0a)
	) name2459 (
		_w3635_,
		_w4335_,
		_w4344_,
		_w4359_,
		_w4360_
	);
	LUT2 #(
		.INIT('h2)
	) name2460 (
		\s12_msel_arb1_state_reg[2]/NET0131 ,
		_w4341_,
		_w4361_
	);
	LUT3 #(
		.INIT('h10)
	) name2461 (
		_w4358_,
		_w4360_,
		_w4361_,
		_w4362_
	);
	LUT3 #(
		.INIT('h01)
	) name2462 (
		_w4343_,
		_w4355_,
		_w4362_,
		_w4363_
	);
	LUT3 #(
		.INIT('h20)
	) name2463 (
		\m2_s12_cyc_o_reg/NET0131 ,
		\rf_conf12_reg[4]/NET0131 ,
		\rf_conf12_reg[5]/NET0131 ,
		_w4364_
	);
	LUT3 #(
		.INIT('h20)
	) name2464 (
		\m3_s12_cyc_o_reg/NET0131 ,
		\rf_conf12_reg[6]/NET0131 ,
		\rf_conf12_reg[7]/NET0131 ,
		_w4365_
	);
	LUT2 #(
		.INIT('h2)
	) name2465 (
		\s12_msel_arb2_state_reg[1]/NET0131 ,
		\s12_msel_arb2_state_reg[2]/NET0131 ,
		_w4366_
	);
	LUT3 #(
		.INIT('h40)
	) name2466 (
		_w4364_,
		_w4365_,
		_w4366_,
		_w4367_
	);
	LUT3 #(
		.INIT('h20)
	) name2467 (
		\m5_s12_cyc_o_reg/NET0131 ,
		\rf_conf12_reg[10]/NET0131 ,
		\rf_conf12_reg[11]/NET0131 ,
		_w4368_
	);
	LUT3 #(
		.INIT('h20)
	) name2468 (
		\m7_s12_cyc_o_reg/NET0131 ,
		\rf_conf12_reg[14]/NET0131 ,
		\rf_conf12_reg[15]/NET0131 ,
		_w4369_
	);
	LUT3 #(
		.INIT('h20)
	) name2469 (
		\m6_s12_cyc_o_reg/NET0131 ,
		\rf_conf12_reg[12]/NET0131 ,
		\rf_conf12_reg[13]/NET0131 ,
		_w4370_
	);
	LUT3 #(
		.INIT('h51)
	) name2470 (
		_w4368_,
		_w4369_,
		_w4370_,
		_w4371_
	);
	LUT3 #(
		.INIT('h20)
	) name2471 (
		\m1_s12_cyc_o_reg/NET0131 ,
		\rf_conf12_reg[2]/NET0131 ,
		\rf_conf12_reg[3]/NET0131 ,
		_w4372_
	);
	LUT3 #(
		.INIT('h20)
	) name2472 (
		\m0_s12_cyc_o_reg/NET0131 ,
		\rf_conf12_reg[0]/NET0131 ,
		\rf_conf12_reg[1]/NET0131 ,
		_w4373_
	);
	LUT2 #(
		.INIT('h1)
	) name2473 (
		_w4370_,
		_w4373_,
		_w4374_
	);
	LUT3 #(
		.INIT('h04)
	) name2474 (
		_w4370_,
		_w4372_,
		_w4373_,
		_w4375_
	);
	LUT3 #(
		.INIT('h20)
	) name2475 (
		\m4_s12_cyc_o_reg/NET0131 ,
		\rf_conf12_reg[8]/NET0131 ,
		\rf_conf12_reg[9]/NET0131 ,
		_w4376_
	);
	LUT2 #(
		.INIT('h1)
	) name2476 (
		_w4364_,
		_w4376_,
		_w4377_
	);
	LUT3 #(
		.INIT('h04)
	) name2477 (
		_w4364_,
		_w4366_,
		_w4376_,
		_w4378_
	);
	LUT4 #(
		.INIT('h0455)
	) name2478 (
		_w4367_,
		_w4371_,
		_w4375_,
		_w4378_,
		_w4379_
	);
	LUT3 #(
		.INIT('h0b)
	) name2479 (
		_w4364_,
		_w4365_,
		_w4372_,
		_w4380_
	);
	LUT2 #(
		.INIT('h1)
	) name2480 (
		\s12_msel_arb2_state_reg[1]/NET0131 ,
		\s12_msel_arb2_state_reg[2]/NET0131 ,
		_w4381_
	);
	LUT2 #(
		.INIT('h4)
	) name2481 (
		_w4373_,
		_w4381_,
		_w4382_
	);
	LUT4 #(
		.INIT('hb0ff)
	) name2482 (
		_w4371_,
		_w4377_,
		_w4380_,
		_w4382_,
		_w4383_
	);
	LUT3 #(
		.INIT('h40)
	) name2483 (
		\s12_msel_arb2_state_reg[0]/NET0131 ,
		_w4379_,
		_w4383_,
		_w4384_
	);
	LUT2 #(
		.INIT('h8)
	) name2484 (
		\s12_msel_arb2_state_reg[1]/NET0131 ,
		\s12_msel_arb2_state_reg[2]/NET0131 ,
		_w4385_
	);
	LUT3 #(
		.INIT('h20)
	) name2485 (
		_w4369_,
		_w4370_,
		_w4385_,
		_w4386_
	);
	LUT3 #(
		.INIT('h04)
	) name2486 (
		_w4364_,
		_w4368_,
		_w4376_,
		_w4387_
	);
	LUT3 #(
		.INIT('h10)
	) name2487 (
		_w4370_,
		_w4373_,
		_w4385_,
		_w4388_
	);
	LUT4 #(
		.INIT('h0233)
	) name2488 (
		_w4380_,
		_w4386_,
		_w4387_,
		_w4388_,
		_w4389_
	);
	LUT2 #(
		.INIT('h4)
	) name2489 (
		\s12_msel_arb2_state_reg[1]/NET0131 ,
		\s12_msel_arb2_state_reg[2]/NET0131 ,
		_w4390_
	);
	LUT3 #(
		.INIT('h20)
	) name2490 (
		_w4368_,
		_w4376_,
		_w4390_,
		_w4391_
	);
	LUT2 #(
		.INIT('h4)
	) name2491 (
		_w4369_,
		_w4373_,
		_w4392_
	);
	LUT4 #(
		.INIT('h000b)
	) name2492 (
		_w4364_,
		_w4365_,
		_w4369_,
		_w4372_,
		_w4393_
	);
	LUT3 #(
		.INIT('h10)
	) name2493 (
		_w4370_,
		_w4376_,
		_w4390_,
		_w4394_
	);
	LUT4 #(
		.INIT('h5455)
	) name2494 (
		_w4391_,
		_w4392_,
		_w4393_,
		_w4394_,
		_w4395_
	);
	LUT2 #(
		.INIT('h8)
	) name2495 (
		_w4389_,
		_w4395_,
		_w4396_
	);
	LUT4 #(
		.INIT('hdf00)
	) name2496 (
		\m0_s12_cyc_o_reg/NET0131 ,
		\rf_conf12_reg[0]/NET0131 ,
		\rf_conf12_reg[1]/NET0131 ,
		\s12_msel_arb2_state_reg[0]/NET0131 ,
		_w4397_
	);
	LUT3 #(
		.INIT('h10)
	) name2497 (
		_w4364_,
		_w4376_,
		_w4397_,
		_w4398_
	);
	LUT3 #(
		.INIT('h20)
	) name2498 (
		\s12_msel_arb2_state_reg[0]/NET0131 ,
		\s12_msel_arb2_state_reg[1]/NET0131 ,
		\s12_msel_arb2_state_reg[2]/NET0131 ,
		_w4399_
	);
	LUT3 #(
		.INIT('h10)
	) name2499 (
		_w4368_,
		_w4370_,
		_w4399_,
		_w4400_
	);
	LUT4 #(
		.INIT('hf100)
	) name2500 (
		_w4392_,
		_w4393_,
		_w4398_,
		_w4400_,
		_w4401_
	);
	LUT3 #(
		.INIT('h08)
	) name2501 (
		_w4384_,
		_w4396_,
		_w4401_,
		_w4402_
	);
	LUT3 #(
		.INIT('hb0)
	) name2502 (
		_w4371_,
		_w4377_,
		_w4380_,
		_w4403_
	);
	LUT3 #(
		.INIT('h02)
	) name2503 (
		\s12_msel_arb2_state_reg[0]/NET0131 ,
		_w4364_,
		_w4376_,
		_w4404_
	);
	LUT2 #(
		.INIT('h8)
	) name2504 (
		_w4374_,
		_w4404_,
		_w4405_
	);
	LUT3 #(
		.INIT('ha2)
	) name2505 (
		_w4381_,
		_w4403_,
		_w4405_,
		_w4406_
	);
	LUT2 #(
		.INIT('h8)
	) name2506 (
		_w4365_,
		_w4366_,
		_w4407_
	);
	LUT4 #(
		.INIT('h0031)
	) name2507 (
		_w4364_,
		_w4370_,
		_w4372_,
		_w4373_,
		_w4408_
	);
	LUT2 #(
		.INIT('h2)
	) name2508 (
		_w4366_,
		_w4376_,
		_w4409_
	);
	LUT4 #(
		.INIT('h0233)
	) name2509 (
		_w4371_,
		_w4407_,
		_w4408_,
		_w4409_,
		_w4410_
	);
	LUT3 #(
		.INIT('h2a)
	) name2510 (
		\s12_msel_arb2_state_reg[0]/NET0131 ,
		_w4368_,
		_w4390_,
		_w4411_
	);
	LUT2 #(
		.INIT('h8)
	) name2511 (
		_w4410_,
		_w4411_,
		_w4412_
	);
	LUT4 #(
		.INIT('hdf00)
	) name2512 (
		\m6_s12_cyc_o_reg/NET0131 ,
		\rf_conf12_reg[12]/NET0131 ,
		\rf_conf12_reg[13]/NET0131 ,
		\s12_msel_arb2_state_reg[0]/NET0131 ,
		_w4413_
	);
	LUT4 #(
		.INIT('h3233)
	) name2513 (
		_w4364_,
		_w4369_,
		_w4376_,
		_w4413_,
		_w4414_
	);
	LUT4 #(
		.INIT('h0d0f)
	) name2514 (
		_w4380_,
		_w4387_,
		_w4392_,
		_w4414_,
		_w4415_
	);
	LUT3 #(
		.INIT('h13)
	) name2515 (
		_w4385_,
		_w4401_,
		_w4415_,
		_w4416_
	);
	LUT3 #(
		.INIT('h40)
	) name2516 (
		_w4406_,
		_w4412_,
		_w4416_,
		_w4417_
	);
	LUT2 #(
		.INIT('h1)
	) name2517 (
		_w4402_,
		_w4417_,
		_w4418_
	);
	LUT2 #(
		.INIT('h2)
	) name2518 (
		\s12_msel_arb3_state_reg[1]/NET0131 ,
		\s12_msel_arb3_state_reg[2]/NET0131 ,
		_w4419_
	);
	LUT2 #(
		.INIT('h4)
	) name2519 (
		_w3255_,
		_w4419_,
		_w4420_
	);
	LUT2 #(
		.INIT('h1)
	) name2520 (
		_w3237_,
		_w3244_,
		_w4421_
	);
	LUT3 #(
		.INIT('hae)
	) name2521 (
		_w3237_,
		_w3244_,
		_w3245_,
		_w4422_
	);
	LUT2 #(
		.INIT('h1)
	) name2522 (
		_w3249_,
		_w3260_,
		_w4423_
	);
	LUT2 #(
		.INIT('h1)
	) name2523 (
		_w3245_,
		_w3250_,
		_w4424_
	);
	LUT4 #(
		.INIT('h7577)
	) name2524 (
		_w4420_,
		_w4422_,
		_w4423_,
		_w4424_,
		_w4425_
	);
	LUT3 #(
		.INIT('h0d)
	) name2525 (
		_w3247_,
		_w3248_,
		_w3249_,
		_w4426_
	);
	LUT4 #(
		.INIT('h00f2)
	) name2526 (
		_w3247_,
		_w3248_,
		_w3249_,
		_w3250_,
		_w4427_
	);
	LUT3 #(
		.INIT('h10)
	) name2527 (
		\s12_msel_arb3_state_reg[0]/NET0131 ,
		\s12_msel_arb3_state_reg[1]/NET0131 ,
		\s12_msel_arb3_state_reg[2]/NET0131 ,
		_w4428_
	);
	LUT4 #(
		.INIT('h2300)
	) name2528 (
		_w3237_,
		_w3238_,
		_w3245_,
		_w4428_,
		_w4429_
	);
	LUT3 #(
		.INIT('hd0)
	) name2529 (
		_w4421_,
		_w4427_,
		_w4429_,
		_w4430_
	);
	LUT3 #(
		.INIT('h0e)
	) name2530 (
		_w3238_,
		_w4425_,
		_w4430_,
		_w4431_
	);
	LUT2 #(
		.INIT('h1)
	) name2531 (
		\s12_msel_arb3_state_reg[1]/NET0131 ,
		\s12_msel_arb3_state_reg[2]/NET0131 ,
		_w4432_
	);
	LUT4 #(
		.INIT('h0080)
	) name2532 (
		\m0_s12_cyc_o_reg/NET0131 ,
		\rf_conf12_reg[0]/NET0131 ,
		\rf_conf12_reg[1]/NET0131 ,
		\s12_msel_arb3_state_reg[0]/NET0131 ,
		_w4433_
	);
	LUT2 #(
		.INIT('h2)
	) name2533 (
		_w4432_,
		_w4433_,
		_w4434_
	);
	LUT2 #(
		.INIT('h1)
	) name2534 (
		_w3238_,
		_w3248_,
		_w4435_
	);
	LUT4 #(
		.INIT('h4fcf)
	) name2535 (
		_w4422_,
		_w4426_,
		_w4434_,
		_w4435_,
		_w4436_
	);
	LUT3 #(
		.INIT('h20)
	) name2536 (
		_w3247_,
		_w3255_,
		_w4419_,
		_w4437_
	);
	LUT3 #(
		.INIT('h20)
	) name2537 (
		\s12_msel_arb3_state_reg[0]/NET0131 ,
		\s12_msel_arb3_state_reg[1]/NET0131 ,
		\s12_msel_arb3_state_reg[2]/NET0131 ,
		_w4438_
	);
	LUT2 #(
		.INIT('h8)
	) name2538 (
		_w3237_,
		_w4438_,
		_w4439_
	);
	LUT2 #(
		.INIT('h1)
	) name2539 (
		_w4437_,
		_w4439_,
		_w4440_
	);
	LUT2 #(
		.INIT('h8)
	) name2540 (
		_w4436_,
		_w4440_,
		_w4441_
	);
	LUT3 #(
		.INIT('h02)
	) name2541 (
		\s12_msel_arb3_state_reg[0]/NET0131 ,
		\s12_msel_arb3_state_reg[1]/NET0131 ,
		\s12_msel_arb3_state_reg[2]/NET0131 ,
		_w4442_
	);
	LUT4 #(
		.INIT('h0100)
	) name2542 (
		_w3238_,
		_w3248_,
		_w3250_,
		_w4442_,
		_w4443_
	);
	LUT2 #(
		.INIT('h4)
	) name2543 (
		_w3237_,
		_w4438_,
		_w4444_
	);
	LUT2 #(
		.INIT('h1)
	) name2544 (
		_w4443_,
		_w4444_,
		_w4445_
	);
	LUT2 #(
		.INIT('h4)
	) name2545 (
		_w3244_,
		_w3250_,
		_w4446_
	);
	LUT4 #(
		.INIT('h0051)
	) name2546 (
		_w3244_,
		_w3247_,
		_w3248_,
		_w3249_,
		_w4447_
	);
	LUT4 #(
		.INIT('h7f00)
	) name2547 (
		\m0_s12_cyc_o_reg/NET0131 ,
		\rf_conf12_reg[0]/NET0131 ,
		\rf_conf12_reg[1]/NET0131 ,
		\s12_msel_arb3_state_reg[0]/NET0131 ,
		_w4448_
	);
	LUT3 #(
		.INIT('h10)
	) name2548 (
		_w3238_,
		_w3248_,
		_w4448_,
		_w4449_
	);
	LUT4 #(
		.INIT('h0054)
	) name2549 (
		_w4443_,
		_w4446_,
		_w4447_,
		_w4449_,
		_w4450_
	);
	LUT3 #(
		.INIT('h01)
	) name2550 (
		_w3245_,
		_w4445_,
		_w4450_,
		_w4451_
	);
	LUT4 #(
		.INIT('h007f)
	) name2551 (
		\m5_s12_cyc_o_reg/NET0131 ,
		\rf_conf12_reg[10]/NET0131 ,
		\rf_conf12_reg[11]/NET0131 ,
		\s12_msel_arb3_state_reg[0]/NET0131 ,
		_w4452_
	);
	LUT4 #(
		.INIT('h0001)
	) name2552 (
		_w3238_,
		_w3248_,
		_w3250_,
		_w4452_,
		_w4453_
	);
	LUT3 #(
		.INIT('h0e)
	) name2553 (
		_w4446_,
		_w4447_,
		_w4453_,
		_w4454_
	);
	LUT4 #(
		.INIT('h0080)
	) name2554 (
		\m6_s12_cyc_o_reg/NET0131 ,
		\rf_conf12_reg[12]/NET0131 ,
		\rf_conf12_reg[13]/NET0131 ,
		\s12_msel_arb3_state_reg[0]/NET0131 ,
		_w4455_
	);
	LUT3 #(
		.INIT('h10)
	) name2555 (
		_w3237_,
		_w3244_,
		_w3245_,
		_w4456_
	);
	LUT4 #(
		.INIT('h020a)
	) name2556 (
		_w3263_,
		_w4426_,
		_w4455_,
		_w4456_,
		_w4457_
	);
	LUT2 #(
		.INIT('h4)
	) name2557 (
		_w4454_,
		_w4457_,
		_w4458_
	);
	LUT4 #(
		.INIT('hfff7)
	) name2558 (
		_w4431_,
		_w4441_,
		_w4451_,
		_w4458_,
		_w4459_
	);
	LUT2 #(
		.INIT('h4)
	) name2559 (
		_w2344_,
		_w2352_,
		_w4460_
	);
	LUT3 #(
		.INIT('h04)
	) name2560 (
		_w2340_,
		_w2342_,
		_w2343_,
		_w4461_
	);
	LUT4 #(
		.INIT('hfd00)
	) name2561 (
		\m4_s13_cyc_o_reg/NET0131 ,
		\rf_conf13_reg[8]/NET0131 ,
		\rf_conf13_reg[9]/NET0131 ,
		\s13_msel_arb0_state_reg[0]/NET0131 ,
		_w4462_
	);
	LUT3 #(
		.INIT('h10)
	) name2562 (
		_w2343_,
		_w2345_,
		_w4462_,
		_w4463_
	);
	LUT3 #(
		.INIT('hf2)
	) name2563 (
		_w2339_,
		_w2340_,
		_w2347_,
		_w4464_
	);
	LUT4 #(
		.INIT('h000d)
	) name2564 (
		_w2339_,
		_w2340_,
		_w2344_,
		_w2347_,
		_w4465_
	);
	LUT4 #(
		.INIT('h5455)
	) name2565 (
		_w4460_,
		_w4461_,
		_w4463_,
		_w4465_,
		_w4466_
	);
	LUT2 #(
		.INIT('h8)
	) name2566 (
		_w2366_,
		_w4466_,
		_w4467_
	);
	LUT2 #(
		.INIT('h8)
	) name2567 (
		\s13_msel_arb0_state_reg[1]/NET0131 ,
		\s13_msel_arb0_state_reg[2]/NET0131 ,
		_w4468_
	);
	LUT2 #(
		.INIT('h2)
	) name2568 (
		_w2347_,
		_w2352_,
		_w4469_
	);
	LUT3 #(
		.INIT('h51)
	) name2569 (
		_w2344_,
		_w2347_,
		_w2352_,
		_w4470_
	);
	LUT4 #(
		.INIT('h2232)
	) name2570 (
		_w2344_,
		_w2345_,
		_w2347_,
		_w2352_,
		_w4471_
	);
	LUT2 #(
		.INIT('h1)
	) name2571 (
		_w2340_,
		_w2352_,
		_w4472_
	);
	LUT4 #(
		.INIT('h00fd)
	) name2572 (
		\m5_s13_cyc_o_reg/NET0131 ,
		\rf_conf13_reg[10]/NET0131 ,
		\rf_conf13_reg[11]/NET0131 ,
		\s13_msel_arb0_state_reg[0]/NET0131 ,
		_w4473_
	);
	LUT3 #(
		.INIT('h01)
	) name2573 (
		_w2340_,
		_w2352_,
		_w4473_,
		_w4474_
	);
	LUT2 #(
		.INIT('h4)
	) name2574 (
		_w2339_,
		_w2343_,
		_w4475_
	);
	LUT3 #(
		.INIT('h0b)
	) name2575 (
		_w2339_,
		_w2343_,
		_w2345_,
		_w4476_
	);
	LUT4 #(
		.INIT('h0111)
	) name2576 (
		_w2342_,
		_w4471_,
		_w4474_,
		_w4476_,
		_w4477_
	);
	LUT4 #(
		.INIT('h1101)
	) name2577 (
		_w2339_,
		_w2342_,
		_w2344_,
		_w2345_,
		_w4478_
	);
	LUT4 #(
		.INIT('hfd00)
	) name2578 (
		\m2_s13_cyc_o_reg/NET0131 ,
		\rf_conf13_reg[4]/NET0131 ,
		\rf_conf13_reg[5]/NET0131 ,
		\s13_msel_arb0_state_reg[0]/NET0131 ,
		_w4479_
	);
	LUT4 #(
		.INIT('h0e0f)
	) name2579 (
		_w2343_,
		_w2345_,
		_w2347_,
		_w4479_,
		_w4480_
	);
	LUT2 #(
		.INIT('h2)
	) name2580 (
		\s13_msel_arb0_state_reg[1]/NET0131 ,
		\s13_msel_arb0_state_reg[2]/NET0131 ,
		_w4481_
	);
	LUT3 #(
		.INIT('hd0)
	) name2581 (
		_w2340_,
		_w2347_,
		_w4481_,
		_w4482_
	);
	LUT4 #(
		.INIT('h1f00)
	) name2582 (
		_w4475_,
		_w4478_,
		_w4480_,
		_w4482_,
		_w4483_
	);
	LUT3 #(
		.INIT('h0d)
	) name2583 (
		_w4468_,
		_w4477_,
		_w4483_,
		_w4484_
	);
	LUT3 #(
		.INIT('h8a)
	) name2584 (
		\s13_msel_arb0_state_reg[0]/NET0131 ,
		_w4467_,
		_w4484_,
		_w4485_
	);
	LUT3 #(
		.INIT('h02)
	) name2585 (
		\s13_msel_arb0_state_reg[0]/NET0131 ,
		_w2343_,
		_w2345_,
		_w4486_
	);
	LUT4 #(
		.INIT('h55fd)
	) name2586 (
		_w4472_,
		_w4475_,
		_w4478_,
		_w4486_,
		_w4487_
	);
	LUT3 #(
		.INIT('h8c)
	) name2587 (
		_w4469_,
		_w4481_,
		_w4487_,
		_w4488_
	);
	LUT3 #(
		.INIT('h20)
	) name2588 (
		_w2342_,
		_w2343_,
		_w4468_,
		_w4489_
	);
	LUT3 #(
		.INIT('h10)
	) name2589 (
		_w2343_,
		_w2345_,
		_w4468_,
		_w4490_
	);
	LUT4 #(
		.INIT('h020f)
	) name2590 (
		_w4470_,
		_w4474_,
		_w4489_,
		_w4490_,
		_w4491_
	);
	LUT3 #(
		.INIT('h20)
	) name2591 (
		_w2344_,
		_w2345_,
		_w2366_,
		_w4492_
	);
	LUT2 #(
		.INIT('h1)
	) name2592 (
		_w2340_,
		_w2343_,
		_w4493_
	);
	LUT4 #(
		.INIT('h00fd)
	) name2593 (
		\m7_s13_cyc_o_reg/NET0131 ,
		\rf_conf13_reg[14]/NET0131 ,
		\rf_conf13_reg[15]/NET0131 ,
		\s13_msel_arb0_state_reg[0]/NET0131 ,
		_w4494_
	);
	LUT3 #(
		.INIT('h01)
	) name2594 (
		_w2340_,
		_w2343_,
		_w4494_,
		_w4495_
	);
	LUT3 #(
		.INIT('h10)
	) name2595 (
		_w2345_,
		_w2352_,
		_w2366_,
		_w4496_
	);
	LUT4 #(
		.INIT('h0133)
	) name2596 (
		_w4464_,
		_w4492_,
		_w4495_,
		_w4496_,
		_w4497_
	);
	LUT2 #(
		.INIT('h8)
	) name2597 (
		_w4491_,
		_w4497_,
		_w4498_
	);
	LUT3 #(
		.INIT('h02)
	) name2598 (
		\s13_msel_arb0_state_reg[0]/NET0131 ,
		_w2345_,
		_w2352_,
		_w4499_
	);
	LUT3 #(
		.INIT('h80)
	) name2599 (
		_w2369_,
		_w4493_,
		_w4499_,
		_w4500_
	);
	LUT3 #(
		.INIT('h04)
	) name2600 (
		_w2345_,
		_w2347_,
		_w2352_,
		_w4501_
	);
	LUT4 #(
		.INIT('h0002)
	) name2601 (
		\m4_s13_cyc_o_reg/NET0131 ,
		\rf_conf13_reg[8]/NET0131 ,
		\rf_conf13_reg[9]/NET0131 ,
		\s13_msel_arb0_state_reg[0]/NET0131 ,
		_w4502_
	);
	LUT4 #(
		.INIT('h00b0)
	) name2602 (
		_w2339_,
		_w2343_,
		_w2369_,
		_w4502_,
		_w4503_
	);
	LUT3 #(
		.INIT('hd0)
	) name2603 (
		_w4478_,
		_w4501_,
		_w4503_,
		_w4504_
	);
	LUT2 #(
		.INIT('h1)
	) name2604 (
		_w4500_,
		_w4504_,
		_w4505_
	);
	LUT4 #(
		.INIT('hba00)
	) name2605 (
		\s13_msel_arb0_state_reg[0]/NET0131 ,
		_w4488_,
		_w4498_,
		_w4505_,
		_w4506_
	);
	LUT2 #(
		.INIT('hb)
	) name2606 (
		_w4485_,
		_w4506_,
		_w4507_
	);
	LUT3 #(
		.INIT('h23)
	) name2607 (
		_w3645_,
		_w3647_,
		_w3657_,
		_w4508_
	);
	LUT4 #(
		.INIT('h2232)
	) name2608 (
		_w3645_,
		_w3647_,
		_w3656_,
		_w3657_,
		_w4509_
	);
	LUT2 #(
		.INIT('h1)
	) name2609 (
		_w3647_,
		_w3657_,
		_w4510_
	);
	LUT4 #(
		.INIT('h0004)
	) name2610 (
		_w3647_,
		_w3653_,
		_w3654_,
		_w3657_,
		_w4511_
	);
	LUT2 #(
		.INIT('h2)
	) name2611 (
		\s13_msel_arb1_state_reg[1]/NET0131 ,
		\s13_msel_arb1_state_reg[2]/NET0131 ,
		_w4512_
	);
	LUT2 #(
		.INIT('h4)
	) name2612 (
		_w3650_,
		_w4512_,
		_w4513_
	);
	LUT4 #(
		.INIT('hfe00)
	) name2613 (
		_w3651_,
		_w4509_,
		_w4511_,
		_w4513_,
		_w4514_
	);
	LUT3 #(
		.INIT('hdc)
	) name2614 (
		_w3645_,
		_w3647_,
		_w3657_,
		_w4515_
	);
	LUT2 #(
		.INIT('h2)
	) name2615 (
		_w3654_,
		_w3656_,
		_w4516_
	);
	LUT2 #(
		.INIT('h4)
	) name2616 (
		_w3650_,
		_w3651_,
		_w4517_
	);
	LUT4 #(
		.INIT('h000b)
	) name2617 (
		_w3650_,
		_w3651_,
		_w3653_,
		_w3656_,
		_w4518_
	);
	LUT4 #(
		.INIT('hf700)
	) name2618 (
		\m0_s13_cyc_o_reg/NET0131 ,
		\rf_conf13_reg[0]/NET0131 ,
		\rf_conf13_reg[1]/NET0131 ,
		\s13_msel_arb1_state_reg[0]/NET0131 ,
		_w4519_
	);
	LUT4 #(
		.INIT('hd0dd)
	) name2619 (
		_w3645_,
		_w3647_,
		_w3650_,
		_w4519_,
		_w4520_
	);
	LUT4 #(
		.INIT('h0155)
	) name2620 (
		_w4515_,
		_w4516_,
		_w4518_,
		_w4520_,
		_w4521_
	);
	LUT2 #(
		.INIT('h4)
	) name2621 (
		\s13_msel_arb1_state_reg[1]/NET0131 ,
		\s13_msel_arb1_state_reg[2]/NET0131 ,
		_w4522_
	);
	LUT4 #(
		.INIT('habbb)
	) name2622 (
		\s13_msel_arb1_state_reg[0]/NET0131 ,
		_w4514_,
		_w4521_,
		_w4522_,
		_w4523_
	);
	LUT4 #(
		.INIT('hff0d)
	) name2623 (
		\s13_msel_arb1_state_reg[0]/NET0131 ,
		_w3650_,
		_w3653_,
		_w3654_,
		_w4524_
	);
	LUT4 #(
		.INIT('h1101)
	) name2624 (
		_w3651_,
		_w4509_,
		_w4510_,
		_w4524_,
		_w4525_
	);
	LUT2 #(
		.INIT('h2)
	) name2625 (
		_w4512_,
		_w4525_,
		_w4526_
	);
	LUT2 #(
		.INIT('h1)
	) name2626 (
		\s13_msel_arb1_state_reg[1]/NET0131 ,
		\s13_msel_arb1_state_reg[2]/NET0131 ,
		_w4527_
	);
	LUT3 #(
		.INIT('h0b)
	) name2627 (
		_w3650_,
		_w3651_,
		_w3653_,
		_w4528_
	);
	LUT3 #(
		.INIT('h02)
	) name2628 (
		_w3645_,
		_w3647_,
		_w3650_,
		_w4529_
	);
	LUT3 #(
		.INIT('h01)
	) name2629 (
		_w3647_,
		_w3650_,
		_w3657_,
		_w4530_
	);
	LUT2 #(
		.INIT('h1)
	) name2630 (
		_w3656_,
		_w4519_,
		_w4531_
	);
	LUT4 #(
		.INIT('h2202)
	) name2631 (
		_w4528_,
		_w4529_,
		_w4530_,
		_w4531_,
		_w4532_
	);
	LUT4 #(
		.INIT('h5455)
	) name2632 (
		_w3645_,
		_w3647_,
		_w3650_,
		_w4519_,
		_w4533_
	);
	LUT3 #(
		.INIT('hb0)
	) name2633 (
		_w3645_,
		_w3657_,
		_w4522_,
		_w4534_
	);
	LUT4 #(
		.INIT('h1f00)
	) name2634 (
		_w4516_,
		_w4518_,
		_w4533_,
		_w4534_,
		_w4535_
	);
	LUT3 #(
		.INIT('h0d)
	) name2635 (
		_w4527_,
		_w4532_,
		_w4535_,
		_w4536_
	);
	LUT3 #(
		.INIT('h8a)
	) name2636 (
		\s13_msel_arb1_state_reg[0]/NET0131 ,
		_w4526_,
		_w4536_,
		_w4537_
	);
	LUT4 #(
		.INIT('h0008)
	) name2637 (
		\m6_s13_cyc_o_reg/NET0131 ,
		\rf_conf13_reg[12]/NET0131 ,
		\rf_conf13_reg[13]/NET0131 ,
		\s13_msel_arb1_state_reg[0]/NET0131 ,
		_w4538_
	);
	LUT2 #(
		.INIT('h8)
	) name2638 (
		\s13_msel_arb1_state_reg[1]/NET0131 ,
		\s13_msel_arb1_state_reg[2]/NET0131 ,
		_w4539_
	);
	LUT2 #(
		.INIT('h4)
	) name2639 (
		_w4538_,
		_w4539_,
		_w4540_
	);
	LUT3 #(
		.INIT('h20)
	) name2640 (
		_w3656_,
		_w4538_,
		_w4539_,
		_w4541_
	);
	LUT4 #(
		.INIT('hf700)
	) name2641 (
		\m2_s13_cyc_o_reg/NET0131 ,
		\rf_conf13_reg[4]/NET0131 ,
		\rf_conf13_reg[5]/NET0131 ,
		\s13_msel_arb1_state_reg[0]/NET0131 ,
		_w4542_
	);
	LUT3 #(
		.INIT('h10)
	) name2642 (
		_w3647_,
		_w3657_,
		_w4542_,
		_w4543_
	);
	LUT4 #(
		.INIT('hf0d0)
	) name2643 (
		_w4528_,
		_w4529_,
		_w4540_,
		_w4543_,
		_w4544_
	);
	LUT3 #(
		.INIT('h32)
	) name2644 (
		_w3645_,
		_w3650_,
		_w3656_,
		_w4545_
	);
	LUT4 #(
		.INIT('h0105)
	) name2645 (
		_w3653_,
		_w4508_,
		_w4517_,
		_w4545_,
		_w4546_
	);
	LUT3 #(
		.INIT('h01)
	) name2646 (
		\s13_msel_arb1_state_reg[0]/NET0131 ,
		\s13_msel_arb1_state_reg[1]/NET0131 ,
		\s13_msel_arb1_state_reg[2]/NET0131 ,
		_w4547_
	);
	LUT4 #(
		.INIT('hbabb)
	) name2647 (
		_w3654_,
		_w4544_,
		_w4546_,
		_w4547_,
		_w4548_
	);
	LUT2 #(
		.INIT('h4)
	) name2648 (
		_w4541_,
		_w4548_,
		_w4549_
	);
	LUT3 #(
		.INIT('hdf)
	) name2649 (
		_w4523_,
		_w4537_,
		_w4549_,
		_w4550_
	);
	LUT3 #(
		.INIT('h20)
	) name2650 (
		\m4_s13_cyc_o_reg/NET0131 ,
		\rf_conf13_reg[8]/NET0131 ,
		\rf_conf13_reg[9]/NET0131 ,
		_w4551_
	);
	LUT3 #(
		.INIT('h20)
	) name2651 (
		\m7_s13_cyc_o_reg/NET0131 ,
		\rf_conf13_reg[14]/NET0131 ,
		\rf_conf13_reg[15]/NET0131 ,
		_w4552_
	);
	LUT3 #(
		.INIT('h20)
	) name2652 (
		\m0_s13_cyc_o_reg/NET0131 ,
		\rf_conf13_reg[0]/NET0131 ,
		\rf_conf13_reg[1]/NET0131 ,
		_w4553_
	);
	LUT2 #(
		.INIT('h4)
	) name2653 (
		_w4552_,
		_w4553_,
		_w4554_
	);
	LUT3 #(
		.INIT('h20)
	) name2654 (
		\m3_s13_cyc_o_reg/NET0131 ,
		\rf_conf13_reg[6]/NET0131 ,
		\rf_conf13_reg[7]/NET0131 ,
		_w4555_
	);
	LUT3 #(
		.INIT('h20)
	) name2655 (
		\m2_s13_cyc_o_reg/NET0131 ,
		\rf_conf13_reg[4]/NET0131 ,
		\rf_conf13_reg[5]/NET0131 ,
		_w4556_
	);
	LUT3 #(
		.INIT('h20)
	) name2656 (
		\m1_s13_cyc_o_reg/NET0131 ,
		\rf_conf13_reg[2]/NET0131 ,
		\rf_conf13_reg[3]/NET0131 ,
		_w4557_
	);
	LUT4 #(
		.INIT('h0051)
	) name2657 (
		_w4552_,
		_w4555_,
		_w4556_,
		_w4557_,
		_w4558_
	);
	LUT3 #(
		.INIT('h20)
	) name2658 (
		\m5_s13_cyc_o_reg/NET0131 ,
		\rf_conf13_reg[10]/NET0131 ,
		\rf_conf13_reg[11]/NET0131 ,
		_w4559_
	);
	LUT3 #(
		.INIT('h20)
	) name2659 (
		\m6_s13_cyc_o_reg/NET0131 ,
		\rf_conf13_reg[12]/NET0131 ,
		\rf_conf13_reg[13]/NET0131 ,
		_w4560_
	);
	LUT3 #(
		.INIT('h8a)
	) name2660 (
		\s13_msel_arb2_state_reg[0]/NET0131 ,
		_w4559_,
		_w4560_,
		_w4561_
	);
	LUT4 #(
		.INIT('hf100)
	) name2661 (
		_w4554_,
		_w4558_,
		_w4559_,
		_w4561_,
		_w4562_
	);
	LUT2 #(
		.INIT('h1)
	) name2662 (
		_w4553_,
		_w4560_,
		_w4563_
	);
	LUT4 #(
		.INIT('hdf00)
	) name2663 (
		\m2_s13_cyc_o_reg/NET0131 ,
		\rf_conf13_reg[4]/NET0131 ,
		\rf_conf13_reg[5]/NET0131 ,
		\s13_msel_arb2_state_reg[0]/NET0131 ,
		_w4564_
	);
	LUT4 #(
		.INIT('h3030)
	) name2664 (
		_w4553_,
		_w4559_,
		_w4560_,
		_w4564_,
		_w4565_
	);
	LUT4 #(
		.INIT('h3233)
	) name2665 (
		_w4553_,
		_w4559_,
		_w4560_,
		_w4564_,
		_w4566_
	);
	LUT4 #(
		.INIT('h010f)
	) name2666 (
		_w4554_,
		_w4558_,
		_w4565_,
		_w4566_,
		_w4567_
	);
	LUT2 #(
		.INIT('h4)
	) name2667 (
		\s13_msel_arb2_state_reg[1]/NET0131 ,
		\s13_msel_arb2_state_reg[2]/NET0131 ,
		_w4568_
	);
	LUT4 #(
		.INIT('hd000)
	) name2668 (
		_w4551_,
		_w4562_,
		_w4567_,
		_w4568_,
		_w4569_
	);
	LUT2 #(
		.INIT('h8)
	) name2669 (
		\s13_msel_arb2_state_reg[1]/NET0131 ,
		\s13_msel_arb2_state_reg[2]/NET0131 ,
		_w4570_
	);
	LUT3 #(
		.INIT('h20)
	) name2670 (
		_w4552_,
		_w4560_,
		_w4570_,
		_w4571_
	);
	LUT3 #(
		.INIT('h0d)
	) name2671 (
		_w4555_,
		_w4556_,
		_w4557_,
		_w4572_
	);
	LUT4 #(
		.INIT('h00df)
	) name2672 (
		\m5_s13_cyc_o_reg/NET0131 ,
		\rf_conf13_reg[10]/NET0131 ,
		\rf_conf13_reg[11]/NET0131 ,
		\s13_msel_arb2_state_reg[0]/NET0131 ,
		_w4573_
	);
	LUT3 #(
		.INIT('h01)
	) name2673 (
		_w4551_,
		_w4556_,
		_w4573_,
		_w4574_
	);
	LUT3 #(
		.INIT('h10)
	) name2674 (
		_w4553_,
		_w4560_,
		_w4570_,
		_w4575_
	);
	LUT4 #(
		.INIT('h0455)
	) name2675 (
		_w4571_,
		_w4572_,
		_w4574_,
		_w4575_,
		_w4576_
	);
	LUT2 #(
		.INIT('h1)
	) name2676 (
		\s13_msel_arb2_state_reg[1]/NET0131 ,
		\s13_msel_arb2_state_reg[2]/NET0131 ,
		_w4577_
	);
	LUT3 #(
		.INIT('h40)
	) name2677 (
		_w4553_,
		_w4557_,
		_w4577_,
		_w4578_
	);
	LUT2 #(
		.INIT('h2)
	) name2678 (
		_w4551_,
		_w4555_,
		_w4579_
	);
	LUT4 #(
		.INIT('h0301)
	) name2679 (
		_w4552_,
		_w4555_,
		_w4559_,
		_w4560_,
		_w4580_
	);
	LUT3 #(
		.INIT('h10)
	) name2680 (
		_w4553_,
		_w4556_,
		_w4577_,
		_w4581_
	);
	LUT4 #(
		.INIT('h5455)
	) name2681 (
		_w4578_,
		_w4579_,
		_w4580_,
		_w4581_,
		_w4582_
	);
	LUT3 #(
		.INIT('h15)
	) name2682 (
		\s13_msel_arb2_state_reg[0]/NET0131 ,
		_w4576_,
		_w4582_,
		_w4583_
	);
	LUT3 #(
		.INIT('h80)
	) name2683 (
		\s13_msel_arb2_state_reg[0]/NET0131 ,
		_w4557_,
		_w4577_,
		_w4584_
	);
	LUT3 #(
		.INIT('h45)
	) name2684 (
		_w4553_,
		_w4559_,
		_w4560_,
		_w4585_
	);
	LUT4 #(
		.INIT('h0eee)
	) name2685 (
		_w4554_,
		_w4558_,
		_w4574_,
		_w4585_,
		_w4586_
	);
	LUT3 #(
		.INIT('h80)
	) name2686 (
		\s13_msel_arb2_state_reg[0]/NET0131 ,
		\s13_msel_arb2_state_reg[1]/NET0131 ,
		\s13_msel_arb2_state_reg[2]/NET0131 ,
		_w4587_
	);
	LUT3 #(
		.INIT('h45)
	) name2687 (
		_w4584_,
		_w4586_,
		_w4587_,
		_w4588_
	);
	LUT3 #(
		.INIT('h40)
	) name2688 (
		_w4557_,
		_w4564_,
		_w4577_,
		_w4589_
	);
	LUT4 #(
		.INIT('h0020)
	) name2689 (
		\m2_s13_cyc_o_reg/NET0131 ,
		\rf_conf13_reg[4]/NET0131 ,
		\rf_conf13_reg[5]/NET0131 ,
		\s13_msel_arb2_state_reg[0]/NET0131 ,
		_w4590_
	);
	LUT2 #(
		.INIT('h2)
	) name2690 (
		\s13_msel_arb2_state_reg[1]/NET0131 ,
		\s13_msel_arb2_state_reg[2]/NET0131 ,
		_w4591_
	);
	LUT2 #(
		.INIT('h4)
	) name2691 (
		_w4590_,
		_w4591_,
		_w4592_
	);
	LUT4 #(
		.INIT('h1110)
	) name2692 (
		_w4579_,
		_w4580_,
		_w4589_,
		_w4592_,
		_w4593_
	);
	LUT3 #(
		.INIT('h40)
	) name2693 (
		_w4551_,
		_w4563_,
		_w4589_,
		_w4594_
	);
	LUT4 #(
		.INIT('hfafb)
	) name2694 (
		_w4553_,
		_w4557_,
		_w4560_,
		_w4564_,
		_w4595_
	);
	LUT3 #(
		.INIT('h10)
	) name2695 (
		_w4551_,
		_w4590_,
		_w4591_,
		_w4596_
	);
	LUT2 #(
		.INIT('h4)
	) name2696 (
		_w4595_,
		_w4596_,
		_w4597_
	);
	LUT3 #(
		.INIT('h01)
	) name2697 (
		_w4593_,
		_w4594_,
		_w4597_,
		_w4598_
	);
	LUT4 #(
		.INIT('hefff)
	) name2698 (
		_w4569_,
		_w4583_,
		_w4588_,
		_w4598_,
		_w4599_
	);
	LUT2 #(
		.INIT('h2)
	) name2699 (
		\s13_msel_arb3_state_reg[1]/NET0131 ,
		\s13_msel_arb3_state_reg[2]/NET0131 ,
		_w4600_
	);
	LUT2 #(
		.INIT('h4)
	) name2700 (
		_w2961_,
		_w4600_,
		_w4601_
	);
	LUT2 #(
		.INIT('h1)
	) name2701 (
		_w2943_,
		_w2950_,
		_w4602_
	);
	LUT3 #(
		.INIT('hae)
	) name2702 (
		_w2943_,
		_w2950_,
		_w2951_,
		_w4603_
	);
	LUT2 #(
		.INIT('h1)
	) name2703 (
		_w2955_,
		_w2966_,
		_w4604_
	);
	LUT2 #(
		.INIT('h1)
	) name2704 (
		_w2951_,
		_w2956_,
		_w4605_
	);
	LUT4 #(
		.INIT('h7577)
	) name2705 (
		_w4601_,
		_w4603_,
		_w4604_,
		_w4605_,
		_w4606_
	);
	LUT3 #(
		.INIT('h0d)
	) name2706 (
		_w2953_,
		_w2954_,
		_w2955_,
		_w4607_
	);
	LUT4 #(
		.INIT('h00f2)
	) name2707 (
		_w2953_,
		_w2954_,
		_w2955_,
		_w2956_,
		_w4608_
	);
	LUT3 #(
		.INIT('h10)
	) name2708 (
		\s13_msel_arb3_state_reg[0]/NET0131 ,
		\s13_msel_arb3_state_reg[1]/NET0131 ,
		\s13_msel_arb3_state_reg[2]/NET0131 ,
		_w4609_
	);
	LUT4 #(
		.INIT('h2300)
	) name2709 (
		_w2943_,
		_w2944_,
		_w2951_,
		_w4609_,
		_w4610_
	);
	LUT3 #(
		.INIT('hd0)
	) name2710 (
		_w4602_,
		_w4608_,
		_w4610_,
		_w4611_
	);
	LUT3 #(
		.INIT('h0e)
	) name2711 (
		_w2944_,
		_w4606_,
		_w4611_,
		_w4612_
	);
	LUT2 #(
		.INIT('h1)
	) name2712 (
		\s13_msel_arb3_state_reg[1]/NET0131 ,
		\s13_msel_arb3_state_reg[2]/NET0131 ,
		_w4613_
	);
	LUT4 #(
		.INIT('h0080)
	) name2713 (
		\m0_s13_cyc_o_reg/NET0131 ,
		\rf_conf13_reg[0]/NET0131 ,
		\rf_conf13_reg[1]/NET0131 ,
		\s13_msel_arb3_state_reg[0]/NET0131 ,
		_w4614_
	);
	LUT2 #(
		.INIT('h2)
	) name2714 (
		_w4613_,
		_w4614_,
		_w4615_
	);
	LUT2 #(
		.INIT('h1)
	) name2715 (
		_w2944_,
		_w2954_,
		_w4616_
	);
	LUT4 #(
		.INIT('h4fcf)
	) name2716 (
		_w4603_,
		_w4607_,
		_w4615_,
		_w4616_,
		_w4617_
	);
	LUT3 #(
		.INIT('h20)
	) name2717 (
		_w2953_,
		_w2961_,
		_w4600_,
		_w4618_
	);
	LUT3 #(
		.INIT('h20)
	) name2718 (
		\s13_msel_arb3_state_reg[0]/NET0131 ,
		\s13_msel_arb3_state_reg[1]/NET0131 ,
		\s13_msel_arb3_state_reg[2]/NET0131 ,
		_w4619_
	);
	LUT2 #(
		.INIT('h8)
	) name2719 (
		_w2943_,
		_w4619_,
		_w4620_
	);
	LUT2 #(
		.INIT('h1)
	) name2720 (
		_w4618_,
		_w4620_,
		_w4621_
	);
	LUT2 #(
		.INIT('h8)
	) name2721 (
		_w4617_,
		_w4621_,
		_w4622_
	);
	LUT3 #(
		.INIT('h02)
	) name2722 (
		\s13_msel_arb3_state_reg[0]/NET0131 ,
		\s13_msel_arb3_state_reg[1]/NET0131 ,
		\s13_msel_arb3_state_reg[2]/NET0131 ,
		_w4623_
	);
	LUT4 #(
		.INIT('h0100)
	) name2723 (
		_w2944_,
		_w2954_,
		_w2956_,
		_w4623_,
		_w4624_
	);
	LUT2 #(
		.INIT('h4)
	) name2724 (
		_w2943_,
		_w4619_,
		_w4625_
	);
	LUT2 #(
		.INIT('h1)
	) name2725 (
		_w4624_,
		_w4625_,
		_w4626_
	);
	LUT2 #(
		.INIT('h4)
	) name2726 (
		_w2950_,
		_w2956_,
		_w4627_
	);
	LUT4 #(
		.INIT('h0051)
	) name2727 (
		_w2950_,
		_w2953_,
		_w2954_,
		_w2955_,
		_w4628_
	);
	LUT4 #(
		.INIT('h7f00)
	) name2728 (
		\m0_s13_cyc_o_reg/NET0131 ,
		\rf_conf13_reg[0]/NET0131 ,
		\rf_conf13_reg[1]/NET0131 ,
		\s13_msel_arb3_state_reg[0]/NET0131 ,
		_w4629_
	);
	LUT3 #(
		.INIT('h10)
	) name2729 (
		_w2944_,
		_w2954_,
		_w4629_,
		_w4630_
	);
	LUT4 #(
		.INIT('h0054)
	) name2730 (
		_w4624_,
		_w4627_,
		_w4628_,
		_w4630_,
		_w4631_
	);
	LUT3 #(
		.INIT('h01)
	) name2731 (
		_w2951_,
		_w4626_,
		_w4631_,
		_w4632_
	);
	LUT4 #(
		.INIT('h007f)
	) name2732 (
		\m5_s13_cyc_o_reg/NET0131 ,
		\rf_conf13_reg[10]/NET0131 ,
		\rf_conf13_reg[11]/NET0131 ,
		\s13_msel_arb3_state_reg[0]/NET0131 ,
		_w4633_
	);
	LUT4 #(
		.INIT('h0001)
	) name2733 (
		_w2944_,
		_w2954_,
		_w2956_,
		_w4633_,
		_w4634_
	);
	LUT3 #(
		.INIT('h0e)
	) name2734 (
		_w4627_,
		_w4628_,
		_w4634_,
		_w4635_
	);
	LUT4 #(
		.INIT('h0080)
	) name2735 (
		\m6_s13_cyc_o_reg/NET0131 ,
		\rf_conf13_reg[12]/NET0131 ,
		\rf_conf13_reg[13]/NET0131 ,
		\s13_msel_arb3_state_reg[0]/NET0131 ,
		_w4636_
	);
	LUT3 #(
		.INIT('h10)
	) name2736 (
		_w2943_,
		_w2950_,
		_w2951_,
		_w4637_
	);
	LUT4 #(
		.INIT('h020a)
	) name2737 (
		_w2969_,
		_w4607_,
		_w4636_,
		_w4637_,
		_w4638_
	);
	LUT2 #(
		.INIT('h4)
	) name2738 (
		_w4635_,
		_w4638_,
		_w4639_
	);
	LUT4 #(
		.INIT('hfff7)
	) name2739 (
		_w4612_,
		_w4622_,
		_w4632_,
		_w4639_,
		_w4640_
	);
	LUT2 #(
		.INIT('h4)
	) name2740 (
		_w2381_,
		_w2389_,
		_w4641_
	);
	LUT3 #(
		.INIT('h04)
	) name2741 (
		_w2377_,
		_w2379_,
		_w2380_,
		_w4642_
	);
	LUT4 #(
		.INIT('hfd00)
	) name2742 (
		\m4_s14_cyc_o_reg/NET0131 ,
		\rf_conf14_reg[8]/NET0131 ,
		\rf_conf14_reg[9]/NET0131 ,
		\s14_msel_arb0_state_reg[0]/NET0131 ,
		_w4643_
	);
	LUT3 #(
		.INIT('h10)
	) name2743 (
		_w2380_,
		_w2382_,
		_w4643_,
		_w4644_
	);
	LUT3 #(
		.INIT('hf2)
	) name2744 (
		_w2376_,
		_w2377_,
		_w2384_,
		_w4645_
	);
	LUT4 #(
		.INIT('h000d)
	) name2745 (
		_w2376_,
		_w2377_,
		_w2381_,
		_w2384_,
		_w4646_
	);
	LUT4 #(
		.INIT('h5455)
	) name2746 (
		_w4641_,
		_w4642_,
		_w4644_,
		_w4646_,
		_w4647_
	);
	LUT2 #(
		.INIT('h8)
	) name2747 (
		_w2403_,
		_w4647_,
		_w4648_
	);
	LUT2 #(
		.INIT('h8)
	) name2748 (
		\s14_msel_arb0_state_reg[1]/NET0131 ,
		\s14_msel_arb0_state_reg[2]/NET0131 ,
		_w4649_
	);
	LUT2 #(
		.INIT('h2)
	) name2749 (
		_w2384_,
		_w2389_,
		_w4650_
	);
	LUT3 #(
		.INIT('h51)
	) name2750 (
		_w2381_,
		_w2384_,
		_w2389_,
		_w4651_
	);
	LUT4 #(
		.INIT('h2232)
	) name2751 (
		_w2381_,
		_w2382_,
		_w2384_,
		_w2389_,
		_w4652_
	);
	LUT2 #(
		.INIT('h1)
	) name2752 (
		_w2377_,
		_w2389_,
		_w4653_
	);
	LUT4 #(
		.INIT('h00fd)
	) name2753 (
		\m5_s14_cyc_o_reg/NET0131 ,
		\rf_conf14_reg[10]/NET0131 ,
		\rf_conf14_reg[11]/NET0131 ,
		\s14_msel_arb0_state_reg[0]/NET0131 ,
		_w4654_
	);
	LUT3 #(
		.INIT('h01)
	) name2754 (
		_w2377_,
		_w2389_,
		_w4654_,
		_w4655_
	);
	LUT2 #(
		.INIT('h4)
	) name2755 (
		_w2376_,
		_w2380_,
		_w4656_
	);
	LUT3 #(
		.INIT('h0b)
	) name2756 (
		_w2376_,
		_w2380_,
		_w2382_,
		_w4657_
	);
	LUT4 #(
		.INIT('h0111)
	) name2757 (
		_w2379_,
		_w4652_,
		_w4655_,
		_w4657_,
		_w4658_
	);
	LUT4 #(
		.INIT('h1101)
	) name2758 (
		_w2376_,
		_w2379_,
		_w2381_,
		_w2382_,
		_w4659_
	);
	LUT4 #(
		.INIT('hfd00)
	) name2759 (
		\m2_s14_cyc_o_reg/NET0131 ,
		\rf_conf14_reg[4]/NET0131 ,
		\rf_conf14_reg[5]/NET0131 ,
		\s14_msel_arb0_state_reg[0]/NET0131 ,
		_w4660_
	);
	LUT4 #(
		.INIT('h0e0f)
	) name2760 (
		_w2380_,
		_w2382_,
		_w2384_,
		_w4660_,
		_w4661_
	);
	LUT2 #(
		.INIT('h2)
	) name2761 (
		\s14_msel_arb0_state_reg[1]/NET0131 ,
		\s14_msel_arb0_state_reg[2]/NET0131 ,
		_w4662_
	);
	LUT3 #(
		.INIT('hd0)
	) name2762 (
		_w2377_,
		_w2384_,
		_w4662_,
		_w4663_
	);
	LUT4 #(
		.INIT('h1f00)
	) name2763 (
		_w4656_,
		_w4659_,
		_w4661_,
		_w4663_,
		_w4664_
	);
	LUT3 #(
		.INIT('h0d)
	) name2764 (
		_w4649_,
		_w4658_,
		_w4664_,
		_w4665_
	);
	LUT3 #(
		.INIT('h8a)
	) name2765 (
		\s14_msel_arb0_state_reg[0]/NET0131 ,
		_w4648_,
		_w4665_,
		_w4666_
	);
	LUT3 #(
		.INIT('h02)
	) name2766 (
		\s14_msel_arb0_state_reg[0]/NET0131 ,
		_w2380_,
		_w2382_,
		_w4667_
	);
	LUT4 #(
		.INIT('h55fd)
	) name2767 (
		_w4653_,
		_w4656_,
		_w4659_,
		_w4667_,
		_w4668_
	);
	LUT3 #(
		.INIT('h8c)
	) name2768 (
		_w4650_,
		_w4662_,
		_w4668_,
		_w4669_
	);
	LUT3 #(
		.INIT('h20)
	) name2769 (
		_w2379_,
		_w2380_,
		_w4649_,
		_w4670_
	);
	LUT3 #(
		.INIT('h10)
	) name2770 (
		_w2380_,
		_w2382_,
		_w4649_,
		_w4671_
	);
	LUT4 #(
		.INIT('h020f)
	) name2771 (
		_w4651_,
		_w4655_,
		_w4670_,
		_w4671_,
		_w4672_
	);
	LUT3 #(
		.INIT('h20)
	) name2772 (
		_w2381_,
		_w2382_,
		_w2403_,
		_w4673_
	);
	LUT2 #(
		.INIT('h1)
	) name2773 (
		_w2377_,
		_w2380_,
		_w4674_
	);
	LUT4 #(
		.INIT('h00fd)
	) name2774 (
		\m7_s14_cyc_o_reg/NET0131 ,
		\rf_conf14_reg[14]/NET0131 ,
		\rf_conf14_reg[15]/NET0131 ,
		\s14_msel_arb0_state_reg[0]/NET0131 ,
		_w4675_
	);
	LUT3 #(
		.INIT('h01)
	) name2775 (
		_w2377_,
		_w2380_,
		_w4675_,
		_w4676_
	);
	LUT3 #(
		.INIT('h10)
	) name2776 (
		_w2382_,
		_w2389_,
		_w2403_,
		_w4677_
	);
	LUT4 #(
		.INIT('h0133)
	) name2777 (
		_w4645_,
		_w4673_,
		_w4676_,
		_w4677_,
		_w4678_
	);
	LUT2 #(
		.INIT('h8)
	) name2778 (
		_w4672_,
		_w4678_,
		_w4679_
	);
	LUT3 #(
		.INIT('h02)
	) name2779 (
		\s14_msel_arb0_state_reg[0]/NET0131 ,
		_w2382_,
		_w2389_,
		_w4680_
	);
	LUT3 #(
		.INIT('h80)
	) name2780 (
		_w2406_,
		_w4674_,
		_w4680_,
		_w4681_
	);
	LUT3 #(
		.INIT('h04)
	) name2781 (
		_w2382_,
		_w2384_,
		_w2389_,
		_w4682_
	);
	LUT4 #(
		.INIT('h0002)
	) name2782 (
		\m4_s14_cyc_o_reg/NET0131 ,
		\rf_conf14_reg[8]/NET0131 ,
		\rf_conf14_reg[9]/NET0131 ,
		\s14_msel_arb0_state_reg[0]/NET0131 ,
		_w4683_
	);
	LUT4 #(
		.INIT('h00b0)
	) name2783 (
		_w2376_,
		_w2380_,
		_w2406_,
		_w4683_,
		_w4684_
	);
	LUT3 #(
		.INIT('hd0)
	) name2784 (
		_w4659_,
		_w4682_,
		_w4684_,
		_w4685_
	);
	LUT2 #(
		.INIT('h1)
	) name2785 (
		_w4681_,
		_w4685_,
		_w4686_
	);
	LUT4 #(
		.INIT('hba00)
	) name2786 (
		\s14_msel_arb0_state_reg[0]/NET0131 ,
		_w4669_,
		_w4679_,
		_w4686_,
		_w4687_
	);
	LUT2 #(
		.INIT('hb)
	) name2787 (
		_w4666_,
		_w4687_,
		_w4688_
	);
	LUT2 #(
		.INIT('h2)
	) name2788 (
		_w3673_,
		_w3678_,
		_w4689_
	);
	LUT4 #(
		.INIT('h000b)
	) name2789 (
		_w3670_,
		_w3671_,
		_w3674_,
		_w3678_,
		_w4690_
	);
	LUT2 #(
		.INIT('h1)
	) name2790 (
		\s14_msel_arb1_state_reg[1]/NET0131 ,
		\s14_msel_arb1_state_reg[2]/NET0131 ,
		_w4691_
	);
	LUT4 #(
		.INIT('h0d00)
	) name2791 (
		_w3682_,
		_w3683_,
		_w3688_,
		_w4691_,
		_w4692_
	);
	LUT4 #(
		.INIT('hab00)
	) name2792 (
		_w3683_,
		_w4689_,
		_w4690_,
		_w4692_,
		_w4693_
	);
	LUT2 #(
		.INIT('h2)
	) name2793 (
		\s14_msel_arb1_state_reg[1]/NET0131 ,
		\s14_msel_arb1_state_reg[2]/NET0131 ,
		_w4694_
	);
	LUT3 #(
		.INIT('h20)
	) name2794 (
		_w3678_,
		_w3682_,
		_w4694_,
		_w4695_
	);
	LUT3 #(
		.INIT('h0b)
	) name2795 (
		_w3670_,
		_w3671_,
		_w3674_,
		_w4696_
	);
	LUT2 #(
		.INIT('h1)
	) name2796 (
		_w3670_,
		_w3688_,
		_w4697_
	);
	LUT4 #(
		.INIT('h00f7)
	) name2797 (
		\m1_s14_cyc_o_reg/NET0131 ,
		\rf_conf14_reg[2]/NET0131 ,
		\rf_conf14_reg[3]/NET0131 ,
		\s14_msel_arb1_state_reg[0]/NET0131 ,
		_w4698_
	);
	LUT3 #(
		.INIT('h01)
	) name2798 (
		_w3670_,
		_w3688_,
		_w4698_,
		_w4699_
	);
	LUT3 #(
		.INIT('h10)
	) name2799 (
		_w3673_,
		_w3682_,
		_w4694_,
		_w4700_
	);
	LUT4 #(
		.INIT('h0455)
	) name2800 (
		_w4695_,
		_w4696_,
		_w4699_,
		_w4700_,
		_w4701_
	);
	LUT2 #(
		.INIT('h4)
	) name2801 (
		_w3673_,
		_w3676_,
		_w4702_
	);
	LUT3 #(
		.INIT('h0d)
	) name2802 (
		_w3678_,
		_w3682_,
		_w3683_,
		_w4703_
	);
	LUT4 #(
		.INIT('haf2f)
	) name2803 (
		_w4696_,
		_w4697_,
		_w4702_,
		_w4703_,
		_w4704_
	);
	LUT4 #(
		.INIT('h4555)
	) name2804 (
		\s14_msel_arb1_state_reg[0]/NET0131 ,
		_w4693_,
		_w4701_,
		_w4704_,
		_w4705_
	);
	LUT4 #(
		.INIT('hf700)
	) name2805 (
		\m0_s14_cyc_o_reg/NET0131 ,
		\rf_conf14_reg[0]/NET0131 ,
		\rf_conf14_reg[1]/NET0131 ,
		\s14_msel_arb1_state_reg[0]/NET0131 ,
		_w4706_
	);
	LUT3 #(
		.INIT('h01)
	) name2806 (
		_w3670_,
		_w3673_,
		_w3682_,
		_w4707_
	);
	LUT4 #(
		.INIT('h0100)
	) name2807 (
		_w3670_,
		_w3673_,
		_w3682_,
		_w4706_,
		_w4708_
	);
	LUT4 #(
		.INIT('h0008)
	) name2808 (
		\m6_s14_cyc_o_reg/NET0131 ,
		\rf_conf14_reg[12]/NET0131 ,
		\rf_conf14_reg[13]/NET0131 ,
		\s14_msel_arb1_state_reg[0]/NET0131 ,
		_w4709_
	);
	LUT2 #(
		.INIT('h2)
	) name2809 (
		_w3671_,
		_w4709_,
		_w4710_
	);
	LUT3 #(
		.INIT('h04)
	) name2810 (
		_w3673_,
		_w3674_,
		_w3682_,
		_w4711_
	);
	LUT2 #(
		.INIT('h1)
	) name2811 (
		_w3688_,
		_w4709_,
		_w4712_
	);
	LUT4 #(
		.INIT('h0233)
	) name2812 (
		_w4703_,
		_w4710_,
		_w4711_,
		_w4712_,
		_w4713_
	);
	LUT2 #(
		.INIT('h8)
	) name2813 (
		\s14_msel_arb1_state_reg[1]/NET0131 ,
		\s14_msel_arb1_state_reg[2]/NET0131 ,
		_w4714_
	);
	LUT3 #(
		.INIT('hb0)
	) name2814 (
		_w4708_,
		_w4713_,
		_w4714_,
		_w4715_
	);
	LUT3 #(
		.INIT('h20)
	) name2815 (
		\s14_msel_arb1_state_reg[0]/NET0131 ,
		\s14_msel_arb1_state_reg[1]/NET0131 ,
		\s14_msel_arb1_state_reg[2]/NET0131 ,
		_w4716_
	);
	LUT4 #(
		.INIT('h00a2)
	) name2816 (
		_w4696_,
		_w4697_,
		_w4703_,
		_w4708_,
		_w4717_
	);
	LUT2 #(
		.INIT('h2)
	) name2817 (
		_w4716_,
		_w4717_,
		_w4718_
	);
	LUT2 #(
		.INIT('h1)
	) name2818 (
		_w3671_,
		_w4706_,
		_w4719_
	);
	LUT4 #(
		.INIT('h0a02)
	) name2819 (
		_w4703_,
		_w4707_,
		_w4711_,
		_w4719_,
		_w4720_
	);
	LUT3 #(
		.INIT('h02)
	) name2820 (
		\s14_msel_arb1_state_reg[0]/NET0131 ,
		\s14_msel_arb1_state_reg[1]/NET0131 ,
		\s14_msel_arb1_state_reg[2]/NET0131 ,
		_w4721_
	);
	LUT3 #(
		.INIT('h51)
	) name2821 (
		_w3673_,
		_w3682_,
		_w3683_,
		_w4722_
	);
	LUT4 #(
		.INIT('h0eee)
	) name2822 (
		_w4689_,
		_w4690_,
		_w4699_,
		_w4722_,
		_w4723_
	);
	LUT3 #(
		.INIT('h08)
	) name2823 (
		\s14_msel_arb1_state_reg[0]/NET0131 ,
		\s14_msel_arb1_state_reg[1]/NET0131 ,
		\s14_msel_arb1_state_reg[2]/NET0131 ,
		_w4724_
	);
	LUT4 #(
		.INIT('hb0bb)
	) name2824 (
		_w4720_,
		_w4721_,
		_w4723_,
		_w4724_,
		_w4725_
	);
	LUT4 #(
		.INIT('hfeff)
	) name2825 (
		_w4705_,
		_w4715_,
		_w4718_,
		_w4725_,
		_w4726_
	);
	LUT2 #(
		.INIT('h2)
	) name2826 (
		\s14_msel_arb2_state_reg[1]/NET0131 ,
		\s14_msel_arb2_state_reg[2]/NET0131 ,
		_w4727_
	);
	LUT2 #(
		.INIT('h4)
	) name2827 (
		_w2991_,
		_w4727_,
		_w4728_
	);
	LUT2 #(
		.INIT('h1)
	) name2828 (
		_w2973_,
		_w2980_,
		_w4729_
	);
	LUT3 #(
		.INIT('hae)
	) name2829 (
		_w2973_,
		_w2980_,
		_w2981_,
		_w4730_
	);
	LUT2 #(
		.INIT('h1)
	) name2830 (
		_w2985_,
		_w2996_,
		_w4731_
	);
	LUT2 #(
		.INIT('h1)
	) name2831 (
		_w2981_,
		_w2986_,
		_w4732_
	);
	LUT4 #(
		.INIT('h7577)
	) name2832 (
		_w4728_,
		_w4730_,
		_w4731_,
		_w4732_,
		_w4733_
	);
	LUT3 #(
		.INIT('h0d)
	) name2833 (
		_w2983_,
		_w2984_,
		_w2985_,
		_w4734_
	);
	LUT4 #(
		.INIT('h00f2)
	) name2834 (
		_w2983_,
		_w2984_,
		_w2985_,
		_w2986_,
		_w4735_
	);
	LUT3 #(
		.INIT('h10)
	) name2835 (
		\s14_msel_arb2_state_reg[0]/NET0131 ,
		\s14_msel_arb2_state_reg[1]/NET0131 ,
		\s14_msel_arb2_state_reg[2]/NET0131 ,
		_w4736_
	);
	LUT4 #(
		.INIT('h2300)
	) name2836 (
		_w2973_,
		_w2974_,
		_w2981_,
		_w4736_,
		_w4737_
	);
	LUT3 #(
		.INIT('hd0)
	) name2837 (
		_w4729_,
		_w4735_,
		_w4737_,
		_w4738_
	);
	LUT3 #(
		.INIT('h0e)
	) name2838 (
		_w2974_,
		_w4733_,
		_w4738_,
		_w4739_
	);
	LUT2 #(
		.INIT('h1)
	) name2839 (
		\s14_msel_arb2_state_reg[1]/NET0131 ,
		\s14_msel_arb2_state_reg[2]/NET0131 ,
		_w4740_
	);
	LUT4 #(
		.INIT('h0020)
	) name2840 (
		\m0_s14_cyc_o_reg/NET0131 ,
		\rf_conf14_reg[0]/NET0131 ,
		\rf_conf14_reg[1]/NET0131 ,
		\s14_msel_arb2_state_reg[0]/NET0131 ,
		_w4741_
	);
	LUT2 #(
		.INIT('h2)
	) name2841 (
		_w4740_,
		_w4741_,
		_w4742_
	);
	LUT2 #(
		.INIT('h1)
	) name2842 (
		_w2974_,
		_w2984_,
		_w4743_
	);
	LUT4 #(
		.INIT('h4fcf)
	) name2843 (
		_w4730_,
		_w4734_,
		_w4742_,
		_w4743_,
		_w4744_
	);
	LUT3 #(
		.INIT('h20)
	) name2844 (
		_w2983_,
		_w2991_,
		_w4727_,
		_w4745_
	);
	LUT3 #(
		.INIT('h20)
	) name2845 (
		\s14_msel_arb2_state_reg[0]/NET0131 ,
		\s14_msel_arb2_state_reg[1]/NET0131 ,
		\s14_msel_arb2_state_reg[2]/NET0131 ,
		_w4746_
	);
	LUT2 #(
		.INIT('h8)
	) name2846 (
		_w2973_,
		_w4746_,
		_w4747_
	);
	LUT2 #(
		.INIT('h1)
	) name2847 (
		_w4745_,
		_w4747_,
		_w4748_
	);
	LUT2 #(
		.INIT('h8)
	) name2848 (
		_w4744_,
		_w4748_,
		_w4749_
	);
	LUT3 #(
		.INIT('h02)
	) name2849 (
		\s14_msel_arb2_state_reg[0]/NET0131 ,
		\s14_msel_arb2_state_reg[1]/NET0131 ,
		\s14_msel_arb2_state_reg[2]/NET0131 ,
		_w4750_
	);
	LUT4 #(
		.INIT('h0100)
	) name2850 (
		_w2974_,
		_w2984_,
		_w2986_,
		_w4750_,
		_w4751_
	);
	LUT2 #(
		.INIT('h4)
	) name2851 (
		_w2973_,
		_w4746_,
		_w4752_
	);
	LUT2 #(
		.INIT('h1)
	) name2852 (
		_w4751_,
		_w4752_,
		_w4753_
	);
	LUT2 #(
		.INIT('h4)
	) name2853 (
		_w2980_,
		_w2986_,
		_w4754_
	);
	LUT4 #(
		.INIT('h0051)
	) name2854 (
		_w2980_,
		_w2983_,
		_w2984_,
		_w2985_,
		_w4755_
	);
	LUT4 #(
		.INIT('hdf00)
	) name2855 (
		\m0_s14_cyc_o_reg/NET0131 ,
		\rf_conf14_reg[0]/NET0131 ,
		\rf_conf14_reg[1]/NET0131 ,
		\s14_msel_arb2_state_reg[0]/NET0131 ,
		_w4756_
	);
	LUT3 #(
		.INIT('h10)
	) name2856 (
		_w2974_,
		_w2984_,
		_w4756_,
		_w4757_
	);
	LUT4 #(
		.INIT('h0054)
	) name2857 (
		_w4751_,
		_w4754_,
		_w4755_,
		_w4757_,
		_w4758_
	);
	LUT3 #(
		.INIT('h01)
	) name2858 (
		_w2981_,
		_w4753_,
		_w4758_,
		_w4759_
	);
	LUT4 #(
		.INIT('h00df)
	) name2859 (
		\m5_s14_cyc_o_reg/NET0131 ,
		\rf_conf14_reg[10]/NET0131 ,
		\rf_conf14_reg[11]/NET0131 ,
		\s14_msel_arb2_state_reg[0]/NET0131 ,
		_w4760_
	);
	LUT4 #(
		.INIT('h0001)
	) name2860 (
		_w2974_,
		_w2984_,
		_w2986_,
		_w4760_,
		_w4761_
	);
	LUT3 #(
		.INIT('h0e)
	) name2861 (
		_w4754_,
		_w4755_,
		_w4761_,
		_w4762_
	);
	LUT4 #(
		.INIT('h0020)
	) name2862 (
		\m6_s14_cyc_o_reg/NET0131 ,
		\rf_conf14_reg[12]/NET0131 ,
		\rf_conf14_reg[13]/NET0131 ,
		\s14_msel_arb2_state_reg[0]/NET0131 ,
		_w4763_
	);
	LUT3 #(
		.INIT('h10)
	) name2863 (
		_w2973_,
		_w2980_,
		_w2981_,
		_w4764_
	);
	LUT4 #(
		.INIT('h020a)
	) name2864 (
		_w2999_,
		_w4734_,
		_w4763_,
		_w4764_,
		_w4765_
	);
	LUT2 #(
		.INIT('h4)
	) name2865 (
		_w4762_,
		_w4765_,
		_w4766_
	);
	LUT4 #(
		.INIT('hfff7)
	) name2866 (
		_w4739_,
		_w4749_,
		_w4759_,
		_w4766_,
		_w4767_
	);
	LUT3 #(
		.INIT('hdc)
	) name2867 (
		_w3270_,
		_w3271_,
		_w3281_,
		_w4768_
	);
	LUT2 #(
		.INIT('h4)
	) name2868 (
		_w3273_,
		_w3275_,
		_w4769_
	);
	LUT4 #(
		.INIT('h000d)
	) name2869 (
		_w3268_,
		_w3269_,
		_w3273_,
		_w3274_,
		_w4770_
	);
	LUT4 #(
		.INIT('h7f00)
	) name2870 (
		\m6_s14_cyc_o_reg/NET0131 ,
		\rf_conf14_reg[12]/NET0131 ,
		\rf_conf14_reg[13]/NET0131 ,
		\s14_msel_arb3_state_reg[0]/NET0131 ,
		_w4771_
	);
	LUT4 #(
		.INIT('ha2f3)
	) name2871 (
		_w3269_,
		_w3270_,
		_w3271_,
		_w4771_,
		_w4772_
	);
	LUT4 #(
		.INIT('h0155)
	) name2872 (
		_w4768_,
		_w4769_,
		_w4770_,
		_w4772_,
		_w4773_
	);
	LUT2 #(
		.INIT('h8)
	) name2873 (
		_w3293_,
		_w4773_,
		_w4774_
	);
	LUT2 #(
		.INIT('h1)
	) name2874 (
		\s14_msel_arb3_state_reg[1]/NET0131 ,
		\s14_msel_arb3_state_reg[2]/NET0131 ,
		_w4775_
	);
	LUT3 #(
		.INIT('h20)
	) name2875 (
		_w3268_,
		_w3269_,
		_w4775_,
		_w4776_
	);
	LUT2 #(
		.INIT('h4)
	) name2876 (
		_w3270_,
		_w3281_,
		_w4777_
	);
	LUT4 #(
		.INIT('h1101)
	) name2877 (
		_w3270_,
		_w3273_,
		_w3274_,
		_w3275_,
		_w4778_
	);
	LUT3 #(
		.INIT('h10)
	) name2878 (
		_w3269_,
		_w3271_,
		_w4775_,
		_w4779_
	);
	LUT4 #(
		.INIT('h5455)
	) name2879 (
		_w4776_,
		_w4777_,
		_w4778_,
		_w4779_,
		_w4780_
	);
	LUT3 #(
		.INIT('h08)
	) name2880 (
		_w3267_,
		_w3273_,
		_w3281_,
		_w4781_
	);
	LUT3 #(
		.INIT('h0d)
	) name2881 (
		_w3268_,
		_w3269_,
		_w3274_,
		_w4782_
	);
	LUT3 #(
		.INIT('h04)
	) name2882 (
		_w3269_,
		_w3270_,
		_w3271_,
		_w4783_
	);
	LUT3 #(
		.INIT('h02)
	) name2883 (
		_w3267_,
		_w3275_,
		_w3281_,
		_w4784_
	);
	LUT4 #(
		.INIT('h0455)
	) name2884 (
		_w4781_,
		_w4782_,
		_w4783_,
		_w4784_,
		_w4785_
	);
	LUT3 #(
		.INIT('h40)
	) name2885 (
		\s14_msel_arb3_state_reg[0]/NET0131 ,
		_w4780_,
		_w4785_,
		_w4786_
	);
	LUT3 #(
		.INIT('h51)
	) name2886 (
		_w3275_,
		_w4782_,
		_w4783_,
		_w4787_
	);
	LUT4 #(
		.INIT('h0001)
	) name2887 (
		_w3269_,
		_w3271_,
		_w3275_,
		_w3281_,
		_w4788_
	);
	LUT2 #(
		.INIT('h1)
	) name2888 (
		_w3273_,
		_w4788_,
		_w4789_
	);
	LUT3 #(
		.INIT('h2a)
	) name2889 (
		\s14_msel_arb3_state_reg[0]/NET0131 ,
		_w3270_,
		_w3293_,
		_w4790_
	);
	LUT4 #(
		.INIT('h7500)
	) name2890 (
		_w3267_,
		_w4787_,
		_w4789_,
		_w4790_,
		_w4791_
	);
	LUT3 #(
		.INIT('h0b)
	) name2891 (
		_w4774_,
		_w4786_,
		_w4791_,
		_w4792_
	);
	LUT2 #(
		.INIT('h4)
	) name2892 (
		_w3268_,
		_w3271_,
		_w4793_
	);
	LUT4 #(
		.INIT('h5455)
	) name2893 (
		_w3268_,
		_w3269_,
		_w3281_,
		_w4771_,
		_w4794_
	);
	LUT4 #(
		.INIT('h010f)
	) name2894 (
		_w4777_,
		_w4778_,
		_w4793_,
		_w4794_,
		_w4795_
	);
	LUT3 #(
		.INIT('h02)
	) name2895 (
		\s14_msel_arb3_state_reg[0]/NET0131 ,
		\s14_msel_arb3_state_reg[1]/NET0131 ,
		\s14_msel_arb3_state_reg[2]/NET0131 ,
		_w4796_
	);
	LUT2 #(
		.INIT('h8)
	) name2896 (
		_w4795_,
		_w4796_,
		_w4797_
	);
	LUT2 #(
		.INIT('h1)
	) name2897 (
		_w3273_,
		_w4771_,
		_w4798_
	);
	LUT3 #(
		.INIT('h01)
	) name2898 (
		_w3269_,
		_w3271_,
		_w3281_,
		_w4799_
	);
	LUT4 #(
		.INIT('h2022)
	) name2899 (
		_w4782_,
		_w4783_,
		_w4798_,
		_w4799_,
		_w4800_
	);
	LUT4 #(
		.INIT('h0080)
	) name2900 (
		\m6_s14_cyc_o_reg/NET0131 ,
		\rf_conf14_reg[12]/NET0131 ,
		\rf_conf14_reg[13]/NET0131 ,
		\s14_msel_arb3_state_reg[0]/NET0131 ,
		_w4801_
	);
	LUT2 #(
		.INIT('h2)
	) name2901 (
		_w3279_,
		_w4801_,
		_w4802_
	);
	LUT3 #(
		.INIT('h10)
	) name2902 (
		_w3269_,
		_w3271_,
		_w4771_,
		_w4803_
	);
	LUT3 #(
		.INIT('h08)
	) name2903 (
		\s14_msel_arb3_state_reg[0]/NET0131 ,
		\s14_msel_arb3_state_reg[1]/NET0131 ,
		\s14_msel_arb3_state_reg[2]/NET0131 ,
		_w4804_
	);
	LUT3 #(
		.INIT('h10)
	) name2904 (
		_w3270_,
		_w3281_,
		_w4804_,
		_w4805_
	);
	LUT4 #(
		.INIT('hf100)
	) name2905 (
		_w4769_,
		_w4770_,
		_w4803_,
		_w4805_,
		_w4806_
	);
	LUT3 #(
		.INIT('h0b)
	) name2906 (
		_w4800_,
		_w4802_,
		_w4806_,
		_w4807_
	);
	LUT2 #(
		.INIT('h4)
	) name2907 (
		_w4797_,
		_w4807_,
		_w4808_
	);
	LUT2 #(
		.INIT('hb)
	) name2908 (
		_w4792_,
		_w4808_,
		_w4809_
	);
	LUT3 #(
		.INIT('hf4)
	) name2909 (
		_w2880_,
		_w2881_,
		_w2885_,
		_w4810_
	);
	LUT4 #(
		.INIT('h000b)
	) name2910 (
		_w2880_,
		_w2881_,
		_w2885_,
		_w2886_,
		_w4811_
	);
	LUT2 #(
		.INIT('h1)
	) name2911 (
		_w2879_,
		_w2880_,
		_w4812_
	);
	LUT4 #(
		.INIT('hf700)
	) name2912 (
		\m4_s15_cyc_o_reg/NET0131 ,
		\rf_conf15_reg[8]/NET0131 ,
		\rf_conf15_reg[9]/NET0131 ,
		\s15_msel_arb1_state_reg[0]/NET0131 ,
		_w4813_
	);
	LUT4 #(
		.INIT('h0302)
	) name2913 (
		_w2878_,
		_w2879_,
		_w2880_,
		_w4813_,
		_w4814_
	);
	LUT4 #(
		.INIT('h00a2)
	) name2914 (
		\s15_msel_arb1_state_reg[2]/NET0131 ,
		_w2884_,
		_w2886_,
		_w2937_,
		_w4815_
	);
	LUT4 #(
		.INIT('h5100)
	) name2915 (
		\s15_msel_arb1_state_reg[1]/NET0131 ,
		_w4811_,
		_w4814_,
		_w4815_,
		_w4816_
	);
	LUT4 #(
		.INIT('h0008)
	) name2916 (
		\m1_s15_cyc_o_reg/NET0131 ,
		\rf_conf15_reg[2]/NET0131 ,
		\rf_conf15_reg[3]/NET0131 ,
		\s15_msel_arb1_state_reg[2]/NET0131 ,
		_w4817_
	);
	LUT3 #(
		.INIT('h51)
	) name2917 (
		_w2878_,
		_w2886_,
		_w2887_,
		_w4818_
	);
	LUT4 #(
		.INIT('h00f7)
	) name2918 (
		\m7_s15_cyc_o_reg/NET0131 ,
		\rf_conf15_reg[14]/NET0131 ,
		\rf_conf15_reg[15]/NET0131 ,
		\s15_msel_arb1_state_reg[0]/NET0131 ,
		_w4819_
	);
	LUT3 #(
		.INIT('h01)
	) name2919 (
		_w2884_,
		_w2887_,
		_w4819_,
		_w4820_
	);
	LUT4 #(
		.INIT('h00f7)
	) name2920 (
		\m2_s15_cyc_o_reg/NET0131 ,
		\rf_conf15_reg[4]/NET0131 ,
		\rf_conf15_reg[5]/NET0131 ,
		\s15_msel_arb1_state_reg[2]/NET0131 ,
		_w4821_
	);
	LUT4 #(
		.INIT('h0455)
	) name2921 (
		_w4817_,
		_w4818_,
		_w4820_,
		_w4821_,
		_w4822_
	);
	LUT4 #(
		.INIT('h0008)
	) name2922 (
		\m0_s15_cyc_o_reg/NET0131 ,
		\rf_conf15_reg[0]/NET0131 ,
		\rf_conf15_reg[1]/NET0131 ,
		\s15_msel_arb1_state_reg[0]/NET0131 ,
		_w4823_
	);
	LUT3 #(
		.INIT('h02)
	) name2923 (
		_w2880_,
		_w2881_,
		_w2885_,
		_w4824_
	);
	LUT4 #(
		.INIT('h0105)
	) name2924 (
		\s15_msel_arb1_state_reg[1]/NET0131 ,
		_w4818_,
		_w4823_,
		_w4824_,
		_w4825_
	);
	LUT3 #(
		.INIT('h45)
	) name2925 (
		_w4816_,
		_w4822_,
		_w4825_,
		_w4826_
	);
	LUT4 #(
		.INIT('h5504)
	) name2926 (
		_w2878_,
		_w2884_,
		_w2886_,
		_w2887_,
		_w4827_
	);
	LUT2 #(
		.INIT('h1)
	) name2927 (
		_w2878_,
		_w2886_,
		_w4828_
	);
	LUT4 #(
		.INIT('h0008)
	) name2928 (
		\m2_s15_cyc_o_reg/NET0131 ,
		\rf_conf15_reg[4]/NET0131 ,
		\rf_conf15_reg[5]/NET0131 ,
		\s15_msel_arb1_state_reg[0]/NET0131 ,
		_w4829_
	);
	LUT2 #(
		.INIT('h1)
	) name2929 (
		\s15_msel_arb1_state_reg[2]/NET0131 ,
		_w4829_,
		_w4830_
	);
	LUT4 #(
		.INIT('h2300)
	) name2930 (
		_w4810_,
		_w4827_,
		_w4828_,
		_w4830_,
		_w4831_
	);
	LUT4 #(
		.INIT('h0008)
	) name2931 (
		\m6_s15_cyc_o_reg/NET0131 ,
		\rf_conf15_reg[12]/NET0131 ,
		\rf_conf15_reg[13]/NET0131 ,
		\s15_msel_arb1_state_reg[0]/NET0131 ,
		_w4832_
	);
	LUT2 #(
		.INIT('h2)
	) name2932 (
		\s15_msel_arb1_state_reg[2]/NET0131 ,
		_w4832_,
		_w4833_
	);
	LUT4 #(
		.INIT('h51ff)
	) name2933 (
		_w4810_,
		_w4812_,
		_w4818_,
		_w4833_,
		_w4834_
	);
	LUT4 #(
		.INIT('h0100)
	) name2934 (
		_w2879_,
		_w2880_,
		_w2884_,
		_w4813_,
		_w4835_
	);
	LUT4 #(
		.INIT('haa8a)
	) name2935 (
		\s15_msel_arb1_state_reg[1]/NET0131 ,
		_w4831_,
		_w4834_,
		_w4835_,
		_w4836_
	);
	LUT2 #(
		.INIT('hd)
	) name2936 (
		_w4826_,
		_w4836_,
		_w4837_
	);
	LUT3 #(
		.INIT('h0b)
	) name2937 (
		_w2894_,
		_w2895_,
		_w2900_,
		_w4838_
	);
	LUT4 #(
		.INIT('haa20)
	) name2938 (
		\s15_msel_arb2_state_reg[2]/NET0131 ,
		_w2894_,
		_w2895_,
		_w2900_,
		_w4839_
	);
	LUT3 #(
		.INIT('h45)
	) name2939 (
		_w2891_,
		_w2898_,
		_w2899_,
		_w4840_
	);
	LUT3 #(
		.INIT('h02)
	) name2940 (
		\s15_msel_arb2_state_reg[2]/NET0131 ,
		_w2892_,
		_w2894_,
		_w4841_
	);
	LUT3 #(
		.INIT('h45)
	) name2941 (
		_w4839_,
		_w4840_,
		_w4841_,
		_w4842_
	);
	LUT4 #(
		.INIT('h4544)
	) name2942 (
		_w2901_,
		_w4839_,
		_w4840_,
		_w4841_,
		_w4843_
	);
	LUT4 #(
		.INIT('h4544)
	) name2943 (
		\s15_msel_arb2_state_reg[2]/NET0131 ,
		_w2891_,
		_w2898_,
		_w2899_,
		_w4844_
	);
	LUT3 #(
		.INIT('h01)
	) name2944 (
		\s15_msel_arb2_state_reg[2]/NET0131 ,
		_w2898_,
		_w2901_,
		_w4845_
	);
	LUT3 #(
		.INIT('h23)
	) name2945 (
		_w4838_,
		_w4844_,
		_w4845_,
		_w4846_
	);
	LUT4 #(
		.INIT('h5150)
	) name2946 (
		_w2892_,
		_w4838_,
		_w4844_,
		_w4845_,
		_w4847_
	);
	LUT3 #(
		.INIT('h01)
	) name2947 (
		\s15_msel_arb2_state_reg[0]/NET0131 ,
		_w4843_,
		_w4847_,
		_w4848_
	);
	LUT4 #(
		.INIT('h0001)
	) name2948 (
		_w2892_,
		_w2894_,
		_w2898_,
		_w2901_,
		_w4849_
	);
	LUT2 #(
		.INIT('h2)
	) name2949 (
		\s15_msel_arb2_state_reg[0]/NET0131 ,
		_w4849_,
		_w4850_
	);
	LUT4 #(
		.INIT('h2aaa)
	) name2950 (
		\s15_msel_arb2_state_reg[1]/NET0131 ,
		_w4842_,
		_w4846_,
		_w4850_,
		_w4851_
	);
	LUT2 #(
		.INIT('h4)
	) name2951 (
		_w4848_,
		_w4851_,
		_w4852_
	);
	LUT3 #(
		.INIT('h04)
	) name2952 (
		_w2898_,
		_w2900_,
		_w2901_,
		_w4853_
	);
	LUT3 #(
		.INIT('h02)
	) name2953 (
		\s15_msel_arb2_state_reg[0]/NET0131 ,
		_w2898_,
		_w2901_,
		_w4854_
	);
	LUT3 #(
		.INIT('h02)
	) name2954 (
		_w4840_,
		_w4853_,
		_w4854_,
		_w4855_
	);
	LUT4 #(
		.INIT('h4044)
	) name2955 (
		_w2891_,
		_w2894_,
		_w2898_,
		_w2899_,
		_w4856_
	);
	LUT3 #(
		.INIT('h01)
	) name2956 (
		\s15_msel_arb2_state_reg[2]/NET0131 ,
		_w2892_,
		_w2895_,
		_w4857_
	);
	LUT3 #(
		.INIT('hb0)
	) name2957 (
		_w4853_,
		_w4856_,
		_w4857_,
		_w4858_
	);
	LUT4 #(
		.INIT('h00df)
	) name2958 (
		\m1_s15_cyc_o_reg/NET0131 ,
		\rf_conf15_reg[2]/NET0131 ,
		\rf_conf15_reg[3]/NET0131 ,
		\s15_msel_arb2_state_reg[2]/NET0131 ,
		_w4859_
	);
	LUT4 #(
		.INIT('hdf00)
	) name2959 (
		\m5_s15_cyc_o_reg/NET0131 ,
		\rf_conf15_reg[10]/NET0131 ,
		\rf_conf15_reg[11]/NET0131 ,
		\s15_msel_arb2_state_reg[2]/NET0131 ,
		_w4860_
	);
	LUT2 #(
		.INIT('h1)
	) name2960 (
		_w4859_,
		_w4860_,
		_w4861_
	);
	LUT4 #(
		.INIT('h1b11)
	) name2961 (
		\s15_msel_arb2_state_reg[2]/NET0131 ,
		_w2895_,
		_w2899_,
		_w2901_,
		_w4862_
	);
	LUT3 #(
		.INIT('h02)
	) name2962 (
		_w2891_,
		_w2892_,
		_w2894_,
		_w4863_
	);
	LUT4 #(
		.INIT('hdf00)
	) name2963 (
		\m4_s15_cyc_o_reg/NET0131 ,
		\rf_conf15_reg[8]/NET0131 ,
		\rf_conf15_reg[9]/NET0131 ,
		\s15_msel_arb2_state_reg[0]/NET0131 ,
		_w4864_
	);
	LUT3 #(
		.INIT('h10)
	) name2964 (
		_w2892_,
		_w2894_,
		_w4864_,
		_w4865_
	);
	LUT4 #(
		.INIT('h0002)
	) name2965 (
		_w4838_,
		_w4861_,
		_w4863_,
		_w4865_,
		_w4866_
	);
	LUT4 #(
		.INIT('hbbb0)
	) name2966 (
		_w4855_,
		_w4858_,
		_w4862_,
		_w4866_,
		_w4867_
	);
	LUT2 #(
		.INIT('h2)
	) name2967 (
		\s15_msel_arb2_state_reg[0]/NET0131 ,
		\s15_msel_arb2_state_reg[1]/NET0131 ,
		_w4868_
	);
	LUT2 #(
		.INIT('h1)
	) name2968 (
		\s15_msel_arb2_state_reg[0]/NET0131 ,
		\s15_msel_arb2_state_reg[1]/NET0131 ,
		_w4869_
	);
	LUT3 #(
		.INIT('h10)
	) name2969 (
		\s15_msel_arb2_state_reg[0]/NET0131 ,
		\s15_msel_arb2_state_reg[1]/NET0131 ,
		\s15_msel_arb2_state_reg[2]/NET0131 ,
		_w4870_
	);
	LUT4 #(
		.INIT('h0020)
	) name2970 (
		\m4_s15_cyc_o_reg/NET0131 ,
		\rf_conf15_reg[8]/NET0131 ,
		\rf_conf15_reg[9]/NET0131 ,
		\s15_msel_arb2_state_reg[0]/NET0131 ,
		_w4871_
	);
	LUT3 #(
		.INIT('h0e)
	) name2971 (
		_w2898_,
		_w2899_,
		_w4871_,
		_w4872_
	);
	LUT4 #(
		.INIT('hfa10)
	) name2972 (
		_w2898_,
		_w2899_,
		_w2901_,
		_w4871_,
		_w4873_
	);
	LUT3 #(
		.INIT('h02)
	) name2973 (
		\s15_msel_arb2_state_reg[0]/NET0131 ,
		_w2892_,
		_w2894_,
		_w4874_
	);
	LUT4 #(
		.INIT('h0002)
	) name2974 (
		_w4838_,
		_w4863_,
		_w4872_,
		_w4874_,
		_w4875_
	);
	LUT3 #(
		.INIT('h02)
	) name2975 (
		_w4870_,
		_w4873_,
		_w4875_,
		_w4876_
	);
	LUT4 #(
		.INIT('h0020)
	) name2976 (
		\m0_s15_cyc_o_reg/NET0131 ,
		\rf_conf15_reg[0]/NET0131 ,
		\rf_conf15_reg[1]/NET0131 ,
		\s15_msel_arb2_state_reg[0]/NET0131 ,
		_w4877_
	);
	LUT3 #(
		.INIT('h0e)
	) name2977 (
		_w2894_,
		_w2895_,
		_w4877_,
		_w4878_
	);
	LUT4 #(
		.INIT('hee02)
	) name2978 (
		_w2892_,
		_w2894_,
		_w2895_,
		_w4877_,
		_w4879_
	);
	LUT4 #(
		.INIT('h0002)
	) name2979 (
		_w4840_,
		_w4853_,
		_w4854_,
		_w4878_,
		_w4880_
	);
	LUT3 #(
		.INIT('h01)
	) name2980 (
		\s15_msel_arb2_state_reg[0]/NET0131 ,
		\s15_msel_arb2_state_reg[1]/NET0131 ,
		\s15_msel_arb2_state_reg[2]/NET0131 ,
		_w4881_
	);
	LUT3 #(
		.INIT('h10)
	) name2981 (
		_w4879_,
		_w4880_,
		_w4881_,
		_w4882_
	);
	LUT4 #(
		.INIT('h000b)
	) name2982 (
		_w4867_,
		_w4868_,
		_w4876_,
		_w4882_,
		_w4883_
	);
	LUT2 #(
		.INIT('hb)
	) name2983 (
		_w4852_,
		_w4883_,
		_w4884_
	);
	LUT4 #(
		.INIT('h0020)
	) name2984 (
		\m6_s15_cyc_o_reg/NET0131 ,
		\rf_conf15_reg[12]/NET0131 ,
		\rf_conf15_reg[13]/NET0131 ,
		\s15_msel_arb2_state_reg[0]/NET0131 ,
		_w4885_
	);
	LUT3 #(
		.INIT('h32)
	) name2985 (
		_w2900_,
		_w4869_,
		_w4885_,
		_w4886_
	);
	LUT3 #(
		.INIT('he0)
	) name2986 (
		_w2899_,
		_w2901_,
		_w4868_,
		_w4887_
	);
	LUT4 #(
		.INIT('haaa8)
	) name2987 (
		\s15_msel_arb2_state_reg[2]/NET0131 ,
		_w2897_,
		_w4886_,
		_w4887_,
		_w4888_
	);
	LUT4 #(
		.INIT('h00df)
	) name2988 (
		\m3_s15_cyc_o_reg/NET0131 ,
		\rf_conf15_reg[6]/NET0131 ,
		\rf_conf15_reg[7]/NET0131 ,
		\s15_msel_arb2_state_reg[2]/NET0131 ,
		_w4889_
	);
	LUT2 #(
		.INIT('h1)
	) name2989 (
		_w4870_,
		_w4889_,
		_w4890_
	);
	LUT3 #(
		.INIT('h01)
	) name2990 (
		_w2892_,
		_w2895_,
		_w4877_,
		_w4891_
	);
	LUT4 #(
		.INIT('h0020)
	) name2991 (
		\m2_s15_cyc_o_reg/NET0131 ,
		\rf_conf15_reg[4]/NET0131 ,
		\rf_conf15_reg[5]/NET0131 ,
		\s15_msel_arb2_state_reg[0]/NET0131 ,
		_w4892_
	);
	LUT3 #(
		.INIT('h31)
	) name2992 (
		\s15_msel_arb2_state_reg[1]/NET0131 ,
		_w4870_,
		_w4892_,
		_w4893_
	);
	LUT4 #(
		.INIT('h1011)
	) name2993 (
		_w2903_,
		_w4890_,
		_w4891_,
		_w4893_,
		_w4894_
	);
	LUT2 #(
		.INIT('he)
	) name2994 (
		_w4888_,
		_w4894_,
		_w4895_
	);
	LUT2 #(
		.INIT('h2)
	) name2995 (
		_w2908_,
		_w2912_,
		_w4896_
	);
	LUT4 #(
		.INIT('h000d)
	) name2996 (
		_w2905_,
		_w2906_,
		_w2909_,
		_w2912_,
		_w4897_
	);
	LUT2 #(
		.INIT('h1)
	) name2997 (
		_w4896_,
		_w4897_,
		_w4898_
	);
	LUT3 #(
		.INIT('ha2)
	) name2998 (
		\s15_msel_arb3_state_reg[2]/NET0131 ,
		_w2913_,
		_w2915_,
		_w4899_
	);
	LUT4 #(
		.INIT('h0a02)
	) name2999 (
		\s15_msel_arb3_state_reg[2]/NET0131 ,
		_w2913_,
		_w2914_,
		_w2915_,
		_w4900_
	);
	LUT4 #(
		.INIT('hab00)
	) name3000 (
		_w2915_,
		_w4896_,
		_w4897_,
		_w4900_,
		_w4901_
	);
	LUT2 #(
		.INIT('h4)
	) name3001 (
		\s15_msel_arb3_state_reg[1]/NET0131 ,
		_w4901_,
		_w4902_
	);
	LUT4 #(
		.INIT('hab00)
	) name3002 (
		_w2915_,
		_w4896_,
		_w4897_,
		_w4899_,
		_w4903_
	);
	LUT3 #(
		.INIT('h0d)
	) name3003 (
		_w2905_,
		_w2906_,
		_w2909_,
		_w4904_
	);
	LUT4 #(
		.INIT('h5504)
	) name3004 (
		\s15_msel_arb3_state_reg[2]/NET0131 ,
		_w2905_,
		_w2906_,
		_w2909_,
		_w4905_
	);
	LUT3 #(
		.INIT('hf2)
	) name3005 (
		_w2912_,
		_w2913_,
		_w2915_,
		_w4906_
	);
	LUT2 #(
		.INIT('h1)
	) name3006 (
		_w2906_,
		_w2914_,
		_w4907_
	);
	LUT3 #(
		.INIT('h01)
	) name3007 (
		\s15_msel_arb3_state_reg[2]/NET0131 ,
		_w2906_,
		_w2914_,
		_w4908_
	);
	LUT3 #(
		.INIT('h15)
	) name3008 (
		_w4905_,
		_w4906_,
		_w4908_,
		_w4909_
	);
	LUT3 #(
		.INIT('h02)
	) name3009 (
		\s15_msel_arb3_state_reg[0]/NET0131 ,
		_w2908_,
		_w2913_,
		_w4910_
	);
	LUT2 #(
		.INIT('h8)
	) name3010 (
		_w4907_,
		_w4910_,
		_w4911_
	);
	LUT2 #(
		.INIT('h2)
	) name3011 (
		\s15_msel_arb3_state_reg[0]/NET0131 ,
		\s15_msel_arb3_state_reg[1]/NET0131 ,
		_w4912_
	);
	LUT4 #(
		.INIT('hfb00)
	) name3012 (
		_w4903_,
		_w4909_,
		_w4911_,
		_w4912_,
		_w4913_
	);
	LUT2 #(
		.INIT('h1)
	) name3013 (
		_w4902_,
		_w4913_,
		_w4914_
	);
	LUT4 #(
		.INIT('h007f)
	) name3014 (
		\m0_s15_cyc_o_reg/NET0131 ,
		\rf_conf15_reg[0]/NET0131 ,
		\rf_conf15_reg[1]/NET0131 ,
		\s15_msel_arb3_state_reg[1]/NET0131 ,
		_w4915_
	);
	LUT4 #(
		.INIT('hea00)
	) name3015 (
		_w4905_,
		_w4906_,
		_w4908_,
		_w4915_,
		_w4916_
	);
	LUT2 #(
		.INIT('h4)
	) name3016 (
		\s15_msel_arb3_state_reg[0]/NET0131 ,
		_w4916_,
		_w4917_
	);
	LUT3 #(
		.INIT('h04)
	) name3017 (
		_w2908_,
		_w2909_,
		_w2913_,
		_w4918_
	);
	LUT4 #(
		.INIT('hccc8)
	) name3018 (
		_w4906_,
		_w4907_,
		_w4910_,
		_w4918_,
		_w4919_
	);
	LUT4 #(
		.INIT('h0080)
	) name3019 (
		\m2_s15_cyc_o_reg/NET0131 ,
		\rf_conf15_reg[4]/NET0131 ,
		\rf_conf15_reg[5]/NET0131 ,
		\s15_msel_arb3_state_reg[0]/NET0131 ,
		_w4920_
	);
	LUT4 #(
		.INIT('h5501)
	) name3020 (
		\s15_msel_arb3_state_reg[2]/NET0131 ,
		_w2905_,
		_w2906_,
		_w4920_,
		_w4921_
	);
	LUT2 #(
		.INIT('h4)
	) name3021 (
		_w4919_,
		_w4921_,
		_w4922_
	);
	LUT4 #(
		.INIT('h0080)
	) name3022 (
		\m6_s15_cyc_o_reg/NET0131 ,
		\rf_conf15_reg[12]/NET0131 ,
		\rf_conf15_reg[13]/NET0131 ,
		\s15_msel_arb3_state_reg[0]/NET0131 ,
		_w4923_
	);
	LUT4 #(
		.INIT('haa02)
	) name3023 (
		\s15_msel_arb3_state_reg[2]/NET0131 ,
		_w2912_,
		_w2913_,
		_w4923_,
		_w4924_
	);
	LUT2 #(
		.INIT('h2)
	) name3024 (
		\s15_msel_arb3_state_reg[1]/NET0131 ,
		_w4924_,
		_w4925_
	);
	LUT4 #(
		.INIT('h007f)
	) name3025 (
		\m5_s15_cyc_o_reg/NET0131 ,
		\rf_conf15_reg[10]/NET0131 ,
		\rf_conf15_reg[11]/NET0131 ,
		\s15_msel_arb3_state_reg[0]/NET0131 ,
		_w4926_
	);
	LUT3 #(
		.INIT('h01)
	) name3026 (
		_w2906_,
		_w2914_,
		_w4926_,
		_w4927_
	);
	LUT3 #(
		.INIT('h02)
	) name3027 (
		\s15_msel_arb3_state_reg[1]/NET0131 ,
		_w2908_,
		_w2913_,
		_w4928_
	);
	LUT3 #(
		.INIT('hd0)
	) name3028 (
		_w4904_,
		_w4927_,
		_w4928_,
		_w4929_
	);
	LUT3 #(
		.INIT('h54)
	) name3029 (
		\s15_msel_arb3_state_reg[0]/NET0131 ,
		_w4925_,
		_w4929_,
		_w4930_
	);
	LUT3 #(
		.INIT('h45)
	) name3030 (
		_w4917_,
		_w4922_,
		_w4930_,
		_w4931_
	);
	LUT3 #(
		.INIT('h51)
	) name3031 (
		_w2908_,
		_w2913_,
		_w2915_,
		_w4932_
	);
	LUT3 #(
		.INIT('h2a)
	) name3032 (
		\s15_msel_arb3_state_reg[2]/NET0131 ,
		_w4927_,
		_w4932_,
		_w4933_
	);
	LUT2 #(
		.INIT('h4)
	) name3033 (
		_w4898_,
		_w4933_,
		_w4934_
	);
	LUT3 #(
		.INIT('h54)
	) name3034 (
		_w2914_,
		_w4906_,
		_w4918_,
		_w4935_
	);
	LUT3 #(
		.INIT('h2a)
	) name3035 (
		_w2923_,
		_w4907_,
		_w4910_,
		_w4936_
	);
	LUT3 #(
		.INIT('h8a)
	) name3036 (
		_w2922_,
		_w4935_,
		_w4936_,
		_w4937_
	);
	LUT2 #(
		.INIT('h4)
	) name3037 (
		_w4934_,
		_w4937_,
		_w4938_
	);
	LUT3 #(
		.INIT('hf7)
	) name3038 (
		_w4914_,
		_w4931_,
		_w4938_,
		_w4939_
	);
	LUT2 #(
		.INIT('h4)
	) name3039 (
		_w2649_,
		_w2654_,
		_w4940_
	);
	LUT4 #(
		.INIT('h000d)
	) name3040 (
		_w2644_,
		_w2645_,
		_w2649_,
		_w2653_,
		_w4941_
	);
	LUT3 #(
		.INIT('h01)
	) name3041 (
		_w2645_,
		_w2647_,
		_w2654_,
		_w4942_
	);
	LUT4 #(
		.INIT('h00fd)
	) name3042 (
		\m5_s1_cyc_o_reg/NET0131 ,
		\rf_conf1_reg[10]/NET0131 ,
		\rf_conf1_reg[11]/NET0131 ,
		\s1_msel_arb0_state_reg[0]/NET0131 ,
		_w4943_
	);
	LUT3 #(
		.INIT('hce)
	) name3043 (
		\s1_msel_arb0_state_reg[0]/NET0131 ,
		_w2648_,
		_w2650_,
		_w4944_
	);
	LUT4 #(
		.INIT('h0eee)
	) name3044 (
		_w4940_,
		_w4941_,
		_w4942_,
		_w4944_,
		_w4945_
	);
	LUT3 #(
		.INIT('hae)
	) name3045 (
		_w2648_,
		_w2649_,
		_w2650_,
		_w4946_
	);
	LUT2 #(
		.INIT('h4)
	) name3046 (
		\s1_msel_arb0_state_reg[1]/NET0131 ,
		\s1_msel_arb0_state_reg[2]/NET0131 ,
		_w4947_
	);
	LUT4 #(
		.INIT('h0002)
	) name3047 (
		\m1_s1_cyc_o_reg/NET0131 ,
		\rf_conf1_reg[2]/NET0131 ,
		\rf_conf1_reg[3]/NET0131 ,
		\s1_msel_arb0_state_reg[1]/NET0131 ,
		_w4948_
	);
	LUT2 #(
		.INIT('h1)
	) name3048 (
		_w4947_,
		_w4948_,
		_w4949_
	);
	LUT3 #(
		.INIT('h23)
	) name3049 (
		_w2644_,
		_w2645_,
		_w2647_,
		_w4950_
	);
	LUT4 #(
		.INIT('h00dc)
	) name3050 (
		_w2644_,
		_w2645_,
		_w2647_,
		_w2653_,
		_w4951_
	);
	LUT3 #(
		.INIT('ha8)
	) name3051 (
		\s1_msel_arb0_state_reg[2]/NET0131 ,
		_w2650_,
		_w2654_,
		_w4952_
	);
	LUT4 #(
		.INIT('hdddc)
	) name3052 (
		_w4946_,
		_w4949_,
		_w4951_,
		_w4952_,
		_w4953_
	);
	LUT4 #(
		.INIT('h08aa)
	) name3053 (
		\s1_msel_arb0_state_reg[0]/NET0131 ,
		_w2677_,
		_w4945_,
		_w4953_,
		_w4954_
	);
	LUT3 #(
		.INIT('h02)
	) name3054 (
		\s1_msel_arb0_state_reg[0]/NET0131 ,
		_w2650_,
		_w2654_,
		_w4955_
	);
	LUT2 #(
		.INIT('h1)
	) name3055 (
		_w2645_,
		_w2647_,
		_w4956_
	);
	LUT3 #(
		.INIT('h80)
	) name3056 (
		_w2672_,
		_w4955_,
		_w4956_,
		_w4957_
	);
	LUT3 #(
		.INIT('h04)
	) name3057 (
		_w2650_,
		_w2653_,
		_w2654_,
		_w4958_
	);
	LUT4 #(
		.INIT('h1101)
	) name3058 (
		_w2644_,
		_w2648_,
		_w2649_,
		_w2650_,
		_w4959_
	);
	LUT4 #(
		.INIT('h0002)
	) name3059 (
		\m2_s1_cyc_o_reg/NET0131 ,
		\rf_conf1_reg[4]/NET0131 ,
		\rf_conf1_reg[5]/NET0131 ,
		\s1_msel_arb0_state_reg[0]/NET0131 ,
		_w4960_
	);
	LUT4 #(
		.INIT('h00b0)
	) name3060 (
		_w2644_,
		_w2647_,
		_w2672_,
		_w4960_,
		_w4961_
	);
	LUT3 #(
		.INIT('hb0)
	) name3061 (
		_w4958_,
		_w4959_,
		_w4961_,
		_w4962_
	);
	LUT2 #(
		.INIT('h1)
	) name3062 (
		_w4957_,
		_w4962_,
		_w4963_
	);
	LUT4 #(
		.INIT('h00f2)
	) name3063 (
		_w2644_,
		_w2645_,
		_w2653_,
		_w2654_,
		_w4964_
	);
	LUT3 #(
		.INIT('ha8)
	) name3064 (
		\s1_msel_arb0_state_reg[2]/NET0131 ,
		_w2647_,
		_w2650_,
		_w4965_
	);
	LUT3 #(
		.INIT('h54)
	) name3065 (
		\s1_msel_arb0_state_reg[2]/NET0131 ,
		_w2645_,
		_w2654_,
		_w4966_
	);
	LUT4 #(
		.INIT('h4454)
	) name3066 (
		_w2647_,
		_w2648_,
		_w2649_,
		_w2650_,
		_w4967_
	);
	LUT4 #(
		.INIT('hd0dd)
	) name3067 (
		_w4964_,
		_w4965_,
		_w4966_,
		_w4967_,
		_w4968_
	);
	LUT2 #(
		.INIT('h1)
	) name3068 (
		\s1_msel_arb0_state_reg[0]/NET0131 ,
		\s1_msel_arb0_state_reg[1]/NET0131 ,
		_w4969_
	);
	LUT3 #(
		.INIT('h02)
	) name3069 (
		\s1_msel_arb0_state_reg[0]/NET0131 ,
		\s1_msel_arb0_state_reg[1]/NET0131 ,
		\s1_msel_arb0_state_reg[2]/NET0131 ,
		_w4970_
	);
	LUT2 #(
		.INIT('h4)
	) name3070 (
		_w2653_,
		_w4970_,
		_w4971_
	);
	LUT4 #(
		.INIT('h8a00)
	) name3071 (
		_w4950_,
		_w4955_,
		_w4959_,
		_w4971_,
		_w4972_
	);
	LUT4 #(
		.INIT('h0001)
	) name3072 (
		_w2645_,
		_w2647_,
		_w2654_,
		_w4943_,
		_w4973_
	);
	LUT3 #(
		.INIT('h40)
	) name3073 (
		\s1_msel_arb0_state_reg[0]/NET0131 ,
		\s1_msel_arb0_state_reg[1]/NET0131 ,
		\s1_msel_arb0_state_reg[2]/NET0131 ,
		_w4974_
	);
	LUT2 #(
		.INIT('h4)
	) name3074 (
		_w2650_,
		_w4974_,
		_w4975_
	);
	LUT4 #(
		.INIT('hf100)
	) name3075 (
		_w4940_,
		_w4941_,
		_w4973_,
		_w4975_,
		_w4976_
	);
	LUT4 #(
		.INIT('h000b)
	) name3076 (
		_w4968_,
		_w4969_,
		_w4972_,
		_w4976_,
		_w4977_
	);
	LUT3 #(
		.INIT('hbf)
	) name3077 (
		_w4954_,
		_w4963_,
		_w4977_,
		_w4978_
	);
	LUT2 #(
		.INIT('h2)
	) name3078 (
		_w3699_,
		_w3704_,
		_w4979_
	);
	LUT4 #(
		.INIT('h000b)
	) name3079 (
		_w3696_,
		_w3697_,
		_w3700_,
		_w3704_,
		_w4980_
	);
	LUT2 #(
		.INIT('h1)
	) name3080 (
		\s1_msel_arb1_state_reg[1]/NET0131 ,
		\s1_msel_arb1_state_reg[2]/NET0131 ,
		_w4981_
	);
	LUT4 #(
		.INIT('h0d00)
	) name3081 (
		_w3708_,
		_w3709_,
		_w3714_,
		_w4981_,
		_w4982_
	);
	LUT4 #(
		.INIT('hab00)
	) name3082 (
		_w3709_,
		_w4979_,
		_w4980_,
		_w4982_,
		_w4983_
	);
	LUT2 #(
		.INIT('h2)
	) name3083 (
		\s1_msel_arb1_state_reg[1]/NET0131 ,
		\s1_msel_arb1_state_reg[2]/NET0131 ,
		_w4984_
	);
	LUT3 #(
		.INIT('h20)
	) name3084 (
		_w3704_,
		_w3708_,
		_w4984_,
		_w4985_
	);
	LUT3 #(
		.INIT('h0b)
	) name3085 (
		_w3696_,
		_w3697_,
		_w3700_,
		_w4986_
	);
	LUT2 #(
		.INIT('h1)
	) name3086 (
		_w3696_,
		_w3714_,
		_w4987_
	);
	LUT4 #(
		.INIT('h00f7)
	) name3087 (
		\m1_s1_cyc_o_reg/NET0131 ,
		\rf_conf1_reg[2]/NET0131 ,
		\rf_conf1_reg[3]/NET0131 ,
		\s1_msel_arb1_state_reg[0]/NET0131 ,
		_w4988_
	);
	LUT3 #(
		.INIT('h01)
	) name3088 (
		_w3696_,
		_w3714_,
		_w4988_,
		_w4989_
	);
	LUT3 #(
		.INIT('h10)
	) name3089 (
		_w3699_,
		_w3708_,
		_w4984_,
		_w4990_
	);
	LUT4 #(
		.INIT('h0455)
	) name3090 (
		_w4985_,
		_w4986_,
		_w4989_,
		_w4990_,
		_w4991_
	);
	LUT2 #(
		.INIT('h4)
	) name3091 (
		_w3699_,
		_w3702_,
		_w4992_
	);
	LUT3 #(
		.INIT('h0d)
	) name3092 (
		_w3704_,
		_w3708_,
		_w3709_,
		_w4993_
	);
	LUT4 #(
		.INIT('haf2f)
	) name3093 (
		_w4986_,
		_w4987_,
		_w4992_,
		_w4993_,
		_w4994_
	);
	LUT4 #(
		.INIT('h4555)
	) name3094 (
		\s1_msel_arb1_state_reg[0]/NET0131 ,
		_w4983_,
		_w4991_,
		_w4994_,
		_w4995_
	);
	LUT4 #(
		.INIT('hf700)
	) name3095 (
		\m0_s1_cyc_o_reg/NET0131 ,
		\rf_conf1_reg[0]/NET0131 ,
		\rf_conf1_reg[1]/NET0131 ,
		\s1_msel_arb1_state_reg[0]/NET0131 ,
		_w4996_
	);
	LUT3 #(
		.INIT('h01)
	) name3096 (
		_w3696_,
		_w3699_,
		_w3708_,
		_w4997_
	);
	LUT4 #(
		.INIT('h0100)
	) name3097 (
		_w3696_,
		_w3699_,
		_w3708_,
		_w4996_,
		_w4998_
	);
	LUT4 #(
		.INIT('h0008)
	) name3098 (
		\m6_s1_cyc_o_reg/NET0131 ,
		\rf_conf1_reg[12]/NET0131 ,
		\rf_conf1_reg[13]/NET0131 ,
		\s1_msel_arb1_state_reg[0]/NET0131 ,
		_w4999_
	);
	LUT2 #(
		.INIT('h2)
	) name3099 (
		_w3697_,
		_w4999_,
		_w5000_
	);
	LUT3 #(
		.INIT('h04)
	) name3100 (
		_w3699_,
		_w3700_,
		_w3708_,
		_w5001_
	);
	LUT2 #(
		.INIT('h1)
	) name3101 (
		_w3714_,
		_w4999_,
		_w5002_
	);
	LUT4 #(
		.INIT('h0233)
	) name3102 (
		_w4993_,
		_w5000_,
		_w5001_,
		_w5002_,
		_w5003_
	);
	LUT2 #(
		.INIT('h8)
	) name3103 (
		\s1_msel_arb1_state_reg[1]/NET0131 ,
		\s1_msel_arb1_state_reg[2]/NET0131 ,
		_w5004_
	);
	LUT3 #(
		.INIT('hb0)
	) name3104 (
		_w4998_,
		_w5003_,
		_w5004_,
		_w5005_
	);
	LUT3 #(
		.INIT('h20)
	) name3105 (
		\s1_msel_arb1_state_reg[0]/NET0131 ,
		\s1_msel_arb1_state_reg[1]/NET0131 ,
		\s1_msel_arb1_state_reg[2]/NET0131 ,
		_w5006_
	);
	LUT4 #(
		.INIT('h00a2)
	) name3106 (
		_w4986_,
		_w4987_,
		_w4993_,
		_w4998_,
		_w5007_
	);
	LUT2 #(
		.INIT('h2)
	) name3107 (
		_w5006_,
		_w5007_,
		_w5008_
	);
	LUT2 #(
		.INIT('h1)
	) name3108 (
		_w3697_,
		_w4996_,
		_w5009_
	);
	LUT4 #(
		.INIT('h0a02)
	) name3109 (
		_w4993_,
		_w4997_,
		_w5001_,
		_w5009_,
		_w5010_
	);
	LUT3 #(
		.INIT('h02)
	) name3110 (
		\s1_msel_arb1_state_reg[0]/NET0131 ,
		\s1_msel_arb1_state_reg[1]/NET0131 ,
		\s1_msel_arb1_state_reg[2]/NET0131 ,
		_w5011_
	);
	LUT3 #(
		.INIT('h51)
	) name3111 (
		_w3699_,
		_w3708_,
		_w3709_,
		_w5012_
	);
	LUT4 #(
		.INIT('h0eee)
	) name3112 (
		_w4979_,
		_w4980_,
		_w4989_,
		_w5012_,
		_w5013_
	);
	LUT3 #(
		.INIT('h08)
	) name3113 (
		\s1_msel_arb1_state_reg[0]/NET0131 ,
		\s1_msel_arb1_state_reg[1]/NET0131 ,
		\s1_msel_arb1_state_reg[2]/NET0131 ,
		_w5014_
	);
	LUT4 #(
		.INIT('hb0bb)
	) name3114 (
		_w5010_,
		_w5011_,
		_w5013_,
		_w5014_,
		_w5015_
	);
	LUT4 #(
		.INIT('hfeff)
	) name3115 (
		_w4995_,
		_w5005_,
		_w5008_,
		_w5015_,
		_w5016_
	);
	LUT2 #(
		.INIT('h4)
	) name3116 (
		\s1_msel_arb2_state_reg[1]/NET0131 ,
		\s1_msel_arb2_state_reg[2]/NET0131 ,
		_w5017_
	);
	LUT3 #(
		.INIT('h20)
	) name3117 (
		_w3299_,
		_w3300_,
		_w5017_,
		_w5018_
	);
	LUT2 #(
		.INIT('h4)
	) name3118 (
		_w3302_,
		_w3314_,
		_w5019_
	);
	LUT2 #(
		.INIT('h2)
	) name3119 (
		_w3305_,
		_w3307_,
		_w5020_
	);
	LUT4 #(
		.INIT('h0051)
	) name3120 (
		_w3302_,
		_w3305_,
		_w3307_,
		_w3310_,
		_w5021_
	);
	LUT3 #(
		.INIT('h10)
	) name3121 (
		_w3300_,
		_w3301_,
		_w5017_,
		_w5022_
	);
	LUT4 #(
		.INIT('h5455)
	) name3122 (
		_w5018_,
		_w5019_,
		_w5021_,
		_w5022_,
		_w5023_
	);
	LUT2 #(
		.INIT('h1)
	) name3123 (
		\s1_msel_arb2_state_reg[0]/NET0131 ,
		_w5023_,
		_w5024_
	);
	LUT2 #(
		.INIT('h1)
	) name3124 (
		_w3300_,
		_w3307_,
		_w5025_
	);
	LUT3 #(
		.INIT('hf2)
	) name3125 (
		_w3300_,
		_w3305_,
		_w3307_,
		_w5026_
	);
	LUT3 #(
		.INIT('h45)
	) name3126 (
		_w3299_,
		_w3301_,
		_w3302_,
		_w5027_
	);
	LUT3 #(
		.INIT('h04)
	) name3127 (
		_w3301_,
		_w3310_,
		_w3314_,
		_w5028_
	);
	LUT3 #(
		.INIT('h02)
	) name3128 (
		\s1_msel_arb2_state_reg[0]/NET0131 ,
		_w3301_,
		_w3314_,
		_w5029_
	);
	LUT4 #(
		.INIT('h0004)
	) name3129 (
		_w5020_,
		_w5027_,
		_w5028_,
		_w5029_,
		_w5030_
	);
	LUT3 #(
		.INIT('h04)
	) name3130 (
		\s1_msel_arb2_state_reg[0]/NET0131 ,
		\s1_msel_arb2_state_reg[1]/NET0131 ,
		\s1_msel_arb2_state_reg[2]/NET0131 ,
		_w5031_
	);
	LUT3 #(
		.INIT('h10)
	) name3131 (
		_w5026_,
		_w5030_,
		_w5031_,
		_w5032_
	);
	LUT2 #(
		.INIT('h1)
	) name3132 (
		_w5024_,
		_w5032_,
		_w5033_
	);
	LUT4 #(
		.INIT('hdf00)
	) name3133 (
		\m6_s1_cyc_o_reg/NET0131 ,
		\rf_conf1_reg[12]/NET0131 ,
		\rf_conf1_reg[13]/NET0131 ,
		\s1_msel_arb2_state_reg[0]/NET0131 ,
		_w5034_
	);
	LUT2 #(
		.INIT('h1)
	) name3134 (
		_w3299_,
		_w5034_,
		_w5035_
	);
	LUT3 #(
		.INIT('h01)
	) name3135 (
		_w3300_,
		_w3307_,
		_w3314_,
		_w5036_
	);
	LUT4 #(
		.INIT('he0ee)
	) name3136 (
		_w5019_,
		_w5021_,
		_w5035_,
		_w5036_,
		_w5037_
	);
	LUT4 #(
		.INIT('h0020)
	) name3137 (
		\m6_s1_cyc_o_reg/NET0131 ,
		\rf_conf1_reg[12]/NET0131 ,
		\rf_conf1_reg[13]/NET0131 ,
		\s1_msel_arb2_state_reg[0]/NET0131 ,
		_w5038_
	);
	LUT2 #(
		.INIT('h8)
	) name3138 (
		\s1_msel_arb2_state_reg[1]/NET0131 ,
		\s1_msel_arb2_state_reg[2]/NET0131 ,
		_w5039_
	);
	LUT2 #(
		.INIT('h4)
	) name3139 (
		_w5038_,
		_w5039_,
		_w5040_
	);
	LUT2 #(
		.INIT('h4)
	) name3140 (
		_w5037_,
		_w5040_,
		_w5041_
	);
	LUT3 #(
		.INIT('h51)
	) name3141 (
		_w3300_,
		_w5027_,
		_w5028_,
		_w5042_
	);
	LUT2 #(
		.INIT('h8)
	) name3142 (
		_w5025_,
		_w5029_,
		_w5043_
	);
	LUT3 #(
		.INIT('h15)
	) name3143 (
		_w3305_,
		_w5025_,
		_w5029_,
		_w5044_
	);
	LUT3 #(
		.INIT('h08)
	) name3144 (
		\s1_msel_arb2_state_reg[0]/NET0131 ,
		\s1_msel_arb2_state_reg[1]/NET0131 ,
		\s1_msel_arb2_state_reg[2]/NET0131 ,
		_w5045_
	);
	LUT3 #(
		.INIT('hb0)
	) name3145 (
		_w5042_,
		_w5044_,
		_w5045_,
		_w5046_
	);
	LUT2 #(
		.INIT('h2)
	) name3146 (
		\s1_msel_arb2_state_reg[0]/NET0131 ,
		\s1_msel_arb2_state_reg[1]/NET0131 ,
		_w5047_
	);
	LUT3 #(
		.INIT('h20)
	) name3147 (
		\s1_msel_arb2_state_reg[0]/NET0131 ,
		\s1_msel_arb2_state_reg[1]/NET0131 ,
		\s1_msel_arb2_state_reg[2]/NET0131 ,
		_w5048_
	);
	LUT3 #(
		.INIT('h01)
	) name3148 (
		_w3301_,
		_w5019_,
		_w5021_,
		_w5049_
	);
	LUT3 #(
		.INIT('h15)
	) name3149 (
		_w3299_,
		_w5025_,
		_w5029_,
		_w5050_
	);
	LUT3 #(
		.INIT('h8a)
	) name3150 (
		_w5048_,
		_w5049_,
		_w5050_,
		_w5051_
	);
	LUT4 #(
		.INIT('h0020)
	) name3151 (
		\m0_s1_cyc_o_reg/NET0131 ,
		\rf_conf1_reg[0]/NET0131 ,
		\rf_conf1_reg[1]/NET0131 ,
		\s1_msel_arb2_state_reg[0]/NET0131 ,
		_w5052_
	);
	LUT4 #(
		.INIT('h00f2)
	) name3152 (
		_w3305_,
		_w3307_,
		_w3310_,
		_w5052_,
		_w5053_
	);
	LUT3 #(
		.INIT('h01)
	) name3153 (
		_w3300_,
		_w3307_,
		_w5052_,
		_w5054_
	);
	LUT3 #(
		.INIT('h23)
	) name3154 (
		_w5027_,
		_w5053_,
		_w5054_,
		_w5055_
	);
	LUT2 #(
		.INIT('h1)
	) name3155 (
		\s1_msel_arb2_state_reg[1]/NET0131 ,
		\s1_msel_arb2_state_reg[2]/NET0131 ,
		_w5056_
	);
	LUT3 #(
		.INIT('hb0)
	) name3156 (
		_w5043_,
		_w5055_,
		_w5056_,
		_w5057_
	);
	LUT4 #(
		.INIT('h0001)
	) name3157 (
		_w5041_,
		_w5046_,
		_w5051_,
		_w5057_,
		_w5058_
	);
	LUT2 #(
		.INIT('h7)
	) name3158 (
		_w5033_,
		_w5058_,
		_w5059_
	);
	LUT3 #(
		.INIT('hdc)
	) name3159 (
		_w3324_,
		_w3325_,
		_w3335_,
		_w5060_
	);
	LUT2 #(
		.INIT('h4)
	) name3160 (
		_w3327_,
		_w3329_,
		_w5061_
	);
	LUT4 #(
		.INIT('h000d)
	) name3161 (
		_w3322_,
		_w3323_,
		_w3327_,
		_w3328_,
		_w5062_
	);
	LUT4 #(
		.INIT('h7f00)
	) name3162 (
		\m6_s1_cyc_o_reg/NET0131 ,
		\rf_conf1_reg[12]/NET0131 ,
		\rf_conf1_reg[13]/NET0131 ,
		\s1_msel_arb3_state_reg[0]/NET0131 ,
		_w5063_
	);
	LUT4 #(
		.INIT('ha2f3)
	) name3163 (
		_w3323_,
		_w3324_,
		_w3325_,
		_w5063_,
		_w5064_
	);
	LUT4 #(
		.INIT('h0155)
	) name3164 (
		_w5060_,
		_w5061_,
		_w5062_,
		_w5064_,
		_w5065_
	);
	LUT2 #(
		.INIT('h8)
	) name3165 (
		_w3347_,
		_w5065_,
		_w5066_
	);
	LUT2 #(
		.INIT('h1)
	) name3166 (
		\s1_msel_arb3_state_reg[1]/NET0131 ,
		\s1_msel_arb3_state_reg[2]/NET0131 ,
		_w5067_
	);
	LUT3 #(
		.INIT('h20)
	) name3167 (
		_w3322_,
		_w3323_,
		_w5067_,
		_w5068_
	);
	LUT2 #(
		.INIT('h4)
	) name3168 (
		_w3324_,
		_w3335_,
		_w5069_
	);
	LUT4 #(
		.INIT('h1101)
	) name3169 (
		_w3324_,
		_w3327_,
		_w3328_,
		_w3329_,
		_w5070_
	);
	LUT3 #(
		.INIT('h10)
	) name3170 (
		_w3323_,
		_w3325_,
		_w5067_,
		_w5071_
	);
	LUT4 #(
		.INIT('h5455)
	) name3171 (
		_w5068_,
		_w5069_,
		_w5070_,
		_w5071_,
		_w5072_
	);
	LUT3 #(
		.INIT('h08)
	) name3172 (
		_w3321_,
		_w3327_,
		_w3335_,
		_w5073_
	);
	LUT3 #(
		.INIT('h0d)
	) name3173 (
		_w3322_,
		_w3323_,
		_w3328_,
		_w5074_
	);
	LUT3 #(
		.INIT('h04)
	) name3174 (
		_w3323_,
		_w3324_,
		_w3325_,
		_w5075_
	);
	LUT3 #(
		.INIT('h02)
	) name3175 (
		_w3321_,
		_w3329_,
		_w3335_,
		_w5076_
	);
	LUT4 #(
		.INIT('h0455)
	) name3176 (
		_w5073_,
		_w5074_,
		_w5075_,
		_w5076_,
		_w5077_
	);
	LUT3 #(
		.INIT('h40)
	) name3177 (
		\s1_msel_arb3_state_reg[0]/NET0131 ,
		_w5072_,
		_w5077_,
		_w5078_
	);
	LUT3 #(
		.INIT('h51)
	) name3178 (
		_w3329_,
		_w5074_,
		_w5075_,
		_w5079_
	);
	LUT4 #(
		.INIT('h0001)
	) name3179 (
		_w3323_,
		_w3325_,
		_w3329_,
		_w3335_,
		_w5080_
	);
	LUT2 #(
		.INIT('h1)
	) name3180 (
		_w3327_,
		_w5080_,
		_w5081_
	);
	LUT3 #(
		.INIT('h2a)
	) name3181 (
		\s1_msel_arb3_state_reg[0]/NET0131 ,
		_w3324_,
		_w3347_,
		_w5082_
	);
	LUT4 #(
		.INIT('h7500)
	) name3182 (
		_w3321_,
		_w5079_,
		_w5081_,
		_w5082_,
		_w5083_
	);
	LUT3 #(
		.INIT('h0b)
	) name3183 (
		_w5066_,
		_w5078_,
		_w5083_,
		_w5084_
	);
	LUT2 #(
		.INIT('h4)
	) name3184 (
		_w3322_,
		_w3325_,
		_w5085_
	);
	LUT4 #(
		.INIT('h5455)
	) name3185 (
		_w3322_,
		_w3323_,
		_w3335_,
		_w5063_,
		_w5086_
	);
	LUT4 #(
		.INIT('h010f)
	) name3186 (
		_w5069_,
		_w5070_,
		_w5085_,
		_w5086_,
		_w5087_
	);
	LUT3 #(
		.INIT('h02)
	) name3187 (
		\s1_msel_arb3_state_reg[0]/NET0131 ,
		\s1_msel_arb3_state_reg[1]/NET0131 ,
		\s1_msel_arb3_state_reg[2]/NET0131 ,
		_w5088_
	);
	LUT2 #(
		.INIT('h8)
	) name3188 (
		_w5087_,
		_w5088_,
		_w5089_
	);
	LUT2 #(
		.INIT('h1)
	) name3189 (
		_w3327_,
		_w5063_,
		_w5090_
	);
	LUT3 #(
		.INIT('h01)
	) name3190 (
		_w3323_,
		_w3325_,
		_w3335_,
		_w5091_
	);
	LUT4 #(
		.INIT('h2022)
	) name3191 (
		_w5074_,
		_w5075_,
		_w5090_,
		_w5091_,
		_w5092_
	);
	LUT4 #(
		.INIT('h0080)
	) name3192 (
		\m6_s1_cyc_o_reg/NET0131 ,
		\rf_conf1_reg[12]/NET0131 ,
		\rf_conf1_reg[13]/NET0131 ,
		\s1_msel_arb3_state_reg[0]/NET0131 ,
		_w5093_
	);
	LUT2 #(
		.INIT('h2)
	) name3193 (
		_w3333_,
		_w5093_,
		_w5094_
	);
	LUT3 #(
		.INIT('h10)
	) name3194 (
		_w3323_,
		_w3325_,
		_w5063_,
		_w5095_
	);
	LUT3 #(
		.INIT('h08)
	) name3195 (
		\s1_msel_arb3_state_reg[0]/NET0131 ,
		\s1_msel_arb3_state_reg[1]/NET0131 ,
		\s1_msel_arb3_state_reg[2]/NET0131 ,
		_w5096_
	);
	LUT3 #(
		.INIT('h10)
	) name3196 (
		_w3324_,
		_w3335_,
		_w5096_,
		_w5097_
	);
	LUT4 #(
		.INIT('hf100)
	) name3197 (
		_w5061_,
		_w5062_,
		_w5095_,
		_w5097_,
		_w5098_
	);
	LUT3 #(
		.INIT('h0b)
	) name3198 (
		_w5092_,
		_w5094_,
		_w5098_,
		_w5099_
	);
	LUT2 #(
		.INIT('h4)
	) name3199 (
		_w5089_,
		_w5099_,
		_w5100_
	);
	LUT2 #(
		.INIT('hb)
	) name3200 (
		_w5084_,
		_w5100_,
		_w5101_
	);
	LUT2 #(
		.INIT('h4)
	) name3201 (
		_w2688_,
		_w2693_,
		_w5102_
	);
	LUT4 #(
		.INIT('h000d)
	) name3202 (
		_w2683_,
		_w2684_,
		_w2688_,
		_w2692_,
		_w5103_
	);
	LUT3 #(
		.INIT('h01)
	) name3203 (
		_w2684_,
		_w2686_,
		_w2693_,
		_w5104_
	);
	LUT4 #(
		.INIT('h00fd)
	) name3204 (
		\m5_s2_cyc_o_reg/NET0131 ,
		\rf_conf2_reg[10]/NET0131 ,
		\rf_conf2_reg[11]/NET0131 ,
		\s2_msel_arb0_state_reg[0]/NET0131 ,
		_w5105_
	);
	LUT3 #(
		.INIT('hce)
	) name3205 (
		\s2_msel_arb0_state_reg[0]/NET0131 ,
		_w2687_,
		_w2689_,
		_w5106_
	);
	LUT4 #(
		.INIT('h0eee)
	) name3206 (
		_w5102_,
		_w5103_,
		_w5104_,
		_w5106_,
		_w5107_
	);
	LUT3 #(
		.INIT('hae)
	) name3207 (
		_w2687_,
		_w2688_,
		_w2689_,
		_w5108_
	);
	LUT2 #(
		.INIT('h4)
	) name3208 (
		\s2_msel_arb0_state_reg[1]/NET0131 ,
		\s2_msel_arb0_state_reg[2]/NET0131 ,
		_w5109_
	);
	LUT4 #(
		.INIT('h0002)
	) name3209 (
		\m1_s2_cyc_o_reg/NET0131 ,
		\rf_conf2_reg[2]/NET0131 ,
		\rf_conf2_reg[3]/NET0131 ,
		\s2_msel_arb0_state_reg[1]/NET0131 ,
		_w5110_
	);
	LUT2 #(
		.INIT('h1)
	) name3210 (
		_w5109_,
		_w5110_,
		_w5111_
	);
	LUT3 #(
		.INIT('h23)
	) name3211 (
		_w2683_,
		_w2684_,
		_w2686_,
		_w5112_
	);
	LUT4 #(
		.INIT('h00dc)
	) name3212 (
		_w2683_,
		_w2684_,
		_w2686_,
		_w2692_,
		_w5113_
	);
	LUT3 #(
		.INIT('ha8)
	) name3213 (
		\s2_msel_arb0_state_reg[2]/NET0131 ,
		_w2689_,
		_w2693_,
		_w5114_
	);
	LUT4 #(
		.INIT('hdddc)
	) name3214 (
		_w5108_,
		_w5111_,
		_w5113_,
		_w5114_,
		_w5115_
	);
	LUT4 #(
		.INIT('h08aa)
	) name3215 (
		\s2_msel_arb0_state_reg[0]/NET0131 ,
		_w2716_,
		_w5107_,
		_w5115_,
		_w5116_
	);
	LUT3 #(
		.INIT('h02)
	) name3216 (
		\s2_msel_arb0_state_reg[0]/NET0131 ,
		_w2689_,
		_w2693_,
		_w5117_
	);
	LUT2 #(
		.INIT('h1)
	) name3217 (
		_w2684_,
		_w2686_,
		_w5118_
	);
	LUT3 #(
		.INIT('h80)
	) name3218 (
		_w2711_,
		_w5117_,
		_w5118_,
		_w5119_
	);
	LUT3 #(
		.INIT('h04)
	) name3219 (
		_w2689_,
		_w2692_,
		_w2693_,
		_w5120_
	);
	LUT4 #(
		.INIT('h1101)
	) name3220 (
		_w2683_,
		_w2687_,
		_w2688_,
		_w2689_,
		_w5121_
	);
	LUT4 #(
		.INIT('h0002)
	) name3221 (
		\m2_s2_cyc_o_reg/NET0131 ,
		\rf_conf2_reg[4]/NET0131 ,
		\rf_conf2_reg[5]/NET0131 ,
		\s2_msel_arb0_state_reg[0]/NET0131 ,
		_w5122_
	);
	LUT4 #(
		.INIT('h00b0)
	) name3222 (
		_w2683_,
		_w2686_,
		_w2711_,
		_w5122_,
		_w5123_
	);
	LUT3 #(
		.INIT('hb0)
	) name3223 (
		_w5120_,
		_w5121_,
		_w5123_,
		_w5124_
	);
	LUT2 #(
		.INIT('h1)
	) name3224 (
		_w5119_,
		_w5124_,
		_w5125_
	);
	LUT4 #(
		.INIT('h00f2)
	) name3225 (
		_w2683_,
		_w2684_,
		_w2692_,
		_w2693_,
		_w5126_
	);
	LUT3 #(
		.INIT('ha8)
	) name3226 (
		\s2_msel_arb0_state_reg[2]/NET0131 ,
		_w2686_,
		_w2689_,
		_w5127_
	);
	LUT3 #(
		.INIT('h54)
	) name3227 (
		\s2_msel_arb0_state_reg[2]/NET0131 ,
		_w2684_,
		_w2693_,
		_w5128_
	);
	LUT4 #(
		.INIT('h4454)
	) name3228 (
		_w2686_,
		_w2687_,
		_w2688_,
		_w2689_,
		_w5129_
	);
	LUT4 #(
		.INIT('hd0dd)
	) name3229 (
		_w5126_,
		_w5127_,
		_w5128_,
		_w5129_,
		_w5130_
	);
	LUT2 #(
		.INIT('h1)
	) name3230 (
		\s2_msel_arb0_state_reg[0]/NET0131 ,
		\s2_msel_arb0_state_reg[1]/NET0131 ,
		_w5131_
	);
	LUT3 #(
		.INIT('h02)
	) name3231 (
		\s2_msel_arb0_state_reg[0]/NET0131 ,
		\s2_msel_arb0_state_reg[1]/NET0131 ,
		\s2_msel_arb0_state_reg[2]/NET0131 ,
		_w5132_
	);
	LUT2 #(
		.INIT('h4)
	) name3232 (
		_w2692_,
		_w5132_,
		_w5133_
	);
	LUT4 #(
		.INIT('h8a00)
	) name3233 (
		_w5112_,
		_w5117_,
		_w5121_,
		_w5133_,
		_w5134_
	);
	LUT4 #(
		.INIT('h0001)
	) name3234 (
		_w2684_,
		_w2686_,
		_w2693_,
		_w5105_,
		_w5135_
	);
	LUT3 #(
		.INIT('h40)
	) name3235 (
		\s2_msel_arb0_state_reg[0]/NET0131 ,
		\s2_msel_arb0_state_reg[1]/NET0131 ,
		\s2_msel_arb0_state_reg[2]/NET0131 ,
		_w5136_
	);
	LUT2 #(
		.INIT('h4)
	) name3236 (
		_w2689_,
		_w5136_,
		_w5137_
	);
	LUT4 #(
		.INIT('hf100)
	) name3237 (
		_w5102_,
		_w5103_,
		_w5135_,
		_w5137_,
		_w5138_
	);
	LUT4 #(
		.INIT('h000b)
	) name3238 (
		_w5130_,
		_w5131_,
		_w5134_,
		_w5138_,
		_w5139_
	);
	LUT3 #(
		.INIT('hbf)
	) name3239 (
		_w5116_,
		_w5125_,
		_w5139_,
		_w5140_
	);
	LUT3 #(
		.INIT('h23)
	) name3240 (
		_w3722_,
		_w3724_,
		_w3734_,
		_w5141_
	);
	LUT4 #(
		.INIT('h2232)
	) name3241 (
		_w3722_,
		_w3724_,
		_w3733_,
		_w3734_,
		_w5142_
	);
	LUT2 #(
		.INIT('h1)
	) name3242 (
		_w3724_,
		_w3734_,
		_w5143_
	);
	LUT4 #(
		.INIT('h0004)
	) name3243 (
		_w3724_,
		_w3730_,
		_w3731_,
		_w3734_,
		_w5144_
	);
	LUT2 #(
		.INIT('h2)
	) name3244 (
		\s2_msel_arb1_state_reg[1]/NET0131 ,
		\s2_msel_arb1_state_reg[2]/NET0131 ,
		_w5145_
	);
	LUT2 #(
		.INIT('h4)
	) name3245 (
		_w3727_,
		_w5145_,
		_w5146_
	);
	LUT4 #(
		.INIT('hfe00)
	) name3246 (
		_w3728_,
		_w5142_,
		_w5144_,
		_w5146_,
		_w5147_
	);
	LUT3 #(
		.INIT('hdc)
	) name3247 (
		_w3722_,
		_w3724_,
		_w3734_,
		_w5148_
	);
	LUT2 #(
		.INIT('h2)
	) name3248 (
		_w3731_,
		_w3733_,
		_w5149_
	);
	LUT2 #(
		.INIT('h4)
	) name3249 (
		_w3727_,
		_w3728_,
		_w5150_
	);
	LUT4 #(
		.INIT('h000b)
	) name3250 (
		_w3727_,
		_w3728_,
		_w3730_,
		_w3733_,
		_w5151_
	);
	LUT4 #(
		.INIT('hf700)
	) name3251 (
		\m0_s2_cyc_o_reg/NET0131 ,
		\rf_conf2_reg[0]/NET0131 ,
		\rf_conf2_reg[1]/NET0131 ,
		\s2_msel_arb1_state_reg[0]/NET0131 ,
		_w5152_
	);
	LUT4 #(
		.INIT('hd0dd)
	) name3252 (
		_w3722_,
		_w3724_,
		_w3727_,
		_w5152_,
		_w5153_
	);
	LUT4 #(
		.INIT('h0155)
	) name3253 (
		_w5148_,
		_w5149_,
		_w5151_,
		_w5153_,
		_w5154_
	);
	LUT2 #(
		.INIT('h4)
	) name3254 (
		\s2_msel_arb1_state_reg[1]/NET0131 ,
		\s2_msel_arb1_state_reg[2]/NET0131 ,
		_w5155_
	);
	LUT4 #(
		.INIT('habbb)
	) name3255 (
		\s2_msel_arb1_state_reg[0]/NET0131 ,
		_w5147_,
		_w5154_,
		_w5155_,
		_w5156_
	);
	LUT4 #(
		.INIT('hff0d)
	) name3256 (
		\s2_msel_arb1_state_reg[0]/NET0131 ,
		_w3727_,
		_w3730_,
		_w3731_,
		_w5157_
	);
	LUT4 #(
		.INIT('h1101)
	) name3257 (
		_w3728_,
		_w5142_,
		_w5143_,
		_w5157_,
		_w5158_
	);
	LUT2 #(
		.INIT('h2)
	) name3258 (
		_w5145_,
		_w5158_,
		_w5159_
	);
	LUT2 #(
		.INIT('h1)
	) name3259 (
		\s2_msel_arb1_state_reg[1]/NET0131 ,
		\s2_msel_arb1_state_reg[2]/NET0131 ,
		_w5160_
	);
	LUT3 #(
		.INIT('h0b)
	) name3260 (
		_w3727_,
		_w3728_,
		_w3730_,
		_w5161_
	);
	LUT3 #(
		.INIT('h02)
	) name3261 (
		_w3722_,
		_w3724_,
		_w3727_,
		_w5162_
	);
	LUT3 #(
		.INIT('h01)
	) name3262 (
		_w3724_,
		_w3727_,
		_w3734_,
		_w5163_
	);
	LUT2 #(
		.INIT('h1)
	) name3263 (
		_w3733_,
		_w5152_,
		_w5164_
	);
	LUT4 #(
		.INIT('h2202)
	) name3264 (
		_w5161_,
		_w5162_,
		_w5163_,
		_w5164_,
		_w5165_
	);
	LUT4 #(
		.INIT('h5455)
	) name3265 (
		_w3722_,
		_w3724_,
		_w3727_,
		_w5152_,
		_w5166_
	);
	LUT3 #(
		.INIT('hb0)
	) name3266 (
		_w3722_,
		_w3734_,
		_w5155_,
		_w5167_
	);
	LUT4 #(
		.INIT('h1f00)
	) name3267 (
		_w5149_,
		_w5151_,
		_w5166_,
		_w5167_,
		_w5168_
	);
	LUT3 #(
		.INIT('h0d)
	) name3268 (
		_w5160_,
		_w5165_,
		_w5168_,
		_w5169_
	);
	LUT3 #(
		.INIT('h8a)
	) name3269 (
		\s2_msel_arb1_state_reg[0]/NET0131 ,
		_w5159_,
		_w5169_,
		_w5170_
	);
	LUT4 #(
		.INIT('h0008)
	) name3270 (
		\m6_s2_cyc_o_reg/NET0131 ,
		\rf_conf2_reg[12]/NET0131 ,
		\rf_conf2_reg[13]/NET0131 ,
		\s2_msel_arb1_state_reg[0]/NET0131 ,
		_w5171_
	);
	LUT2 #(
		.INIT('h8)
	) name3271 (
		\s2_msel_arb1_state_reg[1]/NET0131 ,
		\s2_msel_arb1_state_reg[2]/NET0131 ,
		_w5172_
	);
	LUT2 #(
		.INIT('h4)
	) name3272 (
		_w5171_,
		_w5172_,
		_w5173_
	);
	LUT3 #(
		.INIT('h20)
	) name3273 (
		_w3733_,
		_w5171_,
		_w5172_,
		_w5174_
	);
	LUT4 #(
		.INIT('hf700)
	) name3274 (
		\m2_s2_cyc_o_reg/NET0131 ,
		\rf_conf2_reg[4]/NET0131 ,
		\rf_conf2_reg[5]/NET0131 ,
		\s2_msel_arb1_state_reg[0]/NET0131 ,
		_w5175_
	);
	LUT3 #(
		.INIT('h10)
	) name3275 (
		_w3724_,
		_w3734_,
		_w5175_,
		_w5176_
	);
	LUT4 #(
		.INIT('hf0d0)
	) name3276 (
		_w5161_,
		_w5162_,
		_w5173_,
		_w5176_,
		_w5177_
	);
	LUT3 #(
		.INIT('h32)
	) name3277 (
		_w3722_,
		_w3727_,
		_w3733_,
		_w5178_
	);
	LUT4 #(
		.INIT('h0105)
	) name3278 (
		_w3730_,
		_w5141_,
		_w5150_,
		_w5178_,
		_w5179_
	);
	LUT3 #(
		.INIT('h01)
	) name3279 (
		\s2_msel_arb1_state_reg[0]/NET0131 ,
		\s2_msel_arb1_state_reg[1]/NET0131 ,
		\s2_msel_arb1_state_reg[2]/NET0131 ,
		_w5180_
	);
	LUT4 #(
		.INIT('hbabb)
	) name3280 (
		_w3731_,
		_w5177_,
		_w5179_,
		_w5180_,
		_w5181_
	);
	LUT2 #(
		.INIT('h4)
	) name3281 (
		_w5174_,
		_w5181_,
		_w5182_
	);
	LUT3 #(
		.INIT('hdf)
	) name3282 (
		_w5156_,
		_w5170_,
		_w5182_,
		_w5183_
	);
	LUT3 #(
		.INIT('h20)
	) name3283 (
		\m4_s2_cyc_o_reg/NET0131 ,
		\rf_conf2_reg[8]/NET0131 ,
		\rf_conf2_reg[9]/NET0131 ,
		_w5184_
	);
	LUT3 #(
		.INIT('h20)
	) name3284 (
		\m7_s2_cyc_o_reg/NET0131 ,
		\rf_conf2_reg[14]/NET0131 ,
		\rf_conf2_reg[15]/NET0131 ,
		_w5185_
	);
	LUT3 #(
		.INIT('h20)
	) name3285 (
		\m0_s2_cyc_o_reg/NET0131 ,
		\rf_conf2_reg[0]/NET0131 ,
		\rf_conf2_reg[1]/NET0131 ,
		_w5186_
	);
	LUT2 #(
		.INIT('h4)
	) name3286 (
		_w5185_,
		_w5186_,
		_w5187_
	);
	LUT3 #(
		.INIT('h20)
	) name3287 (
		\m3_s2_cyc_o_reg/NET0131 ,
		\rf_conf2_reg[6]/NET0131 ,
		\rf_conf2_reg[7]/NET0131 ,
		_w5188_
	);
	LUT3 #(
		.INIT('h20)
	) name3288 (
		\m2_s2_cyc_o_reg/NET0131 ,
		\rf_conf2_reg[4]/NET0131 ,
		\rf_conf2_reg[5]/NET0131 ,
		_w5189_
	);
	LUT3 #(
		.INIT('h20)
	) name3289 (
		\m1_s2_cyc_o_reg/NET0131 ,
		\rf_conf2_reg[2]/NET0131 ,
		\rf_conf2_reg[3]/NET0131 ,
		_w5190_
	);
	LUT4 #(
		.INIT('h0051)
	) name3290 (
		_w5185_,
		_w5188_,
		_w5189_,
		_w5190_,
		_w5191_
	);
	LUT3 #(
		.INIT('h20)
	) name3291 (
		\m5_s2_cyc_o_reg/NET0131 ,
		\rf_conf2_reg[10]/NET0131 ,
		\rf_conf2_reg[11]/NET0131 ,
		_w5192_
	);
	LUT3 #(
		.INIT('h20)
	) name3292 (
		\m6_s2_cyc_o_reg/NET0131 ,
		\rf_conf2_reg[12]/NET0131 ,
		\rf_conf2_reg[13]/NET0131 ,
		_w5193_
	);
	LUT3 #(
		.INIT('h8a)
	) name3293 (
		\s2_msel_arb2_state_reg[0]/NET0131 ,
		_w5192_,
		_w5193_,
		_w5194_
	);
	LUT4 #(
		.INIT('hf100)
	) name3294 (
		_w5187_,
		_w5191_,
		_w5192_,
		_w5194_,
		_w5195_
	);
	LUT2 #(
		.INIT('h1)
	) name3295 (
		_w5186_,
		_w5193_,
		_w5196_
	);
	LUT4 #(
		.INIT('hdf00)
	) name3296 (
		\m2_s2_cyc_o_reg/NET0131 ,
		\rf_conf2_reg[4]/NET0131 ,
		\rf_conf2_reg[5]/NET0131 ,
		\s2_msel_arb2_state_reg[0]/NET0131 ,
		_w5197_
	);
	LUT4 #(
		.INIT('h3030)
	) name3297 (
		_w5186_,
		_w5192_,
		_w5193_,
		_w5197_,
		_w5198_
	);
	LUT4 #(
		.INIT('h3233)
	) name3298 (
		_w5186_,
		_w5192_,
		_w5193_,
		_w5197_,
		_w5199_
	);
	LUT4 #(
		.INIT('h010f)
	) name3299 (
		_w5187_,
		_w5191_,
		_w5198_,
		_w5199_,
		_w5200_
	);
	LUT2 #(
		.INIT('h4)
	) name3300 (
		\s2_msel_arb2_state_reg[1]/NET0131 ,
		\s2_msel_arb2_state_reg[2]/NET0131 ,
		_w5201_
	);
	LUT4 #(
		.INIT('hd000)
	) name3301 (
		_w5184_,
		_w5195_,
		_w5200_,
		_w5201_,
		_w5202_
	);
	LUT2 #(
		.INIT('h8)
	) name3302 (
		\s2_msel_arb2_state_reg[1]/NET0131 ,
		\s2_msel_arb2_state_reg[2]/NET0131 ,
		_w5203_
	);
	LUT3 #(
		.INIT('h20)
	) name3303 (
		_w5185_,
		_w5193_,
		_w5203_,
		_w5204_
	);
	LUT3 #(
		.INIT('h0d)
	) name3304 (
		_w5188_,
		_w5189_,
		_w5190_,
		_w5205_
	);
	LUT4 #(
		.INIT('h00df)
	) name3305 (
		\m5_s2_cyc_o_reg/NET0131 ,
		\rf_conf2_reg[10]/NET0131 ,
		\rf_conf2_reg[11]/NET0131 ,
		\s2_msel_arb2_state_reg[0]/NET0131 ,
		_w5206_
	);
	LUT3 #(
		.INIT('h01)
	) name3306 (
		_w5184_,
		_w5189_,
		_w5206_,
		_w5207_
	);
	LUT3 #(
		.INIT('h10)
	) name3307 (
		_w5186_,
		_w5193_,
		_w5203_,
		_w5208_
	);
	LUT4 #(
		.INIT('h0455)
	) name3308 (
		_w5204_,
		_w5205_,
		_w5207_,
		_w5208_,
		_w5209_
	);
	LUT2 #(
		.INIT('h1)
	) name3309 (
		\s2_msel_arb2_state_reg[1]/NET0131 ,
		\s2_msel_arb2_state_reg[2]/NET0131 ,
		_w5210_
	);
	LUT3 #(
		.INIT('h40)
	) name3310 (
		_w5186_,
		_w5190_,
		_w5210_,
		_w5211_
	);
	LUT2 #(
		.INIT('h2)
	) name3311 (
		_w5184_,
		_w5188_,
		_w5212_
	);
	LUT4 #(
		.INIT('h0301)
	) name3312 (
		_w5185_,
		_w5188_,
		_w5192_,
		_w5193_,
		_w5213_
	);
	LUT3 #(
		.INIT('h10)
	) name3313 (
		_w5186_,
		_w5189_,
		_w5210_,
		_w5214_
	);
	LUT4 #(
		.INIT('h5455)
	) name3314 (
		_w5211_,
		_w5212_,
		_w5213_,
		_w5214_,
		_w5215_
	);
	LUT3 #(
		.INIT('h15)
	) name3315 (
		\s2_msel_arb2_state_reg[0]/NET0131 ,
		_w5209_,
		_w5215_,
		_w5216_
	);
	LUT3 #(
		.INIT('h80)
	) name3316 (
		\s2_msel_arb2_state_reg[0]/NET0131 ,
		_w5190_,
		_w5210_,
		_w5217_
	);
	LUT3 #(
		.INIT('h45)
	) name3317 (
		_w5186_,
		_w5192_,
		_w5193_,
		_w5218_
	);
	LUT4 #(
		.INIT('h0eee)
	) name3318 (
		_w5187_,
		_w5191_,
		_w5207_,
		_w5218_,
		_w5219_
	);
	LUT3 #(
		.INIT('h80)
	) name3319 (
		\s2_msel_arb2_state_reg[0]/NET0131 ,
		\s2_msel_arb2_state_reg[1]/NET0131 ,
		\s2_msel_arb2_state_reg[2]/NET0131 ,
		_w5220_
	);
	LUT3 #(
		.INIT('h45)
	) name3320 (
		_w5217_,
		_w5219_,
		_w5220_,
		_w5221_
	);
	LUT3 #(
		.INIT('h40)
	) name3321 (
		_w5190_,
		_w5197_,
		_w5210_,
		_w5222_
	);
	LUT4 #(
		.INIT('h0020)
	) name3322 (
		\m2_s2_cyc_o_reg/NET0131 ,
		\rf_conf2_reg[4]/NET0131 ,
		\rf_conf2_reg[5]/NET0131 ,
		\s2_msel_arb2_state_reg[0]/NET0131 ,
		_w5223_
	);
	LUT2 #(
		.INIT('h2)
	) name3323 (
		\s2_msel_arb2_state_reg[1]/NET0131 ,
		\s2_msel_arb2_state_reg[2]/NET0131 ,
		_w5224_
	);
	LUT2 #(
		.INIT('h4)
	) name3324 (
		_w5223_,
		_w5224_,
		_w5225_
	);
	LUT4 #(
		.INIT('h1110)
	) name3325 (
		_w5212_,
		_w5213_,
		_w5222_,
		_w5225_,
		_w5226_
	);
	LUT3 #(
		.INIT('h40)
	) name3326 (
		_w5184_,
		_w5196_,
		_w5222_,
		_w5227_
	);
	LUT4 #(
		.INIT('hfafb)
	) name3327 (
		_w5186_,
		_w5190_,
		_w5193_,
		_w5197_,
		_w5228_
	);
	LUT3 #(
		.INIT('h10)
	) name3328 (
		_w5184_,
		_w5223_,
		_w5224_,
		_w5229_
	);
	LUT2 #(
		.INIT('h4)
	) name3329 (
		_w5228_,
		_w5229_,
		_w5230_
	);
	LUT3 #(
		.INIT('h01)
	) name3330 (
		_w5226_,
		_w5227_,
		_w5230_,
		_w5231_
	);
	LUT4 #(
		.INIT('hefff)
	) name3331 (
		_w5202_,
		_w5216_,
		_w5221_,
		_w5231_,
		_w5232_
	);
	LUT2 #(
		.INIT('h2)
	) name3332 (
		\s2_msel_arb3_state_reg[1]/NET0131 ,
		\s2_msel_arb3_state_reg[2]/NET0131 ,
		_w5233_
	);
	LUT2 #(
		.INIT('h4)
	) name3333 (
		_w3021_,
		_w5233_,
		_w5234_
	);
	LUT2 #(
		.INIT('h1)
	) name3334 (
		_w3003_,
		_w3010_,
		_w5235_
	);
	LUT3 #(
		.INIT('hae)
	) name3335 (
		_w3003_,
		_w3010_,
		_w3011_,
		_w5236_
	);
	LUT2 #(
		.INIT('h1)
	) name3336 (
		_w3015_,
		_w3026_,
		_w5237_
	);
	LUT2 #(
		.INIT('h1)
	) name3337 (
		_w3011_,
		_w3016_,
		_w5238_
	);
	LUT4 #(
		.INIT('h7577)
	) name3338 (
		_w5234_,
		_w5236_,
		_w5237_,
		_w5238_,
		_w5239_
	);
	LUT3 #(
		.INIT('h0d)
	) name3339 (
		_w3013_,
		_w3014_,
		_w3015_,
		_w5240_
	);
	LUT4 #(
		.INIT('h00f2)
	) name3340 (
		_w3013_,
		_w3014_,
		_w3015_,
		_w3016_,
		_w5241_
	);
	LUT3 #(
		.INIT('h10)
	) name3341 (
		\s2_msel_arb3_state_reg[0]/NET0131 ,
		\s2_msel_arb3_state_reg[1]/NET0131 ,
		\s2_msel_arb3_state_reg[2]/NET0131 ,
		_w5242_
	);
	LUT4 #(
		.INIT('h2300)
	) name3342 (
		_w3003_,
		_w3004_,
		_w3011_,
		_w5242_,
		_w5243_
	);
	LUT3 #(
		.INIT('hd0)
	) name3343 (
		_w5235_,
		_w5241_,
		_w5243_,
		_w5244_
	);
	LUT3 #(
		.INIT('h0e)
	) name3344 (
		_w3004_,
		_w5239_,
		_w5244_,
		_w5245_
	);
	LUT2 #(
		.INIT('h1)
	) name3345 (
		\s2_msel_arb3_state_reg[1]/NET0131 ,
		\s2_msel_arb3_state_reg[2]/NET0131 ,
		_w5246_
	);
	LUT4 #(
		.INIT('h0080)
	) name3346 (
		\m0_s2_cyc_o_reg/NET0131 ,
		\rf_conf2_reg[0]/NET0131 ,
		\rf_conf2_reg[1]/NET0131 ,
		\s2_msel_arb3_state_reg[0]/NET0131 ,
		_w5247_
	);
	LUT2 #(
		.INIT('h2)
	) name3347 (
		_w5246_,
		_w5247_,
		_w5248_
	);
	LUT2 #(
		.INIT('h1)
	) name3348 (
		_w3004_,
		_w3014_,
		_w5249_
	);
	LUT4 #(
		.INIT('h4fcf)
	) name3349 (
		_w5236_,
		_w5240_,
		_w5248_,
		_w5249_,
		_w5250_
	);
	LUT3 #(
		.INIT('h20)
	) name3350 (
		_w3013_,
		_w3021_,
		_w5233_,
		_w5251_
	);
	LUT3 #(
		.INIT('h20)
	) name3351 (
		\s2_msel_arb3_state_reg[0]/NET0131 ,
		\s2_msel_arb3_state_reg[1]/NET0131 ,
		\s2_msel_arb3_state_reg[2]/NET0131 ,
		_w5252_
	);
	LUT2 #(
		.INIT('h8)
	) name3352 (
		_w3003_,
		_w5252_,
		_w5253_
	);
	LUT2 #(
		.INIT('h1)
	) name3353 (
		_w5251_,
		_w5253_,
		_w5254_
	);
	LUT2 #(
		.INIT('h8)
	) name3354 (
		_w5250_,
		_w5254_,
		_w5255_
	);
	LUT3 #(
		.INIT('h02)
	) name3355 (
		\s2_msel_arb3_state_reg[0]/NET0131 ,
		\s2_msel_arb3_state_reg[1]/NET0131 ,
		\s2_msel_arb3_state_reg[2]/NET0131 ,
		_w5256_
	);
	LUT4 #(
		.INIT('h0100)
	) name3356 (
		_w3004_,
		_w3014_,
		_w3016_,
		_w5256_,
		_w5257_
	);
	LUT2 #(
		.INIT('h4)
	) name3357 (
		_w3003_,
		_w5252_,
		_w5258_
	);
	LUT2 #(
		.INIT('h1)
	) name3358 (
		_w5257_,
		_w5258_,
		_w5259_
	);
	LUT2 #(
		.INIT('h4)
	) name3359 (
		_w3010_,
		_w3016_,
		_w5260_
	);
	LUT4 #(
		.INIT('h0051)
	) name3360 (
		_w3010_,
		_w3013_,
		_w3014_,
		_w3015_,
		_w5261_
	);
	LUT4 #(
		.INIT('h7f00)
	) name3361 (
		\m0_s2_cyc_o_reg/NET0131 ,
		\rf_conf2_reg[0]/NET0131 ,
		\rf_conf2_reg[1]/NET0131 ,
		\s2_msel_arb3_state_reg[0]/NET0131 ,
		_w5262_
	);
	LUT3 #(
		.INIT('h10)
	) name3362 (
		_w3004_,
		_w3014_,
		_w5262_,
		_w5263_
	);
	LUT4 #(
		.INIT('h0054)
	) name3363 (
		_w5257_,
		_w5260_,
		_w5261_,
		_w5263_,
		_w5264_
	);
	LUT3 #(
		.INIT('h01)
	) name3364 (
		_w3011_,
		_w5259_,
		_w5264_,
		_w5265_
	);
	LUT4 #(
		.INIT('h007f)
	) name3365 (
		\m5_s2_cyc_o_reg/NET0131 ,
		\rf_conf2_reg[10]/NET0131 ,
		\rf_conf2_reg[11]/NET0131 ,
		\s2_msel_arb3_state_reg[0]/NET0131 ,
		_w5266_
	);
	LUT4 #(
		.INIT('h0001)
	) name3366 (
		_w3004_,
		_w3014_,
		_w3016_,
		_w5266_,
		_w5267_
	);
	LUT3 #(
		.INIT('h0e)
	) name3367 (
		_w5260_,
		_w5261_,
		_w5267_,
		_w5268_
	);
	LUT4 #(
		.INIT('h0080)
	) name3368 (
		\m6_s2_cyc_o_reg/NET0131 ,
		\rf_conf2_reg[12]/NET0131 ,
		\rf_conf2_reg[13]/NET0131 ,
		\s2_msel_arb3_state_reg[0]/NET0131 ,
		_w5269_
	);
	LUT3 #(
		.INIT('h10)
	) name3369 (
		_w3003_,
		_w3010_,
		_w3011_,
		_w5270_
	);
	LUT4 #(
		.INIT('h020a)
	) name3370 (
		_w3029_,
		_w5240_,
		_w5269_,
		_w5270_,
		_w5271_
	);
	LUT2 #(
		.INIT('h4)
	) name3371 (
		_w5268_,
		_w5271_,
		_w5272_
	);
	LUT4 #(
		.INIT('hfff7)
	) name3372 (
		_w5245_,
		_w5255_,
		_w5265_,
		_w5272_,
		_w5273_
	);
	LUT2 #(
		.INIT('h4)
	) name3373 (
		_w2464_,
		_w2472_,
		_w5274_
	);
	LUT3 #(
		.INIT('h04)
	) name3374 (
		_w2460_,
		_w2462_,
		_w2463_,
		_w5275_
	);
	LUT4 #(
		.INIT('hfd00)
	) name3375 (
		\m4_s3_cyc_o_reg/NET0131 ,
		\rf_conf3_reg[8]/NET0131 ,
		\rf_conf3_reg[9]/NET0131 ,
		\s3_msel_arb0_state_reg[0]/NET0131 ,
		_w5276_
	);
	LUT3 #(
		.INIT('h10)
	) name3376 (
		_w2463_,
		_w2465_,
		_w5276_,
		_w5277_
	);
	LUT3 #(
		.INIT('hf2)
	) name3377 (
		_w2459_,
		_w2460_,
		_w2467_,
		_w5278_
	);
	LUT4 #(
		.INIT('h000d)
	) name3378 (
		_w2459_,
		_w2460_,
		_w2464_,
		_w2467_,
		_w5279_
	);
	LUT4 #(
		.INIT('h5455)
	) name3379 (
		_w5274_,
		_w5275_,
		_w5277_,
		_w5279_,
		_w5280_
	);
	LUT2 #(
		.INIT('h8)
	) name3380 (
		_w2486_,
		_w5280_,
		_w5281_
	);
	LUT2 #(
		.INIT('h8)
	) name3381 (
		\s3_msel_arb0_state_reg[1]/NET0131 ,
		\s3_msel_arb0_state_reg[2]/NET0131 ,
		_w5282_
	);
	LUT2 #(
		.INIT('h2)
	) name3382 (
		_w2467_,
		_w2472_,
		_w5283_
	);
	LUT3 #(
		.INIT('h51)
	) name3383 (
		_w2464_,
		_w2467_,
		_w2472_,
		_w5284_
	);
	LUT4 #(
		.INIT('h2232)
	) name3384 (
		_w2464_,
		_w2465_,
		_w2467_,
		_w2472_,
		_w5285_
	);
	LUT2 #(
		.INIT('h1)
	) name3385 (
		_w2460_,
		_w2472_,
		_w5286_
	);
	LUT4 #(
		.INIT('h00fd)
	) name3386 (
		\m5_s3_cyc_o_reg/NET0131 ,
		\rf_conf3_reg[10]/NET0131 ,
		\rf_conf3_reg[11]/NET0131 ,
		\s3_msel_arb0_state_reg[0]/NET0131 ,
		_w5287_
	);
	LUT3 #(
		.INIT('h01)
	) name3387 (
		_w2460_,
		_w2472_,
		_w5287_,
		_w5288_
	);
	LUT2 #(
		.INIT('h4)
	) name3388 (
		_w2459_,
		_w2463_,
		_w5289_
	);
	LUT3 #(
		.INIT('h0b)
	) name3389 (
		_w2459_,
		_w2463_,
		_w2465_,
		_w5290_
	);
	LUT4 #(
		.INIT('h0111)
	) name3390 (
		_w2462_,
		_w5285_,
		_w5288_,
		_w5290_,
		_w5291_
	);
	LUT4 #(
		.INIT('h1101)
	) name3391 (
		_w2459_,
		_w2462_,
		_w2464_,
		_w2465_,
		_w5292_
	);
	LUT4 #(
		.INIT('hfd00)
	) name3392 (
		\m2_s3_cyc_o_reg/NET0131 ,
		\rf_conf3_reg[4]/NET0131 ,
		\rf_conf3_reg[5]/NET0131 ,
		\s3_msel_arb0_state_reg[0]/NET0131 ,
		_w5293_
	);
	LUT4 #(
		.INIT('h0e0f)
	) name3393 (
		_w2463_,
		_w2465_,
		_w2467_,
		_w5293_,
		_w5294_
	);
	LUT2 #(
		.INIT('h2)
	) name3394 (
		\s3_msel_arb0_state_reg[1]/NET0131 ,
		\s3_msel_arb0_state_reg[2]/NET0131 ,
		_w5295_
	);
	LUT3 #(
		.INIT('hd0)
	) name3395 (
		_w2460_,
		_w2467_,
		_w5295_,
		_w5296_
	);
	LUT4 #(
		.INIT('h1f00)
	) name3396 (
		_w5289_,
		_w5292_,
		_w5294_,
		_w5296_,
		_w5297_
	);
	LUT3 #(
		.INIT('h0d)
	) name3397 (
		_w5282_,
		_w5291_,
		_w5297_,
		_w5298_
	);
	LUT3 #(
		.INIT('h8a)
	) name3398 (
		\s3_msel_arb0_state_reg[0]/NET0131 ,
		_w5281_,
		_w5298_,
		_w5299_
	);
	LUT3 #(
		.INIT('h02)
	) name3399 (
		\s3_msel_arb0_state_reg[0]/NET0131 ,
		_w2463_,
		_w2465_,
		_w5300_
	);
	LUT4 #(
		.INIT('h55fd)
	) name3400 (
		_w5286_,
		_w5289_,
		_w5292_,
		_w5300_,
		_w5301_
	);
	LUT3 #(
		.INIT('h8c)
	) name3401 (
		_w5283_,
		_w5295_,
		_w5301_,
		_w5302_
	);
	LUT3 #(
		.INIT('h20)
	) name3402 (
		_w2462_,
		_w2463_,
		_w5282_,
		_w5303_
	);
	LUT3 #(
		.INIT('h10)
	) name3403 (
		_w2463_,
		_w2465_,
		_w5282_,
		_w5304_
	);
	LUT4 #(
		.INIT('h020f)
	) name3404 (
		_w5284_,
		_w5288_,
		_w5303_,
		_w5304_,
		_w5305_
	);
	LUT3 #(
		.INIT('h20)
	) name3405 (
		_w2464_,
		_w2465_,
		_w2486_,
		_w5306_
	);
	LUT2 #(
		.INIT('h1)
	) name3406 (
		_w2460_,
		_w2463_,
		_w5307_
	);
	LUT4 #(
		.INIT('h00fd)
	) name3407 (
		\m7_s3_cyc_o_reg/NET0131 ,
		\rf_conf3_reg[14]/NET0131 ,
		\rf_conf3_reg[15]/NET0131 ,
		\s3_msel_arb0_state_reg[0]/NET0131 ,
		_w5308_
	);
	LUT3 #(
		.INIT('h01)
	) name3408 (
		_w2460_,
		_w2463_,
		_w5308_,
		_w5309_
	);
	LUT3 #(
		.INIT('h10)
	) name3409 (
		_w2465_,
		_w2472_,
		_w2486_,
		_w5310_
	);
	LUT4 #(
		.INIT('h0133)
	) name3410 (
		_w5278_,
		_w5306_,
		_w5309_,
		_w5310_,
		_w5311_
	);
	LUT2 #(
		.INIT('h8)
	) name3411 (
		_w5305_,
		_w5311_,
		_w5312_
	);
	LUT3 #(
		.INIT('h02)
	) name3412 (
		\s3_msel_arb0_state_reg[0]/NET0131 ,
		_w2465_,
		_w2472_,
		_w5313_
	);
	LUT3 #(
		.INIT('h80)
	) name3413 (
		_w2489_,
		_w5307_,
		_w5313_,
		_w5314_
	);
	LUT3 #(
		.INIT('h04)
	) name3414 (
		_w2465_,
		_w2467_,
		_w2472_,
		_w5315_
	);
	LUT4 #(
		.INIT('h0002)
	) name3415 (
		\m4_s3_cyc_o_reg/NET0131 ,
		\rf_conf3_reg[8]/NET0131 ,
		\rf_conf3_reg[9]/NET0131 ,
		\s3_msel_arb0_state_reg[0]/NET0131 ,
		_w5316_
	);
	LUT4 #(
		.INIT('h00b0)
	) name3416 (
		_w2459_,
		_w2463_,
		_w2489_,
		_w5316_,
		_w5317_
	);
	LUT3 #(
		.INIT('hd0)
	) name3417 (
		_w5292_,
		_w5315_,
		_w5317_,
		_w5318_
	);
	LUT2 #(
		.INIT('h1)
	) name3418 (
		_w5314_,
		_w5318_,
		_w5319_
	);
	LUT4 #(
		.INIT('hba00)
	) name3419 (
		\s3_msel_arb0_state_reg[0]/NET0131 ,
		_w5302_,
		_w5312_,
		_w5319_,
		_w5320_
	);
	LUT2 #(
		.INIT('hb)
	) name3420 (
		_w5299_,
		_w5320_,
		_w5321_
	);
	LUT2 #(
		.INIT('h4)
	) name3421 (
		_w3756_,
		_w3757_,
		_w5322_
	);
	LUT3 #(
		.INIT('h0b)
	) name3422 (
		_w3756_,
		_w3757_,
		_w3759_,
		_w5323_
	);
	LUT3 #(
		.INIT('h04)
	) name3423 (
		_w3752_,
		_w3753_,
		_w3756_,
		_w5324_
	);
	LUT3 #(
		.INIT('h51)
	) name3424 (
		_w3760_,
		_w5323_,
		_w5324_,
		_w5325_
	);
	LUT4 #(
		.INIT('hf700)
	) name3425 (
		\m0_s3_cyc_o_reg/NET0131 ,
		\rf_conf3_reg[0]/NET0131 ,
		\rf_conf3_reg[1]/NET0131 ,
		\s3_msel_arb1_state_reg[0]/NET0131 ,
		_w5326_
	);
	LUT3 #(
		.INIT('h10)
	) name3426 (
		_w3752_,
		_w3756_,
		_w5326_,
		_w5327_
	);
	LUT4 #(
		.INIT('h5455)
	) name3427 (
		_w3748_,
		_w3752_,
		_w3756_,
		_w5326_,
		_w5328_
	);
	LUT4 #(
		.INIT('hae00)
	) name3428 (
		_w3760_,
		_w5323_,
		_w5324_,
		_w5328_,
		_w5329_
	);
	LUT2 #(
		.INIT('h8)
	) name3429 (
		\s3_msel_arb1_state_reg[1]/NET0131 ,
		\s3_msel_arb1_state_reg[2]/NET0131 ,
		_w5330_
	);
	LUT2 #(
		.INIT('h4)
	) name3430 (
		_w3749_,
		_w5330_,
		_w5331_
	);
	LUT4 #(
		.INIT('h00f4)
	) name3431 (
		_w3756_,
		_w3757_,
		_w3759_,
		_w3760_,
		_w5332_
	);
	LUT2 #(
		.INIT('h1)
	) name3432 (
		_w3748_,
		_w3753_,
		_w5333_
	);
	LUT2 #(
		.INIT('h4)
	) name3433 (
		_w3756_,
		_w5326_,
		_w5334_
	);
	LUT4 #(
		.INIT('h1011)
	) name3434 (
		_w3748_,
		_w3753_,
		_w3756_,
		_w5326_,
		_w5335_
	);
	LUT2 #(
		.INIT('h4)
	) name3435 (
		\s3_msel_arb1_state_reg[1]/NET0131 ,
		\s3_msel_arb1_state_reg[2]/NET0131 ,
		_w5336_
	);
	LUT4 #(
		.INIT('h3100)
	) name3436 (
		_w3749_,
		_w3752_,
		_w3753_,
		_w5336_,
		_w5337_
	);
	LUT3 #(
		.INIT('hb0)
	) name3437 (
		_w5332_,
		_w5335_,
		_w5337_,
		_w5338_
	);
	LUT2 #(
		.INIT('h1)
	) name3438 (
		\s3_msel_arb1_state_reg[1]/NET0131 ,
		\s3_msel_arb1_state_reg[2]/NET0131 ,
		_w5339_
	);
	LUT2 #(
		.INIT('h4)
	) name3439 (
		_w3760_,
		_w5339_,
		_w5340_
	);
	LUT4 #(
		.INIT('h0031)
	) name3440 (
		_w3749_,
		_w3752_,
		_w3753_,
		_w3756_,
		_w5341_
	);
	LUT4 #(
		.INIT('h8faf)
	) name3441 (
		_w5323_,
		_w5333_,
		_w5340_,
		_w5341_,
		_w5342_
	);
	LUT4 #(
		.INIT('h0b00)
	) name3442 (
		_w5329_,
		_w5331_,
		_w5338_,
		_w5342_,
		_w5343_
	);
	LUT4 #(
		.INIT('h1101)
	) name3443 (
		_w3748_,
		_w3753_,
		_w3759_,
		_w3760_,
		_w5344_
	);
	LUT4 #(
		.INIT('h88a8)
	) name3444 (
		_w3747_,
		_w5322_,
		_w5341_,
		_w5344_,
		_w5345_
	);
	LUT4 #(
		.INIT('hf700)
	) name3445 (
		\m3_s3_cyc_o_reg/NET0131 ,
		\rf_conf3_reg[6]/NET0131 ,
		\rf_conf3_reg[7]/NET0131 ,
		\s3_msel_arb1_state_reg[1]/NET0131 ,
		_w5346_
	);
	LUT2 #(
		.INIT('h2)
	) name3446 (
		\s3_msel_arb1_state_reg[0]/NET0131 ,
		_w5346_,
		_w5347_
	);
	LUT4 #(
		.INIT('h0a02)
	) name3447 (
		\s3_msel_arb1_state_reg[0]/NET0131 ,
		_w3749_,
		_w3752_,
		_w3753_,
		_w5348_
	);
	LUT4 #(
		.INIT('h040f)
	) name3448 (
		_w5334_,
		_w5344_,
		_w5347_,
		_w5348_,
		_w5349_
	);
	LUT2 #(
		.INIT('h1)
	) name3449 (
		_w3748_,
		_w5326_,
		_w5350_
	);
	LUT3 #(
		.INIT('h01)
	) name3450 (
		_w3749_,
		_w3752_,
		_w3756_,
		_w5351_
	);
	LUT4 #(
		.INIT('h00f7)
	) name3451 (
		\m1_s3_cyc_o_reg/NET0131 ,
		\rf_conf3_reg[2]/NET0131 ,
		\rf_conf3_reg[3]/NET0131 ,
		\s3_msel_arb1_state_reg[1]/NET0131 ,
		_w5352_
	);
	LUT3 #(
		.INIT('hb0)
	) name3452 (
		_w3756_,
		_w3757_,
		_w5352_,
		_w5353_
	);
	LUT4 #(
		.INIT('h4500)
	) name3453 (
		_w5324_,
		_w5350_,
		_w5351_,
		_w5353_,
		_w5354_
	);
	LUT4 #(
		.INIT('hbbba)
	) name3454 (
		\s3_msel_arb1_state_reg[2]/NET0131 ,
		_w5345_,
		_w5349_,
		_w5354_,
		_w5355_
	);
	LUT4 #(
		.INIT('h0001)
	) name3455 (
		_w3749_,
		_w3752_,
		_w3756_,
		_w3760_,
		_w5356_
	);
	LUT2 #(
		.INIT('h1)
	) name3456 (
		_w3748_,
		_w5356_,
		_w5357_
	);
	LUT3 #(
		.INIT('h80)
	) name3457 (
		\s3_msel_arb1_state_reg[0]/NET0131 ,
		\s3_msel_arb1_state_reg[1]/NET0131 ,
		\s3_msel_arb1_state_reg[2]/NET0131 ,
		_w5358_
	);
	LUT3 #(
		.INIT('h20)
	) name3458 (
		\s3_msel_arb1_state_reg[0]/NET0131 ,
		\s3_msel_arb1_state_reg[1]/NET0131 ,
		\s3_msel_arb1_state_reg[2]/NET0131 ,
		_w5359_
	);
	LUT3 #(
		.INIT('hd0)
	) name3459 (
		_w3749_,
		_w3753_,
		_w5359_,
		_w5360_
	);
	LUT4 #(
		.INIT('hef00)
	) name3460 (
		_w5327_,
		_w5332_,
		_w5333_,
		_w5360_,
		_w5361_
	);
	LUT4 #(
		.INIT('h004f)
	) name3461 (
		_w5325_,
		_w5357_,
		_w5358_,
		_w5361_,
		_w5362_
	);
	LUT4 #(
		.INIT('h1fff)
	) name3462 (
		\s3_msel_arb1_state_reg[0]/NET0131 ,
		_w5343_,
		_w5355_,
		_w5362_,
		_w5363_
	);
	LUT2 #(
		.INIT('h4)
	) name3463 (
		\s3_msel_arb2_state_reg[1]/NET0131 ,
		\s3_msel_arb2_state_reg[2]/NET0131 ,
		_w5364_
	);
	LUT3 #(
		.INIT('h20)
	) name3464 (
		_w3033_,
		_w3034_,
		_w5364_,
		_w5365_
	);
	LUT2 #(
		.INIT('h4)
	) name3465 (
		_w3036_,
		_w3048_,
		_w5366_
	);
	LUT2 #(
		.INIT('h2)
	) name3466 (
		_w3039_,
		_w3041_,
		_w5367_
	);
	LUT4 #(
		.INIT('h0051)
	) name3467 (
		_w3036_,
		_w3039_,
		_w3041_,
		_w3044_,
		_w5368_
	);
	LUT3 #(
		.INIT('h10)
	) name3468 (
		_w3034_,
		_w3035_,
		_w5364_,
		_w5369_
	);
	LUT4 #(
		.INIT('h5455)
	) name3469 (
		_w5365_,
		_w5366_,
		_w5368_,
		_w5369_,
		_w5370_
	);
	LUT2 #(
		.INIT('h1)
	) name3470 (
		\s3_msel_arb2_state_reg[0]/NET0131 ,
		_w5370_,
		_w5371_
	);
	LUT2 #(
		.INIT('h1)
	) name3471 (
		_w3034_,
		_w3041_,
		_w5372_
	);
	LUT3 #(
		.INIT('hf2)
	) name3472 (
		_w3034_,
		_w3039_,
		_w3041_,
		_w5373_
	);
	LUT3 #(
		.INIT('h45)
	) name3473 (
		_w3033_,
		_w3035_,
		_w3036_,
		_w5374_
	);
	LUT3 #(
		.INIT('h04)
	) name3474 (
		_w3035_,
		_w3044_,
		_w3048_,
		_w5375_
	);
	LUT3 #(
		.INIT('h02)
	) name3475 (
		\s3_msel_arb2_state_reg[0]/NET0131 ,
		_w3035_,
		_w3048_,
		_w5376_
	);
	LUT4 #(
		.INIT('h0004)
	) name3476 (
		_w5367_,
		_w5374_,
		_w5375_,
		_w5376_,
		_w5377_
	);
	LUT3 #(
		.INIT('h04)
	) name3477 (
		\s3_msel_arb2_state_reg[0]/NET0131 ,
		\s3_msel_arb2_state_reg[1]/NET0131 ,
		\s3_msel_arb2_state_reg[2]/NET0131 ,
		_w5378_
	);
	LUT3 #(
		.INIT('h10)
	) name3478 (
		_w5373_,
		_w5377_,
		_w5378_,
		_w5379_
	);
	LUT2 #(
		.INIT('h1)
	) name3479 (
		_w5371_,
		_w5379_,
		_w5380_
	);
	LUT4 #(
		.INIT('hdf00)
	) name3480 (
		\m6_s3_cyc_o_reg/NET0131 ,
		\rf_conf3_reg[12]/NET0131 ,
		\rf_conf3_reg[13]/NET0131 ,
		\s3_msel_arb2_state_reg[0]/NET0131 ,
		_w5381_
	);
	LUT2 #(
		.INIT('h1)
	) name3481 (
		_w3033_,
		_w5381_,
		_w5382_
	);
	LUT3 #(
		.INIT('h01)
	) name3482 (
		_w3034_,
		_w3041_,
		_w3048_,
		_w5383_
	);
	LUT4 #(
		.INIT('he0ee)
	) name3483 (
		_w5366_,
		_w5368_,
		_w5382_,
		_w5383_,
		_w5384_
	);
	LUT4 #(
		.INIT('h0020)
	) name3484 (
		\m6_s3_cyc_o_reg/NET0131 ,
		\rf_conf3_reg[12]/NET0131 ,
		\rf_conf3_reg[13]/NET0131 ,
		\s3_msel_arb2_state_reg[0]/NET0131 ,
		_w5385_
	);
	LUT2 #(
		.INIT('h8)
	) name3485 (
		\s3_msel_arb2_state_reg[1]/NET0131 ,
		\s3_msel_arb2_state_reg[2]/NET0131 ,
		_w5386_
	);
	LUT2 #(
		.INIT('h4)
	) name3486 (
		_w5385_,
		_w5386_,
		_w5387_
	);
	LUT2 #(
		.INIT('h4)
	) name3487 (
		_w5384_,
		_w5387_,
		_w5388_
	);
	LUT3 #(
		.INIT('h51)
	) name3488 (
		_w3034_,
		_w5374_,
		_w5375_,
		_w5389_
	);
	LUT2 #(
		.INIT('h8)
	) name3489 (
		_w5372_,
		_w5376_,
		_w5390_
	);
	LUT3 #(
		.INIT('h15)
	) name3490 (
		_w3039_,
		_w5372_,
		_w5376_,
		_w5391_
	);
	LUT3 #(
		.INIT('h08)
	) name3491 (
		\s3_msel_arb2_state_reg[0]/NET0131 ,
		\s3_msel_arb2_state_reg[1]/NET0131 ,
		\s3_msel_arb2_state_reg[2]/NET0131 ,
		_w5392_
	);
	LUT3 #(
		.INIT('hb0)
	) name3492 (
		_w5389_,
		_w5391_,
		_w5392_,
		_w5393_
	);
	LUT2 #(
		.INIT('h2)
	) name3493 (
		\s3_msel_arb2_state_reg[0]/NET0131 ,
		\s3_msel_arb2_state_reg[1]/NET0131 ,
		_w5394_
	);
	LUT3 #(
		.INIT('h20)
	) name3494 (
		\s3_msel_arb2_state_reg[0]/NET0131 ,
		\s3_msel_arb2_state_reg[1]/NET0131 ,
		\s3_msel_arb2_state_reg[2]/NET0131 ,
		_w5395_
	);
	LUT3 #(
		.INIT('h01)
	) name3495 (
		_w3035_,
		_w5366_,
		_w5368_,
		_w5396_
	);
	LUT3 #(
		.INIT('h15)
	) name3496 (
		_w3033_,
		_w5372_,
		_w5376_,
		_w5397_
	);
	LUT3 #(
		.INIT('h8a)
	) name3497 (
		_w5395_,
		_w5396_,
		_w5397_,
		_w5398_
	);
	LUT4 #(
		.INIT('h0020)
	) name3498 (
		\m0_s3_cyc_o_reg/NET0131 ,
		\rf_conf3_reg[0]/NET0131 ,
		\rf_conf3_reg[1]/NET0131 ,
		\s3_msel_arb2_state_reg[0]/NET0131 ,
		_w5399_
	);
	LUT4 #(
		.INIT('h00f2)
	) name3499 (
		_w3039_,
		_w3041_,
		_w3044_,
		_w5399_,
		_w5400_
	);
	LUT3 #(
		.INIT('h01)
	) name3500 (
		_w3034_,
		_w3041_,
		_w5399_,
		_w5401_
	);
	LUT3 #(
		.INIT('h23)
	) name3501 (
		_w5374_,
		_w5400_,
		_w5401_,
		_w5402_
	);
	LUT2 #(
		.INIT('h1)
	) name3502 (
		\s3_msel_arb2_state_reg[1]/NET0131 ,
		\s3_msel_arb2_state_reg[2]/NET0131 ,
		_w5403_
	);
	LUT3 #(
		.INIT('hb0)
	) name3503 (
		_w5390_,
		_w5402_,
		_w5403_,
		_w5404_
	);
	LUT4 #(
		.INIT('h0001)
	) name3504 (
		_w5388_,
		_w5393_,
		_w5398_,
		_w5404_,
		_w5405_
	);
	LUT2 #(
		.INIT('h7)
	) name3505 (
		_w5380_,
		_w5405_,
		_w5406_
	);
	LUT3 #(
		.INIT('hdc)
	) name3506 (
		_w3356_,
		_w3357_,
		_w3367_,
		_w5407_
	);
	LUT2 #(
		.INIT('h4)
	) name3507 (
		_w3359_,
		_w3361_,
		_w5408_
	);
	LUT4 #(
		.INIT('h000d)
	) name3508 (
		_w3354_,
		_w3355_,
		_w3359_,
		_w3360_,
		_w5409_
	);
	LUT4 #(
		.INIT('h7f00)
	) name3509 (
		\m6_s3_cyc_o_reg/NET0131 ,
		\rf_conf3_reg[12]/NET0131 ,
		\rf_conf3_reg[13]/NET0131 ,
		\s3_msel_arb3_state_reg[0]/NET0131 ,
		_w5410_
	);
	LUT4 #(
		.INIT('ha2f3)
	) name3510 (
		_w3355_,
		_w3356_,
		_w3357_,
		_w5410_,
		_w5411_
	);
	LUT4 #(
		.INIT('h0155)
	) name3511 (
		_w5407_,
		_w5408_,
		_w5409_,
		_w5411_,
		_w5412_
	);
	LUT2 #(
		.INIT('h8)
	) name3512 (
		_w3379_,
		_w5412_,
		_w5413_
	);
	LUT2 #(
		.INIT('h1)
	) name3513 (
		\s3_msel_arb3_state_reg[1]/NET0131 ,
		\s3_msel_arb3_state_reg[2]/NET0131 ,
		_w5414_
	);
	LUT3 #(
		.INIT('h20)
	) name3514 (
		_w3354_,
		_w3355_,
		_w5414_,
		_w5415_
	);
	LUT2 #(
		.INIT('h4)
	) name3515 (
		_w3356_,
		_w3367_,
		_w5416_
	);
	LUT4 #(
		.INIT('h1101)
	) name3516 (
		_w3356_,
		_w3359_,
		_w3360_,
		_w3361_,
		_w5417_
	);
	LUT3 #(
		.INIT('h10)
	) name3517 (
		_w3355_,
		_w3357_,
		_w5414_,
		_w5418_
	);
	LUT4 #(
		.INIT('h5455)
	) name3518 (
		_w5415_,
		_w5416_,
		_w5417_,
		_w5418_,
		_w5419_
	);
	LUT3 #(
		.INIT('h08)
	) name3519 (
		_w3353_,
		_w3359_,
		_w3367_,
		_w5420_
	);
	LUT3 #(
		.INIT('h0d)
	) name3520 (
		_w3354_,
		_w3355_,
		_w3360_,
		_w5421_
	);
	LUT3 #(
		.INIT('h04)
	) name3521 (
		_w3355_,
		_w3356_,
		_w3357_,
		_w5422_
	);
	LUT3 #(
		.INIT('h02)
	) name3522 (
		_w3353_,
		_w3361_,
		_w3367_,
		_w5423_
	);
	LUT4 #(
		.INIT('h0455)
	) name3523 (
		_w5420_,
		_w5421_,
		_w5422_,
		_w5423_,
		_w5424_
	);
	LUT3 #(
		.INIT('h40)
	) name3524 (
		\s3_msel_arb3_state_reg[0]/NET0131 ,
		_w5419_,
		_w5424_,
		_w5425_
	);
	LUT3 #(
		.INIT('h51)
	) name3525 (
		_w3361_,
		_w5421_,
		_w5422_,
		_w5426_
	);
	LUT4 #(
		.INIT('h0001)
	) name3526 (
		_w3355_,
		_w3357_,
		_w3361_,
		_w3367_,
		_w5427_
	);
	LUT2 #(
		.INIT('h1)
	) name3527 (
		_w3359_,
		_w5427_,
		_w5428_
	);
	LUT3 #(
		.INIT('h2a)
	) name3528 (
		\s3_msel_arb3_state_reg[0]/NET0131 ,
		_w3356_,
		_w3379_,
		_w5429_
	);
	LUT4 #(
		.INIT('h7500)
	) name3529 (
		_w3353_,
		_w5426_,
		_w5428_,
		_w5429_,
		_w5430_
	);
	LUT3 #(
		.INIT('h0b)
	) name3530 (
		_w5413_,
		_w5425_,
		_w5430_,
		_w5431_
	);
	LUT2 #(
		.INIT('h4)
	) name3531 (
		_w3354_,
		_w3357_,
		_w5432_
	);
	LUT4 #(
		.INIT('h5455)
	) name3532 (
		_w3354_,
		_w3355_,
		_w3367_,
		_w5410_,
		_w5433_
	);
	LUT4 #(
		.INIT('h010f)
	) name3533 (
		_w5416_,
		_w5417_,
		_w5432_,
		_w5433_,
		_w5434_
	);
	LUT3 #(
		.INIT('h02)
	) name3534 (
		\s3_msel_arb3_state_reg[0]/NET0131 ,
		\s3_msel_arb3_state_reg[1]/NET0131 ,
		\s3_msel_arb3_state_reg[2]/NET0131 ,
		_w5435_
	);
	LUT2 #(
		.INIT('h8)
	) name3535 (
		_w5434_,
		_w5435_,
		_w5436_
	);
	LUT2 #(
		.INIT('h1)
	) name3536 (
		_w3359_,
		_w5410_,
		_w5437_
	);
	LUT3 #(
		.INIT('h01)
	) name3537 (
		_w3355_,
		_w3357_,
		_w3367_,
		_w5438_
	);
	LUT4 #(
		.INIT('h2022)
	) name3538 (
		_w5421_,
		_w5422_,
		_w5437_,
		_w5438_,
		_w5439_
	);
	LUT4 #(
		.INIT('h0080)
	) name3539 (
		\m6_s3_cyc_o_reg/NET0131 ,
		\rf_conf3_reg[12]/NET0131 ,
		\rf_conf3_reg[13]/NET0131 ,
		\s3_msel_arb3_state_reg[0]/NET0131 ,
		_w5440_
	);
	LUT2 #(
		.INIT('h2)
	) name3540 (
		_w3365_,
		_w5440_,
		_w5441_
	);
	LUT3 #(
		.INIT('h10)
	) name3541 (
		_w3355_,
		_w3357_,
		_w5410_,
		_w5442_
	);
	LUT3 #(
		.INIT('h08)
	) name3542 (
		\s3_msel_arb3_state_reg[0]/NET0131 ,
		\s3_msel_arb3_state_reg[1]/NET0131 ,
		\s3_msel_arb3_state_reg[2]/NET0131 ,
		_w5443_
	);
	LUT3 #(
		.INIT('h10)
	) name3543 (
		_w3356_,
		_w3367_,
		_w5443_,
		_w5444_
	);
	LUT4 #(
		.INIT('hf100)
	) name3544 (
		_w5408_,
		_w5409_,
		_w5442_,
		_w5444_,
		_w5445_
	);
	LUT3 #(
		.INIT('h0b)
	) name3545 (
		_w5439_,
		_w5441_,
		_w5445_,
		_w5446_
	);
	LUT2 #(
		.INIT('h4)
	) name3546 (
		_w5436_,
		_w5446_,
		_w5447_
	);
	LUT2 #(
		.INIT('hb)
	) name3547 (
		_w5431_,
		_w5447_,
		_w5448_
	);
	LUT2 #(
		.INIT('h4)
	) name3548 (
		_w2501_,
		_w2509_,
		_w5449_
	);
	LUT3 #(
		.INIT('h04)
	) name3549 (
		_w2497_,
		_w2499_,
		_w2500_,
		_w5450_
	);
	LUT4 #(
		.INIT('hfd00)
	) name3550 (
		\m4_s4_cyc_o_reg/NET0131 ,
		\rf_conf4_reg[8]/NET0131 ,
		\rf_conf4_reg[9]/NET0131 ,
		\s4_msel_arb0_state_reg[0]/NET0131 ,
		_w5451_
	);
	LUT3 #(
		.INIT('h10)
	) name3551 (
		_w2500_,
		_w2502_,
		_w5451_,
		_w5452_
	);
	LUT3 #(
		.INIT('hf2)
	) name3552 (
		_w2496_,
		_w2497_,
		_w2504_,
		_w5453_
	);
	LUT4 #(
		.INIT('h000d)
	) name3553 (
		_w2496_,
		_w2497_,
		_w2501_,
		_w2504_,
		_w5454_
	);
	LUT4 #(
		.INIT('h5455)
	) name3554 (
		_w5449_,
		_w5450_,
		_w5452_,
		_w5454_,
		_w5455_
	);
	LUT2 #(
		.INIT('h8)
	) name3555 (
		_w2523_,
		_w5455_,
		_w5456_
	);
	LUT2 #(
		.INIT('h8)
	) name3556 (
		\s4_msel_arb0_state_reg[1]/NET0131 ,
		\s4_msel_arb0_state_reg[2]/NET0131 ,
		_w5457_
	);
	LUT2 #(
		.INIT('h2)
	) name3557 (
		_w2504_,
		_w2509_,
		_w5458_
	);
	LUT3 #(
		.INIT('h51)
	) name3558 (
		_w2501_,
		_w2504_,
		_w2509_,
		_w5459_
	);
	LUT4 #(
		.INIT('h2232)
	) name3559 (
		_w2501_,
		_w2502_,
		_w2504_,
		_w2509_,
		_w5460_
	);
	LUT2 #(
		.INIT('h1)
	) name3560 (
		_w2497_,
		_w2509_,
		_w5461_
	);
	LUT4 #(
		.INIT('h00fd)
	) name3561 (
		\m5_s4_cyc_o_reg/NET0131 ,
		\rf_conf4_reg[10]/NET0131 ,
		\rf_conf4_reg[11]/NET0131 ,
		\s4_msel_arb0_state_reg[0]/NET0131 ,
		_w5462_
	);
	LUT3 #(
		.INIT('h01)
	) name3562 (
		_w2497_,
		_w2509_,
		_w5462_,
		_w5463_
	);
	LUT2 #(
		.INIT('h4)
	) name3563 (
		_w2496_,
		_w2500_,
		_w5464_
	);
	LUT3 #(
		.INIT('h0b)
	) name3564 (
		_w2496_,
		_w2500_,
		_w2502_,
		_w5465_
	);
	LUT4 #(
		.INIT('h0111)
	) name3565 (
		_w2499_,
		_w5460_,
		_w5463_,
		_w5465_,
		_w5466_
	);
	LUT4 #(
		.INIT('h1101)
	) name3566 (
		_w2496_,
		_w2499_,
		_w2501_,
		_w2502_,
		_w5467_
	);
	LUT4 #(
		.INIT('hfd00)
	) name3567 (
		\m2_s4_cyc_o_reg/NET0131 ,
		\rf_conf4_reg[4]/NET0131 ,
		\rf_conf4_reg[5]/NET0131 ,
		\s4_msel_arb0_state_reg[0]/NET0131 ,
		_w5468_
	);
	LUT4 #(
		.INIT('h0e0f)
	) name3568 (
		_w2500_,
		_w2502_,
		_w2504_,
		_w5468_,
		_w5469_
	);
	LUT2 #(
		.INIT('h2)
	) name3569 (
		\s4_msel_arb0_state_reg[1]/NET0131 ,
		\s4_msel_arb0_state_reg[2]/NET0131 ,
		_w5470_
	);
	LUT3 #(
		.INIT('hd0)
	) name3570 (
		_w2497_,
		_w2504_,
		_w5470_,
		_w5471_
	);
	LUT4 #(
		.INIT('h1f00)
	) name3571 (
		_w5464_,
		_w5467_,
		_w5469_,
		_w5471_,
		_w5472_
	);
	LUT3 #(
		.INIT('h0d)
	) name3572 (
		_w5457_,
		_w5466_,
		_w5472_,
		_w5473_
	);
	LUT3 #(
		.INIT('h8a)
	) name3573 (
		\s4_msel_arb0_state_reg[0]/NET0131 ,
		_w5456_,
		_w5473_,
		_w5474_
	);
	LUT3 #(
		.INIT('h02)
	) name3574 (
		\s4_msel_arb0_state_reg[0]/NET0131 ,
		_w2500_,
		_w2502_,
		_w5475_
	);
	LUT4 #(
		.INIT('h55fd)
	) name3575 (
		_w5461_,
		_w5464_,
		_w5467_,
		_w5475_,
		_w5476_
	);
	LUT3 #(
		.INIT('h8c)
	) name3576 (
		_w5458_,
		_w5470_,
		_w5476_,
		_w5477_
	);
	LUT3 #(
		.INIT('h20)
	) name3577 (
		_w2499_,
		_w2500_,
		_w5457_,
		_w5478_
	);
	LUT3 #(
		.INIT('h10)
	) name3578 (
		_w2500_,
		_w2502_,
		_w5457_,
		_w5479_
	);
	LUT4 #(
		.INIT('h020f)
	) name3579 (
		_w5459_,
		_w5463_,
		_w5478_,
		_w5479_,
		_w5480_
	);
	LUT3 #(
		.INIT('h20)
	) name3580 (
		_w2501_,
		_w2502_,
		_w2523_,
		_w5481_
	);
	LUT2 #(
		.INIT('h1)
	) name3581 (
		_w2497_,
		_w2500_,
		_w5482_
	);
	LUT4 #(
		.INIT('h00fd)
	) name3582 (
		\m7_s4_cyc_o_reg/NET0131 ,
		\rf_conf4_reg[14]/NET0131 ,
		\rf_conf4_reg[15]/NET0131 ,
		\s4_msel_arb0_state_reg[0]/NET0131 ,
		_w5483_
	);
	LUT3 #(
		.INIT('h01)
	) name3583 (
		_w2497_,
		_w2500_,
		_w5483_,
		_w5484_
	);
	LUT3 #(
		.INIT('h10)
	) name3584 (
		_w2502_,
		_w2509_,
		_w2523_,
		_w5485_
	);
	LUT4 #(
		.INIT('h0133)
	) name3585 (
		_w5453_,
		_w5481_,
		_w5484_,
		_w5485_,
		_w5486_
	);
	LUT2 #(
		.INIT('h8)
	) name3586 (
		_w5480_,
		_w5486_,
		_w5487_
	);
	LUT3 #(
		.INIT('h02)
	) name3587 (
		\s4_msel_arb0_state_reg[0]/NET0131 ,
		_w2502_,
		_w2509_,
		_w5488_
	);
	LUT3 #(
		.INIT('h80)
	) name3588 (
		_w2526_,
		_w5482_,
		_w5488_,
		_w5489_
	);
	LUT3 #(
		.INIT('h04)
	) name3589 (
		_w2502_,
		_w2504_,
		_w2509_,
		_w5490_
	);
	LUT4 #(
		.INIT('h0002)
	) name3590 (
		\m4_s4_cyc_o_reg/NET0131 ,
		\rf_conf4_reg[8]/NET0131 ,
		\rf_conf4_reg[9]/NET0131 ,
		\s4_msel_arb0_state_reg[0]/NET0131 ,
		_w5491_
	);
	LUT4 #(
		.INIT('h00b0)
	) name3591 (
		_w2496_,
		_w2500_,
		_w2526_,
		_w5491_,
		_w5492_
	);
	LUT3 #(
		.INIT('hd0)
	) name3592 (
		_w5467_,
		_w5490_,
		_w5492_,
		_w5493_
	);
	LUT2 #(
		.INIT('h1)
	) name3593 (
		_w5489_,
		_w5493_,
		_w5494_
	);
	LUT4 #(
		.INIT('hba00)
	) name3594 (
		\s4_msel_arb0_state_reg[0]/NET0131 ,
		_w5477_,
		_w5487_,
		_w5494_,
		_w5495_
	);
	LUT2 #(
		.INIT('hb)
	) name3595 (
		_w5474_,
		_w5495_,
		_w5496_
	);
	LUT2 #(
		.INIT('h2)
	) name3596 (
		_w3779_,
		_w3784_,
		_w5497_
	);
	LUT4 #(
		.INIT('h000b)
	) name3597 (
		_w3776_,
		_w3777_,
		_w3780_,
		_w3784_,
		_w5498_
	);
	LUT2 #(
		.INIT('h1)
	) name3598 (
		\s4_msel_arb1_state_reg[1]/NET0131 ,
		\s4_msel_arb1_state_reg[2]/NET0131 ,
		_w5499_
	);
	LUT4 #(
		.INIT('h0d00)
	) name3599 (
		_w3788_,
		_w3789_,
		_w3794_,
		_w5499_,
		_w5500_
	);
	LUT4 #(
		.INIT('hab00)
	) name3600 (
		_w3789_,
		_w5497_,
		_w5498_,
		_w5500_,
		_w5501_
	);
	LUT2 #(
		.INIT('h2)
	) name3601 (
		\s4_msel_arb1_state_reg[1]/NET0131 ,
		\s4_msel_arb1_state_reg[2]/NET0131 ,
		_w5502_
	);
	LUT3 #(
		.INIT('h20)
	) name3602 (
		_w3784_,
		_w3788_,
		_w5502_,
		_w5503_
	);
	LUT3 #(
		.INIT('h0b)
	) name3603 (
		_w3776_,
		_w3777_,
		_w3780_,
		_w5504_
	);
	LUT2 #(
		.INIT('h1)
	) name3604 (
		_w3776_,
		_w3794_,
		_w5505_
	);
	LUT4 #(
		.INIT('h00f7)
	) name3605 (
		\m1_s4_cyc_o_reg/NET0131 ,
		\rf_conf4_reg[2]/NET0131 ,
		\rf_conf4_reg[3]/NET0131 ,
		\s4_msel_arb1_state_reg[0]/NET0131 ,
		_w5506_
	);
	LUT3 #(
		.INIT('h01)
	) name3606 (
		_w3776_,
		_w3794_,
		_w5506_,
		_w5507_
	);
	LUT3 #(
		.INIT('h10)
	) name3607 (
		_w3779_,
		_w3788_,
		_w5502_,
		_w5508_
	);
	LUT4 #(
		.INIT('h0455)
	) name3608 (
		_w5503_,
		_w5504_,
		_w5507_,
		_w5508_,
		_w5509_
	);
	LUT2 #(
		.INIT('h4)
	) name3609 (
		_w3779_,
		_w3782_,
		_w5510_
	);
	LUT3 #(
		.INIT('h0d)
	) name3610 (
		_w3784_,
		_w3788_,
		_w3789_,
		_w5511_
	);
	LUT4 #(
		.INIT('haf2f)
	) name3611 (
		_w5504_,
		_w5505_,
		_w5510_,
		_w5511_,
		_w5512_
	);
	LUT4 #(
		.INIT('h4555)
	) name3612 (
		\s4_msel_arb1_state_reg[0]/NET0131 ,
		_w5501_,
		_w5509_,
		_w5512_,
		_w5513_
	);
	LUT4 #(
		.INIT('hf700)
	) name3613 (
		\m0_s4_cyc_o_reg/NET0131 ,
		\rf_conf4_reg[0]/NET0131 ,
		\rf_conf4_reg[1]/NET0131 ,
		\s4_msel_arb1_state_reg[0]/NET0131 ,
		_w5514_
	);
	LUT3 #(
		.INIT('h01)
	) name3614 (
		_w3776_,
		_w3779_,
		_w3788_,
		_w5515_
	);
	LUT4 #(
		.INIT('h0100)
	) name3615 (
		_w3776_,
		_w3779_,
		_w3788_,
		_w5514_,
		_w5516_
	);
	LUT4 #(
		.INIT('h0008)
	) name3616 (
		\m6_s4_cyc_o_reg/NET0131 ,
		\rf_conf4_reg[12]/NET0131 ,
		\rf_conf4_reg[13]/NET0131 ,
		\s4_msel_arb1_state_reg[0]/NET0131 ,
		_w5517_
	);
	LUT2 #(
		.INIT('h2)
	) name3617 (
		_w3777_,
		_w5517_,
		_w5518_
	);
	LUT3 #(
		.INIT('h04)
	) name3618 (
		_w3779_,
		_w3780_,
		_w3788_,
		_w5519_
	);
	LUT2 #(
		.INIT('h1)
	) name3619 (
		_w3794_,
		_w5517_,
		_w5520_
	);
	LUT4 #(
		.INIT('h0233)
	) name3620 (
		_w5511_,
		_w5518_,
		_w5519_,
		_w5520_,
		_w5521_
	);
	LUT2 #(
		.INIT('h8)
	) name3621 (
		\s4_msel_arb1_state_reg[1]/NET0131 ,
		\s4_msel_arb1_state_reg[2]/NET0131 ,
		_w5522_
	);
	LUT3 #(
		.INIT('hb0)
	) name3622 (
		_w5516_,
		_w5521_,
		_w5522_,
		_w5523_
	);
	LUT3 #(
		.INIT('h20)
	) name3623 (
		\s4_msel_arb1_state_reg[0]/NET0131 ,
		\s4_msel_arb1_state_reg[1]/NET0131 ,
		\s4_msel_arb1_state_reg[2]/NET0131 ,
		_w5524_
	);
	LUT4 #(
		.INIT('h00a2)
	) name3624 (
		_w5504_,
		_w5505_,
		_w5511_,
		_w5516_,
		_w5525_
	);
	LUT2 #(
		.INIT('h2)
	) name3625 (
		_w5524_,
		_w5525_,
		_w5526_
	);
	LUT2 #(
		.INIT('h1)
	) name3626 (
		_w3777_,
		_w5514_,
		_w5527_
	);
	LUT4 #(
		.INIT('h0a02)
	) name3627 (
		_w5511_,
		_w5515_,
		_w5519_,
		_w5527_,
		_w5528_
	);
	LUT3 #(
		.INIT('h02)
	) name3628 (
		\s4_msel_arb1_state_reg[0]/NET0131 ,
		\s4_msel_arb1_state_reg[1]/NET0131 ,
		\s4_msel_arb1_state_reg[2]/NET0131 ,
		_w5529_
	);
	LUT3 #(
		.INIT('h51)
	) name3629 (
		_w3779_,
		_w3788_,
		_w3789_,
		_w5530_
	);
	LUT4 #(
		.INIT('h0eee)
	) name3630 (
		_w5497_,
		_w5498_,
		_w5507_,
		_w5530_,
		_w5531_
	);
	LUT3 #(
		.INIT('h08)
	) name3631 (
		\s4_msel_arb1_state_reg[0]/NET0131 ,
		\s4_msel_arb1_state_reg[1]/NET0131 ,
		\s4_msel_arb1_state_reg[2]/NET0131 ,
		_w5532_
	);
	LUT4 #(
		.INIT('hb0bb)
	) name3632 (
		_w5528_,
		_w5529_,
		_w5531_,
		_w5532_,
		_w5533_
	);
	LUT4 #(
		.INIT('hfeff)
	) name3633 (
		_w5513_,
		_w5523_,
		_w5526_,
		_w5533_,
		_w5534_
	);
	LUT3 #(
		.INIT('h20)
	) name3634 (
		\m4_s4_cyc_o_reg/NET0131 ,
		\rf_conf4_reg[8]/NET0131 ,
		\rf_conf4_reg[9]/NET0131 ,
		_w5535_
	);
	LUT3 #(
		.INIT('h20)
	) name3635 (
		\m7_s4_cyc_o_reg/NET0131 ,
		\rf_conf4_reg[14]/NET0131 ,
		\rf_conf4_reg[15]/NET0131 ,
		_w5536_
	);
	LUT3 #(
		.INIT('h20)
	) name3636 (
		\m0_s4_cyc_o_reg/NET0131 ,
		\rf_conf4_reg[0]/NET0131 ,
		\rf_conf4_reg[1]/NET0131 ,
		_w5537_
	);
	LUT2 #(
		.INIT('h4)
	) name3637 (
		_w5536_,
		_w5537_,
		_w5538_
	);
	LUT3 #(
		.INIT('h20)
	) name3638 (
		\m3_s4_cyc_o_reg/NET0131 ,
		\rf_conf4_reg[6]/NET0131 ,
		\rf_conf4_reg[7]/NET0131 ,
		_w5539_
	);
	LUT3 #(
		.INIT('h20)
	) name3639 (
		\m2_s4_cyc_o_reg/NET0131 ,
		\rf_conf4_reg[4]/NET0131 ,
		\rf_conf4_reg[5]/NET0131 ,
		_w5540_
	);
	LUT3 #(
		.INIT('h20)
	) name3640 (
		\m1_s4_cyc_o_reg/NET0131 ,
		\rf_conf4_reg[2]/NET0131 ,
		\rf_conf4_reg[3]/NET0131 ,
		_w5541_
	);
	LUT4 #(
		.INIT('h0051)
	) name3641 (
		_w5536_,
		_w5539_,
		_w5540_,
		_w5541_,
		_w5542_
	);
	LUT3 #(
		.INIT('h20)
	) name3642 (
		\m5_s4_cyc_o_reg/NET0131 ,
		\rf_conf4_reg[10]/NET0131 ,
		\rf_conf4_reg[11]/NET0131 ,
		_w5543_
	);
	LUT3 #(
		.INIT('h20)
	) name3643 (
		\m6_s4_cyc_o_reg/NET0131 ,
		\rf_conf4_reg[12]/NET0131 ,
		\rf_conf4_reg[13]/NET0131 ,
		_w5544_
	);
	LUT3 #(
		.INIT('h8a)
	) name3644 (
		\s4_msel_arb2_state_reg[0]/NET0131 ,
		_w5543_,
		_w5544_,
		_w5545_
	);
	LUT4 #(
		.INIT('hf100)
	) name3645 (
		_w5538_,
		_w5542_,
		_w5543_,
		_w5545_,
		_w5546_
	);
	LUT2 #(
		.INIT('h1)
	) name3646 (
		_w5537_,
		_w5544_,
		_w5547_
	);
	LUT4 #(
		.INIT('hdf00)
	) name3647 (
		\m2_s4_cyc_o_reg/NET0131 ,
		\rf_conf4_reg[4]/NET0131 ,
		\rf_conf4_reg[5]/NET0131 ,
		\s4_msel_arb2_state_reg[0]/NET0131 ,
		_w5548_
	);
	LUT4 #(
		.INIT('h3030)
	) name3648 (
		_w5537_,
		_w5543_,
		_w5544_,
		_w5548_,
		_w5549_
	);
	LUT4 #(
		.INIT('h3233)
	) name3649 (
		_w5537_,
		_w5543_,
		_w5544_,
		_w5548_,
		_w5550_
	);
	LUT4 #(
		.INIT('h010f)
	) name3650 (
		_w5538_,
		_w5542_,
		_w5549_,
		_w5550_,
		_w5551_
	);
	LUT2 #(
		.INIT('h4)
	) name3651 (
		\s4_msel_arb2_state_reg[1]/NET0131 ,
		\s4_msel_arb2_state_reg[2]/NET0131 ,
		_w5552_
	);
	LUT4 #(
		.INIT('hd000)
	) name3652 (
		_w5535_,
		_w5546_,
		_w5551_,
		_w5552_,
		_w5553_
	);
	LUT2 #(
		.INIT('h8)
	) name3653 (
		\s4_msel_arb2_state_reg[1]/NET0131 ,
		\s4_msel_arb2_state_reg[2]/NET0131 ,
		_w5554_
	);
	LUT3 #(
		.INIT('h20)
	) name3654 (
		_w5536_,
		_w5544_,
		_w5554_,
		_w5555_
	);
	LUT3 #(
		.INIT('h0d)
	) name3655 (
		_w5539_,
		_w5540_,
		_w5541_,
		_w5556_
	);
	LUT4 #(
		.INIT('h00df)
	) name3656 (
		\m5_s4_cyc_o_reg/NET0131 ,
		\rf_conf4_reg[10]/NET0131 ,
		\rf_conf4_reg[11]/NET0131 ,
		\s4_msel_arb2_state_reg[0]/NET0131 ,
		_w5557_
	);
	LUT3 #(
		.INIT('h01)
	) name3657 (
		_w5535_,
		_w5540_,
		_w5557_,
		_w5558_
	);
	LUT3 #(
		.INIT('h10)
	) name3658 (
		_w5537_,
		_w5544_,
		_w5554_,
		_w5559_
	);
	LUT4 #(
		.INIT('h0455)
	) name3659 (
		_w5555_,
		_w5556_,
		_w5558_,
		_w5559_,
		_w5560_
	);
	LUT2 #(
		.INIT('h1)
	) name3660 (
		\s4_msel_arb2_state_reg[1]/NET0131 ,
		\s4_msel_arb2_state_reg[2]/NET0131 ,
		_w5561_
	);
	LUT3 #(
		.INIT('h40)
	) name3661 (
		_w5537_,
		_w5541_,
		_w5561_,
		_w5562_
	);
	LUT2 #(
		.INIT('h2)
	) name3662 (
		_w5535_,
		_w5539_,
		_w5563_
	);
	LUT4 #(
		.INIT('h0301)
	) name3663 (
		_w5536_,
		_w5539_,
		_w5543_,
		_w5544_,
		_w5564_
	);
	LUT3 #(
		.INIT('h10)
	) name3664 (
		_w5537_,
		_w5540_,
		_w5561_,
		_w5565_
	);
	LUT4 #(
		.INIT('h5455)
	) name3665 (
		_w5562_,
		_w5563_,
		_w5564_,
		_w5565_,
		_w5566_
	);
	LUT3 #(
		.INIT('h15)
	) name3666 (
		\s4_msel_arb2_state_reg[0]/NET0131 ,
		_w5560_,
		_w5566_,
		_w5567_
	);
	LUT3 #(
		.INIT('h80)
	) name3667 (
		\s4_msel_arb2_state_reg[0]/NET0131 ,
		_w5541_,
		_w5561_,
		_w5568_
	);
	LUT3 #(
		.INIT('h45)
	) name3668 (
		_w5537_,
		_w5543_,
		_w5544_,
		_w5569_
	);
	LUT4 #(
		.INIT('h0eee)
	) name3669 (
		_w5538_,
		_w5542_,
		_w5558_,
		_w5569_,
		_w5570_
	);
	LUT3 #(
		.INIT('h80)
	) name3670 (
		\s4_msel_arb2_state_reg[0]/NET0131 ,
		\s4_msel_arb2_state_reg[1]/NET0131 ,
		\s4_msel_arb2_state_reg[2]/NET0131 ,
		_w5571_
	);
	LUT3 #(
		.INIT('h45)
	) name3671 (
		_w5568_,
		_w5570_,
		_w5571_,
		_w5572_
	);
	LUT3 #(
		.INIT('h40)
	) name3672 (
		_w5541_,
		_w5548_,
		_w5561_,
		_w5573_
	);
	LUT4 #(
		.INIT('h0020)
	) name3673 (
		\m2_s4_cyc_o_reg/NET0131 ,
		\rf_conf4_reg[4]/NET0131 ,
		\rf_conf4_reg[5]/NET0131 ,
		\s4_msel_arb2_state_reg[0]/NET0131 ,
		_w5574_
	);
	LUT2 #(
		.INIT('h2)
	) name3674 (
		\s4_msel_arb2_state_reg[1]/NET0131 ,
		\s4_msel_arb2_state_reg[2]/NET0131 ,
		_w5575_
	);
	LUT2 #(
		.INIT('h4)
	) name3675 (
		_w5574_,
		_w5575_,
		_w5576_
	);
	LUT4 #(
		.INIT('h1110)
	) name3676 (
		_w5563_,
		_w5564_,
		_w5573_,
		_w5576_,
		_w5577_
	);
	LUT3 #(
		.INIT('h40)
	) name3677 (
		_w5535_,
		_w5547_,
		_w5573_,
		_w5578_
	);
	LUT4 #(
		.INIT('hfafb)
	) name3678 (
		_w5537_,
		_w5541_,
		_w5544_,
		_w5548_,
		_w5579_
	);
	LUT3 #(
		.INIT('h10)
	) name3679 (
		_w5535_,
		_w5574_,
		_w5575_,
		_w5580_
	);
	LUT2 #(
		.INIT('h4)
	) name3680 (
		_w5579_,
		_w5580_,
		_w5581_
	);
	LUT3 #(
		.INIT('h01)
	) name3681 (
		_w5577_,
		_w5578_,
		_w5581_,
		_w5582_
	);
	LUT4 #(
		.INIT('hefff)
	) name3682 (
		_w5553_,
		_w5567_,
		_w5572_,
		_w5582_,
		_w5583_
	);
	LUT3 #(
		.INIT('hdc)
	) name3683 (
		_w3058_,
		_w3059_,
		_w3069_,
		_w5584_
	);
	LUT2 #(
		.INIT('h4)
	) name3684 (
		_w3061_,
		_w3063_,
		_w5585_
	);
	LUT4 #(
		.INIT('h000d)
	) name3685 (
		_w3056_,
		_w3057_,
		_w3061_,
		_w3062_,
		_w5586_
	);
	LUT4 #(
		.INIT('h7f00)
	) name3686 (
		\m6_s4_cyc_o_reg/NET0131 ,
		\rf_conf4_reg[12]/NET0131 ,
		\rf_conf4_reg[13]/NET0131 ,
		\s4_msel_arb3_state_reg[0]/NET0131 ,
		_w5587_
	);
	LUT4 #(
		.INIT('ha2f3)
	) name3687 (
		_w3057_,
		_w3058_,
		_w3059_,
		_w5587_,
		_w5588_
	);
	LUT4 #(
		.INIT('h0155)
	) name3688 (
		_w5584_,
		_w5585_,
		_w5586_,
		_w5588_,
		_w5589_
	);
	LUT2 #(
		.INIT('h8)
	) name3689 (
		_w3081_,
		_w5589_,
		_w5590_
	);
	LUT2 #(
		.INIT('h1)
	) name3690 (
		\s4_msel_arb3_state_reg[1]/NET0131 ,
		\s4_msel_arb3_state_reg[2]/NET0131 ,
		_w5591_
	);
	LUT3 #(
		.INIT('h20)
	) name3691 (
		_w3056_,
		_w3057_,
		_w5591_,
		_w5592_
	);
	LUT2 #(
		.INIT('h4)
	) name3692 (
		_w3058_,
		_w3069_,
		_w5593_
	);
	LUT4 #(
		.INIT('h1101)
	) name3693 (
		_w3058_,
		_w3061_,
		_w3062_,
		_w3063_,
		_w5594_
	);
	LUT3 #(
		.INIT('h10)
	) name3694 (
		_w3057_,
		_w3059_,
		_w5591_,
		_w5595_
	);
	LUT4 #(
		.INIT('h5455)
	) name3695 (
		_w5592_,
		_w5593_,
		_w5594_,
		_w5595_,
		_w5596_
	);
	LUT3 #(
		.INIT('h08)
	) name3696 (
		_w3055_,
		_w3061_,
		_w3069_,
		_w5597_
	);
	LUT3 #(
		.INIT('h0d)
	) name3697 (
		_w3056_,
		_w3057_,
		_w3062_,
		_w5598_
	);
	LUT3 #(
		.INIT('h04)
	) name3698 (
		_w3057_,
		_w3058_,
		_w3059_,
		_w5599_
	);
	LUT3 #(
		.INIT('h02)
	) name3699 (
		_w3055_,
		_w3063_,
		_w3069_,
		_w5600_
	);
	LUT4 #(
		.INIT('h0455)
	) name3700 (
		_w5597_,
		_w5598_,
		_w5599_,
		_w5600_,
		_w5601_
	);
	LUT3 #(
		.INIT('h40)
	) name3701 (
		\s4_msel_arb3_state_reg[0]/NET0131 ,
		_w5596_,
		_w5601_,
		_w5602_
	);
	LUT3 #(
		.INIT('h51)
	) name3702 (
		_w3063_,
		_w5598_,
		_w5599_,
		_w5603_
	);
	LUT4 #(
		.INIT('h0001)
	) name3703 (
		_w3057_,
		_w3059_,
		_w3063_,
		_w3069_,
		_w5604_
	);
	LUT2 #(
		.INIT('h1)
	) name3704 (
		_w3061_,
		_w5604_,
		_w5605_
	);
	LUT3 #(
		.INIT('h2a)
	) name3705 (
		\s4_msel_arb3_state_reg[0]/NET0131 ,
		_w3058_,
		_w3081_,
		_w5606_
	);
	LUT4 #(
		.INIT('h7500)
	) name3706 (
		_w3055_,
		_w5603_,
		_w5605_,
		_w5606_,
		_w5607_
	);
	LUT3 #(
		.INIT('h0b)
	) name3707 (
		_w5590_,
		_w5602_,
		_w5607_,
		_w5608_
	);
	LUT2 #(
		.INIT('h4)
	) name3708 (
		_w3056_,
		_w3059_,
		_w5609_
	);
	LUT4 #(
		.INIT('h5455)
	) name3709 (
		_w3056_,
		_w3057_,
		_w3069_,
		_w5587_,
		_w5610_
	);
	LUT4 #(
		.INIT('h010f)
	) name3710 (
		_w5593_,
		_w5594_,
		_w5609_,
		_w5610_,
		_w5611_
	);
	LUT3 #(
		.INIT('h02)
	) name3711 (
		\s4_msel_arb3_state_reg[0]/NET0131 ,
		\s4_msel_arb3_state_reg[1]/NET0131 ,
		\s4_msel_arb3_state_reg[2]/NET0131 ,
		_w5612_
	);
	LUT2 #(
		.INIT('h8)
	) name3712 (
		_w5611_,
		_w5612_,
		_w5613_
	);
	LUT2 #(
		.INIT('h1)
	) name3713 (
		_w3061_,
		_w5587_,
		_w5614_
	);
	LUT3 #(
		.INIT('h01)
	) name3714 (
		_w3057_,
		_w3059_,
		_w3069_,
		_w5615_
	);
	LUT4 #(
		.INIT('h2022)
	) name3715 (
		_w5598_,
		_w5599_,
		_w5614_,
		_w5615_,
		_w5616_
	);
	LUT4 #(
		.INIT('h0080)
	) name3716 (
		\m6_s4_cyc_o_reg/NET0131 ,
		\rf_conf4_reg[12]/NET0131 ,
		\rf_conf4_reg[13]/NET0131 ,
		\s4_msel_arb3_state_reg[0]/NET0131 ,
		_w5617_
	);
	LUT2 #(
		.INIT('h2)
	) name3717 (
		_w3067_,
		_w5617_,
		_w5618_
	);
	LUT3 #(
		.INIT('h10)
	) name3718 (
		_w3057_,
		_w3059_,
		_w5587_,
		_w5619_
	);
	LUT3 #(
		.INIT('h08)
	) name3719 (
		\s4_msel_arb3_state_reg[0]/NET0131 ,
		\s4_msel_arb3_state_reg[1]/NET0131 ,
		\s4_msel_arb3_state_reg[2]/NET0131 ,
		_w5620_
	);
	LUT3 #(
		.INIT('h10)
	) name3720 (
		_w3058_,
		_w3069_,
		_w5620_,
		_w5621_
	);
	LUT4 #(
		.INIT('hf100)
	) name3721 (
		_w5585_,
		_w5586_,
		_w5619_,
		_w5621_,
		_w5622_
	);
	LUT3 #(
		.INIT('h0b)
	) name3722 (
		_w5616_,
		_w5618_,
		_w5622_,
		_w5623_
	);
	LUT2 #(
		.INIT('h4)
	) name3723 (
		_w5613_,
		_w5623_,
		_w5624_
	);
	LUT2 #(
		.INIT('hb)
	) name3724 (
		_w5608_,
		_w5624_,
		_w5625_
	);
	LUT2 #(
		.INIT('h4)
	) name3725 (
		_w2538_,
		_w2546_,
		_w5626_
	);
	LUT3 #(
		.INIT('h04)
	) name3726 (
		_w2534_,
		_w2536_,
		_w2537_,
		_w5627_
	);
	LUT4 #(
		.INIT('hfd00)
	) name3727 (
		\m4_s5_cyc_o_reg/NET0131 ,
		\rf_conf5_reg[8]/NET0131 ,
		\rf_conf5_reg[9]/NET0131 ,
		\s5_msel_arb0_state_reg[0]/NET0131 ,
		_w5628_
	);
	LUT3 #(
		.INIT('h10)
	) name3728 (
		_w2537_,
		_w2539_,
		_w5628_,
		_w5629_
	);
	LUT3 #(
		.INIT('hf2)
	) name3729 (
		_w2533_,
		_w2534_,
		_w2541_,
		_w5630_
	);
	LUT4 #(
		.INIT('h000d)
	) name3730 (
		_w2533_,
		_w2534_,
		_w2538_,
		_w2541_,
		_w5631_
	);
	LUT4 #(
		.INIT('h5455)
	) name3731 (
		_w5626_,
		_w5627_,
		_w5629_,
		_w5631_,
		_w5632_
	);
	LUT2 #(
		.INIT('h8)
	) name3732 (
		_w2560_,
		_w5632_,
		_w5633_
	);
	LUT2 #(
		.INIT('h8)
	) name3733 (
		\s5_msel_arb0_state_reg[1]/NET0131 ,
		\s5_msel_arb0_state_reg[2]/NET0131 ,
		_w5634_
	);
	LUT2 #(
		.INIT('h2)
	) name3734 (
		_w2541_,
		_w2546_,
		_w5635_
	);
	LUT3 #(
		.INIT('h51)
	) name3735 (
		_w2538_,
		_w2541_,
		_w2546_,
		_w5636_
	);
	LUT4 #(
		.INIT('h2232)
	) name3736 (
		_w2538_,
		_w2539_,
		_w2541_,
		_w2546_,
		_w5637_
	);
	LUT2 #(
		.INIT('h1)
	) name3737 (
		_w2534_,
		_w2546_,
		_w5638_
	);
	LUT4 #(
		.INIT('h00fd)
	) name3738 (
		\m5_s5_cyc_o_reg/NET0131 ,
		\rf_conf5_reg[10]/NET0131 ,
		\rf_conf5_reg[11]/NET0131 ,
		\s5_msel_arb0_state_reg[0]/NET0131 ,
		_w5639_
	);
	LUT3 #(
		.INIT('h01)
	) name3739 (
		_w2534_,
		_w2546_,
		_w5639_,
		_w5640_
	);
	LUT2 #(
		.INIT('h4)
	) name3740 (
		_w2533_,
		_w2537_,
		_w5641_
	);
	LUT3 #(
		.INIT('h0b)
	) name3741 (
		_w2533_,
		_w2537_,
		_w2539_,
		_w5642_
	);
	LUT4 #(
		.INIT('h0111)
	) name3742 (
		_w2536_,
		_w5637_,
		_w5640_,
		_w5642_,
		_w5643_
	);
	LUT4 #(
		.INIT('h1101)
	) name3743 (
		_w2533_,
		_w2536_,
		_w2538_,
		_w2539_,
		_w5644_
	);
	LUT4 #(
		.INIT('hfd00)
	) name3744 (
		\m2_s5_cyc_o_reg/NET0131 ,
		\rf_conf5_reg[4]/NET0131 ,
		\rf_conf5_reg[5]/NET0131 ,
		\s5_msel_arb0_state_reg[0]/NET0131 ,
		_w5645_
	);
	LUT4 #(
		.INIT('h0e0f)
	) name3745 (
		_w2537_,
		_w2539_,
		_w2541_,
		_w5645_,
		_w5646_
	);
	LUT2 #(
		.INIT('h2)
	) name3746 (
		\s5_msel_arb0_state_reg[1]/NET0131 ,
		\s5_msel_arb0_state_reg[2]/NET0131 ,
		_w5647_
	);
	LUT3 #(
		.INIT('hd0)
	) name3747 (
		_w2534_,
		_w2541_,
		_w5647_,
		_w5648_
	);
	LUT4 #(
		.INIT('h1f00)
	) name3748 (
		_w5641_,
		_w5644_,
		_w5646_,
		_w5648_,
		_w5649_
	);
	LUT3 #(
		.INIT('h0d)
	) name3749 (
		_w5634_,
		_w5643_,
		_w5649_,
		_w5650_
	);
	LUT3 #(
		.INIT('h8a)
	) name3750 (
		\s5_msel_arb0_state_reg[0]/NET0131 ,
		_w5633_,
		_w5650_,
		_w5651_
	);
	LUT3 #(
		.INIT('h02)
	) name3751 (
		\s5_msel_arb0_state_reg[0]/NET0131 ,
		_w2537_,
		_w2539_,
		_w5652_
	);
	LUT4 #(
		.INIT('h55fd)
	) name3752 (
		_w5638_,
		_w5641_,
		_w5644_,
		_w5652_,
		_w5653_
	);
	LUT3 #(
		.INIT('h8c)
	) name3753 (
		_w5635_,
		_w5647_,
		_w5653_,
		_w5654_
	);
	LUT3 #(
		.INIT('h20)
	) name3754 (
		_w2536_,
		_w2537_,
		_w5634_,
		_w5655_
	);
	LUT3 #(
		.INIT('h10)
	) name3755 (
		_w2537_,
		_w2539_,
		_w5634_,
		_w5656_
	);
	LUT4 #(
		.INIT('h020f)
	) name3756 (
		_w5636_,
		_w5640_,
		_w5655_,
		_w5656_,
		_w5657_
	);
	LUT3 #(
		.INIT('h20)
	) name3757 (
		_w2538_,
		_w2539_,
		_w2560_,
		_w5658_
	);
	LUT2 #(
		.INIT('h1)
	) name3758 (
		_w2534_,
		_w2537_,
		_w5659_
	);
	LUT4 #(
		.INIT('h00fd)
	) name3759 (
		\m7_s5_cyc_o_reg/NET0131 ,
		\rf_conf5_reg[14]/NET0131 ,
		\rf_conf5_reg[15]/NET0131 ,
		\s5_msel_arb0_state_reg[0]/NET0131 ,
		_w5660_
	);
	LUT3 #(
		.INIT('h01)
	) name3760 (
		_w2534_,
		_w2537_,
		_w5660_,
		_w5661_
	);
	LUT3 #(
		.INIT('h10)
	) name3761 (
		_w2539_,
		_w2546_,
		_w2560_,
		_w5662_
	);
	LUT4 #(
		.INIT('h0133)
	) name3762 (
		_w5630_,
		_w5658_,
		_w5661_,
		_w5662_,
		_w5663_
	);
	LUT2 #(
		.INIT('h8)
	) name3763 (
		_w5657_,
		_w5663_,
		_w5664_
	);
	LUT3 #(
		.INIT('h02)
	) name3764 (
		\s5_msel_arb0_state_reg[0]/NET0131 ,
		_w2539_,
		_w2546_,
		_w5665_
	);
	LUT3 #(
		.INIT('h80)
	) name3765 (
		_w2563_,
		_w5659_,
		_w5665_,
		_w5666_
	);
	LUT3 #(
		.INIT('h04)
	) name3766 (
		_w2539_,
		_w2541_,
		_w2546_,
		_w5667_
	);
	LUT4 #(
		.INIT('h0002)
	) name3767 (
		\m4_s5_cyc_o_reg/NET0131 ,
		\rf_conf5_reg[8]/NET0131 ,
		\rf_conf5_reg[9]/NET0131 ,
		\s5_msel_arb0_state_reg[0]/NET0131 ,
		_w5668_
	);
	LUT4 #(
		.INIT('h00b0)
	) name3768 (
		_w2533_,
		_w2537_,
		_w2563_,
		_w5668_,
		_w5669_
	);
	LUT3 #(
		.INIT('hd0)
	) name3769 (
		_w5644_,
		_w5667_,
		_w5669_,
		_w5670_
	);
	LUT2 #(
		.INIT('h1)
	) name3770 (
		_w5666_,
		_w5670_,
		_w5671_
	);
	LUT4 #(
		.INIT('hba00)
	) name3771 (
		\s5_msel_arb0_state_reg[0]/NET0131 ,
		_w5654_,
		_w5664_,
		_w5671_,
		_w5672_
	);
	LUT2 #(
		.INIT('hb)
	) name3772 (
		_w5651_,
		_w5672_,
		_w5673_
	);
	LUT3 #(
		.INIT('hf2)
	) name3773 (
		_w3808_,
		_w3809_,
		_w3812_,
		_w5674_
	);
	LUT4 #(
		.INIT('h0008)
	) name3774 (
		\m4_s5_cyc_o_reg/NET0131 ,
		\rf_conf5_reg[8]/NET0131 ,
		\rf_conf5_reg[9]/NET0131 ,
		\s5_msel_arb1_state_reg[0]/NET0131 ,
		_w5675_
	);
	LUT2 #(
		.INIT('h4)
	) name3775 (
		_w5675_,
		_w3818_,
		_w5676_
	);
	LUT2 #(
		.INIT('h8)
	) name3776 (
		_w5674_,
		_w5676_,
		_w5677_
	);
	LUT3 #(
		.INIT('hf2)
	) name3777 (
		_w3802_,
		_w3803_,
		_w3806_,
		_w5678_
	);
	LUT3 #(
		.INIT('h02)
	) name3778 (
		\s5_msel_arb1_state_reg[0]/NET0131 ,
		_w3803_,
		_w3811_,
		_w5679_
	);
	LUT2 #(
		.INIT('h1)
	) name3779 (
		_w3805_,
		_w3809_,
		_w5680_
	);
	LUT4 #(
		.INIT('h0100)
	) name3780 (
		_w3805_,
		_w3809_,
		_w5675_,
		_w3818_,
		_w5681_
	);
	LUT3 #(
		.INIT('he0)
	) name3781 (
		_w5678_,
		_w5679_,
		_w5681_,
		_w5682_
	);
	LUT4 #(
		.INIT('h0031)
	) name3782 (
		_w3803_,
		_w3805_,
		_w3806_,
		_w3809_,
		_w5683_
	);
	LUT4 #(
		.INIT('h4445)
	) name3783 (
		_w3802_,
		_w3811_,
		_w5674_,
		_w5683_,
		_w5684_
	);
	LUT3 #(
		.INIT('h08)
	) name3784 (
		\s5_msel_arb1_state_reg[0]/NET0131 ,
		\s5_msel_arb1_state_reg[1]/NET0131 ,
		\s5_msel_arb1_state_reg[2]/NET0131 ,
		_w5685_
	);
	LUT4 #(
		.INIT('h0001)
	) name3785 (
		_w3802_,
		_w3806_,
		_w3808_,
		_w3812_,
		_w5686_
	);
	LUT2 #(
		.INIT('h4)
	) name3786 (
		_w3803_,
		_w3821_,
		_w5687_
	);
	LUT3 #(
		.INIT('h45)
	) name3787 (
		_w5685_,
		_w5686_,
		_w5687_,
		_w5688_
	);
	LUT4 #(
		.INIT('h1110)
	) name3788 (
		_w5677_,
		_w5682_,
		_w5684_,
		_w5688_,
		_w5689_
	);
	LUT4 #(
		.INIT('h0008)
	) name3789 (
		\m0_s5_cyc_o_reg/NET0131 ,
		\rf_conf5_reg[0]/NET0131 ,
		\rf_conf5_reg[1]/NET0131 ,
		\s5_msel_arb1_state_reg[0]/NET0131 ,
		_w5690_
	);
	LUT4 #(
		.INIT('h00f2)
	) name3790 (
		_w3802_,
		_w3803_,
		_w3806_,
		_w5690_,
		_w5691_
	);
	LUT3 #(
		.INIT('h01)
	) name3791 (
		_w3803_,
		_w3811_,
		_w5690_,
		_w5692_
	);
	LUT3 #(
		.INIT('h13)
	) name3792 (
		_w5674_,
		_w5691_,
		_w5692_,
		_w5693_
	);
	LUT2 #(
		.INIT('h8)
	) name3793 (
		_w5679_,
		_w5680_,
		_w5694_
	);
	LUT3 #(
		.INIT('ha2)
	) name3794 (
		_w3814_,
		_w5693_,
		_w5694_,
		_w5695_
	);
	LUT3 #(
		.INIT('h10)
	) name3795 (
		_w3803_,
		_w3811_,
		_w3812_,
		_w5696_
	);
	LUT3 #(
		.INIT('h54)
	) name3796 (
		_w3805_,
		_w5678_,
		_w5696_,
		_w5697_
	);
	LUT3 #(
		.INIT('h15)
	) name3797 (
		_w3808_,
		_w5679_,
		_w5680_,
		_w5698_
	);
	LUT4 #(
		.INIT('h0008)
	) name3798 (
		\m6_s5_cyc_o_reg/NET0131 ,
		\rf_conf5_reg[12]/NET0131 ,
		\rf_conf5_reg[13]/NET0131 ,
		\s5_msel_arb1_state_reg[0]/NET0131 ,
		_w5699_
	);
	LUT2 #(
		.INIT('h8)
	) name3799 (
		\s5_msel_arb1_state_reg[1]/NET0131 ,
		\s5_msel_arb1_state_reg[2]/NET0131 ,
		_w5700_
	);
	LUT2 #(
		.INIT('h4)
	) name3800 (
		_w5699_,
		_w5700_,
		_w5701_
	);
	LUT3 #(
		.INIT('hb0)
	) name3801 (
		_w5697_,
		_w5698_,
		_w5701_,
		_w5702_
	);
	LUT3 #(
		.INIT('hfd)
	) name3802 (
		_w5689_,
		_w5695_,
		_w5702_,
		_w5703_
	);
	LUT2 #(
		.INIT('h4)
	) name3803 (
		\s5_msel_arb2_state_reg[1]/NET0131 ,
		\s5_msel_arb2_state_reg[2]/NET0131 ,
		_w5704_
	);
	LUT3 #(
		.INIT('h20)
	) name3804 (
		_w3385_,
		_w3386_,
		_w5704_,
		_w5705_
	);
	LUT2 #(
		.INIT('h4)
	) name3805 (
		_w3388_,
		_w3400_,
		_w5706_
	);
	LUT2 #(
		.INIT('h2)
	) name3806 (
		_w3391_,
		_w3393_,
		_w5707_
	);
	LUT4 #(
		.INIT('h0051)
	) name3807 (
		_w3388_,
		_w3391_,
		_w3393_,
		_w3396_,
		_w5708_
	);
	LUT3 #(
		.INIT('h10)
	) name3808 (
		_w3386_,
		_w3387_,
		_w5704_,
		_w5709_
	);
	LUT4 #(
		.INIT('h5455)
	) name3809 (
		_w5705_,
		_w5706_,
		_w5708_,
		_w5709_,
		_w5710_
	);
	LUT2 #(
		.INIT('h1)
	) name3810 (
		\s5_msel_arb2_state_reg[0]/NET0131 ,
		_w5710_,
		_w5711_
	);
	LUT2 #(
		.INIT('h1)
	) name3811 (
		_w3386_,
		_w3393_,
		_w5712_
	);
	LUT3 #(
		.INIT('hf2)
	) name3812 (
		_w3386_,
		_w3391_,
		_w3393_,
		_w5713_
	);
	LUT3 #(
		.INIT('h45)
	) name3813 (
		_w3385_,
		_w3387_,
		_w3388_,
		_w5714_
	);
	LUT3 #(
		.INIT('h04)
	) name3814 (
		_w3387_,
		_w3396_,
		_w3400_,
		_w5715_
	);
	LUT3 #(
		.INIT('h02)
	) name3815 (
		\s5_msel_arb2_state_reg[0]/NET0131 ,
		_w3387_,
		_w3400_,
		_w5716_
	);
	LUT4 #(
		.INIT('h0004)
	) name3816 (
		_w5707_,
		_w5714_,
		_w5715_,
		_w5716_,
		_w5717_
	);
	LUT3 #(
		.INIT('h04)
	) name3817 (
		\s5_msel_arb2_state_reg[0]/NET0131 ,
		\s5_msel_arb2_state_reg[1]/NET0131 ,
		\s5_msel_arb2_state_reg[2]/NET0131 ,
		_w5718_
	);
	LUT3 #(
		.INIT('h10)
	) name3818 (
		_w5713_,
		_w5717_,
		_w5718_,
		_w5719_
	);
	LUT2 #(
		.INIT('h1)
	) name3819 (
		_w5711_,
		_w5719_,
		_w5720_
	);
	LUT4 #(
		.INIT('hdf00)
	) name3820 (
		\m6_s5_cyc_o_reg/NET0131 ,
		\rf_conf5_reg[12]/NET0131 ,
		\rf_conf5_reg[13]/NET0131 ,
		\s5_msel_arb2_state_reg[0]/NET0131 ,
		_w5721_
	);
	LUT2 #(
		.INIT('h1)
	) name3821 (
		_w3385_,
		_w5721_,
		_w5722_
	);
	LUT3 #(
		.INIT('h01)
	) name3822 (
		_w3386_,
		_w3393_,
		_w3400_,
		_w5723_
	);
	LUT4 #(
		.INIT('he0ee)
	) name3823 (
		_w5706_,
		_w5708_,
		_w5722_,
		_w5723_,
		_w5724_
	);
	LUT4 #(
		.INIT('h0020)
	) name3824 (
		\m6_s5_cyc_o_reg/NET0131 ,
		\rf_conf5_reg[12]/NET0131 ,
		\rf_conf5_reg[13]/NET0131 ,
		\s5_msel_arb2_state_reg[0]/NET0131 ,
		_w5725_
	);
	LUT2 #(
		.INIT('h8)
	) name3825 (
		\s5_msel_arb2_state_reg[1]/NET0131 ,
		\s5_msel_arb2_state_reg[2]/NET0131 ,
		_w5726_
	);
	LUT2 #(
		.INIT('h4)
	) name3826 (
		_w5725_,
		_w5726_,
		_w5727_
	);
	LUT2 #(
		.INIT('h4)
	) name3827 (
		_w5724_,
		_w5727_,
		_w5728_
	);
	LUT3 #(
		.INIT('h51)
	) name3828 (
		_w3386_,
		_w5714_,
		_w5715_,
		_w5729_
	);
	LUT2 #(
		.INIT('h8)
	) name3829 (
		_w5712_,
		_w5716_,
		_w5730_
	);
	LUT3 #(
		.INIT('h15)
	) name3830 (
		_w3391_,
		_w5712_,
		_w5716_,
		_w5731_
	);
	LUT3 #(
		.INIT('h08)
	) name3831 (
		\s5_msel_arb2_state_reg[0]/NET0131 ,
		\s5_msel_arb2_state_reg[1]/NET0131 ,
		\s5_msel_arb2_state_reg[2]/NET0131 ,
		_w5732_
	);
	LUT3 #(
		.INIT('hb0)
	) name3832 (
		_w5729_,
		_w5731_,
		_w5732_,
		_w5733_
	);
	LUT2 #(
		.INIT('h2)
	) name3833 (
		\s5_msel_arb2_state_reg[0]/NET0131 ,
		\s5_msel_arb2_state_reg[1]/NET0131 ,
		_w5734_
	);
	LUT3 #(
		.INIT('h20)
	) name3834 (
		\s5_msel_arb2_state_reg[0]/NET0131 ,
		\s5_msel_arb2_state_reg[1]/NET0131 ,
		\s5_msel_arb2_state_reg[2]/NET0131 ,
		_w5735_
	);
	LUT3 #(
		.INIT('h01)
	) name3835 (
		_w3387_,
		_w5706_,
		_w5708_,
		_w5736_
	);
	LUT3 #(
		.INIT('h15)
	) name3836 (
		_w3385_,
		_w5712_,
		_w5716_,
		_w5737_
	);
	LUT3 #(
		.INIT('h8a)
	) name3837 (
		_w5735_,
		_w5736_,
		_w5737_,
		_w5738_
	);
	LUT4 #(
		.INIT('h0020)
	) name3838 (
		\m0_s5_cyc_o_reg/NET0131 ,
		\rf_conf5_reg[0]/NET0131 ,
		\rf_conf5_reg[1]/NET0131 ,
		\s5_msel_arb2_state_reg[0]/NET0131 ,
		_w5739_
	);
	LUT4 #(
		.INIT('h00f2)
	) name3839 (
		_w3391_,
		_w3393_,
		_w3396_,
		_w5739_,
		_w5740_
	);
	LUT3 #(
		.INIT('h01)
	) name3840 (
		_w3386_,
		_w3393_,
		_w5739_,
		_w5741_
	);
	LUT3 #(
		.INIT('h23)
	) name3841 (
		_w5714_,
		_w5740_,
		_w5741_,
		_w5742_
	);
	LUT2 #(
		.INIT('h1)
	) name3842 (
		\s5_msel_arb2_state_reg[1]/NET0131 ,
		\s5_msel_arb2_state_reg[2]/NET0131 ,
		_w5743_
	);
	LUT3 #(
		.INIT('hb0)
	) name3843 (
		_w5730_,
		_w5742_,
		_w5743_,
		_w5744_
	);
	LUT4 #(
		.INIT('h0001)
	) name3844 (
		_w5728_,
		_w5733_,
		_w5738_,
		_w5744_,
		_w5745_
	);
	LUT2 #(
		.INIT('h7)
	) name3845 (
		_w5720_,
		_w5745_,
		_w5746_
	);
	LUT2 #(
		.INIT('h2)
	) name3846 (
		\s5_msel_arb3_state_reg[1]/NET0131 ,
		\s5_msel_arb3_state_reg[2]/NET0131 ,
		_w5747_
	);
	LUT2 #(
		.INIT('h4)
	) name3847 (
		_w3425_,
		_w5747_,
		_w5748_
	);
	LUT2 #(
		.INIT('h1)
	) name3848 (
		_w3407_,
		_w3414_,
		_w5749_
	);
	LUT3 #(
		.INIT('hae)
	) name3849 (
		_w3407_,
		_w3414_,
		_w3415_,
		_w5750_
	);
	LUT2 #(
		.INIT('h1)
	) name3850 (
		_w3419_,
		_w3430_,
		_w5751_
	);
	LUT2 #(
		.INIT('h1)
	) name3851 (
		_w3415_,
		_w3420_,
		_w5752_
	);
	LUT4 #(
		.INIT('h7577)
	) name3852 (
		_w5748_,
		_w5750_,
		_w5751_,
		_w5752_,
		_w5753_
	);
	LUT3 #(
		.INIT('h0d)
	) name3853 (
		_w3417_,
		_w3418_,
		_w3419_,
		_w5754_
	);
	LUT4 #(
		.INIT('h00f2)
	) name3854 (
		_w3417_,
		_w3418_,
		_w3419_,
		_w3420_,
		_w5755_
	);
	LUT3 #(
		.INIT('h10)
	) name3855 (
		\s5_msel_arb3_state_reg[0]/NET0131 ,
		\s5_msel_arb3_state_reg[1]/NET0131 ,
		\s5_msel_arb3_state_reg[2]/NET0131 ,
		_w5756_
	);
	LUT4 #(
		.INIT('h2300)
	) name3856 (
		_w3407_,
		_w3408_,
		_w3415_,
		_w5756_,
		_w5757_
	);
	LUT3 #(
		.INIT('hd0)
	) name3857 (
		_w5749_,
		_w5755_,
		_w5757_,
		_w5758_
	);
	LUT3 #(
		.INIT('h0e)
	) name3858 (
		_w3408_,
		_w5753_,
		_w5758_,
		_w5759_
	);
	LUT2 #(
		.INIT('h1)
	) name3859 (
		\s5_msel_arb3_state_reg[1]/NET0131 ,
		\s5_msel_arb3_state_reg[2]/NET0131 ,
		_w5760_
	);
	LUT4 #(
		.INIT('h0080)
	) name3860 (
		\m0_s5_cyc_o_reg/NET0131 ,
		\rf_conf5_reg[0]/NET0131 ,
		\rf_conf5_reg[1]/NET0131 ,
		\s5_msel_arb3_state_reg[0]/NET0131 ,
		_w5761_
	);
	LUT2 #(
		.INIT('h2)
	) name3861 (
		_w5760_,
		_w5761_,
		_w5762_
	);
	LUT2 #(
		.INIT('h1)
	) name3862 (
		_w3408_,
		_w3418_,
		_w5763_
	);
	LUT4 #(
		.INIT('h4fcf)
	) name3863 (
		_w5750_,
		_w5754_,
		_w5762_,
		_w5763_,
		_w5764_
	);
	LUT3 #(
		.INIT('h20)
	) name3864 (
		_w3417_,
		_w3425_,
		_w5747_,
		_w5765_
	);
	LUT3 #(
		.INIT('h20)
	) name3865 (
		\s5_msel_arb3_state_reg[0]/NET0131 ,
		\s5_msel_arb3_state_reg[1]/NET0131 ,
		\s5_msel_arb3_state_reg[2]/NET0131 ,
		_w5766_
	);
	LUT2 #(
		.INIT('h8)
	) name3866 (
		_w3407_,
		_w5766_,
		_w5767_
	);
	LUT2 #(
		.INIT('h1)
	) name3867 (
		_w5765_,
		_w5767_,
		_w5768_
	);
	LUT2 #(
		.INIT('h8)
	) name3868 (
		_w5764_,
		_w5768_,
		_w5769_
	);
	LUT3 #(
		.INIT('h02)
	) name3869 (
		\s5_msel_arb3_state_reg[0]/NET0131 ,
		\s5_msel_arb3_state_reg[1]/NET0131 ,
		\s5_msel_arb3_state_reg[2]/NET0131 ,
		_w5770_
	);
	LUT4 #(
		.INIT('h0100)
	) name3870 (
		_w3408_,
		_w3418_,
		_w3420_,
		_w5770_,
		_w5771_
	);
	LUT2 #(
		.INIT('h4)
	) name3871 (
		_w3407_,
		_w5766_,
		_w5772_
	);
	LUT2 #(
		.INIT('h1)
	) name3872 (
		_w5771_,
		_w5772_,
		_w5773_
	);
	LUT2 #(
		.INIT('h4)
	) name3873 (
		_w3414_,
		_w3420_,
		_w5774_
	);
	LUT4 #(
		.INIT('h0051)
	) name3874 (
		_w3414_,
		_w3417_,
		_w3418_,
		_w3419_,
		_w5775_
	);
	LUT4 #(
		.INIT('h7f00)
	) name3875 (
		\m0_s5_cyc_o_reg/NET0131 ,
		\rf_conf5_reg[0]/NET0131 ,
		\rf_conf5_reg[1]/NET0131 ,
		\s5_msel_arb3_state_reg[0]/NET0131 ,
		_w5776_
	);
	LUT3 #(
		.INIT('h10)
	) name3876 (
		_w3408_,
		_w3418_,
		_w5776_,
		_w5777_
	);
	LUT4 #(
		.INIT('h0054)
	) name3877 (
		_w5771_,
		_w5774_,
		_w5775_,
		_w5777_,
		_w5778_
	);
	LUT3 #(
		.INIT('h01)
	) name3878 (
		_w3415_,
		_w5773_,
		_w5778_,
		_w5779_
	);
	LUT4 #(
		.INIT('h007f)
	) name3879 (
		\m5_s5_cyc_o_reg/NET0131 ,
		\rf_conf5_reg[10]/NET0131 ,
		\rf_conf5_reg[11]/NET0131 ,
		\s5_msel_arb3_state_reg[0]/NET0131 ,
		_w5780_
	);
	LUT4 #(
		.INIT('h0001)
	) name3880 (
		_w3408_,
		_w3418_,
		_w3420_,
		_w5780_,
		_w5781_
	);
	LUT3 #(
		.INIT('h0e)
	) name3881 (
		_w5774_,
		_w5775_,
		_w5781_,
		_w5782_
	);
	LUT4 #(
		.INIT('h0080)
	) name3882 (
		\m6_s5_cyc_o_reg/NET0131 ,
		\rf_conf5_reg[12]/NET0131 ,
		\rf_conf5_reg[13]/NET0131 ,
		\s5_msel_arb3_state_reg[0]/NET0131 ,
		_w5783_
	);
	LUT3 #(
		.INIT('h10)
	) name3883 (
		_w3407_,
		_w3414_,
		_w3415_,
		_w5784_
	);
	LUT4 #(
		.INIT('h020a)
	) name3884 (
		_w3433_,
		_w5754_,
		_w5783_,
		_w5784_,
		_w5785_
	);
	LUT2 #(
		.INIT('h4)
	) name3885 (
		_w5782_,
		_w5785_,
		_w5786_
	);
	LUT4 #(
		.INIT('hfff7)
	) name3886 (
		_w5759_,
		_w5769_,
		_w5779_,
		_w5786_,
		_w5787_
	);
	LUT2 #(
		.INIT('h4)
	) name3887 (
		_w2575_,
		_w2583_,
		_w5788_
	);
	LUT3 #(
		.INIT('h04)
	) name3888 (
		_w2571_,
		_w2573_,
		_w2574_,
		_w5789_
	);
	LUT4 #(
		.INIT('hfd00)
	) name3889 (
		\m4_s6_cyc_o_reg/NET0131 ,
		\rf_conf6_reg[8]/NET0131 ,
		\rf_conf6_reg[9]/NET0131 ,
		\s6_msel_arb0_state_reg[0]/NET0131 ,
		_w5790_
	);
	LUT3 #(
		.INIT('h10)
	) name3890 (
		_w2574_,
		_w2576_,
		_w5790_,
		_w5791_
	);
	LUT3 #(
		.INIT('hf2)
	) name3891 (
		_w2570_,
		_w2571_,
		_w2578_,
		_w5792_
	);
	LUT4 #(
		.INIT('h000d)
	) name3892 (
		_w2570_,
		_w2571_,
		_w2575_,
		_w2578_,
		_w5793_
	);
	LUT4 #(
		.INIT('h5455)
	) name3893 (
		_w5788_,
		_w5789_,
		_w5791_,
		_w5793_,
		_w5794_
	);
	LUT2 #(
		.INIT('h8)
	) name3894 (
		_w2597_,
		_w5794_,
		_w5795_
	);
	LUT2 #(
		.INIT('h8)
	) name3895 (
		\s6_msel_arb0_state_reg[1]/NET0131 ,
		\s6_msel_arb0_state_reg[2]/NET0131 ,
		_w5796_
	);
	LUT2 #(
		.INIT('h2)
	) name3896 (
		_w2578_,
		_w2583_,
		_w5797_
	);
	LUT3 #(
		.INIT('h51)
	) name3897 (
		_w2575_,
		_w2578_,
		_w2583_,
		_w5798_
	);
	LUT4 #(
		.INIT('h2232)
	) name3898 (
		_w2575_,
		_w2576_,
		_w2578_,
		_w2583_,
		_w5799_
	);
	LUT2 #(
		.INIT('h1)
	) name3899 (
		_w2571_,
		_w2583_,
		_w5800_
	);
	LUT4 #(
		.INIT('h00fd)
	) name3900 (
		\m5_s6_cyc_o_reg/NET0131 ,
		\rf_conf6_reg[10]/NET0131 ,
		\rf_conf6_reg[11]/NET0131 ,
		\s6_msel_arb0_state_reg[0]/NET0131 ,
		_w5801_
	);
	LUT3 #(
		.INIT('h01)
	) name3901 (
		_w2571_,
		_w2583_,
		_w5801_,
		_w5802_
	);
	LUT2 #(
		.INIT('h4)
	) name3902 (
		_w2570_,
		_w2574_,
		_w5803_
	);
	LUT3 #(
		.INIT('h0b)
	) name3903 (
		_w2570_,
		_w2574_,
		_w2576_,
		_w5804_
	);
	LUT4 #(
		.INIT('h0111)
	) name3904 (
		_w2573_,
		_w5799_,
		_w5802_,
		_w5804_,
		_w5805_
	);
	LUT4 #(
		.INIT('h1101)
	) name3905 (
		_w2570_,
		_w2573_,
		_w2575_,
		_w2576_,
		_w5806_
	);
	LUT4 #(
		.INIT('hfd00)
	) name3906 (
		\m2_s6_cyc_o_reg/NET0131 ,
		\rf_conf6_reg[4]/NET0131 ,
		\rf_conf6_reg[5]/NET0131 ,
		\s6_msel_arb0_state_reg[0]/NET0131 ,
		_w5807_
	);
	LUT4 #(
		.INIT('h0e0f)
	) name3907 (
		_w2574_,
		_w2576_,
		_w2578_,
		_w5807_,
		_w5808_
	);
	LUT2 #(
		.INIT('h2)
	) name3908 (
		\s6_msel_arb0_state_reg[1]/NET0131 ,
		\s6_msel_arb0_state_reg[2]/NET0131 ,
		_w5809_
	);
	LUT3 #(
		.INIT('hd0)
	) name3909 (
		_w2571_,
		_w2578_,
		_w5809_,
		_w5810_
	);
	LUT4 #(
		.INIT('h1f00)
	) name3910 (
		_w5803_,
		_w5806_,
		_w5808_,
		_w5810_,
		_w5811_
	);
	LUT3 #(
		.INIT('h0d)
	) name3911 (
		_w5796_,
		_w5805_,
		_w5811_,
		_w5812_
	);
	LUT3 #(
		.INIT('h8a)
	) name3912 (
		\s6_msel_arb0_state_reg[0]/NET0131 ,
		_w5795_,
		_w5812_,
		_w5813_
	);
	LUT3 #(
		.INIT('h02)
	) name3913 (
		\s6_msel_arb0_state_reg[0]/NET0131 ,
		_w2574_,
		_w2576_,
		_w5814_
	);
	LUT4 #(
		.INIT('h55fd)
	) name3914 (
		_w5800_,
		_w5803_,
		_w5806_,
		_w5814_,
		_w5815_
	);
	LUT3 #(
		.INIT('h8c)
	) name3915 (
		_w5797_,
		_w5809_,
		_w5815_,
		_w5816_
	);
	LUT3 #(
		.INIT('h20)
	) name3916 (
		_w2573_,
		_w2574_,
		_w5796_,
		_w5817_
	);
	LUT3 #(
		.INIT('h10)
	) name3917 (
		_w2574_,
		_w2576_,
		_w5796_,
		_w5818_
	);
	LUT4 #(
		.INIT('h020f)
	) name3918 (
		_w5798_,
		_w5802_,
		_w5817_,
		_w5818_,
		_w5819_
	);
	LUT3 #(
		.INIT('h20)
	) name3919 (
		_w2575_,
		_w2576_,
		_w2597_,
		_w5820_
	);
	LUT2 #(
		.INIT('h1)
	) name3920 (
		_w2571_,
		_w2574_,
		_w5821_
	);
	LUT4 #(
		.INIT('h00fd)
	) name3921 (
		\m7_s6_cyc_o_reg/NET0131 ,
		\rf_conf6_reg[14]/NET0131 ,
		\rf_conf6_reg[15]/NET0131 ,
		\s6_msel_arb0_state_reg[0]/NET0131 ,
		_w5822_
	);
	LUT3 #(
		.INIT('h01)
	) name3922 (
		_w2571_,
		_w2574_,
		_w5822_,
		_w5823_
	);
	LUT3 #(
		.INIT('h10)
	) name3923 (
		_w2576_,
		_w2583_,
		_w2597_,
		_w5824_
	);
	LUT4 #(
		.INIT('h0133)
	) name3924 (
		_w5792_,
		_w5820_,
		_w5823_,
		_w5824_,
		_w5825_
	);
	LUT2 #(
		.INIT('h8)
	) name3925 (
		_w5819_,
		_w5825_,
		_w5826_
	);
	LUT3 #(
		.INIT('h02)
	) name3926 (
		\s6_msel_arb0_state_reg[0]/NET0131 ,
		_w2576_,
		_w2583_,
		_w5827_
	);
	LUT3 #(
		.INIT('h80)
	) name3927 (
		_w2600_,
		_w5821_,
		_w5827_,
		_w5828_
	);
	LUT3 #(
		.INIT('h04)
	) name3928 (
		_w2576_,
		_w2578_,
		_w2583_,
		_w5829_
	);
	LUT4 #(
		.INIT('h0002)
	) name3929 (
		\m4_s6_cyc_o_reg/NET0131 ,
		\rf_conf6_reg[8]/NET0131 ,
		\rf_conf6_reg[9]/NET0131 ,
		\s6_msel_arb0_state_reg[0]/NET0131 ,
		_w5830_
	);
	LUT4 #(
		.INIT('h00b0)
	) name3930 (
		_w2570_,
		_w2574_,
		_w2600_,
		_w5830_,
		_w5831_
	);
	LUT3 #(
		.INIT('hd0)
	) name3931 (
		_w5806_,
		_w5829_,
		_w5831_,
		_w5832_
	);
	LUT2 #(
		.INIT('h1)
	) name3932 (
		_w5828_,
		_w5832_,
		_w5833_
	);
	LUT4 #(
		.INIT('hba00)
	) name3933 (
		\s6_msel_arb0_state_reg[0]/NET0131 ,
		_w5816_,
		_w5826_,
		_w5833_,
		_w5834_
	);
	LUT2 #(
		.INIT('hb)
	) name3934 (
		_w5813_,
		_w5834_,
		_w5835_
	);
	LUT3 #(
		.INIT('hf2)
	) name3935 (
		_w3839_,
		_w3840_,
		_w3843_,
		_w5836_
	);
	LUT4 #(
		.INIT('h0008)
	) name3936 (
		\m4_s6_cyc_o_reg/NET0131 ,
		\rf_conf6_reg[8]/NET0131 ,
		\rf_conf6_reg[9]/NET0131 ,
		\s6_msel_arb1_state_reg[0]/NET0131 ,
		_w5837_
	);
	LUT2 #(
		.INIT('h2)
	) name3937 (
		_w3849_,
		_w5837_,
		_w5838_
	);
	LUT2 #(
		.INIT('h8)
	) name3938 (
		_w5836_,
		_w5838_,
		_w5839_
	);
	LUT3 #(
		.INIT('hf2)
	) name3939 (
		_w3833_,
		_w3834_,
		_w3837_,
		_w5840_
	);
	LUT3 #(
		.INIT('h02)
	) name3940 (
		\s6_msel_arb1_state_reg[0]/NET0131 ,
		_w3834_,
		_w3842_,
		_w5841_
	);
	LUT2 #(
		.INIT('h1)
	) name3941 (
		_w3836_,
		_w3840_,
		_w5842_
	);
	LUT4 #(
		.INIT('h0010)
	) name3942 (
		_w3836_,
		_w3840_,
		_w3849_,
		_w5837_,
		_w5843_
	);
	LUT3 #(
		.INIT('he0)
	) name3943 (
		_w5840_,
		_w5841_,
		_w5843_,
		_w5844_
	);
	LUT4 #(
		.INIT('h0031)
	) name3944 (
		_w3834_,
		_w3836_,
		_w3837_,
		_w3840_,
		_w5845_
	);
	LUT4 #(
		.INIT('h4445)
	) name3945 (
		_w3833_,
		_w3842_,
		_w5836_,
		_w5845_,
		_w5846_
	);
	LUT3 #(
		.INIT('h08)
	) name3946 (
		\s6_msel_arb1_state_reg[0]/NET0131 ,
		\s6_msel_arb1_state_reg[1]/NET0131 ,
		\s6_msel_arb1_state_reg[2]/NET0131 ,
		_w5847_
	);
	LUT4 #(
		.INIT('h0001)
	) name3947 (
		_w3833_,
		_w3837_,
		_w3839_,
		_w3843_,
		_w5848_
	);
	LUT2 #(
		.INIT('h4)
	) name3948 (
		_w3834_,
		_w3852_,
		_w5849_
	);
	LUT3 #(
		.INIT('h45)
	) name3949 (
		_w5847_,
		_w5848_,
		_w5849_,
		_w5850_
	);
	LUT4 #(
		.INIT('h1110)
	) name3950 (
		_w5839_,
		_w5844_,
		_w5846_,
		_w5850_,
		_w5851_
	);
	LUT4 #(
		.INIT('h0008)
	) name3951 (
		\m0_s6_cyc_o_reg/NET0131 ,
		\rf_conf6_reg[0]/NET0131 ,
		\rf_conf6_reg[1]/NET0131 ,
		\s6_msel_arb1_state_reg[0]/NET0131 ,
		_w5852_
	);
	LUT4 #(
		.INIT('h00f2)
	) name3952 (
		_w3833_,
		_w3834_,
		_w3837_,
		_w5852_,
		_w5853_
	);
	LUT3 #(
		.INIT('h01)
	) name3953 (
		_w3834_,
		_w3842_,
		_w5852_,
		_w5854_
	);
	LUT3 #(
		.INIT('h13)
	) name3954 (
		_w5836_,
		_w5853_,
		_w5854_,
		_w5855_
	);
	LUT2 #(
		.INIT('h8)
	) name3955 (
		_w5841_,
		_w5842_,
		_w5856_
	);
	LUT3 #(
		.INIT('ha2)
	) name3956 (
		_w3845_,
		_w5855_,
		_w5856_,
		_w5857_
	);
	LUT3 #(
		.INIT('h10)
	) name3957 (
		_w3834_,
		_w3842_,
		_w3843_,
		_w5858_
	);
	LUT3 #(
		.INIT('h54)
	) name3958 (
		_w3836_,
		_w5840_,
		_w5858_,
		_w5859_
	);
	LUT3 #(
		.INIT('h15)
	) name3959 (
		_w3839_,
		_w5841_,
		_w5842_,
		_w5860_
	);
	LUT4 #(
		.INIT('h0008)
	) name3960 (
		\m6_s6_cyc_o_reg/NET0131 ,
		\rf_conf6_reg[12]/NET0131 ,
		\rf_conf6_reg[13]/NET0131 ,
		\s6_msel_arb1_state_reg[0]/NET0131 ,
		_w5861_
	);
	LUT2 #(
		.INIT('h8)
	) name3961 (
		\s6_msel_arb1_state_reg[1]/NET0131 ,
		\s6_msel_arb1_state_reg[2]/NET0131 ,
		_w5862_
	);
	LUT2 #(
		.INIT('h4)
	) name3962 (
		_w5861_,
		_w5862_,
		_w5863_
	);
	LUT3 #(
		.INIT('hb0)
	) name3963 (
		_w5859_,
		_w5860_,
		_w5863_,
		_w5864_
	);
	LUT3 #(
		.INIT('hfd)
	) name3964 (
		_w5851_,
		_w5857_,
		_w5864_,
		_w5865_
	);
	LUT2 #(
		.INIT('h4)
	) name3965 (
		\s6_msel_arb2_state_reg[1]/NET0131 ,
		\s6_msel_arb2_state_reg[2]/NET0131 ,
		_w5866_
	);
	LUT3 #(
		.INIT('h20)
	) name3966 (
		_w3087_,
		_w3088_,
		_w5866_,
		_w5867_
	);
	LUT2 #(
		.INIT('h4)
	) name3967 (
		_w3090_,
		_w3102_,
		_w5868_
	);
	LUT2 #(
		.INIT('h2)
	) name3968 (
		_w3093_,
		_w3095_,
		_w5869_
	);
	LUT4 #(
		.INIT('h0051)
	) name3969 (
		_w3090_,
		_w3093_,
		_w3095_,
		_w3098_,
		_w5870_
	);
	LUT3 #(
		.INIT('h10)
	) name3970 (
		_w3088_,
		_w3089_,
		_w5866_,
		_w5871_
	);
	LUT4 #(
		.INIT('h5455)
	) name3971 (
		_w5867_,
		_w5868_,
		_w5870_,
		_w5871_,
		_w5872_
	);
	LUT2 #(
		.INIT('h1)
	) name3972 (
		\s6_msel_arb2_state_reg[0]/NET0131 ,
		_w5872_,
		_w5873_
	);
	LUT2 #(
		.INIT('h1)
	) name3973 (
		_w3088_,
		_w3095_,
		_w5874_
	);
	LUT3 #(
		.INIT('hf2)
	) name3974 (
		_w3088_,
		_w3093_,
		_w3095_,
		_w5875_
	);
	LUT3 #(
		.INIT('h45)
	) name3975 (
		_w3087_,
		_w3089_,
		_w3090_,
		_w5876_
	);
	LUT3 #(
		.INIT('h04)
	) name3976 (
		_w3089_,
		_w3098_,
		_w3102_,
		_w5877_
	);
	LUT3 #(
		.INIT('h02)
	) name3977 (
		\s6_msel_arb2_state_reg[0]/NET0131 ,
		_w3089_,
		_w3102_,
		_w5878_
	);
	LUT4 #(
		.INIT('h0004)
	) name3978 (
		_w5869_,
		_w5876_,
		_w5877_,
		_w5878_,
		_w5879_
	);
	LUT3 #(
		.INIT('h04)
	) name3979 (
		\s6_msel_arb2_state_reg[0]/NET0131 ,
		\s6_msel_arb2_state_reg[1]/NET0131 ,
		\s6_msel_arb2_state_reg[2]/NET0131 ,
		_w5880_
	);
	LUT3 #(
		.INIT('h10)
	) name3980 (
		_w5875_,
		_w5879_,
		_w5880_,
		_w5881_
	);
	LUT2 #(
		.INIT('h1)
	) name3981 (
		_w5873_,
		_w5881_,
		_w5882_
	);
	LUT4 #(
		.INIT('hdf00)
	) name3982 (
		\m6_s6_cyc_o_reg/NET0131 ,
		\rf_conf6_reg[12]/NET0131 ,
		\rf_conf6_reg[13]/NET0131 ,
		\s6_msel_arb2_state_reg[0]/NET0131 ,
		_w5883_
	);
	LUT2 #(
		.INIT('h1)
	) name3983 (
		_w3087_,
		_w5883_,
		_w5884_
	);
	LUT3 #(
		.INIT('h01)
	) name3984 (
		_w3088_,
		_w3095_,
		_w3102_,
		_w5885_
	);
	LUT4 #(
		.INIT('he0ee)
	) name3985 (
		_w5868_,
		_w5870_,
		_w5884_,
		_w5885_,
		_w5886_
	);
	LUT4 #(
		.INIT('h0020)
	) name3986 (
		\m6_s6_cyc_o_reg/NET0131 ,
		\rf_conf6_reg[12]/NET0131 ,
		\rf_conf6_reg[13]/NET0131 ,
		\s6_msel_arb2_state_reg[0]/NET0131 ,
		_w5887_
	);
	LUT2 #(
		.INIT('h8)
	) name3987 (
		\s6_msel_arb2_state_reg[1]/NET0131 ,
		\s6_msel_arb2_state_reg[2]/NET0131 ,
		_w5888_
	);
	LUT2 #(
		.INIT('h4)
	) name3988 (
		_w5887_,
		_w5888_,
		_w5889_
	);
	LUT2 #(
		.INIT('h4)
	) name3989 (
		_w5886_,
		_w5889_,
		_w5890_
	);
	LUT3 #(
		.INIT('h51)
	) name3990 (
		_w3088_,
		_w5876_,
		_w5877_,
		_w5891_
	);
	LUT2 #(
		.INIT('h8)
	) name3991 (
		_w5874_,
		_w5878_,
		_w5892_
	);
	LUT3 #(
		.INIT('h15)
	) name3992 (
		_w3093_,
		_w5874_,
		_w5878_,
		_w5893_
	);
	LUT3 #(
		.INIT('h08)
	) name3993 (
		\s6_msel_arb2_state_reg[0]/NET0131 ,
		\s6_msel_arb2_state_reg[1]/NET0131 ,
		\s6_msel_arb2_state_reg[2]/NET0131 ,
		_w5894_
	);
	LUT3 #(
		.INIT('hb0)
	) name3994 (
		_w5891_,
		_w5893_,
		_w5894_,
		_w5895_
	);
	LUT2 #(
		.INIT('h2)
	) name3995 (
		\s6_msel_arb2_state_reg[0]/NET0131 ,
		\s6_msel_arb2_state_reg[1]/NET0131 ,
		_w5896_
	);
	LUT3 #(
		.INIT('h20)
	) name3996 (
		\s6_msel_arb2_state_reg[0]/NET0131 ,
		\s6_msel_arb2_state_reg[1]/NET0131 ,
		\s6_msel_arb2_state_reg[2]/NET0131 ,
		_w5897_
	);
	LUT3 #(
		.INIT('h01)
	) name3997 (
		_w3089_,
		_w5868_,
		_w5870_,
		_w5898_
	);
	LUT3 #(
		.INIT('h15)
	) name3998 (
		_w3087_,
		_w5874_,
		_w5878_,
		_w5899_
	);
	LUT3 #(
		.INIT('h8a)
	) name3999 (
		_w5897_,
		_w5898_,
		_w5899_,
		_w5900_
	);
	LUT4 #(
		.INIT('h0020)
	) name4000 (
		\m0_s6_cyc_o_reg/NET0131 ,
		\rf_conf6_reg[0]/NET0131 ,
		\rf_conf6_reg[1]/NET0131 ,
		\s6_msel_arb2_state_reg[0]/NET0131 ,
		_w5901_
	);
	LUT4 #(
		.INIT('h00f2)
	) name4001 (
		_w3093_,
		_w3095_,
		_w3098_,
		_w5901_,
		_w5902_
	);
	LUT3 #(
		.INIT('h01)
	) name4002 (
		_w3088_,
		_w3095_,
		_w5901_,
		_w5903_
	);
	LUT3 #(
		.INIT('h23)
	) name4003 (
		_w5876_,
		_w5902_,
		_w5903_,
		_w5904_
	);
	LUT2 #(
		.INIT('h1)
	) name4004 (
		\s6_msel_arb2_state_reg[1]/NET0131 ,
		\s6_msel_arb2_state_reg[2]/NET0131 ,
		_w5905_
	);
	LUT3 #(
		.INIT('hb0)
	) name4005 (
		_w5892_,
		_w5904_,
		_w5905_,
		_w5906_
	);
	LUT4 #(
		.INIT('h0001)
	) name4006 (
		_w5890_,
		_w5895_,
		_w5900_,
		_w5906_,
		_w5907_
	);
	LUT2 #(
		.INIT('h7)
	) name4007 (
		_w5882_,
		_w5907_,
		_w5908_
	);
	LUT2 #(
		.INIT('h2)
	) name4008 (
		\s6_msel_arb3_state_reg[1]/NET0131 ,
		\s6_msel_arb3_state_reg[2]/NET0131 ,
		_w5909_
	);
	LUT2 #(
		.INIT('h4)
	) name4009 (
		_w3455_,
		_w5909_,
		_w5910_
	);
	LUT2 #(
		.INIT('h1)
	) name4010 (
		_w3437_,
		_w3444_,
		_w5911_
	);
	LUT3 #(
		.INIT('hae)
	) name4011 (
		_w3437_,
		_w3444_,
		_w3445_,
		_w5912_
	);
	LUT2 #(
		.INIT('h1)
	) name4012 (
		_w3449_,
		_w3460_,
		_w5913_
	);
	LUT2 #(
		.INIT('h1)
	) name4013 (
		_w3445_,
		_w3450_,
		_w5914_
	);
	LUT4 #(
		.INIT('h7577)
	) name4014 (
		_w5910_,
		_w5912_,
		_w5913_,
		_w5914_,
		_w5915_
	);
	LUT3 #(
		.INIT('h0d)
	) name4015 (
		_w3447_,
		_w3448_,
		_w3449_,
		_w5916_
	);
	LUT4 #(
		.INIT('h00f2)
	) name4016 (
		_w3447_,
		_w3448_,
		_w3449_,
		_w3450_,
		_w5917_
	);
	LUT3 #(
		.INIT('h10)
	) name4017 (
		\s6_msel_arb3_state_reg[0]/NET0131 ,
		\s6_msel_arb3_state_reg[1]/NET0131 ,
		\s6_msel_arb3_state_reg[2]/NET0131 ,
		_w5918_
	);
	LUT4 #(
		.INIT('h2300)
	) name4018 (
		_w3437_,
		_w3438_,
		_w3445_,
		_w5918_,
		_w5919_
	);
	LUT3 #(
		.INIT('hd0)
	) name4019 (
		_w5911_,
		_w5917_,
		_w5919_,
		_w5920_
	);
	LUT3 #(
		.INIT('h0e)
	) name4020 (
		_w3438_,
		_w5915_,
		_w5920_,
		_w5921_
	);
	LUT2 #(
		.INIT('h1)
	) name4021 (
		\s6_msel_arb3_state_reg[1]/NET0131 ,
		\s6_msel_arb3_state_reg[2]/NET0131 ,
		_w5922_
	);
	LUT4 #(
		.INIT('h0080)
	) name4022 (
		\m0_s6_cyc_o_reg/NET0131 ,
		\rf_conf6_reg[0]/NET0131 ,
		\rf_conf6_reg[1]/NET0131 ,
		\s6_msel_arb3_state_reg[0]/NET0131 ,
		_w5923_
	);
	LUT2 #(
		.INIT('h2)
	) name4023 (
		_w5922_,
		_w5923_,
		_w5924_
	);
	LUT2 #(
		.INIT('h1)
	) name4024 (
		_w3438_,
		_w3448_,
		_w5925_
	);
	LUT4 #(
		.INIT('h4fcf)
	) name4025 (
		_w5912_,
		_w5916_,
		_w5924_,
		_w5925_,
		_w5926_
	);
	LUT3 #(
		.INIT('h20)
	) name4026 (
		_w3447_,
		_w3455_,
		_w5909_,
		_w5927_
	);
	LUT3 #(
		.INIT('h20)
	) name4027 (
		\s6_msel_arb3_state_reg[0]/NET0131 ,
		\s6_msel_arb3_state_reg[1]/NET0131 ,
		\s6_msel_arb3_state_reg[2]/NET0131 ,
		_w5928_
	);
	LUT2 #(
		.INIT('h8)
	) name4028 (
		_w3437_,
		_w5928_,
		_w5929_
	);
	LUT2 #(
		.INIT('h1)
	) name4029 (
		_w5927_,
		_w5929_,
		_w5930_
	);
	LUT2 #(
		.INIT('h8)
	) name4030 (
		_w5926_,
		_w5930_,
		_w5931_
	);
	LUT3 #(
		.INIT('h02)
	) name4031 (
		\s6_msel_arb3_state_reg[0]/NET0131 ,
		\s6_msel_arb3_state_reg[1]/NET0131 ,
		\s6_msel_arb3_state_reg[2]/NET0131 ,
		_w5932_
	);
	LUT4 #(
		.INIT('h0100)
	) name4032 (
		_w3438_,
		_w3448_,
		_w3450_,
		_w5932_,
		_w5933_
	);
	LUT2 #(
		.INIT('h4)
	) name4033 (
		_w3437_,
		_w5928_,
		_w5934_
	);
	LUT2 #(
		.INIT('h1)
	) name4034 (
		_w5933_,
		_w5934_,
		_w5935_
	);
	LUT2 #(
		.INIT('h4)
	) name4035 (
		_w3444_,
		_w3450_,
		_w5936_
	);
	LUT4 #(
		.INIT('h0051)
	) name4036 (
		_w3444_,
		_w3447_,
		_w3448_,
		_w3449_,
		_w5937_
	);
	LUT4 #(
		.INIT('h7f00)
	) name4037 (
		\m0_s6_cyc_o_reg/NET0131 ,
		\rf_conf6_reg[0]/NET0131 ,
		\rf_conf6_reg[1]/NET0131 ,
		\s6_msel_arb3_state_reg[0]/NET0131 ,
		_w5938_
	);
	LUT3 #(
		.INIT('h10)
	) name4038 (
		_w3438_,
		_w3448_,
		_w5938_,
		_w5939_
	);
	LUT4 #(
		.INIT('h0054)
	) name4039 (
		_w5933_,
		_w5936_,
		_w5937_,
		_w5939_,
		_w5940_
	);
	LUT3 #(
		.INIT('h01)
	) name4040 (
		_w3445_,
		_w5935_,
		_w5940_,
		_w5941_
	);
	LUT4 #(
		.INIT('h007f)
	) name4041 (
		\m5_s6_cyc_o_reg/NET0131 ,
		\rf_conf6_reg[10]/NET0131 ,
		\rf_conf6_reg[11]/NET0131 ,
		\s6_msel_arb3_state_reg[0]/NET0131 ,
		_w5942_
	);
	LUT4 #(
		.INIT('h0001)
	) name4042 (
		_w3438_,
		_w3448_,
		_w3450_,
		_w5942_,
		_w5943_
	);
	LUT3 #(
		.INIT('h0e)
	) name4043 (
		_w5936_,
		_w5937_,
		_w5943_,
		_w5944_
	);
	LUT4 #(
		.INIT('h0080)
	) name4044 (
		\m6_s6_cyc_o_reg/NET0131 ,
		\rf_conf6_reg[12]/NET0131 ,
		\rf_conf6_reg[13]/NET0131 ,
		\s6_msel_arb3_state_reg[0]/NET0131 ,
		_w5945_
	);
	LUT3 #(
		.INIT('h10)
	) name4045 (
		_w3437_,
		_w3444_,
		_w3445_,
		_w5946_
	);
	LUT4 #(
		.INIT('h020a)
	) name4046 (
		_w3463_,
		_w5916_,
		_w5945_,
		_w5946_,
		_w5947_
	);
	LUT2 #(
		.INIT('h4)
	) name4047 (
		_w5944_,
		_w5947_,
		_w5948_
	);
	LUT4 #(
		.INIT('hfff7)
	) name4048 (
		_w5921_,
		_w5931_,
		_w5941_,
		_w5948_,
		_w5949_
	);
	LUT2 #(
		.INIT('h4)
	) name4049 (
		_w2727_,
		_w2732_,
		_w5950_
	);
	LUT4 #(
		.INIT('h000d)
	) name4050 (
		_w2722_,
		_w2723_,
		_w2727_,
		_w2731_,
		_w5951_
	);
	LUT3 #(
		.INIT('h01)
	) name4051 (
		_w2723_,
		_w2725_,
		_w2732_,
		_w5952_
	);
	LUT4 #(
		.INIT('h00fd)
	) name4052 (
		\m5_s7_cyc_o_reg/NET0131 ,
		\rf_conf7_reg[10]/NET0131 ,
		\rf_conf7_reg[11]/NET0131 ,
		\s7_msel_arb0_state_reg[0]/NET0131 ,
		_w5953_
	);
	LUT3 #(
		.INIT('hce)
	) name4053 (
		\s7_msel_arb0_state_reg[0]/NET0131 ,
		_w2726_,
		_w2728_,
		_w5954_
	);
	LUT4 #(
		.INIT('h0eee)
	) name4054 (
		_w5950_,
		_w5951_,
		_w5952_,
		_w5954_,
		_w5955_
	);
	LUT3 #(
		.INIT('hae)
	) name4055 (
		_w2726_,
		_w2727_,
		_w2728_,
		_w5956_
	);
	LUT2 #(
		.INIT('h4)
	) name4056 (
		\s7_msel_arb0_state_reg[1]/NET0131 ,
		\s7_msel_arb0_state_reg[2]/NET0131 ,
		_w5957_
	);
	LUT4 #(
		.INIT('h0002)
	) name4057 (
		\m1_s7_cyc_o_reg/NET0131 ,
		\rf_conf7_reg[2]/NET0131 ,
		\rf_conf7_reg[3]/NET0131 ,
		\s7_msel_arb0_state_reg[1]/NET0131 ,
		_w5958_
	);
	LUT2 #(
		.INIT('h1)
	) name4058 (
		_w5957_,
		_w5958_,
		_w5959_
	);
	LUT3 #(
		.INIT('h23)
	) name4059 (
		_w2722_,
		_w2723_,
		_w2725_,
		_w5960_
	);
	LUT4 #(
		.INIT('h00dc)
	) name4060 (
		_w2722_,
		_w2723_,
		_w2725_,
		_w2731_,
		_w5961_
	);
	LUT3 #(
		.INIT('ha8)
	) name4061 (
		\s7_msel_arb0_state_reg[2]/NET0131 ,
		_w2728_,
		_w2732_,
		_w5962_
	);
	LUT4 #(
		.INIT('hdddc)
	) name4062 (
		_w5956_,
		_w5959_,
		_w5961_,
		_w5962_,
		_w5963_
	);
	LUT4 #(
		.INIT('h08aa)
	) name4063 (
		\s7_msel_arb0_state_reg[0]/NET0131 ,
		_w2755_,
		_w5955_,
		_w5963_,
		_w5964_
	);
	LUT3 #(
		.INIT('h02)
	) name4064 (
		\s7_msel_arb0_state_reg[0]/NET0131 ,
		_w2728_,
		_w2732_,
		_w5965_
	);
	LUT2 #(
		.INIT('h1)
	) name4065 (
		_w2723_,
		_w2725_,
		_w5966_
	);
	LUT3 #(
		.INIT('h80)
	) name4066 (
		_w2750_,
		_w5965_,
		_w5966_,
		_w5967_
	);
	LUT3 #(
		.INIT('h04)
	) name4067 (
		_w2728_,
		_w2731_,
		_w2732_,
		_w5968_
	);
	LUT4 #(
		.INIT('h1101)
	) name4068 (
		_w2722_,
		_w2726_,
		_w2727_,
		_w2728_,
		_w5969_
	);
	LUT4 #(
		.INIT('h0002)
	) name4069 (
		\m2_s7_cyc_o_reg/NET0131 ,
		\rf_conf7_reg[4]/NET0131 ,
		\rf_conf7_reg[5]/NET0131 ,
		\s7_msel_arb0_state_reg[0]/NET0131 ,
		_w5970_
	);
	LUT4 #(
		.INIT('h00b0)
	) name4070 (
		_w2722_,
		_w2725_,
		_w2750_,
		_w5970_,
		_w5971_
	);
	LUT3 #(
		.INIT('hb0)
	) name4071 (
		_w5968_,
		_w5969_,
		_w5971_,
		_w5972_
	);
	LUT2 #(
		.INIT('h1)
	) name4072 (
		_w5967_,
		_w5972_,
		_w5973_
	);
	LUT4 #(
		.INIT('h00f2)
	) name4073 (
		_w2722_,
		_w2723_,
		_w2731_,
		_w2732_,
		_w5974_
	);
	LUT3 #(
		.INIT('ha8)
	) name4074 (
		\s7_msel_arb0_state_reg[2]/NET0131 ,
		_w2725_,
		_w2728_,
		_w5975_
	);
	LUT3 #(
		.INIT('h54)
	) name4075 (
		\s7_msel_arb0_state_reg[2]/NET0131 ,
		_w2723_,
		_w2732_,
		_w5976_
	);
	LUT4 #(
		.INIT('h4454)
	) name4076 (
		_w2725_,
		_w2726_,
		_w2727_,
		_w2728_,
		_w5977_
	);
	LUT4 #(
		.INIT('hd0dd)
	) name4077 (
		_w5974_,
		_w5975_,
		_w5976_,
		_w5977_,
		_w5978_
	);
	LUT2 #(
		.INIT('h1)
	) name4078 (
		\s7_msel_arb0_state_reg[0]/NET0131 ,
		\s7_msel_arb0_state_reg[1]/NET0131 ,
		_w5979_
	);
	LUT3 #(
		.INIT('h02)
	) name4079 (
		\s7_msel_arb0_state_reg[0]/NET0131 ,
		\s7_msel_arb0_state_reg[1]/NET0131 ,
		\s7_msel_arb0_state_reg[2]/NET0131 ,
		_w5980_
	);
	LUT2 #(
		.INIT('h4)
	) name4080 (
		_w2731_,
		_w5980_,
		_w5981_
	);
	LUT4 #(
		.INIT('h8a00)
	) name4081 (
		_w5960_,
		_w5965_,
		_w5969_,
		_w5981_,
		_w5982_
	);
	LUT4 #(
		.INIT('h0001)
	) name4082 (
		_w2723_,
		_w2725_,
		_w2732_,
		_w5953_,
		_w5983_
	);
	LUT3 #(
		.INIT('h40)
	) name4083 (
		\s7_msel_arb0_state_reg[0]/NET0131 ,
		\s7_msel_arb0_state_reg[1]/NET0131 ,
		\s7_msel_arb0_state_reg[2]/NET0131 ,
		_w5984_
	);
	LUT2 #(
		.INIT('h4)
	) name4084 (
		_w2728_,
		_w5984_,
		_w5985_
	);
	LUT4 #(
		.INIT('hf100)
	) name4085 (
		_w5950_,
		_w5951_,
		_w5983_,
		_w5985_,
		_w5986_
	);
	LUT4 #(
		.INIT('h000b)
	) name4086 (
		_w5978_,
		_w5979_,
		_w5982_,
		_w5986_,
		_w5987_
	);
	LUT3 #(
		.INIT('hbf)
	) name4087 (
		_w5964_,
		_w5973_,
		_w5987_,
		_w5988_
	);
	LUT2 #(
		.INIT('h2)
	) name4088 (
		_w3867_,
		_w3868_,
		_w5989_
	);
	LUT3 #(
		.INIT('h51)
	) name4089 (
		_w3864_,
		_w3867_,
		_w3868_,
		_w5990_
	);
	LUT3 #(
		.INIT('h04)
	) name4090 (
		_w3868_,
		_w3871_,
		_w3872_,
		_w5991_
	);
	LUT3 #(
		.INIT('h51)
	) name4091 (
		_w3865_,
		_w5990_,
		_w5991_,
		_w5992_
	);
	LUT4 #(
		.INIT('h0001)
	) name4092 (
		_w3865_,
		_w3868_,
		_w3872_,
		_w3875_,
		_w5993_
	);
	LUT3 #(
		.INIT('h02)
	) name4093 (
		\s7_msel_arb1_state_reg[2]/NET0131 ,
		_w3874_,
		_w5993_,
		_w5994_
	);
	LUT4 #(
		.INIT('h00f7)
	) name4094 (
		\m3_s7_cyc_o_reg/NET0131 ,
		\rf_conf7_reg[6]/NET0131 ,
		\rf_conf7_reg[7]/NET0131 ,
		\s7_msel_arb1_state_reg[2]/NET0131 ,
		_w5995_
	);
	LUT2 #(
		.INIT('h2)
	) name4095 (
		_w3886_,
		_w5995_,
		_w5996_
	);
	LUT4 #(
		.INIT('hf700)
	) name4096 (
		\m0_s7_cyc_o_reg/NET0131 ,
		\rf_conf7_reg[0]/NET0131 ,
		\rf_conf7_reg[1]/NET0131 ,
		\s7_msel_arb1_state_reg[0]/NET0131 ,
		_w5997_
	);
	LUT2 #(
		.INIT('h4)
	) name4097 (
		_w3868_,
		_w5997_,
		_w5998_
	);
	LUT2 #(
		.INIT('h1)
	) name4098 (
		_w3871_,
		_w3874_,
		_w5999_
	);
	LUT4 #(
		.INIT('h000d)
	) name4099 (
		_w3864_,
		_w3865_,
		_w3871_,
		_w3874_,
		_w6000_
	);
	LUT3 #(
		.INIT('h23)
	) name4100 (
		_w3871_,
		_w3872_,
		_w3875_,
		_w6001_
	);
	LUT4 #(
		.INIT('h2300)
	) name4101 (
		_w3871_,
		_w3872_,
		_w3875_,
		_w3886_,
		_w6002_
	);
	LUT4 #(
		.INIT('h1055)
	) name4102 (
		_w5996_,
		_w5998_,
		_w6000_,
		_w6002_,
		_w6003_
	);
	LUT3 #(
		.INIT('h0b)
	) name4103 (
		_w5992_,
		_w5994_,
		_w6003_,
		_w6004_
	);
	LUT3 #(
		.INIT('h01)
	) name4104 (
		_w3868_,
		_w3872_,
		_w3875_,
		_w6005_
	);
	LUT2 #(
		.INIT('h1)
	) name4105 (
		_w3874_,
		_w5997_,
		_w6006_
	);
	LUT4 #(
		.INIT('h2202)
	) name4106 (
		_w5990_,
		_w5991_,
		_w6005_,
		_w6006_,
		_w6007_
	);
	LUT2 #(
		.INIT('h1)
	) name4107 (
		\s7_msel_arb1_state_reg[1]/NET0131 ,
		\s7_msel_arb1_state_reg[2]/NET0131 ,
		_w6008_
	);
	LUT3 #(
		.INIT('h02)
	) name4108 (
		\s7_msel_arb1_state_reg[0]/NET0131 ,
		\s7_msel_arb1_state_reg[1]/NET0131 ,
		\s7_msel_arb1_state_reg[2]/NET0131 ,
		_w6009_
	);
	LUT4 #(
		.INIT('h2232)
	) name4109 (
		_w3864_,
		_w3865_,
		_w3867_,
		_w3868_,
		_w6010_
	);
	LUT3 #(
		.INIT('h10)
	) name4110 (
		_w3868_,
		_w3872_,
		_w5997_,
		_w6011_
	);
	LUT2 #(
		.INIT('h4)
	) name4111 (
		\s7_msel_arb1_state_reg[1]/NET0131 ,
		\s7_msel_arb1_state_reg[2]/NET0131 ,
		_w6012_
	);
	LUT3 #(
		.INIT('h20)
	) name4112 (
		\s7_msel_arb1_state_reg[0]/NET0131 ,
		\s7_msel_arb1_state_reg[1]/NET0131 ,
		\s7_msel_arb1_state_reg[2]/NET0131 ,
		_w6013_
	);
	LUT3 #(
		.INIT('hb0)
	) name4113 (
		_w3871_,
		_w3875_,
		_w6013_,
		_w6014_
	);
	LUT4 #(
		.INIT('hfd00)
	) name4114 (
		_w5999_,
		_w6010_,
		_w6011_,
		_w6014_,
		_w6015_
	);
	LUT3 #(
		.INIT('h0b)
	) name4115 (
		_w6007_,
		_w6009_,
		_w6015_,
		_w6016_
	);
	LUT3 #(
		.INIT('h20)
	) name4116 (
		\s7_msel_arb1_state_reg[0]/NET0131 ,
		_w6004_,
		_w6016_,
		_w6017_
	);
	LUT3 #(
		.INIT('h54)
	) name4117 (
		_w3868_,
		_w3871_,
		_w3874_,
		_w6018_
	);
	LUT4 #(
		.INIT('h5444)
	) name4118 (
		\s7_msel_arb1_state_reg[2]/NET0131 ,
		_w5989_,
		_w6001_,
		_w6018_,
		_w6019_
	);
	LUT2 #(
		.INIT('h8)
	) name4119 (
		\s7_msel_arb1_state_reg[1]/NET0131 ,
		_w6019_,
		_w6020_
	);
	LUT4 #(
		.INIT('h0800)
	) name4120 (
		\m7_s7_cyc_o_reg/NET0131 ,
		\rf_conf7_reg[14]/NET0131 ,
		\rf_conf7_reg[15]/NET0131 ,
		\s7_msel_arb1_state_reg[2]/NET0131 ,
		_w6021_
	);
	LUT4 #(
		.INIT('hf700)
	) name4121 (
		\m0_s7_cyc_o_reg/NET0131 ,
		\rf_conf7_reg[0]/NET0131 ,
		\rf_conf7_reg[1]/NET0131 ,
		\s7_msel_arb1_state_reg[2]/NET0131 ,
		_w6022_
	);
	LUT4 #(
		.INIT('h020f)
	) name4122 (
		_w5990_,
		_w5991_,
		_w6021_,
		_w6022_,
		_w6023_
	);
	LUT3 #(
		.INIT('hf1)
	) name4123 (
		\s7_msel_arb1_state_reg[0]/NET0131 ,
		_w3864_,
		_w3865_,
		_w6024_
	);
	LUT3 #(
		.INIT('h01)
	) name4124 (
		\s7_msel_arb1_state_reg[2]/NET0131 ,
		_w3868_,
		_w3872_,
		_w6025_
	);
	LUT2 #(
		.INIT('h4)
	) name4125 (
		_w6024_,
		_w6025_,
		_w6026_
	);
	LUT4 #(
		.INIT('hf700)
	) name4126 (
		\m6_s7_cyc_o_reg/NET0131 ,
		\rf_conf7_reg[12]/NET0131 ,
		\rf_conf7_reg[13]/NET0131 ,
		\s7_msel_arb1_state_reg[1]/NET0131 ,
		_w6027_
	);
	LUT3 #(
		.INIT('hd0)
	) name4127 (
		_w6023_,
		_w6026_,
		_w6027_,
		_w6028_
	);
	LUT2 #(
		.INIT('h1)
	) name4128 (
		_w6020_,
		_w6028_,
		_w6029_
	);
	LUT4 #(
		.INIT('h0203)
	) name4129 (
		_w3868_,
		_w3871_,
		_w3874_,
		_w5997_,
		_w6030_
	);
	LUT4 #(
		.INIT('h2300)
	) name4130 (
		_w3871_,
		_w3872_,
		_w3875_,
		_w6012_,
		_w6031_
	);
	LUT3 #(
		.INIT('hb0)
	) name4131 (
		_w6010_,
		_w6030_,
		_w6031_,
		_w6032_
	);
	LUT2 #(
		.INIT('h4)
	) name4132 (
		_w3865_,
		_w6008_,
		_w6033_
	);
	LUT4 #(
		.INIT('hd500)
	) name4133 (
		_w5990_,
		_w6001_,
		_w6018_,
		_w6033_,
		_w6034_
	);
	LUT2 #(
		.INIT('h1)
	) name4134 (
		_w6032_,
		_w6034_,
		_w6035_
	);
	LUT3 #(
		.INIT('h40)
	) name4135 (
		_w6004_,
		_w6016_,
		_w6035_,
		_w6036_
	);
	LUT3 #(
		.INIT('h15)
	) name4136 (
		_w6017_,
		_w6029_,
		_w6036_,
		_w6037_
	);
	LUT3 #(
		.INIT('h20)
	) name4137 (
		\m2_s7_cyc_o_reg/NET0131 ,
		\rf_conf7_reg[4]/NET0131 ,
		\rf_conf7_reg[5]/NET0131 ,
		_w6038_
	);
	LUT3 #(
		.INIT('h20)
	) name4138 (
		\m3_s7_cyc_o_reg/NET0131 ,
		\rf_conf7_reg[6]/NET0131 ,
		\rf_conf7_reg[7]/NET0131 ,
		_w6039_
	);
	LUT2 #(
		.INIT('h2)
	) name4139 (
		\s7_msel_arb2_state_reg[1]/NET0131 ,
		\s7_msel_arb2_state_reg[2]/NET0131 ,
		_w6040_
	);
	LUT3 #(
		.INIT('h40)
	) name4140 (
		_w6038_,
		_w6039_,
		_w6040_,
		_w6041_
	);
	LUT3 #(
		.INIT('h20)
	) name4141 (
		\m5_s7_cyc_o_reg/NET0131 ,
		\rf_conf7_reg[10]/NET0131 ,
		\rf_conf7_reg[11]/NET0131 ,
		_w6042_
	);
	LUT3 #(
		.INIT('h20)
	) name4142 (
		\m7_s7_cyc_o_reg/NET0131 ,
		\rf_conf7_reg[14]/NET0131 ,
		\rf_conf7_reg[15]/NET0131 ,
		_w6043_
	);
	LUT3 #(
		.INIT('h20)
	) name4143 (
		\m6_s7_cyc_o_reg/NET0131 ,
		\rf_conf7_reg[12]/NET0131 ,
		\rf_conf7_reg[13]/NET0131 ,
		_w6044_
	);
	LUT3 #(
		.INIT('h51)
	) name4144 (
		_w6042_,
		_w6043_,
		_w6044_,
		_w6045_
	);
	LUT3 #(
		.INIT('h20)
	) name4145 (
		\m1_s7_cyc_o_reg/NET0131 ,
		\rf_conf7_reg[2]/NET0131 ,
		\rf_conf7_reg[3]/NET0131 ,
		_w6046_
	);
	LUT3 #(
		.INIT('h20)
	) name4146 (
		\m0_s7_cyc_o_reg/NET0131 ,
		\rf_conf7_reg[0]/NET0131 ,
		\rf_conf7_reg[1]/NET0131 ,
		_w6047_
	);
	LUT2 #(
		.INIT('h1)
	) name4147 (
		_w6044_,
		_w6047_,
		_w6048_
	);
	LUT3 #(
		.INIT('h04)
	) name4148 (
		_w6044_,
		_w6046_,
		_w6047_,
		_w6049_
	);
	LUT3 #(
		.INIT('h20)
	) name4149 (
		\m4_s7_cyc_o_reg/NET0131 ,
		\rf_conf7_reg[8]/NET0131 ,
		\rf_conf7_reg[9]/NET0131 ,
		_w6050_
	);
	LUT2 #(
		.INIT('h1)
	) name4150 (
		_w6038_,
		_w6050_,
		_w6051_
	);
	LUT3 #(
		.INIT('h04)
	) name4151 (
		_w6038_,
		_w6040_,
		_w6050_,
		_w6052_
	);
	LUT4 #(
		.INIT('h0455)
	) name4152 (
		_w6041_,
		_w6045_,
		_w6049_,
		_w6052_,
		_w6053_
	);
	LUT3 #(
		.INIT('h0b)
	) name4153 (
		_w6038_,
		_w6039_,
		_w6046_,
		_w6054_
	);
	LUT2 #(
		.INIT('h1)
	) name4154 (
		\s7_msel_arb2_state_reg[1]/NET0131 ,
		\s7_msel_arb2_state_reg[2]/NET0131 ,
		_w6055_
	);
	LUT2 #(
		.INIT('h4)
	) name4155 (
		_w6047_,
		_w6055_,
		_w6056_
	);
	LUT4 #(
		.INIT('hb0ff)
	) name4156 (
		_w6045_,
		_w6051_,
		_w6054_,
		_w6056_,
		_w6057_
	);
	LUT3 #(
		.INIT('h40)
	) name4157 (
		\s7_msel_arb2_state_reg[0]/NET0131 ,
		_w6053_,
		_w6057_,
		_w6058_
	);
	LUT2 #(
		.INIT('h8)
	) name4158 (
		\s7_msel_arb2_state_reg[1]/NET0131 ,
		\s7_msel_arb2_state_reg[2]/NET0131 ,
		_w6059_
	);
	LUT3 #(
		.INIT('h20)
	) name4159 (
		_w6043_,
		_w6044_,
		_w6059_,
		_w6060_
	);
	LUT3 #(
		.INIT('h04)
	) name4160 (
		_w6038_,
		_w6042_,
		_w6050_,
		_w6061_
	);
	LUT3 #(
		.INIT('h10)
	) name4161 (
		_w6044_,
		_w6047_,
		_w6059_,
		_w6062_
	);
	LUT4 #(
		.INIT('h0233)
	) name4162 (
		_w6054_,
		_w6060_,
		_w6061_,
		_w6062_,
		_w6063_
	);
	LUT2 #(
		.INIT('h4)
	) name4163 (
		\s7_msel_arb2_state_reg[1]/NET0131 ,
		\s7_msel_arb2_state_reg[2]/NET0131 ,
		_w6064_
	);
	LUT3 #(
		.INIT('h20)
	) name4164 (
		_w6042_,
		_w6050_,
		_w6064_,
		_w6065_
	);
	LUT2 #(
		.INIT('h4)
	) name4165 (
		_w6043_,
		_w6047_,
		_w6066_
	);
	LUT4 #(
		.INIT('h000b)
	) name4166 (
		_w6038_,
		_w6039_,
		_w6043_,
		_w6046_,
		_w6067_
	);
	LUT3 #(
		.INIT('h10)
	) name4167 (
		_w6044_,
		_w6050_,
		_w6064_,
		_w6068_
	);
	LUT4 #(
		.INIT('h5455)
	) name4168 (
		_w6065_,
		_w6066_,
		_w6067_,
		_w6068_,
		_w6069_
	);
	LUT2 #(
		.INIT('h8)
	) name4169 (
		_w6063_,
		_w6069_,
		_w6070_
	);
	LUT4 #(
		.INIT('hdf00)
	) name4170 (
		\m0_s7_cyc_o_reg/NET0131 ,
		\rf_conf7_reg[0]/NET0131 ,
		\rf_conf7_reg[1]/NET0131 ,
		\s7_msel_arb2_state_reg[0]/NET0131 ,
		_w6071_
	);
	LUT3 #(
		.INIT('h10)
	) name4171 (
		_w6038_,
		_w6050_,
		_w6071_,
		_w6072_
	);
	LUT3 #(
		.INIT('h20)
	) name4172 (
		\s7_msel_arb2_state_reg[0]/NET0131 ,
		\s7_msel_arb2_state_reg[1]/NET0131 ,
		\s7_msel_arb2_state_reg[2]/NET0131 ,
		_w6073_
	);
	LUT3 #(
		.INIT('h10)
	) name4173 (
		_w6042_,
		_w6044_,
		_w6073_,
		_w6074_
	);
	LUT4 #(
		.INIT('hf100)
	) name4174 (
		_w6066_,
		_w6067_,
		_w6072_,
		_w6074_,
		_w6075_
	);
	LUT3 #(
		.INIT('h08)
	) name4175 (
		_w6058_,
		_w6070_,
		_w6075_,
		_w6076_
	);
	LUT3 #(
		.INIT('hb0)
	) name4176 (
		_w6045_,
		_w6051_,
		_w6054_,
		_w6077_
	);
	LUT3 #(
		.INIT('h02)
	) name4177 (
		\s7_msel_arb2_state_reg[0]/NET0131 ,
		_w6038_,
		_w6050_,
		_w6078_
	);
	LUT2 #(
		.INIT('h8)
	) name4178 (
		_w6048_,
		_w6078_,
		_w6079_
	);
	LUT3 #(
		.INIT('ha2)
	) name4179 (
		_w6055_,
		_w6077_,
		_w6079_,
		_w6080_
	);
	LUT2 #(
		.INIT('h8)
	) name4180 (
		_w6039_,
		_w6040_,
		_w6081_
	);
	LUT4 #(
		.INIT('h0031)
	) name4181 (
		_w6038_,
		_w6044_,
		_w6046_,
		_w6047_,
		_w6082_
	);
	LUT2 #(
		.INIT('h2)
	) name4182 (
		_w6040_,
		_w6050_,
		_w6083_
	);
	LUT4 #(
		.INIT('h0233)
	) name4183 (
		_w6045_,
		_w6081_,
		_w6082_,
		_w6083_,
		_w6084_
	);
	LUT3 #(
		.INIT('h2a)
	) name4184 (
		\s7_msel_arb2_state_reg[0]/NET0131 ,
		_w6042_,
		_w6064_,
		_w6085_
	);
	LUT2 #(
		.INIT('h8)
	) name4185 (
		_w6084_,
		_w6085_,
		_w6086_
	);
	LUT4 #(
		.INIT('hdf00)
	) name4186 (
		\m6_s7_cyc_o_reg/NET0131 ,
		\rf_conf7_reg[12]/NET0131 ,
		\rf_conf7_reg[13]/NET0131 ,
		\s7_msel_arb2_state_reg[0]/NET0131 ,
		_w6087_
	);
	LUT4 #(
		.INIT('h3233)
	) name4187 (
		_w6038_,
		_w6043_,
		_w6050_,
		_w6087_,
		_w6088_
	);
	LUT4 #(
		.INIT('h0d0f)
	) name4188 (
		_w6054_,
		_w6061_,
		_w6066_,
		_w6088_,
		_w6089_
	);
	LUT3 #(
		.INIT('h13)
	) name4189 (
		_w6059_,
		_w6075_,
		_w6089_,
		_w6090_
	);
	LUT3 #(
		.INIT('h40)
	) name4190 (
		_w6080_,
		_w6086_,
		_w6090_,
		_w6091_
	);
	LUT2 #(
		.INIT('h1)
	) name4191 (
		_w6076_,
		_w6091_,
		_w6092_
	);
	LUT2 #(
		.INIT('h2)
	) name4192 (
		\s7_msel_arb3_state_reg[1]/NET0131 ,
		\s7_msel_arb3_state_reg[2]/NET0131 ,
		_w6093_
	);
	LUT2 #(
		.INIT('h4)
	) name4193 (
		_w3485_,
		_w6093_,
		_w6094_
	);
	LUT2 #(
		.INIT('h1)
	) name4194 (
		_w3467_,
		_w3474_,
		_w6095_
	);
	LUT3 #(
		.INIT('hae)
	) name4195 (
		_w3467_,
		_w3474_,
		_w3475_,
		_w6096_
	);
	LUT2 #(
		.INIT('h1)
	) name4196 (
		_w3479_,
		_w3490_,
		_w6097_
	);
	LUT2 #(
		.INIT('h1)
	) name4197 (
		_w3475_,
		_w3480_,
		_w6098_
	);
	LUT4 #(
		.INIT('h7577)
	) name4198 (
		_w6094_,
		_w6096_,
		_w6097_,
		_w6098_,
		_w6099_
	);
	LUT3 #(
		.INIT('h0d)
	) name4199 (
		_w3477_,
		_w3478_,
		_w3479_,
		_w6100_
	);
	LUT4 #(
		.INIT('h00f2)
	) name4200 (
		_w3477_,
		_w3478_,
		_w3479_,
		_w3480_,
		_w6101_
	);
	LUT3 #(
		.INIT('h10)
	) name4201 (
		\s7_msel_arb3_state_reg[0]/NET0131 ,
		\s7_msel_arb3_state_reg[1]/NET0131 ,
		\s7_msel_arb3_state_reg[2]/NET0131 ,
		_w6102_
	);
	LUT4 #(
		.INIT('h2300)
	) name4202 (
		_w3467_,
		_w3468_,
		_w3475_,
		_w6102_,
		_w6103_
	);
	LUT3 #(
		.INIT('hd0)
	) name4203 (
		_w6095_,
		_w6101_,
		_w6103_,
		_w6104_
	);
	LUT3 #(
		.INIT('h0e)
	) name4204 (
		_w3468_,
		_w6099_,
		_w6104_,
		_w6105_
	);
	LUT2 #(
		.INIT('h1)
	) name4205 (
		\s7_msel_arb3_state_reg[1]/NET0131 ,
		\s7_msel_arb3_state_reg[2]/NET0131 ,
		_w6106_
	);
	LUT4 #(
		.INIT('h0080)
	) name4206 (
		\m0_s7_cyc_o_reg/NET0131 ,
		\rf_conf7_reg[0]/NET0131 ,
		\rf_conf7_reg[1]/NET0131 ,
		\s7_msel_arb3_state_reg[0]/NET0131 ,
		_w6107_
	);
	LUT2 #(
		.INIT('h2)
	) name4207 (
		_w6106_,
		_w6107_,
		_w6108_
	);
	LUT2 #(
		.INIT('h1)
	) name4208 (
		_w3468_,
		_w3478_,
		_w6109_
	);
	LUT4 #(
		.INIT('h4fcf)
	) name4209 (
		_w6096_,
		_w6100_,
		_w6108_,
		_w6109_,
		_w6110_
	);
	LUT3 #(
		.INIT('h20)
	) name4210 (
		_w3477_,
		_w3485_,
		_w6093_,
		_w6111_
	);
	LUT3 #(
		.INIT('h20)
	) name4211 (
		\s7_msel_arb3_state_reg[0]/NET0131 ,
		\s7_msel_arb3_state_reg[1]/NET0131 ,
		\s7_msel_arb3_state_reg[2]/NET0131 ,
		_w6112_
	);
	LUT2 #(
		.INIT('h8)
	) name4212 (
		_w3467_,
		_w6112_,
		_w6113_
	);
	LUT2 #(
		.INIT('h1)
	) name4213 (
		_w6111_,
		_w6113_,
		_w6114_
	);
	LUT2 #(
		.INIT('h8)
	) name4214 (
		_w6110_,
		_w6114_,
		_w6115_
	);
	LUT3 #(
		.INIT('h02)
	) name4215 (
		\s7_msel_arb3_state_reg[0]/NET0131 ,
		\s7_msel_arb3_state_reg[1]/NET0131 ,
		\s7_msel_arb3_state_reg[2]/NET0131 ,
		_w6116_
	);
	LUT4 #(
		.INIT('h0100)
	) name4216 (
		_w3468_,
		_w3478_,
		_w3480_,
		_w6116_,
		_w6117_
	);
	LUT2 #(
		.INIT('h4)
	) name4217 (
		_w3467_,
		_w6112_,
		_w6118_
	);
	LUT2 #(
		.INIT('h1)
	) name4218 (
		_w6117_,
		_w6118_,
		_w6119_
	);
	LUT2 #(
		.INIT('h4)
	) name4219 (
		_w3474_,
		_w3480_,
		_w6120_
	);
	LUT4 #(
		.INIT('h0051)
	) name4220 (
		_w3474_,
		_w3477_,
		_w3478_,
		_w3479_,
		_w6121_
	);
	LUT4 #(
		.INIT('h7f00)
	) name4221 (
		\m0_s7_cyc_o_reg/NET0131 ,
		\rf_conf7_reg[0]/NET0131 ,
		\rf_conf7_reg[1]/NET0131 ,
		\s7_msel_arb3_state_reg[0]/NET0131 ,
		_w6122_
	);
	LUT3 #(
		.INIT('h10)
	) name4222 (
		_w3468_,
		_w3478_,
		_w6122_,
		_w6123_
	);
	LUT4 #(
		.INIT('h0054)
	) name4223 (
		_w6117_,
		_w6120_,
		_w6121_,
		_w6123_,
		_w6124_
	);
	LUT3 #(
		.INIT('h01)
	) name4224 (
		_w3475_,
		_w6119_,
		_w6124_,
		_w6125_
	);
	LUT4 #(
		.INIT('h007f)
	) name4225 (
		\m5_s7_cyc_o_reg/NET0131 ,
		\rf_conf7_reg[10]/NET0131 ,
		\rf_conf7_reg[11]/NET0131 ,
		\s7_msel_arb3_state_reg[0]/NET0131 ,
		_w6126_
	);
	LUT4 #(
		.INIT('h0001)
	) name4226 (
		_w3468_,
		_w3478_,
		_w3480_,
		_w6126_,
		_w6127_
	);
	LUT3 #(
		.INIT('h0e)
	) name4227 (
		_w6120_,
		_w6121_,
		_w6127_,
		_w6128_
	);
	LUT4 #(
		.INIT('h0080)
	) name4228 (
		\m6_s7_cyc_o_reg/NET0131 ,
		\rf_conf7_reg[12]/NET0131 ,
		\rf_conf7_reg[13]/NET0131 ,
		\s7_msel_arb3_state_reg[0]/NET0131 ,
		_w6129_
	);
	LUT3 #(
		.INIT('h10)
	) name4229 (
		_w3467_,
		_w3474_,
		_w3475_,
		_w6130_
	);
	LUT4 #(
		.INIT('h020a)
	) name4230 (
		_w3493_,
		_w6100_,
		_w6129_,
		_w6130_,
		_w6131_
	);
	LUT2 #(
		.INIT('h4)
	) name4231 (
		_w6128_,
		_w6131_,
		_w6132_
	);
	LUT4 #(
		.INIT('hfff7)
	) name4232 (
		_w6105_,
		_w6115_,
		_w6125_,
		_w6132_,
		_w6133_
	);
	LUT2 #(
		.INIT('h4)
	) name4233 (
		_w2612_,
		_w2620_,
		_w6134_
	);
	LUT3 #(
		.INIT('h04)
	) name4234 (
		_w2608_,
		_w2610_,
		_w2611_,
		_w6135_
	);
	LUT4 #(
		.INIT('hfd00)
	) name4235 (
		\m4_s8_cyc_o_reg/NET0131 ,
		\rf_conf8_reg[8]/NET0131 ,
		\rf_conf8_reg[9]/NET0131 ,
		\s8_msel_arb0_state_reg[0]/NET0131 ,
		_w6136_
	);
	LUT3 #(
		.INIT('h10)
	) name4236 (
		_w2611_,
		_w2613_,
		_w6136_,
		_w6137_
	);
	LUT3 #(
		.INIT('hf2)
	) name4237 (
		_w2607_,
		_w2608_,
		_w2615_,
		_w6138_
	);
	LUT4 #(
		.INIT('h000d)
	) name4238 (
		_w2607_,
		_w2608_,
		_w2612_,
		_w2615_,
		_w6139_
	);
	LUT4 #(
		.INIT('h5455)
	) name4239 (
		_w6134_,
		_w6135_,
		_w6137_,
		_w6139_,
		_w6140_
	);
	LUT2 #(
		.INIT('h8)
	) name4240 (
		_w2634_,
		_w6140_,
		_w6141_
	);
	LUT2 #(
		.INIT('h8)
	) name4241 (
		\s8_msel_arb0_state_reg[1]/NET0131 ,
		\s8_msel_arb0_state_reg[2]/NET0131 ,
		_w6142_
	);
	LUT2 #(
		.INIT('h2)
	) name4242 (
		_w2615_,
		_w2620_,
		_w6143_
	);
	LUT3 #(
		.INIT('h51)
	) name4243 (
		_w2612_,
		_w2615_,
		_w2620_,
		_w6144_
	);
	LUT4 #(
		.INIT('h2232)
	) name4244 (
		_w2612_,
		_w2613_,
		_w2615_,
		_w2620_,
		_w6145_
	);
	LUT2 #(
		.INIT('h1)
	) name4245 (
		_w2608_,
		_w2620_,
		_w6146_
	);
	LUT4 #(
		.INIT('h00fd)
	) name4246 (
		\m5_s8_cyc_o_reg/NET0131 ,
		\rf_conf8_reg[10]/NET0131 ,
		\rf_conf8_reg[11]/NET0131 ,
		\s8_msel_arb0_state_reg[0]/NET0131 ,
		_w6147_
	);
	LUT3 #(
		.INIT('h01)
	) name4247 (
		_w2608_,
		_w2620_,
		_w6147_,
		_w6148_
	);
	LUT2 #(
		.INIT('h4)
	) name4248 (
		_w2607_,
		_w2611_,
		_w6149_
	);
	LUT3 #(
		.INIT('h0b)
	) name4249 (
		_w2607_,
		_w2611_,
		_w2613_,
		_w6150_
	);
	LUT4 #(
		.INIT('h0111)
	) name4250 (
		_w2610_,
		_w6145_,
		_w6148_,
		_w6150_,
		_w6151_
	);
	LUT4 #(
		.INIT('h1101)
	) name4251 (
		_w2607_,
		_w2610_,
		_w2612_,
		_w2613_,
		_w6152_
	);
	LUT4 #(
		.INIT('hfd00)
	) name4252 (
		\m2_s8_cyc_o_reg/NET0131 ,
		\rf_conf8_reg[4]/NET0131 ,
		\rf_conf8_reg[5]/NET0131 ,
		\s8_msel_arb0_state_reg[0]/NET0131 ,
		_w6153_
	);
	LUT4 #(
		.INIT('h0e0f)
	) name4253 (
		_w2611_,
		_w2613_,
		_w2615_,
		_w6153_,
		_w6154_
	);
	LUT2 #(
		.INIT('h2)
	) name4254 (
		\s8_msel_arb0_state_reg[1]/NET0131 ,
		\s8_msel_arb0_state_reg[2]/NET0131 ,
		_w6155_
	);
	LUT3 #(
		.INIT('hd0)
	) name4255 (
		_w2608_,
		_w2615_,
		_w6155_,
		_w6156_
	);
	LUT4 #(
		.INIT('h1f00)
	) name4256 (
		_w6149_,
		_w6152_,
		_w6154_,
		_w6156_,
		_w6157_
	);
	LUT3 #(
		.INIT('h0d)
	) name4257 (
		_w6142_,
		_w6151_,
		_w6157_,
		_w6158_
	);
	LUT3 #(
		.INIT('h8a)
	) name4258 (
		\s8_msel_arb0_state_reg[0]/NET0131 ,
		_w6141_,
		_w6158_,
		_w6159_
	);
	LUT3 #(
		.INIT('h02)
	) name4259 (
		\s8_msel_arb0_state_reg[0]/NET0131 ,
		_w2611_,
		_w2613_,
		_w6160_
	);
	LUT4 #(
		.INIT('h55fd)
	) name4260 (
		_w6146_,
		_w6149_,
		_w6152_,
		_w6160_,
		_w6161_
	);
	LUT3 #(
		.INIT('h8c)
	) name4261 (
		_w6143_,
		_w6155_,
		_w6161_,
		_w6162_
	);
	LUT3 #(
		.INIT('h20)
	) name4262 (
		_w2610_,
		_w2611_,
		_w6142_,
		_w6163_
	);
	LUT3 #(
		.INIT('h10)
	) name4263 (
		_w2611_,
		_w2613_,
		_w6142_,
		_w6164_
	);
	LUT4 #(
		.INIT('h020f)
	) name4264 (
		_w6144_,
		_w6148_,
		_w6163_,
		_w6164_,
		_w6165_
	);
	LUT3 #(
		.INIT('h20)
	) name4265 (
		_w2612_,
		_w2613_,
		_w2634_,
		_w6166_
	);
	LUT2 #(
		.INIT('h1)
	) name4266 (
		_w2608_,
		_w2611_,
		_w6167_
	);
	LUT4 #(
		.INIT('h00fd)
	) name4267 (
		\m7_s8_cyc_o_reg/NET0131 ,
		\rf_conf8_reg[14]/NET0131 ,
		\rf_conf8_reg[15]/NET0131 ,
		\s8_msel_arb0_state_reg[0]/NET0131 ,
		_w6168_
	);
	LUT3 #(
		.INIT('h01)
	) name4268 (
		_w2608_,
		_w2611_,
		_w6168_,
		_w6169_
	);
	LUT3 #(
		.INIT('h10)
	) name4269 (
		_w2613_,
		_w2620_,
		_w2634_,
		_w6170_
	);
	LUT4 #(
		.INIT('h0133)
	) name4270 (
		_w6138_,
		_w6166_,
		_w6169_,
		_w6170_,
		_w6171_
	);
	LUT2 #(
		.INIT('h8)
	) name4271 (
		_w6165_,
		_w6171_,
		_w6172_
	);
	LUT3 #(
		.INIT('h02)
	) name4272 (
		\s8_msel_arb0_state_reg[0]/NET0131 ,
		_w2613_,
		_w2620_,
		_w6173_
	);
	LUT3 #(
		.INIT('h80)
	) name4273 (
		_w2637_,
		_w6167_,
		_w6173_,
		_w6174_
	);
	LUT3 #(
		.INIT('h04)
	) name4274 (
		_w2613_,
		_w2615_,
		_w2620_,
		_w6175_
	);
	LUT4 #(
		.INIT('h0002)
	) name4275 (
		\m4_s8_cyc_o_reg/NET0131 ,
		\rf_conf8_reg[8]/NET0131 ,
		\rf_conf8_reg[9]/NET0131 ,
		\s8_msel_arb0_state_reg[0]/NET0131 ,
		_w6176_
	);
	LUT4 #(
		.INIT('h00b0)
	) name4276 (
		_w2607_,
		_w2611_,
		_w2637_,
		_w6176_,
		_w6177_
	);
	LUT3 #(
		.INIT('hd0)
	) name4277 (
		_w6152_,
		_w6175_,
		_w6177_,
		_w6178_
	);
	LUT2 #(
		.INIT('h1)
	) name4278 (
		_w6174_,
		_w6178_,
		_w6179_
	);
	LUT4 #(
		.INIT('hba00)
	) name4279 (
		\s8_msel_arb0_state_reg[0]/NET0131 ,
		_w6162_,
		_w6172_,
		_w6179_,
		_w6180_
	);
	LUT2 #(
		.INIT('hb)
	) name4280 (
		_w6159_,
		_w6180_,
		_w6181_
	);
	LUT3 #(
		.INIT('hf2)
	) name4281 (
		_w3896_,
		_w3897_,
		_w3900_,
		_w6182_
	);
	LUT4 #(
		.INIT('h0008)
	) name4282 (
		\m4_s8_cyc_o_reg/NET0131 ,
		\rf_conf8_reg[8]/NET0131 ,
		\rf_conf8_reg[9]/NET0131 ,
		\s8_msel_arb1_state_reg[0]/NET0131 ,
		_w6183_
	);
	LUT2 #(
		.INIT('h2)
	) name4283 (
		_w3906_,
		_w6183_,
		_w6184_
	);
	LUT2 #(
		.INIT('h8)
	) name4284 (
		_w6182_,
		_w6184_,
		_w6185_
	);
	LUT3 #(
		.INIT('hf2)
	) name4285 (
		_w3890_,
		_w3891_,
		_w3894_,
		_w6186_
	);
	LUT3 #(
		.INIT('h02)
	) name4286 (
		\s8_msel_arb1_state_reg[0]/NET0131 ,
		_w3891_,
		_w3899_,
		_w6187_
	);
	LUT2 #(
		.INIT('h1)
	) name4287 (
		_w3893_,
		_w3897_,
		_w6188_
	);
	LUT4 #(
		.INIT('h0010)
	) name4288 (
		_w3893_,
		_w3897_,
		_w3906_,
		_w6183_,
		_w6189_
	);
	LUT3 #(
		.INIT('he0)
	) name4289 (
		_w6186_,
		_w6187_,
		_w6189_,
		_w6190_
	);
	LUT4 #(
		.INIT('h0031)
	) name4290 (
		_w3891_,
		_w3893_,
		_w3894_,
		_w3897_,
		_w6191_
	);
	LUT4 #(
		.INIT('h4445)
	) name4291 (
		_w3890_,
		_w3899_,
		_w6182_,
		_w6191_,
		_w6192_
	);
	LUT3 #(
		.INIT('h08)
	) name4292 (
		\s8_msel_arb1_state_reg[0]/NET0131 ,
		\s8_msel_arb1_state_reg[1]/NET0131 ,
		\s8_msel_arb1_state_reg[2]/NET0131 ,
		_w6193_
	);
	LUT4 #(
		.INIT('h0001)
	) name4293 (
		_w3890_,
		_w3894_,
		_w3896_,
		_w3900_,
		_w6194_
	);
	LUT2 #(
		.INIT('h4)
	) name4294 (
		_w3891_,
		_w3909_,
		_w6195_
	);
	LUT3 #(
		.INIT('h45)
	) name4295 (
		_w6193_,
		_w6194_,
		_w6195_,
		_w6196_
	);
	LUT4 #(
		.INIT('h1110)
	) name4296 (
		_w6185_,
		_w6190_,
		_w6192_,
		_w6196_,
		_w6197_
	);
	LUT4 #(
		.INIT('h0008)
	) name4297 (
		\m0_s8_cyc_o_reg/NET0131 ,
		\rf_conf8_reg[0]/NET0131 ,
		\rf_conf8_reg[1]/NET0131 ,
		\s8_msel_arb1_state_reg[0]/NET0131 ,
		_w6198_
	);
	LUT4 #(
		.INIT('h00f2)
	) name4298 (
		_w3890_,
		_w3891_,
		_w3894_,
		_w6198_,
		_w6199_
	);
	LUT3 #(
		.INIT('h01)
	) name4299 (
		_w3891_,
		_w3899_,
		_w6198_,
		_w6200_
	);
	LUT3 #(
		.INIT('h13)
	) name4300 (
		_w6182_,
		_w6199_,
		_w6200_,
		_w6201_
	);
	LUT2 #(
		.INIT('h8)
	) name4301 (
		_w6187_,
		_w6188_,
		_w6202_
	);
	LUT3 #(
		.INIT('ha2)
	) name4302 (
		_w3902_,
		_w6201_,
		_w6202_,
		_w6203_
	);
	LUT3 #(
		.INIT('h10)
	) name4303 (
		_w3891_,
		_w3899_,
		_w3900_,
		_w6204_
	);
	LUT3 #(
		.INIT('h54)
	) name4304 (
		_w3893_,
		_w6186_,
		_w6204_,
		_w6205_
	);
	LUT3 #(
		.INIT('h15)
	) name4305 (
		_w3896_,
		_w6187_,
		_w6188_,
		_w6206_
	);
	LUT4 #(
		.INIT('h0008)
	) name4306 (
		\m6_s8_cyc_o_reg/NET0131 ,
		\rf_conf8_reg[12]/NET0131 ,
		\rf_conf8_reg[13]/NET0131 ,
		\s8_msel_arb1_state_reg[0]/NET0131 ,
		_w6207_
	);
	LUT2 #(
		.INIT('h8)
	) name4307 (
		\s8_msel_arb1_state_reg[1]/NET0131 ,
		\s8_msel_arb1_state_reg[2]/NET0131 ,
		_w6208_
	);
	LUT2 #(
		.INIT('h4)
	) name4308 (
		_w6207_,
		_w6208_,
		_w6209_
	);
	LUT3 #(
		.INIT('hb0)
	) name4309 (
		_w6205_,
		_w6206_,
		_w6209_,
		_w6210_
	);
	LUT3 #(
		.INIT('hfd)
	) name4310 (
		_w6197_,
		_w6203_,
		_w6210_,
		_w6211_
	);
	LUT2 #(
		.INIT('h4)
	) name4311 (
		\s8_msel_arb2_state_reg[1]/NET0131 ,
		\s8_msel_arb2_state_reg[2]/NET0131 ,
		_w6212_
	);
	LUT3 #(
		.INIT('h20)
	) name4312 (
		_w3109_,
		_w3110_,
		_w6212_,
		_w6213_
	);
	LUT2 #(
		.INIT('h4)
	) name4313 (
		_w3112_,
		_w3124_,
		_w6214_
	);
	LUT2 #(
		.INIT('h2)
	) name4314 (
		_w3115_,
		_w3117_,
		_w6215_
	);
	LUT4 #(
		.INIT('h0051)
	) name4315 (
		_w3112_,
		_w3115_,
		_w3117_,
		_w3120_,
		_w6216_
	);
	LUT3 #(
		.INIT('h10)
	) name4316 (
		_w3110_,
		_w3111_,
		_w6212_,
		_w6217_
	);
	LUT4 #(
		.INIT('h5455)
	) name4317 (
		_w6213_,
		_w6214_,
		_w6216_,
		_w6217_,
		_w6218_
	);
	LUT2 #(
		.INIT('h1)
	) name4318 (
		\s8_msel_arb2_state_reg[0]/NET0131 ,
		_w6218_,
		_w6219_
	);
	LUT2 #(
		.INIT('h1)
	) name4319 (
		_w3110_,
		_w3117_,
		_w6220_
	);
	LUT3 #(
		.INIT('hf2)
	) name4320 (
		_w3110_,
		_w3115_,
		_w3117_,
		_w6221_
	);
	LUT3 #(
		.INIT('h45)
	) name4321 (
		_w3109_,
		_w3111_,
		_w3112_,
		_w6222_
	);
	LUT3 #(
		.INIT('h04)
	) name4322 (
		_w3111_,
		_w3120_,
		_w3124_,
		_w6223_
	);
	LUT3 #(
		.INIT('h02)
	) name4323 (
		\s8_msel_arb2_state_reg[0]/NET0131 ,
		_w3111_,
		_w3124_,
		_w6224_
	);
	LUT4 #(
		.INIT('h0004)
	) name4324 (
		_w6215_,
		_w6222_,
		_w6223_,
		_w6224_,
		_w6225_
	);
	LUT3 #(
		.INIT('h04)
	) name4325 (
		\s8_msel_arb2_state_reg[0]/NET0131 ,
		\s8_msel_arb2_state_reg[1]/NET0131 ,
		\s8_msel_arb2_state_reg[2]/NET0131 ,
		_w6226_
	);
	LUT3 #(
		.INIT('h10)
	) name4326 (
		_w6221_,
		_w6225_,
		_w6226_,
		_w6227_
	);
	LUT2 #(
		.INIT('h1)
	) name4327 (
		_w6219_,
		_w6227_,
		_w6228_
	);
	LUT4 #(
		.INIT('hdf00)
	) name4328 (
		\m6_s8_cyc_o_reg/NET0131 ,
		\rf_conf8_reg[12]/NET0131 ,
		\rf_conf8_reg[13]/NET0131 ,
		\s8_msel_arb2_state_reg[0]/NET0131 ,
		_w6229_
	);
	LUT2 #(
		.INIT('h1)
	) name4329 (
		_w3109_,
		_w6229_,
		_w6230_
	);
	LUT3 #(
		.INIT('h01)
	) name4330 (
		_w3110_,
		_w3117_,
		_w3124_,
		_w6231_
	);
	LUT4 #(
		.INIT('he0ee)
	) name4331 (
		_w6214_,
		_w6216_,
		_w6230_,
		_w6231_,
		_w6232_
	);
	LUT4 #(
		.INIT('h0020)
	) name4332 (
		\m6_s8_cyc_o_reg/NET0131 ,
		\rf_conf8_reg[12]/NET0131 ,
		\rf_conf8_reg[13]/NET0131 ,
		\s8_msel_arb2_state_reg[0]/NET0131 ,
		_w6233_
	);
	LUT2 #(
		.INIT('h8)
	) name4333 (
		\s8_msel_arb2_state_reg[1]/NET0131 ,
		\s8_msel_arb2_state_reg[2]/NET0131 ,
		_w6234_
	);
	LUT2 #(
		.INIT('h4)
	) name4334 (
		_w6233_,
		_w6234_,
		_w6235_
	);
	LUT2 #(
		.INIT('h4)
	) name4335 (
		_w6232_,
		_w6235_,
		_w6236_
	);
	LUT3 #(
		.INIT('h51)
	) name4336 (
		_w3110_,
		_w6222_,
		_w6223_,
		_w6237_
	);
	LUT2 #(
		.INIT('h8)
	) name4337 (
		_w6220_,
		_w6224_,
		_w6238_
	);
	LUT3 #(
		.INIT('h15)
	) name4338 (
		_w3115_,
		_w6220_,
		_w6224_,
		_w6239_
	);
	LUT3 #(
		.INIT('h08)
	) name4339 (
		\s8_msel_arb2_state_reg[0]/NET0131 ,
		\s8_msel_arb2_state_reg[1]/NET0131 ,
		\s8_msel_arb2_state_reg[2]/NET0131 ,
		_w6240_
	);
	LUT3 #(
		.INIT('hb0)
	) name4340 (
		_w6237_,
		_w6239_,
		_w6240_,
		_w6241_
	);
	LUT2 #(
		.INIT('h2)
	) name4341 (
		\s8_msel_arb2_state_reg[0]/NET0131 ,
		\s8_msel_arb2_state_reg[1]/NET0131 ,
		_w6242_
	);
	LUT3 #(
		.INIT('h20)
	) name4342 (
		\s8_msel_arb2_state_reg[0]/NET0131 ,
		\s8_msel_arb2_state_reg[1]/NET0131 ,
		\s8_msel_arb2_state_reg[2]/NET0131 ,
		_w6243_
	);
	LUT3 #(
		.INIT('h01)
	) name4343 (
		_w3111_,
		_w6214_,
		_w6216_,
		_w6244_
	);
	LUT3 #(
		.INIT('h15)
	) name4344 (
		_w3109_,
		_w6220_,
		_w6224_,
		_w6245_
	);
	LUT3 #(
		.INIT('h8a)
	) name4345 (
		_w6243_,
		_w6244_,
		_w6245_,
		_w6246_
	);
	LUT4 #(
		.INIT('h0020)
	) name4346 (
		\m0_s8_cyc_o_reg/NET0131 ,
		\rf_conf8_reg[0]/NET0131 ,
		\rf_conf8_reg[1]/NET0131 ,
		\s8_msel_arb2_state_reg[0]/NET0131 ,
		_w6247_
	);
	LUT4 #(
		.INIT('h00f2)
	) name4347 (
		_w3115_,
		_w3117_,
		_w3120_,
		_w6247_,
		_w6248_
	);
	LUT3 #(
		.INIT('h01)
	) name4348 (
		_w3110_,
		_w3117_,
		_w6247_,
		_w6249_
	);
	LUT3 #(
		.INIT('h23)
	) name4349 (
		_w6222_,
		_w6248_,
		_w6249_,
		_w6250_
	);
	LUT2 #(
		.INIT('h1)
	) name4350 (
		\s8_msel_arb2_state_reg[1]/NET0131 ,
		\s8_msel_arb2_state_reg[2]/NET0131 ,
		_w6251_
	);
	LUT3 #(
		.INIT('hb0)
	) name4351 (
		_w6238_,
		_w6250_,
		_w6251_,
		_w6252_
	);
	LUT4 #(
		.INIT('h0001)
	) name4352 (
		_w6236_,
		_w6241_,
		_w6246_,
		_w6252_,
		_w6253_
	);
	LUT2 #(
		.INIT('h7)
	) name4353 (
		_w6228_,
		_w6253_,
		_w6254_
	);
	LUT3 #(
		.INIT('hdc)
	) name4354 (
		_w3500_,
		_w3501_,
		_w3511_,
		_w6255_
	);
	LUT2 #(
		.INIT('h4)
	) name4355 (
		_w3503_,
		_w3505_,
		_w6256_
	);
	LUT4 #(
		.INIT('h000d)
	) name4356 (
		_w3498_,
		_w3499_,
		_w3503_,
		_w3504_,
		_w6257_
	);
	LUT4 #(
		.INIT('h7f00)
	) name4357 (
		\m6_s8_cyc_o_reg/NET0131 ,
		\rf_conf8_reg[12]/NET0131 ,
		\rf_conf8_reg[13]/NET0131 ,
		\s8_msel_arb3_state_reg[0]/NET0131 ,
		_w6258_
	);
	LUT4 #(
		.INIT('ha2f3)
	) name4358 (
		_w3499_,
		_w3500_,
		_w3501_,
		_w6258_,
		_w6259_
	);
	LUT4 #(
		.INIT('h0155)
	) name4359 (
		_w6255_,
		_w6256_,
		_w6257_,
		_w6259_,
		_w6260_
	);
	LUT2 #(
		.INIT('h8)
	) name4360 (
		_w3523_,
		_w6260_,
		_w6261_
	);
	LUT2 #(
		.INIT('h1)
	) name4361 (
		\s8_msel_arb3_state_reg[1]/NET0131 ,
		\s8_msel_arb3_state_reg[2]/NET0131 ,
		_w6262_
	);
	LUT3 #(
		.INIT('h20)
	) name4362 (
		_w3498_,
		_w3499_,
		_w6262_,
		_w6263_
	);
	LUT2 #(
		.INIT('h4)
	) name4363 (
		_w3500_,
		_w3511_,
		_w6264_
	);
	LUT4 #(
		.INIT('h1101)
	) name4364 (
		_w3500_,
		_w3503_,
		_w3504_,
		_w3505_,
		_w6265_
	);
	LUT3 #(
		.INIT('h10)
	) name4365 (
		_w3499_,
		_w3501_,
		_w6262_,
		_w6266_
	);
	LUT4 #(
		.INIT('h5455)
	) name4366 (
		_w6263_,
		_w6264_,
		_w6265_,
		_w6266_,
		_w6267_
	);
	LUT3 #(
		.INIT('h08)
	) name4367 (
		_w3497_,
		_w3503_,
		_w3511_,
		_w6268_
	);
	LUT3 #(
		.INIT('h0d)
	) name4368 (
		_w3498_,
		_w3499_,
		_w3504_,
		_w6269_
	);
	LUT3 #(
		.INIT('h04)
	) name4369 (
		_w3499_,
		_w3500_,
		_w3501_,
		_w6270_
	);
	LUT3 #(
		.INIT('h02)
	) name4370 (
		_w3497_,
		_w3505_,
		_w3511_,
		_w6271_
	);
	LUT4 #(
		.INIT('h0455)
	) name4371 (
		_w6268_,
		_w6269_,
		_w6270_,
		_w6271_,
		_w6272_
	);
	LUT3 #(
		.INIT('h40)
	) name4372 (
		\s8_msel_arb3_state_reg[0]/NET0131 ,
		_w6267_,
		_w6272_,
		_w6273_
	);
	LUT3 #(
		.INIT('h51)
	) name4373 (
		_w3505_,
		_w6269_,
		_w6270_,
		_w6274_
	);
	LUT4 #(
		.INIT('h0001)
	) name4374 (
		_w3499_,
		_w3501_,
		_w3505_,
		_w3511_,
		_w6275_
	);
	LUT2 #(
		.INIT('h1)
	) name4375 (
		_w3503_,
		_w6275_,
		_w6276_
	);
	LUT3 #(
		.INIT('h2a)
	) name4376 (
		\s8_msel_arb3_state_reg[0]/NET0131 ,
		_w3500_,
		_w3523_,
		_w6277_
	);
	LUT4 #(
		.INIT('h7500)
	) name4377 (
		_w3497_,
		_w6274_,
		_w6276_,
		_w6277_,
		_w6278_
	);
	LUT3 #(
		.INIT('h0b)
	) name4378 (
		_w6261_,
		_w6273_,
		_w6278_,
		_w6279_
	);
	LUT2 #(
		.INIT('h4)
	) name4379 (
		_w3498_,
		_w3501_,
		_w6280_
	);
	LUT4 #(
		.INIT('h5455)
	) name4380 (
		_w3498_,
		_w3499_,
		_w3511_,
		_w6258_,
		_w6281_
	);
	LUT4 #(
		.INIT('h010f)
	) name4381 (
		_w6264_,
		_w6265_,
		_w6280_,
		_w6281_,
		_w6282_
	);
	LUT3 #(
		.INIT('h02)
	) name4382 (
		\s8_msel_arb3_state_reg[0]/NET0131 ,
		\s8_msel_arb3_state_reg[1]/NET0131 ,
		\s8_msel_arb3_state_reg[2]/NET0131 ,
		_w6283_
	);
	LUT2 #(
		.INIT('h8)
	) name4383 (
		_w6282_,
		_w6283_,
		_w6284_
	);
	LUT2 #(
		.INIT('h1)
	) name4384 (
		_w3503_,
		_w6258_,
		_w6285_
	);
	LUT3 #(
		.INIT('h01)
	) name4385 (
		_w3499_,
		_w3501_,
		_w3511_,
		_w6286_
	);
	LUT4 #(
		.INIT('h2022)
	) name4386 (
		_w6269_,
		_w6270_,
		_w6285_,
		_w6286_,
		_w6287_
	);
	LUT4 #(
		.INIT('h0080)
	) name4387 (
		\m6_s8_cyc_o_reg/NET0131 ,
		\rf_conf8_reg[12]/NET0131 ,
		\rf_conf8_reg[13]/NET0131 ,
		\s8_msel_arb3_state_reg[0]/NET0131 ,
		_w6288_
	);
	LUT2 #(
		.INIT('h2)
	) name4388 (
		_w3509_,
		_w6288_,
		_w6289_
	);
	LUT3 #(
		.INIT('h10)
	) name4389 (
		_w3499_,
		_w3501_,
		_w6258_,
		_w6290_
	);
	LUT3 #(
		.INIT('h08)
	) name4390 (
		\s8_msel_arb3_state_reg[0]/NET0131 ,
		\s8_msel_arb3_state_reg[1]/NET0131 ,
		\s8_msel_arb3_state_reg[2]/NET0131 ,
		_w6291_
	);
	LUT3 #(
		.INIT('h10)
	) name4391 (
		_w3500_,
		_w3511_,
		_w6291_,
		_w6292_
	);
	LUT4 #(
		.INIT('hf100)
	) name4392 (
		_w6256_,
		_w6257_,
		_w6290_,
		_w6292_,
		_w6293_
	);
	LUT3 #(
		.INIT('h0b)
	) name4393 (
		_w6287_,
		_w6289_,
		_w6293_,
		_w6294_
	);
	LUT2 #(
		.INIT('h4)
	) name4394 (
		_w6284_,
		_w6294_,
		_w6295_
	);
	LUT2 #(
		.INIT('hb)
	) name4395 (
		_w6279_,
		_w6295_,
		_w6296_
	);
	LUT2 #(
		.INIT('h4)
	) name4396 (
		_w2766_,
		_w2771_,
		_w6297_
	);
	LUT4 #(
		.INIT('h000d)
	) name4397 (
		_w2761_,
		_w2762_,
		_w2766_,
		_w2770_,
		_w6298_
	);
	LUT3 #(
		.INIT('h01)
	) name4398 (
		_w2762_,
		_w2764_,
		_w2771_,
		_w6299_
	);
	LUT4 #(
		.INIT('h00fd)
	) name4399 (
		\m5_s9_cyc_o_reg/NET0131 ,
		\rf_conf9_reg[10]/NET0131 ,
		\rf_conf9_reg[11]/NET0131 ,
		\s9_msel_arb0_state_reg[0]/NET0131 ,
		_w6300_
	);
	LUT3 #(
		.INIT('hce)
	) name4400 (
		\s9_msel_arb0_state_reg[0]/NET0131 ,
		_w2765_,
		_w2767_,
		_w6301_
	);
	LUT4 #(
		.INIT('h0eee)
	) name4401 (
		_w6297_,
		_w6298_,
		_w6299_,
		_w6301_,
		_w6302_
	);
	LUT3 #(
		.INIT('hae)
	) name4402 (
		_w2765_,
		_w2766_,
		_w2767_,
		_w6303_
	);
	LUT2 #(
		.INIT('h4)
	) name4403 (
		\s9_msel_arb0_state_reg[1]/NET0131 ,
		\s9_msel_arb0_state_reg[2]/NET0131 ,
		_w6304_
	);
	LUT4 #(
		.INIT('h0002)
	) name4404 (
		\m1_s9_cyc_o_reg/NET0131 ,
		\rf_conf9_reg[2]/NET0131 ,
		\rf_conf9_reg[3]/NET0131 ,
		\s9_msel_arb0_state_reg[1]/NET0131 ,
		_w6305_
	);
	LUT2 #(
		.INIT('h1)
	) name4405 (
		_w6304_,
		_w6305_,
		_w6306_
	);
	LUT3 #(
		.INIT('h23)
	) name4406 (
		_w2761_,
		_w2762_,
		_w2764_,
		_w6307_
	);
	LUT4 #(
		.INIT('h00dc)
	) name4407 (
		_w2761_,
		_w2762_,
		_w2764_,
		_w2770_,
		_w6308_
	);
	LUT3 #(
		.INIT('ha8)
	) name4408 (
		\s9_msel_arb0_state_reg[2]/NET0131 ,
		_w2767_,
		_w2771_,
		_w6309_
	);
	LUT4 #(
		.INIT('hdddc)
	) name4409 (
		_w6303_,
		_w6306_,
		_w6308_,
		_w6309_,
		_w6310_
	);
	LUT4 #(
		.INIT('h08aa)
	) name4410 (
		\s9_msel_arb0_state_reg[0]/NET0131 ,
		_w2794_,
		_w6302_,
		_w6310_,
		_w6311_
	);
	LUT3 #(
		.INIT('h02)
	) name4411 (
		\s9_msel_arb0_state_reg[0]/NET0131 ,
		_w2767_,
		_w2771_,
		_w6312_
	);
	LUT2 #(
		.INIT('h1)
	) name4412 (
		_w2762_,
		_w2764_,
		_w6313_
	);
	LUT3 #(
		.INIT('h80)
	) name4413 (
		_w2789_,
		_w6312_,
		_w6313_,
		_w6314_
	);
	LUT3 #(
		.INIT('h04)
	) name4414 (
		_w2767_,
		_w2770_,
		_w2771_,
		_w6315_
	);
	LUT4 #(
		.INIT('h1101)
	) name4415 (
		_w2761_,
		_w2765_,
		_w2766_,
		_w2767_,
		_w6316_
	);
	LUT4 #(
		.INIT('h0002)
	) name4416 (
		\m2_s9_cyc_o_reg/NET0131 ,
		\rf_conf9_reg[4]/NET0131 ,
		\rf_conf9_reg[5]/NET0131 ,
		\s9_msel_arb0_state_reg[0]/NET0131 ,
		_w6317_
	);
	LUT4 #(
		.INIT('h00b0)
	) name4417 (
		_w2761_,
		_w2764_,
		_w2789_,
		_w6317_,
		_w6318_
	);
	LUT3 #(
		.INIT('hb0)
	) name4418 (
		_w6315_,
		_w6316_,
		_w6318_,
		_w6319_
	);
	LUT2 #(
		.INIT('h1)
	) name4419 (
		_w6314_,
		_w6319_,
		_w6320_
	);
	LUT4 #(
		.INIT('h00f2)
	) name4420 (
		_w2761_,
		_w2762_,
		_w2770_,
		_w2771_,
		_w6321_
	);
	LUT3 #(
		.INIT('ha8)
	) name4421 (
		\s9_msel_arb0_state_reg[2]/NET0131 ,
		_w2764_,
		_w2767_,
		_w6322_
	);
	LUT3 #(
		.INIT('h54)
	) name4422 (
		\s9_msel_arb0_state_reg[2]/NET0131 ,
		_w2762_,
		_w2771_,
		_w6323_
	);
	LUT4 #(
		.INIT('h4454)
	) name4423 (
		_w2764_,
		_w2765_,
		_w2766_,
		_w2767_,
		_w6324_
	);
	LUT4 #(
		.INIT('hd0dd)
	) name4424 (
		_w6321_,
		_w6322_,
		_w6323_,
		_w6324_,
		_w6325_
	);
	LUT2 #(
		.INIT('h1)
	) name4425 (
		\s9_msel_arb0_state_reg[0]/NET0131 ,
		\s9_msel_arb0_state_reg[1]/NET0131 ,
		_w6326_
	);
	LUT3 #(
		.INIT('h02)
	) name4426 (
		\s9_msel_arb0_state_reg[0]/NET0131 ,
		\s9_msel_arb0_state_reg[1]/NET0131 ,
		\s9_msel_arb0_state_reg[2]/NET0131 ,
		_w6327_
	);
	LUT2 #(
		.INIT('h4)
	) name4427 (
		_w2770_,
		_w6327_,
		_w6328_
	);
	LUT4 #(
		.INIT('h8a00)
	) name4428 (
		_w6307_,
		_w6312_,
		_w6316_,
		_w6328_,
		_w6329_
	);
	LUT4 #(
		.INIT('h0001)
	) name4429 (
		_w2762_,
		_w2764_,
		_w2771_,
		_w6300_,
		_w6330_
	);
	LUT3 #(
		.INIT('h40)
	) name4430 (
		\s9_msel_arb0_state_reg[0]/NET0131 ,
		\s9_msel_arb0_state_reg[1]/NET0131 ,
		\s9_msel_arb0_state_reg[2]/NET0131 ,
		_w6331_
	);
	LUT2 #(
		.INIT('h4)
	) name4431 (
		_w2767_,
		_w6331_,
		_w6332_
	);
	LUT4 #(
		.INIT('hf100)
	) name4432 (
		_w6297_,
		_w6298_,
		_w6330_,
		_w6332_,
		_w6333_
	);
	LUT4 #(
		.INIT('h000b)
	) name4433 (
		_w6325_,
		_w6326_,
		_w6329_,
		_w6333_,
		_w6334_
	);
	LUT3 #(
		.INIT('hbf)
	) name4434 (
		_w6311_,
		_w6320_,
		_w6334_,
		_w6335_
	);
	LUT3 #(
		.INIT('hf2)
	) name4435 (
		_w3927_,
		_w3928_,
		_w3931_,
		_w6336_
	);
	LUT4 #(
		.INIT('h0008)
	) name4436 (
		\m4_s9_cyc_o_reg/NET0131 ,
		\rf_conf9_reg[8]/NET0131 ,
		\rf_conf9_reg[9]/NET0131 ,
		\s9_msel_arb1_state_reg[0]/NET0131 ,
		_w6337_
	);
	LUT2 #(
		.INIT('h2)
	) name4437 (
		_w3937_,
		_w6337_,
		_w6338_
	);
	LUT2 #(
		.INIT('h8)
	) name4438 (
		_w6336_,
		_w6338_,
		_w6339_
	);
	LUT3 #(
		.INIT('hf2)
	) name4439 (
		_w3921_,
		_w3922_,
		_w3925_,
		_w6340_
	);
	LUT3 #(
		.INIT('h02)
	) name4440 (
		\s9_msel_arb1_state_reg[0]/NET0131 ,
		_w3922_,
		_w3930_,
		_w6341_
	);
	LUT2 #(
		.INIT('h1)
	) name4441 (
		_w3924_,
		_w3928_,
		_w6342_
	);
	LUT4 #(
		.INIT('h0010)
	) name4442 (
		_w3924_,
		_w3928_,
		_w3937_,
		_w6337_,
		_w6343_
	);
	LUT3 #(
		.INIT('he0)
	) name4443 (
		_w6340_,
		_w6341_,
		_w6343_,
		_w6344_
	);
	LUT4 #(
		.INIT('h0031)
	) name4444 (
		_w3922_,
		_w3924_,
		_w3925_,
		_w3928_,
		_w6345_
	);
	LUT4 #(
		.INIT('h4445)
	) name4445 (
		_w3921_,
		_w3930_,
		_w6336_,
		_w6345_,
		_w6346_
	);
	LUT3 #(
		.INIT('h08)
	) name4446 (
		\s9_msel_arb1_state_reg[0]/NET0131 ,
		\s9_msel_arb1_state_reg[1]/NET0131 ,
		\s9_msel_arb1_state_reg[2]/NET0131 ,
		_w6347_
	);
	LUT4 #(
		.INIT('h0001)
	) name4447 (
		_w3921_,
		_w3925_,
		_w3927_,
		_w3931_,
		_w6348_
	);
	LUT2 #(
		.INIT('h4)
	) name4448 (
		_w3922_,
		_w3940_,
		_w6349_
	);
	LUT3 #(
		.INIT('h45)
	) name4449 (
		_w6347_,
		_w6348_,
		_w6349_,
		_w6350_
	);
	LUT4 #(
		.INIT('h1110)
	) name4450 (
		_w6339_,
		_w6344_,
		_w6346_,
		_w6350_,
		_w6351_
	);
	LUT4 #(
		.INIT('h0008)
	) name4451 (
		\m0_s9_cyc_o_reg/NET0131 ,
		\rf_conf9_reg[0]/NET0131 ,
		\rf_conf9_reg[1]/NET0131 ,
		\s9_msel_arb1_state_reg[0]/NET0131 ,
		_w6352_
	);
	LUT4 #(
		.INIT('h00f2)
	) name4452 (
		_w3921_,
		_w3922_,
		_w3925_,
		_w6352_,
		_w6353_
	);
	LUT3 #(
		.INIT('h01)
	) name4453 (
		_w3922_,
		_w3930_,
		_w6352_,
		_w6354_
	);
	LUT3 #(
		.INIT('h13)
	) name4454 (
		_w6336_,
		_w6353_,
		_w6354_,
		_w6355_
	);
	LUT2 #(
		.INIT('h8)
	) name4455 (
		_w6341_,
		_w6342_,
		_w6356_
	);
	LUT3 #(
		.INIT('ha2)
	) name4456 (
		_w3933_,
		_w6355_,
		_w6356_,
		_w6357_
	);
	LUT3 #(
		.INIT('h10)
	) name4457 (
		_w3922_,
		_w3930_,
		_w3931_,
		_w6358_
	);
	LUT3 #(
		.INIT('h54)
	) name4458 (
		_w3924_,
		_w6340_,
		_w6358_,
		_w6359_
	);
	LUT3 #(
		.INIT('h15)
	) name4459 (
		_w3927_,
		_w6341_,
		_w6342_,
		_w6360_
	);
	LUT4 #(
		.INIT('h0008)
	) name4460 (
		\m6_s9_cyc_o_reg/NET0131 ,
		\rf_conf9_reg[12]/NET0131 ,
		\rf_conf9_reg[13]/NET0131 ,
		\s9_msel_arb1_state_reg[0]/NET0131 ,
		_w6361_
	);
	LUT2 #(
		.INIT('h8)
	) name4461 (
		\s9_msel_arb1_state_reg[1]/NET0131 ,
		\s9_msel_arb1_state_reg[2]/NET0131 ,
		_w6362_
	);
	LUT2 #(
		.INIT('h4)
	) name4462 (
		_w6361_,
		_w6362_,
		_w6363_
	);
	LUT3 #(
		.INIT('hb0)
	) name4463 (
		_w6359_,
		_w6360_,
		_w6363_,
		_w6364_
	);
	LUT3 #(
		.INIT('hfd)
	) name4464 (
		_w6351_,
		_w6357_,
		_w6364_,
		_w6365_
	);
	LUT3 #(
		.INIT('h20)
	) name4465 (
		\m2_s9_cyc_o_reg/NET0131 ,
		\rf_conf9_reg[4]/NET0131 ,
		\rf_conf9_reg[5]/NET0131 ,
		_w6366_
	);
	LUT3 #(
		.INIT('h20)
	) name4466 (
		\m3_s9_cyc_o_reg/NET0131 ,
		\rf_conf9_reg[6]/NET0131 ,
		\rf_conf9_reg[7]/NET0131 ,
		_w6367_
	);
	LUT2 #(
		.INIT('h2)
	) name4467 (
		\s9_msel_arb2_state_reg[1]/NET0131 ,
		\s9_msel_arb2_state_reg[2]/NET0131 ,
		_w6368_
	);
	LUT3 #(
		.INIT('h40)
	) name4468 (
		_w6366_,
		_w6367_,
		_w6368_,
		_w6369_
	);
	LUT3 #(
		.INIT('h20)
	) name4469 (
		\m5_s9_cyc_o_reg/NET0131 ,
		\rf_conf9_reg[10]/NET0131 ,
		\rf_conf9_reg[11]/NET0131 ,
		_w6370_
	);
	LUT3 #(
		.INIT('h20)
	) name4470 (
		\m7_s9_cyc_o_reg/NET0131 ,
		\rf_conf9_reg[14]/NET0131 ,
		\rf_conf9_reg[15]/NET0131 ,
		_w6371_
	);
	LUT3 #(
		.INIT('h20)
	) name4471 (
		\m6_s9_cyc_o_reg/NET0131 ,
		\rf_conf9_reg[12]/NET0131 ,
		\rf_conf9_reg[13]/NET0131 ,
		_w6372_
	);
	LUT3 #(
		.INIT('h51)
	) name4472 (
		_w6370_,
		_w6371_,
		_w6372_,
		_w6373_
	);
	LUT3 #(
		.INIT('h20)
	) name4473 (
		\m1_s9_cyc_o_reg/NET0131 ,
		\rf_conf9_reg[2]/NET0131 ,
		\rf_conf9_reg[3]/NET0131 ,
		_w6374_
	);
	LUT3 #(
		.INIT('h20)
	) name4474 (
		\m0_s9_cyc_o_reg/NET0131 ,
		\rf_conf9_reg[0]/NET0131 ,
		\rf_conf9_reg[1]/NET0131 ,
		_w6375_
	);
	LUT2 #(
		.INIT('h1)
	) name4475 (
		_w6372_,
		_w6375_,
		_w6376_
	);
	LUT3 #(
		.INIT('h04)
	) name4476 (
		_w6372_,
		_w6374_,
		_w6375_,
		_w6377_
	);
	LUT3 #(
		.INIT('h20)
	) name4477 (
		\m4_s9_cyc_o_reg/NET0131 ,
		\rf_conf9_reg[8]/NET0131 ,
		\rf_conf9_reg[9]/NET0131 ,
		_w6378_
	);
	LUT2 #(
		.INIT('h1)
	) name4478 (
		_w6366_,
		_w6378_,
		_w6379_
	);
	LUT3 #(
		.INIT('h04)
	) name4479 (
		_w6366_,
		_w6368_,
		_w6378_,
		_w6380_
	);
	LUT4 #(
		.INIT('h0455)
	) name4480 (
		_w6369_,
		_w6373_,
		_w6377_,
		_w6380_,
		_w6381_
	);
	LUT3 #(
		.INIT('h0b)
	) name4481 (
		_w6366_,
		_w6367_,
		_w6374_,
		_w6382_
	);
	LUT2 #(
		.INIT('h1)
	) name4482 (
		\s9_msel_arb2_state_reg[1]/NET0131 ,
		\s9_msel_arb2_state_reg[2]/NET0131 ,
		_w6383_
	);
	LUT2 #(
		.INIT('h4)
	) name4483 (
		_w6375_,
		_w6383_,
		_w6384_
	);
	LUT4 #(
		.INIT('hb0ff)
	) name4484 (
		_w6373_,
		_w6379_,
		_w6382_,
		_w6384_,
		_w6385_
	);
	LUT3 #(
		.INIT('h40)
	) name4485 (
		\s9_msel_arb2_state_reg[0]/NET0131 ,
		_w6381_,
		_w6385_,
		_w6386_
	);
	LUT2 #(
		.INIT('h8)
	) name4486 (
		\s9_msel_arb2_state_reg[1]/NET0131 ,
		\s9_msel_arb2_state_reg[2]/NET0131 ,
		_w6387_
	);
	LUT3 #(
		.INIT('h20)
	) name4487 (
		_w6371_,
		_w6372_,
		_w6387_,
		_w6388_
	);
	LUT3 #(
		.INIT('h04)
	) name4488 (
		_w6366_,
		_w6370_,
		_w6378_,
		_w6389_
	);
	LUT3 #(
		.INIT('h10)
	) name4489 (
		_w6372_,
		_w6375_,
		_w6387_,
		_w6390_
	);
	LUT4 #(
		.INIT('h0233)
	) name4490 (
		_w6382_,
		_w6388_,
		_w6389_,
		_w6390_,
		_w6391_
	);
	LUT2 #(
		.INIT('h4)
	) name4491 (
		\s9_msel_arb2_state_reg[1]/NET0131 ,
		\s9_msel_arb2_state_reg[2]/NET0131 ,
		_w6392_
	);
	LUT3 #(
		.INIT('h20)
	) name4492 (
		_w6370_,
		_w6378_,
		_w6392_,
		_w6393_
	);
	LUT2 #(
		.INIT('h4)
	) name4493 (
		_w6371_,
		_w6375_,
		_w6394_
	);
	LUT4 #(
		.INIT('h000b)
	) name4494 (
		_w6366_,
		_w6367_,
		_w6371_,
		_w6374_,
		_w6395_
	);
	LUT3 #(
		.INIT('h10)
	) name4495 (
		_w6372_,
		_w6378_,
		_w6392_,
		_w6396_
	);
	LUT4 #(
		.INIT('h5455)
	) name4496 (
		_w6393_,
		_w6394_,
		_w6395_,
		_w6396_,
		_w6397_
	);
	LUT2 #(
		.INIT('h8)
	) name4497 (
		_w6391_,
		_w6397_,
		_w6398_
	);
	LUT4 #(
		.INIT('hdf00)
	) name4498 (
		\m0_s9_cyc_o_reg/NET0131 ,
		\rf_conf9_reg[0]/NET0131 ,
		\rf_conf9_reg[1]/NET0131 ,
		\s9_msel_arb2_state_reg[0]/NET0131 ,
		_w6399_
	);
	LUT3 #(
		.INIT('h10)
	) name4499 (
		_w6366_,
		_w6378_,
		_w6399_,
		_w6400_
	);
	LUT3 #(
		.INIT('h20)
	) name4500 (
		\s9_msel_arb2_state_reg[0]/NET0131 ,
		\s9_msel_arb2_state_reg[1]/NET0131 ,
		\s9_msel_arb2_state_reg[2]/NET0131 ,
		_w6401_
	);
	LUT3 #(
		.INIT('h10)
	) name4501 (
		_w6370_,
		_w6372_,
		_w6401_,
		_w6402_
	);
	LUT4 #(
		.INIT('hf100)
	) name4502 (
		_w6394_,
		_w6395_,
		_w6400_,
		_w6402_,
		_w6403_
	);
	LUT3 #(
		.INIT('h08)
	) name4503 (
		_w6386_,
		_w6398_,
		_w6403_,
		_w6404_
	);
	LUT3 #(
		.INIT('hb0)
	) name4504 (
		_w6373_,
		_w6379_,
		_w6382_,
		_w6405_
	);
	LUT3 #(
		.INIT('h02)
	) name4505 (
		\s9_msel_arb2_state_reg[0]/NET0131 ,
		_w6366_,
		_w6378_,
		_w6406_
	);
	LUT2 #(
		.INIT('h8)
	) name4506 (
		_w6376_,
		_w6406_,
		_w6407_
	);
	LUT3 #(
		.INIT('ha2)
	) name4507 (
		_w6383_,
		_w6405_,
		_w6407_,
		_w6408_
	);
	LUT2 #(
		.INIT('h8)
	) name4508 (
		_w6367_,
		_w6368_,
		_w6409_
	);
	LUT4 #(
		.INIT('h0031)
	) name4509 (
		_w6366_,
		_w6372_,
		_w6374_,
		_w6375_,
		_w6410_
	);
	LUT2 #(
		.INIT('h2)
	) name4510 (
		_w6368_,
		_w6378_,
		_w6411_
	);
	LUT4 #(
		.INIT('h0233)
	) name4511 (
		_w6373_,
		_w6409_,
		_w6410_,
		_w6411_,
		_w6412_
	);
	LUT3 #(
		.INIT('h2a)
	) name4512 (
		\s9_msel_arb2_state_reg[0]/NET0131 ,
		_w6370_,
		_w6392_,
		_w6413_
	);
	LUT2 #(
		.INIT('h8)
	) name4513 (
		_w6412_,
		_w6413_,
		_w6414_
	);
	LUT4 #(
		.INIT('hdf00)
	) name4514 (
		\m6_s9_cyc_o_reg/NET0131 ,
		\rf_conf9_reg[12]/NET0131 ,
		\rf_conf9_reg[13]/NET0131 ,
		\s9_msel_arb2_state_reg[0]/NET0131 ,
		_w6415_
	);
	LUT4 #(
		.INIT('h3233)
	) name4515 (
		_w6366_,
		_w6371_,
		_w6378_,
		_w6415_,
		_w6416_
	);
	LUT4 #(
		.INIT('h0d0f)
	) name4516 (
		_w6382_,
		_w6389_,
		_w6394_,
		_w6416_,
		_w6417_
	);
	LUT3 #(
		.INIT('h13)
	) name4517 (
		_w6387_,
		_w6403_,
		_w6417_,
		_w6418_
	);
	LUT3 #(
		.INIT('h40)
	) name4518 (
		_w6408_,
		_w6414_,
		_w6418_,
		_w6419_
	);
	LUT2 #(
		.INIT('h1)
	) name4519 (
		_w6404_,
		_w6419_,
		_w6420_
	);
	LUT3 #(
		.INIT('h80)
	) name4520 (
		\m4_s9_cyc_o_reg/NET0131 ,
		\rf_conf9_reg[8]/NET0131 ,
		\rf_conf9_reg[9]/NET0131 ,
		_w6421_
	);
	LUT3 #(
		.INIT('h80)
	) name4521 (
		\m7_s9_cyc_o_reg/NET0131 ,
		\rf_conf9_reg[14]/NET0131 ,
		\rf_conf9_reg[15]/NET0131 ,
		_w6422_
	);
	LUT3 #(
		.INIT('h80)
	) name4522 (
		\m0_s9_cyc_o_reg/NET0131 ,
		\rf_conf9_reg[0]/NET0131 ,
		\rf_conf9_reg[1]/NET0131 ,
		_w6423_
	);
	LUT2 #(
		.INIT('h4)
	) name4523 (
		_w6422_,
		_w6423_,
		_w6424_
	);
	LUT3 #(
		.INIT('h80)
	) name4524 (
		\m3_s9_cyc_o_reg/NET0131 ,
		\rf_conf9_reg[6]/NET0131 ,
		\rf_conf9_reg[7]/NET0131 ,
		_w6425_
	);
	LUT3 #(
		.INIT('h80)
	) name4525 (
		\m2_s9_cyc_o_reg/NET0131 ,
		\rf_conf9_reg[4]/NET0131 ,
		\rf_conf9_reg[5]/NET0131 ,
		_w6426_
	);
	LUT3 #(
		.INIT('h80)
	) name4526 (
		\m1_s9_cyc_o_reg/NET0131 ,
		\rf_conf9_reg[2]/NET0131 ,
		\rf_conf9_reg[3]/NET0131 ,
		_w6427_
	);
	LUT4 #(
		.INIT('h0051)
	) name4527 (
		_w6422_,
		_w6425_,
		_w6426_,
		_w6427_,
		_w6428_
	);
	LUT3 #(
		.INIT('h80)
	) name4528 (
		\m5_s9_cyc_o_reg/NET0131 ,
		\rf_conf9_reg[10]/NET0131 ,
		\rf_conf9_reg[11]/NET0131 ,
		_w6429_
	);
	LUT3 #(
		.INIT('h80)
	) name4529 (
		\m6_s9_cyc_o_reg/NET0131 ,
		\rf_conf9_reg[12]/NET0131 ,
		\rf_conf9_reg[13]/NET0131 ,
		_w6430_
	);
	LUT3 #(
		.INIT('h8a)
	) name4530 (
		\s9_msel_arb3_state_reg[0]/NET0131 ,
		_w6429_,
		_w6430_,
		_w6431_
	);
	LUT4 #(
		.INIT('hf100)
	) name4531 (
		_w6424_,
		_w6428_,
		_w6429_,
		_w6431_,
		_w6432_
	);
	LUT2 #(
		.INIT('h1)
	) name4532 (
		_w6423_,
		_w6430_,
		_w6433_
	);
	LUT4 #(
		.INIT('h7f00)
	) name4533 (
		\m2_s9_cyc_o_reg/NET0131 ,
		\rf_conf9_reg[4]/NET0131 ,
		\rf_conf9_reg[5]/NET0131 ,
		\s9_msel_arb3_state_reg[0]/NET0131 ,
		_w6434_
	);
	LUT4 #(
		.INIT('h3030)
	) name4534 (
		_w6423_,
		_w6429_,
		_w6430_,
		_w6434_,
		_w6435_
	);
	LUT4 #(
		.INIT('h3233)
	) name4535 (
		_w6423_,
		_w6429_,
		_w6430_,
		_w6434_,
		_w6436_
	);
	LUT4 #(
		.INIT('h010f)
	) name4536 (
		_w6424_,
		_w6428_,
		_w6435_,
		_w6436_,
		_w6437_
	);
	LUT2 #(
		.INIT('h4)
	) name4537 (
		\s9_msel_arb3_state_reg[1]/NET0131 ,
		\s9_msel_arb3_state_reg[2]/NET0131 ,
		_w6438_
	);
	LUT4 #(
		.INIT('hd000)
	) name4538 (
		_w6421_,
		_w6432_,
		_w6437_,
		_w6438_,
		_w6439_
	);
	LUT2 #(
		.INIT('h8)
	) name4539 (
		\s9_msel_arb3_state_reg[1]/NET0131 ,
		\s9_msel_arb3_state_reg[2]/NET0131 ,
		_w6440_
	);
	LUT3 #(
		.INIT('h20)
	) name4540 (
		_w6422_,
		_w6430_,
		_w6440_,
		_w6441_
	);
	LUT3 #(
		.INIT('h0d)
	) name4541 (
		_w6425_,
		_w6426_,
		_w6427_,
		_w6442_
	);
	LUT4 #(
		.INIT('h007f)
	) name4542 (
		\m5_s9_cyc_o_reg/NET0131 ,
		\rf_conf9_reg[10]/NET0131 ,
		\rf_conf9_reg[11]/NET0131 ,
		\s9_msel_arb3_state_reg[0]/NET0131 ,
		_w6443_
	);
	LUT3 #(
		.INIT('h01)
	) name4543 (
		_w6421_,
		_w6426_,
		_w6443_,
		_w6444_
	);
	LUT3 #(
		.INIT('h10)
	) name4544 (
		_w6423_,
		_w6430_,
		_w6440_,
		_w6445_
	);
	LUT4 #(
		.INIT('h0455)
	) name4545 (
		_w6441_,
		_w6442_,
		_w6444_,
		_w6445_,
		_w6446_
	);
	LUT2 #(
		.INIT('h1)
	) name4546 (
		\s9_msel_arb3_state_reg[1]/NET0131 ,
		\s9_msel_arb3_state_reg[2]/NET0131 ,
		_w6447_
	);
	LUT3 #(
		.INIT('h40)
	) name4547 (
		_w6423_,
		_w6427_,
		_w6447_,
		_w6448_
	);
	LUT2 #(
		.INIT('h2)
	) name4548 (
		_w6421_,
		_w6425_,
		_w6449_
	);
	LUT4 #(
		.INIT('h0301)
	) name4549 (
		_w6422_,
		_w6425_,
		_w6429_,
		_w6430_,
		_w6450_
	);
	LUT3 #(
		.INIT('h10)
	) name4550 (
		_w6423_,
		_w6426_,
		_w6447_,
		_w6451_
	);
	LUT4 #(
		.INIT('h5455)
	) name4551 (
		_w6448_,
		_w6449_,
		_w6450_,
		_w6451_,
		_w6452_
	);
	LUT3 #(
		.INIT('h15)
	) name4552 (
		\s9_msel_arb3_state_reg[0]/NET0131 ,
		_w6446_,
		_w6452_,
		_w6453_
	);
	LUT3 #(
		.INIT('h80)
	) name4553 (
		\s9_msel_arb3_state_reg[0]/NET0131 ,
		_w6427_,
		_w6447_,
		_w6454_
	);
	LUT3 #(
		.INIT('h45)
	) name4554 (
		_w6423_,
		_w6429_,
		_w6430_,
		_w6455_
	);
	LUT4 #(
		.INIT('h0eee)
	) name4555 (
		_w6424_,
		_w6428_,
		_w6444_,
		_w6455_,
		_w6456_
	);
	LUT3 #(
		.INIT('h80)
	) name4556 (
		\s9_msel_arb3_state_reg[0]/NET0131 ,
		\s9_msel_arb3_state_reg[1]/NET0131 ,
		\s9_msel_arb3_state_reg[2]/NET0131 ,
		_w6457_
	);
	LUT3 #(
		.INIT('h45)
	) name4557 (
		_w6454_,
		_w6456_,
		_w6457_,
		_w6458_
	);
	LUT3 #(
		.INIT('h40)
	) name4558 (
		_w6427_,
		_w6434_,
		_w6447_,
		_w6459_
	);
	LUT4 #(
		.INIT('h0080)
	) name4559 (
		\m2_s9_cyc_o_reg/NET0131 ,
		\rf_conf9_reg[4]/NET0131 ,
		\rf_conf9_reg[5]/NET0131 ,
		\s9_msel_arb3_state_reg[0]/NET0131 ,
		_w6460_
	);
	LUT2 #(
		.INIT('h2)
	) name4560 (
		\s9_msel_arb3_state_reg[1]/NET0131 ,
		\s9_msel_arb3_state_reg[2]/NET0131 ,
		_w6461_
	);
	LUT2 #(
		.INIT('h4)
	) name4561 (
		_w6460_,
		_w6461_,
		_w6462_
	);
	LUT4 #(
		.INIT('h1110)
	) name4562 (
		_w6449_,
		_w6450_,
		_w6459_,
		_w6462_,
		_w6463_
	);
	LUT3 #(
		.INIT('h40)
	) name4563 (
		_w6421_,
		_w6433_,
		_w6459_,
		_w6464_
	);
	LUT4 #(
		.INIT('hfafb)
	) name4564 (
		_w6423_,
		_w6427_,
		_w6430_,
		_w6434_,
		_w6465_
	);
	LUT3 #(
		.INIT('h10)
	) name4565 (
		_w6421_,
		_w6460_,
		_w6461_,
		_w6466_
	);
	LUT2 #(
		.INIT('h4)
	) name4566 (
		_w6465_,
		_w6466_,
		_w6467_
	);
	LUT3 #(
		.INIT('h01)
	) name4567 (
		_w6463_,
		_w6464_,
		_w6467_,
		_w6468_
	);
	LUT4 #(
		.INIT('hefff)
	) name4568 (
		_w6439_,
		_w6453_,
		_w6458_,
		_w6468_,
		_w6469_
	);
	LUT2 #(
		.INIT('h4)
	) name4569 (
		_w2805_,
		_w2810_,
		_w6470_
	);
	LUT4 #(
		.INIT('h000d)
	) name4570 (
		_w2800_,
		_w2801_,
		_w2805_,
		_w2809_,
		_w6471_
	);
	LUT3 #(
		.INIT('h01)
	) name4571 (
		_w2801_,
		_w2803_,
		_w2810_,
		_w6472_
	);
	LUT4 #(
		.INIT('h00fd)
	) name4572 (
		\m5_s0_cyc_o_reg/NET0131 ,
		\rf_conf0_reg[10]/NET0131 ,
		\rf_conf0_reg[11]/NET0131 ,
		\s0_msel_arb0_state_reg[0]/NET0131 ,
		_w6473_
	);
	LUT3 #(
		.INIT('hce)
	) name4573 (
		\s0_msel_arb0_state_reg[0]/NET0131 ,
		_w2804_,
		_w2806_,
		_w6474_
	);
	LUT4 #(
		.INIT('h0eee)
	) name4574 (
		_w6470_,
		_w6471_,
		_w6472_,
		_w6474_,
		_w6475_
	);
	LUT3 #(
		.INIT('hae)
	) name4575 (
		_w2804_,
		_w2805_,
		_w2806_,
		_w6476_
	);
	LUT2 #(
		.INIT('h4)
	) name4576 (
		\s0_msel_arb0_state_reg[1]/NET0131 ,
		\s0_msel_arb0_state_reg[2]/NET0131 ,
		_w6477_
	);
	LUT4 #(
		.INIT('h0002)
	) name4577 (
		\m1_s0_cyc_o_reg/NET0131 ,
		\rf_conf0_reg[2]/NET0131 ,
		\rf_conf0_reg[3]/NET0131 ,
		\s0_msel_arb0_state_reg[1]/NET0131 ,
		_w6478_
	);
	LUT2 #(
		.INIT('h1)
	) name4578 (
		_w6477_,
		_w6478_,
		_w6479_
	);
	LUT3 #(
		.INIT('h23)
	) name4579 (
		_w2800_,
		_w2801_,
		_w2803_,
		_w6480_
	);
	LUT4 #(
		.INIT('h00dc)
	) name4580 (
		_w2800_,
		_w2801_,
		_w2803_,
		_w2809_,
		_w6481_
	);
	LUT3 #(
		.INIT('ha8)
	) name4581 (
		\s0_msel_arb0_state_reg[2]/NET0131 ,
		_w2806_,
		_w2810_,
		_w6482_
	);
	LUT4 #(
		.INIT('hdddc)
	) name4582 (
		_w6476_,
		_w6479_,
		_w6481_,
		_w6482_,
		_w6483_
	);
	LUT4 #(
		.INIT('h08aa)
	) name4583 (
		\s0_msel_arb0_state_reg[0]/NET0131 ,
		_w2833_,
		_w6475_,
		_w6483_,
		_w6484_
	);
	LUT3 #(
		.INIT('h02)
	) name4584 (
		\s0_msel_arb0_state_reg[0]/NET0131 ,
		_w2806_,
		_w2810_,
		_w6485_
	);
	LUT2 #(
		.INIT('h1)
	) name4585 (
		_w2801_,
		_w2803_,
		_w6486_
	);
	LUT3 #(
		.INIT('h80)
	) name4586 (
		_w2828_,
		_w6485_,
		_w6486_,
		_w6487_
	);
	LUT3 #(
		.INIT('h04)
	) name4587 (
		_w2806_,
		_w2809_,
		_w2810_,
		_w6488_
	);
	LUT4 #(
		.INIT('h1101)
	) name4588 (
		_w2800_,
		_w2804_,
		_w2805_,
		_w2806_,
		_w6489_
	);
	LUT4 #(
		.INIT('h0002)
	) name4589 (
		\m2_s0_cyc_o_reg/NET0131 ,
		\rf_conf0_reg[4]/NET0131 ,
		\rf_conf0_reg[5]/NET0131 ,
		\s0_msel_arb0_state_reg[0]/NET0131 ,
		_w6490_
	);
	LUT4 #(
		.INIT('h00b0)
	) name4590 (
		_w2800_,
		_w2803_,
		_w2828_,
		_w6490_,
		_w6491_
	);
	LUT3 #(
		.INIT('hb0)
	) name4591 (
		_w6488_,
		_w6489_,
		_w6491_,
		_w6492_
	);
	LUT2 #(
		.INIT('h1)
	) name4592 (
		_w6487_,
		_w6492_,
		_w6493_
	);
	LUT4 #(
		.INIT('h00f2)
	) name4593 (
		_w2800_,
		_w2801_,
		_w2809_,
		_w2810_,
		_w6494_
	);
	LUT3 #(
		.INIT('ha8)
	) name4594 (
		\s0_msel_arb0_state_reg[2]/NET0131 ,
		_w2803_,
		_w2806_,
		_w6495_
	);
	LUT3 #(
		.INIT('h54)
	) name4595 (
		\s0_msel_arb0_state_reg[2]/NET0131 ,
		_w2801_,
		_w2810_,
		_w6496_
	);
	LUT4 #(
		.INIT('h4454)
	) name4596 (
		_w2803_,
		_w2804_,
		_w2805_,
		_w2806_,
		_w6497_
	);
	LUT4 #(
		.INIT('hd0dd)
	) name4597 (
		_w6494_,
		_w6495_,
		_w6496_,
		_w6497_,
		_w6498_
	);
	LUT2 #(
		.INIT('h1)
	) name4598 (
		\s0_msel_arb0_state_reg[0]/NET0131 ,
		\s0_msel_arb0_state_reg[1]/NET0131 ,
		_w6499_
	);
	LUT3 #(
		.INIT('h02)
	) name4599 (
		\s0_msel_arb0_state_reg[0]/NET0131 ,
		\s0_msel_arb0_state_reg[1]/NET0131 ,
		\s0_msel_arb0_state_reg[2]/NET0131 ,
		_w6500_
	);
	LUT2 #(
		.INIT('h4)
	) name4600 (
		_w2809_,
		_w6500_,
		_w6501_
	);
	LUT4 #(
		.INIT('h8a00)
	) name4601 (
		_w6480_,
		_w6485_,
		_w6489_,
		_w6501_,
		_w6502_
	);
	LUT4 #(
		.INIT('h0001)
	) name4602 (
		_w2801_,
		_w2803_,
		_w2810_,
		_w6473_,
		_w6503_
	);
	LUT3 #(
		.INIT('h40)
	) name4603 (
		\s0_msel_arb0_state_reg[0]/NET0131 ,
		\s0_msel_arb0_state_reg[1]/NET0131 ,
		\s0_msel_arb0_state_reg[2]/NET0131 ,
		_w6504_
	);
	LUT2 #(
		.INIT('h4)
	) name4604 (
		_w2806_,
		_w6504_,
		_w6505_
	);
	LUT4 #(
		.INIT('hf100)
	) name4605 (
		_w6470_,
		_w6471_,
		_w6503_,
		_w6505_,
		_w6506_
	);
	LUT4 #(
		.INIT('h000b)
	) name4606 (
		_w6498_,
		_w6499_,
		_w6502_,
		_w6506_,
		_w6507_
	);
	LUT3 #(
		.INIT('hbf)
	) name4607 (
		_w6484_,
		_w6493_,
		_w6507_,
		_w6508_
	);
	LUT3 #(
		.INIT('hf2)
	) name4608 (
		_w3958_,
		_w3959_,
		_w3962_,
		_w6509_
	);
	LUT4 #(
		.INIT('h0008)
	) name4609 (
		\m4_s0_cyc_o_reg/NET0131 ,
		\rf_conf0_reg[8]/NET0131 ,
		\rf_conf0_reg[9]/NET0131 ,
		\s0_msel_arb1_state_reg[0]/NET0131 ,
		_w6510_
	);
	LUT2 #(
		.INIT('h2)
	) name4610 (
		_w3968_,
		_w6510_,
		_w6511_
	);
	LUT2 #(
		.INIT('h8)
	) name4611 (
		_w6509_,
		_w6511_,
		_w6512_
	);
	LUT3 #(
		.INIT('hf2)
	) name4612 (
		_w3952_,
		_w3953_,
		_w3956_,
		_w6513_
	);
	LUT3 #(
		.INIT('h02)
	) name4613 (
		\s0_msel_arb1_state_reg[0]/NET0131 ,
		_w3953_,
		_w3961_,
		_w6514_
	);
	LUT2 #(
		.INIT('h1)
	) name4614 (
		_w3955_,
		_w3959_,
		_w6515_
	);
	LUT4 #(
		.INIT('h0010)
	) name4615 (
		_w3955_,
		_w3959_,
		_w3968_,
		_w6510_,
		_w6516_
	);
	LUT3 #(
		.INIT('he0)
	) name4616 (
		_w6513_,
		_w6514_,
		_w6516_,
		_w6517_
	);
	LUT4 #(
		.INIT('h0031)
	) name4617 (
		_w3953_,
		_w3955_,
		_w3956_,
		_w3959_,
		_w6518_
	);
	LUT4 #(
		.INIT('h4445)
	) name4618 (
		_w3952_,
		_w3961_,
		_w6509_,
		_w6518_,
		_w6519_
	);
	LUT3 #(
		.INIT('h08)
	) name4619 (
		\s0_msel_arb1_state_reg[0]/NET0131 ,
		\s0_msel_arb1_state_reg[1]/NET0131 ,
		\s0_msel_arb1_state_reg[2]/NET0131 ,
		_w6520_
	);
	LUT4 #(
		.INIT('h0001)
	) name4620 (
		_w3952_,
		_w3956_,
		_w3958_,
		_w3962_,
		_w6521_
	);
	LUT2 #(
		.INIT('h4)
	) name4621 (
		_w3953_,
		_w3971_,
		_w6522_
	);
	LUT3 #(
		.INIT('h45)
	) name4622 (
		_w6520_,
		_w6521_,
		_w6522_,
		_w6523_
	);
	LUT4 #(
		.INIT('h1110)
	) name4623 (
		_w6512_,
		_w6517_,
		_w6519_,
		_w6523_,
		_w6524_
	);
	LUT4 #(
		.INIT('h0008)
	) name4624 (
		\m0_s0_cyc_o_reg/NET0131 ,
		\rf_conf0_reg[0]/NET0131 ,
		\rf_conf0_reg[1]/NET0131 ,
		\s0_msel_arb1_state_reg[0]/NET0131 ,
		_w6525_
	);
	LUT4 #(
		.INIT('h00f2)
	) name4625 (
		_w3952_,
		_w3953_,
		_w3956_,
		_w6525_,
		_w6526_
	);
	LUT3 #(
		.INIT('h01)
	) name4626 (
		_w3953_,
		_w3961_,
		_w6525_,
		_w6527_
	);
	LUT3 #(
		.INIT('h13)
	) name4627 (
		_w6509_,
		_w6526_,
		_w6527_,
		_w6528_
	);
	LUT2 #(
		.INIT('h8)
	) name4628 (
		_w6514_,
		_w6515_,
		_w6529_
	);
	LUT3 #(
		.INIT('ha2)
	) name4629 (
		_w3964_,
		_w6528_,
		_w6529_,
		_w6530_
	);
	LUT3 #(
		.INIT('h10)
	) name4630 (
		_w3953_,
		_w3961_,
		_w3962_,
		_w6531_
	);
	LUT3 #(
		.INIT('h54)
	) name4631 (
		_w3955_,
		_w6513_,
		_w6531_,
		_w6532_
	);
	LUT3 #(
		.INIT('h15)
	) name4632 (
		_w3958_,
		_w6514_,
		_w6515_,
		_w6533_
	);
	LUT4 #(
		.INIT('h0008)
	) name4633 (
		\m6_s0_cyc_o_reg/NET0131 ,
		\rf_conf0_reg[12]/NET0131 ,
		\rf_conf0_reg[13]/NET0131 ,
		\s0_msel_arb1_state_reg[0]/NET0131 ,
		_w6534_
	);
	LUT2 #(
		.INIT('h8)
	) name4634 (
		\s0_msel_arb1_state_reg[1]/NET0131 ,
		\s0_msel_arb1_state_reg[2]/NET0131 ,
		_w6535_
	);
	LUT2 #(
		.INIT('h4)
	) name4635 (
		_w6534_,
		_w6535_,
		_w6536_
	);
	LUT3 #(
		.INIT('hb0)
	) name4636 (
		_w6532_,
		_w6533_,
		_w6536_,
		_w6537_
	);
	LUT3 #(
		.INIT('hfd)
	) name4637 (
		_w6524_,
		_w6530_,
		_w6537_,
		_w6538_
	);
	LUT2 #(
		.INIT('h4)
	) name4638 (
		\s0_msel_arb2_state_reg[1]/NET0131 ,
		\s0_msel_arb2_state_reg[2]/NET0131 ,
		_w6539_
	);
	LUT3 #(
		.INIT('h20)
	) name4639 (
		_w3131_,
		_w3132_,
		_w6539_,
		_w6540_
	);
	LUT2 #(
		.INIT('h4)
	) name4640 (
		_w3134_,
		_w3146_,
		_w6541_
	);
	LUT2 #(
		.INIT('h2)
	) name4641 (
		_w3137_,
		_w3139_,
		_w6542_
	);
	LUT4 #(
		.INIT('h0051)
	) name4642 (
		_w3134_,
		_w3137_,
		_w3139_,
		_w3142_,
		_w6543_
	);
	LUT3 #(
		.INIT('h10)
	) name4643 (
		_w3132_,
		_w3133_,
		_w6539_,
		_w6544_
	);
	LUT4 #(
		.INIT('h5455)
	) name4644 (
		_w6540_,
		_w6541_,
		_w6543_,
		_w6544_,
		_w6545_
	);
	LUT2 #(
		.INIT('h1)
	) name4645 (
		\s0_msel_arb2_state_reg[0]/NET0131 ,
		_w6545_,
		_w6546_
	);
	LUT2 #(
		.INIT('h1)
	) name4646 (
		_w3132_,
		_w3139_,
		_w6547_
	);
	LUT3 #(
		.INIT('hf2)
	) name4647 (
		_w3132_,
		_w3137_,
		_w3139_,
		_w6548_
	);
	LUT3 #(
		.INIT('h45)
	) name4648 (
		_w3131_,
		_w3133_,
		_w3134_,
		_w6549_
	);
	LUT3 #(
		.INIT('h04)
	) name4649 (
		_w3133_,
		_w3142_,
		_w3146_,
		_w6550_
	);
	LUT3 #(
		.INIT('h02)
	) name4650 (
		\s0_msel_arb2_state_reg[0]/NET0131 ,
		_w3133_,
		_w3146_,
		_w6551_
	);
	LUT4 #(
		.INIT('h0004)
	) name4651 (
		_w6542_,
		_w6549_,
		_w6550_,
		_w6551_,
		_w6552_
	);
	LUT3 #(
		.INIT('h04)
	) name4652 (
		\s0_msel_arb2_state_reg[0]/NET0131 ,
		\s0_msel_arb2_state_reg[1]/NET0131 ,
		\s0_msel_arb2_state_reg[2]/NET0131 ,
		_w6553_
	);
	LUT3 #(
		.INIT('h10)
	) name4653 (
		_w6548_,
		_w6552_,
		_w6553_,
		_w6554_
	);
	LUT2 #(
		.INIT('h1)
	) name4654 (
		_w6546_,
		_w6554_,
		_w6555_
	);
	LUT4 #(
		.INIT('hdf00)
	) name4655 (
		\m6_s0_cyc_o_reg/NET0131 ,
		\rf_conf0_reg[12]/NET0131 ,
		\rf_conf0_reg[13]/NET0131 ,
		\s0_msel_arb2_state_reg[0]/NET0131 ,
		_w6556_
	);
	LUT2 #(
		.INIT('h1)
	) name4656 (
		_w3131_,
		_w6556_,
		_w6557_
	);
	LUT3 #(
		.INIT('h01)
	) name4657 (
		_w3132_,
		_w3139_,
		_w3146_,
		_w6558_
	);
	LUT4 #(
		.INIT('he0ee)
	) name4658 (
		_w6541_,
		_w6543_,
		_w6557_,
		_w6558_,
		_w6559_
	);
	LUT4 #(
		.INIT('h0020)
	) name4659 (
		\m6_s0_cyc_o_reg/NET0131 ,
		\rf_conf0_reg[12]/NET0131 ,
		\rf_conf0_reg[13]/NET0131 ,
		\s0_msel_arb2_state_reg[0]/NET0131 ,
		_w6560_
	);
	LUT2 #(
		.INIT('h8)
	) name4660 (
		\s0_msel_arb2_state_reg[1]/NET0131 ,
		\s0_msel_arb2_state_reg[2]/NET0131 ,
		_w6561_
	);
	LUT2 #(
		.INIT('h4)
	) name4661 (
		_w6560_,
		_w6561_,
		_w6562_
	);
	LUT2 #(
		.INIT('h4)
	) name4662 (
		_w6559_,
		_w6562_,
		_w6563_
	);
	LUT3 #(
		.INIT('h51)
	) name4663 (
		_w3132_,
		_w6549_,
		_w6550_,
		_w6564_
	);
	LUT2 #(
		.INIT('h8)
	) name4664 (
		_w6547_,
		_w6551_,
		_w6565_
	);
	LUT3 #(
		.INIT('h15)
	) name4665 (
		_w3137_,
		_w6547_,
		_w6551_,
		_w6566_
	);
	LUT3 #(
		.INIT('h08)
	) name4666 (
		\s0_msel_arb2_state_reg[0]/NET0131 ,
		\s0_msel_arb2_state_reg[1]/NET0131 ,
		\s0_msel_arb2_state_reg[2]/NET0131 ,
		_w6567_
	);
	LUT3 #(
		.INIT('hb0)
	) name4667 (
		_w6564_,
		_w6566_,
		_w6567_,
		_w6568_
	);
	LUT2 #(
		.INIT('h2)
	) name4668 (
		\s0_msel_arb2_state_reg[0]/NET0131 ,
		\s0_msel_arb2_state_reg[1]/NET0131 ,
		_w6569_
	);
	LUT3 #(
		.INIT('h20)
	) name4669 (
		\s0_msel_arb2_state_reg[0]/NET0131 ,
		\s0_msel_arb2_state_reg[1]/NET0131 ,
		\s0_msel_arb2_state_reg[2]/NET0131 ,
		_w6570_
	);
	LUT3 #(
		.INIT('h01)
	) name4670 (
		_w3133_,
		_w6541_,
		_w6543_,
		_w6571_
	);
	LUT3 #(
		.INIT('h15)
	) name4671 (
		_w3131_,
		_w6547_,
		_w6551_,
		_w6572_
	);
	LUT3 #(
		.INIT('h8a)
	) name4672 (
		_w6570_,
		_w6571_,
		_w6572_,
		_w6573_
	);
	LUT4 #(
		.INIT('h0020)
	) name4673 (
		\m0_s0_cyc_o_reg/NET0131 ,
		\rf_conf0_reg[0]/NET0131 ,
		\rf_conf0_reg[1]/NET0131 ,
		\s0_msel_arb2_state_reg[0]/NET0131 ,
		_w6574_
	);
	LUT4 #(
		.INIT('h00f2)
	) name4674 (
		_w3137_,
		_w3139_,
		_w3142_,
		_w6574_,
		_w6575_
	);
	LUT3 #(
		.INIT('h01)
	) name4675 (
		_w3132_,
		_w3139_,
		_w6574_,
		_w6576_
	);
	LUT3 #(
		.INIT('h23)
	) name4676 (
		_w6549_,
		_w6575_,
		_w6576_,
		_w6577_
	);
	LUT2 #(
		.INIT('h1)
	) name4677 (
		\s0_msel_arb2_state_reg[1]/NET0131 ,
		\s0_msel_arb2_state_reg[2]/NET0131 ,
		_w6578_
	);
	LUT3 #(
		.INIT('hb0)
	) name4678 (
		_w6565_,
		_w6577_,
		_w6578_,
		_w6579_
	);
	LUT4 #(
		.INIT('h0001)
	) name4679 (
		_w6563_,
		_w6568_,
		_w6573_,
		_w6579_,
		_w6580_
	);
	LUT2 #(
		.INIT('h7)
	) name4680 (
		_w6555_,
		_w6580_,
		_w6581_
	);
	LUT2 #(
		.INIT('h2)
	) name4681 (
		\s0_msel_arb3_state_reg[1]/NET0131 ,
		\s0_msel_arb3_state_reg[2]/NET0131 ,
		_w6582_
	);
	LUT2 #(
		.INIT('h4)
	) name4682 (
		_w3547_,
		_w6582_,
		_w6583_
	);
	LUT2 #(
		.INIT('h1)
	) name4683 (
		_w3529_,
		_w3536_,
		_w6584_
	);
	LUT3 #(
		.INIT('hae)
	) name4684 (
		_w3529_,
		_w3536_,
		_w3537_,
		_w6585_
	);
	LUT2 #(
		.INIT('h1)
	) name4685 (
		_w3541_,
		_w3552_,
		_w6586_
	);
	LUT2 #(
		.INIT('h1)
	) name4686 (
		_w3537_,
		_w3542_,
		_w6587_
	);
	LUT4 #(
		.INIT('h7577)
	) name4687 (
		_w6583_,
		_w6585_,
		_w6586_,
		_w6587_,
		_w6588_
	);
	LUT3 #(
		.INIT('h0d)
	) name4688 (
		_w3539_,
		_w3540_,
		_w3541_,
		_w6589_
	);
	LUT4 #(
		.INIT('h00f2)
	) name4689 (
		_w3539_,
		_w3540_,
		_w3541_,
		_w3542_,
		_w6590_
	);
	LUT3 #(
		.INIT('h10)
	) name4690 (
		\s0_msel_arb3_state_reg[0]/NET0131 ,
		\s0_msel_arb3_state_reg[1]/NET0131 ,
		\s0_msel_arb3_state_reg[2]/NET0131 ,
		_w6591_
	);
	LUT4 #(
		.INIT('h2300)
	) name4691 (
		_w3529_,
		_w3530_,
		_w3537_,
		_w6591_,
		_w6592_
	);
	LUT3 #(
		.INIT('hd0)
	) name4692 (
		_w6584_,
		_w6590_,
		_w6592_,
		_w6593_
	);
	LUT3 #(
		.INIT('h0e)
	) name4693 (
		_w3530_,
		_w6588_,
		_w6593_,
		_w6594_
	);
	LUT2 #(
		.INIT('h1)
	) name4694 (
		\s0_msel_arb3_state_reg[1]/NET0131 ,
		\s0_msel_arb3_state_reg[2]/NET0131 ,
		_w6595_
	);
	LUT4 #(
		.INIT('h0080)
	) name4695 (
		\m0_s0_cyc_o_reg/NET0131 ,
		\rf_conf0_reg[0]/NET0131 ,
		\rf_conf0_reg[1]/NET0131 ,
		\s0_msel_arb3_state_reg[0]/NET0131 ,
		_w6596_
	);
	LUT2 #(
		.INIT('h2)
	) name4696 (
		_w6595_,
		_w6596_,
		_w6597_
	);
	LUT2 #(
		.INIT('h1)
	) name4697 (
		_w3530_,
		_w3540_,
		_w6598_
	);
	LUT4 #(
		.INIT('h4fcf)
	) name4698 (
		_w6585_,
		_w6589_,
		_w6597_,
		_w6598_,
		_w6599_
	);
	LUT3 #(
		.INIT('h20)
	) name4699 (
		_w3539_,
		_w3547_,
		_w6582_,
		_w6600_
	);
	LUT3 #(
		.INIT('h20)
	) name4700 (
		\s0_msel_arb3_state_reg[0]/NET0131 ,
		\s0_msel_arb3_state_reg[1]/NET0131 ,
		\s0_msel_arb3_state_reg[2]/NET0131 ,
		_w6601_
	);
	LUT2 #(
		.INIT('h8)
	) name4701 (
		_w3529_,
		_w6601_,
		_w6602_
	);
	LUT2 #(
		.INIT('h1)
	) name4702 (
		_w6600_,
		_w6602_,
		_w6603_
	);
	LUT2 #(
		.INIT('h8)
	) name4703 (
		_w6599_,
		_w6603_,
		_w6604_
	);
	LUT3 #(
		.INIT('h02)
	) name4704 (
		\s0_msel_arb3_state_reg[0]/NET0131 ,
		\s0_msel_arb3_state_reg[1]/NET0131 ,
		\s0_msel_arb3_state_reg[2]/NET0131 ,
		_w6605_
	);
	LUT4 #(
		.INIT('h0100)
	) name4705 (
		_w3530_,
		_w3540_,
		_w3542_,
		_w6605_,
		_w6606_
	);
	LUT2 #(
		.INIT('h4)
	) name4706 (
		_w3529_,
		_w6601_,
		_w6607_
	);
	LUT2 #(
		.INIT('h1)
	) name4707 (
		_w6606_,
		_w6607_,
		_w6608_
	);
	LUT2 #(
		.INIT('h4)
	) name4708 (
		_w3536_,
		_w3542_,
		_w6609_
	);
	LUT4 #(
		.INIT('h0051)
	) name4709 (
		_w3536_,
		_w3539_,
		_w3540_,
		_w3541_,
		_w6610_
	);
	LUT4 #(
		.INIT('h7f00)
	) name4710 (
		\m0_s0_cyc_o_reg/NET0131 ,
		\rf_conf0_reg[0]/NET0131 ,
		\rf_conf0_reg[1]/NET0131 ,
		\s0_msel_arb3_state_reg[0]/NET0131 ,
		_w6611_
	);
	LUT3 #(
		.INIT('h10)
	) name4711 (
		_w3530_,
		_w3540_,
		_w6611_,
		_w6612_
	);
	LUT4 #(
		.INIT('h0054)
	) name4712 (
		_w6606_,
		_w6609_,
		_w6610_,
		_w6612_,
		_w6613_
	);
	LUT3 #(
		.INIT('h01)
	) name4713 (
		_w3537_,
		_w6608_,
		_w6613_,
		_w6614_
	);
	LUT4 #(
		.INIT('h007f)
	) name4714 (
		\m5_s0_cyc_o_reg/NET0131 ,
		\rf_conf0_reg[10]/NET0131 ,
		\rf_conf0_reg[11]/NET0131 ,
		\s0_msel_arb3_state_reg[0]/NET0131 ,
		_w6615_
	);
	LUT4 #(
		.INIT('h0001)
	) name4715 (
		_w3530_,
		_w3540_,
		_w3542_,
		_w6615_,
		_w6616_
	);
	LUT3 #(
		.INIT('h0e)
	) name4716 (
		_w6609_,
		_w6610_,
		_w6616_,
		_w6617_
	);
	LUT4 #(
		.INIT('h0080)
	) name4717 (
		\m6_s0_cyc_o_reg/NET0131 ,
		\rf_conf0_reg[12]/NET0131 ,
		\rf_conf0_reg[13]/NET0131 ,
		\s0_msel_arb3_state_reg[0]/NET0131 ,
		_w6618_
	);
	LUT3 #(
		.INIT('h10)
	) name4718 (
		_w3529_,
		_w3536_,
		_w3537_,
		_w6619_
	);
	LUT4 #(
		.INIT('h020a)
	) name4719 (
		_w3555_,
		_w6589_,
		_w6618_,
		_w6619_,
		_w6620_
	);
	LUT2 #(
		.INIT('h4)
	) name4720 (
		_w6617_,
		_w6620_,
		_w6621_
	);
	LUT4 #(
		.INIT('hfff7)
	) name4721 (
		_w6594_,
		_w6604_,
		_w6614_,
		_w6621_,
		_w6622_
	);
	LUT2 #(
		.INIT('h4)
	) name4722 (
		_w2844_,
		_w2849_,
		_w6623_
	);
	LUT4 #(
		.INIT('h000d)
	) name4723 (
		_w2839_,
		_w2840_,
		_w2844_,
		_w2848_,
		_w6624_
	);
	LUT3 #(
		.INIT('h01)
	) name4724 (
		_w2840_,
		_w2842_,
		_w2849_,
		_w6625_
	);
	LUT4 #(
		.INIT('h00fd)
	) name4725 (
		\m5_s10_cyc_o_reg/NET0131 ,
		\rf_conf10_reg[10]/NET0131 ,
		\rf_conf10_reg[11]/NET0131 ,
		\s10_msel_arb0_state_reg[0]/NET0131 ,
		_w6626_
	);
	LUT3 #(
		.INIT('hce)
	) name4726 (
		\s10_msel_arb0_state_reg[0]/NET0131 ,
		_w2843_,
		_w2845_,
		_w6627_
	);
	LUT4 #(
		.INIT('h0eee)
	) name4727 (
		_w6623_,
		_w6624_,
		_w6625_,
		_w6627_,
		_w6628_
	);
	LUT3 #(
		.INIT('hae)
	) name4728 (
		_w2843_,
		_w2844_,
		_w2845_,
		_w6629_
	);
	LUT2 #(
		.INIT('h4)
	) name4729 (
		\s10_msel_arb0_state_reg[1]/NET0131 ,
		\s10_msel_arb0_state_reg[2]/NET0131 ,
		_w6630_
	);
	LUT4 #(
		.INIT('h0002)
	) name4730 (
		\m1_s10_cyc_o_reg/NET0131 ,
		\rf_conf10_reg[2]/NET0131 ,
		\rf_conf10_reg[3]/NET0131 ,
		\s10_msel_arb0_state_reg[1]/NET0131 ,
		_w6631_
	);
	LUT2 #(
		.INIT('h1)
	) name4731 (
		_w6630_,
		_w6631_,
		_w6632_
	);
	LUT3 #(
		.INIT('h23)
	) name4732 (
		_w2839_,
		_w2840_,
		_w2842_,
		_w6633_
	);
	LUT4 #(
		.INIT('h00dc)
	) name4733 (
		_w2839_,
		_w2840_,
		_w2842_,
		_w2848_,
		_w6634_
	);
	LUT3 #(
		.INIT('ha8)
	) name4734 (
		\s10_msel_arb0_state_reg[2]/NET0131 ,
		_w2845_,
		_w2849_,
		_w6635_
	);
	LUT4 #(
		.INIT('hdddc)
	) name4735 (
		_w6629_,
		_w6632_,
		_w6634_,
		_w6635_,
		_w6636_
	);
	LUT4 #(
		.INIT('h08aa)
	) name4736 (
		\s10_msel_arb0_state_reg[0]/NET0131 ,
		_w2872_,
		_w6628_,
		_w6636_,
		_w6637_
	);
	LUT3 #(
		.INIT('h02)
	) name4737 (
		\s10_msel_arb0_state_reg[0]/NET0131 ,
		_w2845_,
		_w2849_,
		_w6638_
	);
	LUT2 #(
		.INIT('h1)
	) name4738 (
		_w2840_,
		_w2842_,
		_w6639_
	);
	LUT3 #(
		.INIT('h80)
	) name4739 (
		_w2867_,
		_w6638_,
		_w6639_,
		_w6640_
	);
	LUT3 #(
		.INIT('h04)
	) name4740 (
		_w2845_,
		_w2848_,
		_w2849_,
		_w6641_
	);
	LUT4 #(
		.INIT('h1101)
	) name4741 (
		_w2839_,
		_w2843_,
		_w2844_,
		_w2845_,
		_w6642_
	);
	LUT4 #(
		.INIT('h0002)
	) name4742 (
		\m2_s10_cyc_o_reg/NET0131 ,
		\rf_conf10_reg[4]/NET0131 ,
		\rf_conf10_reg[5]/NET0131 ,
		\s10_msel_arb0_state_reg[0]/NET0131 ,
		_w6643_
	);
	LUT4 #(
		.INIT('h00b0)
	) name4743 (
		_w2839_,
		_w2842_,
		_w2867_,
		_w6643_,
		_w6644_
	);
	LUT3 #(
		.INIT('hb0)
	) name4744 (
		_w6641_,
		_w6642_,
		_w6644_,
		_w6645_
	);
	LUT2 #(
		.INIT('h1)
	) name4745 (
		_w6640_,
		_w6645_,
		_w6646_
	);
	LUT4 #(
		.INIT('h00f2)
	) name4746 (
		_w2839_,
		_w2840_,
		_w2848_,
		_w2849_,
		_w6647_
	);
	LUT3 #(
		.INIT('ha8)
	) name4747 (
		\s10_msel_arb0_state_reg[2]/NET0131 ,
		_w2842_,
		_w2845_,
		_w6648_
	);
	LUT3 #(
		.INIT('h54)
	) name4748 (
		\s10_msel_arb0_state_reg[2]/NET0131 ,
		_w2840_,
		_w2849_,
		_w6649_
	);
	LUT4 #(
		.INIT('h4454)
	) name4749 (
		_w2842_,
		_w2843_,
		_w2844_,
		_w2845_,
		_w6650_
	);
	LUT4 #(
		.INIT('hd0dd)
	) name4750 (
		_w6647_,
		_w6648_,
		_w6649_,
		_w6650_,
		_w6651_
	);
	LUT2 #(
		.INIT('h1)
	) name4751 (
		\s10_msel_arb0_state_reg[0]/NET0131 ,
		\s10_msel_arb0_state_reg[1]/NET0131 ,
		_w6652_
	);
	LUT3 #(
		.INIT('h02)
	) name4752 (
		\s10_msel_arb0_state_reg[0]/NET0131 ,
		\s10_msel_arb0_state_reg[1]/NET0131 ,
		\s10_msel_arb0_state_reg[2]/NET0131 ,
		_w6653_
	);
	LUT2 #(
		.INIT('h4)
	) name4753 (
		_w2848_,
		_w6653_,
		_w6654_
	);
	LUT4 #(
		.INIT('h8a00)
	) name4754 (
		_w6633_,
		_w6638_,
		_w6642_,
		_w6654_,
		_w6655_
	);
	LUT4 #(
		.INIT('h0001)
	) name4755 (
		_w2840_,
		_w2842_,
		_w2849_,
		_w6626_,
		_w6656_
	);
	LUT3 #(
		.INIT('h40)
	) name4756 (
		\s10_msel_arb0_state_reg[0]/NET0131 ,
		\s10_msel_arb0_state_reg[1]/NET0131 ,
		\s10_msel_arb0_state_reg[2]/NET0131 ,
		_w6657_
	);
	LUT2 #(
		.INIT('h4)
	) name4757 (
		_w2845_,
		_w6657_,
		_w6658_
	);
	LUT4 #(
		.INIT('hf100)
	) name4758 (
		_w6623_,
		_w6624_,
		_w6656_,
		_w6658_,
		_w6659_
	);
	LUT4 #(
		.INIT('h000b)
	) name4759 (
		_w6651_,
		_w6652_,
		_w6655_,
		_w6659_,
		_w6660_
	);
	LUT3 #(
		.INIT('hbf)
	) name4760 (
		_w6637_,
		_w6646_,
		_w6660_,
		_w6661_
	);
	LUT4 #(
		.INIT('h0100)
	) name4761 (
		_w4026_,
		_w4034_,
		_w4035_,
		_w4052_,
		_w6662_
	);
	LUT4 #(
		.INIT('h2223)
	) name4762 (
		\s10_msel_arb2_state_reg[1]/NET0131 ,
		\s10_msel_arb2_state_reg[2]/NET0131 ,
		_w4026_,
		_w4034_,
		_w6663_
	);
	LUT2 #(
		.INIT('h1)
	) name4763 (
		_w4031_,
		_w4032_,
		_w6664_
	);
	LUT4 #(
		.INIT('h0001)
	) name4764 (
		_w4030_,
		_w4031_,
		_w4032_,
		_w4038_,
		_w6665_
	);
	LUT4 #(
		.INIT('hbbab)
	) name4765 (
		_w4027_,
		_w6662_,
		_w6663_,
		_w6665_,
		_w6666_
	);
	LUT4 #(
		.INIT('hfe00)
	) name4766 (
		_w4030_,
		_w4031_,
		_w4032_,
		_w4052_,
		_w6667_
	);
	LUT3 #(
		.INIT('ha2)
	) name4767 (
		\s10_msel_arb2_state_reg[0]/NET0131 ,
		_w6666_,
		_w6667_,
		_w6668_
	);
	LUT2 #(
		.INIT('h2)
	) name4768 (
		\s10_msel_arb2_state_reg[0]/NET0131 ,
		\s10_msel_arb2_state_reg[1]/NET0131 ,
		_w6669_
	);
	LUT2 #(
		.INIT('h1)
	) name4769 (
		_w4026_,
		_w4027_,
		_w6670_
	);
	LUT4 #(
		.INIT('h0001)
	) name4770 (
		_w4026_,
		_w4027_,
		_w4034_,
		_w4035_,
		_w6671_
	);
	LUT4 #(
		.INIT('hdf00)
	) name4771 (
		\m7_s10_cyc_o_reg/NET0131 ,
		\rf_conf10_reg[14]/NET0131 ,
		\rf_conf10_reg[15]/NET0131 ,
		\s10_msel_arb2_state_reg[0]/NET0131 ,
		_w6672_
	);
	LUT3 #(
		.INIT('h45)
	) name4772 (
		_w6669_,
		_w6671_,
		_w6672_,
		_w6673_
	);
	LUT3 #(
		.INIT('h54)
	) name4773 (
		\s10_msel_arb2_state_reg[1]/NET0131 ,
		_w4030_,
		_w4038_,
		_w6674_
	);
	LUT3 #(
		.INIT('h02)
	) name4774 (
		_w6664_,
		_w6671_,
		_w6674_,
		_w6675_
	);
	LUT3 #(
		.INIT('h54)
	) name4775 (
		\s10_msel_arb2_state_reg[1]/NET0131 ,
		_w4034_,
		_w4035_,
		_w6676_
	);
	LUT4 #(
		.INIT('h0010)
	) name4776 (
		\s10_msel_arb2_state_reg[0]/NET0131 ,
		_w6665_,
		_w6670_,
		_w6676_,
		_w6677_
	);
	LUT4 #(
		.INIT('h5d08)
	) name4777 (
		\s10_msel_arb2_state_reg[2]/NET0131 ,
		_w6673_,
		_w6675_,
		_w6677_,
		_w6678_
	);
	LUT2 #(
		.INIT('he)
	) name4778 (
		_w6668_,
		_w6678_,
		_w6679_
	);
	LUT4 #(
		.INIT('h0100)
	) name4779 (
		_w4364_,
		_w4372_,
		_w4373_,
		_w4390_,
		_w6680_
	);
	LUT4 #(
		.INIT('h2223)
	) name4780 (
		\s12_msel_arb2_state_reg[1]/NET0131 ,
		\s12_msel_arb2_state_reg[2]/NET0131 ,
		_w4364_,
		_w4372_,
		_w6681_
	);
	LUT2 #(
		.INIT('h1)
	) name4781 (
		_w4369_,
		_w4370_,
		_w6682_
	);
	LUT4 #(
		.INIT('h0001)
	) name4782 (
		_w4368_,
		_w4369_,
		_w4370_,
		_w4376_,
		_w6683_
	);
	LUT4 #(
		.INIT('hbbab)
	) name4783 (
		_w4365_,
		_w6680_,
		_w6681_,
		_w6683_,
		_w6684_
	);
	LUT4 #(
		.INIT('hfe00)
	) name4784 (
		_w4368_,
		_w4369_,
		_w4370_,
		_w4390_,
		_w6685_
	);
	LUT3 #(
		.INIT('ha2)
	) name4785 (
		\s12_msel_arb2_state_reg[0]/NET0131 ,
		_w6684_,
		_w6685_,
		_w6686_
	);
	LUT2 #(
		.INIT('h2)
	) name4786 (
		\s12_msel_arb2_state_reg[0]/NET0131 ,
		\s12_msel_arb2_state_reg[1]/NET0131 ,
		_w6687_
	);
	LUT2 #(
		.INIT('h1)
	) name4787 (
		_w4364_,
		_w4365_,
		_w6688_
	);
	LUT4 #(
		.INIT('h0001)
	) name4788 (
		_w4364_,
		_w4365_,
		_w4372_,
		_w4373_,
		_w6689_
	);
	LUT4 #(
		.INIT('hdf00)
	) name4789 (
		\m7_s12_cyc_o_reg/NET0131 ,
		\rf_conf12_reg[14]/NET0131 ,
		\rf_conf12_reg[15]/NET0131 ,
		\s12_msel_arb2_state_reg[0]/NET0131 ,
		_w6690_
	);
	LUT3 #(
		.INIT('h45)
	) name4790 (
		_w6687_,
		_w6689_,
		_w6690_,
		_w6691_
	);
	LUT3 #(
		.INIT('h54)
	) name4791 (
		\s12_msel_arb2_state_reg[1]/NET0131 ,
		_w4368_,
		_w4376_,
		_w6692_
	);
	LUT3 #(
		.INIT('h02)
	) name4792 (
		_w6682_,
		_w6689_,
		_w6692_,
		_w6693_
	);
	LUT3 #(
		.INIT('h54)
	) name4793 (
		\s12_msel_arb2_state_reg[1]/NET0131 ,
		_w4372_,
		_w4373_,
		_w6694_
	);
	LUT4 #(
		.INIT('h0010)
	) name4794 (
		\s12_msel_arb2_state_reg[0]/NET0131 ,
		_w6683_,
		_w6688_,
		_w6694_,
		_w6695_
	);
	LUT4 #(
		.INIT('h5d08)
	) name4795 (
		\s12_msel_arb2_state_reg[2]/NET0131 ,
		_w6691_,
		_w6693_,
		_w6695_,
		_w6696_
	);
	LUT2 #(
		.INIT('he)
	) name4796 (
		_w6686_,
		_w6696_,
		_w6697_
	);
	LUT2 #(
		.INIT('h1)
	) name4797 (
		_w4553_,
		_w4557_,
		_w6698_
	);
	LUT2 #(
		.INIT('h1)
	) name4798 (
		_w4555_,
		_w4556_,
		_w6699_
	);
	LUT4 #(
		.INIT('h0001)
	) name4799 (
		_w4553_,
		_w4555_,
		_w4556_,
		_w4557_,
		_w6700_
	);
	LUT4 #(
		.INIT('h0020)
	) name4800 (
		\m4_s13_cyc_o_reg/NET0131 ,
		\rf_conf13_reg[8]/NET0131 ,
		\rf_conf13_reg[9]/NET0131 ,
		\s13_msel_arb2_state_reg[1]/NET0131 ,
		_w6701_
	);
	LUT3 #(
		.INIT('h54)
	) name4801 (
		\s13_msel_arb2_state_reg[0]/NET0131 ,
		_w4560_,
		_w6701_,
		_w6702_
	);
	LUT3 #(
		.INIT('h54)
	) name4802 (
		\s13_msel_arb2_state_reg[1]/NET0131 ,
		_w4559_,
		_w4560_,
		_w6703_
	);
	LUT4 #(
		.INIT('h0001)
	) name4803 (
		_w4552_,
		_w6700_,
		_w6702_,
		_w6703_,
		_w6704_
	);
	LUT4 #(
		.INIT('h00df)
	) name4804 (
		\m3_s13_cyc_o_reg/NET0131 ,
		\rf_conf13_reg[6]/NET0131 ,
		\rf_conf13_reg[7]/NET0131 ,
		\s13_msel_arb2_state_reg[2]/NET0131 ,
		_w6705_
	);
	LUT4 #(
		.INIT('hab00)
	) name4805 (
		\s13_msel_arb2_state_reg[1]/NET0131 ,
		_w4556_,
		_w4557_,
		_w6705_,
		_w6706_
	);
	LUT2 #(
		.INIT('h1)
	) name4806 (
		_w4552_,
		_w4560_,
		_w6707_
	);
	LUT4 #(
		.INIT('h0001)
	) name4807 (
		_w4551_,
		_w4552_,
		_w4559_,
		_w4560_,
		_w6708_
	);
	LUT2 #(
		.INIT('h1)
	) name4808 (
		\s13_msel_arb2_state_reg[0]/NET0131 ,
		\s13_msel_arb2_state_reg[1]/NET0131 ,
		_w6709_
	);
	LUT3 #(
		.INIT('h13)
	) name4809 (
		_w4553_,
		_w4590_,
		_w6709_,
		_w6710_
	);
	LUT3 #(
		.INIT('h20)
	) name4810 (
		_w6706_,
		_w6708_,
		_w6710_,
		_w6711_
	);
	LUT3 #(
		.INIT('hf2)
	) name4811 (
		\s13_msel_arb2_state_reg[2]/NET0131 ,
		_w6704_,
		_w6711_,
		_w6712_
	);
	LUT2 #(
		.INIT('h1)
	) name4812 (
		_w5186_,
		_w5190_,
		_w6713_
	);
	LUT2 #(
		.INIT('h1)
	) name4813 (
		_w5188_,
		_w5189_,
		_w6714_
	);
	LUT4 #(
		.INIT('h0001)
	) name4814 (
		_w5186_,
		_w5188_,
		_w5189_,
		_w5190_,
		_w6715_
	);
	LUT4 #(
		.INIT('h0020)
	) name4815 (
		\m4_s2_cyc_o_reg/NET0131 ,
		\rf_conf2_reg[8]/NET0131 ,
		\rf_conf2_reg[9]/NET0131 ,
		\s2_msel_arb2_state_reg[1]/NET0131 ,
		_w6716_
	);
	LUT3 #(
		.INIT('h54)
	) name4816 (
		\s2_msel_arb2_state_reg[0]/NET0131 ,
		_w5193_,
		_w6716_,
		_w6717_
	);
	LUT3 #(
		.INIT('h54)
	) name4817 (
		\s2_msel_arb2_state_reg[1]/NET0131 ,
		_w5192_,
		_w5193_,
		_w6718_
	);
	LUT4 #(
		.INIT('h0001)
	) name4818 (
		_w5185_,
		_w6715_,
		_w6717_,
		_w6718_,
		_w6719_
	);
	LUT4 #(
		.INIT('h00df)
	) name4819 (
		\m3_s2_cyc_o_reg/NET0131 ,
		\rf_conf2_reg[6]/NET0131 ,
		\rf_conf2_reg[7]/NET0131 ,
		\s2_msel_arb2_state_reg[2]/NET0131 ,
		_w6720_
	);
	LUT4 #(
		.INIT('hab00)
	) name4820 (
		\s2_msel_arb2_state_reg[1]/NET0131 ,
		_w5189_,
		_w5190_,
		_w6720_,
		_w6721_
	);
	LUT2 #(
		.INIT('h1)
	) name4821 (
		_w5185_,
		_w5193_,
		_w6722_
	);
	LUT4 #(
		.INIT('h0001)
	) name4822 (
		_w5184_,
		_w5185_,
		_w5192_,
		_w5193_,
		_w6723_
	);
	LUT2 #(
		.INIT('h1)
	) name4823 (
		\s2_msel_arb2_state_reg[0]/NET0131 ,
		\s2_msel_arb2_state_reg[1]/NET0131 ,
		_w6724_
	);
	LUT3 #(
		.INIT('h13)
	) name4824 (
		_w5186_,
		_w5223_,
		_w6724_,
		_w6725_
	);
	LUT3 #(
		.INIT('h20)
	) name4825 (
		_w6721_,
		_w6723_,
		_w6725_,
		_w6726_
	);
	LUT3 #(
		.INIT('hf2)
	) name4826 (
		\s2_msel_arb2_state_reg[2]/NET0131 ,
		_w6719_,
		_w6726_,
		_w6727_
	);
	LUT2 #(
		.INIT('h1)
	) name4827 (
		_w5537_,
		_w5541_,
		_w6728_
	);
	LUT2 #(
		.INIT('h1)
	) name4828 (
		_w5539_,
		_w5540_,
		_w6729_
	);
	LUT4 #(
		.INIT('h0001)
	) name4829 (
		_w5537_,
		_w5539_,
		_w5540_,
		_w5541_,
		_w6730_
	);
	LUT4 #(
		.INIT('h0020)
	) name4830 (
		\m4_s4_cyc_o_reg/NET0131 ,
		\rf_conf4_reg[8]/NET0131 ,
		\rf_conf4_reg[9]/NET0131 ,
		\s4_msel_arb2_state_reg[1]/NET0131 ,
		_w6731_
	);
	LUT3 #(
		.INIT('h54)
	) name4831 (
		\s4_msel_arb2_state_reg[0]/NET0131 ,
		_w5544_,
		_w6731_,
		_w6732_
	);
	LUT3 #(
		.INIT('h54)
	) name4832 (
		\s4_msel_arb2_state_reg[1]/NET0131 ,
		_w5543_,
		_w5544_,
		_w6733_
	);
	LUT4 #(
		.INIT('h0001)
	) name4833 (
		_w5536_,
		_w6730_,
		_w6732_,
		_w6733_,
		_w6734_
	);
	LUT4 #(
		.INIT('h00df)
	) name4834 (
		\m3_s4_cyc_o_reg/NET0131 ,
		\rf_conf4_reg[6]/NET0131 ,
		\rf_conf4_reg[7]/NET0131 ,
		\s4_msel_arb2_state_reg[2]/NET0131 ,
		_w6735_
	);
	LUT4 #(
		.INIT('hab00)
	) name4835 (
		\s4_msel_arb2_state_reg[1]/NET0131 ,
		_w5540_,
		_w5541_,
		_w6735_,
		_w6736_
	);
	LUT2 #(
		.INIT('h1)
	) name4836 (
		_w5536_,
		_w5544_,
		_w6737_
	);
	LUT4 #(
		.INIT('h0001)
	) name4837 (
		_w5535_,
		_w5536_,
		_w5543_,
		_w5544_,
		_w6738_
	);
	LUT2 #(
		.INIT('h1)
	) name4838 (
		\s4_msel_arb2_state_reg[0]/NET0131 ,
		\s4_msel_arb2_state_reg[1]/NET0131 ,
		_w6739_
	);
	LUT3 #(
		.INIT('h13)
	) name4839 (
		_w5537_,
		_w5574_,
		_w6739_,
		_w6740_
	);
	LUT3 #(
		.INIT('h20)
	) name4840 (
		_w6736_,
		_w6738_,
		_w6740_,
		_w6741_
	);
	LUT3 #(
		.INIT('hf2)
	) name4841 (
		\s4_msel_arb2_state_reg[2]/NET0131 ,
		_w6734_,
		_w6741_,
		_w6742_
	);
	LUT4 #(
		.INIT('h0100)
	) name4842 (
		_w6038_,
		_w6046_,
		_w6047_,
		_w6064_,
		_w6743_
	);
	LUT4 #(
		.INIT('h2223)
	) name4843 (
		\s7_msel_arb2_state_reg[1]/NET0131 ,
		\s7_msel_arb2_state_reg[2]/NET0131 ,
		_w6038_,
		_w6046_,
		_w6744_
	);
	LUT2 #(
		.INIT('h1)
	) name4844 (
		_w6043_,
		_w6044_,
		_w6745_
	);
	LUT4 #(
		.INIT('h0001)
	) name4845 (
		_w6042_,
		_w6043_,
		_w6044_,
		_w6050_,
		_w6746_
	);
	LUT4 #(
		.INIT('hbbab)
	) name4846 (
		_w6039_,
		_w6743_,
		_w6744_,
		_w6746_,
		_w6747_
	);
	LUT4 #(
		.INIT('hfe00)
	) name4847 (
		_w6042_,
		_w6043_,
		_w6044_,
		_w6064_,
		_w6748_
	);
	LUT3 #(
		.INIT('ha2)
	) name4848 (
		\s7_msel_arb2_state_reg[0]/NET0131 ,
		_w6747_,
		_w6748_,
		_w6749_
	);
	LUT2 #(
		.INIT('h2)
	) name4849 (
		\s7_msel_arb2_state_reg[0]/NET0131 ,
		\s7_msel_arb2_state_reg[1]/NET0131 ,
		_w6750_
	);
	LUT2 #(
		.INIT('h1)
	) name4850 (
		_w6038_,
		_w6039_,
		_w6751_
	);
	LUT4 #(
		.INIT('h0001)
	) name4851 (
		_w6038_,
		_w6039_,
		_w6046_,
		_w6047_,
		_w6752_
	);
	LUT4 #(
		.INIT('hdf00)
	) name4852 (
		\m7_s7_cyc_o_reg/NET0131 ,
		\rf_conf7_reg[14]/NET0131 ,
		\rf_conf7_reg[15]/NET0131 ,
		\s7_msel_arb2_state_reg[0]/NET0131 ,
		_w6753_
	);
	LUT3 #(
		.INIT('h45)
	) name4853 (
		_w6750_,
		_w6752_,
		_w6753_,
		_w6754_
	);
	LUT3 #(
		.INIT('h54)
	) name4854 (
		\s7_msel_arb2_state_reg[1]/NET0131 ,
		_w6042_,
		_w6050_,
		_w6755_
	);
	LUT3 #(
		.INIT('h02)
	) name4855 (
		_w6745_,
		_w6752_,
		_w6755_,
		_w6756_
	);
	LUT3 #(
		.INIT('h54)
	) name4856 (
		\s7_msel_arb2_state_reg[1]/NET0131 ,
		_w6046_,
		_w6047_,
		_w6757_
	);
	LUT4 #(
		.INIT('h0010)
	) name4857 (
		\s7_msel_arb2_state_reg[0]/NET0131 ,
		_w6746_,
		_w6751_,
		_w6757_,
		_w6758_
	);
	LUT4 #(
		.INIT('h5d08)
	) name4858 (
		\s7_msel_arb2_state_reg[2]/NET0131 ,
		_w6754_,
		_w6756_,
		_w6758_,
		_w6759_
	);
	LUT2 #(
		.INIT('he)
	) name4859 (
		_w6749_,
		_w6759_,
		_w6760_
	);
	LUT4 #(
		.INIT('h0100)
	) name4860 (
		_w6366_,
		_w6374_,
		_w6375_,
		_w6392_,
		_w6761_
	);
	LUT4 #(
		.INIT('h2223)
	) name4861 (
		\s9_msel_arb2_state_reg[1]/NET0131 ,
		\s9_msel_arb2_state_reg[2]/NET0131 ,
		_w6366_,
		_w6374_,
		_w6762_
	);
	LUT2 #(
		.INIT('h1)
	) name4862 (
		_w6371_,
		_w6372_,
		_w6763_
	);
	LUT4 #(
		.INIT('h0001)
	) name4863 (
		_w6370_,
		_w6371_,
		_w6372_,
		_w6378_,
		_w6764_
	);
	LUT4 #(
		.INIT('hbbab)
	) name4864 (
		_w6367_,
		_w6761_,
		_w6762_,
		_w6764_,
		_w6765_
	);
	LUT4 #(
		.INIT('hfe00)
	) name4865 (
		_w6370_,
		_w6371_,
		_w6372_,
		_w6392_,
		_w6766_
	);
	LUT3 #(
		.INIT('ha2)
	) name4866 (
		\s9_msel_arb2_state_reg[0]/NET0131 ,
		_w6765_,
		_w6766_,
		_w6767_
	);
	LUT2 #(
		.INIT('h2)
	) name4867 (
		\s9_msel_arb2_state_reg[0]/NET0131 ,
		\s9_msel_arb2_state_reg[1]/NET0131 ,
		_w6768_
	);
	LUT2 #(
		.INIT('h1)
	) name4868 (
		_w6366_,
		_w6367_,
		_w6769_
	);
	LUT4 #(
		.INIT('h0001)
	) name4869 (
		_w6366_,
		_w6367_,
		_w6374_,
		_w6375_,
		_w6770_
	);
	LUT4 #(
		.INIT('hdf00)
	) name4870 (
		\m7_s9_cyc_o_reg/NET0131 ,
		\rf_conf9_reg[14]/NET0131 ,
		\rf_conf9_reg[15]/NET0131 ,
		\s9_msel_arb2_state_reg[0]/NET0131 ,
		_w6771_
	);
	LUT3 #(
		.INIT('h45)
	) name4871 (
		_w6768_,
		_w6770_,
		_w6771_,
		_w6772_
	);
	LUT3 #(
		.INIT('h54)
	) name4872 (
		\s9_msel_arb2_state_reg[1]/NET0131 ,
		_w6370_,
		_w6378_,
		_w6773_
	);
	LUT3 #(
		.INIT('h02)
	) name4873 (
		_w6763_,
		_w6770_,
		_w6773_,
		_w6774_
	);
	LUT3 #(
		.INIT('h54)
	) name4874 (
		\s9_msel_arb2_state_reg[1]/NET0131 ,
		_w6374_,
		_w6375_,
		_w6775_
	);
	LUT4 #(
		.INIT('h0010)
	) name4875 (
		\s9_msel_arb2_state_reg[0]/NET0131 ,
		_w6764_,
		_w6769_,
		_w6775_,
		_w6776_
	);
	LUT4 #(
		.INIT('h5d08)
	) name4876 (
		\s9_msel_arb2_state_reg[2]/NET0131 ,
		_w6772_,
		_w6774_,
		_w6776_,
		_w6777_
	);
	LUT2 #(
		.INIT('he)
	) name4877 (
		_w6767_,
		_w6777_,
		_w6778_
	);
	LUT2 #(
		.INIT('h1)
	) name4878 (
		_w6423_,
		_w6427_,
		_w6779_
	);
	LUT2 #(
		.INIT('h1)
	) name4879 (
		_w6425_,
		_w6426_,
		_w6780_
	);
	LUT4 #(
		.INIT('h0001)
	) name4880 (
		_w6423_,
		_w6425_,
		_w6426_,
		_w6427_,
		_w6781_
	);
	LUT4 #(
		.INIT('h0080)
	) name4881 (
		\m4_s9_cyc_o_reg/NET0131 ,
		\rf_conf9_reg[8]/NET0131 ,
		\rf_conf9_reg[9]/NET0131 ,
		\s9_msel_arb3_state_reg[1]/NET0131 ,
		_w6782_
	);
	LUT3 #(
		.INIT('h54)
	) name4882 (
		\s9_msel_arb3_state_reg[0]/NET0131 ,
		_w6430_,
		_w6782_,
		_w6783_
	);
	LUT3 #(
		.INIT('h54)
	) name4883 (
		\s9_msel_arb3_state_reg[1]/NET0131 ,
		_w6429_,
		_w6430_,
		_w6784_
	);
	LUT4 #(
		.INIT('h0001)
	) name4884 (
		_w6422_,
		_w6781_,
		_w6783_,
		_w6784_,
		_w6785_
	);
	LUT4 #(
		.INIT('h007f)
	) name4885 (
		\m3_s9_cyc_o_reg/NET0131 ,
		\rf_conf9_reg[6]/NET0131 ,
		\rf_conf9_reg[7]/NET0131 ,
		\s9_msel_arb3_state_reg[2]/NET0131 ,
		_w6786_
	);
	LUT4 #(
		.INIT('hab00)
	) name4886 (
		\s9_msel_arb3_state_reg[1]/NET0131 ,
		_w6426_,
		_w6427_,
		_w6786_,
		_w6787_
	);
	LUT2 #(
		.INIT('h1)
	) name4887 (
		_w6422_,
		_w6430_,
		_w6788_
	);
	LUT4 #(
		.INIT('h0001)
	) name4888 (
		_w6421_,
		_w6422_,
		_w6429_,
		_w6430_,
		_w6789_
	);
	LUT2 #(
		.INIT('h1)
	) name4889 (
		\s9_msel_arb3_state_reg[0]/NET0131 ,
		\s9_msel_arb3_state_reg[1]/NET0131 ,
		_w6790_
	);
	LUT3 #(
		.INIT('h13)
	) name4890 (
		_w6423_,
		_w6460_,
		_w6790_,
		_w6791_
	);
	LUT3 #(
		.INIT('h20)
	) name4891 (
		_w6787_,
		_w6789_,
		_w6791_,
		_w6792_
	);
	LUT3 #(
		.INIT('hf2)
	) name4892 (
		\s9_msel_arb3_state_reg[2]/NET0131 ,
		_w6785_,
		_w6792_,
		_w6793_
	);
	LUT3 #(
		.INIT('h54)
	) name4893 (
		\s10_msel_arb0_state_reg[1]/NET0131 ,
		_w2843_,
		_w2863_,
		_w6794_
	);
	LUT4 #(
		.INIT('h0001)
	) name4894 (
		_w2839_,
		_w2840_,
		_w2848_,
		_w2849_,
		_w6795_
	);
	LUT2 #(
		.INIT('h8)
	) name4895 (
		\s10_msel_arb0_state_reg[0]/NET0131 ,
		\s10_msel_arb0_state_reg[1]/NET0131 ,
		_w6796_
	);
	LUT3 #(
		.INIT('h51)
	) name4896 (
		_w2844_,
		_w2845_,
		_w6796_,
		_w6797_
	);
	LUT4 #(
		.INIT('ha8aa)
	) name4897 (
		\s10_msel_arb0_state_reg[2]/NET0131 ,
		_w6794_,
		_w6795_,
		_w6797_,
		_w6798_
	);
	LUT4 #(
		.INIT('h0015)
	) name4898 (
		_w2840_,
		_w2849_,
		_w6652_,
		_w6631_,
		_w6799_
	);
	LUT4 #(
		.INIT('h0001)
	) name4899 (
		_w2842_,
		_w2843_,
		_w2844_,
		_w2845_,
		_w6800_
	);
	LUT4 #(
		.INIT('h00fd)
	) name4900 (
		\m3_s10_cyc_o_reg/NET0131 ,
		\rf_conf10_reg[6]/NET0131 ,
		\rf_conf10_reg[7]/NET0131 ,
		\s10_msel_arb0_state_reg[2]/NET0131 ,
		_w6801_
	);
	LUT4 #(
		.INIT('h0e00)
	) name4901 (
		_w6796_,
		_w6799_,
		_w6800_,
		_w6801_,
		_w6802_
	);
	LUT2 #(
		.INIT('he)
	) name4902 (
		_w6798_,
		_w6802_,
		_w6803_
	);
	LUT3 #(
		.INIT('h04)
	) name4903 (
		\s11_msel_arb0_state_reg[0]/NET0131 ,
		\s11_msel_arb0_state_reg[1]/NET0131 ,
		\s11_msel_arb0_state_reg[2]/NET0131 ,
		_w6804_
	);
	LUT4 #(
		.INIT('h0001)
	) name4904 (
		_w2265_,
		_w2266_,
		_w2268_,
		_w2269_,
		_w6805_
	);
	LUT2 #(
		.INIT('h4)
	) name4905 (
		_w2273_,
		_w4143_,
		_w6806_
	);
	LUT3 #(
		.INIT('h45)
	) name4906 (
		_w6804_,
		_w6805_,
		_w6806_,
		_w6807_
	);
	LUT4 #(
		.INIT('h0002)
	) name4907 (
		\m4_s11_cyc_o_reg/NET0131 ,
		\rf_conf11_reg[8]/NET0131 ,
		\rf_conf11_reg[9]/NET0131 ,
		\s11_msel_arb0_state_reg[2]/NET0131 ,
		_w6808_
	);
	LUT4 #(
		.INIT('h0001)
	) name4908 (
		_w2265_,
		_w2268_,
		_w2269_,
		_w6808_,
		_w6809_
	);
	LUT3 #(
		.INIT('h01)
	) name4909 (
		_w2270_,
		_w2273_,
		_w2278_,
		_w6810_
	);
	LUT3 #(
		.INIT('h10)
	) name4910 (
		\s11_msel_arb0_state_reg[1]/NET0131 ,
		_w6809_,
		_w6810_,
		_w6811_
	);
	LUT3 #(
		.INIT('h01)
	) name4911 (
		_w2265_,
		_w2268_,
		_w2269_,
		_w6812_
	);
	LUT4 #(
		.INIT('h0001)
	) name4912 (
		_w2270_,
		_w2271_,
		_w2273_,
		_w2278_,
		_w6813_
	);
	LUT3 #(
		.INIT('ha2)
	) name4913 (
		_w2295_,
		_w6812_,
		_w6813_,
		_w6814_
	);
	LUT3 #(
		.INIT('h10)
	) name4914 (
		_w2273_,
		_w2278_,
		_w4143_,
		_w6815_
	);
	LUT3 #(
		.INIT('h45)
	) name4915 (
		\s11_msel_arb0_state_reg[0]/NET0131 ,
		_w6805_,
		_w6815_,
		_w6816_
	);
	LUT4 #(
		.INIT('h00fd)
	) name4916 (
		_w6807_,
		_w6811_,
		_w6814_,
		_w6816_,
		_w6817_
	);
	LUT4 #(
		.INIT('h0200)
	) name4917 (
		\m6_s11_cyc_o_reg/NET0131 ,
		\rf_conf11_reg[12]/NET0131 ,
		\rf_conf11_reg[13]/NET0131 ,
		\s11_msel_arb0_state_reg[1]/NET0131 ,
		_w6818_
	);
	LUT3 #(
		.INIT('ha8)
	) name4918 (
		\s11_msel_arb0_state_reg[2]/NET0131 ,
		_w6813_,
		_w6818_,
		_w6819_
	);
	LUT4 #(
		.INIT('h0504)
	) name4919 (
		\s11_msel_arb0_state_reg[1]/NET0131 ,
		\s11_msel_arb0_state_reg[2]/NET0131 ,
		_w6805_,
		_w6813_,
		_w6820_
	);
	LUT3 #(
		.INIT('hc8)
	) name4920 (
		_w2268_,
		_w4130_,
		_w6813_,
		_w6821_
	);
	LUT4 #(
		.INIT('h00ab)
	) name4921 (
		\s11_msel_arb0_state_reg[0]/NET0131 ,
		_w6819_,
		_w6820_,
		_w6821_,
		_w6822_
	);
	LUT2 #(
		.INIT('hb)
	) name4922 (
		_w6817_,
		_w6822_,
		_w6823_
	);
	LUT3 #(
		.INIT('h04)
	) name4923 (
		\s12_msel_arb0_state_reg[0]/NET0131 ,
		\s12_msel_arb0_state_reg[1]/NET0131 ,
		\s12_msel_arb0_state_reg[2]/NET0131 ,
		_w6824_
	);
	LUT4 #(
		.INIT('h0001)
	) name4924 (
		_w2302_,
		_w2303_,
		_w2305_,
		_w2306_,
		_w6825_
	);
	LUT2 #(
		.INIT('h4)
	) name4925 (
		_w2310_,
		_w4308_,
		_w6826_
	);
	LUT3 #(
		.INIT('h45)
	) name4926 (
		_w6824_,
		_w6825_,
		_w6826_,
		_w6827_
	);
	LUT4 #(
		.INIT('h0002)
	) name4927 (
		\m4_s12_cyc_o_reg/NET0131 ,
		\rf_conf12_reg[8]/NET0131 ,
		\rf_conf12_reg[9]/NET0131 ,
		\s12_msel_arb0_state_reg[2]/NET0131 ,
		_w6828_
	);
	LUT4 #(
		.INIT('h0001)
	) name4928 (
		_w2302_,
		_w2305_,
		_w2306_,
		_w6828_,
		_w6829_
	);
	LUT3 #(
		.INIT('h01)
	) name4929 (
		_w2307_,
		_w2310_,
		_w2315_,
		_w6830_
	);
	LUT3 #(
		.INIT('h10)
	) name4930 (
		\s12_msel_arb0_state_reg[1]/NET0131 ,
		_w6829_,
		_w6830_,
		_w6831_
	);
	LUT3 #(
		.INIT('h01)
	) name4931 (
		_w2302_,
		_w2305_,
		_w2306_,
		_w6832_
	);
	LUT4 #(
		.INIT('h0001)
	) name4932 (
		_w2307_,
		_w2308_,
		_w2310_,
		_w2315_,
		_w6833_
	);
	LUT3 #(
		.INIT('ha2)
	) name4933 (
		_w2332_,
		_w6832_,
		_w6833_,
		_w6834_
	);
	LUT3 #(
		.INIT('h10)
	) name4934 (
		_w2310_,
		_w2315_,
		_w4308_,
		_w6835_
	);
	LUT3 #(
		.INIT('h45)
	) name4935 (
		\s12_msel_arb0_state_reg[0]/NET0131 ,
		_w6825_,
		_w6835_,
		_w6836_
	);
	LUT4 #(
		.INIT('h00fd)
	) name4936 (
		_w6827_,
		_w6831_,
		_w6834_,
		_w6836_,
		_w6837_
	);
	LUT4 #(
		.INIT('h0200)
	) name4937 (
		\m6_s12_cyc_o_reg/NET0131 ,
		\rf_conf12_reg[12]/NET0131 ,
		\rf_conf12_reg[13]/NET0131 ,
		\s12_msel_arb0_state_reg[1]/NET0131 ,
		_w6838_
	);
	LUT3 #(
		.INIT('ha8)
	) name4938 (
		\s12_msel_arb0_state_reg[2]/NET0131 ,
		_w6833_,
		_w6838_,
		_w6839_
	);
	LUT4 #(
		.INIT('h0504)
	) name4939 (
		\s12_msel_arb0_state_reg[1]/NET0131 ,
		\s12_msel_arb0_state_reg[2]/NET0131 ,
		_w6825_,
		_w6833_,
		_w6840_
	);
	LUT3 #(
		.INIT('hc8)
	) name4940 (
		_w2305_,
		_w4295_,
		_w6833_,
		_w6841_
	);
	LUT4 #(
		.INIT('h00ab)
	) name4941 (
		\s12_msel_arb0_state_reg[0]/NET0131 ,
		_w6839_,
		_w6840_,
		_w6841_,
		_w6842_
	);
	LUT2 #(
		.INIT('hb)
	) name4942 (
		_w6837_,
		_w6842_,
		_w6843_
	);
	LUT3 #(
		.INIT('h04)
	) name4943 (
		\s13_msel_arb0_state_reg[0]/NET0131 ,
		\s13_msel_arb0_state_reg[1]/NET0131 ,
		\s13_msel_arb0_state_reg[2]/NET0131 ,
		_w6844_
	);
	LUT4 #(
		.INIT('h0001)
	) name4944 (
		_w2339_,
		_w2340_,
		_w2342_,
		_w2343_,
		_w6845_
	);
	LUT2 #(
		.INIT('h4)
	) name4945 (
		_w2347_,
		_w4481_,
		_w6846_
	);
	LUT3 #(
		.INIT('h45)
	) name4946 (
		_w6844_,
		_w6845_,
		_w6846_,
		_w6847_
	);
	LUT4 #(
		.INIT('h0002)
	) name4947 (
		\m4_s13_cyc_o_reg/NET0131 ,
		\rf_conf13_reg[8]/NET0131 ,
		\rf_conf13_reg[9]/NET0131 ,
		\s13_msel_arb0_state_reg[2]/NET0131 ,
		_w6848_
	);
	LUT4 #(
		.INIT('h0001)
	) name4948 (
		_w2339_,
		_w2342_,
		_w2343_,
		_w6848_,
		_w6849_
	);
	LUT3 #(
		.INIT('h01)
	) name4949 (
		_w2344_,
		_w2347_,
		_w2352_,
		_w6850_
	);
	LUT3 #(
		.INIT('h10)
	) name4950 (
		\s13_msel_arb0_state_reg[1]/NET0131 ,
		_w6849_,
		_w6850_,
		_w6851_
	);
	LUT3 #(
		.INIT('h01)
	) name4951 (
		_w2339_,
		_w2342_,
		_w2343_,
		_w6852_
	);
	LUT4 #(
		.INIT('h0001)
	) name4952 (
		_w2344_,
		_w2345_,
		_w2347_,
		_w2352_,
		_w6853_
	);
	LUT3 #(
		.INIT('ha2)
	) name4953 (
		_w2369_,
		_w6852_,
		_w6853_,
		_w6854_
	);
	LUT3 #(
		.INIT('h10)
	) name4954 (
		_w2347_,
		_w2352_,
		_w4481_,
		_w6855_
	);
	LUT3 #(
		.INIT('h45)
	) name4955 (
		\s13_msel_arb0_state_reg[0]/NET0131 ,
		_w6845_,
		_w6855_,
		_w6856_
	);
	LUT4 #(
		.INIT('h00fd)
	) name4956 (
		_w6847_,
		_w6851_,
		_w6854_,
		_w6856_,
		_w6857_
	);
	LUT4 #(
		.INIT('h0200)
	) name4957 (
		\m6_s13_cyc_o_reg/NET0131 ,
		\rf_conf13_reg[12]/NET0131 ,
		\rf_conf13_reg[13]/NET0131 ,
		\s13_msel_arb0_state_reg[1]/NET0131 ,
		_w6858_
	);
	LUT3 #(
		.INIT('ha8)
	) name4958 (
		\s13_msel_arb0_state_reg[2]/NET0131 ,
		_w6853_,
		_w6858_,
		_w6859_
	);
	LUT4 #(
		.INIT('h0504)
	) name4959 (
		\s13_msel_arb0_state_reg[1]/NET0131 ,
		\s13_msel_arb0_state_reg[2]/NET0131 ,
		_w6845_,
		_w6853_,
		_w6860_
	);
	LUT3 #(
		.INIT('hc8)
	) name4960 (
		_w2342_,
		_w4468_,
		_w6853_,
		_w6861_
	);
	LUT4 #(
		.INIT('h00ab)
	) name4961 (
		\s13_msel_arb0_state_reg[0]/NET0131 ,
		_w6859_,
		_w6860_,
		_w6861_,
		_w6862_
	);
	LUT2 #(
		.INIT('hb)
	) name4962 (
		_w6857_,
		_w6862_,
		_w6863_
	);
	LUT3 #(
		.INIT('h04)
	) name4963 (
		\s14_msel_arb0_state_reg[0]/NET0131 ,
		\s14_msel_arb0_state_reg[1]/NET0131 ,
		\s14_msel_arb0_state_reg[2]/NET0131 ,
		_w6864_
	);
	LUT4 #(
		.INIT('h0001)
	) name4964 (
		_w2376_,
		_w2377_,
		_w2379_,
		_w2380_,
		_w6865_
	);
	LUT2 #(
		.INIT('h4)
	) name4965 (
		_w2384_,
		_w4662_,
		_w6866_
	);
	LUT3 #(
		.INIT('h45)
	) name4966 (
		_w6864_,
		_w6865_,
		_w6866_,
		_w6867_
	);
	LUT4 #(
		.INIT('h0002)
	) name4967 (
		\m4_s14_cyc_o_reg/NET0131 ,
		\rf_conf14_reg[8]/NET0131 ,
		\rf_conf14_reg[9]/NET0131 ,
		\s14_msel_arb0_state_reg[2]/NET0131 ,
		_w6868_
	);
	LUT4 #(
		.INIT('h0001)
	) name4968 (
		_w2376_,
		_w2379_,
		_w2380_,
		_w6868_,
		_w6869_
	);
	LUT3 #(
		.INIT('h01)
	) name4969 (
		_w2381_,
		_w2384_,
		_w2389_,
		_w6870_
	);
	LUT3 #(
		.INIT('h10)
	) name4970 (
		\s14_msel_arb0_state_reg[1]/NET0131 ,
		_w6869_,
		_w6870_,
		_w6871_
	);
	LUT3 #(
		.INIT('h01)
	) name4971 (
		_w2376_,
		_w2379_,
		_w2380_,
		_w6872_
	);
	LUT4 #(
		.INIT('h0001)
	) name4972 (
		_w2381_,
		_w2382_,
		_w2384_,
		_w2389_,
		_w6873_
	);
	LUT3 #(
		.INIT('ha2)
	) name4973 (
		_w2406_,
		_w6872_,
		_w6873_,
		_w6874_
	);
	LUT3 #(
		.INIT('h10)
	) name4974 (
		_w2384_,
		_w2389_,
		_w4662_,
		_w6875_
	);
	LUT3 #(
		.INIT('h45)
	) name4975 (
		\s14_msel_arb0_state_reg[0]/NET0131 ,
		_w6865_,
		_w6875_,
		_w6876_
	);
	LUT4 #(
		.INIT('h00fd)
	) name4976 (
		_w6867_,
		_w6871_,
		_w6874_,
		_w6876_,
		_w6877_
	);
	LUT4 #(
		.INIT('h0200)
	) name4977 (
		\m6_s14_cyc_o_reg/NET0131 ,
		\rf_conf14_reg[12]/NET0131 ,
		\rf_conf14_reg[13]/NET0131 ,
		\s14_msel_arb0_state_reg[1]/NET0131 ,
		_w6878_
	);
	LUT3 #(
		.INIT('ha8)
	) name4978 (
		\s14_msel_arb0_state_reg[2]/NET0131 ,
		_w6873_,
		_w6878_,
		_w6879_
	);
	LUT4 #(
		.INIT('h0504)
	) name4979 (
		\s14_msel_arb0_state_reg[1]/NET0131 ,
		\s14_msel_arb0_state_reg[2]/NET0131 ,
		_w6865_,
		_w6873_,
		_w6880_
	);
	LUT3 #(
		.INIT('hc8)
	) name4980 (
		_w2379_,
		_w4649_,
		_w6873_,
		_w6881_
	);
	LUT4 #(
		.INIT('h00ab)
	) name4981 (
		\s14_msel_arb0_state_reg[0]/NET0131 ,
		_w6879_,
		_w6880_,
		_w6881_,
		_w6882_
	);
	LUT2 #(
		.INIT('hb)
	) name4982 (
		_w6877_,
		_w6882_,
		_w6883_
	);
	LUT3 #(
		.INIT('h51)
	) name4983 (
		_w2417_,
		_w2424_,
		_w2425_,
		_w6884_
	);
	LUT3 #(
		.INIT('h02)
	) name4984 (
		_w2420_,
		_w2421_,
		_w2425_,
		_w6885_
	);
	LUT4 #(
		.INIT('hfd00)
	) name4985 (
		\m4_s15_cyc_o_reg/NET0131 ,
		\rf_conf15_reg[8]/NET0131 ,
		\rf_conf15_reg[9]/NET0131 ,
		\s15_msel_arb0_state_reg[0]/NET0131 ,
		_w6886_
	);
	LUT3 #(
		.INIT('h10)
	) name4986 (
		_w2421_,
		_w2425_,
		_w6886_,
		_w6887_
	);
	LUT3 #(
		.INIT('h10)
	) name4987 (
		_w2413_,
		_w2416_,
		_w2452_,
		_w6888_
	);
	LUT4 #(
		.INIT('hfd00)
	) name4988 (
		_w6884_,
		_w6885_,
		_w6887_,
		_w6888_,
		_w6889_
	);
	LUT3 #(
		.INIT('h0d)
	) name4989 (
		_w2413_,
		_w2414_,
		_w2420_,
		_w6890_
	);
	LUT3 #(
		.INIT('h10)
	) name4990 (
		_w2414_,
		_w2416_,
		_w2417_,
		_w6891_
	);
	LUT4 #(
		.INIT('hfd00)
	) name4991 (
		\m0_s15_cyc_o_reg/NET0131 ,
		\rf_conf15_reg[0]/NET0131 ,
		\rf_conf15_reg[1]/NET0131 ,
		\s15_msel_arb0_state_reg[0]/NET0131 ,
		_w6892_
	);
	LUT3 #(
		.INIT('h10)
	) name4992 (
		_w2414_,
		_w2416_,
		_w6892_,
		_w6893_
	);
	LUT3 #(
		.INIT('h10)
	) name4993 (
		_w2421_,
		_w2424_,
		_w2448_,
		_w6894_
	);
	LUT4 #(
		.INIT('hfd00)
	) name4994 (
		_w6890_,
		_w6891_,
		_w6893_,
		_w6894_,
		_w6895_
	);
	LUT4 #(
		.INIT('h27ff)
	) name4995 (
		\s15_msel_arb0_state_reg[2]/NET0131 ,
		_w2413_,
		_w2424_,
		_w2447_,
		_w6896_
	);
	LUT2 #(
		.INIT('h8)
	) name4996 (
		_w2455_,
		_w6896_,
		_w6897_
	);
	LUT3 #(
		.INIT('h10)
	) name4997 (
		_w6889_,
		_w6895_,
		_w6897_,
		_w6898_
	);
	LUT2 #(
		.INIT('h4)
	) name4998 (
		_w2413_,
		_w2416_,
		_w6899_
	);
	LUT4 #(
		.INIT('h1101)
	) name4999 (
		_w2413_,
		_w2417_,
		_w2424_,
		_w2425_,
		_w6900_
	);
	LUT4 #(
		.INIT('hfd00)
	) name5000 (
		\m6_s15_cyc_o_reg/NET0131 ,
		\rf_conf15_reg[12]/NET0131 ,
		\rf_conf15_reg[13]/NET0131 ,
		\s15_msel_arb0_state_reg[0]/NET0131 ,
		_w6901_
	);
	LUT3 #(
		.INIT('h10)
	) name5001 (
		_w2421_,
		_w2425_,
		_w6901_,
		_w6902_
	);
	LUT3 #(
		.INIT('h10)
	) name5002 (
		_w2414_,
		_w2420_,
		_w2430_,
		_w6903_
	);
	LUT4 #(
		.INIT('hf100)
	) name5003 (
		_w6899_,
		_w6900_,
		_w6902_,
		_w6903_,
		_w6904_
	);
	LUT2 #(
		.INIT('h2)
	) name5004 (
		_w2421_,
		_w2424_,
		_w6905_
	);
	LUT4 #(
		.INIT('h000d)
	) name5005 (
		_w2413_,
		_w2414_,
		_w2420_,
		_w2424_,
		_w6906_
	);
	LUT4 #(
		.INIT('hfd00)
	) name5006 (
		\m2_s15_cyc_o_reg/NET0131 ,
		\rf_conf15_reg[4]/NET0131 ,
		\rf_conf15_reg[5]/NET0131 ,
		\s15_msel_arb0_state_reg[0]/NET0131 ,
		_w6907_
	);
	LUT3 #(
		.INIT('h10)
	) name5007 (
		_w2414_,
		_w2416_,
		_w6907_,
		_w6908_
	);
	LUT3 #(
		.INIT('h10)
	) name5008 (
		_w2417_,
		_w2425_,
		_w2454_,
		_w6909_
	);
	LUT4 #(
		.INIT('hf100)
	) name5009 (
		_w6905_,
		_w6906_,
		_w6908_,
		_w6909_,
		_w6910_
	);
	LUT2 #(
		.INIT('h1)
	) name5010 (
		_w6904_,
		_w6910_,
		_w6911_
	);
	LUT2 #(
		.INIT('h8)
	) name5011 (
		_w6898_,
		_w6911_,
		_w6912_
	);
	LUT2 #(
		.INIT('h2)
	) name5012 (
		_w2420_,
		_w2421_,
		_w6913_
	);
	LUT2 #(
		.INIT('h1)
	) name5013 (
		_w2414_,
		_w2421_,
		_w6914_
	);
	LUT4 #(
		.INIT('h0e0f)
	) name5014 (
		_w6899_,
		_w6900_,
		_w6913_,
		_w6914_,
		_w6915_
	);
	LUT2 #(
		.INIT('h4)
	) name5015 (
		_w2416_,
		_w2417_,
		_w6916_
	);
	LUT2 #(
		.INIT('h1)
	) name5016 (
		_w2416_,
		_w2425_,
		_w6917_
	);
	LUT4 #(
		.INIT('h0e0f)
	) name5017 (
		_w6905_,
		_w6906_,
		_w6916_,
		_w6917_,
		_w6918_
	);
	LUT4 #(
		.INIT('hfb73)
	) name5018 (
		\s15_msel_arb0_state_reg[2]/NET0131 ,
		_w2444_,
		_w6915_,
		_w6918_,
		_w6919_
	);
	LUT4 #(
		.INIT('h0002)
	) name5019 (
		\m0_s15_cyc_o_reg/NET0131 ,
		\rf_conf15_reg[0]/NET0131 ,
		\rf_conf15_reg[1]/NET0131 ,
		\s15_msel_arb0_state_reg[0]/NET0131 ,
		_w6920_
	);
	LUT3 #(
		.INIT('h0e)
	) name5020 (
		_w2424_,
		_w2425_,
		_w6920_,
		_w6921_
	);
	LUT4 #(
		.INIT('hfa02)
	) name5021 (
		_w2421_,
		_w2424_,
		_w2425_,
		_w6920_,
		_w6922_
	);
	LUT3 #(
		.INIT('h02)
	) name5022 (
		\s15_msel_arb0_state_reg[0]/NET0131 ,
		_w2414_,
		_w2416_,
		_w6923_
	);
	LUT4 #(
		.INIT('h0002)
	) name5023 (
		_w6890_,
		_w6891_,
		_w6921_,
		_w6923_,
		_w6924_
	);
	LUT3 #(
		.INIT('h02)
	) name5024 (
		_w2449_,
		_w6922_,
		_w6924_,
		_w6925_
	);
	LUT4 #(
		.INIT('h0200)
	) name5025 (
		\m4_s15_cyc_o_reg/NET0131 ,
		\rf_conf15_reg[8]/NET0131 ,
		\rf_conf15_reg[9]/NET0131 ,
		\s15_msel_arb0_state_reg[0]/NET0131 ,
		_w6926_
	);
	LUT3 #(
		.INIT('h0d)
	) name5026 (
		_w2413_,
		_w2414_,
		_w6926_,
		_w6927_
	);
	LUT4 #(
		.INIT('h00dc)
	) name5027 (
		_w2413_,
		_w2414_,
		_w2416_,
		_w6926_,
		_w6928_
	);
	LUT3 #(
		.INIT('h02)
	) name5028 (
		\s15_msel_arb0_state_reg[0]/NET0131 ,
		_w2421_,
		_w2425_,
		_w6929_
	);
	LUT4 #(
		.INIT('h0020)
	) name5029 (
		_w6884_,
		_w6885_,
		_w6927_,
		_w6929_,
		_w6930_
	);
	LUT3 #(
		.INIT('h02)
	) name5030 (
		_w2418_,
		_w6928_,
		_w6930_,
		_w6931_
	);
	LUT3 #(
		.INIT('h02)
	) name5031 (
		_w6919_,
		_w6925_,
		_w6931_,
		_w6932_
	);
	LUT2 #(
		.INIT('h7)
	) name5032 (
		_w6912_,
		_w6932_,
		_w6933_
	);
	LUT4 #(
		.INIT('h0001)
	) name5033 (
		_w2413_,
		_w2414_,
		_w2416_,
		_w2417_,
		_w6934_
	);
	LUT4 #(
		.INIT('h00fd)
	) name5034 (
		\m1_s15_cyc_o_reg/NET0131 ,
		\rf_conf15_reg[2]/NET0131 ,
		\rf_conf15_reg[3]/NET0131 ,
		\s15_msel_arb0_state_reg[2]/NET0131 ,
		_w6935_
	);
	LUT4 #(
		.INIT('h0100)
	) name5035 (
		_w2420_,
		_w2421_,
		_w6920_,
		_w6935_,
		_w6936_
	);
	LUT4 #(
		.INIT('h0001)
	) name5036 (
		_w2420_,
		_w2421_,
		_w2424_,
		_w2425_,
		_w6937_
	);
	LUT2 #(
		.INIT('h4)
	) name5037 (
		\s15_msel_arb0_state_reg[0]/NET0131 ,
		\s15_msel_arb0_state_reg[2]/NET0131 ,
		_w6938_
	);
	LUT4 #(
		.INIT('h0abb)
	) name5038 (
		_w6934_,
		_w6936_,
		_w6937_,
		_w6938_,
		_w6939_
	);
	LUT4 #(
		.INIT('h0100)
	) name5039 (
		_w2421_,
		_w2424_,
		_w2425_,
		_w2452_,
		_w6940_
	);
	LUT4 #(
		.INIT('h0002)
	) name5040 (
		\m2_s15_cyc_o_reg/NET0131 ,
		\rf_conf15_reg[4]/NET0131 ,
		\rf_conf15_reg[5]/NET0131 ,
		\s15_msel_arb0_state_reg[0]/NET0131 ,
		_w6941_
	);
	LUT2 #(
		.INIT('h2)
	) name5041 (
		\s15_msel_arb0_state_reg[1]/NET0131 ,
		\s15_msel_arb0_state_reg[2]/NET0131 ,
		_w6942_
	);
	LUT2 #(
		.INIT('h4)
	) name5042 (
		_w6941_,
		_w6942_,
		_w6943_
	);
	LUT4 #(
		.INIT('haeaf)
	) name5043 (
		_w2420_,
		_w6934_,
		_w6940_,
		_w6943_,
		_w6944_
	);
	LUT4 #(
		.INIT('hfe00)
	) name5044 (
		_w2413_,
		_w2416_,
		_w2417_,
		_w2452_,
		_w6945_
	);
	LUT4 #(
		.INIT('h0002)
	) name5045 (
		\m6_s15_cyc_o_reg/NET0131 ,
		\rf_conf15_reg[12]/NET0131 ,
		\rf_conf15_reg[13]/NET0131 ,
		\s15_msel_arb0_state_reg[0]/NET0131 ,
		_w6946_
	);
	LUT2 #(
		.INIT('h1)
	) name5046 (
		_w2417_,
		_w6946_,
		_w6947_
	);
	LUT2 #(
		.INIT('h8)
	) name5047 (
		\s15_msel_arb0_state_reg[1]/NET0131 ,
		\s15_msel_arb0_state_reg[2]/NET0131 ,
		_w6948_
	);
	LUT4 #(
		.INIT('h1033)
	) name5048 (
		_w6937_,
		_w6945_,
		_w6947_,
		_w6948_,
		_w6949_
	);
	LUT4 #(
		.INIT('h1fff)
	) name5049 (
		\s15_msel_arb0_state_reg[1]/NET0131 ,
		_w6939_,
		_w6944_,
		_w6949_,
		_w6950_
	);
	LUT4 #(
		.INIT('h1110)
	) name5050 (
		_w2891_,
		_w2892_,
		_w2898_,
		_w2899_,
		_w6951_
	);
	LUT3 #(
		.INIT('h02)
	) name5051 (
		\s15_msel_arb2_state_reg[2]/NET0131 ,
		_w2900_,
		_w4885_,
		_w6952_
	);
	LUT3 #(
		.INIT('hd0)
	) name5052 (
		_w2896_,
		_w6951_,
		_w6952_,
		_w6953_
	);
	LUT3 #(
		.INIT('ha2)
	) name5053 (
		\s15_msel_arb2_state_reg[1]/NET0131 ,
		_w4889_,
		_w4892_,
		_w6954_
	);
	LUT4 #(
		.INIT('h000e)
	) name5054 (
		_w2894_,
		_w2895_,
		_w2900_,
		_w2901_,
		_w6955_
	);
	LUT3 #(
		.INIT('h02)
	) name5055 (
		\s15_msel_arb2_state_reg[1]/NET0131 ,
		_w2898_,
		_w2899_,
		_w6956_
	);
	LUT3 #(
		.INIT('h45)
	) name5056 (
		_w6954_,
		_w6955_,
		_w6956_,
		_w6957_
	);
	LUT4 #(
		.INIT('h000e)
	) name5057 (
		_w2891_,
		_w2892_,
		_w2894_,
		_w2895_,
		_w6958_
	);
	LUT3 #(
		.INIT('h04)
	) name5058 (
		\s15_msel_arb2_state_reg[1]/NET0131 ,
		_w4860_,
		_w4871_,
		_w6959_
	);
	LUT3 #(
		.INIT('hd0)
	) name5059 (
		_w2902_,
		_w6958_,
		_w6959_,
		_w6960_
	);
	LUT4 #(
		.INIT('h1110)
	) name5060 (
		_w2898_,
		_w2899_,
		_w2900_,
		_w2901_,
		_w6961_
	);
	LUT3 #(
		.INIT('h04)
	) name5061 (
		\s15_msel_arb2_state_reg[1]/NET0131 ,
		_w4859_,
		_w4877_,
		_w6962_
	);
	LUT3 #(
		.INIT('hd0)
	) name5062 (
		_w2893_,
		_w6961_,
		_w6962_,
		_w6963_
	);
	LUT4 #(
		.INIT('hfff1)
	) name5063 (
		_w6953_,
		_w6957_,
		_w6960_,
		_w6963_,
		_w6964_
	);
	LUT4 #(
		.INIT('hfc54)
	) name5064 (
		_w2906_,
		_w2914_,
		_w2915_,
		_w2922_,
		_w6965_
	);
	LUT2 #(
		.INIT('h4)
	) name5065 (
		_w2905_,
		_w6965_,
		_w6966_
	);
	LUT2 #(
		.INIT('h2)
	) name5066 (
		_w2909_,
		_w4920_,
		_w6967_
	);
	LUT4 #(
		.INIT('h7f00)
	) name5067 (
		\m0_s15_cyc_o_reg/NET0131 ,
		\rf_conf15_reg[0]/NET0131 ,
		\rf_conf15_reg[1]/NET0131 ,
		\s15_msel_arb3_state_reg[1]/NET0131 ,
		_w6968_
	);
	LUT3 #(
		.INIT('h0d)
	) name5068 (
		_w2906_,
		_w2922_,
		_w6968_,
		_w6969_
	);
	LUT3 #(
		.INIT('h01)
	) name5069 (
		_w2905_,
		_w2912_,
		_w2913_,
		_w6970_
	);
	LUT3 #(
		.INIT('he0)
	) name5070 (
		_w6967_,
		_w6969_,
		_w6970_,
		_w6971_
	);
	LUT4 #(
		.INIT('heee0)
	) name5071 (
		_w2908_,
		_w2909_,
		_w2920_,
		_w2921_,
		_w6972_
	);
	LUT2 #(
		.INIT('h1)
	) name5072 (
		\s15_msel_arb3_state_reg[2]/NET0131 ,
		_w6972_,
		_w6973_
	);
	LUT3 #(
		.INIT('h10)
	) name5073 (
		_w6966_,
		_w6971_,
		_w6973_,
		_w6974_
	);
	LUT4 #(
		.INIT('h007f)
	) name5074 (
		\m6_s15_cyc_o_reg/NET0131 ,
		\rf_conf15_reg[12]/NET0131 ,
		\rf_conf15_reg[13]/NET0131 ,
		\s15_msel_arb3_state_reg[1]/NET0131 ,
		_w6975_
	);
	LUT3 #(
		.INIT('h0d)
	) name5075 (
		_w2915_,
		_w4923_,
		_w6975_,
		_w6976_
	);
	LUT3 #(
		.INIT('h02)
	) name5076 (
		_w2907_,
		_w2912_,
		_w6976_,
		_w6977_
	);
	LUT3 #(
		.INIT('h10)
	) name5077 (
		_w2905_,
		_w2906_,
		_w2914_,
		_w6978_
	);
	LUT3 #(
		.INIT('hc4)
	) name5078 (
		_w2910_,
		_w2928_,
		_w6978_,
		_w6979_
	);
	LUT4 #(
		.INIT('h002a)
	) name5079 (
		\s15_msel_arb3_state_reg[2]/NET0131 ,
		_w2914_,
		_w2920_,
		_w2926_,
		_w6980_
	);
	LUT3 #(
		.INIT('h10)
	) name5080 (
		_w6977_,
		_w6979_,
		_w6980_,
		_w6981_
	);
	LUT2 #(
		.INIT('he)
	) name5081 (
		_w6974_,
		_w6981_,
		_w6982_
	);
	LUT3 #(
		.INIT('h54)
	) name5082 (
		\s1_msel_arb0_state_reg[1]/NET0131 ,
		_w2648_,
		_w2668_,
		_w6983_
	);
	LUT4 #(
		.INIT('h0001)
	) name5083 (
		_w2644_,
		_w2645_,
		_w2653_,
		_w2654_,
		_w6984_
	);
	LUT2 #(
		.INIT('h8)
	) name5084 (
		\s1_msel_arb0_state_reg[0]/NET0131 ,
		\s1_msel_arb0_state_reg[1]/NET0131 ,
		_w6985_
	);
	LUT3 #(
		.INIT('h51)
	) name5085 (
		_w2649_,
		_w2650_,
		_w6985_,
		_w6986_
	);
	LUT4 #(
		.INIT('ha8aa)
	) name5086 (
		\s1_msel_arb0_state_reg[2]/NET0131 ,
		_w6983_,
		_w6984_,
		_w6986_,
		_w6987_
	);
	LUT4 #(
		.INIT('h0015)
	) name5087 (
		_w2645_,
		_w2654_,
		_w4969_,
		_w4948_,
		_w6988_
	);
	LUT4 #(
		.INIT('h0001)
	) name5088 (
		_w2647_,
		_w2648_,
		_w2649_,
		_w2650_,
		_w6989_
	);
	LUT4 #(
		.INIT('h00fd)
	) name5089 (
		\m3_s1_cyc_o_reg/NET0131 ,
		\rf_conf1_reg[6]/NET0131 ,
		\rf_conf1_reg[7]/NET0131 ,
		\s1_msel_arb0_state_reg[2]/NET0131 ,
		_w6990_
	);
	LUT4 #(
		.INIT('h0e00)
	) name5090 (
		_w6985_,
		_w6988_,
		_w6989_,
		_w6990_,
		_w6991_
	);
	LUT2 #(
		.INIT('he)
	) name5091 (
		_w6987_,
		_w6991_,
		_w6992_
	);
	LUT3 #(
		.INIT('h54)
	) name5092 (
		\s2_msel_arb0_state_reg[1]/NET0131 ,
		_w2687_,
		_w2707_,
		_w6993_
	);
	LUT4 #(
		.INIT('h0001)
	) name5093 (
		_w2683_,
		_w2684_,
		_w2692_,
		_w2693_,
		_w6994_
	);
	LUT2 #(
		.INIT('h8)
	) name5094 (
		\s2_msel_arb0_state_reg[0]/NET0131 ,
		\s2_msel_arb0_state_reg[1]/NET0131 ,
		_w6995_
	);
	LUT3 #(
		.INIT('h51)
	) name5095 (
		_w2688_,
		_w2689_,
		_w6995_,
		_w6996_
	);
	LUT4 #(
		.INIT('ha8aa)
	) name5096 (
		\s2_msel_arb0_state_reg[2]/NET0131 ,
		_w6993_,
		_w6994_,
		_w6996_,
		_w6997_
	);
	LUT4 #(
		.INIT('h0015)
	) name5097 (
		_w2684_,
		_w2693_,
		_w5131_,
		_w5110_,
		_w6998_
	);
	LUT4 #(
		.INIT('h0001)
	) name5098 (
		_w2686_,
		_w2687_,
		_w2688_,
		_w2689_,
		_w6999_
	);
	LUT4 #(
		.INIT('h00fd)
	) name5099 (
		\m3_s2_cyc_o_reg/NET0131 ,
		\rf_conf2_reg[6]/NET0131 ,
		\rf_conf2_reg[7]/NET0131 ,
		\s2_msel_arb0_state_reg[2]/NET0131 ,
		_w7000_
	);
	LUT4 #(
		.INIT('h0e00)
	) name5100 (
		_w6995_,
		_w6998_,
		_w6999_,
		_w7000_,
		_w7001_
	);
	LUT2 #(
		.INIT('he)
	) name5101 (
		_w6997_,
		_w7001_,
		_w7002_
	);
	LUT3 #(
		.INIT('h04)
	) name5102 (
		\s3_msel_arb0_state_reg[0]/NET0131 ,
		\s3_msel_arb0_state_reg[1]/NET0131 ,
		\s3_msel_arb0_state_reg[2]/NET0131 ,
		_w7003_
	);
	LUT4 #(
		.INIT('h0001)
	) name5103 (
		_w2459_,
		_w2460_,
		_w2462_,
		_w2463_,
		_w7004_
	);
	LUT2 #(
		.INIT('h4)
	) name5104 (
		_w2467_,
		_w5295_,
		_w7005_
	);
	LUT3 #(
		.INIT('h45)
	) name5105 (
		_w7003_,
		_w7004_,
		_w7005_,
		_w7006_
	);
	LUT4 #(
		.INIT('h0002)
	) name5106 (
		\m4_s3_cyc_o_reg/NET0131 ,
		\rf_conf3_reg[8]/NET0131 ,
		\rf_conf3_reg[9]/NET0131 ,
		\s3_msel_arb0_state_reg[2]/NET0131 ,
		_w7007_
	);
	LUT4 #(
		.INIT('h0001)
	) name5107 (
		_w2459_,
		_w2462_,
		_w2463_,
		_w7007_,
		_w7008_
	);
	LUT3 #(
		.INIT('h01)
	) name5108 (
		_w2464_,
		_w2467_,
		_w2472_,
		_w7009_
	);
	LUT3 #(
		.INIT('h10)
	) name5109 (
		\s3_msel_arb0_state_reg[1]/NET0131 ,
		_w7008_,
		_w7009_,
		_w7010_
	);
	LUT3 #(
		.INIT('h01)
	) name5110 (
		_w2459_,
		_w2462_,
		_w2463_,
		_w7011_
	);
	LUT4 #(
		.INIT('h0001)
	) name5111 (
		_w2464_,
		_w2465_,
		_w2467_,
		_w2472_,
		_w7012_
	);
	LUT3 #(
		.INIT('ha2)
	) name5112 (
		_w2489_,
		_w7011_,
		_w7012_,
		_w7013_
	);
	LUT3 #(
		.INIT('h10)
	) name5113 (
		_w2467_,
		_w2472_,
		_w5295_,
		_w7014_
	);
	LUT3 #(
		.INIT('h45)
	) name5114 (
		\s3_msel_arb0_state_reg[0]/NET0131 ,
		_w7004_,
		_w7014_,
		_w7015_
	);
	LUT4 #(
		.INIT('h00fd)
	) name5115 (
		_w7006_,
		_w7010_,
		_w7013_,
		_w7015_,
		_w7016_
	);
	LUT4 #(
		.INIT('h0200)
	) name5116 (
		\m6_s3_cyc_o_reg/NET0131 ,
		\rf_conf3_reg[12]/NET0131 ,
		\rf_conf3_reg[13]/NET0131 ,
		\s3_msel_arb0_state_reg[1]/NET0131 ,
		_w7017_
	);
	LUT3 #(
		.INIT('ha8)
	) name5117 (
		\s3_msel_arb0_state_reg[2]/NET0131 ,
		_w7012_,
		_w7017_,
		_w7018_
	);
	LUT4 #(
		.INIT('h0504)
	) name5118 (
		\s3_msel_arb0_state_reg[1]/NET0131 ,
		\s3_msel_arb0_state_reg[2]/NET0131 ,
		_w7004_,
		_w7012_,
		_w7019_
	);
	LUT3 #(
		.INIT('hc8)
	) name5119 (
		_w2462_,
		_w5282_,
		_w7012_,
		_w7020_
	);
	LUT4 #(
		.INIT('h00ab)
	) name5120 (
		\s3_msel_arb0_state_reg[0]/NET0131 ,
		_w7018_,
		_w7019_,
		_w7020_,
		_w7021_
	);
	LUT2 #(
		.INIT('hb)
	) name5121 (
		_w7016_,
		_w7021_,
		_w7022_
	);
	LUT3 #(
		.INIT('h04)
	) name5122 (
		\s4_msel_arb0_state_reg[0]/NET0131 ,
		\s4_msel_arb0_state_reg[1]/NET0131 ,
		\s4_msel_arb0_state_reg[2]/NET0131 ,
		_w7023_
	);
	LUT4 #(
		.INIT('h0001)
	) name5123 (
		_w2496_,
		_w2497_,
		_w2499_,
		_w2500_,
		_w7024_
	);
	LUT2 #(
		.INIT('h4)
	) name5124 (
		_w2504_,
		_w5470_,
		_w7025_
	);
	LUT3 #(
		.INIT('h45)
	) name5125 (
		_w7023_,
		_w7024_,
		_w7025_,
		_w7026_
	);
	LUT4 #(
		.INIT('h0002)
	) name5126 (
		\m4_s4_cyc_o_reg/NET0131 ,
		\rf_conf4_reg[8]/NET0131 ,
		\rf_conf4_reg[9]/NET0131 ,
		\s4_msel_arb0_state_reg[2]/NET0131 ,
		_w7027_
	);
	LUT4 #(
		.INIT('h0001)
	) name5127 (
		_w2496_,
		_w2499_,
		_w2500_,
		_w7027_,
		_w7028_
	);
	LUT3 #(
		.INIT('h01)
	) name5128 (
		_w2501_,
		_w2504_,
		_w2509_,
		_w7029_
	);
	LUT3 #(
		.INIT('h10)
	) name5129 (
		\s4_msel_arb0_state_reg[1]/NET0131 ,
		_w7028_,
		_w7029_,
		_w7030_
	);
	LUT3 #(
		.INIT('h01)
	) name5130 (
		_w2496_,
		_w2499_,
		_w2500_,
		_w7031_
	);
	LUT4 #(
		.INIT('h0001)
	) name5131 (
		_w2501_,
		_w2502_,
		_w2504_,
		_w2509_,
		_w7032_
	);
	LUT3 #(
		.INIT('ha2)
	) name5132 (
		_w2526_,
		_w7031_,
		_w7032_,
		_w7033_
	);
	LUT3 #(
		.INIT('h10)
	) name5133 (
		_w2504_,
		_w2509_,
		_w5470_,
		_w7034_
	);
	LUT3 #(
		.INIT('h45)
	) name5134 (
		\s4_msel_arb0_state_reg[0]/NET0131 ,
		_w7024_,
		_w7034_,
		_w7035_
	);
	LUT4 #(
		.INIT('h00fd)
	) name5135 (
		_w7026_,
		_w7030_,
		_w7033_,
		_w7035_,
		_w7036_
	);
	LUT4 #(
		.INIT('h0200)
	) name5136 (
		\m6_s4_cyc_o_reg/NET0131 ,
		\rf_conf4_reg[12]/NET0131 ,
		\rf_conf4_reg[13]/NET0131 ,
		\s4_msel_arb0_state_reg[1]/NET0131 ,
		_w7037_
	);
	LUT3 #(
		.INIT('ha8)
	) name5137 (
		\s4_msel_arb0_state_reg[2]/NET0131 ,
		_w7032_,
		_w7037_,
		_w7038_
	);
	LUT4 #(
		.INIT('h0504)
	) name5138 (
		\s4_msel_arb0_state_reg[1]/NET0131 ,
		\s4_msel_arb0_state_reg[2]/NET0131 ,
		_w7024_,
		_w7032_,
		_w7039_
	);
	LUT3 #(
		.INIT('hc8)
	) name5139 (
		_w2499_,
		_w5457_,
		_w7032_,
		_w7040_
	);
	LUT4 #(
		.INIT('h00ab)
	) name5140 (
		\s4_msel_arb0_state_reg[0]/NET0131 ,
		_w7038_,
		_w7039_,
		_w7040_,
		_w7041_
	);
	LUT2 #(
		.INIT('hb)
	) name5141 (
		_w7036_,
		_w7041_,
		_w7042_
	);
	LUT3 #(
		.INIT('h04)
	) name5142 (
		\s5_msel_arb0_state_reg[0]/NET0131 ,
		\s5_msel_arb0_state_reg[1]/NET0131 ,
		\s5_msel_arb0_state_reg[2]/NET0131 ,
		_w7043_
	);
	LUT4 #(
		.INIT('h0001)
	) name5143 (
		_w2533_,
		_w2534_,
		_w2536_,
		_w2537_,
		_w7044_
	);
	LUT2 #(
		.INIT('h4)
	) name5144 (
		_w2541_,
		_w5647_,
		_w7045_
	);
	LUT3 #(
		.INIT('h45)
	) name5145 (
		_w7043_,
		_w7044_,
		_w7045_,
		_w7046_
	);
	LUT4 #(
		.INIT('h0002)
	) name5146 (
		\m4_s5_cyc_o_reg/NET0131 ,
		\rf_conf5_reg[8]/NET0131 ,
		\rf_conf5_reg[9]/NET0131 ,
		\s5_msel_arb0_state_reg[2]/NET0131 ,
		_w7047_
	);
	LUT4 #(
		.INIT('h0001)
	) name5147 (
		_w2533_,
		_w2536_,
		_w2537_,
		_w7047_,
		_w7048_
	);
	LUT3 #(
		.INIT('h01)
	) name5148 (
		_w2538_,
		_w2541_,
		_w2546_,
		_w7049_
	);
	LUT3 #(
		.INIT('h10)
	) name5149 (
		\s5_msel_arb0_state_reg[1]/NET0131 ,
		_w7048_,
		_w7049_,
		_w7050_
	);
	LUT3 #(
		.INIT('h01)
	) name5150 (
		_w2533_,
		_w2536_,
		_w2537_,
		_w7051_
	);
	LUT4 #(
		.INIT('h0001)
	) name5151 (
		_w2538_,
		_w2539_,
		_w2541_,
		_w2546_,
		_w7052_
	);
	LUT3 #(
		.INIT('ha2)
	) name5152 (
		_w2563_,
		_w7051_,
		_w7052_,
		_w7053_
	);
	LUT3 #(
		.INIT('h10)
	) name5153 (
		_w2541_,
		_w2546_,
		_w5647_,
		_w7054_
	);
	LUT3 #(
		.INIT('h45)
	) name5154 (
		\s5_msel_arb0_state_reg[0]/NET0131 ,
		_w7044_,
		_w7054_,
		_w7055_
	);
	LUT4 #(
		.INIT('h00fd)
	) name5155 (
		_w7046_,
		_w7050_,
		_w7053_,
		_w7055_,
		_w7056_
	);
	LUT4 #(
		.INIT('h0200)
	) name5156 (
		\m6_s5_cyc_o_reg/NET0131 ,
		\rf_conf5_reg[12]/NET0131 ,
		\rf_conf5_reg[13]/NET0131 ,
		\s5_msel_arb0_state_reg[1]/NET0131 ,
		_w7057_
	);
	LUT3 #(
		.INIT('ha8)
	) name5157 (
		\s5_msel_arb0_state_reg[2]/NET0131 ,
		_w7052_,
		_w7057_,
		_w7058_
	);
	LUT4 #(
		.INIT('h0504)
	) name5158 (
		\s5_msel_arb0_state_reg[1]/NET0131 ,
		\s5_msel_arb0_state_reg[2]/NET0131 ,
		_w7044_,
		_w7052_,
		_w7059_
	);
	LUT3 #(
		.INIT('hc8)
	) name5159 (
		_w2536_,
		_w5634_,
		_w7052_,
		_w7060_
	);
	LUT4 #(
		.INIT('h00ab)
	) name5160 (
		\s5_msel_arb0_state_reg[0]/NET0131 ,
		_w7058_,
		_w7059_,
		_w7060_,
		_w7061_
	);
	LUT2 #(
		.INIT('hb)
	) name5161 (
		_w7056_,
		_w7061_,
		_w7062_
	);
	LUT3 #(
		.INIT('h04)
	) name5162 (
		\s6_msel_arb0_state_reg[0]/NET0131 ,
		\s6_msel_arb0_state_reg[1]/NET0131 ,
		\s6_msel_arb0_state_reg[2]/NET0131 ,
		_w7063_
	);
	LUT4 #(
		.INIT('h0001)
	) name5163 (
		_w2570_,
		_w2571_,
		_w2573_,
		_w2574_,
		_w7064_
	);
	LUT2 #(
		.INIT('h4)
	) name5164 (
		_w2578_,
		_w5809_,
		_w7065_
	);
	LUT3 #(
		.INIT('h45)
	) name5165 (
		_w7063_,
		_w7064_,
		_w7065_,
		_w7066_
	);
	LUT4 #(
		.INIT('h0002)
	) name5166 (
		\m4_s6_cyc_o_reg/NET0131 ,
		\rf_conf6_reg[8]/NET0131 ,
		\rf_conf6_reg[9]/NET0131 ,
		\s6_msel_arb0_state_reg[2]/NET0131 ,
		_w7067_
	);
	LUT4 #(
		.INIT('h0001)
	) name5167 (
		_w2570_,
		_w2573_,
		_w2574_,
		_w7067_,
		_w7068_
	);
	LUT3 #(
		.INIT('h01)
	) name5168 (
		_w2575_,
		_w2578_,
		_w2583_,
		_w7069_
	);
	LUT3 #(
		.INIT('h10)
	) name5169 (
		\s6_msel_arb0_state_reg[1]/NET0131 ,
		_w7068_,
		_w7069_,
		_w7070_
	);
	LUT3 #(
		.INIT('h01)
	) name5170 (
		_w2570_,
		_w2573_,
		_w2574_,
		_w7071_
	);
	LUT4 #(
		.INIT('h0001)
	) name5171 (
		_w2575_,
		_w2576_,
		_w2578_,
		_w2583_,
		_w7072_
	);
	LUT3 #(
		.INIT('ha2)
	) name5172 (
		_w2600_,
		_w7071_,
		_w7072_,
		_w7073_
	);
	LUT3 #(
		.INIT('h10)
	) name5173 (
		_w2578_,
		_w2583_,
		_w5809_,
		_w7074_
	);
	LUT3 #(
		.INIT('h45)
	) name5174 (
		\s6_msel_arb0_state_reg[0]/NET0131 ,
		_w7064_,
		_w7074_,
		_w7075_
	);
	LUT4 #(
		.INIT('h00fd)
	) name5175 (
		_w7066_,
		_w7070_,
		_w7073_,
		_w7075_,
		_w7076_
	);
	LUT4 #(
		.INIT('h0200)
	) name5176 (
		\m6_s6_cyc_o_reg/NET0131 ,
		\rf_conf6_reg[12]/NET0131 ,
		\rf_conf6_reg[13]/NET0131 ,
		\s6_msel_arb0_state_reg[1]/NET0131 ,
		_w7077_
	);
	LUT3 #(
		.INIT('ha8)
	) name5177 (
		\s6_msel_arb0_state_reg[2]/NET0131 ,
		_w7072_,
		_w7077_,
		_w7078_
	);
	LUT4 #(
		.INIT('h0504)
	) name5178 (
		\s6_msel_arb0_state_reg[1]/NET0131 ,
		\s6_msel_arb0_state_reg[2]/NET0131 ,
		_w7064_,
		_w7072_,
		_w7079_
	);
	LUT3 #(
		.INIT('hc8)
	) name5179 (
		_w2573_,
		_w5796_,
		_w7072_,
		_w7080_
	);
	LUT4 #(
		.INIT('h00ab)
	) name5180 (
		\s6_msel_arb0_state_reg[0]/NET0131 ,
		_w7078_,
		_w7079_,
		_w7080_,
		_w7081_
	);
	LUT2 #(
		.INIT('hb)
	) name5181 (
		_w7076_,
		_w7081_,
		_w7082_
	);
	LUT3 #(
		.INIT('h54)
	) name5182 (
		\s7_msel_arb0_state_reg[1]/NET0131 ,
		_w2726_,
		_w2746_,
		_w7083_
	);
	LUT4 #(
		.INIT('h0001)
	) name5183 (
		_w2722_,
		_w2723_,
		_w2731_,
		_w2732_,
		_w7084_
	);
	LUT2 #(
		.INIT('h8)
	) name5184 (
		\s7_msel_arb0_state_reg[0]/NET0131 ,
		\s7_msel_arb0_state_reg[1]/NET0131 ,
		_w7085_
	);
	LUT3 #(
		.INIT('h51)
	) name5185 (
		_w2727_,
		_w2728_,
		_w7085_,
		_w7086_
	);
	LUT4 #(
		.INIT('ha8aa)
	) name5186 (
		\s7_msel_arb0_state_reg[2]/NET0131 ,
		_w7083_,
		_w7084_,
		_w7086_,
		_w7087_
	);
	LUT4 #(
		.INIT('h0015)
	) name5187 (
		_w2723_,
		_w2732_,
		_w5979_,
		_w5958_,
		_w7088_
	);
	LUT4 #(
		.INIT('h0001)
	) name5188 (
		_w2725_,
		_w2726_,
		_w2727_,
		_w2728_,
		_w7089_
	);
	LUT4 #(
		.INIT('h00fd)
	) name5189 (
		\m3_s7_cyc_o_reg/NET0131 ,
		\rf_conf7_reg[6]/NET0131 ,
		\rf_conf7_reg[7]/NET0131 ,
		\s7_msel_arb0_state_reg[2]/NET0131 ,
		_w7090_
	);
	LUT4 #(
		.INIT('h0e00)
	) name5190 (
		_w7085_,
		_w7088_,
		_w7089_,
		_w7090_,
		_w7091_
	);
	LUT2 #(
		.INIT('he)
	) name5191 (
		_w7087_,
		_w7091_,
		_w7092_
	);
	LUT3 #(
		.INIT('h04)
	) name5192 (
		\s8_msel_arb0_state_reg[0]/NET0131 ,
		\s8_msel_arb0_state_reg[1]/NET0131 ,
		\s8_msel_arb0_state_reg[2]/NET0131 ,
		_w7093_
	);
	LUT4 #(
		.INIT('h0001)
	) name5193 (
		_w2607_,
		_w2608_,
		_w2610_,
		_w2611_,
		_w7094_
	);
	LUT2 #(
		.INIT('h4)
	) name5194 (
		_w2615_,
		_w6155_,
		_w7095_
	);
	LUT3 #(
		.INIT('h45)
	) name5195 (
		_w7093_,
		_w7094_,
		_w7095_,
		_w7096_
	);
	LUT4 #(
		.INIT('h0002)
	) name5196 (
		\m4_s8_cyc_o_reg/NET0131 ,
		\rf_conf8_reg[8]/NET0131 ,
		\rf_conf8_reg[9]/NET0131 ,
		\s8_msel_arb0_state_reg[2]/NET0131 ,
		_w7097_
	);
	LUT4 #(
		.INIT('h0001)
	) name5197 (
		_w2607_,
		_w2610_,
		_w2611_,
		_w7097_,
		_w7098_
	);
	LUT3 #(
		.INIT('h01)
	) name5198 (
		_w2612_,
		_w2615_,
		_w2620_,
		_w7099_
	);
	LUT3 #(
		.INIT('h10)
	) name5199 (
		\s8_msel_arb0_state_reg[1]/NET0131 ,
		_w7098_,
		_w7099_,
		_w7100_
	);
	LUT3 #(
		.INIT('h01)
	) name5200 (
		_w2607_,
		_w2610_,
		_w2611_,
		_w7101_
	);
	LUT4 #(
		.INIT('h0001)
	) name5201 (
		_w2612_,
		_w2613_,
		_w2615_,
		_w2620_,
		_w7102_
	);
	LUT3 #(
		.INIT('hd0)
	) name5202 (
		_w7101_,
		_w7102_,
		_w2637_,
		_w7103_
	);
	LUT3 #(
		.INIT('h10)
	) name5203 (
		_w2615_,
		_w2620_,
		_w6155_,
		_w7104_
	);
	LUT3 #(
		.INIT('h45)
	) name5204 (
		\s8_msel_arb0_state_reg[0]/NET0131 ,
		_w7094_,
		_w7104_,
		_w7105_
	);
	LUT4 #(
		.INIT('h00fd)
	) name5205 (
		_w7096_,
		_w7100_,
		_w7103_,
		_w7105_,
		_w7106_
	);
	LUT4 #(
		.INIT('h0200)
	) name5206 (
		\m6_s8_cyc_o_reg/NET0131 ,
		\rf_conf8_reg[12]/NET0131 ,
		\rf_conf8_reg[13]/NET0131 ,
		\s8_msel_arb0_state_reg[1]/NET0131 ,
		_w7107_
	);
	LUT3 #(
		.INIT('ha8)
	) name5207 (
		\s8_msel_arb0_state_reg[2]/NET0131 ,
		_w7102_,
		_w7107_,
		_w7108_
	);
	LUT4 #(
		.INIT('h0504)
	) name5208 (
		\s8_msel_arb0_state_reg[1]/NET0131 ,
		\s8_msel_arb0_state_reg[2]/NET0131 ,
		_w7094_,
		_w7102_,
		_w7109_
	);
	LUT3 #(
		.INIT('hc8)
	) name5209 (
		_w2610_,
		_w6142_,
		_w7102_,
		_w7110_
	);
	LUT4 #(
		.INIT('h00ab)
	) name5210 (
		\s8_msel_arb0_state_reg[0]/NET0131 ,
		_w7108_,
		_w7109_,
		_w7110_,
		_w7111_
	);
	LUT2 #(
		.INIT('hb)
	) name5211 (
		_w7106_,
		_w7111_,
		_w7112_
	);
	LUT3 #(
		.INIT('h54)
	) name5212 (
		\s9_msel_arb0_state_reg[1]/NET0131 ,
		_w2765_,
		_w2785_,
		_w7113_
	);
	LUT4 #(
		.INIT('h0001)
	) name5213 (
		_w2761_,
		_w2762_,
		_w2770_,
		_w2771_,
		_w7114_
	);
	LUT2 #(
		.INIT('h8)
	) name5214 (
		\s9_msel_arb0_state_reg[0]/NET0131 ,
		\s9_msel_arb0_state_reg[1]/NET0131 ,
		_w7115_
	);
	LUT3 #(
		.INIT('h51)
	) name5215 (
		_w2766_,
		_w2767_,
		_w7115_,
		_w7116_
	);
	LUT4 #(
		.INIT('ha8aa)
	) name5216 (
		\s9_msel_arb0_state_reg[2]/NET0131 ,
		_w7113_,
		_w7114_,
		_w7116_,
		_w7117_
	);
	LUT4 #(
		.INIT('h0015)
	) name5217 (
		_w2762_,
		_w2771_,
		_w6326_,
		_w6305_,
		_w7118_
	);
	LUT4 #(
		.INIT('h0001)
	) name5218 (
		_w2764_,
		_w2765_,
		_w2766_,
		_w2767_,
		_w7119_
	);
	LUT4 #(
		.INIT('h00fd)
	) name5219 (
		\m3_s9_cyc_o_reg/NET0131 ,
		\rf_conf9_reg[6]/NET0131 ,
		\rf_conf9_reg[7]/NET0131 ,
		\s9_msel_arb0_state_reg[2]/NET0131 ,
		_w7120_
	);
	LUT4 #(
		.INIT('h0e00)
	) name5220 (
		_w7115_,
		_w7118_,
		_w7119_,
		_w7120_,
		_w7121_
	);
	LUT2 #(
		.INIT('he)
	) name5221 (
		_w7117_,
		_w7121_,
		_w7122_
	);
	LUT3 #(
		.INIT('h54)
	) name5222 (
		\s0_msel_arb0_state_reg[1]/NET0131 ,
		_w2804_,
		_w2824_,
		_w7123_
	);
	LUT4 #(
		.INIT('h0001)
	) name5223 (
		_w2800_,
		_w2801_,
		_w2809_,
		_w2810_,
		_w7124_
	);
	LUT2 #(
		.INIT('h8)
	) name5224 (
		\s0_msel_arb0_state_reg[0]/NET0131 ,
		\s0_msel_arb0_state_reg[1]/NET0131 ,
		_w7125_
	);
	LUT3 #(
		.INIT('h51)
	) name5225 (
		_w2805_,
		_w2806_,
		_w7125_,
		_w7126_
	);
	LUT4 #(
		.INIT('ha8aa)
	) name5226 (
		\s0_msel_arb0_state_reg[2]/NET0131 ,
		_w7123_,
		_w7124_,
		_w7126_,
		_w7127_
	);
	LUT4 #(
		.INIT('h0015)
	) name5227 (
		_w2801_,
		_w2810_,
		_w6499_,
		_w6478_,
		_w7128_
	);
	LUT4 #(
		.INIT('h0001)
	) name5228 (
		_w2803_,
		_w2804_,
		_w2805_,
		_w2806_,
		_w7129_
	);
	LUT4 #(
		.INIT('h00fd)
	) name5229 (
		\m3_s0_cyc_o_reg/NET0131 ,
		\rf_conf0_reg[6]/NET0131 ,
		\rf_conf0_reg[7]/NET0131 ,
		\s0_msel_arb0_state_reg[2]/NET0131 ,
		_w7130_
	);
	LUT4 #(
		.INIT('h0e00)
	) name5230 (
		_w7125_,
		_w7128_,
		_w7129_,
		_w7130_,
		_w7131_
	);
	LUT2 #(
		.INIT('he)
	) name5231 (
		_w7127_,
		_w7131_,
		_w7132_
	);
	LUT3 #(
		.INIT('h54)
	) name5232 (
		\s10_msel_arb2_state_reg[2]/NET0131 ,
		_w4026_,
		_w4027_,
		_w7133_
	);
	LUT4 #(
		.INIT('h1110)
	) name5233 (
		_w4031_,
		_w4032_,
		_w4034_,
		_w4035_,
		_w7134_
	);
	LUT4 #(
		.INIT('h0d0c)
	) name5234 (
		\s10_msel_arb2_state_reg[0]/NET0131 ,
		_w6674_,
		_w7133_,
		_w7134_,
		_w7135_
	);
	LUT3 #(
		.INIT('h01)
	) name5235 (
		\s10_msel_arb2_state_reg[1]/NET0131 ,
		_w4031_,
		_w4032_,
		_w7136_
	);
	LUT2 #(
		.INIT('h8)
	) name5236 (
		_w6670_,
		_w7136_,
		_w7137_
	);
	LUT3 #(
		.INIT('ha8)
	) name5237 (
		\s10_msel_arb2_state_reg[2]/NET0131 ,
		_w4031_,
		_w4032_,
		_w7138_
	);
	LUT4 #(
		.INIT('h1110)
	) name5238 (
		_w4026_,
		_w4027_,
		_w4030_,
		_w4038_,
		_w7139_
	);
	LUT4 #(
		.INIT('h0d0c)
	) name5239 (
		\s10_msel_arb2_state_reg[0]/NET0131 ,
		_w6676_,
		_w7138_,
		_w7139_,
		_w7140_
	);
	LUT2 #(
		.INIT('h8)
	) name5240 (
		_w4031_,
		_w4047_,
		_w7141_
	);
	LUT3 #(
		.INIT('h10)
	) name5241 (
		_w4034_,
		_w4035_,
		_w4047_,
		_w7142_
	);
	LUT4 #(
		.INIT('h080a)
	) name5242 (
		\s10_msel_arb2_state_reg[0]/NET0131 ,
		_w7139_,
		_w7141_,
		_w7142_,
		_w7143_
	);
	LUT4 #(
		.INIT('h0001)
	) name5243 (
		_w7135_,
		_w7137_,
		_w7140_,
		_w7143_,
		_w7144_
	);
	LUT4 #(
		.INIT('h5400)
	) name5244 (
		_w4030_,
		_w4031_,
		_w4032_,
		_w4061_,
		_w7145_
	);
	LUT4 #(
		.INIT('hdf00)
	) name5245 (
		\m4_s10_cyc_o_reg/NET0131 ,
		\rf_conf10_reg[8]/NET0131 ,
		\rf_conf10_reg[9]/NET0131 ,
		\s10_msel_arb2_state_reg[1]/NET0131 ,
		_w7146_
	);
	LUT3 #(
		.INIT('h01)
	) name5246 (
		_w4026_,
		_w4027_,
		_w7146_,
		_w7147_
	);
	LUT4 #(
		.INIT('h0100)
	) name5247 (
		_w4030_,
		_w4034_,
		_w4035_,
		_w4061_,
		_w7148_
	);
	LUT3 #(
		.INIT('h45)
	) name5248 (
		_w7145_,
		_w7147_,
		_w7148_,
		_w7149_
	);
	LUT4 #(
		.INIT('h2000)
	) name5249 (
		\m3_s10_cyc_o_reg/NET0131 ,
		\rf_conf10_reg[6]/NET0131 ,
		\rf_conf10_reg[7]/NET0131 ,
		\s10_msel_arb2_state_reg[1]/NET0131 ,
		_w7150_
	);
	LUT3 #(
		.INIT('h02)
	) name5250 (
		\s10_msel_arb2_state_reg[1]/NET0131 ,
		_w4030_,
		_w4038_,
		_w7151_
	);
	LUT3 #(
		.INIT('h23)
	) name5251 (
		_w7134_,
		_w7150_,
		_w7151_,
		_w7152_
	);
	LUT4 #(
		.INIT('h0054)
	) name5252 (
		_w4030_,
		_w4031_,
		_w4032_,
		_w4038_,
		_w7153_
	);
	LUT4 #(
		.INIT('h00df)
	) name5253 (
		\m1_s10_cyc_o_reg/NET0131 ,
		\rf_conf10_reg[2]/NET0131 ,
		\rf_conf10_reg[3]/NET0131 ,
		\s10_msel_arb2_state_reg[1]/NET0131 ,
		_w7154_
	);
	LUT3 #(
		.INIT('hd0)
	) name5254 (
		_w6670_,
		_w7153_,
		_w7154_,
		_w7155_
	);
	LUT2 #(
		.INIT('h2)
	) name5255 (
		\s10_msel_arb2_state_reg[0]/NET0131 ,
		\s10_msel_arb2_state_reg[2]/NET0131 ,
		_w7156_
	);
	LUT4 #(
		.INIT('h08aa)
	) name5256 (
		_w7149_,
		_w7152_,
		_w7155_,
		_w7156_,
		_w7157_
	);
	LUT2 #(
		.INIT('hb)
	) name5257 (
		_w7144_,
		_w7157_,
		_w7158_
	);
	LUT4 #(
		.INIT('h4447)
	) name5258 (
		\s10_msel_arb3_state_reg[0]/NET0131 ,
		\s10_msel_arb3_state_reg[2]/NET0131 ,
		_w3165_,
		_w4095_,
		_w7159_
	);
	LUT4 #(
		.INIT('h1110)
	) name5259 (
		_w3153_,
		_w3154_,
		_w3160_,
		_w3161_,
		_w7160_
	);
	LUT2 #(
		.INIT('h8)
	) name5260 (
		_w7159_,
		_w7160_,
		_w7161_
	);
	LUT4 #(
		.INIT('hccc8)
	) name5261 (
		\s10_msel_arb3_state_reg[0]/NET0131 ,
		\s10_msel_arb3_state_reg[2]/NET0131 ,
		_w3153_,
		_w3154_,
		_w7162_
	);
	LUT4 #(
		.INIT('h000e)
	) name5262 (
		_w3163_,
		_w3164_,
		_w3165_,
		_w4095_,
		_w7163_
	);
	LUT2 #(
		.INIT('h4)
	) name5263 (
		_w7162_,
		_w7163_,
		_w7164_
	);
	LUT2 #(
		.INIT('h4)
	) name5264 (
		_w3153_,
		_w3156_,
		_w7165_
	);
	LUT4 #(
		.INIT('h000e)
	) name5265 (
		_w3163_,
		_w3164_,
		_w3165_,
		_w3166_,
		_w7166_
	);
	LUT3 #(
		.INIT('hc4)
	) name5266 (
		_w3162_,
		_w7165_,
		_w7166_,
		_w7167_
	);
	LUT4 #(
		.INIT('h5554)
	) name5267 (
		\s10_msel_arb3_state_reg[1]/NET0131 ,
		_w7161_,
		_w7164_,
		_w7167_,
		_w7168_
	);
	LUT3 #(
		.INIT('ha8)
	) name5268 (
		\s10_msel_arb3_state_reg[2]/NET0131 ,
		_w3165_,
		_w3166_,
		_w7169_
	);
	LUT4 #(
		.INIT('h000e)
	) name5269 (
		_w3153_,
		_w3154_,
		_w3163_,
		_w3164_,
		_w7170_
	);
	LUT3 #(
		.INIT('h54)
	) name5270 (
		_w4117_,
		_w7169_,
		_w7170_,
		_w7171_
	);
	LUT3 #(
		.INIT('h0e)
	) name5271 (
		_w3165_,
		_w3166_,
		_w3171_,
		_w7172_
	);
	LUT2 #(
		.INIT('h4)
	) name5272 (
		_w3164_,
		_w4104_,
		_w7173_
	);
	LUT2 #(
		.INIT('h1)
	) name5273 (
		_w3161_,
		_w3163_,
		_w7174_
	);
	LUT3 #(
		.INIT('he0)
	) name5274 (
		_w7172_,
		_w7173_,
		_w7174_,
		_w7175_
	);
	LUT3 #(
		.INIT('h0e)
	) name5275 (
		_w3153_,
		_w3154_,
		_w3163_,
		_w7176_
	);
	LUT3 #(
		.INIT('h2a)
	) name5276 (
		\s10_msel_arb3_state_reg[1]/NET0131 ,
		_w3172_,
		_w7176_,
		_w7177_
	);
	LUT4 #(
		.INIT('hab00)
	) name5277 (
		_w3160_,
		_w7171_,
		_w7175_,
		_w7177_,
		_w7178_
	);
	LUT2 #(
		.INIT('he)
	) name5278 (
		_w7168_,
		_w7178_,
		_w7179_
	);
	LUT4 #(
		.INIT('h0020)
	) name5279 (
		\m2_s11_cyc_o_reg/NET0131 ,
		\rf_conf11_reg[4]/NET0131 ,
		\rf_conf11_reg[5]/NET0131 ,
		\s11_msel_arb2_state_reg[0]/NET0131 ,
		_w7180_
	);
	LUT3 #(
		.INIT('h01)
	) name5280 (
		_w3183_,
		_w3184_,
		_w7180_,
		_w7181_
	);
	LUT4 #(
		.INIT('h2000)
	) name5281 (
		\m3_s11_cyc_o_reg/NET0131 ,
		\rf_conf11_reg[6]/NET0131 ,
		\rf_conf11_reg[7]/NET0131 ,
		\s11_msel_arb2_state_reg[0]/NET0131 ,
		_w7182_
	);
	LUT2 #(
		.INIT('h1)
	) name5282 (
		\s11_msel_arb2_state_reg[2]/NET0131 ,
		_w7182_,
		_w7183_
	);
	LUT4 #(
		.INIT('h00df)
	) name5283 (
		\m2_s11_cyc_o_reg/NET0131 ,
		\rf_conf11_reg[4]/NET0131 ,
		\rf_conf11_reg[5]/NET0131 ,
		\s11_msel_arb2_state_reg[1]/NET0131 ,
		_w7184_
	);
	LUT3 #(
		.INIT('h01)
	) name5284 (
		_w3194_,
		_w3198_,
		_w7184_,
		_w7185_
	);
	LUT4 #(
		.INIT('hcf4f)
	) name5285 (
		_w3187_,
		_w7181_,
		_w7183_,
		_w7185_,
		_w7186_
	);
	LUT4 #(
		.INIT('haaa2)
	) name5286 (
		\s11_msel_arb2_state_reg[1]/NET0131 ,
		\s11_msel_arb2_state_reg[2]/NET0131 ,
		_w3186_,
		_w4223_,
		_w7187_
	);
	LUT4 #(
		.INIT('h000e)
	) name5287 (
		_w3183_,
		_w3184_,
		_w3189_,
		_w3191_,
		_w7188_
	);
	LUT3 #(
		.INIT('h02)
	) name5288 (
		\s11_msel_arb2_state_reg[1]/NET0131 ,
		_w3194_,
		_w3198_,
		_w7189_
	);
	LUT3 #(
		.INIT('h45)
	) name5289 (
		_w7187_,
		_w7188_,
		_w7189_,
		_w7190_
	);
	LUT2 #(
		.INIT('h2)
	) name5290 (
		_w7186_,
		_w7190_,
		_w7191_
	);
	LUT4 #(
		.INIT('h000e)
	) name5291 (
		_w3189_,
		_w3191_,
		_w3194_,
		_w3198_,
		_w7192_
	);
	LUT2 #(
		.INIT('h2)
	) name5292 (
		_w3187_,
		_w7192_,
		_w7193_
	);
	LUT2 #(
		.INIT('h4)
	) name5293 (
		_w3183_,
		_w4233_,
		_w7194_
	);
	LUT3 #(
		.INIT('h54)
	) name5294 (
		\s11_msel_arb2_state_reg[2]/NET0131 ,
		_w3194_,
		_w3198_,
		_w7195_
	);
	LUT2 #(
		.INIT('h1)
	) name5295 (
		\s11_msel_arb2_state_reg[0]/NET0131 ,
		\s11_msel_arb2_state_reg[1]/NET0131 ,
		_w7196_
	);
	LUT3 #(
		.INIT('h10)
	) name5296 (
		_w3183_,
		_w3184_,
		_w7196_,
		_w7197_
	);
	LUT3 #(
		.INIT('h45)
	) name5297 (
		_w7194_,
		_w7195_,
		_w7197_,
		_w7198_
	);
	LUT3 #(
		.INIT('h54)
	) name5298 (
		\s11_msel_arb2_state_reg[1]/NET0131 ,
		_w3194_,
		_w3198_,
		_w7199_
	);
	LUT3 #(
		.INIT('h54)
	) name5299 (
		\s11_msel_arb2_state_reg[0]/NET0131 ,
		_w3189_,
		_w3191_,
		_w7200_
	);
	LUT3 #(
		.INIT('h10)
	) name5300 (
		\s11_msel_arb2_state_reg[2]/NET0131 ,
		_w7199_,
		_w7200_,
		_w7201_
	);
	LUT4 #(
		.INIT('h1110)
	) name5301 (
		_w3183_,
		_w3184_,
		_w3185_,
		_w3186_,
		_w7202_
	);
	LUT3 #(
		.INIT('h10)
	) name5302 (
		\s11_msel_arb2_state_reg[2]/NET0131 ,
		_w3194_,
		_w4232_,
		_w7203_
	);
	LUT3 #(
		.INIT('hd0)
	) name5303 (
		_w3197_,
		_w7202_,
		_w7203_,
		_w7204_
	);
	LUT4 #(
		.INIT('h000e)
	) name5304 (
		_w7193_,
		_w7198_,
		_w7201_,
		_w7204_,
		_w7205_
	);
	LUT2 #(
		.INIT('hb)
	) name5305 (
		_w7191_,
		_w7205_,
		_w7206_
	);
	LUT4 #(
		.INIT('h1110)
	) name5306 (
		_w3206_,
		_w3207_,
		_w3208_,
		_w3209_,
		_w7207_
	);
	LUT3 #(
		.INIT('h54)
	) name5307 (
		\s11_msel_arb3_state_reg[2]/NET0131 ,
		_w3206_,
		_w3219_,
		_w7208_
	);
	LUT4 #(
		.INIT('hafae)
	) name5308 (
		_w3211_,
		_w3214_,
		_w7207_,
		_w7208_,
		_w7209_
	);
	LUT3 #(
		.INIT('he0)
	) name5309 (
		_w3208_,
		_w3209_,
		_w3222_,
		_w7210_
	);
	LUT3 #(
		.INIT('h51)
	) name5310 (
		\s11_msel_arb3_state_reg[1]/NET0131 ,
		_w7209_,
		_w7210_,
		_w7211_
	);
	LUT4 #(
		.INIT('h00a8)
	) name5311 (
		\s11_msel_arb3_state_reg[2]/NET0131 ,
		_w3206_,
		_w3207_,
		_w3212_,
		_w7212_
	);
	LUT3 #(
		.INIT('h0e)
	) name5312 (
		_w3206_,
		_w3207_,
		_w3213_,
		_w7213_
	);
	LUT3 #(
		.INIT('h54)
	) name5313 (
		_w3209_,
		_w3211_,
		_w3219_,
		_w7214_
	);
	LUT2 #(
		.INIT('h1)
	) name5314 (
		_w3208_,
		_w3212_,
		_w7215_
	);
	LUT4 #(
		.INIT('h0155)
	) name5315 (
		_w7212_,
		_w7213_,
		_w7214_,
		_w7215_,
		_w7216_
	);
	LUT4 #(
		.INIT('h007f)
	) name5316 (
		\m3_s11_cyc_o_reg/NET0131 ,
		\rf_conf11_reg[6]/NET0131 ,
		\rf_conf11_reg[7]/NET0131 ,
		\s11_msel_arb3_state_reg[2]/NET0131 ,
		_w7217_
	);
	LUT4 #(
		.INIT('h02aa)
	) name5317 (
		\s11_msel_arb3_state_reg[1]/NET0131 ,
		_w3211_,
		_w3219_,
		_w7217_,
		_w7218_
	);
	LUT2 #(
		.INIT('h8)
	) name5318 (
		_w7216_,
		_w7218_,
		_w7219_
	);
	LUT3 #(
		.INIT('h54)
	) name5319 (
		\s11_msel_arb3_state_reg[1]/NET0131 ,
		_w3211_,
		_w3219_,
		_w7220_
	);
	LUT4 #(
		.INIT('h000e)
	) name5320 (
		_w3206_,
		_w3207_,
		_w3212_,
		_w3213_,
		_w7221_
	);
	LUT4 #(
		.INIT('h1115)
	) name5321 (
		\s11_msel_arb3_state_reg[0]/NET0131 ,
		\s11_msel_arb3_state_reg[2]/NET0131 ,
		_w7220_,
		_w7221_,
		_w7222_
	);
	LUT4 #(
		.INIT('h1110)
	) name5322 (
		_w3208_,
		_w3209_,
		_w3211_,
		_w3219_,
		_w7223_
	);
	LUT3 #(
		.INIT('h54)
	) name5323 (
		\s11_msel_arb3_state_reg[2]/NET0131 ,
		_w3228_,
		_w7223_,
		_w7224_
	);
	LUT3 #(
		.INIT('h02)
	) name5324 (
		\s11_msel_arb3_state_reg[1]/NET0131 ,
		_w3206_,
		_w3207_,
		_w7225_
	);
	LUT4 #(
		.INIT('h0001)
	) name5325 (
		_w3208_,
		_w3209_,
		_w3212_,
		_w3213_,
		_w7226_
	);
	LUT3 #(
		.INIT('h70)
	) name5326 (
		_w3220_,
		_w7225_,
		_w7226_,
		_w7227_
	);
	LUT3 #(
		.INIT('h02)
	) name5327 (
		_w7222_,
		_w7224_,
		_w7227_,
		_w7228_
	);
	LUT4 #(
		.INIT('hffa8)
	) name5328 (
		\s11_msel_arb3_state_reg[0]/NET0131 ,
		_w7211_,
		_w7219_,
		_w7228_,
		_w7229_
	);
	LUT3 #(
		.INIT('h54)
	) name5329 (
		\s12_msel_arb2_state_reg[2]/NET0131 ,
		_w4364_,
		_w4365_,
		_w7230_
	);
	LUT4 #(
		.INIT('h1110)
	) name5330 (
		_w4369_,
		_w4370_,
		_w4372_,
		_w4373_,
		_w7231_
	);
	LUT4 #(
		.INIT('h0d0c)
	) name5331 (
		\s12_msel_arb2_state_reg[0]/NET0131 ,
		_w6692_,
		_w7230_,
		_w7231_,
		_w7232_
	);
	LUT3 #(
		.INIT('h01)
	) name5332 (
		\s12_msel_arb2_state_reg[1]/NET0131 ,
		_w4369_,
		_w4370_,
		_w7233_
	);
	LUT2 #(
		.INIT('h8)
	) name5333 (
		_w6688_,
		_w7233_,
		_w7234_
	);
	LUT3 #(
		.INIT('ha8)
	) name5334 (
		\s12_msel_arb2_state_reg[2]/NET0131 ,
		_w4369_,
		_w4370_,
		_w7235_
	);
	LUT4 #(
		.INIT('h1110)
	) name5335 (
		_w4364_,
		_w4365_,
		_w4368_,
		_w4376_,
		_w7236_
	);
	LUT4 #(
		.INIT('h0d0c)
	) name5336 (
		\s12_msel_arb2_state_reg[0]/NET0131 ,
		_w6694_,
		_w7235_,
		_w7236_,
		_w7237_
	);
	LUT2 #(
		.INIT('h8)
	) name5337 (
		_w4369_,
		_w4385_,
		_w7238_
	);
	LUT3 #(
		.INIT('h10)
	) name5338 (
		_w4372_,
		_w4373_,
		_w4385_,
		_w7239_
	);
	LUT4 #(
		.INIT('h080a)
	) name5339 (
		\s12_msel_arb2_state_reg[0]/NET0131 ,
		_w7236_,
		_w7238_,
		_w7239_,
		_w7240_
	);
	LUT4 #(
		.INIT('h0001)
	) name5340 (
		_w7232_,
		_w7234_,
		_w7237_,
		_w7240_,
		_w7241_
	);
	LUT4 #(
		.INIT('h5400)
	) name5341 (
		_w4368_,
		_w4369_,
		_w4370_,
		_w4399_,
		_w7242_
	);
	LUT4 #(
		.INIT('hdf00)
	) name5342 (
		\m4_s12_cyc_o_reg/NET0131 ,
		\rf_conf12_reg[8]/NET0131 ,
		\rf_conf12_reg[9]/NET0131 ,
		\s12_msel_arb2_state_reg[1]/NET0131 ,
		_w7243_
	);
	LUT3 #(
		.INIT('h01)
	) name5343 (
		_w4364_,
		_w4365_,
		_w7243_,
		_w7244_
	);
	LUT4 #(
		.INIT('h0100)
	) name5344 (
		_w4368_,
		_w4372_,
		_w4373_,
		_w4399_,
		_w7245_
	);
	LUT3 #(
		.INIT('h45)
	) name5345 (
		_w7242_,
		_w7244_,
		_w7245_,
		_w7246_
	);
	LUT4 #(
		.INIT('h2000)
	) name5346 (
		\m3_s12_cyc_o_reg/NET0131 ,
		\rf_conf12_reg[6]/NET0131 ,
		\rf_conf12_reg[7]/NET0131 ,
		\s12_msel_arb2_state_reg[1]/NET0131 ,
		_w7247_
	);
	LUT3 #(
		.INIT('h02)
	) name5347 (
		\s12_msel_arb2_state_reg[1]/NET0131 ,
		_w4368_,
		_w4376_,
		_w7248_
	);
	LUT3 #(
		.INIT('h23)
	) name5348 (
		_w7231_,
		_w7247_,
		_w7248_,
		_w7249_
	);
	LUT4 #(
		.INIT('h0054)
	) name5349 (
		_w4368_,
		_w4369_,
		_w4370_,
		_w4376_,
		_w7250_
	);
	LUT4 #(
		.INIT('h00df)
	) name5350 (
		\m1_s12_cyc_o_reg/NET0131 ,
		\rf_conf12_reg[2]/NET0131 ,
		\rf_conf12_reg[3]/NET0131 ,
		\s12_msel_arb2_state_reg[1]/NET0131 ,
		_w7251_
	);
	LUT3 #(
		.INIT('hd0)
	) name5351 (
		_w6688_,
		_w7250_,
		_w7251_,
		_w7252_
	);
	LUT2 #(
		.INIT('h2)
	) name5352 (
		\s12_msel_arb2_state_reg[0]/NET0131 ,
		\s12_msel_arb2_state_reg[2]/NET0131 ,
		_w7253_
	);
	LUT4 #(
		.INIT('h08aa)
	) name5353 (
		_w7246_,
		_w7249_,
		_w7252_,
		_w7253_,
		_w7254_
	);
	LUT2 #(
		.INIT('hb)
	) name5354 (
		_w7241_,
		_w7254_,
		_w7255_
	);
	LUT4 #(
		.INIT('h4447)
	) name5355 (
		\s12_msel_arb3_state_reg[0]/NET0131 ,
		\s12_msel_arb3_state_reg[2]/NET0131 ,
		_w3249_,
		_w4433_,
		_w7256_
	);
	LUT4 #(
		.INIT('h1110)
	) name5356 (
		_w3237_,
		_w3238_,
		_w3244_,
		_w3245_,
		_w7257_
	);
	LUT2 #(
		.INIT('h8)
	) name5357 (
		_w7256_,
		_w7257_,
		_w7258_
	);
	LUT4 #(
		.INIT('hccc8)
	) name5358 (
		\s12_msel_arb3_state_reg[0]/NET0131 ,
		\s12_msel_arb3_state_reg[2]/NET0131 ,
		_w3237_,
		_w3238_,
		_w7259_
	);
	LUT4 #(
		.INIT('h000e)
	) name5359 (
		_w3247_,
		_w3248_,
		_w3249_,
		_w4433_,
		_w7260_
	);
	LUT2 #(
		.INIT('h4)
	) name5360 (
		_w7259_,
		_w7260_,
		_w7261_
	);
	LUT2 #(
		.INIT('h4)
	) name5361 (
		_w3237_,
		_w3240_,
		_w7262_
	);
	LUT4 #(
		.INIT('h000e)
	) name5362 (
		_w3247_,
		_w3248_,
		_w3249_,
		_w3250_,
		_w7263_
	);
	LUT3 #(
		.INIT('hc4)
	) name5363 (
		_w3246_,
		_w7262_,
		_w7263_,
		_w7264_
	);
	LUT4 #(
		.INIT('h5554)
	) name5364 (
		\s12_msel_arb3_state_reg[1]/NET0131 ,
		_w7258_,
		_w7261_,
		_w7264_,
		_w7265_
	);
	LUT3 #(
		.INIT('ha8)
	) name5365 (
		\s12_msel_arb3_state_reg[2]/NET0131 ,
		_w3249_,
		_w3250_,
		_w7266_
	);
	LUT4 #(
		.INIT('h000e)
	) name5366 (
		_w3237_,
		_w3238_,
		_w3247_,
		_w3248_,
		_w7267_
	);
	LUT3 #(
		.INIT('h54)
	) name5367 (
		_w4455_,
		_w7266_,
		_w7267_,
		_w7268_
	);
	LUT3 #(
		.INIT('h0e)
	) name5368 (
		_w3249_,
		_w3250_,
		_w3255_,
		_w7269_
	);
	LUT2 #(
		.INIT('h4)
	) name5369 (
		_w3248_,
		_w4442_,
		_w7270_
	);
	LUT2 #(
		.INIT('h1)
	) name5370 (
		_w3245_,
		_w3247_,
		_w7271_
	);
	LUT3 #(
		.INIT('he0)
	) name5371 (
		_w7269_,
		_w7270_,
		_w7271_,
		_w7272_
	);
	LUT3 #(
		.INIT('h0e)
	) name5372 (
		_w3237_,
		_w3238_,
		_w3247_,
		_w7273_
	);
	LUT3 #(
		.INIT('h2a)
	) name5373 (
		\s12_msel_arb3_state_reg[1]/NET0131 ,
		_w3256_,
		_w7273_,
		_w7274_
	);
	LUT4 #(
		.INIT('hab00)
	) name5374 (
		_w3244_,
		_w7268_,
		_w7272_,
		_w7274_,
		_w7275_
	);
	LUT2 #(
		.INIT('he)
	) name5375 (
		_w7265_,
		_w7275_,
		_w7276_
	);
	LUT4 #(
		.INIT('h0302)
	) name5376 (
		_w4551_,
		_w4555_,
		_w4556_,
		_w4559_,
		_w7277_
	);
	LUT4 #(
		.INIT('h888c)
	) name5377 (
		\s13_msel_arb2_state_reg[1]/NET0131 ,
		\s13_msel_arb2_state_reg[2]/NET0131 ,
		_w4551_,
		_w4559_,
		_w7278_
	);
	LUT4 #(
		.INIT('h0051)
	) name5378 (
		\s13_msel_arb2_state_reg[0]/NET0131 ,
		\s13_msel_arb2_state_reg[1]/NET0131 ,
		_w7277_,
		_w7278_,
		_w7279_
	);
	LUT3 #(
		.INIT('h02)
	) name5379 (
		\s13_msel_arb2_state_reg[1]/NET0131 ,
		_w4551_,
		_w4559_,
		_w7280_
	);
	LUT3 #(
		.INIT('ha2)
	) name5380 (
		_w6698_,
		_w6699_,
		_w7280_,
		_w7281_
	);
	LUT3 #(
		.INIT('h54)
	) name5381 (
		\s13_msel_arb2_state_reg[2]/NET0131 ,
		_w4555_,
		_w4556_,
		_w7282_
	);
	LUT3 #(
		.INIT('h04)
	) name5382 (
		\s13_msel_arb2_state_reg[0]/NET0131 ,
		_w6707_,
		_w7282_,
		_w7283_
	);
	LUT3 #(
		.INIT('h45)
	) name5383 (
		_w7279_,
		_w7281_,
		_w7283_,
		_w7284_
	);
	LUT3 #(
		.INIT('h54)
	) name5384 (
		\s13_msel_arb2_state_reg[2]/NET0131 ,
		_w4555_,
		_w4560_,
		_w7285_
	);
	LUT4 #(
		.INIT('hafae)
	) name5385 (
		_w4552_,
		_w6698_,
		_w7277_,
		_w7285_,
		_w7286_
	);
	LUT4 #(
		.INIT('h02aa)
	) name5386 (
		\s13_msel_arb2_state_reg[1]/NET0131 ,
		_w4551_,
		_w4559_,
		_w6705_,
		_w7287_
	);
	LUT3 #(
		.INIT('h8a)
	) name5387 (
		\s13_msel_arb2_state_reg[0]/NET0131 ,
		_w4559_,
		_w4568_,
		_w7288_
	);
	LUT4 #(
		.INIT('h0054)
	) name5388 (
		_w4553_,
		_w4555_,
		_w4556_,
		_w4557_,
		_w7289_
	);
	LUT3 #(
		.INIT('h02)
	) name5389 (
		\s13_msel_arb2_state_reg[0]/NET0131 ,
		_w4552_,
		_w4560_,
		_w7290_
	);
	LUT3 #(
		.INIT('h45)
	) name5390 (
		_w7288_,
		_w7289_,
		_w7290_,
		_w7291_
	);
	LUT3 #(
		.INIT('h07)
	) name5391 (
		_w7286_,
		_w7287_,
		_w7291_,
		_w7292_
	);
	LUT4 #(
		.INIT('h0504)
	) name5392 (
		_w4551_,
		_w4552_,
		_w4559_,
		_w4560_,
		_w7293_
	);
	LUT4 #(
		.INIT('h0020)
	) name5393 (
		\m0_s13_cyc_o_reg/NET0131 ,
		\rf_conf13_reg[0]/NET0131 ,
		\rf_conf13_reg[1]/NET0131 ,
		\s13_msel_arb2_state_reg[0]/NET0131 ,
		_w7294_
	);
	LUT3 #(
		.INIT('h04)
	) name5394 (
		_w4557_,
		_w4577_,
		_w7294_,
		_w7295_
	);
	LUT3 #(
		.INIT('hd0)
	) name5395 (
		_w6699_,
		_w7293_,
		_w7295_,
		_w7296_
	);
	LUT3 #(
		.INIT('hf2)
	) name5396 (
		_w7284_,
		_w7292_,
		_w7296_,
		_w7297_
	);
	LUT4 #(
		.INIT('h4447)
	) name5397 (
		\s13_msel_arb3_state_reg[0]/NET0131 ,
		\s13_msel_arb3_state_reg[2]/NET0131 ,
		_w2955_,
		_w4614_,
		_w7298_
	);
	LUT4 #(
		.INIT('h1110)
	) name5398 (
		_w2943_,
		_w2944_,
		_w2950_,
		_w2951_,
		_w7299_
	);
	LUT2 #(
		.INIT('h8)
	) name5399 (
		_w7298_,
		_w7299_,
		_w7300_
	);
	LUT4 #(
		.INIT('hccc8)
	) name5400 (
		\s13_msel_arb3_state_reg[0]/NET0131 ,
		\s13_msel_arb3_state_reg[2]/NET0131 ,
		_w2943_,
		_w2944_,
		_w7301_
	);
	LUT4 #(
		.INIT('h000e)
	) name5401 (
		_w2953_,
		_w2954_,
		_w2955_,
		_w4614_,
		_w7302_
	);
	LUT2 #(
		.INIT('h4)
	) name5402 (
		_w7301_,
		_w7302_,
		_w7303_
	);
	LUT2 #(
		.INIT('h4)
	) name5403 (
		_w2943_,
		_w2946_,
		_w7304_
	);
	LUT4 #(
		.INIT('h000e)
	) name5404 (
		_w2953_,
		_w2954_,
		_w2955_,
		_w2956_,
		_w7305_
	);
	LUT3 #(
		.INIT('hc4)
	) name5405 (
		_w2952_,
		_w7304_,
		_w7305_,
		_w7306_
	);
	LUT4 #(
		.INIT('h5554)
	) name5406 (
		\s13_msel_arb3_state_reg[1]/NET0131 ,
		_w7300_,
		_w7303_,
		_w7306_,
		_w7307_
	);
	LUT3 #(
		.INIT('ha8)
	) name5407 (
		\s13_msel_arb3_state_reg[2]/NET0131 ,
		_w2955_,
		_w2956_,
		_w7308_
	);
	LUT4 #(
		.INIT('h000e)
	) name5408 (
		_w2943_,
		_w2944_,
		_w2953_,
		_w2954_,
		_w7309_
	);
	LUT3 #(
		.INIT('h54)
	) name5409 (
		_w4636_,
		_w7308_,
		_w7309_,
		_w7310_
	);
	LUT3 #(
		.INIT('h0e)
	) name5410 (
		_w2955_,
		_w2956_,
		_w2961_,
		_w7311_
	);
	LUT2 #(
		.INIT('h4)
	) name5411 (
		_w2954_,
		_w4623_,
		_w7312_
	);
	LUT2 #(
		.INIT('h1)
	) name5412 (
		_w2951_,
		_w2953_,
		_w7313_
	);
	LUT3 #(
		.INIT('he0)
	) name5413 (
		_w7311_,
		_w7312_,
		_w7313_,
		_w7314_
	);
	LUT3 #(
		.INIT('h0e)
	) name5414 (
		_w2943_,
		_w2944_,
		_w2953_,
		_w7315_
	);
	LUT3 #(
		.INIT('h2a)
	) name5415 (
		\s13_msel_arb3_state_reg[1]/NET0131 ,
		_w2962_,
		_w7315_,
		_w7316_
	);
	LUT4 #(
		.INIT('hab00)
	) name5416 (
		_w2950_,
		_w7310_,
		_w7314_,
		_w7316_,
		_w7317_
	);
	LUT2 #(
		.INIT('he)
	) name5417 (
		_w7307_,
		_w7317_,
		_w7318_
	);
	LUT4 #(
		.INIT('h4447)
	) name5418 (
		\s14_msel_arb2_state_reg[0]/NET0131 ,
		\s14_msel_arb2_state_reg[2]/NET0131 ,
		_w2985_,
		_w4741_,
		_w7319_
	);
	LUT4 #(
		.INIT('h1110)
	) name5419 (
		_w2973_,
		_w2974_,
		_w2980_,
		_w2981_,
		_w7320_
	);
	LUT2 #(
		.INIT('h8)
	) name5420 (
		_w7319_,
		_w7320_,
		_w7321_
	);
	LUT4 #(
		.INIT('hccc8)
	) name5421 (
		\s14_msel_arb2_state_reg[0]/NET0131 ,
		\s14_msel_arb2_state_reg[2]/NET0131 ,
		_w2973_,
		_w2974_,
		_w7322_
	);
	LUT4 #(
		.INIT('h000e)
	) name5422 (
		_w2983_,
		_w2984_,
		_w2985_,
		_w4741_,
		_w7323_
	);
	LUT2 #(
		.INIT('h4)
	) name5423 (
		_w7322_,
		_w7323_,
		_w7324_
	);
	LUT2 #(
		.INIT('h4)
	) name5424 (
		_w2973_,
		_w2976_,
		_w7325_
	);
	LUT4 #(
		.INIT('h000e)
	) name5425 (
		_w2983_,
		_w2984_,
		_w2985_,
		_w2986_,
		_w7326_
	);
	LUT3 #(
		.INIT('hc4)
	) name5426 (
		_w2982_,
		_w7325_,
		_w7326_,
		_w7327_
	);
	LUT4 #(
		.INIT('h5554)
	) name5427 (
		\s14_msel_arb2_state_reg[1]/NET0131 ,
		_w7321_,
		_w7324_,
		_w7327_,
		_w7328_
	);
	LUT3 #(
		.INIT('ha8)
	) name5428 (
		\s14_msel_arb2_state_reg[2]/NET0131 ,
		_w2985_,
		_w2986_,
		_w7329_
	);
	LUT4 #(
		.INIT('h000e)
	) name5429 (
		_w2973_,
		_w2974_,
		_w2983_,
		_w2984_,
		_w7330_
	);
	LUT3 #(
		.INIT('h54)
	) name5430 (
		_w4763_,
		_w7329_,
		_w7330_,
		_w7331_
	);
	LUT3 #(
		.INIT('h0e)
	) name5431 (
		_w2985_,
		_w2986_,
		_w2991_,
		_w7332_
	);
	LUT2 #(
		.INIT('h4)
	) name5432 (
		_w2984_,
		_w4750_,
		_w7333_
	);
	LUT2 #(
		.INIT('h1)
	) name5433 (
		_w2981_,
		_w2983_,
		_w7334_
	);
	LUT3 #(
		.INIT('he0)
	) name5434 (
		_w7332_,
		_w7333_,
		_w7334_,
		_w7335_
	);
	LUT3 #(
		.INIT('h0e)
	) name5435 (
		_w2973_,
		_w2974_,
		_w2983_,
		_w7336_
	);
	LUT3 #(
		.INIT('h2a)
	) name5436 (
		\s14_msel_arb2_state_reg[1]/NET0131 ,
		_w2992_,
		_w7336_,
		_w7337_
	);
	LUT4 #(
		.INIT('hab00)
	) name5437 (
		_w2980_,
		_w7331_,
		_w7335_,
		_w7337_,
		_w7338_
	);
	LUT2 #(
		.INIT('he)
	) name5438 (
		_w7328_,
		_w7338_,
		_w7339_
	);
	LUT4 #(
		.INIT('h1110)
	) name5439 (
		_w3268_,
		_w3269_,
		_w3270_,
		_w3271_,
		_w7340_
	);
	LUT3 #(
		.INIT('h54)
	) name5440 (
		\s14_msel_arb3_state_reg[2]/NET0131 ,
		_w3268_,
		_w3281_,
		_w7341_
	);
	LUT4 #(
		.INIT('hafae)
	) name5441 (
		_w3273_,
		_w3276_,
		_w7340_,
		_w7341_,
		_w7342_
	);
	LUT3 #(
		.INIT('he0)
	) name5442 (
		_w3270_,
		_w3271_,
		_w3284_,
		_w7343_
	);
	LUT3 #(
		.INIT('h51)
	) name5443 (
		\s14_msel_arb3_state_reg[1]/NET0131 ,
		_w7342_,
		_w7343_,
		_w7344_
	);
	LUT4 #(
		.INIT('h00a8)
	) name5444 (
		\s14_msel_arb3_state_reg[2]/NET0131 ,
		_w3268_,
		_w3269_,
		_w3274_,
		_w7345_
	);
	LUT3 #(
		.INIT('h0e)
	) name5445 (
		_w3268_,
		_w3269_,
		_w3275_,
		_w7346_
	);
	LUT3 #(
		.INIT('h54)
	) name5446 (
		_w3271_,
		_w3273_,
		_w3281_,
		_w7347_
	);
	LUT2 #(
		.INIT('h1)
	) name5447 (
		_w3270_,
		_w3274_,
		_w7348_
	);
	LUT4 #(
		.INIT('h0155)
	) name5448 (
		_w7345_,
		_w7346_,
		_w7347_,
		_w7348_,
		_w7349_
	);
	LUT4 #(
		.INIT('h007f)
	) name5449 (
		\m3_s14_cyc_o_reg/NET0131 ,
		\rf_conf14_reg[6]/NET0131 ,
		\rf_conf14_reg[7]/NET0131 ,
		\s14_msel_arb3_state_reg[2]/NET0131 ,
		_w7350_
	);
	LUT4 #(
		.INIT('h02aa)
	) name5450 (
		\s14_msel_arb3_state_reg[1]/NET0131 ,
		_w3273_,
		_w3281_,
		_w7350_,
		_w7351_
	);
	LUT2 #(
		.INIT('h8)
	) name5451 (
		_w7349_,
		_w7351_,
		_w7352_
	);
	LUT3 #(
		.INIT('h54)
	) name5452 (
		\s14_msel_arb3_state_reg[1]/NET0131 ,
		_w3273_,
		_w3281_,
		_w7353_
	);
	LUT4 #(
		.INIT('h000e)
	) name5453 (
		_w3268_,
		_w3269_,
		_w3274_,
		_w3275_,
		_w7354_
	);
	LUT4 #(
		.INIT('h1115)
	) name5454 (
		\s14_msel_arb3_state_reg[0]/NET0131 ,
		\s14_msel_arb3_state_reg[2]/NET0131 ,
		_w7353_,
		_w7354_,
		_w7355_
	);
	LUT4 #(
		.INIT('h1110)
	) name5455 (
		_w3270_,
		_w3271_,
		_w3273_,
		_w3281_,
		_w7356_
	);
	LUT3 #(
		.INIT('h54)
	) name5456 (
		\s14_msel_arb3_state_reg[2]/NET0131 ,
		_w3290_,
		_w7356_,
		_w7357_
	);
	LUT3 #(
		.INIT('h02)
	) name5457 (
		\s14_msel_arb3_state_reg[1]/NET0131 ,
		_w3268_,
		_w3269_,
		_w7358_
	);
	LUT4 #(
		.INIT('h0001)
	) name5458 (
		_w3270_,
		_w3271_,
		_w3274_,
		_w3275_,
		_w7359_
	);
	LUT3 #(
		.INIT('h70)
	) name5459 (
		_w3282_,
		_w7358_,
		_w7359_,
		_w7360_
	);
	LUT3 #(
		.INIT('h02)
	) name5460 (
		_w7355_,
		_w7357_,
		_w7360_,
		_w7361_
	);
	LUT4 #(
		.INIT('hffa8)
	) name5461 (
		\s14_msel_arb3_state_reg[0]/NET0131 ,
		_w7344_,
		_w7352_,
		_w7361_,
		_w7362_
	);
	LUT4 #(
		.INIT('h0020)
	) name5462 (
		\m2_s1_cyc_o_reg/NET0131 ,
		\rf_conf1_reg[4]/NET0131 ,
		\rf_conf1_reg[5]/NET0131 ,
		\s1_msel_arb2_state_reg[0]/NET0131 ,
		_w7363_
	);
	LUT3 #(
		.INIT('h01)
	) name5463 (
		_w3299_,
		_w3300_,
		_w7363_,
		_w7364_
	);
	LUT4 #(
		.INIT('h2000)
	) name5464 (
		\m3_s1_cyc_o_reg/NET0131 ,
		\rf_conf1_reg[6]/NET0131 ,
		\rf_conf1_reg[7]/NET0131 ,
		\s1_msel_arb2_state_reg[0]/NET0131 ,
		_w7365_
	);
	LUT2 #(
		.INIT('h1)
	) name5465 (
		\s1_msel_arb2_state_reg[2]/NET0131 ,
		_w7365_,
		_w7366_
	);
	LUT4 #(
		.INIT('h00df)
	) name5466 (
		\m2_s1_cyc_o_reg/NET0131 ,
		\rf_conf1_reg[4]/NET0131 ,
		\rf_conf1_reg[5]/NET0131 ,
		\s1_msel_arb2_state_reg[1]/NET0131 ,
		_w7367_
	);
	LUT3 #(
		.INIT('h01)
	) name5467 (
		_w3310_,
		_w3314_,
		_w7367_,
		_w7368_
	);
	LUT4 #(
		.INIT('hcf4f)
	) name5468 (
		_w3303_,
		_w7364_,
		_w7366_,
		_w7368_,
		_w7369_
	);
	LUT4 #(
		.INIT('haaa2)
	) name5469 (
		\s1_msel_arb2_state_reg[1]/NET0131 ,
		\s1_msel_arb2_state_reg[2]/NET0131 ,
		_w3302_,
		_w5038_,
		_w7370_
	);
	LUT4 #(
		.INIT('h000e)
	) name5470 (
		_w3299_,
		_w3300_,
		_w3305_,
		_w3307_,
		_w7371_
	);
	LUT3 #(
		.INIT('h02)
	) name5471 (
		\s1_msel_arb2_state_reg[1]/NET0131 ,
		_w3310_,
		_w3314_,
		_w7372_
	);
	LUT3 #(
		.INIT('h45)
	) name5472 (
		_w7370_,
		_w7371_,
		_w7372_,
		_w7373_
	);
	LUT2 #(
		.INIT('h2)
	) name5473 (
		_w7369_,
		_w7373_,
		_w7374_
	);
	LUT4 #(
		.INIT('h000e)
	) name5474 (
		_w3305_,
		_w3307_,
		_w3310_,
		_w3314_,
		_w7375_
	);
	LUT2 #(
		.INIT('h2)
	) name5475 (
		_w3303_,
		_w7375_,
		_w7376_
	);
	LUT2 #(
		.INIT('h4)
	) name5476 (
		_w3299_,
		_w5048_,
		_w7377_
	);
	LUT3 #(
		.INIT('h54)
	) name5477 (
		\s1_msel_arb2_state_reg[2]/NET0131 ,
		_w3310_,
		_w3314_,
		_w7378_
	);
	LUT2 #(
		.INIT('h1)
	) name5478 (
		\s1_msel_arb2_state_reg[0]/NET0131 ,
		\s1_msel_arb2_state_reg[1]/NET0131 ,
		_w7379_
	);
	LUT3 #(
		.INIT('h10)
	) name5479 (
		_w3299_,
		_w3300_,
		_w7379_,
		_w7380_
	);
	LUT3 #(
		.INIT('h45)
	) name5480 (
		_w7377_,
		_w7378_,
		_w7380_,
		_w7381_
	);
	LUT3 #(
		.INIT('h54)
	) name5481 (
		\s1_msel_arb2_state_reg[1]/NET0131 ,
		_w3310_,
		_w3314_,
		_w7382_
	);
	LUT3 #(
		.INIT('h54)
	) name5482 (
		\s1_msel_arb2_state_reg[0]/NET0131 ,
		_w3305_,
		_w3307_,
		_w7383_
	);
	LUT3 #(
		.INIT('h10)
	) name5483 (
		\s1_msel_arb2_state_reg[2]/NET0131 ,
		_w7382_,
		_w7383_,
		_w7384_
	);
	LUT4 #(
		.INIT('h1110)
	) name5484 (
		_w3299_,
		_w3300_,
		_w3301_,
		_w3302_,
		_w7385_
	);
	LUT3 #(
		.INIT('h10)
	) name5485 (
		\s1_msel_arb2_state_reg[2]/NET0131 ,
		_w3310_,
		_w5047_,
		_w7386_
	);
	LUT3 #(
		.INIT('hd0)
	) name5486 (
		_w3313_,
		_w7385_,
		_w7386_,
		_w7387_
	);
	LUT4 #(
		.INIT('h000e)
	) name5487 (
		_w7376_,
		_w7381_,
		_w7384_,
		_w7387_,
		_w7388_
	);
	LUT2 #(
		.INIT('hb)
	) name5488 (
		_w7374_,
		_w7388_,
		_w7389_
	);
	LUT4 #(
		.INIT('h1110)
	) name5489 (
		_w3322_,
		_w3323_,
		_w3324_,
		_w3325_,
		_w7390_
	);
	LUT3 #(
		.INIT('h54)
	) name5490 (
		\s1_msel_arb3_state_reg[2]/NET0131 ,
		_w3322_,
		_w3335_,
		_w7391_
	);
	LUT4 #(
		.INIT('hafae)
	) name5491 (
		_w3327_,
		_w3330_,
		_w7390_,
		_w7391_,
		_w7392_
	);
	LUT3 #(
		.INIT('he0)
	) name5492 (
		_w3324_,
		_w3325_,
		_w3338_,
		_w7393_
	);
	LUT3 #(
		.INIT('h51)
	) name5493 (
		\s1_msel_arb3_state_reg[1]/NET0131 ,
		_w7392_,
		_w7393_,
		_w7394_
	);
	LUT4 #(
		.INIT('h00a8)
	) name5494 (
		\s1_msel_arb3_state_reg[2]/NET0131 ,
		_w3322_,
		_w3323_,
		_w3328_,
		_w7395_
	);
	LUT3 #(
		.INIT('h0e)
	) name5495 (
		_w3322_,
		_w3323_,
		_w3329_,
		_w7396_
	);
	LUT3 #(
		.INIT('h54)
	) name5496 (
		_w3325_,
		_w3327_,
		_w3335_,
		_w7397_
	);
	LUT2 #(
		.INIT('h1)
	) name5497 (
		_w3324_,
		_w3328_,
		_w7398_
	);
	LUT4 #(
		.INIT('h0155)
	) name5498 (
		_w7395_,
		_w7396_,
		_w7397_,
		_w7398_,
		_w7399_
	);
	LUT4 #(
		.INIT('h007f)
	) name5499 (
		\m3_s1_cyc_o_reg/NET0131 ,
		\rf_conf1_reg[6]/NET0131 ,
		\rf_conf1_reg[7]/NET0131 ,
		\s1_msel_arb3_state_reg[2]/NET0131 ,
		_w7400_
	);
	LUT4 #(
		.INIT('h02aa)
	) name5500 (
		\s1_msel_arb3_state_reg[1]/NET0131 ,
		_w3327_,
		_w3335_,
		_w7400_,
		_w7401_
	);
	LUT2 #(
		.INIT('h8)
	) name5501 (
		_w7399_,
		_w7401_,
		_w7402_
	);
	LUT3 #(
		.INIT('h54)
	) name5502 (
		\s1_msel_arb3_state_reg[1]/NET0131 ,
		_w3327_,
		_w3335_,
		_w7403_
	);
	LUT4 #(
		.INIT('h000e)
	) name5503 (
		_w3322_,
		_w3323_,
		_w3328_,
		_w3329_,
		_w7404_
	);
	LUT4 #(
		.INIT('h1115)
	) name5504 (
		\s1_msel_arb3_state_reg[0]/NET0131 ,
		\s1_msel_arb3_state_reg[2]/NET0131 ,
		_w7403_,
		_w7404_,
		_w7405_
	);
	LUT4 #(
		.INIT('h1110)
	) name5505 (
		_w3324_,
		_w3325_,
		_w3327_,
		_w3335_,
		_w7406_
	);
	LUT3 #(
		.INIT('h54)
	) name5506 (
		\s1_msel_arb3_state_reg[2]/NET0131 ,
		_w3344_,
		_w7406_,
		_w7407_
	);
	LUT3 #(
		.INIT('h02)
	) name5507 (
		\s1_msel_arb3_state_reg[1]/NET0131 ,
		_w3322_,
		_w3323_,
		_w7408_
	);
	LUT4 #(
		.INIT('h0001)
	) name5508 (
		_w3324_,
		_w3325_,
		_w3328_,
		_w3329_,
		_w7409_
	);
	LUT3 #(
		.INIT('h70)
	) name5509 (
		_w3336_,
		_w7408_,
		_w7409_,
		_w7410_
	);
	LUT3 #(
		.INIT('h02)
	) name5510 (
		_w7405_,
		_w7407_,
		_w7410_,
		_w7411_
	);
	LUT4 #(
		.INIT('hffa8)
	) name5511 (
		\s1_msel_arb3_state_reg[0]/NET0131 ,
		_w7394_,
		_w7402_,
		_w7411_,
		_w7412_
	);
	LUT4 #(
		.INIT('h0302)
	) name5512 (
		_w5184_,
		_w5188_,
		_w5189_,
		_w5192_,
		_w7413_
	);
	LUT4 #(
		.INIT('h888c)
	) name5513 (
		\s2_msel_arb2_state_reg[1]/NET0131 ,
		\s2_msel_arb2_state_reg[2]/NET0131 ,
		_w5184_,
		_w5192_,
		_w7414_
	);
	LUT4 #(
		.INIT('h0051)
	) name5514 (
		\s2_msel_arb2_state_reg[0]/NET0131 ,
		\s2_msel_arb2_state_reg[1]/NET0131 ,
		_w7413_,
		_w7414_,
		_w7415_
	);
	LUT3 #(
		.INIT('h02)
	) name5515 (
		\s2_msel_arb2_state_reg[1]/NET0131 ,
		_w5184_,
		_w5192_,
		_w7416_
	);
	LUT3 #(
		.INIT('ha2)
	) name5516 (
		_w6713_,
		_w6714_,
		_w7416_,
		_w7417_
	);
	LUT3 #(
		.INIT('h54)
	) name5517 (
		\s2_msel_arb2_state_reg[2]/NET0131 ,
		_w5188_,
		_w5189_,
		_w7418_
	);
	LUT3 #(
		.INIT('h04)
	) name5518 (
		\s2_msel_arb2_state_reg[0]/NET0131 ,
		_w6722_,
		_w7418_,
		_w7419_
	);
	LUT3 #(
		.INIT('h45)
	) name5519 (
		_w7415_,
		_w7417_,
		_w7419_,
		_w7420_
	);
	LUT3 #(
		.INIT('h54)
	) name5520 (
		\s2_msel_arb2_state_reg[2]/NET0131 ,
		_w5188_,
		_w5193_,
		_w7421_
	);
	LUT4 #(
		.INIT('hafae)
	) name5521 (
		_w5185_,
		_w6713_,
		_w7413_,
		_w7421_,
		_w7422_
	);
	LUT4 #(
		.INIT('h02aa)
	) name5522 (
		\s2_msel_arb2_state_reg[1]/NET0131 ,
		_w5184_,
		_w5192_,
		_w6720_,
		_w7423_
	);
	LUT3 #(
		.INIT('h8a)
	) name5523 (
		\s2_msel_arb2_state_reg[0]/NET0131 ,
		_w5192_,
		_w5201_,
		_w7424_
	);
	LUT4 #(
		.INIT('h0054)
	) name5524 (
		_w5186_,
		_w5188_,
		_w5189_,
		_w5190_,
		_w7425_
	);
	LUT3 #(
		.INIT('h02)
	) name5525 (
		\s2_msel_arb2_state_reg[0]/NET0131 ,
		_w5185_,
		_w5193_,
		_w7426_
	);
	LUT3 #(
		.INIT('h45)
	) name5526 (
		_w7424_,
		_w7425_,
		_w7426_,
		_w7427_
	);
	LUT3 #(
		.INIT('h07)
	) name5527 (
		_w7422_,
		_w7423_,
		_w7427_,
		_w7428_
	);
	LUT4 #(
		.INIT('h0504)
	) name5528 (
		_w5184_,
		_w5185_,
		_w5192_,
		_w5193_,
		_w7429_
	);
	LUT4 #(
		.INIT('h0020)
	) name5529 (
		\m0_s2_cyc_o_reg/NET0131 ,
		\rf_conf2_reg[0]/NET0131 ,
		\rf_conf2_reg[1]/NET0131 ,
		\s2_msel_arb2_state_reg[0]/NET0131 ,
		_w7430_
	);
	LUT3 #(
		.INIT('h04)
	) name5530 (
		_w5190_,
		_w5210_,
		_w7430_,
		_w7431_
	);
	LUT3 #(
		.INIT('hd0)
	) name5531 (
		_w6714_,
		_w7429_,
		_w7431_,
		_w7432_
	);
	LUT3 #(
		.INIT('hf2)
	) name5532 (
		_w7420_,
		_w7428_,
		_w7432_,
		_w7433_
	);
	LUT4 #(
		.INIT('h4447)
	) name5533 (
		\s2_msel_arb3_state_reg[0]/NET0131 ,
		\s2_msel_arb3_state_reg[2]/NET0131 ,
		_w3015_,
		_w5247_,
		_w7434_
	);
	LUT4 #(
		.INIT('h1110)
	) name5534 (
		_w3003_,
		_w3004_,
		_w3010_,
		_w3011_,
		_w7435_
	);
	LUT2 #(
		.INIT('h8)
	) name5535 (
		_w7434_,
		_w7435_,
		_w7436_
	);
	LUT4 #(
		.INIT('hccc8)
	) name5536 (
		\s2_msel_arb3_state_reg[0]/NET0131 ,
		\s2_msel_arb3_state_reg[2]/NET0131 ,
		_w3003_,
		_w3004_,
		_w7437_
	);
	LUT4 #(
		.INIT('h000e)
	) name5537 (
		_w3013_,
		_w3014_,
		_w3015_,
		_w5247_,
		_w7438_
	);
	LUT2 #(
		.INIT('h4)
	) name5538 (
		_w7437_,
		_w7438_,
		_w7439_
	);
	LUT2 #(
		.INIT('h4)
	) name5539 (
		_w3003_,
		_w3006_,
		_w7440_
	);
	LUT4 #(
		.INIT('h000e)
	) name5540 (
		_w3013_,
		_w3014_,
		_w3015_,
		_w3016_,
		_w7441_
	);
	LUT3 #(
		.INIT('hc4)
	) name5541 (
		_w3012_,
		_w7440_,
		_w7441_,
		_w7442_
	);
	LUT4 #(
		.INIT('h5554)
	) name5542 (
		\s2_msel_arb3_state_reg[1]/NET0131 ,
		_w7436_,
		_w7439_,
		_w7442_,
		_w7443_
	);
	LUT3 #(
		.INIT('ha8)
	) name5543 (
		\s2_msel_arb3_state_reg[2]/NET0131 ,
		_w3015_,
		_w3016_,
		_w7444_
	);
	LUT4 #(
		.INIT('h000e)
	) name5544 (
		_w3003_,
		_w3004_,
		_w3013_,
		_w3014_,
		_w7445_
	);
	LUT3 #(
		.INIT('h54)
	) name5545 (
		_w5269_,
		_w7444_,
		_w7445_,
		_w7446_
	);
	LUT3 #(
		.INIT('h0e)
	) name5546 (
		_w3015_,
		_w3016_,
		_w3021_,
		_w7447_
	);
	LUT2 #(
		.INIT('h4)
	) name5547 (
		_w3014_,
		_w5256_,
		_w7448_
	);
	LUT2 #(
		.INIT('h1)
	) name5548 (
		_w3011_,
		_w3013_,
		_w7449_
	);
	LUT3 #(
		.INIT('he0)
	) name5549 (
		_w7447_,
		_w7448_,
		_w7449_,
		_w7450_
	);
	LUT3 #(
		.INIT('h0e)
	) name5550 (
		_w3003_,
		_w3004_,
		_w3013_,
		_w7451_
	);
	LUT3 #(
		.INIT('h2a)
	) name5551 (
		\s2_msel_arb3_state_reg[1]/NET0131 ,
		_w3022_,
		_w7451_,
		_w7452_
	);
	LUT4 #(
		.INIT('hab00)
	) name5552 (
		_w3010_,
		_w7446_,
		_w7450_,
		_w7452_,
		_w7453_
	);
	LUT2 #(
		.INIT('he)
	) name5553 (
		_w7443_,
		_w7453_,
		_w7454_
	);
	LUT4 #(
		.INIT('h0020)
	) name5554 (
		\m2_s3_cyc_o_reg/NET0131 ,
		\rf_conf3_reg[4]/NET0131 ,
		\rf_conf3_reg[5]/NET0131 ,
		\s3_msel_arb2_state_reg[0]/NET0131 ,
		_w7455_
	);
	LUT3 #(
		.INIT('h01)
	) name5555 (
		_w3033_,
		_w3034_,
		_w7455_,
		_w7456_
	);
	LUT4 #(
		.INIT('h2000)
	) name5556 (
		\m3_s3_cyc_o_reg/NET0131 ,
		\rf_conf3_reg[6]/NET0131 ,
		\rf_conf3_reg[7]/NET0131 ,
		\s3_msel_arb2_state_reg[0]/NET0131 ,
		_w7457_
	);
	LUT2 #(
		.INIT('h1)
	) name5557 (
		\s3_msel_arb2_state_reg[2]/NET0131 ,
		_w7457_,
		_w7458_
	);
	LUT4 #(
		.INIT('h00df)
	) name5558 (
		\m2_s3_cyc_o_reg/NET0131 ,
		\rf_conf3_reg[4]/NET0131 ,
		\rf_conf3_reg[5]/NET0131 ,
		\s3_msel_arb2_state_reg[1]/NET0131 ,
		_w7459_
	);
	LUT3 #(
		.INIT('h01)
	) name5559 (
		_w3044_,
		_w3048_,
		_w7459_,
		_w7460_
	);
	LUT4 #(
		.INIT('hcf4f)
	) name5560 (
		_w3037_,
		_w7456_,
		_w7458_,
		_w7460_,
		_w7461_
	);
	LUT4 #(
		.INIT('haaa2)
	) name5561 (
		\s3_msel_arb2_state_reg[1]/NET0131 ,
		\s3_msel_arb2_state_reg[2]/NET0131 ,
		_w3036_,
		_w5385_,
		_w7462_
	);
	LUT4 #(
		.INIT('h000e)
	) name5562 (
		_w3033_,
		_w3034_,
		_w3039_,
		_w3041_,
		_w7463_
	);
	LUT3 #(
		.INIT('h02)
	) name5563 (
		\s3_msel_arb2_state_reg[1]/NET0131 ,
		_w3044_,
		_w3048_,
		_w7464_
	);
	LUT3 #(
		.INIT('h45)
	) name5564 (
		_w7462_,
		_w7463_,
		_w7464_,
		_w7465_
	);
	LUT2 #(
		.INIT('h2)
	) name5565 (
		_w7461_,
		_w7465_,
		_w7466_
	);
	LUT4 #(
		.INIT('h000e)
	) name5566 (
		_w3039_,
		_w3041_,
		_w3044_,
		_w3048_,
		_w7467_
	);
	LUT2 #(
		.INIT('h2)
	) name5567 (
		_w3037_,
		_w7467_,
		_w7468_
	);
	LUT2 #(
		.INIT('h4)
	) name5568 (
		_w3033_,
		_w5395_,
		_w7469_
	);
	LUT3 #(
		.INIT('h54)
	) name5569 (
		\s3_msel_arb2_state_reg[2]/NET0131 ,
		_w3044_,
		_w3048_,
		_w7470_
	);
	LUT2 #(
		.INIT('h1)
	) name5570 (
		\s3_msel_arb2_state_reg[0]/NET0131 ,
		\s3_msel_arb2_state_reg[1]/NET0131 ,
		_w7471_
	);
	LUT3 #(
		.INIT('h10)
	) name5571 (
		_w3033_,
		_w3034_,
		_w7471_,
		_w7472_
	);
	LUT3 #(
		.INIT('h45)
	) name5572 (
		_w7469_,
		_w7470_,
		_w7472_,
		_w7473_
	);
	LUT3 #(
		.INIT('h54)
	) name5573 (
		\s3_msel_arb2_state_reg[1]/NET0131 ,
		_w3044_,
		_w3048_,
		_w7474_
	);
	LUT3 #(
		.INIT('h54)
	) name5574 (
		\s3_msel_arb2_state_reg[0]/NET0131 ,
		_w3039_,
		_w3041_,
		_w7475_
	);
	LUT3 #(
		.INIT('h10)
	) name5575 (
		\s3_msel_arb2_state_reg[2]/NET0131 ,
		_w7474_,
		_w7475_,
		_w7476_
	);
	LUT4 #(
		.INIT('h1110)
	) name5576 (
		_w3033_,
		_w3034_,
		_w3035_,
		_w3036_,
		_w7477_
	);
	LUT3 #(
		.INIT('h10)
	) name5577 (
		\s3_msel_arb2_state_reg[2]/NET0131 ,
		_w3044_,
		_w5394_,
		_w7478_
	);
	LUT3 #(
		.INIT('hd0)
	) name5578 (
		_w3047_,
		_w7477_,
		_w7478_,
		_w7479_
	);
	LUT4 #(
		.INIT('h000e)
	) name5579 (
		_w7468_,
		_w7473_,
		_w7476_,
		_w7479_,
		_w7480_
	);
	LUT2 #(
		.INIT('hb)
	) name5580 (
		_w7466_,
		_w7480_,
		_w7481_
	);
	LUT4 #(
		.INIT('h1110)
	) name5581 (
		_w3354_,
		_w3355_,
		_w3356_,
		_w3357_,
		_w7482_
	);
	LUT3 #(
		.INIT('h54)
	) name5582 (
		\s3_msel_arb3_state_reg[2]/NET0131 ,
		_w3354_,
		_w3367_,
		_w7483_
	);
	LUT4 #(
		.INIT('hafae)
	) name5583 (
		_w3359_,
		_w3362_,
		_w7482_,
		_w7483_,
		_w7484_
	);
	LUT3 #(
		.INIT('he0)
	) name5584 (
		_w3356_,
		_w3357_,
		_w3370_,
		_w7485_
	);
	LUT3 #(
		.INIT('h51)
	) name5585 (
		\s3_msel_arb3_state_reg[1]/NET0131 ,
		_w7484_,
		_w7485_,
		_w7486_
	);
	LUT4 #(
		.INIT('h00a8)
	) name5586 (
		\s3_msel_arb3_state_reg[2]/NET0131 ,
		_w3354_,
		_w3355_,
		_w3360_,
		_w7487_
	);
	LUT3 #(
		.INIT('h0e)
	) name5587 (
		_w3354_,
		_w3355_,
		_w3361_,
		_w7488_
	);
	LUT3 #(
		.INIT('h54)
	) name5588 (
		_w3357_,
		_w3359_,
		_w3367_,
		_w7489_
	);
	LUT2 #(
		.INIT('h1)
	) name5589 (
		_w3356_,
		_w3360_,
		_w7490_
	);
	LUT4 #(
		.INIT('h0155)
	) name5590 (
		_w7487_,
		_w7488_,
		_w7489_,
		_w7490_,
		_w7491_
	);
	LUT4 #(
		.INIT('h007f)
	) name5591 (
		\m3_s3_cyc_o_reg/NET0131 ,
		\rf_conf3_reg[6]/NET0131 ,
		\rf_conf3_reg[7]/NET0131 ,
		\s3_msel_arb3_state_reg[2]/NET0131 ,
		_w7492_
	);
	LUT4 #(
		.INIT('h02aa)
	) name5592 (
		\s3_msel_arb3_state_reg[1]/NET0131 ,
		_w3359_,
		_w3367_,
		_w7492_,
		_w7493_
	);
	LUT2 #(
		.INIT('h8)
	) name5593 (
		_w7491_,
		_w7493_,
		_w7494_
	);
	LUT3 #(
		.INIT('h54)
	) name5594 (
		\s3_msel_arb3_state_reg[1]/NET0131 ,
		_w3359_,
		_w3367_,
		_w7495_
	);
	LUT4 #(
		.INIT('h000e)
	) name5595 (
		_w3354_,
		_w3355_,
		_w3360_,
		_w3361_,
		_w7496_
	);
	LUT4 #(
		.INIT('h1115)
	) name5596 (
		\s3_msel_arb3_state_reg[0]/NET0131 ,
		\s3_msel_arb3_state_reg[2]/NET0131 ,
		_w7495_,
		_w7496_,
		_w7497_
	);
	LUT4 #(
		.INIT('h1110)
	) name5597 (
		_w3356_,
		_w3357_,
		_w3359_,
		_w3367_,
		_w7498_
	);
	LUT3 #(
		.INIT('h54)
	) name5598 (
		\s3_msel_arb3_state_reg[2]/NET0131 ,
		_w3376_,
		_w7498_,
		_w7499_
	);
	LUT3 #(
		.INIT('h02)
	) name5599 (
		\s3_msel_arb3_state_reg[1]/NET0131 ,
		_w3354_,
		_w3355_,
		_w7500_
	);
	LUT4 #(
		.INIT('h0001)
	) name5600 (
		_w3356_,
		_w3357_,
		_w3360_,
		_w3361_,
		_w7501_
	);
	LUT3 #(
		.INIT('h70)
	) name5601 (
		_w3368_,
		_w7500_,
		_w7501_,
		_w7502_
	);
	LUT3 #(
		.INIT('h02)
	) name5602 (
		_w7497_,
		_w7499_,
		_w7502_,
		_w7503_
	);
	LUT4 #(
		.INIT('hffa8)
	) name5603 (
		\s3_msel_arb3_state_reg[0]/NET0131 ,
		_w7486_,
		_w7494_,
		_w7503_,
		_w7504_
	);
	LUT4 #(
		.INIT('h0302)
	) name5604 (
		_w5535_,
		_w5539_,
		_w5540_,
		_w5543_,
		_w7505_
	);
	LUT4 #(
		.INIT('h888c)
	) name5605 (
		\s4_msel_arb2_state_reg[1]/NET0131 ,
		\s4_msel_arb2_state_reg[2]/NET0131 ,
		_w5535_,
		_w5543_,
		_w7506_
	);
	LUT4 #(
		.INIT('h0051)
	) name5606 (
		\s4_msel_arb2_state_reg[0]/NET0131 ,
		\s4_msel_arb2_state_reg[1]/NET0131 ,
		_w7505_,
		_w7506_,
		_w7507_
	);
	LUT3 #(
		.INIT('h02)
	) name5607 (
		\s4_msel_arb2_state_reg[1]/NET0131 ,
		_w5535_,
		_w5543_,
		_w7508_
	);
	LUT3 #(
		.INIT('ha2)
	) name5608 (
		_w6728_,
		_w6729_,
		_w7508_,
		_w7509_
	);
	LUT3 #(
		.INIT('h54)
	) name5609 (
		\s4_msel_arb2_state_reg[2]/NET0131 ,
		_w5539_,
		_w5540_,
		_w7510_
	);
	LUT3 #(
		.INIT('h04)
	) name5610 (
		\s4_msel_arb2_state_reg[0]/NET0131 ,
		_w6737_,
		_w7510_,
		_w7511_
	);
	LUT3 #(
		.INIT('h45)
	) name5611 (
		_w7507_,
		_w7509_,
		_w7511_,
		_w7512_
	);
	LUT3 #(
		.INIT('h54)
	) name5612 (
		\s4_msel_arb2_state_reg[2]/NET0131 ,
		_w5539_,
		_w5544_,
		_w7513_
	);
	LUT4 #(
		.INIT('hafae)
	) name5613 (
		_w5536_,
		_w6728_,
		_w7505_,
		_w7513_,
		_w7514_
	);
	LUT4 #(
		.INIT('h02aa)
	) name5614 (
		\s4_msel_arb2_state_reg[1]/NET0131 ,
		_w5535_,
		_w5543_,
		_w6735_,
		_w7515_
	);
	LUT3 #(
		.INIT('h8a)
	) name5615 (
		\s4_msel_arb2_state_reg[0]/NET0131 ,
		_w5543_,
		_w5552_,
		_w7516_
	);
	LUT4 #(
		.INIT('h0054)
	) name5616 (
		_w5537_,
		_w5539_,
		_w5540_,
		_w5541_,
		_w7517_
	);
	LUT3 #(
		.INIT('h02)
	) name5617 (
		\s4_msel_arb2_state_reg[0]/NET0131 ,
		_w5536_,
		_w5544_,
		_w7518_
	);
	LUT3 #(
		.INIT('h45)
	) name5618 (
		_w7516_,
		_w7517_,
		_w7518_,
		_w7519_
	);
	LUT3 #(
		.INIT('h07)
	) name5619 (
		_w7514_,
		_w7515_,
		_w7519_,
		_w7520_
	);
	LUT4 #(
		.INIT('h0504)
	) name5620 (
		_w5535_,
		_w5536_,
		_w5543_,
		_w5544_,
		_w7521_
	);
	LUT4 #(
		.INIT('h0020)
	) name5621 (
		\m0_s4_cyc_o_reg/NET0131 ,
		\rf_conf4_reg[0]/NET0131 ,
		\rf_conf4_reg[1]/NET0131 ,
		\s4_msel_arb2_state_reg[0]/NET0131 ,
		_w7522_
	);
	LUT3 #(
		.INIT('h04)
	) name5622 (
		_w5541_,
		_w5561_,
		_w7522_,
		_w7523_
	);
	LUT3 #(
		.INIT('hd0)
	) name5623 (
		_w6729_,
		_w7521_,
		_w7523_,
		_w7524_
	);
	LUT3 #(
		.INIT('hf2)
	) name5624 (
		_w7512_,
		_w7520_,
		_w7524_,
		_w7525_
	);
	LUT4 #(
		.INIT('h1110)
	) name5625 (
		_w3056_,
		_w3057_,
		_w3058_,
		_w3059_,
		_w7526_
	);
	LUT3 #(
		.INIT('h54)
	) name5626 (
		\s4_msel_arb3_state_reg[2]/NET0131 ,
		_w3056_,
		_w3069_,
		_w7527_
	);
	LUT4 #(
		.INIT('hafae)
	) name5627 (
		_w3061_,
		_w3064_,
		_w7526_,
		_w7527_,
		_w7528_
	);
	LUT3 #(
		.INIT('he0)
	) name5628 (
		_w3058_,
		_w3059_,
		_w3072_,
		_w7529_
	);
	LUT3 #(
		.INIT('h51)
	) name5629 (
		\s4_msel_arb3_state_reg[1]/NET0131 ,
		_w7528_,
		_w7529_,
		_w7530_
	);
	LUT4 #(
		.INIT('h00a8)
	) name5630 (
		\s4_msel_arb3_state_reg[2]/NET0131 ,
		_w3056_,
		_w3057_,
		_w3062_,
		_w7531_
	);
	LUT3 #(
		.INIT('h0e)
	) name5631 (
		_w3056_,
		_w3057_,
		_w3063_,
		_w7532_
	);
	LUT3 #(
		.INIT('h54)
	) name5632 (
		_w3059_,
		_w3061_,
		_w3069_,
		_w7533_
	);
	LUT2 #(
		.INIT('h1)
	) name5633 (
		_w3058_,
		_w3062_,
		_w7534_
	);
	LUT4 #(
		.INIT('h0155)
	) name5634 (
		_w7531_,
		_w7532_,
		_w7533_,
		_w7534_,
		_w7535_
	);
	LUT4 #(
		.INIT('h007f)
	) name5635 (
		\m3_s4_cyc_o_reg/NET0131 ,
		\rf_conf4_reg[6]/NET0131 ,
		\rf_conf4_reg[7]/NET0131 ,
		\s4_msel_arb3_state_reg[2]/NET0131 ,
		_w7536_
	);
	LUT4 #(
		.INIT('h02aa)
	) name5636 (
		\s4_msel_arb3_state_reg[1]/NET0131 ,
		_w3061_,
		_w3069_,
		_w7536_,
		_w7537_
	);
	LUT2 #(
		.INIT('h8)
	) name5637 (
		_w7535_,
		_w7537_,
		_w7538_
	);
	LUT3 #(
		.INIT('h54)
	) name5638 (
		\s4_msel_arb3_state_reg[1]/NET0131 ,
		_w3061_,
		_w3069_,
		_w7539_
	);
	LUT4 #(
		.INIT('h000e)
	) name5639 (
		_w3056_,
		_w3057_,
		_w3062_,
		_w3063_,
		_w7540_
	);
	LUT4 #(
		.INIT('h1115)
	) name5640 (
		\s4_msel_arb3_state_reg[0]/NET0131 ,
		\s4_msel_arb3_state_reg[2]/NET0131 ,
		_w7539_,
		_w7540_,
		_w7541_
	);
	LUT4 #(
		.INIT('h1110)
	) name5641 (
		_w3058_,
		_w3059_,
		_w3061_,
		_w3069_,
		_w7542_
	);
	LUT3 #(
		.INIT('h54)
	) name5642 (
		\s4_msel_arb3_state_reg[2]/NET0131 ,
		_w3078_,
		_w7542_,
		_w7543_
	);
	LUT3 #(
		.INIT('h02)
	) name5643 (
		\s4_msel_arb3_state_reg[1]/NET0131 ,
		_w3056_,
		_w3057_,
		_w7544_
	);
	LUT4 #(
		.INIT('h0001)
	) name5644 (
		_w3058_,
		_w3059_,
		_w3062_,
		_w3063_,
		_w7545_
	);
	LUT3 #(
		.INIT('h70)
	) name5645 (
		_w3070_,
		_w7544_,
		_w7545_,
		_w7546_
	);
	LUT3 #(
		.INIT('h02)
	) name5646 (
		_w7541_,
		_w7543_,
		_w7546_,
		_w7547_
	);
	LUT4 #(
		.INIT('hffa8)
	) name5647 (
		\s4_msel_arb3_state_reg[0]/NET0131 ,
		_w7530_,
		_w7538_,
		_w7547_,
		_w7548_
	);
	LUT4 #(
		.INIT('h0020)
	) name5648 (
		\m2_s5_cyc_o_reg/NET0131 ,
		\rf_conf5_reg[4]/NET0131 ,
		\rf_conf5_reg[5]/NET0131 ,
		\s5_msel_arb2_state_reg[0]/NET0131 ,
		_w7549_
	);
	LUT3 #(
		.INIT('h01)
	) name5649 (
		_w3385_,
		_w3386_,
		_w7549_,
		_w7550_
	);
	LUT4 #(
		.INIT('h2000)
	) name5650 (
		\m3_s5_cyc_o_reg/NET0131 ,
		\rf_conf5_reg[6]/NET0131 ,
		\rf_conf5_reg[7]/NET0131 ,
		\s5_msel_arb2_state_reg[0]/NET0131 ,
		_w7551_
	);
	LUT2 #(
		.INIT('h1)
	) name5651 (
		\s5_msel_arb2_state_reg[2]/NET0131 ,
		_w7551_,
		_w7552_
	);
	LUT4 #(
		.INIT('h00df)
	) name5652 (
		\m2_s5_cyc_o_reg/NET0131 ,
		\rf_conf5_reg[4]/NET0131 ,
		\rf_conf5_reg[5]/NET0131 ,
		\s5_msel_arb2_state_reg[1]/NET0131 ,
		_w7553_
	);
	LUT3 #(
		.INIT('h01)
	) name5653 (
		_w3396_,
		_w3400_,
		_w7553_,
		_w7554_
	);
	LUT4 #(
		.INIT('hcf4f)
	) name5654 (
		_w3389_,
		_w7550_,
		_w7552_,
		_w7554_,
		_w7555_
	);
	LUT4 #(
		.INIT('haaa2)
	) name5655 (
		\s5_msel_arb2_state_reg[1]/NET0131 ,
		\s5_msel_arb2_state_reg[2]/NET0131 ,
		_w3388_,
		_w5725_,
		_w7556_
	);
	LUT4 #(
		.INIT('h000e)
	) name5656 (
		_w3385_,
		_w3386_,
		_w3391_,
		_w3393_,
		_w7557_
	);
	LUT3 #(
		.INIT('h02)
	) name5657 (
		\s5_msel_arb2_state_reg[1]/NET0131 ,
		_w3396_,
		_w3400_,
		_w7558_
	);
	LUT3 #(
		.INIT('h45)
	) name5658 (
		_w7556_,
		_w7557_,
		_w7558_,
		_w7559_
	);
	LUT2 #(
		.INIT('h2)
	) name5659 (
		_w7555_,
		_w7559_,
		_w7560_
	);
	LUT4 #(
		.INIT('h000e)
	) name5660 (
		_w3391_,
		_w3393_,
		_w3396_,
		_w3400_,
		_w7561_
	);
	LUT2 #(
		.INIT('h2)
	) name5661 (
		_w3389_,
		_w7561_,
		_w7562_
	);
	LUT2 #(
		.INIT('h4)
	) name5662 (
		_w3385_,
		_w5735_,
		_w7563_
	);
	LUT3 #(
		.INIT('h54)
	) name5663 (
		\s5_msel_arb2_state_reg[2]/NET0131 ,
		_w3396_,
		_w3400_,
		_w7564_
	);
	LUT2 #(
		.INIT('h1)
	) name5664 (
		\s5_msel_arb2_state_reg[0]/NET0131 ,
		\s5_msel_arb2_state_reg[1]/NET0131 ,
		_w7565_
	);
	LUT3 #(
		.INIT('h10)
	) name5665 (
		_w3385_,
		_w3386_,
		_w7565_,
		_w7566_
	);
	LUT3 #(
		.INIT('h45)
	) name5666 (
		_w7563_,
		_w7564_,
		_w7566_,
		_w7567_
	);
	LUT3 #(
		.INIT('h54)
	) name5667 (
		\s5_msel_arb2_state_reg[1]/NET0131 ,
		_w3396_,
		_w3400_,
		_w7568_
	);
	LUT3 #(
		.INIT('h54)
	) name5668 (
		\s5_msel_arb2_state_reg[0]/NET0131 ,
		_w3391_,
		_w3393_,
		_w7569_
	);
	LUT3 #(
		.INIT('h10)
	) name5669 (
		\s5_msel_arb2_state_reg[2]/NET0131 ,
		_w7568_,
		_w7569_,
		_w7570_
	);
	LUT4 #(
		.INIT('h1110)
	) name5670 (
		_w3385_,
		_w3386_,
		_w3387_,
		_w3388_,
		_w7571_
	);
	LUT3 #(
		.INIT('h10)
	) name5671 (
		\s5_msel_arb2_state_reg[2]/NET0131 ,
		_w3396_,
		_w5734_,
		_w7572_
	);
	LUT3 #(
		.INIT('hd0)
	) name5672 (
		_w3399_,
		_w7571_,
		_w7572_,
		_w7573_
	);
	LUT4 #(
		.INIT('h000e)
	) name5673 (
		_w7562_,
		_w7567_,
		_w7570_,
		_w7573_,
		_w7574_
	);
	LUT2 #(
		.INIT('hb)
	) name5674 (
		_w7560_,
		_w7574_,
		_w7575_
	);
	LUT4 #(
		.INIT('h4447)
	) name5675 (
		\s5_msel_arb3_state_reg[0]/NET0131 ,
		\s5_msel_arb3_state_reg[2]/NET0131 ,
		_w3419_,
		_w5761_,
		_w7576_
	);
	LUT4 #(
		.INIT('h1110)
	) name5676 (
		_w3407_,
		_w3408_,
		_w3414_,
		_w3415_,
		_w7577_
	);
	LUT2 #(
		.INIT('h8)
	) name5677 (
		_w7576_,
		_w7577_,
		_w7578_
	);
	LUT4 #(
		.INIT('hccc8)
	) name5678 (
		\s5_msel_arb3_state_reg[0]/NET0131 ,
		\s5_msel_arb3_state_reg[2]/NET0131 ,
		_w3407_,
		_w3408_,
		_w7579_
	);
	LUT4 #(
		.INIT('h000e)
	) name5679 (
		_w3417_,
		_w3418_,
		_w3419_,
		_w5761_,
		_w7580_
	);
	LUT2 #(
		.INIT('h4)
	) name5680 (
		_w7579_,
		_w7580_,
		_w7581_
	);
	LUT2 #(
		.INIT('h4)
	) name5681 (
		_w3407_,
		_w3410_,
		_w7582_
	);
	LUT4 #(
		.INIT('h000e)
	) name5682 (
		_w3417_,
		_w3418_,
		_w3419_,
		_w3420_,
		_w7583_
	);
	LUT3 #(
		.INIT('hc4)
	) name5683 (
		_w3416_,
		_w7582_,
		_w7583_,
		_w7584_
	);
	LUT4 #(
		.INIT('h5554)
	) name5684 (
		\s5_msel_arb3_state_reg[1]/NET0131 ,
		_w7578_,
		_w7581_,
		_w7584_,
		_w7585_
	);
	LUT3 #(
		.INIT('ha8)
	) name5685 (
		\s5_msel_arb3_state_reg[2]/NET0131 ,
		_w3419_,
		_w3420_,
		_w7586_
	);
	LUT4 #(
		.INIT('h000e)
	) name5686 (
		_w3407_,
		_w3408_,
		_w3417_,
		_w3418_,
		_w7587_
	);
	LUT3 #(
		.INIT('h54)
	) name5687 (
		_w5783_,
		_w7586_,
		_w7587_,
		_w7588_
	);
	LUT3 #(
		.INIT('h0e)
	) name5688 (
		_w3419_,
		_w3420_,
		_w3425_,
		_w7589_
	);
	LUT2 #(
		.INIT('h4)
	) name5689 (
		_w3418_,
		_w5770_,
		_w7590_
	);
	LUT2 #(
		.INIT('h1)
	) name5690 (
		_w3415_,
		_w3417_,
		_w7591_
	);
	LUT3 #(
		.INIT('he0)
	) name5691 (
		_w7589_,
		_w7590_,
		_w7591_,
		_w7592_
	);
	LUT3 #(
		.INIT('h0e)
	) name5692 (
		_w3407_,
		_w3408_,
		_w3417_,
		_w7593_
	);
	LUT3 #(
		.INIT('h2a)
	) name5693 (
		\s5_msel_arb3_state_reg[1]/NET0131 ,
		_w3426_,
		_w7593_,
		_w7594_
	);
	LUT4 #(
		.INIT('hab00)
	) name5694 (
		_w3414_,
		_w7588_,
		_w7592_,
		_w7594_,
		_w7595_
	);
	LUT2 #(
		.INIT('he)
	) name5695 (
		_w7585_,
		_w7595_,
		_w7596_
	);
	LUT4 #(
		.INIT('h0020)
	) name5696 (
		\m2_s6_cyc_o_reg/NET0131 ,
		\rf_conf6_reg[4]/NET0131 ,
		\rf_conf6_reg[5]/NET0131 ,
		\s6_msel_arb2_state_reg[0]/NET0131 ,
		_w7597_
	);
	LUT3 #(
		.INIT('h01)
	) name5697 (
		_w3087_,
		_w3088_,
		_w7597_,
		_w7598_
	);
	LUT4 #(
		.INIT('h2000)
	) name5698 (
		\m3_s6_cyc_o_reg/NET0131 ,
		\rf_conf6_reg[6]/NET0131 ,
		\rf_conf6_reg[7]/NET0131 ,
		\s6_msel_arb2_state_reg[0]/NET0131 ,
		_w7599_
	);
	LUT2 #(
		.INIT('h1)
	) name5699 (
		\s6_msel_arb2_state_reg[2]/NET0131 ,
		_w7599_,
		_w7600_
	);
	LUT4 #(
		.INIT('h00df)
	) name5700 (
		\m2_s6_cyc_o_reg/NET0131 ,
		\rf_conf6_reg[4]/NET0131 ,
		\rf_conf6_reg[5]/NET0131 ,
		\s6_msel_arb2_state_reg[1]/NET0131 ,
		_w7601_
	);
	LUT3 #(
		.INIT('h01)
	) name5701 (
		_w3098_,
		_w3102_,
		_w7601_,
		_w7602_
	);
	LUT4 #(
		.INIT('hcf4f)
	) name5702 (
		_w3091_,
		_w7598_,
		_w7600_,
		_w7602_,
		_w7603_
	);
	LUT4 #(
		.INIT('haaa2)
	) name5703 (
		\s6_msel_arb2_state_reg[1]/NET0131 ,
		\s6_msel_arb2_state_reg[2]/NET0131 ,
		_w3090_,
		_w5887_,
		_w7604_
	);
	LUT4 #(
		.INIT('h000e)
	) name5704 (
		_w3087_,
		_w3088_,
		_w3093_,
		_w3095_,
		_w7605_
	);
	LUT3 #(
		.INIT('h02)
	) name5705 (
		\s6_msel_arb2_state_reg[1]/NET0131 ,
		_w3098_,
		_w3102_,
		_w7606_
	);
	LUT3 #(
		.INIT('h45)
	) name5706 (
		_w7604_,
		_w7605_,
		_w7606_,
		_w7607_
	);
	LUT2 #(
		.INIT('h2)
	) name5707 (
		_w7603_,
		_w7607_,
		_w7608_
	);
	LUT4 #(
		.INIT('h000e)
	) name5708 (
		_w3093_,
		_w3095_,
		_w3098_,
		_w3102_,
		_w7609_
	);
	LUT2 #(
		.INIT('h2)
	) name5709 (
		_w3091_,
		_w7609_,
		_w7610_
	);
	LUT2 #(
		.INIT('h4)
	) name5710 (
		_w3087_,
		_w5897_,
		_w7611_
	);
	LUT3 #(
		.INIT('h54)
	) name5711 (
		\s6_msel_arb2_state_reg[2]/NET0131 ,
		_w3098_,
		_w3102_,
		_w7612_
	);
	LUT2 #(
		.INIT('h1)
	) name5712 (
		\s6_msel_arb2_state_reg[0]/NET0131 ,
		\s6_msel_arb2_state_reg[1]/NET0131 ,
		_w7613_
	);
	LUT3 #(
		.INIT('h10)
	) name5713 (
		_w3087_,
		_w3088_,
		_w7613_,
		_w7614_
	);
	LUT3 #(
		.INIT('h45)
	) name5714 (
		_w7611_,
		_w7612_,
		_w7614_,
		_w7615_
	);
	LUT3 #(
		.INIT('h54)
	) name5715 (
		\s6_msel_arb2_state_reg[1]/NET0131 ,
		_w3098_,
		_w3102_,
		_w7616_
	);
	LUT3 #(
		.INIT('h54)
	) name5716 (
		\s6_msel_arb2_state_reg[0]/NET0131 ,
		_w3093_,
		_w3095_,
		_w7617_
	);
	LUT3 #(
		.INIT('h10)
	) name5717 (
		\s6_msel_arb2_state_reg[2]/NET0131 ,
		_w7616_,
		_w7617_,
		_w7618_
	);
	LUT4 #(
		.INIT('h1110)
	) name5718 (
		_w3087_,
		_w3088_,
		_w3089_,
		_w3090_,
		_w7619_
	);
	LUT3 #(
		.INIT('h10)
	) name5719 (
		\s6_msel_arb2_state_reg[2]/NET0131 ,
		_w3098_,
		_w5896_,
		_w7620_
	);
	LUT3 #(
		.INIT('hd0)
	) name5720 (
		_w3101_,
		_w7619_,
		_w7620_,
		_w7621_
	);
	LUT4 #(
		.INIT('h000e)
	) name5721 (
		_w7610_,
		_w7615_,
		_w7618_,
		_w7621_,
		_w7622_
	);
	LUT2 #(
		.INIT('hb)
	) name5722 (
		_w7608_,
		_w7622_,
		_w7623_
	);
	LUT4 #(
		.INIT('h4447)
	) name5723 (
		\s6_msel_arb3_state_reg[0]/NET0131 ,
		\s6_msel_arb3_state_reg[2]/NET0131 ,
		_w3449_,
		_w5923_,
		_w7624_
	);
	LUT4 #(
		.INIT('h1110)
	) name5724 (
		_w3437_,
		_w3438_,
		_w3444_,
		_w3445_,
		_w7625_
	);
	LUT2 #(
		.INIT('h8)
	) name5725 (
		_w7624_,
		_w7625_,
		_w7626_
	);
	LUT4 #(
		.INIT('hccc8)
	) name5726 (
		\s6_msel_arb3_state_reg[0]/NET0131 ,
		\s6_msel_arb3_state_reg[2]/NET0131 ,
		_w3437_,
		_w3438_,
		_w7627_
	);
	LUT4 #(
		.INIT('h000e)
	) name5727 (
		_w3447_,
		_w3448_,
		_w3449_,
		_w5923_,
		_w7628_
	);
	LUT2 #(
		.INIT('h4)
	) name5728 (
		_w7627_,
		_w7628_,
		_w7629_
	);
	LUT2 #(
		.INIT('h4)
	) name5729 (
		_w3437_,
		_w3440_,
		_w7630_
	);
	LUT4 #(
		.INIT('h000e)
	) name5730 (
		_w3447_,
		_w3448_,
		_w3449_,
		_w3450_,
		_w7631_
	);
	LUT3 #(
		.INIT('hc4)
	) name5731 (
		_w3446_,
		_w7630_,
		_w7631_,
		_w7632_
	);
	LUT4 #(
		.INIT('h5554)
	) name5732 (
		\s6_msel_arb3_state_reg[1]/NET0131 ,
		_w7626_,
		_w7629_,
		_w7632_,
		_w7633_
	);
	LUT3 #(
		.INIT('ha8)
	) name5733 (
		\s6_msel_arb3_state_reg[2]/NET0131 ,
		_w3449_,
		_w3450_,
		_w7634_
	);
	LUT4 #(
		.INIT('h000e)
	) name5734 (
		_w3437_,
		_w3438_,
		_w3447_,
		_w3448_,
		_w7635_
	);
	LUT3 #(
		.INIT('h54)
	) name5735 (
		_w5945_,
		_w7634_,
		_w7635_,
		_w7636_
	);
	LUT3 #(
		.INIT('h0e)
	) name5736 (
		_w3449_,
		_w3450_,
		_w3455_,
		_w7637_
	);
	LUT2 #(
		.INIT('h4)
	) name5737 (
		_w3448_,
		_w5932_,
		_w7638_
	);
	LUT2 #(
		.INIT('h1)
	) name5738 (
		_w3445_,
		_w3447_,
		_w7639_
	);
	LUT3 #(
		.INIT('he0)
	) name5739 (
		_w7637_,
		_w7638_,
		_w7639_,
		_w7640_
	);
	LUT3 #(
		.INIT('h0e)
	) name5740 (
		_w3437_,
		_w3438_,
		_w3447_,
		_w7641_
	);
	LUT3 #(
		.INIT('h2a)
	) name5741 (
		\s6_msel_arb3_state_reg[1]/NET0131 ,
		_w3456_,
		_w7641_,
		_w7642_
	);
	LUT4 #(
		.INIT('hab00)
	) name5742 (
		_w3444_,
		_w7636_,
		_w7640_,
		_w7642_,
		_w7643_
	);
	LUT2 #(
		.INIT('he)
	) name5743 (
		_w7633_,
		_w7643_,
		_w7644_
	);
	LUT3 #(
		.INIT('h54)
	) name5744 (
		\s7_msel_arb2_state_reg[2]/NET0131 ,
		_w6038_,
		_w6039_,
		_w7645_
	);
	LUT4 #(
		.INIT('h1110)
	) name5745 (
		_w6043_,
		_w6044_,
		_w6046_,
		_w6047_,
		_w7646_
	);
	LUT4 #(
		.INIT('h0d0c)
	) name5746 (
		\s7_msel_arb2_state_reg[0]/NET0131 ,
		_w6755_,
		_w7645_,
		_w7646_,
		_w7647_
	);
	LUT3 #(
		.INIT('h01)
	) name5747 (
		\s7_msel_arb2_state_reg[1]/NET0131 ,
		_w6043_,
		_w6044_,
		_w7648_
	);
	LUT2 #(
		.INIT('h8)
	) name5748 (
		_w6751_,
		_w7648_,
		_w7649_
	);
	LUT3 #(
		.INIT('ha8)
	) name5749 (
		\s7_msel_arb2_state_reg[2]/NET0131 ,
		_w6043_,
		_w6044_,
		_w7650_
	);
	LUT4 #(
		.INIT('h1110)
	) name5750 (
		_w6038_,
		_w6039_,
		_w6042_,
		_w6050_,
		_w7651_
	);
	LUT4 #(
		.INIT('h0d0c)
	) name5751 (
		\s7_msel_arb2_state_reg[0]/NET0131 ,
		_w6757_,
		_w7650_,
		_w7651_,
		_w7652_
	);
	LUT2 #(
		.INIT('h8)
	) name5752 (
		_w6043_,
		_w6059_,
		_w7653_
	);
	LUT3 #(
		.INIT('h10)
	) name5753 (
		_w6046_,
		_w6047_,
		_w6059_,
		_w7654_
	);
	LUT4 #(
		.INIT('h080a)
	) name5754 (
		\s7_msel_arb2_state_reg[0]/NET0131 ,
		_w7651_,
		_w7653_,
		_w7654_,
		_w7655_
	);
	LUT4 #(
		.INIT('h0001)
	) name5755 (
		_w7647_,
		_w7649_,
		_w7652_,
		_w7655_,
		_w7656_
	);
	LUT4 #(
		.INIT('h5400)
	) name5756 (
		_w6042_,
		_w6043_,
		_w6044_,
		_w6073_,
		_w7657_
	);
	LUT4 #(
		.INIT('hdf00)
	) name5757 (
		\m4_s7_cyc_o_reg/NET0131 ,
		\rf_conf7_reg[8]/NET0131 ,
		\rf_conf7_reg[9]/NET0131 ,
		\s7_msel_arb2_state_reg[1]/NET0131 ,
		_w7658_
	);
	LUT3 #(
		.INIT('h01)
	) name5758 (
		_w6038_,
		_w6039_,
		_w7658_,
		_w7659_
	);
	LUT4 #(
		.INIT('h0100)
	) name5759 (
		_w6042_,
		_w6046_,
		_w6047_,
		_w6073_,
		_w7660_
	);
	LUT3 #(
		.INIT('h45)
	) name5760 (
		_w7657_,
		_w7659_,
		_w7660_,
		_w7661_
	);
	LUT4 #(
		.INIT('h2000)
	) name5761 (
		\m3_s7_cyc_o_reg/NET0131 ,
		\rf_conf7_reg[6]/NET0131 ,
		\rf_conf7_reg[7]/NET0131 ,
		\s7_msel_arb2_state_reg[1]/NET0131 ,
		_w7662_
	);
	LUT3 #(
		.INIT('h02)
	) name5762 (
		\s7_msel_arb2_state_reg[1]/NET0131 ,
		_w6042_,
		_w6050_,
		_w7663_
	);
	LUT3 #(
		.INIT('h23)
	) name5763 (
		_w7646_,
		_w7662_,
		_w7663_,
		_w7664_
	);
	LUT4 #(
		.INIT('h0054)
	) name5764 (
		_w6042_,
		_w6043_,
		_w6044_,
		_w6050_,
		_w7665_
	);
	LUT4 #(
		.INIT('h00df)
	) name5765 (
		\m1_s7_cyc_o_reg/NET0131 ,
		\rf_conf7_reg[2]/NET0131 ,
		\rf_conf7_reg[3]/NET0131 ,
		\s7_msel_arb2_state_reg[1]/NET0131 ,
		_w7666_
	);
	LUT3 #(
		.INIT('hd0)
	) name5766 (
		_w6751_,
		_w7665_,
		_w7666_,
		_w7667_
	);
	LUT2 #(
		.INIT('h2)
	) name5767 (
		\s7_msel_arb2_state_reg[0]/NET0131 ,
		\s7_msel_arb2_state_reg[2]/NET0131 ,
		_w7668_
	);
	LUT4 #(
		.INIT('h08aa)
	) name5768 (
		_w7661_,
		_w7664_,
		_w7667_,
		_w7668_,
		_w7669_
	);
	LUT2 #(
		.INIT('hb)
	) name5769 (
		_w7656_,
		_w7669_,
		_w7670_
	);
	LUT4 #(
		.INIT('h4447)
	) name5770 (
		\s7_msel_arb3_state_reg[0]/NET0131 ,
		\s7_msel_arb3_state_reg[2]/NET0131 ,
		_w3479_,
		_w6107_,
		_w7671_
	);
	LUT4 #(
		.INIT('h1110)
	) name5771 (
		_w3467_,
		_w3468_,
		_w3474_,
		_w3475_,
		_w7672_
	);
	LUT2 #(
		.INIT('h8)
	) name5772 (
		_w7671_,
		_w7672_,
		_w7673_
	);
	LUT4 #(
		.INIT('hccc8)
	) name5773 (
		\s7_msel_arb3_state_reg[0]/NET0131 ,
		\s7_msel_arb3_state_reg[2]/NET0131 ,
		_w3467_,
		_w3468_,
		_w7674_
	);
	LUT4 #(
		.INIT('h000e)
	) name5774 (
		_w3477_,
		_w3478_,
		_w3479_,
		_w6107_,
		_w7675_
	);
	LUT2 #(
		.INIT('h4)
	) name5775 (
		_w7674_,
		_w7675_,
		_w7676_
	);
	LUT2 #(
		.INIT('h4)
	) name5776 (
		_w3467_,
		_w3470_,
		_w7677_
	);
	LUT4 #(
		.INIT('h000e)
	) name5777 (
		_w3477_,
		_w3478_,
		_w3479_,
		_w3480_,
		_w7678_
	);
	LUT3 #(
		.INIT('hc4)
	) name5778 (
		_w3476_,
		_w7677_,
		_w7678_,
		_w7679_
	);
	LUT4 #(
		.INIT('h5554)
	) name5779 (
		\s7_msel_arb3_state_reg[1]/NET0131 ,
		_w7673_,
		_w7676_,
		_w7679_,
		_w7680_
	);
	LUT3 #(
		.INIT('ha8)
	) name5780 (
		\s7_msel_arb3_state_reg[2]/NET0131 ,
		_w3479_,
		_w3480_,
		_w7681_
	);
	LUT4 #(
		.INIT('h000e)
	) name5781 (
		_w3467_,
		_w3468_,
		_w3477_,
		_w3478_,
		_w7682_
	);
	LUT3 #(
		.INIT('h54)
	) name5782 (
		_w6129_,
		_w7681_,
		_w7682_,
		_w7683_
	);
	LUT3 #(
		.INIT('h0e)
	) name5783 (
		_w3479_,
		_w3480_,
		_w3485_,
		_w7684_
	);
	LUT2 #(
		.INIT('h4)
	) name5784 (
		_w3478_,
		_w6116_,
		_w7685_
	);
	LUT2 #(
		.INIT('h1)
	) name5785 (
		_w3475_,
		_w3477_,
		_w7686_
	);
	LUT3 #(
		.INIT('he0)
	) name5786 (
		_w7684_,
		_w7685_,
		_w7686_,
		_w7687_
	);
	LUT3 #(
		.INIT('h0e)
	) name5787 (
		_w3467_,
		_w3468_,
		_w3477_,
		_w7688_
	);
	LUT3 #(
		.INIT('h2a)
	) name5788 (
		\s7_msel_arb3_state_reg[1]/NET0131 ,
		_w3486_,
		_w7688_,
		_w7689_
	);
	LUT4 #(
		.INIT('hab00)
	) name5789 (
		_w3474_,
		_w7683_,
		_w7687_,
		_w7689_,
		_w7690_
	);
	LUT2 #(
		.INIT('he)
	) name5790 (
		_w7680_,
		_w7690_,
		_w7691_
	);
	LUT4 #(
		.INIT('h0020)
	) name5791 (
		\m2_s8_cyc_o_reg/NET0131 ,
		\rf_conf8_reg[4]/NET0131 ,
		\rf_conf8_reg[5]/NET0131 ,
		\s8_msel_arb2_state_reg[0]/NET0131 ,
		_w7692_
	);
	LUT3 #(
		.INIT('h01)
	) name5792 (
		_w3109_,
		_w3110_,
		_w7692_,
		_w7693_
	);
	LUT4 #(
		.INIT('h2000)
	) name5793 (
		\m3_s8_cyc_o_reg/NET0131 ,
		\rf_conf8_reg[6]/NET0131 ,
		\rf_conf8_reg[7]/NET0131 ,
		\s8_msel_arb2_state_reg[0]/NET0131 ,
		_w7694_
	);
	LUT2 #(
		.INIT('h1)
	) name5794 (
		\s8_msel_arb2_state_reg[2]/NET0131 ,
		_w7694_,
		_w7695_
	);
	LUT4 #(
		.INIT('h00df)
	) name5795 (
		\m2_s8_cyc_o_reg/NET0131 ,
		\rf_conf8_reg[4]/NET0131 ,
		\rf_conf8_reg[5]/NET0131 ,
		\s8_msel_arb2_state_reg[1]/NET0131 ,
		_w7696_
	);
	LUT3 #(
		.INIT('h01)
	) name5796 (
		_w3120_,
		_w3124_,
		_w7696_,
		_w7697_
	);
	LUT4 #(
		.INIT('hcf4f)
	) name5797 (
		_w3113_,
		_w7693_,
		_w7695_,
		_w7697_,
		_w7698_
	);
	LUT4 #(
		.INIT('haaa2)
	) name5798 (
		\s8_msel_arb2_state_reg[1]/NET0131 ,
		\s8_msel_arb2_state_reg[2]/NET0131 ,
		_w3112_,
		_w6233_,
		_w7699_
	);
	LUT4 #(
		.INIT('h000e)
	) name5799 (
		_w3109_,
		_w3110_,
		_w3115_,
		_w3117_,
		_w7700_
	);
	LUT3 #(
		.INIT('h02)
	) name5800 (
		\s8_msel_arb2_state_reg[1]/NET0131 ,
		_w3120_,
		_w3124_,
		_w7701_
	);
	LUT3 #(
		.INIT('h45)
	) name5801 (
		_w7699_,
		_w7700_,
		_w7701_,
		_w7702_
	);
	LUT2 #(
		.INIT('h2)
	) name5802 (
		_w7698_,
		_w7702_,
		_w7703_
	);
	LUT4 #(
		.INIT('h000e)
	) name5803 (
		_w3115_,
		_w3117_,
		_w3120_,
		_w3124_,
		_w7704_
	);
	LUT2 #(
		.INIT('h2)
	) name5804 (
		_w3113_,
		_w7704_,
		_w7705_
	);
	LUT2 #(
		.INIT('h4)
	) name5805 (
		_w3109_,
		_w6243_,
		_w7706_
	);
	LUT3 #(
		.INIT('h54)
	) name5806 (
		\s8_msel_arb2_state_reg[2]/NET0131 ,
		_w3120_,
		_w3124_,
		_w7707_
	);
	LUT2 #(
		.INIT('h1)
	) name5807 (
		\s8_msel_arb2_state_reg[0]/NET0131 ,
		\s8_msel_arb2_state_reg[1]/NET0131 ,
		_w7708_
	);
	LUT3 #(
		.INIT('h10)
	) name5808 (
		_w3109_,
		_w3110_,
		_w7708_,
		_w7709_
	);
	LUT3 #(
		.INIT('h45)
	) name5809 (
		_w7706_,
		_w7707_,
		_w7709_,
		_w7710_
	);
	LUT3 #(
		.INIT('h54)
	) name5810 (
		\s8_msel_arb2_state_reg[1]/NET0131 ,
		_w3120_,
		_w3124_,
		_w7711_
	);
	LUT3 #(
		.INIT('h54)
	) name5811 (
		\s8_msel_arb2_state_reg[0]/NET0131 ,
		_w3115_,
		_w3117_,
		_w7712_
	);
	LUT3 #(
		.INIT('h10)
	) name5812 (
		\s8_msel_arb2_state_reg[2]/NET0131 ,
		_w7711_,
		_w7712_,
		_w7713_
	);
	LUT4 #(
		.INIT('h1110)
	) name5813 (
		_w3109_,
		_w3110_,
		_w3111_,
		_w3112_,
		_w7714_
	);
	LUT3 #(
		.INIT('h10)
	) name5814 (
		\s8_msel_arb2_state_reg[2]/NET0131 ,
		_w3120_,
		_w6242_,
		_w7715_
	);
	LUT3 #(
		.INIT('hd0)
	) name5815 (
		_w3123_,
		_w7714_,
		_w7715_,
		_w7716_
	);
	LUT4 #(
		.INIT('h000e)
	) name5816 (
		_w7705_,
		_w7710_,
		_w7713_,
		_w7716_,
		_w7717_
	);
	LUT2 #(
		.INIT('hb)
	) name5817 (
		_w7703_,
		_w7717_,
		_w7718_
	);
	LUT4 #(
		.INIT('h1110)
	) name5818 (
		_w3498_,
		_w3499_,
		_w3500_,
		_w3501_,
		_w7719_
	);
	LUT3 #(
		.INIT('h54)
	) name5819 (
		\s8_msel_arb3_state_reg[2]/NET0131 ,
		_w3498_,
		_w3511_,
		_w7720_
	);
	LUT4 #(
		.INIT('hafae)
	) name5820 (
		_w3503_,
		_w3506_,
		_w7719_,
		_w7720_,
		_w7721_
	);
	LUT3 #(
		.INIT('he0)
	) name5821 (
		_w3500_,
		_w3501_,
		_w3514_,
		_w7722_
	);
	LUT3 #(
		.INIT('h51)
	) name5822 (
		\s8_msel_arb3_state_reg[1]/NET0131 ,
		_w7721_,
		_w7722_,
		_w7723_
	);
	LUT4 #(
		.INIT('h00a8)
	) name5823 (
		\s8_msel_arb3_state_reg[2]/NET0131 ,
		_w3498_,
		_w3499_,
		_w3504_,
		_w7724_
	);
	LUT3 #(
		.INIT('h0e)
	) name5824 (
		_w3498_,
		_w3499_,
		_w3505_,
		_w7725_
	);
	LUT3 #(
		.INIT('h54)
	) name5825 (
		_w3501_,
		_w3503_,
		_w3511_,
		_w7726_
	);
	LUT2 #(
		.INIT('h1)
	) name5826 (
		_w3500_,
		_w3504_,
		_w7727_
	);
	LUT4 #(
		.INIT('h0155)
	) name5827 (
		_w7724_,
		_w7725_,
		_w7726_,
		_w7727_,
		_w7728_
	);
	LUT4 #(
		.INIT('h007f)
	) name5828 (
		\m3_s8_cyc_o_reg/NET0131 ,
		\rf_conf8_reg[6]/NET0131 ,
		\rf_conf8_reg[7]/NET0131 ,
		\s8_msel_arb3_state_reg[2]/NET0131 ,
		_w7729_
	);
	LUT4 #(
		.INIT('h02aa)
	) name5829 (
		\s8_msel_arb3_state_reg[1]/NET0131 ,
		_w3503_,
		_w3511_,
		_w7729_,
		_w7730_
	);
	LUT2 #(
		.INIT('h8)
	) name5830 (
		_w7728_,
		_w7730_,
		_w7731_
	);
	LUT3 #(
		.INIT('h54)
	) name5831 (
		\s8_msel_arb3_state_reg[1]/NET0131 ,
		_w3503_,
		_w3511_,
		_w7732_
	);
	LUT4 #(
		.INIT('h000e)
	) name5832 (
		_w3498_,
		_w3499_,
		_w3504_,
		_w3505_,
		_w7733_
	);
	LUT4 #(
		.INIT('h1115)
	) name5833 (
		\s8_msel_arb3_state_reg[0]/NET0131 ,
		\s8_msel_arb3_state_reg[2]/NET0131 ,
		_w7732_,
		_w7733_,
		_w7734_
	);
	LUT4 #(
		.INIT('h1110)
	) name5834 (
		_w3500_,
		_w3501_,
		_w3503_,
		_w3511_,
		_w7735_
	);
	LUT3 #(
		.INIT('h54)
	) name5835 (
		\s8_msel_arb3_state_reg[2]/NET0131 ,
		_w3520_,
		_w7735_,
		_w7736_
	);
	LUT3 #(
		.INIT('h02)
	) name5836 (
		\s8_msel_arb3_state_reg[1]/NET0131 ,
		_w3498_,
		_w3499_,
		_w7737_
	);
	LUT4 #(
		.INIT('h0001)
	) name5837 (
		_w3500_,
		_w3501_,
		_w3504_,
		_w3505_,
		_w7738_
	);
	LUT3 #(
		.INIT('h70)
	) name5838 (
		_w3512_,
		_w7737_,
		_w7738_,
		_w7739_
	);
	LUT3 #(
		.INIT('h02)
	) name5839 (
		_w7734_,
		_w7736_,
		_w7739_,
		_w7740_
	);
	LUT4 #(
		.INIT('hffa8)
	) name5840 (
		\s8_msel_arb3_state_reg[0]/NET0131 ,
		_w7723_,
		_w7731_,
		_w7740_,
		_w7741_
	);
	LUT3 #(
		.INIT('h54)
	) name5841 (
		\s9_msel_arb2_state_reg[2]/NET0131 ,
		_w6366_,
		_w6367_,
		_w7742_
	);
	LUT4 #(
		.INIT('h1110)
	) name5842 (
		_w6371_,
		_w6372_,
		_w6374_,
		_w6375_,
		_w7743_
	);
	LUT4 #(
		.INIT('h0d0c)
	) name5843 (
		\s9_msel_arb2_state_reg[0]/NET0131 ,
		_w6773_,
		_w7742_,
		_w7743_,
		_w7744_
	);
	LUT3 #(
		.INIT('h01)
	) name5844 (
		\s9_msel_arb2_state_reg[1]/NET0131 ,
		_w6371_,
		_w6372_,
		_w7745_
	);
	LUT2 #(
		.INIT('h8)
	) name5845 (
		_w6769_,
		_w7745_,
		_w7746_
	);
	LUT3 #(
		.INIT('ha8)
	) name5846 (
		\s9_msel_arb2_state_reg[2]/NET0131 ,
		_w6371_,
		_w6372_,
		_w7747_
	);
	LUT4 #(
		.INIT('h1110)
	) name5847 (
		_w6366_,
		_w6367_,
		_w6370_,
		_w6378_,
		_w7748_
	);
	LUT4 #(
		.INIT('h0d0c)
	) name5848 (
		\s9_msel_arb2_state_reg[0]/NET0131 ,
		_w6775_,
		_w7747_,
		_w7748_,
		_w7749_
	);
	LUT2 #(
		.INIT('h8)
	) name5849 (
		_w6371_,
		_w6387_,
		_w7750_
	);
	LUT3 #(
		.INIT('h10)
	) name5850 (
		_w6374_,
		_w6375_,
		_w6387_,
		_w7751_
	);
	LUT4 #(
		.INIT('h080a)
	) name5851 (
		\s9_msel_arb2_state_reg[0]/NET0131 ,
		_w7748_,
		_w7750_,
		_w7751_,
		_w7752_
	);
	LUT4 #(
		.INIT('h0001)
	) name5852 (
		_w7744_,
		_w7746_,
		_w7749_,
		_w7752_,
		_w7753_
	);
	LUT4 #(
		.INIT('h5400)
	) name5853 (
		_w6370_,
		_w6371_,
		_w6372_,
		_w6401_,
		_w7754_
	);
	LUT4 #(
		.INIT('hdf00)
	) name5854 (
		\m4_s9_cyc_o_reg/NET0131 ,
		\rf_conf9_reg[8]/NET0131 ,
		\rf_conf9_reg[9]/NET0131 ,
		\s9_msel_arb2_state_reg[1]/NET0131 ,
		_w7755_
	);
	LUT3 #(
		.INIT('h01)
	) name5855 (
		_w6366_,
		_w6367_,
		_w7755_,
		_w7756_
	);
	LUT4 #(
		.INIT('h0100)
	) name5856 (
		_w6370_,
		_w6374_,
		_w6375_,
		_w6401_,
		_w7757_
	);
	LUT3 #(
		.INIT('h45)
	) name5857 (
		_w7754_,
		_w7756_,
		_w7757_,
		_w7758_
	);
	LUT4 #(
		.INIT('h2000)
	) name5858 (
		\m3_s9_cyc_o_reg/NET0131 ,
		\rf_conf9_reg[6]/NET0131 ,
		\rf_conf9_reg[7]/NET0131 ,
		\s9_msel_arb2_state_reg[1]/NET0131 ,
		_w7759_
	);
	LUT3 #(
		.INIT('h02)
	) name5859 (
		\s9_msel_arb2_state_reg[1]/NET0131 ,
		_w6370_,
		_w6378_,
		_w7760_
	);
	LUT3 #(
		.INIT('h23)
	) name5860 (
		_w7743_,
		_w7759_,
		_w7760_,
		_w7761_
	);
	LUT4 #(
		.INIT('h0054)
	) name5861 (
		_w6370_,
		_w6371_,
		_w6372_,
		_w6378_,
		_w7762_
	);
	LUT4 #(
		.INIT('h00df)
	) name5862 (
		\m1_s9_cyc_o_reg/NET0131 ,
		\rf_conf9_reg[2]/NET0131 ,
		\rf_conf9_reg[3]/NET0131 ,
		\s9_msel_arb2_state_reg[1]/NET0131 ,
		_w7763_
	);
	LUT3 #(
		.INIT('hd0)
	) name5863 (
		_w6769_,
		_w7762_,
		_w7763_,
		_w7764_
	);
	LUT2 #(
		.INIT('h2)
	) name5864 (
		\s9_msel_arb2_state_reg[0]/NET0131 ,
		\s9_msel_arb2_state_reg[2]/NET0131 ,
		_w7765_
	);
	LUT4 #(
		.INIT('h08aa)
	) name5865 (
		_w7758_,
		_w7761_,
		_w7764_,
		_w7765_,
		_w7766_
	);
	LUT2 #(
		.INIT('hb)
	) name5866 (
		_w7753_,
		_w7766_,
		_w7767_
	);
	LUT4 #(
		.INIT('h0302)
	) name5867 (
		_w6421_,
		_w6425_,
		_w6426_,
		_w6429_,
		_w7768_
	);
	LUT4 #(
		.INIT('h888c)
	) name5868 (
		\s9_msel_arb3_state_reg[1]/NET0131 ,
		\s9_msel_arb3_state_reg[2]/NET0131 ,
		_w6421_,
		_w6429_,
		_w7769_
	);
	LUT4 #(
		.INIT('h0051)
	) name5869 (
		\s9_msel_arb3_state_reg[0]/NET0131 ,
		\s9_msel_arb3_state_reg[1]/NET0131 ,
		_w7768_,
		_w7769_,
		_w7770_
	);
	LUT3 #(
		.INIT('h02)
	) name5870 (
		\s9_msel_arb3_state_reg[1]/NET0131 ,
		_w6421_,
		_w6429_,
		_w7771_
	);
	LUT3 #(
		.INIT('ha2)
	) name5871 (
		_w6779_,
		_w6780_,
		_w7771_,
		_w7772_
	);
	LUT3 #(
		.INIT('h54)
	) name5872 (
		\s9_msel_arb3_state_reg[2]/NET0131 ,
		_w6425_,
		_w6426_,
		_w7773_
	);
	LUT3 #(
		.INIT('h04)
	) name5873 (
		\s9_msel_arb3_state_reg[0]/NET0131 ,
		_w6788_,
		_w7773_,
		_w7774_
	);
	LUT3 #(
		.INIT('h45)
	) name5874 (
		_w7770_,
		_w7772_,
		_w7774_,
		_w7775_
	);
	LUT3 #(
		.INIT('h54)
	) name5875 (
		\s9_msel_arb3_state_reg[2]/NET0131 ,
		_w6425_,
		_w6430_,
		_w7776_
	);
	LUT4 #(
		.INIT('hafae)
	) name5876 (
		_w6422_,
		_w6779_,
		_w7768_,
		_w7776_,
		_w7777_
	);
	LUT4 #(
		.INIT('h02aa)
	) name5877 (
		\s9_msel_arb3_state_reg[1]/NET0131 ,
		_w6421_,
		_w6429_,
		_w6786_,
		_w7778_
	);
	LUT3 #(
		.INIT('h8a)
	) name5878 (
		\s9_msel_arb3_state_reg[0]/NET0131 ,
		_w6429_,
		_w6438_,
		_w7779_
	);
	LUT4 #(
		.INIT('h0054)
	) name5879 (
		_w6423_,
		_w6425_,
		_w6426_,
		_w6427_,
		_w7780_
	);
	LUT3 #(
		.INIT('h02)
	) name5880 (
		\s9_msel_arb3_state_reg[0]/NET0131 ,
		_w6422_,
		_w6430_,
		_w7781_
	);
	LUT3 #(
		.INIT('h45)
	) name5881 (
		_w7779_,
		_w7780_,
		_w7781_,
		_w7782_
	);
	LUT3 #(
		.INIT('h07)
	) name5882 (
		_w7777_,
		_w7778_,
		_w7782_,
		_w7783_
	);
	LUT4 #(
		.INIT('h0504)
	) name5883 (
		_w6421_,
		_w6422_,
		_w6429_,
		_w6430_,
		_w7784_
	);
	LUT4 #(
		.INIT('h0080)
	) name5884 (
		\m0_s9_cyc_o_reg/NET0131 ,
		\rf_conf9_reg[0]/NET0131 ,
		\rf_conf9_reg[1]/NET0131 ,
		\s9_msel_arb3_state_reg[0]/NET0131 ,
		_w7785_
	);
	LUT3 #(
		.INIT('h04)
	) name5885 (
		_w6427_,
		_w6447_,
		_w7785_,
		_w7786_
	);
	LUT3 #(
		.INIT('hd0)
	) name5886 (
		_w6780_,
		_w7784_,
		_w7786_,
		_w7787_
	);
	LUT3 #(
		.INIT('hf2)
	) name5887 (
		_w7775_,
		_w7783_,
		_w7787_,
		_w7788_
	);
	LUT4 #(
		.INIT('h0020)
	) name5888 (
		\m2_s0_cyc_o_reg/NET0131 ,
		\rf_conf0_reg[4]/NET0131 ,
		\rf_conf0_reg[5]/NET0131 ,
		\s0_msel_arb2_state_reg[0]/NET0131 ,
		_w7789_
	);
	LUT3 #(
		.INIT('h01)
	) name5889 (
		_w3131_,
		_w3132_,
		_w7789_,
		_w7790_
	);
	LUT4 #(
		.INIT('h2000)
	) name5890 (
		\m3_s0_cyc_o_reg/NET0131 ,
		\rf_conf0_reg[6]/NET0131 ,
		\rf_conf0_reg[7]/NET0131 ,
		\s0_msel_arb2_state_reg[0]/NET0131 ,
		_w7791_
	);
	LUT2 #(
		.INIT('h1)
	) name5891 (
		\s0_msel_arb2_state_reg[2]/NET0131 ,
		_w7791_,
		_w7792_
	);
	LUT4 #(
		.INIT('h00df)
	) name5892 (
		\m2_s0_cyc_o_reg/NET0131 ,
		\rf_conf0_reg[4]/NET0131 ,
		\rf_conf0_reg[5]/NET0131 ,
		\s0_msel_arb2_state_reg[1]/NET0131 ,
		_w7793_
	);
	LUT3 #(
		.INIT('h01)
	) name5893 (
		_w3142_,
		_w3146_,
		_w7793_,
		_w7794_
	);
	LUT4 #(
		.INIT('hcf4f)
	) name5894 (
		_w3135_,
		_w7790_,
		_w7792_,
		_w7794_,
		_w7795_
	);
	LUT4 #(
		.INIT('haaa2)
	) name5895 (
		\s0_msel_arb2_state_reg[1]/NET0131 ,
		\s0_msel_arb2_state_reg[2]/NET0131 ,
		_w3134_,
		_w6560_,
		_w7796_
	);
	LUT4 #(
		.INIT('h000e)
	) name5896 (
		_w3131_,
		_w3132_,
		_w3137_,
		_w3139_,
		_w7797_
	);
	LUT3 #(
		.INIT('h02)
	) name5897 (
		\s0_msel_arb2_state_reg[1]/NET0131 ,
		_w3142_,
		_w3146_,
		_w7798_
	);
	LUT3 #(
		.INIT('h45)
	) name5898 (
		_w7796_,
		_w7797_,
		_w7798_,
		_w7799_
	);
	LUT2 #(
		.INIT('h2)
	) name5899 (
		_w7795_,
		_w7799_,
		_w7800_
	);
	LUT4 #(
		.INIT('h000e)
	) name5900 (
		_w3137_,
		_w3139_,
		_w3142_,
		_w3146_,
		_w7801_
	);
	LUT2 #(
		.INIT('h2)
	) name5901 (
		_w3135_,
		_w7801_,
		_w7802_
	);
	LUT2 #(
		.INIT('h4)
	) name5902 (
		_w3131_,
		_w6570_,
		_w7803_
	);
	LUT3 #(
		.INIT('h54)
	) name5903 (
		\s0_msel_arb2_state_reg[2]/NET0131 ,
		_w3142_,
		_w3146_,
		_w7804_
	);
	LUT2 #(
		.INIT('h1)
	) name5904 (
		\s0_msel_arb2_state_reg[0]/NET0131 ,
		\s0_msel_arb2_state_reg[1]/NET0131 ,
		_w7805_
	);
	LUT3 #(
		.INIT('h10)
	) name5905 (
		_w3131_,
		_w3132_,
		_w7805_,
		_w7806_
	);
	LUT3 #(
		.INIT('h45)
	) name5906 (
		_w7803_,
		_w7804_,
		_w7806_,
		_w7807_
	);
	LUT3 #(
		.INIT('h54)
	) name5907 (
		\s0_msel_arb2_state_reg[1]/NET0131 ,
		_w3142_,
		_w3146_,
		_w7808_
	);
	LUT3 #(
		.INIT('h54)
	) name5908 (
		\s0_msel_arb2_state_reg[0]/NET0131 ,
		_w3137_,
		_w3139_,
		_w7809_
	);
	LUT3 #(
		.INIT('h10)
	) name5909 (
		\s0_msel_arb2_state_reg[2]/NET0131 ,
		_w7808_,
		_w7809_,
		_w7810_
	);
	LUT4 #(
		.INIT('h1110)
	) name5910 (
		_w3131_,
		_w3132_,
		_w3133_,
		_w3134_,
		_w7811_
	);
	LUT3 #(
		.INIT('h10)
	) name5911 (
		\s0_msel_arb2_state_reg[2]/NET0131 ,
		_w3142_,
		_w6569_,
		_w7812_
	);
	LUT3 #(
		.INIT('hd0)
	) name5912 (
		_w3145_,
		_w7811_,
		_w7812_,
		_w7813_
	);
	LUT4 #(
		.INIT('h000e)
	) name5913 (
		_w7802_,
		_w7807_,
		_w7810_,
		_w7813_,
		_w7814_
	);
	LUT2 #(
		.INIT('hb)
	) name5914 (
		_w7800_,
		_w7814_,
		_w7815_
	);
	LUT4 #(
		.INIT('h4447)
	) name5915 (
		\s0_msel_arb3_state_reg[0]/NET0131 ,
		\s0_msel_arb3_state_reg[2]/NET0131 ,
		_w3541_,
		_w6596_,
		_w7816_
	);
	LUT4 #(
		.INIT('h1110)
	) name5916 (
		_w3529_,
		_w3530_,
		_w3536_,
		_w3537_,
		_w7817_
	);
	LUT2 #(
		.INIT('h8)
	) name5917 (
		_w7816_,
		_w7817_,
		_w7818_
	);
	LUT4 #(
		.INIT('hccc8)
	) name5918 (
		\s0_msel_arb3_state_reg[0]/NET0131 ,
		\s0_msel_arb3_state_reg[2]/NET0131 ,
		_w3529_,
		_w3530_,
		_w7819_
	);
	LUT4 #(
		.INIT('h000e)
	) name5919 (
		_w3539_,
		_w3540_,
		_w3541_,
		_w6596_,
		_w7820_
	);
	LUT2 #(
		.INIT('h4)
	) name5920 (
		_w7819_,
		_w7820_,
		_w7821_
	);
	LUT2 #(
		.INIT('h4)
	) name5921 (
		_w3529_,
		_w3532_,
		_w7822_
	);
	LUT4 #(
		.INIT('h000e)
	) name5922 (
		_w3539_,
		_w3540_,
		_w3541_,
		_w3542_,
		_w7823_
	);
	LUT3 #(
		.INIT('hc4)
	) name5923 (
		_w3538_,
		_w7822_,
		_w7823_,
		_w7824_
	);
	LUT4 #(
		.INIT('h5554)
	) name5924 (
		\s0_msel_arb3_state_reg[1]/NET0131 ,
		_w7818_,
		_w7821_,
		_w7824_,
		_w7825_
	);
	LUT3 #(
		.INIT('ha8)
	) name5925 (
		\s0_msel_arb3_state_reg[2]/NET0131 ,
		_w3541_,
		_w3542_,
		_w7826_
	);
	LUT4 #(
		.INIT('h000e)
	) name5926 (
		_w3529_,
		_w3530_,
		_w3539_,
		_w3540_,
		_w7827_
	);
	LUT3 #(
		.INIT('h54)
	) name5927 (
		_w6618_,
		_w7826_,
		_w7827_,
		_w7828_
	);
	LUT3 #(
		.INIT('h0e)
	) name5928 (
		_w3541_,
		_w3542_,
		_w3547_,
		_w7829_
	);
	LUT2 #(
		.INIT('h4)
	) name5929 (
		_w3540_,
		_w6605_,
		_w7830_
	);
	LUT2 #(
		.INIT('h1)
	) name5930 (
		_w3537_,
		_w3539_,
		_w7831_
	);
	LUT3 #(
		.INIT('he0)
	) name5931 (
		_w7829_,
		_w7830_,
		_w7831_,
		_w7832_
	);
	LUT3 #(
		.INIT('h0e)
	) name5932 (
		_w3529_,
		_w3530_,
		_w3539_,
		_w7833_
	);
	LUT3 #(
		.INIT('h2a)
	) name5933 (
		\s0_msel_arb3_state_reg[1]/NET0131 ,
		_w3548_,
		_w7833_,
		_w7834_
	);
	LUT4 #(
		.INIT('hab00)
	) name5934 (
		_w3536_,
		_w7828_,
		_w7832_,
		_w7834_,
		_w7835_
	);
	LUT2 #(
		.INIT('he)
	) name5935 (
		_w7825_,
		_w7835_,
		_w7836_
	);
	LUT4 #(
		.INIT('h000e)
	) name5936 (
		_w3564_,
		_w3565_,
		_w3567_,
		_w3568_,
		_w7837_
	);
	LUT3 #(
		.INIT('h02)
	) name5937 (
		\s10_msel_arb1_state_reg[2]/NET0131 ,
		_w3559_,
		_w3561_,
		_w7838_
	);
	LUT4 #(
		.INIT('h5100)
	) name5938 (
		\s10_msel_arb1_state_reg[0]/NET0131 ,
		_w3578_,
		_w7837_,
		_w7838_,
		_w7839_
	);
	LUT4 #(
		.INIT('h000e)
	) name5939 (
		_w3567_,
		_w3568_,
		_w3570_,
		_w3571_,
		_w7840_
	);
	LUT3 #(
		.INIT('h54)
	) name5940 (
		\s10_msel_arb1_state_reg[2]/NET0131 ,
		_w3564_,
		_w3565_,
		_w7841_
	);
	LUT4 #(
		.INIT('h0031)
	) name5941 (
		_w3577_,
		_w7837_,
		_w7840_,
		_w7841_,
		_w7842_
	);
	LUT2 #(
		.INIT('h4)
	) name5942 (
		\s10_msel_arb1_state_reg[0]/NET0131 ,
		\s10_msel_arb1_state_reg[1]/NET0131 ,
		_w7843_
	);
	LUT3 #(
		.INIT('h45)
	) name5943 (
		_w7839_,
		_w7842_,
		_w7843_,
		_w7844_
	);
	LUT4 #(
		.INIT('h000e)
	) name5944 (
		_w3559_,
		_w3561_,
		_w3564_,
		_w3565_,
		_w7845_
	);
	LUT3 #(
		.INIT('h02)
	) name5945 (
		\s10_msel_arb1_state_reg[0]/NET0131 ,
		_w3567_,
		_w3568_,
		_w7846_
	);
	LUT4 #(
		.INIT('hf700)
	) name5946 (
		\m7_s10_cyc_o_reg/NET0131 ,
		\rf_conf10_reg[14]/NET0131 ,
		\rf_conf10_reg[15]/NET0131 ,
		\s10_msel_arb1_state_reg[2]/NET0131 ,
		_w7847_
	);
	LUT2 #(
		.INIT('h4)
	) name5947 (
		_w4013_,
		_w7847_,
		_w7848_
	);
	LUT3 #(
		.INIT('hb0)
	) name5948 (
		_w7845_,
		_w7846_,
		_w7848_,
		_w7849_
	);
	LUT3 #(
		.INIT('h02)
	) name5949 (
		\s10_msel_arb1_state_reg[1]/NET0131 ,
		_w3559_,
		_w3561_,
		_w7850_
	);
	LUT4 #(
		.INIT('h0800)
	) name5950 (
		\m3_s10_cyc_o_reg/NET0131 ,
		\rf_conf10_reg[6]/NET0131 ,
		\rf_conf10_reg[7]/NET0131 ,
		\s10_msel_arb1_state_reg[0]/NET0131 ,
		_w7851_
	);
	LUT3 #(
		.INIT('ha8)
	) name5951 (
		\s10_msel_arb1_state_reg[1]/NET0131 ,
		\s10_msel_arb1_state_reg[2]/NET0131 ,
		_w7851_,
		_w7852_
	);
	LUT3 #(
		.INIT('h0b)
	) name5952 (
		_w7840_,
		_w7850_,
		_w7852_,
		_w7853_
	);
	LUT4 #(
		.INIT('h1110)
	) name5953 (
		_w3559_,
		_w3561_,
		_w3570_,
		_w3571_,
		_w7854_
	);
	LUT3 #(
		.INIT('h10)
	) name5954 (
		_w3567_,
		_w3575_,
		_w4002_,
		_w7855_
	);
	LUT3 #(
		.INIT('hd0)
	) name5955 (
		_w3566_,
		_w7854_,
		_w7855_,
		_w7856_
	);
	LUT3 #(
		.INIT('h20)
	) name5956 (
		\s10_msel_arb1_state_reg[0]/NET0131 ,
		\s10_msel_arb1_state_reg[1]/NET0131 ,
		\s10_msel_arb1_state_reg[2]/NET0131 ,
		_w7857_
	);
	LUT2 #(
		.INIT('h4)
	) name5957 (
		_w3559_,
		_w7857_,
		_w7858_
	);
	LUT3 #(
		.INIT('hd0)
	) name5958 (
		_w3578_,
		_w7837_,
		_w7858_,
		_w7859_
	);
	LUT4 #(
		.INIT('h000e)
	) name5959 (
		_w7849_,
		_w7853_,
		_w7856_,
		_w7859_,
		_w7860_
	);
	LUT2 #(
		.INIT('h7)
	) name5960 (
		_w7844_,
		_w7860_,
		_w7861_
	);
	LUT4 #(
		.INIT('h000e)
	) name5961 (
		_w3587_,
		_w3588_,
		_w3590_,
		_w3591_,
		_w7862_
	);
	LUT4 #(
		.INIT('h00f7)
	) name5962 (
		\m1_s11_cyc_o_reg/NET0131 ,
		\rf_conf11_reg[2]/NET0131 ,
		\rf_conf11_reg[3]/NET0131 ,
		\s11_msel_arb1_state_reg[1]/NET0131 ,
		_w7863_
	);
	LUT2 #(
		.INIT('h4)
	) name5963 (
		_w3598_,
		_w7863_,
		_w7864_
	);
	LUT4 #(
		.INIT('h5100)
	) name5964 (
		\s11_msel_arb1_state_reg[2]/NET0131 ,
		_w3605_,
		_w7862_,
		_w7864_,
		_w7865_
	);
	LUT4 #(
		.INIT('h1110)
	) name5965 (
		_w3587_,
		_w3588_,
		_w3594_,
		_w3601_,
		_w7866_
	);
	LUT3 #(
		.INIT('h02)
	) name5966 (
		\s11_msel_arb1_state_reg[0]/NET0131 ,
		_w3590_,
		_w3591_,
		_w7867_
	);
	LUT4 #(
		.INIT('h0008)
	) name5967 (
		\m2_s11_cyc_o_reg/NET0131 ,
		\rf_conf11_reg[4]/NET0131 ,
		\rf_conf11_reg[5]/NET0131 ,
		\s11_msel_arb1_state_reg[0]/NET0131 ,
		_w7868_
	);
	LUT2 #(
		.INIT('h1)
	) name5968 (
		_w3584_,
		_w7868_,
		_w7869_
	);
	LUT4 #(
		.INIT('h20aa)
	) name5969 (
		_w3585_,
		_w7866_,
		_w7867_,
		_w7869_,
		_w7870_
	);
	LUT2 #(
		.INIT('h1)
	) name5970 (
		_w7865_,
		_w7870_,
		_w7871_
	);
	LUT3 #(
		.INIT('h04)
	) name5971 (
		_w3591_,
		_w4186_,
		_w7866_,
		_w7872_
	);
	LUT4 #(
		.INIT('h0032)
	) name5972 (
		_w3584_,
		_w3594_,
		_w3600_,
		_w3601_,
		_w7873_
	);
	LUT3 #(
		.INIT('h04)
	) name5973 (
		_w3591_,
		_w3609_,
		_w4170_,
		_w7874_
	);
	LUT3 #(
		.INIT('hd0)
	) name5974 (
		_w3589_,
		_w7873_,
		_w7874_,
		_w7875_
	);
	LUT3 #(
		.INIT('hc8)
	) name5975 (
		_w3587_,
		_w3595_,
		_w3612_,
		_w7876_
	);
	LUT4 #(
		.INIT('h0054)
	) name5976 (
		_w3584_,
		_w3590_,
		_w3591_,
		_w3600_,
		_w7877_
	);
	LUT3 #(
		.INIT('h04)
	) name5977 (
		_w3594_,
		_w3595_,
		_w3601_,
		_w7878_
	);
	LUT3 #(
		.INIT('h45)
	) name5978 (
		_w7876_,
		_w7877_,
		_w7878_,
		_w7879_
	);
	LUT3 #(
		.INIT('h10)
	) name5979 (
		_w7872_,
		_w7875_,
		_w7879_,
		_w7880_
	);
	LUT2 #(
		.INIT('h7)
	) name5980 (
		_w7871_,
		_w7880_,
		_w7881_
	);
	LUT4 #(
		.INIT('h000e)
	) name5981 (
		_w3622_,
		_w3623_,
		_w3625_,
		_w3626_,
		_w7882_
	);
	LUT3 #(
		.INIT('h01)
	) name5982 (
		\s12_msel_arb1_state_reg[1]/NET0131 ,
		_w3619_,
		_w3620_,
		_w7883_
	);
	LUT3 #(
		.INIT('hd0)
	) name5983 (
		_w3641_,
		_w7882_,
		_w7883_,
		_w7884_
	);
	LUT2 #(
		.INIT('h4)
	) name5984 (
		\s12_msel_arb1_state_reg[0]/NET0131 ,
		\s12_msel_arb1_state_reg[1]/NET0131 ,
		_w7885_
	);
	LUT3 #(
		.INIT('he0)
	) name5985 (
		_w3630_,
		_w3631_,
		_w7885_,
		_w7886_
	);
	LUT4 #(
		.INIT('h0302)
	) name5986 (
		_w3619_,
		_w3622_,
		_w3623_,
		_w3639_,
		_w7887_
	);
	LUT3 #(
		.INIT('h10)
	) name5987 (
		_w3625_,
		_w3626_,
		_w7885_,
		_w7888_
	);
	LUT3 #(
		.INIT('h45)
	) name5988 (
		_w7886_,
		_w7887_,
		_w7888_,
		_w7889_
	);
	LUT3 #(
		.INIT('h45)
	) name5989 (
		\s12_msel_arb1_state_reg[2]/NET0131 ,
		_w7884_,
		_w7889_,
		_w7890_
	);
	LUT4 #(
		.INIT('h000e)
	) name5990 (
		_w3625_,
		_w3626_,
		_w3630_,
		_w3631_,
		_w7891_
	);
	LUT3 #(
		.INIT('ha2)
	) name5991 (
		_w3624_,
		_w3640_,
		_w7891_,
		_w7892_
	);
	LUT3 #(
		.INIT('h70)
	) name5992 (
		\s12_msel_arb1_state_reg[0]/NET0131 ,
		\s12_msel_arb1_state_reg[1]/NET0131 ,
		\s12_msel_arb1_state_reg[2]/NET0131 ,
		_w7893_
	);
	LUT3 #(
		.INIT('h40)
	) name5993 (
		\s12_msel_arb1_state_reg[0]/NET0131 ,
		\s12_msel_arb1_state_reg[1]/NET0131 ,
		\s12_msel_arb1_state_reg[2]/NET0131 ,
		_w7894_
	);
	LUT4 #(
		.INIT('h0001)
	) name5994 (
		_w3622_,
		_w3623_,
		_w3630_,
		_w3631_,
		_w7895_
	);
	LUT3 #(
		.INIT('h10)
	) name5995 (
		_w3626_,
		_w3636_,
		_w7893_,
		_w7896_
	);
	LUT3 #(
		.INIT('h45)
	) name5996 (
		_w7894_,
		_w7895_,
		_w7896_,
		_w7897_
	);
	LUT3 #(
		.INIT('ha8)
	) name5997 (
		\s12_msel_arb1_state_reg[2]/NET0131 ,
		_w3622_,
		_w3630_,
		_w7898_
	);
	LUT4 #(
		.INIT('hcfce)
	) name5998 (
		_w3627_,
		_w3631_,
		_w7887_,
		_w7898_,
		_w7899_
	);
	LUT4 #(
		.INIT('h0c4c)
	) name5999 (
		_w3619_,
		_w3629_,
		_w3638_,
		_w3639_,
		_w7900_
	);
	LUT4 #(
		.INIT('h0eee)
	) name6000 (
		_w7892_,
		_w7897_,
		_w7899_,
		_w7900_,
		_w7901_
	);
	LUT2 #(
		.INIT('hb)
	) name6001 (
		_w7890_,
		_w7901_,
		_w7902_
	);
	LUT4 #(
		.INIT('h000e)
	) name6002 (
		_w3650_,
		_w3651_,
		_w3653_,
		_w3654_,
		_w7903_
	);
	LUT3 #(
		.INIT('h02)
	) name6003 (
		\s13_msel_arb1_state_reg[2]/NET0131 ,
		_w3645_,
		_w3647_,
		_w7904_
	);
	LUT4 #(
		.INIT('h5100)
	) name6004 (
		\s13_msel_arb1_state_reg[0]/NET0131 ,
		_w3664_,
		_w7903_,
		_w7904_,
		_w7905_
	);
	LUT4 #(
		.INIT('h000e)
	) name6005 (
		_w3653_,
		_w3654_,
		_w3656_,
		_w3657_,
		_w7906_
	);
	LUT3 #(
		.INIT('h54)
	) name6006 (
		\s13_msel_arb1_state_reg[2]/NET0131 ,
		_w3650_,
		_w3651_,
		_w7907_
	);
	LUT4 #(
		.INIT('h0031)
	) name6007 (
		_w3663_,
		_w7903_,
		_w7906_,
		_w7907_,
		_w7908_
	);
	LUT2 #(
		.INIT('h4)
	) name6008 (
		\s13_msel_arb1_state_reg[0]/NET0131 ,
		\s13_msel_arb1_state_reg[1]/NET0131 ,
		_w7909_
	);
	LUT3 #(
		.INIT('h45)
	) name6009 (
		_w7905_,
		_w7908_,
		_w7909_,
		_w7910_
	);
	LUT4 #(
		.INIT('h000e)
	) name6010 (
		_w3645_,
		_w3647_,
		_w3650_,
		_w3651_,
		_w7911_
	);
	LUT3 #(
		.INIT('h02)
	) name6011 (
		\s13_msel_arb1_state_reg[0]/NET0131 ,
		_w3653_,
		_w3654_,
		_w7912_
	);
	LUT4 #(
		.INIT('hf700)
	) name6012 (
		\m7_s13_cyc_o_reg/NET0131 ,
		\rf_conf13_reg[14]/NET0131 ,
		\rf_conf13_reg[15]/NET0131 ,
		\s13_msel_arb1_state_reg[2]/NET0131 ,
		_w7913_
	);
	LUT2 #(
		.INIT('h4)
	) name6013 (
		_w4538_,
		_w7913_,
		_w7914_
	);
	LUT3 #(
		.INIT('hb0)
	) name6014 (
		_w7911_,
		_w7912_,
		_w7914_,
		_w7915_
	);
	LUT3 #(
		.INIT('h02)
	) name6015 (
		\s13_msel_arb1_state_reg[1]/NET0131 ,
		_w3645_,
		_w3647_,
		_w7916_
	);
	LUT4 #(
		.INIT('h0800)
	) name6016 (
		\m3_s13_cyc_o_reg/NET0131 ,
		\rf_conf13_reg[6]/NET0131 ,
		\rf_conf13_reg[7]/NET0131 ,
		\s13_msel_arb1_state_reg[0]/NET0131 ,
		_w7917_
	);
	LUT3 #(
		.INIT('ha8)
	) name6017 (
		\s13_msel_arb1_state_reg[1]/NET0131 ,
		\s13_msel_arb1_state_reg[2]/NET0131 ,
		_w7917_,
		_w7918_
	);
	LUT3 #(
		.INIT('h0b)
	) name6018 (
		_w7906_,
		_w7916_,
		_w7918_,
		_w7919_
	);
	LUT4 #(
		.INIT('h1110)
	) name6019 (
		_w3645_,
		_w3647_,
		_w3656_,
		_w3657_,
		_w7920_
	);
	LUT3 #(
		.INIT('h10)
	) name6020 (
		_w3653_,
		_w3661_,
		_w4527_,
		_w7921_
	);
	LUT3 #(
		.INIT('hd0)
	) name6021 (
		_w3652_,
		_w7920_,
		_w7921_,
		_w7922_
	);
	LUT3 #(
		.INIT('h20)
	) name6022 (
		\s13_msel_arb1_state_reg[0]/NET0131 ,
		\s13_msel_arb1_state_reg[1]/NET0131 ,
		\s13_msel_arb1_state_reg[2]/NET0131 ,
		_w7923_
	);
	LUT2 #(
		.INIT('h4)
	) name6023 (
		_w3645_,
		_w7923_,
		_w7924_
	);
	LUT3 #(
		.INIT('hd0)
	) name6024 (
		_w3664_,
		_w7903_,
		_w7924_,
		_w7925_
	);
	LUT4 #(
		.INIT('h000e)
	) name6025 (
		_w7915_,
		_w7919_,
		_w7922_,
		_w7925_,
		_w7926_
	);
	LUT2 #(
		.INIT('h7)
	) name6026 (
		_w7910_,
		_w7926_,
		_w7927_
	);
	LUT4 #(
		.INIT('h0001)
	) name6027 (
		_w3673_,
		_w3674_,
		_w3683_,
		_w3688_,
		_w7928_
	);
	LUT3 #(
		.INIT('ha8)
	) name6028 (
		\s14_msel_arb1_state_reg[1]/NET0131 ,
		_w4709_,
		_w7928_,
		_w7929_
	);
	LUT3 #(
		.INIT('h10)
	) name6029 (
		_w3673_,
		_w3674_,
		_w4709_,
		_w7930_
	);
	LUT4 #(
		.INIT('h3332)
	) name6030 (
		\s14_msel_arb1_state_reg[0]/NET0131 ,
		\s14_msel_arb1_state_reg[1]/NET0131 ,
		_w3673_,
		_w3674_,
		_w7931_
	);
	LUT4 #(
		.INIT('h000e)
	) name6031 (
		_w3678_,
		_w3682_,
		_w3683_,
		_w3688_,
		_w7932_
	);
	LUT4 #(
		.INIT('h3031)
	) name6032 (
		_w3671_,
		_w7930_,
		_w7931_,
		_w7932_,
		_w7933_
	);
	LUT3 #(
		.INIT('h8a)
	) name6033 (
		\s14_msel_arb1_state_reg[2]/NET0131 ,
		_w7929_,
		_w7933_,
		_w7934_
	);
	LUT4 #(
		.INIT('h0100)
	) name6034 (
		_w3673_,
		_w3674_,
		_w3688_,
		_w4694_,
		_w7935_
	);
	LUT2 #(
		.INIT('h4)
	) name6035 (
		_w3683_,
		_w7935_,
		_w7936_
	);
	LUT4 #(
		.INIT('h000e)
	) name6036 (
		_w3670_,
		_w3671_,
		_w3673_,
		_w3674_,
		_w7937_
	);
	LUT3 #(
		.INIT('h10)
	) name6037 (
		_w3681_,
		_w3683_,
		_w4691_,
		_w7938_
	);
	LUT3 #(
		.INIT('hd0)
	) name6038 (
		_w3689_,
		_w7937_,
		_w7938_,
		_w7939_
	);
	LUT2 #(
		.INIT('h1)
	) name6039 (
		_w3678_,
		_w3685_,
		_w7940_
	);
	LUT3 #(
		.INIT('h8a)
	) name6040 (
		_w4694_,
		_w7937_,
		_w7940_,
		_w7941_
	);
	LUT2 #(
		.INIT('h4)
	) name6041 (
		_w3674_,
		_w4716_,
		_w7942_
	);
	LUT3 #(
		.INIT('hd0)
	) name6042 (
		_w3672_,
		_w7932_,
		_w7942_,
		_w7943_
	);
	LUT4 #(
		.INIT('h0001)
	) name6043 (
		_w7936_,
		_w7939_,
		_w7941_,
		_w7943_,
		_w7944_
	);
	LUT2 #(
		.INIT('hb)
	) name6044 (
		_w7934_,
		_w7944_,
		_w7945_
	);
	LUT4 #(
		.INIT('h1110)
	) name6045 (
		_w2878_,
		_w2879_,
		_w2886_,
		_w2887_,
		_w7946_
	);
	LUT3 #(
		.INIT('hc4)
	) name6046 (
		_w2882_,
		_w2939_,
		_w7946_,
		_w7947_
	);
	LUT4 #(
		.INIT('h00f7)
	) name6047 (
		\m3_s15_cyc_o_reg/NET0131 ,
		\rf_conf15_reg[6]/NET0131 ,
		\rf_conf15_reg[7]/NET0131 ,
		\s15_msel_arb1_state_reg[2]/NET0131 ,
		_w7948_
	);
	LUT2 #(
		.INIT('h2)
	) name6048 (
		\s15_msel_arb1_state_reg[1]/NET0131 ,
		_w7948_,
		_w7949_
	);
	LUT4 #(
		.INIT('h000e)
	) name6049 (
		_w2880_,
		_w2881_,
		_w2884_,
		_w2885_,
		_w7950_
	);
	LUT3 #(
		.INIT('h02)
	) name6050 (
		\s15_msel_arb1_state_reg[1]/NET0131 ,
		_w2886_,
		_w2887_,
		_w7951_
	);
	LUT3 #(
		.INIT('h45)
	) name6051 (
		_w7949_,
		_w7950_,
		_w7951_,
		_w7952_
	);
	LUT3 #(
		.INIT('h02)
	) name6052 (
		\s15_msel_arb1_state_reg[0]/NET0131 ,
		_w7947_,
		_w7952_,
		_w7953_
	);
	LUT4 #(
		.INIT('h0800)
	) name6053 (
		\m5_s15_cyc_o_reg/NET0131 ,
		\rf_conf15_reg[10]/NET0131 ,
		\rf_conf15_reg[11]/NET0131 ,
		\s15_msel_arb1_state_reg[2]/NET0131 ,
		_w7954_
	);
	LUT4 #(
		.INIT('h000e)
	) name6054 (
		_w2878_,
		_w2879_,
		_w2880_,
		_w2881_,
		_w7955_
	);
	LUT3 #(
		.INIT('h02)
	) name6055 (
		\s15_msel_arb1_state_reg[2]/NET0131 ,
		_w2884_,
		_w2885_,
		_w7956_
	);
	LUT4 #(
		.INIT('h1011)
	) name6056 (
		\s15_msel_arb1_state_reg[1]/NET0131 ,
		_w7954_,
		_w7955_,
		_w7956_,
		_w7957_
	);
	LUT4 #(
		.INIT('h000e)
	) name6057 (
		_w2884_,
		_w2885_,
		_w2886_,
		_w2887_,
		_w7958_
	);
	LUT3 #(
		.INIT('h01)
	) name6058 (
		\s15_msel_arb1_state_reg[2]/NET0131 ,
		_w2878_,
		_w2879_,
		_w7959_
	);
	LUT4 #(
		.INIT('h2022)
	) name6059 (
		\s15_msel_arb1_state_reg[0]/NET0131 ,
		_w4817_,
		_w7958_,
		_w7959_,
		_w7960_
	);
	LUT2 #(
		.INIT('h8)
	) name6060 (
		_w7957_,
		_w7960_,
		_w7961_
	);
	LUT3 #(
		.INIT('h54)
	) name6061 (
		\s15_msel_arb1_state_reg[1]/NET0131 ,
		_w2880_,
		_w2881_,
		_w7962_
	);
	LUT4 #(
		.INIT('h4445)
	) name6062 (
		\s15_msel_arb1_state_reg[0]/NET0131 ,
		\s15_msel_arb1_state_reg[2]/NET0131 ,
		_w7946_,
		_w7962_,
		_w7963_
	);
	LUT2 #(
		.INIT('h4)
	) name6063 (
		\s15_msel_arb1_state_reg[1]/NET0131 ,
		\s15_msel_arb1_state_reg[2]/NET0131 ,
		_w7964_
	);
	LUT3 #(
		.INIT('he0)
	) name6064 (
		_w2886_,
		_w2887_,
		_w7964_,
		_w7965_
	);
	LUT3 #(
		.INIT('h07)
	) name6065 (
		\s15_msel_arb1_state_reg[2]/NET0131 ,
		_w7950_,
		_w7965_,
		_w7966_
	);
	LUT3 #(
		.INIT('h02)
	) name6066 (
		\s15_msel_arb1_state_reg[1]/NET0131 ,
		_w2880_,
		_w2881_,
		_w7967_
	);
	LUT4 #(
		.INIT('h0001)
	) name6067 (
		_w2878_,
		_w2879_,
		_w2884_,
		_w2885_,
		_w7968_
	);
	LUT3 #(
		.INIT('h70)
	) name6068 (
		_w2888_,
		_w7967_,
		_w7968_,
		_w7969_
	);
	LUT3 #(
		.INIT('h08)
	) name6069 (
		_w7963_,
		_w7966_,
		_w7969_,
		_w7970_
	);
	LUT3 #(
		.INIT('hfe)
	) name6070 (
		_w7953_,
		_w7961_,
		_w7970_,
		_w7971_
	);
	LUT4 #(
		.INIT('h0001)
	) name6071 (
		_w3699_,
		_w3700_,
		_w3709_,
		_w3714_,
		_w7972_
	);
	LUT3 #(
		.INIT('ha8)
	) name6072 (
		\s1_msel_arb1_state_reg[1]/NET0131 ,
		_w4999_,
		_w7972_,
		_w7973_
	);
	LUT3 #(
		.INIT('h10)
	) name6073 (
		_w3699_,
		_w3700_,
		_w4999_,
		_w7974_
	);
	LUT4 #(
		.INIT('h3332)
	) name6074 (
		\s1_msel_arb1_state_reg[0]/NET0131 ,
		\s1_msel_arb1_state_reg[1]/NET0131 ,
		_w3699_,
		_w3700_,
		_w7975_
	);
	LUT4 #(
		.INIT('h000e)
	) name6075 (
		_w3704_,
		_w3708_,
		_w3709_,
		_w3714_,
		_w7976_
	);
	LUT4 #(
		.INIT('h3031)
	) name6076 (
		_w3697_,
		_w7974_,
		_w7975_,
		_w7976_,
		_w7977_
	);
	LUT3 #(
		.INIT('h8a)
	) name6077 (
		\s1_msel_arb1_state_reg[2]/NET0131 ,
		_w7973_,
		_w7977_,
		_w7978_
	);
	LUT4 #(
		.INIT('h0100)
	) name6078 (
		_w3699_,
		_w3700_,
		_w3714_,
		_w4984_,
		_w7979_
	);
	LUT2 #(
		.INIT('h4)
	) name6079 (
		_w3709_,
		_w7979_,
		_w7980_
	);
	LUT4 #(
		.INIT('h000e)
	) name6080 (
		_w3696_,
		_w3697_,
		_w3699_,
		_w3700_,
		_w7981_
	);
	LUT3 #(
		.INIT('h10)
	) name6081 (
		_w3707_,
		_w3709_,
		_w4981_,
		_w7982_
	);
	LUT3 #(
		.INIT('hd0)
	) name6082 (
		_w3715_,
		_w7981_,
		_w7982_,
		_w7983_
	);
	LUT2 #(
		.INIT('h1)
	) name6083 (
		_w3704_,
		_w3711_,
		_w7984_
	);
	LUT3 #(
		.INIT('h8a)
	) name6084 (
		_w4984_,
		_w7981_,
		_w7984_,
		_w7985_
	);
	LUT2 #(
		.INIT('h4)
	) name6085 (
		_w3700_,
		_w5006_,
		_w7986_
	);
	LUT3 #(
		.INIT('hd0)
	) name6086 (
		_w3698_,
		_w7976_,
		_w7986_,
		_w7987_
	);
	LUT4 #(
		.INIT('h0001)
	) name6087 (
		_w7980_,
		_w7983_,
		_w7985_,
		_w7987_,
		_w7988_
	);
	LUT2 #(
		.INIT('hb)
	) name6088 (
		_w7978_,
		_w7988_,
		_w7989_
	);
	LUT4 #(
		.INIT('h000e)
	) name6089 (
		_w3727_,
		_w3728_,
		_w3730_,
		_w3731_,
		_w7990_
	);
	LUT3 #(
		.INIT('h02)
	) name6090 (
		\s2_msel_arb1_state_reg[2]/NET0131 ,
		_w3722_,
		_w3724_,
		_w7991_
	);
	LUT4 #(
		.INIT('h5100)
	) name6091 (
		\s2_msel_arb1_state_reg[0]/NET0131 ,
		_w3741_,
		_w7990_,
		_w7991_,
		_w7992_
	);
	LUT4 #(
		.INIT('h000e)
	) name6092 (
		_w3730_,
		_w3731_,
		_w3733_,
		_w3734_,
		_w7993_
	);
	LUT3 #(
		.INIT('h54)
	) name6093 (
		\s2_msel_arb1_state_reg[2]/NET0131 ,
		_w3727_,
		_w3728_,
		_w7994_
	);
	LUT4 #(
		.INIT('h0031)
	) name6094 (
		_w3740_,
		_w7990_,
		_w7993_,
		_w7994_,
		_w7995_
	);
	LUT2 #(
		.INIT('h4)
	) name6095 (
		\s2_msel_arb1_state_reg[0]/NET0131 ,
		\s2_msel_arb1_state_reg[1]/NET0131 ,
		_w7996_
	);
	LUT3 #(
		.INIT('h45)
	) name6096 (
		_w7992_,
		_w7995_,
		_w7996_,
		_w7997_
	);
	LUT4 #(
		.INIT('h000e)
	) name6097 (
		_w3722_,
		_w3724_,
		_w3727_,
		_w3728_,
		_w7998_
	);
	LUT3 #(
		.INIT('h02)
	) name6098 (
		\s2_msel_arb1_state_reg[0]/NET0131 ,
		_w3730_,
		_w3731_,
		_w7999_
	);
	LUT4 #(
		.INIT('hf700)
	) name6099 (
		\m7_s2_cyc_o_reg/NET0131 ,
		\rf_conf2_reg[14]/NET0131 ,
		\rf_conf2_reg[15]/NET0131 ,
		\s2_msel_arb1_state_reg[2]/NET0131 ,
		_w8000_
	);
	LUT2 #(
		.INIT('h4)
	) name6100 (
		_w5171_,
		_w8000_,
		_w8001_
	);
	LUT3 #(
		.INIT('hb0)
	) name6101 (
		_w7998_,
		_w7999_,
		_w8001_,
		_w8002_
	);
	LUT3 #(
		.INIT('h02)
	) name6102 (
		\s2_msel_arb1_state_reg[1]/NET0131 ,
		_w3722_,
		_w3724_,
		_w8003_
	);
	LUT4 #(
		.INIT('h0800)
	) name6103 (
		\m3_s2_cyc_o_reg/NET0131 ,
		\rf_conf2_reg[6]/NET0131 ,
		\rf_conf2_reg[7]/NET0131 ,
		\s2_msel_arb1_state_reg[0]/NET0131 ,
		_w8004_
	);
	LUT3 #(
		.INIT('ha8)
	) name6104 (
		\s2_msel_arb1_state_reg[1]/NET0131 ,
		\s2_msel_arb1_state_reg[2]/NET0131 ,
		_w8004_,
		_w8005_
	);
	LUT3 #(
		.INIT('h0b)
	) name6105 (
		_w7993_,
		_w8003_,
		_w8005_,
		_w8006_
	);
	LUT4 #(
		.INIT('h1110)
	) name6106 (
		_w3722_,
		_w3724_,
		_w3733_,
		_w3734_,
		_w8007_
	);
	LUT3 #(
		.INIT('h10)
	) name6107 (
		_w3730_,
		_w3738_,
		_w5160_,
		_w8008_
	);
	LUT3 #(
		.INIT('hd0)
	) name6108 (
		_w3729_,
		_w8007_,
		_w8008_,
		_w8009_
	);
	LUT3 #(
		.INIT('h20)
	) name6109 (
		\s2_msel_arb1_state_reg[0]/NET0131 ,
		\s2_msel_arb1_state_reg[1]/NET0131 ,
		\s2_msel_arb1_state_reg[2]/NET0131 ,
		_w8010_
	);
	LUT2 #(
		.INIT('h4)
	) name6110 (
		_w3722_,
		_w8010_,
		_w8011_
	);
	LUT3 #(
		.INIT('hd0)
	) name6111 (
		_w3741_,
		_w7990_,
		_w8011_,
		_w8012_
	);
	LUT4 #(
		.INIT('h000e)
	) name6112 (
		_w8002_,
		_w8006_,
		_w8009_,
		_w8012_,
		_w8013_
	);
	LUT2 #(
		.INIT('h7)
	) name6113 (
		_w7997_,
		_w8013_,
		_w8014_
	);
	LUT2 #(
		.INIT('h1)
	) name6114 (
		_w3759_,
		_w3765_,
		_w8015_
	);
	LUT2 #(
		.INIT('h1)
	) name6115 (
		_w3751_,
		_w8015_,
		_w8016_
	);
	LUT4 #(
		.INIT('h0001)
	) name6116 (
		_w3748_,
		_w3749_,
		_w3756_,
		_w3757_,
		_w8017_
	);
	LUT3 #(
		.INIT('h54)
	) name6117 (
		\s3_msel_arb1_state_reg[2]/NET0131 ,
		_w3756_,
		_w3757_,
		_w8018_
	);
	LUT3 #(
		.INIT('h32)
	) name6118 (
		_w3754_,
		_w8017_,
		_w8018_,
		_w8019_
	);
	LUT3 #(
		.INIT('h45)
	) name6119 (
		\s3_msel_arb1_state_reg[1]/NET0131 ,
		_w8016_,
		_w8019_,
		_w8020_
	);
	LUT4 #(
		.INIT('hf700)
	) name6120 (
		\m7_s3_cyc_o_reg/NET0131 ,
		\rf_conf3_reg[14]/NET0131 ,
		\rf_conf3_reg[15]/NET0131 ,
		\s3_msel_arb1_state_reg[1]/NET0131 ,
		_w8021_
	);
	LUT2 #(
		.INIT('h1)
	) name6121 (
		_w5336_,
		_w8021_,
		_w8022_
	);
	LUT4 #(
		.INIT('h000e)
	) name6122 (
		_w3752_,
		_w3753_,
		_w3756_,
		_w3757_,
		_w8023_
	);
	LUT3 #(
		.INIT('h01)
	) name6123 (
		_w3759_,
		_w3760_,
		_w5336_,
		_w8024_
	);
	LUT4 #(
		.INIT('h2022)
	) name6124 (
		\s3_msel_arb1_state_reg[0]/NET0131 ,
		_w8022_,
		_w8023_,
		_w8024_,
		_w8025_
	);
	LUT2 #(
		.INIT('h2)
	) name6125 (
		\s3_msel_arb1_state_reg[1]/NET0131 ,
		\s3_msel_arb1_state_reg[2]/NET0131 ,
		_w8026_
	);
	LUT2 #(
		.INIT('h4)
	) name6126 (
		_w3749_,
		_w8021_,
		_w8027_
	);
	LUT4 #(
		.INIT('h020f)
	) name6127 (
		_w3761_,
		_w8023_,
		_w8026_,
		_w8027_,
		_w8028_
	);
	LUT2 #(
		.INIT('h4)
	) name6128 (
		_w8025_,
		_w8028_,
		_w8029_
	);
	LUT4 #(
		.INIT('h1110)
	) name6129 (
		_w3748_,
		_w3749_,
		_w3759_,
		_w3760_,
		_w8030_
	);
	LUT2 #(
		.INIT('h4)
	) name6130 (
		_w3752_,
		_w8026_,
		_w8031_
	);
	LUT3 #(
		.INIT('h10)
	) name6131 (
		_w3753_,
		_w8030_,
		_w8031_,
		_w8032_
	);
	LUT4 #(
		.INIT('h000e)
	) name6132 (
		_w3756_,
		_w3757_,
		_w3759_,
		_w3760_,
		_w8033_
	);
	LUT2 #(
		.INIT('h4)
	) name6133 (
		_w3753_,
		_w5359_,
		_w8034_
	);
	LUT3 #(
		.INIT('hd0)
	) name6134 (
		_w3750_,
		_w8033_,
		_w8034_,
		_w8035_
	);
	LUT4 #(
		.INIT('h0800)
	) name6135 (
		\m3_s3_cyc_o_reg/NET0131 ,
		\rf_conf3_reg[6]/NET0131 ,
		\rf_conf3_reg[7]/NET0131 ,
		\s3_msel_arb1_state_reg[1]/NET0131 ,
		_w8036_
	);
	LUT2 #(
		.INIT('h1)
	) name6136 (
		_w3747_,
		_w8036_,
		_w8037_
	);
	LUT2 #(
		.INIT('h2)
	) name6137 (
		_w8018_,
		_w8037_,
		_w8038_
	);
	LUT3 #(
		.INIT('h01)
	) name6138 (
		_w8032_,
		_w8035_,
		_w8038_,
		_w8039_
	);
	LUT3 #(
		.INIT('h4f)
	) name6139 (
		_w8020_,
		_w8029_,
		_w8039_,
		_w8040_
	);
	LUT4 #(
		.INIT('h0001)
	) name6140 (
		_w3779_,
		_w3780_,
		_w3789_,
		_w3794_,
		_w8041_
	);
	LUT3 #(
		.INIT('ha8)
	) name6141 (
		\s4_msel_arb1_state_reg[1]/NET0131 ,
		_w5517_,
		_w8041_,
		_w8042_
	);
	LUT3 #(
		.INIT('h10)
	) name6142 (
		_w3779_,
		_w3780_,
		_w5517_,
		_w8043_
	);
	LUT4 #(
		.INIT('h3332)
	) name6143 (
		\s4_msel_arb1_state_reg[0]/NET0131 ,
		\s4_msel_arb1_state_reg[1]/NET0131 ,
		_w3779_,
		_w3780_,
		_w8044_
	);
	LUT4 #(
		.INIT('h000e)
	) name6144 (
		_w3784_,
		_w3788_,
		_w3789_,
		_w3794_,
		_w8045_
	);
	LUT4 #(
		.INIT('h3031)
	) name6145 (
		_w3777_,
		_w8043_,
		_w8044_,
		_w8045_,
		_w8046_
	);
	LUT3 #(
		.INIT('h8a)
	) name6146 (
		\s4_msel_arb1_state_reg[2]/NET0131 ,
		_w8042_,
		_w8046_,
		_w8047_
	);
	LUT4 #(
		.INIT('h0100)
	) name6147 (
		_w3779_,
		_w3780_,
		_w3794_,
		_w5502_,
		_w8048_
	);
	LUT2 #(
		.INIT('h4)
	) name6148 (
		_w3789_,
		_w8048_,
		_w8049_
	);
	LUT4 #(
		.INIT('h000e)
	) name6149 (
		_w3776_,
		_w3777_,
		_w3779_,
		_w3780_,
		_w8050_
	);
	LUT3 #(
		.INIT('h10)
	) name6150 (
		_w3787_,
		_w3789_,
		_w5499_,
		_w8051_
	);
	LUT3 #(
		.INIT('hd0)
	) name6151 (
		_w3795_,
		_w8050_,
		_w8051_,
		_w8052_
	);
	LUT2 #(
		.INIT('h1)
	) name6152 (
		_w3784_,
		_w3791_,
		_w8053_
	);
	LUT3 #(
		.INIT('h8a)
	) name6153 (
		_w5502_,
		_w8050_,
		_w8053_,
		_w8054_
	);
	LUT2 #(
		.INIT('h4)
	) name6154 (
		_w3780_,
		_w5524_,
		_w8055_
	);
	LUT3 #(
		.INIT('hd0)
	) name6155 (
		_w3778_,
		_w8045_,
		_w8055_,
		_w8056_
	);
	LUT4 #(
		.INIT('h0001)
	) name6156 (
		_w8049_,
		_w8052_,
		_w8054_,
		_w8056_,
		_w8057_
	);
	LUT2 #(
		.INIT('hb)
	) name6157 (
		_w8047_,
		_w8057_,
		_w8058_
	);
	LUT3 #(
		.INIT('h54)
	) name6158 (
		\s5_msel_arb1_state_reg[2]/NET0131 ,
		_w3811_,
		_w3812_,
		_w8059_
	);
	LUT4 #(
		.INIT('h000e)
	) name6159 (
		_w3805_,
		_w3806_,
		_w3808_,
		_w3809_,
		_w8060_
	);
	LUT3 #(
		.INIT('ha8)
	) name6160 (
		_w3824_,
		_w8059_,
		_w8060_,
		_w8061_
	);
	LUT3 #(
		.INIT('ha8)
	) name6161 (
		\s5_msel_arb1_state_reg[2]/NET0131 ,
		_w3805_,
		_w3806_,
		_w8062_
	);
	LUT4 #(
		.INIT('h1110)
	) name6162 (
		_w3802_,
		_w3803_,
		_w3811_,
		_w3812_,
		_w8063_
	);
	LUT2 #(
		.INIT('h1)
	) name6163 (
		_w3808_,
		_w5699_,
		_w8064_
	);
	LUT4 #(
		.INIT('h02aa)
	) name6164 (
		\s5_msel_arb1_state_reg[1]/NET0131 ,
		_w8062_,
		_w8063_,
		_w8064_,
		_w8065_
	);
	LUT4 #(
		.INIT('h000e)
	) name6165 (
		_w3808_,
		_w3809_,
		_w3811_,
		_w3812_,
		_w8066_
	);
	LUT3 #(
		.INIT('h04)
	) name6166 (
		_w3806_,
		_w3814_,
		_w5690_,
		_w8067_
	);
	LUT3 #(
		.INIT('hd0)
	) name6167 (
		_w3804_,
		_w8066_,
		_w8067_,
		_w8068_
	);
	LUT4 #(
		.INIT('h000e)
	) name6168 (
		_w3802_,
		_w3803_,
		_w3805_,
		_w3806_,
		_w8069_
	);
	LUT3 #(
		.INIT('h10)
	) name6169 (
		_w3812_,
		_w5675_,
		_w3818_,
		_w8070_
	);
	LUT3 #(
		.INIT('hd0)
	) name6170 (
		_w3810_,
		_w8069_,
		_w8070_,
		_w8071_
	);
	LUT4 #(
		.INIT('hfff4)
	) name6171 (
		_w8061_,
		_w8065_,
		_w8068_,
		_w8071_,
		_w8072_
	);
	LUT3 #(
		.INIT('h54)
	) name6172 (
		\s6_msel_arb1_state_reg[2]/NET0131 ,
		_w3842_,
		_w3843_,
		_w8073_
	);
	LUT4 #(
		.INIT('h000e)
	) name6173 (
		_w3836_,
		_w3837_,
		_w3839_,
		_w3840_,
		_w8074_
	);
	LUT3 #(
		.INIT('ha8)
	) name6174 (
		_w3855_,
		_w8073_,
		_w8074_,
		_w8075_
	);
	LUT3 #(
		.INIT('ha8)
	) name6175 (
		\s6_msel_arb1_state_reg[2]/NET0131 ,
		_w3836_,
		_w3837_,
		_w8076_
	);
	LUT4 #(
		.INIT('h1110)
	) name6176 (
		_w3833_,
		_w3834_,
		_w3842_,
		_w3843_,
		_w8077_
	);
	LUT2 #(
		.INIT('h1)
	) name6177 (
		_w3839_,
		_w5861_,
		_w8078_
	);
	LUT4 #(
		.INIT('h02aa)
	) name6178 (
		\s6_msel_arb1_state_reg[1]/NET0131 ,
		_w8076_,
		_w8077_,
		_w8078_,
		_w8079_
	);
	LUT4 #(
		.INIT('h000e)
	) name6179 (
		_w3839_,
		_w3840_,
		_w3842_,
		_w3843_,
		_w8080_
	);
	LUT3 #(
		.INIT('h04)
	) name6180 (
		_w3837_,
		_w3845_,
		_w5852_,
		_w8081_
	);
	LUT3 #(
		.INIT('hd0)
	) name6181 (
		_w3835_,
		_w8080_,
		_w8081_,
		_w8082_
	);
	LUT4 #(
		.INIT('h000e)
	) name6182 (
		_w3833_,
		_w3834_,
		_w3836_,
		_w3837_,
		_w8083_
	);
	LUT3 #(
		.INIT('h04)
	) name6183 (
		_w3843_,
		_w3849_,
		_w5837_,
		_w8084_
	);
	LUT3 #(
		.INIT('hd0)
	) name6184 (
		_w3841_,
		_w8083_,
		_w8084_,
		_w8085_
	);
	LUT4 #(
		.INIT('hfff4)
	) name6185 (
		_w8075_,
		_w8079_,
		_w8082_,
		_w8085_,
		_w8086_
	);
	LUT4 #(
		.INIT('h000e)
	) name6186 (
		_w3864_,
		_w3865_,
		_w3874_,
		_w3875_,
		_w8087_
	);
	LUT4 #(
		.INIT('h0008)
	) name6187 (
		\m2_s7_cyc_o_reg/NET0131 ,
		\rf_conf7_reg[4]/NET0131 ,
		\rf_conf7_reg[5]/NET0131 ,
		\s7_msel_arb1_state_reg[0]/NET0131 ,
		_w8088_
	);
	LUT2 #(
		.INIT('h2)
	) name6188 (
		_w5995_,
		_w8088_,
		_w8089_
	);
	LUT3 #(
		.INIT('hd0)
	) name6189 (
		_w3873_,
		_w8087_,
		_w8089_,
		_w8090_
	);
	LUT4 #(
		.INIT('h1110)
	) name6190 (
		_w3867_,
		_w3868_,
		_w3871_,
		_w3872_,
		_w8091_
	);
	LUT2 #(
		.INIT('h4)
	) name6191 (
		_w3879_,
		_w3882_,
		_w8092_
	);
	LUT3 #(
		.INIT('hd0)
	) name6192 (
		_w3866_,
		_w8091_,
		_w8092_,
		_w8093_
	);
	LUT3 #(
		.INIT('ha8)
	) name6193 (
		\s7_msel_arb1_state_reg[1]/NET0131 ,
		_w8090_,
		_w8093_,
		_w8094_
	);
	LUT4 #(
		.INIT('h1110)
	) name6194 (
		_w3871_,
		_w3872_,
		_w3874_,
		_w3875_,
		_w8095_
	);
	LUT3 #(
		.INIT('h01)
	) name6195 (
		\s7_msel_arb1_state_reg[2]/NET0131 ,
		_w3864_,
		_w3884_,
		_w8096_
	);
	LUT3 #(
		.INIT('hd0)
	) name6196 (
		_w3869_,
		_w8095_,
		_w8096_,
		_w8097_
	);
	LUT4 #(
		.INIT('h0008)
	) name6197 (
		\m4_s7_cyc_o_reg/NET0131 ,
		\rf_conf7_reg[8]/NET0131 ,
		\rf_conf7_reg[9]/NET0131 ,
		\s7_msel_arb1_state_reg[0]/NET0131 ,
		_w8098_
	);
	LUT4 #(
		.INIT('hf700)
	) name6198 (
		\m5_s7_cyc_o_reg/NET0131 ,
		\rf_conf7_reg[10]/NET0131 ,
		\rf_conf7_reg[11]/NET0131 ,
		\s7_msel_arb1_state_reg[2]/NET0131 ,
		_w8099_
	);
	LUT3 #(
		.INIT('h45)
	) name6199 (
		\s7_msel_arb1_state_reg[1]/NET0131 ,
		_w8098_,
		_w8099_,
		_w8100_
	);
	LUT4 #(
		.INIT('h1110)
	) name6200 (
		_w3864_,
		_w3865_,
		_w3867_,
		_w3868_,
		_w8101_
	);
	LUT3 #(
		.INIT('h01)
	) name6201 (
		\s7_msel_arb1_state_reg[1]/NET0131 ,
		_w3874_,
		_w3875_,
		_w8102_
	);
	LUT3 #(
		.INIT('h45)
	) name6202 (
		_w8100_,
		_w8101_,
		_w8102_,
		_w8103_
	);
	LUT2 #(
		.INIT('h1)
	) name6203 (
		_w8097_,
		_w8103_,
		_w8104_
	);
	LUT2 #(
		.INIT('h1)
	) name6204 (
		_w8094_,
		_w8104_,
		_w8105_
	);
	LUT3 #(
		.INIT('h54)
	) name6205 (
		\s8_msel_arb1_state_reg[2]/NET0131 ,
		_w3899_,
		_w3900_,
		_w8106_
	);
	LUT4 #(
		.INIT('h000e)
	) name6206 (
		_w3893_,
		_w3894_,
		_w3896_,
		_w3897_,
		_w8107_
	);
	LUT3 #(
		.INIT('ha8)
	) name6207 (
		_w3912_,
		_w8106_,
		_w8107_,
		_w8108_
	);
	LUT3 #(
		.INIT('ha8)
	) name6208 (
		\s8_msel_arb1_state_reg[2]/NET0131 ,
		_w3893_,
		_w3894_,
		_w8109_
	);
	LUT4 #(
		.INIT('h1110)
	) name6209 (
		_w3890_,
		_w3891_,
		_w3899_,
		_w3900_,
		_w8110_
	);
	LUT2 #(
		.INIT('h1)
	) name6210 (
		_w3896_,
		_w6207_,
		_w8111_
	);
	LUT4 #(
		.INIT('h02aa)
	) name6211 (
		\s8_msel_arb1_state_reg[1]/NET0131 ,
		_w8109_,
		_w8110_,
		_w8111_,
		_w8112_
	);
	LUT4 #(
		.INIT('h000e)
	) name6212 (
		_w3896_,
		_w3897_,
		_w3899_,
		_w3900_,
		_w8113_
	);
	LUT3 #(
		.INIT('h04)
	) name6213 (
		_w3894_,
		_w3902_,
		_w6198_,
		_w8114_
	);
	LUT3 #(
		.INIT('hd0)
	) name6214 (
		_w3892_,
		_w8113_,
		_w8114_,
		_w8115_
	);
	LUT4 #(
		.INIT('h000e)
	) name6215 (
		_w3890_,
		_w3891_,
		_w3893_,
		_w3894_,
		_w8116_
	);
	LUT3 #(
		.INIT('h04)
	) name6216 (
		_w3900_,
		_w3906_,
		_w6183_,
		_w8117_
	);
	LUT3 #(
		.INIT('hd0)
	) name6217 (
		_w3898_,
		_w8116_,
		_w8117_,
		_w8118_
	);
	LUT4 #(
		.INIT('hfff4)
	) name6218 (
		_w8108_,
		_w8112_,
		_w8115_,
		_w8118_,
		_w8119_
	);
	LUT3 #(
		.INIT('h54)
	) name6219 (
		\s9_msel_arb1_state_reg[2]/NET0131 ,
		_w3930_,
		_w3931_,
		_w8120_
	);
	LUT4 #(
		.INIT('h000e)
	) name6220 (
		_w3924_,
		_w3925_,
		_w3927_,
		_w3928_,
		_w8121_
	);
	LUT3 #(
		.INIT('ha8)
	) name6221 (
		_w3943_,
		_w8120_,
		_w8121_,
		_w8122_
	);
	LUT3 #(
		.INIT('ha8)
	) name6222 (
		\s9_msel_arb1_state_reg[2]/NET0131 ,
		_w3924_,
		_w3925_,
		_w8123_
	);
	LUT4 #(
		.INIT('h1110)
	) name6223 (
		_w3921_,
		_w3922_,
		_w3930_,
		_w3931_,
		_w8124_
	);
	LUT2 #(
		.INIT('h1)
	) name6224 (
		_w3927_,
		_w6361_,
		_w8125_
	);
	LUT4 #(
		.INIT('h02aa)
	) name6225 (
		\s9_msel_arb1_state_reg[1]/NET0131 ,
		_w8123_,
		_w8124_,
		_w8125_,
		_w8126_
	);
	LUT4 #(
		.INIT('h000e)
	) name6226 (
		_w3927_,
		_w3928_,
		_w3930_,
		_w3931_,
		_w8127_
	);
	LUT3 #(
		.INIT('h04)
	) name6227 (
		_w3925_,
		_w3933_,
		_w6352_,
		_w8128_
	);
	LUT3 #(
		.INIT('hd0)
	) name6228 (
		_w3923_,
		_w8127_,
		_w8128_,
		_w8129_
	);
	LUT4 #(
		.INIT('h000e)
	) name6229 (
		_w3921_,
		_w3922_,
		_w3924_,
		_w3925_,
		_w8130_
	);
	LUT3 #(
		.INIT('h04)
	) name6230 (
		_w3931_,
		_w3937_,
		_w6337_,
		_w8131_
	);
	LUT3 #(
		.INIT('hd0)
	) name6231 (
		_w3929_,
		_w8130_,
		_w8131_,
		_w8132_
	);
	LUT4 #(
		.INIT('hfff4)
	) name6232 (
		_w8122_,
		_w8126_,
		_w8129_,
		_w8132_,
		_w8133_
	);
	LUT3 #(
		.INIT('h54)
	) name6233 (
		\s0_msel_arb1_state_reg[2]/NET0131 ,
		_w3961_,
		_w3962_,
		_w8134_
	);
	LUT4 #(
		.INIT('h000e)
	) name6234 (
		_w3955_,
		_w3956_,
		_w3958_,
		_w3959_,
		_w8135_
	);
	LUT3 #(
		.INIT('ha8)
	) name6235 (
		_w3974_,
		_w8134_,
		_w8135_,
		_w8136_
	);
	LUT3 #(
		.INIT('ha8)
	) name6236 (
		\s0_msel_arb1_state_reg[2]/NET0131 ,
		_w3955_,
		_w3956_,
		_w8137_
	);
	LUT4 #(
		.INIT('h1110)
	) name6237 (
		_w3952_,
		_w3953_,
		_w3961_,
		_w3962_,
		_w8138_
	);
	LUT2 #(
		.INIT('h1)
	) name6238 (
		_w3958_,
		_w6534_,
		_w8139_
	);
	LUT4 #(
		.INIT('h02aa)
	) name6239 (
		\s0_msel_arb1_state_reg[1]/NET0131 ,
		_w8137_,
		_w8138_,
		_w8139_,
		_w8140_
	);
	LUT4 #(
		.INIT('h000e)
	) name6240 (
		_w3958_,
		_w3959_,
		_w3961_,
		_w3962_,
		_w8141_
	);
	LUT3 #(
		.INIT('h04)
	) name6241 (
		_w3956_,
		_w3964_,
		_w6525_,
		_w8142_
	);
	LUT3 #(
		.INIT('hd0)
	) name6242 (
		_w3954_,
		_w8141_,
		_w8142_,
		_w8143_
	);
	LUT4 #(
		.INIT('h000e)
	) name6243 (
		_w3952_,
		_w3953_,
		_w3955_,
		_w3956_,
		_w8144_
	);
	LUT3 #(
		.INIT('h04)
	) name6244 (
		_w3962_,
		_w3968_,
		_w6510_,
		_w8145_
	);
	LUT3 #(
		.INIT('hd0)
	) name6245 (
		_w3960_,
		_w8144_,
		_w8145_,
		_w8146_
	);
	LUT4 #(
		.INIT('hfff4)
	) name6246 (
		_w8136_,
		_w8140_,
		_w8143_,
		_w8146_,
		_w8147_
	);
	LUT3 #(
		.INIT('h54)
	) name6247 (
		rst_i_pad,
		\s15_msel_pri_out_reg[1]/NET0131 ,
		\s15_next_reg/P0001 ,
		_w8148_
	);
	LUT3 #(
		.INIT('h70)
	) name6248 (
		_w2904_,
		_w2917_,
		_w8148_,
		_w8149_
	);
	LUT3 #(
		.INIT('h2a)
	) name6249 (
		\m7_data_i[0]_pad ,
		_w1901_,
		_w1902_,
		_w8150_
	);
	LUT3 #(
		.INIT('h2a)
	) name6250 (
		\m6_data_i[0]_pad ,
		_w1908_,
		_w1909_,
		_w8151_
	);
	LUT4 #(
		.INIT('h153f)
	) name6251 (
		_w1907_,
		_w1918_,
		_w8150_,
		_w8151_,
		_w8152_
	);
	LUT3 #(
		.INIT('h2a)
	) name6252 (
		\m5_data_i[0]_pad ,
		_w1901_,
		_w1902_,
		_w8153_
	);
	LUT3 #(
		.INIT('h80)
	) name6253 (
		\m0_data_i[0]_pad ,
		_w1908_,
		_w1909_,
		_w8154_
	);
	LUT4 #(
		.INIT('h153f)
	) name6254 (
		_w1914_,
		_w1920_,
		_w8153_,
		_w8154_,
		_w8155_
	);
	LUT3 #(
		.INIT('h80)
	) name6255 (
		\m4_data_i[0]_pad ,
		_w1908_,
		_w1909_,
		_w8156_
	);
	LUT3 #(
		.INIT('h80)
	) name6256 (
		\m1_data_i[0]_pad ,
		_w1901_,
		_w1902_,
		_w8157_
	);
	LUT4 #(
		.INIT('h135f)
	) name6257 (
		_w1907_,
		_w1920_,
		_w8156_,
		_w8157_,
		_w8158_
	);
	LUT3 #(
		.INIT('h80)
	) name6258 (
		\m3_data_i[0]_pad ,
		_w1901_,
		_w1902_,
		_w8159_
	);
	LUT3 #(
		.INIT('h2a)
	) name6259 (
		\m2_data_i[0]_pad ,
		_w1908_,
		_w1909_,
		_w8160_
	);
	LUT4 #(
		.INIT('h153f)
	) name6260 (
		_w1914_,
		_w1918_,
		_w8159_,
		_w8160_,
		_w8161_
	);
	LUT4 #(
		.INIT('h8000)
	) name6261 (
		_w8152_,
		_w8155_,
		_w8158_,
		_w8161_,
		_w8162_
	);
	LUT4 #(
		.INIT('h7fff)
	) name6262 (
		_w8152_,
		_w8155_,
		_w8158_,
		_w8161_,
		_w8163_
	);
	LUT4 #(
		.INIT('h2aea)
	) name6263 (
		\rf_conf0_reg[0]/NET0131 ,
		\rf_rf_we_reg/P0001 ,
		_w1979_,
		_w8162_,
		_w8164_
	);
	LUT3 #(
		.INIT('h2a)
	) name6264 (
		\m7_data_i[10]_pad ,
		_w1901_,
		_w1902_,
		_w8165_
	);
	LUT3 #(
		.INIT('h2a)
	) name6265 (
		\m6_data_i[10]_pad ,
		_w1908_,
		_w1909_,
		_w8166_
	);
	LUT4 #(
		.INIT('h153f)
	) name6266 (
		_w1907_,
		_w1918_,
		_w8165_,
		_w8166_,
		_w8167_
	);
	LUT3 #(
		.INIT('h2a)
	) name6267 (
		\m5_data_i[10]_pad ,
		_w1901_,
		_w1902_,
		_w8168_
	);
	LUT3 #(
		.INIT('h2a)
	) name6268 (
		\m2_data_i[10]_pad ,
		_w1908_,
		_w1909_,
		_w8169_
	);
	LUT4 #(
		.INIT('h153f)
	) name6269 (
		_w1914_,
		_w1920_,
		_w8168_,
		_w8169_,
		_w8170_
	);
	LUT3 #(
		.INIT('h80)
	) name6270 (
		\m4_data_i[10]_pad ,
		_w1908_,
		_w1909_,
		_w8171_
	);
	LUT3 #(
		.INIT('h80)
	) name6271 (
		\m3_data_i[10]_pad ,
		_w1901_,
		_w1902_,
		_w8172_
	);
	LUT4 #(
		.INIT('h135f)
	) name6272 (
		_w1907_,
		_w1918_,
		_w8171_,
		_w8172_,
		_w8173_
	);
	LUT3 #(
		.INIT('h80)
	) name6273 (
		\m1_data_i[10]_pad ,
		_w1901_,
		_w1902_,
		_w8174_
	);
	LUT3 #(
		.INIT('h80)
	) name6274 (
		\m0_data_i[10]_pad ,
		_w1908_,
		_w1909_,
		_w8175_
	);
	LUT4 #(
		.INIT('h153f)
	) name6275 (
		_w1914_,
		_w1920_,
		_w8174_,
		_w8175_,
		_w8176_
	);
	LUT4 #(
		.INIT('h8000)
	) name6276 (
		_w8167_,
		_w8170_,
		_w8173_,
		_w8176_,
		_w8177_
	);
	LUT4 #(
		.INIT('h7fff)
	) name6277 (
		_w8167_,
		_w8170_,
		_w8173_,
		_w8176_,
		_w8178_
	);
	LUT4 #(
		.INIT('h2aea)
	) name6278 (
		\rf_conf0_reg[10]/NET0131 ,
		\rf_rf_we_reg/P0001 ,
		_w1979_,
		_w8177_,
		_w8179_
	);
	LUT3 #(
		.INIT('h2a)
	) name6279 (
		\m7_data_i[11]_pad ,
		_w1901_,
		_w1902_,
		_w8180_
	);
	LUT3 #(
		.INIT('h2a)
	) name6280 (
		\m6_data_i[11]_pad ,
		_w1908_,
		_w1909_,
		_w8181_
	);
	LUT4 #(
		.INIT('h153f)
	) name6281 (
		_w1907_,
		_w1918_,
		_w8180_,
		_w8181_,
		_w8182_
	);
	LUT3 #(
		.INIT('h2a)
	) name6282 (
		\m5_data_i[11]_pad ,
		_w1901_,
		_w1902_,
		_w8183_
	);
	LUT3 #(
		.INIT('h2a)
	) name6283 (
		\m2_data_i[11]_pad ,
		_w1908_,
		_w1909_,
		_w8184_
	);
	LUT4 #(
		.INIT('h153f)
	) name6284 (
		_w1914_,
		_w1920_,
		_w8183_,
		_w8184_,
		_w8185_
	);
	LUT3 #(
		.INIT('h80)
	) name6285 (
		\m4_data_i[11]_pad ,
		_w1908_,
		_w1909_,
		_w8186_
	);
	LUT3 #(
		.INIT('h80)
	) name6286 (
		\m3_data_i[11]_pad ,
		_w1901_,
		_w1902_,
		_w8187_
	);
	LUT4 #(
		.INIT('h135f)
	) name6287 (
		_w1907_,
		_w1918_,
		_w8186_,
		_w8187_,
		_w8188_
	);
	LUT3 #(
		.INIT('h80)
	) name6288 (
		\m1_data_i[11]_pad ,
		_w1901_,
		_w1902_,
		_w8189_
	);
	LUT3 #(
		.INIT('h80)
	) name6289 (
		\m0_data_i[11]_pad ,
		_w1908_,
		_w1909_,
		_w8190_
	);
	LUT4 #(
		.INIT('h153f)
	) name6290 (
		_w1914_,
		_w1920_,
		_w8189_,
		_w8190_,
		_w8191_
	);
	LUT4 #(
		.INIT('h8000)
	) name6291 (
		_w8182_,
		_w8185_,
		_w8188_,
		_w8191_,
		_w8192_
	);
	LUT4 #(
		.INIT('h7fff)
	) name6292 (
		_w8182_,
		_w8185_,
		_w8188_,
		_w8191_,
		_w8193_
	);
	LUT4 #(
		.INIT('h2aea)
	) name6293 (
		\rf_conf0_reg[11]/NET0131 ,
		\rf_rf_we_reg/P0001 ,
		_w1979_,
		_w8192_,
		_w8194_
	);
	LUT3 #(
		.INIT('h2a)
	) name6294 (
		\m7_data_i[12]_pad ,
		_w1901_,
		_w1902_,
		_w8195_
	);
	LUT3 #(
		.INIT('h2a)
	) name6295 (
		\m6_data_i[12]_pad ,
		_w1908_,
		_w1909_,
		_w8196_
	);
	LUT4 #(
		.INIT('h153f)
	) name6296 (
		_w1907_,
		_w1918_,
		_w8195_,
		_w8196_,
		_w8197_
	);
	LUT3 #(
		.INIT('h2a)
	) name6297 (
		\m5_data_i[12]_pad ,
		_w1901_,
		_w1902_,
		_w8198_
	);
	LUT3 #(
		.INIT('h2a)
	) name6298 (
		\m2_data_i[12]_pad ,
		_w1908_,
		_w1909_,
		_w8199_
	);
	LUT4 #(
		.INIT('h153f)
	) name6299 (
		_w1914_,
		_w1920_,
		_w8198_,
		_w8199_,
		_w8200_
	);
	LUT3 #(
		.INIT('h80)
	) name6300 (
		\m4_data_i[12]_pad ,
		_w1908_,
		_w1909_,
		_w8201_
	);
	LUT3 #(
		.INIT('h80)
	) name6301 (
		\m3_data_i[12]_pad ,
		_w1901_,
		_w1902_,
		_w8202_
	);
	LUT4 #(
		.INIT('h135f)
	) name6302 (
		_w1907_,
		_w1918_,
		_w8201_,
		_w8202_,
		_w8203_
	);
	LUT3 #(
		.INIT('h80)
	) name6303 (
		\m1_data_i[12]_pad ,
		_w1901_,
		_w1902_,
		_w8204_
	);
	LUT3 #(
		.INIT('h80)
	) name6304 (
		\m0_data_i[12]_pad ,
		_w1908_,
		_w1909_,
		_w8205_
	);
	LUT4 #(
		.INIT('h153f)
	) name6305 (
		_w1914_,
		_w1920_,
		_w8204_,
		_w8205_,
		_w8206_
	);
	LUT4 #(
		.INIT('h8000)
	) name6306 (
		_w8197_,
		_w8200_,
		_w8203_,
		_w8206_,
		_w8207_
	);
	LUT4 #(
		.INIT('h7fff)
	) name6307 (
		_w8197_,
		_w8200_,
		_w8203_,
		_w8206_,
		_w8208_
	);
	LUT4 #(
		.INIT('h2aea)
	) name6308 (
		\rf_conf0_reg[12]/NET0131 ,
		\rf_rf_we_reg/P0001 ,
		_w1979_,
		_w8207_,
		_w8209_
	);
	LUT3 #(
		.INIT('h2a)
	) name6309 (
		\m7_data_i[13]_pad ,
		_w1901_,
		_w1902_,
		_w8210_
	);
	LUT3 #(
		.INIT('h2a)
	) name6310 (
		\m6_data_i[13]_pad ,
		_w1908_,
		_w1909_,
		_w8211_
	);
	LUT4 #(
		.INIT('h153f)
	) name6311 (
		_w1907_,
		_w1918_,
		_w8210_,
		_w8211_,
		_w8212_
	);
	LUT3 #(
		.INIT('h2a)
	) name6312 (
		\m5_data_i[13]_pad ,
		_w1901_,
		_w1902_,
		_w8213_
	);
	LUT3 #(
		.INIT('h2a)
	) name6313 (
		\m2_data_i[13]_pad ,
		_w1908_,
		_w1909_,
		_w8214_
	);
	LUT4 #(
		.INIT('h153f)
	) name6314 (
		_w1914_,
		_w1920_,
		_w8213_,
		_w8214_,
		_w8215_
	);
	LUT3 #(
		.INIT('h80)
	) name6315 (
		\m4_data_i[13]_pad ,
		_w1908_,
		_w1909_,
		_w8216_
	);
	LUT3 #(
		.INIT('h80)
	) name6316 (
		\m3_data_i[13]_pad ,
		_w1901_,
		_w1902_,
		_w8217_
	);
	LUT4 #(
		.INIT('h135f)
	) name6317 (
		_w1907_,
		_w1918_,
		_w8216_,
		_w8217_,
		_w8218_
	);
	LUT3 #(
		.INIT('h80)
	) name6318 (
		\m1_data_i[13]_pad ,
		_w1901_,
		_w1902_,
		_w8219_
	);
	LUT3 #(
		.INIT('h80)
	) name6319 (
		\m0_data_i[13]_pad ,
		_w1908_,
		_w1909_,
		_w8220_
	);
	LUT4 #(
		.INIT('h153f)
	) name6320 (
		_w1914_,
		_w1920_,
		_w8219_,
		_w8220_,
		_w8221_
	);
	LUT4 #(
		.INIT('h8000)
	) name6321 (
		_w8212_,
		_w8215_,
		_w8218_,
		_w8221_,
		_w8222_
	);
	LUT4 #(
		.INIT('h7fff)
	) name6322 (
		_w8212_,
		_w8215_,
		_w8218_,
		_w8221_,
		_w8223_
	);
	LUT4 #(
		.INIT('h2aea)
	) name6323 (
		\rf_conf0_reg[13]/NET0131 ,
		\rf_rf_we_reg/P0001 ,
		_w1979_,
		_w8222_,
		_w8224_
	);
	LUT3 #(
		.INIT('h2a)
	) name6324 (
		\m7_data_i[14]_pad ,
		_w1901_,
		_w1902_,
		_w8225_
	);
	LUT3 #(
		.INIT('h2a)
	) name6325 (
		\m6_data_i[14]_pad ,
		_w1908_,
		_w1909_,
		_w8226_
	);
	LUT4 #(
		.INIT('h153f)
	) name6326 (
		_w1907_,
		_w1918_,
		_w8225_,
		_w8226_,
		_w8227_
	);
	LUT3 #(
		.INIT('h2a)
	) name6327 (
		\m5_data_i[14]_pad ,
		_w1901_,
		_w1902_,
		_w8228_
	);
	LUT3 #(
		.INIT('h2a)
	) name6328 (
		\m2_data_i[14]_pad ,
		_w1908_,
		_w1909_,
		_w8229_
	);
	LUT4 #(
		.INIT('h153f)
	) name6329 (
		_w1914_,
		_w1920_,
		_w8228_,
		_w8229_,
		_w8230_
	);
	LUT3 #(
		.INIT('h80)
	) name6330 (
		\m4_data_i[14]_pad ,
		_w1908_,
		_w1909_,
		_w8231_
	);
	LUT3 #(
		.INIT('h80)
	) name6331 (
		\m3_data_i[14]_pad ,
		_w1901_,
		_w1902_,
		_w8232_
	);
	LUT4 #(
		.INIT('h135f)
	) name6332 (
		_w1907_,
		_w1918_,
		_w8231_,
		_w8232_,
		_w8233_
	);
	LUT3 #(
		.INIT('h80)
	) name6333 (
		\m1_data_i[14]_pad ,
		_w1901_,
		_w1902_,
		_w8234_
	);
	LUT3 #(
		.INIT('h80)
	) name6334 (
		\m0_data_i[14]_pad ,
		_w1908_,
		_w1909_,
		_w8235_
	);
	LUT4 #(
		.INIT('h153f)
	) name6335 (
		_w1914_,
		_w1920_,
		_w8234_,
		_w8235_,
		_w8236_
	);
	LUT4 #(
		.INIT('h8000)
	) name6336 (
		_w8227_,
		_w8230_,
		_w8233_,
		_w8236_,
		_w8237_
	);
	LUT4 #(
		.INIT('h7fff)
	) name6337 (
		_w8227_,
		_w8230_,
		_w8233_,
		_w8236_,
		_w8238_
	);
	LUT4 #(
		.INIT('h2aea)
	) name6338 (
		\rf_conf0_reg[14]/NET0131 ,
		\rf_rf_we_reg/P0001 ,
		_w1979_,
		_w8237_,
		_w8239_
	);
	LUT3 #(
		.INIT('h2a)
	) name6339 (
		\m7_data_i[15]_pad ,
		_w1901_,
		_w1902_,
		_w8240_
	);
	LUT3 #(
		.INIT('h2a)
	) name6340 (
		\m6_data_i[15]_pad ,
		_w1908_,
		_w1909_,
		_w8241_
	);
	LUT4 #(
		.INIT('h153f)
	) name6341 (
		_w1907_,
		_w1918_,
		_w8240_,
		_w8241_,
		_w8242_
	);
	LUT3 #(
		.INIT('h2a)
	) name6342 (
		\m5_data_i[15]_pad ,
		_w1901_,
		_w1902_,
		_w8243_
	);
	LUT3 #(
		.INIT('h80)
	) name6343 (
		\m0_data_i[15]_pad ,
		_w1908_,
		_w1909_,
		_w8244_
	);
	LUT4 #(
		.INIT('h153f)
	) name6344 (
		_w1914_,
		_w1920_,
		_w8243_,
		_w8244_,
		_w8245_
	);
	LUT3 #(
		.INIT('h80)
	) name6345 (
		\m4_data_i[15]_pad ,
		_w1908_,
		_w1909_,
		_w8246_
	);
	LUT3 #(
		.INIT('h80)
	) name6346 (
		\m1_data_i[15]_pad ,
		_w1901_,
		_w1902_,
		_w8247_
	);
	LUT4 #(
		.INIT('h135f)
	) name6347 (
		_w1907_,
		_w1920_,
		_w8246_,
		_w8247_,
		_w8248_
	);
	LUT3 #(
		.INIT('h80)
	) name6348 (
		\m3_data_i[15]_pad ,
		_w1901_,
		_w1902_,
		_w8249_
	);
	LUT3 #(
		.INIT('h2a)
	) name6349 (
		\m2_data_i[15]_pad ,
		_w1908_,
		_w1909_,
		_w8250_
	);
	LUT4 #(
		.INIT('h153f)
	) name6350 (
		_w1914_,
		_w1918_,
		_w8249_,
		_w8250_,
		_w8251_
	);
	LUT4 #(
		.INIT('h8000)
	) name6351 (
		_w8242_,
		_w8245_,
		_w8248_,
		_w8251_,
		_w8252_
	);
	LUT4 #(
		.INIT('h7fff)
	) name6352 (
		_w8242_,
		_w8245_,
		_w8248_,
		_w8251_,
		_w8253_
	);
	LUT4 #(
		.INIT('h2aea)
	) name6353 (
		\rf_conf0_reg[15]/NET0131 ,
		\rf_rf_we_reg/P0001 ,
		_w1979_,
		_w8252_,
		_w8254_
	);
	LUT3 #(
		.INIT('h2a)
	) name6354 (
		\m7_data_i[1]_pad ,
		_w1901_,
		_w1902_,
		_w8255_
	);
	LUT3 #(
		.INIT('h2a)
	) name6355 (
		\m6_data_i[1]_pad ,
		_w1908_,
		_w1909_,
		_w8256_
	);
	LUT4 #(
		.INIT('h153f)
	) name6356 (
		_w1907_,
		_w1918_,
		_w8255_,
		_w8256_,
		_w8257_
	);
	LUT3 #(
		.INIT('h2a)
	) name6357 (
		\m5_data_i[1]_pad ,
		_w1901_,
		_w1902_,
		_w8258_
	);
	LUT3 #(
		.INIT('h80)
	) name6358 (
		\m0_data_i[1]_pad ,
		_w1908_,
		_w1909_,
		_w8259_
	);
	LUT4 #(
		.INIT('h153f)
	) name6359 (
		_w1914_,
		_w1920_,
		_w8258_,
		_w8259_,
		_w8260_
	);
	LUT3 #(
		.INIT('h80)
	) name6360 (
		\m4_data_i[1]_pad ,
		_w1908_,
		_w1909_,
		_w8261_
	);
	LUT3 #(
		.INIT('h80)
	) name6361 (
		\m1_data_i[1]_pad ,
		_w1901_,
		_w1902_,
		_w8262_
	);
	LUT4 #(
		.INIT('h135f)
	) name6362 (
		_w1907_,
		_w1920_,
		_w8261_,
		_w8262_,
		_w8263_
	);
	LUT3 #(
		.INIT('h80)
	) name6363 (
		\m3_data_i[1]_pad ,
		_w1901_,
		_w1902_,
		_w8264_
	);
	LUT3 #(
		.INIT('h2a)
	) name6364 (
		\m2_data_i[1]_pad ,
		_w1908_,
		_w1909_,
		_w8265_
	);
	LUT4 #(
		.INIT('h153f)
	) name6365 (
		_w1914_,
		_w1918_,
		_w8264_,
		_w8265_,
		_w8266_
	);
	LUT4 #(
		.INIT('h8000)
	) name6366 (
		_w8257_,
		_w8260_,
		_w8263_,
		_w8266_,
		_w8267_
	);
	LUT4 #(
		.INIT('h7fff)
	) name6367 (
		_w8257_,
		_w8260_,
		_w8263_,
		_w8266_,
		_w8268_
	);
	LUT4 #(
		.INIT('h2aea)
	) name6368 (
		\rf_conf0_reg[1]/NET0131 ,
		\rf_rf_we_reg/P0001 ,
		_w1979_,
		_w8267_,
		_w8269_
	);
	LUT3 #(
		.INIT('h2a)
	) name6369 (
		\m7_data_i[2]_pad ,
		_w1901_,
		_w1902_,
		_w8270_
	);
	LUT3 #(
		.INIT('h2a)
	) name6370 (
		\m6_data_i[2]_pad ,
		_w1908_,
		_w1909_,
		_w8271_
	);
	LUT4 #(
		.INIT('h153f)
	) name6371 (
		_w1907_,
		_w1918_,
		_w8270_,
		_w8271_,
		_w8272_
	);
	LUT3 #(
		.INIT('h2a)
	) name6372 (
		\m5_data_i[2]_pad ,
		_w1901_,
		_w1902_,
		_w8273_
	);
	LUT3 #(
		.INIT('h2a)
	) name6373 (
		\m2_data_i[2]_pad ,
		_w1908_,
		_w1909_,
		_w8274_
	);
	LUT4 #(
		.INIT('h153f)
	) name6374 (
		_w1914_,
		_w1920_,
		_w8273_,
		_w8274_,
		_w8275_
	);
	LUT3 #(
		.INIT('h80)
	) name6375 (
		\m4_data_i[2]_pad ,
		_w1908_,
		_w1909_,
		_w8276_
	);
	LUT3 #(
		.INIT('h80)
	) name6376 (
		\m3_data_i[2]_pad ,
		_w1901_,
		_w1902_,
		_w8277_
	);
	LUT4 #(
		.INIT('h135f)
	) name6377 (
		_w1907_,
		_w1918_,
		_w8276_,
		_w8277_,
		_w8278_
	);
	LUT3 #(
		.INIT('h80)
	) name6378 (
		\m1_data_i[2]_pad ,
		_w1901_,
		_w1902_,
		_w8279_
	);
	LUT3 #(
		.INIT('h80)
	) name6379 (
		\m0_data_i[2]_pad ,
		_w1908_,
		_w1909_,
		_w8280_
	);
	LUT4 #(
		.INIT('h153f)
	) name6380 (
		_w1914_,
		_w1920_,
		_w8279_,
		_w8280_,
		_w8281_
	);
	LUT4 #(
		.INIT('h8000)
	) name6381 (
		_w8272_,
		_w8275_,
		_w8278_,
		_w8281_,
		_w8282_
	);
	LUT4 #(
		.INIT('h7fff)
	) name6382 (
		_w8272_,
		_w8275_,
		_w8278_,
		_w8281_,
		_w8283_
	);
	LUT4 #(
		.INIT('h2aea)
	) name6383 (
		\rf_conf0_reg[2]/NET0131 ,
		\rf_rf_we_reg/P0001 ,
		_w1979_,
		_w8282_,
		_w8284_
	);
	LUT3 #(
		.INIT('h2a)
	) name6384 (
		\m7_data_i[3]_pad ,
		_w1901_,
		_w1902_,
		_w8285_
	);
	LUT3 #(
		.INIT('h2a)
	) name6385 (
		\m6_data_i[3]_pad ,
		_w1908_,
		_w1909_,
		_w8286_
	);
	LUT4 #(
		.INIT('h153f)
	) name6386 (
		_w1907_,
		_w1918_,
		_w8285_,
		_w8286_,
		_w8287_
	);
	LUT3 #(
		.INIT('h2a)
	) name6387 (
		\m5_data_i[3]_pad ,
		_w1901_,
		_w1902_,
		_w8288_
	);
	LUT3 #(
		.INIT('h2a)
	) name6388 (
		\m2_data_i[3]_pad ,
		_w1908_,
		_w1909_,
		_w8289_
	);
	LUT4 #(
		.INIT('h153f)
	) name6389 (
		_w1914_,
		_w1920_,
		_w8288_,
		_w8289_,
		_w8290_
	);
	LUT3 #(
		.INIT('h80)
	) name6390 (
		\m4_data_i[3]_pad ,
		_w1908_,
		_w1909_,
		_w8291_
	);
	LUT3 #(
		.INIT('h80)
	) name6391 (
		\m3_data_i[3]_pad ,
		_w1901_,
		_w1902_,
		_w8292_
	);
	LUT4 #(
		.INIT('h135f)
	) name6392 (
		_w1907_,
		_w1918_,
		_w8291_,
		_w8292_,
		_w8293_
	);
	LUT3 #(
		.INIT('h80)
	) name6393 (
		\m1_data_i[3]_pad ,
		_w1901_,
		_w1902_,
		_w8294_
	);
	LUT3 #(
		.INIT('h80)
	) name6394 (
		\m0_data_i[3]_pad ,
		_w1908_,
		_w1909_,
		_w8295_
	);
	LUT4 #(
		.INIT('h153f)
	) name6395 (
		_w1914_,
		_w1920_,
		_w8294_,
		_w8295_,
		_w8296_
	);
	LUT4 #(
		.INIT('h8000)
	) name6396 (
		_w8287_,
		_w8290_,
		_w8293_,
		_w8296_,
		_w8297_
	);
	LUT4 #(
		.INIT('h7fff)
	) name6397 (
		_w8287_,
		_w8290_,
		_w8293_,
		_w8296_,
		_w8298_
	);
	LUT4 #(
		.INIT('h2aea)
	) name6398 (
		\rf_conf0_reg[3]/NET0131 ,
		\rf_rf_we_reg/P0001 ,
		_w1979_,
		_w8297_,
		_w8299_
	);
	LUT3 #(
		.INIT('h2a)
	) name6399 (
		\m7_data_i[4]_pad ,
		_w1901_,
		_w1902_,
		_w8300_
	);
	LUT3 #(
		.INIT('h2a)
	) name6400 (
		\m6_data_i[4]_pad ,
		_w1908_,
		_w1909_,
		_w8301_
	);
	LUT4 #(
		.INIT('h153f)
	) name6401 (
		_w1907_,
		_w1918_,
		_w8300_,
		_w8301_,
		_w8302_
	);
	LUT3 #(
		.INIT('h2a)
	) name6402 (
		\m5_data_i[4]_pad ,
		_w1901_,
		_w1902_,
		_w8303_
	);
	LUT3 #(
		.INIT('h2a)
	) name6403 (
		\m2_data_i[4]_pad ,
		_w1908_,
		_w1909_,
		_w8304_
	);
	LUT4 #(
		.INIT('h153f)
	) name6404 (
		_w1914_,
		_w1920_,
		_w8303_,
		_w8304_,
		_w8305_
	);
	LUT3 #(
		.INIT('h80)
	) name6405 (
		\m4_data_i[4]_pad ,
		_w1908_,
		_w1909_,
		_w8306_
	);
	LUT3 #(
		.INIT('h80)
	) name6406 (
		\m3_data_i[4]_pad ,
		_w1901_,
		_w1902_,
		_w8307_
	);
	LUT4 #(
		.INIT('h135f)
	) name6407 (
		_w1907_,
		_w1918_,
		_w8306_,
		_w8307_,
		_w8308_
	);
	LUT3 #(
		.INIT('h80)
	) name6408 (
		\m1_data_i[4]_pad ,
		_w1901_,
		_w1902_,
		_w8309_
	);
	LUT3 #(
		.INIT('h80)
	) name6409 (
		\m0_data_i[4]_pad ,
		_w1908_,
		_w1909_,
		_w8310_
	);
	LUT4 #(
		.INIT('h153f)
	) name6410 (
		_w1914_,
		_w1920_,
		_w8309_,
		_w8310_,
		_w8311_
	);
	LUT4 #(
		.INIT('h8000)
	) name6411 (
		_w8302_,
		_w8305_,
		_w8308_,
		_w8311_,
		_w8312_
	);
	LUT4 #(
		.INIT('h7fff)
	) name6412 (
		_w8302_,
		_w8305_,
		_w8308_,
		_w8311_,
		_w8313_
	);
	LUT4 #(
		.INIT('h2aea)
	) name6413 (
		\rf_conf0_reg[4]/NET0131 ,
		\rf_rf_we_reg/P0001 ,
		_w1979_,
		_w8312_,
		_w8314_
	);
	LUT3 #(
		.INIT('h80)
	) name6414 (
		\m3_data_i[5]_pad ,
		_w1901_,
		_w1902_,
		_w8315_
	);
	LUT3 #(
		.INIT('h2a)
	) name6415 (
		\m2_data_i[5]_pad ,
		_w1908_,
		_w1909_,
		_w8316_
	);
	LUT4 #(
		.INIT('h153f)
	) name6416 (
		_w1914_,
		_w1918_,
		_w8315_,
		_w8316_,
		_w8317_
	);
	LUT3 #(
		.INIT('h2a)
	) name6417 (
		\m5_data_i[5]_pad ,
		_w1901_,
		_w1902_,
		_w8318_
	);
	LUT3 #(
		.INIT('h80)
	) name6418 (
		\m0_data_i[5]_pad ,
		_w1908_,
		_w1909_,
		_w8319_
	);
	LUT4 #(
		.INIT('h153f)
	) name6419 (
		_w1914_,
		_w1920_,
		_w8318_,
		_w8319_,
		_w8320_
	);
	LUT3 #(
		.INIT('h80)
	) name6420 (
		\m4_data_i[5]_pad ,
		_w1908_,
		_w1909_,
		_w8321_
	);
	LUT3 #(
		.INIT('h80)
	) name6421 (
		\m1_data_i[5]_pad ,
		_w1901_,
		_w1902_,
		_w8322_
	);
	LUT4 #(
		.INIT('h135f)
	) name6422 (
		_w1907_,
		_w1920_,
		_w8321_,
		_w8322_,
		_w8323_
	);
	LUT3 #(
		.INIT('h2a)
	) name6423 (
		\m7_data_i[5]_pad ,
		_w1901_,
		_w1902_,
		_w8324_
	);
	LUT3 #(
		.INIT('h2a)
	) name6424 (
		\m6_data_i[5]_pad ,
		_w1908_,
		_w1909_,
		_w8325_
	);
	LUT4 #(
		.INIT('h153f)
	) name6425 (
		_w1907_,
		_w1918_,
		_w8324_,
		_w8325_,
		_w8326_
	);
	LUT4 #(
		.INIT('h8000)
	) name6426 (
		_w8317_,
		_w8320_,
		_w8323_,
		_w8326_,
		_w8327_
	);
	LUT4 #(
		.INIT('h7fff)
	) name6427 (
		_w8317_,
		_w8320_,
		_w8323_,
		_w8326_,
		_w8328_
	);
	LUT4 #(
		.INIT('h2aea)
	) name6428 (
		\rf_conf0_reg[5]/NET0131 ,
		\rf_rf_we_reg/P0001 ,
		_w1979_,
		_w8327_,
		_w8329_
	);
	LUT3 #(
		.INIT('h2a)
	) name6429 (
		\m7_data_i[6]_pad ,
		_w1901_,
		_w1902_,
		_w8330_
	);
	LUT3 #(
		.INIT('h2a)
	) name6430 (
		\m6_data_i[6]_pad ,
		_w1908_,
		_w1909_,
		_w8331_
	);
	LUT4 #(
		.INIT('h153f)
	) name6431 (
		_w1907_,
		_w1918_,
		_w8330_,
		_w8331_,
		_w8332_
	);
	LUT3 #(
		.INIT('h2a)
	) name6432 (
		\m5_data_i[6]_pad ,
		_w1901_,
		_w1902_,
		_w8333_
	);
	LUT3 #(
		.INIT('h2a)
	) name6433 (
		\m2_data_i[6]_pad ,
		_w1908_,
		_w1909_,
		_w8334_
	);
	LUT4 #(
		.INIT('h153f)
	) name6434 (
		_w1914_,
		_w1920_,
		_w8333_,
		_w8334_,
		_w8335_
	);
	LUT3 #(
		.INIT('h80)
	) name6435 (
		\m4_data_i[6]_pad ,
		_w1908_,
		_w1909_,
		_w8336_
	);
	LUT3 #(
		.INIT('h80)
	) name6436 (
		\m3_data_i[6]_pad ,
		_w1901_,
		_w1902_,
		_w8337_
	);
	LUT4 #(
		.INIT('h135f)
	) name6437 (
		_w1907_,
		_w1918_,
		_w8336_,
		_w8337_,
		_w8338_
	);
	LUT3 #(
		.INIT('h80)
	) name6438 (
		\m1_data_i[6]_pad ,
		_w1901_,
		_w1902_,
		_w8339_
	);
	LUT3 #(
		.INIT('h80)
	) name6439 (
		\m0_data_i[6]_pad ,
		_w1908_,
		_w1909_,
		_w8340_
	);
	LUT4 #(
		.INIT('h153f)
	) name6440 (
		_w1914_,
		_w1920_,
		_w8339_,
		_w8340_,
		_w8341_
	);
	LUT4 #(
		.INIT('h8000)
	) name6441 (
		_w8332_,
		_w8335_,
		_w8338_,
		_w8341_,
		_w8342_
	);
	LUT4 #(
		.INIT('h7fff)
	) name6442 (
		_w8332_,
		_w8335_,
		_w8338_,
		_w8341_,
		_w8343_
	);
	LUT4 #(
		.INIT('h2aea)
	) name6443 (
		\rf_conf0_reg[6]/NET0131 ,
		\rf_rf_we_reg/P0001 ,
		_w1979_,
		_w8342_,
		_w8344_
	);
	LUT3 #(
		.INIT('h2a)
	) name6444 (
		\m7_data_i[7]_pad ,
		_w1901_,
		_w1902_,
		_w8345_
	);
	LUT3 #(
		.INIT('h2a)
	) name6445 (
		\m6_data_i[7]_pad ,
		_w1908_,
		_w1909_,
		_w8346_
	);
	LUT4 #(
		.INIT('h153f)
	) name6446 (
		_w1907_,
		_w1918_,
		_w8345_,
		_w8346_,
		_w8347_
	);
	LUT3 #(
		.INIT('h2a)
	) name6447 (
		\m5_data_i[7]_pad ,
		_w1901_,
		_w1902_,
		_w8348_
	);
	LUT3 #(
		.INIT('h2a)
	) name6448 (
		\m2_data_i[7]_pad ,
		_w1908_,
		_w1909_,
		_w8349_
	);
	LUT4 #(
		.INIT('h153f)
	) name6449 (
		_w1914_,
		_w1920_,
		_w8348_,
		_w8349_,
		_w8350_
	);
	LUT3 #(
		.INIT('h80)
	) name6450 (
		\m4_data_i[7]_pad ,
		_w1908_,
		_w1909_,
		_w8351_
	);
	LUT3 #(
		.INIT('h80)
	) name6451 (
		\m3_data_i[7]_pad ,
		_w1901_,
		_w1902_,
		_w8352_
	);
	LUT4 #(
		.INIT('h135f)
	) name6452 (
		_w1907_,
		_w1918_,
		_w8351_,
		_w8352_,
		_w8353_
	);
	LUT3 #(
		.INIT('h80)
	) name6453 (
		\m1_data_i[7]_pad ,
		_w1901_,
		_w1902_,
		_w8354_
	);
	LUT3 #(
		.INIT('h80)
	) name6454 (
		\m0_data_i[7]_pad ,
		_w1908_,
		_w1909_,
		_w8355_
	);
	LUT4 #(
		.INIT('h153f)
	) name6455 (
		_w1914_,
		_w1920_,
		_w8354_,
		_w8355_,
		_w8356_
	);
	LUT4 #(
		.INIT('h8000)
	) name6456 (
		_w8347_,
		_w8350_,
		_w8353_,
		_w8356_,
		_w8357_
	);
	LUT4 #(
		.INIT('h7fff)
	) name6457 (
		_w8347_,
		_w8350_,
		_w8353_,
		_w8356_,
		_w8358_
	);
	LUT4 #(
		.INIT('h2aea)
	) name6458 (
		\rf_conf0_reg[7]/NET0131 ,
		\rf_rf_we_reg/P0001 ,
		_w1979_,
		_w8357_,
		_w8359_
	);
	LUT3 #(
		.INIT('h2a)
	) name6459 (
		\m7_data_i[8]_pad ,
		_w1901_,
		_w1902_,
		_w8360_
	);
	LUT3 #(
		.INIT('h2a)
	) name6460 (
		\m6_data_i[8]_pad ,
		_w1908_,
		_w1909_,
		_w8361_
	);
	LUT4 #(
		.INIT('h153f)
	) name6461 (
		_w1907_,
		_w1918_,
		_w8360_,
		_w8361_,
		_w8362_
	);
	LUT3 #(
		.INIT('h2a)
	) name6462 (
		\m5_data_i[8]_pad ,
		_w1901_,
		_w1902_,
		_w8363_
	);
	LUT3 #(
		.INIT('h80)
	) name6463 (
		\m0_data_i[8]_pad ,
		_w1908_,
		_w1909_,
		_w8364_
	);
	LUT4 #(
		.INIT('h153f)
	) name6464 (
		_w1914_,
		_w1920_,
		_w8363_,
		_w8364_,
		_w8365_
	);
	LUT3 #(
		.INIT('h80)
	) name6465 (
		\m4_data_i[8]_pad ,
		_w1908_,
		_w1909_,
		_w8366_
	);
	LUT3 #(
		.INIT('h80)
	) name6466 (
		\m1_data_i[8]_pad ,
		_w1901_,
		_w1902_,
		_w8367_
	);
	LUT4 #(
		.INIT('h135f)
	) name6467 (
		_w1907_,
		_w1920_,
		_w8366_,
		_w8367_,
		_w8368_
	);
	LUT3 #(
		.INIT('h80)
	) name6468 (
		\m3_data_i[8]_pad ,
		_w1901_,
		_w1902_,
		_w8369_
	);
	LUT3 #(
		.INIT('h2a)
	) name6469 (
		\m2_data_i[8]_pad ,
		_w1908_,
		_w1909_,
		_w8370_
	);
	LUT4 #(
		.INIT('h153f)
	) name6470 (
		_w1914_,
		_w1918_,
		_w8369_,
		_w8370_,
		_w8371_
	);
	LUT4 #(
		.INIT('h8000)
	) name6471 (
		_w8362_,
		_w8365_,
		_w8368_,
		_w8371_,
		_w8372_
	);
	LUT4 #(
		.INIT('h7fff)
	) name6472 (
		_w8362_,
		_w8365_,
		_w8368_,
		_w8371_,
		_w8373_
	);
	LUT4 #(
		.INIT('h2aea)
	) name6473 (
		\rf_conf0_reg[8]/NET0131 ,
		\rf_rf_we_reg/P0001 ,
		_w1979_,
		_w8372_,
		_w8374_
	);
	LUT3 #(
		.INIT('h2a)
	) name6474 (
		\m5_data_i[9]_pad ,
		_w1901_,
		_w1902_,
		_w8375_
	);
	LUT3 #(
		.INIT('h80)
	) name6475 (
		\m4_data_i[9]_pad ,
		_w1908_,
		_w1909_,
		_w8376_
	);
	LUT4 #(
		.INIT('h153f)
	) name6476 (
		_w1907_,
		_w1920_,
		_w8375_,
		_w8376_,
		_w8377_
	);
	LUT3 #(
		.INIT('h2a)
	) name6477 (
		\m7_data_i[9]_pad ,
		_w1901_,
		_w1902_,
		_w8378_
	);
	LUT3 #(
		.INIT('h80)
	) name6478 (
		\m0_data_i[9]_pad ,
		_w1908_,
		_w1909_,
		_w8379_
	);
	LUT4 #(
		.INIT('h153f)
	) name6479 (
		_w1914_,
		_w1918_,
		_w8378_,
		_w8379_,
		_w8380_
	);
	LUT3 #(
		.INIT('h2a)
	) name6480 (
		\m6_data_i[9]_pad ,
		_w1908_,
		_w1909_,
		_w8381_
	);
	LUT3 #(
		.INIT('h80)
	) name6481 (
		\m1_data_i[9]_pad ,
		_w1901_,
		_w1902_,
		_w8382_
	);
	LUT4 #(
		.INIT('h135f)
	) name6482 (
		_w1907_,
		_w1920_,
		_w8381_,
		_w8382_,
		_w8383_
	);
	LUT3 #(
		.INIT('h80)
	) name6483 (
		\m3_data_i[9]_pad ,
		_w1901_,
		_w1902_,
		_w8384_
	);
	LUT3 #(
		.INIT('h2a)
	) name6484 (
		\m2_data_i[9]_pad ,
		_w1908_,
		_w1909_,
		_w8385_
	);
	LUT4 #(
		.INIT('h153f)
	) name6485 (
		_w1914_,
		_w1918_,
		_w8384_,
		_w8385_,
		_w8386_
	);
	LUT4 #(
		.INIT('h8000)
	) name6486 (
		_w8377_,
		_w8380_,
		_w8383_,
		_w8386_,
		_w8387_
	);
	LUT4 #(
		.INIT('h7fff)
	) name6487 (
		_w8377_,
		_w8380_,
		_w8383_,
		_w8386_,
		_w8388_
	);
	LUT4 #(
		.INIT('h2aea)
	) name6488 (
		\rf_conf0_reg[9]/NET0131 ,
		\rf_rf_we_reg/P0001 ,
		_w1979_,
		_w8387_,
		_w8389_
	);
	LUT4 #(
		.INIT('h2aea)
	) name6489 (
		\rf_conf10_reg[0]/NET0131 ,
		\rf_rf_we_reg/P0001 ,
		_w1990_,
		_w8162_,
		_w8390_
	);
	LUT4 #(
		.INIT('h2aea)
	) name6490 (
		\rf_conf10_reg[10]/NET0131 ,
		\rf_rf_we_reg/P0001 ,
		_w1990_,
		_w8177_,
		_w8391_
	);
	LUT4 #(
		.INIT('h2aea)
	) name6491 (
		\rf_conf10_reg[11]/NET0131 ,
		\rf_rf_we_reg/P0001 ,
		_w1990_,
		_w8192_,
		_w8392_
	);
	LUT4 #(
		.INIT('h2aea)
	) name6492 (
		\rf_conf10_reg[12]/NET0131 ,
		\rf_rf_we_reg/P0001 ,
		_w1990_,
		_w8207_,
		_w8393_
	);
	LUT4 #(
		.INIT('h2aea)
	) name6493 (
		\rf_conf10_reg[13]/NET0131 ,
		\rf_rf_we_reg/P0001 ,
		_w1990_,
		_w8222_,
		_w8394_
	);
	LUT4 #(
		.INIT('h2aea)
	) name6494 (
		\rf_conf10_reg[15]/NET0131 ,
		\rf_rf_we_reg/P0001 ,
		_w1990_,
		_w8252_,
		_w8395_
	);
	LUT4 #(
		.INIT('h2aea)
	) name6495 (
		\rf_conf10_reg[1]/NET0131 ,
		\rf_rf_we_reg/P0001 ,
		_w1990_,
		_w8267_,
		_w8396_
	);
	LUT4 #(
		.INIT('h2aea)
	) name6496 (
		\rf_conf10_reg[14]/NET0131 ,
		\rf_rf_we_reg/P0001 ,
		_w1990_,
		_w8237_,
		_w8397_
	);
	LUT4 #(
		.INIT('h2aea)
	) name6497 (
		\rf_conf10_reg[2]/NET0131 ,
		\rf_rf_we_reg/P0001 ,
		_w1990_,
		_w8282_,
		_w8398_
	);
	LUT4 #(
		.INIT('h2aea)
	) name6498 (
		\rf_conf10_reg[3]/NET0131 ,
		\rf_rf_we_reg/P0001 ,
		_w1990_,
		_w8297_,
		_w8399_
	);
	LUT4 #(
		.INIT('h2aea)
	) name6499 (
		\rf_conf10_reg[4]/NET0131 ,
		\rf_rf_we_reg/P0001 ,
		_w1990_,
		_w8312_,
		_w8400_
	);
	LUT4 #(
		.INIT('h2aea)
	) name6500 (
		\rf_conf10_reg[5]/NET0131 ,
		\rf_rf_we_reg/P0001 ,
		_w1990_,
		_w8327_,
		_w8401_
	);
	LUT4 #(
		.INIT('h2aea)
	) name6501 (
		\rf_conf10_reg[6]/NET0131 ,
		\rf_rf_we_reg/P0001 ,
		_w1990_,
		_w8342_,
		_w8402_
	);
	LUT4 #(
		.INIT('h2aea)
	) name6502 (
		\rf_conf10_reg[7]/NET0131 ,
		\rf_rf_we_reg/P0001 ,
		_w1990_,
		_w8357_,
		_w8403_
	);
	LUT4 #(
		.INIT('h2aea)
	) name6503 (
		\rf_conf10_reg[8]/NET0131 ,
		\rf_rf_we_reg/P0001 ,
		_w1990_,
		_w8372_,
		_w8404_
	);
	LUT4 #(
		.INIT('h2aea)
	) name6504 (
		\rf_conf10_reg[9]/NET0131 ,
		\rf_rf_we_reg/P0001 ,
		_w1990_,
		_w8387_,
		_w8405_
	);
	LUT4 #(
		.INIT('h2aea)
	) name6505 (
		\rf_conf11_reg[0]/NET0131 ,
		\rf_rf_we_reg/P0001 ,
		_w1987_,
		_w8162_,
		_w8406_
	);
	LUT4 #(
		.INIT('h2aea)
	) name6506 (
		\rf_conf11_reg[10]/NET0131 ,
		\rf_rf_we_reg/P0001 ,
		_w1987_,
		_w8177_,
		_w8407_
	);
	LUT4 #(
		.INIT('h2aea)
	) name6507 (
		\rf_conf11_reg[12]/NET0131 ,
		\rf_rf_we_reg/P0001 ,
		_w1987_,
		_w8207_,
		_w8408_
	);
	LUT4 #(
		.INIT('h2aea)
	) name6508 (
		\rf_conf11_reg[11]/NET0131 ,
		\rf_rf_we_reg/P0001 ,
		_w1987_,
		_w8192_,
		_w8409_
	);
	LUT4 #(
		.INIT('h2aea)
	) name6509 (
		\rf_conf11_reg[13]/NET0131 ,
		\rf_rf_we_reg/P0001 ,
		_w1987_,
		_w8222_,
		_w8410_
	);
	LUT4 #(
		.INIT('h2aea)
	) name6510 (
		\rf_conf11_reg[14]/NET0131 ,
		\rf_rf_we_reg/P0001 ,
		_w1987_,
		_w8237_,
		_w8411_
	);
	LUT4 #(
		.INIT('h2aea)
	) name6511 (
		\rf_conf11_reg[15]/NET0131 ,
		\rf_rf_we_reg/P0001 ,
		_w1987_,
		_w8252_,
		_w8412_
	);
	LUT4 #(
		.INIT('h2aea)
	) name6512 (
		\rf_conf11_reg[1]/NET0131 ,
		\rf_rf_we_reg/P0001 ,
		_w1987_,
		_w8267_,
		_w8413_
	);
	LUT4 #(
		.INIT('h2aea)
	) name6513 (
		\rf_conf11_reg[2]/NET0131 ,
		\rf_rf_we_reg/P0001 ,
		_w1987_,
		_w8282_,
		_w8414_
	);
	LUT4 #(
		.INIT('h2aea)
	) name6514 (
		\rf_conf11_reg[3]/NET0131 ,
		\rf_rf_we_reg/P0001 ,
		_w1987_,
		_w8297_,
		_w8415_
	);
	LUT4 #(
		.INIT('h2aea)
	) name6515 (
		\rf_conf11_reg[4]/NET0131 ,
		\rf_rf_we_reg/P0001 ,
		_w1987_,
		_w8312_,
		_w8416_
	);
	LUT4 #(
		.INIT('h2aea)
	) name6516 (
		\rf_conf11_reg[5]/NET0131 ,
		\rf_rf_we_reg/P0001 ,
		_w1987_,
		_w8327_,
		_w8417_
	);
	LUT4 #(
		.INIT('h2aea)
	) name6517 (
		\rf_conf11_reg[6]/NET0131 ,
		\rf_rf_we_reg/P0001 ,
		_w1987_,
		_w8342_,
		_w8418_
	);
	LUT4 #(
		.INIT('h2aea)
	) name6518 (
		\rf_conf11_reg[7]/NET0131 ,
		\rf_rf_we_reg/P0001 ,
		_w1987_,
		_w8357_,
		_w8419_
	);
	LUT4 #(
		.INIT('h2aea)
	) name6519 (
		\rf_conf11_reg[8]/NET0131 ,
		\rf_rf_we_reg/P0001 ,
		_w1987_,
		_w8372_,
		_w8420_
	);
	LUT4 #(
		.INIT('h2aea)
	) name6520 (
		\rf_conf11_reg[9]/NET0131 ,
		\rf_rf_we_reg/P0001 ,
		_w1987_,
		_w8387_,
		_w8421_
	);
	LUT4 #(
		.INIT('h2aea)
	) name6521 (
		\rf_conf12_reg[0]/NET0131 ,
		\rf_rf_we_reg/P0001 ,
		_w1973_,
		_w8162_,
		_w8422_
	);
	LUT4 #(
		.INIT('h2aea)
	) name6522 (
		\rf_conf12_reg[10]/NET0131 ,
		\rf_rf_we_reg/P0001 ,
		_w1973_,
		_w8177_,
		_w8423_
	);
	LUT4 #(
		.INIT('h2aea)
	) name6523 (
		\rf_conf12_reg[11]/NET0131 ,
		\rf_rf_we_reg/P0001 ,
		_w1973_,
		_w8192_,
		_w8424_
	);
	LUT4 #(
		.INIT('h2aea)
	) name6524 (
		\rf_conf12_reg[12]/NET0131 ,
		\rf_rf_we_reg/P0001 ,
		_w1973_,
		_w8207_,
		_w8425_
	);
	LUT4 #(
		.INIT('h2aea)
	) name6525 (
		\rf_conf12_reg[13]/NET0131 ,
		\rf_rf_we_reg/P0001 ,
		_w1973_,
		_w8222_,
		_w8426_
	);
	LUT4 #(
		.INIT('h2aea)
	) name6526 (
		\rf_conf12_reg[14]/NET0131 ,
		\rf_rf_we_reg/P0001 ,
		_w1973_,
		_w8237_,
		_w8427_
	);
	LUT4 #(
		.INIT('h2aea)
	) name6527 (
		\rf_conf12_reg[15]/NET0131 ,
		\rf_rf_we_reg/P0001 ,
		_w1973_,
		_w8252_,
		_w8428_
	);
	LUT4 #(
		.INIT('h2aea)
	) name6528 (
		\rf_conf12_reg[1]/NET0131 ,
		\rf_rf_we_reg/P0001 ,
		_w1973_,
		_w8267_,
		_w8429_
	);
	LUT4 #(
		.INIT('h2aea)
	) name6529 (
		\rf_conf12_reg[2]/NET0131 ,
		\rf_rf_we_reg/P0001 ,
		_w1973_,
		_w8282_,
		_w8430_
	);
	LUT4 #(
		.INIT('h2aea)
	) name6530 (
		\rf_conf12_reg[3]/NET0131 ,
		\rf_rf_we_reg/P0001 ,
		_w1973_,
		_w8297_,
		_w8431_
	);
	LUT4 #(
		.INIT('h2aea)
	) name6531 (
		\rf_conf12_reg[4]/NET0131 ,
		\rf_rf_we_reg/P0001 ,
		_w1973_,
		_w8312_,
		_w8432_
	);
	LUT4 #(
		.INIT('h2aea)
	) name6532 (
		\rf_conf12_reg[5]/NET0131 ,
		\rf_rf_we_reg/P0001 ,
		_w1973_,
		_w8327_,
		_w8433_
	);
	LUT4 #(
		.INIT('h2aea)
	) name6533 (
		\rf_conf12_reg[6]/NET0131 ,
		\rf_rf_we_reg/P0001 ,
		_w1973_,
		_w8342_,
		_w8434_
	);
	LUT4 #(
		.INIT('h2aea)
	) name6534 (
		\rf_conf12_reg[7]/NET0131 ,
		\rf_rf_we_reg/P0001 ,
		_w1973_,
		_w8357_,
		_w8435_
	);
	LUT4 #(
		.INIT('h2aea)
	) name6535 (
		\rf_conf12_reg[8]/NET0131 ,
		\rf_rf_we_reg/P0001 ,
		_w1973_,
		_w8372_,
		_w8436_
	);
	LUT4 #(
		.INIT('h2aea)
	) name6536 (
		\rf_conf12_reg[9]/NET0131 ,
		\rf_rf_we_reg/P0001 ,
		_w1973_,
		_w8387_,
		_w8437_
	);
	LUT4 #(
		.INIT('h2aea)
	) name6537 (
		\rf_conf13_reg[0]/NET0131 ,
		\rf_rf_we_reg/P0001 ,
		_w1992_,
		_w8162_,
		_w8438_
	);
	LUT4 #(
		.INIT('h2aea)
	) name6538 (
		\rf_conf13_reg[11]/NET0131 ,
		\rf_rf_we_reg/P0001 ,
		_w1992_,
		_w8192_,
		_w8439_
	);
	LUT4 #(
		.INIT('h2aea)
	) name6539 (
		\rf_conf13_reg[10]/NET0131 ,
		\rf_rf_we_reg/P0001 ,
		_w1992_,
		_w8177_,
		_w8440_
	);
	LUT4 #(
		.INIT('h2aea)
	) name6540 (
		\rf_conf13_reg[12]/NET0131 ,
		\rf_rf_we_reg/P0001 ,
		_w1992_,
		_w8207_,
		_w8441_
	);
	LUT4 #(
		.INIT('h2aea)
	) name6541 (
		\rf_conf13_reg[13]/NET0131 ,
		\rf_rf_we_reg/P0001 ,
		_w1992_,
		_w8222_,
		_w8442_
	);
	LUT4 #(
		.INIT('h2aea)
	) name6542 (
		\rf_conf13_reg[14]/NET0131 ,
		\rf_rf_we_reg/P0001 ,
		_w1992_,
		_w8237_,
		_w8443_
	);
	LUT4 #(
		.INIT('h2aea)
	) name6543 (
		\rf_conf13_reg[15]/NET0131 ,
		\rf_rf_we_reg/P0001 ,
		_w1992_,
		_w8252_,
		_w8444_
	);
	LUT4 #(
		.INIT('h2aea)
	) name6544 (
		\rf_conf13_reg[1]/NET0131 ,
		\rf_rf_we_reg/P0001 ,
		_w1992_,
		_w8267_,
		_w8445_
	);
	LUT4 #(
		.INIT('h2aea)
	) name6545 (
		\rf_conf13_reg[2]/NET0131 ,
		\rf_rf_we_reg/P0001 ,
		_w1992_,
		_w8282_,
		_w8446_
	);
	LUT4 #(
		.INIT('h2aea)
	) name6546 (
		\rf_conf13_reg[3]/NET0131 ,
		\rf_rf_we_reg/P0001 ,
		_w1992_,
		_w8297_,
		_w8447_
	);
	LUT4 #(
		.INIT('h2aea)
	) name6547 (
		\rf_conf13_reg[4]/NET0131 ,
		\rf_rf_we_reg/P0001 ,
		_w1992_,
		_w8312_,
		_w8448_
	);
	LUT4 #(
		.INIT('h2aea)
	) name6548 (
		\rf_conf13_reg[5]/NET0131 ,
		\rf_rf_we_reg/P0001 ,
		_w1992_,
		_w8327_,
		_w8449_
	);
	LUT4 #(
		.INIT('h2aea)
	) name6549 (
		\rf_conf13_reg[6]/NET0131 ,
		\rf_rf_we_reg/P0001 ,
		_w1992_,
		_w8342_,
		_w8450_
	);
	LUT4 #(
		.INIT('h2aea)
	) name6550 (
		\rf_conf13_reg[7]/NET0131 ,
		\rf_rf_we_reg/P0001 ,
		_w1992_,
		_w8357_,
		_w8451_
	);
	LUT4 #(
		.INIT('h2aea)
	) name6551 (
		\rf_conf13_reg[8]/NET0131 ,
		\rf_rf_we_reg/P0001 ,
		_w1992_,
		_w8372_,
		_w8452_
	);
	LUT4 #(
		.INIT('h2aea)
	) name6552 (
		\rf_conf13_reg[9]/NET0131 ,
		\rf_rf_we_reg/P0001 ,
		_w1992_,
		_w8387_,
		_w8453_
	);
	LUT4 #(
		.INIT('h2aea)
	) name6553 (
		\rf_conf14_reg[0]/NET0131 ,
		\rf_rf_we_reg/P0001 ,
		_w1974_,
		_w8162_,
		_w8454_
	);
	LUT4 #(
		.INIT('h2aea)
	) name6554 (
		\rf_conf14_reg[10]/NET0131 ,
		\rf_rf_we_reg/P0001 ,
		_w1974_,
		_w8177_,
		_w8455_
	);
	LUT4 #(
		.INIT('h2aea)
	) name6555 (
		\rf_conf14_reg[11]/NET0131 ,
		\rf_rf_we_reg/P0001 ,
		_w1974_,
		_w8192_,
		_w8456_
	);
	LUT4 #(
		.INIT('h2aea)
	) name6556 (
		\rf_conf14_reg[13]/NET0131 ,
		\rf_rf_we_reg/P0001 ,
		_w1974_,
		_w8222_,
		_w8457_
	);
	LUT4 #(
		.INIT('h2aea)
	) name6557 (
		\rf_conf14_reg[14]/NET0131 ,
		\rf_rf_we_reg/P0001 ,
		_w1974_,
		_w8237_,
		_w8458_
	);
	LUT4 #(
		.INIT('h2aea)
	) name6558 (
		\rf_conf14_reg[12]/NET0131 ,
		\rf_rf_we_reg/P0001 ,
		_w1974_,
		_w8207_,
		_w8459_
	);
	LUT4 #(
		.INIT('h2aea)
	) name6559 (
		\rf_conf14_reg[15]/NET0131 ,
		\rf_rf_we_reg/P0001 ,
		_w1974_,
		_w8252_,
		_w8460_
	);
	LUT4 #(
		.INIT('h2aea)
	) name6560 (
		\rf_conf14_reg[1]/NET0131 ,
		\rf_rf_we_reg/P0001 ,
		_w1974_,
		_w8267_,
		_w8461_
	);
	LUT4 #(
		.INIT('h2aea)
	) name6561 (
		\rf_conf14_reg[2]/NET0131 ,
		\rf_rf_we_reg/P0001 ,
		_w1974_,
		_w8282_,
		_w8462_
	);
	LUT4 #(
		.INIT('h2aea)
	) name6562 (
		\rf_conf14_reg[3]/NET0131 ,
		\rf_rf_we_reg/P0001 ,
		_w1974_,
		_w8297_,
		_w8463_
	);
	LUT4 #(
		.INIT('h2aea)
	) name6563 (
		\rf_conf14_reg[5]/NET0131 ,
		\rf_rf_we_reg/P0001 ,
		_w1974_,
		_w8327_,
		_w8464_
	);
	LUT4 #(
		.INIT('h2aea)
	) name6564 (
		\rf_conf14_reg[4]/NET0131 ,
		\rf_rf_we_reg/P0001 ,
		_w1974_,
		_w8312_,
		_w8465_
	);
	LUT4 #(
		.INIT('h2aea)
	) name6565 (
		\rf_conf14_reg[6]/NET0131 ,
		\rf_rf_we_reg/P0001 ,
		_w1974_,
		_w8342_,
		_w8466_
	);
	LUT4 #(
		.INIT('h2aea)
	) name6566 (
		\rf_conf14_reg[7]/NET0131 ,
		\rf_rf_we_reg/P0001 ,
		_w1974_,
		_w8357_,
		_w8467_
	);
	LUT4 #(
		.INIT('h2aea)
	) name6567 (
		\rf_conf14_reg[8]/NET0131 ,
		\rf_rf_we_reg/P0001 ,
		_w1974_,
		_w8372_,
		_w8468_
	);
	LUT4 #(
		.INIT('h2aea)
	) name6568 (
		\rf_conf14_reg[9]/NET0131 ,
		\rf_rf_we_reg/P0001 ,
		_w1974_,
		_w8387_,
		_w8469_
	);
	LUT4 #(
		.INIT('h2aea)
	) name6569 (
		\rf_conf15_reg[0]/NET0131 ,
		\rf_rf_we_reg/P0001 ,
		_w1993_,
		_w8162_,
		_w8470_
	);
	LUT4 #(
		.INIT('h2aea)
	) name6570 (
		\rf_conf15_reg[10]/NET0131 ,
		\rf_rf_we_reg/P0001 ,
		_w1993_,
		_w8177_,
		_w8471_
	);
	LUT4 #(
		.INIT('h2aea)
	) name6571 (
		\rf_conf15_reg[11]/NET0131 ,
		\rf_rf_we_reg/P0001 ,
		_w1993_,
		_w8192_,
		_w8472_
	);
	LUT4 #(
		.INIT('h2aea)
	) name6572 (
		\rf_conf15_reg[12]/NET0131 ,
		\rf_rf_we_reg/P0001 ,
		_w1993_,
		_w8207_,
		_w8473_
	);
	LUT4 #(
		.INIT('h2aea)
	) name6573 (
		\rf_conf15_reg[13]/NET0131 ,
		\rf_rf_we_reg/P0001 ,
		_w1993_,
		_w8222_,
		_w8474_
	);
	LUT4 #(
		.INIT('h2aea)
	) name6574 (
		\rf_conf15_reg[14]/NET0131 ,
		\rf_rf_we_reg/P0001 ,
		_w1993_,
		_w8237_,
		_w8475_
	);
	LUT4 #(
		.INIT('h2aea)
	) name6575 (
		\rf_conf15_reg[15]/NET0131 ,
		\rf_rf_we_reg/P0001 ,
		_w1993_,
		_w8252_,
		_w8476_
	);
	LUT4 #(
		.INIT('h2aea)
	) name6576 (
		\rf_conf15_reg[1]/NET0131 ,
		\rf_rf_we_reg/P0001 ,
		_w1993_,
		_w8267_,
		_w8477_
	);
	LUT4 #(
		.INIT('h2aea)
	) name6577 (
		\rf_conf15_reg[2]/NET0131 ,
		\rf_rf_we_reg/P0001 ,
		_w1993_,
		_w8282_,
		_w8478_
	);
	LUT4 #(
		.INIT('h2aea)
	) name6578 (
		\rf_conf15_reg[3]/NET0131 ,
		\rf_rf_we_reg/P0001 ,
		_w1993_,
		_w8297_,
		_w8479_
	);
	LUT4 #(
		.INIT('h2aea)
	) name6579 (
		\rf_conf15_reg[4]/NET0131 ,
		\rf_rf_we_reg/P0001 ,
		_w1993_,
		_w8312_,
		_w8480_
	);
	LUT4 #(
		.INIT('h2aea)
	) name6580 (
		\rf_conf15_reg[5]/NET0131 ,
		\rf_rf_we_reg/P0001 ,
		_w1993_,
		_w8327_,
		_w8481_
	);
	LUT4 #(
		.INIT('h2aea)
	) name6581 (
		\rf_conf15_reg[6]/NET0131 ,
		\rf_rf_we_reg/P0001 ,
		_w1993_,
		_w8342_,
		_w8482_
	);
	LUT4 #(
		.INIT('h2aea)
	) name6582 (
		\rf_conf15_reg[8]/NET0131 ,
		\rf_rf_we_reg/P0001 ,
		_w1993_,
		_w8372_,
		_w8483_
	);
	LUT4 #(
		.INIT('h2aea)
	) name6583 (
		\rf_conf15_reg[7]/NET0131 ,
		\rf_rf_we_reg/P0001 ,
		_w1993_,
		_w8357_,
		_w8484_
	);
	LUT4 #(
		.INIT('h2aea)
	) name6584 (
		\rf_conf15_reg[9]/NET0131 ,
		\rf_rf_we_reg/P0001 ,
		_w1993_,
		_w8387_,
		_w8485_
	);
	LUT4 #(
		.INIT('h2aea)
	) name6585 (
		\rf_conf1_reg[0]/NET0131 ,
		\rf_rf_we_reg/P0001 ,
		_w1977_,
		_w8162_,
		_w8486_
	);
	LUT4 #(
		.INIT('h2aea)
	) name6586 (
		\rf_conf1_reg[10]/NET0131 ,
		\rf_rf_we_reg/P0001 ,
		_w1977_,
		_w8177_,
		_w8487_
	);
	LUT4 #(
		.INIT('h2aea)
	) name6587 (
		\rf_conf1_reg[11]/NET0131 ,
		\rf_rf_we_reg/P0001 ,
		_w1977_,
		_w8192_,
		_w8488_
	);
	LUT4 #(
		.INIT('h2aea)
	) name6588 (
		\rf_conf1_reg[13]/NET0131 ,
		\rf_rf_we_reg/P0001 ,
		_w1977_,
		_w8222_,
		_w8489_
	);
	LUT4 #(
		.INIT('h2aea)
	) name6589 (
		\rf_conf1_reg[12]/NET0131 ,
		\rf_rf_we_reg/P0001 ,
		_w1977_,
		_w8207_,
		_w8490_
	);
	LUT4 #(
		.INIT('h2aea)
	) name6590 (
		\rf_conf1_reg[14]/NET0131 ,
		\rf_rf_we_reg/P0001 ,
		_w1977_,
		_w8237_,
		_w8491_
	);
	LUT4 #(
		.INIT('h2aea)
	) name6591 (
		\rf_conf1_reg[15]/NET0131 ,
		\rf_rf_we_reg/P0001 ,
		_w1977_,
		_w8252_,
		_w8492_
	);
	LUT4 #(
		.INIT('h2aea)
	) name6592 (
		\rf_conf1_reg[1]/NET0131 ,
		\rf_rf_we_reg/P0001 ,
		_w1977_,
		_w8267_,
		_w8493_
	);
	LUT4 #(
		.INIT('h2aea)
	) name6593 (
		\rf_conf1_reg[2]/NET0131 ,
		\rf_rf_we_reg/P0001 ,
		_w1977_,
		_w8282_,
		_w8494_
	);
	LUT4 #(
		.INIT('h2aea)
	) name6594 (
		\rf_conf1_reg[3]/NET0131 ,
		\rf_rf_we_reg/P0001 ,
		_w1977_,
		_w8297_,
		_w8495_
	);
	LUT4 #(
		.INIT('h2aea)
	) name6595 (
		\rf_conf1_reg[4]/NET0131 ,
		\rf_rf_we_reg/P0001 ,
		_w1977_,
		_w8312_,
		_w8496_
	);
	LUT4 #(
		.INIT('h2aea)
	) name6596 (
		\rf_conf1_reg[5]/NET0131 ,
		\rf_rf_we_reg/P0001 ,
		_w1977_,
		_w8327_,
		_w8497_
	);
	LUT4 #(
		.INIT('h2aea)
	) name6597 (
		\rf_conf1_reg[6]/NET0131 ,
		\rf_rf_we_reg/P0001 ,
		_w1977_,
		_w8342_,
		_w8498_
	);
	LUT4 #(
		.INIT('h2aea)
	) name6598 (
		\rf_conf1_reg[7]/NET0131 ,
		\rf_rf_we_reg/P0001 ,
		_w1977_,
		_w8357_,
		_w8499_
	);
	LUT4 #(
		.INIT('h2aea)
	) name6599 (
		\rf_conf1_reg[8]/NET0131 ,
		\rf_rf_we_reg/P0001 ,
		_w1977_,
		_w8372_,
		_w8500_
	);
	LUT4 #(
		.INIT('h2aea)
	) name6600 (
		\rf_conf1_reg[9]/NET0131 ,
		\rf_rf_we_reg/P0001 ,
		_w1977_,
		_w8387_,
		_w8501_
	);
	LUT4 #(
		.INIT('h2aea)
	) name6601 (
		\rf_conf2_reg[0]/NET0131 ,
		\rf_rf_we_reg/P0001 ,
		_w1976_,
		_w8162_,
		_w8502_
	);
	LUT4 #(
		.INIT('h2aea)
	) name6602 (
		\rf_conf2_reg[10]/NET0131 ,
		\rf_rf_we_reg/P0001 ,
		_w1976_,
		_w8177_,
		_w8503_
	);
	LUT4 #(
		.INIT('h2aea)
	) name6603 (
		\rf_conf2_reg[11]/NET0131 ,
		\rf_rf_we_reg/P0001 ,
		_w1976_,
		_w8192_,
		_w8504_
	);
	LUT4 #(
		.INIT('h2aea)
	) name6604 (
		\rf_conf2_reg[12]/NET0131 ,
		\rf_rf_we_reg/P0001 ,
		_w1976_,
		_w8207_,
		_w8505_
	);
	LUT4 #(
		.INIT('h2aea)
	) name6605 (
		\rf_conf2_reg[13]/NET0131 ,
		\rf_rf_we_reg/P0001 ,
		_w1976_,
		_w8222_,
		_w8506_
	);
	LUT4 #(
		.INIT('h2aea)
	) name6606 (
		\rf_conf2_reg[14]/NET0131 ,
		\rf_rf_we_reg/P0001 ,
		_w1976_,
		_w8237_,
		_w8507_
	);
	LUT4 #(
		.INIT('h2aea)
	) name6607 (
		\rf_conf2_reg[1]/NET0131 ,
		\rf_rf_we_reg/P0001 ,
		_w1976_,
		_w8267_,
		_w8508_
	);
	LUT4 #(
		.INIT('h2aea)
	) name6608 (
		\rf_conf2_reg[15]/NET0131 ,
		\rf_rf_we_reg/P0001 ,
		_w1976_,
		_w8252_,
		_w8509_
	);
	LUT4 #(
		.INIT('h2aea)
	) name6609 (
		\rf_conf2_reg[2]/NET0131 ,
		\rf_rf_we_reg/P0001 ,
		_w1976_,
		_w8282_,
		_w8510_
	);
	LUT4 #(
		.INIT('h2aea)
	) name6610 (
		\rf_conf2_reg[3]/NET0131 ,
		\rf_rf_we_reg/P0001 ,
		_w1976_,
		_w8297_,
		_w8511_
	);
	LUT4 #(
		.INIT('h2aea)
	) name6611 (
		\rf_conf2_reg[4]/NET0131 ,
		\rf_rf_we_reg/P0001 ,
		_w1976_,
		_w8312_,
		_w8512_
	);
	LUT4 #(
		.INIT('h2aea)
	) name6612 (
		\rf_conf2_reg[5]/NET0131 ,
		\rf_rf_we_reg/P0001 ,
		_w1976_,
		_w8327_,
		_w8513_
	);
	LUT4 #(
		.INIT('h2aea)
	) name6613 (
		\rf_conf2_reg[6]/NET0131 ,
		\rf_rf_we_reg/P0001 ,
		_w1976_,
		_w8342_,
		_w8514_
	);
	LUT4 #(
		.INIT('h2aea)
	) name6614 (
		\rf_conf2_reg[7]/NET0131 ,
		\rf_rf_we_reg/P0001 ,
		_w1976_,
		_w8357_,
		_w8515_
	);
	LUT4 #(
		.INIT('h2aea)
	) name6615 (
		\rf_conf2_reg[8]/NET0131 ,
		\rf_rf_we_reg/P0001 ,
		_w1976_,
		_w8372_,
		_w8516_
	);
	LUT4 #(
		.INIT('h2aea)
	) name6616 (
		\rf_conf2_reg[9]/NET0131 ,
		\rf_rf_we_reg/P0001 ,
		_w1976_,
		_w8387_,
		_w8517_
	);
	LUT4 #(
		.INIT('h2aea)
	) name6617 (
		\rf_conf3_reg[0]/NET0131 ,
		\rf_rf_we_reg/P0001 ,
		_w1971_,
		_w8162_,
		_w8518_
	);
	LUT4 #(
		.INIT('h2aea)
	) name6618 (
		\rf_conf3_reg[10]/NET0131 ,
		\rf_rf_we_reg/P0001 ,
		_w1971_,
		_w8177_,
		_w8519_
	);
	LUT4 #(
		.INIT('h2aea)
	) name6619 (
		\rf_conf3_reg[11]/NET0131 ,
		\rf_rf_we_reg/P0001 ,
		_w1971_,
		_w8192_,
		_w8520_
	);
	LUT4 #(
		.INIT('h2aea)
	) name6620 (
		\rf_conf3_reg[12]/NET0131 ,
		\rf_rf_we_reg/P0001 ,
		_w1971_,
		_w8207_,
		_w8521_
	);
	LUT4 #(
		.INIT('h2aea)
	) name6621 (
		\rf_conf3_reg[13]/NET0131 ,
		\rf_rf_we_reg/P0001 ,
		_w1971_,
		_w8222_,
		_w8522_
	);
	LUT4 #(
		.INIT('h2aea)
	) name6622 (
		\rf_conf3_reg[14]/NET0131 ,
		\rf_rf_we_reg/P0001 ,
		_w1971_,
		_w8237_,
		_w8523_
	);
	LUT4 #(
		.INIT('h2aea)
	) name6623 (
		\rf_conf3_reg[15]/NET0131 ,
		\rf_rf_we_reg/P0001 ,
		_w1971_,
		_w8252_,
		_w8524_
	);
	LUT4 #(
		.INIT('h2aea)
	) name6624 (
		\rf_conf3_reg[1]/NET0131 ,
		\rf_rf_we_reg/P0001 ,
		_w1971_,
		_w8267_,
		_w8525_
	);
	LUT4 #(
		.INIT('h2aea)
	) name6625 (
		\rf_conf3_reg[2]/NET0131 ,
		\rf_rf_we_reg/P0001 ,
		_w1971_,
		_w8282_,
		_w8526_
	);
	LUT4 #(
		.INIT('h2aea)
	) name6626 (
		\rf_conf3_reg[4]/NET0131 ,
		\rf_rf_we_reg/P0001 ,
		_w1971_,
		_w8312_,
		_w8527_
	);
	LUT4 #(
		.INIT('h2aea)
	) name6627 (
		\rf_conf3_reg[3]/NET0131 ,
		\rf_rf_we_reg/P0001 ,
		_w1971_,
		_w8297_,
		_w8528_
	);
	LUT4 #(
		.INIT('h2aea)
	) name6628 (
		\rf_conf3_reg[5]/NET0131 ,
		\rf_rf_we_reg/P0001 ,
		_w1971_,
		_w8327_,
		_w8529_
	);
	LUT4 #(
		.INIT('h2aea)
	) name6629 (
		\rf_conf3_reg[6]/NET0131 ,
		\rf_rf_we_reg/P0001 ,
		_w1971_,
		_w8342_,
		_w8530_
	);
	LUT4 #(
		.INIT('h2aea)
	) name6630 (
		\rf_conf3_reg[7]/NET0131 ,
		\rf_rf_we_reg/P0001 ,
		_w1971_,
		_w8357_,
		_w8531_
	);
	LUT4 #(
		.INIT('h2aea)
	) name6631 (
		\rf_conf3_reg[8]/NET0131 ,
		\rf_rf_we_reg/P0001 ,
		_w1971_,
		_w8372_,
		_w8532_
	);
	LUT4 #(
		.INIT('h2aea)
	) name6632 (
		\rf_conf3_reg[9]/NET0131 ,
		\rf_rf_we_reg/P0001 ,
		_w1971_,
		_w8387_,
		_w8533_
	);
	LUT4 #(
		.INIT('h2aea)
	) name6633 (
		\rf_conf4_reg[0]/NET0131 ,
		\rf_rf_we_reg/P0001 ,
		_w1980_,
		_w8162_,
		_w8534_
	);
	LUT4 #(
		.INIT('h2aea)
	) name6634 (
		\rf_conf4_reg[10]/NET0131 ,
		\rf_rf_we_reg/P0001 ,
		_w1980_,
		_w8177_,
		_w8535_
	);
	LUT4 #(
		.INIT('h2aea)
	) name6635 (
		\rf_conf4_reg[11]/NET0131 ,
		\rf_rf_we_reg/P0001 ,
		_w1980_,
		_w8192_,
		_w8536_
	);
	LUT4 #(
		.INIT('h2aea)
	) name6636 (
		\rf_conf4_reg[12]/NET0131 ,
		\rf_rf_we_reg/P0001 ,
		_w1980_,
		_w8207_,
		_w8537_
	);
	LUT4 #(
		.INIT('h2aea)
	) name6637 (
		\rf_conf4_reg[13]/NET0131 ,
		\rf_rf_we_reg/P0001 ,
		_w1980_,
		_w8222_,
		_w8538_
	);
	LUT4 #(
		.INIT('h2aea)
	) name6638 (
		\rf_conf4_reg[14]/NET0131 ,
		\rf_rf_we_reg/P0001 ,
		_w1980_,
		_w8237_,
		_w8539_
	);
	LUT4 #(
		.INIT('h2aea)
	) name6639 (
		\rf_conf4_reg[15]/NET0131 ,
		\rf_rf_we_reg/P0001 ,
		_w1980_,
		_w8252_,
		_w8540_
	);
	LUT4 #(
		.INIT('h2aea)
	) name6640 (
		\rf_conf4_reg[1]/NET0131 ,
		\rf_rf_we_reg/P0001 ,
		_w1980_,
		_w8267_,
		_w8541_
	);
	LUT4 #(
		.INIT('h2aea)
	) name6641 (
		\rf_conf4_reg[2]/NET0131 ,
		\rf_rf_we_reg/P0001 ,
		_w1980_,
		_w8282_,
		_w8542_
	);
	LUT4 #(
		.INIT('h2aea)
	) name6642 (
		\rf_conf4_reg[3]/NET0131 ,
		\rf_rf_we_reg/P0001 ,
		_w1980_,
		_w8297_,
		_w8543_
	);
	LUT4 #(
		.INIT('h2aea)
	) name6643 (
		\rf_conf4_reg[4]/NET0131 ,
		\rf_rf_we_reg/P0001 ,
		_w1980_,
		_w8312_,
		_w8544_
	);
	LUT4 #(
		.INIT('h2aea)
	) name6644 (
		\rf_conf4_reg[5]/NET0131 ,
		\rf_rf_we_reg/P0001 ,
		_w1980_,
		_w8327_,
		_w8545_
	);
	LUT4 #(
		.INIT('h2aea)
	) name6645 (
		\rf_conf4_reg[6]/NET0131 ,
		\rf_rf_we_reg/P0001 ,
		_w1980_,
		_w8342_,
		_w8546_
	);
	LUT4 #(
		.INIT('h2aea)
	) name6646 (
		\rf_conf4_reg[7]/NET0131 ,
		\rf_rf_we_reg/P0001 ,
		_w1980_,
		_w8357_,
		_w8547_
	);
	LUT4 #(
		.INIT('h2aea)
	) name6647 (
		\rf_conf4_reg[8]/NET0131 ,
		\rf_rf_we_reg/P0001 ,
		_w1980_,
		_w8372_,
		_w8548_
	);
	LUT4 #(
		.INIT('h2aea)
	) name6648 (
		\rf_conf4_reg[9]/NET0131 ,
		\rf_rf_we_reg/P0001 ,
		_w1980_,
		_w8387_,
		_w8549_
	);
	LUT4 #(
		.INIT('h2aea)
	) name6649 (
		\rf_conf5_reg[0]/NET0131 ,
		\rf_rf_we_reg/P0001 ,
		_w1970_,
		_w8162_,
		_w8550_
	);
	LUT4 #(
		.INIT('h2aea)
	) name6650 (
		\rf_conf5_reg[10]/NET0131 ,
		\rf_rf_we_reg/P0001 ,
		_w1970_,
		_w8177_,
		_w8551_
	);
	LUT4 #(
		.INIT('h2aea)
	) name6651 (
		\rf_conf5_reg[11]/NET0131 ,
		\rf_rf_we_reg/P0001 ,
		_w1970_,
		_w8192_,
		_w8552_
	);
	LUT4 #(
		.INIT('h2aea)
	) name6652 (
		\rf_conf5_reg[12]/NET0131 ,
		\rf_rf_we_reg/P0001 ,
		_w1970_,
		_w8207_,
		_w8553_
	);
	LUT4 #(
		.INIT('h2aea)
	) name6653 (
		\rf_conf5_reg[13]/NET0131 ,
		\rf_rf_we_reg/P0001 ,
		_w1970_,
		_w8222_,
		_w8554_
	);
	LUT4 #(
		.INIT('h2aea)
	) name6654 (
		\rf_conf5_reg[14]/NET0131 ,
		\rf_rf_we_reg/P0001 ,
		_w1970_,
		_w8237_,
		_w8555_
	);
	LUT4 #(
		.INIT('h2aea)
	) name6655 (
		\rf_conf5_reg[15]/NET0131 ,
		\rf_rf_we_reg/P0001 ,
		_w1970_,
		_w8252_,
		_w8556_
	);
	LUT4 #(
		.INIT('h2aea)
	) name6656 (
		\rf_conf5_reg[1]/NET0131 ,
		\rf_rf_we_reg/P0001 ,
		_w1970_,
		_w8267_,
		_w8557_
	);
	LUT4 #(
		.INIT('h2aea)
	) name6657 (
		\rf_conf5_reg[3]/NET0131 ,
		\rf_rf_we_reg/P0001 ,
		_w1970_,
		_w8297_,
		_w8558_
	);
	LUT4 #(
		.INIT('h2aea)
	) name6658 (
		\rf_conf5_reg[2]/NET0131 ,
		\rf_rf_we_reg/P0001 ,
		_w1970_,
		_w8282_,
		_w8559_
	);
	LUT4 #(
		.INIT('h2aea)
	) name6659 (
		\rf_conf5_reg[4]/NET0131 ,
		\rf_rf_we_reg/P0001 ,
		_w1970_,
		_w8312_,
		_w8560_
	);
	LUT4 #(
		.INIT('h2aea)
	) name6660 (
		\rf_conf5_reg[5]/NET0131 ,
		\rf_rf_we_reg/P0001 ,
		_w1970_,
		_w8327_,
		_w8561_
	);
	LUT4 #(
		.INIT('h2aea)
	) name6661 (
		\rf_conf5_reg[6]/NET0131 ,
		\rf_rf_we_reg/P0001 ,
		_w1970_,
		_w8342_,
		_w8562_
	);
	LUT4 #(
		.INIT('h2aea)
	) name6662 (
		\rf_conf5_reg[7]/NET0131 ,
		\rf_rf_we_reg/P0001 ,
		_w1970_,
		_w8357_,
		_w8563_
	);
	LUT4 #(
		.INIT('h2aea)
	) name6663 (
		\rf_conf5_reg[8]/NET0131 ,
		\rf_rf_we_reg/P0001 ,
		_w1970_,
		_w8372_,
		_w8564_
	);
	LUT4 #(
		.INIT('h2aea)
	) name6664 (
		\rf_conf5_reg[9]/NET0131 ,
		\rf_rf_we_reg/P0001 ,
		_w1970_,
		_w8387_,
		_w8565_
	);
	LUT4 #(
		.INIT('h2aea)
	) name6665 (
		\rf_conf6_reg[0]/NET0131 ,
		\rf_rf_we_reg/P0001 ,
		_w1983_,
		_w8162_,
		_w8566_
	);
	LUT4 #(
		.INIT('h2aea)
	) name6666 (
		\rf_conf6_reg[10]/NET0131 ,
		\rf_rf_we_reg/P0001 ,
		_w1983_,
		_w8177_,
		_w8567_
	);
	LUT4 #(
		.INIT('h2aea)
	) name6667 (
		\rf_conf6_reg[11]/NET0131 ,
		\rf_rf_we_reg/P0001 ,
		_w1983_,
		_w8192_,
		_w8568_
	);
	LUT4 #(
		.INIT('h2aea)
	) name6668 (
		\rf_conf6_reg[12]/NET0131 ,
		\rf_rf_we_reg/P0001 ,
		_w1983_,
		_w8207_,
		_w8569_
	);
	LUT4 #(
		.INIT('h2aea)
	) name6669 (
		\rf_conf6_reg[13]/NET0131 ,
		\rf_rf_we_reg/P0001 ,
		_w1983_,
		_w8222_,
		_w8570_
	);
	LUT4 #(
		.INIT('h2aea)
	) name6670 (
		\rf_conf6_reg[14]/NET0131 ,
		\rf_rf_we_reg/P0001 ,
		_w1983_,
		_w8237_,
		_w8571_
	);
	LUT4 #(
		.INIT('h2aea)
	) name6671 (
		\rf_conf6_reg[15]/NET0131 ,
		\rf_rf_we_reg/P0001 ,
		_w1983_,
		_w8252_,
		_w8572_
	);
	LUT4 #(
		.INIT('h2aea)
	) name6672 (
		\rf_conf6_reg[1]/NET0131 ,
		\rf_rf_we_reg/P0001 ,
		_w1983_,
		_w8267_,
		_w8573_
	);
	LUT4 #(
		.INIT('h2aea)
	) name6673 (
		\rf_conf6_reg[2]/NET0131 ,
		\rf_rf_we_reg/P0001 ,
		_w1983_,
		_w8282_,
		_w8574_
	);
	LUT4 #(
		.INIT('h2aea)
	) name6674 (
		\rf_conf6_reg[3]/NET0131 ,
		\rf_rf_we_reg/P0001 ,
		_w1983_,
		_w8297_,
		_w8575_
	);
	LUT4 #(
		.INIT('h2aea)
	) name6675 (
		\rf_conf6_reg[4]/NET0131 ,
		\rf_rf_we_reg/P0001 ,
		_w1983_,
		_w8312_,
		_w8576_
	);
	LUT4 #(
		.INIT('h2aea)
	) name6676 (
		\rf_conf6_reg[5]/NET0131 ,
		\rf_rf_we_reg/P0001 ,
		_w1983_,
		_w8327_,
		_w8577_
	);
	LUT4 #(
		.INIT('h2aea)
	) name6677 (
		\rf_conf6_reg[6]/NET0131 ,
		\rf_rf_we_reg/P0001 ,
		_w1983_,
		_w8342_,
		_w8578_
	);
	LUT4 #(
		.INIT('h2aea)
	) name6678 (
		\rf_conf6_reg[7]/NET0131 ,
		\rf_rf_we_reg/P0001 ,
		_w1983_,
		_w8357_,
		_w8579_
	);
	LUT4 #(
		.INIT('h2aea)
	) name6679 (
		\rf_conf6_reg[8]/NET0131 ,
		\rf_rf_we_reg/P0001 ,
		_w1983_,
		_w8372_,
		_w8580_
	);
	LUT4 #(
		.INIT('h2aea)
	) name6680 (
		\rf_conf6_reg[9]/NET0131 ,
		\rf_rf_we_reg/P0001 ,
		_w1983_,
		_w8387_,
		_w8581_
	);
	LUT4 #(
		.INIT('h2aea)
	) name6681 (
		\rf_conf7_reg[0]/NET0131 ,
		\rf_rf_we_reg/P0001 ,
		_w1984_,
		_w8162_,
		_w8582_
	);
	LUT4 #(
		.INIT('h2aea)
	) name6682 (
		\rf_conf7_reg[11]/NET0131 ,
		\rf_rf_we_reg/P0001 ,
		_w1984_,
		_w8192_,
		_w8583_
	);
	LUT4 #(
		.INIT('h2aea)
	) name6683 (
		\rf_conf7_reg[10]/NET0131 ,
		\rf_rf_we_reg/P0001 ,
		_w1984_,
		_w8177_,
		_w8584_
	);
	LUT4 #(
		.INIT('h2aea)
	) name6684 (
		\rf_conf7_reg[12]/NET0131 ,
		\rf_rf_we_reg/P0001 ,
		_w1984_,
		_w8207_,
		_w8585_
	);
	LUT4 #(
		.INIT('h2aea)
	) name6685 (
		\rf_conf7_reg[13]/NET0131 ,
		\rf_rf_we_reg/P0001 ,
		_w1984_,
		_w8222_,
		_w8586_
	);
	LUT4 #(
		.INIT('h2aea)
	) name6686 (
		\rf_conf7_reg[14]/NET0131 ,
		\rf_rf_we_reg/P0001 ,
		_w1984_,
		_w8237_,
		_w8587_
	);
	LUT4 #(
		.INIT('h2aea)
	) name6687 (
		\rf_conf7_reg[15]/NET0131 ,
		\rf_rf_we_reg/P0001 ,
		_w1984_,
		_w8252_,
		_w8588_
	);
	LUT4 #(
		.INIT('h2aea)
	) name6688 (
		\rf_conf7_reg[1]/NET0131 ,
		\rf_rf_we_reg/P0001 ,
		_w1984_,
		_w8267_,
		_w8589_
	);
	LUT4 #(
		.INIT('h2aea)
	) name6689 (
		\rf_conf7_reg[2]/NET0131 ,
		\rf_rf_we_reg/P0001 ,
		_w1984_,
		_w8282_,
		_w8590_
	);
	LUT4 #(
		.INIT('h2aea)
	) name6690 (
		\rf_conf7_reg[3]/NET0131 ,
		\rf_rf_we_reg/P0001 ,
		_w1984_,
		_w8297_,
		_w8591_
	);
	LUT4 #(
		.INIT('h2aea)
	) name6691 (
		\rf_conf7_reg[4]/NET0131 ,
		\rf_rf_we_reg/P0001 ,
		_w1984_,
		_w8312_,
		_w8592_
	);
	LUT4 #(
		.INIT('h2aea)
	) name6692 (
		\rf_conf7_reg[5]/NET0131 ,
		\rf_rf_we_reg/P0001 ,
		_w1984_,
		_w8327_,
		_w8593_
	);
	LUT4 #(
		.INIT('h2aea)
	) name6693 (
		\rf_conf7_reg[6]/NET0131 ,
		\rf_rf_we_reg/P0001 ,
		_w1984_,
		_w8342_,
		_w8594_
	);
	LUT4 #(
		.INIT('h2aea)
	) name6694 (
		\rf_conf7_reg[7]/NET0131 ,
		\rf_rf_we_reg/P0001 ,
		_w1984_,
		_w8357_,
		_w8595_
	);
	LUT4 #(
		.INIT('h2aea)
	) name6695 (
		\rf_conf7_reg[8]/NET0131 ,
		\rf_rf_we_reg/P0001 ,
		_w1984_,
		_w8372_,
		_w8596_
	);
	LUT4 #(
		.INIT('h2aea)
	) name6696 (
		\rf_conf7_reg[9]/NET0131 ,
		\rf_rf_we_reg/P0001 ,
		_w1984_,
		_w8387_,
		_w8597_
	);
	LUT4 #(
		.INIT('h2aea)
	) name6697 (
		\rf_conf8_reg[0]/NET0131 ,
		\rf_rf_we_reg/P0001 ,
		_w1986_,
		_w8162_,
		_w8598_
	);
	LUT4 #(
		.INIT('h2aea)
	) name6698 (
		\rf_conf8_reg[10]/NET0131 ,
		\rf_rf_we_reg/P0001 ,
		_w1986_,
		_w8177_,
		_w8599_
	);
	LUT4 #(
		.INIT('h2aea)
	) name6699 (
		\rf_conf8_reg[11]/NET0131 ,
		\rf_rf_we_reg/P0001 ,
		_w1986_,
		_w8192_,
		_w8600_
	);
	LUT4 #(
		.INIT('h2aea)
	) name6700 (
		\rf_conf8_reg[12]/NET0131 ,
		\rf_rf_we_reg/P0001 ,
		_w1986_,
		_w8207_,
		_w8601_
	);
	LUT4 #(
		.INIT('h2aea)
	) name6701 (
		\rf_conf8_reg[13]/NET0131 ,
		\rf_rf_we_reg/P0001 ,
		_w1986_,
		_w8222_,
		_w8602_
	);
	LUT4 #(
		.INIT('h2aea)
	) name6702 (
		\rf_conf8_reg[14]/NET0131 ,
		\rf_rf_we_reg/P0001 ,
		_w1986_,
		_w8237_,
		_w8603_
	);
	LUT4 #(
		.INIT('h2aea)
	) name6703 (
		\rf_conf8_reg[15]/NET0131 ,
		\rf_rf_we_reg/P0001 ,
		_w1986_,
		_w8252_,
		_w8604_
	);
	LUT4 #(
		.INIT('h2aea)
	) name6704 (
		\rf_conf8_reg[1]/NET0131 ,
		\rf_rf_we_reg/P0001 ,
		_w1986_,
		_w8267_,
		_w8605_
	);
	LUT4 #(
		.INIT('h2aea)
	) name6705 (
		\rf_conf8_reg[2]/NET0131 ,
		\rf_rf_we_reg/P0001 ,
		_w1986_,
		_w8282_,
		_w8606_
	);
	LUT4 #(
		.INIT('h2aea)
	) name6706 (
		\rf_conf8_reg[3]/NET0131 ,
		\rf_rf_we_reg/P0001 ,
		_w1986_,
		_w8297_,
		_w8607_
	);
	LUT4 #(
		.INIT('h2aea)
	) name6707 (
		\rf_conf8_reg[5]/NET0131 ,
		\rf_rf_we_reg/P0001 ,
		_w1986_,
		_w8327_,
		_w8608_
	);
	LUT4 #(
		.INIT('h2aea)
	) name6708 (
		\rf_conf8_reg[4]/NET0131 ,
		\rf_rf_we_reg/P0001 ,
		_w1986_,
		_w8312_,
		_w8609_
	);
	LUT4 #(
		.INIT('h2aea)
	) name6709 (
		\rf_conf8_reg[6]/NET0131 ,
		\rf_rf_we_reg/P0001 ,
		_w1986_,
		_w8342_,
		_w8610_
	);
	LUT4 #(
		.INIT('h2aea)
	) name6710 (
		\rf_conf8_reg[7]/NET0131 ,
		\rf_rf_we_reg/P0001 ,
		_w1986_,
		_w8357_,
		_w8611_
	);
	LUT4 #(
		.INIT('h2aea)
	) name6711 (
		\rf_conf8_reg[8]/NET0131 ,
		\rf_rf_we_reg/P0001 ,
		_w1986_,
		_w8372_,
		_w8612_
	);
	LUT4 #(
		.INIT('h2aea)
	) name6712 (
		\rf_conf8_reg[9]/NET0131 ,
		\rf_rf_we_reg/P0001 ,
		_w1986_,
		_w8387_,
		_w8613_
	);
	LUT4 #(
		.INIT('h2aea)
	) name6713 (
		\rf_conf9_reg[0]/NET0131 ,
		\rf_rf_we_reg/P0001 ,
		_w1989_,
		_w8162_,
		_w8614_
	);
	LUT4 #(
		.INIT('h2aea)
	) name6714 (
		\rf_conf9_reg[10]/NET0131 ,
		\rf_rf_we_reg/P0001 ,
		_w1989_,
		_w8177_,
		_w8615_
	);
	LUT4 #(
		.INIT('h2aea)
	) name6715 (
		\rf_conf9_reg[11]/NET0131 ,
		\rf_rf_we_reg/P0001 ,
		_w1989_,
		_w8192_,
		_w8616_
	);
	LUT4 #(
		.INIT('h2aea)
	) name6716 (
		\rf_conf9_reg[12]/NET0131 ,
		\rf_rf_we_reg/P0001 ,
		_w1989_,
		_w8207_,
		_w8617_
	);
	LUT4 #(
		.INIT('h2aea)
	) name6717 (
		\rf_conf9_reg[13]/NET0131 ,
		\rf_rf_we_reg/P0001 ,
		_w1989_,
		_w8222_,
		_w8618_
	);
	LUT4 #(
		.INIT('h2aea)
	) name6718 (
		\rf_conf9_reg[14]/NET0131 ,
		\rf_rf_we_reg/P0001 ,
		_w1989_,
		_w8237_,
		_w8619_
	);
	LUT4 #(
		.INIT('h2aea)
	) name6719 (
		\rf_conf9_reg[15]/NET0131 ,
		\rf_rf_we_reg/P0001 ,
		_w1989_,
		_w8252_,
		_w8620_
	);
	LUT4 #(
		.INIT('h2aea)
	) name6720 (
		\rf_conf9_reg[1]/NET0131 ,
		\rf_rf_we_reg/P0001 ,
		_w1989_,
		_w8267_,
		_w8621_
	);
	LUT4 #(
		.INIT('h2aea)
	) name6721 (
		\rf_conf9_reg[2]/NET0131 ,
		\rf_rf_we_reg/P0001 ,
		_w1989_,
		_w8282_,
		_w8622_
	);
	LUT4 #(
		.INIT('h2aea)
	) name6722 (
		\rf_conf9_reg[3]/NET0131 ,
		\rf_rf_we_reg/P0001 ,
		_w1989_,
		_w8297_,
		_w8623_
	);
	LUT4 #(
		.INIT('h2aea)
	) name6723 (
		\rf_conf9_reg[4]/NET0131 ,
		\rf_rf_we_reg/P0001 ,
		_w1989_,
		_w8312_,
		_w8624_
	);
	LUT4 #(
		.INIT('h2aea)
	) name6724 (
		\rf_conf9_reg[5]/NET0131 ,
		\rf_rf_we_reg/P0001 ,
		_w1989_,
		_w8327_,
		_w8625_
	);
	LUT4 #(
		.INIT('h2aea)
	) name6725 (
		\rf_conf9_reg[6]/NET0131 ,
		\rf_rf_we_reg/P0001 ,
		_w1989_,
		_w8342_,
		_w8626_
	);
	LUT4 #(
		.INIT('h2aea)
	) name6726 (
		\rf_conf9_reg[7]/NET0131 ,
		\rf_rf_we_reg/P0001 ,
		_w1989_,
		_w8357_,
		_w8627_
	);
	LUT4 #(
		.INIT('h2aea)
	) name6727 (
		\rf_conf9_reg[8]/NET0131 ,
		\rf_rf_we_reg/P0001 ,
		_w1989_,
		_w8372_,
		_w8628_
	);
	LUT4 #(
		.INIT('h2aea)
	) name6728 (
		\rf_conf9_reg[9]/NET0131 ,
		\rf_rf_we_reg/P0001 ,
		_w1989_,
		_w8387_,
		_w8629_
	);
	LUT4 #(
		.INIT('h0001)
	) name6729 (
		\rf_rf_ack_reg/P0001 ,
		_w2016_,
		_w2029_,
		_w2043_,
		_w8630_
	);
	LUT2 #(
		.INIT('h8)
	) name6730 (
		_w2097_,
		_w8630_,
		_w8631_
	);
	LUT3 #(
		.INIT('h2a)
	) name6731 (
		\m7_we_i_pad ,
		_w1901_,
		_w1902_,
		_w8632_
	);
	LUT3 #(
		.INIT('h2a)
	) name6732 (
		\m6_we_i_pad ,
		_w1908_,
		_w1909_,
		_w8633_
	);
	LUT4 #(
		.INIT('h153f)
	) name6733 (
		_w1907_,
		_w1918_,
		_w8632_,
		_w8633_,
		_w8634_
	);
	LUT3 #(
		.INIT('h2a)
	) name6734 (
		\m5_we_i_pad ,
		_w1901_,
		_w1902_,
		_w8635_
	);
	LUT3 #(
		.INIT('h2a)
	) name6735 (
		\m2_we_i_pad ,
		_w1908_,
		_w1909_,
		_w8636_
	);
	LUT4 #(
		.INIT('h153f)
	) name6736 (
		_w1914_,
		_w1920_,
		_w8635_,
		_w8636_,
		_w8637_
	);
	LUT3 #(
		.INIT('h80)
	) name6737 (
		\m4_we_i_pad ,
		_w1908_,
		_w1909_,
		_w8638_
	);
	LUT3 #(
		.INIT('h80)
	) name6738 (
		\m3_we_i_pad ,
		_w1901_,
		_w1902_,
		_w8639_
	);
	LUT4 #(
		.INIT('h135f)
	) name6739 (
		_w1907_,
		_w1918_,
		_w8638_,
		_w8639_,
		_w8640_
	);
	LUT3 #(
		.INIT('h80)
	) name6740 (
		\m1_we_i_pad ,
		_w1901_,
		_w1902_,
		_w8641_
	);
	LUT3 #(
		.INIT('h80)
	) name6741 (
		\m0_we_i_pad ,
		_w1908_,
		_w1909_,
		_w8642_
	);
	LUT4 #(
		.INIT('h153f)
	) name6742 (
		_w1914_,
		_w1920_,
		_w8641_,
		_w8642_,
		_w8643_
	);
	LUT4 #(
		.INIT('h8000)
	) name6743 (
		_w8634_,
		_w8637_,
		_w8640_,
		_w8643_,
		_w8644_
	);
	LUT4 #(
		.INIT('h7fff)
	) name6744 (
		_w8634_,
		_w8637_,
		_w8640_,
		_w8643_,
		_w8645_
	);
	LUT2 #(
		.INIT('h1)
	) name6745 (
		\rf_rf_we_reg/P0001 ,
		_w8644_,
		_w8646_
	);
	LUT3 #(
		.INIT('h80)
	) name6746 (
		_w2046_,
		_w2097_,
		_w8646_,
		_w8647_
	);
	LUT4 #(
		.INIT('hf35f)
	) name6747 (
		\s4_msel_arb1_state_reg[1]/NET0131 ,
		\s4_msel_arb2_state_reg[1]/NET0131 ,
		\s4_msel_pri_out_reg[0]/NET0131 ,
		\s4_msel_pri_out_reg[1]/NET0131 ,
		_w8648_
	);
	LUT4 #(
		.INIT('h3ff5)
	) name6748 (
		\s4_msel_arb0_state_reg[1]/NET0131 ,
		\s4_msel_arb3_state_reg[1]/NET0131 ,
		\s4_msel_pri_out_reg[0]/NET0131 ,
		\s4_msel_pri_out_reg[1]/NET0131 ,
		_w8649_
	);
	LUT2 #(
		.INIT('h8)
	) name6749 (
		_w8648_,
		_w8649_,
		_w8650_
	);
	LUT4 #(
		.INIT('h3ff5)
	) name6750 (
		\s4_msel_arb0_state_reg[2]/NET0131 ,
		\s4_msel_arb3_state_reg[2]/NET0131 ,
		\s4_msel_pri_out_reg[0]/NET0131 ,
		\s4_msel_pri_out_reg[1]/NET0131 ,
		_w8651_
	);
	LUT4 #(
		.INIT('hf35f)
	) name6751 (
		\s4_msel_arb1_state_reg[2]/NET0131 ,
		\s4_msel_arb2_state_reg[2]/NET0131 ,
		\s4_msel_pri_out_reg[0]/NET0131 ,
		\s4_msel_pri_out_reg[1]/NET0131 ,
		_w8652_
	);
	LUT2 #(
		.INIT('h8)
	) name6752 (
		_w8651_,
		_w8652_,
		_w8653_
	);
	LUT4 #(
		.INIT('h0888)
	) name6753 (
		_w8648_,
		_w8649_,
		_w8651_,
		_w8652_,
		_w8654_
	);
	LUT4 #(
		.INIT('hf35f)
	) name6754 (
		\s4_msel_arb1_state_reg[0]/NET0131 ,
		\s4_msel_arb2_state_reg[0]/NET0131 ,
		\s4_msel_pri_out_reg[0]/NET0131 ,
		\s4_msel_pri_out_reg[1]/NET0131 ,
		_w8655_
	);
	LUT4 #(
		.INIT('h3ff5)
	) name6755 (
		\s4_msel_arb0_state_reg[0]/NET0131 ,
		\s4_msel_arb3_state_reg[0]/NET0131 ,
		\s4_msel_pri_out_reg[0]/NET0131 ,
		\s4_msel_pri_out_reg[1]/NET0131 ,
		_w8656_
	);
	LUT2 #(
		.INIT('h8)
	) name6756 (
		\m5_s4_cyc_o_reg/NET0131 ,
		\s4_m5_cyc_r_reg/P0001 ,
		_w8657_
	);
	LUT3 #(
		.INIT('h70)
	) name6757 (
		_w8655_,
		_w8656_,
		_w8657_,
		_w8658_
	);
	LUT2 #(
		.INIT('h8)
	) name6758 (
		\m4_s4_cyc_o_reg/NET0131 ,
		\s4_m4_cyc_r_reg/P0001 ,
		_w8659_
	);
	LUT3 #(
		.INIT('h80)
	) name6759 (
		_w8655_,
		_w8656_,
		_w8659_,
		_w8660_
	);
	LUT3 #(
		.INIT('h57)
	) name6760 (
		_w8654_,
		_w8658_,
		_w8660_,
		_w8661_
	);
	LUT4 #(
		.INIT('h8000)
	) name6761 (
		_w8648_,
		_w8649_,
		_w8651_,
		_w8652_,
		_w8662_
	);
	LUT2 #(
		.INIT('h8)
	) name6762 (
		\m1_s4_cyc_o_reg/NET0131 ,
		\s4_m1_cyc_r_reg/P0001 ,
		_w8663_
	);
	LUT3 #(
		.INIT('h70)
	) name6763 (
		_w8655_,
		_w8656_,
		_w8663_,
		_w8664_
	);
	LUT2 #(
		.INIT('h8)
	) name6764 (
		\m0_s4_cyc_o_reg/NET0131 ,
		\s4_m0_cyc_r_reg/P0001 ,
		_w8665_
	);
	LUT3 #(
		.INIT('h80)
	) name6765 (
		_w8655_,
		_w8656_,
		_w8665_,
		_w8666_
	);
	LUT3 #(
		.INIT('h57)
	) name6766 (
		_w8662_,
		_w8664_,
		_w8666_,
		_w8667_
	);
	LUT4 #(
		.INIT('h7000)
	) name6767 (
		_w8648_,
		_w8649_,
		_w8651_,
		_w8652_,
		_w8668_
	);
	LUT2 #(
		.INIT('h8)
	) name6768 (
		\m3_s4_cyc_o_reg/NET0131 ,
		\s4_m3_cyc_r_reg/P0001 ,
		_w8669_
	);
	LUT3 #(
		.INIT('h70)
	) name6769 (
		_w8655_,
		_w8656_,
		_w8669_,
		_w8670_
	);
	LUT2 #(
		.INIT('h8)
	) name6770 (
		\m2_s4_cyc_o_reg/NET0131 ,
		\s4_m2_cyc_r_reg/P0001 ,
		_w8671_
	);
	LUT3 #(
		.INIT('h80)
	) name6771 (
		_w8655_,
		_w8656_,
		_w8671_,
		_w8672_
	);
	LUT3 #(
		.INIT('h57)
	) name6772 (
		_w8668_,
		_w8670_,
		_w8672_,
		_w8673_
	);
	LUT4 #(
		.INIT('h0777)
	) name6773 (
		_w8648_,
		_w8649_,
		_w8651_,
		_w8652_,
		_w8674_
	);
	LUT2 #(
		.INIT('h8)
	) name6774 (
		\m7_s4_cyc_o_reg/NET0131 ,
		\s4_m7_cyc_r_reg/P0001 ,
		_w8675_
	);
	LUT3 #(
		.INIT('h70)
	) name6775 (
		_w8655_,
		_w8656_,
		_w8675_,
		_w8676_
	);
	LUT2 #(
		.INIT('h8)
	) name6776 (
		\m6_s4_cyc_o_reg/NET0131 ,
		\s4_m6_cyc_r_reg/P0001 ,
		_w8677_
	);
	LUT3 #(
		.INIT('h80)
	) name6777 (
		_w8655_,
		_w8656_,
		_w8677_,
		_w8678_
	);
	LUT3 #(
		.INIT('h57)
	) name6778 (
		_w8674_,
		_w8676_,
		_w8678_,
		_w8679_
	);
	LUT4 #(
		.INIT('h8000)
	) name6779 (
		_w8661_,
		_w8667_,
		_w8673_,
		_w8679_,
		_w8680_
	);
	LUT4 #(
		.INIT('h7fff)
	) name6780 (
		_w8661_,
		_w8667_,
		_w8673_,
		_w8679_,
		_w8681_
	);
	LUT2 #(
		.INIT('h8)
	) name6781 (
		_w3569_,
		_w3579_,
		_w8682_
	);
	LUT3 #(
		.INIT('h80)
	) name6782 (
		\s10_next_reg/P0001 ,
		_w6665_,
		_w6671_,
		_w8683_
	);
	LUT2 #(
		.INIT('h8)
	) name6783 (
		_w3167_,
		_w3170_,
		_w8684_
	);
	LUT4 #(
		.INIT('hd111)
	) name6784 (
		\s10_msel_pri_out_reg[0]/NET0131 ,
		\s10_next_reg/P0001 ,
		_w3167_,
		_w3170_,
		_w8685_
	);
	LUT4 #(
		.INIT('h1055)
	) name6785 (
		rst_i_pad,
		_w8682_,
		_w8683_,
		_w8685_,
		_w8686_
	);
	LUT2 #(
		.INIT('h8)
	) name6786 (
		_w3592_,
		_w3608_,
		_w8687_
	);
	LUT3 #(
		.INIT('h80)
	) name6787 (
		\s11_next_reg/P0001 ,
		_w3188_,
		_w3199_,
		_w8688_
	);
	LUT2 #(
		.INIT('h8)
	) name6788 (
		_w3210_,
		_w3221_,
		_w8689_
	);
	LUT4 #(
		.INIT('hd111)
	) name6789 (
		\s11_msel_pri_out_reg[0]/NET0131 ,
		\s11_next_reg/P0001 ,
		_w3210_,
		_w3221_,
		_w8690_
	);
	LUT4 #(
		.INIT('h1055)
	) name6790 (
		rst_i_pad,
		_w8687_,
		_w8688_,
		_w8690_,
		_w8691_
	);
	LUT4 #(
		.INIT('hf35f)
	) name6791 (
		\s5_msel_arb1_state_reg[1]/NET0131 ,
		\s5_msel_arb2_state_reg[1]/NET0131 ,
		\s5_msel_pri_out_reg[0]/NET0131 ,
		\s5_msel_pri_out_reg[1]/NET0131 ,
		_w8692_
	);
	LUT4 #(
		.INIT('h3ff5)
	) name6792 (
		\s5_msel_arb0_state_reg[1]/NET0131 ,
		\s5_msel_arb3_state_reg[1]/NET0131 ,
		\s5_msel_pri_out_reg[0]/NET0131 ,
		\s5_msel_pri_out_reg[1]/NET0131 ,
		_w8693_
	);
	LUT2 #(
		.INIT('h8)
	) name6793 (
		_w8692_,
		_w8693_,
		_w8694_
	);
	LUT4 #(
		.INIT('hf35f)
	) name6794 (
		\s5_msel_arb1_state_reg[2]/NET0131 ,
		\s5_msel_arb2_state_reg[2]/NET0131 ,
		\s5_msel_pri_out_reg[0]/NET0131 ,
		\s5_msel_pri_out_reg[1]/NET0131 ,
		_w8695_
	);
	LUT4 #(
		.INIT('h3ff5)
	) name6795 (
		\s5_msel_arb0_state_reg[2]/NET0131 ,
		\s5_msel_arb3_state_reg[2]/NET0131 ,
		\s5_msel_pri_out_reg[0]/NET0131 ,
		\s5_msel_pri_out_reg[1]/NET0131 ,
		_w8696_
	);
	LUT2 #(
		.INIT('h8)
	) name6796 (
		_w8695_,
		_w8696_,
		_w8697_
	);
	LUT4 #(
		.INIT('h7000)
	) name6797 (
		_w8692_,
		_w8693_,
		_w8695_,
		_w8696_,
		_w8698_
	);
	LUT4 #(
		.INIT('hf35f)
	) name6798 (
		\s5_msel_arb1_state_reg[0]/NET0131 ,
		\s5_msel_arb2_state_reg[0]/NET0131 ,
		\s5_msel_pri_out_reg[0]/NET0131 ,
		\s5_msel_pri_out_reg[1]/NET0131 ,
		_w8699_
	);
	LUT4 #(
		.INIT('h3ff5)
	) name6799 (
		\s5_msel_arb0_state_reg[0]/NET0131 ,
		\s5_msel_arb3_state_reg[0]/NET0131 ,
		\s5_msel_pri_out_reg[0]/NET0131 ,
		\s5_msel_pri_out_reg[1]/NET0131 ,
		_w8700_
	);
	LUT2 #(
		.INIT('h8)
	) name6800 (
		\m3_s5_cyc_o_reg/NET0131 ,
		\s5_m3_cyc_r_reg/P0001 ,
		_w8701_
	);
	LUT3 #(
		.INIT('h70)
	) name6801 (
		_w8699_,
		_w8700_,
		_w8701_,
		_w8702_
	);
	LUT2 #(
		.INIT('h8)
	) name6802 (
		\m2_s5_cyc_o_reg/NET0131 ,
		\s5_m2_cyc_r_reg/P0001 ,
		_w8703_
	);
	LUT3 #(
		.INIT('h80)
	) name6803 (
		_w8699_,
		_w8700_,
		_w8703_,
		_w8704_
	);
	LUT3 #(
		.INIT('h57)
	) name6804 (
		_w8698_,
		_w8702_,
		_w8704_,
		_w8705_
	);
	LUT4 #(
		.INIT('h0888)
	) name6805 (
		_w8692_,
		_w8693_,
		_w8695_,
		_w8696_,
		_w8706_
	);
	LUT2 #(
		.INIT('h8)
	) name6806 (
		\m5_s5_cyc_o_reg/NET0131 ,
		\s5_m5_cyc_r_reg/P0001 ,
		_w8707_
	);
	LUT3 #(
		.INIT('h70)
	) name6807 (
		_w8699_,
		_w8700_,
		_w8707_,
		_w8708_
	);
	LUT2 #(
		.INIT('h8)
	) name6808 (
		\m4_s5_cyc_o_reg/NET0131 ,
		\s5_m4_cyc_r_reg/P0001 ,
		_w8709_
	);
	LUT3 #(
		.INIT('h80)
	) name6809 (
		_w8699_,
		_w8700_,
		_w8709_,
		_w8710_
	);
	LUT3 #(
		.INIT('h57)
	) name6810 (
		_w8706_,
		_w8708_,
		_w8710_,
		_w8711_
	);
	LUT4 #(
		.INIT('h0777)
	) name6811 (
		_w8692_,
		_w8693_,
		_w8695_,
		_w8696_,
		_w8712_
	);
	LUT2 #(
		.INIT('h8)
	) name6812 (
		\m7_s5_cyc_o_reg/NET0131 ,
		\s5_m7_cyc_r_reg/P0001 ,
		_w8713_
	);
	LUT3 #(
		.INIT('h70)
	) name6813 (
		_w8699_,
		_w8700_,
		_w8713_,
		_w8714_
	);
	LUT2 #(
		.INIT('h8)
	) name6814 (
		\m6_s5_cyc_o_reg/NET0131 ,
		\s5_m6_cyc_r_reg/P0001 ,
		_w8715_
	);
	LUT3 #(
		.INIT('h80)
	) name6815 (
		_w8699_,
		_w8700_,
		_w8715_,
		_w8716_
	);
	LUT3 #(
		.INIT('h57)
	) name6816 (
		_w8712_,
		_w8714_,
		_w8716_,
		_w8717_
	);
	LUT4 #(
		.INIT('h8000)
	) name6817 (
		_w8692_,
		_w8693_,
		_w8695_,
		_w8696_,
		_w8718_
	);
	LUT2 #(
		.INIT('h8)
	) name6818 (
		\m1_s5_cyc_o_reg/NET0131 ,
		\s5_m1_cyc_r_reg/P0001 ,
		_w8719_
	);
	LUT3 #(
		.INIT('h70)
	) name6819 (
		_w8699_,
		_w8700_,
		_w8719_,
		_w8720_
	);
	LUT2 #(
		.INIT('h8)
	) name6820 (
		\m0_s5_cyc_o_reg/NET0131 ,
		\s5_m0_cyc_r_reg/P0001 ,
		_w8721_
	);
	LUT3 #(
		.INIT('h80)
	) name6821 (
		_w8699_,
		_w8700_,
		_w8721_,
		_w8722_
	);
	LUT3 #(
		.INIT('h57)
	) name6822 (
		_w8718_,
		_w8720_,
		_w8722_,
		_w8723_
	);
	LUT4 #(
		.INIT('h8000)
	) name6823 (
		_w8705_,
		_w8711_,
		_w8717_,
		_w8723_,
		_w8724_
	);
	LUT4 #(
		.INIT('h7fff)
	) name6824 (
		_w8705_,
		_w8711_,
		_w8717_,
		_w8723_,
		_w8725_
	);
	LUT2 #(
		.INIT('h8)
	) name6825 (
		_w3628_,
		_w3642_,
		_w8726_
	);
	LUT3 #(
		.INIT('h80)
	) name6826 (
		\s12_next_reg/P0001 ,
		_w6683_,
		_w6689_,
		_w8727_
	);
	LUT2 #(
		.INIT('h8)
	) name6827 (
		_w3251_,
		_w3254_,
		_w8728_
	);
	LUT4 #(
		.INIT('hd111)
	) name6828 (
		\s12_msel_pri_out_reg[0]/NET0131 ,
		\s12_next_reg/P0001 ,
		_w3251_,
		_w3254_,
		_w8729_
	);
	LUT4 #(
		.INIT('h1055)
	) name6829 (
		rst_i_pad,
		_w8726_,
		_w8727_,
		_w8729_,
		_w8730_
	);
	LUT2 #(
		.INIT('h8)
	) name6830 (
		_w3655_,
		_w3665_,
		_w8731_
	);
	LUT3 #(
		.INIT('h80)
	) name6831 (
		\s13_next_reg/P0001 ,
		_w6700_,
		_w6708_,
		_w8732_
	);
	LUT2 #(
		.INIT('h8)
	) name6832 (
		_w2957_,
		_w2960_,
		_w8733_
	);
	LUT4 #(
		.INIT('hd111)
	) name6833 (
		\s13_msel_pri_out_reg[0]/NET0131 ,
		\s13_next_reg/P0001 ,
		_w2957_,
		_w2960_,
		_w8734_
	);
	LUT4 #(
		.INIT('h1055)
	) name6834 (
		rst_i_pad,
		_w8731_,
		_w8732_,
		_w8734_,
		_w8735_
	);
	LUT4 #(
		.INIT('h3ff5)
	) name6835 (
		\s6_msel_arb0_state_reg[1]/NET0131 ,
		\s6_msel_arb3_state_reg[1]/NET0131 ,
		\s6_msel_pri_out_reg[0]/NET0131 ,
		\s6_msel_pri_out_reg[1]/NET0131 ,
		_w8736_
	);
	LUT4 #(
		.INIT('hf35f)
	) name6836 (
		\s6_msel_arb1_state_reg[1]/NET0131 ,
		\s6_msel_arb2_state_reg[1]/NET0131 ,
		\s6_msel_pri_out_reg[0]/NET0131 ,
		\s6_msel_pri_out_reg[1]/NET0131 ,
		_w8737_
	);
	LUT2 #(
		.INIT('h8)
	) name6837 (
		_w8736_,
		_w8737_,
		_w8738_
	);
	LUT4 #(
		.INIT('h3ff5)
	) name6838 (
		\s6_msel_arb0_state_reg[2]/NET0131 ,
		\s6_msel_arb3_state_reg[2]/NET0131 ,
		\s6_msel_pri_out_reg[0]/NET0131 ,
		\s6_msel_pri_out_reg[1]/NET0131 ,
		_w8739_
	);
	LUT4 #(
		.INIT('hf35f)
	) name6839 (
		\s6_msel_arb1_state_reg[2]/NET0131 ,
		\s6_msel_arb2_state_reg[2]/NET0131 ,
		\s6_msel_pri_out_reg[0]/NET0131 ,
		\s6_msel_pri_out_reg[1]/NET0131 ,
		_w8740_
	);
	LUT2 #(
		.INIT('h8)
	) name6840 (
		_w8739_,
		_w8740_,
		_w8741_
	);
	LUT4 #(
		.INIT('h8000)
	) name6841 (
		_w8736_,
		_w8737_,
		_w8739_,
		_w8740_,
		_w8742_
	);
	LUT4 #(
		.INIT('hf3f5)
	) name6842 (
		\s6_msel_arb0_state_reg[0]/NET0131 ,
		\s6_msel_arb2_state_reg[0]/NET0131 ,
		\s6_msel_pri_out_reg[0]/NET0131 ,
		\s6_msel_pri_out_reg[1]/NET0131 ,
		_w8743_
	);
	LUT4 #(
		.INIT('h3f5f)
	) name6843 (
		\s6_msel_arb1_state_reg[0]/NET0131 ,
		\s6_msel_arb3_state_reg[0]/NET0131 ,
		\s6_msel_pri_out_reg[0]/NET0131 ,
		\s6_msel_pri_out_reg[1]/NET0131 ,
		_w8744_
	);
	LUT2 #(
		.INIT('h8)
	) name6844 (
		\m1_s6_cyc_o_reg/NET0131 ,
		\s6_m1_cyc_r_reg/P0001 ,
		_w8745_
	);
	LUT3 #(
		.INIT('h70)
	) name6845 (
		_w8743_,
		_w8744_,
		_w8745_,
		_w8746_
	);
	LUT2 #(
		.INIT('h8)
	) name6846 (
		\m0_s6_cyc_o_reg/NET0131 ,
		\s6_m0_cyc_r_reg/P0001 ,
		_w8747_
	);
	LUT3 #(
		.INIT('h80)
	) name6847 (
		_w8743_,
		_w8744_,
		_w8747_,
		_w8748_
	);
	LUT3 #(
		.INIT('h57)
	) name6848 (
		_w8742_,
		_w8746_,
		_w8748_,
		_w8749_
	);
	LUT4 #(
		.INIT('h7000)
	) name6849 (
		_w8736_,
		_w8737_,
		_w8739_,
		_w8740_,
		_w8750_
	);
	LUT2 #(
		.INIT('h8)
	) name6850 (
		\m3_s6_cyc_o_reg/NET0131 ,
		\s6_m3_cyc_r_reg/P0001 ,
		_w8751_
	);
	LUT3 #(
		.INIT('h70)
	) name6851 (
		_w8743_,
		_w8744_,
		_w8751_,
		_w8752_
	);
	LUT2 #(
		.INIT('h8)
	) name6852 (
		\m2_s6_cyc_o_reg/NET0131 ,
		\s6_m2_cyc_r_reg/P0001 ,
		_w8753_
	);
	LUT3 #(
		.INIT('h80)
	) name6853 (
		_w8743_,
		_w8744_,
		_w8753_,
		_w8754_
	);
	LUT3 #(
		.INIT('h57)
	) name6854 (
		_w8750_,
		_w8752_,
		_w8754_,
		_w8755_
	);
	LUT4 #(
		.INIT('h0777)
	) name6855 (
		_w8736_,
		_w8737_,
		_w8739_,
		_w8740_,
		_w8756_
	);
	LUT2 #(
		.INIT('h8)
	) name6856 (
		\m7_s6_cyc_o_reg/NET0131 ,
		\s6_m7_cyc_r_reg/P0001 ,
		_w8757_
	);
	LUT3 #(
		.INIT('h70)
	) name6857 (
		_w8743_,
		_w8744_,
		_w8757_,
		_w8758_
	);
	LUT2 #(
		.INIT('h8)
	) name6858 (
		\m6_s6_cyc_o_reg/NET0131 ,
		\s6_m6_cyc_r_reg/P0001 ,
		_w8759_
	);
	LUT3 #(
		.INIT('h80)
	) name6859 (
		_w8743_,
		_w8744_,
		_w8759_,
		_w8760_
	);
	LUT3 #(
		.INIT('h57)
	) name6860 (
		_w8756_,
		_w8758_,
		_w8760_,
		_w8761_
	);
	LUT4 #(
		.INIT('h0888)
	) name6861 (
		_w8736_,
		_w8737_,
		_w8739_,
		_w8740_,
		_w8762_
	);
	LUT2 #(
		.INIT('h8)
	) name6862 (
		\m5_s6_cyc_o_reg/NET0131 ,
		\s6_m5_cyc_r_reg/P0001 ,
		_w8763_
	);
	LUT3 #(
		.INIT('h70)
	) name6863 (
		_w8743_,
		_w8744_,
		_w8763_,
		_w8764_
	);
	LUT2 #(
		.INIT('h8)
	) name6864 (
		\m4_s6_cyc_o_reg/NET0131 ,
		\s6_m4_cyc_r_reg/P0001 ,
		_w8765_
	);
	LUT3 #(
		.INIT('h80)
	) name6865 (
		_w8743_,
		_w8744_,
		_w8765_,
		_w8766_
	);
	LUT3 #(
		.INIT('h57)
	) name6866 (
		_w8762_,
		_w8764_,
		_w8766_,
		_w8767_
	);
	LUT4 #(
		.INIT('h8000)
	) name6867 (
		_w8749_,
		_w8755_,
		_w8761_,
		_w8767_,
		_w8768_
	);
	LUT4 #(
		.INIT('h7fff)
	) name6868 (
		_w8749_,
		_w8755_,
		_w8761_,
		_w8767_,
		_w8769_
	);
	LUT2 #(
		.INIT('h8)
	) name6869 (
		_w3675_,
		_w3690_,
		_w8770_
	);
	LUT3 #(
		.INIT('h80)
	) name6870 (
		\s14_next_reg/P0001 ,
		_w2987_,
		_w2990_,
		_w8771_
	);
	LUT2 #(
		.INIT('h8)
	) name6871 (
		_w3272_,
		_w3283_,
		_w8772_
	);
	LUT4 #(
		.INIT('hd111)
	) name6872 (
		\s14_msel_pri_out_reg[0]/NET0131 ,
		\s14_next_reg/P0001 ,
		_w3272_,
		_w3283_,
		_w8773_
	);
	LUT4 #(
		.INIT('h1055)
	) name6873 (
		rst_i_pad,
		_w8770_,
		_w8771_,
		_w8773_,
		_w8774_
	);
	LUT4 #(
		.INIT('h3ff5)
	) name6874 (
		\s7_msel_arb0_state_reg[1]/NET0131 ,
		\s7_msel_arb3_state_reg[1]/NET0131 ,
		\s7_msel_pri_out_reg[0]/NET0131 ,
		\s7_msel_pri_out_reg[1]/NET0131 ,
		_w8775_
	);
	LUT4 #(
		.INIT('hf35f)
	) name6875 (
		\s7_msel_arb1_state_reg[1]/NET0131 ,
		\s7_msel_arb2_state_reg[1]/NET0131 ,
		\s7_msel_pri_out_reg[0]/NET0131 ,
		\s7_msel_pri_out_reg[1]/NET0131 ,
		_w8776_
	);
	LUT2 #(
		.INIT('h8)
	) name6876 (
		_w8775_,
		_w8776_,
		_w8777_
	);
	LUT4 #(
		.INIT('hf35f)
	) name6877 (
		\s7_msel_arb1_state_reg[2]/NET0131 ,
		\s7_msel_arb2_state_reg[2]/NET0131 ,
		\s7_msel_pri_out_reg[0]/NET0131 ,
		\s7_msel_pri_out_reg[1]/NET0131 ,
		_w8778_
	);
	LUT4 #(
		.INIT('h3ff5)
	) name6878 (
		\s7_msel_arb0_state_reg[2]/NET0131 ,
		\s7_msel_arb3_state_reg[2]/NET0131 ,
		\s7_msel_pri_out_reg[0]/NET0131 ,
		\s7_msel_pri_out_reg[1]/NET0131 ,
		_w8779_
	);
	LUT2 #(
		.INIT('h8)
	) name6879 (
		_w8778_,
		_w8779_,
		_w8780_
	);
	LUT4 #(
		.INIT('h0777)
	) name6880 (
		_w8775_,
		_w8776_,
		_w8778_,
		_w8779_,
		_w8781_
	);
	LUT4 #(
		.INIT('hf35f)
	) name6881 (
		\s7_msel_arb1_state_reg[0]/NET0131 ,
		\s7_msel_arb2_state_reg[0]/NET0131 ,
		\s7_msel_pri_out_reg[0]/NET0131 ,
		\s7_msel_pri_out_reg[1]/NET0131 ,
		_w8782_
	);
	LUT4 #(
		.INIT('h3ff5)
	) name6882 (
		\s7_msel_arb0_state_reg[0]/NET0131 ,
		\s7_msel_arb3_state_reg[0]/NET0131 ,
		\s7_msel_pri_out_reg[0]/NET0131 ,
		\s7_msel_pri_out_reg[1]/NET0131 ,
		_w8783_
	);
	LUT2 #(
		.INIT('h8)
	) name6883 (
		\m7_s7_cyc_o_reg/NET0131 ,
		\s7_m7_cyc_r_reg/P0001 ,
		_w8784_
	);
	LUT3 #(
		.INIT('h70)
	) name6884 (
		_w8782_,
		_w8783_,
		_w8784_,
		_w8785_
	);
	LUT2 #(
		.INIT('h8)
	) name6885 (
		\m6_s7_cyc_o_reg/NET0131 ,
		\s7_m6_cyc_r_reg/P0001 ,
		_w8786_
	);
	LUT3 #(
		.INIT('h80)
	) name6886 (
		_w8782_,
		_w8783_,
		_w8786_,
		_w8787_
	);
	LUT3 #(
		.INIT('h57)
	) name6887 (
		_w8781_,
		_w8785_,
		_w8787_,
		_w8788_
	);
	LUT4 #(
		.INIT('h8000)
	) name6888 (
		_w8775_,
		_w8776_,
		_w8778_,
		_w8779_,
		_w8789_
	);
	LUT2 #(
		.INIT('h8)
	) name6889 (
		\m1_s7_cyc_o_reg/NET0131 ,
		\s7_m1_cyc_r_reg/P0001 ,
		_w8790_
	);
	LUT3 #(
		.INIT('h70)
	) name6890 (
		_w8782_,
		_w8783_,
		_w8790_,
		_w8791_
	);
	LUT2 #(
		.INIT('h8)
	) name6891 (
		\m0_s7_cyc_o_reg/NET0131 ,
		\s7_m0_cyc_r_reg/P0001 ,
		_w8792_
	);
	LUT3 #(
		.INIT('h80)
	) name6892 (
		_w8782_,
		_w8783_,
		_w8792_,
		_w8793_
	);
	LUT3 #(
		.INIT('h57)
	) name6893 (
		_w8789_,
		_w8791_,
		_w8793_,
		_w8794_
	);
	LUT4 #(
		.INIT('h7000)
	) name6894 (
		_w8775_,
		_w8776_,
		_w8778_,
		_w8779_,
		_w8795_
	);
	LUT2 #(
		.INIT('h8)
	) name6895 (
		\m3_s7_cyc_o_reg/NET0131 ,
		\s7_m3_cyc_r_reg/P0001 ,
		_w8796_
	);
	LUT3 #(
		.INIT('h70)
	) name6896 (
		_w8782_,
		_w8783_,
		_w8796_,
		_w8797_
	);
	LUT2 #(
		.INIT('h8)
	) name6897 (
		\m2_s7_cyc_o_reg/NET0131 ,
		\s7_m2_cyc_r_reg/P0001 ,
		_w8798_
	);
	LUT3 #(
		.INIT('h80)
	) name6898 (
		_w8782_,
		_w8783_,
		_w8798_,
		_w8799_
	);
	LUT3 #(
		.INIT('h57)
	) name6899 (
		_w8795_,
		_w8797_,
		_w8799_,
		_w8800_
	);
	LUT4 #(
		.INIT('h0888)
	) name6900 (
		_w8775_,
		_w8776_,
		_w8778_,
		_w8779_,
		_w8801_
	);
	LUT2 #(
		.INIT('h8)
	) name6901 (
		\m5_s7_cyc_o_reg/NET0131 ,
		\s7_m5_cyc_r_reg/P0001 ,
		_w8802_
	);
	LUT3 #(
		.INIT('h70)
	) name6902 (
		_w8782_,
		_w8783_,
		_w8802_,
		_w8803_
	);
	LUT2 #(
		.INIT('h8)
	) name6903 (
		\m4_s7_cyc_o_reg/NET0131 ,
		\s7_m4_cyc_r_reg/P0001 ,
		_w8804_
	);
	LUT3 #(
		.INIT('h80)
	) name6904 (
		_w8782_,
		_w8783_,
		_w8804_,
		_w8805_
	);
	LUT3 #(
		.INIT('h57)
	) name6905 (
		_w8801_,
		_w8803_,
		_w8805_,
		_w8806_
	);
	LUT4 #(
		.INIT('h8000)
	) name6906 (
		_w8788_,
		_w8794_,
		_w8800_,
		_w8806_,
		_w8807_
	);
	LUT4 #(
		.INIT('h7fff)
	) name6907 (
		_w8788_,
		_w8794_,
		_w8800_,
		_w8806_,
		_w8808_
	);
	LUT2 #(
		.INIT('h8)
	) name6908 (
		_w3701_,
		_w3716_,
		_w8809_
	);
	LUT3 #(
		.INIT('h80)
	) name6909 (
		\s1_next_reg/P0001 ,
		_w3304_,
		_w3315_,
		_w8810_
	);
	LUT2 #(
		.INIT('h8)
	) name6910 (
		_w3326_,
		_w3337_,
		_w8811_
	);
	LUT4 #(
		.INIT('hd111)
	) name6911 (
		\s1_msel_pri_out_reg[0]/NET0131 ,
		\s1_next_reg/P0001 ,
		_w3326_,
		_w3337_,
		_w8812_
	);
	LUT4 #(
		.INIT('h1055)
	) name6912 (
		rst_i_pad,
		_w8809_,
		_w8810_,
		_w8812_,
		_w8813_
	);
	LUT4 #(
		.INIT('hf35f)
	) name6913 (
		\s8_msel_arb1_state_reg[1]/NET0131 ,
		\s8_msel_arb2_state_reg[1]/NET0131 ,
		\s8_msel_pri_out_reg[0]/NET0131 ,
		\s8_msel_pri_out_reg[1]/NET0131 ,
		_w8814_
	);
	LUT4 #(
		.INIT('h3ff5)
	) name6914 (
		\s8_msel_arb0_state_reg[1]/NET0131 ,
		\s8_msel_arb3_state_reg[1]/NET0131 ,
		\s8_msel_pri_out_reg[0]/NET0131 ,
		\s8_msel_pri_out_reg[1]/NET0131 ,
		_w8815_
	);
	LUT2 #(
		.INIT('h8)
	) name6915 (
		_w8814_,
		_w8815_,
		_w8816_
	);
	LUT4 #(
		.INIT('hf35f)
	) name6916 (
		\s8_msel_arb1_state_reg[2]/NET0131 ,
		\s8_msel_arb2_state_reg[2]/NET0131 ,
		\s8_msel_pri_out_reg[0]/NET0131 ,
		\s8_msel_pri_out_reg[1]/NET0131 ,
		_w8817_
	);
	LUT4 #(
		.INIT('h3ff5)
	) name6917 (
		\s8_msel_arb0_state_reg[2]/NET0131 ,
		\s8_msel_arb3_state_reg[2]/NET0131 ,
		\s8_msel_pri_out_reg[0]/NET0131 ,
		\s8_msel_pri_out_reg[1]/NET0131 ,
		_w8818_
	);
	LUT2 #(
		.INIT('h8)
	) name6918 (
		_w8817_,
		_w8818_,
		_w8819_
	);
	LUT4 #(
		.INIT('h8000)
	) name6919 (
		_w8814_,
		_w8815_,
		_w8817_,
		_w8818_,
		_w8820_
	);
	LUT4 #(
		.INIT('hf35f)
	) name6920 (
		\s8_msel_arb1_state_reg[0]/NET0131 ,
		\s8_msel_arb2_state_reg[0]/NET0131 ,
		\s8_msel_pri_out_reg[0]/NET0131 ,
		\s8_msel_pri_out_reg[1]/NET0131 ,
		_w8821_
	);
	LUT4 #(
		.INIT('h3ff5)
	) name6921 (
		\s8_msel_arb0_state_reg[0]/NET0131 ,
		\s8_msel_arb3_state_reg[0]/NET0131 ,
		\s8_msel_pri_out_reg[0]/NET0131 ,
		\s8_msel_pri_out_reg[1]/NET0131 ,
		_w8822_
	);
	LUT2 #(
		.INIT('h8)
	) name6922 (
		\m1_s8_cyc_o_reg/NET0131 ,
		\s8_m1_cyc_r_reg/P0001 ,
		_w8823_
	);
	LUT3 #(
		.INIT('h70)
	) name6923 (
		_w8821_,
		_w8822_,
		_w8823_,
		_w8824_
	);
	LUT2 #(
		.INIT('h8)
	) name6924 (
		\m0_s8_cyc_o_reg/NET0131 ,
		\s8_m0_cyc_r_reg/P0001 ,
		_w8825_
	);
	LUT3 #(
		.INIT('h80)
	) name6925 (
		_w8821_,
		_w8822_,
		_w8825_,
		_w8826_
	);
	LUT3 #(
		.INIT('h57)
	) name6926 (
		_w8820_,
		_w8824_,
		_w8826_,
		_w8827_
	);
	LUT4 #(
		.INIT('h7000)
	) name6927 (
		_w8814_,
		_w8815_,
		_w8817_,
		_w8818_,
		_w8828_
	);
	LUT2 #(
		.INIT('h8)
	) name6928 (
		\m3_s8_cyc_o_reg/NET0131 ,
		\s8_m3_cyc_r_reg/P0001 ,
		_w8829_
	);
	LUT3 #(
		.INIT('h70)
	) name6929 (
		_w8821_,
		_w8822_,
		_w8829_,
		_w8830_
	);
	LUT2 #(
		.INIT('h8)
	) name6930 (
		\m2_s8_cyc_o_reg/NET0131 ,
		\s8_m2_cyc_r_reg/P0001 ,
		_w8831_
	);
	LUT3 #(
		.INIT('h80)
	) name6931 (
		_w8821_,
		_w8822_,
		_w8831_,
		_w8832_
	);
	LUT3 #(
		.INIT('h57)
	) name6932 (
		_w8828_,
		_w8830_,
		_w8832_,
		_w8833_
	);
	LUT4 #(
		.INIT('h0777)
	) name6933 (
		_w8814_,
		_w8815_,
		_w8817_,
		_w8818_,
		_w8834_
	);
	LUT2 #(
		.INIT('h8)
	) name6934 (
		\m7_s8_cyc_o_reg/NET0131 ,
		\s8_m7_cyc_r_reg/P0001 ,
		_w8835_
	);
	LUT3 #(
		.INIT('h70)
	) name6935 (
		_w8821_,
		_w8822_,
		_w8835_,
		_w8836_
	);
	LUT2 #(
		.INIT('h8)
	) name6936 (
		\m6_s8_cyc_o_reg/NET0131 ,
		\s8_m6_cyc_r_reg/P0001 ,
		_w8837_
	);
	LUT3 #(
		.INIT('h80)
	) name6937 (
		_w8821_,
		_w8822_,
		_w8837_,
		_w8838_
	);
	LUT3 #(
		.INIT('h57)
	) name6938 (
		_w8834_,
		_w8836_,
		_w8838_,
		_w8839_
	);
	LUT4 #(
		.INIT('h0888)
	) name6939 (
		_w8814_,
		_w8815_,
		_w8817_,
		_w8818_,
		_w8840_
	);
	LUT2 #(
		.INIT('h8)
	) name6940 (
		\m5_s8_cyc_o_reg/NET0131 ,
		\s8_m5_cyc_r_reg/P0001 ,
		_w8841_
	);
	LUT3 #(
		.INIT('h70)
	) name6941 (
		_w8821_,
		_w8822_,
		_w8841_,
		_w8842_
	);
	LUT2 #(
		.INIT('h8)
	) name6942 (
		\m4_s8_cyc_o_reg/NET0131 ,
		\s8_m4_cyc_r_reg/P0001 ,
		_w8843_
	);
	LUT3 #(
		.INIT('h80)
	) name6943 (
		_w8821_,
		_w8822_,
		_w8843_,
		_w8844_
	);
	LUT3 #(
		.INIT('h57)
	) name6944 (
		_w8840_,
		_w8842_,
		_w8844_,
		_w8845_
	);
	LUT4 #(
		.INIT('h8000)
	) name6945 (
		_w8827_,
		_w8833_,
		_w8839_,
		_w8845_,
		_w8846_
	);
	LUT4 #(
		.INIT('h7fff)
	) name6946 (
		_w8827_,
		_w8833_,
		_w8839_,
		_w8845_,
		_w8847_
	);
	LUT2 #(
		.INIT('h8)
	) name6947 (
		_w3732_,
		_w3742_,
		_w8848_
	);
	LUT3 #(
		.INIT('h80)
	) name6948 (
		\s2_next_reg/P0001 ,
		_w6715_,
		_w6723_,
		_w8849_
	);
	LUT2 #(
		.INIT('h8)
	) name6949 (
		_w3017_,
		_w3020_,
		_w8850_
	);
	LUT4 #(
		.INIT('hd111)
	) name6950 (
		\s2_msel_pri_out_reg[0]/NET0131 ,
		\s2_next_reg/P0001 ,
		_w3017_,
		_w3020_,
		_w8851_
	);
	LUT4 #(
		.INIT('h1055)
	) name6951 (
		rst_i_pad,
		_w8848_,
		_w8849_,
		_w8851_,
		_w8852_
	);
	LUT2 #(
		.INIT('h8)
	) name6952 (
		_w3755_,
		_w3771_,
		_w8853_
	);
	LUT3 #(
		.INIT('h80)
	) name6953 (
		\s3_next_reg/P0001 ,
		_w3038_,
		_w3049_,
		_w8854_
	);
	LUT2 #(
		.INIT('h8)
	) name6954 (
		_w3358_,
		_w3369_,
		_w8855_
	);
	LUT4 #(
		.INIT('hd111)
	) name6955 (
		\s3_msel_pri_out_reg[0]/NET0131 ,
		\s3_next_reg/P0001 ,
		_w3358_,
		_w3369_,
		_w8856_
	);
	LUT4 #(
		.INIT('h1055)
	) name6956 (
		rst_i_pad,
		_w8853_,
		_w8854_,
		_w8856_,
		_w8857_
	);
	LUT4 #(
		.INIT('hf35f)
	) name6957 (
		\s9_msel_arb1_state_reg[1]/NET0131 ,
		\s9_msel_arb2_state_reg[1]/NET0131 ,
		\s9_msel_pri_out_reg[0]/NET0131 ,
		\s9_msel_pri_out_reg[1]/NET0131 ,
		_w8858_
	);
	LUT4 #(
		.INIT('h3ff5)
	) name6958 (
		\s9_msel_arb0_state_reg[1]/NET0131 ,
		\s9_msel_arb3_state_reg[1]/NET0131 ,
		\s9_msel_pri_out_reg[0]/NET0131 ,
		\s9_msel_pri_out_reg[1]/NET0131 ,
		_w8859_
	);
	LUT2 #(
		.INIT('h8)
	) name6959 (
		_w8858_,
		_w8859_,
		_w8860_
	);
	LUT4 #(
		.INIT('hf35f)
	) name6960 (
		\s9_msel_arb1_state_reg[2]/NET0131 ,
		\s9_msel_arb2_state_reg[2]/NET0131 ,
		\s9_msel_pri_out_reg[0]/NET0131 ,
		\s9_msel_pri_out_reg[1]/NET0131 ,
		_w8861_
	);
	LUT4 #(
		.INIT('h3ff5)
	) name6961 (
		\s9_msel_arb0_state_reg[2]/NET0131 ,
		\s9_msel_arb3_state_reg[2]/NET0131 ,
		\s9_msel_pri_out_reg[0]/NET0131 ,
		\s9_msel_pri_out_reg[1]/NET0131 ,
		_w8862_
	);
	LUT2 #(
		.INIT('h8)
	) name6962 (
		_w8861_,
		_w8862_,
		_w8863_
	);
	LUT4 #(
		.INIT('h7000)
	) name6963 (
		_w8858_,
		_w8859_,
		_w8861_,
		_w8862_,
		_w8864_
	);
	LUT4 #(
		.INIT('hf35f)
	) name6964 (
		\s9_msel_arb1_state_reg[0]/NET0131 ,
		\s9_msel_arb2_state_reg[0]/NET0131 ,
		\s9_msel_pri_out_reg[0]/NET0131 ,
		\s9_msel_pri_out_reg[1]/NET0131 ,
		_w8865_
	);
	LUT4 #(
		.INIT('h3ff5)
	) name6965 (
		\s9_msel_arb0_state_reg[0]/NET0131 ,
		\s9_msel_arb3_state_reg[0]/NET0131 ,
		\s9_msel_pri_out_reg[0]/NET0131 ,
		\s9_msel_pri_out_reg[1]/NET0131 ,
		_w8866_
	);
	LUT2 #(
		.INIT('h8)
	) name6966 (
		\m3_s9_cyc_o_reg/NET0131 ,
		\s9_m3_cyc_r_reg/P0001 ,
		_w8867_
	);
	LUT3 #(
		.INIT('h70)
	) name6967 (
		_w8865_,
		_w8866_,
		_w8867_,
		_w8868_
	);
	LUT2 #(
		.INIT('h8)
	) name6968 (
		\m2_s9_cyc_o_reg/NET0131 ,
		\s9_m2_cyc_r_reg/P0001 ,
		_w8869_
	);
	LUT3 #(
		.INIT('h80)
	) name6969 (
		_w8865_,
		_w8866_,
		_w8869_,
		_w8870_
	);
	LUT3 #(
		.INIT('h57)
	) name6970 (
		_w8864_,
		_w8868_,
		_w8870_,
		_w8871_
	);
	LUT4 #(
		.INIT('h8000)
	) name6971 (
		_w8858_,
		_w8859_,
		_w8861_,
		_w8862_,
		_w8872_
	);
	LUT2 #(
		.INIT('h8)
	) name6972 (
		\m1_s9_cyc_o_reg/NET0131 ,
		\s9_m1_cyc_r_reg/P0001 ,
		_w8873_
	);
	LUT3 #(
		.INIT('h70)
	) name6973 (
		_w8865_,
		_w8866_,
		_w8873_,
		_w8874_
	);
	LUT2 #(
		.INIT('h8)
	) name6974 (
		\m0_s9_cyc_o_reg/NET0131 ,
		\s9_m0_cyc_r_reg/P0001 ,
		_w8875_
	);
	LUT3 #(
		.INIT('h80)
	) name6975 (
		_w8865_,
		_w8866_,
		_w8875_,
		_w8876_
	);
	LUT3 #(
		.INIT('h57)
	) name6976 (
		_w8872_,
		_w8874_,
		_w8876_,
		_w8877_
	);
	LUT4 #(
		.INIT('h0777)
	) name6977 (
		_w8858_,
		_w8859_,
		_w8861_,
		_w8862_,
		_w8878_
	);
	LUT2 #(
		.INIT('h8)
	) name6978 (
		\m7_s9_cyc_o_reg/NET0131 ,
		\s9_m7_cyc_r_reg/P0001 ,
		_w8879_
	);
	LUT3 #(
		.INIT('h70)
	) name6979 (
		_w8865_,
		_w8866_,
		_w8879_,
		_w8880_
	);
	LUT2 #(
		.INIT('h8)
	) name6980 (
		\m6_s9_cyc_o_reg/NET0131 ,
		\s9_m6_cyc_r_reg/P0001 ,
		_w8881_
	);
	LUT3 #(
		.INIT('h80)
	) name6981 (
		_w8865_,
		_w8866_,
		_w8881_,
		_w8882_
	);
	LUT3 #(
		.INIT('h57)
	) name6982 (
		_w8878_,
		_w8880_,
		_w8882_,
		_w8883_
	);
	LUT4 #(
		.INIT('h0888)
	) name6983 (
		_w8858_,
		_w8859_,
		_w8861_,
		_w8862_,
		_w8884_
	);
	LUT2 #(
		.INIT('h8)
	) name6984 (
		\m5_s9_cyc_o_reg/NET0131 ,
		\s9_m5_cyc_r_reg/P0001 ,
		_w8885_
	);
	LUT3 #(
		.INIT('h70)
	) name6985 (
		_w8865_,
		_w8866_,
		_w8885_,
		_w8886_
	);
	LUT2 #(
		.INIT('h8)
	) name6986 (
		\m4_s9_cyc_o_reg/NET0131 ,
		\s9_m4_cyc_r_reg/P0001 ,
		_w8887_
	);
	LUT3 #(
		.INIT('h80)
	) name6987 (
		_w8865_,
		_w8866_,
		_w8887_,
		_w8888_
	);
	LUT3 #(
		.INIT('h57)
	) name6988 (
		_w8884_,
		_w8886_,
		_w8888_,
		_w8889_
	);
	LUT4 #(
		.INIT('h8000)
	) name6989 (
		_w8871_,
		_w8877_,
		_w8883_,
		_w8889_,
		_w8890_
	);
	LUT4 #(
		.INIT('h7fff)
	) name6990 (
		_w8871_,
		_w8877_,
		_w8883_,
		_w8889_,
		_w8891_
	);
	LUT2 #(
		.INIT('h8)
	) name6991 (
		_w3781_,
		_w3796_,
		_w8892_
	);
	LUT3 #(
		.INIT('h80)
	) name6992 (
		\s4_next_reg/P0001 ,
		_w6730_,
		_w6738_,
		_w8893_
	);
	LUT2 #(
		.INIT('h8)
	) name6993 (
		_w3060_,
		_w3071_,
		_w8894_
	);
	LUT4 #(
		.INIT('hd111)
	) name6994 (
		\s4_msel_pri_out_reg[0]/NET0131 ,
		\s4_next_reg/P0001 ,
		_w3060_,
		_w3071_,
		_w8895_
	);
	LUT4 #(
		.INIT('h1055)
	) name6995 (
		rst_i_pad,
		_w8892_,
		_w8893_,
		_w8895_,
		_w8896_
	);
	LUT3 #(
		.INIT('h80)
	) name6996 (
		\s5_next_reg/P0001 ,
		_w3390_,
		_w3401_,
		_w8897_
	);
	LUT4 #(
		.INIT('h0001)
	) name6997 (
		_w3802_,
		_w3803_,
		_w3805_,
		_w3806_,
		_w8898_
	);
	LUT2 #(
		.INIT('h8)
	) name6998 (
		_w3813_,
		_w8898_,
		_w8899_
	);
	LUT2 #(
		.INIT('h8)
	) name6999 (
		_w3421_,
		_w3424_,
		_w8900_
	);
	LUT4 #(
		.INIT('hd111)
	) name7000 (
		\s5_msel_pri_out_reg[0]/NET0131 ,
		\s5_next_reg/P0001 ,
		_w3421_,
		_w3424_,
		_w8901_
	);
	LUT4 #(
		.INIT('h0455)
	) name7001 (
		rst_i_pad,
		_w8897_,
		_w8899_,
		_w8901_,
		_w8902_
	);
	LUT4 #(
		.INIT('h3ff5)
	) name7002 (
		\s10_msel_arb0_state_reg[1]/NET0131 ,
		\s10_msel_arb3_state_reg[1]/NET0131 ,
		\s10_msel_pri_out_reg[0]/NET0131 ,
		\s10_msel_pri_out_reg[1]/NET0131 ,
		_w8903_
	);
	LUT4 #(
		.INIT('hf35f)
	) name7003 (
		\s10_msel_arb1_state_reg[1]/NET0131 ,
		\s10_msel_arb2_state_reg[1]/NET0131 ,
		\s10_msel_pri_out_reg[0]/NET0131 ,
		\s10_msel_pri_out_reg[1]/NET0131 ,
		_w8904_
	);
	LUT2 #(
		.INIT('h8)
	) name7004 (
		_w8903_,
		_w8904_,
		_w8905_
	);
	LUT4 #(
		.INIT('h3ff5)
	) name7005 (
		\s10_msel_arb0_state_reg[2]/NET0131 ,
		\s10_msel_arb3_state_reg[2]/NET0131 ,
		\s10_msel_pri_out_reg[0]/NET0131 ,
		\s10_msel_pri_out_reg[1]/NET0131 ,
		_w8906_
	);
	LUT4 #(
		.INIT('hf35f)
	) name7006 (
		\s10_msel_arb1_state_reg[2]/NET0131 ,
		\s10_msel_arb2_state_reg[2]/NET0131 ,
		\s10_msel_pri_out_reg[0]/NET0131 ,
		\s10_msel_pri_out_reg[1]/NET0131 ,
		_w8907_
	);
	LUT2 #(
		.INIT('h8)
	) name7007 (
		_w8906_,
		_w8907_,
		_w8908_
	);
	LUT4 #(
		.INIT('h7000)
	) name7008 (
		_w8903_,
		_w8904_,
		_w8906_,
		_w8907_,
		_w8909_
	);
	LUT4 #(
		.INIT('h3ff5)
	) name7009 (
		\s10_msel_arb0_state_reg[0]/NET0131 ,
		\s10_msel_arb3_state_reg[0]/NET0131 ,
		\s10_msel_pri_out_reg[0]/NET0131 ,
		\s10_msel_pri_out_reg[1]/NET0131 ,
		_w8910_
	);
	LUT4 #(
		.INIT('hf35f)
	) name7010 (
		\s10_msel_arb1_state_reg[0]/NET0131 ,
		\s10_msel_arb2_state_reg[0]/NET0131 ,
		\s10_msel_pri_out_reg[0]/NET0131 ,
		\s10_msel_pri_out_reg[1]/NET0131 ,
		_w8911_
	);
	LUT2 #(
		.INIT('h8)
	) name7011 (
		\m3_s10_cyc_o_reg/NET0131 ,
		\s10_m3_cyc_r_reg/P0001 ,
		_w8912_
	);
	LUT3 #(
		.INIT('h70)
	) name7012 (
		_w8910_,
		_w8911_,
		_w8912_,
		_w8913_
	);
	LUT2 #(
		.INIT('h8)
	) name7013 (
		\m2_s10_cyc_o_reg/NET0131 ,
		\s10_m2_cyc_r_reg/P0001 ,
		_w8914_
	);
	LUT3 #(
		.INIT('h80)
	) name7014 (
		_w8910_,
		_w8911_,
		_w8914_,
		_w8915_
	);
	LUT3 #(
		.INIT('h57)
	) name7015 (
		_w8909_,
		_w8913_,
		_w8915_,
		_w8916_
	);
	LUT4 #(
		.INIT('h0777)
	) name7016 (
		_w8903_,
		_w8904_,
		_w8906_,
		_w8907_,
		_w8917_
	);
	LUT2 #(
		.INIT('h8)
	) name7017 (
		\m7_s10_cyc_o_reg/NET0131 ,
		\s10_m7_cyc_r_reg/P0001 ,
		_w8918_
	);
	LUT3 #(
		.INIT('h70)
	) name7018 (
		_w8910_,
		_w8911_,
		_w8918_,
		_w8919_
	);
	LUT2 #(
		.INIT('h8)
	) name7019 (
		\m6_s10_cyc_o_reg/NET0131 ,
		\s10_m6_cyc_r_reg/P0001 ,
		_w8920_
	);
	LUT3 #(
		.INIT('h80)
	) name7020 (
		_w8910_,
		_w8911_,
		_w8920_,
		_w8921_
	);
	LUT3 #(
		.INIT('h57)
	) name7021 (
		_w8917_,
		_w8919_,
		_w8921_,
		_w8922_
	);
	LUT4 #(
		.INIT('h8000)
	) name7022 (
		_w8903_,
		_w8904_,
		_w8906_,
		_w8907_,
		_w8923_
	);
	LUT2 #(
		.INIT('h8)
	) name7023 (
		\m1_s10_cyc_o_reg/NET0131 ,
		\s10_m1_cyc_r_reg/P0001 ,
		_w8924_
	);
	LUT3 #(
		.INIT('h70)
	) name7024 (
		_w8910_,
		_w8911_,
		_w8924_,
		_w8925_
	);
	LUT2 #(
		.INIT('h8)
	) name7025 (
		\m0_s10_cyc_o_reg/NET0131 ,
		\s10_m0_cyc_r_reg/P0001 ,
		_w8926_
	);
	LUT3 #(
		.INIT('h80)
	) name7026 (
		_w8910_,
		_w8911_,
		_w8926_,
		_w8927_
	);
	LUT3 #(
		.INIT('h57)
	) name7027 (
		_w8923_,
		_w8925_,
		_w8927_,
		_w8928_
	);
	LUT4 #(
		.INIT('h0888)
	) name7028 (
		_w8903_,
		_w8904_,
		_w8906_,
		_w8907_,
		_w8929_
	);
	LUT2 #(
		.INIT('h8)
	) name7029 (
		\m5_s10_cyc_o_reg/NET0131 ,
		\s10_m5_cyc_r_reg/P0001 ,
		_w8930_
	);
	LUT3 #(
		.INIT('h70)
	) name7030 (
		_w8910_,
		_w8911_,
		_w8930_,
		_w8931_
	);
	LUT2 #(
		.INIT('h8)
	) name7031 (
		\m4_s10_cyc_o_reg/NET0131 ,
		\s10_m4_cyc_r_reg/P0001 ,
		_w8932_
	);
	LUT3 #(
		.INIT('h80)
	) name7032 (
		_w8910_,
		_w8911_,
		_w8932_,
		_w8933_
	);
	LUT3 #(
		.INIT('h57)
	) name7033 (
		_w8929_,
		_w8931_,
		_w8933_,
		_w8934_
	);
	LUT4 #(
		.INIT('h8000)
	) name7034 (
		_w8916_,
		_w8922_,
		_w8928_,
		_w8934_,
		_w8935_
	);
	LUT4 #(
		.INIT('h7fff)
	) name7035 (
		_w8916_,
		_w8922_,
		_w8928_,
		_w8934_,
		_w8936_
	);
	LUT3 #(
		.INIT('h80)
	) name7036 (
		\s6_next_reg/P0001 ,
		_w3092_,
		_w3103_,
		_w8937_
	);
	LUT4 #(
		.INIT('h0001)
	) name7037 (
		_w3833_,
		_w3834_,
		_w3836_,
		_w3837_,
		_w8938_
	);
	LUT2 #(
		.INIT('h8)
	) name7038 (
		_w3844_,
		_w8938_,
		_w8939_
	);
	LUT2 #(
		.INIT('h8)
	) name7039 (
		_w3451_,
		_w3454_,
		_w8940_
	);
	LUT4 #(
		.INIT('hd111)
	) name7040 (
		\s6_msel_pri_out_reg[0]/NET0131 ,
		\s6_next_reg/P0001 ,
		_w3451_,
		_w3454_,
		_w8941_
	);
	LUT4 #(
		.INIT('h0455)
	) name7041 (
		rst_i_pad,
		_w8937_,
		_w8939_,
		_w8941_,
		_w8942_
	);
	LUT2 #(
		.INIT('h8)
	) name7042 (
		_w3870_,
		_w3876_,
		_w8943_
	);
	LUT3 #(
		.INIT('h80)
	) name7043 (
		\s7_next_reg/P0001 ,
		_w6746_,
		_w6752_,
		_w8944_
	);
	LUT2 #(
		.INIT('h8)
	) name7044 (
		_w3481_,
		_w3484_,
		_w8945_
	);
	LUT4 #(
		.INIT('hd111)
	) name7045 (
		\s7_msel_pri_out_reg[0]/NET0131 ,
		\s7_next_reg/P0001 ,
		_w3481_,
		_w3484_,
		_w8946_
	);
	LUT4 #(
		.INIT('h1055)
	) name7046 (
		rst_i_pad,
		_w8943_,
		_w8944_,
		_w8946_,
		_w8947_
	);
	LUT4 #(
		.INIT('hf35f)
	) name7047 (
		\s11_msel_arb1_state_reg[1]/NET0131 ,
		\s11_msel_arb2_state_reg[1]/NET0131 ,
		\s11_msel_pri_out_reg[0]/NET0131 ,
		\s11_msel_pri_out_reg[1]/NET0131 ,
		_w8948_
	);
	LUT4 #(
		.INIT('h3ff5)
	) name7048 (
		\s11_msel_arb0_state_reg[1]/NET0131 ,
		\s11_msel_arb3_state_reg[1]/NET0131 ,
		\s11_msel_pri_out_reg[0]/NET0131 ,
		\s11_msel_pri_out_reg[1]/NET0131 ,
		_w8949_
	);
	LUT2 #(
		.INIT('h8)
	) name7049 (
		_w8948_,
		_w8949_,
		_w8950_
	);
	LUT4 #(
		.INIT('hf35f)
	) name7050 (
		\s11_msel_arb1_state_reg[2]/NET0131 ,
		\s11_msel_arb2_state_reg[2]/NET0131 ,
		\s11_msel_pri_out_reg[0]/NET0131 ,
		\s11_msel_pri_out_reg[1]/NET0131 ,
		_w8951_
	);
	LUT4 #(
		.INIT('h3ff5)
	) name7051 (
		\s11_msel_arb0_state_reg[2]/NET0131 ,
		\s11_msel_arb3_state_reg[2]/NET0131 ,
		\s11_msel_pri_out_reg[0]/NET0131 ,
		\s11_msel_pri_out_reg[1]/NET0131 ,
		_w8952_
	);
	LUT2 #(
		.INIT('h8)
	) name7052 (
		_w8951_,
		_w8952_,
		_w8953_
	);
	LUT4 #(
		.INIT('h0888)
	) name7053 (
		_w8948_,
		_w8949_,
		_w8951_,
		_w8952_,
		_w8954_
	);
	LUT4 #(
		.INIT('hf35f)
	) name7054 (
		\s11_msel_arb1_state_reg[0]/NET0131 ,
		\s11_msel_arb2_state_reg[0]/NET0131 ,
		\s11_msel_pri_out_reg[0]/NET0131 ,
		\s11_msel_pri_out_reg[1]/NET0131 ,
		_w8955_
	);
	LUT4 #(
		.INIT('h3ff5)
	) name7055 (
		\s11_msel_arb0_state_reg[0]/NET0131 ,
		\s11_msel_arb3_state_reg[0]/NET0131 ,
		\s11_msel_pri_out_reg[0]/NET0131 ,
		\s11_msel_pri_out_reg[1]/NET0131 ,
		_w8956_
	);
	LUT2 #(
		.INIT('h8)
	) name7056 (
		\m5_s11_cyc_o_reg/NET0131 ,
		\s11_m5_cyc_r_reg/P0001 ,
		_w8957_
	);
	LUT3 #(
		.INIT('h70)
	) name7057 (
		_w8955_,
		_w8956_,
		_w8957_,
		_w8958_
	);
	LUT2 #(
		.INIT('h8)
	) name7058 (
		\m4_s11_cyc_o_reg/NET0131 ,
		\s11_m4_cyc_r_reg/P0001 ,
		_w8959_
	);
	LUT3 #(
		.INIT('h80)
	) name7059 (
		_w8955_,
		_w8956_,
		_w8959_,
		_w8960_
	);
	LUT3 #(
		.INIT('h57)
	) name7060 (
		_w8954_,
		_w8958_,
		_w8960_,
		_w8961_
	);
	LUT4 #(
		.INIT('h8000)
	) name7061 (
		_w8948_,
		_w8949_,
		_w8951_,
		_w8952_,
		_w8962_
	);
	LUT2 #(
		.INIT('h8)
	) name7062 (
		\m1_s11_cyc_o_reg/NET0131 ,
		\s11_m1_cyc_r_reg/P0001 ,
		_w8963_
	);
	LUT3 #(
		.INIT('h70)
	) name7063 (
		_w8955_,
		_w8956_,
		_w8963_,
		_w8964_
	);
	LUT2 #(
		.INIT('h8)
	) name7064 (
		\m0_s11_cyc_o_reg/NET0131 ,
		\s11_m0_cyc_r_reg/P0001 ,
		_w8965_
	);
	LUT3 #(
		.INIT('h80)
	) name7065 (
		_w8955_,
		_w8956_,
		_w8965_,
		_w8966_
	);
	LUT3 #(
		.INIT('h57)
	) name7066 (
		_w8962_,
		_w8964_,
		_w8966_,
		_w8967_
	);
	LUT4 #(
		.INIT('h0777)
	) name7067 (
		_w8948_,
		_w8949_,
		_w8951_,
		_w8952_,
		_w8968_
	);
	LUT2 #(
		.INIT('h8)
	) name7068 (
		\m7_s11_cyc_o_reg/NET0131 ,
		\s11_m7_cyc_r_reg/P0001 ,
		_w8969_
	);
	LUT3 #(
		.INIT('h70)
	) name7069 (
		_w8955_,
		_w8956_,
		_w8969_,
		_w8970_
	);
	LUT2 #(
		.INIT('h8)
	) name7070 (
		\m6_s11_cyc_o_reg/NET0131 ,
		\s11_m6_cyc_r_reg/P0001 ,
		_w8971_
	);
	LUT3 #(
		.INIT('h80)
	) name7071 (
		_w8955_,
		_w8956_,
		_w8971_,
		_w8972_
	);
	LUT3 #(
		.INIT('h57)
	) name7072 (
		_w8968_,
		_w8970_,
		_w8972_,
		_w8973_
	);
	LUT4 #(
		.INIT('h7000)
	) name7073 (
		_w8948_,
		_w8949_,
		_w8951_,
		_w8952_,
		_w8974_
	);
	LUT2 #(
		.INIT('h8)
	) name7074 (
		\m3_s11_cyc_o_reg/NET0131 ,
		\s11_m3_cyc_r_reg/P0001 ,
		_w8975_
	);
	LUT3 #(
		.INIT('h70)
	) name7075 (
		_w8955_,
		_w8956_,
		_w8975_,
		_w8976_
	);
	LUT2 #(
		.INIT('h8)
	) name7076 (
		\m2_s11_cyc_o_reg/NET0131 ,
		\s11_m2_cyc_r_reg/P0001 ,
		_w8977_
	);
	LUT3 #(
		.INIT('h80)
	) name7077 (
		_w8955_,
		_w8956_,
		_w8977_,
		_w8978_
	);
	LUT3 #(
		.INIT('h57)
	) name7078 (
		_w8974_,
		_w8976_,
		_w8978_,
		_w8979_
	);
	LUT4 #(
		.INIT('h8000)
	) name7079 (
		_w8961_,
		_w8967_,
		_w8973_,
		_w8979_,
		_w8980_
	);
	LUT4 #(
		.INIT('h7fff)
	) name7080 (
		_w8961_,
		_w8967_,
		_w8973_,
		_w8979_,
		_w8981_
	);
	LUT4 #(
		.INIT('hf35f)
	) name7081 (
		\s0_msel_arb1_state_reg[1]/NET0131 ,
		\s0_msel_arb2_state_reg[1]/NET0131 ,
		\s0_msel_pri_out_reg[0]/NET0131 ,
		\s0_msel_pri_out_reg[1]/NET0131 ,
		_w8982_
	);
	LUT4 #(
		.INIT('h3ff5)
	) name7082 (
		\s0_msel_arb0_state_reg[1]/NET0131 ,
		\s0_msel_arb3_state_reg[1]/NET0131 ,
		\s0_msel_pri_out_reg[0]/NET0131 ,
		\s0_msel_pri_out_reg[1]/NET0131 ,
		_w8983_
	);
	LUT2 #(
		.INIT('h8)
	) name7083 (
		_w8982_,
		_w8983_,
		_w8984_
	);
	LUT4 #(
		.INIT('hf35f)
	) name7084 (
		\s0_msel_arb1_state_reg[2]/NET0131 ,
		\s0_msel_arb2_state_reg[2]/NET0131 ,
		\s0_msel_pri_out_reg[0]/NET0131 ,
		\s0_msel_pri_out_reg[1]/NET0131 ,
		_w8985_
	);
	LUT4 #(
		.INIT('h3ff5)
	) name7085 (
		\s0_msel_arb0_state_reg[2]/NET0131 ,
		\s0_msel_arb3_state_reg[2]/NET0131 ,
		\s0_msel_pri_out_reg[0]/NET0131 ,
		\s0_msel_pri_out_reg[1]/NET0131 ,
		_w8986_
	);
	LUT2 #(
		.INIT('h8)
	) name7086 (
		_w8985_,
		_w8986_,
		_w8987_
	);
	LUT4 #(
		.INIT('h0777)
	) name7087 (
		_w8982_,
		_w8983_,
		_w8985_,
		_w8986_,
		_w8988_
	);
	LUT4 #(
		.INIT('h3ff5)
	) name7088 (
		\s0_msel_arb0_state_reg[0]/NET0131 ,
		\s0_msel_arb3_state_reg[0]/NET0131 ,
		\s0_msel_pri_out_reg[0]/NET0131 ,
		\s0_msel_pri_out_reg[1]/NET0131 ,
		_w8989_
	);
	LUT4 #(
		.INIT('hf35f)
	) name7089 (
		\s0_msel_arb1_state_reg[0]/NET0131 ,
		\s0_msel_arb2_state_reg[0]/NET0131 ,
		\s0_msel_pri_out_reg[0]/NET0131 ,
		\s0_msel_pri_out_reg[1]/NET0131 ,
		_w8990_
	);
	LUT2 #(
		.INIT('h8)
	) name7090 (
		\m7_s0_cyc_o_reg/NET0131 ,
		\s0_m7_cyc_r_reg/P0001 ,
		_w8991_
	);
	LUT3 #(
		.INIT('h70)
	) name7091 (
		_w8989_,
		_w8990_,
		_w8991_,
		_w8992_
	);
	LUT2 #(
		.INIT('h8)
	) name7092 (
		\m6_s0_cyc_o_reg/NET0131 ,
		\s0_m6_cyc_r_reg/P0001 ,
		_w8993_
	);
	LUT3 #(
		.INIT('h80)
	) name7093 (
		_w8989_,
		_w8990_,
		_w8993_,
		_w8994_
	);
	LUT3 #(
		.INIT('h57)
	) name7094 (
		_w8988_,
		_w8992_,
		_w8994_,
		_w8995_
	);
	LUT4 #(
		.INIT('h0888)
	) name7095 (
		_w8982_,
		_w8983_,
		_w8985_,
		_w8986_,
		_w8996_
	);
	LUT2 #(
		.INIT('h8)
	) name7096 (
		\m5_s0_cyc_o_reg/NET0131 ,
		\s0_m5_cyc_r_reg/P0001 ,
		_w8997_
	);
	LUT3 #(
		.INIT('h70)
	) name7097 (
		_w8989_,
		_w8990_,
		_w8997_,
		_w8998_
	);
	LUT2 #(
		.INIT('h8)
	) name7098 (
		\m4_s0_cyc_o_reg/NET0131 ,
		\s0_m4_cyc_r_reg/P0001 ,
		_w8999_
	);
	LUT3 #(
		.INIT('h80)
	) name7099 (
		_w8989_,
		_w8990_,
		_w8999_,
		_w9000_
	);
	LUT3 #(
		.INIT('h57)
	) name7100 (
		_w8996_,
		_w8998_,
		_w9000_,
		_w9001_
	);
	LUT4 #(
		.INIT('h7000)
	) name7101 (
		_w8982_,
		_w8983_,
		_w8985_,
		_w8986_,
		_w9002_
	);
	LUT2 #(
		.INIT('h8)
	) name7102 (
		\m3_s0_cyc_o_reg/NET0131 ,
		\s0_m3_cyc_r_reg/P0001 ,
		_w9003_
	);
	LUT3 #(
		.INIT('h70)
	) name7103 (
		_w8989_,
		_w8990_,
		_w9003_,
		_w9004_
	);
	LUT2 #(
		.INIT('h8)
	) name7104 (
		\m2_s0_cyc_o_reg/NET0131 ,
		\s0_m2_cyc_r_reg/P0001 ,
		_w9005_
	);
	LUT3 #(
		.INIT('h80)
	) name7105 (
		_w8989_,
		_w8990_,
		_w9005_,
		_w9006_
	);
	LUT3 #(
		.INIT('h57)
	) name7106 (
		_w9002_,
		_w9004_,
		_w9006_,
		_w9007_
	);
	LUT4 #(
		.INIT('h8000)
	) name7107 (
		_w8982_,
		_w8983_,
		_w8985_,
		_w8986_,
		_w9008_
	);
	LUT2 #(
		.INIT('h8)
	) name7108 (
		\m1_s0_cyc_o_reg/NET0131 ,
		\s0_m1_cyc_r_reg/P0001 ,
		_w9009_
	);
	LUT3 #(
		.INIT('h70)
	) name7109 (
		_w8989_,
		_w8990_,
		_w9009_,
		_w9010_
	);
	LUT2 #(
		.INIT('h8)
	) name7110 (
		\m0_s0_cyc_o_reg/NET0131 ,
		\s0_m0_cyc_r_reg/P0001 ,
		_w9011_
	);
	LUT3 #(
		.INIT('h80)
	) name7111 (
		_w8989_,
		_w8990_,
		_w9011_,
		_w9012_
	);
	LUT3 #(
		.INIT('h57)
	) name7112 (
		_w9008_,
		_w9010_,
		_w9012_,
		_w9013_
	);
	LUT4 #(
		.INIT('h8000)
	) name7113 (
		_w8995_,
		_w9001_,
		_w9007_,
		_w9013_,
		_w9014_
	);
	LUT4 #(
		.INIT('h7fff)
	) name7114 (
		_w8995_,
		_w9001_,
		_w9007_,
		_w9013_,
		_w9015_
	);
	LUT3 #(
		.INIT('h80)
	) name7115 (
		\s8_next_reg/P0001 ,
		_w3114_,
		_w3125_,
		_w9016_
	);
	LUT4 #(
		.INIT('h0001)
	) name7116 (
		_w3890_,
		_w3891_,
		_w3893_,
		_w3894_,
		_w9017_
	);
	LUT2 #(
		.INIT('h8)
	) name7117 (
		_w3901_,
		_w9017_,
		_w9018_
	);
	LUT2 #(
		.INIT('h8)
	) name7118 (
		_w3502_,
		_w3513_,
		_w9019_
	);
	LUT4 #(
		.INIT('hd111)
	) name7119 (
		\s8_msel_pri_out_reg[0]/NET0131 ,
		\s8_next_reg/P0001 ,
		_w3502_,
		_w3513_,
		_w9020_
	);
	LUT4 #(
		.INIT('h0455)
	) name7120 (
		rst_i_pad,
		_w9016_,
		_w9018_,
		_w9020_,
		_w9021_
	);
	LUT4 #(
		.INIT('hf35f)
	) name7121 (
		\s12_msel_arb1_state_reg[1]/NET0131 ,
		\s12_msel_arb2_state_reg[1]/NET0131 ,
		\s12_msel_pri_out_reg[0]/NET0131 ,
		\s12_msel_pri_out_reg[1]/NET0131 ,
		_w9022_
	);
	LUT4 #(
		.INIT('h3ff5)
	) name7122 (
		\s12_msel_arb0_state_reg[1]/NET0131 ,
		\s12_msel_arb3_state_reg[1]/NET0131 ,
		\s12_msel_pri_out_reg[0]/NET0131 ,
		\s12_msel_pri_out_reg[1]/NET0131 ,
		_w9023_
	);
	LUT2 #(
		.INIT('h8)
	) name7123 (
		_w9022_,
		_w9023_,
		_w9024_
	);
	LUT4 #(
		.INIT('hf3f5)
	) name7124 (
		\s12_msel_arb0_state_reg[2]/NET0131 ,
		\s12_msel_arb2_state_reg[2]/NET0131 ,
		\s12_msel_pri_out_reg[0]/NET0131 ,
		\s12_msel_pri_out_reg[1]/NET0131 ,
		_w9025_
	);
	LUT4 #(
		.INIT('h3f5f)
	) name7125 (
		\s12_msel_arb1_state_reg[2]/NET0131 ,
		\s12_msel_arb3_state_reg[2]/NET0131 ,
		\s12_msel_pri_out_reg[0]/NET0131 ,
		\s12_msel_pri_out_reg[1]/NET0131 ,
		_w9026_
	);
	LUT2 #(
		.INIT('h8)
	) name7126 (
		_w9025_,
		_w9026_,
		_w9027_
	);
	LUT4 #(
		.INIT('h7000)
	) name7127 (
		_w9022_,
		_w9023_,
		_w9025_,
		_w9026_,
		_w9028_
	);
	LUT4 #(
		.INIT('hf35f)
	) name7128 (
		\s12_msel_arb1_state_reg[0]/NET0131 ,
		\s12_msel_arb2_state_reg[0]/NET0131 ,
		\s12_msel_pri_out_reg[0]/NET0131 ,
		\s12_msel_pri_out_reg[1]/NET0131 ,
		_w9029_
	);
	LUT4 #(
		.INIT('h3ff5)
	) name7129 (
		\s12_msel_arb0_state_reg[0]/NET0131 ,
		\s12_msel_arb3_state_reg[0]/NET0131 ,
		\s12_msel_pri_out_reg[0]/NET0131 ,
		\s12_msel_pri_out_reg[1]/NET0131 ,
		_w9030_
	);
	LUT2 #(
		.INIT('h8)
	) name7130 (
		\m3_s12_cyc_o_reg/NET0131 ,
		\s12_m3_cyc_r_reg/P0001 ,
		_w9031_
	);
	LUT3 #(
		.INIT('h70)
	) name7131 (
		_w9029_,
		_w9030_,
		_w9031_,
		_w9032_
	);
	LUT2 #(
		.INIT('h8)
	) name7132 (
		\m2_s12_cyc_o_reg/NET0131 ,
		\s12_m2_cyc_r_reg/P0001 ,
		_w9033_
	);
	LUT3 #(
		.INIT('h80)
	) name7133 (
		_w9029_,
		_w9030_,
		_w9033_,
		_w9034_
	);
	LUT3 #(
		.INIT('h57)
	) name7134 (
		_w9028_,
		_w9032_,
		_w9034_,
		_w9035_
	);
	LUT4 #(
		.INIT('h0777)
	) name7135 (
		_w9022_,
		_w9023_,
		_w9025_,
		_w9026_,
		_w9036_
	);
	LUT2 #(
		.INIT('h8)
	) name7136 (
		\m7_s12_cyc_o_reg/NET0131 ,
		\s12_m7_cyc_r_reg/P0001 ,
		_w9037_
	);
	LUT3 #(
		.INIT('h70)
	) name7137 (
		_w9029_,
		_w9030_,
		_w9037_,
		_w9038_
	);
	LUT2 #(
		.INIT('h8)
	) name7138 (
		\m6_s12_cyc_o_reg/NET0131 ,
		\s12_m6_cyc_r_reg/P0001 ,
		_w9039_
	);
	LUT3 #(
		.INIT('h80)
	) name7139 (
		_w9029_,
		_w9030_,
		_w9039_,
		_w9040_
	);
	LUT3 #(
		.INIT('h57)
	) name7140 (
		_w9036_,
		_w9038_,
		_w9040_,
		_w9041_
	);
	LUT4 #(
		.INIT('h0888)
	) name7141 (
		_w9022_,
		_w9023_,
		_w9025_,
		_w9026_,
		_w9042_
	);
	LUT2 #(
		.INIT('h8)
	) name7142 (
		\m5_s12_cyc_o_reg/NET0131 ,
		\s12_m5_cyc_r_reg/P0001 ,
		_w9043_
	);
	LUT3 #(
		.INIT('h70)
	) name7143 (
		_w9029_,
		_w9030_,
		_w9043_,
		_w9044_
	);
	LUT2 #(
		.INIT('h8)
	) name7144 (
		\m4_s12_cyc_o_reg/NET0131 ,
		\s12_m4_cyc_r_reg/P0001 ,
		_w9045_
	);
	LUT3 #(
		.INIT('h80)
	) name7145 (
		_w9029_,
		_w9030_,
		_w9045_,
		_w9046_
	);
	LUT3 #(
		.INIT('h57)
	) name7146 (
		_w9042_,
		_w9044_,
		_w9046_,
		_w9047_
	);
	LUT4 #(
		.INIT('h8000)
	) name7147 (
		_w9022_,
		_w9023_,
		_w9025_,
		_w9026_,
		_w9048_
	);
	LUT2 #(
		.INIT('h8)
	) name7148 (
		\m1_s12_cyc_o_reg/NET0131 ,
		\s12_m1_cyc_r_reg/P0001 ,
		_w9049_
	);
	LUT3 #(
		.INIT('h70)
	) name7149 (
		_w9029_,
		_w9030_,
		_w9049_,
		_w9050_
	);
	LUT2 #(
		.INIT('h8)
	) name7150 (
		\m0_s12_cyc_o_reg/NET0131 ,
		\s12_m0_cyc_r_reg/P0001 ,
		_w9051_
	);
	LUT3 #(
		.INIT('h80)
	) name7151 (
		_w9029_,
		_w9030_,
		_w9051_,
		_w9052_
	);
	LUT3 #(
		.INIT('h57)
	) name7152 (
		_w9048_,
		_w9050_,
		_w9052_,
		_w9053_
	);
	LUT4 #(
		.INIT('h8000)
	) name7153 (
		_w9035_,
		_w9041_,
		_w9047_,
		_w9053_,
		_w9054_
	);
	LUT4 #(
		.INIT('h7fff)
	) name7154 (
		_w9035_,
		_w9041_,
		_w9047_,
		_w9053_,
		_w9055_
	);
	LUT3 #(
		.INIT('h80)
	) name7155 (
		\s9_next_reg/P0001 ,
		_w6764_,
		_w6770_,
		_w9056_
	);
	LUT4 #(
		.INIT('h0001)
	) name7156 (
		_w3921_,
		_w3922_,
		_w3924_,
		_w3925_,
		_w9057_
	);
	LUT2 #(
		.INIT('h8)
	) name7157 (
		_w3932_,
		_w9057_,
		_w9058_
	);
	LUT2 #(
		.INIT('h8)
	) name7158 (
		_w6781_,
		_w6789_,
		_w9059_
	);
	LUT4 #(
		.INIT('hd111)
	) name7159 (
		\s9_msel_pri_out_reg[0]/NET0131 ,
		\s9_next_reg/P0001 ,
		_w6781_,
		_w6789_,
		_w9060_
	);
	LUT4 #(
		.INIT('h0455)
	) name7160 (
		rst_i_pad,
		_w9056_,
		_w9058_,
		_w9060_,
		_w9061_
	);
	LUT4 #(
		.INIT('hf35f)
	) name7161 (
		\s13_msel_arb1_state_reg[1]/NET0131 ,
		\s13_msel_arb2_state_reg[1]/NET0131 ,
		\s13_msel_pri_out_reg[0]/NET0131 ,
		\s13_msel_pri_out_reg[1]/NET0131 ,
		_w9062_
	);
	LUT4 #(
		.INIT('h3ff5)
	) name7162 (
		\s13_msel_arb0_state_reg[1]/NET0131 ,
		\s13_msel_arb3_state_reg[1]/NET0131 ,
		\s13_msel_pri_out_reg[0]/NET0131 ,
		\s13_msel_pri_out_reg[1]/NET0131 ,
		_w9063_
	);
	LUT2 #(
		.INIT('h8)
	) name7163 (
		_w9062_,
		_w9063_,
		_w9064_
	);
	LUT4 #(
		.INIT('h3ff5)
	) name7164 (
		\s13_msel_arb0_state_reg[2]/NET0131 ,
		\s13_msel_arb3_state_reg[2]/NET0131 ,
		\s13_msel_pri_out_reg[0]/NET0131 ,
		\s13_msel_pri_out_reg[1]/NET0131 ,
		_w9065_
	);
	LUT4 #(
		.INIT('hf35f)
	) name7165 (
		\s13_msel_arb1_state_reg[2]/NET0131 ,
		\s13_msel_arb2_state_reg[2]/NET0131 ,
		\s13_msel_pri_out_reg[0]/NET0131 ,
		\s13_msel_pri_out_reg[1]/NET0131 ,
		_w9066_
	);
	LUT2 #(
		.INIT('h8)
	) name7166 (
		_w9065_,
		_w9066_,
		_w9067_
	);
	LUT4 #(
		.INIT('h0777)
	) name7167 (
		_w9062_,
		_w9063_,
		_w9065_,
		_w9066_,
		_w9068_
	);
	LUT4 #(
		.INIT('hf35f)
	) name7168 (
		\s13_msel_arb1_state_reg[0]/NET0131 ,
		\s13_msel_arb2_state_reg[0]/NET0131 ,
		\s13_msel_pri_out_reg[0]/NET0131 ,
		\s13_msel_pri_out_reg[1]/NET0131 ,
		_w9069_
	);
	LUT4 #(
		.INIT('h3ff5)
	) name7169 (
		\s13_msel_arb0_state_reg[0]/NET0131 ,
		\s13_msel_arb3_state_reg[0]/NET0131 ,
		\s13_msel_pri_out_reg[0]/NET0131 ,
		\s13_msel_pri_out_reg[1]/NET0131 ,
		_w9070_
	);
	LUT2 #(
		.INIT('h8)
	) name7170 (
		\m7_s13_cyc_o_reg/NET0131 ,
		\s13_m7_cyc_r_reg/P0001 ,
		_w9071_
	);
	LUT3 #(
		.INIT('h70)
	) name7171 (
		_w9069_,
		_w9070_,
		_w9071_,
		_w9072_
	);
	LUT2 #(
		.INIT('h8)
	) name7172 (
		\m6_s13_cyc_o_reg/NET0131 ,
		\s13_m6_cyc_r_reg/P0001 ,
		_w9073_
	);
	LUT3 #(
		.INIT('h80)
	) name7173 (
		_w9069_,
		_w9070_,
		_w9073_,
		_w9074_
	);
	LUT3 #(
		.INIT('h57)
	) name7174 (
		_w9068_,
		_w9072_,
		_w9074_,
		_w9075_
	);
	LUT4 #(
		.INIT('h8000)
	) name7175 (
		_w9062_,
		_w9063_,
		_w9065_,
		_w9066_,
		_w9076_
	);
	LUT2 #(
		.INIT('h8)
	) name7176 (
		\m1_s13_cyc_o_reg/NET0131 ,
		\s13_m1_cyc_r_reg/P0001 ,
		_w9077_
	);
	LUT3 #(
		.INIT('h70)
	) name7177 (
		_w9069_,
		_w9070_,
		_w9077_,
		_w9078_
	);
	LUT2 #(
		.INIT('h8)
	) name7178 (
		\m0_s13_cyc_o_reg/NET0131 ,
		\s13_m0_cyc_r_reg/P0001 ,
		_w9079_
	);
	LUT3 #(
		.INIT('h80)
	) name7179 (
		_w9069_,
		_w9070_,
		_w9079_,
		_w9080_
	);
	LUT3 #(
		.INIT('h57)
	) name7180 (
		_w9076_,
		_w9078_,
		_w9080_,
		_w9081_
	);
	LUT4 #(
		.INIT('h7000)
	) name7181 (
		_w9062_,
		_w9063_,
		_w9065_,
		_w9066_,
		_w9082_
	);
	LUT2 #(
		.INIT('h8)
	) name7182 (
		\m3_s13_cyc_o_reg/NET0131 ,
		\s13_m3_cyc_r_reg/P0001 ,
		_w9083_
	);
	LUT3 #(
		.INIT('h70)
	) name7183 (
		_w9069_,
		_w9070_,
		_w9083_,
		_w9084_
	);
	LUT2 #(
		.INIT('h8)
	) name7184 (
		\m2_s13_cyc_o_reg/NET0131 ,
		\s13_m2_cyc_r_reg/P0001 ,
		_w9085_
	);
	LUT3 #(
		.INIT('h80)
	) name7185 (
		_w9069_,
		_w9070_,
		_w9085_,
		_w9086_
	);
	LUT3 #(
		.INIT('h57)
	) name7186 (
		_w9082_,
		_w9084_,
		_w9086_,
		_w9087_
	);
	LUT4 #(
		.INIT('h0888)
	) name7187 (
		_w9062_,
		_w9063_,
		_w9065_,
		_w9066_,
		_w9088_
	);
	LUT2 #(
		.INIT('h8)
	) name7188 (
		\m5_s13_cyc_o_reg/NET0131 ,
		\s13_m5_cyc_r_reg/P0001 ,
		_w9089_
	);
	LUT3 #(
		.INIT('h70)
	) name7189 (
		_w9069_,
		_w9070_,
		_w9089_,
		_w9090_
	);
	LUT2 #(
		.INIT('h8)
	) name7190 (
		\m4_s13_cyc_o_reg/NET0131 ,
		\s13_m4_cyc_r_reg/P0001 ,
		_w9091_
	);
	LUT3 #(
		.INIT('h80)
	) name7191 (
		_w9069_,
		_w9070_,
		_w9091_,
		_w9092_
	);
	LUT3 #(
		.INIT('h57)
	) name7192 (
		_w9088_,
		_w9090_,
		_w9092_,
		_w9093_
	);
	LUT4 #(
		.INIT('h8000)
	) name7193 (
		_w9075_,
		_w9081_,
		_w9087_,
		_w9093_,
		_w9094_
	);
	LUT4 #(
		.INIT('h7fff)
	) name7194 (
		_w9075_,
		_w9081_,
		_w9087_,
		_w9093_,
		_w9095_
	);
	LUT4 #(
		.INIT('hf35f)
	) name7195 (
		\s1_msel_arb1_state_reg[1]/NET0131 ,
		\s1_msel_arb2_state_reg[1]/NET0131 ,
		\s1_msel_pri_out_reg[0]/NET0131 ,
		\s1_msel_pri_out_reg[1]/NET0131 ,
		_w9096_
	);
	LUT4 #(
		.INIT('h3ff5)
	) name7196 (
		\s1_msel_arb0_state_reg[1]/NET0131 ,
		\s1_msel_arb3_state_reg[1]/NET0131 ,
		\s1_msel_pri_out_reg[0]/NET0131 ,
		\s1_msel_pri_out_reg[1]/NET0131 ,
		_w9097_
	);
	LUT2 #(
		.INIT('h8)
	) name7197 (
		_w9096_,
		_w9097_,
		_w9098_
	);
	LUT4 #(
		.INIT('h3ff5)
	) name7198 (
		\s1_msel_arb0_state_reg[2]/NET0131 ,
		\s1_msel_arb3_state_reg[2]/NET0131 ,
		\s1_msel_pri_out_reg[0]/NET0131 ,
		\s1_msel_pri_out_reg[1]/NET0131 ,
		_w9099_
	);
	LUT4 #(
		.INIT('hf35f)
	) name7199 (
		\s1_msel_arb1_state_reg[2]/NET0131 ,
		\s1_msel_arb2_state_reg[2]/NET0131 ,
		\s1_msel_pri_out_reg[0]/NET0131 ,
		\s1_msel_pri_out_reg[1]/NET0131 ,
		_w9100_
	);
	LUT2 #(
		.INIT('h8)
	) name7200 (
		_w9099_,
		_w9100_,
		_w9101_
	);
	LUT4 #(
		.INIT('h0777)
	) name7201 (
		_w9096_,
		_w9097_,
		_w9099_,
		_w9100_,
		_w9102_
	);
	LUT4 #(
		.INIT('hf35f)
	) name7202 (
		\s1_msel_arb1_state_reg[0]/NET0131 ,
		\s1_msel_arb2_state_reg[0]/NET0131 ,
		\s1_msel_pri_out_reg[0]/NET0131 ,
		\s1_msel_pri_out_reg[1]/NET0131 ,
		_w9103_
	);
	LUT4 #(
		.INIT('h3ff5)
	) name7203 (
		\s1_msel_arb0_state_reg[0]/NET0131 ,
		\s1_msel_arb3_state_reg[0]/NET0131 ,
		\s1_msel_pri_out_reg[0]/NET0131 ,
		\s1_msel_pri_out_reg[1]/NET0131 ,
		_w9104_
	);
	LUT2 #(
		.INIT('h8)
	) name7204 (
		\m7_s1_cyc_o_reg/NET0131 ,
		\s1_m7_cyc_r_reg/P0001 ,
		_w9105_
	);
	LUT3 #(
		.INIT('h70)
	) name7205 (
		_w9103_,
		_w9104_,
		_w9105_,
		_w9106_
	);
	LUT2 #(
		.INIT('h8)
	) name7206 (
		\m6_s1_cyc_o_reg/NET0131 ,
		\s1_m6_cyc_r_reg/P0001 ,
		_w9107_
	);
	LUT3 #(
		.INIT('h80)
	) name7207 (
		_w9103_,
		_w9104_,
		_w9107_,
		_w9108_
	);
	LUT3 #(
		.INIT('h57)
	) name7208 (
		_w9102_,
		_w9106_,
		_w9108_,
		_w9109_
	);
	LUT4 #(
		.INIT('h7000)
	) name7209 (
		_w9096_,
		_w9097_,
		_w9099_,
		_w9100_,
		_w9110_
	);
	LUT2 #(
		.INIT('h8)
	) name7210 (
		\m3_s1_cyc_o_reg/NET0131 ,
		\s1_m3_cyc_r_reg/P0001 ,
		_w9111_
	);
	LUT3 #(
		.INIT('h70)
	) name7211 (
		_w9103_,
		_w9104_,
		_w9111_,
		_w9112_
	);
	LUT2 #(
		.INIT('h8)
	) name7212 (
		\m2_s1_cyc_o_reg/NET0131 ,
		\s1_m2_cyc_r_reg/P0001 ,
		_w9113_
	);
	LUT3 #(
		.INIT('h80)
	) name7213 (
		_w9103_,
		_w9104_,
		_w9113_,
		_w9114_
	);
	LUT3 #(
		.INIT('h57)
	) name7214 (
		_w9110_,
		_w9112_,
		_w9114_,
		_w9115_
	);
	LUT4 #(
		.INIT('h0888)
	) name7215 (
		_w9096_,
		_w9097_,
		_w9099_,
		_w9100_,
		_w9116_
	);
	LUT2 #(
		.INIT('h8)
	) name7216 (
		\m5_s1_cyc_o_reg/NET0131 ,
		\s1_m5_cyc_r_reg/P0001 ,
		_w9117_
	);
	LUT3 #(
		.INIT('h70)
	) name7217 (
		_w9103_,
		_w9104_,
		_w9117_,
		_w9118_
	);
	LUT2 #(
		.INIT('h8)
	) name7218 (
		\m4_s1_cyc_o_reg/NET0131 ,
		\s1_m4_cyc_r_reg/P0001 ,
		_w9119_
	);
	LUT3 #(
		.INIT('h80)
	) name7219 (
		_w9103_,
		_w9104_,
		_w9119_,
		_w9120_
	);
	LUT3 #(
		.INIT('h57)
	) name7220 (
		_w9116_,
		_w9118_,
		_w9120_,
		_w9121_
	);
	LUT4 #(
		.INIT('h8000)
	) name7221 (
		_w9096_,
		_w9097_,
		_w9099_,
		_w9100_,
		_w9122_
	);
	LUT2 #(
		.INIT('h8)
	) name7222 (
		\m1_s1_cyc_o_reg/NET0131 ,
		\s1_m1_cyc_r_reg/P0001 ,
		_w9123_
	);
	LUT3 #(
		.INIT('h70)
	) name7223 (
		_w9103_,
		_w9104_,
		_w9123_,
		_w9124_
	);
	LUT2 #(
		.INIT('h8)
	) name7224 (
		\m0_s1_cyc_o_reg/NET0131 ,
		\s1_m0_cyc_r_reg/P0001 ,
		_w9125_
	);
	LUT3 #(
		.INIT('h80)
	) name7225 (
		_w9103_,
		_w9104_,
		_w9125_,
		_w9126_
	);
	LUT3 #(
		.INIT('h57)
	) name7226 (
		_w9122_,
		_w9124_,
		_w9126_,
		_w9127_
	);
	LUT4 #(
		.INIT('h8000)
	) name7227 (
		_w9109_,
		_w9115_,
		_w9121_,
		_w9127_,
		_w9128_
	);
	LUT4 #(
		.INIT('h7fff)
	) name7228 (
		_w9109_,
		_w9115_,
		_w9121_,
		_w9127_,
		_w9129_
	);
	LUT4 #(
		.INIT('hf35f)
	) name7229 (
		\s14_msel_arb1_state_reg[2]/NET0131 ,
		\s14_msel_arb2_state_reg[2]/NET0131 ,
		\s14_msel_pri_out_reg[0]/NET0131 ,
		\s14_msel_pri_out_reg[1]/NET0131 ,
		_w9130_
	);
	LUT4 #(
		.INIT('h3ff5)
	) name7230 (
		\s14_msel_arb0_state_reg[2]/NET0131 ,
		\s14_msel_arb3_state_reg[2]/NET0131 ,
		\s14_msel_pri_out_reg[0]/NET0131 ,
		\s14_msel_pri_out_reg[1]/NET0131 ,
		_w9131_
	);
	LUT2 #(
		.INIT('h8)
	) name7231 (
		_w9130_,
		_w9131_,
		_w9132_
	);
	LUT4 #(
		.INIT('hf35f)
	) name7232 (
		\s14_msel_arb1_state_reg[1]/NET0131 ,
		\s14_msel_arb2_state_reg[1]/NET0131 ,
		\s14_msel_pri_out_reg[0]/NET0131 ,
		\s14_msel_pri_out_reg[1]/NET0131 ,
		_w9133_
	);
	LUT4 #(
		.INIT('h3ff5)
	) name7233 (
		\s14_msel_arb0_state_reg[1]/NET0131 ,
		\s14_msel_arb3_state_reg[1]/NET0131 ,
		\s14_msel_pri_out_reg[0]/NET0131 ,
		\s14_msel_pri_out_reg[1]/NET0131 ,
		_w9134_
	);
	LUT2 #(
		.INIT('h8)
	) name7234 (
		_w9133_,
		_w9134_,
		_w9135_
	);
	LUT4 #(
		.INIT('h8000)
	) name7235 (
		_w9130_,
		_w9131_,
		_w9133_,
		_w9134_,
		_w9136_
	);
	LUT4 #(
		.INIT('hf35f)
	) name7236 (
		\s14_msel_arb1_state_reg[0]/NET0131 ,
		\s14_msel_arb2_state_reg[0]/NET0131 ,
		\s14_msel_pri_out_reg[0]/NET0131 ,
		\s14_msel_pri_out_reg[1]/NET0131 ,
		_w9137_
	);
	LUT4 #(
		.INIT('h3ff5)
	) name7237 (
		\s14_msel_arb0_state_reg[0]/NET0131 ,
		\s14_msel_arb3_state_reg[0]/NET0131 ,
		\s14_msel_pri_out_reg[0]/NET0131 ,
		\s14_msel_pri_out_reg[1]/NET0131 ,
		_w9138_
	);
	LUT2 #(
		.INIT('h8)
	) name7238 (
		\m1_s14_cyc_o_reg/NET0131 ,
		\s14_m1_cyc_r_reg/P0001 ,
		_w9139_
	);
	LUT3 #(
		.INIT('h70)
	) name7239 (
		_w9137_,
		_w9138_,
		_w9139_,
		_w9140_
	);
	LUT2 #(
		.INIT('h8)
	) name7240 (
		\m0_s14_cyc_o_reg/NET0131 ,
		\s14_m0_cyc_r_reg/P0001 ,
		_w9141_
	);
	LUT3 #(
		.INIT('h80)
	) name7241 (
		_w9137_,
		_w9138_,
		_w9141_,
		_w9142_
	);
	LUT3 #(
		.INIT('h57)
	) name7242 (
		_w9136_,
		_w9140_,
		_w9142_,
		_w9143_
	);
	LUT4 #(
		.INIT('h0888)
	) name7243 (
		_w9130_,
		_w9131_,
		_w9133_,
		_w9134_,
		_w9144_
	);
	LUT2 #(
		.INIT('h8)
	) name7244 (
		\m3_s14_cyc_o_reg/NET0131 ,
		\s14_m3_cyc_r_reg/P0001 ,
		_w9145_
	);
	LUT3 #(
		.INIT('h70)
	) name7245 (
		_w9137_,
		_w9138_,
		_w9145_,
		_w9146_
	);
	LUT2 #(
		.INIT('h8)
	) name7246 (
		\m2_s14_cyc_o_reg/NET0131 ,
		\s14_m2_cyc_r_reg/P0001 ,
		_w9147_
	);
	LUT3 #(
		.INIT('h80)
	) name7247 (
		_w9137_,
		_w9138_,
		_w9147_,
		_w9148_
	);
	LUT3 #(
		.INIT('h57)
	) name7248 (
		_w9144_,
		_w9146_,
		_w9148_,
		_w9149_
	);
	LUT4 #(
		.INIT('h0777)
	) name7249 (
		_w9130_,
		_w9131_,
		_w9133_,
		_w9134_,
		_w9150_
	);
	LUT2 #(
		.INIT('h8)
	) name7250 (
		\m7_s14_cyc_o_reg/NET0131 ,
		\s14_m7_cyc_r_reg/P0001 ,
		_w9151_
	);
	LUT3 #(
		.INIT('h70)
	) name7251 (
		_w9137_,
		_w9138_,
		_w9151_,
		_w9152_
	);
	LUT2 #(
		.INIT('h8)
	) name7252 (
		\m6_s14_cyc_o_reg/NET0131 ,
		\s14_m6_cyc_r_reg/P0001 ,
		_w9153_
	);
	LUT3 #(
		.INIT('h80)
	) name7253 (
		_w9137_,
		_w9138_,
		_w9153_,
		_w9154_
	);
	LUT3 #(
		.INIT('h57)
	) name7254 (
		_w9150_,
		_w9152_,
		_w9154_,
		_w9155_
	);
	LUT4 #(
		.INIT('h7000)
	) name7255 (
		_w9130_,
		_w9131_,
		_w9133_,
		_w9134_,
		_w9156_
	);
	LUT2 #(
		.INIT('h8)
	) name7256 (
		\m5_s14_cyc_o_reg/NET0131 ,
		\s14_m5_cyc_r_reg/P0001 ,
		_w9157_
	);
	LUT3 #(
		.INIT('h70)
	) name7257 (
		_w9137_,
		_w9138_,
		_w9157_,
		_w9158_
	);
	LUT2 #(
		.INIT('h8)
	) name7258 (
		\m4_s14_cyc_o_reg/NET0131 ,
		\s14_m4_cyc_r_reg/P0001 ,
		_w9159_
	);
	LUT3 #(
		.INIT('h80)
	) name7259 (
		_w9137_,
		_w9138_,
		_w9159_,
		_w9160_
	);
	LUT3 #(
		.INIT('h57)
	) name7260 (
		_w9156_,
		_w9158_,
		_w9160_,
		_w9161_
	);
	LUT4 #(
		.INIT('h8000)
	) name7261 (
		_w9143_,
		_w9149_,
		_w9155_,
		_w9161_,
		_w9162_
	);
	LUT4 #(
		.INIT('h7fff)
	) name7262 (
		_w9143_,
		_w9149_,
		_w9155_,
		_w9161_,
		_w9163_
	);
	LUT4 #(
		.INIT('hf35f)
	) name7263 (
		\s2_msel_arb1_state_reg[1]/NET0131 ,
		\s2_msel_arb2_state_reg[1]/NET0131 ,
		\s2_msel_pri_out_reg[0]/NET0131 ,
		\s2_msel_pri_out_reg[1]/NET0131 ,
		_w9164_
	);
	LUT4 #(
		.INIT('h3ff5)
	) name7264 (
		\s2_msel_arb0_state_reg[1]/NET0131 ,
		\s2_msel_arb3_state_reg[1]/NET0131 ,
		\s2_msel_pri_out_reg[0]/NET0131 ,
		\s2_msel_pri_out_reg[1]/NET0131 ,
		_w9165_
	);
	LUT2 #(
		.INIT('h8)
	) name7265 (
		_w9164_,
		_w9165_,
		_w9166_
	);
	LUT4 #(
		.INIT('hf35f)
	) name7266 (
		\s2_msel_arb1_state_reg[2]/NET0131 ,
		\s2_msel_arb2_state_reg[2]/NET0131 ,
		\s2_msel_pri_out_reg[0]/NET0131 ,
		\s2_msel_pri_out_reg[1]/NET0131 ,
		_w9167_
	);
	LUT4 #(
		.INIT('h3ff5)
	) name7267 (
		\s2_msel_arb0_state_reg[2]/NET0131 ,
		\s2_msel_arb3_state_reg[2]/NET0131 ,
		\s2_msel_pri_out_reg[0]/NET0131 ,
		\s2_msel_pri_out_reg[1]/NET0131 ,
		_w9168_
	);
	LUT2 #(
		.INIT('h8)
	) name7268 (
		_w9167_,
		_w9168_,
		_w9169_
	);
	LUT4 #(
		.INIT('h0888)
	) name7269 (
		_w9164_,
		_w9165_,
		_w9167_,
		_w9168_,
		_w9170_
	);
	LUT4 #(
		.INIT('hf35f)
	) name7270 (
		\s2_msel_arb1_state_reg[0]/NET0131 ,
		\s2_msel_arb2_state_reg[0]/NET0131 ,
		\s2_msel_pri_out_reg[0]/NET0131 ,
		\s2_msel_pri_out_reg[1]/NET0131 ,
		_w9171_
	);
	LUT4 #(
		.INIT('h3ff5)
	) name7271 (
		\s2_msel_arb0_state_reg[0]/NET0131 ,
		\s2_msel_arb3_state_reg[0]/NET0131 ,
		\s2_msel_pri_out_reg[0]/NET0131 ,
		\s2_msel_pri_out_reg[1]/NET0131 ,
		_w9172_
	);
	LUT2 #(
		.INIT('h8)
	) name7272 (
		\m5_s2_cyc_o_reg/NET0131 ,
		\s2_m5_cyc_r_reg/P0001 ,
		_w9173_
	);
	LUT3 #(
		.INIT('h70)
	) name7273 (
		_w9171_,
		_w9172_,
		_w9173_,
		_w9174_
	);
	LUT2 #(
		.INIT('h8)
	) name7274 (
		\m4_s2_cyc_o_reg/NET0131 ,
		\s2_m4_cyc_r_reg/P0001 ,
		_w9175_
	);
	LUT3 #(
		.INIT('h80)
	) name7275 (
		_w9171_,
		_w9172_,
		_w9175_,
		_w9176_
	);
	LUT3 #(
		.INIT('h57)
	) name7276 (
		_w9170_,
		_w9174_,
		_w9176_,
		_w9177_
	);
	LUT4 #(
		.INIT('h8000)
	) name7277 (
		_w9164_,
		_w9165_,
		_w9167_,
		_w9168_,
		_w9178_
	);
	LUT2 #(
		.INIT('h8)
	) name7278 (
		\m1_s2_cyc_o_reg/NET0131 ,
		\s2_m1_cyc_r_reg/P0001 ,
		_w9179_
	);
	LUT3 #(
		.INIT('h70)
	) name7279 (
		_w9171_,
		_w9172_,
		_w9179_,
		_w9180_
	);
	LUT2 #(
		.INIT('h8)
	) name7280 (
		\m0_s2_cyc_o_reg/NET0131 ,
		\s2_m0_cyc_r_reg/P0001 ,
		_w9181_
	);
	LUT3 #(
		.INIT('h80)
	) name7281 (
		_w9171_,
		_w9172_,
		_w9181_,
		_w9182_
	);
	LUT3 #(
		.INIT('h57)
	) name7282 (
		_w9178_,
		_w9180_,
		_w9182_,
		_w9183_
	);
	LUT4 #(
		.INIT('h0777)
	) name7283 (
		_w9164_,
		_w9165_,
		_w9167_,
		_w9168_,
		_w9184_
	);
	LUT2 #(
		.INIT('h8)
	) name7284 (
		\m7_s2_cyc_o_reg/NET0131 ,
		\s2_m7_cyc_r_reg/P0001 ,
		_w9185_
	);
	LUT3 #(
		.INIT('h70)
	) name7285 (
		_w9171_,
		_w9172_,
		_w9185_,
		_w9186_
	);
	LUT2 #(
		.INIT('h8)
	) name7286 (
		\m6_s2_cyc_o_reg/NET0131 ,
		\s2_m6_cyc_r_reg/P0001 ,
		_w9187_
	);
	LUT3 #(
		.INIT('h80)
	) name7287 (
		_w9171_,
		_w9172_,
		_w9187_,
		_w9188_
	);
	LUT3 #(
		.INIT('h57)
	) name7288 (
		_w9184_,
		_w9186_,
		_w9188_,
		_w9189_
	);
	LUT4 #(
		.INIT('h7000)
	) name7289 (
		_w9164_,
		_w9165_,
		_w9167_,
		_w9168_,
		_w9190_
	);
	LUT2 #(
		.INIT('h8)
	) name7290 (
		\m3_s2_cyc_o_reg/NET0131 ,
		\s2_m3_cyc_r_reg/P0001 ,
		_w9191_
	);
	LUT3 #(
		.INIT('h70)
	) name7291 (
		_w9171_,
		_w9172_,
		_w9191_,
		_w9192_
	);
	LUT2 #(
		.INIT('h8)
	) name7292 (
		\m2_s2_cyc_o_reg/NET0131 ,
		\s2_m2_cyc_r_reg/P0001 ,
		_w9193_
	);
	LUT3 #(
		.INIT('h80)
	) name7293 (
		_w9171_,
		_w9172_,
		_w9193_,
		_w9194_
	);
	LUT3 #(
		.INIT('h57)
	) name7294 (
		_w9190_,
		_w9192_,
		_w9194_,
		_w9195_
	);
	LUT4 #(
		.INIT('h8000)
	) name7295 (
		_w9177_,
		_w9183_,
		_w9189_,
		_w9195_,
		_w9196_
	);
	LUT4 #(
		.INIT('h7fff)
	) name7296 (
		_w9177_,
		_w9183_,
		_w9189_,
		_w9195_,
		_w9197_
	);
	LUT4 #(
		.INIT('hf35f)
	) name7297 (
		\s3_msel_arb1_state_reg[1]/NET0131 ,
		\s3_msel_arb2_state_reg[1]/NET0131 ,
		\s3_msel_pri_out_reg[0]/NET0131 ,
		\s3_msel_pri_out_reg[1]/NET0131 ,
		_w9198_
	);
	LUT4 #(
		.INIT('h3ff5)
	) name7298 (
		\s3_msel_arb0_state_reg[1]/NET0131 ,
		\s3_msel_arb3_state_reg[1]/NET0131 ,
		\s3_msel_pri_out_reg[0]/NET0131 ,
		\s3_msel_pri_out_reg[1]/NET0131 ,
		_w9199_
	);
	LUT2 #(
		.INIT('h8)
	) name7299 (
		_w9198_,
		_w9199_,
		_w9200_
	);
	LUT4 #(
		.INIT('hf35f)
	) name7300 (
		\s3_msel_arb1_state_reg[2]/NET0131 ,
		\s3_msel_arb2_state_reg[2]/NET0131 ,
		\s3_msel_pri_out_reg[0]/NET0131 ,
		\s3_msel_pri_out_reg[1]/NET0131 ,
		_w9201_
	);
	LUT4 #(
		.INIT('h3ff5)
	) name7301 (
		\s3_msel_arb0_state_reg[2]/NET0131 ,
		\s3_msel_arb3_state_reg[2]/NET0131 ,
		\s3_msel_pri_out_reg[0]/NET0131 ,
		\s3_msel_pri_out_reg[1]/NET0131 ,
		_w9202_
	);
	LUT2 #(
		.INIT('h8)
	) name7302 (
		_w9201_,
		_w9202_,
		_w9203_
	);
	LUT4 #(
		.INIT('h0888)
	) name7303 (
		_w9198_,
		_w9199_,
		_w9201_,
		_w9202_,
		_w9204_
	);
	LUT4 #(
		.INIT('hf35f)
	) name7304 (
		\s3_msel_arb1_state_reg[0]/NET0131 ,
		\s3_msel_arb2_state_reg[0]/NET0131 ,
		\s3_msel_pri_out_reg[0]/NET0131 ,
		\s3_msel_pri_out_reg[1]/NET0131 ,
		_w9205_
	);
	LUT4 #(
		.INIT('h3ff5)
	) name7305 (
		\s3_msel_arb0_state_reg[0]/NET0131 ,
		\s3_msel_arb3_state_reg[0]/NET0131 ,
		\s3_msel_pri_out_reg[0]/NET0131 ,
		\s3_msel_pri_out_reg[1]/NET0131 ,
		_w9206_
	);
	LUT2 #(
		.INIT('h8)
	) name7306 (
		\m5_s3_cyc_o_reg/NET0131 ,
		\s3_m5_cyc_r_reg/P0001 ,
		_w9207_
	);
	LUT3 #(
		.INIT('h70)
	) name7307 (
		_w9205_,
		_w9206_,
		_w9207_,
		_w9208_
	);
	LUT2 #(
		.INIT('h8)
	) name7308 (
		\m4_s3_cyc_o_reg/NET0131 ,
		\s3_m4_cyc_r_reg/P0001 ,
		_w9209_
	);
	LUT3 #(
		.INIT('h80)
	) name7309 (
		_w9205_,
		_w9206_,
		_w9209_,
		_w9210_
	);
	LUT3 #(
		.INIT('h57)
	) name7310 (
		_w9204_,
		_w9208_,
		_w9210_,
		_w9211_
	);
	LUT4 #(
		.INIT('h7000)
	) name7311 (
		_w9198_,
		_w9199_,
		_w9201_,
		_w9202_,
		_w9212_
	);
	LUT2 #(
		.INIT('h8)
	) name7312 (
		\m3_s3_cyc_o_reg/NET0131 ,
		\s3_m3_cyc_r_reg/P0001 ,
		_w9213_
	);
	LUT3 #(
		.INIT('h70)
	) name7313 (
		_w9205_,
		_w9206_,
		_w9213_,
		_w9214_
	);
	LUT2 #(
		.INIT('h8)
	) name7314 (
		\m2_s3_cyc_o_reg/NET0131 ,
		\s3_m2_cyc_r_reg/P0001 ,
		_w9215_
	);
	LUT3 #(
		.INIT('h80)
	) name7315 (
		_w9205_,
		_w9206_,
		_w9215_,
		_w9216_
	);
	LUT3 #(
		.INIT('h57)
	) name7316 (
		_w9212_,
		_w9214_,
		_w9216_,
		_w9217_
	);
	LUT4 #(
		.INIT('h0777)
	) name7317 (
		_w9198_,
		_w9199_,
		_w9201_,
		_w9202_,
		_w9218_
	);
	LUT2 #(
		.INIT('h8)
	) name7318 (
		\m7_s3_cyc_o_reg/NET0131 ,
		\s3_m7_cyc_r_reg/P0001 ,
		_w9219_
	);
	LUT3 #(
		.INIT('h70)
	) name7319 (
		_w9205_,
		_w9206_,
		_w9219_,
		_w9220_
	);
	LUT2 #(
		.INIT('h8)
	) name7320 (
		\m6_s3_cyc_o_reg/NET0131 ,
		\s3_m6_cyc_r_reg/P0001 ,
		_w9221_
	);
	LUT3 #(
		.INIT('h80)
	) name7321 (
		_w9205_,
		_w9206_,
		_w9221_,
		_w9222_
	);
	LUT3 #(
		.INIT('h57)
	) name7322 (
		_w9218_,
		_w9220_,
		_w9222_,
		_w9223_
	);
	LUT4 #(
		.INIT('h8000)
	) name7323 (
		_w9198_,
		_w9199_,
		_w9201_,
		_w9202_,
		_w9224_
	);
	LUT2 #(
		.INIT('h8)
	) name7324 (
		\m1_s3_cyc_o_reg/NET0131 ,
		\s3_m1_cyc_r_reg/P0001 ,
		_w9225_
	);
	LUT3 #(
		.INIT('h70)
	) name7325 (
		_w9205_,
		_w9206_,
		_w9225_,
		_w9226_
	);
	LUT2 #(
		.INIT('h8)
	) name7326 (
		\m0_s3_cyc_o_reg/NET0131 ,
		\s3_m0_cyc_r_reg/P0001 ,
		_w9227_
	);
	LUT3 #(
		.INIT('h80)
	) name7327 (
		_w9205_,
		_w9206_,
		_w9227_,
		_w9228_
	);
	LUT3 #(
		.INIT('h57)
	) name7328 (
		_w9224_,
		_w9226_,
		_w9228_,
		_w9229_
	);
	LUT4 #(
		.INIT('h8000)
	) name7329 (
		_w9211_,
		_w9217_,
		_w9223_,
		_w9229_,
		_w9230_
	);
	LUT4 #(
		.INIT('h7fff)
	) name7330 (
		_w9211_,
		_w9217_,
		_w9223_,
		_w9229_,
		_w9231_
	);
	LUT3 #(
		.INIT('h80)
	) name7331 (
		\s0_next_reg/P0001 ,
		_w3136_,
		_w3147_,
		_w9232_
	);
	LUT4 #(
		.INIT('h0001)
	) name7332 (
		_w3952_,
		_w3953_,
		_w3955_,
		_w3956_,
		_w9233_
	);
	LUT2 #(
		.INIT('h8)
	) name7333 (
		_w3963_,
		_w9233_,
		_w9234_
	);
	LUT2 #(
		.INIT('h8)
	) name7334 (
		_w3543_,
		_w3546_,
		_w9235_
	);
	LUT4 #(
		.INIT('hd111)
	) name7335 (
		\s0_msel_pri_out_reg[0]/NET0131 ,
		\s0_next_reg/P0001 ,
		_w3543_,
		_w3546_,
		_w9236_
	);
	LUT4 #(
		.INIT('h0455)
	) name7336 (
		rst_i_pad,
		_w9232_,
		_w9234_,
		_w9236_,
		_w9237_
	);
	LUT3 #(
		.INIT('h54)
	) name7337 (
		rst_i_pad,
		\s10_msel_pri_out_reg[1]/NET0131 ,
		\s10_next_reg/P0001 ,
		_w9238_
	);
	LUT3 #(
		.INIT('h70)
	) name7338 (
		_w8683_,
		_w8684_,
		_w9238_,
		_w9239_
	);
	LUT3 #(
		.INIT('h54)
	) name7339 (
		rst_i_pad,
		\s11_msel_pri_out_reg[1]/NET0131 ,
		\s11_next_reg/P0001 ,
		_w9240_
	);
	LUT3 #(
		.INIT('h70)
	) name7340 (
		_w8688_,
		_w8689_,
		_w9240_,
		_w9241_
	);
	LUT3 #(
		.INIT('h54)
	) name7341 (
		rst_i_pad,
		\s12_msel_pri_out_reg[1]/NET0131 ,
		\s12_next_reg/P0001 ,
		_w9242_
	);
	LUT3 #(
		.INIT('h70)
	) name7342 (
		_w8727_,
		_w8728_,
		_w9242_,
		_w9243_
	);
	LUT3 #(
		.INIT('h54)
	) name7343 (
		rst_i_pad,
		\s13_msel_pri_out_reg[1]/NET0131 ,
		\s13_next_reg/P0001 ,
		_w9244_
	);
	LUT3 #(
		.INIT('h70)
	) name7344 (
		_w8732_,
		_w8733_,
		_w9244_,
		_w9245_
	);
	LUT3 #(
		.INIT('h54)
	) name7345 (
		rst_i_pad,
		\s14_msel_pri_out_reg[1]/NET0131 ,
		\s14_next_reg/P0001 ,
		_w9246_
	);
	LUT3 #(
		.INIT('h70)
	) name7346 (
		_w8771_,
		_w8772_,
		_w9246_,
		_w9247_
	);
	LUT3 #(
		.INIT('h54)
	) name7347 (
		rst_i_pad,
		\s1_msel_pri_out_reg[1]/NET0131 ,
		\s1_next_reg/P0001 ,
		_w9248_
	);
	LUT3 #(
		.INIT('h70)
	) name7348 (
		_w8810_,
		_w8811_,
		_w9248_,
		_w9249_
	);
	LUT3 #(
		.INIT('h54)
	) name7349 (
		rst_i_pad,
		\s2_msel_pri_out_reg[1]/NET0131 ,
		\s2_next_reg/P0001 ,
		_w9250_
	);
	LUT3 #(
		.INIT('h70)
	) name7350 (
		_w8849_,
		_w8850_,
		_w9250_,
		_w9251_
	);
	LUT3 #(
		.INIT('h54)
	) name7351 (
		rst_i_pad,
		\s3_msel_pri_out_reg[1]/NET0131 ,
		\s3_next_reg/P0001 ,
		_w9252_
	);
	LUT3 #(
		.INIT('h70)
	) name7352 (
		_w8854_,
		_w8855_,
		_w9252_,
		_w9253_
	);
	LUT3 #(
		.INIT('h54)
	) name7353 (
		rst_i_pad,
		\s4_msel_pri_out_reg[1]/NET0131 ,
		\s4_next_reg/P0001 ,
		_w9254_
	);
	LUT3 #(
		.INIT('h70)
	) name7354 (
		_w8893_,
		_w8894_,
		_w9254_,
		_w9255_
	);
	LUT3 #(
		.INIT('h54)
	) name7355 (
		rst_i_pad,
		\s5_msel_pri_out_reg[1]/NET0131 ,
		\s5_next_reg/P0001 ,
		_w9256_
	);
	LUT3 #(
		.INIT('h70)
	) name7356 (
		_w8897_,
		_w8900_,
		_w9256_,
		_w9257_
	);
	LUT3 #(
		.INIT('h54)
	) name7357 (
		rst_i_pad,
		\s6_msel_pri_out_reg[1]/NET0131 ,
		\s6_next_reg/P0001 ,
		_w9258_
	);
	LUT3 #(
		.INIT('h70)
	) name7358 (
		_w8937_,
		_w8940_,
		_w9258_,
		_w9259_
	);
	LUT3 #(
		.INIT('h54)
	) name7359 (
		rst_i_pad,
		\s7_msel_pri_out_reg[1]/NET0131 ,
		\s7_next_reg/P0001 ,
		_w9260_
	);
	LUT3 #(
		.INIT('h70)
	) name7360 (
		_w8944_,
		_w8945_,
		_w9260_,
		_w9261_
	);
	LUT3 #(
		.INIT('h54)
	) name7361 (
		rst_i_pad,
		\s8_msel_pri_out_reg[1]/NET0131 ,
		\s8_next_reg/P0001 ,
		_w9262_
	);
	LUT3 #(
		.INIT('h70)
	) name7362 (
		_w9016_,
		_w9019_,
		_w9262_,
		_w9263_
	);
	LUT3 #(
		.INIT('h54)
	) name7363 (
		rst_i_pad,
		\s9_msel_pri_out_reg[1]/NET0131 ,
		\s9_next_reg/P0001 ,
		_w9264_
	);
	LUT3 #(
		.INIT('h70)
	) name7364 (
		_w9056_,
		_w9059_,
		_w9264_,
		_w9265_
	);
	LUT3 #(
		.INIT('h54)
	) name7365 (
		rst_i_pad,
		\s0_msel_pri_out_reg[1]/NET0131 ,
		\s0_next_reg/P0001 ,
		_w9266_
	);
	LUT3 #(
		.INIT('h70)
	) name7366 (
		_w9232_,
		_w9235_,
		_w9266_,
		_w9267_
	);
	LUT3 #(
		.INIT('h08)
	) name7367 (
		\m5_cyc_i_pad ,
		\m5_s1_cyc_o_reg/NET0131 ,
		\m5_stb_i_pad ,
		_w9268_
	);
	LUT4 #(
		.INIT('h0002)
	) name7368 (
		\m5_addr_i[28]_pad ,
		\m5_addr_i[29]_pad ,
		\m5_addr_i[30]_pad ,
		\m5_addr_i[31]_pad ,
		_w9269_
	);
	LUT2 #(
		.INIT('h8)
	) name7369 (
		\m5_cyc_i_pad ,
		\m5_stb_i_pad ,
		_w9270_
	);
	LUT3 #(
		.INIT('hea)
	) name7370 (
		_w9268_,
		_w9269_,
		_w9270_,
		_w9271_
	);
	LUT3 #(
		.INIT('h08)
	) name7371 (
		\m0_cyc_i_pad ,
		\m0_s0_cyc_o_reg/NET0131 ,
		\m0_stb_i_pad ,
		_w9272_
	);
	LUT4 #(
		.INIT('h0001)
	) name7372 (
		\m0_addr_i[28]_pad ,
		\m0_addr_i[29]_pad ,
		\m0_addr_i[30]_pad ,
		\m0_addr_i[31]_pad ,
		_w9273_
	);
	LUT2 #(
		.INIT('h8)
	) name7373 (
		\m0_cyc_i_pad ,
		\m0_stb_i_pad ,
		_w9274_
	);
	LUT3 #(
		.INIT('hea)
	) name7374 (
		_w9272_,
		_w9273_,
		_w9274_,
		_w9275_
	);
	LUT3 #(
		.INIT('h08)
	) name7375 (
		\m0_cyc_i_pad ,
		\m0_s1_cyc_o_reg/NET0131 ,
		\m0_stb_i_pad ,
		_w9276_
	);
	LUT4 #(
		.INIT('h0002)
	) name7376 (
		\m0_addr_i[28]_pad ,
		\m0_addr_i[29]_pad ,
		\m0_addr_i[30]_pad ,
		\m0_addr_i[31]_pad ,
		_w9277_
	);
	LUT3 #(
		.INIT('hec)
	) name7377 (
		_w9274_,
		_w9276_,
		_w9277_,
		_w9278_
	);
	LUT3 #(
		.INIT('h08)
	) name7378 (
		\m1_cyc_i_pad ,
		\m1_s0_cyc_o_reg/NET0131 ,
		\m1_stb_i_pad ,
		_w9279_
	);
	LUT4 #(
		.INIT('h0001)
	) name7379 (
		\m1_addr_i[28]_pad ,
		\m1_addr_i[29]_pad ,
		\m1_addr_i[30]_pad ,
		\m1_addr_i[31]_pad ,
		_w9280_
	);
	LUT2 #(
		.INIT('h8)
	) name7380 (
		\m1_cyc_i_pad ,
		\m1_stb_i_pad ,
		_w9281_
	);
	LUT3 #(
		.INIT('hea)
	) name7381 (
		_w9279_,
		_w9280_,
		_w9281_,
		_w9282_
	);
	LUT3 #(
		.INIT('h08)
	) name7382 (
		\m2_cyc_i_pad ,
		\m2_s0_cyc_o_reg/NET0131 ,
		\m2_stb_i_pad ,
		_w9283_
	);
	LUT4 #(
		.INIT('h0001)
	) name7383 (
		\m2_addr_i[28]_pad ,
		\m2_addr_i[29]_pad ,
		\m2_addr_i[30]_pad ,
		\m2_addr_i[31]_pad ,
		_w9284_
	);
	LUT2 #(
		.INIT('h8)
	) name7384 (
		\m2_cyc_i_pad ,
		\m2_stb_i_pad ,
		_w9285_
	);
	LUT3 #(
		.INIT('hea)
	) name7385 (
		_w9283_,
		_w9284_,
		_w9285_,
		_w9286_
	);
	LUT3 #(
		.INIT('h08)
	) name7386 (
		\m2_cyc_i_pad ,
		\m2_s1_cyc_o_reg/NET0131 ,
		\m2_stb_i_pad ,
		_w9287_
	);
	LUT4 #(
		.INIT('h0002)
	) name7387 (
		\m2_addr_i[28]_pad ,
		\m2_addr_i[29]_pad ,
		\m2_addr_i[30]_pad ,
		\m2_addr_i[31]_pad ,
		_w9288_
	);
	LUT3 #(
		.INIT('hec)
	) name7388 (
		_w9285_,
		_w9287_,
		_w9288_,
		_w9289_
	);
	LUT3 #(
		.INIT('h08)
	) name7389 (
		\m3_cyc_i_pad ,
		\m3_s0_cyc_o_reg/NET0131 ,
		\m3_stb_i_pad ,
		_w9290_
	);
	LUT4 #(
		.INIT('h0001)
	) name7390 (
		\m3_addr_i[28]_pad ,
		\m3_addr_i[29]_pad ,
		\m3_addr_i[30]_pad ,
		\m3_addr_i[31]_pad ,
		_w9291_
	);
	LUT2 #(
		.INIT('h8)
	) name7391 (
		\m3_cyc_i_pad ,
		\m3_stb_i_pad ,
		_w9292_
	);
	LUT3 #(
		.INIT('hea)
	) name7392 (
		_w9290_,
		_w9291_,
		_w9292_,
		_w9293_
	);
	LUT3 #(
		.INIT('h08)
	) name7393 (
		\m3_cyc_i_pad ,
		\m3_s1_cyc_o_reg/NET0131 ,
		\m3_stb_i_pad ,
		_w9294_
	);
	LUT4 #(
		.INIT('h0002)
	) name7394 (
		\m3_addr_i[28]_pad ,
		\m3_addr_i[29]_pad ,
		\m3_addr_i[30]_pad ,
		\m3_addr_i[31]_pad ,
		_w9295_
	);
	LUT3 #(
		.INIT('hec)
	) name7395 (
		_w9292_,
		_w9294_,
		_w9295_,
		_w9296_
	);
	LUT3 #(
		.INIT('h08)
	) name7396 (
		\m4_cyc_i_pad ,
		\m4_s0_cyc_o_reg/NET0131 ,
		\m4_stb_i_pad ,
		_w9297_
	);
	LUT4 #(
		.INIT('h0001)
	) name7397 (
		\m4_addr_i[28]_pad ,
		\m4_addr_i[29]_pad ,
		\m4_addr_i[30]_pad ,
		\m4_addr_i[31]_pad ,
		_w9298_
	);
	LUT2 #(
		.INIT('h8)
	) name7398 (
		\m4_cyc_i_pad ,
		\m4_stb_i_pad ,
		_w9299_
	);
	LUT3 #(
		.INIT('hea)
	) name7399 (
		_w9297_,
		_w9298_,
		_w9299_,
		_w9300_
	);
	LUT3 #(
		.INIT('h08)
	) name7400 (
		\m4_cyc_i_pad ,
		\m4_s1_cyc_o_reg/NET0131 ,
		\m4_stb_i_pad ,
		_w9301_
	);
	LUT4 #(
		.INIT('h0002)
	) name7401 (
		\m4_addr_i[28]_pad ,
		\m4_addr_i[29]_pad ,
		\m4_addr_i[30]_pad ,
		\m4_addr_i[31]_pad ,
		_w9302_
	);
	LUT3 #(
		.INIT('hec)
	) name7402 (
		_w9299_,
		_w9301_,
		_w9302_,
		_w9303_
	);
	LUT3 #(
		.INIT('h08)
	) name7403 (
		\m5_cyc_i_pad ,
		\m5_s0_cyc_o_reg/NET0131 ,
		\m5_stb_i_pad ,
		_w9304_
	);
	LUT4 #(
		.INIT('h0001)
	) name7404 (
		\m5_addr_i[28]_pad ,
		\m5_addr_i[29]_pad ,
		\m5_addr_i[30]_pad ,
		\m5_addr_i[31]_pad ,
		_w9305_
	);
	LUT3 #(
		.INIT('hec)
	) name7405 (
		_w9270_,
		_w9304_,
		_w9305_,
		_w9306_
	);
	LUT3 #(
		.INIT('h08)
	) name7406 (
		\m6_cyc_i_pad ,
		\m6_s0_cyc_o_reg/NET0131 ,
		\m6_stb_i_pad ,
		_w9307_
	);
	LUT4 #(
		.INIT('h0001)
	) name7407 (
		\m6_addr_i[28]_pad ,
		\m6_addr_i[29]_pad ,
		\m6_addr_i[30]_pad ,
		\m6_addr_i[31]_pad ,
		_w9308_
	);
	LUT2 #(
		.INIT('h8)
	) name7408 (
		\m6_cyc_i_pad ,
		\m6_stb_i_pad ,
		_w9309_
	);
	LUT3 #(
		.INIT('hea)
	) name7409 (
		_w9307_,
		_w9308_,
		_w9309_,
		_w9310_
	);
	LUT3 #(
		.INIT('h08)
	) name7410 (
		\m6_cyc_i_pad ,
		\m6_s1_cyc_o_reg/NET0131 ,
		\m6_stb_i_pad ,
		_w9311_
	);
	LUT4 #(
		.INIT('h0002)
	) name7411 (
		\m6_addr_i[28]_pad ,
		\m6_addr_i[29]_pad ,
		\m6_addr_i[30]_pad ,
		\m6_addr_i[31]_pad ,
		_w9312_
	);
	LUT3 #(
		.INIT('hec)
	) name7412 (
		_w9309_,
		_w9311_,
		_w9312_,
		_w9313_
	);
	LUT3 #(
		.INIT('h08)
	) name7413 (
		\m7_cyc_i_pad ,
		\m7_s0_cyc_o_reg/NET0131 ,
		\m7_stb_i_pad ,
		_w9314_
	);
	LUT4 #(
		.INIT('h0001)
	) name7414 (
		\m7_addr_i[28]_pad ,
		\m7_addr_i[29]_pad ,
		\m7_addr_i[30]_pad ,
		\m7_addr_i[31]_pad ,
		_w9315_
	);
	LUT2 #(
		.INIT('h8)
	) name7415 (
		\m7_cyc_i_pad ,
		\m7_stb_i_pad ,
		_w9316_
	);
	LUT3 #(
		.INIT('hea)
	) name7416 (
		_w9314_,
		_w9315_,
		_w9316_,
		_w9317_
	);
	LUT3 #(
		.INIT('h08)
	) name7417 (
		\m7_cyc_i_pad ,
		\m7_s1_cyc_o_reg/NET0131 ,
		\m7_stb_i_pad ,
		_w9318_
	);
	LUT4 #(
		.INIT('h0002)
	) name7418 (
		\m7_addr_i[28]_pad ,
		\m7_addr_i[29]_pad ,
		\m7_addr_i[30]_pad ,
		\m7_addr_i[31]_pad ,
		_w9319_
	);
	LUT3 #(
		.INIT('hec)
	) name7419 (
		_w9316_,
		_w9318_,
		_w9319_,
		_w9320_
	);
	LUT3 #(
		.INIT('h08)
	) name7420 (
		\m1_cyc_i_pad ,
		\m1_s1_cyc_o_reg/NET0131 ,
		\m1_stb_i_pad ,
		_w9321_
	);
	LUT4 #(
		.INIT('h0002)
	) name7421 (
		\m1_addr_i[28]_pad ,
		\m1_addr_i[29]_pad ,
		\m1_addr_i[30]_pad ,
		\m1_addr_i[31]_pad ,
		_w9322_
	);
	LUT3 #(
		.INIT('hec)
	) name7422 (
		_w9281_,
		_w9321_,
		_w9322_,
		_w9323_
	);
	LUT3 #(
		.INIT('h08)
	) name7423 (
		\m5_cyc_i_pad ,
		\m5_s15_cyc_o_reg/NET0131 ,
		\m5_stb_i_pad ,
		_w9324_
	);
	LUT3 #(
		.INIT('hf8)
	) name7424 (
		_w2064_,
		_w9270_,
		_w9324_,
		_w9325_
	);
	LUT3 #(
		.INIT('h08)
	) name7425 (
		\m7_cyc_i_pad ,
		\m7_s9_cyc_o_reg/NET0131 ,
		\m7_stb_i_pad ,
		_w9326_
	);
	LUT4 #(
		.INIT('h0200)
	) name7426 (
		\m7_addr_i[28]_pad ,
		\m7_addr_i[29]_pad ,
		\m7_addr_i[30]_pad ,
		\m7_addr_i[31]_pad ,
		_w9327_
	);
	LUT3 #(
		.INIT('hec)
	) name7427 (
		_w9316_,
		_w9326_,
		_w9327_,
		_w9328_
	);
	LUT3 #(
		.INIT('h08)
	) name7428 (
		\m7_cyc_i_pad ,
		\m7_s7_cyc_o_reg/NET0131 ,
		\m7_stb_i_pad ,
		_w9329_
	);
	LUT4 #(
		.INIT('h0080)
	) name7429 (
		\m7_addr_i[28]_pad ,
		\m7_addr_i[29]_pad ,
		\m7_addr_i[30]_pad ,
		\m7_addr_i[31]_pad ,
		_w9330_
	);
	LUT3 #(
		.INIT('hec)
	) name7430 (
		_w9316_,
		_w9329_,
		_w9330_,
		_w9331_
	);
	LUT3 #(
		.INIT('h08)
	) name7431 (
		\m7_cyc_i_pad ,
		\m7_s5_cyc_o_reg/NET0131 ,
		\m7_stb_i_pad ,
		_w9332_
	);
	LUT4 #(
		.INIT('h0020)
	) name7432 (
		\m7_addr_i[28]_pad ,
		\m7_addr_i[29]_pad ,
		\m7_addr_i[30]_pad ,
		\m7_addr_i[31]_pad ,
		_w9333_
	);
	LUT3 #(
		.INIT('hec)
	) name7433 (
		_w9316_,
		_w9332_,
		_w9333_,
		_w9334_
	);
	LUT3 #(
		.INIT('h08)
	) name7434 (
		\m6_cyc_i_pad ,
		\m6_s6_cyc_o_reg/NET0131 ,
		\m6_stb_i_pad ,
		_w9335_
	);
	LUT4 #(
		.INIT('h0040)
	) name7435 (
		\m6_addr_i[28]_pad ,
		\m6_addr_i[29]_pad ,
		\m6_addr_i[30]_pad ,
		\m6_addr_i[31]_pad ,
		_w9336_
	);
	LUT3 #(
		.INIT('hec)
	) name7436 (
		_w9309_,
		_w9335_,
		_w9336_,
		_w9337_
	);
	LUT3 #(
		.INIT('h08)
	) name7437 (
		\m7_cyc_i_pad ,
		\m7_s12_cyc_o_reg/NET0131 ,
		\m7_stb_i_pad ,
		_w9338_
	);
	LUT4 #(
		.INIT('h1000)
	) name7438 (
		\m7_addr_i[28]_pad ,
		\m7_addr_i[29]_pad ,
		\m7_addr_i[30]_pad ,
		\m7_addr_i[31]_pad ,
		_w9339_
	);
	LUT3 #(
		.INIT('hec)
	) name7439 (
		_w9316_,
		_w9338_,
		_w9339_,
		_w9340_
	);
	LUT3 #(
		.INIT('h08)
	) name7440 (
		\m6_cyc_i_pad ,
		\m6_s8_cyc_o_reg/NET0131 ,
		\m6_stb_i_pad ,
		_w9341_
	);
	LUT4 #(
		.INIT('h0100)
	) name7441 (
		\m6_addr_i[28]_pad ,
		\m6_addr_i[29]_pad ,
		\m6_addr_i[30]_pad ,
		\m6_addr_i[31]_pad ,
		_w9342_
	);
	LUT3 #(
		.INIT('hec)
	) name7442 (
		_w9309_,
		_w9341_,
		_w9342_,
		_w9343_
	);
	LUT3 #(
		.INIT('h08)
	) name7443 (
		\m5_cyc_i_pad ,
		\m5_s7_cyc_o_reg/NET0131 ,
		\m5_stb_i_pad ,
		_w9344_
	);
	LUT4 #(
		.INIT('h0080)
	) name7444 (
		\m5_addr_i[28]_pad ,
		\m5_addr_i[29]_pad ,
		\m5_addr_i[30]_pad ,
		\m5_addr_i[31]_pad ,
		_w9345_
	);
	LUT3 #(
		.INIT('hec)
	) name7445 (
		_w9270_,
		_w9344_,
		_w9345_,
		_w9346_
	);
	LUT3 #(
		.INIT('h08)
	) name7446 (
		\m5_cyc_i_pad ,
		\m5_s14_cyc_o_reg/NET0131 ,
		\m5_stb_i_pad ,
		_w9347_
	);
	LUT4 #(
		.INIT('h4000)
	) name7447 (
		\m5_addr_i[28]_pad ,
		\m5_addr_i[29]_pad ,
		\m5_addr_i[30]_pad ,
		\m5_addr_i[31]_pad ,
		_w9348_
	);
	LUT3 #(
		.INIT('hec)
	) name7448 (
		_w9270_,
		_w9347_,
		_w9348_,
		_w9349_
	);
	LUT3 #(
		.INIT('h08)
	) name7449 (
		\m5_cyc_i_pad ,
		\m5_s3_cyc_o_reg/NET0131 ,
		\m5_stb_i_pad ,
		_w9350_
	);
	LUT4 #(
		.INIT('h0008)
	) name7450 (
		\m5_addr_i[28]_pad ,
		\m5_addr_i[29]_pad ,
		\m5_addr_i[30]_pad ,
		\m5_addr_i[31]_pad ,
		_w9351_
	);
	LUT3 #(
		.INIT('hec)
	) name7451 (
		_w9270_,
		_w9350_,
		_w9351_,
		_w9352_
	);
	LUT3 #(
		.INIT('h08)
	) name7452 (
		\m5_cyc_i_pad ,
		\m5_s12_cyc_o_reg/NET0131 ,
		\m5_stb_i_pad ,
		_w9353_
	);
	LUT4 #(
		.INIT('h1000)
	) name7453 (
		\m5_addr_i[28]_pad ,
		\m5_addr_i[29]_pad ,
		\m5_addr_i[30]_pad ,
		\m5_addr_i[31]_pad ,
		_w9354_
	);
	LUT3 #(
		.INIT('hec)
	) name7454 (
		_w9270_,
		_w9353_,
		_w9354_,
		_w9355_
	);
	LUT3 #(
		.INIT('h08)
	) name7455 (
		\m4_cyc_i_pad ,
		\m4_s9_cyc_o_reg/NET0131 ,
		\m4_stb_i_pad ,
		_w9356_
	);
	LUT4 #(
		.INIT('h0200)
	) name7456 (
		\m4_addr_i[28]_pad ,
		\m4_addr_i[29]_pad ,
		\m4_addr_i[30]_pad ,
		\m4_addr_i[31]_pad ,
		_w9357_
	);
	LUT3 #(
		.INIT('hec)
	) name7457 (
		_w9299_,
		_w9356_,
		_w9357_,
		_w9358_
	);
	LUT3 #(
		.INIT('h08)
	) name7458 (
		\m4_cyc_i_pad ,
		\m4_s8_cyc_o_reg/NET0131 ,
		\m4_stb_i_pad ,
		_w9359_
	);
	LUT4 #(
		.INIT('h0100)
	) name7459 (
		\m4_addr_i[28]_pad ,
		\m4_addr_i[29]_pad ,
		\m4_addr_i[30]_pad ,
		\m4_addr_i[31]_pad ,
		_w9360_
	);
	LUT3 #(
		.INIT('hec)
	) name7460 (
		_w9299_,
		_w9359_,
		_w9360_,
		_w9361_
	);
	LUT3 #(
		.INIT('h08)
	) name7461 (
		\m4_cyc_i_pad ,
		\m4_s6_cyc_o_reg/NET0131 ,
		\m4_stb_i_pad ,
		_w9362_
	);
	LUT4 #(
		.INIT('h0040)
	) name7462 (
		\m4_addr_i[28]_pad ,
		\m4_addr_i[29]_pad ,
		\m4_addr_i[30]_pad ,
		\m4_addr_i[31]_pad ,
		_w9363_
	);
	LUT3 #(
		.INIT('hec)
	) name7463 (
		_w9299_,
		_w9362_,
		_w9363_,
		_w9364_
	);
	LUT3 #(
		.INIT('h08)
	) name7464 (
		\m4_cyc_i_pad ,
		\m4_s4_cyc_o_reg/NET0131 ,
		\m4_stb_i_pad ,
		_w9365_
	);
	LUT4 #(
		.INIT('h0010)
	) name7465 (
		\m4_addr_i[28]_pad ,
		\m4_addr_i[29]_pad ,
		\m4_addr_i[30]_pad ,
		\m4_addr_i[31]_pad ,
		_w9366_
	);
	LUT3 #(
		.INIT('hec)
	) name7466 (
		_w9299_,
		_w9365_,
		_w9366_,
		_w9367_
	);
	LUT3 #(
		.INIT('h08)
	) name7467 (
		\m4_cyc_i_pad ,
		\m4_s13_cyc_o_reg/NET0131 ,
		\m4_stb_i_pad ,
		_w9368_
	);
	LUT4 #(
		.INIT('h2000)
	) name7468 (
		\m4_addr_i[28]_pad ,
		\m4_addr_i[29]_pad ,
		\m4_addr_i[30]_pad ,
		\m4_addr_i[31]_pad ,
		_w9369_
	);
	LUT3 #(
		.INIT('hec)
	) name7469 (
		_w9299_,
		_w9368_,
		_w9369_,
		_w9370_
	);
	LUT3 #(
		.INIT('h08)
	) name7470 (
		\m4_cyc_i_pad ,
		\m4_s11_cyc_o_reg/NET0131 ,
		\m4_stb_i_pad ,
		_w9371_
	);
	LUT4 #(
		.INIT('h0800)
	) name7471 (
		\m4_addr_i[28]_pad ,
		\m4_addr_i[29]_pad ,
		\m4_addr_i[30]_pad ,
		\m4_addr_i[31]_pad ,
		_w9372_
	);
	LUT3 #(
		.INIT('hec)
	) name7472 (
		_w9299_,
		_w9371_,
		_w9372_,
		_w9373_
	);
	LUT3 #(
		.INIT('h08)
	) name7473 (
		\m3_cyc_i_pad ,
		\m3_s7_cyc_o_reg/NET0131 ,
		\m3_stb_i_pad ,
		_w9374_
	);
	LUT4 #(
		.INIT('h0080)
	) name7474 (
		\m3_addr_i[28]_pad ,
		\m3_addr_i[29]_pad ,
		\m3_addr_i[30]_pad ,
		\m3_addr_i[31]_pad ,
		_w9375_
	);
	LUT3 #(
		.INIT('hec)
	) name7475 (
		_w9292_,
		_w9374_,
		_w9375_,
		_w9376_
	);
	LUT3 #(
		.INIT('h08)
	) name7476 (
		\m3_cyc_i_pad ,
		\m3_s6_cyc_o_reg/NET0131 ,
		\m3_stb_i_pad ,
		_w9377_
	);
	LUT4 #(
		.INIT('h0040)
	) name7477 (
		\m3_addr_i[28]_pad ,
		\m3_addr_i[29]_pad ,
		\m3_addr_i[30]_pad ,
		\m3_addr_i[31]_pad ,
		_w9378_
	);
	LUT3 #(
		.INIT('hec)
	) name7478 (
		_w9292_,
		_w9377_,
		_w9378_,
		_w9379_
	);
	LUT3 #(
		.INIT('h08)
	) name7479 (
		\m0_cyc_i_pad ,
		\m0_s10_cyc_o_reg/NET0131 ,
		\m0_stb_i_pad ,
		_w9380_
	);
	LUT4 #(
		.INIT('h0400)
	) name7480 (
		\m0_addr_i[28]_pad ,
		\m0_addr_i[29]_pad ,
		\m0_addr_i[30]_pad ,
		\m0_addr_i[31]_pad ,
		_w9381_
	);
	LUT3 #(
		.INIT('hec)
	) name7481 (
		_w9274_,
		_w9380_,
		_w9381_,
		_w9382_
	);
	LUT3 #(
		.INIT('h08)
	) name7482 (
		\m0_cyc_i_pad ,
		\m0_s11_cyc_o_reg/NET0131 ,
		\m0_stb_i_pad ,
		_w9383_
	);
	LUT4 #(
		.INIT('h0800)
	) name7483 (
		\m0_addr_i[28]_pad ,
		\m0_addr_i[29]_pad ,
		\m0_addr_i[30]_pad ,
		\m0_addr_i[31]_pad ,
		_w9384_
	);
	LUT3 #(
		.INIT('hec)
	) name7484 (
		_w9274_,
		_w9383_,
		_w9384_,
		_w9385_
	);
	LUT3 #(
		.INIT('h08)
	) name7485 (
		\m3_cyc_i_pad ,
		\m3_s5_cyc_o_reg/NET0131 ,
		\m3_stb_i_pad ,
		_w9386_
	);
	LUT4 #(
		.INIT('h0020)
	) name7486 (
		\m3_addr_i[28]_pad ,
		\m3_addr_i[29]_pad ,
		\m3_addr_i[30]_pad ,
		\m3_addr_i[31]_pad ,
		_w9387_
	);
	LUT3 #(
		.INIT('hec)
	) name7487 (
		_w9292_,
		_w9386_,
		_w9387_,
		_w9388_
	);
	LUT3 #(
		.INIT('h08)
	) name7488 (
		\m0_cyc_i_pad ,
		\m0_s14_cyc_o_reg/NET0131 ,
		\m0_stb_i_pad ,
		_w9389_
	);
	LUT4 #(
		.INIT('h4000)
	) name7489 (
		\m0_addr_i[28]_pad ,
		\m0_addr_i[29]_pad ,
		\m0_addr_i[30]_pad ,
		\m0_addr_i[31]_pad ,
		_w9390_
	);
	LUT3 #(
		.INIT('hec)
	) name7490 (
		_w9274_,
		_w9389_,
		_w9390_,
		_w9391_
	);
	LUT3 #(
		.INIT('h08)
	) name7491 (
		\m0_cyc_i_pad ,
		\m0_s15_cyc_o_reg/NET0131 ,
		\m0_stb_i_pad ,
		_w9392_
	);
	LUT3 #(
		.INIT('hf8)
	) name7492 (
		_w2049_,
		_w9274_,
		_w9392_,
		_w9393_
	);
	LUT3 #(
		.INIT('h08)
	) name7493 (
		\m0_cyc_i_pad ,
		\m0_s2_cyc_o_reg/NET0131 ,
		\m0_stb_i_pad ,
		_w9394_
	);
	LUT4 #(
		.INIT('h0004)
	) name7494 (
		\m0_addr_i[28]_pad ,
		\m0_addr_i[29]_pad ,
		\m0_addr_i[30]_pad ,
		\m0_addr_i[31]_pad ,
		_w9395_
	);
	LUT3 #(
		.INIT('hec)
	) name7495 (
		_w9274_,
		_w9394_,
		_w9395_,
		_w9396_
	);
	LUT3 #(
		.INIT('h08)
	) name7496 (
		\m0_cyc_i_pad ,
		\m0_s3_cyc_o_reg/NET0131 ,
		\m0_stb_i_pad ,
		_w9397_
	);
	LUT4 #(
		.INIT('h0008)
	) name7497 (
		\m0_addr_i[28]_pad ,
		\m0_addr_i[29]_pad ,
		\m0_addr_i[30]_pad ,
		\m0_addr_i[31]_pad ,
		_w9398_
	);
	LUT3 #(
		.INIT('hec)
	) name7498 (
		_w9274_,
		_w9397_,
		_w9398_,
		_w9399_
	);
	LUT3 #(
		.INIT('h08)
	) name7499 (
		\m0_cyc_i_pad ,
		\m0_s5_cyc_o_reg/NET0131 ,
		\m0_stb_i_pad ,
		_w9400_
	);
	LUT4 #(
		.INIT('h0020)
	) name7500 (
		\m0_addr_i[28]_pad ,
		\m0_addr_i[29]_pad ,
		\m0_addr_i[30]_pad ,
		\m0_addr_i[31]_pad ,
		_w9401_
	);
	LUT3 #(
		.INIT('hec)
	) name7501 (
		_w9274_,
		_w9400_,
		_w9401_,
		_w9402_
	);
	LUT3 #(
		.INIT('h08)
	) name7502 (
		\m0_cyc_i_pad ,
		\m0_s6_cyc_o_reg/NET0131 ,
		\m0_stb_i_pad ,
		_w9403_
	);
	LUT4 #(
		.INIT('h0040)
	) name7503 (
		\m0_addr_i[28]_pad ,
		\m0_addr_i[29]_pad ,
		\m0_addr_i[30]_pad ,
		\m0_addr_i[31]_pad ,
		_w9404_
	);
	LUT3 #(
		.INIT('hec)
	) name7504 (
		_w9274_,
		_w9403_,
		_w9404_,
		_w9405_
	);
	LUT3 #(
		.INIT('h08)
	) name7505 (
		\m0_cyc_i_pad ,
		\m0_s7_cyc_o_reg/NET0131 ,
		\m0_stb_i_pad ,
		_w9406_
	);
	LUT4 #(
		.INIT('h0080)
	) name7506 (
		\m0_addr_i[28]_pad ,
		\m0_addr_i[29]_pad ,
		\m0_addr_i[30]_pad ,
		\m0_addr_i[31]_pad ,
		_w9407_
	);
	LUT3 #(
		.INIT('hec)
	) name7507 (
		_w9274_,
		_w9406_,
		_w9407_,
		_w9408_
	);
	LUT3 #(
		.INIT('h08)
	) name7508 (
		\m0_cyc_i_pad ,
		\m0_s8_cyc_o_reg/NET0131 ,
		\m0_stb_i_pad ,
		_w9409_
	);
	LUT4 #(
		.INIT('h0100)
	) name7509 (
		\m0_addr_i[28]_pad ,
		\m0_addr_i[29]_pad ,
		\m0_addr_i[30]_pad ,
		\m0_addr_i[31]_pad ,
		_w9410_
	);
	LUT3 #(
		.INIT('hec)
	) name7510 (
		_w9274_,
		_w9409_,
		_w9410_,
		_w9411_
	);
	LUT3 #(
		.INIT('h08)
	) name7511 (
		\m1_cyc_i_pad ,
		\m1_s10_cyc_o_reg/NET0131 ,
		\m1_stb_i_pad ,
		_w9412_
	);
	LUT4 #(
		.INIT('h0400)
	) name7512 (
		\m1_addr_i[28]_pad ,
		\m1_addr_i[29]_pad ,
		\m1_addr_i[30]_pad ,
		\m1_addr_i[31]_pad ,
		_w9413_
	);
	LUT3 #(
		.INIT('hec)
	) name7513 (
		_w9281_,
		_w9412_,
		_w9413_,
		_w9414_
	);
	LUT3 #(
		.INIT('h08)
	) name7514 (
		\m3_cyc_i_pad ,
		\m3_s3_cyc_o_reg/NET0131 ,
		\m3_stb_i_pad ,
		_w9415_
	);
	LUT4 #(
		.INIT('h0008)
	) name7515 (
		\m3_addr_i[28]_pad ,
		\m3_addr_i[29]_pad ,
		\m3_addr_i[30]_pad ,
		\m3_addr_i[31]_pad ,
		_w9416_
	);
	LUT3 #(
		.INIT('hec)
	) name7516 (
		_w9292_,
		_w9415_,
		_w9416_,
		_w9417_
	);
	LUT3 #(
		.INIT('h08)
	) name7517 (
		\m1_cyc_i_pad ,
		\m1_s13_cyc_o_reg/NET0131 ,
		\m1_stb_i_pad ,
		_w9418_
	);
	LUT4 #(
		.INIT('h2000)
	) name7518 (
		\m1_addr_i[28]_pad ,
		\m1_addr_i[29]_pad ,
		\m1_addr_i[30]_pad ,
		\m1_addr_i[31]_pad ,
		_w9419_
	);
	LUT3 #(
		.INIT('hec)
	) name7519 (
		_w9281_,
		_w9418_,
		_w9419_,
		_w9420_
	);
	LUT3 #(
		.INIT('h08)
	) name7520 (
		\m1_cyc_i_pad ,
		\m1_s14_cyc_o_reg/NET0131 ,
		\m1_stb_i_pad ,
		_w9421_
	);
	LUT4 #(
		.INIT('h4000)
	) name7521 (
		\m1_addr_i[28]_pad ,
		\m1_addr_i[29]_pad ,
		\m1_addr_i[30]_pad ,
		\m1_addr_i[31]_pad ,
		_w9422_
	);
	LUT3 #(
		.INIT('hec)
	) name7522 (
		_w9281_,
		_w9421_,
		_w9422_,
		_w9423_
	);
	LUT3 #(
		.INIT('h08)
	) name7523 (
		\m1_cyc_i_pad ,
		\m1_s15_cyc_o_reg/NET0131 ,
		\m1_stb_i_pad ,
		_w9424_
	);
	LUT3 #(
		.INIT('hf8)
	) name7524 (
		_w2047_,
		_w9281_,
		_w9424_,
		_w9425_
	);
	LUT3 #(
		.INIT('h08)
	) name7525 (
		\m1_cyc_i_pad ,
		\m1_s2_cyc_o_reg/NET0131 ,
		\m1_stb_i_pad ,
		_w9426_
	);
	LUT4 #(
		.INIT('h0004)
	) name7526 (
		\m1_addr_i[28]_pad ,
		\m1_addr_i[29]_pad ,
		\m1_addr_i[30]_pad ,
		\m1_addr_i[31]_pad ,
		_w9427_
	);
	LUT3 #(
		.INIT('hec)
	) name7527 (
		_w9281_,
		_w9426_,
		_w9427_,
		_w9428_
	);
	LUT3 #(
		.INIT('h08)
	) name7528 (
		\m1_cyc_i_pad ,
		\m1_s3_cyc_o_reg/NET0131 ,
		\m1_stb_i_pad ,
		_w9429_
	);
	LUT4 #(
		.INIT('h0008)
	) name7529 (
		\m1_addr_i[28]_pad ,
		\m1_addr_i[29]_pad ,
		\m1_addr_i[30]_pad ,
		\m1_addr_i[31]_pad ,
		_w9430_
	);
	LUT3 #(
		.INIT('hec)
	) name7530 (
		_w9281_,
		_w9429_,
		_w9430_,
		_w9431_
	);
	LUT3 #(
		.INIT('h08)
	) name7531 (
		\m1_cyc_i_pad ,
		\m1_s4_cyc_o_reg/NET0131 ,
		\m1_stb_i_pad ,
		_w9432_
	);
	LUT4 #(
		.INIT('h0010)
	) name7532 (
		\m1_addr_i[28]_pad ,
		\m1_addr_i[29]_pad ,
		\m1_addr_i[30]_pad ,
		\m1_addr_i[31]_pad ,
		_w9433_
	);
	LUT3 #(
		.INIT('hec)
	) name7533 (
		_w9281_,
		_w9432_,
		_w9433_,
		_w9434_
	);
	LUT3 #(
		.INIT('h08)
	) name7534 (
		\m1_cyc_i_pad ,
		\m1_s5_cyc_o_reg/NET0131 ,
		\m1_stb_i_pad ,
		_w9435_
	);
	LUT4 #(
		.INIT('h0020)
	) name7535 (
		\m1_addr_i[28]_pad ,
		\m1_addr_i[29]_pad ,
		\m1_addr_i[30]_pad ,
		\m1_addr_i[31]_pad ,
		_w9436_
	);
	LUT3 #(
		.INIT('hec)
	) name7536 (
		_w9281_,
		_w9435_,
		_w9436_,
		_w9437_
	);
	LUT3 #(
		.INIT('h08)
	) name7537 (
		\m1_cyc_i_pad ,
		\m1_s6_cyc_o_reg/NET0131 ,
		\m1_stb_i_pad ,
		_w9438_
	);
	LUT4 #(
		.INIT('h0040)
	) name7538 (
		\m1_addr_i[28]_pad ,
		\m1_addr_i[29]_pad ,
		\m1_addr_i[30]_pad ,
		\m1_addr_i[31]_pad ,
		_w9439_
	);
	LUT3 #(
		.INIT('hec)
	) name7539 (
		_w9281_,
		_w9438_,
		_w9439_,
		_w9440_
	);
	LUT3 #(
		.INIT('h08)
	) name7540 (
		\m1_cyc_i_pad ,
		\m1_s7_cyc_o_reg/NET0131 ,
		\m1_stb_i_pad ,
		_w9441_
	);
	LUT4 #(
		.INIT('h0080)
	) name7541 (
		\m1_addr_i[28]_pad ,
		\m1_addr_i[29]_pad ,
		\m1_addr_i[30]_pad ,
		\m1_addr_i[31]_pad ,
		_w9442_
	);
	LUT3 #(
		.INIT('hec)
	) name7542 (
		_w9281_,
		_w9441_,
		_w9442_,
		_w9443_
	);
	LUT3 #(
		.INIT('h08)
	) name7543 (
		\m1_cyc_i_pad ,
		\m1_s8_cyc_o_reg/NET0131 ,
		\m1_stb_i_pad ,
		_w9444_
	);
	LUT4 #(
		.INIT('h0100)
	) name7544 (
		\m1_addr_i[28]_pad ,
		\m1_addr_i[29]_pad ,
		\m1_addr_i[30]_pad ,
		\m1_addr_i[31]_pad ,
		_w9445_
	);
	LUT3 #(
		.INIT('hec)
	) name7545 (
		_w9281_,
		_w9444_,
		_w9445_,
		_w9446_
	);
	LUT3 #(
		.INIT('h08)
	) name7546 (
		\m1_cyc_i_pad ,
		\m1_s9_cyc_o_reg/NET0131 ,
		\m1_stb_i_pad ,
		_w9447_
	);
	LUT4 #(
		.INIT('h0200)
	) name7547 (
		\m1_addr_i[28]_pad ,
		\m1_addr_i[29]_pad ,
		\m1_addr_i[30]_pad ,
		\m1_addr_i[31]_pad ,
		_w9448_
	);
	LUT3 #(
		.INIT('hec)
	) name7548 (
		_w9281_,
		_w9447_,
		_w9448_,
		_w9449_
	);
	LUT3 #(
		.INIT('h08)
	) name7549 (
		\m2_cyc_i_pad ,
		\m2_s10_cyc_o_reg/NET0131 ,
		\m2_stb_i_pad ,
		_w9450_
	);
	LUT4 #(
		.INIT('h0400)
	) name7550 (
		\m2_addr_i[28]_pad ,
		\m2_addr_i[29]_pad ,
		\m2_addr_i[30]_pad ,
		\m2_addr_i[31]_pad ,
		_w9451_
	);
	LUT3 #(
		.INIT('hec)
	) name7551 (
		_w9285_,
		_w9450_,
		_w9451_,
		_w9452_
	);
	LUT3 #(
		.INIT('h08)
	) name7552 (
		\m2_cyc_i_pad ,
		\m2_s11_cyc_o_reg/NET0131 ,
		\m2_stb_i_pad ,
		_w9453_
	);
	LUT4 #(
		.INIT('h0800)
	) name7553 (
		\m2_addr_i[28]_pad ,
		\m2_addr_i[29]_pad ,
		\m2_addr_i[30]_pad ,
		\m2_addr_i[31]_pad ,
		_w9454_
	);
	LUT3 #(
		.INIT('hec)
	) name7554 (
		_w9285_,
		_w9453_,
		_w9454_,
		_w9455_
	);
	LUT3 #(
		.INIT('h08)
	) name7555 (
		\m2_cyc_i_pad ,
		\m2_s12_cyc_o_reg/NET0131 ,
		\m2_stb_i_pad ,
		_w9456_
	);
	LUT4 #(
		.INIT('h1000)
	) name7556 (
		\m2_addr_i[28]_pad ,
		\m2_addr_i[29]_pad ,
		\m2_addr_i[30]_pad ,
		\m2_addr_i[31]_pad ,
		_w9457_
	);
	LUT3 #(
		.INIT('hec)
	) name7557 (
		_w9285_,
		_w9456_,
		_w9457_,
		_w9458_
	);
	LUT3 #(
		.INIT('h08)
	) name7558 (
		\m2_cyc_i_pad ,
		\m2_s15_cyc_o_reg/NET0131 ,
		\m2_stb_i_pad ,
		_w9459_
	);
	LUT3 #(
		.INIT('hf8)
	) name7559 (
		_w2057_,
		_w9285_,
		_w9459_,
		_w9460_
	);
	LUT3 #(
		.INIT('h08)
	) name7560 (
		\m2_cyc_i_pad ,
		\m2_s2_cyc_o_reg/NET0131 ,
		\m2_stb_i_pad ,
		_w9461_
	);
	LUT4 #(
		.INIT('h0004)
	) name7561 (
		\m2_addr_i[28]_pad ,
		\m2_addr_i[29]_pad ,
		\m2_addr_i[30]_pad ,
		\m2_addr_i[31]_pad ,
		_w9462_
	);
	LUT3 #(
		.INIT('hec)
	) name7562 (
		_w9285_,
		_w9461_,
		_w9462_,
		_w9463_
	);
	LUT3 #(
		.INIT('h08)
	) name7563 (
		\m2_cyc_i_pad ,
		\m2_s3_cyc_o_reg/NET0131 ,
		\m2_stb_i_pad ,
		_w9464_
	);
	LUT4 #(
		.INIT('h0008)
	) name7564 (
		\m2_addr_i[28]_pad ,
		\m2_addr_i[29]_pad ,
		\m2_addr_i[30]_pad ,
		\m2_addr_i[31]_pad ,
		_w9465_
	);
	LUT3 #(
		.INIT('hec)
	) name7565 (
		_w9285_,
		_w9464_,
		_w9465_,
		_w9466_
	);
	LUT3 #(
		.INIT('h08)
	) name7566 (
		\m2_cyc_i_pad ,
		\m2_s4_cyc_o_reg/NET0131 ,
		\m2_stb_i_pad ,
		_w9467_
	);
	LUT4 #(
		.INIT('h0010)
	) name7567 (
		\m2_addr_i[28]_pad ,
		\m2_addr_i[29]_pad ,
		\m2_addr_i[30]_pad ,
		\m2_addr_i[31]_pad ,
		_w9468_
	);
	LUT3 #(
		.INIT('hec)
	) name7568 (
		_w9285_,
		_w9467_,
		_w9468_,
		_w9469_
	);
	LUT3 #(
		.INIT('h08)
	) name7569 (
		\m2_cyc_i_pad ,
		\m2_s5_cyc_o_reg/NET0131 ,
		\m2_stb_i_pad ,
		_w9470_
	);
	LUT4 #(
		.INIT('h0020)
	) name7570 (
		\m2_addr_i[28]_pad ,
		\m2_addr_i[29]_pad ,
		\m2_addr_i[30]_pad ,
		\m2_addr_i[31]_pad ,
		_w9471_
	);
	LUT3 #(
		.INIT('hec)
	) name7571 (
		_w9285_,
		_w9470_,
		_w9471_,
		_w9472_
	);
	LUT3 #(
		.INIT('h08)
	) name7572 (
		\m2_cyc_i_pad ,
		\m2_s6_cyc_o_reg/NET0131 ,
		\m2_stb_i_pad ,
		_w9473_
	);
	LUT4 #(
		.INIT('h0040)
	) name7573 (
		\m2_addr_i[28]_pad ,
		\m2_addr_i[29]_pad ,
		\m2_addr_i[30]_pad ,
		\m2_addr_i[31]_pad ,
		_w9474_
	);
	LUT3 #(
		.INIT('hec)
	) name7574 (
		_w9285_,
		_w9473_,
		_w9474_,
		_w9475_
	);
	LUT3 #(
		.INIT('h08)
	) name7575 (
		\m2_cyc_i_pad ,
		\m2_s9_cyc_o_reg/NET0131 ,
		\m2_stb_i_pad ,
		_w9476_
	);
	LUT4 #(
		.INIT('h0200)
	) name7576 (
		\m2_addr_i[28]_pad ,
		\m2_addr_i[29]_pad ,
		\m2_addr_i[30]_pad ,
		\m2_addr_i[31]_pad ,
		_w9477_
	);
	LUT3 #(
		.INIT('hec)
	) name7577 (
		_w9285_,
		_w9476_,
		_w9477_,
		_w9478_
	);
	LUT3 #(
		.INIT('h08)
	) name7578 (
		\m3_cyc_i_pad ,
		\m3_s10_cyc_o_reg/NET0131 ,
		\m3_stb_i_pad ,
		_w9479_
	);
	LUT4 #(
		.INIT('h0400)
	) name7579 (
		\m3_addr_i[28]_pad ,
		\m3_addr_i[29]_pad ,
		\m3_addr_i[30]_pad ,
		\m3_addr_i[31]_pad ,
		_w9480_
	);
	LUT3 #(
		.INIT('hec)
	) name7580 (
		_w9292_,
		_w9479_,
		_w9480_,
		_w9481_
	);
	LUT3 #(
		.INIT('h08)
	) name7581 (
		\m3_cyc_i_pad ,
		\m3_s11_cyc_o_reg/NET0131 ,
		\m3_stb_i_pad ,
		_w9482_
	);
	LUT4 #(
		.INIT('h0800)
	) name7582 (
		\m3_addr_i[28]_pad ,
		\m3_addr_i[29]_pad ,
		\m3_addr_i[30]_pad ,
		\m3_addr_i[31]_pad ,
		_w9483_
	);
	LUT3 #(
		.INIT('hec)
	) name7583 (
		_w9292_,
		_w9482_,
		_w9483_,
		_w9484_
	);
	LUT3 #(
		.INIT('h08)
	) name7584 (
		\m3_cyc_i_pad ,
		\m3_s12_cyc_o_reg/NET0131 ,
		\m3_stb_i_pad ,
		_w9485_
	);
	LUT4 #(
		.INIT('h1000)
	) name7585 (
		\m3_addr_i[28]_pad ,
		\m3_addr_i[29]_pad ,
		\m3_addr_i[30]_pad ,
		\m3_addr_i[31]_pad ,
		_w9486_
	);
	LUT3 #(
		.INIT('hec)
	) name7586 (
		_w9292_,
		_w9485_,
		_w9486_,
		_w9487_
	);
	LUT3 #(
		.INIT('h08)
	) name7587 (
		\m3_cyc_i_pad ,
		\m3_s13_cyc_o_reg/NET0131 ,
		\m3_stb_i_pad ,
		_w9488_
	);
	LUT4 #(
		.INIT('h2000)
	) name7588 (
		\m3_addr_i[28]_pad ,
		\m3_addr_i[29]_pad ,
		\m3_addr_i[30]_pad ,
		\m3_addr_i[31]_pad ,
		_w9489_
	);
	LUT3 #(
		.INIT('hec)
	) name7589 (
		_w9292_,
		_w9488_,
		_w9489_,
		_w9490_
	);
	LUT3 #(
		.INIT('h08)
	) name7590 (
		\m3_cyc_i_pad ,
		\m3_s15_cyc_o_reg/NET0131 ,
		\m3_stb_i_pad ,
		_w9491_
	);
	LUT3 #(
		.INIT('hf8)
	) name7591 (
		_w2059_,
		_w9292_,
		_w9491_,
		_w9492_
	);
	LUT3 #(
		.INIT('h08)
	) name7592 (
		\m3_cyc_i_pad ,
		\m3_s2_cyc_o_reg/NET0131 ,
		\m3_stb_i_pad ,
		_w9493_
	);
	LUT4 #(
		.INIT('h0004)
	) name7593 (
		\m3_addr_i[28]_pad ,
		\m3_addr_i[29]_pad ,
		\m3_addr_i[30]_pad ,
		\m3_addr_i[31]_pad ,
		_w9494_
	);
	LUT3 #(
		.INIT('hec)
	) name7594 (
		_w9292_,
		_w9493_,
		_w9494_,
		_w9495_
	);
	LUT3 #(
		.INIT('h08)
	) name7595 (
		\m3_cyc_i_pad ,
		\m3_s14_cyc_o_reg/NET0131 ,
		\m3_stb_i_pad ,
		_w9496_
	);
	LUT4 #(
		.INIT('h4000)
	) name7596 (
		\m3_addr_i[28]_pad ,
		\m3_addr_i[29]_pad ,
		\m3_addr_i[30]_pad ,
		\m3_addr_i[31]_pad ,
		_w9497_
	);
	LUT3 #(
		.INIT('hec)
	) name7597 (
		_w9292_,
		_w9496_,
		_w9497_,
		_w9498_
	);
	LUT3 #(
		.INIT('h08)
	) name7598 (
		\m3_cyc_i_pad ,
		\m3_s4_cyc_o_reg/NET0131 ,
		\m3_stb_i_pad ,
		_w9499_
	);
	LUT4 #(
		.INIT('h0010)
	) name7599 (
		\m3_addr_i[28]_pad ,
		\m3_addr_i[29]_pad ,
		\m3_addr_i[30]_pad ,
		\m3_addr_i[31]_pad ,
		_w9500_
	);
	LUT3 #(
		.INIT('hec)
	) name7600 (
		_w9292_,
		_w9499_,
		_w9500_,
		_w9501_
	);
	LUT3 #(
		.INIT('h08)
	) name7601 (
		\m3_cyc_i_pad ,
		\m3_s8_cyc_o_reg/NET0131 ,
		\m3_stb_i_pad ,
		_w9502_
	);
	LUT4 #(
		.INIT('h0100)
	) name7602 (
		\m3_addr_i[28]_pad ,
		\m3_addr_i[29]_pad ,
		\m3_addr_i[30]_pad ,
		\m3_addr_i[31]_pad ,
		_w9503_
	);
	LUT3 #(
		.INIT('hec)
	) name7603 (
		_w9292_,
		_w9502_,
		_w9503_,
		_w9504_
	);
	LUT3 #(
		.INIT('h08)
	) name7604 (
		\m3_cyc_i_pad ,
		\m3_s9_cyc_o_reg/NET0131 ,
		\m3_stb_i_pad ,
		_w9505_
	);
	LUT4 #(
		.INIT('h0200)
	) name7605 (
		\m3_addr_i[28]_pad ,
		\m3_addr_i[29]_pad ,
		\m3_addr_i[30]_pad ,
		\m3_addr_i[31]_pad ,
		_w9506_
	);
	LUT3 #(
		.INIT('hec)
	) name7606 (
		_w9292_,
		_w9505_,
		_w9506_,
		_w9507_
	);
	LUT3 #(
		.INIT('h08)
	) name7607 (
		\m4_cyc_i_pad ,
		\m4_s10_cyc_o_reg/NET0131 ,
		\m4_stb_i_pad ,
		_w9508_
	);
	LUT4 #(
		.INIT('h0400)
	) name7608 (
		\m4_addr_i[28]_pad ,
		\m4_addr_i[29]_pad ,
		\m4_addr_i[30]_pad ,
		\m4_addr_i[31]_pad ,
		_w9509_
	);
	LUT3 #(
		.INIT('hec)
	) name7609 (
		_w9299_,
		_w9508_,
		_w9509_,
		_w9510_
	);
	LUT3 #(
		.INIT('h08)
	) name7610 (
		\m4_cyc_i_pad ,
		\m4_s12_cyc_o_reg/NET0131 ,
		\m4_stb_i_pad ,
		_w9511_
	);
	LUT4 #(
		.INIT('h1000)
	) name7611 (
		\m4_addr_i[28]_pad ,
		\m4_addr_i[29]_pad ,
		\m4_addr_i[30]_pad ,
		\m4_addr_i[31]_pad ,
		_w9512_
	);
	LUT3 #(
		.INIT('hec)
	) name7612 (
		_w9299_,
		_w9511_,
		_w9512_,
		_w9513_
	);
	LUT3 #(
		.INIT('h08)
	) name7613 (
		\m4_cyc_i_pad ,
		\m4_s14_cyc_o_reg/NET0131 ,
		\m4_stb_i_pad ,
		_w9514_
	);
	LUT4 #(
		.INIT('h4000)
	) name7614 (
		\m4_addr_i[28]_pad ,
		\m4_addr_i[29]_pad ,
		\m4_addr_i[30]_pad ,
		\m4_addr_i[31]_pad ,
		_w9515_
	);
	LUT3 #(
		.INIT('hec)
	) name7615 (
		_w9299_,
		_w9514_,
		_w9515_,
		_w9516_
	);
	LUT3 #(
		.INIT('h08)
	) name7616 (
		\m4_cyc_i_pad ,
		\m4_s15_cyc_o_reg/NET0131 ,
		\m4_stb_i_pad ,
		_w9517_
	);
	LUT3 #(
		.INIT('hf8)
	) name7617 (
		_w2062_,
		_w9299_,
		_w9517_,
		_w9518_
	);
	LUT3 #(
		.INIT('h08)
	) name7618 (
		\m4_cyc_i_pad ,
		\m4_s2_cyc_o_reg/NET0131 ,
		\m4_stb_i_pad ,
		_w9519_
	);
	LUT4 #(
		.INIT('h0004)
	) name7619 (
		\m4_addr_i[28]_pad ,
		\m4_addr_i[29]_pad ,
		\m4_addr_i[30]_pad ,
		\m4_addr_i[31]_pad ,
		_w9520_
	);
	LUT3 #(
		.INIT('hec)
	) name7620 (
		_w9299_,
		_w9519_,
		_w9520_,
		_w9521_
	);
	LUT3 #(
		.INIT('h08)
	) name7621 (
		\m4_cyc_i_pad ,
		\m4_s3_cyc_o_reg/NET0131 ,
		\m4_stb_i_pad ,
		_w9522_
	);
	LUT4 #(
		.INIT('h0008)
	) name7622 (
		\m4_addr_i[28]_pad ,
		\m4_addr_i[29]_pad ,
		\m4_addr_i[30]_pad ,
		\m4_addr_i[31]_pad ,
		_w9523_
	);
	LUT3 #(
		.INIT('hec)
	) name7623 (
		_w9299_,
		_w9522_,
		_w9523_,
		_w9524_
	);
	LUT3 #(
		.INIT('h08)
	) name7624 (
		\m4_cyc_i_pad ,
		\m4_s5_cyc_o_reg/NET0131 ,
		\m4_stb_i_pad ,
		_w9525_
	);
	LUT4 #(
		.INIT('h0020)
	) name7625 (
		\m4_addr_i[28]_pad ,
		\m4_addr_i[29]_pad ,
		\m4_addr_i[30]_pad ,
		\m4_addr_i[31]_pad ,
		_w9526_
	);
	LUT3 #(
		.INIT('hec)
	) name7626 (
		_w9299_,
		_w9525_,
		_w9526_,
		_w9527_
	);
	LUT3 #(
		.INIT('h08)
	) name7627 (
		\m4_cyc_i_pad ,
		\m4_s7_cyc_o_reg/NET0131 ,
		\m4_stb_i_pad ,
		_w9528_
	);
	LUT4 #(
		.INIT('h0080)
	) name7628 (
		\m4_addr_i[28]_pad ,
		\m4_addr_i[29]_pad ,
		\m4_addr_i[30]_pad ,
		\m4_addr_i[31]_pad ,
		_w9529_
	);
	LUT3 #(
		.INIT('hec)
	) name7629 (
		_w9299_,
		_w9528_,
		_w9529_,
		_w9530_
	);
	LUT3 #(
		.INIT('h08)
	) name7630 (
		\m5_cyc_i_pad ,
		\m5_s10_cyc_o_reg/NET0131 ,
		\m5_stb_i_pad ,
		_w9531_
	);
	LUT4 #(
		.INIT('h0400)
	) name7631 (
		\m5_addr_i[28]_pad ,
		\m5_addr_i[29]_pad ,
		\m5_addr_i[30]_pad ,
		\m5_addr_i[31]_pad ,
		_w9532_
	);
	LUT3 #(
		.INIT('hec)
	) name7632 (
		_w9270_,
		_w9531_,
		_w9532_,
		_w9533_
	);
	LUT3 #(
		.INIT('h08)
	) name7633 (
		\m5_cyc_i_pad ,
		\m5_s11_cyc_o_reg/NET0131 ,
		\m5_stb_i_pad ,
		_w9534_
	);
	LUT4 #(
		.INIT('h0800)
	) name7634 (
		\m5_addr_i[28]_pad ,
		\m5_addr_i[29]_pad ,
		\m5_addr_i[30]_pad ,
		\m5_addr_i[31]_pad ,
		_w9535_
	);
	LUT3 #(
		.INIT('hec)
	) name7635 (
		_w9270_,
		_w9534_,
		_w9535_,
		_w9536_
	);
	LUT3 #(
		.INIT('h08)
	) name7636 (
		\m5_cyc_i_pad ,
		\m5_s13_cyc_o_reg/NET0131 ,
		\m5_stb_i_pad ,
		_w9537_
	);
	LUT4 #(
		.INIT('h2000)
	) name7637 (
		\m5_addr_i[28]_pad ,
		\m5_addr_i[29]_pad ,
		\m5_addr_i[30]_pad ,
		\m5_addr_i[31]_pad ,
		_w9538_
	);
	LUT3 #(
		.INIT('hec)
	) name7638 (
		_w9270_,
		_w9537_,
		_w9538_,
		_w9539_
	);
	LUT3 #(
		.INIT('h08)
	) name7639 (
		\m5_cyc_i_pad ,
		\m5_s2_cyc_o_reg/NET0131 ,
		\m5_stb_i_pad ,
		_w9540_
	);
	LUT4 #(
		.INIT('h0004)
	) name7640 (
		\m5_addr_i[28]_pad ,
		\m5_addr_i[29]_pad ,
		\m5_addr_i[30]_pad ,
		\m5_addr_i[31]_pad ,
		_w9541_
	);
	LUT3 #(
		.INIT('hec)
	) name7641 (
		_w9270_,
		_w9540_,
		_w9541_,
		_w9542_
	);
	LUT3 #(
		.INIT('h08)
	) name7642 (
		\m5_cyc_i_pad ,
		\m5_s4_cyc_o_reg/NET0131 ,
		\m5_stb_i_pad ,
		_w9543_
	);
	LUT4 #(
		.INIT('h0010)
	) name7643 (
		\m5_addr_i[28]_pad ,
		\m5_addr_i[29]_pad ,
		\m5_addr_i[30]_pad ,
		\m5_addr_i[31]_pad ,
		_w9544_
	);
	LUT3 #(
		.INIT('hec)
	) name7644 (
		_w9270_,
		_w9543_,
		_w9544_,
		_w9545_
	);
	LUT3 #(
		.INIT('h08)
	) name7645 (
		\m5_cyc_i_pad ,
		\m5_s5_cyc_o_reg/NET0131 ,
		\m5_stb_i_pad ,
		_w9546_
	);
	LUT4 #(
		.INIT('h0020)
	) name7646 (
		\m5_addr_i[28]_pad ,
		\m5_addr_i[29]_pad ,
		\m5_addr_i[30]_pad ,
		\m5_addr_i[31]_pad ,
		_w9547_
	);
	LUT3 #(
		.INIT('hec)
	) name7647 (
		_w9270_,
		_w9546_,
		_w9547_,
		_w9548_
	);
	LUT3 #(
		.INIT('h08)
	) name7648 (
		\m5_cyc_i_pad ,
		\m5_s6_cyc_o_reg/NET0131 ,
		\m5_stb_i_pad ,
		_w9549_
	);
	LUT4 #(
		.INIT('h0040)
	) name7649 (
		\m5_addr_i[28]_pad ,
		\m5_addr_i[29]_pad ,
		\m5_addr_i[30]_pad ,
		\m5_addr_i[31]_pad ,
		_w9550_
	);
	LUT3 #(
		.INIT('hec)
	) name7650 (
		_w9270_,
		_w9549_,
		_w9550_,
		_w9551_
	);
	LUT3 #(
		.INIT('h08)
	) name7651 (
		\m5_cyc_i_pad ,
		\m5_s8_cyc_o_reg/NET0131 ,
		\m5_stb_i_pad ,
		_w9552_
	);
	LUT4 #(
		.INIT('h0100)
	) name7652 (
		\m5_addr_i[28]_pad ,
		\m5_addr_i[29]_pad ,
		\m5_addr_i[30]_pad ,
		\m5_addr_i[31]_pad ,
		_w9553_
	);
	LUT3 #(
		.INIT('hec)
	) name7653 (
		_w9270_,
		_w9552_,
		_w9553_,
		_w9554_
	);
	LUT3 #(
		.INIT('h08)
	) name7654 (
		\m5_cyc_i_pad ,
		\m5_s9_cyc_o_reg/NET0131 ,
		\m5_stb_i_pad ,
		_w9555_
	);
	LUT4 #(
		.INIT('h0200)
	) name7655 (
		\m5_addr_i[28]_pad ,
		\m5_addr_i[29]_pad ,
		\m5_addr_i[30]_pad ,
		\m5_addr_i[31]_pad ,
		_w9556_
	);
	LUT3 #(
		.INIT('hec)
	) name7656 (
		_w9270_,
		_w9555_,
		_w9556_,
		_w9557_
	);
	LUT3 #(
		.INIT('h08)
	) name7657 (
		\m6_cyc_i_pad ,
		\m6_s10_cyc_o_reg/NET0131 ,
		\m6_stb_i_pad ,
		_w9558_
	);
	LUT4 #(
		.INIT('h0400)
	) name7658 (
		\m6_addr_i[28]_pad ,
		\m6_addr_i[29]_pad ,
		\m6_addr_i[30]_pad ,
		\m6_addr_i[31]_pad ,
		_w9559_
	);
	LUT3 #(
		.INIT('hec)
	) name7659 (
		_w9309_,
		_w9558_,
		_w9559_,
		_w9560_
	);
	LUT3 #(
		.INIT('h08)
	) name7660 (
		\m6_cyc_i_pad ,
		\m6_s11_cyc_o_reg/NET0131 ,
		\m6_stb_i_pad ,
		_w9561_
	);
	LUT4 #(
		.INIT('h0800)
	) name7661 (
		\m6_addr_i[28]_pad ,
		\m6_addr_i[29]_pad ,
		\m6_addr_i[30]_pad ,
		\m6_addr_i[31]_pad ,
		_w9562_
	);
	LUT3 #(
		.INIT('hec)
	) name7662 (
		_w9309_,
		_w9561_,
		_w9562_,
		_w9563_
	);
	LUT3 #(
		.INIT('h08)
	) name7663 (
		\m6_cyc_i_pad ,
		\m6_s12_cyc_o_reg/NET0131 ,
		\m6_stb_i_pad ,
		_w9564_
	);
	LUT4 #(
		.INIT('h1000)
	) name7664 (
		\m6_addr_i[28]_pad ,
		\m6_addr_i[29]_pad ,
		\m6_addr_i[30]_pad ,
		\m6_addr_i[31]_pad ,
		_w9565_
	);
	LUT3 #(
		.INIT('hec)
	) name7665 (
		_w9309_,
		_w9564_,
		_w9565_,
		_w9566_
	);
	LUT3 #(
		.INIT('h08)
	) name7666 (
		\m6_cyc_i_pad ,
		\m6_s13_cyc_o_reg/NET0131 ,
		\m6_stb_i_pad ,
		_w9567_
	);
	LUT4 #(
		.INIT('h2000)
	) name7667 (
		\m6_addr_i[28]_pad ,
		\m6_addr_i[29]_pad ,
		\m6_addr_i[30]_pad ,
		\m6_addr_i[31]_pad ,
		_w9568_
	);
	LUT3 #(
		.INIT('hec)
	) name7668 (
		_w9309_,
		_w9567_,
		_w9568_,
		_w9569_
	);
	LUT3 #(
		.INIT('h08)
	) name7669 (
		\m6_cyc_i_pad ,
		\m6_s14_cyc_o_reg/NET0131 ,
		\m6_stb_i_pad ,
		_w9570_
	);
	LUT4 #(
		.INIT('h4000)
	) name7670 (
		\m6_addr_i[28]_pad ,
		\m6_addr_i[29]_pad ,
		\m6_addr_i[30]_pad ,
		\m6_addr_i[31]_pad ,
		_w9571_
	);
	LUT3 #(
		.INIT('hec)
	) name7671 (
		_w9309_,
		_w9570_,
		_w9571_,
		_w9572_
	);
	LUT3 #(
		.INIT('h08)
	) name7672 (
		\m6_cyc_i_pad ,
		\m6_s15_cyc_o_reg/NET0131 ,
		\m6_stb_i_pad ,
		_w9573_
	);
	LUT3 #(
		.INIT('hf8)
	) name7673 (
		_w2054_,
		_w9309_,
		_w9573_,
		_w9574_
	);
	LUT3 #(
		.INIT('h08)
	) name7674 (
		\m6_cyc_i_pad ,
		\m6_s2_cyc_o_reg/NET0131 ,
		\m6_stb_i_pad ,
		_w9575_
	);
	LUT4 #(
		.INIT('h0004)
	) name7675 (
		\m6_addr_i[28]_pad ,
		\m6_addr_i[29]_pad ,
		\m6_addr_i[30]_pad ,
		\m6_addr_i[31]_pad ,
		_w9576_
	);
	LUT3 #(
		.INIT('hec)
	) name7676 (
		_w9309_,
		_w9575_,
		_w9576_,
		_w9577_
	);
	LUT3 #(
		.INIT('h08)
	) name7677 (
		\m6_cyc_i_pad ,
		\m6_s3_cyc_o_reg/NET0131 ,
		\m6_stb_i_pad ,
		_w9578_
	);
	LUT4 #(
		.INIT('h0008)
	) name7678 (
		\m6_addr_i[28]_pad ,
		\m6_addr_i[29]_pad ,
		\m6_addr_i[30]_pad ,
		\m6_addr_i[31]_pad ,
		_w9579_
	);
	LUT3 #(
		.INIT('hec)
	) name7679 (
		_w9309_,
		_w9578_,
		_w9579_,
		_w9580_
	);
	LUT3 #(
		.INIT('h08)
	) name7680 (
		\m6_cyc_i_pad ,
		\m6_s4_cyc_o_reg/NET0131 ,
		\m6_stb_i_pad ,
		_w9581_
	);
	LUT4 #(
		.INIT('h0010)
	) name7681 (
		\m6_addr_i[28]_pad ,
		\m6_addr_i[29]_pad ,
		\m6_addr_i[30]_pad ,
		\m6_addr_i[31]_pad ,
		_w9582_
	);
	LUT3 #(
		.INIT('hec)
	) name7682 (
		_w9309_,
		_w9581_,
		_w9582_,
		_w9583_
	);
	LUT3 #(
		.INIT('h08)
	) name7683 (
		\m6_cyc_i_pad ,
		\m6_s5_cyc_o_reg/NET0131 ,
		\m6_stb_i_pad ,
		_w9584_
	);
	LUT4 #(
		.INIT('h0020)
	) name7684 (
		\m6_addr_i[28]_pad ,
		\m6_addr_i[29]_pad ,
		\m6_addr_i[30]_pad ,
		\m6_addr_i[31]_pad ,
		_w9585_
	);
	LUT3 #(
		.INIT('hec)
	) name7685 (
		_w9309_,
		_w9584_,
		_w9585_,
		_w9586_
	);
	LUT3 #(
		.INIT('h08)
	) name7686 (
		\m6_cyc_i_pad ,
		\m6_s7_cyc_o_reg/NET0131 ,
		\m6_stb_i_pad ,
		_w9587_
	);
	LUT4 #(
		.INIT('h0080)
	) name7687 (
		\m6_addr_i[28]_pad ,
		\m6_addr_i[29]_pad ,
		\m6_addr_i[30]_pad ,
		\m6_addr_i[31]_pad ,
		_w9588_
	);
	LUT3 #(
		.INIT('hec)
	) name7688 (
		_w9309_,
		_w9587_,
		_w9588_,
		_w9589_
	);
	LUT3 #(
		.INIT('h08)
	) name7689 (
		\m6_cyc_i_pad ,
		\m6_s9_cyc_o_reg/NET0131 ,
		\m6_stb_i_pad ,
		_w9590_
	);
	LUT4 #(
		.INIT('h0200)
	) name7690 (
		\m6_addr_i[28]_pad ,
		\m6_addr_i[29]_pad ,
		\m6_addr_i[30]_pad ,
		\m6_addr_i[31]_pad ,
		_w9591_
	);
	LUT3 #(
		.INIT('hec)
	) name7691 (
		_w9309_,
		_w9590_,
		_w9591_,
		_w9592_
	);
	LUT3 #(
		.INIT('h08)
	) name7692 (
		\m7_cyc_i_pad ,
		\m7_s10_cyc_o_reg/NET0131 ,
		\m7_stb_i_pad ,
		_w9593_
	);
	LUT4 #(
		.INIT('h0400)
	) name7693 (
		\m7_addr_i[28]_pad ,
		\m7_addr_i[29]_pad ,
		\m7_addr_i[30]_pad ,
		\m7_addr_i[31]_pad ,
		_w9594_
	);
	LUT3 #(
		.INIT('hec)
	) name7694 (
		_w9316_,
		_w9593_,
		_w9594_,
		_w9595_
	);
	LUT3 #(
		.INIT('h08)
	) name7695 (
		\m7_cyc_i_pad ,
		\m7_s11_cyc_o_reg/NET0131 ,
		\m7_stb_i_pad ,
		_w9596_
	);
	LUT4 #(
		.INIT('h0800)
	) name7696 (
		\m7_addr_i[28]_pad ,
		\m7_addr_i[29]_pad ,
		\m7_addr_i[30]_pad ,
		\m7_addr_i[31]_pad ,
		_w9597_
	);
	LUT3 #(
		.INIT('hec)
	) name7697 (
		_w9316_,
		_w9596_,
		_w9597_,
		_w9598_
	);
	LUT3 #(
		.INIT('h08)
	) name7698 (
		\m7_cyc_i_pad ,
		\m7_s13_cyc_o_reg/NET0131 ,
		\m7_stb_i_pad ,
		_w9599_
	);
	LUT4 #(
		.INIT('h2000)
	) name7699 (
		\m7_addr_i[28]_pad ,
		\m7_addr_i[29]_pad ,
		\m7_addr_i[30]_pad ,
		\m7_addr_i[31]_pad ,
		_w9600_
	);
	LUT3 #(
		.INIT('hec)
	) name7700 (
		_w9316_,
		_w9599_,
		_w9600_,
		_w9601_
	);
	LUT3 #(
		.INIT('h08)
	) name7701 (
		\m7_cyc_i_pad ,
		\m7_s14_cyc_o_reg/NET0131 ,
		\m7_stb_i_pad ,
		_w9602_
	);
	LUT4 #(
		.INIT('h4000)
	) name7702 (
		\m7_addr_i[28]_pad ,
		\m7_addr_i[29]_pad ,
		\m7_addr_i[30]_pad ,
		\m7_addr_i[31]_pad ,
		_w9603_
	);
	LUT3 #(
		.INIT('hec)
	) name7703 (
		_w9316_,
		_w9602_,
		_w9603_,
		_w9604_
	);
	LUT3 #(
		.INIT('h08)
	) name7704 (
		\m7_cyc_i_pad ,
		\m7_s15_cyc_o_reg/NET0131 ,
		\m7_stb_i_pad ,
		_w9605_
	);
	LUT3 #(
		.INIT('hf8)
	) name7705 (
		_w2052_,
		_w9316_,
		_w9605_,
		_w9606_
	);
	LUT3 #(
		.INIT('h08)
	) name7706 (
		\m7_cyc_i_pad ,
		\m7_s2_cyc_o_reg/NET0131 ,
		\m7_stb_i_pad ,
		_w9607_
	);
	LUT4 #(
		.INIT('h0004)
	) name7707 (
		\m7_addr_i[28]_pad ,
		\m7_addr_i[29]_pad ,
		\m7_addr_i[30]_pad ,
		\m7_addr_i[31]_pad ,
		_w9608_
	);
	LUT3 #(
		.INIT('hec)
	) name7708 (
		_w9316_,
		_w9607_,
		_w9608_,
		_w9609_
	);
	LUT3 #(
		.INIT('h08)
	) name7709 (
		\m7_cyc_i_pad ,
		\m7_s3_cyc_o_reg/NET0131 ,
		\m7_stb_i_pad ,
		_w9610_
	);
	LUT4 #(
		.INIT('h0008)
	) name7710 (
		\m7_addr_i[28]_pad ,
		\m7_addr_i[29]_pad ,
		\m7_addr_i[30]_pad ,
		\m7_addr_i[31]_pad ,
		_w9611_
	);
	LUT3 #(
		.INIT('hec)
	) name7711 (
		_w9316_,
		_w9610_,
		_w9611_,
		_w9612_
	);
	LUT3 #(
		.INIT('h08)
	) name7712 (
		\m7_cyc_i_pad ,
		\m7_s4_cyc_o_reg/NET0131 ,
		\m7_stb_i_pad ,
		_w9613_
	);
	LUT4 #(
		.INIT('h0010)
	) name7713 (
		\m7_addr_i[28]_pad ,
		\m7_addr_i[29]_pad ,
		\m7_addr_i[30]_pad ,
		\m7_addr_i[31]_pad ,
		_w9614_
	);
	LUT3 #(
		.INIT('hec)
	) name7714 (
		_w9316_,
		_w9613_,
		_w9614_,
		_w9615_
	);
	LUT3 #(
		.INIT('h08)
	) name7715 (
		\m7_cyc_i_pad ,
		\m7_s6_cyc_o_reg/NET0131 ,
		\m7_stb_i_pad ,
		_w9616_
	);
	LUT4 #(
		.INIT('h0040)
	) name7716 (
		\m7_addr_i[28]_pad ,
		\m7_addr_i[29]_pad ,
		\m7_addr_i[30]_pad ,
		\m7_addr_i[31]_pad ,
		_w9617_
	);
	LUT3 #(
		.INIT('hec)
	) name7717 (
		_w9316_,
		_w9616_,
		_w9617_,
		_w9618_
	);
	LUT3 #(
		.INIT('h08)
	) name7718 (
		\m2_cyc_i_pad ,
		\m2_s8_cyc_o_reg/NET0131 ,
		\m2_stb_i_pad ,
		_w9619_
	);
	LUT4 #(
		.INIT('h0100)
	) name7719 (
		\m2_addr_i[28]_pad ,
		\m2_addr_i[29]_pad ,
		\m2_addr_i[30]_pad ,
		\m2_addr_i[31]_pad ,
		_w9620_
	);
	LUT3 #(
		.INIT('hec)
	) name7720 (
		_w9285_,
		_w9619_,
		_w9620_,
		_w9621_
	);
	LUT3 #(
		.INIT('h08)
	) name7721 (
		\m7_cyc_i_pad ,
		\m7_s8_cyc_o_reg/NET0131 ,
		\m7_stb_i_pad ,
		_w9622_
	);
	LUT4 #(
		.INIT('h0100)
	) name7722 (
		\m7_addr_i[28]_pad ,
		\m7_addr_i[29]_pad ,
		\m7_addr_i[30]_pad ,
		\m7_addr_i[31]_pad ,
		_w9623_
	);
	LUT3 #(
		.INIT('hec)
	) name7723 (
		_w9316_,
		_w9622_,
		_w9623_,
		_w9624_
	);
	LUT3 #(
		.INIT('h08)
	) name7724 (
		\m2_cyc_i_pad ,
		\m2_s7_cyc_o_reg/NET0131 ,
		\m2_stb_i_pad ,
		_w9625_
	);
	LUT4 #(
		.INIT('h0080)
	) name7725 (
		\m2_addr_i[28]_pad ,
		\m2_addr_i[29]_pad ,
		\m2_addr_i[30]_pad ,
		\m2_addr_i[31]_pad ,
		_w9626_
	);
	LUT3 #(
		.INIT('hec)
	) name7726 (
		_w9285_,
		_w9625_,
		_w9626_,
		_w9627_
	);
	LUT3 #(
		.INIT('h08)
	) name7727 (
		\m2_cyc_i_pad ,
		\m2_s13_cyc_o_reg/NET0131 ,
		\m2_stb_i_pad ,
		_w9628_
	);
	LUT4 #(
		.INIT('h2000)
	) name7728 (
		\m2_addr_i[28]_pad ,
		\m2_addr_i[29]_pad ,
		\m2_addr_i[30]_pad ,
		\m2_addr_i[31]_pad ,
		_w9629_
	);
	LUT3 #(
		.INIT('hec)
	) name7729 (
		_w9285_,
		_w9628_,
		_w9629_,
		_w9630_
	);
	LUT3 #(
		.INIT('h08)
	) name7730 (
		\m2_cyc_i_pad ,
		\m2_s14_cyc_o_reg/NET0131 ,
		\m2_stb_i_pad ,
		_w9631_
	);
	LUT4 #(
		.INIT('h4000)
	) name7731 (
		\m2_addr_i[28]_pad ,
		\m2_addr_i[29]_pad ,
		\m2_addr_i[30]_pad ,
		\m2_addr_i[31]_pad ,
		_w9632_
	);
	LUT3 #(
		.INIT('hec)
	) name7732 (
		_w9285_,
		_w9631_,
		_w9632_,
		_w9633_
	);
	LUT3 #(
		.INIT('h08)
	) name7733 (
		\m1_cyc_i_pad ,
		\m1_s12_cyc_o_reg/NET0131 ,
		\m1_stb_i_pad ,
		_w9634_
	);
	LUT4 #(
		.INIT('h1000)
	) name7734 (
		\m1_addr_i[28]_pad ,
		\m1_addr_i[29]_pad ,
		\m1_addr_i[30]_pad ,
		\m1_addr_i[31]_pad ,
		_w9635_
	);
	LUT3 #(
		.INIT('hec)
	) name7735 (
		_w9281_,
		_w9634_,
		_w9635_,
		_w9636_
	);
	LUT3 #(
		.INIT('h08)
	) name7736 (
		\m1_cyc_i_pad ,
		\m1_s11_cyc_o_reg/NET0131 ,
		\m1_stb_i_pad ,
		_w9637_
	);
	LUT4 #(
		.INIT('h0800)
	) name7737 (
		\m1_addr_i[28]_pad ,
		\m1_addr_i[29]_pad ,
		\m1_addr_i[30]_pad ,
		\m1_addr_i[31]_pad ,
		_w9638_
	);
	LUT3 #(
		.INIT('hec)
	) name7738 (
		_w9281_,
		_w9637_,
		_w9638_,
		_w9639_
	);
	LUT3 #(
		.INIT('h08)
	) name7739 (
		\m0_cyc_i_pad ,
		\m0_s9_cyc_o_reg/NET0131 ,
		\m0_stb_i_pad ,
		_w9640_
	);
	LUT4 #(
		.INIT('h0200)
	) name7740 (
		\m0_addr_i[28]_pad ,
		\m0_addr_i[29]_pad ,
		\m0_addr_i[30]_pad ,
		\m0_addr_i[31]_pad ,
		_w9641_
	);
	LUT3 #(
		.INIT('hec)
	) name7741 (
		_w9274_,
		_w9640_,
		_w9641_,
		_w9642_
	);
	LUT3 #(
		.INIT('h08)
	) name7742 (
		\m0_cyc_i_pad ,
		\m0_s4_cyc_o_reg/NET0131 ,
		\m0_stb_i_pad ,
		_w9643_
	);
	LUT4 #(
		.INIT('h0010)
	) name7743 (
		\m0_addr_i[28]_pad ,
		\m0_addr_i[29]_pad ,
		\m0_addr_i[30]_pad ,
		\m0_addr_i[31]_pad ,
		_w9644_
	);
	LUT3 #(
		.INIT('hec)
	) name7744 (
		_w9274_,
		_w9643_,
		_w9644_,
		_w9645_
	);
	LUT3 #(
		.INIT('h08)
	) name7745 (
		\m0_cyc_i_pad ,
		\m0_s13_cyc_o_reg/NET0131 ,
		\m0_stb_i_pad ,
		_w9646_
	);
	LUT4 #(
		.INIT('h2000)
	) name7746 (
		\m0_addr_i[28]_pad ,
		\m0_addr_i[29]_pad ,
		\m0_addr_i[30]_pad ,
		\m0_addr_i[31]_pad ,
		_w9647_
	);
	LUT3 #(
		.INIT('hec)
	) name7747 (
		_w9274_,
		_w9646_,
		_w9647_,
		_w9648_
	);
	LUT3 #(
		.INIT('h08)
	) name7748 (
		\m0_cyc_i_pad ,
		\m0_s12_cyc_o_reg/NET0131 ,
		\m0_stb_i_pad ,
		_w9649_
	);
	LUT4 #(
		.INIT('h1000)
	) name7749 (
		\m0_addr_i[28]_pad ,
		\m0_addr_i[29]_pad ,
		\m0_addr_i[30]_pad ,
		\m0_addr_i[31]_pad ,
		_w9650_
	);
	LUT3 #(
		.INIT('hec)
	) name7750 (
		_w9274_,
		_w9649_,
		_w9650_,
		_w9651_
	);
	LUT3 #(
		.INIT('h15)
	) name7751 (
		\s15_ack_i_pad ,
		_w2046_,
		_w2097_,
		_w9652_
	);
	LUT3 #(
		.INIT('h80)
	) name7752 (
		_w1908_,
		_w1909_,
		_w2049_,
		_w9653_
	);
	LUT2 #(
		.INIT('h8)
	) name7753 (
		_w1914_,
		_w9653_,
		_w9654_
	);
	LUT3 #(
		.INIT('h70)
	) name7754 (
		_w2097_,
		_w8630_,
		_w9654_,
		_w9655_
	);
	LUT4 #(
		.INIT('h8000)
	) name7755 (
		\s14_ack_i_pad ,
		_w9137_,
		_w9138_,
		_w9390_,
		_w9656_
	);
	LUT4 #(
		.INIT('h8000)
	) name7756 (
		\s3_ack_i_pad ,
		_w9205_,
		_w9206_,
		_w9398_,
		_w9657_
	);
	LUT4 #(
		.INIT('h135f)
	) name7757 (
		_w9136_,
		_w9224_,
		_w9656_,
		_w9657_,
		_w9658_
	);
	LUT4 #(
		.INIT('h8000)
	) name7758 (
		\s1_ack_i_pad ,
		_w9103_,
		_w9104_,
		_w9277_,
		_w9659_
	);
	LUT4 #(
		.INIT('h8000)
	) name7759 (
		\s4_ack_i_pad ,
		_w8655_,
		_w8656_,
		_w9644_,
		_w9660_
	);
	LUT4 #(
		.INIT('h153f)
	) name7760 (
		_w8662_,
		_w9122_,
		_w9659_,
		_w9660_,
		_w9661_
	);
	LUT4 #(
		.INIT('h8000)
	) name7761 (
		\s10_ack_i_pad ,
		_w8910_,
		_w8911_,
		_w9381_,
		_w9662_
	);
	LUT4 #(
		.INIT('h8000)
	) name7762 (
		\s2_ack_i_pad ,
		_w9171_,
		_w9172_,
		_w9395_,
		_w9663_
	);
	LUT4 #(
		.INIT('h135f)
	) name7763 (
		_w8923_,
		_w9178_,
		_w9662_,
		_w9663_,
		_w9664_
	);
	LUT4 #(
		.INIT('h8000)
	) name7764 (
		\s13_ack_i_pad ,
		_w9069_,
		_w9070_,
		_w9647_,
		_w9665_
	);
	LUT4 #(
		.INIT('h8000)
	) name7765 (
		\s0_ack_i_pad ,
		_w8989_,
		_w8990_,
		_w9273_,
		_w9666_
	);
	LUT4 #(
		.INIT('h153f)
	) name7766 (
		_w9008_,
		_w9076_,
		_w9665_,
		_w9666_,
		_w9667_
	);
	LUT4 #(
		.INIT('h8000)
	) name7767 (
		_w9658_,
		_w9661_,
		_w9664_,
		_w9667_,
		_w9668_
	);
	LUT4 #(
		.INIT('h8000)
	) name7768 (
		\s6_ack_i_pad ,
		_w8743_,
		_w8744_,
		_w9404_,
		_w9669_
	);
	LUT2 #(
		.INIT('h8)
	) name7769 (
		_w8742_,
		_w9669_,
		_w9670_
	);
	LUT4 #(
		.INIT('h8000)
	) name7770 (
		\s11_ack_i_pad ,
		_w8955_,
		_w8956_,
		_w9384_,
		_w9671_
	);
	LUT4 #(
		.INIT('h8000)
	) name7771 (
		\s9_ack_i_pad ,
		_w8865_,
		_w8866_,
		_w9641_,
		_w9672_
	);
	LUT4 #(
		.INIT('h153f)
	) name7772 (
		_w8872_,
		_w8962_,
		_w9671_,
		_w9672_,
		_w9673_
	);
	LUT4 #(
		.INIT('h8000)
	) name7773 (
		\s7_ack_i_pad ,
		_w8782_,
		_w8783_,
		_w9407_,
		_w9674_
	);
	LUT4 #(
		.INIT('h8000)
	) name7774 (
		\s12_ack_i_pad ,
		_w9029_,
		_w9030_,
		_w9650_,
		_w9675_
	);
	LUT4 #(
		.INIT('h135f)
	) name7775 (
		_w8789_,
		_w9048_,
		_w9674_,
		_w9675_,
		_w9676_
	);
	LUT4 #(
		.INIT('h8000)
	) name7776 (
		\s5_ack_i_pad ,
		_w8699_,
		_w8700_,
		_w9401_,
		_w9677_
	);
	LUT4 #(
		.INIT('h8000)
	) name7777 (
		\s8_ack_i_pad ,
		_w8821_,
		_w8822_,
		_w9410_,
		_w9678_
	);
	LUT4 #(
		.INIT('h135f)
	) name7778 (
		_w8718_,
		_w8820_,
		_w9677_,
		_w9678_,
		_w9679_
	);
	LUT4 #(
		.INIT('h4000)
	) name7779 (
		_w9670_,
		_w9673_,
		_w9676_,
		_w9679_,
		_w9680_
	);
	LUT2 #(
		.INIT('h8)
	) name7780 (
		_w9668_,
		_w9680_,
		_w9681_
	);
	LUT3 #(
		.INIT('h4f)
	) name7781 (
		_w9652_,
		_w9655_,
		_w9681_,
		_w9682_
	);
	LUT4 #(
		.INIT('h0002)
	) name7782 (
		\rf_rf_dout_reg[0]/P0001 ,
		_w2016_,
		_w2029_,
		_w2043_,
		_w9683_
	);
	LUT3 #(
		.INIT('h80)
	) name7783 (
		_w2049_,
		_w2097_,
		_w9683_,
		_w9684_
	);
	LUT2 #(
		.INIT('h8)
	) name7784 (
		\s15_data_i[0]_pad ,
		_w2049_,
		_w9685_
	);
	LUT3 #(
		.INIT('h70)
	) name7785 (
		_w2046_,
		_w2097_,
		_w9685_,
		_w9686_
	);
	LUT4 #(
		.INIT('h135f)
	) name7786 (
		\s1_data_i[0]_pad ,
		\s8_data_i[0]_pad ,
		_w9277_,
		_w9410_,
		_w9687_
	);
	LUT4 #(
		.INIT('h153f)
	) name7787 (
		\s4_data_i[0]_pad ,
		\s6_data_i[0]_pad ,
		_w9404_,
		_w9644_,
		_w9688_
	);
	LUT4 #(
		.INIT('h135f)
	) name7788 (
		\s5_data_i[0]_pad ,
		\s9_data_i[0]_pad ,
		_w9401_,
		_w9641_,
		_w9689_
	);
	LUT4 #(
		.INIT('h135f)
	) name7789 (
		\s10_data_i[0]_pad ,
		\s7_data_i[0]_pad ,
		_w9381_,
		_w9407_,
		_w9690_
	);
	LUT4 #(
		.INIT('h8000)
	) name7790 (
		_w9687_,
		_w9688_,
		_w9689_,
		_w9690_,
		_w9691_
	);
	LUT2 #(
		.INIT('h8)
	) name7791 (
		\s11_data_i[0]_pad ,
		_w9384_,
		_w9692_
	);
	LUT4 #(
		.INIT('h135f)
	) name7792 (
		\s14_data_i[0]_pad ,
		\s3_data_i[0]_pad ,
		_w9390_,
		_w9398_,
		_w9693_
	);
	LUT4 #(
		.INIT('h153f)
	) name7793 (
		\s12_data_i[0]_pad ,
		\s2_data_i[0]_pad ,
		_w9395_,
		_w9650_,
		_w9694_
	);
	LUT4 #(
		.INIT('h135f)
	) name7794 (
		\s0_data_i[0]_pad ,
		\s13_data_i[0]_pad ,
		_w9273_,
		_w9647_,
		_w9695_
	);
	LUT4 #(
		.INIT('h4000)
	) name7795 (
		_w9692_,
		_w9693_,
		_w9694_,
		_w9695_,
		_w9696_
	);
	LUT2 #(
		.INIT('h8)
	) name7796 (
		_w9691_,
		_w9696_,
		_w9697_
	);
	LUT3 #(
		.INIT('hef)
	) name7797 (
		_w9684_,
		_w9686_,
		_w9697_,
		_w9698_
	);
	LUT4 #(
		.INIT('h0002)
	) name7798 (
		\rf_rf_dout_reg[10]/P0001 ,
		_w2016_,
		_w2029_,
		_w2043_,
		_w9699_
	);
	LUT3 #(
		.INIT('h80)
	) name7799 (
		_w2049_,
		_w2097_,
		_w9699_,
		_w9700_
	);
	LUT2 #(
		.INIT('h8)
	) name7800 (
		\s15_data_i[10]_pad ,
		_w2049_,
		_w9701_
	);
	LUT3 #(
		.INIT('h70)
	) name7801 (
		_w2046_,
		_w2097_,
		_w9701_,
		_w9702_
	);
	LUT4 #(
		.INIT('h135f)
	) name7802 (
		\s1_data_i[10]_pad ,
		\s8_data_i[10]_pad ,
		_w9277_,
		_w9410_,
		_w9703_
	);
	LUT4 #(
		.INIT('h153f)
	) name7803 (
		\s4_data_i[10]_pad ,
		\s6_data_i[10]_pad ,
		_w9404_,
		_w9644_,
		_w9704_
	);
	LUT4 #(
		.INIT('h135f)
	) name7804 (
		\s5_data_i[10]_pad ,
		\s9_data_i[10]_pad ,
		_w9401_,
		_w9641_,
		_w9705_
	);
	LUT4 #(
		.INIT('h135f)
	) name7805 (
		\s10_data_i[10]_pad ,
		\s7_data_i[10]_pad ,
		_w9381_,
		_w9407_,
		_w9706_
	);
	LUT4 #(
		.INIT('h8000)
	) name7806 (
		_w9703_,
		_w9704_,
		_w9705_,
		_w9706_,
		_w9707_
	);
	LUT2 #(
		.INIT('h8)
	) name7807 (
		\s11_data_i[10]_pad ,
		_w9384_,
		_w9708_
	);
	LUT4 #(
		.INIT('h135f)
	) name7808 (
		\s14_data_i[10]_pad ,
		\s3_data_i[10]_pad ,
		_w9390_,
		_w9398_,
		_w9709_
	);
	LUT4 #(
		.INIT('h153f)
	) name7809 (
		\s12_data_i[10]_pad ,
		\s2_data_i[10]_pad ,
		_w9395_,
		_w9650_,
		_w9710_
	);
	LUT4 #(
		.INIT('h135f)
	) name7810 (
		\s0_data_i[10]_pad ,
		\s13_data_i[10]_pad ,
		_w9273_,
		_w9647_,
		_w9711_
	);
	LUT4 #(
		.INIT('h4000)
	) name7811 (
		_w9708_,
		_w9709_,
		_w9710_,
		_w9711_,
		_w9712_
	);
	LUT2 #(
		.INIT('h8)
	) name7812 (
		_w9707_,
		_w9712_,
		_w9713_
	);
	LUT3 #(
		.INIT('hef)
	) name7813 (
		_w9700_,
		_w9702_,
		_w9713_,
		_w9714_
	);
	LUT4 #(
		.INIT('h0002)
	) name7814 (
		\rf_rf_dout_reg[11]/P0001 ,
		_w2016_,
		_w2029_,
		_w2043_,
		_w9715_
	);
	LUT3 #(
		.INIT('h80)
	) name7815 (
		_w2049_,
		_w2097_,
		_w9715_,
		_w9716_
	);
	LUT2 #(
		.INIT('h8)
	) name7816 (
		\s15_data_i[11]_pad ,
		_w2049_,
		_w9717_
	);
	LUT3 #(
		.INIT('h70)
	) name7817 (
		_w2046_,
		_w2097_,
		_w9717_,
		_w9718_
	);
	LUT4 #(
		.INIT('h135f)
	) name7818 (
		\s1_data_i[11]_pad ,
		\s8_data_i[11]_pad ,
		_w9277_,
		_w9410_,
		_w9719_
	);
	LUT4 #(
		.INIT('h153f)
	) name7819 (
		\s4_data_i[11]_pad ,
		\s6_data_i[11]_pad ,
		_w9404_,
		_w9644_,
		_w9720_
	);
	LUT4 #(
		.INIT('h135f)
	) name7820 (
		\s5_data_i[11]_pad ,
		\s9_data_i[11]_pad ,
		_w9401_,
		_w9641_,
		_w9721_
	);
	LUT4 #(
		.INIT('h135f)
	) name7821 (
		\s10_data_i[11]_pad ,
		\s7_data_i[11]_pad ,
		_w9381_,
		_w9407_,
		_w9722_
	);
	LUT4 #(
		.INIT('h8000)
	) name7822 (
		_w9719_,
		_w9720_,
		_w9721_,
		_w9722_,
		_w9723_
	);
	LUT2 #(
		.INIT('h8)
	) name7823 (
		\s11_data_i[11]_pad ,
		_w9384_,
		_w9724_
	);
	LUT4 #(
		.INIT('h135f)
	) name7824 (
		\s14_data_i[11]_pad ,
		\s3_data_i[11]_pad ,
		_w9390_,
		_w9398_,
		_w9725_
	);
	LUT4 #(
		.INIT('h153f)
	) name7825 (
		\s12_data_i[11]_pad ,
		\s2_data_i[11]_pad ,
		_w9395_,
		_w9650_,
		_w9726_
	);
	LUT4 #(
		.INIT('h135f)
	) name7826 (
		\s0_data_i[11]_pad ,
		\s13_data_i[11]_pad ,
		_w9273_,
		_w9647_,
		_w9727_
	);
	LUT4 #(
		.INIT('h4000)
	) name7827 (
		_w9724_,
		_w9725_,
		_w9726_,
		_w9727_,
		_w9728_
	);
	LUT2 #(
		.INIT('h8)
	) name7828 (
		_w9723_,
		_w9728_,
		_w9729_
	);
	LUT3 #(
		.INIT('hef)
	) name7829 (
		_w9716_,
		_w9718_,
		_w9729_,
		_w9730_
	);
	LUT4 #(
		.INIT('h0002)
	) name7830 (
		\rf_rf_dout_reg[12]/P0001 ,
		_w2016_,
		_w2029_,
		_w2043_,
		_w9731_
	);
	LUT3 #(
		.INIT('h80)
	) name7831 (
		_w2049_,
		_w2097_,
		_w9731_,
		_w9732_
	);
	LUT2 #(
		.INIT('h8)
	) name7832 (
		\s15_data_i[12]_pad ,
		_w2049_,
		_w9733_
	);
	LUT3 #(
		.INIT('h70)
	) name7833 (
		_w2046_,
		_w2097_,
		_w9733_,
		_w9734_
	);
	LUT4 #(
		.INIT('h135f)
	) name7834 (
		\s1_data_i[12]_pad ,
		\s8_data_i[12]_pad ,
		_w9277_,
		_w9410_,
		_w9735_
	);
	LUT4 #(
		.INIT('h153f)
	) name7835 (
		\s4_data_i[12]_pad ,
		\s6_data_i[12]_pad ,
		_w9404_,
		_w9644_,
		_w9736_
	);
	LUT4 #(
		.INIT('h135f)
	) name7836 (
		\s5_data_i[12]_pad ,
		\s9_data_i[12]_pad ,
		_w9401_,
		_w9641_,
		_w9737_
	);
	LUT4 #(
		.INIT('h135f)
	) name7837 (
		\s10_data_i[12]_pad ,
		\s7_data_i[12]_pad ,
		_w9381_,
		_w9407_,
		_w9738_
	);
	LUT4 #(
		.INIT('h8000)
	) name7838 (
		_w9735_,
		_w9736_,
		_w9737_,
		_w9738_,
		_w9739_
	);
	LUT2 #(
		.INIT('h8)
	) name7839 (
		\s11_data_i[12]_pad ,
		_w9384_,
		_w9740_
	);
	LUT4 #(
		.INIT('h135f)
	) name7840 (
		\s14_data_i[12]_pad ,
		\s3_data_i[12]_pad ,
		_w9390_,
		_w9398_,
		_w9741_
	);
	LUT4 #(
		.INIT('h153f)
	) name7841 (
		\s12_data_i[12]_pad ,
		\s2_data_i[12]_pad ,
		_w9395_,
		_w9650_,
		_w9742_
	);
	LUT4 #(
		.INIT('h135f)
	) name7842 (
		\s0_data_i[12]_pad ,
		\s13_data_i[12]_pad ,
		_w9273_,
		_w9647_,
		_w9743_
	);
	LUT4 #(
		.INIT('h4000)
	) name7843 (
		_w9740_,
		_w9741_,
		_w9742_,
		_w9743_,
		_w9744_
	);
	LUT2 #(
		.INIT('h8)
	) name7844 (
		_w9739_,
		_w9744_,
		_w9745_
	);
	LUT3 #(
		.INIT('hef)
	) name7845 (
		_w9732_,
		_w9734_,
		_w9745_,
		_w9746_
	);
	LUT4 #(
		.INIT('h0002)
	) name7846 (
		\rf_rf_dout_reg[13]/P0001 ,
		_w2016_,
		_w2029_,
		_w2043_,
		_w9747_
	);
	LUT3 #(
		.INIT('h80)
	) name7847 (
		_w2049_,
		_w2097_,
		_w9747_,
		_w9748_
	);
	LUT2 #(
		.INIT('h8)
	) name7848 (
		\s15_data_i[13]_pad ,
		_w2049_,
		_w9749_
	);
	LUT3 #(
		.INIT('h70)
	) name7849 (
		_w2046_,
		_w2097_,
		_w9749_,
		_w9750_
	);
	LUT4 #(
		.INIT('h135f)
	) name7850 (
		\s1_data_i[13]_pad ,
		\s8_data_i[13]_pad ,
		_w9277_,
		_w9410_,
		_w9751_
	);
	LUT4 #(
		.INIT('h153f)
	) name7851 (
		\s4_data_i[13]_pad ,
		\s6_data_i[13]_pad ,
		_w9404_,
		_w9644_,
		_w9752_
	);
	LUT4 #(
		.INIT('h135f)
	) name7852 (
		\s5_data_i[13]_pad ,
		\s9_data_i[13]_pad ,
		_w9401_,
		_w9641_,
		_w9753_
	);
	LUT4 #(
		.INIT('h135f)
	) name7853 (
		\s10_data_i[13]_pad ,
		\s7_data_i[13]_pad ,
		_w9381_,
		_w9407_,
		_w9754_
	);
	LUT4 #(
		.INIT('h8000)
	) name7854 (
		_w9751_,
		_w9752_,
		_w9753_,
		_w9754_,
		_w9755_
	);
	LUT2 #(
		.INIT('h8)
	) name7855 (
		\s11_data_i[13]_pad ,
		_w9384_,
		_w9756_
	);
	LUT4 #(
		.INIT('h135f)
	) name7856 (
		\s14_data_i[13]_pad ,
		\s3_data_i[13]_pad ,
		_w9390_,
		_w9398_,
		_w9757_
	);
	LUT4 #(
		.INIT('h153f)
	) name7857 (
		\s12_data_i[13]_pad ,
		\s2_data_i[13]_pad ,
		_w9395_,
		_w9650_,
		_w9758_
	);
	LUT4 #(
		.INIT('h135f)
	) name7858 (
		\s0_data_i[13]_pad ,
		\s13_data_i[13]_pad ,
		_w9273_,
		_w9647_,
		_w9759_
	);
	LUT4 #(
		.INIT('h4000)
	) name7859 (
		_w9756_,
		_w9757_,
		_w9758_,
		_w9759_,
		_w9760_
	);
	LUT2 #(
		.INIT('h8)
	) name7860 (
		_w9755_,
		_w9760_,
		_w9761_
	);
	LUT3 #(
		.INIT('hef)
	) name7861 (
		_w9748_,
		_w9750_,
		_w9761_,
		_w9762_
	);
	LUT4 #(
		.INIT('h0002)
	) name7862 (
		\rf_rf_dout_reg[14]/P0001 ,
		_w2016_,
		_w2029_,
		_w2043_,
		_w9763_
	);
	LUT3 #(
		.INIT('h80)
	) name7863 (
		_w2049_,
		_w2097_,
		_w9763_,
		_w9764_
	);
	LUT2 #(
		.INIT('h8)
	) name7864 (
		\s15_data_i[14]_pad ,
		_w2049_,
		_w9765_
	);
	LUT3 #(
		.INIT('h70)
	) name7865 (
		_w2046_,
		_w2097_,
		_w9765_,
		_w9766_
	);
	LUT4 #(
		.INIT('h135f)
	) name7866 (
		\s1_data_i[14]_pad ,
		\s8_data_i[14]_pad ,
		_w9277_,
		_w9410_,
		_w9767_
	);
	LUT4 #(
		.INIT('h153f)
	) name7867 (
		\s4_data_i[14]_pad ,
		\s6_data_i[14]_pad ,
		_w9404_,
		_w9644_,
		_w9768_
	);
	LUT4 #(
		.INIT('h135f)
	) name7868 (
		\s5_data_i[14]_pad ,
		\s9_data_i[14]_pad ,
		_w9401_,
		_w9641_,
		_w9769_
	);
	LUT4 #(
		.INIT('h135f)
	) name7869 (
		\s10_data_i[14]_pad ,
		\s7_data_i[14]_pad ,
		_w9381_,
		_w9407_,
		_w9770_
	);
	LUT4 #(
		.INIT('h8000)
	) name7870 (
		_w9767_,
		_w9768_,
		_w9769_,
		_w9770_,
		_w9771_
	);
	LUT2 #(
		.INIT('h8)
	) name7871 (
		\s11_data_i[14]_pad ,
		_w9384_,
		_w9772_
	);
	LUT4 #(
		.INIT('h135f)
	) name7872 (
		\s14_data_i[14]_pad ,
		\s3_data_i[14]_pad ,
		_w9390_,
		_w9398_,
		_w9773_
	);
	LUT4 #(
		.INIT('h153f)
	) name7873 (
		\s12_data_i[14]_pad ,
		\s2_data_i[14]_pad ,
		_w9395_,
		_w9650_,
		_w9774_
	);
	LUT4 #(
		.INIT('h135f)
	) name7874 (
		\s0_data_i[14]_pad ,
		\s13_data_i[14]_pad ,
		_w9273_,
		_w9647_,
		_w9775_
	);
	LUT4 #(
		.INIT('h4000)
	) name7875 (
		_w9772_,
		_w9773_,
		_w9774_,
		_w9775_,
		_w9776_
	);
	LUT2 #(
		.INIT('h8)
	) name7876 (
		_w9771_,
		_w9776_,
		_w9777_
	);
	LUT3 #(
		.INIT('hef)
	) name7877 (
		_w9764_,
		_w9766_,
		_w9777_,
		_w9778_
	);
	LUT4 #(
		.INIT('h0002)
	) name7878 (
		\rf_rf_dout_reg[15]/P0001 ,
		_w2016_,
		_w2029_,
		_w2043_,
		_w9779_
	);
	LUT3 #(
		.INIT('h80)
	) name7879 (
		_w2049_,
		_w2097_,
		_w9779_,
		_w9780_
	);
	LUT2 #(
		.INIT('h8)
	) name7880 (
		\s15_data_i[15]_pad ,
		_w2049_,
		_w9781_
	);
	LUT3 #(
		.INIT('h70)
	) name7881 (
		_w2046_,
		_w2097_,
		_w9781_,
		_w9782_
	);
	LUT4 #(
		.INIT('h135f)
	) name7882 (
		\s1_data_i[15]_pad ,
		\s8_data_i[15]_pad ,
		_w9277_,
		_w9410_,
		_w9783_
	);
	LUT4 #(
		.INIT('h153f)
	) name7883 (
		\s4_data_i[15]_pad ,
		\s6_data_i[15]_pad ,
		_w9404_,
		_w9644_,
		_w9784_
	);
	LUT4 #(
		.INIT('h135f)
	) name7884 (
		\s5_data_i[15]_pad ,
		\s9_data_i[15]_pad ,
		_w9401_,
		_w9641_,
		_w9785_
	);
	LUT4 #(
		.INIT('h135f)
	) name7885 (
		\s10_data_i[15]_pad ,
		\s7_data_i[15]_pad ,
		_w9381_,
		_w9407_,
		_w9786_
	);
	LUT4 #(
		.INIT('h8000)
	) name7886 (
		_w9783_,
		_w9784_,
		_w9785_,
		_w9786_,
		_w9787_
	);
	LUT2 #(
		.INIT('h8)
	) name7887 (
		\s11_data_i[15]_pad ,
		_w9384_,
		_w9788_
	);
	LUT4 #(
		.INIT('h135f)
	) name7888 (
		\s14_data_i[15]_pad ,
		\s3_data_i[15]_pad ,
		_w9390_,
		_w9398_,
		_w9789_
	);
	LUT4 #(
		.INIT('h153f)
	) name7889 (
		\s12_data_i[15]_pad ,
		\s2_data_i[15]_pad ,
		_w9395_,
		_w9650_,
		_w9790_
	);
	LUT4 #(
		.INIT('h135f)
	) name7890 (
		\s0_data_i[15]_pad ,
		\s13_data_i[15]_pad ,
		_w9273_,
		_w9647_,
		_w9791_
	);
	LUT4 #(
		.INIT('h4000)
	) name7891 (
		_w9788_,
		_w9789_,
		_w9790_,
		_w9791_,
		_w9792_
	);
	LUT2 #(
		.INIT('h8)
	) name7892 (
		_w9787_,
		_w9792_,
		_w9793_
	);
	LUT3 #(
		.INIT('hef)
	) name7893 (
		_w9780_,
		_w9782_,
		_w9793_,
		_w9794_
	);
	LUT2 #(
		.INIT('h8)
	) name7894 (
		\s15_data_i[16]_pad ,
		_w2049_,
		_w9795_
	);
	LUT4 #(
		.INIT('h135f)
	) name7895 (
		\s1_data_i[16]_pad ,
		\s8_data_i[16]_pad ,
		_w9277_,
		_w9410_,
		_w9796_
	);
	LUT4 #(
		.INIT('h153f)
	) name7896 (
		\s4_data_i[16]_pad ,
		\s6_data_i[16]_pad ,
		_w9404_,
		_w9644_,
		_w9797_
	);
	LUT4 #(
		.INIT('h135f)
	) name7897 (
		\s5_data_i[16]_pad ,
		\s9_data_i[16]_pad ,
		_w9401_,
		_w9641_,
		_w9798_
	);
	LUT4 #(
		.INIT('h135f)
	) name7898 (
		\s10_data_i[16]_pad ,
		\s7_data_i[16]_pad ,
		_w9381_,
		_w9407_,
		_w9799_
	);
	LUT4 #(
		.INIT('h8000)
	) name7899 (
		_w9796_,
		_w9797_,
		_w9798_,
		_w9799_,
		_w9800_
	);
	LUT2 #(
		.INIT('h8)
	) name7900 (
		\s11_data_i[16]_pad ,
		_w9384_,
		_w9801_
	);
	LUT4 #(
		.INIT('h135f)
	) name7901 (
		\s14_data_i[16]_pad ,
		\s3_data_i[16]_pad ,
		_w9390_,
		_w9398_,
		_w9802_
	);
	LUT4 #(
		.INIT('h153f)
	) name7902 (
		\s12_data_i[16]_pad ,
		\s2_data_i[16]_pad ,
		_w9395_,
		_w9650_,
		_w9803_
	);
	LUT4 #(
		.INIT('h135f)
	) name7903 (
		\s0_data_i[16]_pad ,
		\s13_data_i[16]_pad ,
		_w9273_,
		_w9647_,
		_w9804_
	);
	LUT4 #(
		.INIT('h4000)
	) name7904 (
		_w9801_,
		_w9802_,
		_w9803_,
		_w9804_,
		_w9805_
	);
	LUT2 #(
		.INIT('h8)
	) name7905 (
		_w9800_,
		_w9805_,
		_w9806_
	);
	LUT4 #(
		.INIT('h70ff)
	) name7906 (
		_w2046_,
		_w2097_,
		_w9795_,
		_w9806_,
		_w9807_
	);
	LUT2 #(
		.INIT('h8)
	) name7907 (
		\s15_data_i[17]_pad ,
		_w2049_,
		_w9808_
	);
	LUT4 #(
		.INIT('h135f)
	) name7908 (
		\s1_data_i[17]_pad ,
		\s8_data_i[17]_pad ,
		_w9277_,
		_w9410_,
		_w9809_
	);
	LUT4 #(
		.INIT('h153f)
	) name7909 (
		\s4_data_i[17]_pad ,
		\s6_data_i[17]_pad ,
		_w9404_,
		_w9644_,
		_w9810_
	);
	LUT4 #(
		.INIT('h135f)
	) name7910 (
		\s5_data_i[17]_pad ,
		\s9_data_i[17]_pad ,
		_w9401_,
		_w9641_,
		_w9811_
	);
	LUT4 #(
		.INIT('h135f)
	) name7911 (
		\s10_data_i[17]_pad ,
		\s7_data_i[17]_pad ,
		_w9381_,
		_w9407_,
		_w9812_
	);
	LUT4 #(
		.INIT('h8000)
	) name7912 (
		_w9809_,
		_w9810_,
		_w9811_,
		_w9812_,
		_w9813_
	);
	LUT2 #(
		.INIT('h8)
	) name7913 (
		\s11_data_i[17]_pad ,
		_w9384_,
		_w9814_
	);
	LUT4 #(
		.INIT('h135f)
	) name7914 (
		\s14_data_i[17]_pad ,
		\s3_data_i[17]_pad ,
		_w9390_,
		_w9398_,
		_w9815_
	);
	LUT4 #(
		.INIT('h153f)
	) name7915 (
		\s12_data_i[17]_pad ,
		\s2_data_i[17]_pad ,
		_w9395_,
		_w9650_,
		_w9816_
	);
	LUT4 #(
		.INIT('h135f)
	) name7916 (
		\s0_data_i[17]_pad ,
		\s13_data_i[17]_pad ,
		_w9273_,
		_w9647_,
		_w9817_
	);
	LUT4 #(
		.INIT('h4000)
	) name7917 (
		_w9814_,
		_w9815_,
		_w9816_,
		_w9817_,
		_w9818_
	);
	LUT2 #(
		.INIT('h8)
	) name7918 (
		_w9813_,
		_w9818_,
		_w9819_
	);
	LUT4 #(
		.INIT('h70ff)
	) name7919 (
		_w2046_,
		_w2097_,
		_w9808_,
		_w9819_,
		_w9820_
	);
	LUT2 #(
		.INIT('h8)
	) name7920 (
		\s15_data_i[18]_pad ,
		_w2049_,
		_w9821_
	);
	LUT4 #(
		.INIT('h135f)
	) name7921 (
		\s1_data_i[18]_pad ,
		\s8_data_i[18]_pad ,
		_w9277_,
		_w9410_,
		_w9822_
	);
	LUT4 #(
		.INIT('h153f)
	) name7922 (
		\s4_data_i[18]_pad ,
		\s6_data_i[18]_pad ,
		_w9404_,
		_w9644_,
		_w9823_
	);
	LUT4 #(
		.INIT('h135f)
	) name7923 (
		\s5_data_i[18]_pad ,
		\s9_data_i[18]_pad ,
		_w9401_,
		_w9641_,
		_w9824_
	);
	LUT4 #(
		.INIT('h135f)
	) name7924 (
		\s10_data_i[18]_pad ,
		\s7_data_i[18]_pad ,
		_w9381_,
		_w9407_,
		_w9825_
	);
	LUT4 #(
		.INIT('h8000)
	) name7925 (
		_w9822_,
		_w9823_,
		_w9824_,
		_w9825_,
		_w9826_
	);
	LUT2 #(
		.INIT('h8)
	) name7926 (
		\s11_data_i[18]_pad ,
		_w9384_,
		_w9827_
	);
	LUT4 #(
		.INIT('h135f)
	) name7927 (
		\s14_data_i[18]_pad ,
		\s3_data_i[18]_pad ,
		_w9390_,
		_w9398_,
		_w9828_
	);
	LUT4 #(
		.INIT('h153f)
	) name7928 (
		\s12_data_i[18]_pad ,
		\s2_data_i[18]_pad ,
		_w9395_,
		_w9650_,
		_w9829_
	);
	LUT4 #(
		.INIT('h135f)
	) name7929 (
		\s0_data_i[18]_pad ,
		\s13_data_i[18]_pad ,
		_w9273_,
		_w9647_,
		_w9830_
	);
	LUT4 #(
		.INIT('h4000)
	) name7930 (
		_w9827_,
		_w9828_,
		_w9829_,
		_w9830_,
		_w9831_
	);
	LUT2 #(
		.INIT('h8)
	) name7931 (
		_w9826_,
		_w9831_,
		_w9832_
	);
	LUT4 #(
		.INIT('h70ff)
	) name7932 (
		_w2046_,
		_w2097_,
		_w9821_,
		_w9832_,
		_w9833_
	);
	LUT2 #(
		.INIT('h8)
	) name7933 (
		\s15_data_i[19]_pad ,
		_w2049_,
		_w9834_
	);
	LUT4 #(
		.INIT('h135f)
	) name7934 (
		\s1_data_i[19]_pad ,
		\s8_data_i[19]_pad ,
		_w9277_,
		_w9410_,
		_w9835_
	);
	LUT4 #(
		.INIT('h153f)
	) name7935 (
		\s4_data_i[19]_pad ,
		\s6_data_i[19]_pad ,
		_w9404_,
		_w9644_,
		_w9836_
	);
	LUT4 #(
		.INIT('h135f)
	) name7936 (
		\s5_data_i[19]_pad ,
		\s9_data_i[19]_pad ,
		_w9401_,
		_w9641_,
		_w9837_
	);
	LUT4 #(
		.INIT('h135f)
	) name7937 (
		\s10_data_i[19]_pad ,
		\s7_data_i[19]_pad ,
		_w9381_,
		_w9407_,
		_w9838_
	);
	LUT4 #(
		.INIT('h8000)
	) name7938 (
		_w9835_,
		_w9836_,
		_w9837_,
		_w9838_,
		_w9839_
	);
	LUT2 #(
		.INIT('h8)
	) name7939 (
		\s11_data_i[19]_pad ,
		_w9384_,
		_w9840_
	);
	LUT4 #(
		.INIT('h135f)
	) name7940 (
		\s14_data_i[19]_pad ,
		\s3_data_i[19]_pad ,
		_w9390_,
		_w9398_,
		_w9841_
	);
	LUT4 #(
		.INIT('h153f)
	) name7941 (
		\s12_data_i[19]_pad ,
		\s2_data_i[19]_pad ,
		_w9395_,
		_w9650_,
		_w9842_
	);
	LUT4 #(
		.INIT('h135f)
	) name7942 (
		\s0_data_i[19]_pad ,
		\s13_data_i[19]_pad ,
		_w9273_,
		_w9647_,
		_w9843_
	);
	LUT4 #(
		.INIT('h4000)
	) name7943 (
		_w9840_,
		_w9841_,
		_w9842_,
		_w9843_,
		_w9844_
	);
	LUT2 #(
		.INIT('h8)
	) name7944 (
		_w9839_,
		_w9844_,
		_w9845_
	);
	LUT4 #(
		.INIT('h70ff)
	) name7945 (
		_w2046_,
		_w2097_,
		_w9834_,
		_w9845_,
		_w9846_
	);
	LUT4 #(
		.INIT('h0002)
	) name7946 (
		\rf_rf_dout_reg[1]/P0001 ,
		_w2016_,
		_w2029_,
		_w2043_,
		_w9847_
	);
	LUT3 #(
		.INIT('h80)
	) name7947 (
		_w2049_,
		_w2097_,
		_w9847_,
		_w9848_
	);
	LUT2 #(
		.INIT('h8)
	) name7948 (
		\s15_data_i[1]_pad ,
		_w2049_,
		_w9849_
	);
	LUT3 #(
		.INIT('h70)
	) name7949 (
		_w2046_,
		_w2097_,
		_w9849_,
		_w9850_
	);
	LUT4 #(
		.INIT('h135f)
	) name7950 (
		\s1_data_i[1]_pad ,
		\s8_data_i[1]_pad ,
		_w9277_,
		_w9410_,
		_w9851_
	);
	LUT4 #(
		.INIT('h153f)
	) name7951 (
		\s4_data_i[1]_pad ,
		\s6_data_i[1]_pad ,
		_w9404_,
		_w9644_,
		_w9852_
	);
	LUT4 #(
		.INIT('h135f)
	) name7952 (
		\s5_data_i[1]_pad ,
		\s9_data_i[1]_pad ,
		_w9401_,
		_w9641_,
		_w9853_
	);
	LUT4 #(
		.INIT('h135f)
	) name7953 (
		\s10_data_i[1]_pad ,
		\s7_data_i[1]_pad ,
		_w9381_,
		_w9407_,
		_w9854_
	);
	LUT4 #(
		.INIT('h8000)
	) name7954 (
		_w9851_,
		_w9852_,
		_w9853_,
		_w9854_,
		_w9855_
	);
	LUT2 #(
		.INIT('h8)
	) name7955 (
		\s11_data_i[1]_pad ,
		_w9384_,
		_w9856_
	);
	LUT4 #(
		.INIT('h135f)
	) name7956 (
		\s14_data_i[1]_pad ,
		\s3_data_i[1]_pad ,
		_w9390_,
		_w9398_,
		_w9857_
	);
	LUT4 #(
		.INIT('h153f)
	) name7957 (
		\s12_data_i[1]_pad ,
		\s2_data_i[1]_pad ,
		_w9395_,
		_w9650_,
		_w9858_
	);
	LUT4 #(
		.INIT('h135f)
	) name7958 (
		\s0_data_i[1]_pad ,
		\s13_data_i[1]_pad ,
		_w9273_,
		_w9647_,
		_w9859_
	);
	LUT4 #(
		.INIT('h4000)
	) name7959 (
		_w9856_,
		_w9857_,
		_w9858_,
		_w9859_,
		_w9860_
	);
	LUT2 #(
		.INIT('h8)
	) name7960 (
		_w9855_,
		_w9860_,
		_w9861_
	);
	LUT3 #(
		.INIT('hef)
	) name7961 (
		_w9848_,
		_w9850_,
		_w9861_,
		_w9862_
	);
	LUT2 #(
		.INIT('h8)
	) name7962 (
		\s15_data_i[20]_pad ,
		_w2049_,
		_w9863_
	);
	LUT4 #(
		.INIT('h135f)
	) name7963 (
		\s1_data_i[20]_pad ,
		\s8_data_i[20]_pad ,
		_w9277_,
		_w9410_,
		_w9864_
	);
	LUT4 #(
		.INIT('h153f)
	) name7964 (
		\s4_data_i[20]_pad ,
		\s6_data_i[20]_pad ,
		_w9404_,
		_w9644_,
		_w9865_
	);
	LUT4 #(
		.INIT('h135f)
	) name7965 (
		\s5_data_i[20]_pad ,
		\s9_data_i[20]_pad ,
		_w9401_,
		_w9641_,
		_w9866_
	);
	LUT4 #(
		.INIT('h135f)
	) name7966 (
		\s10_data_i[20]_pad ,
		\s7_data_i[20]_pad ,
		_w9381_,
		_w9407_,
		_w9867_
	);
	LUT4 #(
		.INIT('h8000)
	) name7967 (
		_w9864_,
		_w9865_,
		_w9866_,
		_w9867_,
		_w9868_
	);
	LUT2 #(
		.INIT('h8)
	) name7968 (
		\s11_data_i[20]_pad ,
		_w9384_,
		_w9869_
	);
	LUT4 #(
		.INIT('h135f)
	) name7969 (
		\s14_data_i[20]_pad ,
		\s3_data_i[20]_pad ,
		_w9390_,
		_w9398_,
		_w9870_
	);
	LUT4 #(
		.INIT('h153f)
	) name7970 (
		\s12_data_i[20]_pad ,
		\s2_data_i[20]_pad ,
		_w9395_,
		_w9650_,
		_w9871_
	);
	LUT4 #(
		.INIT('h135f)
	) name7971 (
		\s0_data_i[20]_pad ,
		\s13_data_i[20]_pad ,
		_w9273_,
		_w9647_,
		_w9872_
	);
	LUT4 #(
		.INIT('h4000)
	) name7972 (
		_w9869_,
		_w9870_,
		_w9871_,
		_w9872_,
		_w9873_
	);
	LUT2 #(
		.INIT('h8)
	) name7973 (
		_w9868_,
		_w9873_,
		_w9874_
	);
	LUT4 #(
		.INIT('h70ff)
	) name7974 (
		_w2046_,
		_w2097_,
		_w9863_,
		_w9874_,
		_w9875_
	);
	LUT2 #(
		.INIT('h8)
	) name7975 (
		\s15_data_i[21]_pad ,
		_w2049_,
		_w9876_
	);
	LUT4 #(
		.INIT('h135f)
	) name7976 (
		\s1_data_i[21]_pad ,
		\s8_data_i[21]_pad ,
		_w9277_,
		_w9410_,
		_w9877_
	);
	LUT4 #(
		.INIT('h153f)
	) name7977 (
		\s4_data_i[21]_pad ,
		\s6_data_i[21]_pad ,
		_w9404_,
		_w9644_,
		_w9878_
	);
	LUT4 #(
		.INIT('h135f)
	) name7978 (
		\s5_data_i[21]_pad ,
		\s9_data_i[21]_pad ,
		_w9401_,
		_w9641_,
		_w9879_
	);
	LUT4 #(
		.INIT('h135f)
	) name7979 (
		\s10_data_i[21]_pad ,
		\s7_data_i[21]_pad ,
		_w9381_,
		_w9407_,
		_w9880_
	);
	LUT4 #(
		.INIT('h8000)
	) name7980 (
		_w9877_,
		_w9878_,
		_w9879_,
		_w9880_,
		_w9881_
	);
	LUT2 #(
		.INIT('h8)
	) name7981 (
		\s11_data_i[21]_pad ,
		_w9384_,
		_w9882_
	);
	LUT4 #(
		.INIT('h135f)
	) name7982 (
		\s14_data_i[21]_pad ,
		\s3_data_i[21]_pad ,
		_w9390_,
		_w9398_,
		_w9883_
	);
	LUT4 #(
		.INIT('h153f)
	) name7983 (
		\s12_data_i[21]_pad ,
		\s2_data_i[21]_pad ,
		_w9395_,
		_w9650_,
		_w9884_
	);
	LUT4 #(
		.INIT('h135f)
	) name7984 (
		\s0_data_i[21]_pad ,
		\s13_data_i[21]_pad ,
		_w9273_,
		_w9647_,
		_w9885_
	);
	LUT4 #(
		.INIT('h4000)
	) name7985 (
		_w9882_,
		_w9883_,
		_w9884_,
		_w9885_,
		_w9886_
	);
	LUT2 #(
		.INIT('h8)
	) name7986 (
		_w9881_,
		_w9886_,
		_w9887_
	);
	LUT4 #(
		.INIT('h70ff)
	) name7987 (
		_w2046_,
		_w2097_,
		_w9876_,
		_w9887_,
		_w9888_
	);
	LUT2 #(
		.INIT('h8)
	) name7988 (
		\s15_data_i[22]_pad ,
		_w2049_,
		_w9889_
	);
	LUT4 #(
		.INIT('h135f)
	) name7989 (
		\s1_data_i[22]_pad ,
		\s8_data_i[22]_pad ,
		_w9277_,
		_w9410_,
		_w9890_
	);
	LUT4 #(
		.INIT('h153f)
	) name7990 (
		\s4_data_i[22]_pad ,
		\s6_data_i[22]_pad ,
		_w9404_,
		_w9644_,
		_w9891_
	);
	LUT4 #(
		.INIT('h135f)
	) name7991 (
		\s5_data_i[22]_pad ,
		\s9_data_i[22]_pad ,
		_w9401_,
		_w9641_,
		_w9892_
	);
	LUT4 #(
		.INIT('h135f)
	) name7992 (
		\s10_data_i[22]_pad ,
		\s7_data_i[22]_pad ,
		_w9381_,
		_w9407_,
		_w9893_
	);
	LUT4 #(
		.INIT('h8000)
	) name7993 (
		_w9890_,
		_w9891_,
		_w9892_,
		_w9893_,
		_w9894_
	);
	LUT2 #(
		.INIT('h8)
	) name7994 (
		\s11_data_i[22]_pad ,
		_w9384_,
		_w9895_
	);
	LUT4 #(
		.INIT('h135f)
	) name7995 (
		\s14_data_i[22]_pad ,
		\s3_data_i[22]_pad ,
		_w9390_,
		_w9398_,
		_w9896_
	);
	LUT4 #(
		.INIT('h153f)
	) name7996 (
		\s12_data_i[22]_pad ,
		\s2_data_i[22]_pad ,
		_w9395_,
		_w9650_,
		_w9897_
	);
	LUT4 #(
		.INIT('h135f)
	) name7997 (
		\s0_data_i[22]_pad ,
		\s13_data_i[22]_pad ,
		_w9273_,
		_w9647_,
		_w9898_
	);
	LUT4 #(
		.INIT('h4000)
	) name7998 (
		_w9895_,
		_w9896_,
		_w9897_,
		_w9898_,
		_w9899_
	);
	LUT2 #(
		.INIT('h8)
	) name7999 (
		_w9894_,
		_w9899_,
		_w9900_
	);
	LUT4 #(
		.INIT('h70ff)
	) name8000 (
		_w2046_,
		_w2097_,
		_w9889_,
		_w9900_,
		_w9901_
	);
	LUT2 #(
		.INIT('h8)
	) name8001 (
		\s15_data_i[23]_pad ,
		_w2049_,
		_w9902_
	);
	LUT4 #(
		.INIT('h135f)
	) name8002 (
		\s1_data_i[23]_pad ,
		\s8_data_i[23]_pad ,
		_w9277_,
		_w9410_,
		_w9903_
	);
	LUT4 #(
		.INIT('h153f)
	) name8003 (
		\s4_data_i[23]_pad ,
		\s6_data_i[23]_pad ,
		_w9404_,
		_w9644_,
		_w9904_
	);
	LUT4 #(
		.INIT('h135f)
	) name8004 (
		\s5_data_i[23]_pad ,
		\s9_data_i[23]_pad ,
		_w9401_,
		_w9641_,
		_w9905_
	);
	LUT4 #(
		.INIT('h135f)
	) name8005 (
		\s10_data_i[23]_pad ,
		\s7_data_i[23]_pad ,
		_w9381_,
		_w9407_,
		_w9906_
	);
	LUT4 #(
		.INIT('h8000)
	) name8006 (
		_w9903_,
		_w9904_,
		_w9905_,
		_w9906_,
		_w9907_
	);
	LUT2 #(
		.INIT('h8)
	) name8007 (
		\s11_data_i[23]_pad ,
		_w9384_,
		_w9908_
	);
	LUT4 #(
		.INIT('h135f)
	) name8008 (
		\s14_data_i[23]_pad ,
		\s3_data_i[23]_pad ,
		_w9390_,
		_w9398_,
		_w9909_
	);
	LUT4 #(
		.INIT('h153f)
	) name8009 (
		\s12_data_i[23]_pad ,
		\s2_data_i[23]_pad ,
		_w9395_,
		_w9650_,
		_w9910_
	);
	LUT4 #(
		.INIT('h135f)
	) name8010 (
		\s0_data_i[23]_pad ,
		\s13_data_i[23]_pad ,
		_w9273_,
		_w9647_,
		_w9911_
	);
	LUT4 #(
		.INIT('h4000)
	) name8011 (
		_w9908_,
		_w9909_,
		_w9910_,
		_w9911_,
		_w9912_
	);
	LUT2 #(
		.INIT('h8)
	) name8012 (
		_w9907_,
		_w9912_,
		_w9913_
	);
	LUT4 #(
		.INIT('h70ff)
	) name8013 (
		_w2046_,
		_w2097_,
		_w9902_,
		_w9913_,
		_w9914_
	);
	LUT2 #(
		.INIT('h8)
	) name8014 (
		\s15_data_i[24]_pad ,
		_w2049_,
		_w9915_
	);
	LUT4 #(
		.INIT('h135f)
	) name8015 (
		\s1_data_i[24]_pad ,
		\s8_data_i[24]_pad ,
		_w9277_,
		_w9410_,
		_w9916_
	);
	LUT4 #(
		.INIT('h153f)
	) name8016 (
		\s4_data_i[24]_pad ,
		\s6_data_i[24]_pad ,
		_w9404_,
		_w9644_,
		_w9917_
	);
	LUT4 #(
		.INIT('h135f)
	) name8017 (
		\s5_data_i[24]_pad ,
		\s9_data_i[24]_pad ,
		_w9401_,
		_w9641_,
		_w9918_
	);
	LUT4 #(
		.INIT('h135f)
	) name8018 (
		\s10_data_i[24]_pad ,
		\s7_data_i[24]_pad ,
		_w9381_,
		_w9407_,
		_w9919_
	);
	LUT4 #(
		.INIT('h8000)
	) name8019 (
		_w9916_,
		_w9917_,
		_w9918_,
		_w9919_,
		_w9920_
	);
	LUT2 #(
		.INIT('h8)
	) name8020 (
		\s11_data_i[24]_pad ,
		_w9384_,
		_w9921_
	);
	LUT4 #(
		.INIT('h135f)
	) name8021 (
		\s14_data_i[24]_pad ,
		\s3_data_i[24]_pad ,
		_w9390_,
		_w9398_,
		_w9922_
	);
	LUT4 #(
		.INIT('h153f)
	) name8022 (
		\s12_data_i[24]_pad ,
		\s2_data_i[24]_pad ,
		_w9395_,
		_w9650_,
		_w9923_
	);
	LUT4 #(
		.INIT('h135f)
	) name8023 (
		\s0_data_i[24]_pad ,
		\s13_data_i[24]_pad ,
		_w9273_,
		_w9647_,
		_w9924_
	);
	LUT4 #(
		.INIT('h4000)
	) name8024 (
		_w9921_,
		_w9922_,
		_w9923_,
		_w9924_,
		_w9925_
	);
	LUT2 #(
		.INIT('h8)
	) name8025 (
		_w9920_,
		_w9925_,
		_w9926_
	);
	LUT4 #(
		.INIT('h70ff)
	) name8026 (
		_w2046_,
		_w2097_,
		_w9915_,
		_w9926_,
		_w9927_
	);
	LUT2 #(
		.INIT('h8)
	) name8027 (
		\s15_data_i[25]_pad ,
		_w2049_,
		_w9928_
	);
	LUT4 #(
		.INIT('h135f)
	) name8028 (
		\s1_data_i[25]_pad ,
		\s8_data_i[25]_pad ,
		_w9277_,
		_w9410_,
		_w9929_
	);
	LUT4 #(
		.INIT('h153f)
	) name8029 (
		\s4_data_i[25]_pad ,
		\s6_data_i[25]_pad ,
		_w9404_,
		_w9644_,
		_w9930_
	);
	LUT4 #(
		.INIT('h135f)
	) name8030 (
		\s5_data_i[25]_pad ,
		\s9_data_i[25]_pad ,
		_w9401_,
		_w9641_,
		_w9931_
	);
	LUT4 #(
		.INIT('h135f)
	) name8031 (
		\s10_data_i[25]_pad ,
		\s7_data_i[25]_pad ,
		_w9381_,
		_w9407_,
		_w9932_
	);
	LUT4 #(
		.INIT('h8000)
	) name8032 (
		_w9929_,
		_w9930_,
		_w9931_,
		_w9932_,
		_w9933_
	);
	LUT2 #(
		.INIT('h8)
	) name8033 (
		\s11_data_i[25]_pad ,
		_w9384_,
		_w9934_
	);
	LUT4 #(
		.INIT('h135f)
	) name8034 (
		\s14_data_i[25]_pad ,
		\s3_data_i[25]_pad ,
		_w9390_,
		_w9398_,
		_w9935_
	);
	LUT4 #(
		.INIT('h153f)
	) name8035 (
		\s12_data_i[25]_pad ,
		\s2_data_i[25]_pad ,
		_w9395_,
		_w9650_,
		_w9936_
	);
	LUT4 #(
		.INIT('h135f)
	) name8036 (
		\s0_data_i[25]_pad ,
		\s13_data_i[25]_pad ,
		_w9273_,
		_w9647_,
		_w9937_
	);
	LUT4 #(
		.INIT('h4000)
	) name8037 (
		_w9934_,
		_w9935_,
		_w9936_,
		_w9937_,
		_w9938_
	);
	LUT2 #(
		.INIT('h8)
	) name8038 (
		_w9933_,
		_w9938_,
		_w9939_
	);
	LUT4 #(
		.INIT('h70ff)
	) name8039 (
		_w2046_,
		_w2097_,
		_w9928_,
		_w9939_,
		_w9940_
	);
	LUT2 #(
		.INIT('h8)
	) name8040 (
		\s15_data_i[26]_pad ,
		_w2049_,
		_w9941_
	);
	LUT4 #(
		.INIT('h135f)
	) name8041 (
		\s1_data_i[26]_pad ,
		\s8_data_i[26]_pad ,
		_w9277_,
		_w9410_,
		_w9942_
	);
	LUT4 #(
		.INIT('h153f)
	) name8042 (
		\s4_data_i[26]_pad ,
		\s6_data_i[26]_pad ,
		_w9404_,
		_w9644_,
		_w9943_
	);
	LUT4 #(
		.INIT('h135f)
	) name8043 (
		\s5_data_i[26]_pad ,
		\s9_data_i[26]_pad ,
		_w9401_,
		_w9641_,
		_w9944_
	);
	LUT4 #(
		.INIT('h135f)
	) name8044 (
		\s10_data_i[26]_pad ,
		\s7_data_i[26]_pad ,
		_w9381_,
		_w9407_,
		_w9945_
	);
	LUT4 #(
		.INIT('h8000)
	) name8045 (
		_w9942_,
		_w9943_,
		_w9944_,
		_w9945_,
		_w9946_
	);
	LUT2 #(
		.INIT('h8)
	) name8046 (
		\s11_data_i[26]_pad ,
		_w9384_,
		_w9947_
	);
	LUT4 #(
		.INIT('h135f)
	) name8047 (
		\s14_data_i[26]_pad ,
		\s3_data_i[26]_pad ,
		_w9390_,
		_w9398_,
		_w9948_
	);
	LUT4 #(
		.INIT('h153f)
	) name8048 (
		\s12_data_i[26]_pad ,
		\s2_data_i[26]_pad ,
		_w9395_,
		_w9650_,
		_w9949_
	);
	LUT4 #(
		.INIT('h135f)
	) name8049 (
		\s0_data_i[26]_pad ,
		\s13_data_i[26]_pad ,
		_w9273_,
		_w9647_,
		_w9950_
	);
	LUT4 #(
		.INIT('h4000)
	) name8050 (
		_w9947_,
		_w9948_,
		_w9949_,
		_w9950_,
		_w9951_
	);
	LUT2 #(
		.INIT('h8)
	) name8051 (
		_w9946_,
		_w9951_,
		_w9952_
	);
	LUT4 #(
		.INIT('h70ff)
	) name8052 (
		_w2046_,
		_w2097_,
		_w9941_,
		_w9952_,
		_w9953_
	);
	LUT2 #(
		.INIT('h8)
	) name8053 (
		\s15_data_i[27]_pad ,
		_w2049_,
		_w9954_
	);
	LUT4 #(
		.INIT('h135f)
	) name8054 (
		\s1_data_i[27]_pad ,
		\s8_data_i[27]_pad ,
		_w9277_,
		_w9410_,
		_w9955_
	);
	LUT4 #(
		.INIT('h153f)
	) name8055 (
		\s4_data_i[27]_pad ,
		\s6_data_i[27]_pad ,
		_w9404_,
		_w9644_,
		_w9956_
	);
	LUT4 #(
		.INIT('h135f)
	) name8056 (
		\s5_data_i[27]_pad ,
		\s9_data_i[27]_pad ,
		_w9401_,
		_w9641_,
		_w9957_
	);
	LUT4 #(
		.INIT('h135f)
	) name8057 (
		\s10_data_i[27]_pad ,
		\s7_data_i[27]_pad ,
		_w9381_,
		_w9407_,
		_w9958_
	);
	LUT4 #(
		.INIT('h8000)
	) name8058 (
		_w9955_,
		_w9956_,
		_w9957_,
		_w9958_,
		_w9959_
	);
	LUT2 #(
		.INIT('h8)
	) name8059 (
		\s11_data_i[27]_pad ,
		_w9384_,
		_w9960_
	);
	LUT4 #(
		.INIT('h135f)
	) name8060 (
		\s14_data_i[27]_pad ,
		\s3_data_i[27]_pad ,
		_w9390_,
		_w9398_,
		_w9961_
	);
	LUT4 #(
		.INIT('h153f)
	) name8061 (
		\s12_data_i[27]_pad ,
		\s2_data_i[27]_pad ,
		_w9395_,
		_w9650_,
		_w9962_
	);
	LUT4 #(
		.INIT('h135f)
	) name8062 (
		\s0_data_i[27]_pad ,
		\s13_data_i[27]_pad ,
		_w9273_,
		_w9647_,
		_w9963_
	);
	LUT4 #(
		.INIT('h4000)
	) name8063 (
		_w9960_,
		_w9961_,
		_w9962_,
		_w9963_,
		_w9964_
	);
	LUT2 #(
		.INIT('h8)
	) name8064 (
		_w9959_,
		_w9964_,
		_w9965_
	);
	LUT4 #(
		.INIT('h70ff)
	) name8065 (
		_w2046_,
		_w2097_,
		_w9954_,
		_w9965_,
		_w9966_
	);
	LUT2 #(
		.INIT('h8)
	) name8066 (
		\s15_data_i[28]_pad ,
		_w2049_,
		_w9967_
	);
	LUT4 #(
		.INIT('h135f)
	) name8067 (
		\s1_data_i[28]_pad ,
		\s8_data_i[28]_pad ,
		_w9277_,
		_w9410_,
		_w9968_
	);
	LUT4 #(
		.INIT('h153f)
	) name8068 (
		\s4_data_i[28]_pad ,
		\s6_data_i[28]_pad ,
		_w9404_,
		_w9644_,
		_w9969_
	);
	LUT4 #(
		.INIT('h135f)
	) name8069 (
		\s5_data_i[28]_pad ,
		\s9_data_i[28]_pad ,
		_w9401_,
		_w9641_,
		_w9970_
	);
	LUT4 #(
		.INIT('h135f)
	) name8070 (
		\s10_data_i[28]_pad ,
		\s7_data_i[28]_pad ,
		_w9381_,
		_w9407_,
		_w9971_
	);
	LUT4 #(
		.INIT('h8000)
	) name8071 (
		_w9968_,
		_w9969_,
		_w9970_,
		_w9971_,
		_w9972_
	);
	LUT2 #(
		.INIT('h8)
	) name8072 (
		\s11_data_i[28]_pad ,
		_w9384_,
		_w9973_
	);
	LUT4 #(
		.INIT('h135f)
	) name8073 (
		\s14_data_i[28]_pad ,
		\s3_data_i[28]_pad ,
		_w9390_,
		_w9398_,
		_w9974_
	);
	LUT4 #(
		.INIT('h153f)
	) name8074 (
		\s12_data_i[28]_pad ,
		\s2_data_i[28]_pad ,
		_w9395_,
		_w9650_,
		_w9975_
	);
	LUT4 #(
		.INIT('h135f)
	) name8075 (
		\s0_data_i[28]_pad ,
		\s13_data_i[28]_pad ,
		_w9273_,
		_w9647_,
		_w9976_
	);
	LUT4 #(
		.INIT('h4000)
	) name8076 (
		_w9973_,
		_w9974_,
		_w9975_,
		_w9976_,
		_w9977_
	);
	LUT2 #(
		.INIT('h8)
	) name8077 (
		_w9972_,
		_w9977_,
		_w9978_
	);
	LUT4 #(
		.INIT('h70ff)
	) name8078 (
		_w2046_,
		_w2097_,
		_w9967_,
		_w9978_,
		_w9979_
	);
	LUT2 #(
		.INIT('h8)
	) name8079 (
		\s15_data_i[29]_pad ,
		_w2049_,
		_w9980_
	);
	LUT4 #(
		.INIT('h135f)
	) name8080 (
		\s1_data_i[29]_pad ,
		\s8_data_i[29]_pad ,
		_w9277_,
		_w9410_,
		_w9981_
	);
	LUT4 #(
		.INIT('h153f)
	) name8081 (
		\s4_data_i[29]_pad ,
		\s6_data_i[29]_pad ,
		_w9404_,
		_w9644_,
		_w9982_
	);
	LUT4 #(
		.INIT('h135f)
	) name8082 (
		\s5_data_i[29]_pad ,
		\s9_data_i[29]_pad ,
		_w9401_,
		_w9641_,
		_w9983_
	);
	LUT4 #(
		.INIT('h135f)
	) name8083 (
		\s10_data_i[29]_pad ,
		\s7_data_i[29]_pad ,
		_w9381_,
		_w9407_,
		_w9984_
	);
	LUT4 #(
		.INIT('h8000)
	) name8084 (
		_w9981_,
		_w9982_,
		_w9983_,
		_w9984_,
		_w9985_
	);
	LUT2 #(
		.INIT('h8)
	) name8085 (
		\s11_data_i[29]_pad ,
		_w9384_,
		_w9986_
	);
	LUT4 #(
		.INIT('h135f)
	) name8086 (
		\s14_data_i[29]_pad ,
		\s3_data_i[29]_pad ,
		_w9390_,
		_w9398_,
		_w9987_
	);
	LUT4 #(
		.INIT('h153f)
	) name8087 (
		\s12_data_i[29]_pad ,
		\s2_data_i[29]_pad ,
		_w9395_,
		_w9650_,
		_w9988_
	);
	LUT4 #(
		.INIT('h135f)
	) name8088 (
		\s0_data_i[29]_pad ,
		\s13_data_i[29]_pad ,
		_w9273_,
		_w9647_,
		_w9989_
	);
	LUT4 #(
		.INIT('h4000)
	) name8089 (
		_w9986_,
		_w9987_,
		_w9988_,
		_w9989_,
		_w9990_
	);
	LUT2 #(
		.INIT('h8)
	) name8090 (
		_w9985_,
		_w9990_,
		_w9991_
	);
	LUT4 #(
		.INIT('h70ff)
	) name8091 (
		_w2046_,
		_w2097_,
		_w9980_,
		_w9991_,
		_w9992_
	);
	LUT4 #(
		.INIT('h0002)
	) name8092 (
		\rf_rf_dout_reg[2]/P0001 ,
		_w2016_,
		_w2029_,
		_w2043_,
		_w9993_
	);
	LUT3 #(
		.INIT('h80)
	) name8093 (
		_w2049_,
		_w2097_,
		_w9993_,
		_w9994_
	);
	LUT2 #(
		.INIT('h8)
	) name8094 (
		\s15_data_i[2]_pad ,
		_w2049_,
		_w9995_
	);
	LUT3 #(
		.INIT('h70)
	) name8095 (
		_w2046_,
		_w2097_,
		_w9995_,
		_w9996_
	);
	LUT4 #(
		.INIT('h135f)
	) name8096 (
		\s1_data_i[2]_pad ,
		\s8_data_i[2]_pad ,
		_w9277_,
		_w9410_,
		_w9997_
	);
	LUT4 #(
		.INIT('h153f)
	) name8097 (
		\s4_data_i[2]_pad ,
		\s6_data_i[2]_pad ,
		_w9404_,
		_w9644_,
		_w9998_
	);
	LUT4 #(
		.INIT('h135f)
	) name8098 (
		\s5_data_i[2]_pad ,
		\s9_data_i[2]_pad ,
		_w9401_,
		_w9641_,
		_w9999_
	);
	LUT4 #(
		.INIT('h135f)
	) name8099 (
		\s10_data_i[2]_pad ,
		\s7_data_i[2]_pad ,
		_w9381_,
		_w9407_,
		_w10000_
	);
	LUT4 #(
		.INIT('h8000)
	) name8100 (
		_w9997_,
		_w9998_,
		_w9999_,
		_w10000_,
		_w10001_
	);
	LUT2 #(
		.INIT('h8)
	) name8101 (
		\s11_data_i[2]_pad ,
		_w9384_,
		_w10002_
	);
	LUT4 #(
		.INIT('h135f)
	) name8102 (
		\s14_data_i[2]_pad ,
		\s3_data_i[2]_pad ,
		_w9390_,
		_w9398_,
		_w10003_
	);
	LUT4 #(
		.INIT('h153f)
	) name8103 (
		\s12_data_i[2]_pad ,
		\s2_data_i[2]_pad ,
		_w9395_,
		_w9650_,
		_w10004_
	);
	LUT4 #(
		.INIT('h135f)
	) name8104 (
		\s0_data_i[2]_pad ,
		\s13_data_i[2]_pad ,
		_w9273_,
		_w9647_,
		_w10005_
	);
	LUT4 #(
		.INIT('h4000)
	) name8105 (
		_w10002_,
		_w10003_,
		_w10004_,
		_w10005_,
		_w10006_
	);
	LUT2 #(
		.INIT('h8)
	) name8106 (
		_w10001_,
		_w10006_,
		_w10007_
	);
	LUT3 #(
		.INIT('hef)
	) name8107 (
		_w9994_,
		_w9996_,
		_w10007_,
		_w10008_
	);
	LUT2 #(
		.INIT('h8)
	) name8108 (
		\s15_data_i[30]_pad ,
		_w2049_,
		_w10009_
	);
	LUT4 #(
		.INIT('h135f)
	) name8109 (
		\s1_data_i[30]_pad ,
		\s8_data_i[30]_pad ,
		_w9277_,
		_w9410_,
		_w10010_
	);
	LUT4 #(
		.INIT('h153f)
	) name8110 (
		\s4_data_i[30]_pad ,
		\s6_data_i[30]_pad ,
		_w9404_,
		_w9644_,
		_w10011_
	);
	LUT4 #(
		.INIT('h135f)
	) name8111 (
		\s5_data_i[30]_pad ,
		\s9_data_i[30]_pad ,
		_w9401_,
		_w9641_,
		_w10012_
	);
	LUT4 #(
		.INIT('h135f)
	) name8112 (
		\s10_data_i[30]_pad ,
		\s7_data_i[30]_pad ,
		_w9381_,
		_w9407_,
		_w10013_
	);
	LUT4 #(
		.INIT('h8000)
	) name8113 (
		_w10010_,
		_w10011_,
		_w10012_,
		_w10013_,
		_w10014_
	);
	LUT2 #(
		.INIT('h8)
	) name8114 (
		\s11_data_i[30]_pad ,
		_w9384_,
		_w10015_
	);
	LUT4 #(
		.INIT('h135f)
	) name8115 (
		\s14_data_i[30]_pad ,
		\s3_data_i[30]_pad ,
		_w9390_,
		_w9398_,
		_w10016_
	);
	LUT4 #(
		.INIT('h153f)
	) name8116 (
		\s12_data_i[30]_pad ,
		\s2_data_i[30]_pad ,
		_w9395_,
		_w9650_,
		_w10017_
	);
	LUT4 #(
		.INIT('h135f)
	) name8117 (
		\s0_data_i[30]_pad ,
		\s13_data_i[30]_pad ,
		_w9273_,
		_w9647_,
		_w10018_
	);
	LUT4 #(
		.INIT('h4000)
	) name8118 (
		_w10015_,
		_w10016_,
		_w10017_,
		_w10018_,
		_w10019_
	);
	LUT2 #(
		.INIT('h8)
	) name8119 (
		_w10014_,
		_w10019_,
		_w10020_
	);
	LUT4 #(
		.INIT('h70ff)
	) name8120 (
		_w2046_,
		_w2097_,
		_w10009_,
		_w10020_,
		_w10021_
	);
	LUT2 #(
		.INIT('h8)
	) name8121 (
		\s15_data_i[31]_pad ,
		_w2049_,
		_w10022_
	);
	LUT4 #(
		.INIT('h135f)
	) name8122 (
		\s1_data_i[31]_pad ,
		\s8_data_i[31]_pad ,
		_w9277_,
		_w9410_,
		_w10023_
	);
	LUT4 #(
		.INIT('h153f)
	) name8123 (
		\s4_data_i[31]_pad ,
		\s6_data_i[31]_pad ,
		_w9404_,
		_w9644_,
		_w10024_
	);
	LUT4 #(
		.INIT('h135f)
	) name8124 (
		\s5_data_i[31]_pad ,
		\s9_data_i[31]_pad ,
		_w9401_,
		_w9641_,
		_w10025_
	);
	LUT4 #(
		.INIT('h135f)
	) name8125 (
		\s10_data_i[31]_pad ,
		\s7_data_i[31]_pad ,
		_w9381_,
		_w9407_,
		_w10026_
	);
	LUT4 #(
		.INIT('h8000)
	) name8126 (
		_w10023_,
		_w10024_,
		_w10025_,
		_w10026_,
		_w10027_
	);
	LUT2 #(
		.INIT('h8)
	) name8127 (
		\s11_data_i[31]_pad ,
		_w9384_,
		_w10028_
	);
	LUT4 #(
		.INIT('h135f)
	) name8128 (
		\s14_data_i[31]_pad ,
		\s3_data_i[31]_pad ,
		_w9390_,
		_w9398_,
		_w10029_
	);
	LUT4 #(
		.INIT('h153f)
	) name8129 (
		\s12_data_i[31]_pad ,
		\s2_data_i[31]_pad ,
		_w9395_,
		_w9650_,
		_w10030_
	);
	LUT4 #(
		.INIT('h135f)
	) name8130 (
		\s0_data_i[31]_pad ,
		\s13_data_i[31]_pad ,
		_w9273_,
		_w9647_,
		_w10031_
	);
	LUT4 #(
		.INIT('h4000)
	) name8131 (
		_w10028_,
		_w10029_,
		_w10030_,
		_w10031_,
		_w10032_
	);
	LUT2 #(
		.INIT('h8)
	) name8132 (
		_w10027_,
		_w10032_,
		_w10033_
	);
	LUT4 #(
		.INIT('h70ff)
	) name8133 (
		_w2046_,
		_w2097_,
		_w10022_,
		_w10033_,
		_w10034_
	);
	LUT4 #(
		.INIT('h0002)
	) name8134 (
		\rf_rf_dout_reg[3]/P0001 ,
		_w2016_,
		_w2029_,
		_w2043_,
		_w10035_
	);
	LUT3 #(
		.INIT('h80)
	) name8135 (
		_w2049_,
		_w2097_,
		_w10035_,
		_w10036_
	);
	LUT2 #(
		.INIT('h8)
	) name8136 (
		\s15_data_i[3]_pad ,
		_w2049_,
		_w10037_
	);
	LUT3 #(
		.INIT('h70)
	) name8137 (
		_w2046_,
		_w2097_,
		_w10037_,
		_w10038_
	);
	LUT4 #(
		.INIT('h135f)
	) name8138 (
		\s1_data_i[3]_pad ,
		\s8_data_i[3]_pad ,
		_w9277_,
		_w9410_,
		_w10039_
	);
	LUT4 #(
		.INIT('h153f)
	) name8139 (
		\s4_data_i[3]_pad ,
		\s6_data_i[3]_pad ,
		_w9404_,
		_w9644_,
		_w10040_
	);
	LUT4 #(
		.INIT('h135f)
	) name8140 (
		\s5_data_i[3]_pad ,
		\s9_data_i[3]_pad ,
		_w9401_,
		_w9641_,
		_w10041_
	);
	LUT4 #(
		.INIT('h135f)
	) name8141 (
		\s10_data_i[3]_pad ,
		\s7_data_i[3]_pad ,
		_w9381_,
		_w9407_,
		_w10042_
	);
	LUT4 #(
		.INIT('h8000)
	) name8142 (
		_w10039_,
		_w10040_,
		_w10041_,
		_w10042_,
		_w10043_
	);
	LUT2 #(
		.INIT('h8)
	) name8143 (
		\s11_data_i[3]_pad ,
		_w9384_,
		_w10044_
	);
	LUT4 #(
		.INIT('h135f)
	) name8144 (
		\s14_data_i[3]_pad ,
		\s3_data_i[3]_pad ,
		_w9390_,
		_w9398_,
		_w10045_
	);
	LUT4 #(
		.INIT('h153f)
	) name8145 (
		\s12_data_i[3]_pad ,
		\s2_data_i[3]_pad ,
		_w9395_,
		_w9650_,
		_w10046_
	);
	LUT4 #(
		.INIT('h135f)
	) name8146 (
		\s0_data_i[3]_pad ,
		\s13_data_i[3]_pad ,
		_w9273_,
		_w9647_,
		_w10047_
	);
	LUT4 #(
		.INIT('h4000)
	) name8147 (
		_w10044_,
		_w10045_,
		_w10046_,
		_w10047_,
		_w10048_
	);
	LUT2 #(
		.INIT('h8)
	) name8148 (
		_w10043_,
		_w10048_,
		_w10049_
	);
	LUT3 #(
		.INIT('hef)
	) name8149 (
		_w10036_,
		_w10038_,
		_w10049_,
		_w10050_
	);
	LUT4 #(
		.INIT('h0002)
	) name8150 (
		\rf_rf_dout_reg[4]/P0001 ,
		_w2016_,
		_w2029_,
		_w2043_,
		_w10051_
	);
	LUT3 #(
		.INIT('h80)
	) name8151 (
		_w2049_,
		_w2097_,
		_w10051_,
		_w10052_
	);
	LUT2 #(
		.INIT('h8)
	) name8152 (
		\s15_data_i[4]_pad ,
		_w2049_,
		_w10053_
	);
	LUT3 #(
		.INIT('h70)
	) name8153 (
		_w2046_,
		_w2097_,
		_w10053_,
		_w10054_
	);
	LUT4 #(
		.INIT('h135f)
	) name8154 (
		\s1_data_i[4]_pad ,
		\s8_data_i[4]_pad ,
		_w9277_,
		_w9410_,
		_w10055_
	);
	LUT4 #(
		.INIT('h153f)
	) name8155 (
		\s4_data_i[4]_pad ,
		\s6_data_i[4]_pad ,
		_w9404_,
		_w9644_,
		_w10056_
	);
	LUT4 #(
		.INIT('h135f)
	) name8156 (
		\s5_data_i[4]_pad ,
		\s9_data_i[4]_pad ,
		_w9401_,
		_w9641_,
		_w10057_
	);
	LUT4 #(
		.INIT('h135f)
	) name8157 (
		\s10_data_i[4]_pad ,
		\s7_data_i[4]_pad ,
		_w9381_,
		_w9407_,
		_w10058_
	);
	LUT4 #(
		.INIT('h8000)
	) name8158 (
		_w10055_,
		_w10056_,
		_w10057_,
		_w10058_,
		_w10059_
	);
	LUT2 #(
		.INIT('h8)
	) name8159 (
		\s11_data_i[4]_pad ,
		_w9384_,
		_w10060_
	);
	LUT4 #(
		.INIT('h135f)
	) name8160 (
		\s14_data_i[4]_pad ,
		\s3_data_i[4]_pad ,
		_w9390_,
		_w9398_,
		_w10061_
	);
	LUT4 #(
		.INIT('h153f)
	) name8161 (
		\s12_data_i[4]_pad ,
		\s2_data_i[4]_pad ,
		_w9395_,
		_w9650_,
		_w10062_
	);
	LUT4 #(
		.INIT('h135f)
	) name8162 (
		\s0_data_i[4]_pad ,
		\s13_data_i[4]_pad ,
		_w9273_,
		_w9647_,
		_w10063_
	);
	LUT4 #(
		.INIT('h4000)
	) name8163 (
		_w10060_,
		_w10061_,
		_w10062_,
		_w10063_,
		_w10064_
	);
	LUT2 #(
		.INIT('h8)
	) name8164 (
		_w10059_,
		_w10064_,
		_w10065_
	);
	LUT3 #(
		.INIT('hef)
	) name8165 (
		_w10052_,
		_w10054_,
		_w10065_,
		_w10066_
	);
	LUT4 #(
		.INIT('h0002)
	) name8166 (
		\rf_rf_dout_reg[5]/P0001 ,
		_w2016_,
		_w2029_,
		_w2043_,
		_w10067_
	);
	LUT3 #(
		.INIT('h80)
	) name8167 (
		_w2049_,
		_w2097_,
		_w10067_,
		_w10068_
	);
	LUT2 #(
		.INIT('h8)
	) name8168 (
		\s15_data_i[5]_pad ,
		_w2049_,
		_w10069_
	);
	LUT3 #(
		.INIT('h70)
	) name8169 (
		_w2046_,
		_w2097_,
		_w10069_,
		_w10070_
	);
	LUT4 #(
		.INIT('h135f)
	) name8170 (
		\s1_data_i[5]_pad ,
		\s8_data_i[5]_pad ,
		_w9277_,
		_w9410_,
		_w10071_
	);
	LUT4 #(
		.INIT('h153f)
	) name8171 (
		\s4_data_i[5]_pad ,
		\s6_data_i[5]_pad ,
		_w9404_,
		_w9644_,
		_w10072_
	);
	LUT4 #(
		.INIT('h135f)
	) name8172 (
		\s5_data_i[5]_pad ,
		\s9_data_i[5]_pad ,
		_w9401_,
		_w9641_,
		_w10073_
	);
	LUT4 #(
		.INIT('h135f)
	) name8173 (
		\s10_data_i[5]_pad ,
		\s7_data_i[5]_pad ,
		_w9381_,
		_w9407_,
		_w10074_
	);
	LUT4 #(
		.INIT('h8000)
	) name8174 (
		_w10071_,
		_w10072_,
		_w10073_,
		_w10074_,
		_w10075_
	);
	LUT2 #(
		.INIT('h8)
	) name8175 (
		\s11_data_i[5]_pad ,
		_w9384_,
		_w10076_
	);
	LUT4 #(
		.INIT('h135f)
	) name8176 (
		\s14_data_i[5]_pad ,
		\s3_data_i[5]_pad ,
		_w9390_,
		_w9398_,
		_w10077_
	);
	LUT4 #(
		.INIT('h153f)
	) name8177 (
		\s12_data_i[5]_pad ,
		\s2_data_i[5]_pad ,
		_w9395_,
		_w9650_,
		_w10078_
	);
	LUT4 #(
		.INIT('h135f)
	) name8178 (
		\s0_data_i[5]_pad ,
		\s13_data_i[5]_pad ,
		_w9273_,
		_w9647_,
		_w10079_
	);
	LUT4 #(
		.INIT('h4000)
	) name8179 (
		_w10076_,
		_w10077_,
		_w10078_,
		_w10079_,
		_w10080_
	);
	LUT2 #(
		.INIT('h8)
	) name8180 (
		_w10075_,
		_w10080_,
		_w10081_
	);
	LUT3 #(
		.INIT('hef)
	) name8181 (
		_w10068_,
		_w10070_,
		_w10081_,
		_w10082_
	);
	LUT4 #(
		.INIT('h0002)
	) name8182 (
		\rf_rf_dout_reg[6]/P0001 ,
		_w2016_,
		_w2029_,
		_w2043_,
		_w10083_
	);
	LUT3 #(
		.INIT('h80)
	) name8183 (
		_w2049_,
		_w2097_,
		_w10083_,
		_w10084_
	);
	LUT2 #(
		.INIT('h8)
	) name8184 (
		\s15_data_i[6]_pad ,
		_w2049_,
		_w10085_
	);
	LUT3 #(
		.INIT('h70)
	) name8185 (
		_w2046_,
		_w2097_,
		_w10085_,
		_w10086_
	);
	LUT4 #(
		.INIT('h135f)
	) name8186 (
		\s1_data_i[6]_pad ,
		\s8_data_i[6]_pad ,
		_w9277_,
		_w9410_,
		_w10087_
	);
	LUT4 #(
		.INIT('h153f)
	) name8187 (
		\s4_data_i[6]_pad ,
		\s6_data_i[6]_pad ,
		_w9404_,
		_w9644_,
		_w10088_
	);
	LUT4 #(
		.INIT('h135f)
	) name8188 (
		\s5_data_i[6]_pad ,
		\s9_data_i[6]_pad ,
		_w9401_,
		_w9641_,
		_w10089_
	);
	LUT4 #(
		.INIT('h135f)
	) name8189 (
		\s10_data_i[6]_pad ,
		\s7_data_i[6]_pad ,
		_w9381_,
		_w9407_,
		_w10090_
	);
	LUT4 #(
		.INIT('h8000)
	) name8190 (
		_w10087_,
		_w10088_,
		_w10089_,
		_w10090_,
		_w10091_
	);
	LUT2 #(
		.INIT('h8)
	) name8191 (
		\s11_data_i[6]_pad ,
		_w9384_,
		_w10092_
	);
	LUT4 #(
		.INIT('h135f)
	) name8192 (
		\s14_data_i[6]_pad ,
		\s3_data_i[6]_pad ,
		_w9390_,
		_w9398_,
		_w10093_
	);
	LUT4 #(
		.INIT('h153f)
	) name8193 (
		\s12_data_i[6]_pad ,
		\s2_data_i[6]_pad ,
		_w9395_,
		_w9650_,
		_w10094_
	);
	LUT4 #(
		.INIT('h135f)
	) name8194 (
		\s0_data_i[6]_pad ,
		\s13_data_i[6]_pad ,
		_w9273_,
		_w9647_,
		_w10095_
	);
	LUT4 #(
		.INIT('h4000)
	) name8195 (
		_w10092_,
		_w10093_,
		_w10094_,
		_w10095_,
		_w10096_
	);
	LUT2 #(
		.INIT('h8)
	) name8196 (
		_w10091_,
		_w10096_,
		_w10097_
	);
	LUT3 #(
		.INIT('hef)
	) name8197 (
		_w10084_,
		_w10086_,
		_w10097_,
		_w10098_
	);
	LUT4 #(
		.INIT('h0002)
	) name8198 (
		\rf_rf_dout_reg[7]/P0001 ,
		_w2016_,
		_w2029_,
		_w2043_,
		_w10099_
	);
	LUT3 #(
		.INIT('h80)
	) name8199 (
		_w2049_,
		_w2097_,
		_w10099_,
		_w10100_
	);
	LUT2 #(
		.INIT('h8)
	) name8200 (
		\s15_data_i[7]_pad ,
		_w2049_,
		_w10101_
	);
	LUT3 #(
		.INIT('h70)
	) name8201 (
		_w2046_,
		_w2097_,
		_w10101_,
		_w10102_
	);
	LUT4 #(
		.INIT('h135f)
	) name8202 (
		\s1_data_i[7]_pad ,
		\s8_data_i[7]_pad ,
		_w9277_,
		_w9410_,
		_w10103_
	);
	LUT4 #(
		.INIT('h153f)
	) name8203 (
		\s4_data_i[7]_pad ,
		\s6_data_i[7]_pad ,
		_w9404_,
		_w9644_,
		_w10104_
	);
	LUT4 #(
		.INIT('h135f)
	) name8204 (
		\s5_data_i[7]_pad ,
		\s9_data_i[7]_pad ,
		_w9401_,
		_w9641_,
		_w10105_
	);
	LUT4 #(
		.INIT('h135f)
	) name8205 (
		\s10_data_i[7]_pad ,
		\s7_data_i[7]_pad ,
		_w9381_,
		_w9407_,
		_w10106_
	);
	LUT4 #(
		.INIT('h8000)
	) name8206 (
		_w10103_,
		_w10104_,
		_w10105_,
		_w10106_,
		_w10107_
	);
	LUT2 #(
		.INIT('h8)
	) name8207 (
		\s11_data_i[7]_pad ,
		_w9384_,
		_w10108_
	);
	LUT4 #(
		.INIT('h135f)
	) name8208 (
		\s14_data_i[7]_pad ,
		\s3_data_i[7]_pad ,
		_w9390_,
		_w9398_,
		_w10109_
	);
	LUT4 #(
		.INIT('h153f)
	) name8209 (
		\s12_data_i[7]_pad ,
		\s2_data_i[7]_pad ,
		_w9395_,
		_w9650_,
		_w10110_
	);
	LUT4 #(
		.INIT('h135f)
	) name8210 (
		\s0_data_i[7]_pad ,
		\s13_data_i[7]_pad ,
		_w9273_,
		_w9647_,
		_w10111_
	);
	LUT4 #(
		.INIT('h4000)
	) name8211 (
		_w10108_,
		_w10109_,
		_w10110_,
		_w10111_,
		_w10112_
	);
	LUT2 #(
		.INIT('h8)
	) name8212 (
		_w10107_,
		_w10112_,
		_w10113_
	);
	LUT3 #(
		.INIT('hef)
	) name8213 (
		_w10100_,
		_w10102_,
		_w10113_,
		_w10114_
	);
	LUT4 #(
		.INIT('h0002)
	) name8214 (
		\rf_rf_dout_reg[8]/P0001 ,
		_w2016_,
		_w2029_,
		_w2043_,
		_w10115_
	);
	LUT3 #(
		.INIT('h80)
	) name8215 (
		_w2049_,
		_w2097_,
		_w10115_,
		_w10116_
	);
	LUT2 #(
		.INIT('h8)
	) name8216 (
		\s15_data_i[8]_pad ,
		_w2049_,
		_w10117_
	);
	LUT3 #(
		.INIT('h70)
	) name8217 (
		_w2046_,
		_w2097_,
		_w10117_,
		_w10118_
	);
	LUT4 #(
		.INIT('h135f)
	) name8218 (
		\s1_data_i[8]_pad ,
		\s8_data_i[8]_pad ,
		_w9277_,
		_w9410_,
		_w10119_
	);
	LUT4 #(
		.INIT('h153f)
	) name8219 (
		\s4_data_i[8]_pad ,
		\s6_data_i[8]_pad ,
		_w9404_,
		_w9644_,
		_w10120_
	);
	LUT4 #(
		.INIT('h135f)
	) name8220 (
		\s5_data_i[8]_pad ,
		\s9_data_i[8]_pad ,
		_w9401_,
		_w9641_,
		_w10121_
	);
	LUT4 #(
		.INIT('h135f)
	) name8221 (
		\s10_data_i[8]_pad ,
		\s7_data_i[8]_pad ,
		_w9381_,
		_w9407_,
		_w10122_
	);
	LUT4 #(
		.INIT('h8000)
	) name8222 (
		_w10119_,
		_w10120_,
		_w10121_,
		_w10122_,
		_w10123_
	);
	LUT2 #(
		.INIT('h8)
	) name8223 (
		\s11_data_i[8]_pad ,
		_w9384_,
		_w10124_
	);
	LUT4 #(
		.INIT('h135f)
	) name8224 (
		\s14_data_i[8]_pad ,
		\s3_data_i[8]_pad ,
		_w9390_,
		_w9398_,
		_w10125_
	);
	LUT4 #(
		.INIT('h153f)
	) name8225 (
		\s12_data_i[8]_pad ,
		\s2_data_i[8]_pad ,
		_w9395_,
		_w9650_,
		_w10126_
	);
	LUT4 #(
		.INIT('h135f)
	) name8226 (
		\s0_data_i[8]_pad ,
		\s13_data_i[8]_pad ,
		_w9273_,
		_w9647_,
		_w10127_
	);
	LUT4 #(
		.INIT('h4000)
	) name8227 (
		_w10124_,
		_w10125_,
		_w10126_,
		_w10127_,
		_w10128_
	);
	LUT2 #(
		.INIT('h8)
	) name8228 (
		_w10123_,
		_w10128_,
		_w10129_
	);
	LUT3 #(
		.INIT('hef)
	) name8229 (
		_w10116_,
		_w10118_,
		_w10129_,
		_w10130_
	);
	LUT4 #(
		.INIT('h0002)
	) name8230 (
		\rf_rf_dout_reg[9]/P0001 ,
		_w2016_,
		_w2029_,
		_w2043_,
		_w10131_
	);
	LUT3 #(
		.INIT('h80)
	) name8231 (
		_w2049_,
		_w2097_,
		_w10131_,
		_w10132_
	);
	LUT2 #(
		.INIT('h8)
	) name8232 (
		\s15_data_i[9]_pad ,
		_w2049_,
		_w10133_
	);
	LUT3 #(
		.INIT('h70)
	) name8233 (
		_w2046_,
		_w2097_,
		_w10133_,
		_w10134_
	);
	LUT4 #(
		.INIT('h135f)
	) name8234 (
		\s1_data_i[9]_pad ,
		\s8_data_i[9]_pad ,
		_w9277_,
		_w9410_,
		_w10135_
	);
	LUT4 #(
		.INIT('h153f)
	) name8235 (
		\s4_data_i[9]_pad ,
		\s6_data_i[9]_pad ,
		_w9404_,
		_w9644_,
		_w10136_
	);
	LUT4 #(
		.INIT('h135f)
	) name8236 (
		\s5_data_i[9]_pad ,
		\s9_data_i[9]_pad ,
		_w9401_,
		_w9641_,
		_w10137_
	);
	LUT4 #(
		.INIT('h135f)
	) name8237 (
		\s10_data_i[9]_pad ,
		\s7_data_i[9]_pad ,
		_w9381_,
		_w9407_,
		_w10138_
	);
	LUT4 #(
		.INIT('h8000)
	) name8238 (
		_w10135_,
		_w10136_,
		_w10137_,
		_w10138_,
		_w10139_
	);
	LUT2 #(
		.INIT('h8)
	) name8239 (
		\s11_data_i[9]_pad ,
		_w9384_,
		_w10140_
	);
	LUT4 #(
		.INIT('h135f)
	) name8240 (
		\s14_data_i[9]_pad ,
		\s3_data_i[9]_pad ,
		_w9390_,
		_w9398_,
		_w10141_
	);
	LUT4 #(
		.INIT('h153f)
	) name8241 (
		\s12_data_i[9]_pad ,
		\s2_data_i[9]_pad ,
		_w9395_,
		_w9650_,
		_w10142_
	);
	LUT4 #(
		.INIT('h135f)
	) name8242 (
		\s0_data_i[9]_pad ,
		\s13_data_i[9]_pad ,
		_w9273_,
		_w9647_,
		_w10143_
	);
	LUT4 #(
		.INIT('h4000)
	) name8243 (
		_w10140_,
		_w10141_,
		_w10142_,
		_w10143_,
		_w10144_
	);
	LUT2 #(
		.INIT('h8)
	) name8244 (
		_w10139_,
		_w10144_,
		_w10145_
	);
	LUT3 #(
		.INIT('hef)
	) name8245 (
		_w10132_,
		_w10134_,
		_w10145_,
		_w10146_
	);
	LUT3 #(
		.INIT('h80)
	) name8246 (
		\s15_err_i_pad ,
		_w1914_,
		_w9653_,
		_w10147_
	);
	LUT4 #(
		.INIT('h8000)
	) name8247 (
		\s0_err_i_pad ,
		_w8989_,
		_w8990_,
		_w9273_,
		_w10148_
	);
	LUT4 #(
		.INIT('h8000)
	) name8248 (
		\s8_err_i_pad ,
		_w8821_,
		_w8822_,
		_w9410_,
		_w10149_
	);
	LUT4 #(
		.INIT('h153f)
	) name8249 (
		_w8820_,
		_w9008_,
		_w10148_,
		_w10149_,
		_w10150_
	);
	LUT4 #(
		.INIT('h8000)
	) name8250 (
		\s3_err_i_pad ,
		_w9205_,
		_w9206_,
		_w9398_,
		_w10151_
	);
	LUT4 #(
		.INIT('h8000)
	) name8251 (
		\s14_err_i_pad ,
		_w9137_,
		_w9138_,
		_w9390_,
		_w10152_
	);
	LUT4 #(
		.INIT('h153f)
	) name8252 (
		_w9136_,
		_w9224_,
		_w10151_,
		_w10152_,
		_w10153_
	);
	LUT4 #(
		.INIT('h8000)
	) name8253 (
		\s7_err_i_pad ,
		_w8782_,
		_w8783_,
		_w9407_,
		_w10154_
	);
	LUT4 #(
		.INIT('h8000)
	) name8254 (
		\s5_err_i_pad ,
		_w8699_,
		_w8700_,
		_w9401_,
		_w10155_
	);
	LUT4 #(
		.INIT('h153f)
	) name8255 (
		_w8718_,
		_w8789_,
		_w10154_,
		_w10155_,
		_w10156_
	);
	LUT4 #(
		.INIT('h8000)
	) name8256 (
		\s12_err_i_pad ,
		_w9029_,
		_w9030_,
		_w9650_,
		_w10157_
	);
	LUT4 #(
		.INIT('h8000)
	) name8257 (
		\s13_err_i_pad ,
		_w9069_,
		_w9070_,
		_w9647_,
		_w10158_
	);
	LUT4 #(
		.INIT('h135f)
	) name8258 (
		_w9048_,
		_w9076_,
		_w10157_,
		_w10158_,
		_w10159_
	);
	LUT4 #(
		.INIT('h8000)
	) name8259 (
		_w10150_,
		_w10153_,
		_w10156_,
		_w10159_,
		_w10160_
	);
	LUT4 #(
		.INIT('h8000)
	) name8260 (
		\s4_err_i_pad ,
		_w8655_,
		_w8656_,
		_w9644_,
		_w10161_
	);
	LUT2 #(
		.INIT('h8)
	) name8261 (
		_w8662_,
		_w10161_,
		_w10162_
	);
	LUT4 #(
		.INIT('h8000)
	) name8262 (
		\s1_err_i_pad ,
		_w9103_,
		_w9104_,
		_w9277_,
		_w10163_
	);
	LUT4 #(
		.INIT('h8000)
	) name8263 (
		\s6_err_i_pad ,
		_w8743_,
		_w8744_,
		_w9404_,
		_w10164_
	);
	LUT4 #(
		.INIT('h153f)
	) name8264 (
		_w8742_,
		_w9122_,
		_w10163_,
		_w10164_,
		_w10165_
	);
	LUT4 #(
		.INIT('h8000)
	) name8265 (
		\s9_err_i_pad ,
		_w8865_,
		_w8866_,
		_w9641_,
		_w10166_
	);
	LUT4 #(
		.INIT('h8000)
	) name8266 (
		\s10_err_i_pad ,
		_w8910_,
		_w8911_,
		_w9381_,
		_w10167_
	);
	LUT4 #(
		.INIT('h135f)
	) name8267 (
		_w8872_,
		_w8923_,
		_w10166_,
		_w10167_,
		_w10168_
	);
	LUT4 #(
		.INIT('h8000)
	) name8268 (
		\s11_err_i_pad ,
		_w8955_,
		_w8956_,
		_w9384_,
		_w10169_
	);
	LUT4 #(
		.INIT('h8000)
	) name8269 (
		\s2_err_i_pad ,
		_w9171_,
		_w9172_,
		_w9395_,
		_w10170_
	);
	LUT4 #(
		.INIT('h135f)
	) name8270 (
		_w8962_,
		_w9178_,
		_w10169_,
		_w10170_,
		_w10171_
	);
	LUT4 #(
		.INIT('h4000)
	) name8271 (
		_w10162_,
		_w10165_,
		_w10168_,
		_w10171_,
		_w10172_
	);
	LUT2 #(
		.INIT('h8)
	) name8272 (
		_w10160_,
		_w10172_,
		_w10173_
	);
	LUT4 #(
		.INIT('h70ff)
	) name8273 (
		_w2046_,
		_w2097_,
		_w10147_,
		_w10173_,
		_w10174_
	);
	LUT3 #(
		.INIT('h80)
	) name8274 (
		\s15_rty_i_pad ,
		_w1914_,
		_w9653_,
		_w10175_
	);
	LUT4 #(
		.INIT('h8000)
	) name8275 (
		\s6_rty_i_pad ,
		_w8743_,
		_w8744_,
		_w9404_,
		_w10176_
	);
	LUT4 #(
		.INIT('h8000)
	) name8276 (
		\s12_rty_i_pad ,
		_w9029_,
		_w9030_,
		_w9650_,
		_w10177_
	);
	LUT4 #(
		.INIT('h135f)
	) name8277 (
		_w8742_,
		_w9048_,
		_w10176_,
		_w10177_,
		_w10178_
	);
	LUT4 #(
		.INIT('h8000)
	) name8278 (
		\s3_rty_i_pad ,
		_w9205_,
		_w9206_,
		_w9398_,
		_w10179_
	);
	LUT4 #(
		.INIT('h8000)
	) name8279 (
		\s11_rty_i_pad ,
		_w8955_,
		_w8956_,
		_w9384_,
		_w10180_
	);
	LUT4 #(
		.INIT('h153f)
	) name8280 (
		_w8962_,
		_w9224_,
		_w10179_,
		_w10180_,
		_w10181_
	);
	LUT4 #(
		.INIT('h8000)
	) name8281 (
		\s10_rty_i_pad ,
		_w8910_,
		_w8911_,
		_w9381_,
		_w10182_
	);
	LUT4 #(
		.INIT('h8000)
	) name8282 (
		\s5_rty_i_pad ,
		_w8699_,
		_w8700_,
		_w9401_,
		_w10183_
	);
	LUT4 #(
		.INIT('h153f)
	) name8283 (
		_w8718_,
		_w8923_,
		_w10182_,
		_w10183_,
		_w10184_
	);
	LUT4 #(
		.INIT('h8000)
	) name8284 (
		\s8_rty_i_pad ,
		_w8821_,
		_w8822_,
		_w9410_,
		_w10185_
	);
	LUT4 #(
		.INIT('h8000)
	) name8285 (
		\s13_rty_i_pad ,
		_w9069_,
		_w9070_,
		_w9647_,
		_w10186_
	);
	LUT4 #(
		.INIT('h135f)
	) name8286 (
		_w8820_,
		_w9076_,
		_w10185_,
		_w10186_,
		_w10187_
	);
	LUT4 #(
		.INIT('h8000)
	) name8287 (
		_w10178_,
		_w10181_,
		_w10184_,
		_w10187_,
		_w10188_
	);
	LUT4 #(
		.INIT('h8000)
	) name8288 (
		\s7_rty_i_pad ,
		_w8782_,
		_w8783_,
		_w9407_,
		_w10189_
	);
	LUT2 #(
		.INIT('h8)
	) name8289 (
		_w8789_,
		_w10189_,
		_w10190_
	);
	LUT4 #(
		.INIT('h8000)
	) name8290 (
		\s1_rty_i_pad ,
		_w9103_,
		_w9104_,
		_w9277_,
		_w10191_
	);
	LUT4 #(
		.INIT('h8000)
	) name8291 (
		\s9_rty_i_pad ,
		_w8865_,
		_w8866_,
		_w9641_,
		_w10192_
	);
	LUT4 #(
		.INIT('h153f)
	) name8292 (
		_w8872_,
		_w9122_,
		_w10191_,
		_w10192_,
		_w10193_
	);
	LUT4 #(
		.INIT('h8000)
	) name8293 (
		\s0_rty_i_pad ,
		_w8989_,
		_w8990_,
		_w9273_,
		_w10194_
	);
	LUT4 #(
		.INIT('h8000)
	) name8294 (
		\s4_rty_i_pad ,
		_w8655_,
		_w8656_,
		_w9644_,
		_w10195_
	);
	LUT4 #(
		.INIT('h153f)
	) name8295 (
		_w8662_,
		_w9008_,
		_w10194_,
		_w10195_,
		_w10196_
	);
	LUT4 #(
		.INIT('h8000)
	) name8296 (
		\s14_rty_i_pad ,
		_w9137_,
		_w9138_,
		_w9390_,
		_w10197_
	);
	LUT4 #(
		.INIT('h8000)
	) name8297 (
		\s2_rty_i_pad ,
		_w9171_,
		_w9172_,
		_w9395_,
		_w10198_
	);
	LUT4 #(
		.INIT('h135f)
	) name8298 (
		_w9136_,
		_w9178_,
		_w10197_,
		_w10198_,
		_w10199_
	);
	LUT4 #(
		.INIT('h4000)
	) name8299 (
		_w10190_,
		_w10193_,
		_w10196_,
		_w10199_,
		_w10200_
	);
	LUT2 #(
		.INIT('h8)
	) name8300 (
		_w10188_,
		_w10200_,
		_w10201_
	);
	LUT4 #(
		.INIT('h70ff)
	) name8301 (
		_w2046_,
		_w2097_,
		_w10175_,
		_w10201_,
		_w10202_
	);
	LUT3 #(
		.INIT('h80)
	) name8302 (
		_w1901_,
		_w1902_,
		_w2047_,
		_w10203_
	);
	LUT2 #(
		.INIT('h8)
	) name8303 (
		_w1920_,
		_w10203_,
		_w10204_
	);
	LUT3 #(
		.INIT('h70)
	) name8304 (
		_w2097_,
		_w8630_,
		_w10204_,
		_w10205_
	);
	LUT4 #(
		.INIT('h2a00)
	) name8305 (
		\s5_ack_i_pad ,
		_w8699_,
		_w8700_,
		_w9436_,
		_w10206_
	);
	LUT4 #(
		.INIT('h2a00)
	) name8306 (
		\s1_ack_i_pad ,
		_w9103_,
		_w9104_,
		_w9322_,
		_w10207_
	);
	LUT4 #(
		.INIT('h135f)
	) name8307 (
		_w8718_,
		_w9122_,
		_w10206_,
		_w10207_,
		_w10208_
	);
	LUT4 #(
		.INIT('h2a00)
	) name8308 (
		\s12_ack_i_pad ,
		_w9029_,
		_w9030_,
		_w9635_,
		_w10209_
	);
	LUT4 #(
		.INIT('h2a00)
	) name8309 (
		\s10_ack_i_pad ,
		_w8910_,
		_w8911_,
		_w9413_,
		_w10210_
	);
	LUT4 #(
		.INIT('h153f)
	) name8310 (
		_w8923_,
		_w9048_,
		_w10209_,
		_w10210_,
		_w10211_
	);
	LUT4 #(
		.INIT('h2a00)
	) name8311 (
		\s7_ack_i_pad ,
		_w8782_,
		_w8783_,
		_w9442_,
		_w10212_
	);
	LUT4 #(
		.INIT('h2a00)
	) name8312 (
		\s14_ack_i_pad ,
		_w9137_,
		_w9138_,
		_w9422_,
		_w10213_
	);
	LUT4 #(
		.INIT('h135f)
	) name8313 (
		_w8789_,
		_w9136_,
		_w10212_,
		_w10213_,
		_w10214_
	);
	LUT4 #(
		.INIT('h2a00)
	) name8314 (
		\s13_ack_i_pad ,
		_w9069_,
		_w9070_,
		_w9419_,
		_w10215_
	);
	LUT4 #(
		.INIT('h2a00)
	) name8315 (
		\s9_ack_i_pad ,
		_w8865_,
		_w8866_,
		_w9448_,
		_w10216_
	);
	LUT4 #(
		.INIT('h153f)
	) name8316 (
		_w8872_,
		_w9076_,
		_w10215_,
		_w10216_,
		_w10217_
	);
	LUT4 #(
		.INIT('h8000)
	) name8317 (
		_w10208_,
		_w10211_,
		_w10214_,
		_w10217_,
		_w10218_
	);
	LUT4 #(
		.INIT('h2a00)
	) name8318 (
		\s3_ack_i_pad ,
		_w9205_,
		_w9206_,
		_w9430_,
		_w10219_
	);
	LUT2 #(
		.INIT('h8)
	) name8319 (
		_w9224_,
		_w10219_,
		_w10220_
	);
	LUT4 #(
		.INIT('h2a00)
	) name8320 (
		\s11_ack_i_pad ,
		_w8955_,
		_w8956_,
		_w9638_,
		_w10221_
	);
	LUT4 #(
		.INIT('h2a00)
	) name8321 (
		\s6_ack_i_pad ,
		_w8743_,
		_w8744_,
		_w9439_,
		_w10222_
	);
	LUT4 #(
		.INIT('h153f)
	) name8322 (
		_w8742_,
		_w8962_,
		_w10221_,
		_w10222_,
		_w10223_
	);
	LUT4 #(
		.INIT('h2a00)
	) name8323 (
		\s4_ack_i_pad ,
		_w8655_,
		_w8656_,
		_w9433_,
		_w10224_
	);
	LUT4 #(
		.INIT('h2a00)
	) name8324 (
		\s0_ack_i_pad ,
		_w8989_,
		_w8990_,
		_w9280_,
		_w10225_
	);
	LUT4 #(
		.INIT('h135f)
	) name8325 (
		_w8662_,
		_w9008_,
		_w10224_,
		_w10225_,
		_w10226_
	);
	LUT4 #(
		.INIT('h2a00)
	) name8326 (
		\s2_ack_i_pad ,
		_w9171_,
		_w9172_,
		_w9427_,
		_w10227_
	);
	LUT4 #(
		.INIT('h2a00)
	) name8327 (
		\s8_ack_i_pad ,
		_w8821_,
		_w8822_,
		_w9445_,
		_w10228_
	);
	LUT4 #(
		.INIT('h153f)
	) name8328 (
		_w8820_,
		_w9178_,
		_w10227_,
		_w10228_,
		_w10229_
	);
	LUT4 #(
		.INIT('h4000)
	) name8329 (
		_w10220_,
		_w10223_,
		_w10226_,
		_w10229_,
		_w10230_
	);
	LUT2 #(
		.INIT('h8)
	) name8330 (
		_w10218_,
		_w10230_,
		_w10231_
	);
	LUT3 #(
		.INIT('h4f)
	) name8331 (
		_w9652_,
		_w10205_,
		_w10231_,
		_w10232_
	);
	LUT3 #(
		.INIT('h80)
	) name8332 (
		_w2047_,
		_w2097_,
		_w9683_,
		_w10233_
	);
	LUT2 #(
		.INIT('h8)
	) name8333 (
		\s15_data_i[0]_pad ,
		_w2047_,
		_w10234_
	);
	LUT3 #(
		.INIT('h70)
	) name8334 (
		_w2046_,
		_w2097_,
		_w10234_,
		_w10235_
	);
	LUT4 #(
		.INIT('h153f)
	) name8335 (
		\s12_data_i[0]_pad ,
		\s1_data_i[0]_pad ,
		_w9322_,
		_w9635_,
		_w10236_
	);
	LUT4 #(
		.INIT('h135f)
	) name8336 (
		\s0_data_i[0]_pad ,
		\s10_data_i[0]_pad ,
		_w9280_,
		_w9413_,
		_w10237_
	);
	LUT4 #(
		.INIT('h135f)
	) name8337 (
		\s3_data_i[0]_pad ,
		\s4_data_i[0]_pad ,
		_w9430_,
		_w9433_,
		_w10238_
	);
	LUT4 #(
		.INIT('h135f)
	) name8338 (
		\s6_data_i[0]_pad ,
		\s9_data_i[0]_pad ,
		_w9439_,
		_w9448_,
		_w10239_
	);
	LUT4 #(
		.INIT('h8000)
	) name8339 (
		_w10236_,
		_w10237_,
		_w10238_,
		_w10239_,
		_w10240_
	);
	LUT2 #(
		.INIT('h8)
	) name8340 (
		\s14_data_i[0]_pad ,
		_w9422_,
		_w10241_
	);
	LUT4 #(
		.INIT('h153f)
	) name8341 (
		\s11_data_i[0]_pad ,
		\s7_data_i[0]_pad ,
		_w9442_,
		_w9638_,
		_w10242_
	);
	LUT4 #(
		.INIT('h135f)
	) name8342 (
		\s5_data_i[0]_pad ,
		\s8_data_i[0]_pad ,
		_w9436_,
		_w9445_,
		_w10243_
	);
	LUT4 #(
		.INIT('h135f)
	) name8343 (
		\s13_data_i[0]_pad ,
		\s2_data_i[0]_pad ,
		_w9419_,
		_w9427_,
		_w10244_
	);
	LUT4 #(
		.INIT('h4000)
	) name8344 (
		_w10241_,
		_w10242_,
		_w10243_,
		_w10244_,
		_w10245_
	);
	LUT2 #(
		.INIT('h8)
	) name8345 (
		_w10240_,
		_w10245_,
		_w10246_
	);
	LUT3 #(
		.INIT('hef)
	) name8346 (
		_w10233_,
		_w10235_,
		_w10246_,
		_w10247_
	);
	LUT3 #(
		.INIT('h80)
	) name8347 (
		_w2047_,
		_w2097_,
		_w9699_,
		_w10248_
	);
	LUT2 #(
		.INIT('h8)
	) name8348 (
		\s15_data_i[10]_pad ,
		_w2047_,
		_w10249_
	);
	LUT3 #(
		.INIT('h70)
	) name8349 (
		_w2046_,
		_w2097_,
		_w10249_,
		_w10250_
	);
	LUT4 #(
		.INIT('h153f)
	) name8350 (
		\s12_data_i[10]_pad ,
		\s1_data_i[10]_pad ,
		_w9322_,
		_w9635_,
		_w10251_
	);
	LUT4 #(
		.INIT('h135f)
	) name8351 (
		\s0_data_i[10]_pad ,
		\s10_data_i[10]_pad ,
		_w9280_,
		_w9413_,
		_w10252_
	);
	LUT4 #(
		.INIT('h135f)
	) name8352 (
		\s3_data_i[10]_pad ,
		\s4_data_i[10]_pad ,
		_w9430_,
		_w9433_,
		_w10253_
	);
	LUT4 #(
		.INIT('h135f)
	) name8353 (
		\s6_data_i[10]_pad ,
		\s9_data_i[10]_pad ,
		_w9439_,
		_w9448_,
		_w10254_
	);
	LUT4 #(
		.INIT('h8000)
	) name8354 (
		_w10251_,
		_w10252_,
		_w10253_,
		_w10254_,
		_w10255_
	);
	LUT2 #(
		.INIT('h8)
	) name8355 (
		\s14_data_i[10]_pad ,
		_w9422_,
		_w10256_
	);
	LUT4 #(
		.INIT('h153f)
	) name8356 (
		\s11_data_i[10]_pad ,
		\s7_data_i[10]_pad ,
		_w9442_,
		_w9638_,
		_w10257_
	);
	LUT4 #(
		.INIT('h135f)
	) name8357 (
		\s5_data_i[10]_pad ,
		\s8_data_i[10]_pad ,
		_w9436_,
		_w9445_,
		_w10258_
	);
	LUT4 #(
		.INIT('h135f)
	) name8358 (
		\s13_data_i[10]_pad ,
		\s2_data_i[10]_pad ,
		_w9419_,
		_w9427_,
		_w10259_
	);
	LUT4 #(
		.INIT('h4000)
	) name8359 (
		_w10256_,
		_w10257_,
		_w10258_,
		_w10259_,
		_w10260_
	);
	LUT2 #(
		.INIT('h8)
	) name8360 (
		_w10255_,
		_w10260_,
		_w10261_
	);
	LUT3 #(
		.INIT('hef)
	) name8361 (
		_w10248_,
		_w10250_,
		_w10261_,
		_w10262_
	);
	LUT3 #(
		.INIT('h80)
	) name8362 (
		_w2047_,
		_w2097_,
		_w9715_,
		_w10263_
	);
	LUT2 #(
		.INIT('h8)
	) name8363 (
		\s15_data_i[11]_pad ,
		_w2047_,
		_w10264_
	);
	LUT3 #(
		.INIT('h70)
	) name8364 (
		_w2046_,
		_w2097_,
		_w10264_,
		_w10265_
	);
	LUT4 #(
		.INIT('h153f)
	) name8365 (
		\s14_data_i[11]_pad ,
		\s1_data_i[11]_pad ,
		_w9322_,
		_w9422_,
		_w10266_
	);
	LUT4 #(
		.INIT('h135f)
	) name8366 (
		\s10_data_i[11]_pad ,
		\s7_data_i[11]_pad ,
		_w9413_,
		_w9442_,
		_w10267_
	);
	LUT4 #(
		.INIT('h135f)
	) name8367 (
		\s2_data_i[11]_pad ,
		\s5_data_i[11]_pad ,
		_w9427_,
		_w9436_,
		_w10268_
	);
	LUT4 #(
		.INIT('h135f)
	) name8368 (
		\s0_data_i[11]_pad ,
		\s6_data_i[11]_pad ,
		_w9280_,
		_w9439_,
		_w10269_
	);
	LUT4 #(
		.INIT('h8000)
	) name8369 (
		_w10266_,
		_w10267_,
		_w10268_,
		_w10269_,
		_w10270_
	);
	LUT2 #(
		.INIT('h8)
	) name8370 (
		\s11_data_i[11]_pad ,
		_w9638_,
		_w10271_
	);
	LUT4 #(
		.INIT('h135f)
	) name8371 (
		\s4_data_i[11]_pad ,
		\s8_data_i[11]_pad ,
		_w9433_,
		_w9445_,
		_w10272_
	);
	LUT4 #(
		.INIT('h153f)
	) name8372 (
		\s12_data_i[11]_pad ,
		\s3_data_i[11]_pad ,
		_w9430_,
		_w9635_,
		_w10273_
	);
	LUT4 #(
		.INIT('h135f)
	) name8373 (
		\s13_data_i[11]_pad ,
		\s9_data_i[11]_pad ,
		_w9419_,
		_w9448_,
		_w10274_
	);
	LUT4 #(
		.INIT('h4000)
	) name8374 (
		_w10271_,
		_w10272_,
		_w10273_,
		_w10274_,
		_w10275_
	);
	LUT2 #(
		.INIT('h8)
	) name8375 (
		_w10270_,
		_w10275_,
		_w10276_
	);
	LUT3 #(
		.INIT('hef)
	) name8376 (
		_w10263_,
		_w10265_,
		_w10276_,
		_w10277_
	);
	LUT3 #(
		.INIT('h80)
	) name8377 (
		_w2047_,
		_w2097_,
		_w9731_,
		_w10278_
	);
	LUT2 #(
		.INIT('h8)
	) name8378 (
		\s15_data_i[12]_pad ,
		_w2047_,
		_w10279_
	);
	LUT3 #(
		.INIT('h70)
	) name8379 (
		_w2046_,
		_w2097_,
		_w10279_,
		_w10280_
	);
	LUT4 #(
		.INIT('h153f)
	) name8380 (
		\s12_data_i[12]_pad ,
		\s1_data_i[12]_pad ,
		_w9322_,
		_w9635_,
		_w10281_
	);
	LUT4 #(
		.INIT('h135f)
	) name8381 (
		\s0_data_i[12]_pad ,
		\s10_data_i[12]_pad ,
		_w9280_,
		_w9413_,
		_w10282_
	);
	LUT4 #(
		.INIT('h135f)
	) name8382 (
		\s3_data_i[12]_pad ,
		\s4_data_i[12]_pad ,
		_w9430_,
		_w9433_,
		_w10283_
	);
	LUT4 #(
		.INIT('h135f)
	) name8383 (
		\s6_data_i[12]_pad ,
		\s9_data_i[12]_pad ,
		_w9439_,
		_w9448_,
		_w10284_
	);
	LUT4 #(
		.INIT('h8000)
	) name8384 (
		_w10281_,
		_w10282_,
		_w10283_,
		_w10284_,
		_w10285_
	);
	LUT2 #(
		.INIT('h8)
	) name8385 (
		\s14_data_i[12]_pad ,
		_w9422_,
		_w10286_
	);
	LUT4 #(
		.INIT('h153f)
	) name8386 (
		\s11_data_i[12]_pad ,
		\s7_data_i[12]_pad ,
		_w9442_,
		_w9638_,
		_w10287_
	);
	LUT4 #(
		.INIT('h135f)
	) name8387 (
		\s5_data_i[12]_pad ,
		\s8_data_i[12]_pad ,
		_w9436_,
		_w9445_,
		_w10288_
	);
	LUT4 #(
		.INIT('h135f)
	) name8388 (
		\s13_data_i[12]_pad ,
		\s2_data_i[12]_pad ,
		_w9419_,
		_w9427_,
		_w10289_
	);
	LUT4 #(
		.INIT('h4000)
	) name8389 (
		_w10286_,
		_w10287_,
		_w10288_,
		_w10289_,
		_w10290_
	);
	LUT2 #(
		.INIT('h8)
	) name8390 (
		_w10285_,
		_w10290_,
		_w10291_
	);
	LUT3 #(
		.INIT('hef)
	) name8391 (
		_w10278_,
		_w10280_,
		_w10291_,
		_w10292_
	);
	LUT3 #(
		.INIT('h80)
	) name8392 (
		_w2047_,
		_w2097_,
		_w9747_,
		_w10293_
	);
	LUT2 #(
		.INIT('h8)
	) name8393 (
		\s15_data_i[13]_pad ,
		_w2047_,
		_w10294_
	);
	LUT3 #(
		.INIT('h70)
	) name8394 (
		_w2046_,
		_w2097_,
		_w10294_,
		_w10295_
	);
	LUT4 #(
		.INIT('h153f)
	) name8395 (
		\s12_data_i[13]_pad ,
		\s1_data_i[13]_pad ,
		_w9322_,
		_w9635_,
		_w10296_
	);
	LUT4 #(
		.INIT('h135f)
	) name8396 (
		\s0_data_i[13]_pad ,
		\s10_data_i[13]_pad ,
		_w9280_,
		_w9413_,
		_w10297_
	);
	LUT4 #(
		.INIT('h135f)
	) name8397 (
		\s3_data_i[13]_pad ,
		\s4_data_i[13]_pad ,
		_w9430_,
		_w9433_,
		_w10298_
	);
	LUT4 #(
		.INIT('h135f)
	) name8398 (
		\s6_data_i[13]_pad ,
		\s9_data_i[13]_pad ,
		_w9439_,
		_w9448_,
		_w10299_
	);
	LUT4 #(
		.INIT('h8000)
	) name8399 (
		_w10296_,
		_w10297_,
		_w10298_,
		_w10299_,
		_w10300_
	);
	LUT2 #(
		.INIT('h8)
	) name8400 (
		\s14_data_i[13]_pad ,
		_w9422_,
		_w10301_
	);
	LUT4 #(
		.INIT('h153f)
	) name8401 (
		\s11_data_i[13]_pad ,
		\s7_data_i[13]_pad ,
		_w9442_,
		_w9638_,
		_w10302_
	);
	LUT4 #(
		.INIT('h135f)
	) name8402 (
		\s5_data_i[13]_pad ,
		\s8_data_i[13]_pad ,
		_w9436_,
		_w9445_,
		_w10303_
	);
	LUT4 #(
		.INIT('h135f)
	) name8403 (
		\s13_data_i[13]_pad ,
		\s2_data_i[13]_pad ,
		_w9419_,
		_w9427_,
		_w10304_
	);
	LUT4 #(
		.INIT('h4000)
	) name8404 (
		_w10301_,
		_w10302_,
		_w10303_,
		_w10304_,
		_w10305_
	);
	LUT2 #(
		.INIT('h8)
	) name8405 (
		_w10300_,
		_w10305_,
		_w10306_
	);
	LUT3 #(
		.INIT('hef)
	) name8406 (
		_w10293_,
		_w10295_,
		_w10306_,
		_w10307_
	);
	LUT3 #(
		.INIT('h80)
	) name8407 (
		_w2047_,
		_w2097_,
		_w9763_,
		_w10308_
	);
	LUT2 #(
		.INIT('h8)
	) name8408 (
		\s15_data_i[14]_pad ,
		_w2047_,
		_w10309_
	);
	LUT3 #(
		.INIT('h70)
	) name8409 (
		_w2046_,
		_w2097_,
		_w10309_,
		_w10310_
	);
	LUT4 #(
		.INIT('h153f)
	) name8410 (
		\s12_data_i[14]_pad ,
		\s1_data_i[14]_pad ,
		_w9322_,
		_w9635_,
		_w10311_
	);
	LUT4 #(
		.INIT('h135f)
	) name8411 (
		\s0_data_i[14]_pad ,
		\s10_data_i[14]_pad ,
		_w9280_,
		_w9413_,
		_w10312_
	);
	LUT4 #(
		.INIT('h135f)
	) name8412 (
		\s3_data_i[14]_pad ,
		\s4_data_i[14]_pad ,
		_w9430_,
		_w9433_,
		_w10313_
	);
	LUT4 #(
		.INIT('h135f)
	) name8413 (
		\s6_data_i[14]_pad ,
		\s9_data_i[14]_pad ,
		_w9439_,
		_w9448_,
		_w10314_
	);
	LUT4 #(
		.INIT('h8000)
	) name8414 (
		_w10311_,
		_w10312_,
		_w10313_,
		_w10314_,
		_w10315_
	);
	LUT2 #(
		.INIT('h8)
	) name8415 (
		\s14_data_i[14]_pad ,
		_w9422_,
		_w10316_
	);
	LUT4 #(
		.INIT('h153f)
	) name8416 (
		\s11_data_i[14]_pad ,
		\s7_data_i[14]_pad ,
		_w9442_,
		_w9638_,
		_w10317_
	);
	LUT4 #(
		.INIT('h135f)
	) name8417 (
		\s5_data_i[14]_pad ,
		\s8_data_i[14]_pad ,
		_w9436_,
		_w9445_,
		_w10318_
	);
	LUT4 #(
		.INIT('h135f)
	) name8418 (
		\s13_data_i[14]_pad ,
		\s2_data_i[14]_pad ,
		_w9419_,
		_w9427_,
		_w10319_
	);
	LUT4 #(
		.INIT('h4000)
	) name8419 (
		_w10316_,
		_w10317_,
		_w10318_,
		_w10319_,
		_w10320_
	);
	LUT2 #(
		.INIT('h8)
	) name8420 (
		_w10315_,
		_w10320_,
		_w10321_
	);
	LUT3 #(
		.INIT('hef)
	) name8421 (
		_w10308_,
		_w10310_,
		_w10321_,
		_w10322_
	);
	LUT3 #(
		.INIT('h80)
	) name8422 (
		_w2047_,
		_w2097_,
		_w9779_,
		_w10323_
	);
	LUT2 #(
		.INIT('h8)
	) name8423 (
		\s15_data_i[15]_pad ,
		_w2047_,
		_w10324_
	);
	LUT3 #(
		.INIT('h70)
	) name8424 (
		_w2046_,
		_w2097_,
		_w10324_,
		_w10325_
	);
	LUT4 #(
		.INIT('h153f)
	) name8425 (
		\s12_data_i[15]_pad ,
		\s1_data_i[15]_pad ,
		_w9322_,
		_w9635_,
		_w10326_
	);
	LUT4 #(
		.INIT('h135f)
	) name8426 (
		\s0_data_i[15]_pad ,
		\s10_data_i[15]_pad ,
		_w9280_,
		_w9413_,
		_w10327_
	);
	LUT4 #(
		.INIT('h135f)
	) name8427 (
		\s3_data_i[15]_pad ,
		\s4_data_i[15]_pad ,
		_w9430_,
		_w9433_,
		_w10328_
	);
	LUT4 #(
		.INIT('h135f)
	) name8428 (
		\s6_data_i[15]_pad ,
		\s9_data_i[15]_pad ,
		_w9439_,
		_w9448_,
		_w10329_
	);
	LUT4 #(
		.INIT('h8000)
	) name8429 (
		_w10326_,
		_w10327_,
		_w10328_,
		_w10329_,
		_w10330_
	);
	LUT2 #(
		.INIT('h8)
	) name8430 (
		\s14_data_i[15]_pad ,
		_w9422_,
		_w10331_
	);
	LUT4 #(
		.INIT('h153f)
	) name8431 (
		\s11_data_i[15]_pad ,
		\s7_data_i[15]_pad ,
		_w9442_,
		_w9638_,
		_w10332_
	);
	LUT4 #(
		.INIT('h135f)
	) name8432 (
		\s5_data_i[15]_pad ,
		\s8_data_i[15]_pad ,
		_w9436_,
		_w9445_,
		_w10333_
	);
	LUT4 #(
		.INIT('h135f)
	) name8433 (
		\s13_data_i[15]_pad ,
		\s2_data_i[15]_pad ,
		_w9419_,
		_w9427_,
		_w10334_
	);
	LUT4 #(
		.INIT('h4000)
	) name8434 (
		_w10331_,
		_w10332_,
		_w10333_,
		_w10334_,
		_w10335_
	);
	LUT2 #(
		.INIT('h8)
	) name8435 (
		_w10330_,
		_w10335_,
		_w10336_
	);
	LUT3 #(
		.INIT('hef)
	) name8436 (
		_w10323_,
		_w10325_,
		_w10336_,
		_w10337_
	);
	LUT2 #(
		.INIT('h8)
	) name8437 (
		\s15_data_i[16]_pad ,
		_w2047_,
		_w10338_
	);
	LUT4 #(
		.INIT('h135f)
	) name8438 (
		\s1_data_i[16]_pad ,
		\s8_data_i[16]_pad ,
		_w9322_,
		_w9445_,
		_w10339_
	);
	LUT4 #(
		.INIT('h135f)
	) name8439 (
		\s0_data_i[16]_pad ,
		\s7_data_i[16]_pad ,
		_w9280_,
		_w9442_,
		_w10340_
	);
	LUT4 #(
		.INIT('h135f)
	) name8440 (
		\s3_data_i[16]_pad ,
		\s9_data_i[16]_pad ,
		_w9430_,
		_w9448_,
		_w10341_
	);
	LUT4 #(
		.INIT('h135f)
	) name8441 (
		\s10_data_i[16]_pad ,
		\s4_data_i[16]_pad ,
		_w9413_,
		_w9433_,
		_w10342_
	);
	LUT4 #(
		.INIT('h8000)
	) name8442 (
		_w10339_,
		_w10340_,
		_w10341_,
		_w10342_,
		_w10343_
	);
	LUT2 #(
		.INIT('h8)
	) name8443 (
		\s11_data_i[16]_pad ,
		_w9638_,
		_w10344_
	);
	LUT4 #(
		.INIT('h135f)
	) name8444 (
		\s14_data_i[16]_pad ,
		\s2_data_i[16]_pad ,
		_w9422_,
		_w9427_,
		_w10345_
	);
	LUT4 #(
		.INIT('h153f)
	) name8445 (
		\s12_data_i[16]_pad ,
		\s5_data_i[16]_pad ,
		_w9436_,
		_w9635_,
		_w10346_
	);
	LUT4 #(
		.INIT('h135f)
	) name8446 (
		\s13_data_i[16]_pad ,
		\s6_data_i[16]_pad ,
		_w9419_,
		_w9439_,
		_w10347_
	);
	LUT4 #(
		.INIT('h4000)
	) name8447 (
		_w10344_,
		_w10345_,
		_w10346_,
		_w10347_,
		_w10348_
	);
	LUT2 #(
		.INIT('h8)
	) name8448 (
		_w10343_,
		_w10348_,
		_w10349_
	);
	LUT4 #(
		.INIT('h70ff)
	) name8449 (
		_w2046_,
		_w2097_,
		_w10338_,
		_w10349_,
		_w10350_
	);
	LUT2 #(
		.INIT('h8)
	) name8450 (
		\s15_data_i[17]_pad ,
		_w2047_,
		_w10351_
	);
	LUT4 #(
		.INIT('h135f)
	) name8451 (
		\s1_data_i[17]_pad ,
		\s8_data_i[17]_pad ,
		_w9322_,
		_w9445_,
		_w10352_
	);
	LUT4 #(
		.INIT('h135f)
	) name8452 (
		\s4_data_i[17]_pad ,
		\s6_data_i[17]_pad ,
		_w9433_,
		_w9439_,
		_w10353_
	);
	LUT4 #(
		.INIT('h135f)
	) name8453 (
		\s3_data_i[17]_pad ,
		\s9_data_i[17]_pad ,
		_w9430_,
		_w9448_,
		_w10354_
	);
	LUT4 #(
		.INIT('h135f)
	) name8454 (
		\s10_data_i[17]_pad ,
		\s7_data_i[17]_pad ,
		_w9413_,
		_w9442_,
		_w10355_
	);
	LUT4 #(
		.INIT('h8000)
	) name8455 (
		_w10352_,
		_w10353_,
		_w10354_,
		_w10355_,
		_w10356_
	);
	LUT2 #(
		.INIT('h8)
	) name8456 (
		\s11_data_i[17]_pad ,
		_w9638_,
		_w10357_
	);
	LUT4 #(
		.INIT('h135f)
	) name8457 (
		\s14_data_i[17]_pad ,
		\s2_data_i[17]_pad ,
		_w9422_,
		_w9427_,
		_w10358_
	);
	LUT4 #(
		.INIT('h153f)
	) name8458 (
		\s12_data_i[17]_pad ,
		\s5_data_i[17]_pad ,
		_w9436_,
		_w9635_,
		_w10359_
	);
	LUT4 #(
		.INIT('h135f)
	) name8459 (
		\s0_data_i[17]_pad ,
		\s13_data_i[17]_pad ,
		_w9280_,
		_w9419_,
		_w10360_
	);
	LUT4 #(
		.INIT('h4000)
	) name8460 (
		_w10357_,
		_w10358_,
		_w10359_,
		_w10360_,
		_w10361_
	);
	LUT2 #(
		.INIT('h8)
	) name8461 (
		_w10356_,
		_w10361_,
		_w10362_
	);
	LUT4 #(
		.INIT('h70ff)
	) name8462 (
		_w2046_,
		_w2097_,
		_w10351_,
		_w10362_,
		_w10363_
	);
	LUT2 #(
		.INIT('h8)
	) name8463 (
		\s15_data_i[18]_pad ,
		_w2047_,
		_w10364_
	);
	LUT4 #(
		.INIT('h135f)
	) name8464 (
		\s1_data_i[18]_pad ,
		\s8_data_i[18]_pad ,
		_w9322_,
		_w9445_,
		_w10365_
	);
	LUT4 #(
		.INIT('h135f)
	) name8465 (
		\s0_data_i[18]_pad ,
		\s7_data_i[18]_pad ,
		_w9280_,
		_w9442_,
		_w10366_
	);
	LUT4 #(
		.INIT('h135f)
	) name8466 (
		\s3_data_i[18]_pad ,
		\s9_data_i[18]_pad ,
		_w9430_,
		_w9448_,
		_w10367_
	);
	LUT4 #(
		.INIT('h135f)
	) name8467 (
		\s10_data_i[18]_pad ,
		\s4_data_i[18]_pad ,
		_w9413_,
		_w9433_,
		_w10368_
	);
	LUT4 #(
		.INIT('h8000)
	) name8468 (
		_w10365_,
		_w10366_,
		_w10367_,
		_w10368_,
		_w10369_
	);
	LUT2 #(
		.INIT('h8)
	) name8469 (
		\s11_data_i[18]_pad ,
		_w9638_,
		_w10370_
	);
	LUT4 #(
		.INIT('h135f)
	) name8470 (
		\s14_data_i[18]_pad ,
		\s2_data_i[18]_pad ,
		_w9422_,
		_w9427_,
		_w10371_
	);
	LUT4 #(
		.INIT('h153f)
	) name8471 (
		\s12_data_i[18]_pad ,
		\s5_data_i[18]_pad ,
		_w9436_,
		_w9635_,
		_w10372_
	);
	LUT4 #(
		.INIT('h135f)
	) name8472 (
		\s13_data_i[18]_pad ,
		\s6_data_i[18]_pad ,
		_w9419_,
		_w9439_,
		_w10373_
	);
	LUT4 #(
		.INIT('h4000)
	) name8473 (
		_w10370_,
		_w10371_,
		_w10372_,
		_w10373_,
		_w10374_
	);
	LUT2 #(
		.INIT('h8)
	) name8474 (
		_w10369_,
		_w10374_,
		_w10375_
	);
	LUT4 #(
		.INIT('h70ff)
	) name8475 (
		_w2046_,
		_w2097_,
		_w10364_,
		_w10375_,
		_w10376_
	);
	LUT2 #(
		.INIT('h8)
	) name8476 (
		\s15_data_i[19]_pad ,
		_w2047_,
		_w10377_
	);
	LUT4 #(
		.INIT('h135f)
	) name8477 (
		\s1_data_i[19]_pad ,
		\s8_data_i[19]_pad ,
		_w9322_,
		_w9445_,
		_w10378_
	);
	LUT4 #(
		.INIT('h135f)
	) name8478 (
		\s4_data_i[19]_pad ,
		\s6_data_i[19]_pad ,
		_w9433_,
		_w9439_,
		_w10379_
	);
	LUT4 #(
		.INIT('h135f)
	) name8479 (
		\s3_data_i[19]_pad ,
		\s9_data_i[19]_pad ,
		_w9430_,
		_w9448_,
		_w10380_
	);
	LUT4 #(
		.INIT('h135f)
	) name8480 (
		\s10_data_i[19]_pad ,
		\s7_data_i[19]_pad ,
		_w9413_,
		_w9442_,
		_w10381_
	);
	LUT4 #(
		.INIT('h8000)
	) name8481 (
		_w10378_,
		_w10379_,
		_w10380_,
		_w10381_,
		_w10382_
	);
	LUT2 #(
		.INIT('h8)
	) name8482 (
		\s11_data_i[19]_pad ,
		_w9638_,
		_w10383_
	);
	LUT4 #(
		.INIT('h135f)
	) name8483 (
		\s14_data_i[19]_pad ,
		\s2_data_i[19]_pad ,
		_w9422_,
		_w9427_,
		_w10384_
	);
	LUT4 #(
		.INIT('h153f)
	) name8484 (
		\s12_data_i[19]_pad ,
		\s5_data_i[19]_pad ,
		_w9436_,
		_w9635_,
		_w10385_
	);
	LUT4 #(
		.INIT('h135f)
	) name8485 (
		\s0_data_i[19]_pad ,
		\s13_data_i[19]_pad ,
		_w9280_,
		_w9419_,
		_w10386_
	);
	LUT4 #(
		.INIT('h4000)
	) name8486 (
		_w10383_,
		_w10384_,
		_w10385_,
		_w10386_,
		_w10387_
	);
	LUT2 #(
		.INIT('h8)
	) name8487 (
		_w10382_,
		_w10387_,
		_w10388_
	);
	LUT4 #(
		.INIT('h70ff)
	) name8488 (
		_w2046_,
		_w2097_,
		_w10377_,
		_w10388_,
		_w10389_
	);
	LUT3 #(
		.INIT('h80)
	) name8489 (
		_w2047_,
		_w2097_,
		_w9847_,
		_w10390_
	);
	LUT2 #(
		.INIT('h8)
	) name8490 (
		\s15_data_i[1]_pad ,
		_w2047_,
		_w10391_
	);
	LUT3 #(
		.INIT('h70)
	) name8491 (
		_w2046_,
		_w2097_,
		_w10391_,
		_w10392_
	);
	LUT4 #(
		.INIT('h153f)
	) name8492 (
		\s12_data_i[1]_pad ,
		\s1_data_i[1]_pad ,
		_w9322_,
		_w9635_,
		_w10393_
	);
	LUT4 #(
		.INIT('h135f)
	) name8493 (
		\s0_data_i[1]_pad ,
		\s10_data_i[1]_pad ,
		_w9280_,
		_w9413_,
		_w10394_
	);
	LUT4 #(
		.INIT('h135f)
	) name8494 (
		\s3_data_i[1]_pad ,
		\s4_data_i[1]_pad ,
		_w9430_,
		_w9433_,
		_w10395_
	);
	LUT4 #(
		.INIT('h135f)
	) name8495 (
		\s6_data_i[1]_pad ,
		\s9_data_i[1]_pad ,
		_w9439_,
		_w9448_,
		_w10396_
	);
	LUT4 #(
		.INIT('h8000)
	) name8496 (
		_w10393_,
		_w10394_,
		_w10395_,
		_w10396_,
		_w10397_
	);
	LUT2 #(
		.INIT('h8)
	) name8497 (
		\s14_data_i[1]_pad ,
		_w9422_,
		_w10398_
	);
	LUT4 #(
		.INIT('h153f)
	) name8498 (
		\s11_data_i[1]_pad ,
		\s7_data_i[1]_pad ,
		_w9442_,
		_w9638_,
		_w10399_
	);
	LUT4 #(
		.INIT('h135f)
	) name8499 (
		\s5_data_i[1]_pad ,
		\s8_data_i[1]_pad ,
		_w9436_,
		_w9445_,
		_w10400_
	);
	LUT4 #(
		.INIT('h135f)
	) name8500 (
		\s13_data_i[1]_pad ,
		\s2_data_i[1]_pad ,
		_w9419_,
		_w9427_,
		_w10401_
	);
	LUT4 #(
		.INIT('h4000)
	) name8501 (
		_w10398_,
		_w10399_,
		_w10400_,
		_w10401_,
		_w10402_
	);
	LUT2 #(
		.INIT('h8)
	) name8502 (
		_w10397_,
		_w10402_,
		_w10403_
	);
	LUT3 #(
		.INIT('hef)
	) name8503 (
		_w10390_,
		_w10392_,
		_w10403_,
		_w10404_
	);
	LUT2 #(
		.INIT('h8)
	) name8504 (
		\s15_data_i[20]_pad ,
		_w2047_,
		_w10405_
	);
	LUT4 #(
		.INIT('h135f)
	) name8505 (
		\s1_data_i[20]_pad ,
		\s8_data_i[20]_pad ,
		_w9322_,
		_w9445_,
		_w10406_
	);
	LUT4 #(
		.INIT('h135f)
	) name8506 (
		\s4_data_i[20]_pad ,
		\s6_data_i[20]_pad ,
		_w9433_,
		_w9439_,
		_w10407_
	);
	LUT4 #(
		.INIT('h135f)
	) name8507 (
		\s3_data_i[20]_pad ,
		\s9_data_i[20]_pad ,
		_w9430_,
		_w9448_,
		_w10408_
	);
	LUT4 #(
		.INIT('h135f)
	) name8508 (
		\s10_data_i[20]_pad ,
		\s7_data_i[20]_pad ,
		_w9413_,
		_w9442_,
		_w10409_
	);
	LUT4 #(
		.INIT('h8000)
	) name8509 (
		_w10406_,
		_w10407_,
		_w10408_,
		_w10409_,
		_w10410_
	);
	LUT2 #(
		.INIT('h8)
	) name8510 (
		\s11_data_i[20]_pad ,
		_w9638_,
		_w10411_
	);
	LUT4 #(
		.INIT('h135f)
	) name8511 (
		\s14_data_i[20]_pad ,
		\s2_data_i[20]_pad ,
		_w9422_,
		_w9427_,
		_w10412_
	);
	LUT4 #(
		.INIT('h153f)
	) name8512 (
		\s12_data_i[20]_pad ,
		\s5_data_i[20]_pad ,
		_w9436_,
		_w9635_,
		_w10413_
	);
	LUT4 #(
		.INIT('h135f)
	) name8513 (
		\s0_data_i[20]_pad ,
		\s13_data_i[20]_pad ,
		_w9280_,
		_w9419_,
		_w10414_
	);
	LUT4 #(
		.INIT('h4000)
	) name8514 (
		_w10411_,
		_w10412_,
		_w10413_,
		_w10414_,
		_w10415_
	);
	LUT2 #(
		.INIT('h8)
	) name8515 (
		_w10410_,
		_w10415_,
		_w10416_
	);
	LUT4 #(
		.INIT('h70ff)
	) name8516 (
		_w2046_,
		_w2097_,
		_w10405_,
		_w10416_,
		_w10417_
	);
	LUT2 #(
		.INIT('h8)
	) name8517 (
		\s15_data_i[21]_pad ,
		_w2047_,
		_w10418_
	);
	LUT4 #(
		.INIT('h135f)
	) name8518 (
		\s1_data_i[21]_pad ,
		\s8_data_i[21]_pad ,
		_w9322_,
		_w9445_,
		_w10419_
	);
	LUT4 #(
		.INIT('h135f)
	) name8519 (
		\s4_data_i[21]_pad ,
		\s6_data_i[21]_pad ,
		_w9433_,
		_w9439_,
		_w10420_
	);
	LUT4 #(
		.INIT('h135f)
	) name8520 (
		\s3_data_i[21]_pad ,
		\s9_data_i[21]_pad ,
		_w9430_,
		_w9448_,
		_w10421_
	);
	LUT4 #(
		.INIT('h135f)
	) name8521 (
		\s10_data_i[21]_pad ,
		\s7_data_i[21]_pad ,
		_w9413_,
		_w9442_,
		_w10422_
	);
	LUT4 #(
		.INIT('h8000)
	) name8522 (
		_w10419_,
		_w10420_,
		_w10421_,
		_w10422_,
		_w10423_
	);
	LUT2 #(
		.INIT('h8)
	) name8523 (
		\s11_data_i[21]_pad ,
		_w9638_,
		_w10424_
	);
	LUT4 #(
		.INIT('h135f)
	) name8524 (
		\s14_data_i[21]_pad ,
		\s2_data_i[21]_pad ,
		_w9422_,
		_w9427_,
		_w10425_
	);
	LUT4 #(
		.INIT('h153f)
	) name8525 (
		\s12_data_i[21]_pad ,
		\s5_data_i[21]_pad ,
		_w9436_,
		_w9635_,
		_w10426_
	);
	LUT4 #(
		.INIT('h135f)
	) name8526 (
		\s0_data_i[21]_pad ,
		\s13_data_i[21]_pad ,
		_w9280_,
		_w9419_,
		_w10427_
	);
	LUT4 #(
		.INIT('h4000)
	) name8527 (
		_w10424_,
		_w10425_,
		_w10426_,
		_w10427_,
		_w10428_
	);
	LUT2 #(
		.INIT('h8)
	) name8528 (
		_w10423_,
		_w10428_,
		_w10429_
	);
	LUT4 #(
		.INIT('h70ff)
	) name8529 (
		_w2046_,
		_w2097_,
		_w10418_,
		_w10429_,
		_w10430_
	);
	LUT2 #(
		.INIT('h8)
	) name8530 (
		\s15_data_i[22]_pad ,
		_w2047_,
		_w10431_
	);
	LUT4 #(
		.INIT('h135f)
	) name8531 (
		\s1_data_i[22]_pad ,
		\s8_data_i[22]_pad ,
		_w9322_,
		_w9445_,
		_w10432_
	);
	LUT4 #(
		.INIT('h135f)
	) name8532 (
		\s4_data_i[22]_pad ,
		\s6_data_i[22]_pad ,
		_w9433_,
		_w9439_,
		_w10433_
	);
	LUT4 #(
		.INIT('h135f)
	) name8533 (
		\s3_data_i[22]_pad ,
		\s9_data_i[22]_pad ,
		_w9430_,
		_w9448_,
		_w10434_
	);
	LUT4 #(
		.INIT('h135f)
	) name8534 (
		\s10_data_i[22]_pad ,
		\s7_data_i[22]_pad ,
		_w9413_,
		_w9442_,
		_w10435_
	);
	LUT4 #(
		.INIT('h8000)
	) name8535 (
		_w10432_,
		_w10433_,
		_w10434_,
		_w10435_,
		_w10436_
	);
	LUT2 #(
		.INIT('h8)
	) name8536 (
		\s11_data_i[22]_pad ,
		_w9638_,
		_w10437_
	);
	LUT4 #(
		.INIT('h135f)
	) name8537 (
		\s14_data_i[22]_pad ,
		\s2_data_i[22]_pad ,
		_w9422_,
		_w9427_,
		_w10438_
	);
	LUT4 #(
		.INIT('h153f)
	) name8538 (
		\s12_data_i[22]_pad ,
		\s5_data_i[22]_pad ,
		_w9436_,
		_w9635_,
		_w10439_
	);
	LUT4 #(
		.INIT('h135f)
	) name8539 (
		\s0_data_i[22]_pad ,
		\s13_data_i[22]_pad ,
		_w9280_,
		_w9419_,
		_w10440_
	);
	LUT4 #(
		.INIT('h4000)
	) name8540 (
		_w10437_,
		_w10438_,
		_w10439_,
		_w10440_,
		_w10441_
	);
	LUT2 #(
		.INIT('h8)
	) name8541 (
		_w10436_,
		_w10441_,
		_w10442_
	);
	LUT4 #(
		.INIT('h70ff)
	) name8542 (
		_w2046_,
		_w2097_,
		_w10431_,
		_w10442_,
		_w10443_
	);
	LUT2 #(
		.INIT('h8)
	) name8543 (
		\s15_data_i[23]_pad ,
		_w2047_,
		_w10444_
	);
	LUT4 #(
		.INIT('h153f)
	) name8544 (
		\s12_data_i[23]_pad ,
		\s1_data_i[23]_pad ,
		_w9322_,
		_w9635_,
		_w10445_
	);
	LUT4 #(
		.INIT('h135f)
	) name8545 (
		\s4_data_i[23]_pad ,
		\s6_data_i[23]_pad ,
		_w9433_,
		_w9439_,
		_w10446_
	);
	LUT4 #(
		.INIT('h135f)
	) name8546 (
		\s3_data_i[23]_pad ,
		\s9_data_i[23]_pad ,
		_w9430_,
		_w9448_,
		_w10447_
	);
	LUT4 #(
		.INIT('h135f)
	) name8547 (
		\s10_data_i[23]_pad ,
		\s7_data_i[23]_pad ,
		_w9413_,
		_w9442_,
		_w10448_
	);
	LUT4 #(
		.INIT('h8000)
	) name8548 (
		_w10445_,
		_w10446_,
		_w10447_,
		_w10448_,
		_w10449_
	);
	LUT2 #(
		.INIT('h8)
	) name8549 (
		\s14_data_i[23]_pad ,
		_w9422_,
		_w10450_
	);
	LUT4 #(
		.INIT('h153f)
	) name8550 (
		\s11_data_i[23]_pad ,
		\s2_data_i[23]_pad ,
		_w9427_,
		_w9638_,
		_w10451_
	);
	LUT4 #(
		.INIT('h135f)
	) name8551 (
		\s5_data_i[23]_pad ,
		\s8_data_i[23]_pad ,
		_w9436_,
		_w9445_,
		_w10452_
	);
	LUT4 #(
		.INIT('h135f)
	) name8552 (
		\s0_data_i[23]_pad ,
		\s13_data_i[23]_pad ,
		_w9280_,
		_w9419_,
		_w10453_
	);
	LUT4 #(
		.INIT('h4000)
	) name8553 (
		_w10450_,
		_w10451_,
		_w10452_,
		_w10453_,
		_w10454_
	);
	LUT2 #(
		.INIT('h8)
	) name8554 (
		_w10449_,
		_w10454_,
		_w10455_
	);
	LUT4 #(
		.INIT('h70ff)
	) name8555 (
		_w2046_,
		_w2097_,
		_w10444_,
		_w10455_,
		_w10456_
	);
	LUT2 #(
		.INIT('h8)
	) name8556 (
		\s15_data_i[24]_pad ,
		_w2047_,
		_w10457_
	);
	LUT4 #(
		.INIT('h135f)
	) name8557 (
		\s1_data_i[24]_pad ,
		\s8_data_i[24]_pad ,
		_w9322_,
		_w9445_,
		_w10458_
	);
	LUT4 #(
		.INIT('h135f)
	) name8558 (
		\s4_data_i[24]_pad ,
		\s6_data_i[24]_pad ,
		_w9433_,
		_w9439_,
		_w10459_
	);
	LUT4 #(
		.INIT('h135f)
	) name8559 (
		\s3_data_i[24]_pad ,
		\s9_data_i[24]_pad ,
		_w9430_,
		_w9448_,
		_w10460_
	);
	LUT4 #(
		.INIT('h135f)
	) name8560 (
		\s10_data_i[24]_pad ,
		\s7_data_i[24]_pad ,
		_w9413_,
		_w9442_,
		_w10461_
	);
	LUT4 #(
		.INIT('h8000)
	) name8561 (
		_w10458_,
		_w10459_,
		_w10460_,
		_w10461_,
		_w10462_
	);
	LUT2 #(
		.INIT('h8)
	) name8562 (
		\s11_data_i[24]_pad ,
		_w9638_,
		_w10463_
	);
	LUT4 #(
		.INIT('h135f)
	) name8563 (
		\s14_data_i[24]_pad ,
		\s2_data_i[24]_pad ,
		_w9422_,
		_w9427_,
		_w10464_
	);
	LUT4 #(
		.INIT('h153f)
	) name8564 (
		\s12_data_i[24]_pad ,
		\s5_data_i[24]_pad ,
		_w9436_,
		_w9635_,
		_w10465_
	);
	LUT4 #(
		.INIT('h135f)
	) name8565 (
		\s0_data_i[24]_pad ,
		\s13_data_i[24]_pad ,
		_w9280_,
		_w9419_,
		_w10466_
	);
	LUT4 #(
		.INIT('h4000)
	) name8566 (
		_w10463_,
		_w10464_,
		_w10465_,
		_w10466_,
		_w10467_
	);
	LUT2 #(
		.INIT('h8)
	) name8567 (
		_w10462_,
		_w10467_,
		_w10468_
	);
	LUT4 #(
		.INIT('h70ff)
	) name8568 (
		_w2046_,
		_w2097_,
		_w10457_,
		_w10468_,
		_w10469_
	);
	LUT2 #(
		.INIT('h8)
	) name8569 (
		\s15_data_i[25]_pad ,
		_w2047_,
		_w10470_
	);
	LUT4 #(
		.INIT('h135f)
	) name8570 (
		\s1_data_i[25]_pad ,
		\s8_data_i[25]_pad ,
		_w9322_,
		_w9445_,
		_w10471_
	);
	LUT4 #(
		.INIT('h135f)
	) name8571 (
		\s4_data_i[25]_pad ,
		\s6_data_i[25]_pad ,
		_w9433_,
		_w9439_,
		_w10472_
	);
	LUT4 #(
		.INIT('h135f)
	) name8572 (
		\s3_data_i[25]_pad ,
		\s9_data_i[25]_pad ,
		_w9430_,
		_w9448_,
		_w10473_
	);
	LUT4 #(
		.INIT('h135f)
	) name8573 (
		\s10_data_i[25]_pad ,
		\s7_data_i[25]_pad ,
		_w9413_,
		_w9442_,
		_w10474_
	);
	LUT4 #(
		.INIT('h8000)
	) name8574 (
		_w10471_,
		_w10472_,
		_w10473_,
		_w10474_,
		_w10475_
	);
	LUT2 #(
		.INIT('h8)
	) name8575 (
		\s11_data_i[25]_pad ,
		_w9638_,
		_w10476_
	);
	LUT4 #(
		.INIT('h135f)
	) name8576 (
		\s14_data_i[25]_pad ,
		\s2_data_i[25]_pad ,
		_w9422_,
		_w9427_,
		_w10477_
	);
	LUT4 #(
		.INIT('h153f)
	) name8577 (
		\s12_data_i[25]_pad ,
		\s5_data_i[25]_pad ,
		_w9436_,
		_w9635_,
		_w10478_
	);
	LUT4 #(
		.INIT('h135f)
	) name8578 (
		\s0_data_i[25]_pad ,
		\s13_data_i[25]_pad ,
		_w9280_,
		_w9419_,
		_w10479_
	);
	LUT4 #(
		.INIT('h4000)
	) name8579 (
		_w10476_,
		_w10477_,
		_w10478_,
		_w10479_,
		_w10480_
	);
	LUT2 #(
		.INIT('h8)
	) name8580 (
		_w10475_,
		_w10480_,
		_w10481_
	);
	LUT4 #(
		.INIT('h70ff)
	) name8581 (
		_w2046_,
		_w2097_,
		_w10470_,
		_w10481_,
		_w10482_
	);
	LUT2 #(
		.INIT('h8)
	) name8582 (
		\s15_data_i[26]_pad ,
		_w2047_,
		_w10483_
	);
	LUT4 #(
		.INIT('h135f)
	) name8583 (
		\s1_data_i[26]_pad ,
		\s8_data_i[26]_pad ,
		_w9322_,
		_w9445_,
		_w10484_
	);
	LUT4 #(
		.INIT('h135f)
	) name8584 (
		\s4_data_i[26]_pad ,
		\s6_data_i[26]_pad ,
		_w9433_,
		_w9439_,
		_w10485_
	);
	LUT4 #(
		.INIT('h135f)
	) name8585 (
		\s3_data_i[26]_pad ,
		\s9_data_i[26]_pad ,
		_w9430_,
		_w9448_,
		_w10486_
	);
	LUT4 #(
		.INIT('h135f)
	) name8586 (
		\s10_data_i[26]_pad ,
		\s7_data_i[26]_pad ,
		_w9413_,
		_w9442_,
		_w10487_
	);
	LUT4 #(
		.INIT('h8000)
	) name8587 (
		_w10484_,
		_w10485_,
		_w10486_,
		_w10487_,
		_w10488_
	);
	LUT2 #(
		.INIT('h8)
	) name8588 (
		\s11_data_i[26]_pad ,
		_w9638_,
		_w10489_
	);
	LUT4 #(
		.INIT('h135f)
	) name8589 (
		\s14_data_i[26]_pad ,
		\s2_data_i[26]_pad ,
		_w9422_,
		_w9427_,
		_w10490_
	);
	LUT4 #(
		.INIT('h153f)
	) name8590 (
		\s12_data_i[26]_pad ,
		\s5_data_i[26]_pad ,
		_w9436_,
		_w9635_,
		_w10491_
	);
	LUT4 #(
		.INIT('h135f)
	) name8591 (
		\s0_data_i[26]_pad ,
		\s13_data_i[26]_pad ,
		_w9280_,
		_w9419_,
		_w10492_
	);
	LUT4 #(
		.INIT('h4000)
	) name8592 (
		_w10489_,
		_w10490_,
		_w10491_,
		_w10492_,
		_w10493_
	);
	LUT2 #(
		.INIT('h8)
	) name8593 (
		_w10488_,
		_w10493_,
		_w10494_
	);
	LUT4 #(
		.INIT('h70ff)
	) name8594 (
		_w2046_,
		_w2097_,
		_w10483_,
		_w10494_,
		_w10495_
	);
	LUT2 #(
		.INIT('h8)
	) name8595 (
		\s15_data_i[27]_pad ,
		_w2047_,
		_w10496_
	);
	LUT4 #(
		.INIT('h135f)
	) name8596 (
		\s1_data_i[27]_pad ,
		\s8_data_i[27]_pad ,
		_w9322_,
		_w9445_,
		_w10497_
	);
	LUT4 #(
		.INIT('h135f)
	) name8597 (
		\s4_data_i[27]_pad ,
		\s6_data_i[27]_pad ,
		_w9433_,
		_w9439_,
		_w10498_
	);
	LUT4 #(
		.INIT('h135f)
	) name8598 (
		\s3_data_i[27]_pad ,
		\s9_data_i[27]_pad ,
		_w9430_,
		_w9448_,
		_w10499_
	);
	LUT4 #(
		.INIT('h135f)
	) name8599 (
		\s10_data_i[27]_pad ,
		\s7_data_i[27]_pad ,
		_w9413_,
		_w9442_,
		_w10500_
	);
	LUT4 #(
		.INIT('h8000)
	) name8600 (
		_w10497_,
		_w10498_,
		_w10499_,
		_w10500_,
		_w10501_
	);
	LUT2 #(
		.INIT('h8)
	) name8601 (
		\s11_data_i[27]_pad ,
		_w9638_,
		_w10502_
	);
	LUT4 #(
		.INIT('h135f)
	) name8602 (
		\s14_data_i[27]_pad ,
		\s2_data_i[27]_pad ,
		_w9422_,
		_w9427_,
		_w10503_
	);
	LUT4 #(
		.INIT('h153f)
	) name8603 (
		\s12_data_i[27]_pad ,
		\s5_data_i[27]_pad ,
		_w9436_,
		_w9635_,
		_w10504_
	);
	LUT4 #(
		.INIT('h135f)
	) name8604 (
		\s0_data_i[27]_pad ,
		\s13_data_i[27]_pad ,
		_w9280_,
		_w9419_,
		_w10505_
	);
	LUT4 #(
		.INIT('h4000)
	) name8605 (
		_w10502_,
		_w10503_,
		_w10504_,
		_w10505_,
		_w10506_
	);
	LUT2 #(
		.INIT('h8)
	) name8606 (
		_w10501_,
		_w10506_,
		_w10507_
	);
	LUT4 #(
		.INIT('h70ff)
	) name8607 (
		_w2046_,
		_w2097_,
		_w10496_,
		_w10507_,
		_w10508_
	);
	LUT2 #(
		.INIT('h8)
	) name8608 (
		\s15_data_i[28]_pad ,
		_w2047_,
		_w10509_
	);
	LUT4 #(
		.INIT('h135f)
	) name8609 (
		\s1_data_i[28]_pad ,
		\s8_data_i[28]_pad ,
		_w9322_,
		_w9445_,
		_w10510_
	);
	LUT4 #(
		.INIT('h135f)
	) name8610 (
		\s4_data_i[28]_pad ,
		\s9_data_i[28]_pad ,
		_w9433_,
		_w9448_,
		_w10511_
	);
	LUT4 #(
		.INIT('h135f)
	) name8611 (
		\s3_data_i[28]_pad ,
		\s6_data_i[28]_pad ,
		_w9430_,
		_w9439_,
		_w10512_
	);
	LUT4 #(
		.INIT('h135f)
	) name8612 (
		\s10_data_i[28]_pad ,
		\s7_data_i[28]_pad ,
		_w9413_,
		_w9442_,
		_w10513_
	);
	LUT4 #(
		.INIT('h8000)
	) name8613 (
		_w10510_,
		_w10511_,
		_w10512_,
		_w10513_,
		_w10514_
	);
	LUT2 #(
		.INIT('h8)
	) name8614 (
		\s11_data_i[28]_pad ,
		_w9638_,
		_w10515_
	);
	LUT4 #(
		.INIT('h135f)
	) name8615 (
		\s14_data_i[28]_pad ,
		\s2_data_i[28]_pad ,
		_w9422_,
		_w9427_,
		_w10516_
	);
	LUT4 #(
		.INIT('h153f)
	) name8616 (
		\s12_data_i[28]_pad ,
		\s5_data_i[28]_pad ,
		_w9436_,
		_w9635_,
		_w10517_
	);
	LUT4 #(
		.INIT('h135f)
	) name8617 (
		\s0_data_i[28]_pad ,
		\s13_data_i[28]_pad ,
		_w9280_,
		_w9419_,
		_w10518_
	);
	LUT4 #(
		.INIT('h4000)
	) name8618 (
		_w10515_,
		_w10516_,
		_w10517_,
		_w10518_,
		_w10519_
	);
	LUT2 #(
		.INIT('h8)
	) name8619 (
		_w10514_,
		_w10519_,
		_w10520_
	);
	LUT4 #(
		.INIT('h70ff)
	) name8620 (
		_w2046_,
		_w2097_,
		_w10509_,
		_w10520_,
		_w10521_
	);
	LUT2 #(
		.INIT('h8)
	) name8621 (
		\s15_data_i[29]_pad ,
		_w2047_,
		_w10522_
	);
	LUT4 #(
		.INIT('h135f)
	) name8622 (
		\s1_data_i[29]_pad ,
		\s8_data_i[29]_pad ,
		_w9322_,
		_w9445_,
		_w10523_
	);
	LUT4 #(
		.INIT('h135f)
	) name8623 (
		\s4_data_i[29]_pad ,
		\s6_data_i[29]_pad ,
		_w9433_,
		_w9439_,
		_w10524_
	);
	LUT4 #(
		.INIT('h135f)
	) name8624 (
		\s3_data_i[29]_pad ,
		\s9_data_i[29]_pad ,
		_w9430_,
		_w9448_,
		_w10525_
	);
	LUT4 #(
		.INIT('h135f)
	) name8625 (
		\s10_data_i[29]_pad ,
		\s7_data_i[29]_pad ,
		_w9413_,
		_w9442_,
		_w10526_
	);
	LUT4 #(
		.INIT('h8000)
	) name8626 (
		_w10523_,
		_w10524_,
		_w10525_,
		_w10526_,
		_w10527_
	);
	LUT2 #(
		.INIT('h8)
	) name8627 (
		\s11_data_i[29]_pad ,
		_w9638_,
		_w10528_
	);
	LUT4 #(
		.INIT('h135f)
	) name8628 (
		\s14_data_i[29]_pad ,
		\s2_data_i[29]_pad ,
		_w9422_,
		_w9427_,
		_w10529_
	);
	LUT4 #(
		.INIT('h153f)
	) name8629 (
		\s12_data_i[29]_pad ,
		\s5_data_i[29]_pad ,
		_w9436_,
		_w9635_,
		_w10530_
	);
	LUT4 #(
		.INIT('h135f)
	) name8630 (
		\s0_data_i[29]_pad ,
		\s13_data_i[29]_pad ,
		_w9280_,
		_w9419_,
		_w10531_
	);
	LUT4 #(
		.INIT('h4000)
	) name8631 (
		_w10528_,
		_w10529_,
		_w10530_,
		_w10531_,
		_w10532_
	);
	LUT2 #(
		.INIT('h8)
	) name8632 (
		_w10527_,
		_w10532_,
		_w10533_
	);
	LUT4 #(
		.INIT('h70ff)
	) name8633 (
		_w2046_,
		_w2097_,
		_w10522_,
		_w10533_,
		_w10534_
	);
	LUT3 #(
		.INIT('h80)
	) name8634 (
		_w2047_,
		_w2097_,
		_w9993_,
		_w10535_
	);
	LUT2 #(
		.INIT('h8)
	) name8635 (
		\s15_data_i[2]_pad ,
		_w2047_,
		_w10536_
	);
	LUT3 #(
		.INIT('h70)
	) name8636 (
		_w2046_,
		_w2097_,
		_w10536_,
		_w10537_
	);
	LUT4 #(
		.INIT('h153f)
	) name8637 (
		\s12_data_i[2]_pad ,
		\s1_data_i[2]_pad ,
		_w9322_,
		_w9635_,
		_w10538_
	);
	LUT4 #(
		.INIT('h135f)
	) name8638 (
		\s0_data_i[2]_pad ,
		\s10_data_i[2]_pad ,
		_w9280_,
		_w9413_,
		_w10539_
	);
	LUT4 #(
		.INIT('h135f)
	) name8639 (
		\s3_data_i[2]_pad ,
		\s4_data_i[2]_pad ,
		_w9430_,
		_w9433_,
		_w10540_
	);
	LUT4 #(
		.INIT('h135f)
	) name8640 (
		\s6_data_i[2]_pad ,
		\s9_data_i[2]_pad ,
		_w9439_,
		_w9448_,
		_w10541_
	);
	LUT4 #(
		.INIT('h8000)
	) name8641 (
		_w10538_,
		_w10539_,
		_w10540_,
		_w10541_,
		_w10542_
	);
	LUT2 #(
		.INIT('h8)
	) name8642 (
		\s14_data_i[2]_pad ,
		_w9422_,
		_w10543_
	);
	LUT4 #(
		.INIT('h153f)
	) name8643 (
		\s11_data_i[2]_pad ,
		\s7_data_i[2]_pad ,
		_w9442_,
		_w9638_,
		_w10544_
	);
	LUT4 #(
		.INIT('h135f)
	) name8644 (
		\s5_data_i[2]_pad ,
		\s8_data_i[2]_pad ,
		_w9436_,
		_w9445_,
		_w10545_
	);
	LUT4 #(
		.INIT('h135f)
	) name8645 (
		\s13_data_i[2]_pad ,
		\s2_data_i[2]_pad ,
		_w9419_,
		_w9427_,
		_w10546_
	);
	LUT4 #(
		.INIT('h4000)
	) name8646 (
		_w10543_,
		_w10544_,
		_w10545_,
		_w10546_,
		_w10547_
	);
	LUT2 #(
		.INIT('h8)
	) name8647 (
		_w10542_,
		_w10547_,
		_w10548_
	);
	LUT3 #(
		.INIT('hef)
	) name8648 (
		_w10535_,
		_w10537_,
		_w10548_,
		_w10549_
	);
	LUT2 #(
		.INIT('h8)
	) name8649 (
		\s15_data_i[30]_pad ,
		_w2047_,
		_w10550_
	);
	LUT4 #(
		.INIT('h135f)
	) name8650 (
		\s1_data_i[30]_pad ,
		\s8_data_i[30]_pad ,
		_w9322_,
		_w9445_,
		_w10551_
	);
	LUT4 #(
		.INIT('h135f)
	) name8651 (
		\s4_data_i[30]_pad ,
		\s6_data_i[30]_pad ,
		_w9433_,
		_w9439_,
		_w10552_
	);
	LUT4 #(
		.INIT('h135f)
	) name8652 (
		\s3_data_i[30]_pad ,
		\s9_data_i[30]_pad ,
		_w9430_,
		_w9448_,
		_w10553_
	);
	LUT4 #(
		.INIT('h135f)
	) name8653 (
		\s10_data_i[30]_pad ,
		\s7_data_i[30]_pad ,
		_w9413_,
		_w9442_,
		_w10554_
	);
	LUT4 #(
		.INIT('h8000)
	) name8654 (
		_w10551_,
		_w10552_,
		_w10553_,
		_w10554_,
		_w10555_
	);
	LUT2 #(
		.INIT('h8)
	) name8655 (
		\s11_data_i[30]_pad ,
		_w9638_,
		_w10556_
	);
	LUT4 #(
		.INIT('h135f)
	) name8656 (
		\s14_data_i[30]_pad ,
		\s2_data_i[30]_pad ,
		_w9422_,
		_w9427_,
		_w10557_
	);
	LUT4 #(
		.INIT('h153f)
	) name8657 (
		\s12_data_i[30]_pad ,
		\s5_data_i[30]_pad ,
		_w9436_,
		_w9635_,
		_w10558_
	);
	LUT4 #(
		.INIT('h135f)
	) name8658 (
		\s0_data_i[30]_pad ,
		\s13_data_i[30]_pad ,
		_w9280_,
		_w9419_,
		_w10559_
	);
	LUT4 #(
		.INIT('h4000)
	) name8659 (
		_w10556_,
		_w10557_,
		_w10558_,
		_w10559_,
		_w10560_
	);
	LUT2 #(
		.INIT('h8)
	) name8660 (
		_w10555_,
		_w10560_,
		_w10561_
	);
	LUT4 #(
		.INIT('h70ff)
	) name8661 (
		_w2046_,
		_w2097_,
		_w10550_,
		_w10561_,
		_w10562_
	);
	LUT2 #(
		.INIT('h8)
	) name8662 (
		\s15_data_i[31]_pad ,
		_w2047_,
		_w10563_
	);
	LUT4 #(
		.INIT('h135f)
	) name8663 (
		\s1_data_i[31]_pad ,
		\s8_data_i[31]_pad ,
		_w9322_,
		_w9445_,
		_w10564_
	);
	LUT4 #(
		.INIT('h135f)
	) name8664 (
		\s4_data_i[31]_pad ,
		\s6_data_i[31]_pad ,
		_w9433_,
		_w9439_,
		_w10565_
	);
	LUT4 #(
		.INIT('h135f)
	) name8665 (
		\s3_data_i[31]_pad ,
		\s9_data_i[31]_pad ,
		_w9430_,
		_w9448_,
		_w10566_
	);
	LUT4 #(
		.INIT('h135f)
	) name8666 (
		\s10_data_i[31]_pad ,
		\s7_data_i[31]_pad ,
		_w9413_,
		_w9442_,
		_w10567_
	);
	LUT4 #(
		.INIT('h8000)
	) name8667 (
		_w10564_,
		_w10565_,
		_w10566_,
		_w10567_,
		_w10568_
	);
	LUT2 #(
		.INIT('h8)
	) name8668 (
		\s11_data_i[31]_pad ,
		_w9638_,
		_w10569_
	);
	LUT4 #(
		.INIT('h135f)
	) name8669 (
		\s14_data_i[31]_pad ,
		\s2_data_i[31]_pad ,
		_w9422_,
		_w9427_,
		_w10570_
	);
	LUT4 #(
		.INIT('h153f)
	) name8670 (
		\s12_data_i[31]_pad ,
		\s5_data_i[31]_pad ,
		_w9436_,
		_w9635_,
		_w10571_
	);
	LUT4 #(
		.INIT('h135f)
	) name8671 (
		\s0_data_i[31]_pad ,
		\s13_data_i[31]_pad ,
		_w9280_,
		_w9419_,
		_w10572_
	);
	LUT4 #(
		.INIT('h4000)
	) name8672 (
		_w10569_,
		_w10570_,
		_w10571_,
		_w10572_,
		_w10573_
	);
	LUT2 #(
		.INIT('h8)
	) name8673 (
		_w10568_,
		_w10573_,
		_w10574_
	);
	LUT4 #(
		.INIT('h70ff)
	) name8674 (
		_w2046_,
		_w2097_,
		_w10563_,
		_w10574_,
		_w10575_
	);
	LUT3 #(
		.INIT('h80)
	) name8675 (
		_w2047_,
		_w2097_,
		_w10035_,
		_w10576_
	);
	LUT2 #(
		.INIT('h8)
	) name8676 (
		\s15_data_i[3]_pad ,
		_w2047_,
		_w10577_
	);
	LUT3 #(
		.INIT('h70)
	) name8677 (
		_w2046_,
		_w2097_,
		_w10577_,
		_w10578_
	);
	LUT4 #(
		.INIT('h153f)
	) name8678 (
		\s12_data_i[3]_pad ,
		\s1_data_i[3]_pad ,
		_w9322_,
		_w9635_,
		_w10579_
	);
	LUT4 #(
		.INIT('h135f)
	) name8679 (
		\s7_data_i[3]_pad ,
		\s9_data_i[3]_pad ,
		_w9442_,
		_w9448_,
		_w10580_
	);
	LUT4 #(
		.INIT('h135f)
	) name8680 (
		\s3_data_i[3]_pad ,
		\s6_data_i[3]_pad ,
		_w9430_,
		_w9439_,
		_w10581_
	);
	LUT4 #(
		.INIT('h135f)
	) name8681 (
		\s10_data_i[3]_pad ,
		\s13_data_i[3]_pad ,
		_w9413_,
		_w9419_,
		_w10582_
	);
	LUT4 #(
		.INIT('h8000)
	) name8682 (
		_w10579_,
		_w10580_,
		_w10581_,
		_w10582_,
		_w10583_
	);
	LUT2 #(
		.INIT('h8)
	) name8683 (
		\s14_data_i[3]_pad ,
		_w9422_,
		_w10584_
	);
	LUT4 #(
		.INIT('h153f)
	) name8684 (
		\s11_data_i[3]_pad ,
		\s2_data_i[3]_pad ,
		_w9427_,
		_w9638_,
		_w10585_
	);
	LUT4 #(
		.INIT('h135f)
	) name8685 (
		\s5_data_i[3]_pad ,
		\s8_data_i[3]_pad ,
		_w9436_,
		_w9445_,
		_w10586_
	);
	LUT4 #(
		.INIT('h135f)
	) name8686 (
		\s0_data_i[3]_pad ,
		\s4_data_i[3]_pad ,
		_w9280_,
		_w9433_,
		_w10587_
	);
	LUT4 #(
		.INIT('h4000)
	) name8687 (
		_w10584_,
		_w10585_,
		_w10586_,
		_w10587_,
		_w10588_
	);
	LUT2 #(
		.INIT('h8)
	) name8688 (
		_w10583_,
		_w10588_,
		_w10589_
	);
	LUT3 #(
		.INIT('hef)
	) name8689 (
		_w10576_,
		_w10578_,
		_w10589_,
		_w10590_
	);
	LUT3 #(
		.INIT('h80)
	) name8690 (
		_w2047_,
		_w2097_,
		_w10051_,
		_w10591_
	);
	LUT2 #(
		.INIT('h8)
	) name8691 (
		\s15_data_i[4]_pad ,
		_w2047_,
		_w10592_
	);
	LUT3 #(
		.INIT('h70)
	) name8692 (
		_w2046_,
		_w2097_,
		_w10592_,
		_w10593_
	);
	LUT4 #(
		.INIT('h153f)
	) name8693 (
		\s12_data_i[4]_pad ,
		\s1_data_i[4]_pad ,
		_w9322_,
		_w9635_,
		_w10594_
	);
	LUT4 #(
		.INIT('h135f)
	) name8694 (
		\s0_data_i[4]_pad ,
		\s10_data_i[4]_pad ,
		_w9280_,
		_w9413_,
		_w10595_
	);
	LUT4 #(
		.INIT('h135f)
	) name8695 (
		\s3_data_i[4]_pad ,
		\s4_data_i[4]_pad ,
		_w9430_,
		_w9433_,
		_w10596_
	);
	LUT4 #(
		.INIT('h135f)
	) name8696 (
		\s6_data_i[4]_pad ,
		\s9_data_i[4]_pad ,
		_w9439_,
		_w9448_,
		_w10597_
	);
	LUT4 #(
		.INIT('h8000)
	) name8697 (
		_w10594_,
		_w10595_,
		_w10596_,
		_w10597_,
		_w10598_
	);
	LUT2 #(
		.INIT('h8)
	) name8698 (
		\s14_data_i[4]_pad ,
		_w9422_,
		_w10599_
	);
	LUT4 #(
		.INIT('h153f)
	) name8699 (
		\s11_data_i[4]_pad ,
		\s7_data_i[4]_pad ,
		_w9442_,
		_w9638_,
		_w10600_
	);
	LUT4 #(
		.INIT('h135f)
	) name8700 (
		\s5_data_i[4]_pad ,
		\s8_data_i[4]_pad ,
		_w9436_,
		_w9445_,
		_w10601_
	);
	LUT4 #(
		.INIT('h135f)
	) name8701 (
		\s13_data_i[4]_pad ,
		\s2_data_i[4]_pad ,
		_w9419_,
		_w9427_,
		_w10602_
	);
	LUT4 #(
		.INIT('h4000)
	) name8702 (
		_w10599_,
		_w10600_,
		_w10601_,
		_w10602_,
		_w10603_
	);
	LUT2 #(
		.INIT('h8)
	) name8703 (
		_w10598_,
		_w10603_,
		_w10604_
	);
	LUT3 #(
		.INIT('hef)
	) name8704 (
		_w10591_,
		_w10593_,
		_w10604_,
		_w10605_
	);
	LUT3 #(
		.INIT('h80)
	) name8705 (
		_w2047_,
		_w2097_,
		_w10067_,
		_w10606_
	);
	LUT2 #(
		.INIT('h8)
	) name8706 (
		\s15_data_i[5]_pad ,
		_w2047_,
		_w10607_
	);
	LUT3 #(
		.INIT('h70)
	) name8707 (
		_w2046_,
		_w2097_,
		_w10607_,
		_w10608_
	);
	LUT4 #(
		.INIT('h153f)
	) name8708 (
		\s14_data_i[5]_pad ,
		\s1_data_i[5]_pad ,
		_w9322_,
		_w9422_,
		_w10609_
	);
	LUT4 #(
		.INIT('h135f)
	) name8709 (
		\s10_data_i[5]_pad ,
		\s7_data_i[5]_pad ,
		_w9413_,
		_w9442_,
		_w10610_
	);
	LUT4 #(
		.INIT('h135f)
	) name8710 (
		\s2_data_i[5]_pad ,
		\s5_data_i[5]_pad ,
		_w9427_,
		_w9436_,
		_w10611_
	);
	LUT4 #(
		.INIT('h135f)
	) name8711 (
		\s0_data_i[5]_pad ,
		\s6_data_i[5]_pad ,
		_w9280_,
		_w9439_,
		_w10612_
	);
	LUT4 #(
		.INIT('h8000)
	) name8712 (
		_w10609_,
		_w10610_,
		_w10611_,
		_w10612_,
		_w10613_
	);
	LUT2 #(
		.INIT('h8)
	) name8713 (
		\s11_data_i[5]_pad ,
		_w9638_,
		_w10614_
	);
	LUT4 #(
		.INIT('h135f)
	) name8714 (
		\s4_data_i[5]_pad ,
		\s8_data_i[5]_pad ,
		_w9433_,
		_w9445_,
		_w10615_
	);
	LUT4 #(
		.INIT('h153f)
	) name8715 (
		\s12_data_i[5]_pad ,
		\s3_data_i[5]_pad ,
		_w9430_,
		_w9635_,
		_w10616_
	);
	LUT4 #(
		.INIT('h135f)
	) name8716 (
		\s13_data_i[5]_pad ,
		\s9_data_i[5]_pad ,
		_w9419_,
		_w9448_,
		_w10617_
	);
	LUT4 #(
		.INIT('h4000)
	) name8717 (
		_w10614_,
		_w10615_,
		_w10616_,
		_w10617_,
		_w10618_
	);
	LUT2 #(
		.INIT('h8)
	) name8718 (
		_w10613_,
		_w10618_,
		_w10619_
	);
	LUT3 #(
		.INIT('hef)
	) name8719 (
		_w10606_,
		_w10608_,
		_w10619_,
		_w10620_
	);
	LUT3 #(
		.INIT('h80)
	) name8720 (
		_w2047_,
		_w2097_,
		_w10083_,
		_w10621_
	);
	LUT2 #(
		.INIT('h8)
	) name8721 (
		\s15_data_i[6]_pad ,
		_w2047_,
		_w10622_
	);
	LUT3 #(
		.INIT('h70)
	) name8722 (
		_w2046_,
		_w2097_,
		_w10622_,
		_w10623_
	);
	LUT4 #(
		.INIT('h153f)
	) name8723 (
		\s12_data_i[6]_pad ,
		\s1_data_i[6]_pad ,
		_w9322_,
		_w9635_,
		_w10624_
	);
	LUT4 #(
		.INIT('h135f)
	) name8724 (
		\s0_data_i[6]_pad ,
		\s10_data_i[6]_pad ,
		_w9280_,
		_w9413_,
		_w10625_
	);
	LUT4 #(
		.INIT('h135f)
	) name8725 (
		\s3_data_i[6]_pad ,
		\s4_data_i[6]_pad ,
		_w9430_,
		_w9433_,
		_w10626_
	);
	LUT4 #(
		.INIT('h135f)
	) name8726 (
		\s6_data_i[6]_pad ,
		\s9_data_i[6]_pad ,
		_w9439_,
		_w9448_,
		_w10627_
	);
	LUT4 #(
		.INIT('h8000)
	) name8727 (
		_w10624_,
		_w10625_,
		_w10626_,
		_w10627_,
		_w10628_
	);
	LUT2 #(
		.INIT('h8)
	) name8728 (
		\s14_data_i[6]_pad ,
		_w9422_,
		_w10629_
	);
	LUT4 #(
		.INIT('h153f)
	) name8729 (
		\s11_data_i[6]_pad ,
		\s7_data_i[6]_pad ,
		_w9442_,
		_w9638_,
		_w10630_
	);
	LUT4 #(
		.INIT('h135f)
	) name8730 (
		\s5_data_i[6]_pad ,
		\s8_data_i[6]_pad ,
		_w9436_,
		_w9445_,
		_w10631_
	);
	LUT4 #(
		.INIT('h135f)
	) name8731 (
		\s13_data_i[6]_pad ,
		\s2_data_i[6]_pad ,
		_w9419_,
		_w9427_,
		_w10632_
	);
	LUT4 #(
		.INIT('h4000)
	) name8732 (
		_w10629_,
		_w10630_,
		_w10631_,
		_w10632_,
		_w10633_
	);
	LUT2 #(
		.INIT('h8)
	) name8733 (
		_w10628_,
		_w10633_,
		_w10634_
	);
	LUT3 #(
		.INIT('hef)
	) name8734 (
		_w10621_,
		_w10623_,
		_w10634_,
		_w10635_
	);
	LUT3 #(
		.INIT('h80)
	) name8735 (
		_w2047_,
		_w2097_,
		_w10099_,
		_w10636_
	);
	LUT2 #(
		.INIT('h8)
	) name8736 (
		\s15_data_i[7]_pad ,
		_w2047_,
		_w10637_
	);
	LUT3 #(
		.INIT('h70)
	) name8737 (
		_w2046_,
		_w2097_,
		_w10637_,
		_w10638_
	);
	LUT4 #(
		.INIT('h153f)
	) name8738 (
		\s12_data_i[7]_pad ,
		\s1_data_i[7]_pad ,
		_w9322_,
		_w9635_,
		_w10639_
	);
	LUT4 #(
		.INIT('h135f)
	) name8739 (
		\s0_data_i[7]_pad ,
		\s10_data_i[7]_pad ,
		_w9280_,
		_w9413_,
		_w10640_
	);
	LUT4 #(
		.INIT('h135f)
	) name8740 (
		\s3_data_i[7]_pad ,
		\s4_data_i[7]_pad ,
		_w9430_,
		_w9433_,
		_w10641_
	);
	LUT4 #(
		.INIT('h135f)
	) name8741 (
		\s6_data_i[7]_pad ,
		\s9_data_i[7]_pad ,
		_w9439_,
		_w9448_,
		_w10642_
	);
	LUT4 #(
		.INIT('h8000)
	) name8742 (
		_w10639_,
		_w10640_,
		_w10641_,
		_w10642_,
		_w10643_
	);
	LUT2 #(
		.INIT('h8)
	) name8743 (
		\s14_data_i[7]_pad ,
		_w9422_,
		_w10644_
	);
	LUT4 #(
		.INIT('h153f)
	) name8744 (
		\s11_data_i[7]_pad ,
		\s7_data_i[7]_pad ,
		_w9442_,
		_w9638_,
		_w10645_
	);
	LUT4 #(
		.INIT('h135f)
	) name8745 (
		\s5_data_i[7]_pad ,
		\s8_data_i[7]_pad ,
		_w9436_,
		_w9445_,
		_w10646_
	);
	LUT4 #(
		.INIT('h135f)
	) name8746 (
		\s13_data_i[7]_pad ,
		\s2_data_i[7]_pad ,
		_w9419_,
		_w9427_,
		_w10647_
	);
	LUT4 #(
		.INIT('h4000)
	) name8747 (
		_w10644_,
		_w10645_,
		_w10646_,
		_w10647_,
		_w10648_
	);
	LUT2 #(
		.INIT('h8)
	) name8748 (
		_w10643_,
		_w10648_,
		_w10649_
	);
	LUT3 #(
		.INIT('hef)
	) name8749 (
		_w10636_,
		_w10638_,
		_w10649_,
		_w10650_
	);
	LUT3 #(
		.INIT('h80)
	) name8750 (
		_w2047_,
		_w2097_,
		_w10115_,
		_w10651_
	);
	LUT2 #(
		.INIT('h8)
	) name8751 (
		\s15_data_i[8]_pad ,
		_w2047_,
		_w10652_
	);
	LUT3 #(
		.INIT('h70)
	) name8752 (
		_w2046_,
		_w2097_,
		_w10652_,
		_w10653_
	);
	LUT4 #(
		.INIT('h153f)
	) name8753 (
		\s12_data_i[8]_pad ,
		\s1_data_i[8]_pad ,
		_w9322_,
		_w9635_,
		_w10654_
	);
	LUT4 #(
		.INIT('h135f)
	) name8754 (
		\s0_data_i[8]_pad ,
		\s10_data_i[8]_pad ,
		_w9280_,
		_w9413_,
		_w10655_
	);
	LUT4 #(
		.INIT('h135f)
	) name8755 (
		\s3_data_i[8]_pad ,
		\s4_data_i[8]_pad ,
		_w9430_,
		_w9433_,
		_w10656_
	);
	LUT4 #(
		.INIT('h135f)
	) name8756 (
		\s6_data_i[8]_pad ,
		\s9_data_i[8]_pad ,
		_w9439_,
		_w9448_,
		_w10657_
	);
	LUT4 #(
		.INIT('h8000)
	) name8757 (
		_w10654_,
		_w10655_,
		_w10656_,
		_w10657_,
		_w10658_
	);
	LUT2 #(
		.INIT('h8)
	) name8758 (
		\s14_data_i[8]_pad ,
		_w9422_,
		_w10659_
	);
	LUT4 #(
		.INIT('h153f)
	) name8759 (
		\s11_data_i[8]_pad ,
		\s7_data_i[8]_pad ,
		_w9442_,
		_w9638_,
		_w10660_
	);
	LUT4 #(
		.INIT('h135f)
	) name8760 (
		\s5_data_i[8]_pad ,
		\s8_data_i[8]_pad ,
		_w9436_,
		_w9445_,
		_w10661_
	);
	LUT4 #(
		.INIT('h135f)
	) name8761 (
		\s13_data_i[8]_pad ,
		\s2_data_i[8]_pad ,
		_w9419_,
		_w9427_,
		_w10662_
	);
	LUT4 #(
		.INIT('h4000)
	) name8762 (
		_w10659_,
		_w10660_,
		_w10661_,
		_w10662_,
		_w10663_
	);
	LUT2 #(
		.INIT('h8)
	) name8763 (
		_w10658_,
		_w10663_,
		_w10664_
	);
	LUT3 #(
		.INIT('hef)
	) name8764 (
		_w10651_,
		_w10653_,
		_w10664_,
		_w10665_
	);
	LUT3 #(
		.INIT('h80)
	) name8765 (
		_w2047_,
		_w2097_,
		_w10131_,
		_w10666_
	);
	LUT2 #(
		.INIT('h8)
	) name8766 (
		\s15_data_i[9]_pad ,
		_w2047_,
		_w10667_
	);
	LUT3 #(
		.INIT('h70)
	) name8767 (
		_w2046_,
		_w2097_,
		_w10667_,
		_w10668_
	);
	LUT4 #(
		.INIT('h135f)
	) name8768 (
		\s1_data_i[9]_pad ,
		\s8_data_i[9]_pad ,
		_w9322_,
		_w9445_,
		_w10669_
	);
	LUT4 #(
		.INIT('h135f)
	) name8769 (
		\s0_data_i[9]_pad ,
		\s10_data_i[9]_pad ,
		_w9280_,
		_w9413_,
		_w10670_
	);
	LUT4 #(
		.INIT('h135f)
	) name8770 (
		\s3_data_i[9]_pad ,
		\s4_data_i[9]_pad ,
		_w9430_,
		_w9433_,
		_w10671_
	);
	LUT4 #(
		.INIT('h135f)
	) name8771 (
		\s6_data_i[9]_pad ,
		\s9_data_i[9]_pad ,
		_w9439_,
		_w9448_,
		_w10672_
	);
	LUT4 #(
		.INIT('h8000)
	) name8772 (
		_w10669_,
		_w10670_,
		_w10671_,
		_w10672_,
		_w10673_
	);
	LUT2 #(
		.INIT('h8)
	) name8773 (
		\s11_data_i[9]_pad ,
		_w9638_,
		_w10674_
	);
	LUT4 #(
		.INIT('h135f)
	) name8774 (
		\s14_data_i[9]_pad ,
		\s7_data_i[9]_pad ,
		_w9422_,
		_w9442_,
		_w10675_
	);
	LUT4 #(
		.INIT('h153f)
	) name8775 (
		\s12_data_i[9]_pad ,
		\s5_data_i[9]_pad ,
		_w9436_,
		_w9635_,
		_w10676_
	);
	LUT4 #(
		.INIT('h135f)
	) name8776 (
		\s13_data_i[9]_pad ,
		\s2_data_i[9]_pad ,
		_w9419_,
		_w9427_,
		_w10677_
	);
	LUT4 #(
		.INIT('h4000)
	) name8777 (
		_w10674_,
		_w10675_,
		_w10676_,
		_w10677_,
		_w10678_
	);
	LUT2 #(
		.INIT('h8)
	) name8778 (
		_w10673_,
		_w10678_,
		_w10679_
	);
	LUT3 #(
		.INIT('hef)
	) name8779 (
		_w10666_,
		_w10668_,
		_w10679_,
		_w10680_
	);
	LUT3 #(
		.INIT('h80)
	) name8780 (
		\s15_err_i_pad ,
		_w1920_,
		_w10203_,
		_w10681_
	);
	LUT4 #(
		.INIT('h2a00)
	) name8781 (
		\s14_err_i_pad ,
		_w9137_,
		_w9138_,
		_w9422_,
		_w10682_
	);
	LUT4 #(
		.INIT('h2a00)
	) name8782 (
		\s8_err_i_pad ,
		_w8821_,
		_w8822_,
		_w9445_,
		_w10683_
	);
	LUT4 #(
		.INIT('h153f)
	) name8783 (
		_w8820_,
		_w9136_,
		_w10682_,
		_w10683_,
		_w10684_
	);
	LUT4 #(
		.INIT('h2a00)
	) name8784 (
		\s9_err_i_pad ,
		_w8865_,
		_w8866_,
		_w9448_,
		_w10685_
	);
	LUT4 #(
		.INIT('h2a00)
	) name8785 (
		\s0_err_i_pad ,
		_w8989_,
		_w8990_,
		_w9280_,
		_w10686_
	);
	LUT4 #(
		.INIT('h135f)
	) name8786 (
		_w8872_,
		_w9008_,
		_w10685_,
		_w10686_,
		_w10687_
	);
	LUT4 #(
		.INIT('h2a00)
	) name8787 (
		\s6_err_i_pad ,
		_w8743_,
		_w8744_,
		_w9439_,
		_w10688_
	);
	LUT4 #(
		.INIT('h2a00)
	) name8788 (
		\s10_err_i_pad ,
		_w8910_,
		_w8911_,
		_w9413_,
		_w10689_
	);
	LUT4 #(
		.INIT('h135f)
	) name8789 (
		_w8742_,
		_w8923_,
		_w10688_,
		_w10689_,
		_w10690_
	);
	LUT4 #(
		.INIT('h2a00)
	) name8790 (
		\s4_err_i_pad ,
		_w8655_,
		_w8656_,
		_w9433_,
		_w10691_
	);
	LUT4 #(
		.INIT('h2a00)
	) name8791 (
		\s13_err_i_pad ,
		_w9069_,
		_w9070_,
		_w9419_,
		_w10692_
	);
	LUT4 #(
		.INIT('h135f)
	) name8792 (
		_w8662_,
		_w9076_,
		_w10691_,
		_w10692_,
		_w10693_
	);
	LUT4 #(
		.INIT('h8000)
	) name8793 (
		_w10684_,
		_w10687_,
		_w10690_,
		_w10693_,
		_w10694_
	);
	LUT4 #(
		.INIT('h2a00)
	) name8794 (
		\s12_err_i_pad ,
		_w9029_,
		_w9030_,
		_w9635_,
		_w10695_
	);
	LUT2 #(
		.INIT('h8)
	) name8795 (
		_w9048_,
		_w10695_,
		_w10696_
	);
	LUT4 #(
		.INIT('h2a00)
	) name8796 (
		\s5_err_i_pad ,
		_w8699_,
		_w8700_,
		_w9436_,
		_w10697_
	);
	LUT4 #(
		.INIT('h2a00)
	) name8797 (
		\s7_err_i_pad ,
		_w8782_,
		_w8783_,
		_w9442_,
		_w10698_
	);
	LUT4 #(
		.INIT('h135f)
	) name8798 (
		_w8718_,
		_w8789_,
		_w10697_,
		_w10698_,
		_w10699_
	);
	LUT4 #(
		.INIT('h2a00)
	) name8799 (
		\s1_err_i_pad ,
		_w9103_,
		_w9104_,
		_w9322_,
		_w10700_
	);
	LUT4 #(
		.INIT('h2a00)
	) name8800 (
		\s2_err_i_pad ,
		_w9171_,
		_w9172_,
		_w9427_,
		_w10701_
	);
	LUT4 #(
		.INIT('h135f)
	) name8801 (
		_w9122_,
		_w9178_,
		_w10700_,
		_w10701_,
		_w10702_
	);
	LUT4 #(
		.INIT('h2a00)
	) name8802 (
		\s11_err_i_pad ,
		_w8955_,
		_w8956_,
		_w9638_,
		_w10703_
	);
	LUT4 #(
		.INIT('h2a00)
	) name8803 (
		\s3_err_i_pad ,
		_w9205_,
		_w9206_,
		_w9430_,
		_w10704_
	);
	LUT4 #(
		.INIT('h135f)
	) name8804 (
		_w8962_,
		_w9224_,
		_w10703_,
		_w10704_,
		_w10705_
	);
	LUT4 #(
		.INIT('h4000)
	) name8805 (
		_w10696_,
		_w10699_,
		_w10702_,
		_w10705_,
		_w10706_
	);
	LUT2 #(
		.INIT('h8)
	) name8806 (
		_w10694_,
		_w10706_,
		_w10707_
	);
	LUT4 #(
		.INIT('h70ff)
	) name8807 (
		_w2046_,
		_w2097_,
		_w10681_,
		_w10707_,
		_w10708_
	);
	LUT3 #(
		.INIT('h80)
	) name8808 (
		\s15_rty_i_pad ,
		_w1920_,
		_w10203_,
		_w10709_
	);
	LUT4 #(
		.INIT('h2a00)
	) name8809 (
		\s5_rty_i_pad ,
		_w8699_,
		_w8700_,
		_w9436_,
		_w10710_
	);
	LUT4 #(
		.INIT('h2a00)
	) name8810 (
		\s12_rty_i_pad ,
		_w9029_,
		_w9030_,
		_w9635_,
		_w10711_
	);
	LUT4 #(
		.INIT('h135f)
	) name8811 (
		_w8718_,
		_w9048_,
		_w10710_,
		_w10711_,
		_w10712_
	);
	LUT4 #(
		.INIT('h2a00)
	) name8812 (
		\s6_rty_i_pad ,
		_w8743_,
		_w8744_,
		_w9439_,
		_w10713_
	);
	LUT4 #(
		.INIT('h2a00)
	) name8813 (
		\s9_rty_i_pad ,
		_w8865_,
		_w8866_,
		_w9448_,
		_w10714_
	);
	LUT4 #(
		.INIT('h135f)
	) name8814 (
		_w8742_,
		_w8872_,
		_w10713_,
		_w10714_,
		_w10715_
	);
	LUT4 #(
		.INIT('h2a00)
	) name8815 (
		\s0_rty_i_pad ,
		_w8989_,
		_w8990_,
		_w9280_,
		_w10716_
	);
	LUT4 #(
		.INIT('h2a00)
	) name8816 (
		\s7_rty_i_pad ,
		_w8782_,
		_w8783_,
		_w9442_,
		_w10717_
	);
	LUT4 #(
		.INIT('h153f)
	) name8817 (
		_w8789_,
		_w9008_,
		_w10716_,
		_w10717_,
		_w10718_
	);
	LUT4 #(
		.INIT('h2a00)
	) name8818 (
		\s10_rty_i_pad ,
		_w8910_,
		_w8911_,
		_w9413_,
		_w10719_
	);
	LUT4 #(
		.INIT('h2a00)
	) name8819 (
		\s13_rty_i_pad ,
		_w9069_,
		_w9070_,
		_w9419_,
		_w10720_
	);
	LUT4 #(
		.INIT('h135f)
	) name8820 (
		_w8923_,
		_w9076_,
		_w10719_,
		_w10720_,
		_w10721_
	);
	LUT4 #(
		.INIT('h8000)
	) name8821 (
		_w10712_,
		_w10715_,
		_w10718_,
		_w10721_,
		_w10722_
	);
	LUT4 #(
		.INIT('h2a00)
	) name8822 (
		\s3_rty_i_pad ,
		_w9205_,
		_w9206_,
		_w9430_,
		_w10723_
	);
	LUT2 #(
		.INIT('h8)
	) name8823 (
		_w9224_,
		_w10723_,
		_w10724_
	);
	LUT4 #(
		.INIT('h2a00)
	) name8824 (
		\s2_rty_i_pad ,
		_w9171_,
		_w9172_,
		_w9427_,
		_w10725_
	);
	LUT4 #(
		.INIT('h2a00)
	) name8825 (
		\s4_rty_i_pad ,
		_w8655_,
		_w8656_,
		_w9433_,
		_w10726_
	);
	LUT4 #(
		.INIT('h153f)
	) name8826 (
		_w8662_,
		_w9178_,
		_w10725_,
		_w10726_,
		_w10727_
	);
	LUT4 #(
		.INIT('h2a00)
	) name8827 (
		\s8_rty_i_pad ,
		_w8821_,
		_w8822_,
		_w9445_,
		_w10728_
	);
	LUT4 #(
		.INIT('h2a00)
	) name8828 (
		\s11_rty_i_pad ,
		_w8955_,
		_w8956_,
		_w9638_,
		_w10729_
	);
	LUT4 #(
		.INIT('h135f)
	) name8829 (
		_w8820_,
		_w8962_,
		_w10728_,
		_w10729_,
		_w10730_
	);
	LUT4 #(
		.INIT('h2a00)
	) name8830 (
		\s14_rty_i_pad ,
		_w9137_,
		_w9138_,
		_w9422_,
		_w10731_
	);
	LUT4 #(
		.INIT('h2a00)
	) name8831 (
		\s1_rty_i_pad ,
		_w9103_,
		_w9104_,
		_w9322_,
		_w10732_
	);
	LUT4 #(
		.INIT('h153f)
	) name8832 (
		_w9122_,
		_w9136_,
		_w10731_,
		_w10732_,
		_w10733_
	);
	LUT4 #(
		.INIT('h4000)
	) name8833 (
		_w10724_,
		_w10727_,
		_w10730_,
		_w10733_,
		_w10734_
	);
	LUT2 #(
		.INIT('h8)
	) name8834 (
		_w10722_,
		_w10734_,
		_w10735_
	);
	LUT4 #(
		.INIT('h70ff)
	) name8835 (
		_w2046_,
		_w2097_,
		_w10709_,
		_w10735_,
		_w10736_
	);
	LUT3 #(
		.INIT('h70)
	) name8836 (
		_w1908_,
		_w1909_,
		_w2057_,
		_w10737_
	);
	LUT2 #(
		.INIT('h8)
	) name8837 (
		_w1914_,
		_w10737_,
		_w10738_
	);
	LUT3 #(
		.INIT('h70)
	) name8838 (
		_w2097_,
		_w8630_,
		_w10738_,
		_w10739_
	);
	LUT4 #(
		.INIT('h8000)
	) name8839 (
		\s11_ack_i_pad ,
		_w8955_,
		_w8956_,
		_w9454_,
		_w10740_
	);
	LUT4 #(
		.INIT('h8000)
	) name8840 (
		\s3_ack_i_pad ,
		_w9205_,
		_w9206_,
		_w9465_,
		_w10741_
	);
	LUT4 #(
		.INIT('h135f)
	) name8841 (
		_w8974_,
		_w9212_,
		_w10740_,
		_w10741_,
		_w10742_
	);
	LUT4 #(
		.INIT('h8000)
	) name8842 (
		\s1_ack_i_pad ,
		_w9103_,
		_w9104_,
		_w9288_,
		_w10743_
	);
	LUT4 #(
		.INIT('h8000)
	) name8843 (
		\s7_ack_i_pad ,
		_w8782_,
		_w8783_,
		_w9626_,
		_w10744_
	);
	LUT4 #(
		.INIT('h153f)
	) name8844 (
		_w8795_,
		_w9110_,
		_w10743_,
		_w10744_,
		_w10745_
	);
	LUT4 #(
		.INIT('h8000)
	) name8845 (
		\s10_ack_i_pad ,
		_w8910_,
		_w8911_,
		_w9451_,
		_w10746_
	);
	LUT4 #(
		.INIT('h8000)
	) name8846 (
		\s2_ack_i_pad ,
		_w9171_,
		_w9172_,
		_w9462_,
		_w10747_
	);
	LUT4 #(
		.INIT('h135f)
	) name8847 (
		_w8909_,
		_w9190_,
		_w10746_,
		_w10747_,
		_w10748_
	);
	LUT4 #(
		.INIT('h8000)
	) name8848 (
		\s13_ack_i_pad ,
		_w9069_,
		_w9070_,
		_w9629_,
		_w10749_
	);
	LUT4 #(
		.INIT('h8000)
	) name8849 (
		\s6_ack_i_pad ,
		_w8743_,
		_w8744_,
		_w9474_,
		_w10750_
	);
	LUT4 #(
		.INIT('h153f)
	) name8850 (
		_w8750_,
		_w9082_,
		_w10749_,
		_w10750_,
		_w10751_
	);
	LUT4 #(
		.INIT('h8000)
	) name8851 (
		_w10742_,
		_w10745_,
		_w10748_,
		_w10751_,
		_w10752_
	);
	LUT4 #(
		.INIT('h8000)
	) name8852 (
		\s8_ack_i_pad ,
		_w8821_,
		_w8822_,
		_w9620_,
		_w10753_
	);
	LUT2 #(
		.INIT('h8)
	) name8853 (
		_w8828_,
		_w10753_,
		_w10754_
	);
	LUT4 #(
		.INIT('h8000)
	) name8854 (
		\s14_ack_i_pad ,
		_w9137_,
		_w9138_,
		_w9632_,
		_w10755_
	);
	LUT4 #(
		.INIT('h8000)
	) name8855 (
		\s9_ack_i_pad ,
		_w8865_,
		_w8866_,
		_w9477_,
		_w10756_
	);
	LUT4 #(
		.INIT('h153f)
	) name8856 (
		_w8864_,
		_w9144_,
		_w10755_,
		_w10756_,
		_w10757_
	);
	LUT4 #(
		.INIT('h8000)
	) name8857 (
		\s4_ack_i_pad ,
		_w8655_,
		_w8656_,
		_w9468_,
		_w10758_
	);
	LUT4 #(
		.INIT('h8000)
	) name8858 (
		\s0_ack_i_pad ,
		_w8989_,
		_w8990_,
		_w9284_,
		_w10759_
	);
	LUT4 #(
		.INIT('h135f)
	) name8859 (
		_w8668_,
		_w9002_,
		_w10758_,
		_w10759_,
		_w10760_
	);
	LUT4 #(
		.INIT('h8000)
	) name8860 (
		\s5_ack_i_pad ,
		_w8699_,
		_w8700_,
		_w9471_,
		_w10761_
	);
	LUT4 #(
		.INIT('h8000)
	) name8861 (
		\s12_ack_i_pad ,
		_w9029_,
		_w9030_,
		_w9457_,
		_w10762_
	);
	LUT4 #(
		.INIT('h135f)
	) name8862 (
		_w8698_,
		_w9028_,
		_w10761_,
		_w10762_,
		_w10763_
	);
	LUT4 #(
		.INIT('h4000)
	) name8863 (
		_w10754_,
		_w10757_,
		_w10760_,
		_w10763_,
		_w10764_
	);
	LUT2 #(
		.INIT('h8)
	) name8864 (
		_w10752_,
		_w10764_,
		_w10765_
	);
	LUT3 #(
		.INIT('h4f)
	) name8865 (
		_w9652_,
		_w10739_,
		_w10765_,
		_w10766_
	);
	LUT3 #(
		.INIT('h80)
	) name8866 (
		_w2057_,
		_w2097_,
		_w9683_,
		_w10767_
	);
	LUT2 #(
		.INIT('h8)
	) name8867 (
		\s15_data_i[0]_pad ,
		_w2057_,
		_w10768_
	);
	LUT3 #(
		.INIT('h70)
	) name8868 (
		_w2046_,
		_w2097_,
		_w10768_,
		_w10769_
	);
	LUT4 #(
		.INIT('h153f)
	) name8869 (
		\s13_data_i[0]_pad ,
		\s2_data_i[0]_pad ,
		_w9462_,
		_w9629_,
		_w10770_
	);
	LUT4 #(
		.INIT('h135f)
	) name8870 (
		\s3_data_i[0]_pad ,
		\s7_data_i[0]_pad ,
		_w9465_,
		_w9626_,
		_w10771_
	);
	LUT4 #(
		.INIT('h135f)
	) name8871 (
		\s11_data_i[0]_pad ,
		\s5_data_i[0]_pad ,
		_w9454_,
		_w9471_,
		_w10772_
	);
	LUT4 #(
		.INIT('h153f)
	) name8872 (
		\s14_data_i[0]_pad ,
		\s8_data_i[0]_pad ,
		_w9620_,
		_w9632_,
		_w10773_
	);
	LUT4 #(
		.INIT('h8000)
	) name8873 (
		_w10770_,
		_w10771_,
		_w10772_,
		_w10773_,
		_w10774_
	);
	LUT2 #(
		.INIT('h8)
	) name8874 (
		\s1_data_i[0]_pad ,
		_w9288_,
		_w10775_
	);
	LUT4 #(
		.INIT('h135f)
	) name8875 (
		\s12_data_i[0]_pad ,
		\s4_data_i[0]_pad ,
		_w9457_,
		_w9468_,
		_w10776_
	);
	LUT4 #(
		.INIT('h135f)
	) name8876 (
		\s10_data_i[0]_pad ,
		\s9_data_i[0]_pad ,
		_w9451_,
		_w9477_,
		_w10777_
	);
	LUT4 #(
		.INIT('h135f)
	) name8877 (
		\s0_data_i[0]_pad ,
		\s6_data_i[0]_pad ,
		_w9284_,
		_w9474_,
		_w10778_
	);
	LUT4 #(
		.INIT('h4000)
	) name8878 (
		_w10775_,
		_w10776_,
		_w10777_,
		_w10778_,
		_w10779_
	);
	LUT2 #(
		.INIT('h8)
	) name8879 (
		_w10774_,
		_w10779_,
		_w10780_
	);
	LUT3 #(
		.INIT('hef)
	) name8880 (
		_w10767_,
		_w10769_,
		_w10780_,
		_w10781_
	);
	LUT3 #(
		.INIT('h80)
	) name8881 (
		_w2057_,
		_w2097_,
		_w9699_,
		_w10782_
	);
	LUT2 #(
		.INIT('h8)
	) name8882 (
		\s15_data_i[10]_pad ,
		_w2057_,
		_w10783_
	);
	LUT3 #(
		.INIT('h70)
	) name8883 (
		_w2046_,
		_w2097_,
		_w10783_,
		_w10784_
	);
	LUT4 #(
		.INIT('h153f)
	) name8884 (
		\s13_data_i[10]_pad ,
		\s8_data_i[10]_pad ,
		_w9620_,
		_w9629_,
		_w10785_
	);
	LUT4 #(
		.INIT('h153f)
	) name8885 (
		\s10_data_i[10]_pad ,
		\s1_data_i[10]_pad ,
		_w9288_,
		_w9451_,
		_w10786_
	);
	LUT4 #(
		.INIT('h135f)
	) name8886 (
		\s5_data_i[10]_pad ,
		\s6_data_i[10]_pad ,
		_w9471_,
		_w9474_,
		_w10787_
	);
	LUT4 #(
		.INIT('h135f)
	) name8887 (
		\s2_data_i[10]_pad ,
		\s7_data_i[10]_pad ,
		_w9462_,
		_w9626_,
		_w10788_
	);
	LUT4 #(
		.INIT('h8000)
	) name8888 (
		_w10785_,
		_w10786_,
		_w10787_,
		_w10788_,
		_w10789_
	);
	LUT2 #(
		.INIT('h8)
	) name8889 (
		\s11_data_i[10]_pad ,
		_w9454_,
		_w10790_
	);
	LUT4 #(
		.INIT('h135f)
	) name8890 (
		\s3_data_i[10]_pad ,
		\s4_data_i[10]_pad ,
		_w9465_,
		_w9468_,
		_w10791_
	);
	LUT4 #(
		.INIT('h135f)
	) name8891 (
		\s12_data_i[10]_pad ,
		\s14_data_i[10]_pad ,
		_w9457_,
		_w9632_,
		_w10792_
	);
	LUT4 #(
		.INIT('h135f)
	) name8892 (
		\s0_data_i[10]_pad ,
		\s9_data_i[10]_pad ,
		_w9284_,
		_w9477_,
		_w10793_
	);
	LUT4 #(
		.INIT('h4000)
	) name8893 (
		_w10790_,
		_w10791_,
		_w10792_,
		_w10793_,
		_w10794_
	);
	LUT2 #(
		.INIT('h8)
	) name8894 (
		_w10789_,
		_w10794_,
		_w10795_
	);
	LUT3 #(
		.INIT('hef)
	) name8895 (
		_w10782_,
		_w10784_,
		_w10795_,
		_w10796_
	);
	LUT3 #(
		.INIT('h80)
	) name8896 (
		_w2057_,
		_w2097_,
		_w9715_,
		_w10797_
	);
	LUT2 #(
		.INIT('h8)
	) name8897 (
		\s15_data_i[11]_pad ,
		_w2057_,
		_w10798_
	);
	LUT3 #(
		.INIT('h70)
	) name8898 (
		_w2046_,
		_w2097_,
		_w10798_,
		_w10799_
	);
	LUT4 #(
		.INIT('h153f)
	) name8899 (
		\s13_data_i[11]_pad ,
		\s8_data_i[11]_pad ,
		_w9620_,
		_w9629_,
		_w10800_
	);
	LUT4 #(
		.INIT('h153f)
	) name8900 (
		\s10_data_i[11]_pad ,
		\s1_data_i[11]_pad ,
		_w9288_,
		_w9451_,
		_w10801_
	);
	LUT4 #(
		.INIT('h135f)
	) name8901 (
		\s5_data_i[11]_pad ,
		\s6_data_i[11]_pad ,
		_w9471_,
		_w9474_,
		_w10802_
	);
	LUT4 #(
		.INIT('h135f)
	) name8902 (
		\s2_data_i[11]_pad ,
		\s7_data_i[11]_pad ,
		_w9462_,
		_w9626_,
		_w10803_
	);
	LUT4 #(
		.INIT('h8000)
	) name8903 (
		_w10800_,
		_w10801_,
		_w10802_,
		_w10803_,
		_w10804_
	);
	LUT2 #(
		.INIT('h8)
	) name8904 (
		\s11_data_i[11]_pad ,
		_w9454_,
		_w10805_
	);
	LUT4 #(
		.INIT('h135f)
	) name8905 (
		\s3_data_i[11]_pad ,
		\s4_data_i[11]_pad ,
		_w9465_,
		_w9468_,
		_w10806_
	);
	LUT4 #(
		.INIT('h135f)
	) name8906 (
		\s12_data_i[11]_pad ,
		\s14_data_i[11]_pad ,
		_w9457_,
		_w9632_,
		_w10807_
	);
	LUT4 #(
		.INIT('h135f)
	) name8907 (
		\s0_data_i[11]_pad ,
		\s9_data_i[11]_pad ,
		_w9284_,
		_w9477_,
		_w10808_
	);
	LUT4 #(
		.INIT('h4000)
	) name8908 (
		_w10805_,
		_w10806_,
		_w10807_,
		_w10808_,
		_w10809_
	);
	LUT2 #(
		.INIT('h8)
	) name8909 (
		_w10804_,
		_w10809_,
		_w10810_
	);
	LUT3 #(
		.INIT('hef)
	) name8910 (
		_w10797_,
		_w10799_,
		_w10810_,
		_w10811_
	);
	LUT3 #(
		.INIT('h80)
	) name8911 (
		_w2057_,
		_w2097_,
		_w9731_,
		_w10812_
	);
	LUT2 #(
		.INIT('h8)
	) name8912 (
		\s15_data_i[12]_pad ,
		_w2057_,
		_w10813_
	);
	LUT3 #(
		.INIT('h70)
	) name8913 (
		_w2046_,
		_w2097_,
		_w10813_,
		_w10814_
	);
	LUT4 #(
		.INIT('h153f)
	) name8914 (
		\s13_data_i[12]_pad ,
		\s8_data_i[12]_pad ,
		_w9620_,
		_w9629_,
		_w10815_
	);
	LUT4 #(
		.INIT('h153f)
	) name8915 (
		\s10_data_i[12]_pad ,
		\s1_data_i[12]_pad ,
		_w9288_,
		_w9451_,
		_w10816_
	);
	LUT4 #(
		.INIT('h135f)
	) name8916 (
		\s5_data_i[12]_pad ,
		\s6_data_i[12]_pad ,
		_w9471_,
		_w9474_,
		_w10817_
	);
	LUT4 #(
		.INIT('h135f)
	) name8917 (
		\s2_data_i[12]_pad ,
		\s7_data_i[12]_pad ,
		_w9462_,
		_w9626_,
		_w10818_
	);
	LUT4 #(
		.INIT('h8000)
	) name8918 (
		_w10815_,
		_w10816_,
		_w10817_,
		_w10818_,
		_w10819_
	);
	LUT2 #(
		.INIT('h8)
	) name8919 (
		\s11_data_i[12]_pad ,
		_w9454_,
		_w10820_
	);
	LUT4 #(
		.INIT('h135f)
	) name8920 (
		\s3_data_i[12]_pad ,
		\s4_data_i[12]_pad ,
		_w9465_,
		_w9468_,
		_w10821_
	);
	LUT4 #(
		.INIT('h135f)
	) name8921 (
		\s12_data_i[12]_pad ,
		\s14_data_i[12]_pad ,
		_w9457_,
		_w9632_,
		_w10822_
	);
	LUT4 #(
		.INIT('h135f)
	) name8922 (
		\s0_data_i[12]_pad ,
		\s9_data_i[12]_pad ,
		_w9284_,
		_w9477_,
		_w10823_
	);
	LUT4 #(
		.INIT('h4000)
	) name8923 (
		_w10820_,
		_w10821_,
		_w10822_,
		_w10823_,
		_w10824_
	);
	LUT2 #(
		.INIT('h8)
	) name8924 (
		_w10819_,
		_w10824_,
		_w10825_
	);
	LUT3 #(
		.INIT('hef)
	) name8925 (
		_w10812_,
		_w10814_,
		_w10825_,
		_w10826_
	);
	LUT3 #(
		.INIT('h80)
	) name8926 (
		_w2057_,
		_w2097_,
		_w9747_,
		_w10827_
	);
	LUT2 #(
		.INIT('h8)
	) name8927 (
		\s15_data_i[13]_pad ,
		_w2057_,
		_w10828_
	);
	LUT3 #(
		.INIT('h70)
	) name8928 (
		_w2046_,
		_w2097_,
		_w10828_,
		_w10829_
	);
	LUT4 #(
		.INIT('h135f)
	) name8929 (
		\s1_data_i[13]_pad ,
		\s8_data_i[13]_pad ,
		_w9288_,
		_w9620_,
		_w10830_
	);
	LUT4 #(
		.INIT('h135f)
	) name8930 (
		\s4_data_i[13]_pad ,
		\s6_data_i[13]_pad ,
		_w9468_,
		_w9474_,
		_w10831_
	);
	LUT4 #(
		.INIT('h135f)
	) name8931 (
		\s5_data_i[13]_pad ,
		\s9_data_i[13]_pad ,
		_w9471_,
		_w9477_,
		_w10832_
	);
	LUT4 #(
		.INIT('h135f)
	) name8932 (
		\s10_data_i[13]_pad ,
		\s7_data_i[13]_pad ,
		_w9451_,
		_w9626_,
		_w10833_
	);
	LUT4 #(
		.INIT('h8000)
	) name8933 (
		_w10830_,
		_w10831_,
		_w10832_,
		_w10833_,
		_w10834_
	);
	LUT2 #(
		.INIT('h8)
	) name8934 (
		\s11_data_i[13]_pad ,
		_w9454_,
		_w10835_
	);
	LUT4 #(
		.INIT('h153f)
	) name8935 (
		\s13_data_i[13]_pad ,
		\s3_data_i[13]_pad ,
		_w9465_,
		_w9629_,
		_w10836_
	);
	LUT4 #(
		.INIT('h135f)
	) name8936 (
		\s12_data_i[13]_pad ,
		\s14_data_i[13]_pad ,
		_w9457_,
		_w9632_,
		_w10837_
	);
	LUT4 #(
		.INIT('h135f)
	) name8937 (
		\s0_data_i[13]_pad ,
		\s2_data_i[13]_pad ,
		_w9284_,
		_w9462_,
		_w10838_
	);
	LUT4 #(
		.INIT('h4000)
	) name8938 (
		_w10835_,
		_w10836_,
		_w10837_,
		_w10838_,
		_w10839_
	);
	LUT2 #(
		.INIT('h8)
	) name8939 (
		_w10834_,
		_w10839_,
		_w10840_
	);
	LUT3 #(
		.INIT('hef)
	) name8940 (
		_w10827_,
		_w10829_,
		_w10840_,
		_w10841_
	);
	LUT3 #(
		.INIT('h80)
	) name8941 (
		_w2057_,
		_w2097_,
		_w9763_,
		_w10842_
	);
	LUT2 #(
		.INIT('h8)
	) name8942 (
		\s15_data_i[14]_pad ,
		_w2057_,
		_w10843_
	);
	LUT3 #(
		.INIT('h70)
	) name8943 (
		_w2046_,
		_w2097_,
		_w10843_,
		_w10844_
	);
	LUT4 #(
		.INIT('h135f)
	) name8944 (
		\s12_data_i[14]_pad ,
		\s13_data_i[14]_pad ,
		_w9457_,
		_w9629_,
		_w10845_
	);
	LUT4 #(
		.INIT('h153f)
	) name8945 (
		\s10_data_i[14]_pad ,
		\s1_data_i[14]_pad ,
		_w9288_,
		_w9451_,
		_w10846_
	);
	LUT4 #(
		.INIT('h135f)
	) name8946 (
		\s0_data_i[14]_pad ,
		\s5_data_i[14]_pad ,
		_w9284_,
		_w9471_,
		_w10847_
	);
	LUT4 #(
		.INIT('h135f)
	) name8947 (
		\s2_data_i[14]_pad ,
		\s4_data_i[14]_pad ,
		_w9462_,
		_w9468_,
		_w10848_
	);
	LUT4 #(
		.INIT('h8000)
	) name8948 (
		_w10845_,
		_w10846_,
		_w10847_,
		_w10848_,
		_w10849_
	);
	LUT2 #(
		.INIT('h8)
	) name8949 (
		\s14_data_i[14]_pad ,
		_w9632_,
		_w10850_
	);
	LUT4 #(
		.INIT('h135f)
	) name8950 (
		\s3_data_i[14]_pad ,
		\s7_data_i[14]_pad ,
		_w9465_,
		_w9626_,
		_w10851_
	);
	LUT4 #(
		.INIT('h135f)
	) name8951 (
		\s11_data_i[14]_pad ,
		\s8_data_i[14]_pad ,
		_w9454_,
		_w9620_,
		_w10852_
	);
	LUT4 #(
		.INIT('h135f)
	) name8952 (
		\s6_data_i[14]_pad ,
		\s9_data_i[14]_pad ,
		_w9474_,
		_w9477_,
		_w10853_
	);
	LUT4 #(
		.INIT('h4000)
	) name8953 (
		_w10850_,
		_w10851_,
		_w10852_,
		_w10853_,
		_w10854_
	);
	LUT2 #(
		.INIT('h8)
	) name8954 (
		_w10849_,
		_w10854_,
		_w10855_
	);
	LUT3 #(
		.INIT('hef)
	) name8955 (
		_w10842_,
		_w10844_,
		_w10855_,
		_w10856_
	);
	LUT3 #(
		.INIT('h80)
	) name8956 (
		_w2057_,
		_w2097_,
		_w9779_,
		_w10857_
	);
	LUT2 #(
		.INIT('h8)
	) name8957 (
		\s15_data_i[15]_pad ,
		_w2057_,
		_w10858_
	);
	LUT3 #(
		.INIT('h70)
	) name8958 (
		_w2046_,
		_w2097_,
		_w10858_,
		_w10859_
	);
	LUT4 #(
		.INIT('h135f)
	) name8959 (
		\s12_data_i[15]_pad ,
		\s13_data_i[15]_pad ,
		_w9457_,
		_w9629_,
		_w10860_
	);
	LUT4 #(
		.INIT('h135f)
	) name8960 (
		\s10_data_i[15]_pad ,
		\s3_data_i[15]_pad ,
		_w9451_,
		_w9465_,
		_w10861_
	);
	LUT4 #(
		.INIT('h135f)
	) name8961 (
		\s0_data_i[15]_pad ,
		\s2_data_i[15]_pad ,
		_w9284_,
		_w9462_,
		_w10862_
	);
	LUT4 #(
		.INIT('h135f)
	) name8962 (
		\s4_data_i[15]_pad ,
		\s5_data_i[15]_pad ,
		_w9468_,
		_w9471_,
		_w10863_
	);
	LUT4 #(
		.INIT('h8000)
	) name8963 (
		_w10860_,
		_w10861_,
		_w10862_,
		_w10863_,
		_w10864_
	);
	LUT2 #(
		.INIT('h8)
	) name8964 (
		\s14_data_i[15]_pad ,
		_w9632_,
		_w10865_
	);
	LUT4 #(
		.INIT('h135f)
	) name8965 (
		\s1_data_i[15]_pad ,
		\s7_data_i[15]_pad ,
		_w9288_,
		_w9626_,
		_w10866_
	);
	LUT4 #(
		.INIT('h135f)
	) name8966 (
		\s11_data_i[15]_pad ,
		\s8_data_i[15]_pad ,
		_w9454_,
		_w9620_,
		_w10867_
	);
	LUT4 #(
		.INIT('h135f)
	) name8967 (
		\s6_data_i[15]_pad ,
		\s9_data_i[15]_pad ,
		_w9474_,
		_w9477_,
		_w10868_
	);
	LUT4 #(
		.INIT('h4000)
	) name8968 (
		_w10865_,
		_w10866_,
		_w10867_,
		_w10868_,
		_w10869_
	);
	LUT2 #(
		.INIT('h8)
	) name8969 (
		_w10864_,
		_w10869_,
		_w10870_
	);
	LUT3 #(
		.INIT('hef)
	) name8970 (
		_w10857_,
		_w10859_,
		_w10870_,
		_w10871_
	);
	LUT2 #(
		.INIT('h8)
	) name8971 (
		\s15_data_i[16]_pad ,
		_w2057_,
		_w10872_
	);
	LUT4 #(
		.INIT('h135f)
	) name8972 (
		\s12_data_i[16]_pad ,
		\s13_data_i[16]_pad ,
		_w9457_,
		_w9629_,
		_w10873_
	);
	LUT4 #(
		.INIT('h135f)
	) name8973 (
		\s10_data_i[16]_pad ,
		\s3_data_i[16]_pad ,
		_w9451_,
		_w9465_,
		_w10874_
	);
	LUT4 #(
		.INIT('h135f)
	) name8974 (
		\s2_data_i[16]_pad ,
		\s6_data_i[16]_pad ,
		_w9462_,
		_w9474_,
		_w10875_
	);
	LUT4 #(
		.INIT('h135f)
	) name8975 (
		\s5_data_i[16]_pad ,
		\s7_data_i[16]_pad ,
		_w9471_,
		_w9626_,
		_w10876_
	);
	LUT4 #(
		.INIT('h8000)
	) name8976 (
		_w10873_,
		_w10874_,
		_w10875_,
		_w10876_,
		_w10877_
	);
	LUT2 #(
		.INIT('h8)
	) name8977 (
		\s14_data_i[16]_pad ,
		_w9632_,
		_w10878_
	);
	LUT4 #(
		.INIT('h135f)
	) name8978 (
		\s1_data_i[16]_pad ,
		\s4_data_i[16]_pad ,
		_w9288_,
		_w9468_,
		_w10879_
	);
	LUT4 #(
		.INIT('h135f)
	) name8979 (
		\s11_data_i[16]_pad ,
		\s8_data_i[16]_pad ,
		_w9454_,
		_w9620_,
		_w10880_
	);
	LUT4 #(
		.INIT('h135f)
	) name8980 (
		\s0_data_i[16]_pad ,
		\s9_data_i[16]_pad ,
		_w9284_,
		_w9477_,
		_w10881_
	);
	LUT4 #(
		.INIT('h4000)
	) name8981 (
		_w10878_,
		_w10879_,
		_w10880_,
		_w10881_,
		_w10882_
	);
	LUT2 #(
		.INIT('h8)
	) name8982 (
		_w10877_,
		_w10882_,
		_w10883_
	);
	LUT4 #(
		.INIT('h70ff)
	) name8983 (
		_w2046_,
		_w2097_,
		_w10872_,
		_w10883_,
		_w10884_
	);
	LUT2 #(
		.INIT('h8)
	) name8984 (
		\s15_data_i[17]_pad ,
		_w2057_,
		_w10885_
	);
	LUT4 #(
		.INIT('h135f)
	) name8985 (
		\s12_data_i[17]_pad ,
		\s13_data_i[17]_pad ,
		_w9457_,
		_w9629_,
		_w10886_
	);
	LUT4 #(
		.INIT('h153f)
	) name8986 (
		\s10_data_i[17]_pad ,
		\s1_data_i[17]_pad ,
		_w9288_,
		_w9451_,
		_w10887_
	);
	LUT4 #(
		.INIT('h135f)
	) name8987 (
		\s5_data_i[17]_pad ,
		\s6_data_i[17]_pad ,
		_w9471_,
		_w9474_,
		_w10888_
	);
	LUT4 #(
		.INIT('h135f)
	) name8988 (
		\s2_data_i[17]_pad ,
		\s7_data_i[17]_pad ,
		_w9462_,
		_w9626_,
		_w10889_
	);
	LUT4 #(
		.INIT('h8000)
	) name8989 (
		_w10886_,
		_w10887_,
		_w10888_,
		_w10889_,
		_w10890_
	);
	LUT2 #(
		.INIT('h8)
	) name8990 (
		\s14_data_i[17]_pad ,
		_w9632_,
		_w10891_
	);
	LUT4 #(
		.INIT('h135f)
	) name8991 (
		\s3_data_i[17]_pad ,
		\s4_data_i[17]_pad ,
		_w9465_,
		_w9468_,
		_w10892_
	);
	LUT4 #(
		.INIT('h135f)
	) name8992 (
		\s11_data_i[17]_pad ,
		\s8_data_i[17]_pad ,
		_w9454_,
		_w9620_,
		_w10893_
	);
	LUT4 #(
		.INIT('h135f)
	) name8993 (
		\s0_data_i[17]_pad ,
		\s9_data_i[17]_pad ,
		_w9284_,
		_w9477_,
		_w10894_
	);
	LUT4 #(
		.INIT('h4000)
	) name8994 (
		_w10891_,
		_w10892_,
		_w10893_,
		_w10894_,
		_w10895_
	);
	LUT2 #(
		.INIT('h8)
	) name8995 (
		_w10890_,
		_w10895_,
		_w10896_
	);
	LUT4 #(
		.INIT('h70ff)
	) name8996 (
		_w2046_,
		_w2097_,
		_w10885_,
		_w10896_,
		_w10897_
	);
	LUT2 #(
		.INIT('h8)
	) name8997 (
		\s15_data_i[18]_pad ,
		_w2057_,
		_w10898_
	);
	LUT4 #(
		.INIT('h135f)
	) name8998 (
		\s12_data_i[18]_pad ,
		\s13_data_i[18]_pad ,
		_w9457_,
		_w9629_,
		_w10899_
	);
	LUT4 #(
		.INIT('h153f)
	) name8999 (
		\s10_data_i[18]_pad ,
		\s1_data_i[18]_pad ,
		_w9288_,
		_w9451_,
		_w10900_
	);
	LUT4 #(
		.INIT('h135f)
	) name9000 (
		\s5_data_i[18]_pad ,
		\s6_data_i[18]_pad ,
		_w9471_,
		_w9474_,
		_w10901_
	);
	LUT4 #(
		.INIT('h135f)
	) name9001 (
		\s2_data_i[18]_pad ,
		\s7_data_i[18]_pad ,
		_w9462_,
		_w9626_,
		_w10902_
	);
	LUT4 #(
		.INIT('h8000)
	) name9002 (
		_w10899_,
		_w10900_,
		_w10901_,
		_w10902_,
		_w10903_
	);
	LUT2 #(
		.INIT('h8)
	) name9003 (
		\s14_data_i[18]_pad ,
		_w9632_,
		_w10904_
	);
	LUT4 #(
		.INIT('h135f)
	) name9004 (
		\s3_data_i[18]_pad ,
		\s4_data_i[18]_pad ,
		_w9465_,
		_w9468_,
		_w10905_
	);
	LUT4 #(
		.INIT('h135f)
	) name9005 (
		\s11_data_i[18]_pad ,
		\s8_data_i[18]_pad ,
		_w9454_,
		_w9620_,
		_w10906_
	);
	LUT4 #(
		.INIT('h135f)
	) name9006 (
		\s0_data_i[18]_pad ,
		\s9_data_i[18]_pad ,
		_w9284_,
		_w9477_,
		_w10907_
	);
	LUT4 #(
		.INIT('h4000)
	) name9007 (
		_w10904_,
		_w10905_,
		_w10906_,
		_w10907_,
		_w10908_
	);
	LUT2 #(
		.INIT('h8)
	) name9008 (
		_w10903_,
		_w10908_,
		_w10909_
	);
	LUT4 #(
		.INIT('h70ff)
	) name9009 (
		_w2046_,
		_w2097_,
		_w10898_,
		_w10909_,
		_w10910_
	);
	LUT2 #(
		.INIT('h8)
	) name9010 (
		\s15_data_i[19]_pad ,
		_w2057_,
		_w10911_
	);
	LUT4 #(
		.INIT('h135f)
	) name9011 (
		\s12_data_i[19]_pad ,
		\s13_data_i[19]_pad ,
		_w9457_,
		_w9629_,
		_w10912_
	);
	LUT4 #(
		.INIT('h153f)
	) name9012 (
		\s10_data_i[19]_pad ,
		\s1_data_i[19]_pad ,
		_w9288_,
		_w9451_,
		_w10913_
	);
	LUT4 #(
		.INIT('h135f)
	) name9013 (
		\s5_data_i[19]_pad ,
		\s6_data_i[19]_pad ,
		_w9471_,
		_w9474_,
		_w10914_
	);
	LUT4 #(
		.INIT('h135f)
	) name9014 (
		\s2_data_i[19]_pad ,
		\s7_data_i[19]_pad ,
		_w9462_,
		_w9626_,
		_w10915_
	);
	LUT4 #(
		.INIT('h8000)
	) name9015 (
		_w10912_,
		_w10913_,
		_w10914_,
		_w10915_,
		_w10916_
	);
	LUT2 #(
		.INIT('h8)
	) name9016 (
		\s14_data_i[19]_pad ,
		_w9632_,
		_w10917_
	);
	LUT4 #(
		.INIT('h135f)
	) name9017 (
		\s3_data_i[19]_pad ,
		\s4_data_i[19]_pad ,
		_w9465_,
		_w9468_,
		_w10918_
	);
	LUT4 #(
		.INIT('h135f)
	) name9018 (
		\s11_data_i[19]_pad ,
		\s8_data_i[19]_pad ,
		_w9454_,
		_w9620_,
		_w10919_
	);
	LUT4 #(
		.INIT('h135f)
	) name9019 (
		\s0_data_i[19]_pad ,
		\s9_data_i[19]_pad ,
		_w9284_,
		_w9477_,
		_w10920_
	);
	LUT4 #(
		.INIT('h4000)
	) name9020 (
		_w10917_,
		_w10918_,
		_w10919_,
		_w10920_,
		_w10921_
	);
	LUT2 #(
		.INIT('h8)
	) name9021 (
		_w10916_,
		_w10921_,
		_w10922_
	);
	LUT4 #(
		.INIT('h70ff)
	) name9022 (
		_w2046_,
		_w2097_,
		_w10911_,
		_w10922_,
		_w10923_
	);
	LUT3 #(
		.INIT('h80)
	) name9023 (
		_w2057_,
		_w2097_,
		_w9847_,
		_w10924_
	);
	LUT2 #(
		.INIT('h8)
	) name9024 (
		\s15_data_i[1]_pad ,
		_w2057_,
		_w10925_
	);
	LUT3 #(
		.INIT('h70)
	) name9025 (
		_w2046_,
		_w2097_,
		_w10925_,
		_w10926_
	);
	LUT4 #(
		.INIT('h135f)
	) name9026 (
		\s10_data_i[1]_pad ,
		\s8_data_i[1]_pad ,
		_w9451_,
		_w9620_,
		_w10927_
	);
	LUT4 #(
		.INIT('h135f)
	) name9027 (
		\s1_data_i[1]_pad ,
		\s4_data_i[1]_pad ,
		_w9288_,
		_w9468_,
		_w10928_
	);
	LUT4 #(
		.INIT('h135f)
	) name9028 (
		\s0_data_i[1]_pad ,
		\s5_data_i[1]_pad ,
		_w9284_,
		_w9471_,
		_w10929_
	);
	LUT4 #(
		.INIT('h153f)
	) name9029 (
		\s13_data_i[1]_pad ,
		\s2_data_i[1]_pad ,
		_w9462_,
		_w9629_,
		_w10930_
	);
	LUT4 #(
		.INIT('h8000)
	) name9030 (
		_w10927_,
		_w10928_,
		_w10929_,
		_w10930_,
		_w10931_
	);
	LUT2 #(
		.INIT('h8)
	) name9031 (
		\s11_data_i[1]_pad ,
		_w9454_,
		_w10932_
	);
	LUT4 #(
		.INIT('h135f)
	) name9032 (
		\s3_data_i[1]_pad ,
		\s7_data_i[1]_pad ,
		_w9465_,
		_w9626_,
		_w10933_
	);
	LUT4 #(
		.INIT('h135f)
	) name9033 (
		\s12_data_i[1]_pad ,
		\s14_data_i[1]_pad ,
		_w9457_,
		_w9632_,
		_w10934_
	);
	LUT4 #(
		.INIT('h135f)
	) name9034 (
		\s6_data_i[1]_pad ,
		\s9_data_i[1]_pad ,
		_w9474_,
		_w9477_,
		_w10935_
	);
	LUT4 #(
		.INIT('h4000)
	) name9035 (
		_w10932_,
		_w10933_,
		_w10934_,
		_w10935_,
		_w10936_
	);
	LUT2 #(
		.INIT('h8)
	) name9036 (
		_w10931_,
		_w10936_,
		_w10937_
	);
	LUT3 #(
		.INIT('hef)
	) name9037 (
		_w10924_,
		_w10926_,
		_w10937_,
		_w10938_
	);
	LUT2 #(
		.INIT('h8)
	) name9038 (
		\s15_data_i[20]_pad ,
		_w2057_,
		_w10939_
	);
	LUT4 #(
		.INIT('h135f)
	) name9039 (
		\s12_data_i[20]_pad ,
		\s13_data_i[20]_pad ,
		_w9457_,
		_w9629_,
		_w10940_
	);
	LUT4 #(
		.INIT('h153f)
	) name9040 (
		\s10_data_i[20]_pad ,
		\s1_data_i[20]_pad ,
		_w9288_,
		_w9451_,
		_w10941_
	);
	LUT4 #(
		.INIT('h135f)
	) name9041 (
		\s5_data_i[20]_pad ,
		\s6_data_i[20]_pad ,
		_w9471_,
		_w9474_,
		_w10942_
	);
	LUT4 #(
		.INIT('h135f)
	) name9042 (
		\s2_data_i[20]_pad ,
		\s7_data_i[20]_pad ,
		_w9462_,
		_w9626_,
		_w10943_
	);
	LUT4 #(
		.INIT('h8000)
	) name9043 (
		_w10940_,
		_w10941_,
		_w10942_,
		_w10943_,
		_w10944_
	);
	LUT2 #(
		.INIT('h8)
	) name9044 (
		\s14_data_i[20]_pad ,
		_w9632_,
		_w10945_
	);
	LUT4 #(
		.INIT('h135f)
	) name9045 (
		\s3_data_i[20]_pad ,
		\s4_data_i[20]_pad ,
		_w9465_,
		_w9468_,
		_w10946_
	);
	LUT4 #(
		.INIT('h135f)
	) name9046 (
		\s11_data_i[20]_pad ,
		\s8_data_i[20]_pad ,
		_w9454_,
		_w9620_,
		_w10947_
	);
	LUT4 #(
		.INIT('h135f)
	) name9047 (
		\s0_data_i[20]_pad ,
		\s9_data_i[20]_pad ,
		_w9284_,
		_w9477_,
		_w10948_
	);
	LUT4 #(
		.INIT('h4000)
	) name9048 (
		_w10945_,
		_w10946_,
		_w10947_,
		_w10948_,
		_w10949_
	);
	LUT2 #(
		.INIT('h8)
	) name9049 (
		_w10944_,
		_w10949_,
		_w10950_
	);
	LUT4 #(
		.INIT('h70ff)
	) name9050 (
		_w2046_,
		_w2097_,
		_w10939_,
		_w10950_,
		_w10951_
	);
	LUT2 #(
		.INIT('h8)
	) name9051 (
		\s15_data_i[21]_pad ,
		_w2057_,
		_w10952_
	);
	LUT4 #(
		.INIT('h135f)
	) name9052 (
		\s12_data_i[21]_pad ,
		\s13_data_i[21]_pad ,
		_w9457_,
		_w9629_,
		_w10953_
	);
	LUT4 #(
		.INIT('h153f)
	) name9053 (
		\s10_data_i[21]_pad ,
		\s1_data_i[21]_pad ,
		_w9288_,
		_w9451_,
		_w10954_
	);
	LUT4 #(
		.INIT('h135f)
	) name9054 (
		\s5_data_i[21]_pad ,
		\s6_data_i[21]_pad ,
		_w9471_,
		_w9474_,
		_w10955_
	);
	LUT4 #(
		.INIT('h135f)
	) name9055 (
		\s2_data_i[21]_pad ,
		\s7_data_i[21]_pad ,
		_w9462_,
		_w9626_,
		_w10956_
	);
	LUT4 #(
		.INIT('h8000)
	) name9056 (
		_w10953_,
		_w10954_,
		_w10955_,
		_w10956_,
		_w10957_
	);
	LUT2 #(
		.INIT('h8)
	) name9057 (
		\s14_data_i[21]_pad ,
		_w9632_,
		_w10958_
	);
	LUT4 #(
		.INIT('h135f)
	) name9058 (
		\s3_data_i[21]_pad ,
		\s4_data_i[21]_pad ,
		_w9465_,
		_w9468_,
		_w10959_
	);
	LUT4 #(
		.INIT('h135f)
	) name9059 (
		\s11_data_i[21]_pad ,
		\s8_data_i[21]_pad ,
		_w9454_,
		_w9620_,
		_w10960_
	);
	LUT4 #(
		.INIT('h135f)
	) name9060 (
		\s0_data_i[21]_pad ,
		\s9_data_i[21]_pad ,
		_w9284_,
		_w9477_,
		_w10961_
	);
	LUT4 #(
		.INIT('h4000)
	) name9061 (
		_w10958_,
		_w10959_,
		_w10960_,
		_w10961_,
		_w10962_
	);
	LUT2 #(
		.INIT('h8)
	) name9062 (
		_w10957_,
		_w10962_,
		_w10963_
	);
	LUT4 #(
		.INIT('h70ff)
	) name9063 (
		_w2046_,
		_w2097_,
		_w10952_,
		_w10963_,
		_w10964_
	);
	LUT2 #(
		.INIT('h8)
	) name9064 (
		\s15_data_i[22]_pad ,
		_w2057_,
		_w10965_
	);
	LUT4 #(
		.INIT('h135f)
	) name9065 (
		\s12_data_i[22]_pad ,
		\s13_data_i[22]_pad ,
		_w9457_,
		_w9629_,
		_w10966_
	);
	LUT4 #(
		.INIT('h153f)
	) name9066 (
		\s10_data_i[22]_pad ,
		\s1_data_i[22]_pad ,
		_w9288_,
		_w9451_,
		_w10967_
	);
	LUT4 #(
		.INIT('h135f)
	) name9067 (
		\s5_data_i[22]_pad ,
		\s6_data_i[22]_pad ,
		_w9471_,
		_w9474_,
		_w10968_
	);
	LUT4 #(
		.INIT('h135f)
	) name9068 (
		\s2_data_i[22]_pad ,
		\s7_data_i[22]_pad ,
		_w9462_,
		_w9626_,
		_w10969_
	);
	LUT4 #(
		.INIT('h8000)
	) name9069 (
		_w10966_,
		_w10967_,
		_w10968_,
		_w10969_,
		_w10970_
	);
	LUT2 #(
		.INIT('h8)
	) name9070 (
		\s14_data_i[22]_pad ,
		_w9632_,
		_w10971_
	);
	LUT4 #(
		.INIT('h135f)
	) name9071 (
		\s3_data_i[22]_pad ,
		\s4_data_i[22]_pad ,
		_w9465_,
		_w9468_,
		_w10972_
	);
	LUT4 #(
		.INIT('h135f)
	) name9072 (
		\s11_data_i[22]_pad ,
		\s8_data_i[22]_pad ,
		_w9454_,
		_w9620_,
		_w10973_
	);
	LUT4 #(
		.INIT('h135f)
	) name9073 (
		\s0_data_i[22]_pad ,
		\s9_data_i[22]_pad ,
		_w9284_,
		_w9477_,
		_w10974_
	);
	LUT4 #(
		.INIT('h4000)
	) name9074 (
		_w10971_,
		_w10972_,
		_w10973_,
		_w10974_,
		_w10975_
	);
	LUT2 #(
		.INIT('h8)
	) name9075 (
		_w10970_,
		_w10975_,
		_w10976_
	);
	LUT4 #(
		.INIT('h70ff)
	) name9076 (
		_w2046_,
		_w2097_,
		_w10965_,
		_w10976_,
		_w10977_
	);
	LUT2 #(
		.INIT('h8)
	) name9077 (
		\s15_data_i[23]_pad ,
		_w2057_,
		_w10978_
	);
	LUT4 #(
		.INIT('h135f)
	) name9078 (
		\s12_data_i[23]_pad ,
		\s13_data_i[23]_pad ,
		_w9457_,
		_w9629_,
		_w10979_
	);
	LUT4 #(
		.INIT('h153f)
	) name9079 (
		\s10_data_i[23]_pad ,
		\s1_data_i[23]_pad ,
		_w9288_,
		_w9451_,
		_w10980_
	);
	LUT4 #(
		.INIT('h135f)
	) name9080 (
		\s5_data_i[23]_pad ,
		\s6_data_i[23]_pad ,
		_w9471_,
		_w9474_,
		_w10981_
	);
	LUT4 #(
		.INIT('h135f)
	) name9081 (
		\s2_data_i[23]_pad ,
		\s7_data_i[23]_pad ,
		_w9462_,
		_w9626_,
		_w10982_
	);
	LUT4 #(
		.INIT('h8000)
	) name9082 (
		_w10979_,
		_w10980_,
		_w10981_,
		_w10982_,
		_w10983_
	);
	LUT2 #(
		.INIT('h8)
	) name9083 (
		\s14_data_i[23]_pad ,
		_w9632_,
		_w10984_
	);
	LUT4 #(
		.INIT('h135f)
	) name9084 (
		\s3_data_i[23]_pad ,
		\s4_data_i[23]_pad ,
		_w9465_,
		_w9468_,
		_w10985_
	);
	LUT4 #(
		.INIT('h135f)
	) name9085 (
		\s11_data_i[23]_pad ,
		\s8_data_i[23]_pad ,
		_w9454_,
		_w9620_,
		_w10986_
	);
	LUT4 #(
		.INIT('h135f)
	) name9086 (
		\s0_data_i[23]_pad ,
		\s9_data_i[23]_pad ,
		_w9284_,
		_w9477_,
		_w10987_
	);
	LUT4 #(
		.INIT('h4000)
	) name9087 (
		_w10984_,
		_w10985_,
		_w10986_,
		_w10987_,
		_w10988_
	);
	LUT2 #(
		.INIT('h8)
	) name9088 (
		_w10983_,
		_w10988_,
		_w10989_
	);
	LUT4 #(
		.INIT('h70ff)
	) name9089 (
		_w2046_,
		_w2097_,
		_w10978_,
		_w10989_,
		_w10990_
	);
	LUT2 #(
		.INIT('h8)
	) name9090 (
		\s15_data_i[24]_pad ,
		_w2057_,
		_w10991_
	);
	LUT4 #(
		.INIT('h135f)
	) name9091 (
		\s12_data_i[24]_pad ,
		\s13_data_i[24]_pad ,
		_w9457_,
		_w9629_,
		_w10992_
	);
	LUT4 #(
		.INIT('h153f)
	) name9092 (
		\s10_data_i[24]_pad ,
		\s1_data_i[24]_pad ,
		_w9288_,
		_w9451_,
		_w10993_
	);
	LUT4 #(
		.INIT('h135f)
	) name9093 (
		\s5_data_i[24]_pad ,
		\s6_data_i[24]_pad ,
		_w9471_,
		_w9474_,
		_w10994_
	);
	LUT4 #(
		.INIT('h135f)
	) name9094 (
		\s2_data_i[24]_pad ,
		\s7_data_i[24]_pad ,
		_w9462_,
		_w9626_,
		_w10995_
	);
	LUT4 #(
		.INIT('h8000)
	) name9095 (
		_w10992_,
		_w10993_,
		_w10994_,
		_w10995_,
		_w10996_
	);
	LUT2 #(
		.INIT('h8)
	) name9096 (
		\s14_data_i[24]_pad ,
		_w9632_,
		_w10997_
	);
	LUT4 #(
		.INIT('h135f)
	) name9097 (
		\s3_data_i[24]_pad ,
		\s4_data_i[24]_pad ,
		_w9465_,
		_w9468_,
		_w10998_
	);
	LUT4 #(
		.INIT('h135f)
	) name9098 (
		\s11_data_i[24]_pad ,
		\s8_data_i[24]_pad ,
		_w9454_,
		_w9620_,
		_w10999_
	);
	LUT4 #(
		.INIT('h135f)
	) name9099 (
		\s0_data_i[24]_pad ,
		\s9_data_i[24]_pad ,
		_w9284_,
		_w9477_,
		_w11000_
	);
	LUT4 #(
		.INIT('h4000)
	) name9100 (
		_w10997_,
		_w10998_,
		_w10999_,
		_w11000_,
		_w11001_
	);
	LUT2 #(
		.INIT('h8)
	) name9101 (
		_w10996_,
		_w11001_,
		_w11002_
	);
	LUT4 #(
		.INIT('h70ff)
	) name9102 (
		_w2046_,
		_w2097_,
		_w10991_,
		_w11002_,
		_w11003_
	);
	LUT2 #(
		.INIT('h8)
	) name9103 (
		\s15_data_i[25]_pad ,
		_w2057_,
		_w11004_
	);
	LUT4 #(
		.INIT('h135f)
	) name9104 (
		\s12_data_i[25]_pad ,
		\s13_data_i[25]_pad ,
		_w9457_,
		_w9629_,
		_w11005_
	);
	LUT4 #(
		.INIT('h153f)
	) name9105 (
		\s10_data_i[25]_pad ,
		\s1_data_i[25]_pad ,
		_w9288_,
		_w9451_,
		_w11006_
	);
	LUT4 #(
		.INIT('h135f)
	) name9106 (
		\s5_data_i[25]_pad ,
		\s6_data_i[25]_pad ,
		_w9471_,
		_w9474_,
		_w11007_
	);
	LUT4 #(
		.INIT('h135f)
	) name9107 (
		\s2_data_i[25]_pad ,
		\s7_data_i[25]_pad ,
		_w9462_,
		_w9626_,
		_w11008_
	);
	LUT4 #(
		.INIT('h8000)
	) name9108 (
		_w11005_,
		_w11006_,
		_w11007_,
		_w11008_,
		_w11009_
	);
	LUT2 #(
		.INIT('h8)
	) name9109 (
		\s14_data_i[25]_pad ,
		_w9632_,
		_w11010_
	);
	LUT4 #(
		.INIT('h135f)
	) name9110 (
		\s3_data_i[25]_pad ,
		\s4_data_i[25]_pad ,
		_w9465_,
		_w9468_,
		_w11011_
	);
	LUT4 #(
		.INIT('h135f)
	) name9111 (
		\s11_data_i[25]_pad ,
		\s8_data_i[25]_pad ,
		_w9454_,
		_w9620_,
		_w11012_
	);
	LUT4 #(
		.INIT('h135f)
	) name9112 (
		\s0_data_i[25]_pad ,
		\s9_data_i[25]_pad ,
		_w9284_,
		_w9477_,
		_w11013_
	);
	LUT4 #(
		.INIT('h4000)
	) name9113 (
		_w11010_,
		_w11011_,
		_w11012_,
		_w11013_,
		_w11014_
	);
	LUT2 #(
		.INIT('h8)
	) name9114 (
		_w11009_,
		_w11014_,
		_w11015_
	);
	LUT4 #(
		.INIT('h70ff)
	) name9115 (
		_w2046_,
		_w2097_,
		_w11004_,
		_w11015_,
		_w11016_
	);
	LUT2 #(
		.INIT('h8)
	) name9116 (
		\s15_data_i[26]_pad ,
		_w2057_,
		_w11017_
	);
	LUT4 #(
		.INIT('h135f)
	) name9117 (
		\s12_data_i[26]_pad ,
		\s13_data_i[26]_pad ,
		_w9457_,
		_w9629_,
		_w11018_
	);
	LUT4 #(
		.INIT('h153f)
	) name9118 (
		\s10_data_i[26]_pad ,
		\s1_data_i[26]_pad ,
		_w9288_,
		_w9451_,
		_w11019_
	);
	LUT4 #(
		.INIT('h135f)
	) name9119 (
		\s5_data_i[26]_pad ,
		\s6_data_i[26]_pad ,
		_w9471_,
		_w9474_,
		_w11020_
	);
	LUT4 #(
		.INIT('h135f)
	) name9120 (
		\s2_data_i[26]_pad ,
		\s7_data_i[26]_pad ,
		_w9462_,
		_w9626_,
		_w11021_
	);
	LUT4 #(
		.INIT('h8000)
	) name9121 (
		_w11018_,
		_w11019_,
		_w11020_,
		_w11021_,
		_w11022_
	);
	LUT2 #(
		.INIT('h8)
	) name9122 (
		\s14_data_i[26]_pad ,
		_w9632_,
		_w11023_
	);
	LUT4 #(
		.INIT('h135f)
	) name9123 (
		\s3_data_i[26]_pad ,
		\s4_data_i[26]_pad ,
		_w9465_,
		_w9468_,
		_w11024_
	);
	LUT4 #(
		.INIT('h135f)
	) name9124 (
		\s11_data_i[26]_pad ,
		\s8_data_i[26]_pad ,
		_w9454_,
		_w9620_,
		_w11025_
	);
	LUT4 #(
		.INIT('h135f)
	) name9125 (
		\s0_data_i[26]_pad ,
		\s9_data_i[26]_pad ,
		_w9284_,
		_w9477_,
		_w11026_
	);
	LUT4 #(
		.INIT('h4000)
	) name9126 (
		_w11023_,
		_w11024_,
		_w11025_,
		_w11026_,
		_w11027_
	);
	LUT2 #(
		.INIT('h8)
	) name9127 (
		_w11022_,
		_w11027_,
		_w11028_
	);
	LUT4 #(
		.INIT('h70ff)
	) name9128 (
		_w2046_,
		_w2097_,
		_w11017_,
		_w11028_,
		_w11029_
	);
	LUT2 #(
		.INIT('h8)
	) name9129 (
		\s15_data_i[27]_pad ,
		_w2057_,
		_w11030_
	);
	LUT4 #(
		.INIT('h135f)
	) name9130 (
		\s12_data_i[27]_pad ,
		\s13_data_i[27]_pad ,
		_w9457_,
		_w9629_,
		_w11031_
	);
	LUT4 #(
		.INIT('h153f)
	) name9131 (
		\s10_data_i[27]_pad ,
		\s1_data_i[27]_pad ,
		_w9288_,
		_w9451_,
		_w11032_
	);
	LUT4 #(
		.INIT('h135f)
	) name9132 (
		\s5_data_i[27]_pad ,
		\s6_data_i[27]_pad ,
		_w9471_,
		_w9474_,
		_w11033_
	);
	LUT4 #(
		.INIT('h135f)
	) name9133 (
		\s2_data_i[27]_pad ,
		\s7_data_i[27]_pad ,
		_w9462_,
		_w9626_,
		_w11034_
	);
	LUT4 #(
		.INIT('h8000)
	) name9134 (
		_w11031_,
		_w11032_,
		_w11033_,
		_w11034_,
		_w11035_
	);
	LUT2 #(
		.INIT('h8)
	) name9135 (
		\s14_data_i[27]_pad ,
		_w9632_,
		_w11036_
	);
	LUT4 #(
		.INIT('h135f)
	) name9136 (
		\s3_data_i[27]_pad ,
		\s4_data_i[27]_pad ,
		_w9465_,
		_w9468_,
		_w11037_
	);
	LUT4 #(
		.INIT('h135f)
	) name9137 (
		\s11_data_i[27]_pad ,
		\s8_data_i[27]_pad ,
		_w9454_,
		_w9620_,
		_w11038_
	);
	LUT4 #(
		.INIT('h135f)
	) name9138 (
		\s0_data_i[27]_pad ,
		\s9_data_i[27]_pad ,
		_w9284_,
		_w9477_,
		_w11039_
	);
	LUT4 #(
		.INIT('h4000)
	) name9139 (
		_w11036_,
		_w11037_,
		_w11038_,
		_w11039_,
		_w11040_
	);
	LUT2 #(
		.INIT('h8)
	) name9140 (
		_w11035_,
		_w11040_,
		_w11041_
	);
	LUT4 #(
		.INIT('h70ff)
	) name9141 (
		_w2046_,
		_w2097_,
		_w11030_,
		_w11041_,
		_w11042_
	);
	LUT2 #(
		.INIT('h8)
	) name9142 (
		\s15_data_i[28]_pad ,
		_w2057_,
		_w11043_
	);
	LUT4 #(
		.INIT('h135f)
	) name9143 (
		\s12_data_i[28]_pad ,
		\s13_data_i[28]_pad ,
		_w9457_,
		_w9629_,
		_w11044_
	);
	LUT4 #(
		.INIT('h153f)
	) name9144 (
		\s10_data_i[28]_pad ,
		\s1_data_i[28]_pad ,
		_w9288_,
		_w9451_,
		_w11045_
	);
	LUT4 #(
		.INIT('h135f)
	) name9145 (
		\s5_data_i[28]_pad ,
		\s6_data_i[28]_pad ,
		_w9471_,
		_w9474_,
		_w11046_
	);
	LUT4 #(
		.INIT('h135f)
	) name9146 (
		\s2_data_i[28]_pad ,
		\s7_data_i[28]_pad ,
		_w9462_,
		_w9626_,
		_w11047_
	);
	LUT4 #(
		.INIT('h8000)
	) name9147 (
		_w11044_,
		_w11045_,
		_w11046_,
		_w11047_,
		_w11048_
	);
	LUT2 #(
		.INIT('h8)
	) name9148 (
		\s14_data_i[28]_pad ,
		_w9632_,
		_w11049_
	);
	LUT4 #(
		.INIT('h135f)
	) name9149 (
		\s3_data_i[28]_pad ,
		\s4_data_i[28]_pad ,
		_w9465_,
		_w9468_,
		_w11050_
	);
	LUT4 #(
		.INIT('h135f)
	) name9150 (
		\s11_data_i[28]_pad ,
		\s8_data_i[28]_pad ,
		_w9454_,
		_w9620_,
		_w11051_
	);
	LUT4 #(
		.INIT('h135f)
	) name9151 (
		\s0_data_i[28]_pad ,
		\s9_data_i[28]_pad ,
		_w9284_,
		_w9477_,
		_w11052_
	);
	LUT4 #(
		.INIT('h4000)
	) name9152 (
		_w11049_,
		_w11050_,
		_w11051_,
		_w11052_,
		_w11053_
	);
	LUT2 #(
		.INIT('h8)
	) name9153 (
		_w11048_,
		_w11053_,
		_w11054_
	);
	LUT4 #(
		.INIT('h70ff)
	) name9154 (
		_w2046_,
		_w2097_,
		_w11043_,
		_w11054_,
		_w11055_
	);
	LUT2 #(
		.INIT('h8)
	) name9155 (
		\s15_data_i[29]_pad ,
		_w2057_,
		_w11056_
	);
	LUT4 #(
		.INIT('h135f)
	) name9156 (
		\s12_data_i[29]_pad ,
		\s13_data_i[29]_pad ,
		_w9457_,
		_w9629_,
		_w11057_
	);
	LUT4 #(
		.INIT('h153f)
	) name9157 (
		\s10_data_i[29]_pad ,
		\s1_data_i[29]_pad ,
		_w9288_,
		_w9451_,
		_w11058_
	);
	LUT4 #(
		.INIT('h135f)
	) name9158 (
		\s5_data_i[29]_pad ,
		\s6_data_i[29]_pad ,
		_w9471_,
		_w9474_,
		_w11059_
	);
	LUT4 #(
		.INIT('h135f)
	) name9159 (
		\s2_data_i[29]_pad ,
		\s7_data_i[29]_pad ,
		_w9462_,
		_w9626_,
		_w11060_
	);
	LUT4 #(
		.INIT('h8000)
	) name9160 (
		_w11057_,
		_w11058_,
		_w11059_,
		_w11060_,
		_w11061_
	);
	LUT2 #(
		.INIT('h8)
	) name9161 (
		\s14_data_i[29]_pad ,
		_w9632_,
		_w11062_
	);
	LUT4 #(
		.INIT('h135f)
	) name9162 (
		\s3_data_i[29]_pad ,
		\s4_data_i[29]_pad ,
		_w9465_,
		_w9468_,
		_w11063_
	);
	LUT4 #(
		.INIT('h135f)
	) name9163 (
		\s11_data_i[29]_pad ,
		\s8_data_i[29]_pad ,
		_w9454_,
		_w9620_,
		_w11064_
	);
	LUT4 #(
		.INIT('h135f)
	) name9164 (
		\s0_data_i[29]_pad ,
		\s9_data_i[29]_pad ,
		_w9284_,
		_w9477_,
		_w11065_
	);
	LUT4 #(
		.INIT('h4000)
	) name9165 (
		_w11062_,
		_w11063_,
		_w11064_,
		_w11065_,
		_w11066_
	);
	LUT2 #(
		.INIT('h8)
	) name9166 (
		_w11061_,
		_w11066_,
		_w11067_
	);
	LUT4 #(
		.INIT('h70ff)
	) name9167 (
		_w2046_,
		_w2097_,
		_w11056_,
		_w11067_,
		_w11068_
	);
	LUT3 #(
		.INIT('h80)
	) name9168 (
		_w2057_,
		_w2097_,
		_w9993_,
		_w11069_
	);
	LUT2 #(
		.INIT('h8)
	) name9169 (
		\s15_data_i[2]_pad ,
		_w2057_,
		_w11070_
	);
	LUT3 #(
		.INIT('h70)
	) name9170 (
		_w2046_,
		_w2097_,
		_w11070_,
		_w11071_
	);
	LUT4 #(
		.INIT('h135f)
	) name9171 (
		\s1_data_i[2]_pad ,
		\s8_data_i[2]_pad ,
		_w9288_,
		_w9620_,
		_w11072_
	);
	LUT4 #(
		.INIT('h135f)
	) name9172 (
		\s4_data_i[2]_pad ,
		\s6_data_i[2]_pad ,
		_w9468_,
		_w9474_,
		_w11073_
	);
	LUT4 #(
		.INIT('h135f)
	) name9173 (
		\s5_data_i[2]_pad ,
		\s9_data_i[2]_pad ,
		_w9471_,
		_w9477_,
		_w11074_
	);
	LUT4 #(
		.INIT('h135f)
	) name9174 (
		\s10_data_i[2]_pad ,
		\s7_data_i[2]_pad ,
		_w9451_,
		_w9626_,
		_w11075_
	);
	LUT4 #(
		.INIT('h8000)
	) name9175 (
		_w11072_,
		_w11073_,
		_w11074_,
		_w11075_,
		_w11076_
	);
	LUT2 #(
		.INIT('h8)
	) name9176 (
		\s11_data_i[2]_pad ,
		_w9454_,
		_w11077_
	);
	LUT4 #(
		.INIT('h153f)
	) name9177 (
		\s13_data_i[2]_pad ,
		\s3_data_i[2]_pad ,
		_w9465_,
		_w9629_,
		_w11078_
	);
	LUT4 #(
		.INIT('h135f)
	) name9178 (
		\s12_data_i[2]_pad ,
		\s14_data_i[2]_pad ,
		_w9457_,
		_w9632_,
		_w11079_
	);
	LUT4 #(
		.INIT('h135f)
	) name9179 (
		\s0_data_i[2]_pad ,
		\s2_data_i[2]_pad ,
		_w9284_,
		_w9462_,
		_w11080_
	);
	LUT4 #(
		.INIT('h4000)
	) name9180 (
		_w11077_,
		_w11078_,
		_w11079_,
		_w11080_,
		_w11081_
	);
	LUT2 #(
		.INIT('h8)
	) name9181 (
		_w11076_,
		_w11081_,
		_w11082_
	);
	LUT3 #(
		.INIT('hef)
	) name9182 (
		_w11069_,
		_w11071_,
		_w11082_,
		_w11083_
	);
	LUT2 #(
		.INIT('h8)
	) name9183 (
		\s15_data_i[30]_pad ,
		_w2057_,
		_w11084_
	);
	LUT4 #(
		.INIT('h135f)
	) name9184 (
		\s12_data_i[30]_pad ,
		\s13_data_i[30]_pad ,
		_w9457_,
		_w9629_,
		_w11085_
	);
	LUT4 #(
		.INIT('h153f)
	) name9185 (
		\s10_data_i[30]_pad ,
		\s1_data_i[30]_pad ,
		_w9288_,
		_w9451_,
		_w11086_
	);
	LUT4 #(
		.INIT('h135f)
	) name9186 (
		\s5_data_i[30]_pad ,
		\s6_data_i[30]_pad ,
		_w9471_,
		_w9474_,
		_w11087_
	);
	LUT4 #(
		.INIT('h135f)
	) name9187 (
		\s2_data_i[30]_pad ,
		\s7_data_i[30]_pad ,
		_w9462_,
		_w9626_,
		_w11088_
	);
	LUT4 #(
		.INIT('h8000)
	) name9188 (
		_w11085_,
		_w11086_,
		_w11087_,
		_w11088_,
		_w11089_
	);
	LUT2 #(
		.INIT('h8)
	) name9189 (
		\s14_data_i[30]_pad ,
		_w9632_,
		_w11090_
	);
	LUT4 #(
		.INIT('h135f)
	) name9190 (
		\s3_data_i[30]_pad ,
		\s4_data_i[30]_pad ,
		_w9465_,
		_w9468_,
		_w11091_
	);
	LUT4 #(
		.INIT('h135f)
	) name9191 (
		\s11_data_i[30]_pad ,
		\s8_data_i[30]_pad ,
		_w9454_,
		_w9620_,
		_w11092_
	);
	LUT4 #(
		.INIT('h135f)
	) name9192 (
		\s0_data_i[30]_pad ,
		\s9_data_i[30]_pad ,
		_w9284_,
		_w9477_,
		_w11093_
	);
	LUT4 #(
		.INIT('h4000)
	) name9193 (
		_w11090_,
		_w11091_,
		_w11092_,
		_w11093_,
		_w11094_
	);
	LUT2 #(
		.INIT('h8)
	) name9194 (
		_w11089_,
		_w11094_,
		_w11095_
	);
	LUT4 #(
		.INIT('h70ff)
	) name9195 (
		_w2046_,
		_w2097_,
		_w11084_,
		_w11095_,
		_w11096_
	);
	LUT2 #(
		.INIT('h8)
	) name9196 (
		\s15_data_i[31]_pad ,
		_w2057_,
		_w11097_
	);
	LUT4 #(
		.INIT('h135f)
	) name9197 (
		\s12_data_i[31]_pad ,
		\s13_data_i[31]_pad ,
		_w9457_,
		_w9629_,
		_w11098_
	);
	LUT4 #(
		.INIT('h153f)
	) name9198 (
		\s10_data_i[31]_pad ,
		\s1_data_i[31]_pad ,
		_w9288_,
		_w9451_,
		_w11099_
	);
	LUT4 #(
		.INIT('h135f)
	) name9199 (
		\s5_data_i[31]_pad ,
		\s6_data_i[31]_pad ,
		_w9471_,
		_w9474_,
		_w11100_
	);
	LUT4 #(
		.INIT('h135f)
	) name9200 (
		\s2_data_i[31]_pad ,
		\s7_data_i[31]_pad ,
		_w9462_,
		_w9626_,
		_w11101_
	);
	LUT4 #(
		.INIT('h8000)
	) name9201 (
		_w11098_,
		_w11099_,
		_w11100_,
		_w11101_,
		_w11102_
	);
	LUT2 #(
		.INIT('h8)
	) name9202 (
		\s14_data_i[31]_pad ,
		_w9632_,
		_w11103_
	);
	LUT4 #(
		.INIT('h135f)
	) name9203 (
		\s3_data_i[31]_pad ,
		\s4_data_i[31]_pad ,
		_w9465_,
		_w9468_,
		_w11104_
	);
	LUT4 #(
		.INIT('h135f)
	) name9204 (
		\s11_data_i[31]_pad ,
		\s8_data_i[31]_pad ,
		_w9454_,
		_w9620_,
		_w11105_
	);
	LUT4 #(
		.INIT('h135f)
	) name9205 (
		\s0_data_i[31]_pad ,
		\s9_data_i[31]_pad ,
		_w9284_,
		_w9477_,
		_w11106_
	);
	LUT4 #(
		.INIT('h4000)
	) name9206 (
		_w11103_,
		_w11104_,
		_w11105_,
		_w11106_,
		_w11107_
	);
	LUT2 #(
		.INIT('h8)
	) name9207 (
		_w11102_,
		_w11107_,
		_w11108_
	);
	LUT4 #(
		.INIT('h70ff)
	) name9208 (
		_w2046_,
		_w2097_,
		_w11097_,
		_w11108_,
		_w11109_
	);
	LUT3 #(
		.INIT('h80)
	) name9209 (
		_w2057_,
		_w2097_,
		_w10035_,
		_w11110_
	);
	LUT2 #(
		.INIT('h8)
	) name9210 (
		\s15_data_i[3]_pad ,
		_w2057_,
		_w11111_
	);
	LUT3 #(
		.INIT('h70)
	) name9211 (
		_w2046_,
		_w2097_,
		_w11111_,
		_w11112_
	);
	LUT4 #(
		.INIT('h153f)
	) name9212 (
		\s13_data_i[3]_pad ,
		\s8_data_i[3]_pad ,
		_w9620_,
		_w9629_,
		_w11113_
	);
	LUT4 #(
		.INIT('h153f)
	) name9213 (
		\s10_data_i[3]_pad ,
		\s1_data_i[3]_pad ,
		_w9288_,
		_w9451_,
		_w11114_
	);
	LUT4 #(
		.INIT('h135f)
	) name9214 (
		\s5_data_i[3]_pad ,
		\s6_data_i[3]_pad ,
		_w9471_,
		_w9474_,
		_w11115_
	);
	LUT4 #(
		.INIT('h135f)
	) name9215 (
		\s2_data_i[3]_pad ,
		\s7_data_i[3]_pad ,
		_w9462_,
		_w9626_,
		_w11116_
	);
	LUT4 #(
		.INIT('h8000)
	) name9216 (
		_w11113_,
		_w11114_,
		_w11115_,
		_w11116_,
		_w11117_
	);
	LUT2 #(
		.INIT('h8)
	) name9217 (
		\s11_data_i[3]_pad ,
		_w9454_,
		_w11118_
	);
	LUT4 #(
		.INIT('h135f)
	) name9218 (
		\s3_data_i[3]_pad ,
		\s4_data_i[3]_pad ,
		_w9465_,
		_w9468_,
		_w11119_
	);
	LUT4 #(
		.INIT('h135f)
	) name9219 (
		\s12_data_i[3]_pad ,
		\s14_data_i[3]_pad ,
		_w9457_,
		_w9632_,
		_w11120_
	);
	LUT4 #(
		.INIT('h135f)
	) name9220 (
		\s0_data_i[3]_pad ,
		\s9_data_i[3]_pad ,
		_w9284_,
		_w9477_,
		_w11121_
	);
	LUT4 #(
		.INIT('h4000)
	) name9221 (
		_w11118_,
		_w11119_,
		_w11120_,
		_w11121_,
		_w11122_
	);
	LUT2 #(
		.INIT('h8)
	) name9222 (
		_w11117_,
		_w11122_,
		_w11123_
	);
	LUT3 #(
		.INIT('hef)
	) name9223 (
		_w11110_,
		_w11112_,
		_w11123_,
		_w11124_
	);
	LUT3 #(
		.INIT('h80)
	) name9224 (
		_w2057_,
		_w2097_,
		_w10051_,
		_w11125_
	);
	LUT2 #(
		.INIT('h8)
	) name9225 (
		\s15_data_i[4]_pad ,
		_w2057_,
		_w11126_
	);
	LUT3 #(
		.INIT('h70)
	) name9226 (
		_w2046_,
		_w2097_,
		_w11126_,
		_w11127_
	);
	LUT4 #(
		.INIT('h153f)
	) name9227 (
		\s13_data_i[4]_pad ,
		\s2_data_i[4]_pad ,
		_w9462_,
		_w9629_,
		_w11128_
	);
	LUT4 #(
		.INIT('h135f)
	) name9228 (
		\s3_data_i[4]_pad ,
		\s7_data_i[4]_pad ,
		_w9465_,
		_w9626_,
		_w11129_
	);
	LUT4 #(
		.INIT('h135f)
	) name9229 (
		\s11_data_i[4]_pad ,
		\s5_data_i[4]_pad ,
		_w9454_,
		_w9471_,
		_w11130_
	);
	LUT4 #(
		.INIT('h153f)
	) name9230 (
		\s14_data_i[4]_pad ,
		\s8_data_i[4]_pad ,
		_w9620_,
		_w9632_,
		_w11131_
	);
	LUT4 #(
		.INIT('h8000)
	) name9231 (
		_w11128_,
		_w11129_,
		_w11130_,
		_w11131_,
		_w11132_
	);
	LUT2 #(
		.INIT('h8)
	) name9232 (
		\s1_data_i[4]_pad ,
		_w9288_,
		_w11133_
	);
	LUT4 #(
		.INIT('h135f)
	) name9233 (
		\s12_data_i[4]_pad ,
		\s4_data_i[4]_pad ,
		_w9457_,
		_w9468_,
		_w11134_
	);
	LUT4 #(
		.INIT('h135f)
	) name9234 (
		\s10_data_i[4]_pad ,
		\s9_data_i[4]_pad ,
		_w9451_,
		_w9477_,
		_w11135_
	);
	LUT4 #(
		.INIT('h135f)
	) name9235 (
		\s0_data_i[4]_pad ,
		\s6_data_i[4]_pad ,
		_w9284_,
		_w9474_,
		_w11136_
	);
	LUT4 #(
		.INIT('h4000)
	) name9236 (
		_w11133_,
		_w11134_,
		_w11135_,
		_w11136_,
		_w11137_
	);
	LUT2 #(
		.INIT('h8)
	) name9237 (
		_w11132_,
		_w11137_,
		_w11138_
	);
	LUT3 #(
		.INIT('hef)
	) name9238 (
		_w11125_,
		_w11127_,
		_w11138_,
		_w11139_
	);
	LUT3 #(
		.INIT('h80)
	) name9239 (
		_w2057_,
		_w2097_,
		_w10067_,
		_w11140_
	);
	LUT2 #(
		.INIT('h8)
	) name9240 (
		\s15_data_i[5]_pad ,
		_w2057_,
		_w11141_
	);
	LUT3 #(
		.INIT('h70)
	) name9241 (
		_w2046_,
		_w2097_,
		_w11141_,
		_w11142_
	);
	LUT4 #(
		.INIT('h153f)
	) name9242 (
		\s13_data_i[5]_pad ,
		\s8_data_i[5]_pad ,
		_w9620_,
		_w9629_,
		_w11143_
	);
	LUT4 #(
		.INIT('h153f)
	) name9243 (
		\s10_data_i[5]_pad ,
		\s1_data_i[5]_pad ,
		_w9288_,
		_w9451_,
		_w11144_
	);
	LUT4 #(
		.INIT('h135f)
	) name9244 (
		\s5_data_i[5]_pad ,
		\s6_data_i[5]_pad ,
		_w9471_,
		_w9474_,
		_w11145_
	);
	LUT4 #(
		.INIT('h135f)
	) name9245 (
		\s2_data_i[5]_pad ,
		\s7_data_i[5]_pad ,
		_w9462_,
		_w9626_,
		_w11146_
	);
	LUT4 #(
		.INIT('h8000)
	) name9246 (
		_w11143_,
		_w11144_,
		_w11145_,
		_w11146_,
		_w11147_
	);
	LUT2 #(
		.INIT('h8)
	) name9247 (
		\s11_data_i[5]_pad ,
		_w9454_,
		_w11148_
	);
	LUT4 #(
		.INIT('h135f)
	) name9248 (
		\s3_data_i[5]_pad ,
		\s4_data_i[5]_pad ,
		_w9465_,
		_w9468_,
		_w11149_
	);
	LUT4 #(
		.INIT('h135f)
	) name9249 (
		\s12_data_i[5]_pad ,
		\s14_data_i[5]_pad ,
		_w9457_,
		_w9632_,
		_w11150_
	);
	LUT4 #(
		.INIT('h135f)
	) name9250 (
		\s0_data_i[5]_pad ,
		\s9_data_i[5]_pad ,
		_w9284_,
		_w9477_,
		_w11151_
	);
	LUT4 #(
		.INIT('h4000)
	) name9251 (
		_w11148_,
		_w11149_,
		_w11150_,
		_w11151_,
		_w11152_
	);
	LUT2 #(
		.INIT('h8)
	) name9252 (
		_w11147_,
		_w11152_,
		_w11153_
	);
	LUT3 #(
		.INIT('hef)
	) name9253 (
		_w11140_,
		_w11142_,
		_w11153_,
		_w11154_
	);
	LUT3 #(
		.INIT('h80)
	) name9254 (
		_w2057_,
		_w2097_,
		_w10083_,
		_w11155_
	);
	LUT2 #(
		.INIT('h8)
	) name9255 (
		\s15_data_i[6]_pad ,
		_w2057_,
		_w11156_
	);
	LUT3 #(
		.INIT('h70)
	) name9256 (
		_w2046_,
		_w2097_,
		_w11156_,
		_w11157_
	);
	LUT4 #(
		.INIT('h153f)
	) name9257 (
		\s13_data_i[6]_pad ,
		\s8_data_i[6]_pad ,
		_w9620_,
		_w9629_,
		_w11158_
	);
	LUT4 #(
		.INIT('h153f)
	) name9258 (
		\s10_data_i[6]_pad ,
		\s1_data_i[6]_pad ,
		_w9288_,
		_w9451_,
		_w11159_
	);
	LUT4 #(
		.INIT('h135f)
	) name9259 (
		\s5_data_i[6]_pad ,
		\s6_data_i[6]_pad ,
		_w9471_,
		_w9474_,
		_w11160_
	);
	LUT4 #(
		.INIT('h135f)
	) name9260 (
		\s2_data_i[6]_pad ,
		\s7_data_i[6]_pad ,
		_w9462_,
		_w9626_,
		_w11161_
	);
	LUT4 #(
		.INIT('h8000)
	) name9261 (
		_w11158_,
		_w11159_,
		_w11160_,
		_w11161_,
		_w11162_
	);
	LUT2 #(
		.INIT('h8)
	) name9262 (
		\s11_data_i[6]_pad ,
		_w9454_,
		_w11163_
	);
	LUT4 #(
		.INIT('h135f)
	) name9263 (
		\s3_data_i[6]_pad ,
		\s4_data_i[6]_pad ,
		_w9465_,
		_w9468_,
		_w11164_
	);
	LUT4 #(
		.INIT('h135f)
	) name9264 (
		\s12_data_i[6]_pad ,
		\s14_data_i[6]_pad ,
		_w9457_,
		_w9632_,
		_w11165_
	);
	LUT4 #(
		.INIT('h135f)
	) name9265 (
		\s0_data_i[6]_pad ,
		\s9_data_i[6]_pad ,
		_w9284_,
		_w9477_,
		_w11166_
	);
	LUT4 #(
		.INIT('h4000)
	) name9266 (
		_w11163_,
		_w11164_,
		_w11165_,
		_w11166_,
		_w11167_
	);
	LUT2 #(
		.INIT('h8)
	) name9267 (
		_w11162_,
		_w11167_,
		_w11168_
	);
	LUT3 #(
		.INIT('hef)
	) name9268 (
		_w11155_,
		_w11157_,
		_w11168_,
		_w11169_
	);
	LUT3 #(
		.INIT('h80)
	) name9269 (
		_w2057_,
		_w2097_,
		_w10099_,
		_w11170_
	);
	LUT2 #(
		.INIT('h8)
	) name9270 (
		\s15_data_i[7]_pad ,
		_w2057_,
		_w11171_
	);
	LUT3 #(
		.INIT('h70)
	) name9271 (
		_w2046_,
		_w2097_,
		_w11171_,
		_w11172_
	);
	LUT4 #(
		.INIT('h153f)
	) name9272 (
		\s13_data_i[7]_pad ,
		\s2_data_i[7]_pad ,
		_w9462_,
		_w9629_,
		_w11173_
	);
	LUT4 #(
		.INIT('h135f)
	) name9273 (
		\s3_data_i[7]_pad ,
		\s7_data_i[7]_pad ,
		_w9465_,
		_w9626_,
		_w11174_
	);
	LUT4 #(
		.INIT('h135f)
	) name9274 (
		\s11_data_i[7]_pad ,
		\s5_data_i[7]_pad ,
		_w9454_,
		_w9471_,
		_w11175_
	);
	LUT4 #(
		.INIT('h153f)
	) name9275 (
		\s14_data_i[7]_pad ,
		\s8_data_i[7]_pad ,
		_w9620_,
		_w9632_,
		_w11176_
	);
	LUT4 #(
		.INIT('h8000)
	) name9276 (
		_w11173_,
		_w11174_,
		_w11175_,
		_w11176_,
		_w11177_
	);
	LUT2 #(
		.INIT('h8)
	) name9277 (
		\s1_data_i[7]_pad ,
		_w9288_,
		_w11178_
	);
	LUT4 #(
		.INIT('h135f)
	) name9278 (
		\s12_data_i[7]_pad ,
		\s4_data_i[7]_pad ,
		_w9457_,
		_w9468_,
		_w11179_
	);
	LUT4 #(
		.INIT('h135f)
	) name9279 (
		\s10_data_i[7]_pad ,
		\s9_data_i[7]_pad ,
		_w9451_,
		_w9477_,
		_w11180_
	);
	LUT4 #(
		.INIT('h135f)
	) name9280 (
		\s0_data_i[7]_pad ,
		\s6_data_i[7]_pad ,
		_w9284_,
		_w9474_,
		_w11181_
	);
	LUT4 #(
		.INIT('h4000)
	) name9281 (
		_w11178_,
		_w11179_,
		_w11180_,
		_w11181_,
		_w11182_
	);
	LUT2 #(
		.INIT('h8)
	) name9282 (
		_w11177_,
		_w11182_,
		_w11183_
	);
	LUT3 #(
		.INIT('hef)
	) name9283 (
		_w11170_,
		_w11172_,
		_w11183_,
		_w11184_
	);
	LUT3 #(
		.INIT('h80)
	) name9284 (
		_w2057_,
		_w2097_,
		_w10115_,
		_w11185_
	);
	LUT2 #(
		.INIT('h8)
	) name9285 (
		\s15_data_i[8]_pad ,
		_w2057_,
		_w11186_
	);
	LUT3 #(
		.INIT('h70)
	) name9286 (
		_w2046_,
		_w2097_,
		_w11186_,
		_w11187_
	);
	LUT4 #(
		.INIT('h153f)
	) name9287 (
		\s13_data_i[8]_pad ,
		\s8_data_i[8]_pad ,
		_w9620_,
		_w9629_,
		_w11188_
	);
	LUT4 #(
		.INIT('h153f)
	) name9288 (
		\s10_data_i[8]_pad ,
		\s1_data_i[8]_pad ,
		_w9288_,
		_w9451_,
		_w11189_
	);
	LUT4 #(
		.INIT('h135f)
	) name9289 (
		\s5_data_i[8]_pad ,
		\s6_data_i[8]_pad ,
		_w9471_,
		_w9474_,
		_w11190_
	);
	LUT4 #(
		.INIT('h135f)
	) name9290 (
		\s2_data_i[8]_pad ,
		\s7_data_i[8]_pad ,
		_w9462_,
		_w9626_,
		_w11191_
	);
	LUT4 #(
		.INIT('h8000)
	) name9291 (
		_w11188_,
		_w11189_,
		_w11190_,
		_w11191_,
		_w11192_
	);
	LUT2 #(
		.INIT('h8)
	) name9292 (
		\s11_data_i[8]_pad ,
		_w9454_,
		_w11193_
	);
	LUT4 #(
		.INIT('h135f)
	) name9293 (
		\s3_data_i[8]_pad ,
		\s4_data_i[8]_pad ,
		_w9465_,
		_w9468_,
		_w11194_
	);
	LUT4 #(
		.INIT('h135f)
	) name9294 (
		\s12_data_i[8]_pad ,
		\s14_data_i[8]_pad ,
		_w9457_,
		_w9632_,
		_w11195_
	);
	LUT4 #(
		.INIT('h135f)
	) name9295 (
		\s0_data_i[8]_pad ,
		\s9_data_i[8]_pad ,
		_w9284_,
		_w9477_,
		_w11196_
	);
	LUT4 #(
		.INIT('h4000)
	) name9296 (
		_w11193_,
		_w11194_,
		_w11195_,
		_w11196_,
		_w11197_
	);
	LUT2 #(
		.INIT('h8)
	) name9297 (
		_w11192_,
		_w11197_,
		_w11198_
	);
	LUT3 #(
		.INIT('hef)
	) name9298 (
		_w11185_,
		_w11187_,
		_w11198_,
		_w11199_
	);
	LUT3 #(
		.INIT('h80)
	) name9299 (
		_w2057_,
		_w2097_,
		_w10131_,
		_w11200_
	);
	LUT2 #(
		.INIT('h8)
	) name9300 (
		\s15_data_i[9]_pad ,
		_w2057_,
		_w11201_
	);
	LUT3 #(
		.INIT('h70)
	) name9301 (
		_w2046_,
		_w2097_,
		_w11201_,
		_w11202_
	);
	LUT4 #(
		.INIT('h153f)
	) name9302 (
		\s13_data_i[9]_pad ,
		\s2_data_i[9]_pad ,
		_w9462_,
		_w9629_,
		_w11203_
	);
	LUT4 #(
		.INIT('h135f)
	) name9303 (
		\s3_data_i[9]_pad ,
		\s7_data_i[9]_pad ,
		_w9465_,
		_w9626_,
		_w11204_
	);
	LUT4 #(
		.INIT('h135f)
	) name9304 (
		\s11_data_i[9]_pad ,
		\s5_data_i[9]_pad ,
		_w9454_,
		_w9471_,
		_w11205_
	);
	LUT4 #(
		.INIT('h153f)
	) name9305 (
		\s14_data_i[9]_pad ,
		\s8_data_i[9]_pad ,
		_w9620_,
		_w9632_,
		_w11206_
	);
	LUT4 #(
		.INIT('h8000)
	) name9306 (
		_w11203_,
		_w11204_,
		_w11205_,
		_w11206_,
		_w11207_
	);
	LUT2 #(
		.INIT('h8)
	) name9307 (
		\s1_data_i[9]_pad ,
		_w9288_,
		_w11208_
	);
	LUT4 #(
		.INIT('h135f)
	) name9308 (
		\s12_data_i[9]_pad ,
		\s4_data_i[9]_pad ,
		_w9457_,
		_w9468_,
		_w11209_
	);
	LUT4 #(
		.INIT('h135f)
	) name9309 (
		\s10_data_i[9]_pad ,
		\s9_data_i[9]_pad ,
		_w9451_,
		_w9477_,
		_w11210_
	);
	LUT4 #(
		.INIT('h135f)
	) name9310 (
		\s0_data_i[9]_pad ,
		\s6_data_i[9]_pad ,
		_w9284_,
		_w9474_,
		_w11211_
	);
	LUT4 #(
		.INIT('h4000)
	) name9311 (
		_w11208_,
		_w11209_,
		_w11210_,
		_w11211_,
		_w11212_
	);
	LUT2 #(
		.INIT('h8)
	) name9312 (
		_w11207_,
		_w11212_,
		_w11213_
	);
	LUT3 #(
		.INIT('hef)
	) name9313 (
		_w11200_,
		_w11202_,
		_w11213_,
		_w11214_
	);
	LUT3 #(
		.INIT('h80)
	) name9314 (
		\s15_err_i_pad ,
		_w1914_,
		_w10737_,
		_w11215_
	);
	LUT4 #(
		.INIT('h8000)
	) name9315 (
		\s11_err_i_pad ,
		_w8955_,
		_w8956_,
		_w9454_,
		_w11216_
	);
	LUT4 #(
		.INIT('h8000)
	) name9316 (
		\s3_err_i_pad ,
		_w9205_,
		_w9206_,
		_w9465_,
		_w11217_
	);
	LUT4 #(
		.INIT('h135f)
	) name9317 (
		_w8974_,
		_w9212_,
		_w11216_,
		_w11217_,
		_w11218_
	);
	LUT4 #(
		.INIT('h8000)
	) name9318 (
		\s9_err_i_pad ,
		_w8865_,
		_w8866_,
		_w9477_,
		_w11219_
	);
	LUT4 #(
		.INIT('h8000)
	) name9319 (
		\s0_err_i_pad ,
		_w8989_,
		_w8990_,
		_w9284_,
		_w11220_
	);
	LUT4 #(
		.INIT('h135f)
	) name9320 (
		_w8864_,
		_w9002_,
		_w11219_,
		_w11220_,
		_w11221_
	);
	LUT4 #(
		.INIT('h8000)
	) name9321 (
		\s6_err_i_pad ,
		_w8743_,
		_w8744_,
		_w9474_,
		_w11222_
	);
	LUT4 #(
		.INIT('h8000)
	) name9322 (
		\s10_err_i_pad ,
		_w8910_,
		_w8911_,
		_w9451_,
		_w11223_
	);
	LUT4 #(
		.INIT('h135f)
	) name9323 (
		_w8750_,
		_w8909_,
		_w11222_,
		_w11223_,
		_w11224_
	);
	LUT4 #(
		.INIT('h8000)
	) name9324 (
		\s4_err_i_pad ,
		_w8655_,
		_w8656_,
		_w9468_,
		_w11225_
	);
	LUT4 #(
		.INIT('h8000)
	) name9325 (
		\s13_err_i_pad ,
		_w9069_,
		_w9070_,
		_w9629_,
		_w11226_
	);
	LUT4 #(
		.INIT('h135f)
	) name9326 (
		_w8668_,
		_w9082_,
		_w11225_,
		_w11226_,
		_w11227_
	);
	LUT4 #(
		.INIT('h8000)
	) name9327 (
		_w11218_,
		_w11221_,
		_w11224_,
		_w11227_,
		_w11228_
	);
	LUT4 #(
		.INIT('h8000)
	) name9328 (
		\s8_err_i_pad ,
		_w8821_,
		_w8822_,
		_w9620_,
		_w11229_
	);
	LUT2 #(
		.INIT('h8)
	) name9329 (
		_w8828_,
		_w11229_,
		_w11230_
	);
	LUT4 #(
		.INIT('h8000)
	) name9330 (
		\s2_err_i_pad ,
		_w9171_,
		_w9172_,
		_w9462_,
		_w11231_
	);
	LUT4 #(
		.INIT('h8000)
	) name9331 (
		\s7_err_i_pad ,
		_w8782_,
		_w8783_,
		_w9626_,
		_w11232_
	);
	LUT4 #(
		.INIT('h153f)
	) name9332 (
		_w8795_,
		_w9190_,
		_w11231_,
		_w11232_,
		_w11233_
	);
	LUT4 #(
		.INIT('h8000)
	) name9333 (
		\s12_err_i_pad ,
		_w9029_,
		_w9030_,
		_w9457_,
		_w11234_
	);
	LUT4 #(
		.INIT('h8000)
	) name9334 (
		\s14_err_i_pad ,
		_w9137_,
		_w9138_,
		_w9632_,
		_w11235_
	);
	LUT4 #(
		.INIT('h135f)
	) name9335 (
		_w9028_,
		_w9144_,
		_w11234_,
		_w11235_,
		_w11236_
	);
	LUT4 #(
		.INIT('h8000)
	) name9336 (
		\s5_err_i_pad ,
		_w8699_,
		_w8700_,
		_w9471_,
		_w11237_
	);
	LUT4 #(
		.INIT('h8000)
	) name9337 (
		\s1_err_i_pad ,
		_w9103_,
		_w9104_,
		_w9288_,
		_w11238_
	);
	LUT4 #(
		.INIT('h135f)
	) name9338 (
		_w8698_,
		_w9110_,
		_w11237_,
		_w11238_,
		_w11239_
	);
	LUT4 #(
		.INIT('h4000)
	) name9339 (
		_w11230_,
		_w11233_,
		_w11236_,
		_w11239_,
		_w11240_
	);
	LUT2 #(
		.INIT('h8)
	) name9340 (
		_w11228_,
		_w11240_,
		_w11241_
	);
	LUT4 #(
		.INIT('h70ff)
	) name9341 (
		_w2046_,
		_w2097_,
		_w11215_,
		_w11241_,
		_w11242_
	);
	LUT3 #(
		.INIT('h80)
	) name9342 (
		\s15_rty_i_pad ,
		_w1914_,
		_w10737_,
		_w11243_
	);
	LUT4 #(
		.INIT('h8000)
	) name9343 (
		\s11_rty_i_pad ,
		_w8955_,
		_w8956_,
		_w9454_,
		_w11244_
	);
	LUT4 #(
		.INIT('h8000)
	) name9344 (
		\s3_rty_i_pad ,
		_w9205_,
		_w9206_,
		_w9465_,
		_w11245_
	);
	LUT4 #(
		.INIT('h135f)
	) name9345 (
		_w8974_,
		_w9212_,
		_w11244_,
		_w11245_,
		_w11246_
	);
	LUT4 #(
		.INIT('h8000)
	) name9346 (
		\s6_rty_i_pad ,
		_w8743_,
		_w8744_,
		_w9474_,
		_w11247_
	);
	LUT4 #(
		.INIT('h8000)
	) name9347 (
		\s0_rty_i_pad ,
		_w8989_,
		_w8990_,
		_w9284_,
		_w11248_
	);
	LUT4 #(
		.INIT('h135f)
	) name9348 (
		_w8750_,
		_w9002_,
		_w11247_,
		_w11248_,
		_w11249_
	);
	LUT4 #(
		.INIT('h8000)
	) name9349 (
		\s9_rty_i_pad ,
		_w8865_,
		_w8866_,
		_w9477_,
		_w11250_
	);
	LUT4 #(
		.INIT('h8000)
	) name9350 (
		\s7_rty_i_pad ,
		_w8782_,
		_w8783_,
		_w9626_,
		_w11251_
	);
	LUT4 #(
		.INIT('h153f)
	) name9351 (
		_w8795_,
		_w8864_,
		_w11250_,
		_w11251_,
		_w11252_
	);
	LUT4 #(
		.INIT('h8000)
	) name9352 (
		\s4_rty_i_pad ,
		_w8655_,
		_w8656_,
		_w9468_,
		_w11253_
	);
	LUT4 #(
		.INIT('h8000)
	) name9353 (
		\s13_rty_i_pad ,
		_w9069_,
		_w9070_,
		_w9629_,
		_w11254_
	);
	LUT4 #(
		.INIT('h135f)
	) name9354 (
		_w8668_,
		_w9082_,
		_w11253_,
		_w11254_,
		_w11255_
	);
	LUT4 #(
		.INIT('h8000)
	) name9355 (
		_w11246_,
		_w11249_,
		_w11252_,
		_w11255_,
		_w11256_
	);
	LUT4 #(
		.INIT('h8000)
	) name9356 (
		\s8_rty_i_pad ,
		_w8821_,
		_w8822_,
		_w9620_,
		_w11257_
	);
	LUT2 #(
		.INIT('h8)
	) name9357 (
		_w8828_,
		_w11257_,
		_w11258_
	);
	LUT4 #(
		.INIT('h8000)
	) name9358 (
		\s2_rty_i_pad ,
		_w9171_,
		_w9172_,
		_w9462_,
		_w11259_
	);
	LUT4 #(
		.INIT('h8000)
	) name9359 (
		\s10_rty_i_pad ,
		_w8910_,
		_w8911_,
		_w9451_,
		_w11260_
	);
	LUT4 #(
		.INIT('h153f)
	) name9360 (
		_w8909_,
		_w9190_,
		_w11259_,
		_w11260_,
		_w11261_
	);
	LUT4 #(
		.INIT('h8000)
	) name9361 (
		\s12_rty_i_pad ,
		_w9029_,
		_w9030_,
		_w9457_,
		_w11262_
	);
	LUT4 #(
		.INIT('h8000)
	) name9362 (
		\s14_rty_i_pad ,
		_w9137_,
		_w9138_,
		_w9632_,
		_w11263_
	);
	LUT4 #(
		.INIT('h135f)
	) name9363 (
		_w9028_,
		_w9144_,
		_w11262_,
		_w11263_,
		_w11264_
	);
	LUT4 #(
		.INIT('h8000)
	) name9364 (
		\s5_rty_i_pad ,
		_w8699_,
		_w8700_,
		_w9471_,
		_w11265_
	);
	LUT4 #(
		.INIT('h8000)
	) name9365 (
		\s1_rty_i_pad ,
		_w9103_,
		_w9104_,
		_w9288_,
		_w11266_
	);
	LUT4 #(
		.INIT('h135f)
	) name9366 (
		_w8698_,
		_w9110_,
		_w11265_,
		_w11266_,
		_w11267_
	);
	LUT4 #(
		.INIT('h4000)
	) name9367 (
		_w11258_,
		_w11261_,
		_w11264_,
		_w11267_,
		_w11268_
	);
	LUT2 #(
		.INIT('h8)
	) name9368 (
		_w11256_,
		_w11268_,
		_w11269_
	);
	LUT4 #(
		.INIT('h70ff)
	) name9369 (
		_w2046_,
		_w2097_,
		_w11243_,
		_w11269_,
		_w11270_
	);
	LUT3 #(
		.INIT('h80)
	) name9370 (
		_w1901_,
		_w1902_,
		_w2059_,
		_w11271_
	);
	LUT2 #(
		.INIT('h8)
	) name9371 (
		_w1918_,
		_w11271_,
		_w11272_
	);
	LUT3 #(
		.INIT('h70)
	) name9372 (
		_w2097_,
		_w8630_,
		_w11272_,
		_w11273_
	);
	LUT4 #(
		.INIT('h2a00)
	) name9373 (
		\s5_ack_i_pad ,
		_w8699_,
		_w8700_,
		_w9387_,
		_w11274_
	);
	LUT4 #(
		.INIT('h2a00)
	) name9374 (
		\s1_ack_i_pad ,
		_w9103_,
		_w9104_,
		_w9295_,
		_w11275_
	);
	LUT4 #(
		.INIT('h135f)
	) name9375 (
		_w8698_,
		_w9110_,
		_w11274_,
		_w11275_,
		_w11276_
	);
	LUT4 #(
		.INIT('h2a00)
	) name9376 (
		\s8_ack_i_pad ,
		_w8821_,
		_w8822_,
		_w9503_,
		_w11277_
	);
	LUT4 #(
		.INIT('h2a00)
	) name9377 (
		\s10_ack_i_pad ,
		_w8910_,
		_w8911_,
		_w9480_,
		_w11278_
	);
	LUT4 #(
		.INIT('h135f)
	) name9378 (
		_w8828_,
		_w8909_,
		_w11277_,
		_w11278_,
		_w11279_
	);
	LUT4 #(
		.INIT('h2a00)
	) name9379 (
		\s7_ack_i_pad ,
		_w8782_,
		_w8783_,
		_w9375_,
		_w11280_
	);
	LUT4 #(
		.INIT('h2a00)
	) name9380 (
		\s11_ack_i_pad ,
		_w8955_,
		_w8956_,
		_w9483_,
		_w11281_
	);
	LUT4 #(
		.INIT('h135f)
	) name9381 (
		_w8795_,
		_w8974_,
		_w11280_,
		_w11281_,
		_w11282_
	);
	LUT4 #(
		.INIT('h2a00)
	) name9382 (
		\s13_ack_i_pad ,
		_w9069_,
		_w9070_,
		_w9489_,
		_w11283_
	);
	LUT4 #(
		.INIT('h2a00)
	) name9383 (
		\s9_ack_i_pad ,
		_w8865_,
		_w8866_,
		_w9506_,
		_w11284_
	);
	LUT4 #(
		.INIT('h153f)
	) name9384 (
		_w8864_,
		_w9082_,
		_w11283_,
		_w11284_,
		_w11285_
	);
	LUT4 #(
		.INIT('h8000)
	) name9385 (
		_w11276_,
		_w11279_,
		_w11282_,
		_w11285_,
		_w11286_
	);
	LUT4 #(
		.INIT('h2a00)
	) name9386 (
		\s3_ack_i_pad ,
		_w9205_,
		_w9206_,
		_w9416_,
		_w11287_
	);
	LUT2 #(
		.INIT('h8)
	) name9387 (
		_w9212_,
		_w11287_,
		_w11288_
	);
	LUT4 #(
		.INIT('h2a00)
	) name9388 (
		\s14_ack_i_pad ,
		_w9137_,
		_w9138_,
		_w9497_,
		_w11289_
	);
	LUT4 #(
		.INIT('h2a00)
	) name9389 (
		\s6_ack_i_pad ,
		_w8743_,
		_w8744_,
		_w9378_,
		_w11290_
	);
	LUT4 #(
		.INIT('h153f)
	) name9390 (
		_w8750_,
		_w9144_,
		_w11289_,
		_w11290_,
		_w11291_
	);
	LUT4 #(
		.INIT('h2a00)
	) name9391 (
		\s4_ack_i_pad ,
		_w8655_,
		_w8656_,
		_w9500_,
		_w11292_
	);
	LUT4 #(
		.INIT('h2a00)
	) name9392 (
		\s0_ack_i_pad ,
		_w8989_,
		_w8990_,
		_w9291_,
		_w11293_
	);
	LUT4 #(
		.INIT('h135f)
	) name9393 (
		_w8668_,
		_w9002_,
		_w11292_,
		_w11293_,
		_w11294_
	);
	LUT4 #(
		.INIT('h2a00)
	) name9394 (
		\s2_ack_i_pad ,
		_w9171_,
		_w9172_,
		_w9494_,
		_w11295_
	);
	LUT4 #(
		.INIT('h2a00)
	) name9395 (
		\s12_ack_i_pad ,
		_w9029_,
		_w9030_,
		_w9486_,
		_w11296_
	);
	LUT4 #(
		.INIT('h153f)
	) name9396 (
		_w9028_,
		_w9190_,
		_w11295_,
		_w11296_,
		_w11297_
	);
	LUT4 #(
		.INIT('h4000)
	) name9397 (
		_w11288_,
		_w11291_,
		_w11294_,
		_w11297_,
		_w11298_
	);
	LUT2 #(
		.INIT('h8)
	) name9398 (
		_w11286_,
		_w11298_,
		_w11299_
	);
	LUT3 #(
		.INIT('h4f)
	) name9399 (
		_w9652_,
		_w11273_,
		_w11299_,
		_w11300_
	);
	LUT3 #(
		.INIT('h80)
	) name9400 (
		_w2059_,
		_w2097_,
		_w9683_,
		_w11301_
	);
	LUT2 #(
		.INIT('h8)
	) name9401 (
		\s15_data_i[0]_pad ,
		_w2059_,
		_w11302_
	);
	LUT3 #(
		.INIT('h70)
	) name9402 (
		_w2046_,
		_w2097_,
		_w11302_,
		_w11303_
	);
	LUT4 #(
		.INIT('h135f)
	) name9403 (
		\s1_data_i[0]_pad ,
		\s8_data_i[0]_pad ,
		_w9295_,
		_w9503_,
		_w11304_
	);
	LUT4 #(
		.INIT('h153f)
	) name9404 (
		\s4_data_i[0]_pad ,
		\s6_data_i[0]_pad ,
		_w9378_,
		_w9500_,
		_w11305_
	);
	LUT4 #(
		.INIT('h135f)
	) name9405 (
		\s5_data_i[0]_pad ,
		\s9_data_i[0]_pad ,
		_w9387_,
		_w9506_,
		_w11306_
	);
	LUT4 #(
		.INIT('h153f)
	) name9406 (
		\s10_data_i[0]_pad ,
		\s7_data_i[0]_pad ,
		_w9375_,
		_w9480_,
		_w11307_
	);
	LUT4 #(
		.INIT('h8000)
	) name9407 (
		_w11304_,
		_w11305_,
		_w11306_,
		_w11307_,
		_w11308_
	);
	LUT2 #(
		.INIT('h8)
	) name9408 (
		\s11_data_i[0]_pad ,
		_w9483_,
		_w11309_
	);
	LUT4 #(
		.INIT('h153f)
	) name9409 (
		\s13_data_i[0]_pad ,
		\s3_data_i[0]_pad ,
		_w9416_,
		_w9489_,
		_w11310_
	);
	LUT4 #(
		.INIT('h135f)
	) name9410 (
		\s12_data_i[0]_pad ,
		\s14_data_i[0]_pad ,
		_w9486_,
		_w9497_,
		_w11311_
	);
	LUT4 #(
		.INIT('h135f)
	) name9411 (
		\s0_data_i[0]_pad ,
		\s2_data_i[0]_pad ,
		_w9291_,
		_w9494_,
		_w11312_
	);
	LUT4 #(
		.INIT('h4000)
	) name9412 (
		_w11309_,
		_w11310_,
		_w11311_,
		_w11312_,
		_w11313_
	);
	LUT2 #(
		.INIT('h8)
	) name9413 (
		_w11308_,
		_w11313_,
		_w11314_
	);
	LUT3 #(
		.INIT('hef)
	) name9414 (
		_w11301_,
		_w11303_,
		_w11314_,
		_w11315_
	);
	LUT3 #(
		.INIT('h80)
	) name9415 (
		_w2059_,
		_w2097_,
		_w9699_,
		_w11316_
	);
	LUT2 #(
		.INIT('h8)
	) name9416 (
		\s15_data_i[10]_pad ,
		_w2059_,
		_w11317_
	);
	LUT3 #(
		.INIT('h70)
	) name9417 (
		_w2046_,
		_w2097_,
		_w11317_,
		_w11318_
	);
	LUT4 #(
		.INIT('h135f)
	) name9418 (
		\s13_data_i[10]_pad ,
		\s8_data_i[10]_pad ,
		_w9489_,
		_w9503_,
		_w11319_
	);
	LUT4 #(
		.INIT('h153f)
	) name9419 (
		\s10_data_i[10]_pad ,
		\s1_data_i[10]_pad ,
		_w9295_,
		_w9480_,
		_w11320_
	);
	LUT4 #(
		.INIT('h153f)
	) name9420 (
		\s5_data_i[10]_pad ,
		\s6_data_i[10]_pad ,
		_w9378_,
		_w9387_,
		_w11321_
	);
	LUT4 #(
		.INIT('h153f)
	) name9421 (
		\s2_data_i[10]_pad ,
		\s7_data_i[10]_pad ,
		_w9375_,
		_w9494_,
		_w11322_
	);
	LUT4 #(
		.INIT('h8000)
	) name9422 (
		_w11319_,
		_w11320_,
		_w11321_,
		_w11322_,
		_w11323_
	);
	LUT2 #(
		.INIT('h8)
	) name9423 (
		\s11_data_i[10]_pad ,
		_w9483_,
		_w11324_
	);
	LUT4 #(
		.INIT('h135f)
	) name9424 (
		\s3_data_i[10]_pad ,
		\s4_data_i[10]_pad ,
		_w9416_,
		_w9500_,
		_w11325_
	);
	LUT4 #(
		.INIT('h135f)
	) name9425 (
		\s12_data_i[10]_pad ,
		\s14_data_i[10]_pad ,
		_w9486_,
		_w9497_,
		_w11326_
	);
	LUT4 #(
		.INIT('h135f)
	) name9426 (
		\s0_data_i[10]_pad ,
		\s9_data_i[10]_pad ,
		_w9291_,
		_w9506_,
		_w11327_
	);
	LUT4 #(
		.INIT('h4000)
	) name9427 (
		_w11324_,
		_w11325_,
		_w11326_,
		_w11327_,
		_w11328_
	);
	LUT2 #(
		.INIT('h8)
	) name9428 (
		_w11323_,
		_w11328_,
		_w11329_
	);
	LUT3 #(
		.INIT('hef)
	) name9429 (
		_w11316_,
		_w11318_,
		_w11329_,
		_w11330_
	);
	LUT3 #(
		.INIT('h80)
	) name9430 (
		_w2059_,
		_w2097_,
		_w9715_,
		_w11331_
	);
	LUT2 #(
		.INIT('h8)
	) name9431 (
		\s15_data_i[11]_pad ,
		_w2059_,
		_w11332_
	);
	LUT3 #(
		.INIT('h70)
	) name9432 (
		_w2046_,
		_w2097_,
		_w11332_,
		_w11333_
	);
	LUT4 #(
		.INIT('h135f)
	) name9433 (
		\s13_data_i[11]_pad ,
		\s8_data_i[11]_pad ,
		_w9489_,
		_w9503_,
		_w11334_
	);
	LUT4 #(
		.INIT('h153f)
	) name9434 (
		\s10_data_i[11]_pad ,
		\s1_data_i[11]_pad ,
		_w9295_,
		_w9480_,
		_w11335_
	);
	LUT4 #(
		.INIT('h153f)
	) name9435 (
		\s5_data_i[11]_pad ,
		\s6_data_i[11]_pad ,
		_w9378_,
		_w9387_,
		_w11336_
	);
	LUT4 #(
		.INIT('h153f)
	) name9436 (
		\s2_data_i[11]_pad ,
		\s7_data_i[11]_pad ,
		_w9375_,
		_w9494_,
		_w11337_
	);
	LUT4 #(
		.INIT('h8000)
	) name9437 (
		_w11334_,
		_w11335_,
		_w11336_,
		_w11337_,
		_w11338_
	);
	LUT2 #(
		.INIT('h8)
	) name9438 (
		\s11_data_i[11]_pad ,
		_w9483_,
		_w11339_
	);
	LUT4 #(
		.INIT('h135f)
	) name9439 (
		\s3_data_i[11]_pad ,
		\s4_data_i[11]_pad ,
		_w9416_,
		_w9500_,
		_w11340_
	);
	LUT4 #(
		.INIT('h135f)
	) name9440 (
		\s12_data_i[11]_pad ,
		\s14_data_i[11]_pad ,
		_w9486_,
		_w9497_,
		_w11341_
	);
	LUT4 #(
		.INIT('h135f)
	) name9441 (
		\s0_data_i[11]_pad ,
		\s9_data_i[11]_pad ,
		_w9291_,
		_w9506_,
		_w11342_
	);
	LUT4 #(
		.INIT('h4000)
	) name9442 (
		_w11339_,
		_w11340_,
		_w11341_,
		_w11342_,
		_w11343_
	);
	LUT2 #(
		.INIT('h8)
	) name9443 (
		_w11338_,
		_w11343_,
		_w11344_
	);
	LUT3 #(
		.INIT('hef)
	) name9444 (
		_w11331_,
		_w11333_,
		_w11344_,
		_w11345_
	);
	LUT3 #(
		.INIT('h80)
	) name9445 (
		_w2059_,
		_w2097_,
		_w9731_,
		_w11346_
	);
	LUT2 #(
		.INIT('h8)
	) name9446 (
		\s15_data_i[12]_pad ,
		_w2059_,
		_w11347_
	);
	LUT3 #(
		.INIT('h70)
	) name9447 (
		_w2046_,
		_w2097_,
		_w11347_,
		_w11348_
	);
	LUT4 #(
		.INIT('h135f)
	) name9448 (
		\s13_data_i[12]_pad ,
		\s8_data_i[12]_pad ,
		_w9489_,
		_w9503_,
		_w11349_
	);
	LUT4 #(
		.INIT('h153f)
	) name9449 (
		\s10_data_i[12]_pad ,
		\s1_data_i[12]_pad ,
		_w9295_,
		_w9480_,
		_w11350_
	);
	LUT4 #(
		.INIT('h153f)
	) name9450 (
		\s5_data_i[12]_pad ,
		\s6_data_i[12]_pad ,
		_w9378_,
		_w9387_,
		_w11351_
	);
	LUT4 #(
		.INIT('h153f)
	) name9451 (
		\s2_data_i[12]_pad ,
		\s7_data_i[12]_pad ,
		_w9375_,
		_w9494_,
		_w11352_
	);
	LUT4 #(
		.INIT('h8000)
	) name9452 (
		_w11349_,
		_w11350_,
		_w11351_,
		_w11352_,
		_w11353_
	);
	LUT2 #(
		.INIT('h8)
	) name9453 (
		\s11_data_i[12]_pad ,
		_w9483_,
		_w11354_
	);
	LUT4 #(
		.INIT('h135f)
	) name9454 (
		\s3_data_i[12]_pad ,
		\s4_data_i[12]_pad ,
		_w9416_,
		_w9500_,
		_w11355_
	);
	LUT4 #(
		.INIT('h135f)
	) name9455 (
		\s12_data_i[12]_pad ,
		\s14_data_i[12]_pad ,
		_w9486_,
		_w9497_,
		_w11356_
	);
	LUT4 #(
		.INIT('h135f)
	) name9456 (
		\s0_data_i[12]_pad ,
		\s9_data_i[12]_pad ,
		_w9291_,
		_w9506_,
		_w11357_
	);
	LUT4 #(
		.INIT('h4000)
	) name9457 (
		_w11354_,
		_w11355_,
		_w11356_,
		_w11357_,
		_w11358_
	);
	LUT2 #(
		.INIT('h8)
	) name9458 (
		_w11353_,
		_w11358_,
		_w11359_
	);
	LUT3 #(
		.INIT('hef)
	) name9459 (
		_w11346_,
		_w11348_,
		_w11359_,
		_w11360_
	);
	LUT3 #(
		.INIT('h80)
	) name9460 (
		_w2059_,
		_w2097_,
		_w9747_,
		_w11361_
	);
	LUT2 #(
		.INIT('h8)
	) name9461 (
		\s15_data_i[13]_pad ,
		_w2059_,
		_w11362_
	);
	LUT3 #(
		.INIT('h70)
	) name9462 (
		_w2046_,
		_w2097_,
		_w11362_,
		_w11363_
	);
	LUT4 #(
		.INIT('h135f)
	) name9463 (
		\s1_data_i[13]_pad ,
		\s8_data_i[13]_pad ,
		_w9295_,
		_w9503_,
		_w11364_
	);
	LUT4 #(
		.INIT('h153f)
	) name9464 (
		\s4_data_i[13]_pad ,
		\s6_data_i[13]_pad ,
		_w9378_,
		_w9500_,
		_w11365_
	);
	LUT4 #(
		.INIT('h135f)
	) name9465 (
		\s5_data_i[13]_pad ,
		\s9_data_i[13]_pad ,
		_w9387_,
		_w9506_,
		_w11366_
	);
	LUT4 #(
		.INIT('h153f)
	) name9466 (
		\s10_data_i[13]_pad ,
		\s7_data_i[13]_pad ,
		_w9375_,
		_w9480_,
		_w11367_
	);
	LUT4 #(
		.INIT('h8000)
	) name9467 (
		_w11364_,
		_w11365_,
		_w11366_,
		_w11367_,
		_w11368_
	);
	LUT2 #(
		.INIT('h8)
	) name9468 (
		\s11_data_i[13]_pad ,
		_w9483_,
		_w11369_
	);
	LUT4 #(
		.INIT('h153f)
	) name9469 (
		\s13_data_i[13]_pad ,
		\s3_data_i[13]_pad ,
		_w9416_,
		_w9489_,
		_w11370_
	);
	LUT4 #(
		.INIT('h135f)
	) name9470 (
		\s12_data_i[13]_pad ,
		\s14_data_i[13]_pad ,
		_w9486_,
		_w9497_,
		_w11371_
	);
	LUT4 #(
		.INIT('h135f)
	) name9471 (
		\s0_data_i[13]_pad ,
		\s2_data_i[13]_pad ,
		_w9291_,
		_w9494_,
		_w11372_
	);
	LUT4 #(
		.INIT('h4000)
	) name9472 (
		_w11369_,
		_w11370_,
		_w11371_,
		_w11372_,
		_w11373_
	);
	LUT2 #(
		.INIT('h8)
	) name9473 (
		_w11368_,
		_w11373_,
		_w11374_
	);
	LUT3 #(
		.INIT('hef)
	) name9474 (
		_w11361_,
		_w11363_,
		_w11374_,
		_w11375_
	);
	LUT3 #(
		.INIT('h80)
	) name9475 (
		_w2059_,
		_w2097_,
		_w9763_,
		_w11376_
	);
	LUT2 #(
		.INIT('h8)
	) name9476 (
		\s15_data_i[14]_pad ,
		_w2059_,
		_w11377_
	);
	LUT3 #(
		.INIT('h70)
	) name9477 (
		_w2046_,
		_w2097_,
		_w11377_,
		_w11378_
	);
	LUT4 #(
		.INIT('h135f)
	) name9478 (
		\s4_data_i[14]_pad ,
		\s8_data_i[14]_pad ,
		_w9500_,
		_w9503_,
		_w11379_
	);
	LUT4 #(
		.INIT('h135f)
	) name9479 (
		\s1_data_i[14]_pad ,
		\s7_data_i[14]_pad ,
		_w9295_,
		_w9375_,
		_w11380_
	);
	LUT4 #(
		.INIT('h153f)
	) name9480 (
		\s5_data_i[14]_pad ,
		\s6_data_i[14]_pad ,
		_w9378_,
		_w9387_,
		_w11381_
	);
	LUT4 #(
		.INIT('h135f)
	) name9481 (
		\s13_data_i[14]_pad ,
		\s2_data_i[14]_pad ,
		_w9489_,
		_w9494_,
		_w11382_
	);
	LUT4 #(
		.INIT('h8000)
	) name9482 (
		_w11379_,
		_w11380_,
		_w11381_,
		_w11382_,
		_w11383_
	);
	LUT2 #(
		.INIT('h8)
	) name9483 (
		\s11_data_i[14]_pad ,
		_w9483_,
		_w11384_
	);
	LUT4 #(
		.INIT('h153f)
	) name9484 (
		\s10_data_i[14]_pad ,
		\s3_data_i[14]_pad ,
		_w9416_,
		_w9480_,
		_w11385_
	);
	LUT4 #(
		.INIT('h135f)
	) name9485 (
		\s12_data_i[14]_pad ,
		\s14_data_i[14]_pad ,
		_w9486_,
		_w9497_,
		_w11386_
	);
	LUT4 #(
		.INIT('h135f)
	) name9486 (
		\s0_data_i[14]_pad ,
		\s9_data_i[14]_pad ,
		_w9291_,
		_w9506_,
		_w11387_
	);
	LUT4 #(
		.INIT('h4000)
	) name9487 (
		_w11384_,
		_w11385_,
		_w11386_,
		_w11387_,
		_w11388_
	);
	LUT2 #(
		.INIT('h8)
	) name9488 (
		_w11383_,
		_w11388_,
		_w11389_
	);
	LUT3 #(
		.INIT('hef)
	) name9489 (
		_w11376_,
		_w11378_,
		_w11389_,
		_w11390_
	);
	LUT3 #(
		.INIT('h80)
	) name9490 (
		_w2059_,
		_w2097_,
		_w9779_,
		_w11391_
	);
	LUT2 #(
		.INIT('h8)
	) name9491 (
		\s15_data_i[15]_pad ,
		_w2059_,
		_w11392_
	);
	LUT3 #(
		.INIT('h70)
	) name9492 (
		_w2046_,
		_w2097_,
		_w11392_,
		_w11393_
	);
	LUT4 #(
		.INIT('h135f)
	) name9493 (
		\s1_data_i[15]_pad ,
		\s8_data_i[15]_pad ,
		_w9295_,
		_w9503_,
		_w11394_
	);
	LUT4 #(
		.INIT('h153f)
	) name9494 (
		\s4_data_i[15]_pad ,
		\s6_data_i[15]_pad ,
		_w9378_,
		_w9500_,
		_w11395_
	);
	LUT4 #(
		.INIT('h135f)
	) name9495 (
		\s5_data_i[15]_pad ,
		\s9_data_i[15]_pad ,
		_w9387_,
		_w9506_,
		_w11396_
	);
	LUT4 #(
		.INIT('h153f)
	) name9496 (
		\s10_data_i[15]_pad ,
		\s7_data_i[15]_pad ,
		_w9375_,
		_w9480_,
		_w11397_
	);
	LUT4 #(
		.INIT('h8000)
	) name9497 (
		_w11394_,
		_w11395_,
		_w11396_,
		_w11397_,
		_w11398_
	);
	LUT2 #(
		.INIT('h8)
	) name9498 (
		\s11_data_i[15]_pad ,
		_w9483_,
		_w11399_
	);
	LUT4 #(
		.INIT('h153f)
	) name9499 (
		\s13_data_i[15]_pad ,
		\s3_data_i[15]_pad ,
		_w9416_,
		_w9489_,
		_w11400_
	);
	LUT4 #(
		.INIT('h135f)
	) name9500 (
		\s12_data_i[15]_pad ,
		\s14_data_i[15]_pad ,
		_w9486_,
		_w9497_,
		_w11401_
	);
	LUT4 #(
		.INIT('h135f)
	) name9501 (
		\s0_data_i[15]_pad ,
		\s2_data_i[15]_pad ,
		_w9291_,
		_w9494_,
		_w11402_
	);
	LUT4 #(
		.INIT('h4000)
	) name9502 (
		_w11399_,
		_w11400_,
		_w11401_,
		_w11402_,
		_w11403_
	);
	LUT2 #(
		.INIT('h8)
	) name9503 (
		_w11398_,
		_w11403_,
		_w11404_
	);
	LUT3 #(
		.INIT('hef)
	) name9504 (
		_w11391_,
		_w11393_,
		_w11404_,
		_w11405_
	);
	LUT2 #(
		.INIT('h8)
	) name9505 (
		\s15_data_i[16]_pad ,
		_w2059_,
		_w11406_
	);
	LUT4 #(
		.INIT('h135f)
	) name9506 (
		\s12_data_i[16]_pad ,
		\s13_data_i[16]_pad ,
		_w9486_,
		_w9489_,
		_w11407_
	);
	LUT4 #(
		.INIT('h153f)
	) name9507 (
		\s10_data_i[16]_pad ,
		\s1_data_i[16]_pad ,
		_w9295_,
		_w9480_,
		_w11408_
	);
	LUT4 #(
		.INIT('h153f)
	) name9508 (
		\s5_data_i[16]_pad ,
		\s6_data_i[16]_pad ,
		_w9378_,
		_w9387_,
		_w11409_
	);
	LUT4 #(
		.INIT('h153f)
	) name9509 (
		\s2_data_i[16]_pad ,
		\s7_data_i[16]_pad ,
		_w9375_,
		_w9494_,
		_w11410_
	);
	LUT4 #(
		.INIT('h8000)
	) name9510 (
		_w11407_,
		_w11408_,
		_w11409_,
		_w11410_,
		_w11411_
	);
	LUT2 #(
		.INIT('h8)
	) name9511 (
		\s14_data_i[16]_pad ,
		_w9497_,
		_w11412_
	);
	LUT4 #(
		.INIT('h135f)
	) name9512 (
		\s3_data_i[16]_pad ,
		\s4_data_i[16]_pad ,
		_w9416_,
		_w9500_,
		_w11413_
	);
	LUT4 #(
		.INIT('h135f)
	) name9513 (
		\s11_data_i[16]_pad ,
		\s8_data_i[16]_pad ,
		_w9483_,
		_w9503_,
		_w11414_
	);
	LUT4 #(
		.INIT('h135f)
	) name9514 (
		\s0_data_i[16]_pad ,
		\s9_data_i[16]_pad ,
		_w9291_,
		_w9506_,
		_w11415_
	);
	LUT4 #(
		.INIT('h4000)
	) name9515 (
		_w11412_,
		_w11413_,
		_w11414_,
		_w11415_,
		_w11416_
	);
	LUT2 #(
		.INIT('h8)
	) name9516 (
		_w11411_,
		_w11416_,
		_w11417_
	);
	LUT4 #(
		.INIT('h70ff)
	) name9517 (
		_w2046_,
		_w2097_,
		_w11406_,
		_w11417_,
		_w11418_
	);
	LUT2 #(
		.INIT('h8)
	) name9518 (
		\s15_data_i[17]_pad ,
		_w2059_,
		_w11419_
	);
	LUT4 #(
		.INIT('h135f)
	) name9519 (
		\s12_data_i[17]_pad ,
		\s13_data_i[17]_pad ,
		_w9486_,
		_w9489_,
		_w11420_
	);
	LUT4 #(
		.INIT('h153f)
	) name9520 (
		\s10_data_i[17]_pad ,
		\s1_data_i[17]_pad ,
		_w9295_,
		_w9480_,
		_w11421_
	);
	LUT4 #(
		.INIT('h153f)
	) name9521 (
		\s5_data_i[17]_pad ,
		\s6_data_i[17]_pad ,
		_w9378_,
		_w9387_,
		_w11422_
	);
	LUT4 #(
		.INIT('h153f)
	) name9522 (
		\s2_data_i[17]_pad ,
		\s7_data_i[17]_pad ,
		_w9375_,
		_w9494_,
		_w11423_
	);
	LUT4 #(
		.INIT('h8000)
	) name9523 (
		_w11420_,
		_w11421_,
		_w11422_,
		_w11423_,
		_w11424_
	);
	LUT2 #(
		.INIT('h8)
	) name9524 (
		\s14_data_i[17]_pad ,
		_w9497_,
		_w11425_
	);
	LUT4 #(
		.INIT('h135f)
	) name9525 (
		\s3_data_i[17]_pad ,
		\s4_data_i[17]_pad ,
		_w9416_,
		_w9500_,
		_w11426_
	);
	LUT4 #(
		.INIT('h135f)
	) name9526 (
		\s11_data_i[17]_pad ,
		\s8_data_i[17]_pad ,
		_w9483_,
		_w9503_,
		_w11427_
	);
	LUT4 #(
		.INIT('h135f)
	) name9527 (
		\s0_data_i[17]_pad ,
		\s9_data_i[17]_pad ,
		_w9291_,
		_w9506_,
		_w11428_
	);
	LUT4 #(
		.INIT('h4000)
	) name9528 (
		_w11425_,
		_w11426_,
		_w11427_,
		_w11428_,
		_w11429_
	);
	LUT2 #(
		.INIT('h8)
	) name9529 (
		_w11424_,
		_w11429_,
		_w11430_
	);
	LUT4 #(
		.INIT('h70ff)
	) name9530 (
		_w2046_,
		_w2097_,
		_w11419_,
		_w11430_,
		_w11431_
	);
	LUT2 #(
		.INIT('h8)
	) name9531 (
		\s15_data_i[18]_pad ,
		_w2059_,
		_w11432_
	);
	LUT4 #(
		.INIT('h135f)
	) name9532 (
		\s12_data_i[18]_pad ,
		\s13_data_i[18]_pad ,
		_w9486_,
		_w9489_,
		_w11433_
	);
	LUT4 #(
		.INIT('h153f)
	) name9533 (
		\s10_data_i[18]_pad ,
		\s1_data_i[18]_pad ,
		_w9295_,
		_w9480_,
		_w11434_
	);
	LUT4 #(
		.INIT('h153f)
	) name9534 (
		\s5_data_i[18]_pad ,
		\s6_data_i[18]_pad ,
		_w9378_,
		_w9387_,
		_w11435_
	);
	LUT4 #(
		.INIT('h153f)
	) name9535 (
		\s2_data_i[18]_pad ,
		\s7_data_i[18]_pad ,
		_w9375_,
		_w9494_,
		_w11436_
	);
	LUT4 #(
		.INIT('h8000)
	) name9536 (
		_w11433_,
		_w11434_,
		_w11435_,
		_w11436_,
		_w11437_
	);
	LUT2 #(
		.INIT('h8)
	) name9537 (
		\s14_data_i[18]_pad ,
		_w9497_,
		_w11438_
	);
	LUT4 #(
		.INIT('h135f)
	) name9538 (
		\s3_data_i[18]_pad ,
		\s4_data_i[18]_pad ,
		_w9416_,
		_w9500_,
		_w11439_
	);
	LUT4 #(
		.INIT('h135f)
	) name9539 (
		\s11_data_i[18]_pad ,
		\s8_data_i[18]_pad ,
		_w9483_,
		_w9503_,
		_w11440_
	);
	LUT4 #(
		.INIT('h135f)
	) name9540 (
		\s0_data_i[18]_pad ,
		\s9_data_i[18]_pad ,
		_w9291_,
		_w9506_,
		_w11441_
	);
	LUT4 #(
		.INIT('h4000)
	) name9541 (
		_w11438_,
		_w11439_,
		_w11440_,
		_w11441_,
		_w11442_
	);
	LUT2 #(
		.INIT('h8)
	) name9542 (
		_w11437_,
		_w11442_,
		_w11443_
	);
	LUT4 #(
		.INIT('h70ff)
	) name9543 (
		_w2046_,
		_w2097_,
		_w11432_,
		_w11443_,
		_w11444_
	);
	LUT2 #(
		.INIT('h8)
	) name9544 (
		\s15_data_i[19]_pad ,
		_w2059_,
		_w11445_
	);
	LUT4 #(
		.INIT('h135f)
	) name9545 (
		\s12_data_i[19]_pad ,
		\s13_data_i[19]_pad ,
		_w9486_,
		_w9489_,
		_w11446_
	);
	LUT4 #(
		.INIT('h153f)
	) name9546 (
		\s10_data_i[19]_pad ,
		\s1_data_i[19]_pad ,
		_w9295_,
		_w9480_,
		_w11447_
	);
	LUT4 #(
		.INIT('h153f)
	) name9547 (
		\s5_data_i[19]_pad ,
		\s6_data_i[19]_pad ,
		_w9378_,
		_w9387_,
		_w11448_
	);
	LUT4 #(
		.INIT('h153f)
	) name9548 (
		\s2_data_i[19]_pad ,
		\s7_data_i[19]_pad ,
		_w9375_,
		_w9494_,
		_w11449_
	);
	LUT4 #(
		.INIT('h8000)
	) name9549 (
		_w11446_,
		_w11447_,
		_w11448_,
		_w11449_,
		_w11450_
	);
	LUT2 #(
		.INIT('h8)
	) name9550 (
		\s14_data_i[19]_pad ,
		_w9497_,
		_w11451_
	);
	LUT4 #(
		.INIT('h135f)
	) name9551 (
		\s3_data_i[19]_pad ,
		\s4_data_i[19]_pad ,
		_w9416_,
		_w9500_,
		_w11452_
	);
	LUT4 #(
		.INIT('h135f)
	) name9552 (
		\s11_data_i[19]_pad ,
		\s8_data_i[19]_pad ,
		_w9483_,
		_w9503_,
		_w11453_
	);
	LUT4 #(
		.INIT('h135f)
	) name9553 (
		\s0_data_i[19]_pad ,
		\s9_data_i[19]_pad ,
		_w9291_,
		_w9506_,
		_w11454_
	);
	LUT4 #(
		.INIT('h4000)
	) name9554 (
		_w11451_,
		_w11452_,
		_w11453_,
		_w11454_,
		_w11455_
	);
	LUT2 #(
		.INIT('h8)
	) name9555 (
		_w11450_,
		_w11455_,
		_w11456_
	);
	LUT4 #(
		.INIT('h70ff)
	) name9556 (
		_w2046_,
		_w2097_,
		_w11445_,
		_w11456_,
		_w11457_
	);
	LUT3 #(
		.INIT('h80)
	) name9557 (
		_w2059_,
		_w2097_,
		_w9847_,
		_w11458_
	);
	LUT2 #(
		.INIT('h8)
	) name9558 (
		\s15_data_i[1]_pad ,
		_w2059_,
		_w11459_
	);
	LUT3 #(
		.INIT('h70)
	) name9559 (
		_w2046_,
		_w2097_,
		_w11459_,
		_w11460_
	);
	LUT4 #(
		.INIT('h135f)
	) name9560 (
		\s1_data_i[1]_pad ,
		\s8_data_i[1]_pad ,
		_w9295_,
		_w9503_,
		_w11461_
	);
	LUT4 #(
		.INIT('h153f)
	) name9561 (
		\s4_data_i[1]_pad ,
		\s6_data_i[1]_pad ,
		_w9378_,
		_w9500_,
		_w11462_
	);
	LUT4 #(
		.INIT('h135f)
	) name9562 (
		\s5_data_i[1]_pad ,
		\s9_data_i[1]_pad ,
		_w9387_,
		_w9506_,
		_w11463_
	);
	LUT4 #(
		.INIT('h153f)
	) name9563 (
		\s10_data_i[1]_pad ,
		\s7_data_i[1]_pad ,
		_w9375_,
		_w9480_,
		_w11464_
	);
	LUT4 #(
		.INIT('h8000)
	) name9564 (
		_w11461_,
		_w11462_,
		_w11463_,
		_w11464_,
		_w11465_
	);
	LUT2 #(
		.INIT('h8)
	) name9565 (
		\s11_data_i[1]_pad ,
		_w9483_,
		_w11466_
	);
	LUT4 #(
		.INIT('h153f)
	) name9566 (
		\s13_data_i[1]_pad ,
		\s3_data_i[1]_pad ,
		_w9416_,
		_w9489_,
		_w11467_
	);
	LUT4 #(
		.INIT('h135f)
	) name9567 (
		\s12_data_i[1]_pad ,
		\s14_data_i[1]_pad ,
		_w9486_,
		_w9497_,
		_w11468_
	);
	LUT4 #(
		.INIT('h135f)
	) name9568 (
		\s0_data_i[1]_pad ,
		\s2_data_i[1]_pad ,
		_w9291_,
		_w9494_,
		_w11469_
	);
	LUT4 #(
		.INIT('h4000)
	) name9569 (
		_w11466_,
		_w11467_,
		_w11468_,
		_w11469_,
		_w11470_
	);
	LUT2 #(
		.INIT('h8)
	) name9570 (
		_w11465_,
		_w11470_,
		_w11471_
	);
	LUT3 #(
		.INIT('hef)
	) name9571 (
		_w11458_,
		_w11460_,
		_w11471_,
		_w11472_
	);
	LUT2 #(
		.INIT('h8)
	) name9572 (
		\s15_data_i[20]_pad ,
		_w2059_,
		_w11473_
	);
	LUT4 #(
		.INIT('h135f)
	) name9573 (
		\s12_data_i[20]_pad ,
		\s13_data_i[20]_pad ,
		_w9486_,
		_w9489_,
		_w11474_
	);
	LUT4 #(
		.INIT('h153f)
	) name9574 (
		\s10_data_i[20]_pad ,
		\s1_data_i[20]_pad ,
		_w9295_,
		_w9480_,
		_w11475_
	);
	LUT4 #(
		.INIT('h153f)
	) name9575 (
		\s5_data_i[20]_pad ,
		\s6_data_i[20]_pad ,
		_w9378_,
		_w9387_,
		_w11476_
	);
	LUT4 #(
		.INIT('h153f)
	) name9576 (
		\s2_data_i[20]_pad ,
		\s7_data_i[20]_pad ,
		_w9375_,
		_w9494_,
		_w11477_
	);
	LUT4 #(
		.INIT('h8000)
	) name9577 (
		_w11474_,
		_w11475_,
		_w11476_,
		_w11477_,
		_w11478_
	);
	LUT2 #(
		.INIT('h8)
	) name9578 (
		\s14_data_i[20]_pad ,
		_w9497_,
		_w11479_
	);
	LUT4 #(
		.INIT('h135f)
	) name9579 (
		\s3_data_i[20]_pad ,
		\s4_data_i[20]_pad ,
		_w9416_,
		_w9500_,
		_w11480_
	);
	LUT4 #(
		.INIT('h135f)
	) name9580 (
		\s11_data_i[20]_pad ,
		\s8_data_i[20]_pad ,
		_w9483_,
		_w9503_,
		_w11481_
	);
	LUT4 #(
		.INIT('h135f)
	) name9581 (
		\s0_data_i[20]_pad ,
		\s9_data_i[20]_pad ,
		_w9291_,
		_w9506_,
		_w11482_
	);
	LUT4 #(
		.INIT('h4000)
	) name9582 (
		_w11479_,
		_w11480_,
		_w11481_,
		_w11482_,
		_w11483_
	);
	LUT2 #(
		.INIT('h8)
	) name9583 (
		_w11478_,
		_w11483_,
		_w11484_
	);
	LUT4 #(
		.INIT('h70ff)
	) name9584 (
		_w2046_,
		_w2097_,
		_w11473_,
		_w11484_,
		_w11485_
	);
	LUT2 #(
		.INIT('h8)
	) name9585 (
		\s15_data_i[21]_pad ,
		_w2059_,
		_w11486_
	);
	LUT4 #(
		.INIT('h135f)
	) name9586 (
		\s12_data_i[21]_pad ,
		\s13_data_i[21]_pad ,
		_w9486_,
		_w9489_,
		_w11487_
	);
	LUT4 #(
		.INIT('h153f)
	) name9587 (
		\s10_data_i[21]_pad ,
		\s1_data_i[21]_pad ,
		_w9295_,
		_w9480_,
		_w11488_
	);
	LUT4 #(
		.INIT('h153f)
	) name9588 (
		\s5_data_i[21]_pad ,
		\s6_data_i[21]_pad ,
		_w9378_,
		_w9387_,
		_w11489_
	);
	LUT4 #(
		.INIT('h153f)
	) name9589 (
		\s2_data_i[21]_pad ,
		\s7_data_i[21]_pad ,
		_w9375_,
		_w9494_,
		_w11490_
	);
	LUT4 #(
		.INIT('h8000)
	) name9590 (
		_w11487_,
		_w11488_,
		_w11489_,
		_w11490_,
		_w11491_
	);
	LUT2 #(
		.INIT('h8)
	) name9591 (
		\s14_data_i[21]_pad ,
		_w9497_,
		_w11492_
	);
	LUT4 #(
		.INIT('h135f)
	) name9592 (
		\s3_data_i[21]_pad ,
		\s4_data_i[21]_pad ,
		_w9416_,
		_w9500_,
		_w11493_
	);
	LUT4 #(
		.INIT('h135f)
	) name9593 (
		\s11_data_i[21]_pad ,
		\s8_data_i[21]_pad ,
		_w9483_,
		_w9503_,
		_w11494_
	);
	LUT4 #(
		.INIT('h135f)
	) name9594 (
		\s0_data_i[21]_pad ,
		\s9_data_i[21]_pad ,
		_w9291_,
		_w9506_,
		_w11495_
	);
	LUT4 #(
		.INIT('h4000)
	) name9595 (
		_w11492_,
		_w11493_,
		_w11494_,
		_w11495_,
		_w11496_
	);
	LUT2 #(
		.INIT('h8)
	) name9596 (
		_w11491_,
		_w11496_,
		_w11497_
	);
	LUT4 #(
		.INIT('h70ff)
	) name9597 (
		_w2046_,
		_w2097_,
		_w11486_,
		_w11497_,
		_w11498_
	);
	LUT2 #(
		.INIT('h8)
	) name9598 (
		\s15_data_i[22]_pad ,
		_w2059_,
		_w11499_
	);
	LUT4 #(
		.INIT('h135f)
	) name9599 (
		\s12_data_i[22]_pad ,
		\s13_data_i[22]_pad ,
		_w9486_,
		_w9489_,
		_w11500_
	);
	LUT4 #(
		.INIT('h153f)
	) name9600 (
		\s10_data_i[22]_pad ,
		\s1_data_i[22]_pad ,
		_w9295_,
		_w9480_,
		_w11501_
	);
	LUT4 #(
		.INIT('h153f)
	) name9601 (
		\s5_data_i[22]_pad ,
		\s6_data_i[22]_pad ,
		_w9378_,
		_w9387_,
		_w11502_
	);
	LUT4 #(
		.INIT('h153f)
	) name9602 (
		\s2_data_i[22]_pad ,
		\s7_data_i[22]_pad ,
		_w9375_,
		_w9494_,
		_w11503_
	);
	LUT4 #(
		.INIT('h8000)
	) name9603 (
		_w11500_,
		_w11501_,
		_w11502_,
		_w11503_,
		_w11504_
	);
	LUT2 #(
		.INIT('h8)
	) name9604 (
		\s14_data_i[22]_pad ,
		_w9497_,
		_w11505_
	);
	LUT4 #(
		.INIT('h135f)
	) name9605 (
		\s3_data_i[22]_pad ,
		\s4_data_i[22]_pad ,
		_w9416_,
		_w9500_,
		_w11506_
	);
	LUT4 #(
		.INIT('h135f)
	) name9606 (
		\s11_data_i[22]_pad ,
		\s8_data_i[22]_pad ,
		_w9483_,
		_w9503_,
		_w11507_
	);
	LUT4 #(
		.INIT('h135f)
	) name9607 (
		\s0_data_i[22]_pad ,
		\s9_data_i[22]_pad ,
		_w9291_,
		_w9506_,
		_w11508_
	);
	LUT4 #(
		.INIT('h4000)
	) name9608 (
		_w11505_,
		_w11506_,
		_w11507_,
		_w11508_,
		_w11509_
	);
	LUT2 #(
		.INIT('h8)
	) name9609 (
		_w11504_,
		_w11509_,
		_w11510_
	);
	LUT4 #(
		.INIT('h70ff)
	) name9610 (
		_w2046_,
		_w2097_,
		_w11499_,
		_w11510_,
		_w11511_
	);
	LUT2 #(
		.INIT('h8)
	) name9611 (
		\s15_data_i[23]_pad ,
		_w2059_,
		_w11512_
	);
	LUT4 #(
		.INIT('h135f)
	) name9612 (
		\s12_data_i[23]_pad ,
		\s13_data_i[23]_pad ,
		_w9486_,
		_w9489_,
		_w11513_
	);
	LUT4 #(
		.INIT('h153f)
	) name9613 (
		\s10_data_i[23]_pad ,
		\s1_data_i[23]_pad ,
		_w9295_,
		_w9480_,
		_w11514_
	);
	LUT4 #(
		.INIT('h153f)
	) name9614 (
		\s5_data_i[23]_pad ,
		\s6_data_i[23]_pad ,
		_w9378_,
		_w9387_,
		_w11515_
	);
	LUT4 #(
		.INIT('h153f)
	) name9615 (
		\s2_data_i[23]_pad ,
		\s7_data_i[23]_pad ,
		_w9375_,
		_w9494_,
		_w11516_
	);
	LUT4 #(
		.INIT('h8000)
	) name9616 (
		_w11513_,
		_w11514_,
		_w11515_,
		_w11516_,
		_w11517_
	);
	LUT2 #(
		.INIT('h8)
	) name9617 (
		\s14_data_i[23]_pad ,
		_w9497_,
		_w11518_
	);
	LUT4 #(
		.INIT('h135f)
	) name9618 (
		\s3_data_i[23]_pad ,
		\s4_data_i[23]_pad ,
		_w9416_,
		_w9500_,
		_w11519_
	);
	LUT4 #(
		.INIT('h135f)
	) name9619 (
		\s11_data_i[23]_pad ,
		\s8_data_i[23]_pad ,
		_w9483_,
		_w9503_,
		_w11520_
	);
	LUT4 #(
		.INIT('h135f)
	) name9620 (
		\s0_data_i[23]_pad ,
		\s9_data_i[23]_pad ,
		_w9291_,
		_w9506_,
		_w11521_
	);
	LUT4 #(
		.INIT('h4000)
	) name9621 (
		_w11518_,
		_w11519_,
		_w11520_,
		_w11521_,
		_w11522_
	);
	LUT2 #(
		.INIT('h8)
	) name9622 (
		_w11517_,
		_w11522_,
		_w11523_
	);
	LUT4 #(
		.INIT('h70ff)
	) name9623 (
		_w2046_,
		_w2097_,
		_w11512_,
		_w11523_,
		_w11524_
	);
	LUT2 #(
		.INIT('h8)
	) name9624 (
		\s15_data_i[24]_pad ,
		_w2059_,
		_w11525_
	);
	LUT4 #(
		.INIT('h135f)
	) name9625 (
		\s12_data_i[24]_pad ,
		\s13_data_i[24]_pad ,
		_w9486_,
		_w9489_,
		_w11526_
	);
	LUT4 #(
		.INIT('h153f)
	) name9626 (
		\s10_data_i[24]_pad ,
		\s1_data_i[24]_pad ,
		_w9295_,
		_w9480_,
		_w11527_
	);
	LUT4 #(
		.INIT('h153f)
	) name9627 (
		\s5_data_i[24]_pad ,
		\s6_data_i[24]_pad ,
		_w9378_,
		_w9387_,
		_w11528_
	);
	LUT4 #(
		.INIT('h153f)
	) name9628 (
		\s2_data_i[24]_pad ,
		\s7_data_i[24]_pad ,
		_w9375_,
		_w9494_,
		_w11529_
	);
	LUT4 #(
		.INIT('h8000)
	) name9629 (
		_w11526_,
		_w11527_,
		_w11528_,
		_w11529_,
		_w11530_
	);
	LUT2 #(
		.INIT('h8)
	) name9630 (
		\s14_data_i[24]_pad ,
		_w9497_,
		_w11531_
	);
	LUT4 #(
		.INIT('h135f)
	) name9631 (
		\s3_data_i[24]_pad ,
		\s4_data_i[24]_pad ,
		_w9416_,
		_w9500_,
		_w11532_
	);
	LUT4 #(
		.INIT('h135f)
	) name9632 (
		\s11_data_i[24]_pad ,
		\s8_data_i[24]_pad ,
		_w9483_,
		_w9503_,
		_w11533_
	);
	LUT4 #(
		.INIT('h135f)
	) name9633 (
		\s0_data_i[24]_pad ,
		\s9_data_i[24]_pad ,
		_w9291_,
		_w9506_,
		_w11534_
	);
	LUT4 #(
		.INIT('h4000)
	) name9634 (
		_w11531_,
		_w11532_,
		_w11533_,
		_w11534_,
		_w11535_
	);
	LUT2 #(
		.INIT('h8)
	) name9635 (
		_w11530_,
		_w11535_,
		_w11536_
	);
	LUT4 #(
		.INIT('h70ff)
	) name9636 (
		_w2046_,
		_w2097_,
		_w11525_,
		_w11536_,
		_w11537_
	);
	LUT2 #(
		.INIT('h8)
	) name9637 (
		\s15_data_i[25]_pad ,
		_w2059_,
		_w11538_
	);
	LUT4 #(
		.INIT('h135f)
	) name9638 (
		\s12_data_i[25]_pad ,
		\s13_data_i[25]_pad ,
		_w9486_,
		_w9489_,
		_w11539_
	);
	LUT4 #(
		.INIT('h153f)
	) name9639 (
		\s10_data_i[25]_pad ,
		\s1_data_i[25]_pad ,
		_w9295_,
		_w9480_,
		_w11540_
	);
	LUT4 #(
		.INIT('h153f)
	) name9640 (
		\s5_data_i[25]_pad ,
		\s6_data_i[25]_pad ,
		_w9378_,
		_w9387_,
		_w11541_
	);
	LUT4 #(
		.INIT('h153f)
	) name9641 (
		\s2_data_i[25]_pad ,
		\s7_data_i[25]_pad ,
		_w9375_,
		_w9494_,
		_w11542_
	);
	LUT4 #(
		.INIT('h8000)
	) name9642 (
		_w11539_,
		_w11540_,
		_w11541_,
		_w11542_,
		_w11543_
	);
	LUT2 #(
		.INIT('h8)
	) name9643 (
		\s14_data_i[25]_pad ,
		_w9497_,
		_w11544_
	);
	LUT4 #(
		.INIT('h135f)
	) name9644 (
		\s3_data_i[25]_pad ,
		\s4_data_i[25]_pad ,
		_w9416_,
		_w9500_,
		_w11545_
	);
	LUT4 #(
		.INIT('h135f)
	) name9645 (
		\s11_data_i[25]_pad ,
		\s8_data_i[25]_pad ,
		_w9483_,
		_w9503_,
		_w11546_
	);
	LUT4 #(
		.INIT('h135f)
	) name9646 (
		\s0_data_i[25]_pad ,
		\s9_data_i[25]_pad ,
		_w9291_,
		_w9506_,
		_w11547_
	);
	LUT4 #(
		.INIT('h4000)
	) name9647 (
		_w11544_,
		_w11545_,
		_w11546_,
		_w11547_,
		_w11548_
	);
	LUT2 #(
		.INIT('h8)
	) name9648 (
		_w11543_,
		_w11548_,
		_w11549_
	);
	LUT4 #(
		.INIT('h70ff)
	) name9649 (
		_w2046_,
		_w2097_,
		_w11538_,
		_w11549_,
		_w11550_
	);
	LUT2 #(
		.INIT('h8)
	) name9650 (
		\s15_data_i[26]_pad ,
		_w2059_,
		_w11551_
	);
	LUT4 #(
		.INIT('h135f)
	) name9651 (
		\s12_data_i[26]_pad ,
		\s13_data_i[26]_pad ,
		_w9486_,
		_w9489_,
		_w11552_
	);
	LUT4 #(
		.INIT('h153f)
	) name9652 (
		\s10_data_i[26]_pad ,
		\s1_data_i[26]_pad ,
		_w9295_,
		_w9480_,
		_w11553_
	);
	LUT4 #(
		.INIT('h153f)
	) name9653 (
		\s5_data_i[26]_pad ,
		\s6_data_i[26]_pad ,
		_w9378_,
		_w9387_,
		_w11554_
	);
	LUT4 #(
		.INIT('h153f)
	) name9654 (
		\s2_data_i[26]_pad ,
		\s7_data_i[26]_pad ,
		_w9375_,
		_w9494_,
		_w11555_
	);
	LUT4 #(
		.INIT('h8000)
	) name9655 (
		_w11552_,
		_w11553_,
		_w11554_,
		_w11555_,
		_w11556_
	);
	LUT2 #(
		.INIT('h8)
	) name9656 (
		\s14_data_i[26]_pad ,
		_w9497_,
		_w11557_
	);
	LUT4 #(
		.INIT('h135f)
	) name9657 (
		\s3_data_i[26]_pad ,
		\s4_data_i[26]_pad ,
		_w9416_,
		_w9500_,
		_w11558_
	);
	LUT4 #(
		.INIT('h135f)
	) name9658 (
		\s11_data_i[26]_pad ,
		\s8_data_i[26]_pad ,
		_w9483_,
		_w9503_,
		_w11559_
	);
	LUT4 #(
		.INIT('h135f)
	) name9659 (
		\s0_data_i[26]_pad ,
		\s9_data_i[26]_pad ,
		_w9291_,
		_w9506_,
		_w11560_
	);
	LUT4 #(
		.INIT('h4000)
	) name9660 (
		_w11557_,
		_w11558_,
		_w11559_,
		_w11560_,
		_w11561_
	);
	LUT2 #(
		.INIT('h8)
	) name9661 (
		_w11556_,
		_w11561_,
		_w11562_
	);
	LUT4 #(
		.INIT('h70ff)
	) name9662 (
		_w2046_,
		_w2097_,
		_w11551_,
		_w11562_,
		_w11563_
	);
	LUT2 #(
		.INIT('h8)
	) name9663 (
		\s15_data_i[27]_pad ,
		_w2059_,
		_w11564_
	);
	LUT4 #(
		.INIT('h135f)
	) name9664 (
		\s12_data_i[27]_pad ,
		\s13_data_i[27]_pad ,
		_w9486_,
		_w9489_,
		_w11565_
	);
	LUT4 #(
		.INIT('h153f)
	) name9665 (
		\s10_data_i[27]_pad ,
		\s1_data_i[27]_pad ,
		_w9295_,
		_w9480_,
		_w11566_
	);
	LUT4 #(
		.INIT('h153f)
	) name9666 (
		\s5_data_i[27]_pad ,
		\s6_data_i[27]_pad ,
		_w9378_,
		_w9387_,
		_w11567_
	);
	LUT4 #(
		.INIT('h153f)
	) name9667 (
		\s2_data_i[27]_pad ,
		\s7_data_i[27]_pad ,
		_w9375_,
		_w9494_,
		_w11568_
	);
	LUT4 #(
		.INIT('h8000)
	) name9668 (
		_w11565_,
		_w11566_,
		_w11567_,
		_w11568_,
		_w11569_
	);
	LUT2 #(
		.INIT('h8)
	) name9669 (
		\s14_data_i[27]_pad ,
		_w9497_,
		_w11570_
	);
	LUT4 #(
		.INIT('h135f)
	) name9670 (
		\s3_data_i[27]_pad ,
		\s4_data_i[27]_pad ,
		_w9416_,
		_w9500_,
		_w11571_
	);
	LUT4 #(
		.INIT('h135f)
	) name9671 (
		\s11_data_i[27]_pad ,
		\s8_data_i[27]_pad ,
		_w9483_,
		_w9503_,
		_w11572_
	);
	LUT4 #(
		.INIT('h135f)
	) name9672 (
		\s0_data_i[27]_pad ,
		\s9_data_i[27]_pad ,
		_w9291_,
		_w9506_,
		_w11573_
	);
	LUT4 #(
		.INIT('h4000)
	) name9673 (
		_w11570_,
		_w11571_,
		_w11572_,
		_w11573_,
		_w11574_
	);
	LUT2 #(
		.INIT('h8)
	) name9674 (
		_w11569_,
		_w11574_,
		_w11575_
	);
	LUT4 #(
		.INIT('h70ff)
	) name9675 (
		_w2046_,
		_w2097_,
		_w11564_,
		_w11575_,
		_w11576_
	);
	LUT2 #(
		.INIT('h8)
	) name9676 (
		\s15_data_i[28]_pad ,
		_w2059_,
		_w11577_
	);
	LUT4 #(
		.INIT('h135f)
	) name9677 (
		\s12_data_i[28]_pad ,
		\s13_data_i[28]_pad ,
		_w9486_,
		_w9489_,
		_w11578_
	);
	LUT4 #(
		.INIT('h153f)
	) name9678 (
		\s10_data_i[28]_pad ,
		\s1_data_i[28]_pad ,
		_w9295_,
		_w9480_,
		_w11579_
	);
	LUT4 #(
		.INIT('h153f)
	) name9679 (
		\s5_data_i[28]_pad ,
		\s6_data_i[28]_pad ,
		_w9378_,
		_w9387_,
		_w11580_
	);
	LUT4 #(
		.INIT('h153f)
	) name9680 (
		\s2_data_i[28]_pad ,
		\s7_data_i[28]_pad ,
		_w9375_,
		_w9494_,
		_w11581_
	);
	LUT4 #(
		.INIT('h8000)
	) name9681 (
		_w11578_,
		_w11579_,
		_w11580_,
		_w11581_,
		_w11582_
	);
	LUT2 #(
		.INIT('h8)
	) name9682 (
		\s14_data_i[28]_pad ,
		_w9497_,
		_w11583_
	);
	LUT4 #(
		.INIT('h135f)
	) name9683 (
		\s3_data_i[28]_pad ,
		\s4_data_i[28]_pad ,
		_w9416_,
		_w9500_,
		_w11584_
	);
	LUT4 #(
		.INIT('h135f)
	) name9684 (
		\s11_data_i[28]_pad ,
		\s8_data_i[28]_pad ,
		_w9483_,
		_w9503_,
		_w11585_
	);
	LUT4 #(
		.INIT('h135f)
	) name9685 (
		\s0_data_i[28]_pad ,
		\s9_data_i[28]_pad ,
		_w9291_,
		_w9506_,
		_w11586_
	);
	LUT4 #(
		.INIT('h4000)
	) name9686 (
		_w11583_,
		_w11584_,
		_w11585_,
		_w11586_,
		_w11587_
	);
	LUT2 #(
		.INIT('h8)
	) name9687 (
		_w11582_,
		_w11587_,
		_w11588_
	);
	LUT4 #(
		.INIT('h70ff)
	) name9688 (
		_w2046_,
		_w2097_,
		_w11577_,
		_w11588_,
		_w11589_
	);
	LUT2 #(
		.INIT('h8)
	) name9689 (
		\s15_data_i[29]_pad ,
		_w2059_,
		_w11590_
	);
	LUT4 #(
		.INIT('h135f)
	) name9690 (
		\s12_data_i[29]_pad ,
		\s13_data_i[29]_pad ,
		_w9486_,
		_w9489_,
		_w11591_
	);
	LUT4 #(
		.INIT('h153f)
	) name9691 (
		\s10_data_i[29]_pad ,
		\s1_data_i[29]_pad ,
		_w9295_,
		_w9480_,
		_w11592_
	);
	LUT4 #(
		.INIT('h153f)
	) name9692 (
		\s5_data_i[29]_pad ,
		\s6_data_i[29]_pad ,
		_w9378_,
		_w9387_,
		_w11593_
	);
	LUT4 #(
		.INIT('h153f)
	) name9693 (
		\s2_data_i[29]_pad ,
		\s7_data_i[29]_pad ,
		_w9375_,
		_w9494_,
		_w11594_
	);
	LUT4 #(
		.INIT('h8000)
	) name9694 (
		_w11591_,
		_w11592_,
		_w11593_,
		_w11594_,
		_w11595_
	);
	LUT2 #(
		.INIT('h8)
	) name9695 (
		\s14_data_i[29]_pad ,
		_w9497_,
		_w11596_
	);
	LUT4 #(
		.INIT('h135f)
	) name9696 (
		\s3_data_i[29]_pad ,
		\s4_data_i[29]_pad ,
		_w9416_,
		_w9500_,
		_w11597_
	);
	LUT4 #(
		.INIT('h135f)
	) name9697 (
		\s11_data_i[29]_pad ,
		\s8_data_i[29]_pad ,
		_w9483_,
		_w9503_,
		_w11598_
	);
	LUT4 #(
		.INIT('h135f)
	) name9698 (
		\s0_data_i[29]_pad ,
		\s9_data_i[29]_pad ,
		_w9291_,
		_w9506_,
		_w11599_
	);
	LUT4 #(
		.INIT('h4000)
	) name9699 (
		_w11596_,
		_w11597_,
		_w11598_,
		_w11599_,
		_w11600_
	);
	LUT2 #(
		.INIT('h8)
	) name9700 (
		_w11595_,
		_w11600_,
		_w11601_
	);
	LUT4 #(
		.INIT('h70ff)
	) name9701 (
		_w2046_,
		_w2097_,
		_w11590_,
		_w11601_,
		_w11602_
	);
	LUT3 #(
		.INIT('h80)
	) name9702 (
		_w2059_,
		_w2097_,
		_w9993_,
		_w11603_
	);
	LUT2 #(
		.INIT('h8)
	) name9703 (
		\s15_data_i[2]_pad ,
		_w2059_,
		_w11604_
	);
	LUT3 #(
		.INIT('h70)
	) name9704 (
		_w2046_,
		_w2097_,
		_w11604_,
		_w11605_
	);
	LUT4 #(
		.INIT('h135f)
	) name9705 (
		\s1_data_i[2]_pad ,
		\s8_data_i[2]_pad ,
		_w9295_,
		_w9503_,
		_w11606_
	);
	LUT4 #(
		.INIT('h153f)
	) name9706 (
		\s4_data_i[2]_pad ,
		\s6_data_i[2]_pad ,
		_w9378_,
		_w9500_,
		_w11607_
	);
	LUT4 #(
		.INIT('h135f)
	) name9707 (
		\s5_data_i[2]_pad ,
		\s9_data_i[2]_pad ,
		_w9387_,
		_w9506_,
		_w11608_
	);
	LUT4 #(
		.INIT('h153f)
	) name9708 (
		\s10_data_i[2]_pad ,
		\s7_data_i[2]_pad ,
		_w9375_,
		_w9480_,
		_w11609_
	);
	LUT4 #(
		.INIT('h8000)
	) name9709 (
		_w11606_,
		_w11607_,
		_w11608_,
		_w11609_,
		_w11610_
	);
	LUT2 #(
		.INIT('h8)
	) name9710 (
		\s11_data_i[2]_pad ,
		_w9483_,
		_w11611_
	);
	LUT4 #(
		.INIT('h153f)
	) name9711 (
		\s13_data_i[2]_pad ,
		\s3_data_i[2]_pad ,
		_w9416_,
		_w9489_,
		_w11612_
	);
	LUT4 #(
		.INIT('h135f)
	) name9712 (
		\s12_data_i[2]_pad ,
		\s14_data_i[2]_pad ,
		_w9486_,
		_w9497_,
		_w11613_
	);
	LUT4 #(
		.INIT('h135f)
	) name9713 (
		\s0_data_i[2]_pad ,
		\s2_data_i[2]_pad ,
		_w9291_,
		_w9494_,
		_w11614_
	);
	LUT4 #(
		.INIT('h4000)
	) name9714 (
		_w11611_,
		_w11612_,
		_w11613_,
		_w11614_,
		_w11615_
	);
	LUT2 #(
		.INIT('h8)
	) name9715 (
		_w11610_,
		_w11615_,
		_w11616_
	);
	LUT3 #(
		.INIT('hef)
	) name9716 (
		_w11603_,
		_w11605_,
		_w11616_,
		_w11617_
	);
	LUT2 #(
		.INIT('h8)
	) name9717 (
		\s15_data_i[30]_pad ,
		_w2059_,
		_w11618_
	);
	LUT4 #(
		.INIT('h135f)
	) name9718 (
		\s12_data_i[30]_pad ,
		\s13_data_i[30]_pad ,
		_w9486_,
		_w9489_,
		_w11619_
	);
	LUT4 #(
		.INIT('h153f)
	) name9719 (
		\s10_data_i[30]_pad ,
		\s1_data_i[30]_pad ,
		_w9295_,
		_w9480_,
		_w11620_
	);
	LUT4 #(
		.INIT('h153f)
	) name9720 (
		\s5_data_i[30]_pad ,
		\s6_data_i[30]_pad ,
		_w9378_,
		_w9387_,
		_w11621_
	);
	LUT4 #(
		.INIT('h153f)
	) name9721 (
		\s2_data_i[30]_pad ,
		\s7_data_i[30]_pad ,
		_w9375_,
		_w9494_,
		_w11622_
	);
	LUT4 #(
		.INIT('h8000)
	) name9722 (
		_w11619_,
		_w11620_,
		_w11621_,
		_w11622_,
		_w11623_
	);
	LUT2 #(
		.INIT('h8)
	) name9723 (
		\s14_data_i[30]_pad ,
		_w9497_,
		_w11624_
	);
	LUT4 #(
		.INIT('h135f)
	) name9724 (
		\s3_data_i[30]_pad ,
		\s4_data_i[30]_pad ,
		_w9416_,
		_w9500_,
		_w11625_
	);
	LUT4 #(
		.INIT('h135f)
	) name9725 (
		\s11_data_i[30]_pad ,
		\s8_data_i[30]_pad ,
		_w9483_,
		_w9503_,
		_w11626_
	);
	LUT4 #(
		.INIT('h135f)
	) name9726 (
		\s0_data_i[30]_pad ,
		\s9_data_i[30]_pad ,
		_w9291_,
		_w9506_,
		_w11627_
	);
	LUT4 #(
		.INIT('h4000)
	) name9727 (
		_w11624_,
		_w11625_,
		_w11626_,
		_w11627_,
		_w11628_
	);
	LUT2 #(
		.INIT('h8)
	) name9728 (
		_w11623_,
		_w11628_,
		_w11629_
	);
	LUT4 #(
		.INIT('h70ff)
	) name9729 (
		_w2046_,
		_w2097_,
		_w11618_,
		_w11629_,
		_w11630_
	);
	LUT2 #(
		.INIT('h8)
	) name9730 (
		\s15_data_i[31]_pad ,
		_w2059_,
		_w11631_
	);
	LUT4 #(
		.INIT('h135f)
	) name9731 (
		\s12_data_i[31]_pad ,
		\s13_data_i[31]_pad ,
		_w9486_,
		_w9489_,
		_w11632_
	);
	LUT4 #(
		.INIT('h153f)
	) name9732 (
		\s10_data_i[31]_pad ,
		\s1_data_i[31]_pad ,
		_w9295_,
		_w9480_,
		_w11633_
	);
	LUT4 #(
		.INIT('h153f)
	) name9733 (
		\s5_data_i[31]_pad ,
		\s6_data_i[31]_pad ,
		_w9378_,
		_w9387_,
		_w11634_
	);
	LUT4 #(
		.INIT('h153f)
	) name9734 (
		\s2_data_i[31]_pad ,
		\s7_data_i[31]_pad ,
		_w9375_,
		_w9494_,
		_w11635_
	);
	LUT4 #(
		.INIT('h8000)
	) name9735 (
		_w11632_,
		_w11633_,
		_w11634_,
		_w11635_,
		_w11636_
	);
	LUT2 #(
		.INIT('h8)
	) name9736 (
		\s14_data_i[31]_pad ,
		_w9497_,
		_w11637_
	);
	LUT4 #(
		.INIT('h135f)
	) name9737 (
		\s3_data_i[31]_pad ,
		\s4_data_i[31]_pad ,
		_w9416_,
		_w9500_,
		_w11638_
	);
	LUT4 #(
		.INIT('h135f)
	) name9738 (
		\s11_data_i[31]_pad ,
		\s8_data_i[31]_pad ,
		_w9483_,
		_w9503_,
		_w11639_
	);
	LUT4 #(
		.INIT('h135f)
	) name9739 (
		\s0_data_i[31]_pad ,
		\s9_data_i[31]_pad ,
		_w9291_,
		_w9506_,
		_w11640_
	);
	LUT4 #(
		.INIT('h4000)
	) name9740 (
		_w11637_,
		_w11638_,
		_w11639_,
		_w11640_,
		_w11641_
	);
	LUT2 #(
		.INIT('h8)
	) name9741 (
		_w11636_,
		_w11641_,
		_w11642_
	);
	LUT4 #(
		.INIT('h70ff)
	) name9742 (
		_w2046_,
		_w2097_,
		_w11631_,
		_w11642_,
		_w11643_
	);
	LUT3 #(
		.INIT('h80)
	) name9743 (
		_w2059_,
		_w2097_,
		_w10035_,
		_w11644_
	);
	LUT2 #(
		.INIT('h8)
	) name9744 (
		\s15_data_i[3]_pad ,
		_w2059_,
		_w11645_
	);
	LUT3 #(
		.INIT('h70)
	) name9745 (
		_w2046_,
		_w2097_,
		_w11645_,
		_w11646_
	);
	LUT4 #(
		.INIT('h135f)
	) name9746 (
		\s13_data_i[3]_pad ,
		\s8_data_i[3]_pad ,
		_w9489_,
		_w9503_,
		_w11647_
	);
	LUT4 #(
		.INIT('h153f)
	) name9747 (
		\s10_data_i[3]_pad ,
		\s1_data_i[3]_pad ,
		_w9295_,
		_w9480_,
		_w11648_
	);
	LUT4 #(
		.INIT('h153f)
	) name9748 (
		\s5_data_i[3]_pad ,
		\s6_data_i[3]_pad ,
		_w9378_,
		_w9387_,
		_w11649_
	);
	LUT4 #(
		.INIT('h153f)
	) name9749 (
		\s2_data_i[3]_pad ,
		\s7_data_i[3]_pad ,
		_w9375_,
		_w9494_,
		_w11650_
	);
	LUT4 #(
		.INIT('h8000)
	) name9750 (
		_w11647_,
		_w11648_,
		_w11649_,
		_w11650_,
		_w11651_
	);
	LUT2 #(
		.INIT('h8)
	) name9751 (
		\s11_data_i[3]_pad ,
		_w9483_,
		_w11652_
	);
	LUT4 #(
		.INIT('h135f)
	) name9752 (
		\s3_data_i[3]_pad ,
		\s4_data_i[3]_pad ,
		_w9416_,
		_w9500_,
		_w11653_
	);
	LUT4 #(
		.INIT('h135f)
	) name9753 (
		\s12_data_i[3]_pad ,
		\s14_data_i[3]_pad ,
		_w9486_,
		_w9497_,
		_w11654_
	);
	LUT4 #(
		.INIT('h135f)
	) name9754 (
		\s0_data_i[3]_pad ,
		\s9_data_i[3]_pad ,
		_w9291_,
		_w9506_,
		_w11655_
	);
	LUT4 #(
		.INIT('h4000)
	) name9755 (
		_w11652_,
		_w11653_,
		_w11654_,
		_w11655_,
		_w11656_
	);
	LUT2 #(
		.INIT('h8)
	) name9756 (
		_w11651_,
		_w11656_,
		_w11657_
	);
	LUT3 #(
		.INIT('hef)
	) name9757 (
		_w11644_,
		_w11646_,
		_w11657_,
		_w11658_
	);
	LUT3 #(
		.INIT('h80)
	) name9758 (
		_w2059_,
		_w2097_,
		_w10051_,
		_w11659_
	);
	LUT2 #(
		.INIT('h8)
	) name9759 (
		\s15_data_i[4]_pad ,
		_w2059_,
		_w11660_
	);
	LUT3 #(
		.INIT('h70)
	) name9760 (
		_w2046_,
		_w2097_,
		_w11660_,
		_w11661_
	);
	LUT4 #(
		.INIT('h135f)
	) name9761 (
		\s4_data_i[4]_pad ,
		\s8_data_i[4]_pad ,
		_w9500_,
		_w9503_,
		_w11662_
	);
	LUT4 #(
		.INIT('h135f)
	) name9762 (
		\s1_data_i[4]_pad ,
		\s7_data_i[4]_pad ,
		_w9295_,
		_w9375_,
		_w11663_
	);
	LUT4 #(
		.INIT('h153f)
	) name9763 (
		\s5_data_i[4]_pad ,
		\s6_data_i[4]_pad ,
		_w9378_,
		_w9387_,
		_w11664_
	);
	LUT4 #(
		.INIT('h135f)
	) name9764 (
		\s13_data_i[4]_pad ,
		\s2_data_i[4]_pad ,
		_w9489_,
		_w9494_,
		_w11665_
	);
	LUT4 #(
		.INIT('h8000)
	) name9765 (
		_w11662_,
		_w11663_,
		_w11664_,
		_w11665_,
		_w11666_
	);
	LUT2 #(
		.INIT('h8)
	) name9766 (
		\s11_data_i[4]_pad ,
		_w9483_,
		_w11667_
	);
	LUT4 #(
		.INIT('h153f)
	) name9767 (
		\s10_data_i[4]_pad ,
		\s3_data_i[4]_pad ,
		_w9416_,
		_w9480_,
		_w11668_
	);
	LUT4 #(
		.INIT('h135f)
	) name9768 (
		\s12_data_i[4]_pad ,
		\s14_data_i[4]_pad ,
		_w9486_,
		_w9497_,
		_w11669_
	);
	LUT4 #(
		.INIT('h135f)
	) name9769 (
		\s0_data_i[4]_pad ,
		\s9_data_i[4]_pad ,
		_w9291_,
		_w9506_,
		_w11670_
	);
	LUT4 #(
		.INIT('h4000)
	) name9770 (
		_w11667_,
		_w11668_,
		_w11669_,
		_w11670_,
		_w11671_
	);
	LUT2 #(
		.INIT('h8)
	) name9771 (
		_w11666_,
		_w11671_,
		_w11672_
	);
	LUT3 #(
		.INIT('hef)
	) name9772 (
		_w11659_,
		_w11661_,
		_w11672_,
		_w11673_
	);
	LUT3 #(
		.INIT('h80)
	) name9773 (
		_w2059_,
		_w2097_,
		_w10067_,
		_w11674_
	);
	LUT2 #(
		.INIT('h8)
	) name9774 (
		\s15_data_i[5]_pad ,
		_w2059_,
		_w11675_
	);
	LUT3 #(
		.INIT('h70)
	) name9775 (
		_w2046_,
		_w2097_,
		_w11675_,
		_w11676_
	);
	LUT4 #(
		.INIT('h135f)
	) name9776 (
		\s13_data_i[5]_pad ,
		\s8_data_i[5]_pad ,
		_w9489_,
		_w9503_,
		_w11677_
	);
	LUT4 #(
		.INIT('h153f)
	) name9777 (
		\s10_data_i[5]_pad ,
		\s1_data_i[5]_pad ,
		_w9295_,
		_w9480_,
		_w11678_
	);
	LUT4 #(
		.INIT('h153f)
	) name9778 (
		\s5_data_i[5]_pad ,
		\s6_data_i[5]_pad ,
		_w9378_,
		_w9387_,
		_w11679_
	);
	LUT4 #(
		.INIT('h153f)
	) name9779 (
		\s2_data_i[5]_pad ,
		\s7_data_i[5]_pad ,
		_w9375_,
		_w9494_,
		_w11680_
	);
	LUT4 #(
		.INIT('h8000)
	) name9780 (
		_w11677_,
		_w11678_,
		_w11679_,
		_w11680_,
		_w11681_
	);
	LUT2 #(
		.INIT('h8)
	) name9781 (
		\s11_data_i[5]_pad ,
		_w9483_,
		_w11682_
	);
	LUT4 #(
		.INIT('h135f)
	) name9782 (
		\s3_data_i[5]_pad ,
		\s4_data_i[5]_pad ,
		_w9416_,
		_w9500_,
		_w11683_
	);
	LUT4 #(
		.INIT('h135f)
	) name9783 (
		\s12_data_i[5]_pad ,
		\s14_data_i[5]_pad ,
		_w9486_,
		_w9497_,
		_w11684_
	);
	LUT4 #(
		.INIT('h135f)
	) name9784 (
		\s0_data_i[5]_pad ,
		\s9_data_i[5]_pad ,
		_w9291_,
		_w9506_,
		_w11685_
	);
	LUT4 #(
		.INIT('h4000)
	) name9785 (
		_w11682_,
		_w11683_,
		_w11684_,
		_w11685_,
		_w11686_
	);
	LUT2 #(
		.INIT('h8)
	) name9786 (
		_w11681_,
		_w11686_,
		_w11687_
	);
	LUT3 #(
		.INIT('hef)
	) name9787 (
		_w11674_,
		_w11676_,
		_w11687_,
		_w11688_
	);
	LUT3 #(
		.INIT('h80)
	) name9788 (
		_w2059_,
		_w2097_,
		_w10083_,
		_w11689_
	);
	LUT2 #(
		.INIT('h8)
	) name9789 (
		\s15_data_i[6]_pad ,
		_w2059_,
		_w11690_
	);
	LUT3 #(
		.INIT('h70)
	) name9790 (
		_w2046_,
		_w2097_,
		_w11690_,
		_w11691_
	);
	LUT4 #(
		.INIT('h135f)
	) name9791 (
		\s13_data_i[6]_pad ,
		\s8_data_i[6]_pad ,
		_w9489_,
		_w9503_,
		_w11692_
	);
	LUT4 #(
		.INIT('h153f)
	) name9792 (
		\s10_data_i[6]_pad ,
		\s1_data_i[6]_pad ,
		_w9295_,
		_w9480_,
		_w11693_
	);
	LUT4 #(
		.INIT('h153f)
	) name9793 (
		\s5_data_i[6]_pad ,
		\s6_data_i[6]_pad ,
		_w9378_,
		_w9387_,
		_w11694_
	);
	LUT4 #(
		.INIT('h153f)
	) name9794 (
		\s2_data_i[6]_pad ,
		\s7_data_i[6]_pad ,
		_w9375_,
		_w9494_,
		_w11695_
	);
	LUT4 #(
		.INIT('h8000)
	) name9795 (
		_w11692_,
		_w11693_,
		_w11694_,
		_w11695_,
		_w11696_
	);
	LUT2 #(
		.INIT('h8)
	) name9796 (
		\s11_data_i[6]_pad ,
		_w9483_,
		_w11697_
	);
	LUT4 #(
		.INIT('h135f)
	) name9797 (
		\s3_data_i[6]_pad ,
		\s4_data_i[6]_pad ,
		_w9416_,
		_w9500_,
		_w11698_
	);
	LUT4 #(
		.INIT('h135f)
	) name9798 (
		\s12_data_i[6]_pad ,
		\s14_data_i[6]_pad ,
		_w9486_,
		_w9497_,
		_w11699_
	);
	LUT4 #(
		.INIT('h135f)
	) name9799 (
		\s0_data_i[6]_pad ,
		\s9_data_i[6]_pad ,
		_w9291_,
		_w9506_,
		_w11700_
	);
	LUT4 #(
		.INIT('h4000)
	) name9800 (
		_w11697_,
		_w11698_,
		_w11699_,
		_w11700_,
		_w11701_
	);
	LUT2 #(
		.INIT('h8)
	) name9801 (
		_w11696_,
		_w11701_,
		_w11702_
	);
	LUT3 #(
		.INIT('hef)
	) name9802 (
		_w11689_,
		_w11691_,
		_w11702_,
		_w11703_
	);
	LUT3 #(
		.INIT('h80)
	) name9803 (
		_w2059_,
		_w2097_,
		_w10099_,
		_w11704_
	);
	LUT2 #(
		.INIT('h8)
	) name9804 (
		\s15_data_i[7]_pad ,
		_w2059_,
		_w11705_
	);
	LUT3 #(
		.INIT('h70)
	) name9805 (
		_w2046_,
		_w2097_,
		_w11705_,
		_w11706_
	);
	LUT4 #(
		.INIT('h135f)
	) name9806 (
		\s13_data_i[7]_pad ,
		\s2_data_i[7]_pad ,
		_w9489_,
		_w9494_,
		_w11707_
	);
	LUT4 #(
		.INIT('h153f)
	) name9807 (
		\s11_data_i[7]_pad ,
		\s6_data_i[7]_pad ,
		_w9378_,
		_w9483_,
		_w11708_
	);
	LUT4 #(
		.INIT('h135f)
	) name9808 (
		\s3_data_i[7]_pad ,
		\s4_data_i[7]_pad ,
		_w9416_,
		_w9500_,
		_w11709_
	);
	LUT4 #(
		.INIT('h153f)
	) name9809 (
		\s12_data_i[7]_pad ,
		\s7_data_i[7]_pad ,
		_w9375_,
		_w9486_,
		_w11710_
	);
	LUT4 #(
		.INIT('h8000)
	) name9810 (
		_w11707_,
		_w11708_,
		_w11709_,
		_w11710_,
		_w11711_
	);
	LUT2 #(
		.INIT('h8)
	) name9811 (
		\s1_data_i[7]_pad ,
		_w9295_,
		_w11712_
	);
	LUT4 #(
		.INIT('h135f)
	) name9812 (
		\s0_data_i[7]_pad ,
		\s8_data_i[7]_pad ,
		_w9291_,
		_w9503_,
		_w11713_
	);
	LUT4 #(
		.INIT('h135f)
	) name9813 (
		\s10_data_i[7]_pad ,
		\s9_data_i[7]_pad ,
		_w9480_,
		_w9506_,
		_w11714_
	);
	LUT4 #(
		.INIT('h153f)
	) name9814 (
		\s14_data_i[7]_pad ,
		\s5_data_i[7]_pad ,
		_w9387_,
		_w9497_,
		_w11715_
	);
	LUT4 #(
		.INIT('h4000)
	) name9815 (
		_w11712_,
		_w11713_,
		_w11714_,
		_w11715_,
		_w11716_
	);
	LUT2 #(
		.INIT('h8)
	) name9816 (
		_w11711_,
		_w11716_,
		_w11717_
	);
	LUT3 #(
		.INIT('hef)
	) name9817 (
		_w11704_,
		_w11706_,
		_w11717_,
		_w11718_
	);
	LUT3 #(
		.INIT('h80)
	) name9818 (
		_w2059_,
		_w2097_,
		_w10115_,
		_w11719_
	);
	LUT2 #(
		.INIT('h8)
	) name9819 (
		\s15_data_i[8]_pad ,
		_w2059_,
		_w11720_
	);
	LUT3 #(
		.INIT('h70)
	) name9820 (
		_w2046_,
		_w2097_,
		_w11720_,
		_w11721_
	);
	LUT4 #(
		.INIT('h135f)
	) name9821 (
		\s13_data_i[8]_pad ,
		\s8_data_i[8]_pad ,
		_w9489_,
		_w9503_,
		_w11722_
	);
	LUT4 #(
		.INIT('h153f)
	) name9822 (
		\s10_data_i[8]_pad ,
		\s1_data_i[8]_pad ,
		_w9295_,
		_w9480_,
		_w11723_
	);
	LUT4 #(
		.INIT('h153f)
	) name9823 (
		\s5_data_i[8]_pad ,
		\s6_data_i[8]_pad ,
		_w9378_,
		_w9387_,
		_w11724_
	);
	LUT4 #(
		.INIT('h153f)
	) name9824 (
		\s2_data_i[8]_pad ,
		\s7_data_i[8]_pad ,
		_w9375_,
		_w9494_,
		_w11725_
	);
	LUT4 #(
		.INIT('h8000)
	) name9825 (
		_w11722_,
		_w11723_,
		_w11724_,
		_w11725_,
		_w11726_
	);
	LUT2 #(
		.INIT('h8)
	) name9826 (
		\s11_data_i[8]_pad ,
		_w9483_,
		_w11727_
	);
	LUT4 #(
		.INIT('h135f)
	) name9827 (
		\s3_data_i[8]_pad ,
		\s4_data_i[8]_pad ,
		_w9416_,
		_w9500_,
		_w11728_
	);
	LUT4 #(
		.INIT('h135f)
	) name9828 (
		\s12_data_i[8]_pad ,
		\s14_data_i[8]_pad ,
		_w9486_,
		_w9497_,
		_w11729_
	);
	LUT4 #(
		.INIT('h135f)
	) name9829 (
		\s0_data_i[8]_pad ,
		\s9_data_i[8]_pad ,
		_w9291_,
		_w9506_,
		_w11730_
	);
	LUT4 #(
		.INIT('h4000)
	) name9830 (
		_w11727_,
		_w11728_,
		_w11729_,
		_w11730_,
		_w11731_
	);
	LUT2 #(
		.INIT('h8)
	) name9831 (
		_w11726_,
		_w11731_,
		_w11732_
	);
	LUT3 #(
		.INIT('hef)
	) name9832 (
		_w11719_,
		_w11721_,
		_w11732_,
		_w11733_
	);
	LUT3 #(
		.INIT('h80)
	) name9833 (
		_w2059_,
		_w2097_,
		_w10131_,
		_w11734_
	);
	LUT2 #(
		.INIT('h8)
	) name9834 (
		\s15_data_i[9]_pad ,
		_w2059_,
		_w11735_
	);
	LUT3 #(
		.INIT('h70)
	) name9835 (
		_w2046_,
		_w2097_,
		_w11735_,
		_w11736_
	);
	LUT4 #(
		.INIT('h135f)
	) name9836 (
		\s13_data_i[9]_pad ,
		\s2_data_i[9]_pad ,
		_w9489_,
		_w9494_,
		_w11737_
	);
	LUT4 #(
		.INIT('h153f)
	) name9837 (
		\s11_data_i[9]_pad ,
		\s6_data_i[9]_pad ,
		_w9378_,
		_w9483_,
		_w11738_
	);
	LUT4 #(
		.INIT('h135f)
	) name9838 (
		\s3_data_i[9]_pad ,
		\s4_data_i[9]_pad ,
		_w9416_,
		_w9500_,
		_w11739_
	);
	LUT4 #(
		.INIT('h153f)
	) name9839 (
		\s12_data_i[9]_pad ,
		\s7_data_i[9]_pad ,
		_w9375_,
		_w9486_,
		_w11740_
	);
	LUT4 #(
		.INIT('h8000)
	) name9840 (
		_w11737_,
		_w11738_,
		_w11739_,
		_w11740_,
		_w11741_
	);
	LUT2 #(
		.INIT('h8)
	) name9841 (
		\s1_data_i[9]_pad ,
		_w9295_,
		_w11742_
	);
	LUT4 #(
		.INIT('h135f)
	) name9842 (
		\s0_data_i[9]_pad ,
		\s8_data_i[9]_pad ,
		_w9291_,
		_w9503_,
		_w11743_
	);
	LUT4 #(
		.INIT('h135f)
	) name9843 (
		\s10_data_i[9]_pad ,
		\s9_data_i[9]_pad ,
		_w9480_,
		_w9506_,
		_w11744_
	);
	LUT4 #(
		.INIT('h153f)
	) name9844 (
		\s14_data_i[9]_pad ,
		\s5_data_i[9]_pad ,
		_w9387_,
		_w9497_,
		_w11745_
	);
	LUT4 #(
		.INIT('h4000)
	) name9845 (
		_w11742_,
		_w11743_,
		_w11744_,
		_w11745_,
		_w11746_
	);
	LUT2 #(
		.INIT('h8)
	) name9846 (
		_w11741_,
		_w11746_,
		_w11747_
	);
	LUT3 #(
		.INIT('hef)
	) name9847 (
		_w11734_,
		_w11736_,
		_w11747_,
		_w11748_
	);
	LUT3 #(
		.INIT('h80)
	) name9848 (
		\s15_err_i_pad ,
		_w1918_,
		_w11271_,
		_w11749_
	);
	LUT4 #(
		.INIT('h2a00)
	) name9849 (
		\s14_err_i_pad ,
		_w9137_,
		_w9138_,
		_w9497_,
		_w11750_
	);
	LUT4 #(
		.INIT('h2a00)
	) name9850 (
		\s3_err_i_pad ,
		_w9205_,
		_w9206_,
		_w9416_,
		_w11751_
	);
	LUT4 #(
		.INIT('h135f)
	) name9851 (
		_w9144_,
		_w9212_,
		_w11750_,
		_w11751_,
		_w11752_
	);
	LUT4 #(
		.INIT('h2a00)
	) name9852 (
		\s13_err_i_pad ,
		_w9069_,
		_w9070_,
		_w9489_,
		_w11753_
	);
	LUT4 #(
		.INIT('h2a00)
	) name9853 (
		\s6_err_i_pad ,
		_w8743_,
		_w8744_,
		_w9378_,
		_w11754_
	);
	LUT4 #(
		.INIT('h153f)
	) name9854 (
		_w8750_,
		_w9082_,
		_w11753_,
		_w11754_,
		_w11755_
	);
	LUT4 #(
		.INIT('h2a00)
	) name9855 (
		\s0_err_i_pad ,
		_w8989_,
		_w8990_,
		_w9291_,
		_w11756_
	);
	LUT4 #(
		.INIT('h2a00)
	) name9856 (
		\s10_err_i_pad ,
		_w8910_,
		_w8911_,
		_w9480_,
		_w11757_
	);
	LUT4 #(
		.INIT('h153f)
	) name9857 (
		_w8909_,
		_w9002_,
		_w11756_,
		_w11757_,
		_w11758_
	);
	LUT4 #(
		.INIT('h2a00)
	) name9858 (
		\s9_err_i_pad ,
		_w8865_,
		_w8866_,
		_w9506_,
		_w11759_
	);
	LUT4 #(
		.INIT('h2a00)
	) name9859 (
		\s7_err_i_pad ,
		_w8782_,
		_w8783_,
		_w9375_,
		_w11760_
	);
	LUT4 #(
		.INIT('h153f)
	) name9860 (
		_w8795_,
		_w8864_,
		_w11759_,
		_w11760_,
		_w11761_
	);
	LUT4 #(
		.INIT('h8000)
	) name9861 (
		_w11752_,
		_w11755_,
		_w11758_,
		_w11761_,
		_w11762_
	);
	LUT4 #(
		.INIT('h2a00)
	) name9862 (
		\s12_err_i_pad ,
		_w9029_,
		_w9030_,
		_w9486_,
		_w11763_
	);
	LUT2 #(
		.INIT('h8)
	) name9863 (
		_w9028_,
		_w11763_,
		_w11764_
	);
	LUT4 #(
		.INIT('h2a00)
	) name9864 (
		\s11_err_i_pad ,
		_w8955_,
		_w8956_,
		_w9483_,
		_w11765_
	);
	LUT4 #(
		.INIT('h2a00)
	) name9865 (
		\s4_err_i_pad ,
		_w8655_,
		_w8656_,
		_w9500_,
		_w11766_
	);
	LUT4 #(
		.INIT('h153f)
	) name9866 (
		_w8668_,
		_w8974_,
		_w11765_,
		_w11766_,
		_w11767_
	);
	LUT4 #(
		.INIT('h2a00)
	) name9867 (
		\s1_err_i_pad ,
		_w9103_,
		_w9104_,
		_w9295_,
		_w11768_
	);
	LUT4 #(
		.INIT('h2a00)
	) name9868 (
		\s2_err_i_pad ,
		_w9171_,
		_w9172_,
		_w9494_,
		_w11769_
	);
	LUT4 #(
		.INIT('h135f)
	) name9869 (
		_w9110_,
		_w9190_,
		_w11768_,
		_w11769_,
		_w11770_
	);
	LUT4 #(
		.INIT('h2a00)
	) name9870 (
		\s5_err_i_pad ,
		_w8699_,
		_w8700_,
		_w9387_,
		_w11771_
	);
	LUT4 #(
		.INIT('h2a00)
	) name9871 (
		\s8_err_i_pad ,
		_w8821_,
		_w8822_,
		_w9503_,
		_w11772_
	);
	LUT4 #(
		.INIT('h135f)
	) name9872 (
		_w8698_,
		_w8828_,
		_w11771_,
		_w11772_,
		_w11773_
	);
	LUT4 #(
		.INIT('h4000)
	) name9873 (
		_w11764_,
		_w11767_,
		_w11770_,
		_w11773_,
		_w11774_
	);
	LUT2 #(
		.INIT('h8)
	) name9874 (
		_w11762_,
		_w11774_,
		_w11775_
	);
	LUT4 #(
		.INIT('h70ff)
	) name9875 (
		_w2046_,
		_w2097_,
		_w11749_,
		_w11775_,
		_w11776_
	);
	LUT3 #(
		.INIT('h80)
	) name9876 (
		\s15_rty_i_pad ,
		_w1918_,
		_w11271_,
		_w11777_
	);
	LUT4 #(
		.INIT('h2a00)
	) name9877 (
		\s11_rty_i_pad ,
		_w8955_,
		_w8956_,
		_w9483_,
		_w11778_
	);
	LUT4 #(
		.INIT('h2a00)
	) name9878 (
		\s3_rty_i_pad ,
		_w9205_,
		_w9206_,
		_w9416_,
		_w11779_
	);
	LUT4 #(
		.INIT('h135f)
	) name9879 (
		_w8974_,
		_w9212_,
		_w11778_,
		_w11779_,
		_w11780_
	);
	LUT4 #(
		.INIT('h2a00)
	) name9880 (
		\s13_rty_i_pad ,
		_w9069_,
		_w9070_,
		_w9489_,
		_w11781_
	);
	LUT4 #(
		.INIT('h2a00)
	) name9881 (
		\s0_rty_i_pad ,
		_w8989_,
		_w8990_,
		_w9291_,
		_w11782_
	);
	LUT4 #(
		.INIT('h153f)
	) name9882 (
		_w9002_,
		_w9082_,
		_w11781_,
		_w11782_,
		_w11783_
	);
	LUT4 #(
		.INIT('h2a00)
	) name9883 (
		\s6_rty_i_pad ,
		_w8743_,
		_w8744_,
		_w9378_,
		_w11784_
	);
	LUT4 #(
		.INIT('h2a00)
	) name9884 (
		\s10_rty_i_pad ,
		_w8910_,
		_w8911_,
		_w9480_,
		_w11785_
	);
	LUT4 #(
		.INIT('h135f)
	) name9885 (
		_w8750_,
		_w8909_,
		_w11784_,
		_w11785_,
		_w11786_
	);
	LUT4 #(
		.INIT('h2a00)
	) name9886 (
		\s9_rty_i_pad ,
		_w8865_,
		_w8866_,
		_w9506_,
		_w11787_
	);
	LUT4 #(
		.INIT('h2a00)
	) name9887 (
		\s4_rty_i_pad ,
		_w8655_,
		_w8656_,
		_w9500_,
		_w11788_
	);
	LUT4 #(
		.INIT('h153f)
	) name9888 (
		_w8668_,
		_w8864_,
		_w11787_,
		_w11788_,
		_w11789_
	);
	LUT4 #(
		.INIT('h8000)
	) name9889 (
		_w11780_,
		_w11783_,
		_w11786_,
		_w11789_,
		_w11790_
	);
	LUT4 #(
		.INIT('h2a00)
	) name9890 (
		\s8_rty_i_pad ,
		_w8821_,
		_w8822_,
		_w9503_,
		_w11791_
	);
	LUT2 #(
		.INIT('h8)
	) name9891 (
		_w8828_,
		_w11791_,
		_w11792_
	);
	LUT4 #(
		.INIT('h2a00)
	) name9892 (
		\s14_rty_i_pad ,
		_w9137_,
		_w9138_,
		_w9497_,
		_w11793_
	);
	LUT4 #(
		.INIT('h2a00)
	) name9893 (
		\s7_rty_i_pad ,
		_w8782_,
		_w8783_,
		_w9375_,
		_w11794_
	);
	LUT4 #(
		.INIT('h153f)
	) name9894 (
		_w8795_,
		_w9144_,
		_w11793_,
		_w11794_,
		_w11795_
	);
	LUT4 #(
		.INIT('h2a00)
	) name9895 (
		\s1_rty_i_pad ,
		_w9103_,
		_w9104_,
		_w9295_,
		_w11796_
	);
	LUT4 #(
		.INIT('h2a00)
	) name9896 (
		\s2_rty_i_pad ,
		_w9171_,
		_w9172_,
		_w9494_,
		_w11797_
	);
	LUT4 #(
		.INIT('h135f)
	) name9897 (
		_w9110_,
		_w9190_,
		_w11796_,
		_w11797_,
		_w11798_
	);
	LUT4 #(
		.INIT('h2a00)
	) name9898 (
		\s5_rty_i_pad ,
		_w8699_,
		_w8700_,
		_w9387_,
		_w11799_
	);
	LUT4 #(
		.INIT('h2a00)
	) name9899 (
		\s12_rty_i_pad ,
		_w9029_,
		_w9030_,
		_w9486_,
		_w11800_
	);
	LUT4 #(
		.INIT('h135f)
	) name9900 (
		_w8698_,
		_w9028_,
		_w11799_,
		_w11800_,
		_w11801_
	);
	LUT4 #(
		.INIT('h4000)
	) name9901 (
		_w11792_,
		_w11795_,
		_w11798_,
		_w11801_,
		_w11802_
	);
	LUT2 #(
		.INIT('h8)
	) name9902 (
		_w11790_,
		_w11802_,
		_w11803_
	);
	LUT4 #(
		.INIT('h70ff)
	) name9903 (
		_w2046_,
		_w2097_,
		_w11777_,
		_w11803_,
		_w11804_
	);
	LUT3 #(
		.INIT('h80)
	) name9904 (
		_w1908_,
		_w1909_,
		_w2062_,
		_w11805_
	);
	LUT2 #(
		.INIT('h8)
	) name9905 (
		_w1907_,
		_w11805_,
		_w11806_
	);
	LUT3 #(
		.INIT('h70)
	) name9906 (
		_w2097_,
		_w8630_,
		_w11806_,
		_w11807_
	);
	LUT4 #(
		.INIT('h8000)
	) name9907 (
		\s14_ack_i_pad ,
		_w9137_,
		_w9138_,
		_w9515_,
		_w11808_
	);
	LUT4 #(
		.INIT('h8000)
	) name9908 (
		\s3_ack_i_pad ,
		_w9205_,
		_w9206_,
		_w9523_,
		_w11809_
	);
	LUT4 #(
		.INIT('h135f)
	) name9909 (
		_w9156_,
		_w9204_,
		_w11808_,
		_w11809_,
		_w11810_
	);
	LUT4 #(
		.INIT('h8000)
	) name9910 (
		\s8_ack_i_pad ,
		_w8821_,
		_w8822_,
		_w9360_,
		_w11811_
	);
	LUT4 #(
		.INIT('h8000)
	) name9911 (
		\s7_ack_i_pad ,
		_w8782_,
		_w8783_,
		_w9529_,
		_w11812_
	);
	LUT4 #(
		.INIT('h153f)
	) name9912 (
		_w8801_,
		_w8840_,
		_w11811_,
		_w11812_,
		_w11813_
	);
	LUT4 #(
		.INIT('h8000)
	) name9913 (
		\s10_ack_i_pad ,
		_w8910_,
		_w8911_,
		_w9509_,
		_w11814_
	);
	LUT4 #(
		.INIT('h8000)
	) name9914 (
		\s11_ack_i_pad ,
		_w8955_,
		_w8956_,
		_w9372_,
		_w11815_
	);
	LUT4 #(
		.INIT('h135f)
	) name9915 (
		_w8929_,
		_w8954_,
		_w11814_,
		_w11815_,
		_w11816_
	);
	LUT4 #(
		.INIT('h8000)
	) name9916 (
		\s13_ack_i_pad ,
		_w9069_,
		_w9070_,
		_w9369_,
		_w11817_
	);
	LUT4 #(
		.INIT('h8000)
	) name9917 (
		\s6_ack_i_pad ,
		_w8743_,
		_w8744_,
		_w9363_,
		_w11818_
	);
	LUT4 #(
		.INIT('h153f)
	) name9918 (
		_w8762_,
		_w9088_,
		_w11817_,
		_w11818_,
		_w11819_
	);
	LUT4 #(
		.INIT('h8000)
	) name9919 (
		_w11810_,
		_w11813_,
		_w11816_,
		_w11819_,
		_w11820_
	);
	LUT4 #(
		.INIT('h8000)
	) name9920 (
		\s12_ack_i_pad ,
		_w9029_,
		_w9030_,
		_w9512_,
		_w11821_
	);
	LUT2 #(
		.INIT('h8)
	) name9921 (
		_w9042_,
		_w11821_,
		_w11822_
	);
	LUT4 #(
		.INIT('h8000)
	) name9922 (
		\s2_ack_i_pad ,
		_w9171_,
		_w9172_,
		_w9520_,
		_w11823_
	);
	LUT4 #(
		.INIT('h8000)
	) name9923 (
		\s9_ack_i_pad ,
		_w8865_,
		_w8866_,
		_w9357_,
		_w11824_
	);
	LUT4 #(
		.INIT('h153f)
	) name9924 (
		_w8884_,
		_w9170_,
		_w11823_,
		_w11824_,
		_w11825_
	);
	LUT4 #(
		.INIT('h8000)
	) name9925 (
		\s4_ack_i_pad ,
		_w8655_,
		_w8656_,
		_w9366_,
		_w11826_
	);
	LUT4 #(
		.INIT('h8000)
	) name9926 (
		\s0_ack_i_pad ,
		_w8989_,
		_w8990_,
		_w9298_,
		_w11827_
	);
	LUT4 #(
		.INIT('h135f)
	) name9927 (
		_w8654_,
		_w8996_,
		_w11826_,
		_w11827_,
		_w11828_
	);
	LUT4 #(
		.INIT('h8000)
	) name9928 (
		\s5_ack_i_pad ,
		_w8699_,
		_w8700_,
		_w9526_,
		_w11829_
	);
	LUT4 #(
		.INIT('h8000)
	) name9929 (
		\s1_ack_i_pad ,
		_w9103_,
		_w9104_,
		_w9302_,
		_w11830_
	);
	LUT4 #(
		.INIT('h135f)
	) name9930 (
		_w8706_,
		_w9116_,
		_w11829_,
		_w11830_,
		_w11831_
	);
	LUT4 #(
		.INIT('h4000)
	) name9931 (
		_w11822_,
		_w11825_,
		_w11828_,
		_w11831_,
		_w11832_
	);
	LUT2 #(
		.INIT('h8)
	) name9932 (
		_w11820_,
		_w11832_,
		_w11833_
	);
	LUT3 #(
		.INIT('h4f)
	) name9933 (
		_w9652_,
		_w11807_,
		_w11833_,
		_w11834_
	);
	LUT3 #(
		.INIT('h80)
	) name9934 (
		_w2062_,
		_w2097_,
		_w9683_,
		_w11835_
	);
	LUT2 #(
		.INIT('h8)
	) name9935 (
		\s15_data_i[0]_pad ,
		_w2062_,
		_w11836_
	);
	LUT3 #(
		.INIT('h70)
	) name9936 (
		_w2046_,
		_w2097_,
		_w11836_,
		_w11837_
	);
	LUT4 #(
		.INIT('h135f)
	) name9937 (
		\s1_data_i[0]_pad ,
		\s8_data_i[0]_pad ,
		_w9302_,
		_w9360_,
		_w11838_
	);
	LUT4 #(
		.INIT('h153f)
	) name9938 (
		\s4_data_i[0]_pad ,
		\s6_data_i[0]_pad ,
		_w9363_,
		_w9366_,
		_w11839_
	);
	LUT4 #(
		.INIT('h153f)
	) name9939 (
		\s3_data_i[0]_pad ,
		\s9_data_i[0]_pad ,
		_w9357_,
		_w9523_,
		_w11840_
	);
	LUT4 #(
		.INIT('h135f)
	) name9940 (
		\s10_data_i[0]_pad ,
		\s7_data_i[0]_pad ,
		_w9509_,
		_w9529_,
		_w11841_
	);
	LUT4 #(
		.INIT('h8000)
	) name9941 (
		_w11838_,
		_w11839_,
		_w11840_,
		_w11841_,
		_w11842_
	);
	LUT2 #(
		.INIT('h8)
	) name9942 (
		\s11_data_i[0]_pad ,
		_w9372_,
		_w11843_
	);
	LUT4 #(
		.INIT('h135f)
	) name9943 (
		\s14_data_i[0]_pad ,
		\s2_data_i[0]_pad ,
		_w9515_,
		_w9520_,
		_w11844_
	);
	LUT4 #(
		.INIT('h135f)
	) name9944 (
		\s12_data_i[0]_pad ,
		\s5_data_i[0]_pad ,
		_w9512_,
		_w9526_,
		_w11845_
	);
	LUT4 #(
		.INIT('h135f)
	) name9945 (
		\s0_data_i[0]_pad ,
		\s13_data_i[0]_pad ,
		_w9298_,
		_w9369_,
		_w11846_
	);
	LUT4 #(
		.INIT('h4000)
	) name9946 (
		_w11843_,
		_w11844_,
		_w11845_,
		_w11846_,
		_w11847_
	);
	LUT2 #(
		.INIT('h8)
	) name9947 (
		_w11842_,
		_w11847_,
		_w11848_
	);
	LUT3 #(
		.INIT('hef)
	) name9948 (
		_w11835_,
		_w11837_,
		_w11848_,
		_w11849_
	);
	LUT3 #(
		.INIT('h80)
	) name9949 (
		_w2062_,
		_w2097_,
		_w9699_,
		_w11850_
	);
	LUT2 #(
		.INIT('h8)
	) name9950 (
		\s15_data_i[10]_pad ,
		_w2062_,
		_w11851_
	);
	LUT3 #(
		.INIT('h70)
	) name9951 (
		_w2046_,
		_w2097_,
		_w11851_,
		_w11852_
	);
	LUT4 #(
		.INIT('h135f)
	) name9952 (
		\s1_data_i[10]_pad ,
		\s8_data_i[10]_pad ,
		_w9302_,
		_w9360_,
		_w11853_
	);
	LUT4 #(
		.INIT('h153f)
	) name9953 (
		\s4_data_i[10]_pad ,
		\s6_data_i[10]_pad ,
		_w9363_,
		_w9366_,
		_w11854_
	);
	LUT4 #(
		.INIT('h153f)
	) name9954 (
		\s3_data_i[10]_pad ,
		\s9_data_i[10]_pad ,
		_w9357_,
		_w9523_,
		_w11855_
	);
	LUT4 #(
		.INIT('h135f)
	) name9955 (
		\s10_data_i[10]_pad ,
		\s7_data_i[10]_pad ,
		_w9509_,
		_w9529_,
		_w11856_
	);
	LUT4 #(
		.INIT('h8000)
	) name9956 (
		_w11853_,
		_w11854_,
		_w11855_,
		_w11856_,
		_w11857_
	);
	LUT2 #(
		.INIT('h8)
	) name9957 (
		\s11_data_i[10]_pad ,
		_w9372_,
		_w11858_
	);
	LUT4 #(
		.INIT('h135f)
	) name9958 (
		\s14_data_i[10]_pad ,
		\s2_data_i[10]_pad ,
		_w9515_,
		_w9520_,
		_w11859_
	);
	LUT4 #(
		.INIT('h135f)
	) name9959 (
		\s12_data_i[10]_pad ,
		\s5_data_i[10]_pad ,
		_w9512_,
		_w9526_,
		_w11860_
	);
	LUT4 #(
		.INIT('h135f)
	) name9960 (
		\s0_data_i[10]_pad ,
		\s13_data_i[10]_pad ,
		_w9298_,
		_w9369_,
		_w11861_
	);
	LUT4 #(
		.INIT('h4000)
	) name9961 (
		_w11858_,
		_w11859_,
		_w11860_,
		_w11861_,
		_w11862_
	);
	LUT2 #(
		.INIT('h8)
	) name9962 (
		_w11857_,
		_w11862_,
		_w11863_
	);
	LUT3 #(
		.INIT('hef)
	) name9963 (
		_w11850_,
		_w11852_,
		_w11863_,
		_w11864_
	);
	LUT3 #(
		.INIT('h80)
	) name9964 (
		_w2062_,
		_w2097_,
		_w9715_,
		_w11865_
	);
	LUT2 #(
		.INIT('h8)
	) name9965 (
		\s15_data_i[11]_pad ,
		_w2062_,
		_w11866_
	);
	LUT3 #(
		.INIT('h70)
	) name9966 (
		_w2046_,
		_w2097_,
		_w11866_,
		_w11867_
	);
	LUT4 #(
		.INIT('h135f)
	) name9967 (
		\s1_data_i[11]_pad ,
		\s8_data_i[11]_pad ,
		_w9302_,
		_w9360_,
		_w11868_
	);
	LUT4 #(
		.INIT('h153f)
	) name9968 (
		\s4_data_i[11]_pad ,
		\s6_data_i[11]_pad ,
		_w9363_,
		_w9366_,
		_w11869_
	);
	LUT4 #(
		.INIT('h153f)
	) name9969 (
		\s3_data_i[11]_pad ,
		\s9_data_i[11]_pad ,
		_w9357_,
		_w9523_,
		_w11870_
	);
	LUT4 #(
		.INIT('h135f)
	) name9970 (
		\s10_data_i[11]_pad ,
		\s7_data_i[11]_pad ,
		_w9509_,
		_w9529_,
		_w11871_
	);
	LUT4 #(
		.INIT('h8000)
	) name9971 (
		_w11868_,
		_w11869_,
		_w11870_,
		_w11871_,
		_w11872_
	);
	LUT2 #(
		.INIT('h8)
	) name9972 (
		\s11_data_i[11]_pad ,
		_w9372_,
		_w11873_
	);
	LUT4 #(
		.INIT('h135f)
	) name9973 (
		\s14_data_i[11]_pad ,
		\s2_data_i[11]_pad ,
		_w9515_,
		_w9520_,
		_w11874_
	);
	LUT4 #(
		.INIT('h135f)
	) name9974 (
		\s12_data_i[11]_pad ,
		\s5_data_i[11]_pad ,
		_w9512_,
		_w9526_,
		_w11875_
	);
	LUT4 #(
		.INIT('h135f)
	) name9975 (
		\s0_data_i[11]_pad ,
		\s13_data_i[11]_pad ,
		_w9298_,
		_w9369_,
		_w11876_
	);
	LUT4 #(
		.INIT('h4000)
	) name9976 (
		_w11873_,
		_w11874_,
		_w11875_,
		_w11876_,
		_w11877_
	);
	LUT2 #(
		.INIT('h8)
	) name9977 (
		_w11872_,
		_w11877_,
		_w11878_
	);
	LUT3 #(
		.INIT('hef)
	) name9978 (
		_w11865_,
		_w11867_,
		_w11878_,
		_w11879_
	);
	LUT3 #(
		.INIT('h80)
	) name9979 (
		_w2062_,
		_w2097_,
		_w9731_,
		_w11880_
	);
	LUT2 #(
		.INIT('h8)
	) name9980 (
		\s15_data_i[12]_pad ,
		_w2062_,
		_w11881_
	);
	LUT3 #(
		.INIT('h70)
	) name9981 (
		_w2046_,
		_w2097_,
		_w11881_,
		_w11882_
	);
	LUT4 #(
		.INIT('h135f)
	) name9982 (
		\s1_data_i[12]_pad ,
		\s8_data_i[12]_pad ,
		_w9302_,
		_w9360_,
		_w11883_
	);
	LUT4 #(
		.INIT('h153f)
	) name9983 (
		\s4_data_i[12]_pad ,
		\s6_data_i[12]_pad ,
		_w9363_,
		_w9366_,
		_w11884_
	);
	LUT4 #(
		.INIT('h153f)
	) name9984 (
		\s3_data_i[12]_pad ,
		\s9_data_i[12]_pad ,
		_w9357_,
		_w9523_,
		_w11885_
	);
	LUT4 #(
		.INIT('h135f)
	) name9985 (
		\s10_data_i[12]_pad ,
		\s7_data_i[12]_pad ,
		_w9509_,
		_w9529_,
		_w11886_
	);
	LUT4 #(
		.INIT('h8000)
	) name9986 (
		_w11883_,
		_w11884_,
		_w11885_,
		_w11886_,
		_w11887_
	);
	LUT2 #(
		.INIT('h8)
	) name9987 (
		\s11_data_i[12]_pad ,
		_w9372_,
		_w11888_
	);
	LUT4 #(
		.INIT('h135f)
	) name9988 (
		\s14_data_i[12]_pad ,
		\s2_data_i[12]_pad ,
		_w9515_,
		_w9520_,
		_w11889_
	);
	LUT4 #(
		.INIT('h135f)
	) name9989 (
		\s12_data_i[12]_pad ,
		\s5_data_i[12]_pad ,
		_w9512_,
		_w9526_,
		_w11890_
	);
	LUT4 #(
		.INIT('h135f)
	) name9990 (
		\s0_data_i[12]_pad ,
		\s13_data_i[12]_pad ,
		_w9298_,
		_w9369_,
		_w11891_
	);
	LUT4 #(
		.INIT('h4000)
	) name9991 (
		_w11888_,
		_w11889_,
		_w11890_,
		_w11891_,
		_w11892_
	);
	LUT2 #(
		.INIT('h8)
	) name9992 (
		_w11887_,
		_w11892_,
		_w11893_
	);
	LUT3 #(
		.INIT('hef)
	) name9993 (
		_w11880_,
		_w11882_,
		_w11893_,
		_w11894_
	);
	LUT3 #(
		.INIT('h80)
	) name9994 (
		_w2062_,
		_w2097_,
		_w9747_,
		_w11895_
	);
	LUT2 #(
		.INIT('h8)
	) name9995 (
		\s15_data_i[13]_pad ,
		_w2062_,
		_w11896_
	);
	LUT3 #(
		.INIT('h70)
	) name9996 (
		_w2046_,
		_w2097_,
		_w11896_,
		_w11897_
	);
	LUT4 #(
		.INIT('h135f)
	) name9997 (
		\s1_data_i[13]_pad ,
		\s8_data_i[13]_pad ,
		_w9302_,
		_w9360_,
		_w11898_
	);
	LUT4 #(
		.INIT('h153f)
	) name9998 (
		\s4_data_i[13]_pad ,
		\s6_data_i[13]_pad ,
		_w9363_,
		_w9366_,
		_w11899_
	);
	LUT4 #(
		.INIT('h153f)
	) name9999 (
		\s3_data_i[13]_pad ,
		\s9_data_i[13]_pad ,
		_w9357_,
		_w9523_,
		_w11900_
	);
	LUT4 #(
		.INIT('h135f)
	) name10000 (
		\s10_data_i[13]_pad ,
		\s7_data_i[13]_pad ,
		_w9509_,
		_w9529_,
		_w11901_
	);
	LUT4 #(
		.INIT('h8000)
	) name10001 (
		_w11898_,
		_w11899_,
		_w11900_,
		_w11901_,
		_w11902_
	);
	LUT2 #(
		.INIT('h8)
	) name10002 (
		\s11_data_i[13]_pad ,
		_w9372_,
		_w11903_
	);
	LUT4 #(
		.INIT('h135f)
	) name10003 (
		\s14_data_i[13]_pad ,
		\s2_data_i[13]_pad ,
		_w9515_,
		_w9520_,
		_w11904_
	);
	LUT4 #(
		.INIT('h135f)
	) name10004 (
		\s12_data_i[13]_pad ,
		\s5_data_i[13]_pad ,
		_w9512_,
		_w9526_,
		_w11905_
	);
	LUT4 #(
		.INIT('h135f)
	) name10005 (
		\s0_data_i[13]_pad ,
		\s13_data_i[13]_pad ,
		_w9298_,
		_w9369_,
		_w11906_
	);
	LUT4 #(
		.INIT('h4000)
	) name10006 (
		_w11903_,
		_w11904_,
		_w11905_,
		_w11906_,
		_w11907_
	);
	LUT2 #(
		.INIT('h8)
	) name10007 (
		_w11902_,
		_w11907_,
		_w11908_
	);
	LUT3 #(
		.INIT('hef)
	) name10008 (
		_w11895_,
		_w11897_,
		_w11908_,
		_w11909_
	);
	LUT3 #(
		.INIT('h80)
	) name10009 (
		_w2062_,
		_w2097_,
		_w9763_,
		_w11910_
	);
	LUT2 #(
		.INIT('h8)
	) name10010 (
		\s15_data_i[14]_pad ,
		_w2062_,
		_w11911_
	);
	LUT3 #(
		.INIT('h70)
	) name10011 (
		_w2046_,
		_w2097_,
		_w11911_,
		_w11912_
	);
	LUT4 #(
		.INIT('h135f)
	) name10012 (
		\s1_data_i[14]_pad ,
		\s8_data_i[14]_pad ,
		_w9302_,
		_w9360_,
		_w11913_
	);
	LUT4 #(
		.INIT('h135f)
	) name10013 (
		\s0_data_i[14]_pad ,
		\s10_data_i[14]_pad ,
		_w9298_,
		_w9509_,
		_w11914_
	);
	LUT4 #(
		.INIT('h153f)
	) name10014 (
		\s3_data_i[14]_pad ,
		\s6_data_i[14]_pad ,
		_w9363_,
		_w9523_,
		_w11915_
	);
	LUT4 #(
		.INIT('h135f)
	) name10015 (
		\s4_data_i[14]_pad ,
		\s7_data_i[14]_pad ,
		_w9366_,
		_w9529_,
		_w11916_
	);
	LUT4 #(
		.INIT('h8000)
	) name10016 (
		_w11913_,
		_w11914_,
		_w11915_,
		_w11916_,
		_w11917_
	);
	LUT2 #(
		.INIT('h8)
	) name10017 (
		\s11_data_i[14]_pad ,
		_w9372_,
		_w11918_
	);
	LUT4 #(
		.INIT('h135f)
	) name10018 (
		\s14_data_i[14]_pad ,
		\s2_data_i[14]_pad ,
		_w9515_,
		_w9520_,
		_w11919_
	);
	LUT4 #(
		.INIT('h135f)
	) name10019 (
		\s12_data_i[14]_pad ,
		\s5_data_i[14]_pad ,
		_w9512_,
		_w9526_,
		_w11920_
	);
	LUT4 #(
		.INIT('h153f)
	) name10020 (
		\s13_data_i[14]_pad ,
		\s9_data_i[14]_pad ,
		_w9357_,
		_w9369_,
		_w11921_
	);
	LUT4 #(
		.INIT('h4000)
	) name10021 (
		_w11918_,
		_w11919_,
		_w11920_,
		_w11921_,
		_w11922_
	);
	LUT2 #(
		.INIT('h8)
	) name10022 (
		_w11917_,
		_w11922_,
		_w11923_
	);
	LUT3 #(
		.INIT('hef)
	) name10023 (
		_w11910_,
		_w11912_,
		_w11923_,
		_w11924_
	);
	LUT3 #(
		.INIT('h80)
	) name10024 (
		_w2062_,
		_w2097_,
		_w9779_,
		_w11925_
	);
	LUT2 #(
		.INIT('h8)
	) name10025 (
		\s15_data_i[15]_pad ,
		_w2062_,
		_w11926_
	);
	LUT3 #(
		.INIT('h70)
	) name10026 (
		_w2046_,
		_w2097_,
		_w11926_,
		_w11927_
	);
	LUT4 #(
		.INIT('h135f)
	) name10027 (
		\s1_data_i[15]_pad ,
		\s8_data_i[15]_pad ,
		_w9302_,
		_w9360_,
		_w11928_
	);
	LUT4 #(
		.INIT('h153f)
	) name10028 (
		\s4_data_i[15]_pad ,
		\s6_data_i[15]_pad ,
		_w9363_,
		_w9366_,
		_w11929_
	);
	LUT4 #(
		.INIT('h153f)
	) name10029 (
		\s3_data_i[15]_pad ,
		\s9_data_i[15]_pad ,
		_w9357_,
		_w9523_,
		_w11930_
	);
	LUT4 #(
		.INIT('h135f)
	) name10030 (
		\s10_data_i[15]_pad ,
		\s7_data_i[15]_pad ,
		_w9509_,
		_w9529_,
		_w11931_
	);
	LUT4 #(
		.INIT('h8000)
	) name10031 (
		_w11928_,
		_w11929_,
		_w11930_,
		_w11931_,
		_w11932_
	);
	LUT2 #(
		.INIT('h8)
	) name10032 (
		\s11_data_i[15]_pad ,
		_w9372_,
		_w11933_
	);
	LUT4 #(
		.INIT('h135f)
	) name10033 (
		\s14_data_i[15]_pad ,
		\s2_data_i[15]_pad ,
		_w9515_,
		_w9520_,
		_w11934_
	);
	LUT4 #(
		.INIT('h135f)
	) name10034 (
		\s12_data_i[15]_pad ,
		\s5_data_i[15]_pad ,
		_w9512_,
		_w9526_,
		_w11935_
	);
	LUT4 #(
		.INIT('h135f)
	) name10035 (
		\s0_data_i[15]_pad ,
		\s13_data_i[15]_pad ,
		_w9298_,
		_w9369_,
		_w11936_
	);
	LUT4 #(
		.INIT('h4000)
	) name10036 (
		_w11933_,
		_w11934_,
		_w11935_,
		_w11936_,
		_w11937_
	);
	LUT2 #(
		.INIT('h8)
	) name10037 (
		_w11932_,
		_w11937_,
		_w11938_
	);
	LUT3 #(
		.INIT('hef)
	) name10038 (
		_w11925_,
		_w11927_,
		_w11938_,
		_w11939_
	);
	LUT2 #(
		.INIT('h8)
	) name10039 (
		\s15_data_i[16]_pad ,
		_w2062_,
		_w11940_
	);
	LUT4 #(
		.INIT('h135f)
	) name10040 (
		\s1_data_i[16]_pad ,
		\s8_data_i[16]_pad ,
		_w9302_,
		_w9360_,
		_w11941_
	);
	LUT4 #(
		.INIT('h153f)
	) name10041 (
		\s4_data_i[16]_pad ,
		\s6_data_i[16]_pad ,
		_w9363_,
		_w9366_,
		_w11942_
	);
	LUT4 #(
		.INIT('h153f)
	) name10042 (
		\s3_data_i[16]_pad ,
		\s9_data_i[16]_pad ,
		_w9357_,
		_w9523_,
		_w11943_
	);
	LUT4 #(
		.INIT('h135f)
	) name10043 (
		\s10_data_i[16]_pad ,
		\s7_data_i[16]_pad ,
		_w9509_,
		_w9529_,
		_w11944_
	);
	LUT4 #(
		.INIT('h8000)
	) name10044 (
		_w11941_,
		_w11942_,
		_w11943_,
		_w11944_,
		_w11945_
	);
	LUT2 #(
		.INIT('h8)
	) name10045 (
		\s11_data_i[16]_pad ,
		_w9372_,
		_w11946_
	);
	LUT4 #(
		.INIT('h135f)
	) name10046 (
		\s14_data_i[16]_pad ,
		\s2_data_i[16]_pad ,
		_w9515_,
		_w9520_,
		_w11947_
	);
	LUT4 #(
		.INIT('h135f)
	) name10047 (
		\s12_data_i[16]_pad ,
		\s5_data_i[16]_pad ,
		_w9512_,
		_w9526_,
		_w11948_
	);
	LUT4 #(
		.INIT('h135f)
	) name10048 (
		\s0_data_i[16]_pad ,
		\s13_data_i[16]_pad ,
		_w9298_,
		_w9369_,
		_w11949_
	);
	LUT4 #(
		.INIT('h4000)
	) name10049 (
		_w11946_,
		_w11947_,
		_w11948_,
		_w11949_,
		_w11950_
	);
	LUT2 #(
		.INIT('h8)
	) name10050 (
		_w11945_,
		_w11950_,
		_w11951_
	);
	LUT4 #(
		.INIT('h70ff)
	) name10051 (
		_w2046_,
		_w2097_,
		_w11940_,
		_w11951_,
		_w11952_
	);
	LUT2 #(
		.INIT('h8)
	) name10052 (
		\s15_data_i[17]_pad ,
		_w2062_,
		_w11953_
	);
	LUT4 #(
		.INIT('h135f)
	) name10053 (
		\s1_data_i[17]_pad ,
		\s8_data_i[17]_pad ,
		_w9302_,
		_w9360_,
		_w11954_
	);
	LUT4 #(
		.INIT('h153f)
	) name10054 (
		\s4_data_i[17]_pad ,
		\s6_data_i[17]_pad ,
		_w9363_,
		_w9366_,
		_w11955_
	);
	LUT4 #(
		.INIT('h153f)
	) name10055 (
		\s3_data_i[17]_pad ,
		\s9_data_i[17]_pad ,
		_w9357_,
		_w9523_,
		_w11956_
	);
	LUT4 #(
		.INIT('h135f)
	) name10056 (
		\s10_data_i[17]_pad ,
		\s7_data_i[17]_pad ,
		_w9509_,
		_w9529_,
		_w11957_
	);
	LUT4 #(
		.INIT('h8000)
	) name10057 (
		_w11954_,
		_w11955_,
		_w11956_,
		_w11957_,
		_w11958_
	);
	LUT2 #(
		.INIT('h8)
	) name10058 (
		\s11_data_i[17]_pad ,
		_w9372_,
		_w11959_
	);
	LUT4 #(
		.INIT('h135f)
	) name10059 (
		\s14_data_i[17]_pad ,
		\s2_data_i[17]_pad ,
		_w9515_,
		_w9520_,
		_w11960_
	);
	LUT4 #(
		.INIT('h135f)
	) name10060 (
		\s12_data_i[17]_pad ,
		\s5_data_i[17]_pad ,
		_w9512_,
		_w9526_,
		_w11961_
	);
	LUT4 #(
		.INIT('h135f)
	) name10061 (
		\s0_data_i[17]_pad ,
		\s13_data_i[17]_pad ,
		_w9298_,
		_w9369_,
		_w11962_
	);
	LUT4 #(
		.INIT('h4000)
	) name10062 (
		_w11959_,
		_w11960_,
		_w11961_,
		_w11962_,
		_w11963_
	);
	LUT2 #(
		.INIT('h8)
	) name10063 (
		_w11958_,
		_w11963_,
		_w11964_
	);
	LUT4 #(
		.INIT('h70ff)
	) name10064 (
		_w2046_,
		_w2097_,
		_w11953_,
		_w11964_,
		_w11965_
	);
	LUT2 #(
		.INIT('h8)
	) name10065 (
		\s15_data_i[18]_pad ,
		_w2062_,
		_w11966_
	);
	LUT4 #(
		.INIT('h153f)
	) name10066 (
		\s12_data_i[18]_pad ,
		\s1_data_i[18]_pad ,
		_w9302_,
		_w9512_,
		_w11967_
	);
	LUT4 #(
		.INIT('h153f)
	) name10067 (
		\s4_data_i[18]_pad ,
		\s6_data_i[18]_pad ,
		_w9363_,
		_w9366_,
		_w11968_
	);
	LUT4 #(
		.INIT('h153f)
	) name10068 (
		\s3_data_i[18]_pad ,
		\s9_data_i[18]_pad ,
		_w9357_,
		_w9523_,
		_w11969_
	);
	LUT4 #(
		.INIT('h135f)
	) name10069 (
		\s10_data_i[18]_pad ,
		\s7_data_i[18]_pad ,
		_w9509_,
		_w9529_,
		_w11970_
	);
	LUT4 #(
		.INIT('h8000)
	) name10070 (
		_w11967_,
		_w11968_,
		_w11969_,
		_w11970_,
		_w11971_
	);
	LUT2 #(
		.INIT('h8)
	) name10071 (
		\s14_data_i[18]_pad ,
		_w9515_,
		_w11972_
	);
	LUT4 #(
		.INIT('h135f)
	) name10072 (
		\s11_data_i[18]_pad ,
		\s2_data_i[18]_pad ,
		_w9372_,
		_w9520_,
		_w11973_
	);
	LUT4 #(
		.INIT('h153f)
	) name10073 (
		\s5_data_i[18]_pad ,
		\s8_data_i[18]_pad ,
		_w9360_,
		_w9526_,
		_w11974_
	);
	LUT4 #(
		.INIT('h135f)
	) name10074 (
		\s0_data_i[18]_pad ,
		\s13_data_i[18]_pad ,
		_w9298_,
		_w9369_,
		_w11975_
	);
	LUT4 #(
		.INIT('h4000)
	) name10075 (
		_w11972_,
		_w11973_,
		_w11974_,
		_w11975_,
		_w11976_
	);
	LUT2 #(
		.INIT('h8)
	) name10076 (
		_w11971_,
		_w11976_,
		_w11977_
	);
	LUT4 #(
		.INIT('h70ff)
	) name10077 (
		_w2046_,
		_w2097_,
		_w11966_,
		_w11977_,
		_w11978_
	);
	LUT2 #(
		.INIT('h8)
	) name10078 (
		\s15_data_i[19]_pad ,
		_w2062_,
		_w11979_
	);
	LUT4 #(
		.INIT('h135f)
	) name10079 (
		\s1_data_i[19]_pad ,
		\s8_data_i[19]_pad ,
		_w9302_,
		_w9360_,
		_w11980_
	);
	LUT4 #(
		.INIT('h153f)
	) name10080 (
		\s4_data_i[19]_pad ,
		\s6_data_i[19]_pad ,
		_w9363_,
		_w9366_,
		_w11981_
	);
	LUT4 #(
		.INIT('h153f)
	) name10081 (
		\s3_data_i[19]_pad ,
		\s9_data_i[19]_pad ,
		_w9357_,
		_w9523_,
		_w11982_
	);
	LUT4 #(
		.INIT('h135f)
	) name10082 (
		\s10_data_i[19]_pad ,
		\s7_data_i[19]_pad ,
		_w9509_,
		_w9529_,
		_w11983_
	);
	LUT4 #(
		.INIT('h8000)
	) name10083 (
		_w11980_,
		_w11981_,
		_w11982_,
		_w11983_,
		_w11984_
	);
	LUT2 #(
		.INIT('h8)
	) name10084 (
		\s11_data_i[19]_pad ,
		_w9372_,
		_w11985_
	);
	LUT4 #(
		.INIT('h135f)
	) name10085 (
		\s14_data_i[19]_pad ,
		\s2_data_i[19]_pad ,
		_w9515_,
		_w9520_,
		_w11986_
	);
	LUT4 #(
		.INIT('h135f)
	) name10086 (
		\s12_data_i[19]_pad ,
		\s5_data_i[19]_pad ,
		_w9512_,
		_w9526_,
		_w11987_
	);
	LUT4 #(
		.INIT('h135f)
	) name10087 (
		\s0_data_i[19]_pad ,
		\s13_data_i[19]_pad ,
		_w9298_,
		_w9369_,
		_w11988_
	);
	LUT4 #(
		.INIT('h4000)
	) name10088 (
		_w11985_,
		_w11986_,
		_w11987_,
		_w11988_,
		_w11989_
	);
	LUT2 #(
		.INIT('h8)
	) name10089 (
		_w11984_,
		_w11989_,
		_w11990_
	);
	LUT4 #(
		.INIT('h70ff)
	) name10090 (
		_w2046_,
		_w2097_,
		_w11979_,
		_w11990_,
		_w11991_
	);
	LUT3 #(
		.INIT('h80)
	) name10091 (
		_w2062_,
		_w2097_,
		_w9847_,
		_w11992_
	);
	LUT2 #(
		.INIT('h8)
	) name10092 (
		\s15_data_i[1]_pad ,
		_w2062_,
		_w11993_
	);
	LUT3 #(
		.INIT('h70)
	) name10093 (
		_w2046_,
		_w2097_,
		_w11993_,
		_w11994_
	);
	LUT4 #(
		.INIT('h135f)
	) name10094 (
		\s1_data_i[1]_pad ,
		\s8_data_i[1]_pad ,
		_w9302_,
		_w9360_,
		_w11995_
	);
	LUT4 #(
		.INIT('h153f)
	) name10095 (
		\s4_data_i[1]_pad ,
		\s6_data_i[1]_pad ,
		_w9363_,
		_w9366_,
		_w11996_
	);
	LUT4 #(
		.INIT('h153f)
	) name10096 (
		\s3_data_i[1]_pad ,
		\s9_data_i[1]_pad ,
		_w9357_,
		_w9523_,
		_w11997_
	);
	LUT4 #(
		.INIT('h135f)
	) name10097 (
		\s10_data_i[1]_pad ,
		\s7_data_i[1]_pad ,
		_w9509_,
		_w9529_,
		_w11998_
	);
	LUT4 #(
		.INIT('h8000)
	) name10098 (
		_w11995_,
		_w11996_,
		_w11997_,
		_w11998_,
		_w11999_
	);
	LUT2 #(
		.INIT('h8)
	) name10099 (
		\s11_data_i[1]_pad ,
		_w9372_,
		_w12000_
	);
	LUT4 #(
		.INIT('h135f)
	) name10100 (
		\s14_data_i[1]_pad ,
		\s2_data_i[1]_pad ,
		_w9515_,
		_w9520_,
		_w12001_
	);
	LUT4 #(
		.INIT('h135f)
	) name10101 (
		\s12_data_i[1]_pad ,
		\s5_data_i[1]_pad ,
		_w9512_,
		_w9526_,
		_w12002_
	);
	LUT4 #(
		.INIT('h135f)
	) name10102 (
		\s0_data_i[1]_pad ,
		\s13_data_i[1]_pad ,
		_w9298_,
		_w9369_,
		_w12003_
	);
	LUT4 #(
		.INIT('h4000)
	) name10103 (
		_w12000_,
		_w12001_,
		_w12002_,
		_w12003_,
		_w12004_
	);
	LUT2 #(
		.INIT('h8)
	) name10104 (
		_w11999_,
		_w12004_,
		_w12005_
	);
	LUT3 #(
		.INIT('hef)
	) name10105 (
		_w11992_,
		_w11994_,
		_w12005_,
		_w12006_
	);
	LUT2 #(
		.INIT('h8)
	) name10106 (
		\s15_data_i[20]_pad ,
		_w2062_,
		_w12007_
	);
	LUT4 #(
		.INIT('h135f)
	) name10107 (
		\s1_data_i[20]_pad ,
		\s8_data_i[20]_pad ,
		_w9302_,
		_w9360_,
		_w12008_
	);
	LUT4 #(
		.INIT('h153f)
	) name10108 (
		\s4_data_i[20]_pad ,
		\s6_data_i[20]_pad ,
		_w9363_,
		_w9366_,
		_w12009_
	);
	LUT4 #(
		.INIT('h153f)
	) name10109 (
		\s3_data_i[20]_pad ,
		\s9_data_i[20]_pad ,
		_w9357_,
		_w9523_,
		_w12010_
	);
	LUT4 #(
		.INIT('h135f)
	) name10110 (
		\s10_data_i[20]_pad ,
		\s7_data_i[20]_pad ,
		_w9509_,
		_w9529_,
		_w12011_
	);
	LUT4 #(
		.INIT('h8000)
	) name10111 (
		_w12008_,
		_w12009_,
		_w12010_,
		_w12011_,
		_w12012_
	);
	LUT2 #(
		.INIT('h8)
	) name10112 (
		\s11_data_i[20]_pad ,
		_w9372_,
		_w12013_
	);
	LUT4 #(
		.INIT('h135f)
	) name10113 (
		\s14_data_i[20]_pad ,
		\s2_data_i[20]_pad ,
		_w9515_,
		_w9520_,
		_w12014_
	);
	LUT4 #(
		.INIT('h135f)
	) name10114 (
		\s12_data_i[20]_pad ,
		\s5_data_i[20]_pad ,
		_w9512_,
		_w9526_,
		_w12015_
	);
	LUT4 #(
		.INIT('h135f)
	) name10115 (
		\s0_data_i[20]_pad ,
		\s13_data_i[20]_pad ,
		_w9298_,
		_w9369_,
		_w12016_
	);
	LUT4 #(
		.INIT('h4000)
	) name10116 (
		_w12013_,
		_w12014_,
		_w12015_,
		_w12016_,
		_w12017_
	);
	LUT2 #(
		.INIT('h8)
	) name10117 (
		_w12012_,
		_w12017_,
		_w12018_
	);
	LUT4 #(
		.INIT('h70ff)
	) name10118 (
		_w2046_,
		_w2097_,
		_w12007_,
		_w12018_,
		_w12019_
	);
	LUT2 #(
		.INIT('h8)
	) name10119 (
		\s15_data_i[21]_pad ,
		_w2062_,
		_w12020_
	);
	LUT4 #(
		.INIT('h135f)
	) name10120 (
		\s1_data_i[21]_pad ,
		\s8_data_i[21]_pad ,
		_w9302_,
		_w9360_,
		_w12021_
	);
	LUT4 #(
		.INIT('h153f)
	) name10121 (
		\s4_data_i[21]_pad ,
		\s6_data_i[21]_pad ,
		_w9363_,
		_w9366_,
		_w12022_
	);
	LUT4 #(
		.INIT('h153f)
	) name10122 (
		\s3_data_i[21]_pad ,
		\s9_data_i[21]_pad ,
		_w9357_,
		_w9523_,
		_w12023_
	);
	LUT4 #(
		.INIT('h135f)
	) name10123 (
		\s10_data_i[21]_pad ,
		\s7_data_i[21]_pad ,
		_w9509_,
		_w9529_,
		_w12024_
	);
	LUT4 #(
		.INIT('h8000)
	) name10124 (
		_w12021_,
		_w12022_,
		_w12023_,
		_w12024_,
		_w12025_
	);
	LUT2 #(
		.INIT('h8)
	) name10125 (
		\s11_data_i[21]_pad ,
		_w9372_,
		_w12026_
	);
	LUT4 #(
		.INIT('h135f)
	) name10126 (
		\s14_data_i[21]_pad ,
		\s2_data_i[21]_pad ,
		_w9515_,
		_w9520_,
		_w12027_
	);
	LUT4 #(
		.INIT('h135f)
	) name10127 (
		\s12_data_i[21]_pad ,
		\s5_data_i[21]_pad ,
		_w9512_,
		_w9526_,
		_w12028_
	);
	LUT4 #(
		.INIT('h135f)
	) name10128 (
		\s0_data_i[21]_pad ,
		\s13_data_i[21]_pad ,
		_w9298_,
		_w9369_,
		_w12029_
	);
	LUT4 #(
		.INIT('h4000)
	) name10129 (
		_w12026_,
		_w12027_,
		_w12028_,
		_w12029_,
		_w12030_
	);
	LUT2 #(
		.INIT('h8)
	) name10130 (
		_w12025_,
		_w12030_,
		_w12031_
	);
	LUT4 #(
		.INIT('h70ff)
	) name10131 (
		_w2046_,
		_w2097_,
		_w12020_,
		_w12031_,
		_w12032_
	);
	LUT2 #(
		.INIT('h8)
	) name10132 (
		\s15_data_i[22]_pad ,
		_w2062_,
		_w12033_
	);
	LUT4 #(
		.INIT('h135f)
	) name10133 (
		\s1_data_i[22]_pad ,
		\s8_data_i[22]_pad ,
		_w9302_,
		_w9360_,
		_w12034_
	);
	LUT4 #(
		.INIT('h153f)
	) name10134 (
		\s4_data_i[22]_pad ,
		\s6_data_i[22]_pad ,
		_w9363_,
		_w9366_,
		_w12035_
	);
	LUT4 #(
		.INIT('h153f)
	) name10135 (
		\s3_data_i[22]_pad ,
		\s9_data_i[22]_pad ,
		_w9357_,
		_w9523_,
		_w12036_
	);
	LUT4 #(
		.INIT('h135f)
	) name10136 (
		\s10_data_i[22]_pad ,
		\s7_data_i[22]_pad ,
		_w9509_,
		_w9529_,
		_w12037_
	);
	LUT4 #(
		.INIT('h8000)
	) name10137 (
		_w12034_,
		_w12035_,
		_w12036_,
		_w12037_,
		_w12038_
	);
	LUT2 #(
		.INIT('h8)
	) name10138 (
		\s11_data_i[22]_pad ,
		_w9372_,
		_w12039_
	);
	LUT4 #(
		.INIT('h135f)
	) name10139 (
		\s14_data_i[22]_pad ,
		\s2_data_i[22]_pad ,
		_w9515_,
		_w9520_,
		_w12040_
	);
	LUT4 #(
		.INIT('h135f)
	) name10140 (
		\s12_data_i[22]_pad ,
		\s5_data_i[22]_pad ,
		_w9512_,
		_w9526_,
		_w12041_
	);
	LUT4 #(
		.INIT('h135f)
	) name10141 (
		\s0_data_i[22]_pad ,
		\s13_data_i[22]_pad ,
		_w9298_,
		_w9369_,
		_w12042_
	);
	LUT4 #(
		.INIT('h4000)
	) name10142 (
		_w12039_,
		_w12040_,
		_w12041_,
		_w12042_,
		_w12043_
	);
	LUT2 #(
		.INIT('h8)
	) name10143 (
		_w12038_,
		_w12043_,
		_w12044_
	);
	LUT4 #(
		.INIT('h70ff)
	) name10144 (
		_w2046_,
		_w2097_,
		_w12033_,
		_w12044_,
		_w12045_
	);
	LUT2 #(
		.INIT('h8)
	) name10145 (
		\s15_data_i[23]_pad ,
		_w2062_,
		_w12046_
	);
	LUT4 #(
		.INIT('h135f)
	) name10146 (
		\s1_data_i[23]_pad ,
		\s8_data_i[23]_pad ,
		_w9302_,
		_w9360_,
		_w12047_
	);
	LUT4 #(
		.INIT('h153f)
	) name10147 (
		\s4_data_i[23]_pad ,
		\s6_data_i[23]_pad ,
		_w9363_,
		_w9366_,
		_w12048_
	);
	LUT4 #(
		.INIT('h153f)
	) name10148 (
		\s3_data_i[23]_pad ,
		\s9_data_i[23]_pad ,
		_w9357_,
		_w9523_,
		_w12049_
	);
	LUT4 #(
		.INIT('h135f)
	) name10149 (
		\s10_data_i[23]_pad ,
		\s7_data_i[23]_pad ,
		_w9509_,
		_w9529_,
		_w12050_
	);
	LUT4 #(
		.INIT('h8000)
	) name10150 (
		_w12047_,
		_w12048_,
		_w12049_,
		_w12050_,
		_w12051_
	);
	LUT2 #(
		.INIT('h8)
	) name10151 (
		\s11_data_i[23]_pad ,
		_w9372_,
		_w12052_
	);
	LUT4 #(
		.INIT('h135f)
	) name10152 (
		\s14_data_i[23]_pad ,
		\s2_data_i[23]_pad ,
		_w9515_,
		_w9520_,
		_w12053_
	);
	LUT4 #(
		.INIT('h135f)
	) name10153 (
		\s12_data_i[23]_pad ,
		\s5_data_i[23]_pad ,
		_w9512_,
		_w9526_,
		_w12054_
	);
	LUT4 #(
		.INIT('h135f)
	) name10154 (
		\s0_data_i[23]_pad ,
		\s13_data_i[23]_pad ,
		_w9298_,
		_w9369_,
		_w12055_
	);
	LUT4 #(
		.INIT('h4000)
	) name10155 (
		_w12052_,
		_w12053_,
		_w12054_,
		_w12055_,
		_w12056_
	);
	LUT2 #(
		.INIT('h8)
	) name10156 (
		_w12051_,
		_w12056_,
		_w12057_
	);
	LUT4 #(
		.INIT('h70ff)
	) name10157 (
		_w2046_,
		_w2097_,
		_w12046_,
		_w12057_,
		_w12058_
	);
	LUT2 #(
		.INIT('h8)
	) name10158 (
		\s15_data_i[24]_pad ,
		_w2062_,
		_w12059_
	);
	LUT4 #(
		.INIT('h135f)
	) name10159 (
		\s1_data_i[24]_pad ,
		\s8_data_i[24]_pad ,
		_w9302_,
		_w9360_,
		_w12060_
	);
	LUT4 #(
		.INIT('h153f)
	) name10160 (
		\s4_data_i[24]_pad ,
		\s6_data_i[24]_pad ,
		_w9363_,
		_w9366_,
		_w12061_
	);
	LUT4 #(
		.INIT('h153f)
	) name10161 (
		\s3_data_i[24]_pad ,
		\s9_data_i[24]_pad ,
		_w9357_,
		_w9523_,
		_w12062_
	);
	LUT4 #(
		.INIT('h135f)
	) name10162 (
		\s10_data_i[24]_pad ,
		\s7_data_i[24]_pad ,
		_w9509_,
		_w9529_,
		_w12063_
	);
	LUT4 #(
		.INIT('h8000)
	) name10163 (
		_w12060_,
		_w12061_,
		_w12062_,
		_w12063_,
		_w12064_
	);
	LUT2 #(
		.INIT('h8)
	) name10164 (
		\s11_data_i[24]_pad ,
		_w9372_,
		_w12065_
	);
	LUT4 #(
		.INIT('h135f)
	) name10165 (
		\s14_data_i[24]_pad ,
		\s2_data_i[24]_pad ,
		_w9515_,
		_w9520_,
		_w12066_
	);
	LUT4 #(
		.INIT('h135f)
	) name10166 (
		\s12_data_i[24]_pad ,
		\s5_data_i[24]_pad ,
		_w9512_,
		_w9526_,
		_w12067_
	);
	LUT4 #(
		.INIT('h135f)
	) name10167 (
		\s0_data_i[24]_pad ,
		\s13_data_i[24]_pad ,
		_w9298_,
		_w9369_,
		_w12068_
	);
	LUT4 #(
		.INIT('h4000)
	) name10168 (
		_w12065_,
		_w12066_,
		_w12067_,
		_w12068_,
		_w12069_
	);
	LUT2 #(
		.INIT('h8)
	) name10169 (
		_w12064_,
		_w12069_,
		_w12070_
	);
	LUT4 #(
		.INIT('h70ff)
	) name10170 (
		_w2046_,
		_w2097_,
		_w12059_,
		_w12070_,
		_w12071_
	);
	LUT2 #(
		.INIT('h8)
	) name10171 (
		\s15_data_i[25]_pad ,
		_w2062_,
		_w12072_
	);
	LUT4 #(
		.INIT('h135f)
	) name10172 (
		\s1_data_i[25]_pad ,
		\s8_data_i[25]_pad ,
		_w9302_,
		_w9360_,
		_w12073_
	);
	LUT4 #(
		.INIT('h153f)
	) name10173 (
		\s4_data_i[25]_pad ,
		\s6_data_i[25]_pad ,
		_w9363_,
		_w9366_,
		_w12074_
	);
	LUT4 #(
		.INIT('h153f)
	) name10174 (
		\s3_data_i[25]_pad ,
		\s9_data_i[25]_pad ,
		_w9357_,
		_w9523_,
		_w12075_
	);
	LUT4 #(
		.INIT('h135f)
	) name10175 (
		\s10_data_i[25]_pad ,
		\s7_data_i[25]_pad ,
		_w9509_,
		_w9529_,
		_w12076_
	);
	LUT4 #(
		.INIT('h8000)
	) name10176 (
		_w12073_,
		_w12074_,
		_w12075_,
		_w12076_,
		_w12077_
	);
	LUT2 #(
		.INIT('h8)
	) name10177 (
		\s11_data_i[25]_pad ,
		_w9372_,
		_w12078_
	);
	LUT4 #(
		.INIT('h135f)
	) name10178 (
		\s14_data_i[25]_pad ,
		\s2_data_i[25]_pad ,
		_w9515_,
		_w9520_,
		_w12079_
	);
	LUT4 #(
		.INIT('h135f)
	) name10179 (
		\s12_data_i[25]_pad ,
		\s5_data_i[25]_pad ,
		_w9512_,
		_w9526_,
		_w12080_
	);
	LUT4 #(
		.INIT('h135f)
	) name10180 (
		\s0_data_i[25]_pad ,
		\s13_data_i[25]_pad ,
		_w9298_,
		_w9369_,
		_w12081_
	);
	LUT4 #(
		.INIT('h4000)
	) name10181 (
		_w12078_,
		_w12079_,
		_w12080_,
		_w12081_,
		_w12082_
	);
	LUT2 #(
		.INIT('h8)
	) name10182 (
		_w12077_,
		_w12082_,
		_w12083_
	);
	LUT4 #(
		.INIT('h70ff)
	) name10183 (
		_w2046_,
		_w2097_,
		_w12072_,
		_w12083_,
		_w12084_
	);
	LUT2 #(
		.INIT('h8)
	) name10184 (
		\s15_data_i[26]_pad ,
		_w2062_,
		_w12085_
	);
	LUT4 #(
		.INIT('h135f)
	) name10185 (
		\s1_data_i[26]_pad ,
		\s8_data_i[26]_pad ,
		_w9302_,
		_w9360_,
		_w12086_
	);
	LUT4 #(
		.INIT('h153f)
	) name10186 (
		\s4_data_i[26]_pad ,
		\s6_data_i[26]_pad ,
		_w9363_,
		_w9366_,
		_w12087_
	);
	LUT4 #(
		.INIT('h153f)
	) name10187 (
		\s3_data_i[26]_pad ,
		\s9_data_i[26]_pad ,
		_w9357_,
		_w9523_,
		_w12088_
	);
	LUT4 #(
		.INIT('h135f)
	) name10188 (
		\s10_data_i[26]_pad ,
		\s7_data_i[26]_pad ,
		_w9509_,
		_w9529_,
		_w12089_
	);
	LUT4 #(
		.INIT('h8000)
	) name10189 (
		_w12086_,
		_w12087_,
		_w12088_,
		_w12089_,
		_w12090_
	);
	LUT2 #(
		.INIT('h8)
	) name10190 (
		\s11_data_i[26]_pad ,
		_w9372_,
		_w12091_
	);
	LUT4 #(
		.INIT('h135f)
	) name10191 (
		\s14_data_i[26]_pad ,
		\s2_data_i[26]_pad ,
		_w9515_,
		_w9520_,
		_w12092_
	);
	LUT4 #(
		.INIT('h135f)
	) name10192 (
		\s12_data_i[26]_pad ,
		\s5_data_i[26]_pad ,
		_w9512_,
		_w9526_,
		_w12093_
	);
	LUT4 #(
		.INIT('h135f)
	) name10193 (
		\s0_data_i[26]_pad ,
		\s13_data_i[26]_pad ,
		_w9298_,
		_w9369_,
		_w12094_
	);
	LUT4 #(
		.INIT('h4000)
	) name10194 (
		_w12091_,
		_w12092_,
		_w12093_,
		_w12094_,
		_w12095_
	);
	LUT2 #(
		.INIT('h8)
	) name10195 (
		_w12090_,
		_w12095_,
		_w12096_
	);
	LUT4 #(
		.INIT('h70ff)
	) name10196 (
		_w2046_,
		_w2097_,
		_w12085_,
		_w12096_,
		_w12097_
	);
	LUT2 #(
		.INIT('h8)
	) name10197 (
		\s15_data_i[27]_pad ,
		_w2062_,
		_w12098_
	);
	LUT4 #(
		.INIT('h135f)
	) name10198 (
		\s1_data_i[27]_pad ,
		\s8_data_i[27]_pad ,
		_w9302_,
		_w9360_,
		_w12099_
	);
	LUT4 #(
		.INIT('h153f)
	) name10199 (
		\s4_data_i[27]_pad ,
		\s6_data_i[27]_pad ,
		_w9363_,
		_w9366_,
		_w12100_
	);
	LUT4 #(
		.INIT('h153f)
	) name10200 (
		\s3_data_i[27]_pad ,
		\s9_data_i[27]_pad ,
		_w9357_,
		_w9523_,
		_w12101_
	);
	LUT4 #(
		.INIT('h135f)
	) name10201 (
		\s10_data_i[27]_pad ,
		\s7_data_i[27]_pad ,
		_w9509_,
		_w9529_,
		_w12102_
	);
	LUT4 #(
		.INIT('h8000)
	) name10202 (
		_w12099_,
		_w12100_,
		_w12101_,
		_w12102_,
		_w12103_
	);
	LUT2 #(
		.INIT('h8)
	) name10203 (
		\s11_data_i[27]_pad ,
		_w9372_,
		_w12104_
	);
	LUT4 #(
		.INIT('h135f)
	) name10204 (
		\s14_data_i[27]_pad ,
		\s2_data_i[27]_pad ,
		_w9515_,
		_w9520_,
		_w12105_
	);
	LUT4 #(
		.INIT('h135f)
	) name10205 (
		\s12_data_i[27]_pad ,
		\s5_data_i[27]_pad ,
		_w9512_,
		_w9526_,
		_w12106_
	);
	LUT4 #(
		.INIT('h135f)
	) name10206 (
		\s0_data_i[27]_pad ,
		\s13_data_i[27]_pad ,
		_w9298_,
		_w9369_,
		_w12107_
	);
	LUT4 #(
		.INIT('h4000)
	) name10207 (
		_w12104_,
		_w12105_,
		_w12106_,
		_w12107_,
		_w12108_
	);
	LUT2 #(
		.INIT('h8)
	) name10208 (
		_w12103_,
		_w12108_,
		_w12109_
	);
	LUT4 #(
		.INIT('h70ff)
	) name10209 (
		_w2046_,
		_w2097_,
		_w12098_,
		_w12109_,
		_w12110_
	);
	LUT2 #(
		.INIT('h8)
	) name10210 (
		\s15_data_i[28]_pad ,
		_w2062_,
		_w12111_
	);
	LUT4 #(
		.INIT('h135f)
	) name10211 (
		\s1_data_i[28]_pad ,
		\s8_data_i[28]_pad ,
		_w9302_,
		_w9360_,
		_w12112_
	);
	LUT4 #(
		.INIT('h153f)
	) name10212 (
		\s4_data_i[28]_pad ,
		\s6_data_i[28]_pad ,
		_w9363_,
		_w9366_,
		_w12113_
	);
	LUT4 #(
		.INIT('h153f)
	) name10213 (
		\s3_data_i[28]_pad ,
		\s9_data_i[28]_pad ,
		_w9357_,
		_w9523_,
		_w12114_
	);
	LUT4 #(
		.INIT('h135f)
	) name10214 (
		\s10_data_i[28]_pad ,
		\s7_data_i[28]_pad ,
		_w9509_,
		_w9529_,
		_w12115_
	);
	LUT4 #(
		.INIT('h8000)
	) name10215 (
		_w12112_,
		_w12113_,
		_w12114_,
		_w12115_,
		_w12116_
	);
	LUT2 #(
		.INIT('h8)
	) name10216 (
		\s11_data_i[28]_pad ,
		_w9372_,
		_w12117_
	);
	LUT4 #(
		.INIT('h135f)
	) name10217 (
		\s14_data_i[28]_pad ,
		\s2_data_i[28]_pad ,
		_w9515_,
		_w9520_,
		_w12118_
	);
	LUT4 #(
		.INIT('h135f)
	) name10218 (
		\s12_data_i[28]_pad ,
		\s5_data_i[28]_pad ,
		_w9512_,
		_w9526_,
		_w12119_
	);
	LUT4 #(
		.INIT('h135f)
	) name10219 (
		\s0_data_i[28]_pad ,
		\s13_data_i[28]_pad ,
		_w9298_,
		_w9369_,
		_w12120_
	);
	LUT4 #(
		.INIT('h4000)
	) name10220 (
		_w12117_,
		_w12118_,
		_w12119_,
		_w12120_,
		_w12121_
	);
	LUT2 #(
		.INIT('h8)
	) name10221 (
		_w12116_,
		_w12121_,
		_w12122_
	);
	LUT4 #(
		.INIT('h70ff)
	) name10222 (
		_w2046_,
		_w2097_,
		_w12111_,
		_w12122_,
		_w12123_
	);
	LUT2 #(
		.INIT('h8)
	) name10223 (
		\s15_data_i[29]_pad ,
		_w2062_,
		_w12124_
	);
	LUT4 #(
		.INIT('h135f)
	) name10224 (
		\s1_data_i[29]_pad ,
		\s8_data_i[29]_pad ,
		_w9302_,
		_w9360_,
		_w12125_
	);
	LUT4 #(
		.INIT('h153f)
	) name10225 (
		\s4_data_i[29]_pad ,
		\s6_data_i[29]_pad ,
		_w9363_,
		_w9366_,
		_w12126_
	);
	LUT4 #(
		.INIT('h153f)
	) name10226 (
		\s3_data_i[29]_pad ,
		\s9_data_i[29]_pad ,
		_w9357_,
		_w9523_,
		_w12127_
	);
	LUT4 #(
		.INIT('h135f)
	) name10227 (
		\s10_data_i[29]_pad ,
		\s7_data_i[29]_pad ,
		_w9509_,
		_w9529_,
		_w12128_
	);
	LUT4 #(
		.INIT('h8000)
	) name10228 (
		_w12125_,
		_w12126_,
		_w12127_,
		_w12128_,
		_w12129_
	);
	LUT2 #(
		.INIT('h8)
	) name10229 (
		\s11_data_i[29]_pad ,
		_w9372_,
		_w12130_
	);
	LUT4 #(
		.INIT('h135f)
	) name10230 (
		\s14_data_i[29]_pad ,
		\s2_data_i[29]_pad ,
		_w9515_,
		_w9520_,
		_w12131_
	);
	LUT4 #(
		.INIT('h135f)
	) name10231 (
		\s12_data_i[29]_pad ,
		\s5_data_i[29]_pad ,
		_w9512_,
		_w9526_,
		_w12132_
	);
	LUT4 #(
		.INIT('h135f)
	) name10232 (
		\s0_data_i[29]_pad ,
		\s13_data_i[29]_pad ,
		_w9298_,
		_w9369_,
		_w12133_
	);
	LUT4 #(
		.INIT('h4000)
	) name10233 (
		_w12130_,
		_w12131_,
		_w12132_,
		_w12133_,
		_w12134_
	);
	LUT2 #(
		.INIT('h8)
	) name10234 (
		_w12129_,
		_w12134_,
		_w12135_
	);
	LUT4 #(
		.INIT('h70ff)
	) name10235 (
		_w2046_,
		_w2097_,
		_w12124_,
		_w12135_,
		_w12136_
	);
	LUT3 #(
		.INIT('h80)
	) name10236 (
		_w2062_,
		_w2097_,
		_w9993_,
		_w12137_
	);
	LUT2 #(
		.INIT('h8)
	) name10237 (
		\s15_data_i[2]_pad ,
		_w2062_,
		_w12138_
	);
	LUT3 #(
		.INIT('h70)
	) name10238 (
		_w2046_,
		_w2097_,
		_w12138_,
		_w12139_
	);
	LUT4 #(
		.INIT('h135f)
	) name10239 (
		\s1_data_i[2]_pad ,
		\s8_data_i[2]_pad ,
		_w9302_,
		_w9360_,
		_w12140_
	);
	LUT4 #(
		.INIT('h153f)
	) name10240 (
		\s4_data_i[2]_pad ,
		\s6_data_i[2]_pad ,
		_w9363_,
		_w9366_,
		_w12141_
	);
	LUT4 #(
		.INIT('h153f)
	) name10241 (
		\s3_data_i[2]_pad ,
		\s9_data_i[2]_pad ,
		_w9357_,
		_w9523_,
		_w12142_
	);
	LUT4 #(
		.INIT('h135f)
	) name10242 (
		\s10_data_i[2]_pad ,
		\s7_data_i[2]_pad ,
		_w9509_,
		_w9529_,
		_w12143_
	);
	LUT4 #(
		.INIT('h8000)
	) name10243 (
		_w12140_,
		_w12141_,
		_w12142_,
		_w12143_,
		_w12144_
	);
	LUT2 #(
		.INIT('h8)
	) name10244 (
		\s11_data_i[2]_pad ,
		_w9372_,
		_w12145_
	);
	LUT4 #(
		.INIT('h135f)
	) name10245 (
		\s14_data_i[2]_pad ,
		\s2_data_i[2]_pad ,
		_w9515_,
		_w9520_,
		_w12146_
	);
	LUT4 #(
		.INIT('h135f)
	) name10246 (
		\s12_data_i[2]_pad ,
		\s5_data_i[2]_pad ,
		_w9512_,
		_w9526_,
		_w12147_
	);
	LUT4 #(
		.INIT('h135f)
	) name10247 (
		\s0_data_i[2]_pad ,
		\s13_data_i[2]_pad ,
		_w9298_,
		_w9369_,
		_w12148_
	);
	LUT4 #(
		.INIT('h4000)
	) name10248 (
		_w12145_,
		_w12146_,
		_w12147_,
		_w12148_,
		_w12149_
	);
	LUT2 #(
		.INIT('h8)
	) name10249 (
		_w12144_,
		_w12149_,
		_w12150_
	);
	LUT3 #(
		.INIT('hef)
	) name10250 (
		_w12137_,
		_w12139_,
		_w12150_,
		_w12151_
	);
	LUT2 #(
		.INIT('h8)
	) name10251 (
		\s15_data_i[30]_pad ,
		_w2062_,
		_w12152_
	);
	LUT4 #(
		.INIT('h135f)
	) name10252 (
		\s1_data_i[30]_pad ,
		\s8_data_i[30]_pad ,
		_w9302_,
		_w9360_,
		_w12153_
	);
	LUT4 #(
		.INIT('h153f)
	) name10253 (
		\s4_data_i[30]_pad ,
		\s6_data_i[30]_pad ,
		_w9363_,
		_w9366_,
		_w12154_
	);
	LUT4 #(
		.INIT('h153f)
	) name10254 (
		\s3_data_i[30]_pad ,
		\s9_data_i[30]_pad ,
		_w9357_,
		_w9523_,
		_w12155_
	);
	LUT4 #(
		.INIT('h135f)
	) name10255 (
		\s10_data_i[30]_pad ,
		\s7_data_i[30]_pad ,
		_w9509_,
		_w9529_,
		_w12156_
	);
	LUT4 #(
		.INIT('h8000)
	) name10256 (
		_w12153_,
		_w12154_,
		_w12155_,
		_w12156_,
		_w12157_
	);
	LUT2 #(
		.INIT('h8)
	) name10257 (
		\s11_data_i[30]_pad ,
		_w9372_,
		_w12158_
	);
	LUT4 #(
		.INIT('h135f)
	) name10258 (
		\s14_data_i[30]_pad ,
		\s2_data_i[30]_pad ,
		_w9515_,
		_w9520_,
		_w12159_
	);
	LUT4 #(
		.INIT('h135f)
	) name10259 (
		\s12_data_i[30]_pad ,
		\s5_data_i[30]_pad ,
		_w9512_,
		_w9526_,
		_w12160_
	);
	LUT4 #(
		.INIT('h135f)
	) name10260 (
		\s0_data_i[30]_pad ,
		\s13_data_i[30]_pad ,
		_w9298_,
		_w9369_,
		_w12161_
	);
	LUT4 #(
		.INIT('h4000)
	) name10261 (
		_w12158_,
		_w12159_,
		_w12160_,
		_w12161_,
		_w12162_
	);
	LUT2 #(
		.INIT('h8)
	) name10262 (
		_w12157_,
		_w12162_,
		_w12163_
	);
	LUT4 #(
		.INIT('h70ff)
	) name10263 (
		_w2046_,
		_w2097_,
		_w12152_,
		_w12163_,
		_w12164_
	);
	LUT2 #(
		.INIT('h8)
	) name10264 (
		\s15_data_i[31]_pad ,
		_w2062_,
		_w12165_
	);
	LUT4 #(
		.INIT('h135f)
	) name10265 (
		\s1_data_i[31]_pad ,
		\s8_data_i[31]_pad ,
		_w9302_,
		_w9360_,
		_w12166_
	);
	LUT4 #(
		.INIT('h153f)
	) name10266 (
		\s4_data_i[31]_pad ,
		\s6_data_i[31]_pad ,
		_w9363_,
		_w9366_,
		_w12167_
	);
	LUT4 #(
		.INIT('h153f)
	) name10267 (
		\s3_data_i[31]_pad ,
		\s9_data_i[31]_pad ,
		_w9357_,
		_w9523_,
		_w12168_
	);
	LUT4 #(
		.INIT('h135f)
	) name10268 (
		\s10_data_i[31]_pad ,
		\s7_data_i[31]_pad ,
		_w9509_,
		_w9529_,
		_w12169_
	);
	LUT4 #(
		.INIT('h8000)
	) name10269 (
		_w12166_,
		_w12167_,
		_w12168_,
		_w12169_,
		_w12170_
	);
	LUT2 #(
		.INIT('h8)
	) name10270 (
		\s11_data_i[31]_pad ,
		_w9372_,
		_w12171_
	);
	LUT4 #(
		.INIT('h135f)
	) name10271 (
		\s14_data_i[31]_pad ,
		\s2_data_i[31]_pad ,
		_w9515_,
		_w9520_,
		_w12172_
	);
	LUT4 #(
		.INIT('h135f)
	) name10272 (
		\s12_data_i[31]_pad ,
		\s5_data_i[31]_pad ,
		_w9512_,
		_w9526_,
		_w12173_
	);
	LUT4 #(
		.INIT('h135f)
	) name10273 (
		\s0_data_i[31]_pad ,
		\s13_data_i[31]_pad ,
		_w9298_,
		_w9369_,
		_w12174_
	);
	LUT4 #(
		.INIT('h4000)
	) name10274 (
		_w12171_,
		_w12172_,
		_w12173_,
		_w12174_,
		_w12175_
	);
	LUT2 #(
		.INIT('h8)
	) name10275 (
		_w12170_,
		_w12175_,
		_w12176_
	);
	LUT4 #(
		.INIT('h70ff)
	) name10276 (
		_w2046_,
		_w2097_,
		_w12165_,
		_w12176_,
		_w12177_
	);
	LUT3 #(
		.INIT('h80)
	) name10277 (
		_w2062_,
		_w2097_,
		_w10035_,
		_w12178_
	);
	LUT2 #(
		.INIT('h8)
	) name10278 (
		\s15_data_i[3]_pad ,
		_w2062_,
		_w12179_
	);
	LUT3 #(
		.INIT('h70)
	) name10279 (
		_w2046_,
		_w2097_,
		_w12179_,
		_w12180_
	);
	LUT4 #(
		.INIT('h135f)
	) name10280 (
		\s1_data_i[3]_pad ,
		\s8_data_i[3]_pad ,
		_w9302_,
		_w9360_,
		_w12181_
	);
	LUT4 #(
		.INIT('h153f)
	) name10281 (
		\s4_data_i[3]_pad ,
		\s6_data_i[3]_pad ,
		_w9363_,
		_w9366_,
		_w12182_
	);
	LUT4 #(
		.INIT('h153f)
	) name10282 (
		\s3_data_i[3]_pad ,
		\s9_data_i[3]_pad ,
		_w9357_,
		_w9523_,
		_w12183_
	);
	LUT4 #(
		.INIT('h135f)
	) name10283 (
		\s10_data_i[3]_pad ,
		\s7_data_i[3]_pad ,
		_w9509_,
		_w9529_,
		_w12184_
	);
	LUT4 #(
		.INIT('h8000)
	) name10284 (
		_w12181_,
		_w12182_,
		_w12183_,
		_w12184_,
		_w12185_
	);
	LUT2 #(
		.INIT('h8)
	) name10285 (
		\s11_data_i[3]_pad ,
		_w9372_,
		_w12186_
	);
	LUT4 #(
		.INIT('h135f)
	) name10286 (
		\s14_data_i[3]_pad ,
		\s2_data_i[3]_pad ,
		_w9515_,
		_w9520_,
		_w12187_
	);
	LUT4 #(
		.INIT('h135f)
	) name10287 (
		\s12_data_i[3]_pad ,
		\s5_data_i[3]_pad ,
		_w9512_,
		_w9526_,
		_w12188_
	);
	LUT4 #(
		.INIT('h135f)
	) name10288 (
		\s0_data_i[3]_pad ,
		\s13_data_i[3]_pad ,
		_w9298_,
		_w9369_,
		_w12189_
	);
	LUT4 #(
		.INIT('h4000)
	) name10289 (
		_w12186_,
		_w12187_,
		_w12188_,
		_w12189_,
		_w12190_
	);
	LUT2 #(
		.INIT('h8)
	) name10290 (
		_w12185_,
		_w12190_,
		_w12191_
	);
	LUT3 #(
		.INIT('hef)
	) name10291 (
		_w12178_,
		_w12180_,
		_w12191_,
		_w12192_
	);
	LUT3 #(
		.INIT('h80)
	) name10292 (
		_w2062_,
		_w2097_,
		_w10051_,
		_w12193_
	);
	LUT2 #(
		.INIT('h8)
	) name10293 (
		\s15_data_i[4]_pad ,
		_w2062_,
		_w12194_
	);
	LUT3 #(
		.INIT('h70)
	) name10294 (
		_w2046_,
		_w2097_,
		_w12194_,
		_w12195_
	);
	LUT4 #(
		.INIT('h135f)
	) name10295 (
		\s1_data_i[4]_pad ,
		\s8_data_i[4]_pad ,
		_w9302_,
		_w9360_,
		_w12196_
	);
	LUT4 #(
		.INIT('h153f)
	) name10296 (
		\s4_data_i[4]_pad ,
		\s6_data_i[4]_pad ,
		_w9363_,
		_w9366_,
		_w12197_
	);
	LUT4 #(
		.INIT('h153f)
	) name10297 (
		\s3_data_i[4]_pad ,
		\s9_data_i[4]_pad ,
		_w9357_,
		_w9523_,
		_w12198_
	);
	LUT4 #(
		.INIT('h135f)
	) name10298 (
		\s10_data_i[4]_pad ,
		\s7_data_i[4]_pad ,
		_w9509_,
		_w9529_,
		_w12199_
	);
	LUT4 #(
		.INIT('h8000)
	) name10299 (
		_w12196_,
		_w12197_,
		_w12198_,
		_w12199_,
		_w12200_
	);
	LUT2 #(
		.INIT('h8)
	) name10300 (
		\s11_data_i[4]_pad ,
		_w9372_,
		_w12201_
	);
	LUT4 #(
		.INIT('h135f)
	) name10301 (
		\s14_data_i[4]_pad ,
		\s2_data_i[4]_pad ,
		_w9515_,
		_w9520_,
		_w12202_
	);
	LUT4 #(
		.INIT('h135f)
	) name10302 (
		\s12_data_i[4]_pad ,
		\s5_data_i[4]_pad ,
		_w9512_,
		_w9526_,
		_w12203_
	);
	LUT4 #(
		.INIT('h135f)
	) name10303 (
		\s0_data_i[4]_pad ,
		\s13_data_i[4]_pad ,
		_w9298_,
		_w9369_,
		_w12204_
	);
	LUT4 #(
		.INIT('h4000)
	) name10304 (
		_w12201_,
		_w12202_,
		_w12203_,
		_w12204_,
		_w12205_
	);
	LUT2 #(
		.INIT('h8)
	) name10305 (
		_w12200_,
		_w12205_,
		_w12206_
	);
	LUT3 #(
		.INIT('hef)
	) name10306 (
		_w12193_,
		_w12195_,
		_w12206_,
		_w12207_
	);
	LUT3 #(
		.INIT('h80)
	) name10307 (
		_w2062_,
		_w2097_,
		_w10067_,
		_w12208_
	);
	LUT2 #(
		.INIT('h8)
	) name10308 (
		\s15_data_i[5]_pad ,
		_w2062_,
		_w12209_
	);
	LUT3 #(
		.INIT('h70)
	) name10309 (
		_w2046_,
		_w2097_,
		_w12209_,
		_w12210_
	);
	LUT4 #(
		.INIT('h135f)
	) name10310 (
		\s1_data_i[5]_pad ,
		\s8_data_i[5]_pad ,
		_w9302_,
		_w9360_,
		_w12211_
	);
	LUT4 #(
		.INIT('h153f)
	) name10311 (
		\s4_data_i[5]_pad ,
		\s6_data_i[5]_pad ,
		_w9363_,
		_w9366_,
		_w12212_
	);
	LUT4 #(
		.INIT('h153f)
	) name10312 (
		\s3_data_i[5]_pad ,
		\s9_data_i[5]_pad ,
		_w9357_,
		_w9523_,
		_w12213_
	);
	LUT4 #(
		.INIT('h135f)
	) name10313 (
		\s10_data_i[5]_pad ,
		\s7_data_i[5]_pad ,
		_w9509_,
		_w9529_,
		_w12214_
	);
	LUT4 #(
		.INIT('h8000)
	) name10314 (
		_w12211_,
		_w12212_,
		_w12213_,
		_w12214_,
		_w12215_
	);
	LUT2 #(
		.INIT('h8)
	) name10315 (
		\s11_data_i[5]_pad ,
		_w9372_,
		_w12216_
	);
	LUT4 #(
		.INIT('h135f)
	) name10316 (
		\s14_data_i[5]_pad ,
		\s2_data_i[5]_pad ,
		_w9515_,
		_w9520_,
		_w12217_
	);
	LUT4 #(
		.INIT('h135f)
	) name10317 (
		\s12_data_i[5]_pad ,
		\s5_data_i[5]_pad ,
		_w9512_,
		_w9526_,
		_w12218_
	);
	LUT4 #(
		.INIT('h135f)
	) name10318 (
		\s0_data_i[5]_pad ,
		\s13_data_i[5]_pad ,
		_w9298_,
		_w9369_,
		_w12219_
	);
	LUT4 #(
		.INIT('h4000)
	) name10319 (
		_w12216_,
		_w12217_,
		_w12218_,
		_w12219_,
		_w12220_
	);
	LUT2 #(
		.INIT('h8)
	) name10320 (
		_w12215_,
		_w12220_,
		_w12221_
	);
	LUT3 #(
		.INIT('hef)
	) name10321 (
		_w12208_,
		_w12210_,
		_w12221_,
		_w12222_
	);
	LUT3 #(
		.INIT('h80)
	) name10322 (
		_w2062_,
		_w2097_,
		_w10083_,
		_w12223_
	);
	LUT2 #(
		.INIT('h8)
	) name10323 (
		\s15_data_i[6]_pad ,
		_w2062_,
		_w12224_
	);
	LUT3 #(
		.INIT('h70)
	) name10324 (
		_w2046_,
		_w2097_,
		_w12224_,
		_w12225_
	);
	LUT4 #(
		.INIT('h153f)
	) name10325 (
		\s11_data_i[6]_pad ,
		\s1_data_i[6]_pad ,
		_w9302_,
		_w9372_,
		_w12226_
	);
	LUT4 #(
		.INIT('h153f)
	) name10326 (
		\s4_data_i[6]_pad ,
		\s6_data_i[6]_pad ,
		_w9363_,
		_w9366_,
		_w12227_
	);
	LUT4 #(
		.INIT('h153f)
	) name10327 (
		\s5_data_i[6]_pad ,
		\s9_data_i[6]_pad ,
		_w9357_,
		_w9526_,
		_w12228_
	);
	LUT4 #(
		.INIT('h135f)
	) name10328 (
		\s10_data_i[6]_pad ,
		\s7_data_i[6]_pad ,
		_w9509_,
		_w9529_,
		_w12229_
	);
	LUT4 #(
		.INIT('h8000)
	) name10329 (
		_w12226_,
		_w12227_,
		_w12228_,
		_w12229_,
		_w12230_
	);
	LUT2 #(
		.INIT('h8)
	) name10330 (
		\s12_data_i[6]_pad ,
		_w9512_,
		_w12231_
	);
	LUT4 #(
		.INIT('h135f)
	) name10331 (
		\s2_data_i[6]_pad ,
		\s3_data_i[6]_pad ,
		_w9520_,
		_w9523_,
		_w12232_
	);
	LUT4 #(
		.INIT('h153f)
	) name10332 (
		\s14_data_i[6]_pad ,
		\s8_data_i[6]_pad ,
		_w9360_,
		_w9515_,
		_w12233_
	);
	LUT4 #(
		.INIT('h135f)
	) name10333 (
		\s0_data_i[6]_pad ,
		\s13_data_i[6]_pad ,
		_w9298_,
		_w9369_,
		_w12234_
	);
	LUT4 #(
		.INIT('h4000)
	) name10334 (
		_w12231_,
		_w12232_,
		_w12233_,
		_w12234_,
		_w12235_
	);
	LUT2 #(
		.INIT('h8)
	) name10335 (
		_w12230_,
		_w12235_,
		_w12236_
	);
	LUT3 #(
		.INIT('hef)
	) name10336 (
		_w12223_,
		_w12225_,
		_w12236_,
		_w12237_
	);
	LUT3 #(
		.INIT('h80)
	) name10337 (
		_w2062_,
		_w2097_,
		_w10099_,
		_w12238_
	);
	LUT2 #(
		.INIT('h8)
	) name10338 (
		\s15_data_i[7]_pad ,
		_w2062_,
		_w12239_
	);
	LUT3 #(
		.INIT('h70)
	) name10339 (
		_w2046_,
		_w2097_,
		_w12239_,
		_w12240_
	);
	LUT4 #(
		.INIT('h135f)
	) name10340 (
		\s1_data_i[7]_pad ,
		\s8_data_i[7]_pad ,
		_w9302_,
		_w9360_,
		_w12241_
	);
	LUT4 #(
		.INIT('h153f)
	) name10341 (
		\s4_data_i[7]_pad ,
		\s6_data_i[7]_pad ,
		_w9363_,
		_w9366_,
		_w12242_
	);
	LUT4 #(
		.INIT('h153f)
	) name10342 (
		\s3_data_i[7]_pad ,
		\s9_data_i[7]_pad ,
		_w9357_,
		_w9523_,
		_w12243_
	);
	LUT4 #(
		.INIT('h135f)
	) name10343 (
		\s10_data_i[7]_pad ,
		\s7_data_i[7]_pad ,
		_w9509_,
		_w9529_,
		_w12244_
	);
	LUT4 #(
		.INIT('h8000)
	) name10344 (
		_w12241_,
		_w12242_,
		_w12243_,
		_w12244_,
		_w12245_
	);
	LUT2 #(
		.INIT('h8)
	) name10345 (
		\s11_data_i[7]_pad ,
		_w9372_,
		_w12246_
	);
	LUT4 #(
		.INIT('h135f)
	) name10346 (
		\s14_data_i[7]_pad ,
		\s2_data_i[7]_pad ,
		_w9515_,
		_w9520_,
		_w12247_
	);
	LUT4 #(
		.INIT('h135f)
	) name10347 (
		\s12_data_i[7]_pad ,
		\s5_data_i[7]_pad ,
		_w9512_,
		_w9526_,
		_w12248_
	);
	LUT4 #(
		.INIT('h135f)
	) name10348 (
		\s0_data_i[7]_pad ,
		\s13_data_i[7]_pad ,
		_w9298_,
		_w9369_,
		_w12249_
	);
	LUT4 #(
		.INIT('h4000)
	) name10349 (
		_w12246_,
		_w12247_,
		_w12248_,
		_w12249_,
		_w12250_
	);
	LUT2 #(
		.INIT('h8)
	) name10350 (
		_w12245_,
		_w12250_,
		_w12251_
	);
	LUT3 #(
		.INIT('hef)
	) name10351 (
		_w12238_,
		_w12240_,
		_w12251_,
		_w12252_
	);
	LUT3 #(
		.INIT('h80)
	) name10352 (
		_w2062_,
		_w2097_,
		_w10115_,
		_w12253_
	);
	LUT2 #(
		.INIT('h8)
	) name10353 (
		\s15_data_i[8]_pad ,
		_w2062_,
		_w12254_
	);
	LUT3 #(
		.INIT('h70)
	) name10354 (
		_w2046_,
		_w2097_,
		_w12254_,
		_w12255_
	);
	LUT4 #(
		.INIT('h135f)
	) name10355 (
		\s1_data_i[8]_pad ,
		\s8_data_i[8]_pad ,
		_w9302_,
		_w9360_,
		_w12256_
	);
	LUT4 #(
		.INIT('h153f)
	) name10356 (
		\s4_data_i[8]_pad ,
		\s6_data_i[8]_pad ,
		_w9363_,
		_w9366_,
		_w12257_
	);
	LUT4 #(
		.INIT('h153f)
	) name10357 (
		\s3_data_i[8]_pad ,
		\s9_data_i[8]_pad ,
		_w9357_,
		_w9523_,
		_w12258_
	);
	LUT4 #(
		.INIT('h135f)
	) name10358 (
		\s10_data_i[8]_pad ,
		\s7_data_i[8]_pad ,
		_w9509_,
		_w9529_,
		_w12259_
	);
	LUT4 #(
		.INIT('h8000)
	) name10359 (
		_w12256_,
		_w12257_,
		_w12258_,
		_w12259_,
		_w12260_
	);
	LUT2 #(
		.INIT('h8)
	) name10360 (
		\s11_data_i[8]_pad ,
		_w9372_,
		_w12261_
	);
	LUT4 #(
		.INIT('h135f)
	) name10361 (
		\s14_data_i[8]_pad ,
		\s2_data_i[8]_pad ,
		_w9515_,
		_w9520_,
		_w12262_
	);
	LUT4 #(
		.INIT('h135f)
	) name10362 (
		\s12_data_i[8]_pad ,
		\s5_data_i[8]_pad ,
		_w9512_,
		_w9526_,
		_w12263_
	);
	LUT4 #(
		.INIT('h135f)
	) name10363 (
		\s0_data_i[8]_pad ,
		\s13_data_i[8]_pad ,
		_w9298_,
		_w9369_,
		_w12264_
	);
	LUT4 #(
		.INIT('h4000)
	) name10364 (
		_w12261_,
		_w12262_,
		_w12263_,
		_w12264_,
		_w12265_
	);
	LUT2 #(
		.INIT('h8)
	) name10365 (
		_w12260_,
		_w12265_,
		_w12266_
	);
	LUT3 #(
		.INIT('hef)
	) name10366 (
		_w12253_,
		_w12255_,
		_w12266_,
		_w12267_
	);
	LUT3 #(
		.INIT('h80)
	) name10367 (
		_w2062_,
		_w2097_,
		_w10131_,
		_w12268_
	);
	LUT2 #(
		.INIT('h8)
	) name10368 (
		\s15_data_i[9]_pad ,
		_w2062_,
		_w12269_
	);
	LUT3 #(
		.INIT('h70)
	) name10369 (
		_w2046_,
		_w2097_,
		_w12269_,
		_w12270_
	);
	LUT4 #(
		.INIT('h135f)
	) name10370 (
		\s1_data_i[9]_pad ,
		\s8_data_i[9]_pad ,
		_w9302_,
		_w9360_,
		_w12271_
	);
	LUT4 #(
		.INIT('h153f)
	) name10371 (
		\s4_data_i[9]_pad ,
		\s6_data_i[9]_pad ,
		_w9363_,
		_w9366_,
		_w12272_
	);
	LUT4 #(
		.INIT('h153f)
	) name10372 (
		\s3_data_i[9]_pad ,
		\s9_data_i[9]_pad ,
		_w9357_,
		_w9523_,
		_w12273_
	);
	LUT4 #(
		.INIT('h135f)
	) name10373 (
		\s10_data_i[9]_pad ,
		\s7_data_i[9]_pad ,
		_w9509_,
		_w9529_,
		_w12274_
	);
	LUT4 #(
		.INIT('h8000)
	) name10374 (
		_w12271_,
		_w12272_,
		_w12273_,
		_w12274_,
		_w12275_
	);
	LUT2 #(
		.INIT('h8)
	) name10375 (
		\s11_data_i[9]_pad ,
		_w9372_,
		_w12276_
	);
	LUT4 #(
		.INIT('h135f)
	) name10376 (
		\s14_data_i[9]_pad ,
		\s2_data_i[9]_pad ,
		_w9515_,
		_w9520_,
		_w12277_
	);
	LUT4 #(
		.INIT('h135f)
	) name10377 (
		\s12_data_i[9]_pad ,
		\s5_data_i[9]_pad ,
		_w9512_,
		_w9526_,
		_w12278_
	);
	LUT4 #(
		.INIT('h135f)
	) name10378 (
		\s0_data_i[9]_pad ,
		\s13_data_i[9]_pad ,
		_w9298_,
		_w9369_,
		_w12279_
	);
	LUT4 #(
		.INIT('h4000)
	) name10379 (
		_w12276_,
		_w12277_,
		_w12278_,
		_w12279_,
		_w12280_
	);
	LUT2 #(
		.INIT('h8)
	) name10380 (
		_w12275_,
		_w12280_,
		_w12281_
	);
	LUT3 #(
		.INIT('hef)
	) name10381 (
		_w12268_,
		_w12270_,
		_w12281_,
		_w12282_
	);
	LUT3 #(
		.INIT('h80)
	) name10382 (
		\s15_err_i_pad ,
		_w1907_,
		_w11805_,
		_w12283_
	);
	LUT4 #(
		.INIT('h8000)
	) name10383 (
		\s6_err_i_pad ,
		_w8743_,
		_w8744_,
		_w9363_,
		_w12284_
	);
	LUT4 #(
		.INIT('h8000)
	) name10384 (
		\s1_err_i_pad ,
		_w9103_,
		_w9104_,
		_w9302_,
		_w12285_
	);
	LUT4 #(
		.INIT('h135f)
	) name10385 (
		_w8762_,
		_w9116_,
		_w12284_,
		_w12285_,
		_w12286_
	);
	LUT4 #(
		.INIT('h8000)
	) name10386 (
		\s7_err_i_pad ,
		_w8782_,
		_w8783_,
		_w9529_,
		_w12287_
	);
	LUT4 #(
		.INIT('h8000)
	) name10387 (
		\s3_err_i_pad ,
		_w9205_,
		_w9206_,
		_w9523_,
		_w12288_
	);
	LUT4 #(
		.INIT('h135f)
	) name10388 (
		_w8801_,
		_w9204_,
		_w12287_,
		_w12288_,
		_w12289_
	);
	LUT4 #(
		.INIT('h8000)
	) name10389 (
		\s14_err_i_pad ,
		_w9137_,
		_w9138_,
		_w9515_,
		_w12290_
	);
	LUT4 #(
		.INIT('h8000)
	) name10390 (
		\s13_err_i_pad ,
		_w9069_,
		_w9070_,
		_w9369_,
		_w12291_
	);
	LUT4 #(
		.INIT('h153f)
	) name10391 (
		_w9088_,
		_w9156_,
		_w12290_,
		_w12291_,
		_w12292_
	);
	LUT4 #(
		.INIT('h8000)
	) name10392 (
		\s10_err_i_pad ,
		_w8910_,
		_w8911_,
		_w9509_,
		_w12293_
	);
	LUT4 #(
		.INIT('h8000)
	) name10393 (
		\s9_err_i_pad ,
		_w8865_,
		_w8866_,
		_w9357_,
		_w12294_
	);
	LUT4 #(
		.INIT('h153f)
	) name10394 (
		_w8884_,
		_w8929_,
		_w12293_,
		_w12294_,
		_w12295_
	);
	LUT4 #(
		.INIT('h8000)
	) name10395 (
		_w12286_,
		_w12289_,
		_w12292_,
		_w12295_,
		_w12296_
	);
	LUT4 #(
		.INIT('h8000)
	) name10396 (
		\s0_err_i_pad ,
		_w8989_,
		_w8990_,
		_w9298_,
		_w12297_
	);
	LUT2 #(
		.INIT('h8)
	) name10397 (
		_w8996_,
		_w12297_,
		_w12298_
	);
	LUT4 #(
		.INIT('h8000)
	) name10398 (
		\s11_err_i_pad ,
		_w8955_,
		_w8956_,
		_w9372_,
		_w12299_
	);
	LUT4 #(
		.INIT('h8000)
	) name10399 (
		\s5_err_i_pad ,
		_w8699_,
		_w8700_,
		_w9526_,
		_w12300_
	);
	LUT4 #(
		.INIT('h153f)
	) name10400 (
		_w8706_,
		_w8954_,
		_w12299_,
		_w12300_,
		_w12301_
	);
	LUT4 #(
		.INIT('h8000)
	) name10401 (
		\s12_err_i_pad ,
		_w9029_,
		_w9030_,
		_w9512_,
		_w12302_
	);
	LUT4 #(
		.INIT('h8000)
	) name10402 (
		\s4_err_i_pad ,
		_w8655_,
		_w8656_,
		_w9366_,
		_w12303_
	);
	LUT4 #(
		.INIT('h153f)
	) name10403 (
		_w8654_,
		_w9042_,
		_w12302_,
		_w12303_,
		_w12304_
	);
	LUT4 #(
		.INIT('h8000)
	) name10404 (
		\s2_err_i_pad ,
		_w9171_,
		_w9172_,
		_w9520_,
		_w12305_
	);
	LUT4 #(
		.INIT('h8000)
	) name10405 (
		\s8_err_i_pad ,
		_w8821_,
		_w8822_,
		_w9360_,
		_w12306_
	);
	LUT4 #(
		.INIT('h153f)
	) name10406 (
		_w8840_,
		_w9170_,
		_w12305_,
		_w12306_,
		_w12307_
	);
	LUT4 #(
		.INIT('h4000)
	) name10407 (
		_w12298_,
		_w12301_,
		_w12304_,
		_w12307_,
		_w12308_
	);
	LUT2 #(
		.INIT('h8)
	) name10408 (
		_w12296_,
		_w12308_,
		_w12309_
	);
	LUT4 #(
		.INIT('h70ff)
	) name10409 (
		_w2046_,
		_w2097_,
		_w12283_,
		_w12309_,
		_w12310_
	);
	LUT3 #(
		.INIT('h80)
	) name10410 (
		\s15_rty_i_pad ,
		_w1907_,
		_w11805_,
		_w12311_
	);
	LUT4 #(
		.INIT('h8000)
	) name10411 (
		\s14_rty_i_pad ,
		_w9137_,
		_w9138_,
		_w9515_,
		_w12312_
	);
	LUT4 #(
		.INIT('h8000)
	) name10412 (
		\s1_rty_i_pad ,
		_w9103_,
		_w9104_,
		_w9302_,
		_w12313_
	);
	LUT4 #(
		.INIT('h153f)
	) name10413 (
		_w9116_,
		_w9156_,
		_w12312_,
		_w12313_,
		_w12314_
	);
	LUT4 #(
		.INIT('h8000)
	) name10414 (
		\s10_rty_i_pad ,
		_w8910_,
		_w8911_,
		_w9509_,
		_w12315_
	);
	LUT4 #(
		.INIT('h8000)
	) name10415 (
		\s7_rty_i_pad ,
		_w8782_,
		_w8783_,
		_w9529_,
		_w12316_
	);
	LUT4 #(
		.INIT('h153f)
	) name10416 (
		_w8801_,
		_w8929_,
		_w12315_,
		_w12316_,
		_w12317_
	);
	LUT4 #(
		.INIT('h8000)
	) name10417 (
		\s8_rty_i_pad ,
		_w8821_,
		_w8822_,
		_w9360_,
		_w12318_
	);
	LUT4 #(
		.INIT('h8000)
	) name10418 (
		\s9_rty_i_pad ,
		_w8865_,
		_w8866_,
		_w9357_,
		_w12319_
	);
	LUT4 #(
		.INIT('h135f)
	) name10419 (
		_w8840_,
		_w8884_,
		_w12318_,
		_w12319_,
		_w12320_
	);
	LUT4 #(
		.INIT('h8000)
	) name10420 (
		\s6_rty_i_pad ,
		_w8743_,
		_w8744_,
		_w9363_,
		_w12321_
	);
	LUT4 #(
		.INIT('h8000)
	) name10421 (
		\s13_rty_i_pad ,
		_w9069_,
		_w9070_,
		_w9369_,
		_w12322_
	);
	LUT4 #(
		.INIT('h135f)
	) name10422 (
		_w8762_,
		_w9088_,
		_w12321_,
		_w12322_,
		_w12323_
	);
	LUT4 #(
		.INIT('h8000)
	) name10423 (
		_w12314_,
		_w12317_,
		_w12320_,
		_w12323_,
		_w12324_
	);
	LUT4 #(
		.INIT('h8000)
	) name10424 (
		\s12_rty_i_pad ,
		_w9029_,
		_w9030_,
		_w9512_,
		_w12325_
	);
	LUT2 #(
		.INIT('h8)
	) name10425 (
		_w9042_,
		_w12325_,
		_w12326_
	);
	LUT4 #(
		.INIT('h8000)
	) name10426 (
		\s5_rty_i_pad ,
		_w8699_,
		_w8700_,
		_w9526_,
		_w12327_
	);
	LUT4 #(
		.INIT('h8000)
	) name10427 (
		\s4_rty_i_pad ,
		_w8655_,
		_w8656_,
		_w9366_,
		_w12328_
	);
	LUT4 #(
		.INIT('h153f)
	) name10428 (
		_w8654_,
		_w8706_,
		_w12327_,
		_w12328_,
		_w12329_
	);
	LUT4 #(
		.INIT('h8000)
	) name10429 (
		\s0_rty_i_pad ,
		_w8989_,
		_w8990_,
		_w9298_,
		_w12330_
	);
	LUT4 #(
		.INIT('h8000)
	) name10430 (
		\s11_rty_i_pad ,
		_w8955_,
		_w8956_,
		_w9372_,
		_w12331_
	);
	LUT4 #(
		.INIT('h153f)
	) name10431 (
		_w8954_,
		_w8996_,
		_w12330_,
		_w12331_,
		_w12332_
	);
	LUT4 #(
		.INIT('h8000)
	) name10432 (
		\s2_rty_i_pad ,
		_w9171_,
		_w9172_,
		_w9520_,
		_w12333_
	);
	LUT4 #(
		.INIT('h8000)
	) name10433 (
		\s3_rty_i_pad ,
		_w9205_,
		_w9206_,
		_w9523_,
		_w12334_
	);
	LUT4 #(
		.INIT('h135f)
	) name10434 (
		_w9170_,
		_w9204_,
		_w12333_,
		_w12334_,
		_w12335_
	);
	LUT4 #(
		.INIT('h4000)
	) name10435 (
		_w12326_,
		_w12329_,
		_w12332_,
		_w12335_,
		_w12336_
	);
	LUT2 #(
		.INIT('h8)
	) name10436 (
		_w12324_,
		_w12336_,
		_w12337_
	);
	LUT4 #(
		.INIT('h70ff)
	) name10437 (
		_w2046_,
		_w2097_,
		_w12311_,
		_w12337_,
		_w12338_
	);
	LUT3 #(
		.INIT('h70)
	) name10438 (
		_w1901_,
		_w1902_,
		_w2064_,
		_w12339_
	);
	LUT2 #(
		.INIT('h8)
	) name10439 (
		_w1920_,
		_w12339_,
		_w12340_
	);
	LUT3 #(
		.INIT('h70)
	) name10440 (
		_w2097_,
		_w8630_,
		_w12340_,
		_w12341_
	);
	LUT4 #(
		.INIT('h2a00)
	) name10441 (
		\s11_ack_i_pad ,
		_w8955_,
		_w8956_,
		_w9535_,
		_w12342_
	);
	LUT4 #(
		.INIT('h2a00)
	) name10442 (
		\s3_ack_i_pad ,
		_w9205_,
		_w9206_,
		_w9351_,
		_w12343_
	);
	LUT4 #(
		.INIT('h135f)
	) name10443 (
		_w8954_,
		_w9204_,
		_w12342_,
		_w12343_,
		_w12344_
	);
	LUT4 #(
		.INIT('h2a00)
	) name10444 (
		\s1_ack_i_pad ,
		_w9103_,
		_w9104_,
		_w9269_,
		_w12345_
	);
	LUT4 #(
		.INIT('h2a00)
	) name10445 (
		\s7_ack_i_pad ,
		_w8782_,
		_w8783_,
		_w9345_,
		_w12346_
	);
	LUT4 #(
		.INIT('h153f)
	) name10446 (
		_w8801_,
		_w9116_,
		_w12345_,
		_w12346_,
		_w12347_
	);
	LUT4 #(
		.INIT('h2a00)
	) name10447 (
		\s10_ack_i_pad ,
		_w8910_,
		_w8911_,
		_w9532_,
		_w12348_
	);
	LUT4 #(
		.INIT('h2a00)
	) name10448 (
		\s2_ack_i_pad ,
		_w9171_,
		_w9172_,
		_w9541_,
		_w12349_
	);
	LUT4 #(
		.INIT('h135f)
	) name10449 (
		_w8929_,
		_w9170_,
		_w12348_,
		_w12349_,
		_w12350_
	);
	LUT4 #(
		.INIT('h2a00)
	) name10450 (
		\s13_ack_i_pad ,
		_w9069_,
		_w9070_,
		_w9538_,
		_w12351_
	);
	LUT4 #(
		.INIT('h2a00)
	) name10451 (
		\s6_ack_i_pad ,
		_w8743_,
		_w8744_,
		_w9550_,
		_w12352_
	);
	LUT4 #(
		.INIT('h153f)
	) name10452 (
		_w8762_,
		_w9088_,
		_w12351_,
		_w12352_,
		_w12353_
	);
	LUT4 #(
		.INIT('h8000)
	) name10453 (
		_w12344_,
		_w12347_,
		_w12350_,
		_w12353_,
		_w12354_
	);
	LUT4 #(
		.INIT('h2a00)
	) name10454 (
		\s8_ack_i_pad ,
		_w8821_,
		_w8822_,
		_w9553_,
		_w12355_
	);
	LUT2 #(
		.INIT('h8)
	) name10455 (
		_w8840_,
		_w12355_,
		_w12356_
	);
	LUT4 #(
		.INIT('h2a00)
	) name10456 (
		\s14_ack_i_pad ,
		_w9137_,
		_w9138_,
		_w9348_,
		_w12357_
	);
	LUT4 #(
		.INIT('h2a00)
	) name10457 (
		\s9_ack_i_pad ,
		_w8865_,
		_w8866_,
		_w9556_,
		_w12358_
	);
	LUT4 #(
		.INIT('h153f)
	) name10458 (
		_w8884_,
		_w9156_,
		_w12357_,
		_w12358_,
		_w12359_
	);
	LUT4 #(
		.INIT('h2a00)
	) name10459 (
		\s4_ack_i_pad ,
		_w8655_,
		_w8656_,
		_w9544_,
		_w12360_
	);
	LUT4 #(
		.INIT('h2a00)
	) name10460 (
		\s0_ack_i_pad ,
		_w8989_,
		_w8990_,
		_w9305_,
		_w12361_
	);
	LUT4 #(
		.INIT('h135f)
	) name10461 (
		_w8654_,
		_w8996_,
		_w12360_,
		_w12361_,
		_w12362_
	);
	LUT4 #(
		.INIT('h2a00)
	) name10462 (
		\s5_ack_i_pad ,
		_w8699_,
		_w8700_,
		_w9547_,
		_w12363_
	);
	LUT4 #(
		.INIT('h2a00)
	) name10463 (
		\s12_ack_i_pad ,
		_w9029_,
		_w9030_,
		_w9354_,
		_w12364_
	);
	LUT4 #(
		.INIT('h135f)
	) name10464 (
		_w8706_,
		_w9042_,
		_w12363_,
		_w12364_,
		_w12365_
	);
	LUT4 #(
		.INIT('h4000)
	) name10465 (
		_w12356_,
		_w12359_,
		_w12362_,
		_w12365_,
		_w12366_
	);
	LUT2 #(
		.INIT('h8)
	) name10466 (
		_w12354_,
		_w12366_,
		_w12367_
	);
	LUT3 #(
		.INIT('h4f)
	) name10467 (
		_w9652_,
		_w12341_,
		_w12367_,
		_w12368_
	);
	LUT3 #(
		.INIT('h80)
	) name10468 (
		_w2064_,
		_w2097_,
		_w9683_,
		_w12369_
	);
	LUT2 #(
		.INIT('h8)
	) name10469 (
		\s15_data_i[0]_pad ,
		_w2064_,
		_w12370_
	);
	LUT3 #(
		.INIT('h70)
	) name10470 (
		_w2046_,
		_w2097_,
		_w12370_,
		_w12371_
	);
	LUT4 #(
		.INIT('h153f)
	) name10471 (
		\s12_data_i[0]_pad ,
		\s1_data_i[0]_pad ,
		_w9269_,
		_w9354_,
		_w12372_
	);
	LUT4 #(
		.INIT('h135f)
	) name10472 (
		\s0_data_i[0]_pad ,
		\s10_data_i[0]_pad ,
		_w9305_,
		_w9532_,
		_w12373_
	);
	LUT4 #(
		.INIT('h135f)
	) name10473 (
		\s3_data_i[0]_pad ,
		\s4_data_i[0]_pad ,
		_w9351_,
		_w9544_,
		_w12374_
	);
	LUT4 #(
		.INIT('h135f)
	) name10474 (
		\s6_data_i[0]_pad ,
		\s9_data_i[0]_pad ,
		_w9550_,
		_w9556_,
		_w12375_
	);
	LUT4 #(
		.INIT('h8000)
	) name10475 (
		_w12372_,
		_w12373_,
		_w12374_,
		_w12375_,
		_w12376_
	);
	LUT2 #(
		.INIT('h8)
	) name10476 (
		\s14_data_i[0]_pad ,
		_w9348_,
		_w12377_
	);
	LUT4 #(
		.INIT('h153f)
	) name10477 (
		\s11_data_i[0]_pad ,
		\s7_data_i[0]_pad ,
		_w9345_,
		_w9535_,
		_w12378_
	);
	LUT4 #(
		.INIT('h135f)
	) name10478 (
		\s5_data_i[0]_pad ,
		\s8_data_i[0]_pad ,
		_w9547_,
		_w9553_,
		_w12379_
	);
	LUT4 #(
		.INIT('h135f)
	) name10479 (
		\s13_data_i[0]_pad ,
		\s2_data_i[0]_pad ,
		_w9538_,
		_w9541_,
		_w12380_
	);
	LUT4 #(
		.INIT('h4000)
	) name10480 (
		_w12377_,
		_w12378_,
		_w12379_,
		_w12380_,
		_w12381_
	);
	LUT2 #(
		.INIT('h8)
	) name10481 (
		_w12376_,
		_w12381_,
		_w12382_
	);
	LUT3 #(
		.INIT('hef)
	) name10482 (
		_w12369_,
		_w12371_,
		_w12382_,
		_w12383_
	);
	LUT3 #(
		.INIT('h80)
	) name10483 (
		_w2064_,
		_w2097_,
		_w9699_,
		_w12384_
	);
	LUT2 #(
		.INIT('h8)
	) name10484 (
		\s15_data_i[10]_pad ,
		_w2064_,
		_w12385_
	);
	LUT3 #(
		.INIT('h70)
	) name10485 (
		_w2046_,
		_w2097_,
		_w12385_,
		_w12386_
	);
	LUT4 #(
		.INIT('h153f)
	) name10486 (
		\s12_data_i[10]_pad ,
		\s1_data_i[10]_pad ,
		_w9269_,
		_w9354_,
		_w12387_
	);
	LUT4 #(
		.INIT('h135f)
	) name10487 (
		\s0_data_i[10]_pad ,
		\s10_data_i[10]_pad ,
		_w9305_,
		_w9532_,
		_w12388_
	);
	LUT4 #(
		.INIT('h135f)
	) name10488 (
		\s3_data_i[10]_pad ,
		\s4_data_i[10]_pad ,
		_w9351_,
		_w9544_,
		_w12389_
	);
	LUT4 #(
		.INIT('h135f)
	) name10489 (
		\s6_data_i[10]_pad ,
		\s9_data_i[10]_pad ,
		_w9550_,
		_w9556_,
		_w12390_
	);
	LUT4 #(
		.INIT('h8000)
	) name10490 (
		_w12387_,
		_w12388_,
		_w12389_,
		_w12390_,
		_w12391_
	);
	LUT2 #(
		.INIT('h8)
	) name10491 (
		\s14_data_i[10]_pad ,
		_w9348_,
		_w12392_
	);
	LUT4 #(
		.INIT('h153f)
	) name10492 (
		\s11_data_i[10]_pad ,
		\s7_data_i[10]_pad ,
		_w9345_,
		_w9535_,
		_w12393_
	);
	LUT4 #(
		.INIT('h135f)
	) name10493 (
		\s5_data_i[10]_pad ,
		\s8_data_i[10]_pad ,
		_w9547_,
		_w9553_,
		_w12394_
	);
	LUT4 #(
		.INIT('h135f)
	) name10494 (
		\s13_data_i[10]_pad ,
		\s2_data_i[10]_pad ,
		_w9538_,
		_w9541_,
		_w12395_
	);
	LUT4 #(
		.INIT('h4000)
	) name10495 (
		_w12392_,
		_w12393_,
		_w12394_,
		_w12395_,
		_w12396_
	);
	LUT2 #(
		.INIT('h8)
	) name10496 (
		_w12391_,
		_w12396_,
		_w12397_
	);
	LUT3 #(
		.INIT('hef)
	) name10497 (
		_w12384_,
		_w12386_,
		_w12397_,
		_w12398_
	);
	LUT3 #(
		.INIT('h80)
	) name10498 (
		_w2064_,
		_w2097_,
		_w9715_,
		_w12399_
	);
	LUT2 #(
		.INIT('h8)
	) name10499 (
		\s15_data_i[11]_pad ,
		_w2064_,
		_w12400_
	);
	LUT3 #(
		.INIT('h70)
	) name10500 (
		_w2046_,
		_w2097_,
		_w12400_,
		_w12401_
	);
	LUT4 #(
		.INIT('h135f)
	) name10501 (
		\s1_data_i[11]_pad ,
		\s7_data_i[11]_pad ,
		_w9269_,
		_w9345_,
		_w12402_
	);
	LUT4 #(
		.INIT('h135f)
	) name10502 (
		\s2_data_i[11]_pad ,
		\s5_data_i[11]_pad ,
		_w9541_,
		_w9547_,
		_w12403_
	);
	LUT4 #(
		.INIT('h153f)
	) name10503 (
		\s12_data_i[11]_pad ,
		\s3_data_i[11]_pad ,
		_w9351_,
		_w9354_,
		_w12404_
	);
	LUT4 #(
		.INIT('h135f)
	) name10504 (
		\s14_data_i[11]_pad ,
		\s8_data_i[11]_pad ,
		_w9348_,
		_w9553_,
		_w12405_
	);
	LUT4 #(
		.INIT('h8000)
	) name10505 (
		_w12402_,
		_w12403_,
		_w12404_,
		_w12405_,
		_w12406_
	);
	LUT2 #(
		.INIT('h8)
	) name10506 (
		\s0_data_i[11]_pad ,
		_w9305_,
		_w12407_
	);
	LUT4 #(
		.INIT('h135f)
	) name10507 (
		\s11_data_i[11]_pad ,
		\s13_data_i[11]_pad ,
		_w9535_,
		_w9538_,
		_w12408_
	);
	LUT4 #(
		.INIT('h135f)
	) name10508 (
		\s4_data_i[11]_pad ,
		\s6_data_i[11]_pad ,
		_w9544_,
		_w9550_,
		_w12409_
	);
	LUT4 #(
		.INIT('h135f)
	) name10509 (
		\s10_data_i[11]_pad ,
		\s9_data_i[11]_pad ,
		_w9532_,
		_w9556_,
		_w12410_
	);
	LUT4 #(
		.INIT('h4000)
	) name10510 (
		_w12407_,
		_w12408_,
		_w12409_,
		_w12410_,
		_w12411_
	);
	LUT2 #(
		.INIT('h8)
	) name10511 (
		_w12406_,
		_w12411_,
		_w12412_
	);
	LUT3 #(
		.INIT('hef)
	) name10512 (
		_w12399_,
		_w12401_,
		_w12412_,
		_w12413_
	);
	LUT3 #(
		.INIT('h80)
	) name10513 (
		_w2064_,
		_w2097_,
		_w9731_,
		_w12414_
	);
	LUT2 #(
		.INIT('h8)
	) name10514 (
		\s15_data_i[12]_pad ,
		_w2064_,
		_w12415_
	);
	LUT3 #(
		.INIT('h70)
	) name10515 (
		_w2046_,
		_w2097_,
		_w12415_,
		_w12416_
	);
	LUT4 #(
		.INIT('h153f)
	) name10516 (
		\s12_data_i[12]_pad ,
		\s1_data_i[12]_pad ,
		_w9269_,
		_w9354_,
		_w12417_
	);
	LUT4 #(
		.INIT('h135f)
	) name10517 (
		\s0_data_i[12]_pad ,
		\s10_data_i[12]_pad ,
		_w9305_,
		_w9532_,
		_w12418_
	);
	LUT4 #(
		.INIT('h135f)
	) name10518 (
		\s3_data_i[12]_pad ,
		\s4_data_i[12]_pad ,
		_w9351_,
		_w9544_,
		_w12419_
	);
	LUT4 #(
		.INIT('h135f)
	) name10519 (
		\s6_data_i[12]_pad ,
		\s9_data_i[12]_pad ,
		_w9550_,
		_w9556_,
		_w12420_
	);
	LUT4 #(
		.INIT('h8000)
	) name10520 (
		_w12417_,
		_w12418_,
		_w12419_,
		_w12420_,
		_w12421_
	);
	LUT2 #(
		.INIT('h8)
	) name10521 (
		\s14_data_i[12]_pad ,
		_w9348_,
		_w12422_
	);
	LUT4 #(
		.INIT('h153f)
	) name10522 (
		\s11_data_i[12]_pad ,
		\s7_data_i[12]_pad ,
		_w9345_,
		_w9535_,
		_w12423_
	);
	LUT4 #(
		.INIT('h135f)
	) name10523 (
		\s5_data_i[12]_pad ,
		\s8_data_i[12]_pad ,
		_w9547_,
		_w9553_,
		_w12424_
	);
	LUT4 #(
		.INIT('h135f)
	) name10524 (
		\s13_data_i[12]_pad ,
		\s2_data_i[12]_pad ,
		_w9538_,
		_w9541_,
		_w12425_
	);
	LUT4 #(
		.INIT('h4000)
	) name10525 (
		_w12422_,
		_w12423_,
		_w12424_,
		_w12425_,
		_w12426_
	);
	LUT2 #(
		.INIT('h8)
	) name10526 (
		_w12421_,
		_w12426_,
		_w12427_
	);
	LUT3 #(
		.INIT('hef)
	) name10527 (
		_w12414_,
		_w12416_,
		_w12427_,
		_w12428_
	);
	LUT3 #(
		.INIT('h80)
	) name10528 (
		_w2064_,
		_w2097_,
		_w9747_,
		_w12429_
	);
	LUT2 #(
		.INIT('h8)
	) name10529 (
		\s15_data_i[13]_pad ,
		_w2064_,
		_w12430_
	);
	LUT3 #(
		.INIT('h70)
	) name10530 (
		_w2046_,
		_w2097_,
		_w12430_,
		_w12431_
	);
	LUT4 #(
		.INIT('h153f)
	) name10531 (
		\s12_data_i[13]_pad ,
		\s1_data_i[13]_pad ,
		_w9269_,
		_w9354_,
		_w12432_
	);
	LUT4 #(
		.INIT('h135f)
	) name10532 (
		\s0_data_i[13]_pad ,
		\s10_data_i[13]_pad ,
		_w9305_,
		_w9532_,
		_w12433_
	);
	LUT4 #(
		.INIT('h135f)
	) name10533 (
		\s3_data_i[13]_pad ,
		\s4_data_i[13]_pad ,
		_w9351_,
		_w9544_,
		_w12434_
	);
	LUT4 #(
		.INIT('h135f)
	) name10534 (
		\s6_data_i[13]_pad ,
		\s9_data_i[13]_pad ,
		_w9550_,
		_w9556_,
		_w12435_
	);
	LUT4 #(
		.INIT('h8000)
	) name10535 (
		_w12432_,
		_w12433_,
		_w12434_,
		_w12435_,
		_w12436_
	);
	LUT2 #(
		.INIT('h8)
	) name10536 (
		\s14_data_i[13]_pad ,
		_w9348_,
		_w12437_
	);
	LUT4 #(
		.INIT('h153f)
	) name10537 (
		\s11_data_i[13]_pad ,
		\s7_data_i[13]_pad ,
		_w9345_,
		_w9535_,
		_w12438_
	);
	LUT4 #(
		.INIT('h135f)
	) name10538 (
		\s5_data_i[13]_pad ,
		\s8_data_i[13]_pad ,
		_w9547_,
		_w9553_,
		_w12439_
	);
	LUT4 #(
		.INIT('h135f)
	) name10539 (
		\s13_data_i[13]_pad ,
		\s2_data_i[13]_pad ,
		_w9538_,
		_w9541_,
		_w12440_
	);
	LUT4 #(
		.INIT('h4000)
	) name10540 (
		_w12437_,
		_w12438_,
		_w12439_,
		_w12440_,
		_w12441_
	);
	LUT2 #(
		.INIT('h8)
	) name10541 (
		_w12436_,
		_w12441_,
		_w12442_
	);
	LUT3 #(
		.INIT('hef)
	) name10542 (
		_w12429_,
		_w12431_,
		_w12442_,
		_w12443_
	);
	LUT3 #(
		.INIT('h80)
	) name10543 (
		_w2064_,
		_w2097_,
		_w9763_,
		_w12444_
	);
	LUT2 #(
		.INIT('h8)
	) name10544 (
		\s15_data_i[14]_pad ,
		_w2064_,
		_w12445_
	);
	LUT3 #(
		.INIT('h70)
	) name10545 (
		_w2046_,
		_w2097_,
		_w12445_,
		_w12446_
	);
	LUT4 #(
		.INIT('h153f)
	) name10546 (
		\s12_data_i[14]_pad ,
		\s1_data_i[14]_pad ,
		_w9269_,
		_w9354_,
		_w12447_
	);
	LUT4 #(
		.INIT('h135f)
	) name10547 (
		\s0_data_i[14]_pad ,
		\s10_data_i[14]_pad ,
		_w9305_,
		_w9532_,
		_w12448_
	);
	LUT4 #(
		.INIT('h135f)
	) name10548 (
		\s3_data_i[14]_pad ,
		\s4_data_i[14]_pad ,
		_w9351_,
		_w9544_,
		_w12449_
	);
	LUT4 #(
		.INIT('h135f)
	) name10549 (
		\s6_data_i[14]_pad ,
		\s9_data_i[14]_pad ,
		_w9550_,
		_w9556_,
		_w12450_
	);
	LUT4 #(
		.INIT('h8000)
	) name10550 (
		_w12447_,
		_w12448_,
		_w12449_,
		_w12450_,
		_w12451_
	);
	LUT2 #(
		.INIT('h8)
	) name10551 (
		\s14_data_i[14]_pad ,
		_w9348_,
		_w12452_
	);
	LUT4 #(
		.INIT('h153f)
	) name10552 (
		\s11_data_i[14]_pad ,
		\s7_data_i[14]_pad ,
		_w9345_,
		_w9535_,
		_w12453_
	);
	LUT4 #(
		.INIT('h135f)
	) name10553 (
		\s5_data_i[14]_pad ,
		\s8_data_i[14]_pad ,
		_w9547_,
		_w9553_,
		_w12454_
	);
	LUT4 #(
		.INIT('h135f)
	) name10554 (
		\s13_data_i[14]_pad ,
		\s2_data_i[14]_pad ,
		_w9538_,
		_w9541_,
		_w12455_
	);
	LUT4 #(
		.INIT('h4000)
	) name10555 (
		_w12452_,
		_w12453_,
		_w12454_,
		_w12455_,
		_w12456_
	);
	LUT2 #(
		.INIT('h8)
	) name10556 (
		_w12451_,
		_w12456_,
		_w12457_
	);
	LUT3 #(
		.INIT('hef)
	) name10557 (
		_w12444_,
		_w12446_,
		_w12457_,
		_w12458_
	);
	LUT3 #(
		.INIT('h80)
	) name10558 (
		_w2064_,
		_w2097_,
		_w9779_,
		_w12459_
	);
	LUT2 #(
		.INIT('h8)
	) name10559 (
		\s15_data_i[15]_pad ,
		_w2064_,
		_w12460_
	);
	LUT3 #(
		.INIT('h70)
	) name10560 (
		_w2046_,
		_w2097_,
		_w12460_,
		_w12461_
	);
	LUT4 #(
		.INIT('h153f)
	) name10561 (
		\s12_data_i[15]_pad ,
		\s1_data_i[15]_pad ,
		_w9269_,
		_w9354_,
		_w12462_
	);
	LUT4 #(
		.INIT('h135f)
	) name10562 (
		\s0_data_i[15]_pad ,
		\s10_data_i[15]_pad ,
		_w9305_,
		_w9532_,
		_w12463_
	);
	LUT4 #(
		.INIT('h135f)
	) name10563 (
		\s3_data_i[15]_pad ,
		\s4_data_i[15]_pad ,
		_w9351_,
		_w9544_,
		_w12464_
	);
	LUT4 #(
		.INIT('h135f)
	) name10564 (
		\s6_data_i[15]_pad ,
		\s9_data_i[15]_pad ,
		_w9550_,
		_w9556_,
		_w12465_
	);
	LUT4 #(
		.INIT('h8000)
	) name10565 (
		_w12462_,
		_w12463_,
		_w12464_,
		_w12465_,
		_w12466_
	);
	LUT2 #(
		.INIT('h8)
	) name10566 (
		\s14_data_i[15]_pad ,
		_w9348_,
		_w12467_
	);
	LUT4 #(
		.INIT('h153f)
	) name10567 (
		\s11_data_i[15]_pad ,
		\s7_data_i[15]_pad ,
		_w9345_,
		_w9535_,
		_w12468_
	);
	LUT4 #(
		.INIT('h135f)
	) name10568 (
		\s5_data_i[15]_pad ,
		\s8_data_i[15]_pad ,
		_w9547_,
		_w9553_,
		_w12469_
	);
	LUT4 #(
		.INIT('h135f)
	) name10569 (
		\s13_data_i[15]_pad ,
		\s2_data_i[15]_pad ,
		_w9538_,
		_w9541_,
		_w12470_
	);
	LUT4 #(
		.INIT('h4000)
	) name10570 (
		_w12467_,
		_w12468_,
		_w12469_,
		_w12470_,
		_w12471_
	);
	LUT2 #(
		.INIT('h8)
	) name10571 (
		_w12466_,
		_w12471_,
		_w12472_
	);
	LUT3 #(
		.INIT('hef)
	) name10572 (
		_w12459_,
		_w12461_,
		_w12472_,
		_w12473_
	);
	LUT2 #(
		.INIT('h8)
	) name10573 (
		\s15_data_i[16]_pad ,
		_w2064_,
		_w12474_
	);
	LUT4 #(
		.INIT('h135f)
	) name10574 (
		\s1_data_i[16]_pad ,
		\s8_data_i[16]_pad ,
		_w9269_,
		_w9553_,
		_w12475_
	);
	LUT4 #(
		.INIT('h135f)
	) name10575 (
		\s4_data_i[16]_pad ,
		\s6_data_i[16]_pad ,
		_w9544_,
		_w9550_,
		_w12476_
	);
	LUT4 #(
		.INIT('h135f)
	) name10576 (
		\s3_data_i[16]_pad ,
		\s9_data_i[16]_pad ,
		_w9351_,
		_w9556_,
		_w12477_
	);
	LUT4 #(
		.INIT('h153f)
	) name10577 (
		\s10_data_i[16]_pad ,
		\s7_data_i[16]_pad ,
		_w9345_,
		_w9532_,
		_w12478_
	);
	LUT4 #(
		.INIT('h8000)
	) name10578 (
		_w12475_,
		_w12476_,
		_w12477_,
		_w12478_,
		_w12479_
	);
	LUT2 #(
		.INIT('h8)
	) name10579 (
		\s11_data_i[16]_pad ,
		_w9535_,
		_w12480_
	);
	LUT4 #(
		.INIT('h135f)
	) name10580 (
		\s14_data_i[16]_pad ,
		\s2_data_i[16]_pad ,
		_w9348_,
		_w9541_,
		_w12481_
	);
	LUT4 #(
		.INIT('h135f)
	) name10581 (
		\s12_data_i[16]_pad ,
		\s5_data_i[16]_pad ,
		_w9354_,
		_w9547_,
		_w12482_
	);
	LUT4 #(
		.INIT('h135f)
	) name10582 (
		\s0_data_i[16]_pad ,
		\s13_data_i[16]_pad ,
		_w9305_,
		_w9538_,
		_w12483_
	);
	LUT4 #(
		.INIT('h4000)
	) name10583 (
		_w12480_,
		_w12481_,
		_w12482_,
		_w12483_,
		_w12484_
	);
	LUT2 #(
		.INIT('h8)
	) name10584 (
		_w12479_,
		_w12484_,
		_w12485_
	);
	LUT4 #(
		.INIT('h70ff)
	) name10585 (
		_w2046_,
		_w2097_,
		_w12474_,
		_w12485_,
		_w12486_
	);
	LUT2 #(
		.INIT('h8)
	) name10586 (
		\s15_data_i[17]_pad ,
		_w2064_,
		_w12487_
	);
	LUT4 #(
		.INIT('h135f)
	) name10587 (
		\s1_data_i[17]_pad ,
		\s8_data_i[17]_pad ,
		_w9269_,
		_w9553_,
		_w12488_
	);
	LUT4 #(
		.INIT('h135f)
	) name10588 (
		\s4_data_i[17]_pad ,
		\s6_data_i[17]_pad ,
		_w9544_,
		_w9550_,
		_w12489_
	);
	LUT4 #(
		.INIT('h135f)
	) name10589 (
		\s3_data_i[17]_pad ,
		\s9_data_i[17]_pad ,
		_w9351_,
		_w9556_,
		_w12490_
	);
	LUT4 #(
		.INIT('h153f)
	) name10590 (
		\s10_data_i[17]_pad ,
		\s7_data_i[17]_pad ,
		_w9345_,
		_w9532_,
		_w12491_
	);
	LUT4 #(
		.INIT('h8000)
	) name10591 (
		_w12488_,
		_w12489_,
		_w12490_,
		_w12491_,
		_w12492_
	);
	LUT2 #(
		.INIT('h8)
	) name10592 (
		\s11_data_i[17]_pad ,
		_w9535_,
		_w12493_
	);
	LUT4 #(
		.INIT('h135f)
	) name10593 (
		\s14_data_i[17]_pad ,
		\s2_data_i[17]_pad ,
		_w9348_,
		_w9541_,
		_w12494_
	);
	LUT4 #(
		.INIT('h135f)
	) name10594 (
		\s12_data_i[17]_pad ,
		\s5_data_i[17]_pad ,
		_w9354_,
		_w9547_,
		_w12495_
	);
	LUT4 #(
		.INIT('h135f)
	) name10595 (
		\s0_data_i[17]_pad ,
		\s13_data_i[17]_pad ,
		_w9305_,
		_w9538_,
		_w12496_
	);
	LUT4 #(
		.INIT('h4000)
	) name10596 (
		_w12493_,
		_w12494_,
		_w12495_,
		_w12496_,
		_w12497_
	);
	LUT2 #(
		.INIT('h8)
	) name10597 (
		_w12492_,
		_w12497_,
		_w12498_
	);
	LUT4 #(
		.INIT('h70ff)
	) name10598 (
		_w2046_,
		_w2097_,
		_w12487_,
		_w12498_,
		_w12499_
	);
	LUT2 #(
		.INIT('h8)
	) name10599 (
		\s15_data_i[18]_pad ,
		_w2064_,
		_w12500_
	);
	LUT4 #(
		.INIT('h135f)
	) name10600 (
		\s1_data_i[18]_pad ,
		\s8_data_i[18]_pad ,
		_w9269_,
		_w9553_,
		_w12501_
	);
	LUT4 #(
		.INIT('h135f)
	) name10601 (
		\s4_data_i[18]_pad ,
		\s6_data_i[18]_pad ,
		_w9544_,
		_w9550_,
		_w12502_
	);
	LUT4 #(
		.INIT('h135f)
	) name10602 (
		\s3_data_i[18]_pad ,
		\s9_data_i[18]_pad ,
		_w9351_,
		_w9556_,
		_w12503_
	);
	LUT4 #(
		.INIT('h153f)
	) name10603 (
		\s10_data_i[18]_pad ,
		\s7_data_i[18]_pad ,
		_w9345_,
		_w9532_,
		_w12504_
	);
	LUT4 #(
		.INIT('h8000)
	) name10604 (
		_w12501_,
		_w12502_,
		_w12503_,
		_w12504_,
		_w12505_
	);
	LUT2 #(
		.INIT('h8)
	) name10605 (
		\s11_data_i[18]_pad ,
		_w9535_,
		_w12506_
	);
	LUT4 #(
		.INIT('h135f)
	) name10606 (
		\s14_data_i[18]_pad ,
		\s2_data_i[18]_pad ,
		_w9348_,
		_w9541_,
		_w12507_
	);
	LUT4 #(
		.INIT('h135f)
	) name10607 (
		\s12_data_i[18]_pad ,
		\s5_data_i[18]_pad ,
		_w9354_,
		_w9547_,
		_w12508_
	);
	LUT4 #(
		.INIT('h135f)
	) name10608 (
		\s0_data_i[18]_pad ,
		\s13_data_i[18]_pad ,
		_w9305_,
		_w9538_,
		_w12509_
	);
	LUT4 #(
		.INIT('h4000)
	) name10609 (
		_w12506_,
		_w12507_,
		_w12508_,
		_w12509_,
		_w12510_
	);
	LUT2 #(
		.INIT('h8)
	) name10610 (
		_w12505_,
		_w12510_,
		_w12511_
	);
	LUT4 #(
		.INIT('h70ff)
	) name10611 (
		_w2046_,
		_w2097_,
		_w12500_,
		_w12511_,
		_w12512_
	);
	LUT2 #(
		.INIT('h8)
	) name10612 (
		\s15_data_i[19]_pad ,
		_w2064_,
		_w12513_
	);
	LUT4 #(
		.INIT('h135f)
	) name10613 (
		\s1_data_i[19]_pad ,
		\s8_data_i[19]_pad ,
		_w9269_,
		_w9553_,
		_w12514_
	);
	LUT4 #(
		.INIT('h135f)
	) name10614 (
		\s4_data_i[19]_pad ,
		\s6_data_i[19]_pad ,
		_w9544_,
		_w9550_,
		_w12515_
	);
	LUT4 #(
		.INIT('h135f)
	) name10615 (
		\s3_data_i[19]_pad ,
		\s9_data_i[19]_pad ,
		_w9351_,
		_w9556_,
		_w12516_
	);
	LUT4 #(
		.INIT('h153f)
	) name10616 (
		\s10_data_i[19]_pad ,
		\s7_data_i[19]_pad ,
		_w9345_,
		_w9532_,
		_w12517_
	);
	LUT4 #(
		.INIT('h8000)
	) name10617 (
		_w12514_,
		_w12515_,
		_w12516_,
		_w12517_,
		_w12518_
	);
	LUT2 #(
		.INIT('h8)
	) name10618 (
		\s11_data_i[19]_pad ,
		_w9535_,
		_w12519_
	);
	LUT4 #(
		.INIT('h135f)
	) name10619 (
		\s14_data_i[19]_pad ,
		\s2_data_i[19]_pad ,
		_w9348_,
		_w9541_,
		_w12520_
	);
	LUT4 #(
		.INIT('h135f)
	) name10620 (
		\s12_data_i[19]_pad ,
		\s5_data_i[19]_pad ,
		_w9354_,
		_w9547_,
		_w12521_
	);
	LUT4 #(
		.INIT('h135f)
	) name10621 (
		\s0_data_i[19]_pad ,
		\s13_data_i[19]_pad ,
		_w9305_,
		_w9538_,
		_w12522_
	);
	LUT4 #(
		.INIT('h4000)
	) name10622 (
		_w12519_,
		_w12520_,
		_w12521_,
		_w12522_,
		_w12523_
	);
	LUT2 #(
		.INIT('h8)
	) name10623 (
		_w12518_,
		_w12523_,
		_w12524_
	);
	LUT4 #(
		.INIT('h70ff)
	) name10624 (
		_w2046_,
		_w2097_,
		_w12513_,
		_w12524_,
		_w12525_
	);
	LUT3 #(
		.INIT('h80)
	) name10625 (
		_w2064_,
		_w2097_,
		_w9847_,
		_w12526_
	);
	LUT2 #(
		.INIT('h8)
	) name10626 (
		\s15_data_i[1]_pad ,
		_w2064_,
		_w12527_
	);
	LUT3 #(
		.INIT('h70)
	) name10627 (
		_w2046_,
		_w2097_,
		_w12527_,
		_w12528_
	);
	LUT4 #(
		.INIT('h153f)
	) name10628 (
		\s12_data_i[1]_pad ,
		\s1_data_i[1]_pad ,
		_w9269_,
		_w9354_,
		_w12529_
	);
	LUT4 #(
		.INIT('h135f)
	) name10629 (
		\s0_data_i[1]_pad ,
		\s10_data_i[1]_pad ,
		_w9305_,
		_w9532_,
		_w12530_
	);
	LUT4 #(
		.INIT('h135f)
	) name10630 (
		\s3_data_i[1]_pad ,
		\s4_data_i[1]_pad ,
		_w9351_,
		_w9544_,
		_w12531_
	);
	LUT4 #(
		.INIT('h135f)
	) name10631 (
		\s6_data_i[1]_pad ,
		\s9_data_i[1]_pad ,
		_w9550_,
		_w9556_,
		_w12532_
	);
	LUT4 #(
		.INIT('h8000)
	) name10632 (
		_w12529_,
		_w12530_,
		_w12531_,
		_w12532_,
		_w12533_
	);
	LUT2 #(
		.INIT('h8)
	) name10633 (
		\s14_data_i[1]_pad ,
		_w9348_,
		_w12534_
	);
	LUT4 #(
		.INIT('h153f)
	) name10634 (
		\s11_data_i[1]_pad ,
		\s7_data_i[1]_pad ,
		_w9345_,
		_w9535_,
		_w12535_
	);
	LUT4 #(
		.INIT('h135f)
	) name10635 (
		\s5_data_i[1]_pad ,
		\s8_data_i[1]_pad ,
		_w9547_,
		_w9553_,
		_w12536_
	);
	LUT4 #(
		.INIT('h135f)
	) name10636 (
		\s13_data_i[1]_pad ,
		\s2_data_i[1]_pad ,
		_w9538_,
		_w9541_,
		_w12537_
	);
	LUT4 #(
		.INIT('h4000)
	) name10637 (
		_w12534_,
		_w12535_,
		_w12536_,
		_w12537_,
		_w12538_
	);
	LUT2 #(
		.INIT('h8)
	) name10638 (
		_w12533_,
		_w12538_,
		_w12539_
	);
	LUT3 #(
		.INIT('hef)
	) name10639 (
		_w12526_,
		_w12528_,
		_w12539_,
		_w12540_
	);
	LUT2 #(
		.INIT('h8)
	) name10640 (
		\s15_data_i[20]_pad ,
		_w2064_,
		_w12541_
	);
	LUT4 #(
		.INIT('h135f)
	) name10641 (
		\s1_data_i[20]_pad ,
		\s8_data_i[20]_pad ,
		_w9269_,
		_w9553_,
		_w12542_
	);
	LUT4 #(
		.INIT('h135f)
	) name10642 (
		\s4_data_i[20]_pad ,
		\s6_data_i[20]_pad ,
		_w9544_,
		_w9550_,
		_w12543_
	);
	LUT4 #(
		.INIT('h135f)
	) name10643 (
		\s3_data_i[20]_pad ,
		\s9_data_i[20]_pad ,
		_w9351_,
		_w9556_,
		_w12544_
	);
	LUT4 #(
		.INIT('h153f)
	) name10644 (
		\s10_data_i[20]_pad ,
		\s7_data_i[20]_pad ,
		_w9345_,
		_w9532_,
		_w12545_
	);
	LUT4 #(
		.INIT('h8000)
	) name10645 (
		_w12542_,
		_w12543_,
		_w12544_,
		_w12545_,
		_w12546_
	);
	LUT2 #(
		.INIT('h8)
	) name10646 (
		\s11_data_i[20]_pad ,
		_w9535_,
		_w12547_
	);
	LUT4 #(
		.INIT('h135f)
	) name10647 (
		\s14_data_i[20]_pad ,
		\s2_data_i[20]_pad ,
		_w9348_,
		_w9541_,
		_w12548_
	);
	LUT4 #(
		.INIT('h135f)
	) name10648 (
		\s12_data_i[20]_pad ,
		\s5_data_i[20]_pad ,
		_w9354_,
		_w9547_,
		_w12549_
	);
	LUT4 #(
		.INIT('h135f)
	) name10649 (
		\s0_data_i[20]_pad ,
		\s13_data_i[20]_pad ,
		_w9305_,
		_w9538_,
		_w12550_
	);
	LUT4 #(
		.INIT('h4000)
	) name10650 (
		_w12547_,
		_w12548_,
		_w12549_,
		_w12550_,
		_w12551_
	);
	LUT2 #(
		.INIT('h8)
	) name10651 (
		_w12546_,
		_w12551_,
		_w12552_
	);
	LUT4 #(
		.INIT('h70ff)
	) name10652 (
		_w2046_,
		_w2097_,
		_w12541_,
		_w12552_,
		_w12553_
	);
	LUT2 #(
		.INIT('h8)
	) name10653 (
		\s15_data_i[21]_pad ,
		_w2064_,
		_w12554_
	);
	LUT4 #(
		.INIT('h135f)
	) name10654 (
		\s1_data_i[21]_pad ,
		\s8_data_i[21]_pad ,
		_w9269_,
		_w9553_,
		_w12555_
	);
	LUT4 #(
		.INIT('h135f)
	) name10655 (
		\s4_data_i[21]_pad ,
		\s6_data_i[21]_pad ,
		_w9544_,
		_w9550_,
		_w12556_
	);
	LUT4 #(
		.INIT('h135f)
	) name10656 (
		\s3_data_i[21]_pad ,
		\s9_data_i[21]_pad ,
		_w9351_,
		_w9556_,
		_w12557_
	);
	LUT4 #(
		.INIT('h153f)
	) name10657 (
		\s10_data_i[21]_pad ,
		\s7_data_i[21]_pad ,
		_w9345_,
		_w9532_,
		_w12558_
	);
	LUT4 #(
		.INIT('h8000)
	) name10658 (
		_w12555_,
		_w12556_,
		_w12557_,
		_w12558_,
		_w12559_
	);
	LUT2 #(
		.INIT('h8)
	) name10659 (
		\s11_data_i[21]_pad ,
		_w9535_,
		_w12560_
	);
	LUT4 #(
		.INIT('h135f)
	) name10660 (
		\s14_data_i[21]_pad ,
		\s2_data_i[21]_pad ,
		_w9348_,
		_w9541_,
		_w12561_
	);
	LUT4 #(
		.INIT('h135f)
	) name10661 (
		\s12_data_i[21]_pad ,
		\s5_data_i[21]_pad ,
		_w9354_,
		_w9547_,
		_w12562_
	);
	LUT4 #(
		.INIT('h135f)
	) name10662 (
		\s0_data_i[21]_pad ,
		\s13_data_i[21]_pad ,
		_w9305_,
		_w9538_,
		_w12563_
	);
	LUT4 #(
		.INIT('h4000)
	) name10663 (
		_w12560_,
		_w12561_,
		_w12562_,
		_w12563_,
		_w12564_
	);
	LUT2 #(
		.INIT('h8)
	) name10664 (
		_w12559_,
		_w12564_,
		_w12565_
	);
	LUT4 #(
		.INIT('h70ff)
	) name10665 (
		_w2046_,
		_w2097_,
		_w12554_,
		_w12565_,
		_w12566_
	);
	LUT2 #(
		.INIT('h8)
	) name10666 (
		\s15_data_i[22]_pad ,
		_w2064_,
		_w12567_
	);
	LUT4 #(
		.INIT('h135f)
	) name10667 (
		\s1_data_i[22]_pad ,
		\s8_data_i[22]_pad ,
		_w9269_,
		_w9553_,
		_w12568_
	);
	LUT4 #(
		.INIT('h135f)
	) name10668 (
		\s4_data_i[22]_pad ,
		\s6_data_i[22]_pad ,
		_w9544_,
		_w9550_,
		_w12569_
	);
	LUT4 #(
		.INIT('h135f)
	) name10669 (
		\s3_data_i[22]_pad ,
		\s9_data_i[22]_pad ,
		_w9351_,
		_w9556_,
		_w12570_
	);
	LUT4 #(
		.INIT('h153f)
	) name10670 (
		\s10_data_i[22]_pad ,
		\s7_data_i[22]_pad ,
		_w9345_,
		_w9532_,
		_w12571_
	);
	LUT4 #(
		.INIT('h8000)
	) name10671 (
		_w12568_,
		_w12569_,
		_w12570_,
		_w12571_,
		_w12572_
	);
	LUT2 #(
		.INIT('h8)
	) name10672 (
		\s11_data_i[22]_pad ,
		_w9535_,
		_w12573_
	);
	LUT4 #(
		.INIT('h135f)
	) name10673 (
		\s14_data_i[22]_pad ,
		\s2_data_i[22]_pad ,
		_w9348_,
		_w9541_,
		_w12574_
	);
	LUT4 #(
		.INIT('h135f)
	) name10674 (
		\s12_data_i[22]_pad ,
		\s5_data_i[22]_pad ,
		_w9354_,
		_w9547_,
		_w12575_
	);
	LUT4 #(
		.INIT('h135f)
	) name10675 (
		\s0_data_i[22]_pad ,
		\s13_data_i[22]_pad ,
		_w9305_,
		_w9538_,
		_w12576_
	);
	LUT4 #(
		.INIT('h4000)
	) name10676 (
		_w12573_,
		_w12574_,
		_w12575_,
		_w12576_,
		_w12577_
	);
	LUT2 #(
		.INIT('h8)
	) name10677 (
		_w12572_,
		_w12577_,
		_w12578_
	);
	LUT4 #(
		.INIT('h70ff)
	) name10678 (
		_w2046_,
		_w2097_,
		_w12567_,
		_w12578_,
		_w12579_
	);
	LUT2 #(
		.INIT('h8)
	) name10679 (
		\s15_data_i[23]_pad ,
		_w2064_,
		_w12580_
	);
	LUT4 #(
		.INIT('h135f)
	) name10680 (
		\s1_data_i[23]_pad ,
		\s8_data_i[23]_pad ,
		_w9269_,
		_w9553_,
		_w12581_
	);
	LUT4 #(
		.INIT('h135f)
	) name10681 (
		\s4_data_i[23]_pad ,
		\s6_data_i[23]_pad ,
		_w9544_,
		_w9550_,
		_w12582_
	);
	LUT4 #(
		.INIT('h135f)
	) name10682 (
		\s3_data_i[23]_pad ,
		\s9_data_i[23]_pad ,
		_w9351_,
		_w9556_,
		_w12583_
	);
	LUT4 #(
		.INIT('h153f)
	) name10683 (
		\s10_data_i[23]_pad ,
		\s7_data_i[23]_pad ,
		_w9345_,
		_w9532_,
		_w12584_
	);
	LUT4 #(
		.INIT('h8000)
	) name10684 (
		_w12581_,
		_w12582_,
		_w12583_,
		_w12584_,
		_w12585_
	);
	LUT2 #(
		.INIT('h8)
	) name10685 (
		\s11_data_i[23]_pad ,
		_w9535_,
		_w12586_
	);
	LUT4 #(
		.INIT('h135f)
	) name10686 (
		\s14_data_i[23]_pad ,
		\s2_data_i[23]_pad ,
		_w9348_,
		_w9541_,
		_w12587_
	);
	LUT4 #(
		.INIT('h135f)
	) name10687 (
		\s12_data_i[23]_pad ,
		\s5_data_i[23]_pad ,
		_w9354_,
		_w9547_,
		_w12588_
	);
	LUT4 #(
		.INIT('h135f)
	) name10688 (
		\s0_data_i[23]_pad ,
		\s13_data_i[23]_pad ,
		_w9305_,
		_w9538_,
		_w12589_
	);
	LUT4 #(
		.INIT('h4000)
	) name10689 (
		_w12586_,
		_w12587_,
		_w12588_,
		_w12589_,
		_w12590_
	);
	LUT2 #(
		.INIT('h8)
	) name10690 (
		_w12585_,
		_w12590_,
		_w12591_
	);
	LUT4 #(
		.INIT('h70ff)
	) name10691 (
		_w2046_,
		_w2097_,
		_w12580_,
		_w12591_,
		_w12592_
	);
	LUT2 #(
		.INIT('h8)
	) name10692 (
		\s15_data_i[24]_pad ,
		_w2064_,
		_w12593_
	);
	LUT4 #(
		.INIT('h135f)
	) name10693 (
		\s1_data_i[24]_pad ,
		\s8_data_i[24]_pad ,
		_w9269_,
		_w9553_,
		_w12594_
	);
	LUT4 #(
		.INIT('h135f)
	) name10694 (
		\s4_data_i[24]_pad ,
		\s6_data_i[24]_pad ,
		_w9544_,
		_w9550_,
		_w12595_
	);
	LUT4 #(
		.INIT('h135f)
	) name10695 (
		\s3_data_i[24]_pad ,
		\s9_data_i[24]_pad ,
		_w9351_,
		_w9556_,
		_w12596_
	);
	LUT4 #(
		.INIT('h153f)
	) name10696 (
		\s10_data_i[24]_pad ,
		\s7_data_i[24]_pad ,
		_w9345_,
		_w9532_,
		_w12597_
	);
	LUT4 #(
		.INIT('h8000)
	) name10697 (
		_w12594_,
		_w12595_,
		_w12596_,
		_w12597_,
		_w12598_
	);
	LUT2 #(
		.INIT('h8)
	) name10698 (
		\s11_data_i[24]_pad ,
		_w9535_,
		_w12599_
	);
	LUT4 #(
		.INIT('h135f)
	) name10699 (
		\s14_data_i[24]_pad ,
		\s2_data_i[24]_pad ,
		_w9348_,
		_w9541_,
		_w12600_
	);
	LUT4 #(
		.INIT('h135f)
	) name10700 (
		\s12_data_i[24]_pad ,
		\s5_data_i[24]_pad ,
		_w9354_,
		_w9547_,
		_w12601_
	);
	LUT4 #(
		.INIT('h135f)
	) name10701 (
		\s0_data_i[24]_pad ,
		\s13_data_i[24]_pad ,
		_w9305_,
		_w9538_,
		_w12602_
	);
	LUT4 #(
		.INIT('h4000)
	) name10702 (
		_w12599_,
		_w12600_,
		_w12601_,
		_w12602_,
		_w12603_
	);
	LUT2 #(
		.INIT('h8)
	) name10703 (
		_w12598_,
		_w12603_,
		_w12604_
	);
	LUT4 #(
		.INIT('h70ff)
	) name10704 (
		_w2046_,
		_w2097_,
		_w12593_,
		_w12604_,
		_w12605_
	);
	LUT2 #(
		.INIT('h8)
	) name10705 (
		\s15_data_i[25]_pad ,
		_w2064_,
		_w12606_
	);
	LUT4 #(
		.INIT('h135f)
	) name10706 (
		\s1_data_i[25]_pad ,
		\s8_data_i[25]_pad ,
		_w9269_,
		_w9553_,
		_w12607_
	);
	LUT4 #(
		.INIT('h135f)
	) name10707 (
		\s4_data_i[25]_pad ,
		\s6_data_i[25]_pad ,
		_w9544_,
		_w9550_,
		_w12608_
	);
	LUT4 #(
		.INIT('h135f)
	) name10708 (
		\s3_data_i[25]_pad ,
		\s9_data_i[25]_pad ,
		_w9351_,
		_w9556_,
		_w12609_
	);
	LUT4 #(
		.INIT('h153f)
	) name10709 (
		\s10_data_i[25]_pad ,
		\s7_data_i[25]_pad ,
		_w9345_,
		_w9532_,
		_w12610_
	);
	LUT4 #(
		.INIT('h8000)
	) name10710 (
		_w12607_,
		_w12608_,
		_w12609_,
		_w12610_,
		_w12611_
	);
	LUT2 #(
		.INIT('h8)
	) name10711 (
		\s11_data_i[25]_pad ,
		_w9535_,
		_w12612_
	);
	LUT4 #(
		.INIT('h135f)
	) name10712 (
		\s14_data_i[25]_pad ,
		\s2_data_i[25]_pad ,
		_w9348_,
		_w9541_,
		_w12613_
	);
	LUT4 #(
		.INIT('h135f)
	) name10713 (
		\s12_data_i[25]_pad ,
		\s5_data_i[25]_pad ,
		_w9354_,
		_w9547_,
		_w12614_
	);
	LUT4 #(
		.INIT('h135f)
	) name10714 (
		\s0_data_i[25]_pad ,
		\s13_data_i[25]_pad ,
		_w9305_,
		_w9538_,
		_w12615_
	);
	LUT4 #(
		.INIT('h4000)
	) name10715 (
		_w12612_,
		_w12613_,
		_w12614_,
		_w12615_,
		_w12616_
	);
	LUT2 #(
		.INIT('h8)
	) name10716 (
		_w12611_,
		_w12616_,
		_w12617_
	);
	LUT4 #(
		.INIT('h70ff)
	) name10717 (
		_w2046_,
		_w2097_,
		_w12606_,
		_w12617_,
		_w12618_
	);
	LUT2 #(
		.INIT('h8)
	) name10718 (
		\s15_data_i[26]_pad ,
		_w2064_,
		_w12619_
	);
	LUT4 #(
		.INIT('h135f)
	) name10719 (
		\s1_data_i[26]_pad ,
		\s8_data_i[26]_pad ,
		_w9269_,
		_w9553_,
		_w12620_
	);
	LUT4 #(
		.INIT('h135f)
	) name10720 (
		\s4_data_i[26]_pad ,
		\s6_data_i[26]_pad ,
		_w9544_,
		_w9550_,
		_w12621_
	);
	LUT4 #(
		.INIT('h135f)
	) name10721 (
		\s3_data_i[26]_pad ,
		\s9_data_i[26]_pad ,
		_w9351_,
		_w9556_,
		_w12622_
	);
	LUT4 #(
		.INIT('h153f)
	) name10722 (
		\s10_data_i[26]_pad ,
		\s7_data_i[26]_pad ,
		_w9345_,
		_w9532_,
		_w12623_
	);
	LUT4 #(
		.INIT('h8000)
	) name10723 (
		_w12620_,
		_w12621_,
		_w12622_,
		_w12623_,
		_w12624_
	);
	LUT2 #(
		.INIT('h8)
	) name10724 (
		\s11_data_i[26]_pad ,
		_w9535_,
		_w12625_
	);
	LUT4 #(
		.INIT('h135f)
	) name10725 (
		\s14_data_i[26]_pad ,
		\s2_data_i[26]_pad ,
		_w9348_,
		_w9541_,
		_w12626_
	);
	LUT4 #(
		.INIT('h135f)
	) name10726 (
		\s12_data_i[26]_pad ,
		\s5_data_i[26]_pad ,
		_w9354_,
		_w9547_,
		_w12627_
	);
	LUT4 #(
		.INIT('h135f)
	) name10727 (
		\s0_data_i[26]_pad ,
		\s13_data_i[26]_pad ,
		_w9305_,
		_w9538_,
		_w12628_
	);
	LUT4 #(
		.INIT('h4000)
	) name10728 (
		_w12625_,
		_w12626_,
		_w12627_,
		_w12628_,
		_w12629_
	);
	LUT2 #(
		.INIT('h8)
	) name10729 (
		_w12624_,
		_w12629_,
		_w12630_
	);
	LUT4 #(
		.INIT('h70ff)
	) name10730 (
		_w2046_,
		_w2097_,
		_w12619_,
		_w12630_,
		_w12631_
	);
	LUT2 #(
		.INIT('h8)
	) name10731 (
		\s15_data_i[27]_pad ,
		_w2064_,
		_w12632_
	);
	LUT4 #(
		.INIT('h135f)
	) name10732 (
		\s1_data_i[27]_pad ,
		\s8_data_i[27]_pad ,
		_w9269_,
		_w9553_,
		_w12633_
	);
	LUT4 #(
		.INIT('h135f)
	) name10733 (
		\s4_data_i[27]_pad ,
		\s6_data_i[27]_pad ,
		_w9544_,
		_w9550_,
		_w12634_
	);
	LUT4 #(
		.INIT('h135f)
	) name10734 (
		\s3_data_i[27]_pad ,
		\s9_data_i[27]_pad ,
		_w9351_,
		_w9556_,
		_w12635_
	);
	LUT4 #(
		.INIT('h153f)
	) name10735 (
		\s10_data_i[27]_pad ,
		\s7_data_i[27]_pad ,
		_w9345_,
		_w9532_,
		_w12636_
	);
	LUT4 #(
		.INIT('h8000)
	) name10736 (
		_w12633_,
		_w12634_,
		_w12635_,
		_w12636_,
		_w12637_
	);
	LUT2 #(
		.INIT('h8)
	) name10737 (
		\s11_data_i[27]_pad ,
		_w9535_,
		_w12638_
	);
	LUT4 #(
		.INIT('h135f)
	) name10738 (
		\s14_data_i[27]_pad ,
		\s2_data_i[27]_pad ,
		_w9348_,
		_w9541_,
		_w12639_
	);
	LUT4 #(
		.INIT('h135f)
	) name10739 (
		\s12_data_i[27]_pad ,
		\s5_data_i[27]_pad ,
		_w9354_,
		_w9547_,
		_w12640_
	);
	LUT4 #(
		.INIT('h135f)
	) name10740 (
		\s0_data_i[27]_pad ,
		\s13_data_i[27]_pad ,
		_w9305_,
		_w9538_,
		_w12641_
	);
	LUT4 #(
		.INIT('h4000)
	) name10741 (
		_w12638_,
		_w12639_,
		_w12640_,
		_w12641_,
		_w12642_
	);
	LUT2 #(
		.INIT('h8)
	) name10742 (
		_w12637_,
		_w12642_,
		_w12643_
	);
	LUT4 #(
		.INIT('h70ff)
	) name10743 (
		_w2046_,
		_w2097_,
		_w12632_,
		_w12643_,
		_w12644_
	);
	LUT2 #(
		.INIT('h8)
	) name10744 (
		\s15_data_i[28]_pad ,
		_w2064_,
		_w12645_
	);
	LUT4 #(
		.INIT('h135f)
	) name10745 (
		\s1_data_i[28]_pad ,
		\s8_data_i[28]_pad ,
		_w9269_,
		_w9553_,
		_w12646_
	);
	LUT4 #(
		.INIT('h135f)
	) name10746 (
		\s4_data_i[28]_pad ,
		\s6_data_i[28]_pad ,
		_w9544_,
		_w9550_,
		_w12647_
	);
	LUT4 #(
		.INIT('h135f)
	) name10747 (
		\s3_data_i[28]_pad ,
		\s9_data_i[28]_pad ,
		_w9351_,
		_w9556_,
		_w12648_
	);
	LUT4 #(
		.INIT('h153f)
	) name10748 (
		\s10_data_i[28]_pad ,
		\s7_data_i[28]_pad ,
		_w9345_,
		_w9532_,
		_w12649_
	);
	LUT4 #(
		.INIT('h8000)
	) name10749 (
		_w12646_,
		_w12647_,
		_w12648_,
		_w12649_,
		_w12650_
	);
	LUT2 #(
		.INIT('h8)
	) name10750 (
		\s11_data_i[28]_pad ,
		_w9535_,
		_w12651_
	);
	LUT4 #(
		.INIT('h135f)
	) name10751 (
		\s14_data_i[28]_pad ,
		\s2_data_i[28]_pad ,
		_w9348_,
		_w9541_,
		_w12652_
	);
	LUT4 #(
		.INIT('h135f)
	) name10752 (
		\s12_data_i[28]_pad ,
		\s5_data_i[28]_pad ,
		_w9354_,
		_w9547_,
		_w12653_
	);
	LUT4 #(
		.INIT('h135f)
	) name10753 (
		\s0_data_i[28]_pad ,
		\s13_data_i[28]_pad ,
		_w9305_,
		_w9538_,
		_w12654_
	);
	LUT4 #(
		.INIT('h4000)
	) name10754 (
		_w12651_,
		_w12652_,
		_w12653_,
		_w12654_,
		_w12655_
	);
	LUT2 #(
		.INIT('h8)
	) name10755 (
		_w12650_,
		_w12655_,
		_w12656_
	);
	LUT4 #(
		.INIT('h70ff)
	) name10756 (
		_w2046_,
		_w2097_,
		_w12645_,
		_w12656_,
		_w12657_
	);
	LUT2 #(
		.INIT('h8)
	) name10757 (
		\s15_data_i[29]_pad ,
		_w2064_,
		_w12658_
	);
	LUT4 #(
		.INIT('h135f)
	) name10758 (
		\s1_data_i[29]_pad ,
		\s8_data_i[29]_pad ,
		_w9269_,
		_w9553_,
		_w12659_
	);
	LUT4 #(
		.INIT('h135f)
	) name10759 (
		\s4_data_i[29]_pad ,
		\s6_data_i[29]_pad ,
		_w9544_,
		_w9550_,
		_w12660_
	);
	LUT4 #(
		.INIT('h135f)
	) name10760 (
		\s3_data_i[29]_pad ,
		\s9_data_i[29]_pad ,
		_w9351_,
		_w9556_,
		_w12661_
	);
	LUT4 #(
		.INIT('h153f)
	) name10761 (
		\s10_data_i[29]_pad ,
		\s7_data_i[29]_pad ,
		_w9345_,
		_w9532_,
		_w12662_
	);
	LUT4 #(
		.INIT('h8000)
	) name10762 (
		_w12659_,
		_w12660_,
		_w12661_,
		_w12662_,
		_w12663_
	);
	LUT2 #(
		.INIT('h8)
	) name10763 (
		\s11_data_i[29]_pad ,
		_w9535_,
		_w12664_
	);
	LUT4 #(
		.INIT('h135f)
	) name10764 (
		\s14_data_i[29]_pad ,
		\s2_data_i[29]_pad ,
		_w9348_,
		_w9541_,
		_w12665_
	);
	LUT4 #(
		.INIT('h135f)
	) name10765 (
		\s12_data_i[29]_pad ,
		\s5_data_i[29]_pad ,
		_w9354_,
		_w9547_,
		_w12666_
	);
	LUT4 #(
		.INIT('h135f)
	) name10766 (
		\s0_data_i[29]_pad ,
		\s13_data_i[29]_pad ,
		_w9305_,
		_w9538_,
		_w12667_
	);
	LUT4 #(
		.INIT('h4000)
	) name10767 (
		_w12664_,
		_w12665_,
		_w12666_,
		_w12667_,
		_w12668_
	);
	LUT2 #(
		.INIT('h8)
	) name10768 (
		_w12663_,
		_w12668_,
		_w12669_
	);
	LUT4 #(
		.INIT('h70ff)
	) name10769 (
		_w2046_,
		_w2097_,
		_w12658_,
		_w12669_,
		_w12670_
	);
	LUT3 #(
		.INIT('h80)
	) name10770 (
		_w2064_,
		_w2097_,
		_w9993_,
		_w12671_
	);
	LUT2 #(
		.INIT('h8)
	) name10771 (
		\s15_data_i[2]_pad ,
		_w2064_,
		_w12672_
	);
	LUT3 #(
		.INIT('h70)
	) name10772 (
		_w2046_,
		_w2097_,
		_w12672_,
		_w12673_
	);
	LUT4 #(
		.INIT('h153f)
	) name10773 (
		\s12_data_i[2]_pad ,
		\s1_data_i[2]_pad ,
		_w9269_,
		_w9354_,
		_w12674_
	);
	LUT4 #(
		.INIT('h135f)
	) name10774 (
		\s0_data_i[2]_pad ,
		\s10_data_i[2]_pad ,
		_w9305_,
		_w9532_,
		_w12675_
	);
	LUT4 #(
		.INIT('h135f)
	) name10775 (
		\s3_data_i[2]_pad ,
		\s4_data_i[2]_pad ,
		_w9351_,
		_w9544_,
		_w12676_
	);
	LUT4 #(
		.INIT('h135f)
	) name10776 (
		\s6_data_i[2]_pad ,
		\s9_data_i[2]_pad ,
		_w9550_,
		_w9556_,
		_w12677_
	);
	LUT4 #(
		.INIT('h8000)
	) name10777 (
		_w12674_,
		_w12675_,
		_w12676_,
		_w12677_,
		_w12678_
	);
	LUT2 #(
		.INIT('h8)
	) name10778 (
		\s14_data_i[2]_pad ,
		_w9348_,
		_w12679_
	);
	LUT4 #(
		.INIT('h153f)
	) name10779 (
		\s11_data_i[2]_pad ,
		\s7_data_i[2]_pad ,
		_w9345_,
		_w9535_,
		_w12680_
	);
	LUT4 #(
		.INIT('h135f)
	) name10780 (
		\s5_data_i[2]_pad ,
		\s8_data_i[2]_pad ,
		_w9547_,
		_w9553_,
		_w12681_
	);
	LUT4 #(
		.INIT('h135f)
	) name10781 (
		\s13_data_i[2]_pad ,
		\s2_data_i[2]_pad ,
		_w9538_,
		_w9541_,
		_w12682_
	);
	LUT4 #(
		.INIT('h4000)
	) name10782 (
		_w12679_,
		_w12680_,
		_w12681_,
		_w12682_,
		_w12683_
	);
	LUT2 #(
		.INIT('h8)
	) name10783 (
		_w12678_,
		_w12683_,
		_w12684_
	);
	LUT3 #(
		.INIT('hef)
	) name10784 (
		_w12671_,
		_w12673_,
		_w12684_,
		_w12685_
	);
	LUT2 #(
		.INIT('h8)
	) name10785 (
		\s15_data_i[30]_pad ,
		_w2064_,
		_w12686_
	);
	LUT4 #(
		.INIT('h135f)
	) name10786 (
		\s1_data_i[30]_pad ,
		\s8_data_i[30]_pad ,
		_w9269_,
		_w9553_,
		_w12687_
	);
	LUT4 #(
		.INIT('h135f)
	) name10787 (
		\s4_data_i[30]_pad ,
		\s6_data_i[30]_pad ,
		_w9544_,
		_w9550_,
		_w12688_
	);
	LUT4 #(
		.INIT('h135f)
	) name10788 (
		\s3_data_i[30]_pad ,
		\s9_data_i[30]_pad ,
		_w9351_,
		_w9556_,
		_w12689_
	);
	LUT4 #(
		.INIT('h153f)
	) name10789 (
		\s10_data_i[30]_pad ,
		\s7_data_i[30]_pad ,
		_w9345_,
		_w9532_,
		_w12690_
	);
	LUT4 #(
		.INIT('h8000)
	) name10790 (
		_w12687_,
		_w12688_,
		_w12689_,
		_w12690_,
		_w12691_
	);
	LUT2 #(
		.INIT('h8)
	) name10791 (
		\s11_data_i[30]_pad ,
		_w9535_,
		_w12692_
	);
	LUT4 #(
		.INIT('h135f)
	) name10792 (
		\s14_data_i[30]_pad ,
		\s2_data_i[30]_pad ,
		_w9348_,
		_w9541_,
		_w12693_
	);
	LUT4 #(
		.INIT('h135f)
	) name10793 (
		\s12_data_i[30]_pad ,
		\s5_data_i[30]_pad ,
		_w9354_,
		_w9547_,
		_w12694_
	);
	LUT4 #(
		.INIT('h135f)
	) name10794 (
		\s0_data_i[30]_pad ,
		\s13_data_i[30]_pad ,
		_w9305_,
		_w9538_,
		_w12695_
	);
	LUT4 #(
		.INIT('h4000)
	) name10795 (
		_w12692_,
		_w12693_,
		_w12694_,
		_w12695_,
		_w12696_
	);
	LUT2 #(
		.INIT('h8)
	) name10796 (
		_w12691_,
		_w12696_,
		_w12697_
	);
	LUT4 #(
		.INIT('h70ff)
	) name10797 (
		_w2046_,
		_w2097_,
		_w12686_,
		_w12697_,
		_w12698_
	);
	LUT2 #(
		.INIT('h8)
	) name10798 (
		\s15_data_i[31]_pad ,
		_w2064_,
		_w12699_
	);
	LUT4 #(
		.INIT('h135f)
	) name10799 (
		\s1_data_i[31]_pad ,
		\s8_data_i[31]_pad ,
		_w9269_,
		_w9553_,
		_w12700_
	);
	LUT4 #(
		.INIT('h135f)
	) name10800 (
		\s4_data_i[31]_pad ,
		\s6_data_i[31]_pad ,
		_w9544_,
		_w9550_,
		_w12701_
	);
	LUT4 #(
		.INIT('h135f)
	) name10801 (
		\s3_data_i[31]_pad ,
		\s9_data_i[31]_pad ,
		_w9351_,
		_w9556_,
		_w12702_
	);
	LUT4 #(
		.INIT('h153f)
	) name10802 (
		\s10_data_i[31]_pad ,
		\s7_data_i[31]_pad ,
		_w9345_,
		_w9532_,
		_w12703_
	);
	LUT4 #(
		.INIT('h8000)
	) name10803 (
		_w12700_,
		_w12701_,
		_w12702_,
		_w12703_,
		_w12704_
	);
	LUT2 #(
		.INIT('h8)
	) name10804 (
		\s11_data_i[31]_pad ,
		_w9535_,
		_w12705_
	);
	LUT4 #(
		.INIT('h135f)
	) name10805 (
		\s14_data_i[31]_pad ,
		\s2_data_i[31]_pad ,
		_w9348_,
		_w9541_,
		_w12706_
	);
	LUT4 #(
		.INIT('h135f)
	) name10806 (
		\s12_data_i[31]_pad ,
		\s5_data_i[31]_pad ,
		_w9354_,
		_w9547_,
		_w12707_
	);
	LUT4 #(
		.INIT('h135f)
	) name10807 (
		\s0_data_i[31]_pad ,
		\s13_data_i[31]_pad ,
		_w9305_,
		_w9538_,
		_w12708_
	);
	LUT4 #(
		.INIT('h4000)
	) name10808 (
		_w12705_,
		_w12706_,
		_w12707_,
		_w12708_,
		_w12709_
	);
	LUT2 #(
		.INIT('h8)
	) name10809 (
		_w12704_,
		_w12709_,
		_w12710_
	);
	LUT4 #(
		.INIT('h70ff)
	) name10810 (
		_w2046_,
		_w2097_,
		_w12699_,
		_w12710_,
		_w12711_
	);
	LUT3 #(
		.INIT('h80)
	) name10811 (
		_w2064_,
		_w2097_,
		_w10035_,
		_w12712_
	);
	LUT2 #(
		.INIT('h8)
	) name10812 (
		\s15_data_i[3]_pad ,
		_w2064_,
		_w12713_
	);
	LUT3 #(
		.INIT('h70)
	) name10813 (
		_w2046_,
		_w2097_,
		_w12713_,
		_w12714_
	);
	LUT4 #(
		.INIT('h153f)
	) name10814 (
		\s12_data_i[3]_pad ,
		\s1_data_i[3]_pad ,
		_w9269_,
		_w9354_,
		_w12715_
	);
	LUT4 #(
		.INIT('h135f)
	) name10815 (
		\s4_data_i[3]_pad ,
		\s6_data_i[3]_pad ,
		_w9544_,
		_w9550_,
		_w12716_
	);
	LUT4 #(
		.INIT('h135f)
	) name10816 (
		\s3_data_i[3]_pad ,
		\s9_data_i[3]_pad ,
		_w9351_,
		_w9556_,
		_w12717_
	);
	LUT4 #(
		.INIT('h153f)
	) name10817 (
		\s10_data_i[3]_pad ,
		\s7_data_i[3]_pad ,
		_w9345_,
		_w9532_,
		_w12718_
	);
	LUT4 #(
		.INIT('h8000)
	) name10818 (
		_w12715_,
		_w12716_,
		_w12717_,
		_w12718_,
		_w12719_
	);
	LUT2 #(
		.INIT('h8)
	) name10819 (
		\s14_data_i[3]_pad ,
		_w9348_,
		_w12720_
	);
	LUT4 #(
		.INIT('h135f)
	) name10820 (
		\s11_data_i[3]_pad ,
		\s2_data_i[3]_pad ,
		_w9535_,
		_w9541_,
		_w12721_
	);
	LUT4 #(
		.INIT('h135f)
	) name10821 (
		\s5_data_i[3]_pad ,
		\s8_data_i[3]_pad ,
		_w9547_,
		_w9553_,
		_w12722_
	);
	LUT4 #(
		.INIT('h135f)
	) name10822 (
		\s0_data_i[3]_pad ,
		\s13_data_i[3]_pad ,
		_w9305_,
		_w9538_,
		_w12723_
	);
	LUT4 #(
		.INIT('h4000)
	) name10823 (
		_w12720_,
		_w12721_,
		_w12722_,
		_w12723_,
		_w12724_
	);
	LUT2 #(
		.INIT('h8)
	) name10824 (
		_w12719_,
		_w12724_,
		_w12725_
	);
	LUT3 #(
		.INIT('hef)
	) name10825 (
		_w12712_,
		_w12714_,
		_w12725_,
		_w12726_
	);
	LUT3 #(
		.INIT('h80)
	) name10826 (
		_w2064_,
		_w2097_,
		_w10051_,
		_w12727_
	);
	LUT2 #(
		.INIT('h8)
	) name10827 (
		\s15_data_i[4]_pad ,
		_w2064_,
		_w12728_
	);
	LUT3 #(
		.INIT('h70)
	) name10828 (
		_w2046_,
		_w2097_,
		_w12728_,
		_w12729_
	);
	LUT4 #(
		.INIT('h153f)
	) name10829 (
		\s12_data_i[4]_pad ,
		\s1_data_i[4]_pad ,
		_w9269_,
		_w9354_,
		_w12730_
	);
	LUT4 #(
		.INIT('h135f)
	) name10830 (
		\s0_data_i[4]_pad ,
		\s10_data_i[4]_pad ,
		_w9305_,
		_w9532_,
		_w12731_
	);
	LUT4 #(
		.INIT('h135f)
	) name10831 (
		\s3_data_i[4]_pad ,
		\s4_data_i[4]_pad ,
		_w9351_,
		_w9544_,
		_w12732_
	);
	LUT4 #(
		.INIT('h135f)
	) name10832 (
		\s6_data_i[4]_pad ,
		\s9_data_i[4]_pad ,
		_w9550_,
		_w9556_,
		_w12733_
	);
	LUT4 #(
		.INIT('h8000)
	) name10833 (
		_w12730_,
		_w12731_,
		_w12732_,
		_w12733_,
		_w12734_
	);
	LUT2 #(
		.INIT('h8)
	) name10834 (
		\s14_data_i[4]_pad ,
		_w9348_,
		_w12735_
	);
	LUT4 #(
		.INIT('h153f)
	) name10835 (
		\s11_data_i[4]_pad ,
		\s7_data_i[4]_pad ,
		_w9345_,
		_w9535_,
		_w12736_
	);
	LUT4 #(
		.INIT('h135f)
	) name10836 (
		\s5_data_i[4]_pad ,
		\s8_data_i[4]_pad ,
		_w9547_,
		_w9553_,
		_w12737_
	);
	LUT4 #(
		.INIT('h135f)
	) name10837 (
		\s13_data_i[4]_pad ,
		\s2_data_i[4]_pad ,
		_w9538_,
		_w9541_,
		_w12738_
	);
	LUT4 #(
		.INIT('h4000)
	) name10838 (
		_w12735_,
		_w12736_,
		_w12737_,
		_w12738_,
		_w12739_
	);
	LUT2 #(
		.INIT('h8)
	) name10839 (
		_w12734_,
		_w12739_,
		_w12740_
	);
	LUT3 #(
		.INIT('hef)
	) name10840 (
		_w12727_,
		_w12729_,
		_w12740_,
		_w12741_
	);
	LUT3 #(
		.INIT('h80)
	) name10841 (
		_w2064_,
		_w2097_,
		_w10067_,
		_w12742_
	);
	LUT2 #(
		.INIT('h8)
	) name10842 (
		\s15_data_i[5]_pad ,
		_w2064_,
		_w12743_
	);
	LUT3 #(
		.INIT('h70)
	) name10843 (
		_w2046_,
		_w2097_,
		_w12743_,
		_w12744_
	);
	LUT4 #(
		.INIT('h153f)
	) name10844 (
		\s12_data_i[5]_pad ,
		\s1_data_i[5]_pad ,
		_w9269_,
		_w9354_,
		_w12745_
	);
	LUT4 #(
		.INIT('h135f)
	) name10845 (
		\s7_data_i[5]_pad ,
		\s9_data_i[5]_pad ,
		_w9345_,
		_w9556_,
		_w12746_
	);
	LUT4 #(
		.INIT('h135f)
	) name10846 (
		\s3_data_i[5]_pad ,
		\s6_data_i[5]_pad ,
		_w9351_,
		_w9550_,
		_w12747_
	);
	LUT4 #(
		.INIT('h135f)
	) name10847 (
		\s10_data_i[5]_pad ,
		\s13_data_i[5]_pad ,
		_w9532_,
		_w9538_,
		_w12748_
	);
	LUT4 #(
		.INIT('h8000)
	) name10848 (
		_w12745_,
		_w12746_,
		_w12747_,
		_w12748_,
		_w12749_
	);
	LUT2 #(
		.INIT('h8)
	) name10849 (
		\s14_data_i[5]_pad ,
		_w9348_,
		_w12750_
	);
	LUT4 #(
		.INIT('h135f)
	) name10850 (
		\s11_data_i[5]_pad ,
		\s2_data_i[5]_pad ,
		_w9535_,
		_w9541_,
		_w12751_
	);
	LUT4 #(
		.INIT('h135f)
	) name10851 (
		\s5_data_i[5]_pad ,
		\s8_data_i[5]_pad ,
		_w9547_,
		_w9553_,
		_w12752_
	);
	LUT4 #(
		.INIT('h135f)
	) name10852 (
		\s0_data_i[5]_pad ,
		\s4_data_i[5]_pad ,
		_w9305_,
		_w9544_,
		_w12753_
	);
	LUT4 #(
		.INIT('h4000)
	) name10853 (
		_w12750_,
		_w12751_,
		_w12752_,
		_w12753_,
		_w12754_
	);
	LUT2 #(
		.INIT('h8)
	) name10854 (
		_w12749_,
		_w12754_,
		_w12755_
	);
	LUT3 #(
		.INIT('hef)
	) name10855 (
		_w12742_,
		_w12744_,
		_w12755_,
		_w12756_
	);
	LUT3 #(
		.INIT('h80)
	) name10856 (
		_w2064_,
		_w2097_,
		_w10083_,
		_w12757_
	);
	LUT2 #(
		.INIT('h8)
	) name10857 (
		\s15_data_i[6]_pad ,
		_w2064_,
		_w12758_
	);
	LUT3 #(
		.INIT('h70)
	) name10858 (
		_w2046_,
		_w2097_,
		_w12758_,
		_w12759_
	);
	LUT4 #(
		.INIT('h153f)
	) name10859 (
		\s12_data_i[6]_pad ,
		\s1_data_i[6]_pad ,
		_w9269_,
		_w9354_,
		_w12760_
	);
	LUT4 #(
		.INIT('h135f)
	) name10860 (
		\s0_data_i[6]_pad ,
		\s10_data_i[6]_pad ,
		_w9305_,
		_w9532_,
		_w12761_
	);
	LUT4 #(
		.INIT('h135f)
	) name10861 (
		\s3_data_i[6]_pad ,
		\s4_data_i[6]_pad ,
		_w9351_,
		_w9544_,
		_w12762_
	);
	LUT4 #(
		.INIT('h135f)
	) name10862 (
		\s6_data_i[6]_pad ,
		\s9_data_i[6]_pad ,
		_w9550_,
		_w9556_,
		_w12763_
	);
	LUT4 #(
		.INIT('h8000)
	) name10863 (
		_w12760_,
		_w12761_,
		_w12762_,
		_w12763_,
		_w12764_
	);
	LUT2 #(
		.INIT('h8)
	) name10864 (
		\s14_data_i[6]_pad ,
		_w9348_,
		_w12765_
	);
	LUT4 #(
		.INIT('h153f)
	) name10865 (
		\s11_data_i[6]_pad ,
		\s7_data_i[6]_pad ,
		_w9345_,
		_w9535_,
		_w12766_
	);
	LUT4 #(
		.INIT('h135f)
	) name10866 (
		\s5_data_i[6]_pad ,
		\s8_data_i[6]_pad ,
		_w9547_,
		_w9553_,
		_w12767_
	);
	LUT4 #(
		.INIT('h135f)
	) name10867 (
		\s13_data_i[6]_pad ,
		\s2_data_i[6]_pad ,
		_w9538_,
		_w9541_,
		_w12768_
	);
	LUT4 #(
		.INIT('h4000)
	) name10868 (
		_w12765_,
		_w12766_,
		_w12767_,
		_w12768_,
		_w12769_
	);
	LUT2 #(
		.INIT('h8)
	) name10869 (
		_w12764_,
		_w12769_,
		_w12770_
	);
	LUT3 #(
		.INIT('hef)
	) name10870 (
		_w12757_,
		_w12759_,
		_w12770_,
		_w12771_
	);
	LUT3 #(
		.INIT('h80)
	) name10871 (
		_w2064_,
		_w2097_,
		_w10099_,
		_w12772_
	);
	LUT2 #(
		.INIT('h8)
	) name10872 (
		\s15_data_i[7]_pad ,
		_w2064_,
		_w12773_
	);
	LUT3 #(
		.INIT('h70)
	) name10873 (
		_w2046_,
		_w2097_,
		_w12773_,
		_w12774_
	);
	LUT4 #(
		.INIT('h153f)
	) name10874 (
		\s12_data_i[7]_pad ,
		\s1_data_i[7]_pad ,
		_w9269_,
		_w9354_,
		_w12775_
	);
	LUT4 #(
		.INIT('h135f)
	) name10875 (
		\s0_data_i[7]_pad ,
		\s10_data_i[7]_pad ,
		_w9305_,
		_w9532_,
		_w12776_
	);
	LUT4 #(
		.INIT('h135f)
	) name10876 (
		\s3_data_i[7]_pad ,
		\s4_data_i[7]_pad ,
		_w9351_,
		_w9544_,
		_w12777_
	);
	LUT4 #(
		.INIT('h135f)
	) name10877 (
		\s6_data_i[7]_pad ,
		\s9_data_i[7]_pad ,
		_w9550_,
		_w9556_,
		_w12778_
	);
	LUT4 #(
		.INIT('h8000)
	) name10878 (
		_w12775_,
		_w12776_,
		_w12777_,
		_w12778_,
		_w12779_
	);
	LUT2 #(
		.INIT('h8)
	) name10879 (
		\s14_data_i[7]_pad ,
		_w9348_,
		_w12780_
	);
	LUT4 #(
		.INIT('h153f)
	) name10880 (
		\s11_data_i[7]_pad ,
		\s7_data_i[7]_pad ,
		_w9345_,
		_w9535_,
		_w12781_
	);
	LUT4 #(
		.INIT('h135f)
	) name10881 (
		\s5_data_i[7]_pad ,
		\s8_data_i[7]_pad ,
		_w9547_,
		_w9553_,
		_w12782_
	);
	LUT4 #(
		.INIT('h135f)
	) name10882 (
		\s13_data_i[7]_pad ,
		\s2_data_i[7]_pad ,
		_w9538_,
		_w9541_,
		_w12783_
	);
	LUT4 #(
		.INIT('h4000)
	) name10883 (
		_w12780_,
		_w12781_,
		_w12782_,
		_w12783_,
		_w12784_
	);
	LUT2 #(
		.INIT('h8)
	) name10884 (
		_w12779_,
		_w12784_,
		_w12785_
	);
	LUT3 #(
		.INIT('hef)
	) name10885 (
		_w12772_,
		_w12774_,
		_w12785_,
		_w12786_
	);
	LUT3 #(
		.INIT('h80)
	) name10886 (
		_w2064_,
		_w2097_,
		_w10115_,
		_w12787_
	);
	LUT2 #(
		.INIT('h8)
	) name10887 (
		\s15_data_i[8]_pad ,
		_w2064_,
		_w12788_
	);
	LUT3 #(
		.INIT('h70)
	) name10888 (
		_w2046_,
		_w2097_,
		_w12788_,
		_w12789_
	);
	LUT4 #(
		.INIT('h153f)
	) name10889 (
		\s12_data_i[8]_pad ,
		\s1_data_i[8]_pad ,
		_w9269_,
		_w9354_,
		_w12790_
	);
	LUT4 #(
		.INIT('h135f)
	) name10890 (
		\s0_data_i[8]_pad ,
		\s10_data_i[8]_pad ,
		_w9305_,
		_w9532_,
		_w12791_
	);
	LUT4 #(
		.INIT('h135f)
	) name10891 (
		\s3_data_i[8]_pad ,
		\s4_data_i[8]_pad ,
		_w9351_,
		_w9544_,
		_w12792_
	);
	LUT4 #(
		.INIT('h135f)
	) name10892 (
		\s6_data_i[8]_pad ,
		\s9_data_i[8]_pad ,
		_w9550_,
		_w9556_,
		_w12793_
	);
	LUT4 #(
		.INIT('h8000)
	) name10893 (
		_w12790_,
		_w12791_,
		_w12792_,
		_w12793_,
		_w12794_
	);
	LUT2 #(
		.INIT('h8)
	) name10894 (
		\s14_data_i[8]_pad ,
		_w9348_,
		_w12795_
	);
	LUT4 #(
		.INIT('h153f)
	) name10895 (
		\s11_data_i[8]_pad ,
		\s7_data_i[8]_pad ,
		_w9345_,
		_w9535_,
		_w12796_
	);
	LUT4 #(
		.INIT('h135f)
	) name10896 (
		\s5_data_i[8]_pad ,
		\s8_data_i[8]_pad ,
		_w9547_,
		_w9553_,
		_w12797_
	);
	LUT4 #(
		.INIT('h135f)
	) name10897 (
		\s13_data_i[8]_pad ,
		\s2_data_i[8]_pad ,
		_w9538_,
		_w9541_,
		_w12798_
	);
	LUT4 #(
		.INIT('h4000)
	) name10898 (
		_w12795_,
		_w12796_,
		_w12797_,
		_w12798_,
		_w12799_
	);
	LUT2 #(
		.INIT('h8)
	) name10899 (
		_w12794_,
		_w12799_,
		_w12800_
	);
	LUT3 #(
		.INIT('hef)
	) name10900 (
		_w12787_,
		_w12789_,
		_w12800_,
		_w12801_
	);
	LUT3 #(
		.INIT('h80)
	) name10901 (
		_w2064_,
		_w2097_,
		_w10131_,
		_w12802_
	);
	LUT2 #(
		.INIT('h8)
	) name10902 (
		\s15_data_i[9]_pad ,
		_w2064_,
		_w12803_
	);
	LUT3 #(
		.INIT('h70)
	) name10903 (
		_w2046_,
		_w2097_,
		_w12803_,
		_w12804_
	);
	LUT4 #(
		.INIT('h153f)
	) name10904 (
		\s12_data_i[9]_pad ,
		\s1_data_i[9]_pad ,
		_w9269_,
		_w9354_,
		_w12805_
	);
	LUT4 #(
		.INIT('h135f)
	) name10905 (
		\s0_data_i[9]_pad ,
		\s10_data_i[9]_pad ,
		_w9305_,
		_w9532_,
		_w12806_
	);
	LUT4 #(
		.INIT('h135f)
	) name10906 (
		\s3_data_i[9]_pad ,
		\s4_data_i[9]_pad ,
		_w9351_,
		_w9544_,
		_w12807_
	);
	LUT4 #(
		.INIT('h135f)
	) name10907 (
		\s6_data_i[9]_pad ,
		\s9_data_i[9]_pad ,
		_w9550_,
		_w9556_,
		_w12808_
	);
	LUT4 #(
		.INIT('h8000)
	) name10908 (
		_w12805_,
		_w12806_,
		_w12807_,
		_w12808_,
		_w12809_
	);
	LUT2 #(
		.INIT('h8)
	) name10909 (
		\s14_data_i[9]_pad ,
		_w9348_,
		_w12810_
	);
	LUT4 #(
		.INIT('h153f)
	) name10910 (
		\s11_data_i[9]_pad ,
		\s7_data_i[9]_pad ,
		_w9345_,
		_w9535_,
		_w12811_
	);
	LUT4 #(
		.INIT('h135f)
	) name10911 (
		\s5_data_i[9]_pad ,
		\s8_data_i[9]_pad ,
		_w9547_,
		_w9553_,
		_w12812_
	);
	LUT4 #(
		.INIT('h135f)
	) name10912 (
		\s13_data_i[9]_pad ,
		\s2_data_i[9]_pad ,
		_w9538_,
		_w9541_,
		_w12813_
	);
	LUT4 #(
		.INIT('h4000)
	) name10913 (
		_w12810_,
		_w12811_,
		_w12812_,
		_w12813_,
		_w12814_
	);
	LUT2 #(
		.INIT('h8)
	) name10914 (
		_w12809_,
		_w12814_,
		_w12815_
	);
	LUT3 #(
		.INIT('hef)
	) name10915 (
		_w12802_,
		_w12804_,
		_w12815_,
		_w12816_
	);
	LUT3 #(
		.INIT('h80)
	) name10916 (
		\s15_err_i_pad ,
		_w1920_,
		_w12339_,
		_w12817_
	);
	LUT4 #(
		.INIT('h2a00)
	) name10917 (
		\s6_err_i_pad ,
		_w8743_,
		_w8744_,
		_w9550_,
		_w12818_
	);
	LUT4 #(
		.INIT('h2a00)
	) name10918 (
		\s1_err_i_pad ,
		_w9103_,
		_w9104_,
		_w9269_,
		_w12819_
	);
	LUT4 #(
		.INIT('h135f)
	) name10919 (
		_w8762_,
		_w9116_,
		_w12818_,
		_w12819_,
		_w12820_
	);
	LUT4 #(
		.INIT('h2a00)
	) name10920 (
		\s12_err_i_pad ,
		_w9029_,
		_w9030_,
		_w9354_,
		_w12821_
	);
	LUT4 #(
		.INIT('h2a00)
	) name10921 (
		\s13_err_i_pad ,
		_w9069_,
		_w9070_,
		_w9538_,
		_w12822_
	);
	LUT4 #(
		.INIT('h135f)
	) name10922 (
		_w9042_,
		_w9088_,
		_w12821_,
		_w12822_,
		_w12823_
	);
	LUT4 #(
		.INIT('h2a00)
	) name10923 (
		\s10_err_i_pad ,
		_w8910_,
		_w8911_,
		_w9532_,
		_w12824_
	);
	LUT4 #(
		.INIT('h2a00)
	) name10924 (
		\s5_err_i_pad ,
		_w8699_,
		_w8700_,
		_w9547_,
		_w12825_
	);
	LUT4 #(
		.INIT('h153f)
	) name10925 (
		_w8706_,
		_w8929_,
		_w12824_,
		_w12825_,
		_w12826_
	);
	LUT4 #(
		.INIT('h2a00)
	) name10926 (
		\s8_err_i_pad ,
		_w8821_,
		_w8822_,
		_w9553_,
		_w12827_
	);
	LUT4 #(
		.INIT('h2a00)
	) name10927 (
		\s0_err_i_pad ,
		_w8989_,
		_w8990_,
		_w9305_,
		_w12828_
	);
	LUT4 #(
		.INIT('h135f)
	) name10928 (
		_w8840_,
		_w8996_,
		_w12827_,
		_w12828_,
		_w12829_
	);
	LUT4 #(
		.INIT('h8000)
	) name10929 (
		_w12820_,
		_w12823_,
		_w12826_,
		_w12829_,
		_w12830_
	);
	LUT4 #(
		.INIT('h2a00)
	) name10930 (
		\s7_err_i_pad ,
		_w8782_,
		_w8783_,
		_w9345_,
		_w12831_
	);
	LUT2 #(
		.INIT('h8)
	) name10931 (
		_w8801_,
		_w12831_,
		_w12832_
	);
	LUT4 #(
		.INIT('h2a00)
	) name10932 (
		\s2_err_i_pad ,
		_w9171_,
		_w9172_,
		_w9541_,
		_w12833_
	);
	LUT4 #(
		.INIT('h2a00)
	) name10933 (
		\s4_err_i_pad ,
		_w8655_,
		_w8656_,
		_w9544_,
		_w12834_
	);
	LUT4 #(
		.INIT('h153f)
	) name10934 (
		_w8654_,
		_w9170_,
		_w12833_,
		_w12834_,
		_w12835_
	);
	LUT4 #(
		.INIT('h2a00)
	) name10935 (
		\s9_err_i_pad ,
		_w8865_,
		_w8866_,
		_w9556_,
		_w12836_
	);
	LUT4 #(
		.INIT('h2a00)
	) name10936 (
		\s3_err_i_pad ,
		_w9205_,
		_w9206_,
		_w9351_,
		_w12837_
	);
	LUT4 #(
		.INIT('h135f)
	) name10937 (
		_w8884_,
		_w9204_,
		_w12836_,
		_w12837_,
		_w12838_
	);
	LUT4 #(
		.INIT('h2a00)
	) name10938 (
		\s11_err_i_pad ,
		_w8955_,
		_w8956_,
		_w9535_,
		_w12839_
	);
	LUT4 #(
		.INIT('h2a00)
	) name10939 (
		\s14_err_i_pad ,
		_w9137_,
		_w9138_,
		_w9348_,
		_w12840_
	);
	LUT4 #(
		.INIT('h135f)
	) name10940 (
		_w8954_,
		_w9156_,
		_w12839_,
		_w12840_,
		_w12841_
	);
	LUT4 #(
		.INIT('h4000)
	) name10941 (
		_w12832_,
		_w12835_,
		_w12838_,
		_w12841_,
		_w12842_
	);
	LUT2 #(
		.INIT('h8)
	) name10942 (
		_w12830_,
		_w12842_,
		_w12843_
	);
	LUT4 #(
		.INIT('h70ff)
	) name10943 (
		_w2046_,
		_w2097_,
		_w12817_,
		_w12843_,
		_w12844_
	);
	LUT3 #(
		.INIT('h80)
	) name10944 (
		\s15_rty_i_pad ,
		_w1920_,
		_w12339_,
		_w12845_
	);
	LUT4 #(
		.INIT('h2a00)
	) name10945 (
		\s14_rty_i_pad ,
		_w9137_,
		_w9138_,
		_w9348_,
		_w12846_
	);
	LUT4 #(
		.INIT('h2a00)
	) name10946 (
		\s1_rty_i_pad ,
		_w9103_,
		_w9104_,
		_w9269_,
		_w12847_
	);
	LUT4 #(
		.INIT('h153f)
	) name10947 (
		_w9116_,
		_w9156_,
		_w12846_,
		_w12847_,
		_w12848_
	);
	LUT4 #(
		.INIT('h2a00)
	) name10948 (
		\s13_rty_i_pad ,
		_w9069_,
		_w9070_,
		_w9538_,
		_w12849_
	);
	LUT4 #(
		.INIT('h2a00)
	) name10949 (
		\s9_rty_i_pad ,
		_w8865_,
		_w8866_,
		_w9556_,
		_w12850_
	);
	LUT4 #(
		.INIT('h153f)
	) name10950 (
		_w8884_,
		_w9088_,
		_w12849_,
		_w12850_,
		_w12851_
	);
	LUT4 #(
		.INIT('h2a00)
	) name10951 (
		\s0_rty_i_pad ,
		_w8989_,
		_w8990_,
		_w9305_,
		_w12852_
	);
	LUT4 #(
		.INIT('h2a00)
	) name10952 (
		\s6_rty_i_pad ,
		_w8743_,
		_w8744_,
		_w9550_,
		_w12853_
	);
	LUT4 #(
		.INIT('h153f)
	) name10953 (
		_w8762_,
		_w8996_,
		_w12852_,
		_w12853_,
		_w12854_
	);
	LUT4 #(
		.INIT('h2a00)
	) name10954 (
		\s7_rty_i_pad ,
		_w8782_,
		_w8783_,
		_w9345_,
		_w12855_
	);
	LUT4 #(
		.INIT('h2a00)
	) name10955 (
		\s10_rty_i_pad ,
		_w8910_,
		_w8911_,
		_w9532_,
		_w12856_
	);
	LUT4 #(
		.INIT('h135f)
	) name10956 (
		_w8801_,
		_w8929_,
		_w12855_,
		_w12856_,
		_w12857_
	);
	LUT4 #(
		.INIT('h8000)
	) name10957 (
		_w12848_,
		_w12851_,
		_w12854_,
		_w12857_,
		_w12858_
	);
	LUT4 #(
		.INIT('h2a00)
	) name10958 (
		\s12_rty_i_pad ,
		_w9029_,
		_w9030_,
		_w9354_,
		_w12859_
	);
	LUT2 #(
		.INIT('h8)
	) name10959 (
		_w9042_,
		_w12859_,
		_w12860_
	);
	LUT4 #(
		.INIT('h2a00)
	) name10960 (
		\s11_rty_i_pad ,
		_w8955_,
		_w8956_,
		_w9535_,
		_w12861_
	);
	LUT4 #(
		.INIT('h2a00)
	) name10961 (
		\s4_rty_i_pad ,
		_w8655_,
		_w8656_,
		_w9544_,
		_w12862_
	);
	LUT4 #(
		.INIT('h153f)
	) name10962 (
		_w8654_,
		_w8954_,
		_w12861_,
		_w12862_,
		_w12863_
	);
	LUT4 #(
		.INIT('h2a00)
	) name10963 (
		\s3_rty_i_pad ,
		_w9205_,
		_w9206_,
		_w9351_,
		_w12864_
	);
	LUT4 #(
		.INIT('h2a00)
	) name10964 (
		\s5_rty_i_pad ,
		_w8699_,
		_w8700_,
		_w9547_,
		_w12865_
	);
	LUT4 #(
		.INIT('h153f)
	) name10965 (
		_w8706_,
		_w9204_,
		_w12864_,
		_w12865_,
		_w12866_
	);
	LUT4 #(
		.INIT('h2a00)
	) name10966 (
		\s2_rty_i_pad ,
		_w9171_,
		_w9172_,
		_w9541_,
		_w12867_
	);
	LUT4 #(
		.INIT('h2a00)
	) name10967 (
		\s8_rty_i_pad ,
		_w8821_,
		_w8822_,
		_w9553_,
		_w12868_
	);
	LUT4 #(
		.INIT('h153f)
	) name10968 (
		_w8840_,
		_w9170_,
		_w12867_,
		_w12868_,
		_w12869_
	);
	LUT4 #(
		.INIT('h4000)
	) name10969 (
		_w12860_,
		_w12863_,
		_w12866_,
		_w12869_,
		_w12870_
	);
	LUT2 #(
		.INIT('h8)
	) name10970 (
		_w12858_,
		_w12870_,
		_w12871_
	);
	LUT4 #(
		.INIT('h70ff)
	) name10971 (
		_w2046_,
		_w2097_,
		_w12845_,
		_w12871_,
		_w12872_
	);
	LUT3 #(
		.INIT('h70)
	) name10972 (
		_w1908_,
		_w1909_,
		_w2054_,
		_w12873_
	);
	LUT2 #(
		.INIT('h8)
	) name10973 (
		_w1907_,
		_w12873_,
		_w12874_
	);
	LUT3 #(
		.INIT('h70)
	) name10974 (
		_w2097_,
		_w8630_,
		_w12874_,
		_w12875_
	);
	LUT4 #(
		.INIT('h8000)
	) name10975 (
		\s5_ack_i_pad ,
		_w8699_,
		_w8700_,
		_w9585_,
		_w12876_
	);
	LUT4 #(
		.INIT('h8000)
	) name10976 (
		\s1_ack_i_pad ,
		_w9103_,
		_w9104_,
		_w9312_,
		_w12877_
	);
	LUT4 #(
		.INIT('h135f)
	) name10977 (
		_w8712_,
		_w9102_,
		_w12876_,
		_w12877_,
		_w12878_
	);
	LUT4 #(
		.INIT('h8000)
	) name10978 (
		\s8_ack_i_pad ,
		_w8821_,
		_w8822_,
		_w9342_,
		_w12879_
	);
	LUT4 #(
		.INIT('h8000)
	) name10979 (
		\s4_ack_i_pad ,
		_w8655_,
		_w8656_,
		_w9582_,
		_w12880_
	);
	LUT4 #(
		.INIT('h153f)
	) name10980 (
		_w8674_,
		_w8834_,
		_w12879_,
		_w12880_,
		_w12881_
	);
	LUT4 #(
		.INIT('h8000)
	) name10981 (
		\s6_ack_i_pad ,
		_w8743_,
		_w8744_,
		_w9336_,
		_w12882_
	);
	LUT4 #(
		.INIT('h8000)
	) name10982 (
		\s11_ack_i_pad ,
		_w8955_,
		_w8956_,
		_w9562_,
		_w12883_
	);
	LUT4 #(
		.INIT('h135f)
	) name10983 (
		_w8756_,
		_w8968_,
		_w12882_,
		_w12883_,
		_w12884_
	);
	LUT4 #(
		.INIT('h8000)
	) name10984 (
		\s0_ack_i_pad ,
		_w8989_,
		_w8990_,
		_w9308_,
		_w12885_
	);
	LUT4 #(
		.INIT('h8000)
	) name10985 (
		\s10_ack_i_pad ,
		_w8910_,
		_w8911_,
		_w9559_,
		_w12886_
	);
	LUT4 #(
		.INIT('h153f)
	) name10986 (
		_w8917_,
		_w8988_,
		_w12885_,
		_w12886_,
		_w12887_
	);
	LUT4 #(
		.INIT('h8000)
	) name10987 (
		_w12878_,
		_w12881_,
		_w12884_,
		_w12887_,
		_w12888_
	);
	LUT4 #(
		.INIT('h8000)
	) name10988 (
		\s3_ack_i_pad ,
		_w9205_,
		_w9206_,
		_w9579_,
		_w12889_
	);
	LUT2 #(
		.INIT('h8)
	) name10989 (
		_w9218_,
		_w12889_,
		_w12890_
	);
	LUT4 #(
		.INIT('h8000)
	) name10990 (
		\s14_ack_i_pad ,
		_w9137_,
		_w9138_,
		_w9571_,
		_w12891_
	);
	LUT4 #(
		.INIT('h8000)
	) name10991 (
		\s9_ack_i_pad ,
		_w8865_,
		_w8866_,
		_w9591_,
		_w12892_
	);
	LUT4 #(
		.INIT('h153f)
	) name10992 (
		_w8878_,
		_w9150_,
		_w12891_,
		_w12892_,
		_w12893_
	);
	LUT4 #(
		.INIT('h8000)
	) name10993 (
		\s7_ack_i_pad ,
		_w8782_,
		_w8783_,
		_w9588_,
		_w12894_
	);
	LUT4 #(
		.INIT('h8000)
	) name10994 (
		\s13_ack_i_pad ,
		_w9069_,
		_w9070_,
		_w9568_,
		_w12895_
	);
	LUT4 #(
		.INIT('h135f)
	) name10995 (
		_w8781_,
		_w9068_,
		_w12894_,
		_w12895_,
		_w12896_
	);
	LUT4 #(
		.INIT('h8000)
	) name10996 (
		\s2_ack_i_pad ,
		_w9171_,
		_w9172_,
		_w9576_,
		_w12897_
	);
	LUT4 #(
		.INIT('h8000)
	) name10997 (
		\s12_ack_i_pad ,
		_w9029_,
		_w9030_,
		_w9565_,
		_w12898_
	);
	LUT4 #(
		.INIT('h153f)
	) name10998 (
		_w9036_,
		_w9184_,
		_w12897_,
		_w12898_,
		_w12899_
	);
	LUT4 #(
		.INIT('h4000)
	) name10999 (
		_w12890_,
		_w12893_,
		_w12896_,
		_w12899_,
		_w12900_
	);
	LUT2 #(
		.INIT('h8)
	) name11000 (
		_w12888_,
		_w12900_,
		_w12901_
	);
	LUT3 #(
		.INIT('h4f)
	) name11001 (
		_w9652_,
		_w12875_,
		_w12901_,
		_w12902_
	);
	LUT3 #(
		.INIT('h80)
	) name11002 (
		_w2054_,
		_w2097_,
		_w9683_,
		_w12903_
	);
	LUT2 #(
		.INIT('h8)
	) name11003 (
		\s15_data_i[0]_pad ,
		_w2054_,
		_w12904_
	);
	LUT3 #(
		.INIT('h70)
	) name11004 (
		_w2046_,
		_w2097_,
		_w12904_,
		_w12905_
	);
	LUT4 #(
		.INIT('h153f)
	) name11005 (
		\s12_data_i[0]_pad ,
		\s1_data_i[0]_pad ,
		_w9312_,
		_w9565_,
		_w12906_
	);
	LUT4 #(
		.INIT('h135f)
	) name11006 (
		\s7_data_i[0]_pad ,
		\s9_data_i[0]_pad ,
		_w9588_,
		_w9591_,
		_w12907_
	);
	LUT4 #(
		.INIT('h153f)
	) name11007 (
		\s3_data_i[0]_pad ,
		\s6_data_i[0]_pad ,
		_w9336_,
		_w9579_,
		_w12908_
	);
	LUT4 #(
		.INIT('h135f)
	) name11008 (
		\s10_data_i[0]_pad ,
		\s13_data_i[0]_pad ,
		_w9559_,
		_w9568_,
		_w12909_
	);
	LUT4 #(
		.INIT('h8000)
	) name11009 (
		_w12906_,
		_w12907_,
		_w12908_,
		_w12909_,
		_w12910_
	);
	LUT2 #(
		.INIT('h8)
	) name11010 (
		\s14_data_i[0]_pad ,
		_w9571_,
		_w12911_
	);
	LUT4 #(
		.INIT('h135f)
	) name11011 (
		\s11_data_i[0]_pad ,
		\s2_data_i[0]_pad ,
		_w9562_,
		_w9576_,
		_w12912_
	);
	LUT4 #(
		.INIT('h153f)
	) name11012 (
		\s5_data_i[0]_pad ,
		\s8_data_i[0]_pad ,
		_w9342_,
		_w9585_,
		_w12913_
	);
	LUT4 #(
		.INIT('h135f)
	) name11013 (
		\s0_data_i[0]_pad ,
		\s4_data_i[0]_pad ,
		_w9308_,
		_w9582_,
		_w12914_
	);
	LUT4 #(
		.INIT('h4000)
	) name11014 (
		_w12911_,
		_w12912_,
		_w12913_,
		_w12914_,
		_w12915_
	);
	LUT2 #(
		.INIT('h8)
	) name11015 (
		_w12910_,
		_w12915_,
		_w12916_
	);
	LUT3 #(
		.INIT('hef)
	) name11016 (
		_w12903_,
		_w12905_,
		_w12916_,
		_w12917_
	);
	LUT3 #(
		.INIT('h80)
	) name11017 (
		_w2054_,
		_w2097_,
		_w9699_,
		_w12918_
	);
	LUT2 #(
		.INIT('h8)
	) name11018 (
		\s15_data_i[10]_pad ,
		_w2054_,
		_w12919_
	);
	LUT3 #(
		.INIT('h70)
	) name11019 (
		_w2046_,
		_w2097_,
		_w12919_,
		_w12920_
	);
	LUT4 #(
		.INIT('h153f)
	) name11020 (
		\s12_data_i[10]_pad ,
		\s1_data_i[10]_pad ,
		_w9312_,
		_w9565_,
		_w12921_
	);
	LUT4 #(
		.INIT('h153f)
	) name11021 (
		\s4_data_i[10]_pad ,
		\s6_data_i[10]_pad ,
		_w9336_,
		_w9582_,
		_w12922_
	);
	LUT4 #(
		.INIT('h135f)
	) name11022 (
		\s3_data_i[10]_pad ,
		\s9_data_i[10]_pad ,
		_w9579_,
		_w9591_,
		_w12923_
	);
	LUT4 #(
		.INIT('h135f)
	) name11023 (
		\s10_data_i[10]_pad ,
		\s7_data_i[10]_pad ,
		_w9559_,
		_w9588_,
		_w12924_
	);
	LUT4 #(
		.INIT('h8000)
	) name11024 (
		_w12921_,
		_w12922_,
		_w12923_,
		_w12924_,
		_w12925_
	);
	LUT2 #(
		.INIT('h8)
	) name11025 (
		\s14_data_i[10]_pad ,
		_w9571_,
		_w12926_
	);
	LUT4 #(
		.INIT('h135f)
	) name11026 (
		\s11_data_i[10]_pad ,
		\s2_data_i[10]_pad ,
		_w9562_,
		_w9576_,
		_w12927_
	);
	LUT4 #(
		.INIT('h153f)
	) name11027 (
		\s5_data_i[10]_pad ,
		\s8_data_i[10]_pad ,
		_w9342_,
		_w9585_,
		_w12928_
	);
	LUT4 #(
		.INIT('h135f)
	) name11028 (
		\s0_data_i[10]_pad ,
		\s13_data_i[10]_pad ,
		_w9308_,
		_w9568_,
		_w12929_
	);
	LUT4 #(
		.INIT('h4000)
	) name11029 (
		_w12926_,
		_w12927_,
		_w12928_,
		_w12929_,
		_w12930_
	);
	LUT2 #(
		.INIT('h8)
	) name11030 (
		_w12925_,
		_w12930_,
		_w12931_
	);
	LUT3 #(
		.INIT('hef)
	) name11031 (
		_w12918_,
		_w12920_,
		_w12931_,
		_w12932_
	);
	LUT3 #(
		.INIT('h80)
	) name11032 (
		_w2054_,
		_w2097_,
		_w9715_,
		_w12933_
	);
	LUT2 #(
		.INIT('h8)
	) name11033 (
		\s15_data_i[11]_pad ,
		_w2054_,
		_w12934_
	);
	LUT3 #(
		.INIT('h70)
	) name11034 (
		_w2046_,
		_w2097_,
		_w12934_,
		_w12935_
	);
	LUT4 #(
		.INIT('h153f)
	) name11035 (
		\s12_data_i[11]_pad ,
		\s1_data_i[11]_pad ,
		_w9312_,
		_w9565_,
		_w12936_
	);
	LUT4 #(
		.INIT('h153f)
	) name11036 (
		\s4_data_i[11]_pad ,
		\s6_data_i[11]_pad ,
		_w9336_,
		_w9582_,
		_w12937_
	);
	LUT4 #(
		.INIT('h135f)
	) name11037 (
		\s3_data_i[11]_pad ,
		\s9_data_i[11]_pad ,
		_w9579_,
		_w9591_,
		_w12938_
	);
	LUT4 #(
		.INIT('h135f)
	) name11038 (
		\s10_data_i[11]_pad ,
		\s7_data_i[11]_pad ,
		_w9559_,
		_w9588_,
		_w12939_
	);
	LUT4 #(
		.INIT('h8000)
	) name11039 (
		_w12936_,
		_w12937_,
		_w12938_,
		_w12939_,
		_w12940_
	);
	LUT2 #(
		.INIT('h8)
	) name11040 (
		\s14_data_i[11]_pad ,
		_w9571_,
		_w12941_
	);
	LUT4 #(
		.INIT('h135f)
	) name11041 (
		\s11_data_i[11]_pad ,
		\s2_data_i[11]_pad ,
		_w9562_,
		_w9576_,
		_w12942_
	);
	LUT4 #(
		.INIT('h153f)
	) name11042 (
		\s5_data_i[11]_pad ,
		\s8_data_i[11]_pad ,
		_w9342_,
		_w9585_,
		_w12943_
	);
	LUT4 #(
		.INIT('h135f)
	) name11043 (
		\s0_data_i[11]_pad ,
		\s13_data_i[11]_pad ,
		_w9308_,
		_w9568_,
		_w12944_
	);
	LUT4 #(
		.INIT('h4000)
	) name11044 (
		_w12941_,
		_w12942_,
		_w12943_,
		_w12944_,
		_w12945_
	);
	LUT2 #(
		.INIT('h8)
	) name11045 (
		_w12940_,
		_w12945_,
		_w12946_
	);
	LUT3 #(
		.INIT('hef)
	) name11046 (
		_w12933_,
		_w12935_,
		_w12946_,
		_w12947_
	);
	LUT3 #(
		.INIT('h80)
	) name11047 (
		_w2054_,
		_w2097_,
		_w9731_,
		_w12948_
	);
	LUT2 #(
		.INIT('h8)
	) name11048 (
		\s15_data_i[12]_pad ,
		_w2054_,
		_w12949_
	);
	LUT3 #(
		.INIT('h70)
	) name11049 (
		_w2046_,
		_w2097_,
		_w12949_,
		_w12950_
	);
	LUT4 #(
		.INIT('h153f)
	) name11050 (
		\s12_data_i[12]_pad ,
		\s1_data_i[12]_pad ,
		_w9312_,
		_w9565_,
		_w12951_
	);
	LUT4 #(
		.INIT('h153f)
	) name11051 (
		\s4_data_i[12]_pad ,
		\s6_data_i[12]_pad ,
		_w9336_,
		_w9582_,
		_w12952_
	);
	LUT4 #(
		.INIT('h135f)
	) name11052 (
		\s3_data_i[12]_pad ,
		\s9_data_i[12]_pad ,
		_w9579_,
		_w9591_,
		_w12953_
	);
	LUT4 #(
		.INIT('h135f)
	) name11053 (
		\s10_data_i[12]_pad ,
		\s7_data_i[12]_pad ,
		_w9559_,
		_w9588_,
		_w12954_
	);
	LUT4 #(
		.INIT('h8000)
	) name11054 (
		_w12951_,
		_w12952_,
		_w12953_,
		_w12954_,
		_w12955_
	);
	LUT2 #(
		.INIT('h8)
	) name11055 (
		\s14_data_i[12]_pad ,
		_w9571_,
		_w12956_
	);
	LUT4 #(
		.INIT('h135f)
	) name11056 (
		\s11_data_i[12]_pad ,
		\s2_data_i[12]_pad ,
		_w9562_,
		_w9576_,
		_w12957_
	);
	LUT4 #(
		.INIT('h153f)
	) name11057 (
		\s5_data_i[12]_pad ,
		\s8_data_i[12]_pad ,
		_w9342_,
		_w9585_,
		_w12958_
	);
	LUT4 #(
		.INIT('h135f)
	) name11058 (
		\s0_data_i[12]_pad ,
		\s13_data_i[12]_pad ,
		_w9308_,
		_w9568_,
		_w12959_
	);
	LUT4 #(
		.INIT('h4000)
	) name11059 (
		_w12956_,
		_w12957_,
		_w12958_,
		_w12959_,
		_w12960_
	);
	LUT2 #(
		.INIT('h8)
	) name11060 (
		_w12955_,
		_w12960_,
		_w12961_
	);
	LUT3 #(
		.INIT('hef)
	) name11061 (
		_w12948_,
		_w12950_,
		_w12961_,
		_w12962_
	);
	LUT3 #(
		.INIT('h80)
	) name11062 (
		_w2054_,
		_w2097_,
		_w9747_,
		_w12963_
	);
	LUT2 #(
		.INIT('h8)
	) name11063 (
		\s15_data_i[13]_pad ,
		_w2054_,
		_w12964_
	);
	LUT3 #(
		.INIT('h70)
	) name11064 (
		_w2046_,
		_w2097_,
		_w12964_,
		_w12965_
	);
	LUT4 #(
		.INIT('h153f)
	) name11065 (
		\s12_data_i[13]_pad ,
		\s1_data_i[13]_pad ,
		_w9312_,
		_w9565_,
		_w12966_
	);
	LUT4 #(
		.INIT('h135f)
	) name11066 (
		\s0_data_i[13]_pad ,
		\s10_data_i[13]_pad ,
		_w9308_,
		_w9559_,
		_w12967_
	);
	LUT4 #(
		.INIT('h135f)
	) name11067 (
		\s3_data_i[13]_pad ,
		\s4_data_i[13]_pad ,
		_w9579_,
		_w9582_,
		_w12968_
	);
	LUT4 #(
		.INIT('h135f)
	) name11068 (
		\s6_data_i[13]_pad ,
		\s9_data_i[13]_pad ,
		_w9336_,
		_w9591_,
		_w12969_
	);
	LUT4 #(
		.INIT('h8000)
	) name11069 (
		_w12966_,
		_w12967_,
		_w12968_,
		_w12969_,
		_w12970_
	);
	LUT2 #(
		.INIT('h8)
	) name11070 (
		\s14_data_i[13]_pad ,
		_w9571_,
		_w12971_
	);
	LUT4 #(
		.INIT('h135f)
	) name11071 (
		\s11_data_i[13]_pad ,
		\s7_data_i[13]_pad ,
		_w9562_,
		_w9588_,
		_w12972_
	);
	LUT4 #(
		.INIT('h153f)
	) name11072 (
		\s5_data_i[13]_pad ,
		\s8_data_i[13]_pad ,
		_w9342_,
		_w9585_,
		_w12973_
	);
	LUT4 #(
		.INIT('h135f)
	) name11073 (
		\s13_data_i[13]_pad ,
		\s2_data_i[13]_pad ,
		_w9568_,
		_w9576_,
		_w12974_
	);
	LUT4 #(
		.INIT('h4000)
	) name11074 (
		_w12971_,
		_w12972_,
		_w12973_,
		_w12974_,
		_w12975_
	);
	LUT2 #(
		.INIT('h8)
	) name11075 (
		_w12970_,
		_w12975_,
		_w12976_
	);
	LUT3 #(
		.INIT('hef)
	) name11076 (
		_w12963_,
		_w12965_,
		_w12976_,
		_w12977_
	);
	LUT3 #(
		.INIT('h80)
	) name11077 (
		_w2054_,
		_w2097_,
		_w9763_,
		_w12978_
	);
	LUT2 #(
		.INIT('h8)
	) name11078 (
		\s15_data_i[14]_pad ,
		_w2054_,
		_w12979_
	);
	LUT3 #(
		.INIT('h70)
	) name11079 (
		_w2046_,
		_w2097_,
		_w12979_,
		_w12980_
	);
	LUT4 #(
		.INIT('h153f)
	) name11080 (
		\s12_data_i[14]_pad ,
		\s1_data_i[14]_pad ,
		_w9312_,
		_w9565_,
		_w12981_
	);
	LUT4 #(
		.INIT('h135f)
	) name11081 (
		\s0_data_i[14]_pad ,
		\s7_data_i[14]_pad ,
		_w9308_,
		_w9588_,
		_w12982_
	);
	LUT4 #(
		.INIT('h135f)
	) name11082 (
		\s3_data_i[14]_pad ,
		\s9_data_i[14]_pad ,
		_w9579_,
		_w9591_,
		_w12983_
	);
	LUT4 #(
		.INIT('h135f)
	) name11083 (
		\s10_data_i[14]_pad ,
		\s4_data_i[14]_pad ,
		_w9559_,
		_w9582_,
		_w12984_
	);
	LUT4 #(
		.INIT('h8000)
	) name11084 (
		_w12981_,
		_w12982_,
		_w12983_,
		_w12984_,
		_w12985_
	);
	LUT2 #(
		.INIT('h8)
	) name11085 (
		\s14_data_i[14]_pad ,
		_w9571_,
		_w12986_
	);
	LUT4 #(
		.INIT('h135f)
	) name11086 (
		\s11_data_i[14]_pad ,
		\s2_data_i[14]_pad ,
		_w9562_,
		_w9576_,
		_w12987_
	);
	LUT4 #(
		.INIT('h153f)
	) name11087 (
		\s5_data_i[14]_pad ,
		\s8_data_i[14]_pad ,
		_w9342_,
		_w9585_,
		_w12988_
	);
	LUT4 #(
		.INIT('h153f)
	) name11088 (
		\s13_data_i[14]_pad ,
		\s6_data_i[14]_pad ,
		_w9336_,
		_w9568_,
		_w12989_
	);
	LUT4 #(
		.INIT('h4000)
	) name11089 (
		_w12986_,
		_w12987_,
		_w12988_,
		_w12989_,
		_w12990_
	);
	LUT2 #(
		.INIT('h8)
	) name11090 (
		_w12985_,
		_w12990_,
		_w12991_
	);
	LUT3 #(
		.INIT('hef)
	) name11091 (
		_w12978_,
		_w12980_,
		_w12991_,
		_w12992_
	);
	LUT3 #(
		.INIT('h80)
	) name11092 (
		_w2054_,
		_w2097_,
		_w9779_,
		_w12993_
	);
	LUT2 #(
		.INIT('h8)
	) name11093 (
		\s15_data_i[15]_pad ,
		_w2054_,
		_w12994_
	);
	LUT3 #(
		.INIT('h70)
	) name11094 (
		_w2046_,
		_w2097_,
		_w12994_,
		_w12995_
	);
	LUT4 #(
		.INIT('h153f)
	) name11095 (
		\s12_data_i[15]_pad ,
		\s1_data_i[15]_pad ,
		_w9312_,
		_w9565_,
		_w12996_
	);
	LUT4 #(
		.INIT('h135f)
	) name11096 (
		\s0_data_i[15]_pad ,
		\s10_data_i[15]_pad ,
		_w9308_,
		_w9559_,
		_w12997_
	);
	LUT4 #(
		.INIT('h135f)
	) name11097 (
		\s3_data_i[15]_pad ,
		\s4_data_i[15]_pad ,
		_w9579_,
		_w9582_,
		_w12998_
	);
	LUT4 #(
		.INIT('h135f)
	) name11098 (
		\s6_data_i[15]_pad ,
		\s9_data_i[15]_pad ,
		_w9336_,
		_w9591_,
		_w12999_
	);
	LUT4 #(
		.INIT('h8000)
	) name11099 (
		_w12996_,
		_w12997_,
		_w12998_,
		_w12999_,
		_w13000_
	);
	LUT2 #(
		.INIT('h8)
	) name11100 (
		\s14_data_i[15]_pad ,
		_w9571_,
		_w13001_
	);
	LUT4 #(
		.INIT('h135f)
	) name11101 (
		\s11_data_i[15]_pad ,
		\s7_data_i[15]_pad ,
		_w9562_,
		_w9588_,
		_w13002_
	);
	LUT4 #(
		.INIT('h153f)
	) name11102 (
		\s5_data_i[15]_pad ,
		\s8_data_i[15]_pad ,
		_w9342_,
		_w9585_,
		_w13003_
	);
	LUT4 #(
		.INIT('h135f)
	) name11103 (
		\s13_data_i[15]_pad ,
		\s2_data_i[15]_pad ,
		_w9568_,
		_w9576_,
		_w13004_
	);
	LUT4 #(
		.INIT('h4000)
	) name11104 (
		_w13001_,
		_w13002_,
		_w13003_,
		_w13004_,
		_w13005_
	);
	LUT2 #(
		.INIT('h8)
	) name11105 (
		_w13000_,
		_w13005_,
		_w13006_
	);
	LUT3 #(
		.INIT('hef)
	) name11106 (
		_w12993_,
		_w12995_,
		_w13006_,
		_w13007_
	);
	LUT2 #(
		.INIT('h8)
	) name11107 (
		\s15_data_i[16]_pad ,
		_w2054_,
		_w13008_
	);
	LUT4 #(
		.INIT('h135f)
	) name11108 (
		\s1_data_i[16]_pad ,
		\s8_data_i[16]_pad ,
		_w9312_,
		_w9342_,
		_w13009_
	);
	LUT4 #(
		.INIT('h153f)
	) name11109 (
		\s4_data_i[16]_pad ,
		\s6_data_i[16]_pad ,
		_w9336_,
		_w9582_,
		_w13010_
	);
	LUT4 #(
		.INIT('h135f)
	) name11110 (
		\s3_data_i[16]_pad ,
		\s9_data_i[16]_pad ,
		_w9579_,
		_w9591_,
		_w13011_
	);
	LUT4 #(
		.INIT('h135f)
	) name11111 (
		\s10_data_i[16]_pad ,
		\s7_data_i[16]_pad ,
		_w9559_,
		_w9588_,
		_w13012_
	);
	LUT4 #(
		.INIT('h8000)
	) name11112 (
		_w13009_,
		_w13010_,
		_w13011_,
		_w13012_,
		_w13013_
	);
	LUT2 #(
		.INIT('h8)
	) name11113 (
		\s11_data_i[16]_pad ,
		_w9562_,
		_w13014_
	);
	LUT4 #(
		.INIT('h135f)
	) name11114 (
		\s14_data_i[16]_pad ,
		\s2_data_i[16]_pad ,
		_w9571_,
		_w9576_,
		_w13015_
	);
	LUT4 #(
		.INIT('h135f)
	) name11115 (
		\s12_data_i[16]_pad ,
		\s5_data_i[16]_pad ,
		_w9565_,
		_w9585_,
		_w13016_
	);
	LUT4 #(
		.INIT('h135f)
	) name11116 (
		\s0_data_i[16]_pad ,
		\s13_data_i[16]_pad ,
		_w9308_,
		_w9568_,
		_w13017_
	);
	LUT4 #(
		.INIT('h4000)
	) name11117 (
		_w13014_,
		_w13015_,
		_w13016_,
		_w13017_,
		_w13018_
	);
	LUT2 #(
		.INIT('h8)
	) name11118 (
		_w13013_,
		_w13018_,
		_w13019_
	);
	LUT4 #(
		.INIT('h70ff)
	) name11119 (
		_w2046_,
		_w2097_,
		_w13008_,
		_w13019_,
		_w13020_
	);
	LUT2 #(
		.INIT('h8)
	) name11120 (
		\s15_data_i[17]_pad ,
		_w2054_,
		_w13021_
	);
	LUT4 #(
		.INIT('h135f)
	) name11121 (
		\s1_data_i[17]_pad ,
		\s8_data_i[17]_pad ,
		_w9312_,
		_w9342_,
		_w13022_
	);
	LUT4 #(
		.INIT('h153f)
	) name11122 (
		\s4_data_i[17]_pad ,
		\s6_data_i[17]_pad ,
		_w9336_,
		_w9582_,
		_w13023_
	);
	LUT4 #(
		.INIT('h135f)
	) name11123 (
		\s3_data_i[17]_pad ,
		\s9_data_i[17]_pad ,
		_w9579_,
		_w9591_,
		_w13024_
	);
	LUT4 #(
		.INIT('h135f)
	) name11124 (
		\s10_data_i[17]_pad ,
		\s7_data_i[17]_pad ,
		_w9559_,
		_w9588_,
		_w13025_
	);
	LUT4 #(
		.INIT('h8000)
	) name11125 (
		_w13022_,
		_w13023_,
		_w13024_,
		_w13025_,
		_w13026_
	);
	LUT2 #(
		.INIT('h8)
	) name11126 (
		\s11_data_i[17]_pad ,
		_w9562_,
		_w13027_
	);
	LUT4 #(
		.INIT('h135f)
	) name11127 (
		\s14_data_i[17]_pad ,
		\s2_data_i[17]_pad ,
		_w9571_,
		_w9576_,
		_w13028_
	);
	LUT4 #(
		.INIT('h135f)
	) name11128 (
		\s12_data_i[17]_pad ,
		\s5_data_i[17]_pad ,
		_w9565_,
		_w9585_,
		_w13029_
	);
	LUT4 #(
		.INIT('h135f)
	) name11129 (
		\s0_data_i[17]_pad ,
		\s13_data_i[17]_pad ,
		_w9308_,
		_w9568_,
		_w13030_
	);
	LUT4 #(
		.INIT('h4000)
	) name11130 (
		_w13027_,
		_w13028_,
		_w13029_,
		_w13030_,
		_w13031_
	);
	LUT2 #(
		.INIT('h8)
	) name11131 (
		_w13026_,
		_w13031_,
		_w13032_
	);
	LUT4 #(
		.INIT('h70ff)
	) name11132 (
		_w2046_,
		_w2097_,
		_w13021_,
		_w13032_,
		_w13033_
	);
	LUT2 #(
		.INIT('h8)
	) name11133 (
		\s15_data_i[18]_pad ,
		_w2054_,
		_w13034_
	);
	LUT4 #(
		.INIT('h135f)
	) name11134 (
		\s1_data_i[18]_pad ,
		\s8_data_i[18]_pad ,
		_w9312_,
		_w9342_,
		_w13035_
	);
	LUT4 #(
		.INIT('h153f)
	) name11135 (
		\s4_data_i[18]_pad ,
		\s6_data_i[18]_pad ,
		_w9336_,
		_w9582_,
		_w13036_
	);
	LUT4 #(
		.INIT('h135f)
	) name11136 (
		\s3_data_i[18]_pad ,
		\s9_data_i[18]_pad ,
		_w9579_,
		_w9591_,
		_w13037_
	);
	LUT4 #(
		.INIT('h135f)
	) name11137 (
		\s10_data_i[18]_pad ,
		\s7_data_i[18]_pad ,
		_w9559_,
		_w9588_,
		_w13038_
	);
	LUT4 #(
		.INIT('h8000)
	) name11138 (
		_w13035_,
		_w13036_,
		_w13037_,
		_w13038_,
		_w13039_
	);
	LUT2 #(
		.INIT('h8)
	) name11139 (
		\s11_data_i[18]_pad ,
		_w9562_,
		_w13040_
	);
	LUT4 #(
		.INIT('h135f)
	) name11140 (
		\s14_data_i[18]_pad ,
		\s2_data_i[18]_pad ,
		_w9571_,
		_w9576_,
		_w13041_
	);
	LUT4 #(
		.INIT('h135f)
	) name11141 (
		\s12_data_i[18]_pad ,
		\s5_data_i[18]_pad ,
		_w9565_,
		_w9585_,
		_w13042_
	);
	LUT4 #(
		.INIT('h135f)
	) name11142 (
		\s0_data_i[18]_pad ,
		\s13_data_i[18]_pad ,
		_w9308_,
		_w9568_,
		_w13043_
	);
	LUT4 #(
		.INIT('h4000)
	) name11143 (
		_w13040_,
		_w13041_,
		_w13042_,
		_w13043_,
		_w13044_
	);
	LUT2 #(
		.INIT('h8)
	) name11144 (
		_w13039_,
		_w13044_,
		_w13045_
	);
	LUT4 #(
		.INIT('h70ff)
	) name11145 (
		_w2046_,
		_w2097_,
		_w13034_,
		_w13045_,
		_w13046_
	);
	LUT2 #(
		.INIT('h8)
	) name11146 (
		\s15_data_i[19]_pad ,
		_w2054_,
		_w13047_
	);
	LUT4 #(
		.INIT('h135f)
	) name11147 (
		\s1_data_i[19]_pad ,
		\s8_data_i[19]_pad ,
		_w9312_,
		_w9342_,
		_w13048_
	);
	LUT4 #(
		.INIT('h153f)
	) name11148 (
		\s4_data_i[19]_pad ,
		\s6_data_i[19]_pad ,
		_w9336_,
		_w9582_,
		_w13049_
	);
	LUT4 #(
		.INIT('h135f)
	) name11149 (
		\s3_data_i[19]_pad ,
		\s9_data_i[19]_pad ,
		_w9579_,
		_w9591_,
		_w13050_
	);
	LUT4 #(
		.INIT('h135f)
	) name11150 (
		\s10_data_i[19]_pad ,
		\s7_data_i[19]_pad ,
		_w9559_,
		_w9588_,
		_w13051_
	);
	LUT4 #(
		.INIT('h8000)
	) name11151 (
		_w13048_,
		_w13049_,
		_w13050_,
		_w13051_,
		_w13052_
	);
	LUT2 #(
		.INIT('h8)
	) name11152 (
		\s11_data_i[19]_pad ,
		_w9562_,
		_w13053_
	);
	LUT4 #(
		.INIT('h135f)
	) name11153 (
		\s14_data_i[19]_pad ,
		\s2_data_i[19]_pad ,
		_w9571_,
		_w9576_,
		_w13054_
	);
	LUT4 #(
		.INIT('h135f)
	) name11154 (
		\s12_data_i[19]_pad ,
		\s5_data_i[19]_pad ,
		_w9565_,
		_w9585_,
		_w13055_
	);
	LUT4 #(
		.INIT('h135f)
	) name11155 (
		\s0_data_i[19]_pad ,
		\s13_data_i[19]_pad ,
		_w9308_,
		_w9568_,
		_w13056_
	);
	LUT4 #(
		.INIT('h4000)
	) name11156 (
		_w13053_,
		_w13054_,
		_w13055_,
		_w13056_,
		_w13057_
	);
	LUT2 #(
		.INIT('h8)
	) name11157 (
		_w13052_,
		_w13057_,
		_w13058_
	);
	LUT4 #(
		.INIT('h70ff)
	) name11158 (
		_w2046_,
		_w2097_,
		_w13047_,
		_w13058_,
		_w13059_
	);
	LUT3 #(
		.INIT('h80)
	) name11159 (
		_w2054_,
		_w2097_,
		_w9847_,
		_w13060_
	);
	LUT2 #(
		.INIT('h8)
	) name11160 (
		\s15_data_i[1]_pad ,
		_w2054_,
		_w13061_
	);
	LUT3 #(
		.INIT('h70)
	) name11161 (
		_w2046_,
		_w2097_,
		_w13061_,
		_w13062_
	);
	LUT4 #(
		.INIT('h153f)
	) name11162 (
		\s12_data_i[1]_pad ,
		\s1_data_i[1]_pad ,
		_w9312_,
		_w9565_,
		_w13063_
	);
	LUT4 #(
		.INIT('h135f)
	) name11163 (
		\s0_data_i[1]_pad ,
		\s10_data_i[1]_pad ,
		_w9308_,
		_w9559_,
		_w13064_
	);
	LUT4 #(
		.INIT('h135f)
	) name11164 (
		\s3_data_i[1]_pad ,
		\s4_data_i[1]_pad ,
		_w9579_,
		_w9582_,
		_w13065_
	);
	LUT4 #(
		.INIT('h135f)
	) name11165 (
		\s6_data_i[1]_pad ,
		\s9_data_i[1]_pad ,
		_w9336_,
		_w9591_,
		_w13066_
	);
	LUT4 #(
		.INIT('h8000)
	) name11166 (
		_w13063_,
		_w13064_,
		_w13065_,
		_w13066_,
		_w13067_
	);
	LUT2 #(
		.INIT('h8)
	) name11167 (
		\s14_data_i[1]_pad ,
		_w9571_,
		_w13068_
	);
	LUT4 #(
		.INIT('h135f)
	) name11168 (
		\s11_data_i[1]_pad ,
		\s7_data_i[1]_pad ,
		_w9562_,
		_w9588_,
		_w13069_
	);
	LUT4 #(
		.INIT('h153f)
	) name11169 (
		\s5_data_i[1]_pad ,
		\s8_data_i[1]_pad ,
		_w9342_,
		_w9585_,
		_w13070_
	);
	LUT4 #(
		.INIT('h135f)
	) name11170 (
		\s13_data_i[1]_pad ,
		\s2_data_i[1]_pad ,
		_w9568_,
		_w9576_,
		_w13071_
	);
	LUT4 #(
		.INIT('h4000)
	) name11171 (
		_w13068_,
		_w13069_,
		_w13070_,
		_w13071_,
		_w13072_
	);
	LUT2 #(
		.INIT('h8)
	) name11172 (
		_w13067_,
		_w13072_,
		_w13073_
	);
	LUT3 #(
		.INIT('hef)
	) name11173 (
		_w13060_,
		_w13062_,
		_w13073_,
		_w13074_
	);
	LUT2 #(
		.INIT('h8)
	) name11174 (
		\s15_data_i[20]_pad ,
		_w2054_,
		_w13075_
	);
	LUT4 #(
		.INIT('h135f)
	) name11175 (
		\s1_data_i[20]_pad ,
		\s8_data_i[20]_pad ,
		_w9312_,
		_w9342_,
		_w13076_
	);
	LUT4 #(
		.INIT('h153f)
	) name11176 (
		\s4_data_i[20]_pad ,
		\s6_data_i[20]_pad ,
		_w9336_,
		_w9582_,
		_w13077_
	);
	LUT4 #(
		.INIT('h135f)
	) name11177 (
		\s3_data_i[20]_pad ,
		\s9_data_i[20]_pad ,
		_w9579_,
		_w9591_,
		_w13078_
	);
	LUT4 #(
		.INIT('h135f)
	) name11178 (
		\s10_data_i[20]_pad ,
		\s7_data_i[20]_pad ,
		_w9559_,
		_w9588_,
		_w13079_
	);
	LUT4 #(
		.INIT('h8000)
	) name11179 (
		_w13076_,
		_w13077_,
		_w13078_,
		_w13079_,
		_w13080_
	);
	LUT2 #(
		.INIT('h8)
	) name11180 (
		\s11_data_i[20]_pad ,
		_w9562_,
		_w13081_
	);
	LUT4 #(
		.INIT('h135f)
	) name11181 (
		\s14_data_i[20]_pad ,
		\s2_data_i[20]_pad ,
		_w9571_,
		_w9576_,
		_w13082_
	);
	LUT4 #(
		.INIT('h135f)
	) name11182 (
		\s12_data_i[20]_pad ,
		\s5_data_i[20]_pad ,
		_w9565_,
		_w9585_,
		_w13083_
	);
	LUT4 #(
		.INIT('h135f)
	) name11183 (
		\s0_data_i[20]_pad ,
		\s13_data_i[20]_pad ,
		_w9308_,
		_w9568_,
		_w13084_
	);
	LUT4 #(
		.INIT('h4000)
	) name11184 (
		_w13081_,
		_w13082_,
		_w13083_,
		_w13084_,
		_w13085_
	);
	LUT2 #(
		.INIT('h8)
	) name11185 (
		_w13080_,
		_w13085_,
		_w13086_
	);
	LUT4 #(
		.INIT('h70ff)
	) name11186 (
		_w2046_,
		_w2097_,
		_w13075_,
		_w13086_,
		_w13087_
	);
	LUT2 #(
		.INIT('h8)
	) name11187 (
		\s15_data_i[21]_pad ,
		_w2054_,
		_w13088_
	);
	LUT4 #(
		.INIT('h135f)
	) name11188 (
		\s1_data_i[21]_pad ,
		\s8_data_i[21]_pad ,
		_w9312_,
		_w9342_,
		_w13089_
	);
	LUT4 #(
		.INIT('h153f)
	) name11189 (
		\s4_data_i[21]_pad ,
		\s6_data_i[21]_pad ,
		_w9336_,
		_w9582_,
		_w13090_
	);
	LUT4 #(
		.INIT('h135f)
	) name11190 (
		\s3_data_i[21]_pad ,
		\s9_data_i[21]_pad ,
		_w9579_,
		_w9591_,
		_w13091_
	);
	LUT4 #(
		.INIT('h135f)
	) name11191 (
		\s10_data_i[21]_pad ,
		\s7_data_i[21]_pad ,
		_w9559_,
		_w9588_,
		_w13092_
	);
	LUT4 #(
		.INIT('h8000)
	) name11192 (
		_w13089_,
		_w13090_,
		_w13091_,
		_w13092_,
		_w13093_
	);
	LUT2 #(
		.INIT('h8)
	) name11193 (
		\s11_data_i[21]_pad ,
		_w9562_,
		_w13094_
	);
	LUT4 #(
		.INIT('h135f)
	) name11194 (
		\s14_data_i[21]_pad ,
		\s2_data_i[21]_pad ,
		_w9571_,
		_w9576_,
		_w13095_
	);
	LUT4 #(
		.INIT('h135f)
	) name11195 (
		\s12_data_i[21]_pad ,
		\s5_data_i[21]_pad ,
		_w9565_,
		_w9585_,
		_w13096_
	);
	LUT4 #(
		.INIT('h135f)
	) name11196 (
		\s0_data_i[21]_pad ,
		\s13_data_i[21]_pad ,
		_w9308_,
		_w9568_,
		_w13097_
	);
	LUT4 #(
		.INIT('h4000)
	) name11197 (
		_w13094_,
		_w13095_,
		_w13096_,
		_w13097_,
		_w13098_
	);
	LUT2 #(
		.INIT('h8)
	) name11198 (
		_w13093_,
		_w13098_,
		_w13099_
	);
	LUT4 #(
		.INIT('h70ff)
	) name11199 (
		_w2046_,
		_w2097_,
		_w13088_,
		_w13099_,
		_w13100_
	);
	LUT2 #(
		.INIT('h8)
	) name11200 (
		\s15_data_i[22]_pad ,
		_w2054_,
		_w13101_
	);
	LUT4 #(
		.INIT('h135f)
	) name11201 (
		\s1_data_i[22]_pad ,
		\s8_data_i[22]_pad ,
		_w9312_,
		_w9342_,
		_w13102_
	);
	LUT4 #(
		.INIT('h135f)
	) name11202 (
		\s0_data_i[22]_pad ,
		\s7_data_i[22]_pad ,
		_w9308_,
		_w9588_,
		_w13103_
	);
	LUT4 #(
		.INIT('h135f)
	) name11203 (
		\s3_data_i[22]_pad ,
		\s9_data_i[22]_pad ,
		_w9579_,
		_w9591_,
		_w13104_
	);
	LUT4 #(
		.INIT('h135f)
	) name11204 (
		\s10_data_i[22]_pad ,
		\s4_data_i[22]_pad ,
		_w9559_,
		_w9582_,
		_w13105_
	);
	LUT4 #(
		.INIT('h8000)
	) name11205 (
		_w13102_,
		_w13103_,
		_w13104_,
		_w13105_,
		_w13106_
	);
	LUT2 #(
		.INIT('h8)
	) name11206 (
		\s11_data_i[22]_pad ,
		_w9562_,
		_w13107_
	);
	LUT4 #(
		.INIT('h135f)
	) name11207 (
		\s14_data_i[22]_pad ,
		\s2_data_i[22]_pad ,
		_w9571_,
		_w9576_,
		_w13108_
	);
	LUT4 #(
		.INIT('h135f)
	) name11208 (
		\s12_data_i[22]_pad ,
		\s5_data_i[22]_pad ,
		_w9565_,
		_w9585_,
		_w13109_
	);
	LUT4 #(
		.INIT('h153f)
	) name11209 (
		\s13_data_i[22]_pad ,
		\s6_data_i[22]_pad ,
		_w9336_,
		_w9568_,
		_w13110_
	);
	LUT4 #(
		.INIT('h4000)
	) name11210 (
		_w13107_,
		_w13108_,
		_w13109_,
		_w13110_,
		_w13111_
	);
	LUT2 #(
		.INIT('h8)
	) name11211 (
		_w13106_,
		_w13111_,
		_w13112_
	);
	LUT4 #(
		.INIT('h70ff)
	) name11212 (
		_w2046_,
		_w2097_,
		_w13101_,
		_w13112_,
		_w13113_
	);
	LUT2 #(
		.INIT('h8)
	) name11213 (
		\s15_data_i[23]_pad ,
		_w2054_,
		_w13114_
	);
	LUT4 #(
		.INIT('h135f)
	) name11214 (
		\s1_data_i[23]_pad ,
		\s8_data_i[23]_pad ,
		_w9312_,
		_w9342_,
		_w13115_
	);
	LUT4 #(
		.INIT('h153f)
	) name11215 (
		\s4_data_i[23]_pad ,
		\s6_data_i[23]_pad ,
		_w9336_,
		_w9582_,
		_w13116_
	);
	LUT4 #(
		.INIT('h135f)
	) name11216 (
		\s5_data_i[23]_pad ,
		\s9_data_i[23]_pad ,
		_w9585_,
		_w9591_,
		_w13117_
	);
	LUT4 #(
		.INIT('h135f)
	) name11217 (
		\s10_data_i[23]_pad ,
		\s7_data_i[23]_pad ,
		_w9559_,
		_w9588_,
		_w13118_
	);
	LUT4 #(
		.INIT('h8000)
	) name11218 (
		_w13115_,
		_w13116_,
		_w13117_,
		_w13118_,
		_w13119_
	);
	LUT2 #(
		.INIT('h8)
	) name11219 (
		\s11_data_i[23]_pad ,
		_w9562_,
		_w13120_
	);
	LUT4 #(
		.INIT('h135f)
	) name11220 (
		\s14_data_i[23]_pad ,
		\s3_data_i[23]_pad ,
		_w9571_,
		_w9579_,
		_w13121_
	);
	LUT4 #(
		.INIT('h135f)
	) name11221 (
		\s12_data_i[23]_pad ,
		\s2_data_i[23]_pad ,
		_w9565_,
		_w9576_,
		_w13122_
	);
	LUT4 #(
		.INIT('h135f)
	) name11222 (
		\s0_data_i[23]_pad ,
		\s13_data_i[23]_pad ,
		_w9308_,
		_w9568_,
		_w13123_
	);
	LUT4 #(
		.INIT('h4000)
	) name11223 (
		_w13120_,
		_w13121_,
		_w13122_,
		_w13123_,
		_w13124_
	);
	LUT2 #(
		.INIT('h8)
	) name11224 (
		_w13119_,
		_w13124_,
		_w13125_
	);
	LUT4 #(
		.INIT('h70ff)
	) name11225 (
		_w2046_,
		_w2097_,
		_w13114_,
		_w13125_,
		_w13126_
	);
	LUT2 #(
		.INIT('h8)
	) name11226 (
		\s15_data_i[24]_pad ,
		_w2054_,
		_w13127_
	);
	LUT4 #(
		.INIT('h135f)
	) name11227 (
		\s1_data_i[24]_pad ,
		\s8_data_i[24]_pad ,
		_w9312_,
		_w9342_,
		_w13128_
	);
	LUT4 #(
		.INIT('h153f)
	) name11228 (
		\s4_data_i[24]_pad ,
		\s6_data_i[24]_pad ,
		_w9336_,
		_w9582_,
		_w13129_
	);
	LUT4 #(
		.INIT('h135f)
	) name11229 (
		\s3_data_i[24]_pad ,
		\s9_data_i[24]_pad ,
		_w9579_,
		_w9591_,
		_w13130_
	);
	LUT4 #(
		.INIT('h135f)
	) name11230 (
		\s10_data_i[24]_pad ,
		\s7_data_i[24]_pad ,
		_w9559_,
		_w9588_,
		_w13131_
	);
	LUT4 #(
		.INIT('h8000)
	) name11231 (
		_w13128_,
		_w13129_,
		_w13130_,
		_w13131_,
		_w13132_
	);
	LUT2 #(
		.INIT('h8)
	) name11232 (
		\s11_data_i[24]_pad ,
		_w9562_,
		_w13133_
	);
	LUT4 #(
		.INIT('h135f)
	) name11233 (
		\s14_data_i[24]_pad ,
		\s2_data_i[24]_pad ,
		_w9571_,
		_w9576_,
		_w13134_
	);
	LUT4 #(
		.INIT('h135f)
	) name11234 (
		\s12_data_i[24]_pad ,
		\s5_data_i[24]_pad ,
		_w9565_,
		_w9585_,
		_w13135_
	);
	LUT4 #(
		.INIT('h135f)
	) name11235 (
		\s0_data_i[24]_pad ,
		\s13_data_i[24]_pad ,
		_w9308_,
		_w9568_,
		_w13136_
	);
	LUT4 #(
		.INIT('h4000)
	) name11236 (
		_w13133_,
		_w13134_,
		_w13135_,
		_w13136_,
		_w13137_
	);
	LUT2 #(
		.INIT('h8)
	) name11237 (
		_w13132_,
		_w13137_,
		_w13138_
	);
	LUT4 #(
		.INIT('h70ff)
	) name11238 (
		_w2046_,
		_w2097_,
		_w13127_,
		_w13138_,
		_w13139_
	);
	LUT2 #(
		.INIT('h8)
	) name11239 (
		\s15_data_i[25]_pad ,
		_w2054_,
		_w13140_
	);
	LUT4 #(
		.INIT('h135f)
	) name11240 (
		\s1_data_i[25]_pad ,
		\s8_data_i[25]_pad ,
		_w9312_,
		_w9342_,
		_w13141_
	);
	LUT4 #(
		.INIT('h153f)
	) name11241 (
		\s4_data_i[25]_pad ,
		\s6_data_i[25]_pad ,
		_w9336_,
		_w9582_,
		_w13142_
	);
	LUT4 #(
		.INIT('h135f)
	) name11242 (
		\s3_data_i[25]_pad ,
		\s9_data_i[25]_pad ,
		_w9579_,
		_w9591_,
		_w13143_
	);
	LUT4 #(
		.INIT('h135f)
	) name11243 (
		\s10_data_i[25]_pad ,
		\s7_data_i[25]_pad ,
		_w9559_,
		_w9588_,
		_w13144_
	);
	LUT4 #(
		.INIT('h8000)
	) name11244 (
		_w13141_,
		_w13142_,
		_w13143_,
		_w13144_,
		_w13145_
	);
	LUT2 #(
		.INIT('h8)
	) name11245 (
		\s11_data_i[25]_pad ,
		_w9562_,
		_w13146_
	);
	LUT4 #(
		.INIT('h135f)
	) name11246 (
		\s14_data_i[25]_pad ,
		\s2_data_i[25]_pad ,
		_w9571_,
		_w9576_,
		_w13147_
	);
	LUT4 #(
		.INIT('h135f)
	) name11247 (
		\s12_data_i[25]_pad ,
		\s5_data_i[25]_pad ,
		_w9565_,
		_w9585_,
		_w13148_
	);
	LUT4 #(
		.INIT('h135f)
	) name11248 (
		\s0_data_i[25]_pad ,
		\s13_data_i[25]_pad ,
		_w9308_,
		_w9568_,
		_w13149_
	);
	LUT4 #(
		.INIT('h4000)
	) name11249 (
		_w13146_,
		_w13147_,
		_w13148_,
		_w13149_,
		_w13150_
	);
	LUT2 #(
		.INIT('h8)
	) name11250 (
		_w13145_,
		_w13150_,
		_w13151_
	);
	LUT4 #(
		.INIT('h70ff)
	) name11251 (
		_w2046_,
		_w2097_,
		_w13140_,
		_w13151_,
		_w13152_
	);
	LUT2 #(
		.INIT('h8)
	) name11252 (
		\s15_data_i[26]_pad ,
		_w2054_,
		_w13153_
	);
	LUT4 #(
		.INIT('h135f)
	) name11253 (
		\s1_data_i[26]_pad ,
		\s8_data_i[26]_pad ,
		_w9312_,
		_w9342_,
		_w13154_
	);
	LUT4 #(
		.INIT('h153f)
	) name11254 (
		\s4_data_i[26]_pad ,
		\s6_data_i[26]_pad ,
		_w9336_,
		_w9582_,
		_w13155_
	);
	LUT4 #(
		.INIT('h135f)
	) name11255 (
		\s3_data_i[26]_pad ,
		\s9_data_i[26]_pad ,
		_w9579_,
		_w9591_,
		_w13156_
	);
	LUT4 #(
		.INIT('h135f)
	) name11256 (
		\s10_data_i[26]_pad ,
		\s7_data_i[26]_pad ,
		_w9559_,
		_w9588_,
		_w13157_
	);
	LUT4 #(
		.INIT('h8000)
	) name11257 (
		_w13154_,
		_w13155_,
		_w13156_,
		_w13157_,
		_w13158_
	);
	LUT2 #(
		.INIT('h8)
	) name11258 (
		\s11_data_i[26]_pad ,
		_w9562_,
		_w13159_
	);
	LUT4 #(
		.INIT('h135f)
	) name11259 (
		\s14_data_i[26]_pad ,
		\s2_data_i[26]_pad ,
		_w9571_,
		_w9576_,
		_w13160_
	);
	LUT4 #(
		.INIT('h135f)
	) name11260 (
		\s12_data_i[26]_pad ,
		\s5_data_i[26]_pad ,
		_w9565_,
		_w9585_,
		_w13161_
	);
	LUT4 #(
		.INIT('h135f)
	) name11261 (
		\s0_data_i[26]_pad ,
		\s13_data_i[26]_pad ,
		_w9308_,
		_w9568_,
		_w13162_
	);
	LUT4 #(
		.INIT('h4000)
	) name11262 (
		_w13159_,
		_w13160_,
		_w13161_,
		_w13162_,
		_w13163_
	);
	LUT2 #(
		.INIT('h8)
	) name11263 (
		_w13158_,
		_w13163_,
		_w13164_
	);
	LUT4 #(
		.INIT('h70ff)
	) name11264 (
		_w2046_,
		_w2097_,
		_w13153_,
		_w13164_,
		_w13165_
	);
	LUT2 #(
		.INIT('h8)
	) name11265 (
		\s15_data_i[27]_pad ,
		_w2054_,
		_w13166_
	);
	LUT4 #(
		.INIT('h135f)
	) name11266 (
		\s1_data_i[27]_pad ,
		\s8_data_i[27]_pad ,
		_w9312_,
		_w9342_,
		_w13167_
	);
	LUT4 #(
		.INIT('h153f)
	) name11267 (
		\s4_data_i[27]_pad ,
		\s6_data_i[27]_pad ,
		_w9336_,
		_w9582_,
		_w13168_
	);
	LUT4 #(
		.INIT('h135f)
	) name11268 (
		\s3_data_i[27]_pad ,
		\s9_data_i[27]_pad ,
		_w9579_,
		_w9591_,
		_w13169_
	);
	LUT4 #(
		.INIT('h135f)
	) name11269 (
		\s10_data_i[27]_pad ,
		\s7_data_i[27]_pad ,
		_w9559_,
		_w9588_,
		_w13170_
	);
	LUT4 #(
		.INIT('h8000)
	) name11270 (
		_w13167_,
		_w13168_,
		_w13169_,
		_w13170_,
		_w13171_
	);
	LUT2 #(
		.INIT('h8)
	) name11271 (
		\s11_data_i[27]_pad ,
		_w9562_,
		_w13172_
	);
	LUT4 #(
		.INIT('h135f)
	) name11272 (
		\s14_data_i[27]_pad ,
		\s2_data_i[27]_pad ,
		_w9571_,
		_w9576_,
		_w13173_
	);
	LUT4 #(
		.INIT('h135f)
	) name11273 (
		\s12_data_i[27]_pad ,
		\s5_data_i[27]_pad ,
		_w9565_,
		_w9585_,
		_w13174_
	);
	LUT4 #(
		.INIT('h135f)
	) name11274 (
		\s0_data_i[27]_pad ,
		\s13_data_i[27]_pad ,
		_w9308_,
		_w9568_,
		_w13175_
	);
	LUT4 #(
		.INIT('h4000)
	) name11275 (
		_w13172_,
		_w13173_,
		_w13174_,
		_w13175_,
		_w13176_
	);
	LUT2 #(
		.INIT('h8)
	) name11276 (
		_w13171_,
		_w13176_,
		_w13177_
	);
	LUT4 #(
		.INIT('h70ff)
	) name11277 (
		_w2046_,
		_w2097_,
		_w13166_,
		_w13177_,
		_w13178_
	);
	LUT2 #(
		.INIT('h8)
	) name11278 (
		\s15_data_i[28]_pad ,
		_w2054_,
		_w13179_
	);
	LUT4 #(
		.INIT('h135f)
	) name11279 (
		\s1_data_i[28]_pad ,
		\s8_data_i[28]_pad ,
		_w9312_,
		_w9342_,
		_w13180_
	);
	LUT4 #(
		.INIT('h153f)
	) name11280 (
		\s4_data_i[28]_pad ,
		\s6_data_i[28]_pad ,
		_w9336_,
		_w9582_,
		_w13181_
	);
	LUT4 #(
		.INIT('h135f)
	) name11281 (
		\s3_data_i[28]_pad ,
		\s9_data_i[28]_pad ,
		_w9579_,
		_w9591_,
		_w13182_
	);
	LUT4 #(
		.INIT('h135f)
	) name11282 (
		\s10_data_i[28]_pad ,
		\s7_data_i[28]_pad ,
		_w9559_,
		_w9588_,
		_w13183_
	);
	LUT4 #(
		.INIT('h8000)
	) name11283 (
		_w13180_,
		_w13181_,
		_w13182_,
		_w13183_,
		_w13184_
	);
	LUT2 #(
		.INIT('h8)
	) name11284 (
		\s11_data_i[28]_pad ,
		_w9562_,
		_w13185_
	);
	LUT4 #(
		.INIT('h135f)
	) name11285 (
		\s14_data_i[28]_pad ,
		\s2_data_i[28]_pad ,
		_w9571_,
		_w9576_,
		_w13186_
	);
	LUT4 #(
		.INIT('h135f)
	) name11286 (
		\s12_data_i[28]_pad ,
		\s5_data_i[28]_pad ,
		_w9565_,
		_w9585_,
		_w13187_
	);
	LUT4 #(
		.INIT('h135f)
	) name11287 (
		\s0_data_i[28]_pad ,
		\s13_data_i[28]_pad ,
		_w9308_,
		_w9568_,
		_w13188_
	);
	LUT4 #(
		.INIT('h4000)
	) name11288 (
		_w13185_,
		_w13186_,
		_w13187_,
		_w13188_,
		_w13189_
	);
	LUT2 #(
		.INIT('h8)
	) name11289 (
		_w13184_,
		_w13189_,
		_w13190_
	);
	LUT4 #(
		.INIT('h70ff)
	) name11290 (
		_w2046_,
		_w2097_,
		_w13179_,
		_w13190_,
		_w13191_
	);
	LUT2 #(
		.INIT('h8)
	) name11291 (
		\s15_data_i[29]_pad ,
		_w2054_,
		_w13192_
	);
	LUT4 #(
		.INIT('h135f)
	) name11292 (
		\s1_data_i[29]_pad ,
		\s8_data_i[29]_pad ,
		_w9312_,
		_w9342_,
		_w13193_
	);
	LUT4 #(
		.INIT('h153f)
	) name11293 (
		\s4_data_i[29]_pad ,
		\s6_data_i[29]_pad ,
		_w9336_,
		_w9582_,
		_w13194_
	);
	LUT4 #(
		.INIT('h135f)
	) name11294 (
		\s3_data_i[29]_pad ,
		\s9_data_i[29]_pad ,
		_w9579_,
		_w9591_,
		_w13195_
	);
	LUT4 #(
		.INIT('h135f)
	) name11295 (
		\s10_data_i[29]_pad ,
		\s7_data_i[29]_pad ,
		_w9559_,
		_w9588_,
		_w13196_
	);
	LUT4 #(
		.INIT('h8000)
	) name11296 (
		_w13193_,
		_w13194_,
		_w13195_,
		_w13196_,
		_w13197_
	);
	LUT2 #(
		.INIT('h8)
	) name11297 (
		\s11_data_i[29]_pad ,
		_w9562_,
		_w13198_
	);
	LUT4 #(
		.INIT('h135f)
	) name11298 (
		\s14_data_i[29]_pad ,
		\s2_data_i[29]_pad ,
		_w9571_,
		_w9576_,
		_w13199_
	);
	LUT4 #(
		.INIT('h135f)
	) name11299 (
		\s12_data_i[29]_pad ,
		\s5_data_i[29]_pad ,
		_w9565_,
		_w9585_,
		_w13200_
	);
	LUT4 #(
		.INIT('h135f)
	) name11300 (
		\s0_data_i[29]_pad ,
		\s13_data_i[29]_pad ,
		_w9308_,
		_w9568_,
		_w13201_
	);
	LUT4 #(
		.INIT('h4000)
	) name11301 (
		_w13198_,
		_w13199_,
		_w13200_,
		_w13201_,
		_w13202_
	);
	LUT2 #(
		.INIT('h8)
	) name11302 (
		_w13197_,
		_w13202_,
		_w13203_
	);
	LUT4 #(
		.INIT('h70ff)
	) name11303 (
		_w2046_,
		_w2097_,
		_w13192_,
		_w13203_,
		_w13204_
	);
	LUT3 #(
		.INIT('h80)
	) name11304 (
		_w2054_,
		_w2097_,
		_w9993_,
		_w13205_
	);
	LUT2 #(
		.INIT('h8)
	) name11305 (
		\s15_data_i[2]_pad ,
		_w2054_,
		_w13206_
	);
	LUT3 #(
		.INIT('h70)
	) name11306 (
		_w2046_,
		_w2097_,
		_w13206_,
		_w13207_
	);
	LUT4 #(
		.INIT('h153f)
	) name11307 (
		\s12_data_i[2]_pad ,
		\s1_data_i[2]_pad ,
		_w9312_,
		_w9565_,
		_w13208_
	);
	LUT4 #(
		.INIT('h135f)
	) name11308 (
		\s0_data_i[2]_pad ,
		\s10_data_i[2]_pad ,
		_w9308_,
		_w9559_,
		_w13209_
	);
	LUT4 #(
		.INIT('h135f)
	) name11309 (
		\s3_data_i[2]_pad ,
		\s4_data_i[2]_pad ,
		_w9579_,
		_w9582_,
		_w13210_
	);
	LUT4 #(
		.INIT('h135f)
	) name11310 (
		\s6_data_i[2]_pad ,
		\s9_data_i[2]_pad ,
		_w9336_,
		_w9591_,
		_w13211_
	);
	LUT4 #(
		.INIT('h8000)
	) name11311 (
		_w13208_,
		_w13209_,
		_w13210_,
		_w13211_,
		_w13212_
	);
	LUT2 #(
		.INIT('h8)
	) name11312 (
		\s14_data_i[2]_pad ,
		_w9571_,
		_w13213_
	);
	LUT4 #(
		.INIT('h135f)
	) name11313 (
		\s11_data_i[2]_pad ,
		\s7_data_i[2]_pad ,
		_w9562_,
		_w9588_,
		_w13214_
	);
	LUT4 #(
		.INIT('h153f)
	) name11314 (
		\s5_data_i[2]_pad ,
		\s8_data_i[2]_pad ,
		_w9342_,
		_w9585_,
		_w13215_
	);
	LUT4 #(
		.INIT('h135f)
	) name11315 (
		\s13_data_i[2]_pad ,
		\s2_data_i[2]_pad ,
		_w9568_,
		_w9576_,
		_w13216_
	);
	LUT4 #(
		.INIT('h4000)
	) name11316 (
		_w13213_,
		_w13214_,
		_w13215_,
		_w13216_,
		_w13217_
	);
	LUT2 #(
		.INIT('h8)
	) name11317 (
		_w13212_,
		_w13217_,
		_w13218_
	);
	LUT3 #(
		.INIT('hef)
	) name11318 (
		_w13205_,
		_w13207_,
		_w13218_,
		_w13219_
	);
	LUT2 #(
		.INIT('h8)
	) name11319 (
		\s15_data_i[30]_pad ,
		_w2054_,
		_w13220_
	);
	LUT4 #(
		.INIT('h135f)
	) name11320 (
		\s1_data_i[30]_pad ,
		\s8_data_i[30]_pad ,
		_w9312_,
		_w9342_,
		_w13221_
	);
	LUT4 #(
		.INIT('h153f)
	) name11321 (
		\s4_data_i[30]_pad ,
		\s6_data_i[30]_pad ,
		_w9336_,
		_w9582_,
		_w13222_
	);
	LUT4 #(
		.INIT('h135f)
	) name11322 (
		\s3_data_i[30]_pad ,
		\s9_data_i[30]_pad ,
		_w9579_,
		_w9591_,
		_w13223_
	);
	LUT4 #(
		.INIT('h135f)
	) name11323 (
		\s10_data_i[30]_pad ,
		\s7_data_i[30]_pad ,
		_w9559_,
		_w9588_,
		_w13224_
	);
	LUT4 #(
		.INIT('h8000)
	) name11324 (
		_w13221_,
		_w13222_,
		_w13223_,
		_w13224_,
		_w13225_
	);
	LUT2 #(
		.INIT('h8)
	) name11325 (
		\s11_data_i[30]_pad ,
		_w9562_,
		_w13226_
	);
	LUT4 #(
		.INIT('h135f)
	) name11326 (
		\s14_data_i[30]_pad ,
		\s2_data_i[30]_pad ,
		_w9571_,
		_w9576_,
		_w13227_
	);
	LUT4 #(
		.INIT('h135f)
	) name11327 (
		\s12_data_i[30]_pad ,
		\s5_data_i[30]_pad ,
		_w9565_,
		_w9585_,
		_w13228_
	);
	LUT4 #(
		.INIT('h135f)
	) name11328 (
		\s0_data_i[30]_pad ,
		\s13_data_i[30]_pad ,
		_w9308_,
		_w9568_,
		_w13229_
	);
	LUT4 #(
		.INIT('h4000)
	) name11329 (
		_w13226_,
		_w13227_,
		_w13228_,
		_w13229_,
		_w13230_
	);
	LUT2 #(
		.INIT('h8)
	) name11330 (
		_w13225_,
		_w13230_,
		_w13231_
	);
	LUT4 #(
		.INIT('h70ff)
	) name11331 (
		_w2046_,
		_w2097_,
		_w13220_,
		_w13231_,
		_w13232_
	);
	LUT2 #(
		.INIT('h8)
	) name11332 (
		\s15_data_i[31]_pad ,
		_w2054_,
		_w13233_
	);
	LUT4 #(
		.INIT('h135f)
	) name11333 (
		\s1_data_i[31]_pad ,
		\s8_data_i[31]_pad ,
		_w9312_,
		_w9342_,
		_w13234_
	);
	LUT4 #(
		.INIT('h153f)
	) name11334 (
		\s4_data_i[31]_pad ,
		\s6_data_i[31]_pad ,
		_w9336_,
		_w9582_,
		_w13235_
	);
	LUT4 #(
		.INIT('h135f)
	) name11335 (
		\s3_data_i[31]_pad ,
		\s9_data_i[31]_pad ,
		_w9579_,
		_w9591_,
		_w13236_
	);
	LUT4 #(
		.INIT('h135f)
	) name11336 (
		\s10_data_i[31]_pad ,
		\s7_data_i[31]_pad ,
		_w9559_,
		_w9588_,
		_w13237_
	);
	LUT4 #(
		.INIT('h8000)
	) name11337 (
		_w13234_,
		_w13235_,
		_w13236_,
		_w13237_,
		_w13238_
	);
	LUT2 #(
		.INIT('h8)
	) name11338 (
		\s11_data_i[31]_pad ,
		_w9562_,
		_w13239_
	);
	LUT4 #(
		.INIT('h135f)
	) name11339 (
		\s14_data_i[31]_pad ,
		\s2_data_i[31]_pad ,
		_w9571_,
		_w9576_,
		_w13240_
	);
	LUT4 #(
		.INIT('h135f)
	) name11340 (
		\s12_data_i[31]_pad ,
		\s5_data_i[31]_pad ,
		_w9565_,
		_w9585_,
		_w13241_
	);
	LUT4 #(
		.INIT('h135f)
	) name11341 (
		\s0_data_i[31]_pad ,
		\s13_data_i[31]_pad ,
		_w9308_,
		_w9568_,
		_w13242_
	);
	LUT4 #(
		.INIT('h4000)
	) name11342 (
		_w13239_,
		_w13240_,
		_w13241_,
		_w13242_,
		_w13243_
	);
	LUT2 #(
		.INIT('h8)
	) name11343 (
		_w13238_,
		_w13243_,
		_w13244_
	);
	LUT4 #(
		.INIT('h70ff)
	) name11344 (
		_w2046_,
		_w2097_,
		_w13233_,
		_w13244_,
		_w13245_
	);
	LUT3 #(
		.INIT('h80)
	) name11345 (
		_w2054_,
		_w2097_,
		_w10035_,
		_w13246_
	);
	LUT2 #(
		.INIT('h8)
	) name11346 (
		\s15_data_i[3]_pad ,
		_w2054_,
		_w13247_
	);
	LUT3 #(
		.INIT('h70)
	) name11347 (
		_w2046_,
		_w2097_,
		_w13247_,
		_w13248_
	);
	LUT4 #(
		.INIT('h153f)
	) name11348 (
		\s12_data_i[3]_pad ,
		\s1_data_i[3]_pad ,
		_w9312_,
		_w9565_,
		_w13249_
	);
	LUT4 #(
		.INIT('h153f)
	) name11349 (
		\s4_data_i[3]_pad ,
		\s6_data_i[3]_pad ,
		_w9336_,
		_w9582_,
		_w13250_
	);
	LUT4 #(
		.INIT('h135f)
	) name11350 (
		\s3_data_i[3]_pad ,
		\s9_data_i[3]_pad ,
		_w9579_,
		_w9591_,
		_w13251_
	);
	LUT4 #(
		.INIT('h135f)
	) name11351 (
		\s10_data_i[3]_pad ,
		\s7_data_i[3]_pad ,
		_w9559_,
		_w9588_,
		_w13252_
	);
	LUT4 #(
		.INIT('h8000)
	) name11352 (
		_w13249_,
		_w13250_,
		_w13251_,
		_w13252_,
		_w13253_
	);
	LUT2 #(
		.INIT('h8)
	) name11353 (
		\s14_data_i[3]_pad ,
		_w9571_,
		_w13254_
	);
	LUT4 #(
		.INIT('h135f)
	) name11354 (
		\s11_data_i[3]_pad ,
		\s2_data_i[3]_pad ,
		_w9562_,
		_w9576_,
		_w13255_
	);
	LUT4 #(
		.INIT('h153f)
	) name11355 (
		\s5_data_i[3]_pad ,
		\s8_data_i[3]_pad ,
		_w9342_,
		_w9585_,
		_w13256_
	);
	LUT4 #(
		.INIT('h135f)
	) name11356 (
		\s0_data_i[3]_pad ,
		\s13_data_i[3]_pad ,
		_w9308_,
		_w9568_,
		_w13257_
	);
	LUT4 #(
		.INIT('h4000)
	) name11357 (
		_w13254_,
		_w13255_,
		_w13256_,
		_w13257_,
		_w13258_
	);
	LUT2 #(
		.INIT('h8)
	) name11358 (
		_w13253_,
		_w13258_,
		_w13259_
	);
	LUT3 #(
		.INIT('hef)
	) name11359 (
		_w13246_,
		_w13248_,
		_w13259_,
		_w13260_
	);
	LUT3 #(
		.INIT('h80)
	) name11360 (
		_w2054_,
		_w2097_,
		_w10051_,
		_w13261_
	);
	LUT2 #(
		.INIT('h8)
	) name11361 (
		\s15_data_i[4]_pad ,
		_w2054_,
		_w13262_
	);
	LUT3 #(
		.INIT('h70)
	) name11362 (
		_w2046_,
		_w2097_,
		_w13262_,
		_w13263_
	);
	LUT4 #(
		.INIT('h135f)
	) name11363 (
		\s1_data_i[4]_pad ,
		\s5_data_i[4]_pad ,
		_w9312_,
		_w9585_,
		_w13264_
	);
	LUT4 #(
		.INIT('h135f)
	) name11364 (
		\s14_data_i[4]_pad ,
		\s4_data_i[4]_pad ,
		_w9571_,
		_w9582_,
		_w13265_
	);
	LUT4 #(
		.INIT('h135f)
	) name11365 (
		\s6_data_i[4]_pad ,
		\s8_data_i[4]_pad ,
		_w9336_,
		_w9342_,
		_w13266_
	);
	LUT4 #(
		.INIT('h135f)
	) name11366 (
		\s12_data_i[4]_pad ,
		\s7_data_i[4]_pad ,
		_w9565_,
		_w9588_,
		_w13267_
	);
	LUT4 #(
		.INIT('h8000)
	) name11367 (
		_w13264_,
		_w13265_,
		_w13266_,
		_w13267_,
		_w13268_
	);
	LUT2 #(
		.INIT('h8)
	) name11368 (
		\s9_data_i[4]_pad ,
		_w9591_,
		_w13269_
	);
	LUT4 #(
		.INIT('h135f)
	) name11369 (
		\s2_data_i[4]_pad ,
		\s3_data_i[4]_pad ,
		_w9576_,
		_w9579_,
		_w13270_
	);
	LUT4 #(
		.INIT('h135f)
	) name11370 (
		\s10_data_i[4]_pad ,
		\s11_data_i[4]_pad ,
		_w9559_,
		_w9562_,
		_w13271_
	);
	LUT4 #(
		.INIT('h135f)
	) name11371 (
		\s0_data_i[4]_pad ,
		\s13_data_i[4]_pad ,
		_w9308_,
		_w9568_,
		_w13272_
	);
	LUT4 #(
		.INIT('h4000)
	) name11372 (
		_w13269_,
		_w13270_,
		_w13271_,
		_w13272_,
		_w13273_
	);
	LUT2 #(
		.INIT('h8)
	) name11373 (
		_w13268_,
		_w13273_,
		_w13274_
	);
	LUT3 #(
		.INIT('hef)
	) name11374 (
		_w13261_,
		_w13263_,
		_w13274_,
		_w13275_
	);
	LUT3 #(
		.INIT('h80)
	) name11375 (
		_w2054_,
		_w2097_,
		_w10067_,
		_w13276_
	);
	LUT2 #(
		.INIT('h8)
	) name11376 (
		\s15_data_i[5]_pad ,
		_w2054_,
		_w13277_
	);
	LUT3 #(
		.INIT('h70)
	) name11377 (
		_w2046_,
		_w2097_,
		_w13277_,
		_w13278_
	);
	LUT4 #(
		.INIT('h153f)
	) name11378 (
		\s12_data_i[5]_pad ,
		\s1_data_i[5]_pad ,
		_w9312_,
		_w9565_,
		_w13279_
	);
	LUT4 #(
		.INIT('h153f)
	) name11379 (
		\s4_data_i[5]_pad ,
		\s6_data_i[5]_pad ,
		_w9336_,
		_w9582_,
		_w13280_
	);
	LUT4 #(
		.INIT('h135f)
	) name11380 (
		\s3_data_i[5]_pad ,
		\s9_data_i[5]_pad ,
		_w9579_,
		_w9591_,
		_w13281_
	);
	LUT4 #(
		.INIT('h135f)
	) name11381 (
		\s10_data_i[5]_pad ,
		\s7_data_i[5]_pad ,
		_w9559_,
		_w9588_,
		_w13282_
	);
	LUT4 #(
		.INIT('h8000)
	) name11382 (
		_w13279_,
		_w13280_,
		_w13281_,
		_w13282_,
		_w13283_
	);
	LUT2 #(
		.INIT('h8)
	) name11383 (
		\s14_data_i[5]_pad ,
		_w9571_,
		_w13284_
	);
	LUT4 #(
		.INIT('h135f)
	) name11384 (
		\s11_data_i[5]_pad ,
		\s2_data_i[5]_pad ,
		_w9562_,
		_w9576_,
		_w13285_
	);
	LUT4 #(
		.INIT('h153f)
	) name11385 (
		\s5_data_i[5]_pad ,
		\s8_data_i[5]_pad ,
		_w9342_,
		_w9585_,
		_w13286_
	);
	LUT4 #(
		.INIT('h135f)
	) name11386 (
		\s0_data_i[5]_pad ,
		\s13_data_i[5]_pad ,
		_w9308_,
		_w9568_,
		_w13287_
	);
	LUT4 #(
		.INIT('h4000)
	) name11387 (
		_w13284_,
		_w13285_,
		_w13286_,
		_w13287_,
		_w13288_
	);
	LUT2 #(
		.INIT('h8)
	) name11388 (
		_w13283_,
		_w13288_,
		_w13289_
	);
	LUT3 #(
		.INIT('hef)
	) name11389 (
		_w13276_,
		_w13278_,
		_w13289_,
		_w13290_
	);
	LUT3 #(
		.INIT('h80)
	) name11390 (
		_w2054_,
		_w2097_,
		_w10083_,
		_w13291_
	);
	LUT2 #(
		.INIT('h8)
	) name11391 (
		\s15_data_i[6]_pad ,
		_w2054_,
		_w13292_
	);
	LUT3 #(
		.INIT('h70)
	) name11392 (
		_w2046_,
		_w2097_,
		_w13292_,
		_w13293_
	);
	LUT4 #(
		.INIT('h153f)
	) name11393 (
		\s12_data_i[6]_pad ,
		\s1_data_i[6]_pad ,
		_w9312_,
		_w9565_,
		_w13294_
	);
	LUT4 #(
		.INIT('h153f)
	) name11394 (
		\s4_data_i[6]_pad ,
		\s6_data_i[6]_pad ,
		_w9336_,
		_w9582_,
		_w13295_
	);
	LUT4 #(
		.INIT('h135f)
	) name11395 (
		\s3_data_i[6]_pad ,
		\s9_data_i[6]_pad ,
		_w9579_,
		_w9591_,
		_w13296_
	);
	LUT4 #(
		.INIT('h135f)
	) name11396 (
		\s10_data_i[6]_pad ,
		\s7_data_i[6]_pad ,
		_w9559_,
		_w9588_,
		_w13297_
	);
	LUT4 #(
		.INIT('h8000)
	) name11397 (
		_w13294_,
		_w13295_,
		_w13296_,
		_w13297_,
		_w13298_
	);
	LUT2 #(
		.INIT('h8)
	) name11398 (
		\s14_data_i[6]_pad ,
		_w9571_,
		_w13299_
	);
	LUT4 #(
		.INIT('h135f)
	) name11399 (
		\s11_data_i[6]_pad ,
		\s2_data_i[6]_pad ,
		_w9562_,
		_w9576_,
		_w13300_
	);
	LUT4 #(
		.INIT('h153f)
	) name11400 (
		\s5_data_i[6]_pad ,
		\s8_data_i[6]_pad ,
		_w9342_,
		_w9585_,
		_w13301_
	);
	LUT4 #(
		.INIT('h135f)
	) name11401 (
		\s0_data_i[6]_pad ,
		\s13_data_i[6]_pad ,
		_w9308_,
		_w9568_,
		_w13302_
	);
	LUT4 #(
		.INIT('h4000)
	) name11402 (
		_w13299_,
		_w13300_,
		_w13301_,
		_w13302_,
		_w13303_
	);
	LUT2 #(
		.INIT('h8)
	) name11403 (
		_w13298_,
		_w13303_,
		_w13304_
	);
	LUT3 #(
		.INIT('hef)
	) name11404 (
		_w13291_,
		_w13293_,
		_w13304_,
		_w13305_
	);
	LUT3 #(
		.INIT('h80)
	) name11405 (
		_w2054_,
		_w2097_,
		_w10099_,
		_w13306_
	);
	LUT2 #(
		.INIT('h8)
	) name11406 (
		\s15_data_i[7]_pad ,
		_w2054_,
		_w13307_
	);
	LUT3 #(
		.INIT('h70)
	) name11407 (
		_w2046_,
		_w2097_,
		_w13307_,
		_w13308_
	);
	LUT4 #(
		.INIT('h135f)
	) name11408 (
		\s1_data_i[7]_pad ,
		\s5_data_i[7]_pad ,
		_w9312_,
		_w9585_,
		_w13309_
	);
	LUT4 #(
		.INIT('h135f)
	) name11409 (
		\s14_data_i[7]_pad ,
		\s4_data_i[7]_pad ,
		_w9571_,
		_w9582_,
		_w13310_
	);
	LUT4 #(
		.INIT('h135f)
	) name11410 (
		\s6_data_i[7]_pad ,
		\s8_data_i[7]_pad ,
		_w9336_,
		_w9342_,
		_w13311_
	);
	LUT4 #(
		.INIT('h135f)
	) name11411 (
		\s12_data_i[7]_pad ,
		\s7_data_i[7]_pad ,
		_w9565_,
		_w9588_,
		_w13312_
	);
	LUT4 #(
		.INIT('h8000)
	) name11412 (
		_w13309_,
		_w13310_,
		_w13311_,
		_w13312_,
		_w13313_
	);
	LUT2 #(
		.INIT('h8)
	) name11413 (
		\s9_data_i[7]_pad ,
		_w9591_,
		_w13314_
	);
	LUT4 #(
		.INIT('h135f)
	) name11414 (
		\s2_data_i[7]_pad ,
		\s3_data_i[7]_pad ,
		_w9576_,
		_w9579_,
		_w13315_
	);
	LUT4 #(
		.INIT('h135f)
	) name11415 (
		\s10_data_i[7]_pad ,
		\s11_data_i[7]_pad ,
		_w9559_,
		_w9562_,
		_w13316_
	);
	LUT4 #(
		.INIT('h135f)
	) name11416 (
		\s0_data_i[7]_pad ,
		\s13_data_i[7]_pad ,
		_w9308_,
		_w9568_,
		_w13317_
	);
	LUT4 #(
		.INIT('h4000)
	) name11417 (
		_w13314_,
		_w13315_,
		_w13316_,
		_w13317_,
		_w13318_
	);
	LUT2 #(
		.INIT('h8)
	) name11418 (
		_w13313_,
		_w13318_,
		_w13319_
	);
	LUT3 #(
		.INIT('hef)
	) name11419 (
		_w13306_,
		_w13308_,
		_w13319_,
		_w13320_
	);
	LUT3 #(
		.INIT('h80)
	) name11420 (
		_w2054_,
		_w2097_,
		_w10115_,
		_w13321_
	);
	LUT2 #(
		.INIT('h8)
	) name11421 (
		\s15_data_i[8]_pad ,
		_w2054_,
		_w13322_
	);
	LUT3 #(
		.INIT('h70)
	) name11422 (
		_w2046_,
		_w2097_,
		_w13322_,
		_w13323_
	);
	LUT4 #(
		.INIT('h153f)
	) name11423 (
		\s12_data_i[8]_pad ,
		\s1_data_i[8]_pad ,
		_w9312_,
		_w9565_,
		_w13324_
	);
	LUT4 #(
		.INIT('h153f)
	) name11424 (
		\s4_data_i[8]_pad ,
		\s6_data_i[8]_pad ,
		_w9336_,
		_w9582_,
		_w13325_
	);
	LUT4 #(
		.INIT('h135f)
	) name11425 (
		\s3_data_i[8]_pad ,
		\s9_data_i[8]_pad ,
		_w9579_,
		_w9591_,
		_w13326_
	);
	LUT4 #(
		.INIT('h135f)
	) name11426 (
		\s10_data_i[8]_pad ,
		\s7_data_i[8]_pad ,
		_w9559_,
		_w9588_,
		_w13327_
	);
	LUT4 #(
		.INIT('h8000)
	) name11427 (
		_w13324_,
		_w13325_,
		_w13326_,
		_w13327_,
		_w13328_
	);
	LUT2 #(
		.INIT('h8)
	) name11428 (
		\s14_data_i[8]_pad ,
		_w9571_,
		_w13329_
	);
	LUT4 #(
		.INIT('h135f)
	) name11429 (
		\s11_data_i[8]_pad ,
		\s2_data_i[8]_pad ,
		_w9562_,
		_w9576_,
		_w13330_
	);
	LUT4 #(
		.INIT('h153f)
	) name11430 (
		\s5_data_i[8]_pad ,
		\s8_data_i[8]_pad ,
		_w9342_,
		_w9585_,
		_w13331_
	);
	LUT4 #(
		.INIT('h135f)
	) name11431 (
		\s0_data_i[8]_pad ,
		\s13_data_i[8]_pad ,
		_w9308_,
		_w9568_,
		_w13332_
	);
	LUT4 #(
		.INIT('h4000)
	) name11432 (
		_w13329_,
		_w13330_,
		_w13331_,
		_w13332_,
		_w13333_
	);
	LUT2 #(
		.INIT('h8)
	) name11433 (
		_w13328_,
		_w13333_,
		_w13334_
	);
	LUT3 #(
		.INIT('hef)
	) name11434 (
		_w13321_,
		_w13323_,
		_w13334_,
		_w13335_
	);
	LUT3 #(
		.INIT('h80)
	) name11435 (
		_w2054_,
		_w2097_,
		_w10131_,
		_w13336_
	);
	LUT2 #(
		.INIT('h8)
	) name11436 (
		\s15_data_i[9]_pad ,
		_w2054_,
		_w13337_
	);
	LUT3 #(
		.INIT('h70)
	) name11437 (
		_w2046_,
		_w2097_,
		_w13337_,
		_w13338_
	);
	LUT4 #(
		.INIT('h135f)
	) name11438 (
		\s1_data_i[9]_pad ,
		\s5_data_i[9]_pad ,
		_w9312_,
		_w9585_,
		_w13339_
	);
	LUT4 #(
		.INIT('h135f)
	) name11439 (
		\s14_data_i[9]_pad ,
		\s4_data_i[9]_pad ,
		_w9571_,
		_w9582_,
		_w13340_
	);
	LUT4 #(
		.INIT('h135f)
	) name11440 (
		\s6_data_i[9]_pad ,
		\s8_data_i[9]_pad ,
		_w9336_,
		_w9342_,
		_w13341_
	);
	LUT4 #(
		.INIT('h135f)
	) name11441 (
		\s12_data_i[9]_pad ,
		\s7_data_i[9]_pad ,
		_w9565_,
		_w9588_,
		_w13342_
	);
	LUT4 #(
		.INIT('h8000)
	) name11442 (
		_w13339_,
		_w13340_,
		_w13341_,
		_w13342_,
		_w13343_
	);
	LUT2 #(
		.INIT('h8)
	) name11443 (
		\s9_data_i[9]_pad ,
		_w9591_,
		_w13344_
	);
	LUT4 #(
		.INIT('h135f)
	) name11444 (
		\s2_data_i[9]_pad ,
		\s3_data_i[9]_pad ,
		_w9576_,
		_w9579_,
		_w13345_
	);
	LUT4 #(
		.INIT('h135f)
	) name11445 (
		\s10_data_i[9]_pad ,
		\s11_data_i[9]_pad ,
		_w9559_,
		_w9562_,
		_w13346_
	);
	LUT4 #(
		.INIT('h135f)
	) name11446 (
		\s0_data_i[9]_pad ,
		\s13_data_i[9]_pad ,
		_w9308_,
		_w9568_,
		_w13347_
	);
	LUT4 #(
		.INIT('h4000)
	) name11447 (
		_w13344_,
		_w13345_,
		_w13346_,
		_w13347_,
		_w13348_
	);
	LUT2 #(
		.INIT('h8)
	) name11448 (
		_w13343_,
		_w13348_,
		_w13349_
	);
	LUT3 #(
		.INIT('hef)
	) name11449 (
		_w13336_,
		_w13338_,
		_w13349_,
		_w13350_
	);
	LUT3 #(
		.INIT('h80)
	) name11450 (
		\s15_err_i_pad ,
		_w1907_,
		_w12873_,
		_w13351_
	);
	LUT4 #(
		.INIT('h8000)
	) name11451 (
		\s2_err_i_pad ,
		_w9171_,
		_w9172_,
		_w9576_,
		_w13352_
	);
	LUT4 #(
		.INIT('h8000)
	) name11452 (
		\s12_err_i_pad ,
		_w9029_,
		_w9030_,
		_w9565_,
		_w13353_
	);
	LUT4 #(
		.INIT('h153f)
	) name11453 (
		_w9036_,
		_w9184_,
		_w13352_,
		_w13353_,
		_w13354_
	);
	LUT4 #(
		.INIT('h8000)
	) name11454 (
		\s13_err_i_pad ,
		_w9069_,
		_w9070_,
		_w9568_,
		_w13355_
	);
	LUT4 #(
		.INIT('h8000)
	) name11455 (
		\s9_err_i_pad ,
		_w8865_,
		_w8866_,
		_w9591_,
		_w13356_
	);
	LUT4 #(
		.INIT('h153f)
	) name11456 (
		_w8878_,
		_w9068_,
		_w13355_,
		_w13356_,
		_w13357_
	);
	LUT4 #(
		.INIT('h8000)
	) name11457 (
		\s6_err_i_pad ,
		_w8743_,
		_w8744_,
		_w9336_,
		_w13358_
	);
	LUT4 #(
		.INIT('h8000)
	) name11458 (
		\s4_err_i_pad ,
		_w8655_,
		_w8656_,
		_w9582_,
		_w13359_
	);
	LUT4 #(
		.INIT('h153f)
	) name11459 (
		_w8674_,
		_w8756_,
		_w13358_,
		_w13359_,
		_w13360_
	);
	LUT4 #(
		.INIT('h8000)
	) name11460 (
		\s0_err_i_pad ,
		_w8989_,
		_w8990_,
		_w9308_,
		_w13361_
	);
	LUT4 #(
		.INIT('h8000)
	) name11461 (
		\s10_err_i_pad ,
		_w8910_,
		_w8911_,
		_w9559_,
		_w13362_
	);
	LUT4 #(
		.INIT('h153f)
	) name11462 (
		_w8917_,
		_w8988_,
		_w13361_,
		_w13362_,
		_w13363_
	);
	LUT4 #(
		.INIT('h8000)
	) name11463 (
		_w13354_,
		_w13357_,
		_w13360_,
		_w13363_,
		_w13364_
	);
	LUT4 #(
		.INIT('h8000)
	) name11464 (
		\s1_err_i_pad ,
		_w9103_,
		_w9104_,
		_w9312_,
		_w13365_
	);
	LUT2 #(
		.INIT('h8)
	) name11465 (
		_w9102_,
		_w13365_,
		_w13366_
	);
	LUT4 #(
		.INIT('h8000)
	) name11466 (
		\s11_err_i_pad ,
		_w8955_,
		_w8956_,
		_w9562_,
		_w13367_
	);
	LUT4 #(
		.INIT('h8000)
	) name11467 (
		\s7_err_i_pad ,
		_w8782_,
		_w8783_,
		_w9588_,
		_w13368_
	);
	LUT4 #(
		.INIT('h153f)
	) name11468 (
		_w8781_,
		_w8968_,
		_w13367_,
		_w13368_,
		_w13369_
	);
	LUT4 #(
		.INIT('h8000)
	) name11469 (
		\s3_err_i_pad ,
		_w9205_,
		_w9206_,
		_w9579_,
		_w13370_
	);
	LUT4 #(
		.INIT('h8000)
	) name11470 (
		\s5_err_i_pad ,
		_w8699_,
		_w8700_,
		_w9585_,
		_w13371_
	);
	LUT4 #(
		.INIT('h153f)
	) name11471 (
		_w8712_,
		_w9218_,
		_w13370_,
		_w13371_,
		_w13372_
	);
	LUT4 #(
		.INIT('h8000)
	) name11472 (
		\s14_err_i_pad ,
		_w9137_,
		_w9138_,
		_w9571_,
		_w13373_
	);
	LUT4 #(
		.INIT('h8000)
	) name11473 (
		\s8_err_i_pad ,
		_w8821_,
		_w8822_,
		_w9342_,
		_w13374_
	);
	LUT4 #(
		.INIT('h153f)
	) name11474 (
		_w8834_,
		_w9150_,
		_w13373_,
		_w13374_,
		_w13375_
	);
	LUT4 #(
		.INIT('h4000)
	) name11475 (
		_w13366_,
		_w13369_,
		_w13372_,
		_w13375_,
		_w13376_
	);
	LUT2 #(
		.INIT('h8)
	) name11476 (
		_w13364_,
		_w13376_,
		_w13377_
	);
	LUT4 #(
		.INIT('h70ff)
	) name11477 (
		_w2046_,
		_w2097_,
		_w13351_,
		_w13377_,
		_w13378_
	);
	LUT3 #(
		.INIT('h80)
	) name11478 (
		\s15_rty_i_pad ,
		_w1907_,
		_w12873_,
		_w13379_
	);
	LUT4 #(
		.INIT('h8000)
	) name11479 (
		\s2_rty_i_pad ,
		_w9171_,
		_w9172_,
		_w9576_,
		_w13380_
	);
	LUT4 #(
		.INIT('h8000)
	) name11480 (
		\s3_rty_i_pad ,
		_w9205_,
		_w9206_,
		_w9579_,
		_w13381_
	);
	LUT4 #(
		.INIT('h135f)
	) name11481 (
		_w9184_,
		_w9218_,
		_w13380_,
		_w13381_,
		_w13382_
	);
	LUT4 #(
		.INIT('h8000)
	) name11482 (
		\s13_rty_i_pad ,
		_w9069_,
		_w9070_,
		_w9568_,
		_w13383_
	);
	LUT4 #(
		.INIT('h8000)
	) name11483 (
		\s0_rty_i_pad ,
		_w8989_,
		_w8990_,
		_w9308_,
		_w13384_
	);
	LUT4 #(
		.INIT('h153f)
	) name11484 (
		_w8988_,
		_w9068_,
		_w13383_,
		_w13384_,
		_w13385_
	);
	LUT4 #(
		.INIT('h8000)
	) name11485 (
		\s6_rty_i_pad ,
		_w8743_,
		_w8744_,
		_w9336_,
		_w13386_
	);
	LUT4 #(
		.INIT('h8000)
	) name11486 (
		\s10_rty_i_pad ,
		_w8910_,
		_w8911_,
		_w9559_,
		_w13387_
	);
	LUT4 #(
		.INIT('h135f)
	) name11487 (
		_w8756_,
		_w8917_,
		_w13386_,
		_w13387_,
		_w13388_
	);
	LUT4 #(
		.INIT('h8000)
	) name11488 (
		\s9_rty_i_pad ,
		_w8865_,
		_w8866_,
		_w9591_,
		_w13389_
	);
	LUT4 #(
		.INIT('h8000)
	) name11489 (
		\s4_rty_i_pad ,
		_w8655_,
		_w8656_,
		_w9582_,
		_w13390_
	);
	LUT4 #(
		.INIT('h153f)
	) name11490 (
		_w8674_,
		_w8878_,
		_w13389_,
		_w13390_,
		_w13391_
	);
	LUT4 #(
		.INIT('h8000)
	) name11491 (
		_w13382_,
		_w13385_,
		_w13388_,
		_w13391_,
		_w13392_
	);
	LUT4 #(
		.INIT('h8000)
	) name11492 (
		\s1_rty_i_pad ,
		_w9103_,
		_w9104_,
		_w9312_,
		_w13393_
	);
	LUT2 #(
		.INIT('h8)
	) name11493 (
		_w9102_,
		_w13393_,
		_w13394_
	);
	LUT4 #(
		.INIT('h8000)
	) name11494 (
		\s14_rty_i_pad ,
		_w9137_,
		_w9138_,
		_w9571_,
		_w13395_
	);
	LUT4 #(
		.INIT('h8000)
	) name11495 (
		\s7_rty_i_pad ,
		_w8782_,
		_w8783_,
		_w9588_,
		_w13396_
	);
	LUT4 #(
		.INIT('h153f)
	) name11496 (
		_w8781_,
		_w9150_,
		_w13395_,
		_w13396_,
		_w13397_
	);
	LUT4 #(
		.INIT('h8000)
	) name11497 (
		\s8_rty_i_pad ,
		_w8821_,
		_w8822_,
		_w9342_,
		_w13398_
	);
	LUT4 #(
		.INIT('h8000)
	) name11498 (
		\s11_rty_i_pad ,
		_w8955_,
		_w8956_,
		_w9562_,
		_w13399_
	);
	LUT4 #(
		.INIT('h135f)
	) name11499 (
		_w8834_,
		_w8968_,
		_w13398_,
		_w13399_,
		_w13400_
	);
	LUT4 #(
		.INIT('h8000)
	) name11500 (
		\s5_rty_i_pad ,
		_w8699_,
		_w8700_,
		_w9585_,
		_w13401_
	);
	LUT4 #(
		.INIT('h8000)
	) name11501 (
		\s12_rty_i_pad ,
		_w9029_,
		_w9030_,
		_w9565_,
		_w13402_
	);
	LUT4 #(
		.INIT('h135f)
	) name11502 (
		_w8712_,
		_w9036_,
		_w13401_,
		_w13402_,
		_w13403_
	);
	LUT4 #(
		.INIT('h4000)
	) name11503 (
		_w13394_,
		_w13397_,
		_w13400_,
		_w13403_,
		_w13404_
	);
	LUT2 #(
		.INIT('h8)
	) name11504 (
		_w13392_,
		_w13404_,
		_w13405_
	);
	LUT4 #(
		.INIT('h70ff)
	) name11505 (
		_w2046_,
		_w2097_,
		_w13379_,
		_w13405_,
		_w13406_
	);
	LUT3 #(
		.INIT('h70)
	) name11506 (
		_w1901_,
		_w1902_,
		_w2052_,
		_w13407_
	);
	LUT2 #(
		.INIT('h8)
	) name11507 (
		_w1918_,
		_w13407_,
		_w13408_
	);
	LUT3 #(
		.INIT('h70)
	) name11508 (
		_w2097_,
		_w8630_,
		_w13408_,
		_w13409_
	);
	LUT4 #(
		.INIT('h2a00)
	) name11509 (
		\s5_ack_i_pad ,
		_w8699_,
		_w8700_,
		_w9333_,
		_w13410_
	);
	LUT4 #(
		.INIT('h2a00)
	) name11510 (
		\s8_ack_i_pad ,
		_w8821_,
		_w8822_,
		_w9623_,
		_w13411_
	);
	LUT4 #(
		.INIT('h135f)
	) name11511 (
		_w8712_,
		_w8834_,
		_w13410_,
		_w13411_,
		_w13412_
	);
	LUT4 #(
		.INIT('h2a00)
	) name11512 (
		\s12_ack_i_pad ,
		_w9029_,
		_w9030_,
		_w9339_,
		_w13413_
	);
	LUT4 #(
		.INIT('h2a00)
	) name11513 (
		\s4_ack_i_pad ,
		_w8655_,
		_w8656_,
		_w9614_,
		_w13414_
	);
	LUT4 #(
		.INIT('h153f)
	) name11514 (
		_w8674_,
		_w9036_,
		_w13413_,
		_w13414_,
		_w13415_
	);
	LUT4 #(
		.INIT('h2a00)
	) name11515 (
		\s6_ack_i_pad ,
		_w8743_,
		_w8744_,
		_w9617_,
		_w13416_
	);
	LUT4 #(
		.INIT('h2a00)
	) name11516 (
		\s14_ack_i_pad ,
		_w9137_,
		_w9138_,
		_w9603_,
		_w13417_
	);
	LUT4 #(
		.INIT('h135f)
	) name11517 (
		_w8756_,
		_w9150_,
		_w13416_,
		_w13417_,
		_w13418_
	);
	LUT4 #(
		.INIT('h2a00)
	) name11518 (
		\s0_ack_i_pad ,
		_w8989_,
		_w8990_,
		_w9315_,
		_w13419_
	);
	LUT4 #(
		.INIT('h2a00)
	) name11519 (
		\s10_ack_i_pad ,
		_w8910_,
		_w8911_,
		_w9594_,
		_w13420_
	);
	LUT4 #(
		.INIT('h153f)
	) name11520 (
		_w8917_,
		_w8988_,
		_w13419_,
		_w13420_,
		_w13421_
	);
	LUT4 #(
		.INIT('h8000)
	) name11521 (
		_w13412_,
		_w13415_,
		_w13418_,
		_w13421_,
		_w13422_
	);
	LUT4 #(
		.INIT('h2a00)
	) name11522 (
		\s3_ack_i_pad ,
		_w9205_,
		_w9206_,
		_w9611_,
		_w13423_
	);
	LUT2 #(
		.INIT('h8)
	) name11523 (
		_w9218_,
		_w13423_,
		_w13424_
	);
	LUT4 #(
		.INIT('h2a00)
	) name11524 (
		\s2_ack_i_pad ,
		_w9171_,
		_w9172_,
		_w9608_,
		_w13425_
	);
	LUT4 #(
		.INIT('h2a00)
	) name11525 (
		\s9_ack_i_pad ,
		_w8865_,
		_w8866_,
		_w9327_,
		_w13426_
	);
	LUT4 #(
		.INIT('h153f)
	) name11526 (
		_w8878_,
		_w9184_,
		_w13425_,
		_w13426_,
		_w13427_
	);
	LUT4 #(
		.INIT('h2a00)
	) name11527 (
		\s7_ack_i_pad ,
		_w8782_,
		_w8783_,
		_w9330_,
		_w13428_
	);
	LUT4 #(
		.INIT('h2a00)
	) name11528 (
		\s13_ack_i_pad ,
		_w9069_,
		_w9070_,
		_w9600_,
		_w13429_
	);
	LUT4 #(
		.INIT('h135f)
	) name11529 (
		_w8781_,
		_w9068_,
		_w13428_,
		_w13429_,
		_w13430_
	);
	LUT4 #(
		.INIT('h2a00)
	) name11530 (
		\s11_ack_i_pad ,
		_w8955_,
		_w8956_,
		_w9597_,
		_w13431_
	);
	LUT4 #(
		.INIT('h2a00)
	) name11531 (
		\s1_ack_i_pad ,
		_w9103_,
		_w9104_,
		_w9319_,
		_w13432_
	);
	LUT4 #(
		.INIT('h135f)
	) name11532 (
		_w8968_,
		_w9102_,
		_w13431_,
		_w13432_,
		_w13433_
	);
	LUT4 #(
		.INIT('h4000)
	) name11533 (
		_w13424_,
		_w13427_,
		_w13430_,
		_w13433_,
		_w13434_
	);
	LUT2 #(
		.INIT('h8)
	) name11534 (
		_w13422_,
		_w13434_,
		_w13435_
	);
	LUT3 #(
		.INIT('h4f)
	) name11535 (
		_w9652_,
		_w13409_,
		_w13435_,
		_w13436_
	);
	LUT3 #(
		.INIT('h80)
	) name11536 (
		_w2052_,
		_w2097_,
		_w9683_,
		_w13437_
	);
	LUT2 #(
		.INIT('h8)
	) name11537 (
		\s15_data_i[0]_pad ,
		_w2052_,
		_w13438_
	);
	LUT3 #(
		.INIT('h70)
	) name11538 (
		_w2046_,
		_w2097_,
		_w13438_,
		_w13439_
	);
	LUT4 #(
		.INIT('h135f)
	) name11539 (
		\s1_data_i[0]_pad ,
		\s8_data_i[0]_pad ,
		_w9319_,
		_w9623_,
		_w13440_
	);
	LUT4 #(
		.INIT('h135f)
	) name11540 (
		\s4_data_i[0]_pad ,
		\s6_data_i[0]_pad ,
		_w9614_,
		_w9617_,
		_w13441_
	);
	LUT4 #(
		.INIT('h153f)
	) name11541 (
		\s5_data_i[0]_pad ,
		\s9_data_i[0]_pad ,
		_w9327_,
		_w9333_,
		_w13442_
	);
	LUT4 #(
		.INIT('h153f)
	) name11542 (
		\s10_data_i[0]_pad ,
		\s7_data_i[0]_pad ,
		_w9330_,
		_w9594_,
		_w13443_
	);
	LUT4 #(
		.INIT('h8000)
	) name11543 (
		_w13440_,
		_w13441_,
		_w13442_,
		_w13443_,
		_w13444_
	);
	LUT2 #(
		.INIT('h8)
	) name11544 (
		\s11_data_i[0]_pad ,
		_w9597_,
		_w13445_
	);
	LUT4 #(
		.INIT('h135f)
	) name11545 (
		\s13_data_i[0]_pad ,
		\s3_data_i[0]_pad ,
		_w9600_,
		_w9611_,
		_w13446_
	);
	LUT4 #(
		.INIT('h135f)
	) name11546 (
		\s12_data_i[0]_pad ,
		\s14_data_i[0]_pad ,
		_w9339_,
		_w9603_,
		_w13447_
	);
	LUT4 #(
		.INIT('h135f)
	) name11547 (
		\s0_data_i[0]_pad ,
		\s2_data_i[0]_pad ,
		_w9315_,
		_w9608_,
		_w13448_
	);
	LUT4 #(
		.INIT('h4000)
	) name11548 (
		_w13445_,
		_w13446_,
		_w13447_,
		_w13448_,
		_w13449_
	);
	LUT2 #(
		.INIT('h8)
	) name11549 (
		_w13444_,
		_w13449_,
		_w13450_
	);
	LUT3 #(
		.INIT('hef)
	) name11550 (
		_w13437_,
		_w13439_,
		_w13450_,
		_w13451_
	);
	LUT3 #(
		.INIT('h80)
	) name11551 (
		_w2052_,
		_w2097_,
		_w9699_,
		_w13452_
	);
	LUT2 #(
		.INIT('h8)
	) name11552 (
		\s15_data_i[10]_pad ,
		_w2052_,
		_w13453_
	);
	LUT3 #(
		.INIT('h70)
	) name11553 (
		_w2046_,
		_w2097_,
		_w13453_,
		_w13454_
	);
	LUT4 #(
		.INIT('h135f)
	) name11554 (
		\s1_data_i[10]_pad ,
		\s8_data_i[10]_pad ,
		_w9319_,
		_w9623_,
		_w13455_
	);
	LUT4 #(
		.INIT('h135f)
	) name11555 (
		\s4_data_i[10]_pad ,
		\s6_data_i[10]_pad ,
		_w9614_,
		_w9617_,
		_w13456_
	);
	LUT4 #(
		.INIT('h153f)
	) name11556 (
		\s5_data_i[10]_pad ,
		\s9_data_i[10]_pad ,
		_w9327_,
		_w9333_,
		_w13457_
	);
	LUT4 #(
		.INIT('h153f)
	) name11557 (
		\s10_data_i[10]_pad ,
		\s7_data_i[10]_pad ,
		_w9330_,
		_w9594_,
		_w13458_
	);
	LUT4 #(
		.INIT('h8000)
	) name11558 (
		_w13455_,
		_w13456_,
		_w13457_,
		_w13458_,
		_w13459_
	);
	LUT2 #(
		.INIT('h8)
	) name11559 (
		\s11_data_i[10]_pad ,
		_w9597_,
		_w13460_
	);
	LUT4 #(
		.INIT('h135f)
	) name11560 (
		\s13_data_i[10]_pad ,
		\s3_data_i[10]_pad ,
		_w9600_,
		_w9611_,
		_w13461_
	);
	LUT4 #(
		.INIT('h135f)
	) name11561 (
		\s12_data_i[10]_pad ,
		\s14_data_i[10]_pad ,
		_w9339_,
		_w9603_,
		_w13462_
	);
	LUT4 #(
		.INIT('h135f)
	) name11562 (
		\s0_data_i[10]_pad ,
		\s2_data_i[10]_pad ,
		_w9315_,
		_w9608_,
		_w13463_
	);
	LUT4 #(
		.INIT('h4000)
	) name11563 (
		_w13460_,
		_w13461_,
		_w13462_,
		_w13463_,
		_w13464_
	);
	LUT2 #(
		.INIT('h8)
	) name11564 (
		_w13459_,
		_w13464_,
		_w13465_
	);
	LUT3 #(
		.INIT('hef)
	) name11565 (
		_w13452_,
		_w13454_,
		_w13465_,
		_w13466_
	);
	LUT3 #(
		.INIT('h80)
	) name11566 (
		_w2052_,
		_w2097_,
		_w9715_,
		_w13467_
	);
	LUT2 #(
		.INIT('h8)
	) name11567 (
		\s15_data_i[11]_pad ,
		_w2052_,
		_w13468_
	);
	LUT3 #(
		.INIT('h70)
	) name11568 (
		_w2046_,
		_w2097_,
		_w13468_,
		_w13469_
	);
	LUT4 #(
		.INIT('h135f)
	) name11569 (
		\s1_data_i[11]_pad ,
		\s6_data_i[11]_pad ,
		_w9319_,
		_w9617_,
		_w13470_
	);
	LUT4 #(
		.INIT('h135f)
	) name11570 (
		\s14_data_i[11]_pad ,
		\s8_data_i[11]_pad ,
		_w9603_,
		_w9623_,
		_w13471_
	);
	LUT4 #(
		.INIT('h153f)
	) name11571 (
		\s11_data_i[11]_pad ,
		\s9_data_i[11]_pad ,
		_w9327_,
		_w9597_,
		_w13472_
	);
	LUT4 #(
		.INIT('h153f)
	) name11572 (
		\s12_data_i[11]_pad ,
		\s5_data_i[11]_pad ,
		_w9333_,
		_w9339_,
		_w13473_
	);
	LUT4 #(
		.INIT('h8000)
	) name11573 (
		_w13470_,
		_w13471_,
		_w13472_,
		_w13473_,
		_w13474_
	);
	LUT2 #(
		.INIT('h8)
	) name11574 (
		\s13_data_i[11]_pad ,
		_w9600_,
		_w13475_
	);
	LUT4 #(
		.INIT('h135f)
	) name11575 (
		\s0_data_i[11]_pad ,
		\s3_data_i[11]_pad ,
		_w9315_,
		_w9611_,
		_w13476_
	);
	LUT4 #(
		.INIT('h135f)
	) name11576 (
		\s10_data_i[11]_pad ,
		\s2_data_i[11]_pad ,
		_w9594_,
		_w9608_,
		_w13477_
	);
	LUT4 #(
		.INIT('h153f)
	) name11577 (
		\s4_data_i[11]_pad ,
		\s7_data_i[11]_pad ,
		_w9330_,
		_w9614_,
		_w13478_
	);
	LUT4 #(
		.INIT('h4000)
	) name11578 (
		_w13475_,
		_w13476_,
		_w13477_,
		_w13478_,
		_w13479_
	);
	LUT2 #(
		.INIT('h8)
	) name11579 (
		_w13474_,
		_w13479_,
		_w13480_
	);
	LUT3 #(
		.INIT('hef)
	) name11580 (
		_w13467_,
		_w13469_,
		_w13480_,
		_w13481_
	);
	LUT3 #(
		.INIT('h80)
	) name11581 (
		_w2052_,
		_w2097_,
		_w9731_,
		_w13482_
	);
	LUT2 #(
		.INIT('h8)
	) name11582 (
		\s15_data_i[12]_pad ,
		_w2052_,
		_w13483_
	);
	LUT3 #(
		.INIT('h70)
	) name11583 (
		_w2046_,
		_w2097_,
		_w13483_,
		_w13484_
	);
	LUT4 #(
		.INIT('h135f)
	) name11584 (
		\s1_data_i[12]_pad ,
		\s8_data_i[12]_pad ,
		_w9319_,
		_w9623_,
		_w13485_
	);
	LUT4 #(
		.INIT('h135f)
	) name11585 (
		\s4_data_i[12]_pad ,
		\s6_data_i[12]_pad ,
		_w9614_,
		_w9617_,
		_w13486_
	);
	LUT4 #(
		.INIT('h153f)
	) name11586 (
		\s5_data_i[12]_pad ,
		\s9_data_i[12]_pad ,
		_w9327_,
		_w9333_,
		_w13487_
	);
	LUT4 #(
		.INIT('h153f)
	) name11587 (
		\s10_data_i[12]_pad ,
		\s7_data_i[12]_pad ,
		_w9330_,
		_w9594_,
		_w13488_
	);
	LUT4 #(
		.INIT('h8000)
	) name11588 (
		_w13485_,
		_w13486_,
		_w13487_,
		_w13488_,
		_w13489_
	);
	LUT2 #(
		.INIT('h8)
	) name11589 (
		\s11_data_i[12]_pad ,
		_w9597_,
		_w13490_
	);
	LUT4 #(
		.INIT('h135f)
	) name11590 (
		\s13_data_i[12]_pad ,
		\s3_data_i[12]_pad ,
		_w9600_,
		_w9611_,
		_w13491_
	);
	LUT4 #(
		.INIT('h135f)
	) name11591 (
		\s12_data_i[12]_pad ,
		\s14_data_i[12]_pad ,
		_w9339_,
		_w9603_,
		_w13492_
	);
	LUT4 #(
		.INIT('h135f)
	) name11592 (
		\s0_data_i[12]_pad ,
		\s2_data_i[12]_pad ,
		_w9315_,
		_w9608_,
		_w13493_
	);
	LUT4 #(
		.INIT('h4000)
	) name11593 (
		_w13490_,
		_w13491_,
		_w13492_,
		_w13493_,
		_w13494_
	);
	LUT2 #(
		.INIT('h8)
	) name11594 (
		_w13489_,
		_w13494_,
		_w13495_
	);
	LUT3 #(
		.INIT('hef)
	) name11595 (
		_w13482_,
		_w13484_,
		_w13495_,
		_w13496_
	);
	LUT3 #(
		.INIT('h80)
	) name11596 (
		_w2052_,
		_w2097_,
		_w9747_,
		_w13497_
	);
	LUT2 #(
		.INIT('h8)
	) name11597 (
		\s15_data_i[13]_pad ,
		_w2052_,
		_w13498_
	);
	LUT3 #(
		.INIT('h70)
	) name11598 (
		_w2046_,
		_w2097_,
		_w13498_,
		_w13499_
	);
	LUT4 #(
		.INIT('h135f)
	) name11599 (
		\s1_data_i[13]_pad ,
		\s8_data_i[13]_pad ,
		_w9319_,
		_w9623_,
		_w13500_
	);
	LUT4 #(
		.INIT('h135f)
	) name11600 (
		\s4_data_i[13]_pad ,
		\s6_data_i[13]_pad ,
		_w9614_,
		_w9617_,
		_w13501_
	);
	LUT4 #(
		.INIT('h153f)
	) name11601 (
		\s5_data_i[13]_pad ,
		\s9_data_i[13]_pad ,
		_w9327_,
		_w9333_,
		_w13502_
	);
	LUT4 #(
		.INIT('h153f)
	) name11602 (
		\s10_data_i[13]_pad ,
		\s7_data_i[13]_pad ,
		_w9330_,
		_w9594_,
		_w13503_
	);
	LUT4 #(
		.INIT('h8000)
	) name11603 (
		_w13500_,
		_w13501_,
		_w13502_,
		_w13503_,
		_w13504_
	);
	LUT2 #(
		.INIT('h8)
	) name11604 (
		\s11_data_i[13]_pad ,
		_w9597_,
		_w13505_
	);
	LUT4 #(
		.INIT('h135f)
	) name11605 (
		\s13_data_i[13]_pad ,
		\s3_data_i[13]_pad ,
		_w9600_,
		_w9611_,
		_w13506_
	);
	LUT4 #(
		.INIT('h135f)
	) name11606 (
		\s12_data_i[13]_pad ,
		\s14_data_i[13]_pad ,
		_w9339_,
		_w9603_,
		_w13507_
	);
	LUT4 #(
		.INIT('h135f)
	) name11607 (
		\s0_data_i[13]_pad ,
		\s2_data_i[13]_pad ,
		_w9315_,
		_w9608_,
		_w13508_
	);
	LUT4 #(
		.INIT('h4000)
	) name11608 (
		_w13505_,
		_w13506_,
		_w13507_,
		_w13508_,
		_w13509_
	);
	LUT2 #(
		.INIT('h8)
	) name11609 (
		_w13504_,
		_w13509_,
		_w13510_
	);
	LUT3 #(
		.INIT('hef)
	) name11610 (
		_w13497_,
		_w13499_,
		_w13510_,
		_w13511_
	);
	LUT3 #(
		.INIT('h80)
	) name11611 (
		_w2052_,
		_w2097_,
		_w9763_,
		_w13512_
	);
	LUT2 #(
		.INIT('h8)
	) name11612 (
		\s15_data_i[14]_pad ,
		_w2052_,
		_w13513_
	);
	LUT3 #(
		.INIT('h70)
	) name11613 (
		_w2046_,
		_w2097_,
		_w13513_,
		_w13514_
	);
	LUT4 #(
		.INIT('h135f)
	) name11614 (
		\s1_data_i[14]_pad ,
		\s8_data_i[14]_pad ,
		_w9319_,
		_w9623_,
		_w13515_
	);
	LUT4 #(
		.INIT('h135f)
	) name11615 (
		\s4_data_i[14]_pad ,
		\s6_data_i[14]_pad ,
		_w9614_,
		_w9617_,
		_w13516_
	);
	LUT4 #(
		.INIT('h153f)
	) name11616 (
		\s5_data_i[14]_pad ,
		\s9_data_i[14]_pad ,
		_w9327_,
		_w9333_,
		_w13517_
	);
	LUT4 #(
		.INIT('h153f)
	) name11617 (
		\s10_data_i[14]_pad ,
		\s7_data_i[14]_pad ,
		_w9330_,
		_w9594_,
		_w13518_
	);
	LUT4 #(
		.INIT('h8000)
	) name11618 (
		_w13515_,
		_w13516_,
		_w13517_,
		_w13518_,
		_w13519_
	);
	LUT2 #(
		.INIT('h8)
	) name11619 (
		\s11_data_i[14]_pad ,
		_w9597_,
		_w13520_
	);
	LUT4 #(
		.INIT('h135f)
	) name11620 (
		\s13_data_i[14]_pad ,
		\s3_data_i[14]_pad ,
		_w9600_,
		_w9611_,
		_w13521_
	);
	LUT4 #(
		.INIT('h135f)
	) name11621 (
		\s12_data_i[14]_pad ,
		\s14_data_i[14]_pad ,
		_w9339_,
		_w9603_,
		_w13522_
	);
	LUT4 #(
		.INIT('h135f)
	) name11622 (
		\s0_data_i[14]_pad ,
		\s2_data_i[14]_pad ,
		_w9315_,
		_w9608_,
		_w13523_
	);
	LUT4 #(
		.INIT('h4000)
	) name11623 (
		_w13520_,
		_w13521_,
		_w13522_,
		_w13523_,
		_w13524_
	);
	LUT2 #(
		.INIT('h8)
	) name11624 (
		_w13519_,
		_w13524_,
		_w13525_
	);
	LUT3 #(
		.INIT('hef)
	) name11625 (
		_w13512_,
		_w13514_,
		_w13525_,
		_w13526_
	);
	LUT3 #(
		.INIT('h80)
	) name11626 (
		_w2052_,
		_w2097_,
		_w9779_,
		_w13527_
	);
	LUT2 #(
		.INIT('h8)
	) name11627 (
		\s15_data_i[15]_pad ,
		_w2052_,
		_w13528_
	);
	LUT3 #(
		.INIT('h70)
	) name11628 (
		_w2046_,
		_w2097_,
		_w13528_,
		_w13529_
	);
	LUT4 #(
		.INIT('h135f)
	) name11629 (
		\s1_data_i[15]_pad ,
		\s8_data_i[15]_pad ,
		_w9319_,
		_w9623_,
		_w13530_
	);
	LUT4 #(
		.INIT('h135f)
	) name11630 (
		\s4_data_i[15]_pad ,
		\s6_data_i[15]_pad ,
		_w9614_,
		_w9617_,
		_w13531_
	);
	LUT4 #(
		.INIT('h153f)
	) name11631 (
		\s5_data_i[15]_pad ,
		\s9_data_i[15]_pad ,
		_w9327_,
		_w9333_,
		_w13532_
	);
	LUT4 #(
		.INIT('h153f)
	) name11632 (
		\s10_data_i[15]_pad ,
		\s7_data_i[15]_pad ,
		_w9330_,
		_w9594_,
		_w13533_
	);
	LUT4 #(
		.INIT('h8000)
	) name11633 (
		_w13530_,
		_w13531_,
		_w13532_,
		_w13533_,
		_w13534_
	);
	LUT2 #(
		.INIT('h8)
	) name11634 (
		\s11_data_i[15]_pad ,
		_w9597_,
		_w13535_
	);
	LUT4 #(
		.INIT('h135f)
	) name11635 (
		\s13_data_i[15]_pad ,
		\s3_data_i[15]_pad ,
		_w9600_,
		_w9611_,
		_w13536_
	);
	LUT4 #(
		.INIT('h135f)
	) name11636 (
		\s12_data_i[15]_pad ,
		\s14_data_i[15]_pad ,
		_w9339_,
		_w9603_,
		_w13537_
	);
	LUT4 #(
		.INIT('h135f)
	) name11637 (
		\s0_data_i[15]_pad ,
		\s2_data_i[15]_pad ,
		_w9315_,
		_w9608_,
		_w13538_
	);
	LUT4 #(
		.INIT('h4000)
	) name11638 (
		_w13535_,
		_w13536_,
		_w13537_,
		_w13538_,
		_w13539_
	);
	LUT2 #(
		.INIT('h8)
	) name11639 (
		_w13534_,
		_w13539_,
		_w13540_
	);
	LUT3 #(
		.INIT('hef)
	) name11640 (
		_w13527_,
		_w13529_,
		_w13540_,
		_w13541_
	);
	LUT2 #(
		.INIT('h8)
	) name11641 (
		\s15_data_i[16]_pad ,
		_w2052_,
		_w13542_
	);
	LUT4 #(
		.INIT('h135f)
	) name11642 (
		\s12_data_i[16]_pad ,
		\s13_data_i[16]_pad ,
		_w9339_,
		_w9600_,
		_w13543_
	);
	LUT4 #(
		.INIT('h153f)
	) name11643 (
		\s10_data_i[16]_pad ,
		\s1_data_i[16]_pad ,
		_w9319_,
		_w9594_,
		_w13544_
	);
	LUT4 #(
		.INIT('h135f)
	) name11644 (
		\s5_data_i[16]_pad ,
		\s6_data_i[16]_pad ,
		_w9333_,
		_w9617_,
		_w13545_
	);
	LUT4 #(
		.INIT('h153f)
	) name11645 (
		\s2_data_i[16]_pad ,
		\s7_data_i[16]_pad ,
		_w9330_,
		_w9608_,
		_w13546_
	);
	LUT4 #(
		.INIT('h8000)
	) name11646 (
		_w13543_,
		_w13544_,
		_w13545_,
		_w13546_,
		_w13547_
	);
	LUT2 #(
		.INIT('h8)
	) name11647 (
		\s14_data_i[16]_pad ,
		_w9603_,
		_w13548_
	);
	LUT4 #(
		.INIT('h135f)
	) name11648 (
		\s3_data_i[16]_pad ,
		\s4_data_i[16]_pad ,
		_w9611_,
		_w9614_,
		_w13549_
	);
	LUT4 #(
		.INIT('h135f)
	) name11649 (
		\s11_data_i[16]_pad ,
		\s8_data_i[16]_pad ,
		_w9597_,
		_w9623_,
		_w13550_
	);
	LUT4 #(
		.INIT('h135f)
	) name11650 (
		\s0_data_i[16]_pad ,
		\s9_data_i[16]_pad ,
		_w9315_,
		_w9327_,
		_w13551_
	);
	LUT4 #(
		.INIT('h4000)
	) name11651 (
		_w13548_,
		_w13549_,
		_w13550_,
		_w13551_,
		_w13552_
	);
	LUT2 #(
		.INIT('h8)
	) name11652 (
		_w13547_,
		_w13552_,
		_w13553_
	);
	LUT4 #(
		.INIT('h70ff)
	) name11653 (
		_w2046_,
		_w2097_,
		_w13542_,
		_w13553_,
		_w13554_
	);
	LUT2 #(
		.INIT('h8)
	) name11654 (
		\s15_data_i[17]_pad ,
		_w2052_,
		_w13555_
	);
	LUT4 #(
		.INIT('h135f)
	) name11655 (
		\s12_data_i[17]_pad ,
		\s13_data_i[17]_pad ,
		_w9339_,
		_w9600_,
		_w13556_
	);
	LUT4 #(
		.INIT('h153f)
	) name11656 (
		\s10_data_i[17]_pad ,
		\s1_data_i[17]_pad ,
		_w9319_,
		_w9594_,
		_w13557_
	);
	LUT4 #(
		.INIT('h135f)
	) name11657 (
		\s5_data_i[17]_pad ,
		\s6_data_i[17]_pad ,
		_w9333_,
		_w9617_,
		_w13558_
	);
	LUT4 #(
		.INIT('h153f)
	) name11658 (
		\s2_data_i[17]_pad ,
		\s7_data_i[17]_pad ,
		_w9330_,
		_w9608_,
		_w13559_
	);
	LUT4 #(
		.INIT('h8000)
	) name11659 (
		_w13556_,
		_w13557_,
		_w13558_,
		_w13559_,
		_w13560_
	);
	LUT2 #(
		.INIT('h8)
	) name11660 (
		\s14_data_i[17]_pad ,
		_w9603_,
		_w13561_
	);
	LUT4 #(
		.INIT('h135f)
	) name11661 (
		\s3_data_i[17]_pad ,
		\s4_data_i[17]_pad ,
		_w9611_,
		_w9614_,
		_w13562_
	);
	LUT4 #(
		.INIT('h135f)
	) name11662 (
		\s11_data_i[17]_pad ,
		\s8_data_i[17]_pad ,
		_w9597_,
		_w9623_,
		_w13563_
	);
	LUT4 #(
		.INIT('h135f)
	) name11663 (
		\s0_data_i[17]_pad ,
		\s9_data_i[17]_pad ,
		_w9315_,
		_w9327_,
		_w13564_
	);
	LUT4 #(
		.INIT('h4000)
	) name11664 (
		_w13561_,
		_w13562_,
		_w13563_,
		_w13564_,
		_w13565_
	);
	LUT2 #(
		.INIT('h8)
	) name11665 (
		_w13560_,
		_w13565_,
		_w13566_
	);
	LUT4 #(
		.INIT('h70ff)
	) name11666 (
		_w2046_,
		_w2097_,
		_w13555_,
		_w13566_,
		_w13567_
	);
	LUT2 #(
		.INIT('h8)
	) name11667 (
		\s15_data_i[18]_pad ,
		_w2052_,
		_w13568_
	);
	LUT4 #(
		.INIT('h135f)
	) name11668 (
		\s12_data_i[18]_pad ,
		\s13_data_i[18]_pad ,
		_w9339_,
		_w9600_,
		_w13569_
	);
	LUT4 #(
		.INIT('h153f)
	) name11669 (
		\s10_data_i[18]_pad ,
		\s1_data_i[18]_pad ,
		_w9319_,
		_w9594_,
		_w13570_
	);
	LUT4 #(
		.INIT('h135f)
	) name11670 (
		\s5_data_i[18]_pad ,
		\s6_data_i[18]_pad ,
		_w9333_,
		_w9617_,
		_w13571_
	);
	LUT4 #(
		.INIT('h153f)
	) name11671 (
		\s2_data_i[18]_pad ,
		\s7_data_i[18]_pad ,
		_w9330_,
		_w9608_,
		_w13572_
	);
	LUT4 #(
		.INIT('h8000)
	) name11672 (
		_w13569_,
		_w13570_,
		_w13571_,
		_w13572_,
		_w13573_
	);
	LUT2 #(
		.INIT('h8)
	) name11673 (
		\s14_data_i[18]_pad ,
		_w9603_,
		_w13574_
	);
	LUT4 #(
		.INIT('h135f)
	) name11674 (
		\s3_data_i[18]_pad ,
		\s4_data_i[18]_pad ,
		_w9611_,
		_w9614_,
		_w13575_
	);
	LUT4 #(
		.INIT('h135f)
	) name11675 (
		\s11_data_i[18]_pad ,
		\s8_data_i[18]_pad ,
		_w9597_,
		_w9623_,
		_w13576_
	);
	LUT4 #(
		.INIT('h135f)
	) name11676 (
		\s0_data_i[18]_pad ,
		\s9_data_i[18]_pad ,
		_w9315_,
		_w9327_,
		_w13577_
	);
	LUT4 #(
		.INIT('h4000)
	) name11677 (
		_w13574_,
		_w13575_,
		_w13576_,
		_w13577_,
		_w13578_
	);
	LUT2 #(
		.INIT('h8)
	) name11678 (
		_w13573_,
		_w13578_,
		_w13579_
	);
	LUT4 #(
		.INIT('h70ff)
	) name11679 (
		_w2046_,
		_w2097_,
		_w13568_,
		_w13579_,
		_w13580_
	);
	LUT2 #(
		.INIT('h8)
	) name11680 (
		\s15_data_i[19]_pad ,
		_w2052_,
		_w13581_
	);
	LUT4 #(
		.INIT('h135f)
	) name11681 (
		\s12_data_i[19]_pad ,
		\s13_data_i[19]_pad ,
		_w9339_,
		_w9600_,
		_w13582_
	);
	LUT4 #(
		.INIT('h153f)
	) name11682 (
		\s10_data_i[19]_pad ,
		\s1_data_i[19]_pad ,
		_w9319_,
		_w9594_,
		_w13583_
	);
	LUT4 #(
		.INIT('h135f)
	) name11683 (
		\s5_data_i[19]_pad ,
		\s6_data_i[19]_pad ,
		_w9333_,
		_w9617_,
		_w13584_
	);
	LUT4 #(
		.INIT('h153f)
	) name11684 (
		\s2_data_i[19]_pad ,
		\s7_data_i[19]_pad ,
		_w9330_,
		_w9608_,
		_w13585_
	);
	LUT4 #(
		.INIT('h8000)
	) name11685 (
		_w13582_,
		_w13583_,
		_w13584_,
		_w13585_,
		_w13586_
	);
	LUT2 #(
		.INIT('h8)
	) name11686 (
		\s14_data_i[19]_pad ,
		_w9603_,
		_w13587_
	);
	LUT4 #(
		.INIT('h135f)
	) name11687 (
		\s3_data_i[19]_pad ,
		\s4_data_i[19]_pad ,
		_w9611_,
		_w9614_,
		_w13588_
	);
	LUT4 #(
		.INIT('h135f)
	) name11688 (
		\s11_data_i[19]_pad ,
		\s8_data_i[19]_pad ,
		_w9597_,
		_w9623_,
		_w13589_
	);
	LUT4 #(
		.INIT('h135f)
	) name11689 (
		\s0_data_i[19]_pad ,
		\s9_data_i[19]_pad ,
		_w9315_,
		_w9327_,
		_w13590_
	);
	LUT4 #(
		.INIT('h4000)
	) name11690 (
		_w13587_,
		_w13588_,
		_w13589_,
		_w13590_,
		_w13591_
	);
	LUT2 #(
		.INIT('h8)
	) name11691 (
		_w13586_,
		_w13591_,
		_w13592_
	);
	LUT4 #(
		.INIT('h70ff)
	) name11692 (
		_w2046_,
		_w2097_,
		_w13581_,
		_w13592_,
		_w13593_
	);
	LUT3 #(
		.INIT('h80)
	) name11693 (
		_w2052_,
		_w2097_,
		_w9847_,
		_w13594_
	);
	LUT2 #(
		.INIT('h8)
	) name11694 (
		\s15_data_i[1]_pad ,
		_w2052_,
		_w13595_
	);
	LUT3 #(
		.INIT('h70)
	) name11695 (
		_w2046_,
		_w2097_,
		_w13595_,
		_w13596_
	);
	LUT4 #(
		.INIT('h135f)
	) name11696 (
		\s1_data_i[1]_pad ,
		\s8_data_i[1]_pad ,
		_w9319_,
		_w9623_,
		_w13597_
	);
	LUT4 #(
		.INIT('h135f)
	) name11697 (
		\s4_data_i[1]_pad ,
		\s6_data_i[1]_pad ,
		_w9614_,
		_w9617_,
		_w13598_
	);
	LUT4 #(
		.INIT('h153f)
	) name11698 (
		\s5_data_i[1]_pad ,
		\s9_data_i[1]_pad ,
		_w9327_,
		_w9333_,
		_w13599_
	);
	LUT4 #(
		.INIT('h153f)
	) name11699 (
		\s10_data_i[1]_pad ,
		\s7_data_i[1]_pad ,
		_w9330_,
		_w9594_,
		_w13600_
	);
	LUT4 #(
		.INIT('h8000)
	) name11700 (
		_w13597_,
		_w13598_,
		_w13599_,
		_w13600_,
		_w13601_
	);
	LUT2 #(
		.INIT('h8)
	) name11701 (
		\s11_data_i[1]_pad ,
		_w9597_,
		_w13602_
	);
	LUT4 #(
		.INIT('h135f)
	) name11702 (
		\s13_data_i[1]_pad ,
		\s3_data_i[1]_pad ,
		_w9600_,
		_w9611_,
		_w13603_
	);
	LUT4 #(
		.INIT('h135f)
	) name11703 (
		\s12_data_i[1]_pad ,
		\s14_data_i[1]_pad ,
		_w9339_,
		_w9603_,
		_w13604_
	);
	LUT4 #(
		.INIT('h135f)
	) name11704 (
		\s0_data_i[1]_pad ,
		\s2_data_i[1]_pad ,
		_w9315_,
		_w9608_,
		_w13605_
	);
	LUT4 #(
		.INIT('h4000)
	) name11705 (
		_w13602_,
		_w13603_,
		_w13604_,
		_w13605_,
		_w13606_
	);
	LUT2 #(
		.INIT('h8)
	) name11706 (
		_w13601_,
		_w13606_,
		_w13607_
	);
	LUT3 #(
		.INIT('hef)
	) name11707 (
		_w13594_,
		_w13596_,
		_w13607_,
		_w13608_
	);
	LUT2 #(
		.INIT('h8)
	) name11708 (
		\s15_data_i[20]_pad ,
		_w2052_,
		_w13609_
	);
	LUT4 #(
		.INIT('h135f)
	) name11709 (
		\s12_data_i[20]_pad ,
		\s13_data_i[20]_pad ,
		_w9339_,
		_w9600_,
		_w13610_
	);
	LUT4 #(
		.INIT('h153f)
	) name11710 (
		\s10_data_i[20]_pad ,
		\s1_data_i[20]_pad ,
		_w9319_,
		_w9594_,
		_w13611_
	);
	LUT4 #(
		.INIT('h135f)
	) name11711 (
		\s5_data_i[20]_pad ,
		\s6_data_i[20]_pad ,
		_w9333_,
		_w9617_,
		_w13612_
	);
	LUT4 #(
		.INIT('h153f)
	) name11712 (
		\s2_data_i[20]_pad ,
		\s7_data_i[20]_pad ,
		_w9330_,
		_w9608_,
		_w13613_
	);
	LUT4 #(
		.INIT('h8000)
	) name11713 (
		_w13610_,
		_w13611_,
		_w13612_,
		_w13613_,
		_w13614_
	);
	LUT2 #(
		.INIT('h8)
	) name11714 (
		\s14_data_i[20]_pad ,
		_w9603_,
		_w13615_
	);
	LUT4 #(
		.INIT('h135f)
	) name11715 (
		\s3_data_i[20]_pad ,
		\s4_data_i[20]_pad ,
		_w9611_,
		_w9614_,
		_w13616_
	);
	LUT4 #(
		.INIT('h135f)
	) name11716 (
		\s11_data_i[20]_pad ,
		\s8_data_i[20]_pad ,
		_w9597_,
		_w9623_,
		_w13617_
	);
	LUT4 #(
		.INIT('h135f)
	) name11717 (
		\s0_data_i[20]_pad ,
		\s9_data_i[20]_pad ,
		_w9315_,
		_w9327_,
		_w13618_
	);
	LUT4 #(
		.INIT('h4000)
	) name11718 (
		_w13615_,
		_w13616_,
		_w13617_,
		_w13618_,
		_w13619_
	);
	LUT2 #(
		.INIT('h8)
	) name11719 (
		_w13614_,
		_w13619_,
		_w13620_
	);
	LUT4 #(
		.INIT('h70ff)
	) name11720 (
		_w2046_,
		_w2097_,
		_w13609_,
		_w13620_,
		_w13621_
	);
	LUT2 #(
		.INIT('h8)
	) name11721 (
		\s15_data_i[21]_pad ,
		_w2052_,
		_w13622_
	);
	LUT4 #(
		.INIT('h135f)
	) name11722 (
		\s12_data_i[21]_pad ,
		\s13_data_i[21]_pad ,
		_w9339_,
		_w9600_,
		_w13623_
	);
	LUT4 #(
		.INIT('h153f)
	) name11723 (
		\s10_data_i[21]_pad ,
		\s1_data_i[21]_pad ,
		_w9319_,
		_w9594_,
		_w13624_
	);
	LUT4 #(
		.INIT('h135f)
	) name11724 (
		\s5_data_i[21]_pad ,
		\s6_data_i[21]_pad ,
		_w9333_,
		_w9617_,
		_w13625_
	);
	LUT4 #(
		.INIT('h153f)
	) name11725 (
		\s2_data_i[21]_pad ,
		\s7_data_i[21]_pad ,
		_w9330_,
		_w9608_,
		_w13626_
	);
	LUT4 #(
		.INIT('h8000)
	) name11726 (
		_w13623_,
		_w13624_,
		_w13625_,
		_w13626_,
		_w13627_
	);
	LUT2 #(
		.INIT('h8)
	) name11727 (
		\s14_data_i[21]_pad ,
		_w9603_,
		_w13628_
	);
	LUT4 #(
		.INIT('h135f)
	) name11728 (
		\s3_data_i[21]_pad ,
		\s4_data_i[21]_pad ,
		_w9611_,
		_w9614_,
		_w13629_
	);
	LUT4 #(
		.INIT('h135f)
	) name11729 (
		\s11_data_i[21]_pad ,
		\s8_data_i[21]_pad ,
		_w9597_,
		_w9623_,
		_w13630_
	);
	LUT4 #(
		.INIT('h135f)
	) name11730 (
		\s0_data_i[21]_pad ,
		\s9_data_i[21]_pad ,
		_w9315_,
		_w9327_,
		_w13631_
	);
	LUT4 #(
		.INIT('h4000)
	) name11731 (
		_w13628_,
		_w13629_,
		_w13630_,
		_w13631_,
		_w13632_
	);
	LUT2 #(
		.INIT('h8)
	) name11732 (
		_w13627_,
		_w13632_,
		_w13633_
	);
	LUT4 #(
		.INIT('h70ff)
	) name11733 (
		_w2046_,
		_w2097_,
		_w13622_,
		_w13633_,
		_w13634_
	);
	LUT2 #(
		.INIT('h8)
	) name11734 (
		\s15_data_i[22]_pad ,
		_w2052_,
		_w13635_
	);
	LUT4 #(
		.INIT('h135f)
	) name11735 (
		\s12_data_i[22]_pad ,
		\s13_data_i[22]_pad ,
		_w9339_,
		_w9600_,
		_w13636_
	);
	LUT4 #(
		.INIT('h153f)
	) name11736 (
		\s10_data_i[22]_pad ,
		\s1_data_i[22]_pad ,
		_w9319_,
		_w9594_,
		_w13637_
	);
	LUT4 #(
		.INIT('h135f)
	) name11737 (
		\s5_data_i[22]_pad ,
		\s6_data_i[22]_pad ,
		_w9333_,
		_w9617_,
		_w13638_
	);
	LUT4 #(
		.INIT('h153f)
	) name11738 (
		\s2_data_i[22]_pad ,
		\s7_data_i[22]_pad ,
		_w9330_,
		_w9608_,
		_w13639_
	);
	LUT4 #(
		.INIT('h8000)
	) name11739 (
		_w13636_,
		_w13637_,
		_w13638_,
		_w13639_,
		_w13640_
	);
	LUT2 #(
		.INIT('h8)
	) name11740 (
		\s14_data_i[22]_pad ,
		_w9603_,
		_w13641_
	);
	LUT4 #(
		.INIT('h135f)
	) name11741 (
		\s3_data_i[22]_pad ,
		\s4_data_i[22]_pad ,
		_w9611_,
		_w9614_,
		_w13642_
	);
	LUT4 #(
		.INIT('h135f)
	) name11742 (
		\s11_data_i[22]_pad ,
		\s8_data_i[22]_pad ,
		_w9597_,
		_w9623_,
		_w13643_
	);
	LUT4 #(
		.INIT('h135f)
	) name11743 (
		\s0_data_i[22]_pad ,
		\s9_data_i[22]_pad ,
		_w9315_,
		_w9327_,
		_w13644_
	);
	LUT4 #(
		.INIT('h4000)
	) name11744 (
		_w13641_,
		_w13642_,
		_w13643_,
		_w13644_,
		_w13645_
	);
	LUT2 #(
		.INIT('h8)
	) name11745 (
		_w13640_,
		_w13645_,
		_w13646_
	);
	LUT4 #(
		.INIT('h70ff)
	) name11746 (
		_w2046_,
		_w2097_,
		_w13635_,
		_w13646_,
		_w13647_
	);
	LUT2 #(
		.INIT('h8)
	) name11747 (
		\s15_data_i[23]_pad ,
		_w2052_,
		_w13648_
	);
	LUT4 #(
		.INIT('h135f)
	) name11748 (
		\s12_data_i[23]_pad ,
		\s13_data_i[23]_pad ,
		_w9339_,
		_w9600_,
		_w13649_
	);
	LUT4 #(
		.INIT('h153f)
	) name11749 (
		\s10_data_i[23]_pad ,
		\s1_data_i[23]_pad ,
		_w9319_,
		_w9594_,
		_w13650_
	);
	LUT4 #(
		.INIT('h135f)
	) name11750 (
		\s5_data_i[23]_pad ,
		\s6_data_i[23]_pad ,
		_w9333_,
		_w9617_,
		_w13651_
	);
	LUT4 #(
		.INIT('h153f)
	) name11751 (
		\s2_data_i[23]_pad ,
		\s7_data_i[23]_pad ,
		_w9330_,
		_w9608_,
		_w13652_
	);
	LUT4 #(
		.INIT('h8000)
	) name11752 (
		_w13649_,
		_w13650_,
		_w13651_,
		_w13652_,
		_w13653_
	);
	LUT2 #(
		.INIT('h8)
	) name11753 (
		\s14_data_i[23]_pad ,
		_w9603_,
		_w13654_
	);
	LUT4 #(
		.INIT('h135f)
	) name11754 (
		\s3_data_i[23]_pad ,
		\s4_data_i[23]_pad ,
		_w9611_,
		_w9614_,
		_w13655_
	);
	LUT4 #(
		.INIT('h135f)
	) name11755 (
		\s11_data_i[23]_pad ,
		\s8_data_i[23]_pad ,
		_w9597_,
		_w9623_,
		_w13656_
	);
	LUT4 #(
		.INIT('h135f)
	) name11756 (
		\s0_data_i[23]_pad ,
		\s9_data_i[23]_pad ,
		_w9315_,
		_w9327_,
		_w13657_
	);
	LUT4 #(
		.INIT('h4000)
	) name11757 (
		_w13654_,
		_w13655_,
		_w13656_,
		_w13657_,
		_w13658_
	);
	LUT2 #(
		.INIT('h8)
	) name11758 (
		_w13653_,
		_w13658_,
		_w13659_
	);
	LUT4 #(
		.INIT('h70ff)
	) name11759 (
		_w2046_,
		_w2097_,
		_w13648_,
		_w13659_,
		_w13660_
	);
	LUT2 #(
		.INIT('h8)
	) name11760 (
		\s15_data_i[24]_pad ,
		_w2052_,
		_w13661_
	);
	LUT4 #(
		.INIT('h135f)
	) name11761 (
		\s12_data_i[24]_pad ,
		\s13_data_i[24]_pad ,
		_w9339_,
		_w9600_,
		_w13662_
	);
	LUT4 #(
		.INIT('h153f)
	) name11762 (
		\s10_data_i[24]_pad ,
		\s1_data_i[24]_pad ,
		_w9319_,
		_w9594_,
		_w13663_
	);
	LUT4 #(
		.INIT('h135f)
	) name11763 (
		\s5_data_i[24]_pad ,
		\s6_data_i[24]_pad ,
		_w9333_,
		_w9617_,
		_w13664_
	);
	LUT4 #(
		.INIT('h153f)
	) name11764 (
		\s2_data_i[24]_pad ,
		\s7_data_i[24]_pad ,
		_w9330_,
		_w9608_,
		_w13665_
	);
	LUT4 #(
		.INIT('h8000)
	) name11765 (
		_w13662_,
		_w13663_,
		_w13664_,
		_w13665_,
		_w13666_
	);
	LUT2 #(
		.INIT('h8)
	) name11766 (
		\s14_data_i[24]_pad ,
		_w9603_,
		_w13667_
	);
	LUT4 #(
		.INIT('h135f)
	) name11767 (
		\s3_data_i[24]_pad ,
		\s4_data_i[24]_pad ,
		_w9611_,
		_w9614_,
		_w13668_
	);
	LUT4 #(
		.INIT('h135f)
	) name11768 (
		\s11_data_i[24]_pad ,
		\s8_data_i[24]_pad ,
		_w9597_,
		_w9623_,
		_w13669_
	);
	LUT4 #(
		.INIT('h135f)
	) name11769 (
		\s0_data_i[24]_pad ,
		\s9_data_i[24]_pad ,
		_w9315_,
		_w9327_,
		_w13670_
	);
	LUT4 #(
		.INIT('h4000)
	) name11770 (
		_w13667_,
		_w13668_,
		_w13669_,
		_w13670_,
		_w13671_
	);
	LUT2 #(
		.INIT('h8)
	) name11771 (
		_w13666_,
		_w13671_,
		_w13672_
	);
	LUT4 #(
		.INIT('h70ff)
	) name11772 (
		_w2046_,
		_w2097_,
		_w13661_,
		_w13672_,
		_w13673_
	);
	LUT2 #(
		.INIT('h8)
	) name11773 (
		\s15_data_i[25]_pad ,
		_w2052_,
		_w13674_
	);
	LUT4 #(
		.INIT('h135f)
	) name11774 (
		\s12_data_i[25]_pad ,
		\s13_data_i[25]_pad ,
		_w9339_,
		_w9600_,
		_w13675_
	);
	LUT4 #(
		.INIT('h153f)
	) name11775 (
		\s10_data_i[25]_pad ,
		\s1_data_i[25]_pad ,
		_w9319_,
		_w9594_,
		_w13676_
	);
	LUT4 #(
		.INIT('h135f)
	) name11776 (
		\s5_data_i[25]_pad ,
		\s6_data_i[25]_pad ,
		_w9333_,
		_w9617_,
		_w13677_
	);
	LUT4 #(
		.INIT('h153f)
	) name11777 (
		\s2_data_i[25]_pad ,
		\s7_data_i[25]_pad ,
		_w9330_,
		_w9608_,
		_w13678_
	);
	LUT4 #(
		.INIT('h8000)
	) name11778 (
		_w13675_,
		_w13676_,
		_w13677_,
		_w13678_,
		_w13679_
	);
	LUT2 #(
		.INIT('h8)
	) name11779 (
		\s14_data_i[25]_pad ,
		_w9603_,
		_w13680_
	);
	LUT4 #(
		.INIT('h135f)
	) name11780 (
		\s3_data_i[25]_pad ,
		\s4_data_i[25]_pad ,
		_w9611_,
		_w9614_,
		_w13681_
	);
	LUT4 #(
		.INIT('h135f)
	) name11781 (
		\s11_data_i[25]_pad ,
		\s8_data_i[25]_pad ,
		_w9597_,
		_w9623_,
		_w13682_
	);
	LUT4 #(
		.INIT('h135f)
	) name11782 (
		\s0_data_i[25]_pad ,
		\s9_data_i[25]_pad ,
		_w9315_,
		_w9327_,
		_w13683_
	);
	LUT4 #(
		.INIT('h4000)
	) name11783 (
		_w13680_,
		_w13681_,
		_w13682_,
		_w13683_,
		_w13684_
	);
	LUT2 #(
		.INIT('h8)
	) name11784 (
		_w13679_,
		_w13684_,
		_w13685_
	);
	LUT4 #(
		.INIT('h70ff)
	) name11785 (
		_w2046_,
		_w2097_,
		_w13674_,
		_w13685_,
		_w13686_
	);
	LUT2 #(
		.INIT('h8)
	) name11786 (
		\s15_data_i[26]_pad ,
		_w2052_,
		_w13687_
	);
	LUT4 #(
		.INIT('h135f)
	) name11787 (
		\s12_data_i[26]_pad ,
		\s13_data_i[26]_pad ,
		_w9339_,
		_w9600_,
		_w13688_
	);
	LUT4 #(
		.INIT('h153f)
	) name11788 (
		\s10_data_i[26]_pad ,
		\s1_data_i[26]_pad ,
		_w9319_,
		_w9594_,
		_w13689_
	);
	LUT4 #(
		.INIT('h135f)
	) name11789 (
		\s5_data_i[26]_pad ,
		\s6_data_i[26]_pad ,
		_w9333_,
		_w9617_,
		_w13690_
	);
	LUT4 #(
		.INIT('h153f)
	) name11790 (
		\s2_data_i[26]_pad ,
		\s7_data_i[26]_pad ,
		_w9330_,
		_w9608_,
		_w13691_
	);
	LUT4 #(
		.INIT('h8000)
	) name11791 (
		_w13688_,
		_w13689_,
		_w13690_,
		_w13691_,
		_w13692_
	);
	LUT2 #(
		.INIT('h8)
	) name11792 (
		\s14_data_i[26]_pad ,
		_w9603_,
		_w13693_
	);
	LUT4 #(
		.INIT('h135f)
	) name11793 (
		\s3_data_i[26]_pad ,
		\s4_data_i[26]_pad ,
		_w9611_,
		_w9614_,
		_w13694_
	);
	LUT4 #(
		.INIT('h135f)
	) name11794 (
		\s11_data_i[26]_pad ,
		\s8_data_i[26]_pad ,
		_w9597_,
		_w9623_,
		_w13695_
	);
	LUT4 #(
		.INIT('h135f)
	) name11795 (
		\s0_data_i[26]_pad ,
		\s9_data_i[26]_pad ,
		_w9315_,
		_w9327_,
		_w13696_
	);
	LUT4 #(
		.INIT('h4000)
	) name11796 (
		_w13693_,
		_w13694_,
		_w13695_,
		_w13696_,
		_w13697_
	);
	LUT2 #(
		.INIT('h8)
	) name11797 (
		_w13692_,
		_w13697_,
		_w13698_
	);
	LUT4 #(
		.INIT('h70ff)
	) name11798 (
		_w2046_,
		_w2097_,
		_w13687_,
		_w13698_,
		_w13699_
	);
	LUT2 #(
		.INIT('h8)
	) name11799 (
		\s15_data_i[27]_pad ,
		_w2052_,
		_w13700_
	);
	LUT4 #(
		.INIT('h135f)
	) name11800 (
		\s12_data_i[27]_pad ,
		\s13_data_i[27]_pad ,
		_w9339_,
		_w9600_,
		_w13701_
	);
	LUT4 #(
		.INIT('h153f)
	) name11801 (
		\s10_data_i[27]_pad ,
		\s1_data_i[27]_pad ,
		_w9319_,
		_w9594_,
		_w13702_
	);
	LUT4 #(
		.INIT('h135f)
	) name11802 (
		\s5_data_i[27]_pad ,
		\s6_data_i[27]_pad ,
		_w9333_,
		_w9617_,
		_w13703_
	);
	LUT4 #(
		.INIT('h153f)
	) name11803 (
		\s2_data_i[27]_pad ,
		\s7_data_i[27]_pad ,
		_w9330_,
		_w9608_,
		_w13704_
	);
	LUT4 #(
		.INIT('h8000)
	) name11804 (
		_w13701_,
		_w13702_,
		_w13703_,
		_w13704_,
		_w13705_
	);
	LUT2 #(
		.INIT('h8)
	) name11805 (
		\s14_data_i[27]_pad ,
		_w9603_,
		_w13706_
	);
	LUT4 #(
		.INIT('h135f)
	) name11806 (
		\s3_data_i[27]_pad ,
		\s4_data_i[27]_pad ,
		_w9611_,
		_w9614_,
		_w13707_
	);
	LUT4 #(
		.INIT('h135f)
	) name11807 (
		\s11_data_i[27]_pad ,
		\s8_data_i[27]_pad ,
		_w9597_,
		_w9623_,
		_w13708_
	);
	LUT4 #(
		.INIT('h135f)
	) name11808 (
		\s0_data_i[27]_pad ,
		\s9_data_i[27]_pad ,
		_w9315_,
		_w9327_,
		_w13709_
	);
	LUT4 #(
		.INIT('h4000)
	) name11809 (
		_w13706_,
		_w13707_,
		_w13708_,
		_w13709_,
		_w13710_
	);
	LUT2 #(
		.INIT('h8)
	) name11810 (
		_w13705_,
		_w13710_,
		_w13711_
	);
	LUT4 #(
		.INIT('h70ff)
	) name11811 (
		_w2046_,
		_w2097_,
		_w13700_,
		_w13711_,
		_w13712_
	);
	LUT2 #(
		.INIT('h8)
	) name11812 (
		\s15_data_i[28]_pad ,
		_w2052_,
		_w13713_
	);
	LUT4 #(
		.INIT('h135f)
	) name11813 (
		\s12_data_i[28]_pad ,
		\s13_data_i[28]_pad ,
		_w9339_,
		_w9600_,
		_w13714_
	);
	LUT4 #(
		.INIT('h153f)
	) name11814 (
		\s10_data_i[28]_pad ,
		\s1_data_i[28]_pad ,
		_w9319_,
		_w9594_,
		_w13715_
	);
	LUT4 #(
		.INIT('h135f)
	) name11815 (
		\s5_data_i[28]_pad ,
		\s6_data_i[28]_pad ,
		_w9333_,
		_w9617_,
		_w13716_
	);
	LUT4 #(
		.INIT('h153f)
	) name11816 (
		\s2_data_i[28]_pad ,
		\s7_data_i[28]_pad ,
		_w9330_,
		_w9608_,
		_w13717_
	);
	LUT4 #(
		.INIT('h8000)
	) name11817 (
		_w13714_,
		_w13715_,
		_w13716_,
		_w13717_,
		_w13718_
	);
	LUT2 #(
		.INIT('h8)
	) name11818 (
		\s14_data_i[28]_pad ,
		_w9603_,
		_w13719_
	);
	LUT4 #(
		.INIT('h135f)
	) name11819 (
		\s3_data_i[28]_pad ,
		\s4_data_i[28]_pad ,
		_w9611_,
		_w9614_,
		_w13720_
	);
	LUT4 #(
		.INIT('h135f)
	) name11820 (
		\s11_data_i[28]_pad ,
		\s8_data_i[28]_pad ,
		_w9597_,
		_w9623_,
		_w13721_
	);
	LUT4 #(
		.INIT('h135f)
	) name11821 (
		\s0_data_i[28]_pad ,
		\s9_data_i[28]_pad ,
		_w9315_,
		_w9327_,
		_w13722_
	);
	LUT4 #(
		.INIT('h4000)
	) name11822 (
		_w13719_,
		_w13720_,
		_w13721_,
		_w13722_,
		_w13723_
	);
	LUT2 #(
		.INIT('h8)
	) name11823 (
		_w13718_,
		_w13723_,
		_w13724_
	);
	LUT4 #(
		.INIT('h70ff)
	) name11824 (
		_w2046_,
		_w2097_,
		_w13713_,
		_w13724_,
		_w13725_
	);
	LUT2 #(
		.INIT('h8)
	) name11825 (
		\s15_data_i[29]_pad ,
		_w2052_,
		_w13726_
	);
	LUT4 #(
		.INIT('h135f)
	) name11826 (
		\s12_data_i[29]_pad ,
		\s13_data_i[29]_pad ,
		_w9339_,
		_w9600_,
		_w13727_
	);
	LUT4 #(
		.INIT('h153f)
	) name11827 (
		\s10_data_i[29]_pad ,
		\s1_data_i[29]_pad ,
		_w9319_,
		_w9594_,
		_w13728_
	);
	LUT4 #(
		.INIT('h135f)
	) name11828 (
		\s5_data_i[29]_pad ,
		\s6_data_i[29]_pad ,
		_w9333_,
		_w9617_,
		_w13729_
	);
	LUT4 #(
		.INIT('h153f)
	) name11829 (
		\s2_data_i[29]_pad ,
		\s7_data_i[29]_pad ,
		_w9330_,
		_w9608_,
		_w13730_
	);
	LUT4 #(
		.INIT('h8000)
	) name11830 (
		_w13727_,
		_w13728_,
		_w13729_,
		_w13730_,
		_w13731_
	);
	LUT2 #(
		.INIT('h8)
	) name11831 (
		\s14_data_i[29]_pad ,
		_w9603_,
		_w13732_
	);
	LUT4 #(
		.INIT('h135f)
	) name11832 (
		\s3_data_i[29]_pad ,
		\s4_data_i[29]_pad ,
		_w9611_,
		_w9614_,
		_w13733_
	);
	LUT4 #(
		.INIT('h135f)
	) name11833 (
		\s11_data_i[29]_pad ,
		\s8_data_i[29]_pad ,
		_w9597_,
		_w9623_,
		_w13734_
	);
	LUT4 #(
		.INIT('h135f)
	) name11834 (
		\s0_data_i[29]_pad ,
		\s9_data_i[29]_pad ,
		_w9315_,
		_w9327_,
		_w13735_
	);
	LUT4 #(
		.INIT('h4000)
	) name11835 (
		_w13732_,
		_w13733_,
		_w13734_,
		_w13735_,
		_w13736_
	);
	LUT2 #(
		.INIT('h8)
	) name11836 (
		_w13731_,
		_w13736_,
		_w13737_
	);
	LUT4 #(
		.INIT('h70ff)
	) name11837 (
		_w2046_,
		_w2097_,
		_w13726_,
		_w13737_,
		_w13738_
	);
	LUT3 #(
		.INIT('h80)
	) name11838 (
		_w2052_,
		_w2097_,
		_w9993_,
		_w13739_
	);
	LUT2 #(
		.INIT('h8)
	) name11839 (
		\s15_data_i[2]_pad ,
		_w2052_,
		_w13740_
	);
	LUT3 #(
		.INIT('h70)
	) name11840 (
		_w2046_,
		_w2097_,
		_w13740_,
		_w13741_
	);
	LUT4 #(
		.INIT('h135f)
	) name11841 (
		\s1_data_i[2]_pad ,
		\s8_data_i[2]_pad ,
		_w9319_,
		_w9623_,
		_w13742_
	);
	LUT4 #(
		.INIT('h135f)
	) name11842 (
		\s4_data_i[2]_pad ,
		\s6_data_i[2]_pad ,
		_w9614_,
		_w9617_,
		_w13743_
	);
	LUT4 #(
		.INIT('h153f)
	) name11843 (
		\s5_data_i[2]_pad ,
		\s9_data_i[2]_pad ,
		_w9327_,
		_w9333_,
		_w13744_
	);
	LUT4 #(
		.INIT('h153f)
	) name11844 (
		\s10_data_i[2]_pad ,
		\s7_data_i[2]_pad ,
		_w9330_,
		_w9594_,
		_w13745_
	);
	LUT4 #(
		.INIT('h8000)
	) name11845 (
		_w13742_,
		_w13743_,
		_w13744_,
		_w13745_,
		_w13746_
	);
	LUT2 #(
		.INIT('h8)
	) name11846 (
		\s11_data_i[2]_pad ,
		_w9597_,
		_w13747_
	);
	LUT4 #(
		.INIT('h135f)
	) name11847 (
		\s13_data_i[2]_pad ,
		\s3_data_i[2]_pad ,
		_w9600_,
		_w9611_,
		_w13748_
	);
	LUT4 #(
		.INIT('h135f)
	) name11848 (
		\s12_data_i[2]_pad ,
		\s14_data_i[2]_pad ,
		_w9339_,
		_w9603_,
		_w13749_
	);
	LUT4 #(
		.INIT('h135f)
	) name11849 (
		\s0_data_i[2]_pad ,
		\s2_data_i[2]_pad ,
		_w9315_,
		_w9608_,
		_w13750_
	);
	LUT4 #(
		.INIT('h4000)
	) name11850 (
		_w13747_,
		_w13748_,
		_w13749_,
		_w13750_,
		_w13751_
	);
	LUT2 #(
		.INIT('h8)
	) name11851 (
		_w13746_,
		_w13751_,
		_w13752_
	);
	LUT3 #(
		.INIT('hef)
	) name11852 (
		_w13739_,
		_w13741_,
		_w13752_,
		_w13753_
	);
	LUT2 #(
		.INIT('h8)
	) name11853 (
		\s15_data_i[30]_pad ,
		_w2052_,
		_w13754_
	);
	LUT4 #(
		.INIT('h135f)
	) name11854 (
		\s12_data_i[30]_pad ,
		\s13_data_i[30]_pad ,
		_w9339_,
		_w9600_,
		_w13755_
	);
	LUT4 #(
		.INIT('h153f)
	) name11855 (
		\s10_data_i[30]_pad ,
		\s1_data_i[30]_pad ,
		_w9319_,
		_w9594_,
		_w13756_
	);
	LUT4 #(
		.INIT('h135f)
	) name11856 (
		\s5_data_i[30]_pad ,
		\s6_data_i[30]_pad ,
		_w9333_,
		_w9617_,
		_w13757_
	);
	LUT4 #(
		.INIT('h153f)
	) name11857 (
		\s2_data_i[30]_pad ,
		\s7_data_i[30]_pad ,
		_w9330_,
		_w9608_,
		_w13758_
	);
	LUT4 #(
		.INIT('h8000)
	) name11858 (
		_w13755_,
		_w13756_,
		_w13757_,
		_w13758_,
		_w13759_
	);
	LUT2 #(
		.INIT('h8)
	) name11859 (
		\s14_data_i[30]_pad ,
		_w9603_,
		_w13760_
	);
	LUT4 #(
		.INIT('h135f)
	) name11860 (
		\s3_data_i[30]_pad ,
		\s4_data_i[30]_pad ,
		_w9611_,
		_w9614_,
		_w13761_
	);
	LUT4 #(
		.INIT('h135f)
	) name11861 (
		\s11_data_i[30]_pad ,
		\s8_data_i[30]_pad ,
		_w9597_,
		_w9623_,
		_w13762_
	);
	LUT4 #(
		.INIT('h135f)
	) name11862 (
		\s0_data_i[30]_pad ,
		\s9_data_i[30]_pad ,
		_w9315_,
		_w9327_,
		_w13763_
	);
	LUT4 #(
		.INIT('h4000)
	) name11863 (
		_w13760_,
		_w13761_,
		_w13762_,
		_w13763_,
		_w13764_
	);
	LUT2 #(
		.INIT('h8)
	) name11864 (
		_w13759_,
		_w13764_,
		_w13765_
	);
	LUT4 #(
		.INIT('h70ff)
	) name11865 (
		_w2046_,
		_w2097_,
		_w13754_,
		_w13765_,
		_w13766_
	);
	LUT2 #(
		.INIT('h8)
	) name11866 (
		\s15_data_i[31]_pad ,
		_w2052_,
		_w13767_
	);
	LUT4 #(
		.INIT('h135f)
	) name11867 (
		\s12_data_i[31]_pad ,
		\s13_data_i[31]_pad ,
		_w9339_,
		_w9600_,
		_w13768_
	);
	LUT4 #(
		.INIT('h153f)
	) name11868 (
		\s10_data_i[31]_pad ,
		\s1_data_i[31]_pad ,
		_w9319_,
		_w9594_,
		_w13769_
	);
	LUT4 #(
		.INIT('h135f)
	) name11869 (
		\s5_data_i[31]_pad ,
		\s6_data_i[31]_pad ,
		_w9333_,
		_w9617_,
		_w13770_
	);
	LUT4 #(
		.INIT('h153f)
	) name11870 (
		\s2_data_i[31]_pad ,
		\s7_data_i[31]_pad ,
		_w9330_,
		_w9608_,
		_w13771_
	);
	LUT4 #(
		.INIT('h8000)
	) name11871 (
		_w13768_,
		_w13769_,
		_w13770_,
		_w13771_,
		_w13772_
	);
	LUT2 #(
		.INIT('h8)
	) name11872 (
		\s14_data_i[31]_pad ,
		_w9603_,
		_w13773_
	);
	LUT4 #(
		.INIT('h135f)
	) name11873 (
		\s3_data_i[31]_pad ,
		\s4_data_i[31]_pad ,
		_w9611_,
		_w9614_,
		_w13774_
	);
	LUT4 #(
		.INIT('h135f)
	) name11874 (
		\s11_data_i[31]_pad ,
		\s8_data_i[31]_pad ,
		_w9597_,
		_w9623_,
		_w13775_
	);
	LUT4 #(
		.INIT('h135f)
	) name11875 (
		\s0_data_i[31]_pad ,
		\s9_data_i[31]_pad ,
		_w9315_,
		_w9327_,
		_w13776_
	);
	LUT4 #(
		.INIT('h4000)
	) name11876 (
		_w13773_,
		_w13774_,
		_w13775_,
		_w13776_,
		_w13777_
	);
	LUT2 #(
		.INIT('h8)
	) name11877 (
		_w13772_,
		_w13777_,
		_w13778_
	);
	LUT4 #(
		.INIT('h70ff)
	) name11878 (
		_w2046_,
		_w2097_,
		_w13767_,
		_w13778_,
		_w13779_
	);
	LUT3 #(
		.INIT('h80)
	) name11879 (
		_w2052_,
		_w2097_,
		_w10035_,
		_w13780_
	);
	LUT2 #(
		.INIT('h8)
	) name11880 (
		\s15_data_i[3]_pad ,
		_w2052_,
		_w13781_
	);
	LUT3 #(
		.INIT('h70)
	) name11881 (
		_w2046_,
		_w2097_,
		_w13781_,
		_w13782_
	);
	LUT4 #(
		.INIT('h135f)
	) name11882 (
		\s7_data_i[3]_pad ,
		\s8_data_i[3]_pad ,
		_w9330_,
		_w9623_,
		_w13783_
	);
	LUT4 #(
		.INIT('h153f)
	) name11883 (
		\s10_data_i[3]_pad ,
		\s1_data_i[3]_pad ,
		_w9319_,
		_w9594_,
		_w13784_
	);
	LUT4 #(
		.INIT('h153f)
	) name11884 (
		\s5_data_i[3]_pad ,
		\s9_data_i[3]_pad ,
		_w9327_,
		_w9333_,
		_w13785_
	);
	LUT4 #(
		.INIT('h135f)
	) name11885 (
		\s13_data_i[3]_pad ,
		\s2_data_i[3]_pad ,
		_w9600_,
		_w9608_,
		_w13786_
	);
	LUT4 #(
		.INIT('h8000)
	) name11886 (
		_w13783_,
		_w13784_,
		_w13785_,
		_w13786_,
		_w13787_
	);
	LUT2 #(
		.INIT('h8)
	) name11887 (
		\s11_data_i[3]_pad ,
		_w9597_,
		_w13788_
	);
	LUT4 #(
		.INIT('h135f)
	) name11888 (
		\s3_data_i[3]_pad ,
		\s4_data_i[3]_pad ,
		_w9611_,
		_w9614_,
		_w13789_
	);
	LUT4 #(
		.INIT('h135f)
	) name11889 (
		\s12_data_i[3]_pad ,
		\s14_data_i[3]_pad ,
		_w9339_,
		_w9603_,
		_w13790_
	);
	LUT4 #(
		.INIT('h135f)
	) name11890 (
		\s0_data_i[3]_pad ,
		\s6_data_i[3]_pad ,
		_w9315_,
		_w9617_,
		_w13791_
	);
	LUT4 #(
		.INIT('h4000)
	) name11891 (
		_w13788_,
		_w13789_,
		_w13790_,
		_w13791_,
		_w13792_
	);
	LUT2 #(
		.INIT('h8)
	) name11892 (
		_w13787_,
		_w13792_,
		_w13793_
	);
	LUT3 #(
		.INIT('hef)
	) name11893 (
		_w13780_,
		_w13782_,
		_w13793_,
		_w13794_
	);
	LUT3 #(
		.INIT('h80)
	) name11894 (
		_w2052_,
		_w2097_,
		_w10051_,
		_w13795_
	);
	LUT2 #(
		.INIT('h8)
	) name11895 (
		\s15_data_i[4]_pad ,
		_w2052_,
		_w13796_
	);
	LUT3 #(
		.INIT('h70)
	) name11896 (
		_w2046_,
		_w2097_,
		_w13796_,
		_w13797_
	);
	LUT4 #(
		.INIT('h135f)
	) name11897 (
		\s1_data_i[4]_pad ,
		\s8_data_i[4]_pad ,
		_w9319_,
		_w9623_,
		_w13798_
	);
	LUT4 #(
		.INIT('h135f)
	) name11898 (
		\s4_data_i[4]_pad ,
		\s6_data_i[4]_pad ,
		_w9614_,
		_w9617_,
		_w13799_
	);
	LUT4 #(
		.INIT('h153f)
	) name11899 (
		\s5_data_i[4]_pad ,
		\s9_data_i[4]_pad ,
		_w9327_,
		_w9333_,
		_w13800_
	);
	LUT4 #(
		.INIT('h153f)
	) name11900 (
		\s10_data_i[4]_pad ,
		\s7_data_i[4]_pad ,
		_w9330_,
		_w9594_,
		_w13801_
	);
	LUT4 #(
		.INIT('h8000)
	) name11901 (
		_w13798_,
		_w13799_,
		_w13800_,
		_w13801_,
		_w13802_
	);
	LUT2 #(
		.INIT('h8)
	) name11902 (
		\s11_data_i[4]_pad ,
		_w9597_,
		_w13803_
	);
	LUT4 #(
		.INIT('h135f)
	) name11903 (
		\s13_data_i[4]_pad ,
		\s3_data_i[4]_pad ,
		_w9600_,
		_w9611_,
		_w13804_
	);
	LUT4 #(
		.INIT('h135f)
	) name11904 (
		\s12_data_i[4]_pad ,
		\s14_data_i[4]_pad ,
		_w9339_,
		_w9603_,
		_w13805_
	);
	LUT4 #(
		.INIT('h135f)
	) name11905 (
		\s0_data_i[4]_pad ,
		\s2_data_i[4]_pad ,
		_w9315_,
		_w9608_,
		_w13806_
	);
	LUT4 #(
		.INIT('h4000)
	) name11906 (
		_w13803_,
		_w13804_,
		_w13805_,
		_w13806_,
		_w13807_
	);
	LUT2 #(
		.INIT('h8)
	) name11907 (
		_w13802_,
		_w13807_,
		_w13808_
	);
	LUT3 #(
		.INIT('hef)
	) name11908 (
		_w13795_,
		_w13797_,
		_w13808_,
		_w13809_
	);
	LUT3 #(
		.INIT('h80)
	) name11909 (
		_w2052_,
		_w2097_,
		_w10067_,
		_w13810_
	);
	LUT2 #(
		.INIT('h8)
	) name11910 (
		\s15_data_i[5]_pad ,
		_w2052_,
		_w13811_
	);
	LUT3 #(
		.INIT('h70)
	) name11911 (
		_w2046_,
		_w2097_,
		_w13811_,
		_w13812_
	);
	LUT4 #(
		.INIT('h135f)
	) name11912 (
		\s13_data_i[5]_pad ,
		\s2_data_i[5]_pad ,
		_w9600_,
		_w9608_,
		_w13813_
	);
	LUT4 #(
		.INIT('h135f)
	) name11913 (
		\s12_data_i[5]_pad ,
		\s4_data_i[5]_pad ,
		_w9339_,
		_w9614_,
		_w13814_
	);
	LUT4 #(
		.INIT('h135f)
	) name11914 (
		\s14_data_i[5]_pad ,
		\s3_data_i[5]_pad ,
		_w9603_,
		_w9611_,
		_w13815_
	);
	LUT4 #(
		.INIT('h135f)
	) name11915 (
		\s11_data_i[5]_pad ,
		\s8_data_i[5]_pad ,
		_w9597_,
		_w9623_,
		_w13816_
	);
	LUT4 #(
		.INIT('h8000)
	) name11916 (
		_w13813_,
		_w13814_,
		_w13815_,
		_w13816_,
		_w13817_
	);
	LUT2 #(
		.INIT('h8)
	) name11917 (
		\s1_data_i[5]_pad ,
		_w9319_,
		_w13818_
	);
	LUT4 #(
		.INIT('h153f)
	) name11918 (
		\s5_data_i[5]_pad ,
		\s7_data_i[5]_pad ,
		_w9330_,
		_w9333_,
		_w13819_
	);
	LUT4 #(
		.INIT('h153f)
	) name11919 (
		\s10_data_i[5]_pad ,
		\s9_data_i[5]_pad ,
		_w9327_,
		_w9594_,
		_w13820_
	);
	LUT4 #(
		.INIT('h135f)
	) name11920 (
		\s0_data_i[5]_pad ,
		\s6_data_i[5]_pad ,
		_w9315_,
		_w9617_,
		_w13821_
	);
	LUT4 #(
		.INIT('h4000)
	) name11921 (
		_w13818_,
		_w13819_,
		_w13820_,
		_w13821_,
		_w13822_
	);
	LUT2 #(
		.INIT('h8)
	) name11922 (
		_w13817_,
		_w13822_,
		_w13823_
	);
	LUT3 #(
		.INIT('hef)
	) name11923 (
		_w13810_,
		_w13812_,
		_w13823_,
		_w13824_
	);
	LUT3 #(
		.INIT('h80)
	) name11924 (
		_w2052_,
		_w2097_,
		_w10083_,
		_w13825_
	);
	LUT2 #(
		.INIT('h8)
	) name11925 (
		\s15_data_i[6]_pad ,
		_w2052_,
		_w13826_
	);
	LUT3 #(
		.INIT('h70)
	) name11926 (
		_w2046_,
		_w2097_,
		_w13826_,
		_w13827_
	);
	LUT4 #(
		.INIT('h135f)
	) name11927 (
		\s1_data_i[6]_pad ,
		\s8_data_i[6]_pad ,
		_w9319_,
		_w9623_,
		_w13828_
	);
	LUT4 #(
		.INIT('h135f)
	) name11928 (
		\s4_data_i[6]_pad ,
		\s6_data_i[6]_pad ,
		_w9614_,
		_w9617_,
		_w13829_
	);
	LUT4 #(
		.INIT('h153f)
	) name11929 (
		\s5_data_i[6]_pad ,
		\s9_data_i[6]_pad ,
		_w9327_,
		_w9333_,
		_w13830_
	);
	LUT4 #(
		.INIT('h153f)
	) name11930 (
		\s10_data_i[6]_pad ,
		\s7_data_i[6]_pad ,
		_w9330_,
		_w9594_,
		_w13831_
	);
	LUT4 #(
		.INIT('h8000)
	) name11931 (
		_w13828_,
		_w13829_,
		_w13830_,
		_w13831_,
		_w13832_
	);
	LUT2 #(
		.INIT('h8)
	) name11932 (
		\s11_data_i[6]_pad ,
		_w9597_,
		_w13833_
	);
	LUT4 #(
		.INIT('h135f)
	) name11933 (
		\s13_data_i[6]_pad ,
		\s3_data_i[6]_pad ,
		_w9600_,
		_w9611_,
		_w13834_
	);
	LUT4 #(
		.INIT('h135f)
	) name11934 (
		\s12_data_i[6]_pad ,
		\s14_data_i[6]_pad ,
		_w9339_,
		_w9603_,
		_w13835_
	);
	LUT4 #(
		.INIT('h135f)
	) name11935 (
		\s0_data_i[6]_pad ,
		\s2_data_i[6]_pad ,
		_w9315_,
		_w9608_,
		_w13836_
	);
	LUT4 #(
		.INIT('h4000)
	) name11936 (
		_w13833_,
		_w13834_,
		_w13835_,
		_w13836_,
		_w13837_
	);
	LUT2 #(
		.INIT('h8)
	) name11937 (
		_w13832_,
		_w13837_,
		_w13838_
	);
	LUT3 #(
		.INIT('hef)
	) name11938 (
		_w13825_,
		_w13827_,
		_w13838_,
		_w13839_
	);
	LUT3 #(
		.INIT('h80)
	) name11939 (
		_w2052_,
		_w2097_,
		_w10099_,
		_w13840_
	);
	LUT2 #(
		.INIT('h8)
	) name11940 (
		\s15_data_i[7]_pad ,
		_w2052_,
		_w13841_
	);
	LUT3 #(
		.INIT('h70)
	) name11941 (
		_w2046_,
		_w2097_,
		_w13841_,
		_w13842_
	);
	LUT4 #(
		.INIT('h135f)
	) name11942 (
		\s1_data_i[7]_pad ,
		\s8_data_i[7]_pad ,
		_w9319_,
		_w9623_,
		_w13843_
	);
	LUT4 #(
		.INIT('h135f)
	) name11943 (
		\s4_data_i[7]_pad ,
		\s6_data_i[7]_pad ,
		_w9614_,
		_w9617_,
		_w13844_
	);
	LUT4 #(
		.INIT('h153f)
	) name11944 (
		\s5_data_i[7]_pad ,
		\s9_data_i[7]_pad ,
		_w9327_,
		_w9333_,
		_w13845_
	);
	LUT4 #(
		.INIT('h153f)
	) name11945 (
		\s10_data_i[7]_pad ,
		\s7_data_i[7]_pad ,
		_w9330_,
		_w9594_,
		_w13846_
	);
	LUT4 #(
		.INIT('h8000)
	) name11946 (
		_w13843_,
		_w13844_,
		_w13845_,
		_w13846_,
		_w13847_
	);
	LUT2 #(
		.INIT('h8)
	) name11947 (
		\s11_data_i[7]_pad ,
		_w9597_,
		_w13848_
	);
	LUT4 #(
		.INIT('h135f)
	) name11948 (
		\s13_data_i[7]_pad ,
		\s3_data_i[7]_pad ,
		_w9600_,
		_w9611_,
		_w13849_
	);
	LUT4 #(
		.INIT('h135f)
	) name11949 (
		\s12_data_i[7]_pad ,
		\s14_data_i[7]_pad ,
		_w9339_,
		_w9603_,
		_w13850_
	);
	LUT4 #(
		.INIT('h135f)
	) name11950 (
		\s0_data_i[7]_pad ,
		\s2_data_i[7]_pad ,
		_w9315_,
		_w9608_,
		_w13851_
	);
	LUT4 #(
		.INIT('h4000)
	) name11951 (
		_w13848_,
		_w13849_,
		_w13850_,
		_w13851_,
		_w13852_
	);
	LUT2 #(
		.INIT('h8)
	) name11952 (
		_w13847_,
		_w13852_,
		_w13853_
	);
	LUT3 #(
		.INIT('hef)
	) name11953 (
		_w13840_,
		_w13842_,
		_w13853_,
		_w13854_
	);
	LUT3 #(
		.INIT('h80)
	) name11954 (
		_w2052_,
		_w2097_,
		_w10115_,
		_w13855_
	);
	LUT2 #(
		.INIT('h8)
	) name11955 (
		\s15_data_i[8]_pad ,
		_w2052_,
		_w13856_
	);
	LUT3 #(
		.INIT('h70)
	) name11956 (
		_w2046_,
		_w2097_,
		_w13856_,
		_w13857_
	);
	LUT4 #(
		.INIT('h135f)
	) name11957 (
		\s1_data_i[8]_pad ,
		\s8_data_i[8]_pad ,
		_w9319_,
		_w9623_,
		_w13858_
	);
	LUT4 #(
		.INIT('h135f)
	) name11958 (
		\s4_data_i[8]_pad ,
		\s6_data_i[8]_pad ,
		_w9614_,
		_w9617_,
		_w13859_
	);
	LUT4 #(
		.INIT('h153f)
	) name11959 (
		\s5_data_i[8]_pad ,
		\s9_data_i[8]_pad ,
		_w9327_,
		_w9333_,
		_w13860_
	);
	LUT4 #(
		.INIT('h153f)
	) name11960 (
		\s10_data_i[8]_pad ,
		\s7_data_i[8]_pad ,
		_w9330_,
		_w9594_,
		_w13861_
	);
	LUT4 #(
		.INIT('h8000)
	) name11961 (
		_w13858_,
		_w13859_,
		_w13860_,
		_w13861_,
		_w13862_
	);
	LUT2 #(
		.INIT('h8)
	) name11962 (
		\s11_data_i[8]_pad ,
		_w9597_,
		_w13863_
	);
	LUT4 #(
		.INIT('h135f)
	) name11963 (
		\s13_data_i[8]_pad ,
		\s3_data_i[8]_pad ,
		_w9600_,
		_w9611_,
		_w13864_
	);
	LUT4 #(
		.INIT('h135f)
	) name11964 (
		\s12_data_i[8]_pad ,
		\s14_data_i[8]_pad ,
		_w9339_,
		_w9603_,
		_w13865_
	);
	LUT4 #(
		.INIT('h135f)
	) name11965 (
		\s0_data_i[8]_pad ,
		\s2_data_i[8]_pad ,
		_w9315_,
		_w9608_,
		_w13866_
	);
	LUT4 #(
		.INIT('h4000)
	) name11966 (
		_w13863_,
		_w13864_,
		_w13865_,
		_w13866_,
		_w13867_
	);
	LUT2 #(
		.INIT('h8)
	) name11967 (
		_w13862_,
		_w13867_,
		_w13868_
	);
	LUT3 #(
		.INIT('hef)
	) name11968 (
		_w13855_,
		_w13857_,
		_w13868_,
		_w13869_
	);
	LUT3 #(
		.INIT('h80)
	) name11969 (
		_w2052_,
		_w2097_,
		_w10131_,
		_w13870_
	);
	LUT2 #(
		.INIT('h8)
	) name11970 (
		\s15_data_i[9]_pad ,
		_w2052_,
		_w13871_
	);
	LUT3 #(
		.INIT('h70)
	) name11971 (
		_w2046_,
		_w2097_,
		_w13871_,
		_w13872_
	);
	LUT4 #(
		.INIT('h135f)
	) name11972 (
		\s1_data_i[9]_pad ,
		\s8_data_i[9]_pad ,
		_w9319_,
		_w9623_,
		_w13873_
	);
	LUT4 #(
		.INIT('h135f)
	) name11973 (
		\s4_data_i[9]_pad ,
		\s6_data_i[9]_pad ,
		_w9614_,
		_w9617_,
		_w13874_
	);
	LUT4 #(
		.INIT('h153f)
	) name11974 (
		\s5_data_i[9]_pad ,
		\s9_data_i[9]_pad ,
		_w9327_,
		_w9333_,
		_w13875_
	);
	LUT4 #(
		.INIT('h153f)
	) name11975 (
		\s10_data_i[9]_pad ,
		\s7_data_i[9]_pad ,
		_w9330_,
		_w9594_,
		_w13876_
	);
	LUT4 #(
		.INIT('h8000)
	) name11976 (
		_w13873_,
		_w13874_,
		_w13875_,
		_w13876_,
		_w13877_
	);
	LUT2 #(
		.INIT('h8)
	) name11977 (
		\s11_data_i[9]_pad ,
		_w9597_,
		_w13878_
	);
	LUT4 #(
		.INIT('h135f)
	) name11978 (
		\s13_data_i[9]_pad ,
		\s3_data_i[9]_pad ,
		_w9600_,
		_w9611_,
		_w13879_
	);
	LUT4 #(
		.INIT('h135f)
	) name11979 (
		\s12_data_i[9]_pad ,
		\s14_data_i[9]_pad ,
		_w9339_,
		_w9603_,
		_w13880_
	);
	LUT4 #(
		.INIT('h135f)
	) name11980 (
		\s0_data_i[9]_pad ,
		\s2_data_i[9]_pad ,
		_w9315_,
		_w9608_,
		_w13881_
	);
	LUT4 #(
		.INIT('h4000)
	) name11981 (
		_w13878_,
		_w13879_,
		_w13880_,
		_w13881_,
		_w13882_
	);
	LUT2 #(
		.INIT('h8)
	) name11982 (
		_w13877_,
		_w13882_,
		_w13883_
	);
	LUT3 #(
		.INIT('hef)
	) name11983 (
		_w13870_,
		_w13872_,
		_w13883_,
		_w13884_
	);
	LUT3 #(
		.INIT('h80)
	) name11984 (
		\s15_err_i_pad ,
		_w1918_,
		_w13407_,
		_w13885_
	);
	LUT4 #(
		.INIT('h2a00)
	) name11985 (
		\s11_err_i_pad ,
		_w8955_,
		_w8956_,
		_w9597_,
		_w13886_
	);
	LUT4 #(
		.INIT('h2a00)
	) name11986 (
		\s3_err_i_pad ,
		_w9205_,
		_w9206_,
		_w9611_,
		_w13887_
	);
	LUT4 #(
		.INIT('h135f)
	) name11987 (
		_w8968_,
		_w9218_,
		_w13886_,
		_w13887_,
		_w13888_
	);
	LUT4 #(
		.INIT('h2a00)
	) name11988 (
		\s13_err_i_pad ,
		_w9069_,
		_w9070_,
		_w9600_,
		_w13889_
	);
	LUT4 #(
		.INIT('h2a00)
	) name11989 (
		\s9_err_i_pad ,
		_w8865_,
		_w8866_,
		_w9327_,
		_w13890_
	);
	LUT4 #(
		.INIT('h153f)
	) name11990 (
		_w8878_,
		_w9068_,
		_w13889_,
		_w13890_,
		_w13891_
	);
	LUT4 #(
		.INIT('h2a00)
	) name11991 (
		\s6_err_i_pad ,
		_w8743_,
		_w8744_,
		_w9617_,
		_w13892_
	);
	LUT4 #(
		.INIT('h2a00)
	) name11992 (
		\s0_err_i_pad ,
		_w8989_,
		_w8990_,
		_w9315_,
		_w13893_
	);
	LUT4 #(
		.INIT('h135f)
	) name11993 (
		_w8756_,
		_w8988_,
		_w13892_,
		_w13893_,
		_w13894_
	);
	LUT4 #(
		.INIT('h2a00)
	) name11994 (
		\s4_err_i_pad ,
		_w8655_,
		_w8656_,
		_w9614_,
		_w13895_
	);
	LUT4 #(
		.INIT('h2a00)
	) name11995 (
		\s10_err_i_pad ,
		_w8910_,
		_w8911_,
		_w9594_,
		_w13896_
	);
	LUT4 #(
		.INIT('h135f)
	) name11996 (
		_w8674_,
		_w8917_,
		_w13895_,
		_w13896_,
		_w13897_
	);
	LUT4 #(
		.INIT('h8000)
	) name11997 (
		_w13888_,
		_w13891_,
		_w13894_,
		_w13897_,
		_w13898_
	);
	LUT4 #(
		.INIT('h2a00)
	) name11998 (
		\s8_err_i_pad ,
		_w8821_,
		_w8822_,
		_w9623_,
		_w13899_
	);
	LUT2 #(
		.INIT('h8)
	) name11999 (
		_w8834_,
		_w13899_,
		_w13900_
	);
	LUT4 #(
		.INIT('h2a00)
	) name12000 (
		\s2_err_i_pad ,
		_w9171_,
		_w9172_,
		_w9608_,
		_w13901_
	);
	LUT4 #(
		.INIT('h2a00)
	) name12001 (
		\s7_err_i_pad ,
		_w8782_,
		_w8783_,
		_w9330_,
		_w13902_
	);
	LUT4 #(
		.INIT('h153f)
	) name12002 (
		_w8781_,
		_w9184_,
		_w13901_,
		_w13902_,
		_w13903_
	);
	LUT4 #(
		.INIT('h2a00)
	) name12003 (
		\s12_err_i_pad ,
		_w9029_,
		_w9030_,
		_w9339_,
		_w13904_
	);
	LUT4 #(
		.INIT('h2a00)
	) name12004 (
		\s14_err_i_pad ,
		_w9137_,
		_w9138_,
		_w9603_,
		_w13905_
	);
	LUT4 #(
		.INIT('h135f)
	) name12005 (
		_w9036_,
		_w9150_,
		_w13904_,
		_w13905_,
		_w13906_
	);
	LUT4 #(
		.INIT('h2a00)
	) name12006 (
		\s5_err_i_pad ,
		_w8699_,
		_w8700_,
		_w9333_,
		_w13907_
	);
	LUT4 #(
		.INIT('h2a00)
	) name12007 (
		\s1_err_i_pad ,
		_w9103_,
		_w9104_,
		_w9319_,
		_w13908_
	);
	LUT4 #(
		.INIT('h135f)
	) name12008 (
		_w8712_,
		_w9102_,
		_w13907_,
		_w13908_,
		_w13909_
	);
	LUT4 #(
		.INIT('h4000)
	) name12009 (
		_w13900_,
		_w13903_,
		_w13906_,
		_w13909_,
		_w13910_
	);
	LUT2 #(
		.INIT('h8)
	) name12010 (
		_w13898_,
		_w13910_,
		_w13911_
	);
	LUT4 #(
		.INIT('h70ff)
	) name12011 (
		_w2046_,
		_w2097_,
		_w13885_,
		_w13911_,
		_w13912_
	);
	LUT3 #(
		.INIT('h80)
	) name12012 (
		\s15_rty_i_pad ,
		_w1918_,
		_w13407_,
		_w13913_
	);
	LUT4 #(
		.INIT('h2a00)
	) name12013 (
		\s2_rty_i_pad ,
		_w9171_,
		_w9172_,
		_w9608_,
		_w13914_
	);
	LUT4 #(
		.INIT('h2a00)
	) name12014 (
		\s3_rty_i_pad ,
		_w9205_,
		_w9206_,
		_w9611_,
		_w13915_
	);
	LUT4 #(
		.INIT('h135f)
	) name12015 (
		_w9184_,
		_w9218_,
		_w13914_,
		_w13915_,
		_w13916_
	);
	LUT4 #(
		.INIT('h2a00)
	) name12016 (
		\s13_rty_i_pad ,
		_w9069_,
		_w9070_,
		_w9600_,
		_w13917_
	);
	LUT4 #(
		.INIT('h2a00)
	) name12017 (
		\s9_rty_i_pad ,
		_w8865_,
		_w8866_,
		_w9327_,
		_w13918_
	);
	LUT4 #(
		.INIT('h153f)
	) name12018 (
		_w8878_,
		_w9068_,
		_w13917_,
		_w13918_,
		_w13919_
	);
	LUT4 #(
		.INIT('h2a00)
	) name12019 (
		\s0_rty_i_pad ,
		_w8989_,
		_w8990_,
		_w9315_,
		_w13920_
	);
	LUT4 #(
		.INIT('h2a00)
	) name12020 (
		\s7_rty_i_pad ,
		_w8782_,
		_w8783_,
		_w9330_,
		_w13921_
	);
	LUT4 #(
		.INIT('h153f)
	) name12021 (
		_w8781_,
		_w8988_,
		_w13920_,
		_w13921_,
		_w13922_
	);
	LUT4 #(
		.INIT('h2a00)
	) name12022 (
		\s6_rty_i_pad ,
		_w8743_,
		_w8744_,
		_w9617_,
		_w13923_
	);
	LUT4 #(
		.INIT('h2a00)
	) name12023 (
		\s10_rty_i_pad ,
		_w8910_,
		_w8911_,
		_w9594_,
		_w13924_
	);
	LUT4 #(
		.INIT('h135f)
	) name12024 (
		_w8756_,
		_w8917_,
		_w13923_,
		_w13924_,
		_w13925_
	);
	LUT4 #(
		.INIT('h8000)
	) name12025 (
		_w13916_,
		_w13919_,
		_w13922_,
		_w13925_,
		_w13926_
	);
	LUT4 #(
		.INIT('h2a00)
	) name12026 (
		\s1_rty_i_pad ,
		_w9103_,
		_w9104_,
		_w9319_,
		_w13927_
	);
	LUT2 #(
		.INIT('h8)
	) name12027 (
		_w9102_,
		_w13927_,
		_w13928_
	);
	LUT4 #(
		.INIT('h2a00)
	) name12028 (
		\s11_rty_i_pad ,
		_w8955_,
		_w8956_,
		_w9597_,
		_w13929_
	);
	LUT4 #(
		.INIT('h2a00)
	) name12029 (
		\s4_rty_i_pad ,
		_w8655_,
		_w8656_,
		_w9614_,
		_w13930_
	);
	LUT4 #(
		.INIT('h153f)
	) name12030 (
		_w8674_,
		_w8968_,
		_w13929_,
		_w13930_,
		_w13931_
	);
	LUT4 #(
		.INIT('h2a00)
	) name12031 (
		\s12_rty_i_pad ,
		_w9029_,
		_w9030_,
		_w9339_,
		_w13932_
	);
	LUT4 #(
		.INIT('h2a00)
	) name12032 (
		\s14_rty_i_pad ,
		_w9137_,
		_w9138_,
		_w9603_,
		_w13933_
	);
	LUT4 #(
		.INIT('h135f)
	) name12033 (
		_w9036_,
		_w9150_,
		_w13932_,
		_w13933_,
		_w13934_
	);
	LUT4 #(
		.INIT('h2a00)
	) name12034 (
		\s5_rty_i_pad ,
		_w8699_,
		_w8700_,
		_w9333_,
		_w13935_
	);
	LUT4 #(
		.INIT('h2a00)
	) name12035 (
		\s8_rty_i_pad ,
		_w8821_,
		_w8822_,
		_w9623_,
		_w13936_
	);
	LUT4 #(
		.INIT('h135f)
	) name12036 (
		_w8712_,
		_w8834_,
		_w13935_,
		_w13936_,
		_w13937_
	);
	LUT4 #(
		.INIT('h4000)
	) name12037 (
		_w13928_,
		_w13931_,
		_w13934_,
		_w13937_,
		_w13938_
	);
	LUT2 #(
		.INIT('h8)
	) name12038 (
		_w13926_,
		_w13938_,
		_w13939_
	);
	LUT4 #(
		.INIT('h70ff)
	) name12039 (
		_w2046_,
		_w2097_,
		_w13913_,
		_w13939_,
		_w13940_
	);
	LUT3 #(
		.INIT('h80)
	) name12040 (
		\m2_addr_i[0]_pad ,
		_w8989_,
		_w8990_,
		_w13941_
	);
	LUT3 #(
		.INIT('h2a)
	) name12041 (
		\m3_addr_i[0]_pad ,
		_w8989_,
		_w8990_,
		_w13942_
	);
	LUT3 #(
		.INIT('h57)
	) name12042 (
		_w9002_,
		_w13941_,
		_w13942_,
		_w13943_
	);
	LUT3 #(
		.INIT('h80)
	) name12043 (
		\m0_addr_i[0]_pad ,
		_w8989_,
		_w8990_,
		_w13944_
	);
	LUT3 #(
		.INIT('h2a)
	) name12044 (
		\m7_addr_i[0]_pad ,
		_w8989_,
		_w8990_,
		_w13945_
	);
	LUT4 #(
		.INIT('h6e7f)
	) name12045 (
		_w8984_,
		_w8987_,
		_w13944_,
		_w13945_,
		_w13946_
	);
	LUT3 #(
		.INIT('h2a)
	) name12046 (
		\m1_addr_i[0]_pad ,
		_w8989_,
		_w8990_,
		_w13947_
	);
	LUT3 #(
		.INIT('h80)
	) name12047 (
		\m6_addr_i[0]_pad ,
		_w8989_,
		_w8990_,
		_w13948_
	);
	LUT4 #(
		.INIT('h6e7f)
	) name12048 (
		_w8984_,
		_w8987_,
		_w13947_,
		_w13948_,
		_w13949_
	);
	LUT3 #(
		.INIT('h80)
	) name12049 (
		\m4_addr_i[0]_pad ,
		_w8989_,
		_w8990_,
		_w13950_
	);
	LUT3 #(
		.INIT('h2a)
	) name12050 (
		\m5_addr_i[0]_pad ,
		_w8989_,
		_w8990_,
		_w13951_
	);
	LUT3 #(
		.INIT('h57)
	) name12051 (
		_w8996_,
		_w13950_,
		_w13951_,
		_w13952_
	);
	LUT4 #(
		.INIT('h7fff)
	) name12052 (
		_w13943_,
		_w13946_,
		_w13949_,
		_w13952_,
		_w13953_
	);
	LUT3 #(
		.INIT('h80)
	) name12053 (
		\m2_addr_i[10]_pad ,
		_w8989_,
		_w8990_,
		_w13954_
	);
	LUT3 #(
		.INIT('h2a)
	) name12054 (
		\m3_addr_i[10]_pad ,
		_w8989_,
		_w8990_,
		_w13955_
	);
	LUT3 #(
		.INIT('h57)
	) name12055 (
		_w9002_,
		_w13954_,
		_w13955_,
		_w13956_
	);
	LUT3 #(
		.INIT('h80)
	) name12056 (
		\m0_addr_i[10]_pad ,
		_w8989_,
		_w8990_,
		_w13957_
	);
	LUT3 #(
		.INIT('h2a)
	) name12057 (
		\m5_addr_i[10]_pad ,
		_w8989_,
		_w8990_,
		_w13958_
	);
	LUT4 #(
		.INIT('h5d7f)
	) name12058 (
		_w8984_,
		_w8987_,
		_w13957_,
		_w13958_,
		_w13959_
	);
	LUT3 #(
		.INIT('h2a)
	) name12059 (
		\m1_addr_i[10]_pad ,
		_w8989_,
		_w8990_,
		_w13960_
	);
	LUT3 #(
		.INIT('h80)
	) name12060 (
		\m4_addr_i[10]_pad ,
		_w8989_,
		_w8990_,
		_w13961_
	);
	LUT4 #(
		.INIT('h5d7f)
	) name12061 (
		_w8984_,
		_w8987_,
		_w13960_,
		_w13961_,
		_w13962_
	);
	LUT3 #(
		.INIT('h80)
	) name12062 (
		\m6_addr_i[10]_pad ,
		_w8989_,
		_w8990_,
		_w13963_
	);
	LUT3 #(
		.INIT('h2a)
	) name12063 (
		\m7_addr_i[10]_pad ,
		_w8989_,
		_w8990_,
		_w13964_
	);
	LUT3 #(
		.INIT('h57)
	) name12064 (
		_w8988_,
		_w13963_,
		_w13964_,
		_w13965_
	);
	LUT4 #(
		.INIT('h7fff)
	) name12065 (
		_w13956_,
		_w13959_,
		_w13962_,
		_w13965_,
		_w13966_
	);
	LUT3 #(
		.INIT('h80)
	) name12066 (
		\m2_addr_i[11]_pad ,
		_w8989_,
		_w8990_,
		_w13967_
	);
	LUT3 #(
		.INIT('h2a)
	) name12067 (
		\m3_addr_i[11]_pad ,
		_w8989_,
		_w8990_,
		_w13968_
	);
	LUT3 #(
		.INIT('h57)
	) name12068 (
		_w9002_,
		_w13967_,
		_w13968_,
		_w13969_
	);
	LUT3 #(
		.INIT('h80)
	) name12069 (
		\m6_addr_i[11]_pad ,
		_w8989_,
		_w8990_,
		_w13970_
	);
	LUT3 #(
		.INIT('h2a)
	) name12070 (
		\m1_addr_i[11]_pad ,
		_w8989_,
		_w8990_,
		_w13971_
	);
	LUT4 #(
		.INIT('h67ef)
	) name12071 (
		_w8984_,
		_w8987_,
		_w13970_,
		_w13971_,
		_w13972_
	);
	LUT3 #(
		.INIT('h2a)
	) name12072 (
		\m7_addr_i[11]_pad ,
		_w8989_,
		_w8990_,
		_w13973_
	);
	LUT3 #(
		.INIT('h80)
	) name12073 (
		\m0_addr_i[11]_pad ,
		_w8989_,
		_w8990_,
		_w13974_
	);
	LUT4 #(
		.INIT('h67ef)
	) name12074 (
		_w8984_,
		_w8987_,
		_w13973_,
		_w13974_,
		_w13975_
	);
	LUT3 #(
		.INIT('h80)
	) name12075 (
		\m4_addr_i[11]_pad ,
		_w8989_,
		_w8990_,
		_w13976_
	);
	LUT3 #(
		.INIT('h2a)
	) name12076 (
		\m5_addr_i[11]_pad ,
		_w8989_,
		_w8990_,
		_w13977_
	);
	LUT3 #(
		.INIT('h57)
	) name12077 (
		_w8996_,
		_w13976_,
		_w13977_,
		_w13978_
	);
	LUT4 #(
		.INIT('h7fff)
	) name12078 (
		_w13969_,
		_w13972_,
		_w13975_,
		_w13978_,
		_w13979_
	);
	LUT3 #(
		.INIT('h80)
	) name12079 (
		\m6_addr_i[12]_pad ,
		_w8989_,
		_w8990_,
		_w13980_
	);
	LUT3 #(
		.INIT('h2a)
	) name12080 (
		\m7_addr_i[12]_pad ,
		_w8989_,
		_w8990_,
		_w13981_
	);
	LUT3 #(
		.INIT('h57)
	) name12081 (
		_w8988_,
		_w13980_,
		_w13981_,
		_w13982_
	);
	LUT3 #(
		.INIT('h80)
	) name12082 (
		\m4_addr_i[12]_pad ,
		_w8989_,
		_w8990_,
		_w13983_
	);
	LUT3 #(
		.INIT('h2a)
	) name12083 (
		\m3_addr_i[12]_pad ,
		_w8989_,
		_w8990_,
		_w13984_
	);
	LUT4 #(
		.INIT('h9bdf)
	) name12084 (
		_w8984_,
		_w8987_,
		_w13983_,
		_w13984_,
		_w13985_
	);
	LUT3 #(
		.INIT('h2a)
	) name12085 (
		\m5_addr_i[12]_pad ,
		_w8989_,
		_w8990_,
		_w13986_
	);
	LUT3 #(
		.INIT('h80)
	) name12086 (
		\m2_addr_i[12]_pad ,
		_w8989_,
		_w8990_,
		_w13987_
	);
	LUT4 #(
		.INIT('h9bdf)
	) name12087 (
		_w8984_,
		_w8987_,
		_w13986_,
		_w13987_,
		_w13988_
	);
	LUT3 #(
		.INIT('h80)
	) name12088 (
		\m0_addr_i[12]_pad ,
		_w8989_,
		_w8990_,
		_w13989_
	);
	LUT3 #(
		.INIT('h2a)
	) name12089 (
		\m1_addr_i[12]_pad ,
		_w8989_,
		_w8990_,
		_w13990_
	);
	LUT3 #(
		.INIT('h57)
	) name12090 (
		_w9008_,
		_w13989_,
		_w13990_,
		_w13991_
	);
	LUT4 #(
		.INIT('h7fff)
	) name12091 (
		_w13982_,
		_w13985_,
		_w13988_,
		_w13991_,
		_w13992_
	);
	LUT3 #(
		.INIT('h80)
	) name12092 (
		\m6_addr_i[13]_pad ,
		_w8989_,
		_w8990_,
		_w13993_
	);
	LUT3 #(
		.INIT('h2a)
	) name12093 (
		\m7_addr_i[13]_pad ,
		_w8989_,
		_w8990_,
		_w13994_
	);
	LUT3 #(
		.INIT('h57)
	) name12094 (
		_w8988_,
		_w13993_,
		_w13994_,
		_w13995_
	);
	LUT3 #(
		.INIT('h80)
	) name12095 (
		\m4_addr_i[13]_pad ,
		_w8989_,
		_w8990_,
		_w13996_
	);
	LUT3 #(
		.INIT('h2a)
	) name12096 (
		\m1_addr_i[13]_pad ,
		_w8989_,
		_w8990_,
		_w13997_
	);
	LUT4 #(
		.INIT('h57df)
	) name12097 (
		_w8984_,
		_w8987_,
		_w13996_,
		_w13997_,
		_w13998_
	);
	LUT3 #(
		.INIT('h2a)
	) name12098 (
		\m5_addr_i[13]_pad ,
		_w8989_,
		_w8990_,
		_w13999_
	);
	LUT3 #(
		.INIT('h80)
	) name12099 (
		\m0_addr_i[13]_pad ,
		_w8989_,
		_w8990_,
		_w14000_
	);
	LUT4 #(
		.INIT('h57df)
	) name12100 (
		_w8984_,
		_w8987_,
		_w13999_,
		_w14000_,
		_w14001_
	);
	LUT3 #(
		.INIT('h80)
	) name12101 (
		\m2_addr_i[13]_pad ,
		_w8989_,
		_w8990_,
		_w14002_
	);
	LUT3 #(
		.INIT('h2a)
	) name12102 (
		\m3_addr_i[13]_pad ,
		_w8989_,
		_w8990_,
		_w14003_
	);
	LUT3 #(
		.INIT('h57)
	) name12103 (
		_w9002_,
		_w14002_,
		_w14003_,
		_w14004_
	);
	LUT4 #(
		.INIT('h7fff)
	) name12104 (
		_w13995_,
		_w13998_,
		_w14001_,
		_w14004_,
		_w14005_
	);
	LUT3 #(
		.INIT('h80)
	) name12105 (
		\m4_addr_i[14]_pad ,
		_w8989_,
		_w8990_,
		_w14006_
	);
	LUT3 #(
		.INIT('h2a)
	) name12106 (
		\m5_addr_i[14]_pad ,
		_w8989_,
		_w8990_,
		_w14007_
	);
	LUT3 #(
		.INIT('h57)
	) name12107 (
		_w8996_,
		_w14006_,
		_w14007_,
		_w14008_
	);
	LUT3 #(
		.INIT('h80)
	) name12108 (
		\m6_addr_i[14]_pad ,
		_w8989_,
		_w8990_,
		_w14009_
	);
	LUT3 #(
		.INIT('h2a)
	) name12109 (
		\m1_addr_i[14]_pad ,
		_w8989_,
		_w8990_,
		_w14010_
	);
	LUT4 #(
		.INIT('h67ef)
	) name12110 (
		_w8984_,
		_w8987_,
		_w14009_,
		_w14010_,
		_w14011_
	);
	LUT3 #(
		.INIT('h2a)
	) name12111 (
		\m7_addr_i[14]_pad ,
		_w8989_,
		_w8990_,
		_w14012_
	);
	LUT3 #(
		.INIT('h80)
	) name12112 (
		\m0_addr_i[14]_pad ,
		_w8989_,
		_w8990_,
		_w14013_
	);
	LUT4 #(
		.INIT('h67ef)
	) name12113 (
		_w8984_,
		_w8987_,
		_w14012_,
		_w14013_,
		_w14014_
	);
	LUT3 #(
		.INIT('h80)
	) name12114 (
		\m2_addr_i[14]_pad ,
		_w8989_,
		_w8990_,
		_w14015_
	);
	LUT3 #(
		.INIT('h2a)
	) name12115 (
		\m3_addr_i[14]_pad ,
		_w8989_,
		_w8990_,
		_w14016_
	);
	LUT3 #(
		.INIT('h57)
	) name12116 (
		_w9002_,
		_w14015_,
		_w14016_,
		_w14017_
	);
	LUT4 #(
		.INIT('h7fff)
	) name12117 (
		_w14008_,
		_w14011_,
		_w14014_,
		_w14017_,
		_w14018_
	);
	LUT3 #(
		.INIT('h80)
	) name12118 (
		\m2_addr_i[15]_pad ,
		_w8989_,
		_w8990_,
		_w14019_
	);
	LUT3 #(
		.INIT('h2a)
	) name12119 (
		\m3_addr_i[15]_pad ,
		_w8989_,
		_w8990_,
		_w14020_
	);
	LUT3 #(
		.INIT('h57)
	) name12120 (
		_w9002_,
		_w14019_,
		_w14020_,
		_w14021_
	);
	LUT3 #(
		.INIT('h80)
	) name12121 (
		\m0_addr_i[15]_pad ,
		_w8989_,
		_w8990_,
		_w14022_
	);
	LUT3 #(
		.INIT('h2a)
	) name12122 (
		\m7_addr_i[15]_pad ,
		_w8989_,
		_w8990_,
		_w14023_
	);
	LUT4 #(
		.INIT('h6e7f)
	) name12123 (
		_w8984_,
		_w8987_,
		_w14022_,
		_w14023_,
		_w14024_
	);
	LUT3 #(
		.INIT('h2a)
	) name12124 (
		\m1_addr_i[15]_pad ,
		_w8989_,
		_w8990_,
		_w14025_
	);
	LUT3 #(
		.INIT('h80)
	) name12125 (
		\m6_addr_i[15]_pad ,
		_w8989_,
		_w8990_,
		_w14026_
	);
	LUT4 #(
		.INIT('h6e7f)
	) name12126 (
		_w8984_,
		_w8987_,
		_w14025_,
		_w14026_,
		_w14027_
	);
	LUT3 #(
		.INIT('h80)
	) name12127 (
		\m4_addr_i[15]_pad ,
		_w8989_,
		_w8990_,
		_w14028_
	);
	LUT3 #(
		.INIT('h2a)
	) name12128 (
		\m5_addr_i[15]_pad ,
		_w8989_,
		_w8990_,
		_w14029_
	);
	LUT3 #(
		.INIT('h57)
	) name12129 (
		_w8996_,
		_w14028_,
		_w14029_,
		_w14030_
	);
	LUT4 #(
		.INIT('h7fff)
	) name12130 (
		_w14021_,
		_w14024_,
		_w14027_,
		_w14030_,
		_w14031_
	);
	LUT3 #(
		.INIT('h80)
	) name12131 (
		\m0_addr_i[16]_pad ,
		_w8989_,
		_w8990_,
		_w14032_
	);
	LUT3 #(
		.INIT('h2a)
	) name12132 (
		\m1_addr_i[16]_pad ,
		_w8989_,
		_w8990_,
		_w14033_
	);
	LUT3 #(
		.INIT('h57)
	) name12133 (
		_w9008_,
		_w14032_,
		_w14033_,
		_w14034_
	);
	LUT3 #(
		.INIT('h80)
	) name12134 (
		\m4_addr_i[16]_pad ,
		_w8989_,
		_w8990_,
		_w14035_
	);
	LUT3 #(
		.INIT('h2a)
	) name12135 (
		\m3_addr_i[16]_pad ,
		_w8989_,
		_w8990_,
		_w14036_
	);
	LUT4 #(
		.INIT('h9bdf)
	) name12136 (
		_w8984_,
		_w8987_,
		_w14035_,
		_w14036_,
		_w14037_
	);
	LUT3 #(
		.INIT('h2a)
	) name12137 (
		\m5_addr_i[16]_pad ,
		_w8989_,
		_w8990_,
		_w14038_
	);
	LUT3 #(
		.INIT('h80)
	) name12138 (
		\m2_addr_i[16]_pad ,
		_w8989_,
		_w8990_,
		_w14039_
	);
	LUT4 #(
		.INIT('h9bdf)
	) name12139 (
		_w8984_,
		_w8987_,
		_w14038_,
		_w14039_,
		_w14040_
	);
	LUT3 #(
		.INIT('h80)
	) name12140 (
		\m6_addr_i[16]_pad ,
		_w8989_,
		_w8990_,
		_w14041_
	);
	LUT3 #(
		.INIT('h2a)
	) name12141 (
		\m7_addr_i[16]_pad ,
		_w8989_,
		_w8990_,
		_w14042_
	);
	LUT3 #(
		.INIT('h57)
	) name12142 (
		_w8988_,
		_w14041_,
		_w14042_,
		_w14043_
	);
	LUT4 #(
		.INIT('h7fff)
	) name12143 (
		_w14034_,
		_w14037_,
		_w14040_,
		_w14043_,
		_w14044_
	);
	LUT3 #(
		.INIT('h80)
	) name12144 (
		\m4_addr_i[17]_pad ,
		_w8989_,
		_w8990_,
		_w14045_
	);
	LUT3 #(
		.INIT('h2a)
	) name12145 (
		\m5_addr_i[17]_pad ,
		_w8989_,
		_w8990_,
		_w14046_
	);
	LUT3 #(
		.INIT('h57)
	) name12146 (
		_w8996_,
		_w14045_,
		_w14046_,
		_w14047_
	);
	LUT3 #(
		.INIT('h80)
	) name12147 (
		\m0_addr_i[17]_pad ,
		_w8989_,
		_w8990_,
		_w14048_
	);
	LUT3 #(
		.INIT('h2a)
	) name12148 (
		\m3_addr_i[17]_pad ,
		_w8989_,
		_w8990_,
		_w14049_
	);
	LUT4 #(
		.INIT('h3b7f)
	) name12149 (
		_w8984_,
		_w8987_,
		_w14048_,
		_w14049_,
		_w14050_
	);
	LUT3 #(
		.INIT('h2a)
	) name12150 (
		\m1_addr_i[17]_pad ,
		_w8989_,
		_w8990_,
		_w14051_
	);
	LUT3 #(
		.INIT('h80)
	) name12151 (
		\m2_addr_i[17]_pad ,
		_w8989_,
		_w8990_,
		_w14052_
	);
	LUT4 #(
		.INIT('h3b7f)
	) name12152 (
		_w8984_,
		_w8987_,
		_w14051_,
		_w14052_,
		_w14053_
	);
	LUT3 #(
		.INIT('h80)
	) name12153 (
		\m6_addr_i[17]_pad ,
		_w8989_,
		_w8990_,
		_w14054_
	);
	LUT3 #(
		.INIT('h2a)
	) name12154 (
		\m7_addr_i[17]_pad ,
		_w8989_,
		_w8990_,
		_w14055_
	);
	LUT3 #(
		.INIT('h57)
	) name12155 (
		_w8988_,
		_w14054_,
		_w14055_,
		_w14056_
	);
	LUT4 #(
		.INIT('h7fff)
	) name12156 (
		_w14047_,
		_w14050_,
		_w14053_,
		_w14056_,
		_w14057_
	);
	LUT3 #(
		.INIT('h80)
	) name12157 (
		\m2_addr_i[18]_pad ,
		_w8989_,
		_w8990_,
		_w14058_
	);
	LUT3 #(
		.INIT('h2a)
	) name12158 (
		\m3_addr_i[18]_pad ,
		_w8989_,
		_w8990_,
		_w14059_
	);
	LUT3 #(
		.INIT('h57)
	) name12159 (
		_w9002_,
		_w14058_,
		_w14059_,
		_w14060_
	);
	LUT3 #(
		.INIT('h80)
	) name12160 (
		\m0_addr_i[18]_pad ,
		_w8989_,
		_w8990_,
		_w14061_
	);
	LUT3 #(
		.INIT('h2a)
	) name12161 (
		\m5_addr_i[18]_pad ,
		_w8989_,
		_w8990_,
		_w14062_
	);
	LUT4 #(
		.INIT('h5d7f)
	) name12162 (
		_w8984_,
		_w8987_,
		_w14061_,
		_w14062_,
		_w14063_
	);
	LUT3 #(
		.INIT('h2a)
	) name12163 (
		\m1_addr_i[18]_pad ,
		_w8989_,
		_w8990_,
		_w14064_
	);
	LUT3 #(
		.INIT('h80)
	) name12164 (
		\m4_addr_i[18]_pad ,
		_w8989_,
		_w8990_,
		_w14065_
	);
	LUT4 #(
		.INIT('h5d7f)
	) name12165 (
		_w8984_,
		_w8987_,
		_w14064_,
		_w14065_,
		_w14066_
	);
	LUT3 #(
		.INIT('h80)
	) name12166 (
		\m6_addr_i[18]_pad ,
		_w8989_,
		_w8990_,
		_w14067_
	);
	LUT3 #(
		.INIT('h2a)
	) name12167 (
		\m7_addr_i[18]_pad ,
		_w8989_,
		_w8990_,
		_w14068_
	);
	LUT3 #(
		.INIT('h57)
	) name12168 (
		_w8988_,
		_w14067_,
		_w14068_,
		_w14069_
	);
	LUT4 #(
		.INIT('h7fff)
	) name12169 (
		_w14060_,
		_w14063_,
		_w14066_,
		_w14069_,
		_w14070_
	);
	LUT3 #(
		.INIT('h80)
	) name12170 (
		\m2_addr_i[19]_pad ,
		_w8989_,
		_w8990_,
		_w14071_
	);
	LUT3 #(
		.INIT('h2a)
	) name12171 (
		\m3_addr_i[19]_pad ,
		_w8989_,
		_w8990_,
		_w14072_
	);
	LUT3 #(
		.INIT('h57)
	) name12172 (
		_w9002_,
		_w14071_,
		_w14072_,
		_w14073_
	);
	LUT3 #(
		.INIT('h80)
	) name12173 (
		\m4_addr_i[19]_pad ,
		_w8989_,
		_w8990_,
		_w14074_
	);
	LUT3 #(
		.INIT('h2a)
	) name12174 (
		\m1_addr_i[19]_pad ,
		_w8989_,
		_w8990_,
		_w14075_
	);
	LUT4 #(
		.INIT('h57df)
	) name12175 (
		_w8984_,
		_w8987_,
		_w14074_,
		_w14075_,
		_w14076_
	);
	LUT3 #(
		.INIT('h2a)
	) name12176 (
		\m5_addr_i[19]_pad ,
		_w8989_,
		_w8990_,
		_w14077_
	);
	LUT3 #(
		.INIT('h80)
	) name12177 (
		\m0_addr_i[19]_pad ,
		_w8989_,
		_w8990_,
		_w14078_
	);
	LUT4 #(
		.INIT('h57df)
	) name12178 (
		_w8984_,
		_w8987_,
		_w14077_,
		_w14078_,
		_w14079_
	);
	LUT3 #(
		.INIT('h80)
	) name12179 (
		\m6_addr_i[19]_pad ,
		_w8989_,
		_w8990_,
		_w14080_
	);
	LUT3 #(
		.INIT('h2a)
	) name12180 (
		\m7_addr_i[19]_pad ,
		_w8989_,
		_w8990_,
		_w14081_
	);
	LUT3 #(
		.INIT('h57)
	) name12181 (
		_w8988_,
		_w14080_,
		_w14081_,
		_w14082_
	);
	LUT4 #(
		.INIT('h7fff)
	) name12182 (
		_w14073_,
		_w14076_,
		_w14079_,
		_w14082_,
		_w14083_
	);
	LUT3 #(
		.INIT('h80)
	) name12183 (
		\m0_addr_i[1]_pad ,
		_w8989_,
		_w8990_,
		_w14084_
	);
	LUT3 #(
		.INIT('h2a)
	) name12184 (
		\m1_addr_i[1]_pad ,
		_w8989_,
		_w8990_,
		_w14085_
	);
	LUT3 #(
		.INIT('h57)
	) name12185 (
		_w9008_,
		_w14084_,
		_w14085_,
		_w14086_
	);
	LUT3 #(
		.INIT('h80)
	) name12186 (
		\m6_addr_i[1]_pad ,
		_w8989_,
		_w8990_,
		_w14087_
	);
	LUT3 #(
		.INIT('h2a)
	) name12187 (
		\m3_addr_i[1]_pad ,
		_w8989_,
		_w8990_,
		_w14088_
	);
	LUT4 #(
		.INIT('habef)
	) name12188 (
		_w8984_,
		_w8987_,
		_w14087_,
		_w14088_,
		_w14089_
	);
	LUT3 #(
		.INIT('h2a)
	) name12189 (
		\m7_addr_i[1]_pad ,
		_w8989_,
		_w8990_,
		_w14090_
	);
	LUT3 #(
		.INIT('h80)
	) name12190 (
		\m2_addr_i[1]_pad ,
		_w8989_,
		_w8990_,
		_w14091_
	);
	LUT4 #(
		.INIT('habef)
	) name12191 (
		_w8984_,
		_w8987_,
		_w14090_,
		_w14091_,
		_w14092_
	);
	LUT3 #(
		.INIT('h80)
	) name12192 (
		\m4_addr_i[1]_pad ,
		_w8989_,
		_w8990_,
		_w14093_
	);
	LUT3 #(
		.INIT('h2a)
	) name12193 (
		\m5_addr_i[1]_pad ,
		_w8989_,
		_w8990_,
		_w14094_
	);
	LUT3 #(
		.INIT('h57)
	) name12194 (
		_w8996_,
		_w14093_,
		_w14094_,
		_w14095_
	);
	LUT4 #(
		.INIT('h7fff)
	) name12195 (
		_w14086_,
		_w14089_,
		_w14092_,
		_w14095_,
		_w14096_
	);
	LUT3 #(
		.INIT('h80)
	) name12196 (
		\m6_addr_i[20]_pad ,
		_w8989_,
		_w8990_,
		_w14097_
	);
	LUT3 #(
		.INIT('h2a)
	) name12197 (
		\m7_addr_i[20]_pad ,
		_w8989_,
		_w8990_,
		_w14098_
	);
	LUT3 #(
		.INIT('h57)
	) name12198 (
		_w8988_,
		_w14097_,
		_w14098_,
		_w14099_
	);
	LUT3 #(
		.INIT('h80)
	) name12199 (
		\m4_addr_i[20]_pad ,
		_w8989_,
		_w8990_,
		_w14100_
	);
	LUT3 #(
		.INIT('h2a)
	) name12200 (
		\m1_addr_i[20]_pad ,
		_w8989_,
		_w8990_,
		_w14101_
	);
	LUT4 #(
		.INIT('h57df)
	) name12201 (
		_w8984_,
		_w8987_,
		_w14100_,
		_w14101_,
		_w14102_
	);
	LUT3 #(
		.INIT('h2a)
	) name12202 (
		\m5_addr_i[20]_pad ,
		_w8989_,
		_w8990_,
		_w14103_
	);
	LUT3 #(
		.INIT('h80)
	) name12203 (
		\m0_addr_i[20]_pad ,
		_w8989_,
		_w8990_,
		_w14104_
	);
	LUT4 #(
		.INIT('h57df)
	) name12204 (
		_w8984_,
		_w8987_,
		_w14103_,
		_w14104_,
		_w14105_
	);
	LUT3 #(
		.INIT('h80)
	) name12205 (
		\m2_addr_i[20]_pad ,
		_w8989_,
		_w8990_,
		_w14106_
	);
	LUT3 #(
		.INIT('h2a)
	) name12206 (
		\m3_addr_i[20]_pad ,
		_w8989_,
		_w8990_,
		_w14107_
	);
	LUT3 #(
		.INIT('h57)
	) name12207 (
		_w9002_,
		_w14106_,
		_w14107_,
		_w14108_
	);
	LUT4 #(
		.INIT('h7fff)
	) name12208 (
		_w14099_,
		_w14102_,
		_w14105_,
		_w14108_,
		_w14109_
	);
	LUT3 #(
		.INIT('h80)
	) name12209 (
		\m6_addr_i[21]_pad ,
		_w8989_,
		_w8990_,
		_w14110_
	);
	LUT3 #(
		.INIT('h2a)
	) name12210 (
		\m7_addr_i[21]_pad ,
		_w8989_,
		_w8990_,
		_w14111_
	);
	LUT3 #(
		.INIT('h57)
	) name12211 (
		_w8988_,
		_w14110_,
		_w14111_,
		_w14112_
	);
	LUT3 #(
		.INIT('h80)
	) name12212 (
		\m0_addr_i[21]_pad ,
		_w8989_,
		_w8990_,
		_w14113_
	);
	LUT3 #(
		.INIT('h2a)
	) name12213 (
		\m3_addr_i[21]_pad ,
		_w8989_,
		_w8990_,
		_w14114_
	);
	LUT4 #(
		.INIT('h3b7f)
	) name12214 (
		_w8984_,
		_w8987_,
		_w14113_,
		_w14114_,
		_w14115_
	);
	LUT3 #(
		.INIT('h2a)
	) name12215 (
		\m1_addr_i[21]_pad ,
		_w8989_,
		_w8990_,
		_w14116_
	);
	LUT3 #(
		.INIT('h80)
	) name12216 (
		\m2_addr_i[21]_pad ,
		_w8989_,
		_w8990_,
		_w14117_
	);
	LUT4 #(
		.INIT('h3b7f)
	) name12217 (
		_w8984_,
		_w8987_,
		_w14116_,
		_w14117_,
		_w14118_
	);
	LUT3 #(
		.INIT('h80)
	) name12218 (
		\m4_addr_i[21]_pad ,
		_w8989_,
		_w8990_,
		_w14119_
	);
	LUT3 #(
		.INIT('h2a)
	) name12219 (
		\m5_addr_i[21]_pad ,
		_w8989_,
		_w8990_,
		_w14120_
	);
	LUT3 #(
		.INIT('h57)
	) name12220 (
		_w8996_,
		_w14119_,
		_w14120_,
		_w14121_
	);
	LUT4 #(
		.INIT('h7fff)
	) name12221 (
		_w14112_,
		_w14115_,
		_w14118_,
		_w14121_,
		_w14122_
	);
	LUT3 #(
		.INIT('h80)
	) name12222 (
		\m6_addr_i[22]_pad ,
		_w8989_,
		_w8990_,
		_w14123_
	);
	LUT3 #(
		.INIT('h2a)
	) name12223 (
		\m7_addr_i[22]_pad ,
		_w8989_,
		_w8990_,
		_w14124_
	);
	LUT3 #(
		.INIT('h57)
	) name12224 (
		_w8988_,
		_w14123_,
		_w14124_,
		_w14125_
	);
	LUT3 #(
		.INIT('h80)
	) name12225 (
		\m2_addr_i[22]_pad ,
		_w8989_,
		_w8990_,
		_w14126_
	);
	LUT3 #(
		.INIT('h2a)
	) name12226 (
		\m1_addr_i[22]_pad ,
		_w8989_,
		_w8990_,
		_w14127_
	);
	LUT4 #(
		.INIT('h37bf)
	) name12227 (
		_w8984_,
		_w8987_,
		_w14126_,
		_w14127_,
		_w14128_
	);
	LUT3 #(
		.INIT('h2a)
	) name12228 (
		\m3_addr_i[22]_pad ,
		_w8989_,
		_w8990_,
		_w14129_
	);
	LUT3 #(
		.INIT('h80)
	) name12229 (
		\m0_addr_i[22]_pad ,
		_w8989_,
		_w8990_,
		_w14130_
	);
	LUT4 #(
		.INIT('h37bf)
	) name12230 (
		_w8984_,
		_w8987_,
		_w14129_,
		_w14130_,
		_w14131_
	);
	LUT3 #(
		.INIT('h80)
	) name12231 (
		\m4_addr_i[22]_pad ,
		_w8989_,
		_w8990_,
		_w14132_
	);
	LUT3 #(
		.INIT('h2a)
	) name12232 (
		\m5_addr_i[22]_pad ,
		_w8989_,
		_w8990_,
		_w14133_
	);
	LUT3 #(
		.INIT('h57)
	) name12233 (
		_w8996_,
		_w14132_,
		_w14133_,
		_w14134_
	);
	LUT4 #(
		.INIT('h7fff)
	) name12234 (
		_w14125_,
		_w14128_,
		_w14131_,
		_w14134_,
		_w14135_
	);
	LUT3 #(
		.INIT('h80)
	) name12235 (
		\m4_addr_i[23]_pad ,
		_w8989_,
		_w8990_,
		_w14136_
	);
	LUT3 #(
		.INIT('h2a)
	) name12236 (
		\m5_addr_i[23]_pad ,
		_w8989_,
		_w8990_,
		_w14137_
	);
	LUT3 #(
		.INIT('h57)
	) name12237 (
		_w8996_,
		_w14136_,
		_w14137_,
		_w14138_
	);
	LUT3 #(
		.INIT('h80)
	) name12238 (
		\m0_addr_i[23]_pad ,
		_w8989_,
		_w8990_,
		_w14139_
	);
	LUT3 #(
		.INIT('h2a)
	) name12239 (
		\m7_addr_i[23]_pad ,
		_w8989_,
		_w8990_,
		_w14140_
	);
	LUT4 #(
		.INIT('h6e7f)
	) name12240 (
		_w8984_,
		_w8987_,
		_w14139_,
		_w14140_,
		_w14141_
	);
	LUT3 #(
		.INIT('h2a)
	) name12241 (
		\m1_addr_i[23]_pad ,
		_w8989_,
		_w8990_,
		_w14142_
	);
	LUT3 #(
		.INIT('h80)
	) name12242 (
		\m6_addr_i[23]_pad ,
		_w8989_,
		_w8990_,
		_w14143_
	);
	LUT4 #(
		.INIT('h6e7f)
	) name12243 (
		_w8984_,
		_w8987_,
		_w14142_,
		_w14143_,
		_w14144_
	);
	LUT3 #(
		.INIT('h80)
	) name12244 (
		\m2_addr_i[23]_pad ,
		_w8989_,
		_w8990_,
		_w14145_
	);
	LUT3 #(
		.INIT('h2a)
	) name12245 (
		\m3_addr_i[23]_pad ,
		_w8989_,
		_w8990_,
		_w14146_
	);
	LUT3 #(
		.INIT('h57)
	) name12246 (
		_w9002_,
		_w14145_,
		_w14146_,
		_w14147_
	);
	LUT4 #(
		.INIT('h7fff)
	) name12247 (
		_w14138_,
		_w14141_,
		_w14144_,
		_w14147_,
		_w14148_
	);
	LUT3 #(
		.INIT('h80)
	) name12248 (
		\m0_addr_i[24]_pad ,
		_w8989_,
		_w8990_,
		_w14149_
	);
	LUT3 #(
		.INIT('h2a)
	) name12249 (
		\m7_addr_i[24]_pad ,
		_w8989_,
		_w8990_,
		_w14150_
	);
	LUT4 #(
		.INIT('h6e7f)
	) name12250 (
		_w8984_,
		_w8987_,
		_w14149_,
		_w14150_,
		_w14151_
	);
	LUT3 #(
		.INIT('h2a)
	) name12251 (
		\m1_addr_i[24]_pad ,
		_w8989_,
		_w8990_,
		_w14152_
	);
	LUT3 #(
		.INIT('h80)
	) name12252 (
		\m4_addr_i[24]_pad ,
		_w8989_,
		_w8990_,
		_w14153_
	);
	LUT4 #(
		.INIT('h5d7f)
	) name12253 (
		_w8984_,
		_w8987_,
		_w14152_,
		_w14153_,
		_w14154_
	);
	LUT3 #(
		.INIT('h80)
	) name12254 (
		\m2_addr_i[24]_pad ,
		_w8989_,
		_w8990_,
		_w14155_
	);
	LUT3 #(
		.INIT('h2a)
	) name12255 (
		\m3_addr_i[24]_pad ,
		_w8989_,
		_w8990_,
		_w14156_
	);
	LUT3 #(
		.INIT('h57)
	) name12256 (
		_w9002_,
		_w14155_,
		_w14156_,
		_w14157_
	);
	LUT3 #(
		.INIT('h2a)
	) name12257 (
		\m5_addr_i[24]_pad ,
		_w8989_,
		_w8990_,
		_w14158_
	);
	LUT3 #(
		.INIT('h80)
	) name12258 (
		\m6_addr_i[24]_pad ,
		_w8989_,
		_w8990_,
		_w14159_
	);
	LUT4 #(
		.INIT('hcedf)
	) name12259 (
		_w8984_,
		_w8987_,
		_w14158_,
		_w14159_,
		_w14160_
	);
	LUT4 #(
		.INIT('h7fff)
	) name12260 (
		_w14151_,
		_w14154_,
		_w14157_,
		_w14160_,
		_w14161_
	);
	LUT3 #(
		.INIT('h80)
	) name12261 (
		\m0_addr_i[25]_pad ,
		_w8989_,
		_w8990_,
		_w14162_
	);
	LUT3 #(
		.INIT('h2a)
	) name12262 (
		\m7_addr_i[25]_pad ,
		_w8989_,
		_w8990_,
		_w14163_
	);
	LUT4 #(
		.INIT('h6e7f)
	) name12263 (
		_w8984_,
		_w8987_,
		_w14162_,
		_w14163_,
		_w14164_
	);
	LUT3 #(
		.INIT('h2a)
	) name12264 (
		\m1_addr_i[25]_pad ,
		_w8989_,
		_w8990_,
		_w14165_
	);
	LUT3 #(
		.INIT('h80)
	) name12265 (
		\m4_addr_i[25]_pad ,
		_w8989_,
		_w8990_,
		_w14166_
	);
	LUT4 #(
		.INIT('h5d7f)
	) name12266 (
		_w8984_,
		_w8987_,
		_w14165_,
		_w14166_,
		_w14167_
	);
	LUT3 #(
		.INIT('h80)
	) name12267 (
		\m2_addr_i[25]_pad ,
		_w8989_,
		_w8990_,
		_w14168_
	);
	LUT3 #(
		.INIT('h2a)
	) name12268 (
		\m3_addr_i[25]_pad ,
		_w8989_,
		_w8990_,
		_w14169_
	);
	LUT3 #(
		.INIT('h57)
	) name12269 (
		_w9002_,
		_w14168_,
		_w14169_,
		_w14170_
	);
	LUT3 #(
		.INIT('h2a)
	) name12270 (
		\m5_addr_i[25]_pad ,
		_w8989_,
		_w8990_,
		_w14171_
	);
	LUT3 #(
		.INIT('h80)
	) name12271 (
		\m6_addr_i[25]_pad ,
		_w8989_,
		_w8990_,
		_w14172_
	);
	LUT4 #(
		.INIT('hcedf)
	) name12272 (
		_w8984_,
		_w8987_,
		_w14171_,
		_w14172_,
		_w14173_
	);
	LUT4 #(
		.INIT('h7fff)
	) name12273 (
		_w14164_,
		_w14167_,
		_w14170_,
		_w14173_,
		_w14174_
	);
	LUT3 #(
		.INIT('h2a)
	) name12274 (
		\m1_addr_i[26]_pad ,
		_w8989_,
		_w8990_,
		_w14175_
	);
	LUT3 #(
		.INIT('h80)
	) name12275 (
		\m2_addr_i[26]_pad ,
		_w8989_,
		_w8990_,
		_w14176_
	);
	LUT4 #(
		.INIT('h3b7f)
	) name12276 (
		_w8984_,
		_w8987_,
		_w14175_,
		_w14176_,
		_w14177_
	);
	LUT3 #(
		.INIT('h80)
	) name12277 (
		\m0_addr_i[26]_pad ,
		_w8989_,
		_w8990_,
		_w14178_
	);
	LUT3 #(
		.INIT('h80)
	) name12278 (
		\m4_addr_i[26]_pad ,
		_w8989_,
		_w8990_,
		_w14179_
	);
	LUT4 #(
		.INIT('h5d7f)
	) name12279 (
		_w8984_,
		_w8987_,
		_w14178_,
		_w14179_,
		_w14180_
	);
	LUT3 #(
		.INIT('h2a)
	) name12280 (
		\m7_addr_i[26]_pad ,
		_w8989_,
		_w8990_,
		_w14181_
	);
	LUT3 #(
		.INIT('h2a)
	) name12281 (
		\m3_addr_i[26]_pad ,
		_w8989_,
		_w8990_,
		_w14182_
	);
	LUT4 #(
		.INIT('habef)
	) name12282 (
		_w8984_,
		_w8987_,
		_w14181_,
		_w14182_,
		_w14183_
	);
	LUT3 #(
		.INIT('h2a)
	) name12283 (
		\m5_addr_i[26]_pad ,
		_w8989_,
		_w8990_,
		_w14184_
	);
	LUT3 #(
		.INIT('h80)
	) name12284 (
		\m6_addr_i[26]_pad ,
		_w8989_,
		_w8990_,
		_w14185_
	);
	LUT4 #(
		.INIT('hcedf)
	) name12285 (
		_w8984_,
		_w8987_,
		_w14184_,
		_w14185_,
		_w14186_
	);
	LUT4 #(
		.INIT('h7fff)
	) name12286 (
		_w14177_,
		_w14180_,
		_w14183_,
		_w14186_,
		_w14187_
	);
	LUT3 #(
		.INIT('h2a)
	) name12287 (
		\m1_addr_i[27]_pad ,
		_w8989_,
		_w8990_,
		_w14188_
	);
	LUT3 #(
		.INIT('h80)
	) name12288 (
		\m2_addr_i[27]_pad ,
		_w8989_,
		_w8990_,
		_w14189_
	);
	LUT4 #(
		.INIT('h3b7f)
	) name12289 (
		_w8984_,
		_w8987_,
		_w14188_,
		_w14189_,
		_w14190_
	);
	LUT3 #(
		.INIT('h80)
	) name12290 (
		\m0_addr_i[27]_pad ,
		_w8989_,
		_w8990_,
		_w14191_
	);
	LUT3 #(
		.INIT('h80)
	) name12291 (
		\m6_addr_i[27]_pad ,
		_w8989_,
		_w8990_,
		_w14192_
	);
	LUT4 #(
		.INIT('h6e7f)
	) name12292 (
		_w8984_,
		_w8987_,
		_w14191_,
		_w14192_,
		_w14193_
	);
	LUT3 #(
		.INIT('h2a)
	) name12293 (
		\m7_addr_i[27]_pad ,
		_w8989_,
		_w8990_,
		_w14194_
	);
	LUT3 #(
		.INIT('h2a)
	) name12294 (
		\m5_addr_i[27]_pad ,
		_w8989_,
		_w8990_,
		_w14195_
	);
	LUT4 #(
		.INIT('hcdef)
	) name12295 (
		_w8984_,
		_w8987_,
		_w14194_,
		_w14195_,
		_w14196_
	);
	LUT3 #(
		.INIT('h2a)
	) name12296 (
		\m3_addr_i[27]_pad ,
		_w8989_,
		_w8990_,
		_w14197_
	);
	LUT3 #(
		.INIT('h80)
	) name12297 (
		\m4_addr_i[27]_pad ,
		_w8989_,
		_w8990_,
		_w14198_
	);
	LUT4 #(
		.INIT('h9dbf)
	) name12298 (
		_w8984_,
		_w8987_,
		_w14197_,
		_w14198_,
		_w14199_
	);
	LUT4 #(
		.INIT('h7fff)
	) name12299 (
		_w14190_,
		_w14193_,
		_w14196_,
		_w14199_,
		_w14200_
	);
	LUT3 #(
		.INIT('h2a)
	) name12300 (
		\m1_addr_i[28]_pad ,
		_w8989_,
		_w8990_,
		_w14201_
	);
	LUT3 #(
		.INIT('h80)
	) name12301 (
		\m2_addr_i[28]_pad ,
		_w8989_,
		_w8990_,
		_w14202_
	);
	LUT4 #(
		.INIT('h3b7f)
	) name12302 (
		_w8984_,
		_w8987_,
		_w14201_,
		_w14202_,
		_w14203_
	);
	LUT3 #(
		.INIT('h2a)
	) name12303 (
		\m5_addr_i[28]_pad ,
		_w8989_,
		_w8990_,
		_w14204_
	);
	LUT3 #(
		.INIT('h80)
	) name12304 (
		\m4_addr_i[28]_pad ,
		_w8989_,
		_w8990_,
		_w14205_
	);
	LUT3 #(
		.INIT('h57)
	) name12305 (
		_w8996_,
		_w14204_,
		_w14205_,
		_w14206_
	);
	LUT3 #(
		.INIT('h80)
	) name12306 (
		\m6_addr_i[28]_pad ,
		_w8989_,
		_w8990_,
		_w14207_
	);
	LUT3 #(
		.INIT('h2a)
	) name12307 (
		\m3_addr_i[28]_pad ,
		_w8989_,
		_w8990_,
		_w14208_
	);
	LUT4 #(
		.INIT('habef)
	) name12308 (
		_w8984_,
		_w8987_,
		_w14207_,
		_w14208_,
		_w14209_
	);
	LUT3 #(
		.INIT('h80)
	) name12309 (
		\m0_addr_i[28]_pad ,
		_w8989_,
		_w8990_,
		_w14210_
	);
	LUT3 #(
		.INIT('h2a)
	) name12310 (
		\m7_addr_i[28]_pad ,
		_w8989_,
		_w8990_,
		_w14211_
	);
	LUT4 #(
		.INIT('h6e7f)
	) name12311 (
		_w8984_,
		_w8987_,
		_w14210_,
		_w14211_,
		_w14212_
	);
	LUT4 #(
		.INIT('h7fff)
	) name12312 (
		_w14203_,
		_w14206_,
		_w14209_,
		_w14212_,
		_w14213_
	);
	LUT3 #(
		.INIT('h2a)
	) name12313 (
		\m3_addr_i[29]_pad ,
		_w8989_,
		_w8990_,
		_w14214_
	);
	LUT3 #(
		.INIT('h80)
	) name12314 (
		\m4_addr_i[29]_pad ,
		_w8989_,
		_w8990_,
		_w14215_
	);
	LUT4 #(
		.INIT('h9dbf)
	) name12315 (
		_w8984_,
		_w8987_,
		_w14214_,
		_w14215_,
		_w14216_
	);
	LUT3 #(
		.INIT('h2a)
	) name12316 (
		\m1_addr_i[29]_pad ,
		_w8989_,
		_w8990_,
		_w14217_
	);
	LUT3 #(
		.INIT('h2a)
	) name12317 (
		\m7_addr_i[29]_pad ,
		_w8989_,
		_w8990_,
		_w14218_
	);
	LUT4 #(
		.INIT('h6e7f)
	) name12318 (
		_w8984_,
		_w8987_,
		_w14217_,
		_w14218_,
		_w14219_
	);
	LUT3 #(
		.INIT('h80)
	) name12319 (
		\m2_addr_i[29]_pad ,
		_w8989_,
		_w8990_,
		_w14220_
	);
	LUT3 #(
		.INIT('h80)
	) name12320 (
		\m0_addr_i[29]_pad ,
		_w8989_,
		_w8990_,
		_w14221_
	);
	LUT4 #(
		.INIT('h37bf)
	) name12321 (
		_w8984_,
		_w8987_,
		_w14220_,
		_w14221_,
		_w14222_
	);
	LUT3 #(
		.INIT('h2a)
	) name12322 (
		\m5_addr_i[29]_pad ,
		_w8989_,
		_w8990_,
		_w14223_
	);
	LUT3 #(
		.INIT('h80)
	) name12323 (
		\m6_addr_i[29]_pad ,
		_w8989_,
		_w8990_,
		_w14224_
	);
	LUT4 #(
		.INIT('hcedf)
	) name12324 (
		_w8984_,
		_w8987_,
		_w14223_,
		_w14224_,
		_w14225_
	);
	LUT4 #(
		.INIT('h7fff)
	) name12325 (
		_w14216_,
		_w14219_,
		_w14222_,
		_w14225_,
		_w14226_
	);
	LUT3 #(
		.INIT('h80)
	) name12326 (
		\m2_addr_i[2]_pad ,
		_w8989_,
		_w8990_,
		_w14227_
	);
	LUT3 #(
		.INIT('h2a)
	) name12327 (
		\m3_addr_i[2]_pad ,
		_w8989_,
		_w8990_,
		_w14228_
	);
	LUT3 #(
		.INIT('h57)
	) name12328 (
		_w9002_,
		_w14227_,
		_w14228_,
		_w14229_
	);
	LUT3 #(
		.INIT('h80)
	) name12329 (
		\m0_addr_i[2]_pad ,
		_w8989_,
		_w8990_,
		_w14230_
	);
	LUT3 #(
		.INIT('h2a)
	) name12330 (
		\m7_addr_i[2]_pad ,
		_w8989_,
		_w8990_,
		_w14231_
	);
	LUT4 #(
		.INIT('h6e7f)
	) name12331 (
		_w8984_,
		_w8987_,
		_w14230_,
		_w14231_,
		_w14232_
	);
	LUT3 #(
		.INIT('h2a)
	) name12332 (
		\m1_addr_i[2]_pad ,
		_w8989_,
		_w8990_,
		_w14233_
	);
	LUT3 #(
		.INIT('h80)
	) name12333 (
		\m6_addr_i[2]_pad ,
		_w8989_,
		_w8990_,
		_w14234_
	);
	LUT4 #(
		.INIT('h6e7f)
	) name12334 (
		_w8984_,
		_w8987_,
		_w14233_,
		_w14234_,
		_w14235_
	);
	LUT3 #(
		.INIT('h80)
	) name12335 (
		\m4_addr_i[2]_pad ,
		_w8989_,
		_w8990_,
		_w14236_
	);
	LUT3 #(
		.INIT('h2a)
	) name12336 (
		\m5_addr_i[2]_pad ,
		_w8989_,
		_w8990_,
		_w14237_
	);
	LUT3 #(
		.INIT('h57)
	) name12337 (
		_w8996_,
		_w14236_,
		_w14237_,
		_w14238_
	);
	LUT4 #(
		.INIT('h7fff)
	) name12338 (
		_w14229_,
		_w14232_,
		_w14235_,
		_w14238_,
		_w14239_
	);
	LUT3 #(
		.INIT('h2a)
	) name12339 (
		\m3_addr_i[30]_pad ,
		_w8989_,
		_w8990_,
		_w14240_
	);
	LUT3 #(
		.INIT('h80)
	) name12340 (
		\m4_addr_i[30]_pad ,
		_w8989_,
		_w8990_,
		_w14241_
	);
	LUT4 #(
		.INIT('h9dbf)
	) name12341 (
		_w8984_,
		_w8987_,
		_w14240_,
		_w14241_,
		_w14242_
	);
	LUT3 #(
		.INIT('h80)
	) name12342 (
		\m0_addr_i[30]_pad ,
		_w8989_,
		_w8990_,
		_w14243_
	);
	LUT3 #(
		.INIT('h80)
	) name12343 (
		\m6_addr_i[30]_pad ,
		_w8989_,
		_w8990_,
		_w14244_
	);
	LUT4 #(
		.INIT('h6e7f)
	) name12344 (
		_w8984_,
		_w8987_,
		_w14243_,
		_w14244_,
		_w14245_
	);
	LUT3 #(
		.INIT('h2a)
	) name12345 (
		\m7_addr_i[30]_pad ,
		_w8989_,
		_w8990_,
		_w14246_
	);
	LUT3 #(
		.INIT('h2a)
	) name12346 (
		\m5_addr_i[30]_pad ,
		_w8989_,
		_w8990_,
		_w14247_
	);
	LUT4 #(
		.INIT('hcdef)
	) name12347 (
		_w8984_,
		_w8987_,
		_w14246_,
		_w14247_,
		_w14248_
	);
	LUT3 #(
		.INIT('h2a)
	) name12348 (
		\m1_addr_i[30]_pad ,
		_w8989_,
		_w8990_,
		_w14249_
	);
	LUT3 #(
		.INIT('h80)
	) name12349 (
		\m2_addr_i[30]_pad ,
		_w8989_,
		_w8990_,
		_w14250_
	);
	LUT4 #(
		.INIT('h3b7f)
	) name12350 (
		_w8984_,
		_w8987_,
		_w14249_,
		_w14250_,
		_w14251_
	);
	LUT4 #(
		.INIT('h7fff)
	) name12351 (
		_w14242_,
		_w14245_,
		_w14248_,
		_w14251_,
		_w14252_
	);
	LUT3 #(
		.INIT('h2a)
	) name12352 (
		\m1_addr_i[31]_pad ,
		_w8989_,
		_w8990_,
		_w14253_
	);
	LUT3 #(
		.INIT('h80)
	) name12353 (
		\m2_addr_i[31]_pad ,
		_w8989_,
		_w8990_,
		_w14254_
	);
	LUT4 #(
		.INIT('h3b7f)
	) name12354 (
		_w8984_,
		_w8987_,
		_w14253_,
		_w14254_,
		_w14255_
	);
	LUT3 #(
		.INIT('h80)
	) name12355 (
		\m0_addr_i[31]_pad ,
		_w8989_,
		_w8990_,
		_w14256_
	);
	LUT3 #(
		.INIT('h80)
	) name12356 (
		\m4_addr_i[31]_pad ,
		_w8989_,
		_w8990_,
		_w14257_
	);
	LUT4 #(
		.INIT('h5d7f)
	) name12357 (
		_w8984_,
		_w8987_,
		_w14256_,
		_w14257_,
		_w14258_
	);
	LUT3 #(
		.INIT('h2a)
	) name12358 (
		\m7_addr_i[31]_pad ,
		_w8989_,
		_w8990_,
		_w14259_
	);
	LUT3 #(
		.INIT('h2a)
	) name12359 (
		\m3_addr_i[31]_pad ,
		_w8989_,
		_w8990_,
		_w14260_
	);
	LUT4 #(
		.INIT('habef)
	) name12360 (
		_w8984_,
		_w8987_,
		_w14259_,
		_w14260_,
		_w14261_
	);
	LUT3 #(
		.INIT('h2a)
	) name12361 (
		\m5_addr_i[31]_pad ,
		_w8989_,
		_w8990_,
		_w14262_
	);
	LUT3 #(
		.INIT('h80)
	) name12362 (
		\m6_addr_i[31]_pad ,
		_w8989_,
		_w8990_,
		_w14263_
	);
	LUT4 #(
		.INIT('hcedf)
	) name12363 (
		_w8984_,
		_w8987_,
		_w14262_,
		_w14263_,
		_w14264_
	);
	LUT4 #(
		.INIT('h7fff)
	) name12364 (
		_w14255_,
		_w14258_,
		_w14261_,
		_w14264_,
		_w14265_
	);
	LUT3 #(
		.INIT('h80)
	) name12365 (
		\m2_addr_i[3]_pad ,
		_w8989_,
		_w8990_,
		_w14266_
	);
	LUT3 #(
		.INIT('h2a)
	) name12366 (
		\m3_addr_i[3]_pad ,
		_w8989_,
		_w8990_,
		_w14267_
	);
	LUT3 #(
		.INIT('h57)
	) name12367 (
		_w9002_,
		_w14266_,
		_w14267_,
		_w14268_
	);
	LUT3 #(
		.INIT('h80)
	) name12368 (
		\m0_addr_i[3]_pad ,
		_w8989_,
		_w8990_,
		_w14269_
	);
	LUT3 #(
		.INIT('h2a)
	) name12369 (
		\m7_addr_i[3]_pad ,
		_w8989_,
		_w8990_,
		_w14270_
	);
	LUT4 #(
		.INIT('h6e7f)
	) name12370 (
		_w8984_,
		_w8987_,
		_w14269_,
		_w14270_,
		_w14271_
	);
	LUT3 #(
		.INIT('h2a)
	) name12371 (
		\m1_addr_i[3]_pad ,
		_w8989_,
		_w8990_,
		_w14272_
	);
	LUT3 #(
		.INIT('h80)
	) name12372 (
		\m6_addr_i[3]_pad ,
		_w8989_,
		_w8990_,
		_w14273_
	);
	LUT4 #(
		.INIT('h6e7f)
	) name12373 (
		_w8984_,
		_w8987_,
		_w14272_,
		_w14273_,
		_w14274_
	);
	LUT3 #(
		.INIT('h80)
	) name12374 (
		\m4_addr_i[3]_pad ,
		_w8989_,
		_w8990_,
		_w14275_
	);
	LUT3 #(
		.INIT('h2a)
	) name12375 (
		\m5_addr_i[3]_pad ,
		_w8989_,
		_w8990_,
		_w14276_
	);
	LUT3 #(
		.INIT('h57)
	) name12376 (
		_w8996_,
		_w14275_,
		_w14276_,
		_w14277_
	);
	LUT4 #(
		.INIT('h7fff)
	) name12377 (
		_w14268_,
		_w14271_,
		_w14274_,
		_w14277_,
		_w14278_
	);
	LUT3 #(
		.INIT('h80)
	) name12378 (
		\m2_addr_i[4]_pad ,
		_w8989_,
		_w8990_,
		_w14279_
	);
	LUT3 #(
		.INIT('h2a)
	) name12379 (
		\m3_addr_i[4]_pad ,
		_w8989_,
		_w8990_,
		_w14280_
	);
	LUT3 #(
		.INIT('h57)
	) name12380 (
		_w9002_,
		_w14279_,
		_w14280_,
		_w14281_
	);
	LUT3 #(
		.INIT('h80)
	) name12381 (
		\m0_addr_i[4]_pad ,
		_w8989_,
		_w8990_,
		_w14282_
	);
	LUT3 #(
		.INIT('h2a)
	) name12382 (
		\m7_addr_i[4]_pad ,
		_w8989_,
		_w8990_,
		_w14283_
	);
	LUT4 #(
		.INIT('h6e7f)
	) name12383 (
		_w8984_,
		_w8987_,
		_w14282_,
		_w14283_,
		_w14284_
	);
	LUT3 #(
		.INIT('h2a)
	) name12384 (
		\m1_addr_i[4]_pad ,
		_w8989_,
		_w8990_,
		_w14285_
	);
	LUT3 #(
		.INIT('h80)
	) name12385 (
		\m6_addr_i[4]_pad ,
		_w8989_,
		_w8990_,
		_w14286_
	);
	LUT4 #(
		.INIT('h6e7f)
	) name12386 (
		_w8984_,
		_w8987_,
		_w14285_,
		_w14286_,
		_w14287_
	);
	LUT3 #(
		.INIT('h80)
	) name12387 (
		\m4_addr_i[4]_pad ,
		_w8989_,
		_w8990_,
		_w14288_
	);
	LUT3 #(
		.INIT('h2a)
	) name12388 (
		\m5_addr_i[4]_pad ,
		_w8989_,
		_w8990_,
		_w14289_
	);
	LUT3 #(
		.INIT('h57)
	) name12389 (
		_w8996_,
		_w14288_,
		_w14289_,
		_w14290_
	);
	LUT4 #(
		.INIT('h7fff)
	) name12390 (
		_w14281_,
		_w14284_,
		_w14287_,
		_w14290_,
		_w14291_
	);
	LUT3 #(
		.INIT('h80)
	) name12391 (
		\m2_addr_i[5]_pad ,
		_w8989_,
		_w8990_,
		_w14292_
	);
	LUT3 #(
		.INIT('h2a)
	) name12392 (
		\m3_addr_i[5]_pad ,
		_w8989_,
		_w8990_,
		_w14293_
	);
	LUT3 #(
		.INIT('h57)
	) name12393 (
		_w9002_,
		_w14292_,
		_w14293_,
		_w14294_
	);
	LUT3 #(
		.INIT('h80)
	) name12394 (
		\m0_addr_i[5]_pad ,
		_w8989_,
		_w8990_,
		_w14295_
	);
	LUT3 #(
		.INIT('h2a)
	) name12395 (
		\m7_addr_i[5]_pad ,
		_w8989_,
		_w8990_,
		_w14296_
	);
	LUT4 #(
		.INIT('h6e7f)
	) name12396 (
		_w8984_,
		_w8987_,
		_w14295_,
		_w14296_,
		_w14297_
	);
	LUT3 #(
		.INIT('h2a)
	) name12397 (
		\m1_addr_i[5]_pad ,
		_w8989_,
		_w8990_,
		_w14298_
	);
	LUT3 #(
		.INIT('h80)
	) name12398 (
		\m6_addr_i[5]_pad ,
		_w8989_,
		_w8990_,
		_w14299_
	);
	LUT4 #(
		.INIT('h6e7f)
	) name12399 (
		_w8984_,
		_w8987_,
		_w14298_,
		_w14299_,
		_w14300_
	);
	LUT3 #(
		.INIT('h80)
	) name12400 (
		\m4_addr_i[5]_pad ,
		_w8989_,
		_w8990_,
		_w14301_
	);
	LUT3 #(
		.INIT('h2a)
	) name12401 (
		\m5_addr_i[5]_pad ,
		_w8989_,
		_w8990_,
		_w14302_
	);
	LUT3 #(
		.INIT('h57)
	) name12402 (
		_w8996_,
		_w14301_,
		_w14302_,
		_w14303_
	);
	LUT4 #(
		.INIT('h7fff)
	) name12403 (
		_w14294_,
		_w14297_,
		_w14300_,
		_w14303_,
		_w14304_
	);
	LUT3 #(
		.INIT('h80)
	) name12404 (
		\m2_addr_i[6]_pad ,
		_w8989_,
		_w8990_,
		_w14305_
	);
	LUT3 #(
		.INIT('h2a)
	) name12405 (
		\m3_addr_i[6]_pad ,
		_w8989_,
		_w8990_,
		_w14306_
	);
	LUT3 #(
		.INIT('h57)
	) name12406 (
		_w9002_,
		_w14305_,
		_w14306_,
		_w14307_
	);
	LUT3 #(
		.INIT('h80)
	) name12407 (
		\m0_addr_i[6]_pad ,
		_w8989_,
		_w8990_,
		_w14308_
	);
	LUT3 #(
		.INIT('h2a)
	) name12408 (
		\m7_addr_i[6]_pad ,
		_w8989_,
		_w8990_,
		_w14309_
	);
	LUT4 #(
		.INIT('h6e7f)
	) name12409 (
		_w8984_,
		_w8987_,
		_w14308_,
		_w14309_,
		_w14310_
	);
	LUT3 #(
		.INIT('h2a)
	) name12410 (
		\m1_addr_i[6]_pad ,
		_w8989_,
		_w8990_,
		_w14311_
	);
	LUT3 #(
		.INIT('h80)
	) name12411 (
		\m6_addr_i[6]_pad ,
		_w8989_,
		_w8990_,
		_w14312_
	);
	LUT4 #(
		.INIT('h6e7f)
	) name12412 (
		_w8984_,
		_w8987_,
		_w14311_,
		_w14312_,
		_w14313_
	);
	LUT3 #(
		.INIT('h80)
	) name12413 (
		\m4_addr_i[6]_pad ,
		_w8989_,
		_w8990_,
		_w14314_
	);
	LUT3 #(
		.INIT('h2a)
	) name12414 (
		\m5_addr_i[6]_pad ,
		_w8989_,
		_w8990_,
		_w14315_
	);
	LUT3 #(
		.INIT('h57)
	) name12415 (
		_w8996_,
		_w14314_,
		_w14315_,
		_w14316_
	);
	LUT4 #(
		.INIT('h7fff)
	) name12416 (
		_w14307_,
		_w14310_,
		_w14313_,
		_w14316_,
		_w14317_
	);
	LUT3 #(
		.INIT('h80)
	) name12417 (
		\m2_addr_i[7]_pad ,
		_w8989_,
		_w8990_,
		_w14318_
	);
	LUT3 #(
		.INIT('h2a)
	) name12418 (
		\m3_addr_i[7]_pad ,
		_w8989_,
		_w8990_,
		_w14319_
	);
	LUT3 #(
		.INIT('h57)
	) name12419 (
		_w9002_,
		_w14318_,
		_w14319_,
		_w14320_
	);
	LUT3 #(
		.INIT('h80)
	) name12420 (
		\m0_addr_i[7]_pad ,
		_w8989_,
		_w8990_,
		_w14321_
	);
	LUT3 #(
		.INIT('h2a)
	) name12421 (
		\m7_addr_i[7]_pad ,
		_w8989_,
		_w8990_,
		_w14322_
	);
	LUT4 #(
		.INIT('h6e7f)
	) name12422 (
		_w8984_,
		_w8987_,
		_w14321_,
		_w14322_,
		_w14323_
	);
	LUT3 #(
		.INIT('h2a)
	) name12423 (
		\m1_addr_i[7]_pad ,
		_w8989_,
		_w8990_,
		_w14324_
	);
	LUT3 #(
		.INIT('h80)
	) name12424 (
		\m6_addr_i[7]_pad ,
		_w8989_,
		_w8990_,
		_w14325_
	);
	LUT4 #(
		.INIT('h6e7f)
	) name12425 (
		_w8984_,
		_w8987_,
		_w14324_,
		_w14325_,
		_w14326_
	);
	LUT3 #(
		.INIT('h80)
	) name12426 (
		\m4_addr_i[7]_pad ,
		_w8989_,
		_w8990_,
		_w14327_
	);
	LUT3 #(
		.INIT('h2a)
	) name12427 (
		\m5_addr_i[7]_pad ,
		_w8989_,
		_w8990_,
		_w14328_
	);
	LUT3 #(
		.INIT('h57)
	) name12428 (
		_w8996_,
		_w14327_,
		_w14328_,
		_w14329_
	);
	LUT4 #(
		.INIT('h7fff)
	) name12429 (
		_w14320_,
		_w14323_,
		_w14326_,
		_w14329_,
		_w14330_
	);
	LUT3 #(
		.INIT('h80)
	) name12430 (
		\m0_addr_i[8]_pad ,
		_w8989_,
		_w8990_,
		_w14331_
	);
	LUT3 #(
		.INIT('h2a)
	) name12431 (
		\m1_addr_i[8]_pad ,
		_w8989_,
		_w8990_,
		_w14332_
	);
	LUT3 #(
		.INIT('h57)
	) name12432 (
		_w9008_,
		_w14331_,
		_w14332_,
		_w14333_
	);
	LUT3 #(
		.INIT('h80)
	) name12433 (
		\m6_addr_i[8]_pad ,
		_w8989_,
		_w8990_,
		_w14334_
	);
	LUT3 #(
		.INIT('h2a)
	) name12434 (
		\m3_addr_i[8]_pad ,
		_w8989_,
		_w8990_,
		_w14335_
	);
	LUT4 #(
		.INIT('habef)
	) name12435 (
		_w8984_,
		_w8987_,
		_w14334_,
		_w14335_,
		_w14336_
	);
	LUT3 #(
		.INIT('h2a)
	) name12436 (
		\m7_addr_i[8]_pad ,
		_w8989_,
		_w8990_,
		_w14337_
	);
	LUT3 #(
		.INIT('h80)
	) name12437 (
		\m2_addr_i[8]_pad ,
		_w8989_,
		_w8990_,
		_w14338_
	);
	LUT4 #(
		.INIT('habef)
	) name12438 (
		_w8984_,
		_w8987_,
		_w14337_,
		_w14338_,
		_w14339_
	);
	LUT3 #(
		.INIT('h80)
	) name12439 (
		\m4_addr_i[8]_pad ,
		_w8989_,
		_w8990_,
		_w14340_
	);
	LUT3 #(
		.INIT('h2a)
	) name12440 (
		\m5_addr_i[8]_pad ,
		_w8989_,
		_w8990_,
		_w14341_
	);
	LUT3 #(
		.INIT('h57)
	) name12441 (
		_w8996_,
		_w14340_,
		_w14341_,
		_w14342_
	);
	LUT4 #(
		.INIT('h7fff)
	) name12442 (
		_w14333_,
		_w14336_,
		_w14339_,
		_w14342_,
		_w14343_
	);
	LUT3 #(
		.INIT('h80)
	) name12443 (
		\m0_addr_i[9]_pad ,
		_w8989_,
		_w8990_,
		_w14344_
	);
	LUT3 #(
		.INIT('h2a)
	) name12444 (
		\m1_addr_i[9]_pad ,
		_w8989_,
		_w8990_,
		_w14345_
	);
	LUT3 #(
		.INIT('h57)
	) name12445 (
		_w9008_,
		_w14344_,
		_w14345_,
		_w14346_
	);
	LUT3 #(
		.INIT('h80)
	) name12446 (
		\m4_addr_i[9]_pad ,
		_w8989_,
		_w8990_,
		_w14347_
	);
	LUT3 #(
		.INIT('h2a)
	) name12447 (
		\m3_addr_i[9]_pad ,
		_w8989_,
		_w8990_,
		_w14348_
	);
	LUT4 #(
		.INIT('h9bdf)
	) name12448 (
		_w8984_,
		_w8987_,
		_w14347_,
		_w14348_,
		_w14349_
	);
	LUT3 #(
		.INIT('h2a)
	) name12449 (
		\m5_addr_i[9]_pad ,
		_w8989_,
		_w8990_,
		_w14350_
	);
	LUT3 #(
		.INIT('h80)
	) name12450 (
		\m2_addr_i[9]_pad ,
		_w8989_,
		_w8990_,
		_w14351_
	);
	LUT4 #(
		.INIT('h9bdf)
	) name12451 (
		_w8984_,
		_w8987_,
		_w14350_,
		_w14351_,
		_w14352_
	);
	LUT3 #(
		.INIT('h80)
	) name12452 (
		\m6_addr_i[9]_pad ,
		_w8989_,
		_w8990_,
		_w14353_
	);
	LUT3 #(
		.INIT('h2a)
	) name12453 (
		\m7_addr_i[9]_pad ,
		_w8989_,
		_w8990_,
		_w14354_
	);
	LUT3 #(
		.INIT('h57)
	) name12454 (
		_w8988_,
		_w14353_,
		_w14354_,
		_w14355_
	);
	LUT4 #(
		.INIT('h7fff)
	) name12455 (
		_w14346_,
		_w14349_,
		_w14352_,
		_w14355_,
		_w14356_
	);
	LUT3 #(
		.INIT('h80)
	) name12456 (
		\m0_data_i[0]_pad ,
		_w8989_,
		_w8990_,
		_w14357_
	);
	LUT3 #(
		.INIT('h2a)
	) name12457 (
		\m1_data_i[0]_pad ,
		_w8989_,
		_w8990_,
		_w14358_
	);
	LUT3 #(
		.INIT('h57)
	) name12458 (
		_w9008_,
		_w14357_,
		_w14358_,
		_w14359_
	);
	LUT3 #(
		.INIT('h80)
	) name12459 (
		\m4_data_i[0]_pad ,
		_w8989_,
		_w8990_,
		_w14360_
	);
	LUT3 #(
		.INIT('h2a)
	) name12460 (
		\m3_data_i[0]_pad ,
		_w8989_,
		_w8990_,
		_w14361_
	);
	LUT4 #(
		.INIT('h9bdf)
	) name12461 (
		_w8984_,
		_w8987_,
		_w14360_,
		_w14361_,
		_w14362_
	);
	LUT3 #(
		.INIT('h2a)
	) name12462 (
		\m5_data_i[0]_pad ,
		_w8989_,
		_w8990_,
		_w14363_
	);
	LUT3 #(
		.INIT('h80)
	) name12463 (
		\m2_data_i[0]_pad ,
		_w8989_,
		_w8990_,
		_w14364_
	);
	LUT4 #(
		.INIT('h9bdf)
	) name12464 (
		_w8984_,
		_w8987_,
		_w14363_,
		_w14364_,
		_w14365_
	);
	LUT3 #(
		.INIT('h80)
	) name12465 (
		\m6_data_i[0]_pad ,
		_w8989_,
		_w8990_,
		_w14366_
	);
	LUT3 #(
		.INIT('h2a)
	) name12466 (
		\m7_data_i[0]_pad ,
		_w8989_,
		_w8990_,
		_w14367_
	);
	LUT3 #(
		.INIT('h57)
	) name12467 (
		_w8988_,
		_w14366_,
		_w14367_,
		_w14368_
	);
	LUT4 #(
		.INIT('h7fff)
	) name12468 (
		_w14359_,
		_w14362_,
		_w14365_,
		_w14368_,
		_w14369_
	);
	LUT3 #(
		.INIT('h80)
	) name12469 (
		\m0_data_i[10]_pad ,
		_w8989_,
		_w8990_,
		_w14370_
	);
	LUT3 #(
		.INIT('h2a)
	) name12470 (
		\m1_data_i[10]_pad ,
		_w8989_,
		_w8990_,
		_w14371_
	);
	LUT3 #(
		.INIT('h57)
	) name12471 (
		_w9008_,
		_w14370_,
		_w14371_,
		_w14372_
	);
	LUT3 #(
		.INIT('h80)
	) name12472 (
		\m6_data_i[10]_pad ,
		_w8989_,
		_w8990_,
		_w14373_
	);
	LUT3 #(
		.INIT('h2a)
	) name12473 (
		\m3_data_i[10]_pad ,
		_w8989_,
		_w8990_,
		_w14374_
	);
	LUT4 #(
		.INIT('habef)
	) name12474 (
		_w8984_,
		_w8987_,
		_w14373_,
		_w14374_,
		_w14375_
	);
	LUT3 #(
		.INIT('h2a)
	) name12475 (
		\m7_data_i[10]_pad ,
		_w8989_,
		_w8990_,
		_w14376_
	);
	LUT3 #(
		.INIT('h80)
	) name12476 (
		\m2_data_i[10]_pad ,
		_w8989_,
		_w8990_,
		_w14377_
	);
	LUT4 #(
		.INIT('habef)
	) name12477 (
		_w8984_,
		_w8987_,
		_w14376_,
		_w14377_,
		_w14378_
	);
	LUT3 #(
		.INIT('h80)
	) name12478 (
		\m4_data_i[10]_pad ,
		_w8989_,
		_w8990_,
		_w14379_
	);
	LUT3 #(
		.INIT('h2a)
	) name12479 (
		\m5_data_i[10]_pad ,
		_w8989_,
		_w8990_,
		_w14380_
	);
	LUT3 #(
		.INIT('h57)
	) name12480 (
		_w8996_,
		_w14379_,
		_w14380_,
		_w14381_
	);
	LUT4 #(
		.INIT('h7fff)
	) name12481 (
		_w14372_,
		_w14375_,
		_w14378_,
		_w14381_,
		_w14382_
	);
	LUT3 #(
		.INIT('h80)
	) name12482 (
		\m2_data_i[11]_pad ,
		_w8989_,
		_w8990_,
		_w14383_
	);
	LUT3 #(
		.INIT('h2a)
	) name12483 (
		\m3_data_i[11]_pad ,
		_w8989_,
		_w8990_,
		_w14384_
	);
	LUT3 #(
		.INIT('h57)
	) name12484 (
		_w9002_,
		_w14383_,
		_w14384_,
		_w14385_
	);
	LUT3 #(
		.INIT('h80)
	) name12485 (
		\m6_data_i[11]_pad ,
		_w8989_,
		_w8990_,
		_w14386_
	);
	LUT3 #(
		.INIT('h2a)
	) name12486 (
		\m1_data_i[11]_pad ,
		_w8989_,
		_w8990_,
		_w14387_
	);
	LUT4 #(
		.INIT('h67ef)
	) name12487 (
		_w8984_,
		_w8987_,
		_w14386_,
		_w14387_,
		_w14388_
	);
	LUT3 #(
		.INIT('h2a)
	) name12488 (
		\m7_data_i[11]_pad ,
		_w8989_,
		_w8990_,
		_w14389_
	);
	LUT3 #(
		.INIT('h80)
	) name12489 (
		\m0_data_i[11]_pad ,
		_w8989_,
		_w8990_,
		_w14390_
	);
	LUT4 #(
		.INIT('h67ef)
	) name12490 (
		_w8984_,
		_w8987_,
		_w14389_,
		_w14390_,
		_w14391_
	);
	LUT3 #(
		.INIT('h80)
	) name12491 (
		\m4_data_i[11]_pad ,
		_w8989_,
		_w8990_,
		_w14392_
	);
	LUT3 #(
		.INIT('h2a)
	) name12492 (
		\m5_data_i[11]_pad ,
		_w8989_,
		_w8990_,
		_w14393_
	);
	LUT3 #(
		.INIT('h57)
	) name12493 (
		_w8996_,
		_w14392_,
		_w14393_,
		_w14394_
	);
	LUT4 #(
		.INIT('h7fff)
	) name12494 (
		_w14385_,
		_w14388_,
		_w14391_,
		_w14394_,
		_w14395_
	);
	LUT3 #(
		.INIT('h80)
	) name12495 (
		\m0_data_i[12]_pad ,
		_w8989_,
		_w8990_,
		_w14396_
	);
	LUT3 #(
		.INIT('h2a)
	) name12496 (
		\m1_data_i[12]_pad ,
		_w8989_,
		_w8990_,
		_w14397_
	);
	LUT3 #(
		.INIT('h57)
	) name12497 (
		_w9008_,
		_w14396_,
		_w14397_,
		_w14398_
	);
	LUT3 #(
		.INIT('h80)
	) name12498 (
		\m4_data_i[12]_pad ,
		_w8989_,
		_w8990_,
		_w14399_
	);
	LUT3 #(
		.INIT('h2a)
	) name12499 (
		\m3_data_i[12]_pad ,
		_w8989_,
		_w8990_,
		_w14400_
	);
	LUT4 #(
		.INIT('h9bdf)
	) name12500 (
		_w8984_,
		_w8987_,
		_w14399_,
		_w14400_,
		_w14401_
	);
	LUT3 #(
		.INIT('h2a)
	) name12501 (
		\m5_data_i[12]_pad ,
		_w8989_,
		_w8990_,
		_w14402_
	);
	LUT3 #(
		.INIT('h80)
	) name12502 (
		\m2_data_i[12]_pad ,
		_w8989_,
		_w8990_,
		_w14403_
	);
	LUT4 #(
		.INIT('h9bdf)
	) name12503 (
		_w8984_,
		_w8987_,
		_w14402_,
		_w14403_,
		_w14404_
	);
	LUT3 #(
		.INIT('h80)
	) name12504 (
		\m6_data_i[12]_pad ,
		_w8989_,
		_w8990_,
		_w14405_
	);
	LUT3 #(
		.INIT('h2a)
	) name12505 (
		\m7_data_i[12]_pad ,
		_w8989_,
		_w8990_,
		_w14406_
	);
	LUT3 #(
		.INIT('h57)
	) name12506 (
		_w8988_,
		_w14405_,
		_w14406_,
		_w14407_
	);
	LUT4 #(
		.INIT('h7fff)
	) name12507 (
		_w14398_,
		_w14401_,
		_w14404_,
		_w14407_,
		_w14408_
	);
	LUT3 #(
		.INIT('h80)
	) name12508 (
		\m0_data_i[13]_pad ,
		_w8989_,
		_w8990_,
		_w14409_
	);
	LUT3 #(
		.INIT('h2a)
	) name12509 (
		\m1_data_i[13]_pad ,
		_w8989_,
		_w8990_,
		_w14410_
	);
	LUT3 #(
		.INIT('h57)
	) name12510 (
		_w9008_,
		_w14409_,
		_w14410_,
		_w14411_
	);
	LUT3 #(
		.INIT('h80)
	) name12511 (
		\m2_data_i[13]_pad ,
		_w8989_,
		_w8990_,
		_w14412_
	);
	LUT3 #(
		.INIT('h2a)
	) name12512 (
		\m7_data_i[13]_pad ,
		_w8989_,
		_w8990_,
		_w14413_
	);
	LUT4 #(
		.INIT('haebf)
	) name12513 (
		_w8984_,
		_w8987_,
		_w14412_,
		_w14413_,
		_w14414_
	);
	LUT3 #(
		.INIT('h2a)
	) name12514 (
		\m3_data_i[13]_pad ,
		_w8989_,
		_w8990_,
		_w14415_
	);
	LUT3 #(
		.INIT('h80)
	) name12515 (
		\m6_data_i[13]_pad ,
		_w8989_,
		_w8990_,
		_w14416_
	);
	LUT4 #(
		.INIT('haebf)
	) name12516 (
		_w8984_,
		_w8987_,
		_w14415_,
		_w14416_,
		_w14417_
	);
	LUT3 #(
		.INIT('h80)
	) name12517 (
		\m4_data_i[13]_pad ,
		_w8989_,
		_w8990_,
		_w14418_
	);
	LUT3 #(
		.INIT('h2a)
	) name12518 (
		\m5_data_i[13]_pad ,
		_w8989_,
		_w8990_,
		_w14419_
	);
	LUT3 #(
		.INIT('h57)
	) name12519 (
		_w8996_,
		_w14418_,
		_w14419_,
		_w14420_
	);
	LUT4 #(
		.INIT('h7fff)
	) name12520 (
		_w14411_,
		_w14414_,
		_w14417_,
		_w14420_,
		_w14421_
	);
	LUT3 #(
		.INIT('h80)
	) name12521 (
		\m2_data_i[14]_pad ,
		_w8989_,
		_w8990_,
		_w14422_
	);
	LUT3 #(
		.INIT('h2a)
	) name12522 (
		\m3_data_i[14]_pad ,
		_w8989_,
		_w8990_,
		_w14423_
	);
	LUT3 #(
		.INIT('h57)
	) name12523 (
		_w9002_,
		_w14422_,
		_w14423_,
		_w14424_
	);
	LUT3 #(
		.INIT('h80)
	) name12524 (
		\m6_data_i[14]_pad ,
		_w8989_,
		_w8990_,
		_w14425_
	);
	LUT3 #(
		.INIT('h2a)
	) name12525 (
		\m1_data_i[14]_pad ,
		_w8989_,
		_w8990_,
		_w14426_
	);
	LUT4 #(
		.INIT('h67ef)
	) name12526 (
		_w8984_,
		_w8987_,
		_w14425_,
		_w14426_,
		_w14427_
	);
	LUT3 #(
		.INIT('h2a)
	) name12527 (
		\m7_data_i[14]_pad ,
		_w8989_,
		_w8990_,
		_w14428_
	);
	LUT3 #(
		.INIT('h80)
	) name12528 (
		\m0_data_i[14]_pad ,
		_w8989_,
		_w8990_,
		_w14429_
	);
	LUT4 #(
		.INIT('h67ef)
	) name12529 (
		_w8984_,
		_w8987_,
		_w14428_,
		_w14429_,
		_w14430_
	);
	LUT3 #(
		.INIT('h80)
	) name12530 (
		\m4_data_i[14]_pad ,
		_w8989_,
		_w8990_,
		_w14431_
	);
	LUT3 #(
		.INIT('h2a)
	) name12531 (
		\m5_data_i[14]_pad ,
		_w8989_,
		_w8990_,
		_w14432_
	);
	LUT3 #(
		.INIT('h57)
	) name12532 (
		_w8996_,
		_w14431_,
		_w14432_,
		_w14433_
	);
	LUT4 #(
		.INIT('h7fff)
	) name12533 (
		_w14424_,
		_w14427_,
		_w14430_,
		_w14433_,
		_w14434_
	);
	LUT3 #(
		.INIT('h80)
	) name12534 (
		\m2_data_i[15]_pad ,
		_w8989_,
		_w8990_,
		_w14435_
	);
	LUT3 #(
		.INIT('h2a)
	) name12535 (
		\m3_data_i[15]_pad ,
		_w8989_,
		_w8990_,
		_w14436_
	);
	LUT3 #(
		.INIT('h57)
	) name12536 (
		_w9002_,
		_w14435_,
		_w14436_,
		_w14437_
	);
	LUT3 #(
		.INIT('h80)
	) name12537 (
		\m0_data_i[15]_pad ,
		_w8989_,
		_w8990_,
		_w14438_
	);
	LUT3 #(
		.INIT('h2a)
	) name12538 (
		\m7_data_i[15]_pad ,
		_w8989_,
		_w8990_,
		_w14439_
	);
	LUT4 #(
		.INIT('h6e7f)
	) name12539 (
		_w8984_,
		_w8987_,
		_w14438_,
		_w14439_,
		_w14440_
	);
	LUT3 #(
		.INIT('h2a)
	) name12540 (
		\m1_data_i[15]_pad ,
		_w8989_,
		_w8990_,
		_w14441_
	);
	LUT3 #(
		.INIT('h80)
	) name12541 (
		\m6_data_i[15]_pad ,
		_w8989_,
		_w8990_,
		_w14442_
	);
	LUT4 #(
		.INIT('h6e7f)
	) name12542 (
		_w8984_,
		_w8987_,
		_w14441_,
		_w14442_,
		_w14443_
	);
	LUT3 #(
		.INIT('h80)
	) name12543 (
		\m4_data_i[15]_pad ,
		_w8989_,
		_w8990_,
		_w14444_
	);
	LUT3 #(
		.INIT('h2a)
	) name12544 (
		\m5_data_i[15]_pad ,
		_w8989_,
		_w8990_,
		_w14445_
	);
	LUT3 #(
		.INIT('h57)
	) name12545 (
		_w8996_,
		_w14444_,
		_w14445_,
		_w14446_
	);
	LUT4 #(
		.INIT('h7fff)
	) name12546 (
		_w14437_,
		_w14440_,
		_w14443_,
		_w14446_,
		_w14447_
	);
	LUT3 #(
		.INIT('h80)
	) name12547 (
		\m0_data_i[16]_pad ,
		_w8989_,
		_w8990_,
		_w14448_
	);
	LUT3 #(
		.INIT('h2a)
	) name12548 (
		\m1_data_i[16]_pad ,
		_w8989_,
		_w8990_,
		_w14449_
	);
	LUT3 #(
		.INIT('h57)
	) name12549 (
		_w9008_,
		_w14448_,
		_w14449_,
		_w14450_
	);
	LUT3 #(
		.INIT('h80)
	) name12550 (
		\m4_data_i[16]_pad ,
		_w8989_,
		_w8990_,
		_w14451_
	);
	LUT3 #(
		.INIT('h2a)
	) name12551 (
		\m3_data_i[16]_pad ,
		_w8989_,
		_w8990_,
		_w14452_
	);
	LUT4 #(
		.INIT('h9bdf)
	) name12552 (
		_w8984_,
		_w8987_,
		_w14451_,
		_w14452_,
		_w14453_
	);
	LUT3 #(
		.INIT('h2a)
	) name12553 (
		\m5_data_i[16]_pad ,
		_w8989_,
		_w8990_,
		_w14454_
	);
	LUT3 #(
		.INIT('h80)
	) name12554 (
		\m2_data_i[16]_pad ,
		_w8989_,
		_w8990_,
		_w14455_
	);
	LUT4 #(
		.INIT('h9bdf)
	) name12555 (
		_w8984_,
		_w8987_,
		_w14454_,
		_w14455_,
		_w14456_
	);
	LUT3 #(
		.INIT('h80)
	) name12556 (
		\m6_data_i[16]_pad ,
		_w8989_,
		_w8990_,
		_w14457_
	);
	LUT3 #(
		.INIT('h2a)
	) name12557 (
		\m7_data_i[16]_pad ,
		_w8989_,
		_w8990_,
		_w14458_
	);
	LUT3 #(
		.INIT('h57)
	) name12558 (
		_w8988_,
		_w14457_,
		_w14458_,
		_w14459_
	);
	LUT4 #(
		.INIT('h7fff)
	) name12559 (
		_w14450_,
		_w14453_,
		_w14456_,
		_w14459_,
		_w14460_
	);
	LUT3 #(
		.INIT('h80)
	) name12560 (
		\m2_data_i[17]_pad ,
		_w8989_,
		_w8990_,
		_w14461_
	);
	LUT3 #(
		.INIT('h2a)
	) name12561 (
		\m3_data_i[17]_pad ,
		_w8989_,
		_w8990_,
		_w14462_
	);
	LUT3 #(
		.INIT('h57)
	) name12562 (
		_w9002_,
		_w14461_,
		_w14462_,
		_w14463_
	);
	LUT3 #(
		.INIT('h80)
	) name12563 (
		\m0_data_i[17]_pad ,
		_w8989_,
		_w8990_,
		_w14464_
	);
	LUT3 #(
		.INIT('h2a)
	) name12564 (
		\m7_data_i[17]_pad ,
		_w8989_,
		_w8990_,
		_w14465_
	);
	LUT4 #(
		.INIT('h6e7f)
	) name12565 (
		_w8984_,
		_w8987_,
		_w14464_,
		_w14465_,
		_w14466_
	);
	LUT3 #(
		.INIT('h2a)
	) name12566 (
		\m1_data_i[17]_pad ,
		_w8989_,
		_w8990_,
		_w14467_
	);
	LUT3 #(
		.INIT('h80)
	) name12567 (
		\m6_data_i[17]_pad ,
		_w8989_,
		_w8990_,
		_w14468_
	);
	LUT4 #(
		.INIT('h6e7f)
	) name12568 (
		_w8984_,
		_w8987_,
		_w14467_,
		_w14468_,
		_w14469_
	);
	LUT3 #(
		.INIT('h80)
	) name12569 (
		\m4_data_i[17]_pad ,
		_w8989_,
		_w8990_,
		_w14470_
	);
	LUT3 #(
		.INIT('h2a)
	) name12570 (
		\m5_data_i[17]_pad ,
		_w8989_,
		_w8990_,
		_w14471_
	);
	LUT3 #(
		.INIT('h57)
	) name12571 (
		_w8996_,
		_w14470_,
		_w14471_,
		_w14472_
	);
	LUT4 #(
		.INIT('h7fff)
	) name12572 (
		_w14463_,
		_w14466_,
		_w14469_,
		_w14472_,
		_w14473_
	);
	LUT3 #(
		.INIT('h80)
	) name12573 (
		\m4_data_i[18]_pad ,
		_w8989_,
		_w8990_,
		_w14474_
	);
	LUT3 #(
		.INIT('h2a)
	) name12574 (
		\m5_data_i[18]_pad ,
		_w8989_,
		_w8990_,
		_w14475_
	);
	LUT3 #(
		.INIT('h57)
	) name12575 (
		_w8996_,
		_w14474_,
		_w14475_,
		_w14476_
	);
	LUT3 #(
		.INIT('h80)
	) name12576 (
		\m0_data_i[18]_pad ,
		_w8989_,
		_w8990_,
		_w14477_
	);
	LUT3 #(
		.INIT('h2a)
	) name12577 (
		\m7_data_i[18]_pad ,
		_w8989_,
		_w8990_,
		_w14478_
	);
	LUT4 #(
		.INIT('h6e7f)
	) name12578 (
		_w8984_,
		_w8987_,
		_w14477_,
		_w14478_,
		_w14479_
	);
	LUT3 #(
		.INIT('h2a)
	) name12579 (
		\m1_data_i[18]_pad ,
		_w8989_,
		_w8990_,
		_w14480_
	);
	LUT3 #(
		.INIT('h80)
	) name12580 (
		\m6_data_i[18]_pad ,
		_w8989_,
		_w8990_,
		_w14481_
	);
	LUT4 #(
		.INIT('h6e7f)
	) name12581 (
		_w8984_,
		_w8987_,
		_w14480_,
		_w14481_,
		_w14482_
	);
	LUT3 #(
		.INIT('h80)
	) name12582 (
		\m2_data_i[18]_pad ,
		_w8989_,
		_w8990_,
		_w14483_
	);
	LUT3 #(
		.INIT('h2a)
	) name12583 (
		\m3_data_i[18]_pad ,
		_w8989_,
		_w8990_,
		_w14484_
	);
	LUT3 #(
		.INIT('h57)
	) name12584 (
		_w9002_,
		_w14483_,
		_w14484_,
		_w14485_
	);
	LUT4 #(
		.INIT('h7fff)
	) name12585 (
		_w14476_,
		_w14479_,
		_w14482_,
		_w14485_,
		_w14486_
	);
	LUT3 #(
		.INIT('h80)
	) name12586 (
		\m2_data_i[19]_pad ,
		_w8989_,
		_w8990_,
		_w14487_
	);
	LUT3 #(
		.INIT('h2a)
	) name12587 (
		\m3_data_i[19]_pad ,
		_w8989_,
		_w8990_,
		_w14488_
	);
	LUT3 #(
		.INIT('h57)
	) name12588 (
		_w9002_,
		_w14487_,
		_w14488_,
		_w14489_
	);
	LUT3 #(
		.INIT('h80)
	) name12589 (
		\m0_data_i[19]_pad ,
		_w8989_,
		_w8990_,
		_w14490_
	);
	LUT3 #(
		.INIT('h2a)
	) name12590 (
		\m7_data_i[19]_pad ,
		_w8989_,
		_w8990_,
		_w14491_
	);
	LUT4 #(
		.INIT('h6e7f)
	) name12591 (
		_w8984_,
		_w8987_,
		_w14490_,
		_w14491_,
		_w14492_
	);
	LUT3 #(
		.INIT('h2a)
	) name12592 (
		\m1_data_i[19]_pad ,
		_w8989_,
		_w8990_,
		_w14493_
	);
	LUT3 #(
		.INIT('h80)
	) name12593 (
		\m6_data_i[19]_pad ,
		_w8989_,
		_w8990_,
		_w14494_
	);
	LUT4 #(
		.INIT('h6e7f)
	) name12594 (
		_w8984_,
		_w8987_,
		_w14493_,
		_w14494_,
		_w14495_
	);
	LUT3 #(
		.INIT('h80)
	) name12595 (
		\m4_data_i[19]_pad ,
		_w8989_,
		_w8990_,
		_w14496_
	);
	LUT3 #(
		.INIT('h2a)
	) name12596 (
		\m5_data_i[19]_pad ,
		_w8989_,
		_w8990_,
		_w14497_
	);
	LUT3 #(
		.INIT('h57)
	) name12597 (
		_w8996_,
		_w14496_,
		_w14497_,
		_w14498_
	);
	LUT4 #(
		.INIT('h7fff)
	) name12598 (
		_w14489_,
		_w14492_,
		_w14495_,
		_w14498_,
		_w14499_
	);
	LUT3 #(
		.INIT('h80)
	) name12599 (
		\m4_data_i[1]_pad ,
		_w8989_,
		_w8990_,
		_w14500_
	);
	LUT3 #(
		.INIT('h2a)
	) name12600 (
		\m5_data_i[1]_pad ,
		_w8989_,
		_w8990_,
		_w14501_
	);
	LUT3 #(
		.INIT('h57)
	) name12601 (
		_w8996_,
		_w14500_,
		_w14501_,
		_w14502_
	);
	LUT3 #(
		.INIT('h80)
	) name12602 (
		\m6_data_i[1]_pad ,
		_w8989_,
		_w8990_,
		_w14503_
	);
	LUT3 #(
		.INIT('h2a)
	) name12603 (
		\m1_data_i[1]_pad ,
		_w8989_,
		_w8990_,
		_w14504_
	);
	LUT4 #(
		.INIT('h67ef)
	) name12604 (
		_w8984_,
		_w8987_,
		_w14503_,
		_w14504_,
		_w14505_
	);
	LUT3 #(
		.INIT('h2a)
	) name12605 (
		\m7_data_i[1]_pad ,
		_w8989_,
		_w8990_,
		_w14506_
	);
	LUT3 #(
		.INIT('h80)
	) name12606 (
		\m0_data_i[1]_pad ,
		_w8989_,
		_w8990_,
		_w14507_
	);
	LUT4 #(
		.INIT('h67ef)
	) name12607 (
		_w8984_,
		_w8987_,
		_w14506_,
		_w14507_,
		_w14508_
	);
	LUT3 #(
		.INIT('h80)
	) name12608 (
		\m2_data_i[1]_pad ,
		_w8989_,
		_w8990_,
		_w14509_
	);
	LUT3 #(
		.INIT('h2a)
	) name12609 (
		\m3_data_i[1]_pad ,
		_w8989_,
		_w8990_,
		_w14510_
	);
	LUT3 #(
		.INIT('h57)
	) name12610 (
		_w9002_,
		_w14509_,
		_w14510_,
		_w14511_
	);
	LUT4 #(
		.INIT('h7fff)
	) name12611 (
		_w14502_,
		_w14505_,
		_w14508_,
		_w14511_,
		_w14512_
	);
	LUT3 #(
		.INIT('h80)
	) name12612 (
		\m6_data_i[20]_pad ,
		_w8989_,
		_w8990_,
		_w14513_
	);
	LUT3 #(
		.INIT('h2a)
	) name12613 (
		\m7_data_i[20]_pad ,
		_w8989_,
		_w8990_,
		_w14514_
	);
	LUT3 #(
		.INIT('h57)
	) name12614 (
		_w8988_,
		_w14513_,
		_w14514_,
		_w14515_
	);
	LUT3 #(
		.INIT('h80)
	) name12615 (
		\m2_data_i[20]_pad ,
		_w8989_,
		_w8990_,
		_w14516_
	);
	LUT3 #(
		.INIT('h2a)
	) name12616 (
		\m5_data_i[20]_pad ,
		_w8989_,
		_w8990_,
		_w14517_
	);
	LUT4 #(
		.INIT('h9dbf)
	) name12617 (
		_w8984_,
		_w8987_,
		_w14516_,
		_w14517_,
		_w14518_
	);
	LUT3 #(
		.INIT('h2a)
	) name12618 (
		\m3_data_i[20]_pad ,
		_w8989_,
		_w8990_,
		_w14519_
	);
	LUT3 #(
		.INIT('h80)
	) name12619 (
		\m4_data_i[20]_pad ,
		_w8989_,
		_w8990_,
		_w14520_
	);
	LUT4 #(
		.INIT('h9dbf)
	) name12620 (
		_w8984_,
		_w8987_,
		_w14519_,
		_w14520_,
		_w14521_
	);
	LUT3 #(
		.INIT('h80)
	) name12621 (
		\m0_data_i[20]_pad ,
		_w8989_,
		_w8990_,
		_w14522_
	);
	LUT3 #(
		.INIT('h2a)
	) name12622 (
		\m1_data_i[20]_pad ,
		_w8989_,
		_w8990_,
		_w14523_
	);
	LUT3 #(
		.INIT('h57)
	) name12623 (
		_w9008_,
		_w14522_,
		_w14523_,
		_w14524_
	);
	LUT4 #(
		.INIT('h7fff)
	) name12624 (
		_w14515_,
		_w14518_,
		_w14521_,
		_w14524_,
		_w14525_
	);
	LUT3 #(
		.INIT('h80)
	) name12625 (
		\m6_data_i[21]_pad ,
		_w8989_,
		_w8990_,
		_w14526_
	);
	LUT3 #(
		.INIT('h2a)
	) name12626 (
		\m7_data_i[21]_pad ,
		_w8989_,
		_w8990_,
		_w14527_
	);
	LUT3 #(
		.INIT('h57)
	) name12627 (
		_w8988_,
		_w14526_,
		_w14527_,
		_w14528_
	);
	LUT3 #(
		.INIT('h80)
	) name12628 (
		\m2_data_i[21]_pad ,
		_w8989_,
		_w8990_,
		_w14529_
	);
	LUT3 #(
		.INIT('h2a)
	) name12629 (
		\m5_data_i[21]_pad ,
		_w8989_,
		_w8990_,
		_w14530_
	);
	LUT4 #(
		.INIT('h9dbf)
	) name12630 (
		_w8984_,
		_w8987_,
		_w14529_,
		_w14530_,
		_w14531_
	);
	LUT3 #(
		.INIT('h2a)
	) name12631 (
		\m3_data_i[21]_pad ,
		_w8989_,
		_w8990_,
		_w14532_
	);
	LUT3 #(
		.INIT('h80)
	) name12632 (
		\m4_data_i[21]_pad ,
		_w8989_,
		_w8990_,
		_w14533_
	);
	LUT4 #(
		.INIT('h9dbf)
	) name12633 (
		_w8984_,
		_w8987_,
		_w14532_,
		_w14533_,
		_w14534_
	);
	LUT3 #(
		.INIT('h80)
	) name12634 (
		\m0_data_i[21]_pad ,
		_w8989_,
		_w8990_,
		_w14535_
	);
	LUT3 #(
		.INIT('h2a)
	) name12635 (
		\m1_data_i[21]_pad ,
		_w8989_,
		_w8990_,
		_w14536_
	);
	LUT3 #(
		.INIT('h57)
	) name12636 (
		_w9008_,
		_w14535_,
		_w14536_,
		_w14537_
	);
	LUT4 #(
		.INIT('h7fff)
	) name12637 (
		_w14528_,
		_w14531_,
		_w14534_,
		_w14537_,
		_w14538_
	);
	LUT3 #(
		.INIT('h80)
	) name12638 (
		\m6_data_i[22]_pad ,
		_w8989_,
		_w8990_,
		_w14539_
	);
	LUT3 #(
		.INIT('h2a)
	) name12639 (
		\m7_data_i[22]_pad ,
		_w8989_,
		_w8990_,
		_w14540_
	);
	LUT3 #(
		.INIT('h57)
	) name12640 (
		_w8988_,
		_w14539_,
		_w14540_,
		_w14541_
	);
	LUT3 #(
		.INIT('h80)
	) name12641 (
		\m4_data_i[22]_pad ,
		_w8989_,
		_w8990_,
		_w14542_
	);
	LUT3 #(
		.INIT('h2a)
	) name12642 (
		\m3_data_i[22]_pad ,
		_w8989_,
		_w8990_,
		_w14543_
	);
	LUT4 #(
		.INIT('h9bdf)
	) name12643 (
		_w8984_,
		_w8987_,
		_w14542_,
		_w14543_,
		_w14544_
	);
	LUT3 #(
		.INIT('h2a)
	) name12644 (
		\m5_data_i[22]_pad ,
		_w8989_,
		_w8990_,
		_w14545_
	);
	LUT3 #(
		.INIT('h80)
	) name12645 (
		\m2_data_i[22]_pad ,
		_w8989_,
		_w8990_,
		_w14546_
	);
	LUT4 #(
		.INIT('h9bdf)
	) name12646 (
		_w8984_,
		_w8987_,
		_w14545_,
		_w14546_,
		_w14547_
	);
	LUT3 #(
		.INIT('h80)
	) name12647 (
		\m0_data_i[22]_pad ,
		_w8989_,
		_w8990_,
		_w14548_
	);
	LUT3 #(
		.INIT('h2a)
	) name12648 (
		\m1_data_i[22]_pad ,
		_w8989_,
		_w8990_,
		_w14549_
	);
	LUT3 #(
		.INIT('h57)
	) name12649 (
		_w9008_,
		_w14548_,
		_w14549_,
		_w14550_
	);
	LUT4 #(
		.INIT('h7fff)
	) name12650 (
		_w14541_,
		_w14544_,
		_w14547_,
		_w14550_,
		_w14551_
	);
	LUT3 #(
		.INIT('h80)
	) name12651 (
		\m6_data_i[23]_pad ,
		_w8989_,
		_w8990_,
		_w14552_
	);
	LUT3 #(
		.INIT('h2a)
	) name12652 (
		\m7_data_i[23]_pad ,
		_w8989_,
		_w8990_,
		_w14553_
	);
	LUT3 #(
		.INIT('h57)
	) name12653 (
		_w8988_,
		_w14552_,
		_w14553_,
		_w14554_
	);
	LUT3 #(
		.INIT('h80)
	) name12654 (
		\m4_data_i[23]_pad ,
		_w8989_,
		_w8990_,
		_w14555_
	);
	LUT3 #(
		.INIT('h2a)
	) name12655 (
		\m3_data_i[23]_pad ,
		_w8989_,
		_w8990_,
		_w14556_
	);
	LUT4 #(
		.INIT('h9bdf)
	) name12656 (
		_w8984_,
		_w8987_,
		_w14555_,
		_w14556_,
		_w14557_
	);
	LUT3 #(
		.INIT('h2a)
	) name12657 (
		\m5_data_i[23]_pad ,
		_w8989_,
		_w8990_,
		_w14558_
	);
	LUT3 #(
		.INIT('h80)
	) name12658 (
		\m2_data_i[23]_pad ,
		_w8989_,
		_w8990_,
		_w14559_
	);
	LUT4 #(
		.INIT('h9bdf)
	) name12659 (
		_w8984_,
		_w8987_,
		_w14558_,
		_w14559_,
		_w14560_
	);
	LUT3 #(
		.INIT('h80)
	) name12660 (
		\m0_data_i[23]_pad ,
		_w8989_,
		_w8990_,
		_w14561_
	);
	LUT3 #(
		.INIT('h2a)
	) name12661 (
		\m1_data_i[23]_pad ,
		_w8989_,
		_w8990_,
		_w14562_
	);
	LUT3 #(
		.INIT('h57)
	) name12662 (
		_w9008_,
		_w14561_,
		_w14562_,
		_w14563_
	);
	LUT4 #(
		.INIT('h7fff)
	) name12663 (
		_w14554_,
		_w14557_,
		_w14560_,
		_w14563_,
		_w14564_
	);
	LUT3 #(
		.INIT('h80)
	) name12664 (
		\m0_data_i[24]_pad ,
		_w8989_,
		_w8990_,
		_w14565_
	);
	LUT3 #(
		.INIT('h2a)
	) name12665 (
		\m1_data_i[24]_pad ,
		_w8989_,
		_w8990_,
		_w14566_
	);
	LUT3 #(
		.INIT('h57)
	) name12666 (
		_w9008_,
		_w14565_,
		_w14566_,
		_w14567_
	);
	LUT3 #(
		.INIT('h80)
	) name12667 (
		\m4_data_i[24]_pad ,
		_w8989_,
		_w8990_,
		_w14568_
	);
	LUT3 #(
		.INIT('h2a)
	) name12668 (
		\m7_data_i[24]_pad ,
		_w8989_,
		_w8990_,
		_w14569_
	);
	LUT4 #(
		.INIT('hcedf)
	) name12669 (
		_w8984_,
		_w8987_,
		_w14568_,
		_w14569_,
		_w14570_
	);
	LUT3 #(
		.INIT('h2a)
	) name12670 (
		\m5_data_i[24]_pad ,
		_w8989_,
		_w8990_,
		_w14571_
	);
	LUT3 #(
		.INIT('h80)
	) name12671 (
		\m6_data_i[24]_pad ,
		_w8989_,
		_w8990_,
		_w14572_
	);
	LUT4 #(
		.INIT('hcedf)
	) name12672 (
		_w8984_,
		_w8987_,
		_w14571_,
		_w14572_,
		_w14573_
	);
	LUT3 #(
		.INIT('h80)
	) name12673 (
		\m2_data_i[24]_pad ,
		_w8989_,
		_w8990_,
		_w14574_
	);
	LUT3 #(
		.INIT('h2a)
	) name12674 (
		\m3_data_i[24]_pad ,
		_w8989_,
		_w8990_,
		_w14575_
	);
	LUT3 #(
		.INIT('h57)
	) name12675 (
		_w9002_,
		_w14574_,
		_w14575_,
		_w14576_
	);
	LUT4 #(
		.INIT('h7fff)
	) name12676 (
		_w14567_,
		_w14570_,
		_w14573_,
		_w14576_,
		_w14577_
	);
	LUT3 #(
		.INIT('h80)
	) name12677 (
		\m0_data_i[25]_pad ,
		_w8989_,
		_w8990_,
		_w14578_
	);
	LUT3 #(
		.INIT('h2a)
	) name12678 (
		\m1_data_i[25]_pad ,
		_w8989_,
		_w8990_,
		_w14579_
	);
	LUT3 #(
		.INIT('h57)
	) name12679 (
		_w9008_,
		_w14578_,
		_w14579_,
		_w14580_
	);
	LUT3 #(
		.INIT('h80)
	) name12680 (
		\m6_data_i[25]_pad ,
		_w8989_,
		_w8990_,
		_w14581_
	);
	LUT3 #(
		.INIT('h2a)
	) name12681 (
		\m3_data_i[25]_pad ,
		_w8989_,
		_w8990_,
		_w14582_
	);
	LUT4 #(
		.INIT('habef)
	) name12682 (
		_w8984_,
		_w8987_,
		_w14581_,
		_w14582_,
		_w14583_
	);
	LUT3 #(
		.INIT('h2a)
	) name12683 (
		\m7_data_i[25]_pad ,
		_w8989_,
		_w8990_,
		_w14584_
	);
	LUT3 #(
		.INIT('h80)
	) name12684 (
		\m2_data_i[25]_pad ,
		_w8989_,
		_w8990_,
		_w14585_
	);
	LUT4 #(
		.INIT('habef)
	) name12685 (
		_w8984_,
		_w8987_,
		_w14584_,
		_w14585_,
		_w14586_
	);
	LUT3 #(
		.INIT('h80)
	) name12686 (
		\m4_data_i[25]_pad ,
		_w8989_,
		_w8990_,
		_w14587_
	);
	LUT3 #(
		.INIT('h2a)
	) name12687 (
		\m5_data_i[25]_pad ,
		_w8989_,
		_w8990_,
		_w14588_
	);
	LUT3 #(
		.INIT('h57)
	) name12688 (
		_w8996_,
		_w14587_,
		_w14588_,
		_w14589_
	);
	LUT4 #(
		.INIT('h7fff)
	) name12689 (
		_w14580_,
		_w14583_,
		_w14586_,
		_w14589_,
		_w14590_
	);
	LUT3 #(
		.INIT('h80)
	) name12690 (
		\m6_data_i[26]_pad ,
		_w8989_,
		_w8990_,
		_w14591_
	);
	LUT3 #(
		.INIT('h2a)
	) name12691 (
		\m7_data_i[26]_pad ,
		_w8989_,
		_w8990_,
		_w14592_
	);
	LUT3 #(
		.INIT('h57)
	) name12692 (
		_w8988_,
		_w14591_,
		_w14592_,
		_w14593_
	);
	LUT3 #(
		.INIT('h80)
	) name12693 (
		\m4_data_i[26]_pad ,
		_w8989_,
		_w8990_,
		_w14594_
	);
	LUT3 #(
		.INIT('h2a)
	) name12694 (
		\m1_data_i[26]_pad ,
		_w8989_,
		_w8990_,
		_w14595_
	);
	LUT4 #(
		.INIT('h57df)
	) name12695 (
		_w8984_,
		_w8987_,
		_w14594_,
		_w14595_,
		_w14596_
	);
	LUT3 #(
		.INIT('h2a)
	) name12696 (
		\m5_data_i[26]_pad ,
		_w8989_,
		_w8990_,
		_w14597_
	);
	LUT3 #(
		.INIT('h80)
	) name12697 (
		\m0_data_i[26]_pad ,
		_w8989_,
		_w8990_,
		_w14598_
	);
	LUT4 #(
		.INIT('h57df)
	) name12698 (
		_w8984_,
		_w8987_,
		_w14597_,
		_w14598_,
		_w14599_
	);
	LUT3 #(
		.INIT('h80)
	) name12699 (
		\m2_data_i[26]_pad ,
		_w8989_,
		_w8990_,
		_w14600_
	);
	LUT3 #(
		.INIT('h2a)
	) name12700 (
		\m3_data_i[26]_pad ,
		_w8989_,
		_w8990_,
		_w14601_
	);
	LUT3 #(
		.INIT('h57)
	) name12701 (
		_w9002_,
		_w14600_,
		_w14601_,
		_w14602_
	);
	LUT4 #(
		.INIT('h7fff)
	) name12702 (
		_w14593_,
		_w14596_,
		_w14599_,
		_w14602_,
		_w14603_
	);
	LUT3 #(
		.INIT('h80)
	) name12703 (
		\m6_data_i[27]_pad ,
		_w8989_,
		_w8990_,
		_w14604_
	);
	LUT3 #(
		.INIT('h2a)
	) name12704 (
		\m7_data_i[27]_pad ,
		_w8989_,
		_w8990_,
		_w14605_
	);
	LUT3 #(
		.INIT('h57)
	) name12705 (
		_w8988_,
		_w14604_,
		_w14605_,
		_w14606_
	);
	LUT3 #(
		.INIT('h80)
	) name12706 (
		\m4_data_i[27]_pad ,
		_w8989_,
		_w8990_,
		_w14607_
	);
	LUT3 #(
		.INIT('h2a)
	) name12707 (
		\m3_data_i[27]_pad ,
		_w8989_,
		_w8990_,
		_w14608_
	);
	LUT4 #(
		.INIT('h9bdf)
	) name12708 (
		_w8984_,
		_w8987_,
		_w14607_,
		_w14608_,
		_w14609_
	);
	LUT3 #(
		.INIT('h2a)
	) name12709 (
		\m5_data_i[27]_pad ,
		_w8989_,
		_w8990_,
		_w14610_
	);
	LUT3 #(
		.INIT('h80)
	) name12710 (
		\m2_data_i[27]_pad ,
		_w8989_,
		_w8990_,
		_w14611_
	);
	LUT4 #(
		.INIT('h9bdf)
	) name12711 (
		_w8984_,
		_w8987_,
		_w14610_,
		_w14611_,
		_w14612_
	);
	LUT3 #(
		.INIT('h80)
	) name12712 (
		\m0_data_i[27]_pad ,
		_w8989_,
		_w8990_,
		_w14613_
	);
	LUT3 #(
		.INIT('h2a)
	) name12713 (
		\m1_data_i[27]_pad ,
		_w8989_,
		_w8990_,
		_w14614_
	);
	LUT3 #(
		.INIT('h57)
	) name12714 (
		_w9008_,
		_w14613_,
		_w14614_,
		_w14615_
	);
	LUT4 #(
		.INIT('h7fff)
	) name12715 (
		_w14606_,
		_w14609_,
		_w14612_,
		_w14615_,
		_w14616_
	);
	LUT3 #(
		.INIT('h80)
	) name12716 (
		\m4_data_i[28]_pad ,
		_w8989_,
		_w8990_,
		_w14617_
	);
	LUT3 #(
		.INIT('h2a)
	) name12717 (
		\m5_data_i[28]_pad ,
		_w8989_,
		_w8990_,
		_w14618_
	);
	LUT3 #(
		.INIT('h57)
	) name12718 (
		_w8996_,
		_w14617_,
		_w14618_,
		_w14619_
	);
	LUT3 #(
		.INIT('h80)
	) name12719 (
		\m6_data_i[28]_pad ,
		_w8989_,
		_w8990_,
		_w14620_
	);
	LUT3 #(
		.INIT('h2a)
	) name12720 (
		\m1_data_i[28]_pad ,
		_w8989_,
		_w8990_,
		_w14621_
	);
	LUT4 #(
		.INIT('h67ef)
	) name12721 (
		_w8984_,
		_w8987_,
		_w14620_,
		_w14621_,
		_w14622_
	);
	LUT3 #(
		.INIT('h2a)
	) name12722 (
		\m7_data_i[28]_pad ,
		_w8989_,
		_w8990_,
		_w14623_
	);
	LUT3 #(
		.INIT('h80)
	) name12723 (
		\m0_data_i[28]_pad ,
		_w8989_,
		_w8990_,
		_w14624_
	);
	LUT4 #(
		.INIT('h67ef)
	) name12724 (
		_w8984_,
		_w8987_,
		_w14623_,
		_w14624_,
		_w14625_
	);
	LUT3 #(
		.INIT('h80)
	) name12725 (
		\m2_data_i[28]_pad ,
		_w8989_,
		_w8990_,
		_w14626_
	);
	LUT3 #(
		.INIT('h2a)
	) name12726 (
		\m3_data_i[28]_pad ,
		_w8989_,
		_w8990_,
		_w14627_
	);
	LUT3 #(
		.INIT('h57)
	) name12727 (
		_w9002_,
		_w14626_,
		_w14627_,
		_w14628_
	);
	LUT4 #(
		.INIT('h7fff)
	) name12728 (
		_w14619_,
		_w14622_,
		_w14625_,
		_w14628_,
		_w14629_
	);
	LUT3 #(
		.INIT('h80)
	) name12729 (
		\m6_data_i[29]_pad ,
		_w8989_,
		_w8990_,
		_w14630_
	);
	LUT3 #(
		.INIT('h2a)
	) name12730 (
		\m7_data_i[29]_pad ,
		_w8989_,
		_w8990_,
		_w14631_
	);
	LUT3 #(
		.INIT('h57)
	) name12731 (
		_w8988_,
		_w14630_,
		_w14631_,
		_w14632_
	);
	LUT3 #(
		.INIT('h80)
	) name12732 (
		\m4_data_i[29]_pad ,
		_w8989_,
		_w8990_,
		_w14633_
	);
	LUT3 #(
		.INIT('h2a)
	) name12733 (
		\m3_data_i[29]_pad ,
		_w8989_,
		_w8990_,
		_w14634_
	);
	LUT4 #(
		.INIT('h9bdf)
	) name12734 (
		_w8984_,
		_w8987_,
		_w14633_,
		_w14634_,
		_w14635_
	);
	LUT3 #(
		.INIT('h2a)
	) name12735 (
		\m5_data_i[29]_pad ,
		_w8989_,
		_w8990_,
		_w14636_
	);
	LUT3 #(
		.INIT('h80)
	) name12736 (
		\m2_data_i[29]_pad ,
		_w8989_,
		_w8990_,
		_w14637_
	);
	LUT4 #(
		.INIT('h9bdf)
	) name12737 (
		_w8984_,
		_w8987_,
		_w14636_,
		_w14637_,
		_w14638_
	);
	LUT3 #(
		.INIT('h80)
	) name12738 (
		\m0_data_i[29]_pad ,
		_w8989_,
		_w8990_,
		_w14639_
	);
	LUT3 #(
		.INIT('h2a)
	) name12739 (
		\m1_data_i[29]_pad ,
		_w8989_,
		_w8990_,
		_w14640_
	);
	LUT3 #(
		.INIT('h57)
	) name12740 (
		_w9008_,
		_w14639_,
		_w14640_,
		_w14641_
	);
	LUT4 #(
		.INIT('h7fff)
	) name12741 (
		_w14632_,
		_w14635_,
		_w14638_,
		_w14641_,
		_w14642_
	);
	LUT3 #(
		.INIT('h80)
	) name12742 (
		\m0_data_i[2]_pad ,
		_w8989_,
		_w8990_,
		_w14643_
	);
	LUT3 #(
		.INIT('h2a)
	) name12743 (
		\m1_data_i[2]_pad ,
		_w8989_,
		_w8990_,
		_w14644_
	);
	LUT3 #(
		.INIT('h57)
	) name12744 (
		_w9008_,
		_w14643_,
		_w14644_,
		_w14645_
	);
	LUT3 #(
		.INIT('h80)
	) name12745 (
		\m2_data_i[2]_pad ,
		_w8989_,
		_w8990_,
		_w14646_
	);
	LUT3 #(
		.INIT('h2a)
	) name12746 (
		\m7_data_i[2]_pad ,
		_w8989_,
		_w8990_,
		_w14647_
	);
	LUT4 #(
		.INIT('haebf)
	) name12747 (
		_w8984_,
		_w8987_,
		_w14646_,
		_w14647_,
		_w14648_
	);
	LUT3 #(
		.INIT('h2a)
	) name12748 (
		\m3_data_i[2]_pad ,
		_w8989_,
		_w8990_,
		_w14649_
	);
	LUT3 #(
		.INIT('h80)
	) name12749 (
		\m6_data_i[2]_pad ,
		_w8989_,
		_w8990_,
		_w14650_
	);
	LUT4 #(
		.INIT('haebf)
	) name12750 (
		_w8984_,
		_w8987_,
		_w14649_,
		_w14650_,
		_w14651_
	);
	LUT3 #(
		.INIT('h80)
	) name12751 (
		\m4_data_i[2]_pad ,
		_w8989_,
		_w8990_,
		_w14652_
	);
	LUT3 #(
		.INIT('h2a)
	) name12752 (
		\m5_data_i[2]_pad ,
		_w8989_,
		_w8990_,
		_w14653_
	);
	LUT3 #(
		.INIT('h57)
	) name12753 (
		_w8996_,
		_w14652_,
		_w14653_,
		_w14654_
	);
	LUT4 #(
		.INIT('h7fff)
	) name12754 (
		_w14645_,
		_w14648_,
		_w14651_,
		_w14654_,
		_w14655_
	);
	LUT3 #(
		.INIT('h80)
	) name12755 (
		\m4_data_i[30]_pad ,
		_w8989_,
		_w8990_,
		_w14656_
	);
	LUT3 #(
		.INIT('h2a)
	) name12756 (
		\m5_data_i[30]_pad ,
		_w8989_,
		_w8990_,
		_w14657_
	);
	LUT3 #(
		.INIT('h57)
	) name12757 (
		_w8996_,
		_w14656_,
		_w14657_,
		_w14658_
	);
	LUT3 #(
		.INIT('h80)
	) name12758 (
		\m0_data_i[30]_pad ,
		_w8989_,
		_w8990_,
		_w14659_
	);
	LUT3 #(
		.INIT('h2a)
	) name12759 (
		\m3_data_i[30]_pad ,
		_w8989_,
		_w8990_,
		_w14660_
	);
	LUT4 #(
		.INIT('h3b7f)
	) name12760 (
		_w8984_,
		_w8987_,
		_w14659_,
		_w14660_,
		_w14661_
	);
	LUT3 #(
		.INIT('h2a)
	) name12761 (
		\m1_data_i[30]_pad ,
		_w8989_,
		_w8990_,
		_w14662_
	);
	LUT3 #(
		.INIT('h80)
	) name12762 (
		\m2_data_i[30]_pad ,
		_w8989_,
		_w8990_,
		_w14663_
	);
	LUT4 #(
		.INIT('h3b7f)
	) name12763 (
		_w8984_,
		_w8987_,
		_w14662_,
		_w14663_,
		_w14664_
	);
	LUT3 #(
		.INIT('h80)
	) name12764 (
		\m6_data_i[30]_pad ,
		_w8989_,
		_w8990_,
		_w14665_
	);
	LUT3 #(
		.INIT('h2a)
	) name12765 (
		\m7_data_i[30]_pad ,
		_w8989_,
		_w8990_,
		_w14666_
	);
	LUT3 #(
		.INIT('h57)
	) name12766 (
		_w8988_,
		_w14665_,
		_w14666_,
		_w14667_
	);
	LUT4 #(
		.INIT('h7fff)
	) name12767 (
		_w14658_,
		_w14661_,
		_w14664_,
		_w14667_,
		_w14668_
	);
	LUT3 #(
		.INIT('h80)
	) name12768 (
		\m6_data_i[31]_pad ,
		_w8989_,
		_w8990_,
		_w14669_
	);
	LUT3 #(
		.INIT('h2a)
	) name12769 (
		\m7_data_i[31]_pad ,
		_w8989_,
		_w8990_,
		_w14670_
	);
	LUT3 #(
		.INIT('h57)
	) name12770 (
		_w8988_,
		_w14669_,
		_w14670_,
		_w14671_
	);
	LUT3 #(
		.INIT('h80)
	) name12771 (
		\m4_data_i[31]_pad ,
		_w8989_,
		_w8990_,
		_w14672_
	);
	LUT3 #(
		.INIT('h2a)
	) name12772 (
		\m3_data_i[31]_pad ,
		_w8989_,
		_w8990_,
		_w14673_
	);
	LUT4 #(
		.INIT('h9bdf)
	) name12773 (
		_w8984_,
		_w8987_,
		_w14672_,
		_w14673_,
		_w14674_
	);
	LUT3 #(
		.INIT('h2a)
	) name12774 (
		\m5_data_i[31]_pad ,
		_w8989_,
		_w8990_,
		_w14675_
	);
	LUT3 #(
		.INIT('h80)
	) name12775 (
		\m2_data_i[31]_pad ,
		_w8989_,
		_w8990_,
		_w14676_
	);
	LUT4 #(
		.INIT('h9bdf)
	) name12776 (
		_w8984_,
		_w8987_,
		_w14675_,
		_w14676_,
		_w14677_
	);
	LUT3 #(
		.INIT('h80)
	) name12777 (
		\m0_data_i[31]_pad ,
		_w8989_,
		_w8990_,
		_w14678_
	);
	LUT3 #(
		.INIT('h2a)
	) name12778 (
		\m1_data_i[31]_pad ,
		_w8989_,
		_w8990_,
		_w14679_
	);
	LUT3 #(
		.INIT('h57)
	) name12779 (
		_w9008_,
		_w14678_,
		_w14679_,
		_w14680_
	);
	LUT4 #(
		.INIT('h7fff)
	) name12780 (
		_w14671_,
		_w14674_,
		_w14677_,
		_w14680_,
		_w14681_
	);
	LUT3 #(
		.INIT('h80)
	) name12781 (
		\m0_data_i[3]_pad ,
		_w8989_,
		_w8990_,
		_w14682_
	);
	LUT3 #(
		.INIT('h2a)
	) name12782 (
		\m1_data_i[3]_pad ,
		_w8989_,
		_w8990_,
		_w14683_
	);
	LUT3 #(
		.INIT('h57)
	) name12783 (
		_w9008_,
		_w14682_,
		_w14683_,
		_w14684_
	);
	LUT3 #(
		.INIT('h80)
	) name12784 (
		\m4_data_i[3]_pad ,
		_w8989_,
		_w8990_,
		_w14685_
	);
	LUT3 #(
		.INIT('h2a)
	) name12785 (
		\m3_data_i[3]_pad ,
		_w8989_,
		_w8990_,
		_w14686_
	);
	LUT4 #(
		.INIT('h9bdf)
	) name12786 (
		_w8984_,
		_w8987_,
		_w14685_,
		_w14686_,
		_w14687_
	);
	LUT3 #(
		.INIT('h2a)
	) name12787 (
		\m5_data_i[3]_pad ,
		_w8989_,
		_w8990_,
		_w14688_
	);
	LUT3 #(
		.INIT('h80)
	) name12788 (
		\m2_data_i[3]_pad ,
		_w8989_,
		_w8990_,
		_w14689_
	);
	LUT4 #(
		.INIT('h9bdf)
	) name12789 (
		_w8984_,
		_w8987_,
		_w14688_,
		_w14689_,
		_w14690_
	);
	LUT3 #(
		.INIT('h80)
	) name12790 (
		\m6_data_i[3]_pad ,
		_w8989_,
		_w8990_,
		_w14691_
	);
	LUT3 #(
		.INIT('h2a)
	) name12791 (
		\m7_data_i[3]_pad ,
		_w8989_,
		_w8990_,
		_w14692_
	);
	LUT3 #(
		.INIT('h57)
	) name12792 (
		_w8988_,
		_w14691_,
		_w14692_,
		_w14693_
	);
	LUT4 #(
		.INIT('h7fff)
	) name12793 (
		_w14684_,
		_w14687_,
		_w14690_,
		_w14693_,
		_w14694_
	);
	LUT3 #(
		.INIT('h80)
	) name12794 (
		\m2_data_i[4]_pad ,
		_w8989_,
		_w8990_,
		_w14695_
	);
	LUT3 #(
		.INIT('h2a)
	) name12795 (
		\m3_data_i[4]_pad ,
		_w8989_,
		_w8990_,
		_w14696_
	);
	LUT3 #(
		.INIT('h57)
	) name12796 (
		_w9002_,
		_w14695_,
		_w14696_,
		_w14697_
	);
	LUT3 #(
		.INIT('h80)
	) name12797 (
		\m4_data_i[4]_pad ,
		_w8989_,
		_w8990_,
		_w14698_
	);
	LUT3 #(
		.INIT('h2a)
	) name12798 (
		\m1_data_i[4]_pad ,
		_w8989_,
		_w8990_,
		_w14699_
	);
	LUT4 #(
		.INIT('h57df)
	) name12799 (
		_w8984_,
		_w8987_,
		_w14698_,
		_w14699_,
		_w14700_
	);
	LUT3 #(
		.INIT('h2a)
	) name12800 (
		\m5_data_i[4]_pad ,
		_w8989_,
		_w8990_,
		_w14701_
	);
	LUT3 #(
		.INIT('h80)
	) name12801 (
		\m0_data_i[4]_pad ,
		_w8989_,
		_w8990_,
		_w14702_
	);
	LUT4 #(
		.INIT('h57df)
	) name12802 (
		_w8984_,
		_w8987_,
		_w14701_,
		_w14702_,
		_w14703_
	);
	LUT3 #(
		.INIT('h80)
	) name12803 (
		\m6_data_i[4]_pad ,
		_w8989_,
		_w8990_,
		_w14704_
	);
	LUT3 #(
		.INIT('h2a)
	) name12804 (
		\m7_data_i[4]_pad ,
		_w8989_,
		_w8990_,
		_w14705_
	);
	LUT3 #(
		.INIT('h57)
	) name12805 (
		_w8988_,
		_w14704_,
		_w14705_,
		_w14706_
	);
	LUT4 #(
		.INIT('h7fff)
	) name12806 (
		_w14697_,
		_w14700_,
		_w14703_,
		_w14706_,
		_w14707_
	);
	LUT3 #(
		.INIT('h80)
	) name12807 (
		\m6_data_i[5]_pad ,
		_w8989_,
		_w8990_,
		_w14708_
	);
	LUT3 #(
		.INIT('h2a)
	) name12808 (
		\m7_data_i[5]_pad ,
		_w8989_,
		_w8990_,
		_w14709_
	);
	LUT3 #(
		.INIT('h57)
	) name12809 (
		_w8988_,
		_w14708_,
		_w14709_,
		_w14710_
	);
	LUT3 #(
		.INIT('h80)
	) name12810 (
		\m4_data_i[5]_pad ,
		_w8989_,
		_w8990_,
		_w14711_
	);
	LUT3 #(
		.INIT('h2a)
	) name12811 (
		\m3_data_i[5]_pad ,
		_w8989_,
		_w8990_,
		_w14712_
	);
	LUT4 #(
		.INIT('h9bdf)
	) name12812 (
		_w8984_,
		_w8987_,
		_w14711_,
		_w14712_,
		_w14713_
	);
	LUT3 #(
		.INIT('h2a)
	) name12813 (
		\m5_data_i[5]_pad ,
		_w8989_,
		_w8990_,
		_w14714_
	);
	LUT3 #(
		.INIT('h80)
	) name12814 (
		\m2_data_i[5]_pad ,
		_w8989_,
		_w8990_,
		_w14715_
	);
	LUT4 #(
		.INIT('h9bdf)
	) name12815 (
		_w8984_,
		_w8987_,
		_w14714_,
		_w14715_,
		_w14716_
	);
	LUT3 #(
		.INIT('h80)
	) name12816 (
		\m0_data_i[5]_pad ,
		_w8989_,
		_w8990_,
		_w14717_
	);
	LUT3 #(
		.INIT('h2a)
	) name12817 (
		\m1_data_i[5]_pad ,
		_w8989_,
		_w8990_,
		_w14718_
	);
	LUT3 #(
		.INIT('h57)
	) name12818 (
		_w9008_,
		_w14717_,
		_w14718_,
		_w14719_
	);
	LUT4 #(
		.INIT('h7fff)
	) name12819 (
		_w14710_,
		_w14713_,
		_w14716_,
		_w14719_,
		_w14720_
	);
	LUT3 #(
		.INIT('h80)
	) name12820 (
		\m2_data_i[6]_pad ,
		_w8989_,
		_w8990_,
		_w14721_
	);
	LUT3 #(
		.INIT('h2a)
	) name12821 (
		\m3_data_i[6]_pad ,
		_w8989_,
		_w8990_,
		_w14722_
	);
	LUT3 #(
		.INIT('h57)
	) name12822 (
		_w9002_,
		_w14721_,
		_w14722_,
		_w14723_
	);
	LUT3 #(
		.INIT('h80)
	) name12823 (
		\m6_data_i[6]_pad ,
		_w8989_,
		_w8990_,
		_w14724_
	);
	LUT3 #(
		.INIT('h2a)
	) name12824 (
		\m1_data_i[6]_pad ,
		_w8989_,
		_w8990_,
		_w14725_
	);
	LUT4 #(
		.INIT('h67ef)
	) name12825 (
		_w8984_,
		_w8987_,
		_w14724_,
		_w14725_,
		_w14726_
	);
	LUT3 #(
		.INIT('h2a)
	) name12826 (
		\m7_data_i[6]_pad ,
		_w8989_,
		_w8990_,
		_w14727_
	);
	LUT3 #(
		.INIT('h80)
	) name12827 (
		\m0_data_i[6]_pad ,
		_w8989_,
		_w8990_,
		_w14728_
	);
	LUT4 #(
		.INIT('h67ef)
	) name12828 (
		_w8984_,
		_w8987_,
		_w14727_,
		_w14728_,
		_w14729_
	);
	LUT3 #(
		.INIT('h80)
	) name12829 (
		\m4_data_i[6]_pad ,
		_w8989_,
		_w8990_,
		_w14730_
	);
	LUT3 #(
		.INIT('h2a)
	) name12830 (
		\m5_data_i[6]_pad ,
		_w8989_,
		_w8990_,
		_w14731_
	);
	LUT3 #(
		.INIT('h57)
	) name12831 (
		_w8996_,
		_w14730_,
		_w14731_,
		_w14732_
	);
	LUT4 #(
		.INIT('h7fff)
	) name12832 (
		_w14723_,
		_w14726_,
		_w14729_,
		_w14732_,
		_w14733_
	);
	LUT3 #(
		.INIT('h80)
	) name12833 (
		\m6_data_i[7]_pad ,
		_w8989_,
		_w8990_,
		_w14734_
	);
	LUT3 #(
		.INIT('h2a)
	) name12834 (
		\m7_data_i[7]_pad ,
		_w8989_,
		_w8990_,
		_w14735_
	);
	LUT3 #(
		.INIT('h57)
	) name12835 (
		_w8988_,
		_w14734_,
		_w14735_,
		_w14736_
	);
	LUT3 #(
		.INIT('h80)
	) name12836 (
		\m4_data_i[7]_pad ,
		_w8989_,
		_w8990_,
		_w14737_
	);
	LUT3 #(
		.INIT('h2a)
	) name12837 (
		\m1_data_i[7]_pad ,
		_w8989_,
		_w8990_,
		_w14738_
	);
	LUT4 #(
		.INIT('h57df)
	) name12838 (
		_w8984_,
		_w8987_,
		_w14737_,
		_w14738_,
		_w14739_
	);
	LUT3 #(
		.INIT('h2a)
	) name12839 (
		\m5_data_i[7]_pad ,
		_w8989_,
		_w8990_,
		_w14740_
	);
	LUT3 #(
		.INIT('h80)
	) name12840 (
		\m0_data_i[7]_pad ,
		_w8989_,
		_w8990_,
		_w14741_
	);
	LUT4 #(
		.INIT('h57df)
	) name12841 (
		_w8984_,
		_w8987_,
		_w14740_,
		_w14741_,
		_w14742_
	);
	LUT3 #(
		.INIT('h80)
	) name12842 (
		\m2_data_i[7]_pad ,
		_w8989_,
		_w8990_,
		_w14743_
	);
	LUT3 #(
		.INIT('h2a)
	) name12843 (
		\m3_data_i[7]_pad ,
		_w8989_,
		_w8990_,
		_w14744_
	);
	LUT3 #(
		.INIT('h57)
	) name12844 (
		_w9002_,
		_w14743_,
		_w14744_,
		_w14745_
	);
	LUT4 #(
		.INIT('h7fff)
	) name12845 (
		_w14736_,
		_w14739_,
		_w14742_,
		_w14745_,
		_w14746_
	);
	LUT3 #(
		.INIT('h80)
	) name12846 (
		\m6_data_i[8]_pad ,
		_w8989_,
		_w8990_,
		_w14747_
	);
	LUT3 #(
		.INIT('h2a)
	) name12847 (
		\m7_data_i[8]_pad ,
		_w8989_,
		_w8990_,
		_w14748_
	);
	LUT3 #(
		.INIT('h57)
	) name12848 (
		_w8988_,
		_w14747_,
		_w14748_,
		_w14749_
	);
	LUT3 #(
		.INIT('h80)
	) name12849 (
		\m4_data_i[8]_pad ,
		_w8989_,
		_w8990_,
		_w14750_
	);
	LUT3 #(
		.INIT('h2a)
	) name12850 (
		\m1_data_i[8]_pad ,
		_w8989_,
		_w8990_,
		_w14751_
	);
	LUT4 #(
		.INIT('h57df)
	) name12851 (
		_w8984_,
		_w8987_,
		_w14750_,
		_w14751_,
		_w14752_
	);
	LUT3 #(
		.INIT('h2a)
	) name12852 (
		\m5_data_i[8]_pad ,
		_w8989_,
		_w8990_,
		_w14753_
	);
	LUT3 #(
		.INIT('h80)
	) name12853 (
		\m0_data_i[8]_pad ,
		_w8989_,
		_w8990_,
		_w14754_
	);
	LUT4 #(
		.INIT('h57df)
	) name12854 (
		_w8984_,
		_w8987_,
		_w14753_,
		_w14754_,
		_w14755_
	);
	LUT3 #(
		.INIT('h80)
	) name12855 (
		\m2_data_i[8]_pad ,
		_w8989_,
		_w8990_,
		_w14756_
	);
	LUT3 #(
		.INIT('h2a)
	) name12856 (
		\m3_data_i[8]_pad ,
		_w8989_,
		_w8990_,
		_w14757_
	);
	LUT3 #(
		.INIT('h57)
	) name12857 (
		_w9002_,
		_w14756_,
		_w14757_,
		_w14758_
	);
	LUT4 #(
		.INIT('h7fff)
	) name12858 (
		_w14749_,
		_w14752_,
		_w14755_,
		_w14758_,
		_w14759_
	);
	LUT3 #(
		.INIT('h80)
	) name12859 (
		\m6_data_i[9]_pad ,
		_w8989_,
		_w8990_,
		_w14760_
	);
	LUT3 #(
		.INIT('h2a)
	) name12860 (
		\m7_data_i[9]_pad ,
		_w8989_,
		_w8990_,
		_w14761_
	);
	LUT3 #(
		.INIT('h57)
	) name12861 (
		_w8988_,
		_w14760_,
		_w14761_,
		_w14762_
	);
	LUT3 #(
		.INIT('h80)
	) name12862 (
		\m4_data_i[9]_pad ,
		_w8989_,
		_w8990_,
		_w14763_
	);
	LUT3 #(
		.INIT('h2a)
	) name12863 (
		\m1_data_i[9]_pad ,
		_w8989_,
		_w8990_,
		_w14764_
	);
	LUT4 #(
		.INIT('h57df)
	) name12864 (
		_w8984_,
		_w8987_,
		_w14763_,
		_w14764_,
		_w14765_
	);
	LUT3 #(
		.INIT('h2a)
	) name12865 (
		\m5_data_i[9]_pad ,
		_w8989_,
		_w8990_,
		_w14766_
	);
	LUT3 #(
		.INIT('h80)
	) name12866 (
		\m0_data_i[9]_pad ,
		_w8989_,
		_w8990_,
		_w14767_
	);
	LUT4 #(
		.INIT('h57df)
	) name12867 (
		_w8984_,
		_w8987_,
		_w14766_,
		_w14767_,
		_w14768_
	);
	LUT3 #(
		.INIT('h80)
	) name12868 (
		\m2_data_i[9]_pad ,
		_w8989_,
		_w8990_,
		_w14769_
	);
	LUT3 #(
		.INIT('h2a)
	) name12869 (
		\m3_data_i[9]_pad ,
		_w8989_,
		_w8990_,
		_w14770_
	);
	LUT3 #(
		.INIT('h57)
	) name12870 (
		_w9002_,
		_w14769_,
		_w14770_,
		_w14771_
	);
	LUT4 #(
		.INIT('h7fff)
	) name12871 (
		_w14762_,
		_w14765_,
		_w14768_,
		_w14771_,
		_w14772_
	);
	LUT3 #(
		.INIT('h80)
	) name12872 (
		\m2_sel_i[0]_pad ,
		_w8989_,
		_w8990_,
		_w14773_
	);
	LUT3 #(
		.INIT('h2a)
	) name12873 (
		\m3_sel_i[0]_pad ,
		_w8989_,
		_w8990_,
		_w14774_
	);
	LUT3 #(
		.INIT('h57)
	) name12874 (
		_w9002_,
		_w14773_,
		_w14774_,
		_w14775_
	);
	LUT3 #(
		.INIT('h80)
	) name12875 (
		\m0_sel_i[0]_pad ,
		_w8989_,
		_w8990_,
		_w14776_
	);
	LUT3 #(
		.INIT('h2a)
	) name12876 (
		\m7_sel_i[0]_pad ,
		_w8989_,
		_w8990_,
		_w14777_
	);
	LUT4 #(
		.INIT('h6e7f)
	) name12877 (
		_w8984_,
		_w8987_,
		_w14776_,
		_w14777_,
		_w14778_
	);
	LUT3 #(
		.INIT('h2a)
	) name12878 (
		\m1_sel_i[0]_pad ,
		_w8989_,
		_w8990_,
		_w14779_
	);
	LUT3 #(
		.INIT('h80)
	) name12879 (
		\m6_sel_i[0]_pad ,
		_w8989_,
		_w8990_,
		_w14780_
	);
	LUT4 #(
		.INIT('h6e7f)
	) name12880 (
		_w8984_,
		_w8987_,
		_w14779_,
		_w14780_,
		_w14781_
	);
	LUT3 #(
		.INIT('h80)
	) name12881 (
		\m4_sel_i[0]_pad ,
		_w8989_,
		_w8990_,
		_w14782_
	);
	LUT3 #(
		.INIT('h2a)
	) name12882 (
		\m5_sel_i[0]_pad ,
		_w8989_,
		_w8990_,
		_w14783_
	);
	LUT3 #(
		.INIT('h57)
	) name12883 (
		_w8996_,
		_w14782_,
		_w14783_,
		_w14784_
	);
	LUT4 #(
		.INIT('h7fff)
	) name12884 (
		_w14775_,
		_w14778_,
		_w14781_,
		_w14784_,
		_w14785_
	);
	LUT3 #(
		.INIT('h80)
	) name12885 (
		\m0_sel_i[1]_pad ,
		_w8989_,
		_w8990_,
		_w14786_
	);
	LUT3 #(
		.INIT('h2a)
	) name12886 (
		\m1_sel_i[1]_pad ,
		_w8989_,
		_w8990_,
		_w14787_
	);
	LUT3 #(
		.INIT('h57)
	) name12887 (
		_w9008_,
		_w14786_,
		_w14787_,
		_w14788_
	);
	LUT3 #(
		.INIT('h80)
	) name12888 (
		\m6_sel_i[1]_pad ,
		_w8989_,
		_w8990_,
		_w14789_
	);
	LUT3 #(
		.INIT('h2a)
	) name12889 (
		\m3_sel_i[1]_pad ,
		_w8989_,
		_w8990_,
		_w14790_
	);
	LUT4 #(
		.INIT('habef)
	) name12890 (
		_w8984_,
		_w8987_,
		_w14789_,
		_w14790_,
		_w14791_
	);
	LUT3 #(
		.INIT('h2a)
	) name12891 (
		\m7_sel_i[1]_pad ,
		_w8989_,
		_w8990_,
		_w14792_
	);
	LUT3 #(
		.INIT('h80)
	) name12892 (
		\m2_sel_i[1]_pad ,
		_w8989_,
		_w8990_,
		_w14793_
	);
	LUT4 #(
		.INIT('habef)
	) name12893 (
		_w8984_,
		_w8987_,
		_w14792_,
		_w14793_,
		_w14794_
	);
	LUT3 #(
		.INIT('h80)
	) name12894 (
		\m4_sel_i[1]_pad ,
		_w8989_,
		_w8990_,
		_w14795_
	);
	LUT3 #(
		.INIT('h2a)
	) name12895 (
		\m5_sel_i[1]_pad ,
		_w8989_,
		_w8990_,
		_w14796_
	);
	LUT3 #(
		.INIT('h57)
	) name12896 (
		_w8996_,
		_w14795_,
		_w14796_,
		_w14797_
	);
	LUT4 #(
		.INIT('h7fff)
	) name12897 (
		_w14788_,
		_w14791_,
		_w14794_,
		_w14797_,
		_w14798_
	);
	LUT3 #(
		.INIT('h80)
	) name12898 (
		\m2_sel_i[2]_pad ,
		_w8989_,
		_w8990_,
		_w14799_
	);
	LUT3 #(
		.INIT('h2a)
	) name12899 (
		\m3_sel_i[2]_pad ,
		_w8989_,
		_w8990_,
		_w14800_
	);
	LUT3 #(
		.INIT('h57)
	) name12900 (
		_w9002_,
		_w14799_,
		_w14800_,
		_w14801_
	);
	LUT3 #(
		.INIT('h80)
	) name12901 (
		\m0_sel_i[2]_pad ,
		_w8989_,
		_w8990_,
		_w14802_
	);
	LUT3 #(
		.INIT('h2a)
	) name12902 (
		\m5_sel_i[2]_pad ,
		_w8989_,
		_w8990_,
		_w14803_
	);
	LUT4 #(
		.INIT('h5d7f)
	) name12903 (
		_w8984_,
		_w8987_,
		_w14802_,
		_w14803_,
		_w14804_
	);
	LUT3 #(
		.INIT('h2a)
	) name12904 (
		\m1_sel_i[2]_pad ,
		_w8989_,
		_w8990_,
		_w14805_
	);
	LUT3 #(
		.INIT('h80)
	) name12905 (
		\m4_sel_i[2]_pad ,
		_w8989_,
		_w8990_,
		_w14806_
	);
	LUT4 #(
		.INIT('h5d7f)
	) name12906 (
		_w8984_,
		_w8987_,
		_w14805_,
		_w14806_,
		_w14807_
	);
	LUT3 #(
		.INIT('h80)
	) name12907 (
		\m6_sel_i[2]_pad ,
		_w8989_,
		_w8990_,
		_w14808_
	);
	LUT3 #(
		.INIT('h2a)
	) name12908 (
		\m7_sel_i[2]_pad ,
		_w8989_,
		_w8990_,
		_w14809_
	);
	LUT3 #(
		.INIT('h57)
	) name12909 (
		_w8988_,
		_w14808_,
		_w14809_,
		_w14810_
	);
	LUT4 #(
		.INIT('h7fff)
	) name12910 (
		_w14801_,
		_w14804_,
		_w14807_,
		_w14810_,
		_w14811_
	);
	LUT3 #(
		.INIT('h80)
	) name12911 (
		\m2_sel_i[3]_pad ,
		_w8989_,
		_w8990_,
		_w14812_
	);
	LUT3 #(
		.INIT('h2a)
	) name12912 (
		\m3_sel_i[3]_pad ,
		_w8989_,
		_w8990_,
		_w14813_
	);
	LUT3 #(
		.INIT('h57)
	) name12913 (
		_w9002_,
		_w14812_,
		_w14813_,
		_w14814_
	);
	LUT3 #(
		.INIT('h80)
	) name12914 (
		\m0_sel_i[3]_pad ,
		_w8989_,
		_w8990_,
		_w14815_
	);
	LUT3 #(
		.INIT('h2a)
	) name12915 (
		\m7_sel_i[3]_pad ,
		_w8989_,
		_w8990_,
		_w14816_
	);
	LUT4 #(
		.INIT('h6e7f)
	) name12916 (
		_w8984_,
		_w8987_,
		_w14815_,
		_w14816_,
		_w14817_
	);
	LUT3 #(
		.INIT('h2a)
	) name12917 (
		\m1_sel_i[3]_pad ,
		_w8989_,
		_w8990_,
		_w14818_
	);
	LUT3 #(
		.INIT('h80)
	) name12918 (
		\m6_sel_i[3]_pad ,
		_w8989_,
		_w8990_,
		_w14819_
	);
	LUT4 #(
		.INIT('h6e7f)
	) name12919 (
		_w8984_,
		_w8987_,
		_w14818_,
		_w14819_,
		_w14820_
	);
	LUT3 #(
		.INIT('h80)
	) name12920 (
		\m4_sel_i[3]_pad ,
		_w8989_,
		_w8990_,
		_w14821_
	);
	LUT3 #(
		.INIT('h2a)
	) name12921 (
		\m5_sel_i[3]_pad ,
		_w8989_,
		_w8990_,
		_w14822_
	);
	LUT3 #(
		.INIT('h57)
	) name12922 (
		_w8996_,
		_w14821_,
		_w14822_,
		_w14823_
	);
	LUT4 #(
		.INIT('h7fff)
	) name12923 (
		_w14814_,
		_w14817_,
		_w14820_,
		_w14823_,
		_w14824_
	);
	LUT4 #(
		.INIT('h2a00)
	) name12924 (
		\m1_stb_i_pad ,
		_w8989_,
		_w8990_,
		_w9280_,
		_w14825_
	);
	LUT4 #(
		.INIT('h2a00)
	) name12925 (
		\m7_stb_i_pad ,
		_w8989_,
		_w8990_,
		_w9315_,
		_w14826_
	);
	LUT4 #(
		.INIT('h6e7f)
	) name12926 (
		_w8984_,
		_w8987_,
		_w14825_,
		_w14826_,
		_w14827_
	);
	LUT4 #(
		.INIT('h8000)
	) name12927 (
		\m2_stb_i_pad ,
		_w8989_,
		_w8990_,
		_w9284_,
		_w14828_
	);
	LUT4 #(
		.INIT('h2a00)
	) name12928 (
		\m3_stb_i_pad ,
		_w8989_,
		_w8990_,
		_w9291_,
		_w14829_
	);
	LUT3 #(
		.INIT('h57)
	) name12929 (
		_w9002_,
		_w14828_,
		_w14829_,
		_w14830_
	);
	LUT4 #(
		.INIT('h8000)
	) name12930 (
		\m0_stb_i_pad ,
		_w8989_,
		_w8990_,
		_w9273_,
		_w14831_
	);
	LUT4 #(
		.INIT('h2a00)
	) name12931 (
		\m5_stb_i_pad ,
		_w8989_,
		_w8990_,
		_w9305_,
		_w14832_
	);
	LUT4 #(
		.INIT('h5d7f)
	) name12932 (
		_w8984_,
		_w8987_,
		_w14831_,
		_w14832_,
		_w14833_
	);
	LUT4 #(
		.INIT('h8000)
	) name12933 (
		\m4_stb_i_pad ,
		_w8989_,
		_w8990_,
		_w9298_,
		_w14834_
	);
	LUT4 #(
		.INIT('h8000)
	) name12934 (
		\m6_stb_i_pad ,
		_w8989_,
		_w8990_,
		_w9308_,
		_w14835_
	);
	LUT4 #(
		.INIT('hcedf)
	) name12935 (
		_w8984_,
		_w8987_,
		_w14834_,
		_w14835_,
		_w14836_
	);
	LUT4 #(
		.INIT('h7fff)
	) name12936 (
		_w14827_,
		_w14830_,
		_w14833_,
		_w14836_,
		_w14837_
	);
	LUT3 #(
		.INIT('h80)
	) name12937 (
		\m2_we_i_pad ,
		_w8989_,
		_w8990_,
		_w14838_
	);
	LUT3 #(
		.INIT('h2a)
	) name12938 (
		\m3_we_i_pad ,
		_w8989_,
		_w8990_,
		_w14839_
	);
	LUT3 #(
		.INIT('h57)
	) name12939 (
		_w9002_,
		_w14838_,
		_w14839_,
		_w14840_
	);
	LUT3 #(
		.INIT('h80)
	) name12940 (
		\m0_we_i_pad ,
		_w8989_,
		_w8990_,
		_w14841_
	);
	LUT3 #(
		.INIT('h2a)
	) name12941 (
		\m7_we_i_pad ,
		_w8989_,
		_w8990_,
		_w14842_
	);
	LUT4 #(
		.INIT('h6e7f)
	) name12942 (
		_w8984_,
		_w8987_,
		_w14841_,
		_w14842_,
		_w14843_
	);
	LUT3 #(
		.INIT('h2a)
	) name12943 (
		\m1_we_i_pad ,
		_w8989_,
		_w8990_,
		_w14844_
	);
	LUT3 #(
		.INIT('h80)
	) name12944 (
		\m6_we_i_pad ,
		_w8989_,
		_w8990_,
		_w14845_
	);
	LUT4 #(
		.INIT('h6e7f)
	) name12945 (
		_w8984_,
		_w8987_,
		_w14844_,
		_w14845_,
		_w14846_
	);
	LUT3 #(
		.INIT('h80)
	) name12946 (
		\m4_we_i_pad ,
		_w8989_,
		_w8990_,
		_w14847_
	);
	LUT3 #(
		.INIT('h2a)
	) name12947 (
		\m5_we_i_pad ,
		_w8989_,
		_w8990_,
		_w14848_
	);
	LUT3 #(
		.INIT('h57)
	) name12948 (
		_w8996_,
		_w14847_,
		_w14848_,
		_w14849_
	);
	LUT4 #(
		.INIT('h7fff)
	) name12949 (
		_w14840_,
		_w14843_,
		_w14846_,
		_w14849_,
		_w14850_
	);
	LUT3 #(
		.INIT('h2a)
	) name12950 (
		\m1_addr_i[0]_pad ,
		_w8910_,
		_w8911_,
		_w14851_
	);
	LUT3 #(
		.INIT('h80)
	) name12951 (
		\m2_addr_i[0]_pad ,
		_w8910_,
		_w8911_,
		_w14852_
	);
	LUT4 #(
		.INIT('h3b7f)
	) name12952 (
		_w8905_,
		_w8908_,
		_w14851_,
		_w14852_,
		_w14853_
	);
	LUT3 #(
		.INIT('h80)
	) name12953 (
		\m0_addr_i[0]_pad ,
		_w8910_,
		_w8911_,
		_w14854_
	);
	LUT3 #(
		.INIT('h80)
	) name12954 (
		\m4_addr_i[0]_pad ,
		_w8910_,
		_w8911_,
		_w14855_
	);
	LUT4 #(
		.INIT('h5d7f)
	) name12955 (
		_w8905_,
		_w8908_,
		_w14854_,
		_w14855_,
		_w14856_
	);
	LUT3 #(
		.INIT('h2a)
	) name12956 (
		\m7_addr_i[0]_pad ,
		_w8910_,
		_w8911_,
		_w14857_
	);
	LUT3 #(
		.INIT('h2a)
	) name12957 (
		\m3_addr_i[0]_pad ,
		_w8910_,
		_w8911_,
		_w14858_
	);
	LUT4 #(
		.INIT('habef)
	) name12958 (
		_w8905_,
		_w8908_,
		_w14857_,
		_w14858_,
		_w14859_
	);
	LUT3 #(
		.INIT('h80)
	) name12959 (
		\m6_addr_i[0]_pad ,
		_w8910_,
		_w8911_,
		_w14860_
	);
	LUT3 #(
		.INIT('h2a)
	) name12960 (
		\m5_addr_i[0]_pad ,
		_w8910_,
		_w8911_,
		_w14861_
	);
	LUT4 #(
		.INIT('hcdef)
	) name12961 (
		_w8905_,
		_w8908_,
		_w14860_,
		_w14861_,
		_w14862_
	);
	LUT4 #(
		.INIT('h7fff)
	) name12962 (
		_w14853_,
		_w14856_,
		_w14859_,
		_w14862_,
		_w14863_
	);
	LUT3 #(
		.INIT('h2a)
	) name12963 (
		\m1_addr_i[10]_pad ,
		_w8910_,
		_w8911_,
		_w14864_
	);
	LUT3 #(
		.INIT('h80)
	) name12964 (
		\m2_addr_i[10]_pad ,
		_w8910_,
		_w8911_,
		_w14865_
	);
	LUT4 #(
		.INIT('h3b7f)
	) name12965 (
		_w8905_,
		_w8908_,
		_w14864_,
		_w14865_,
		_w14866_
	);
	LUT3 #(
		.INIT('h80)
	) name12966 (
		\m6_addr_i[10]_pad ,
		_w8910_,
		_w8911_,
		_w14867_
	);
	LUT3 #(
		.INIT('h80)
	) name12967 (
		\m4_addr_i[10]_pad ,
		_w8910_,
		_w8911_,
		_w14868_
	);
	LUT4 #(
		.INIT('hcdef)
	) name12968 (
		_w8905_,
		_w8908_,
		_w14867_,
		_w14868_,
		_w14869_
	);
	LUT3 #(
		.INIT('h2a)
	) name12969 (
		\m5_addr_i[10]_pad ,
		_w8910_,
		_w8911_,
		_w14870_
	);
	LUT3 #(
		.INIT('h2a)
	) name12970 (
		\m3_addr_i[10]_pad ,
		_w8910_,
		_w8911_,
		_w14871_
	);
	LUT4 #(
		.INIT('h9bdf)
	) name12971 (
		_w8905_,
		_w8908_,
		_w14870_,
		_w14871_,
		_w14872_
	);
	LUT3 #(
		.INIT('h80)
	) name12972 (
		\m0_addr_i[10]_pad ,
		_w8910_,
		_w8911_,
		_w14873_
	);
	LUT3 #(
		.INIT('h2a)
	) name12973 (
		\m7_addr_i[10]_pad ,
		_w8910_,
		_w8911_,
		_w14874_
	);
	LUT4 #(
		.INIT('h6e7f)
	) name12974 (
		_w8905_,
		_w8908_,
		_w14873_,
		_w14874_,
		_w14875_
	);
	LUT4 #(
		.INIT('h7fff)
	) name12975 (
		_w14866_,
		_w14869_,
		_w14872_,
		_w14875_,
		_w14876_
	);
	LUT3 #(
		.INIT('h2a)
	) name12976 (
		\m3_addr_i[11]_pad ,
		_w8910_,
		_w8911_,
		_w14877_
	);
	LUT3 #(
		.INIT('h80)
	) name12977 (
		\m4_addr_i[11]_pad ,
		_w8910_,
		_w8911_,
		_w14878_
	);
	LUT4 #(
		.INIT('h9dbf)
	) name12978 (
		_w8905_,
		_w8908_,
		_w14877_,
		_w14878_,
		_w14879_
	);
	LUT3 #(
		.INIT('h80)
	) name12979 (
		\m0_addr_i[11]_pad ,
		_w8910_,
		_w8911_,
		_w14880_
	);
	LUT3 #(
		.INIT('h80)
	) name12980 (
		\m2_addr_i[11]_pad ,
		_w8910_,
		_w8911_,
		_w14881_
	);
	LUT4 #(
		.INIT('h3b7f)
	) name12981 (
		_w8905_,
		_w8908_,
		_w14880_,
		_w14881_,
		_w14882_
	);
	LUT3 #(
		.INIT('h2a)
	) name12982 (
		\m7_addr_i[11]_pad ,
		_w8910_,
		_w8911_,
		_w14883_
	);
	LUT3 #(
		.INIT('h2a)
	) name12983 (
		\m1_addr_i[11]_pad ,
		_w8910_,
		_w8911_,
		_w14884_
	);
	LUT4 #(
		.INIT('h67ef)
	) name12984 (
		_w8905_,
		_w8908_,
		_w14883_,
		_w14884_,
		_w14885_
	);
	LUT3 #(
		.INIT('h80)
	) name12985 (
		\m6_addr_i[11]_pad ,
		_w8910_,
		_w8911_,
		_w14886_
	);
	LUT3 #(
		.INIT('h2a)
	) name12986 (
		\m5_addr_i[11]_pad ,
		_w8910_,
		_w8911_,
		_w14887_
	);
	LUT4 #(
		.INIT('hcdef)
	) name12987 (
		_w8905_,
		_w8908_,
		_w14886_,
		_w14887_,
		_w14888_
	);
	LUT4 #(
		.INIT('h7fff)
	) name12988 (
		_w14879_,
		_w14882_,
		_w14885_,
		_w14888_,
		_w14889_
	);
	LUT3 #(
		.INIT('h2a)
	) name12989 (
		\m1_addr_i[12]_pad ,
		_w8910_,
		_w8911_,
		_w14890_
	);
	LUT3 #(
		.INIT('h80)
	) name12990 (
		\m2_addr_i[12]_pad ,
		_w8910_,
		_w8911_,
		_w14891_
	);
	LUT4 #(
		.INIT('h3b7f)
	) name12991 (
		_w8905_,
		_w8908_,
		_w14890_,
		_w14891_,
		_w14892_
	);
	LUT3 #(
		.INIT('h2a)
	) name12992 (
		\m3_addr_i[12]_pad ,
		_w8910_,
		_w8911_,
		_w14893_
	);
	LUT3 #(
		.INIT('h2a)
	) name12993 (
		\m7_addr_i[12]_pad ,
		_w8910_,
		_w8911_,
		_w14894_
	);
	LUT4 #(
		.INIT('haebf)
	) name12994 (
		_w8905_,
		_w8908_,
		_w14893_,
		_w14894_,
		_w14895_
	);
	LUT3 #(
		.INIT('h80)
	) name12995 (
		\m4_addr_i[12]_pad ,
		_w8910_,
		_w8911_,
		_w14896_
	);
	LUT3 #(
		.INIT('h80)
	) name12996 (
		\m0_addr_i[12]_pad ,
		_w8910_,
		_w8911_,
		_w14897_
	);
	LUT4 #(
		.INIT('h57df)
	) name12997 (
		_w8905_,
		_w8908_,
		_w14896_,
		_w14897_,
		_w14898_
	);
	LUT3 #(
		.INIT('h80)
	) name12998 (
		\m6_addr_i[12]_pad ,
		_w8910_,
		_w8911_,
		_w14899_
	);
	LUT3 #(
		.INIT('h2a)
	) name12999 (
		\m5_addr_i[12]_pad ,
		_w8910_,
		_w8911_,
		_w14900_
	);
	LUT4 #(
		.INIT('hcdef)
	) name13000 (
		_w8905_,
		_w8908_,
		_w14899_,
		_w14900_,
		_w14901_
	);
	LUT4 #(
		.INIT('h7fff)
	) name13001 (
		_w14892_,
		_w14895_,
		_w14898_,
		_w14901_,
		_w14902_
	);
	LUT3 #(
		.INIT('h2a)
	) name13002 (
		\m3_addr_i[13]_pad ,
		_w8910_,
		_w8911_,
		_w14903_
	);
	LUT3 #(
		.INIT('h80)
	) name13003 (
		\m4_addr_i[13]_pad ,
		_w8910_,
		_w8911_,
		_w14904_
	);
	LUT4 #(
		.INIT('h9dbf)
	) name13004 (
		_w8905_,
		_w8908_,
		_w14903_,
		_w14904_,
		_w14905_
	);
	LUT3 #(
		.INIT('h80)
	) name13005 (
		\m0_addr_i[13]_pad ,
		_w8910_,
		_w8911_,
		_w14906_
	);
	LUT3 #(
		.INIT('h2a)
	) name13006 (
		\m5_addr_i[13]_pad ,
		_w8910_,
		_w8911_,
		_w14907_
	);
	LUT4 #(
		.INIT('h5d7f)
	) name13007 (
		_w8905_,
		_w8908_,
		_w14906_,
		_w14907_,
		_w14908_
	);
	LUT3 #(
		.INIT('h2a)
	) name13008 (
		\m7_addr_i[13]_pad ,
		_w8910_,
		_w8911_,
		_w14909_
	);
	LUT3 #(
		.INIT('h80)
	) name13009 (
		\m6_addr_i[13]_pad ,
		_w8910_,
		_w8911_,
		_w14910_
	);
	LUT3 #(
		.INIT('h57)
	) name13010 (
		_w8917_,
		_w14909_,
		_w14910_,
		_w14911_
	);
	LUT3 #(
		.INIT('h2a)
	) name13011 (
		\m1_addr_i[13]_pad ,
		_w8910_,
		_w8911_,
		_w14912_
	);
	LUT3 #(
		.INIT('h80)
	) name13012 (
		\m2_addr_i[13]_pad ,
		_w8910_,
		_w8911_,
		_w14913_
	);
	LUT4 #(
		.INIT('h3b7f)
	) name13013 (
		_w8905_,
		_w8908_,
		_w14912_,
		_w14913_,
		_w14914_
	);
	LUT4 #(
		.INIT('h7fff)
	) name13014 (
		_w14905_,
		_w14908_,
		_w14911_,
		_w14914_,
		_w14915_
	);
	LUT3 #(
		.INIT('h2a)
	) name13015 (
		\m3_addr_i[14]_pad ,
		_w8910_,
		_w8911_,
		_w14916_
	);
	LUT3 #(
		.INIT('h80)
	) name13016 (
		\m4_addr_i[14]_pad ,
		_w8910_,
		_w8911_,
		_w14917_
	);
	LUT4 #(
		.INIT('h9dbf)
	) name13017 (
		_w8905_,
		_w8908_,
		_w14916_,
		_w14917_,
		_w14918_
	);
	LUT3 #(
		.INIT('h2a)
	) name13018 (
		\m1_addr_i[14]_pad ,
		_w8910_,
		_w8911_,
		_w14919_
	);
	LUT3 #(
		.INIT('h2a)
	) name13019 (
		\m5_addr_i[14]_pad ,
		_w8910_,
		_w8911_,
		_w14920_
	);
	LUT4 #(
		.INIT('h5d7f)
	) name13020 (
		_w8905_,
		_w8908_,
		_w14919_,
		_w14920_,
		_w14921_
	);
	LUT3 #(
		.INIT('h80)
	) name13021 (
		\m2_addr_i[14]_pad ,
		_w8910_,
		_w8911_,
		_w14922_
	);
	LUT3 #(
		.INIT('h80)
	) name13022 (
		\m6_addr_i[14]_pad ,
		_w8910_,
		_w8911_,
		_w14923_
	);
	LUT4 #(
		.INIT('haebf)
	) name13023 (
		_w8905_,
		_w8908_,
		_w14922_,
		_w14923_,
		_w14924_
	);
	LUT3 #(
		.INIT('h80)
	) name13024 (
		\m0_addr_i[14]_pad ,
		_w8910_,
		_w8911_,
		_w14925_
	);
	LUT3 #(
		.INIT('h2a)
	) name13025 (
		\m7_addr_i[14]_pad ,
		_w8910_,
		_w8911_,
		_w14926_
	);
	LUT4 #(
		.INIT('h6e7f)
	) name13026 (
		_w8905_,
		_w8908_,
		_w14925_,
		_w14926_,
		_w14927_
	);
	LUT4 #(
		.INIT('h7fff)
	) name13027 (
		_w14918_,
		_w14921_,
		_w14924_,
		_w14927_,
		_w14928_
	);
	LUT3 #(
		.INIT('h2a)
	) name13028 (
		\m1_addr_i[15]_pad ,
		_w8910_,
		_w8911_,
		_w14929_
	);
	LUT3 #(
		.INIT('h80)
	) name13029 (
		\m2_addr_i[15]_pad ,
		_w8910_,
		_w8911_,
		_w14930_
	);
	LUT4 #(
		.INIT('h3b7f)
	) name13030 (
		_w8905_,
		_w8908_,
		_w14929_,
		_w14930_,
		_w14931_
	);
	LUT3 #(
		.INIT('h80)
	) name13031 (
		\m0_addr_i[15]_pad ,
		_w8910_,
		_w8911_,
		_w14932_
	);
	LUT3 #(
		.INIT('h80)
	) name13032 (
		\m4_addr_i[15]_pad ,
		_w8910_,
		_w8911_,
		_w14933_
	);
	LUT4 #(
		.INIT('h5d7f)
	) name13033 (
		_w8905_,
		_w8908_,
		_w14932_,
		_w14933_,
		_w14934_
	);
	LUT3 #(
		.INIT('h2a)
	) name13034 (
		\m7_addr_i[15]_pad ,
		_w8910_,
		_w8911_,
		_w14935_
	);
	LUT3 #(
		.INIT('h2a)
	) name13035 (
		\m3_addr_i[15]_pad ,
		_w8910_,
		_w8911_,
		_w14936_
	);
	LUT4 #(
		.INIT('habef)
	) name13036 (
		_w8905_,
		_w8908_,
		_w14935_,
		_w14936_,
		_w14937_
	);
	LUT3 #(
		.INIT('h80)
	) name13037 (
		\m6_addr_i[15]_pad ,
		_w8910_,
		_w8911_,
		_w14938_
	);
	LUT3 #(
		.INIT('h2a)
	) name13038 (
		\m5_addr_i[15]_pad ,
		_w8910_,
		_w8911_,
		_w14939_
	);
	LUT4 #(
		.INIT('hcdef)
	) name13039 (
		_w8905_,
		_w8908_,
		_w14938_,
		_w14939_,
		_w14940_
	);
	LUT4 #(
		.INIT('h7fff)
	) name13040 (
		_w14931_,
		_w14934_,
		_w14937_,
		_w14940_,
		_w14941_
	);
	LUT3 #(
		.INIT('h80)
	) name13041 (
		\m6_addr_i[16]_pad ,
		_w8910_,
		_w8911_,
		_w14942_
	);
	LUT3 #(
		.INIT('h2a)
	) name13042 (
		\m5_addr_i[16]_pad ,
		_w8910_,
		_w8911_,
		_w14943_
	);
	LUT4 #(
		.INIT('hcdef)
	) name13043 (
		_w8905_,
		_w8908_,
		_w14942_,
		_w14943_,
		_w14944_
	);
	LUT3 #(
		.INIT('h80)
	) name13044 (
		\m0_addr_i[16]_pad ,
		_w8910_,
		_w8911_,
		_w14945_
	);
	LUT3 #(
		.INIT('h80)
	) name13045 (
		\m4_addr_i[16]_pad ,
		_w8910_,
		_w8911_,
		_w14946_
	);
	LUT4 #(
		.INIT('h5d7f)
	) name13046 (
		_w8905_,
		_w8908_,
		_w14945_,
		_w14946_,
		_w14947_
	);
	LUT3 #(
		.INIT('h2a)
	) name13047 (
		\m7_addr_i[16]_pad ,
		_w8910_,
		_w8911_,
		_w14948_
	);
	LUT3 #(
		.INIT('h2a)
	) name13048 (
		\m3_addr_i[16]_pad ,
		_w8910_,
		_w8911_,
		_w14949_
	);
	LUT4 #(
		.INIT('habef)
	) name13049 (
		_w8905_,
		_w8908_,
		_w14948_,
		_w14949_,
		_w14950_
	);
	LUT3 #(
		.INIT('h2a)
	) name13050 (
		\m1_addr_i[16]_pad ,
		_w8910_,
		_w8911_,
		_w14951_
	);
	LUT3 #(
		.INIT('h80)
	) name13051 (
		\m2_addr_i[16]_pad ,
		_w8910_,
		_w8911_,
		_w14952_
	);
	LUT4 #(
		.INIT('h3b7f)
	) name13052 (
		_w8905_,
		_w8908_,
		_w14951_,
		_w14952_,
		_w14953_
	);
	LUT4 #(
		.INIT('h7fff)
	) name13053 (
		_w14944_,
		_w14947_,
		_w14950_,
		_w14953_,
		_w14954_
	);
	LUT3 #(
		.INIT('h80)
	) name13054 (
		\m0_addr_i[17]_pad ,
		_w8910_,
		_w8911_,
		_w14955_
	);
	LUT3 #(
		.INIT('h2a)
	) name13055 (
		\m7_addr_i[17]_pad ,
		_w8910_,
		_w8911_,
		_w14956_
	);
	LUT4 #(
		.INIT('h6e7f)
	) name13056 (
		_w8905_,
		_w8908_,
		_w14955_,
		_w14956_,
		_w14957_
	);
	LUT3 #(
		.INIT('h2a)
	) name13057 (
		\m1_addr_i[17]_pad ,
		_w8910_,
		_w8911_,
		_w14958_
	);
	LUT3 #(
		.INIT('h80)
	) name13058 (
		\m4_addr_i[17]_pad ,
		_w8910_,
		_w8911_,
		_w14959_
	);
	LUT4 #(
		.INIT('h5d7f)
	) name13059 (
		_w8905_,
		_w8908_,
		_w14958_,
		_w14959_,
		_w14960_
	);
	LUT3 #(
		.INIT('h80)
	) name13060 (
		\m2_addr_i[17]_pad ,
		_w8910_,
		_w8911_,
		_w14961_
	);
	LUT3 #(
		.INIT('h2a)
	) name13061 (
		\m3_addr_i[17]_pad ,
		_w8910_,
		_w8911_,
		_w14962_
	);
	LUT3 #(
		.INIT('h57)
	) name13062 (
		_w8909_,
		_w14961_,
		_w14962_,
		_w14963_
	);
	LUT3 #(
		.INIT('h80)
	) name13063 (
		\m6_addr_i[17]_pad ,
		_w8910_,
		_w8911_,
		_w14964_
	);
	LUT3 #(
		.INIT('h2a)
	) name13064 (
		\m5_addr_i[17]_pad ,
		_w8910_,
		_w8911_,
		_w14965_
	);
	LUT4 #(
		.INIT('hcdef)
	) name13065 (
		_w8905_,
		_w8908_,
		_w14964_,
		_w14965_,
		_w14966_
	);
	LUT4 #(
		.INIT('h7fff)
	) name13066 (
		_w14957_,
		_w14960_,
		_w14963_,
		_w14966_,
		_w14967_
	);
	LUT3 #(
		.INIT('h2a)
	) name13067 (
		\m3_addr_i[18]_pad ,
		_w8910_,
		_w8911_,
		_w14968_
	);
	LUT3 #(
		.INIT('h80)
	) name13068 (
		\m4_addr_i[18]_pad ,
		_w8910_,
		_w8911_,
		_w14969_
	);
	LUT4 #(
		.INIT('h9dbf)
	) name13069 (
		_w8905_,
		_w8908_,
		_w14968_,
		_w14969_,
		_w14970_
	);
	LUT3 #(
		.INIT('h2a)
	) name13070 (
		\m1_addr_i[18]_pad ,
		_w8910_,
		_w8911_,
		_w14971_
	);
	LUT3 #(
		.INIT('h2a)
	) name13071 (
		\m5_addr_i[18]_pad ,
		_w8910_,
		_w8911_,
		_w14972_
	);
	LUT4 #(
		.INIT('h5d7f)
	) name13072 (
		_w8905_,
		_w8908_,
		_w14971_,
		_w14972_,
		_w14973_
	);
	LUT3 #(
		.INIT('h80)
	) name13073 (
		\m2_addr_i[18]_pad ,
		_w8910_,
		_w8911_,
		_w14974_
	);
	LUT3 #(
		.INIT('h80)
	) name13074 (
		\m6_addr_i[18]_pad ,
		_w8910_,
		_w8911_,
		_w14975_
	);
	LUT4 #(
		.INIT('haebf)
	) name13075 (
		_w8905_,
		_w8908_,
		_w14974_,
		_w14975_,
		_w14976_
	);
	LUT3 #(
		.INIT('h80)
	) name13076 (
		\m0_addr_i[18]_pad ,
		_w8910_,
		_w8911_,
		_w14977_
	);
	LUT3 #(
		.INIT('h2a)
	) name13077 (
		\m7_addr_i[18]_pad ,
		_w8910_,
		_w8911_,
		_w14978_
	);
	LUT4 #(
		.INIT('h6e7f)
	) name13078 (
		_w8905_,
		_w8908_,
		_w14977_,
		_w14978_,
		_w14979_
	);
	LUT4 #(
		.INIT('h7fff)
	) name13079 (
		_w14970_,
		_w14973_,
		_w14976_,
		_w14979_,
		_w14980_
	);
	LUT3 #(
		.INIT('h80)
	) name13080 (
		\m6_addr_i[19]_pad ,
		_w8910_,
		_w8911_,
		_w14981_
	);
	LUT3 #(
		.INIT('h2a)
	) name13081 (
		\m5_addr_i[19]_pad ,
		_w8910_,
		_w8911_,
		_w14982_
	);
	LUT4 #(
		.INIT('hcdef)
	) name13082 (
		_w8905_,
		_w8908_,
		_w14981_,
		_w14982_,
		_w14983_
	);
	LUT3 #(
		.INIT('h80)
	) name13083 (
		\m0_addr_i[19]_pad ,
		_w8910_,
		_w8911_,
		_w14984_
	);
	LUT3 #(
		.INIT('h80)
	) name13084 (
		\m4_addr_i[19]_pad ,
		_w8910_,
		_w8911_,
		_w14985_
	);
	LUT4 #(
		.INIT('h5d7f)
	) name13085 (
		_w8905_,
		_w8908_,
		_w14984_,
		_w14985_,
		_w14986_
	);
	LUT3 #(
		.INIT('h2a)
	) name13086 (
		\m7_addr_i[19]_pad ,
		_w8910_,
		_w8911_,
		_w14987_
	);
	LUT3 #(
		.INIT('h2a)
	) name13087 (
		\m3_addr_i[19]_pad ,
		_w8910_,
		_w8911_,
		_w14988_
	);
	LUT4 #(
		.INIT('habef)
	) name13088 (
		_w8905_,
		_w8908_,
		_w14987_,
		_w14988_,
		_w14989_
	);
	LUT3 #(
		.INIT('h2a)
	) name13089 (
		\m1_addr_i[19]_pad ,
		_w8910_,
		_w8911_,
		_w14990_
	);
	LUT3 #(
		.INIT('h80)
	) name13090 (
		\m2_addr_i[19]_pad ,
		_w8910_,
		_w8911_,
		_w14991_
	);
	LUT4 #(
		.INIT('h3b7f)
	) name13091 (
		_w8905_,
		_w8908_,
		_w14990_,
		_w14991_,
		_w14992_
	);
	LUT4 #(
		.INIT('h7fff)
	) name13092 (
		_w14983_,
		_w14986_,
		_w14989_,
		_w14992_,
		_w14993_
	);
	LUT3 #(
		.INIT('h80)
	) name13093 (
		\m0_addr_i[1]_pad ,
		_w8910_,
		_w8911_,
		_w14994_
	);
	LUT3 #(
		.INIT('h2a)
	) name13094 (
		\m7_addr_i[1]_pad ,
		_w8910_,
		_w8911_,
		_w14995_
	);
	LUT4 #(
		.INIT('h6e7f)
	) name13095 (
		_w8905_,
		_w8908_,
		_w14994_,
		_w14995_,
		_w14996_
	);
	LUT3 #(
		.INIT('h80)
	) name13096 (
		\m6_addr_i[1]_pad ,
		_w8910_,
		_w8911_,
		_w14997_
	);
	LUT3 #(
		.INIT('h80)
	) name13097 (
		\m2_addr_i[1]_pad ,
		_w8910_,
		_w8911_,
		_w14998_
	);
	LUT4 #(
		.INIT('habef)
	) name13098 (
		_w8905_,
		_w8908_,
		_w14997_,
		_w14998_,
		_w14999_
	);
	LUT3 #(
		.INIT('h2a)
	) name13099 (
		\m5_addr_i[1]_pad ,
		_w8910_,
		_w8911_,
		_w15000_
	);
	LUT3 #(
		.INIT('h2a)
	) name13100 (
		\m1_addr_i[1]_pad ,
		_w8910_,
		_w8911_,
		_w15001_
	);
	LUT4 #(
		.INIT('h57df)
	) name13101 (
		_w8905_,
		_w8908_,
		_w15000_,
		_w15001_,
		_w15002_
	);
	LUT3 #(
		.INIT('h2a)
	) name13102 (
		\m3_addr_i[1]_pad ,
		_w8910_,
		_w8911_,
		_w15003_
	);
	LUT3 #(
		.INIT('h80)
	) name13103 (
		\m4_addr_i[1]_pad ,
		_w8910_,
		_w8911_,
		_w15004_
	);
	LUT4 #(
		.INIT('h9dbf)
	) name13104 (
		_w8905_,
		_w8908_,
		_w15003_,
		_w15004_,
		_w15005_
	);
	LUT4 #(
		.INIT('h7fff)
	) name13105 (
		_w14996_,
		_w14999_,
		_w15002_,
		_w15005_,
		_w15006_
	);
	LUT3 #(
		.INIT('h2a)
	) name13106 (
		\m1_addr_i[20]_pad ,
		_w8910_,
		_w8911_,
		_w15007_
	);
	LUT3 #(
		.INIT('h80)
	) name13107 (
		\m2_addr_i[20]_pad ,
		_w8910_,
		_w8911_,
		_w15008_
	);
	LUT4 #(
		.INIT('h3b7f)
	) name13108 (
		_w8905_,
		_w8908_,
		_w15007_,
		_w15008_,
		_w15009_
	);
	LUT3 #(
		.INIT('h80)
	) name13109 (
		\m0_addr_i[20]_pad ,
		_w8910_,
		_w8911_,
		_w15010_
	);
	LUT3 #(
		.INIT('h80)
	) name13110 (
		\m4_addr_i[20]_pad ,
		_w8910_,
		_w8911_,
		_w15011_
	);
	LUT4 #(
		.INIT('h5d7f)
	) name13111 (
		_w8905_,
		_w8908_,
		_w15010_,
		_w15011_,
		_w15012_
	);
	LUT3 #(
		.INIT('h2a)
	) name13112 (
		\m7_addr_i[20]_pad ,
		_w8910_,
		_w8911_,
		_w15013_
	);
	LUT3 #(
		.INIT('h2a)
	) name13113 (
		\m3_addr_i[20]_pad ,
		_w8910_,
		_w8911_,
		_w15014_
	);
	LUT4 #(
		.INIT('habef)
	) name13114 (
		_w8905_,
		_w8908_,
		_w15013_,
		_w15014_,
		_w15015_
	);
	LUT3 #(
		.INIT('h80)
	) name13115 (
		\m6_addr_i[20]_pad ,
		_w8910_,
		_w8911_,
		_w15016_
	);
	LUT3 #(
		.INIT('h2a)
	) name13116 (
		\m5_addr_i[20]_pad ,
		_w8910_,
		_w8911_,
		_w15017_
	);
	LUT4 #(
		.INIT('hcdef)
	) name13117 (
		_w8905_,
		_w8908_,
		_w15016_,
		_w15017_,
		_w15018_
	);
	LUT4 #(
		.INIT('h7fff)
	) name13118 (
		_w15009_,
		_w15012_,
		_w15015_,
		_w15018_,
		_w15019_
	);
	LUT3 #(
		.INIT('h2a)
	) name13119 (
		\m3_addr_i[21]_pad ,
		_w8910_,
		_w8911_,
		_w15020_
	);
	LUT3 #(
		.INIT('h80)
	) name13120 (
		\m4_addr_i[21]_pad ,
		_w8910_,
		_w8911_,
		_w15021_
	);
	LUT4 #(
		.INIT('h9dbf)
	) name13121 (
		_w8905_,
		_w8908_,
		_w15020_,
		_w15021_,
		_w15022_
	);
	LUT3 #(
		.INIT('h2a)
	) name13122 (
		\m1_addr_i[21]_pad ,
		_w8910_,
		_w8911_,
		_w15023_
	);
	LUT3 #(
		.INIT('h2a)
	) name13123 (
		\m7_addr_i[21]_pad ,
		_w8910_,
		_w8911_,
		_w15024_
	);
	LUT4 #(
		.INIT('h6e7f)
	) name13124 (
		_w8905_,
		_w8908_,
		_w15023_,
		_w15024_,
		_w15025_
	);
	LUT3 #(
		.INIT('h80)
	) name13125 (
		\m2_addr_i[21]_pad ,
		_w8910_,
		_w8911_,
		_w15026_
	);
	LUT3 #(
		.INIT('h80)
	) name13126 (
		\m0_addr_i[21]_pad ,
		_w8910_,
		_w8911_,
		_w15027_
	);
	LUT4 #(
		.INIT('h37bf)
	) name13127 (
		_w8905_,
		_w8908_,
		_w15026_,
		_w15027_,
		_w15028_
	);
	LUT3 #(
		.INIT('h80)
	) name13128 (
		\m6_addr_i[21]_pad ,
		_w8910_,
		_w8911_,
		_w15029_
	);
	LUT3 #(
		.INIT('h2a)
	) name13129 (
		\m5_addr_i[21]_pad ,
		_w8910_,
		_w8911_,
		_w15030_
	);
	LUT4 #(
		.INIT('hcdef)
	) name13130 (
		_w8905_,
		_w8908_,
		_w15029_,
		_w15030_,
		_w15031_
	);
	LUT4 #(
		.INIT('h7fff)
	) name13131 (
		_w15022_,
		_w15025_,
		_w15028_,
		_w15031_,
		_w15032_
	);
	LUT3 #(
		.INIT('h2a)
	) name13132 (
		\m1_addr_i[22]_pad ,
		_w8910_,
		_w8911_,
		_w15033_
	);
	LUT3 #(
		.INIT('h80)
	) name13133 (
		\m2_addr_i[22]_pad ,
		_w8910_,
		_w8911_,
		_w15034_
	);
	LUT4 #(
		.INIT('h3b7f)
	) name13134 (
		_w8905_,
		_w8908_,
		_w15033_,
		_w15034_,
		_w15035_
	);
	LUT3 #(
		.INIT('h80)
	) name13135 (
		\m0_addr_i[22]_pad ,
		_w8910_,
		_w8911_,
		_w15036_
	);
	LUT3 #(
		.INIT('h80)
	) name13136 (
		\m4_addr_i[22]_pad ,
		_w8910_,
		_w8911_,
		_w15037_
	);
	LUT4 #(
		.INIT('h5d7f)
	) name13137 (
		_w8905_,
		_w8908_,
		_w15036_,
		_w15037_,
		_w15038_
	);
	LUT3 #(
		.INIT('h2a)
	) name13138 (
		\m7_addr_i[22]_pad ,
		_w8910_,
		_w8911_,
		_w15039_
	);
	LUT3 #(
		.INIT('h2a)
	) name13139 (
		\m3_addr_i[22]_pad ,
		_w8910_,
		_w8911_,
		_w15040_
	);
	LUT4 #(
		.INIT('habef)
	) name13140 (
		_w8905_,
		_w8908_,
		_w15039_,
		_w15040_,
		_w15041_
	);
	LUT3 #(
		.INIT('h80)
	) name13141 (
		\m6_addr_i[22]_pad ,
		_w8910_,
		_w8911_,
		_w15042_
	);
	LUT3 #(
		.INIT('h2a)
	) name13142 (
		\m5_addr_i[22]_pad ,
		_w8910_,
		_w8911_,
		_w15043_
	);
	LUT4 #(
		.INIT('hcdef)
	) name13143 (
		_w8905_,
		_w8908_,
		_w15042_,
		_w15043_,
		_w15044_
	);
	LUT4 #(
		.INIT('h7fff)
	) name13144 (
		_w15035_,
		_w15038_,
		_w15041_,
		_w15044_,
		_w15045_
	);
	LUT3 #(
		.INIT('h2a)
	) name13145 (
		\m1_addr_i[23]_pad ,
		_w8910_,
		_w8911_,
		_w15046_
	);
	LUT3 #(
		.INIT('h80)
	) name13146 (
		\m2_addr_i[23]_pad ,
		_w8910_,
		_w8911_,
		_w15047_
	);
	LUT4 #(
		.INIT('h3b7f)
	) name13147 (
		_w8905_,
		_w8908_,
		_w15046_,
		_w15047_,
		_w15048_
	);
	LUT3 #(
		.INIT('h80)
	) name13148 (
		\m0_addr_i[23]_pad ,
		_w8910_,
		_w8911_,
		_w15049_
	);
	LUT3 #(
		.INIT('h80)
	) name13149 (
		\m4_addr_i[23]_pad ,
		_w8910_,
		_w8911_,
		_w15050_
	);
	LUT4 #(
		.INIT('h5d7f)
	) name13150 (
		_w8905_,
		_w8908_,
		_w15049_,
		_w15050_,
		_w15051_
	);
	LUT3 #(
		.INIT('h2a)
	) name13151 (
		\m7_addr_i[23]_pad ,
		_w8910_,
		_w8911_,
		_w15052_
	);
	LUT3 #(
		.INIT('h2a)
	) name13152 (
		\m3_addr_i[23]_pad ,
		_w8910_,
		_w8911_,
		_w15053_
	);
	LUT4 #(
		.INIT('habef)
	) name13153 (
		_w8905_,
		_w8908_,
		_w15052_,
		_w15053_,
		_w15054_
	);
	LUT3 #(
		.INIT('h80)
	) name13154 (
		\m6_addr_i[23]_pad ,
		_w8910_,
		_w8911_,
		_w15055_
	);
	LUT3 #(
		.INIT('h2a)
	) name13155 (
		\m5_addr_i[23]_pad ,
		_w8910_,
		_w8911_,
		_w15056_
	);
	LUT4 #(
		.INIT('hcdef)
	) name13156 (
		_w8905_,
		_w8908_,
		_w15055_,
		_w15056_,
		_w15057_
	);
	LUT4 #(
		.INIT('h7fff)
	) name13157 (
		_w15048_,
		_w15051_,
		_w15054_,
		_w15057_,
		_w15058_
	);
	LUT3 #(
		.INIT('h2a)
	) name13158 (
		\m3_addr_i[24]_pad ,
		_w8910_,
		_w8911_,
		_w15059_
	);
	LUT3 #(
		.INIT('h80)
	) name13159 (
		\m4_addr_i[24]_pad ,
		_w8910_,
		_w8911_,
		_w15060_
	);
	LUT4 #(
		.INIT('h9dbf)
	) name13160 (
		_w8905_,
		_w8908_,
		_w15059_,
		_w15060_,
		_w15061_
	);
	LUT3 #(
		.INIT('h2a)
	) name13161 (
		\m5_addr_i[24]_pad ,
		_w8910_,
		_w8911_,
		_w15062_
	);
	LUT3 #(
		.INIT('h2a)
	) name13162 (
		\m7_addr_i[24]_pad ,
		_w8910_,
		_w8911_,
		_w15063_
	);
	LUT4 #(
		.INIT('hcedf)
	) name13163 (
		_w8905_,
		_w8908_,
		_w15062_,
		_w15063_,
		_w15064_
	);
	LUT3 #(
		.INIT('h80)
	) name13164 (
		\m6_addr_i[24]_pad ,
		_w8910_,
		_w8911_,
		_w15065_
	);
	LUT3 #(
		.INIT('h80)
	) name13165 (
		\m0_addr_i[24]_pad ,
		_w8910_,
		_w8911_,
		_w15066_
	);
	LUT4 #(
		.INIT('h67ef)
	) name13166 (
		_w8905_,
		_w8908_,
		_w15065_,
		_w15066_,
		_w15067_
	);
	LUT3 #(
		.INIT('h2a)
	) name13167 (
		\m1_addr_i[24]_pad ,
		_w8910_,
		_w8911_,
		_w15068_
	);
	LUT3 #(
		.INIT('h80)
	) name13168 (
		\m2_addr_i[24]_pad ,
		_w8910_,
		_w8911_,
		_w15069_
	);
	LUT4 #(
		.INIT('h3b7f)
	) name13169 (
		_w8905_,
		_w8908_,
		_w15068_,
		_w15069_,
		_w15070_
	);
	LUT4 #(
		.INIT('h7fff)
	) name13170 (
		_w15061_,
		_w15064_,
		_w15067_,
		_w15070_,
		_w15071_
	);
	LUT3 #(
		.INIT('h80)
	) name13171 (
		\m0_addr_i[25]_pad ,
		_w8910_,
		_w8911_,
		_w15072_
	);
	LUT3 #(
		.INIT('h2a)
	) name13172 (
		\m7_addr_i[25]_pad ,
		_w8910_,
		_w8911_,
		_w15073_
	);
	LUT4 #(
		.INIT('h6e7f)
	) name13173 (
		_w8905_,
		_w8908_,
		_w15072_,
		_w15073_,
		_w15074_
	);
	LUT3 #(
		.INIT('h2a)
	) name13174 (
		\m1_addr_i[25]_pad ,
		_w8910_,
		_w8911_,
		_w15075_
	);
	LUT3 #(
		.INIT('h80)
	) name13175 (
		\m4_addr_i[25]_pad ,
		_w8910_,
		_w8911_,
		_w15076_
	);
	LUT4 #(
		.INIT('h5d7f)
	) name13176 (
		_w8905_,
		_w8908_,
		_w15075_,
		_w15076_,
		_w15077_
	);
	LUT3 #(
		.INIT('h80)
	) name13177 (
		\m2_addr_i[25]_pad ,
		_w8910_,
		_w8911_,
		_w15078_
	);
	LUT3 #(
		.INIT('h2a)
	) name13178 (
		\m3_addr_i[25]_pad ,
		_w8910_,
		_w8911_,
		_w15079_
	);
	LUT3 #(
		.INIT('h57)
	) name13179 (
		_w8909_,
		_w15078_,
		_w15079_,
		_w15080_
	);
	LUT3 #(
		.INIT('h2a)
	) name13180 (
		\m5_addr_i[25]_pad ,
		_w8910_,
		_w8911_,
		_w15081_
	);
	LUT3 #(
		.INIT('h80)
	) name13181 (
		\m6_addr_i[25]_pad ,
		_w8910_,
		_w8911_,
		_w15082_
	);
	LUT4 #(
		.INIT('hcedf)
	) name13182 (
		_w8905_,
		_w8908_,
		_w15081_,
		_w15082_,
		_w15083_
	);
	LUT4 #(
		.INIT('h7fff)
	) name13183 (
		_w15074_,
		_w15077_,
		_w15080_,
		_w15083_,
		_w15084_
	);
	LUT3 #(
		.INIT('h80)
	) name13184 (
		\m0_addr_i[26]_pad ,
		_w8910_,
		_w8911_,
		_w15085_
	);
	LUT3 #(
		.INIT('h2a)
	) name13185 (
		\m7_addr_i[26]_pad ,
		_w8910_,
		_w8911_,
		_w15086_
	);
	LUT4 #(
		.INIT('h6e7f)
	) name13186 (
		_w8905_,
		_w8908_,
		_w15085_,
		_w15086_,
		_w15087_
	);
	LUT3 #(
		.INIT('h2a)
	) name13187 (
		\m5_addr_i[26]_pad ,
		_w8910_,
		_w8911_,
		_w15088_
	);
	LUT3 #(
		.INIT('h80)
	) name13188 (
		\m2_addr_i[26]_pad ,
		_w8910_,
		_w8911_,
		_w15089_
	);
	LUT4 #(
		.INIT('h9bdf)
	) name13189 (
		_w8905_,
		_w8908_,
		_w15088_,
		_w15089_,
		_w15090_
	);
	LUT3 #(
		.INIT('h80)
	) name13190 (
		\m6_addr_i[26]_pad ,
		_w8910_,
		_w8911_,
		_w15091_
	);
	LUT3 #(
		.INIT('h2a)
	) name13191 (
		\m1_addr_i[26]_pad ,
		_w8910_,
		_w8911_,
		_w15092_
	);
	LUT4 #(
		.INIT('h67ef)
	) name13192 (
		_w8905_,
		_w8908_,
		_w15091_,
		_w15092_,
		_w15093_
	);
	LUT3 #(
		.INIT('h2a)
	) name13193 (
		\m3_addr_i[26]_pad ,
		_w8910_,
		_w8911_,
		_w15094_
	);
	LUT3 #(
		.INIT('h80)
	) name13194 (
		\m4_addr_i[26]_pad ,
		_w8910_,
		_w8911_,
		_w15095_
	);
	LUT4 #(
		.INIT('h9dbf)
	) name13195 (
		_w8905_,
		_w8908_,
		_w15094_,
		_w15095_,
		_w15096_
	);
	LUT4 #(
		.INIT('h7fff)
	) name13196 (
		_w15087_,
		_w15090_,
		_w15093_,
		_w15096_,
		_w15097_
	);
	LUT3 #(
		.INIT('h80)
	) name13197 (
		\m0_addr_i[27]_pad ,
		_w8910_,
		_w8911_,
		_w15098_
	);
	LUT3 #(
		.INIT('h2a)
	) name13198 (
		\m7_addr_i[27]_pad ,
		_w8910_,
		_w8911_,
		_w15099_
	);
	LUT4 #(
		.INIT('h6e7f)
	) name13199 (
		_w8905_,
		_w8908_,
		_w15098_,
		_w15099_,
		_w15100_
	);
	LUT3 #(
		.INIT('h2a)
	) name13200 (
		\m1_addr_i[27]_pad ,
		_w8910_,
		_w8911_,
		_w15101_
	);
	LUT3 #(
		.INIT('h80)
	) name13201 (
		\m4_addr_i[27]_pad ,
		_w8910_,
		_w8911_,
		_w15102_
	);
	LUT4 #(
		.INIT('h5d7f)
	) name13202 (
		_w8905_,
		_w8908_,
		_w15101_,
		_w15102_,
		_w15103_
	);
	LUT3 #(
		.INIT('h80)
	) name13203 (
		\m2_addr_i[27]_pad ,
		_w8910_,
		_w8911_,
		_w15104_
	);
	LUT3 #(
		.INIT('h2a)
	) name13204 (
		\m3_addr_i[27]_pad ,
		_w8910_,
		_w8911_,
		_w15105_
	);
	LUT3 #(
		.INIT('h57)
	) name13205 (
		_w8909_,
		_w15104_,
		_w15105_,
		_w15106_
	);
	LUT3 #(
		.INIT('h2a)
	) name13206 (
		\m5_addr_i[27]_pad ,
		_w8910_,
		_w8911_,
		_w15107_
	);
	LUT3 #(
		.INIT('h80)
	) name13207 (
		\m6_addr_i[27]_pad ,
		_w8910_,
		_w8911_,
		_w15108_
	);
	LUT4 #(
		.INIT('hcedf)
	) name13208 (
		_w8905_,
		_w8908_,
		_w15107_,
		_w15108_,
		_w15109_
	);
	LUT4 #(
		.INIT('h7fff)
	) name13209 (
		_w15100_,
		_w15103_,
		_w15106_,
		_w15109_,
		_w15110_
	);
	LUT3 #(
		.INIT('h2a)
	) name13210 (
		\m3_addr_i[28]_pad ,
		_w8910_,
		_w8911_,
		_w15111_
	);
	LUT3 #(
		.INIT('h80)
	) name13211 (
		\m4_addr_i[28]_pad ,
		_w8910_,
		_w8911_,
		_w15112_
	);
	LUT4 #(
		.INIT('h9dbf)
	) name13212 (
		_w8905_,
		_w8908_,
		_w15111_,
		_w15112_,
		_w15113_
	);
	LUT3 #(
		.INIT('h2a)
	) name13213 (
		\m5_addr_i[28]_pad ,
		_w8910_,
		_w8911_,
		_w15114_
	);
	LUT3 #(
		.INIT('h2a)
	) name13214 (
		\m7_addr_i[28]_pad ,
		_w8910_,
		_w8911_,
		_w15115_
	);
	LUT4 #(
		.INIT('hcedf)
	) name13215 (
		_w8905_,
		_w8908_,
		_w15114_,
		_w15115_,
		_w15116_
	);
	LUT3 #(
		.INIT('h80)
	) name13216 (
		\m6_addr_i[28]_pad ,
		_w8910_,
		_w8911_,
		_w15117_
	);
	LUT3 #(
		.INIT('h80)
	) name13217 (
		\m0_addr_i[28]_pad ,
		_w8910_,
		_w8911_,
		_w15118_
	);
	LUT4 #(
		.INIT('h67ef)
	) name13218 (
		_w8905_,
		_w8908_,
		_w15117_,
		_w15118_,
		_w15119_
	);
	LUT3 #(
		.INIT('h2a)
	) name13219 (
		\m1_addr_i[28]_pad ,
		_w8910_,
		_w8911_,
		_w15120_
	);
	LUT3 #(
		.INIT('h80)
	) name13220 (
		\m2_addr_i[28]_pad ,
		_w8910_,
		_w8911_,
		_w15121_
	);
	LUT4 #(
		.INIT('h3b7f)
	) name13221 (
		_w8905_,
		_w8908_,
		_w15120_,
		_w15121_,
		_w15122_
	);
	LUT4 #(
		.INIT('h7fff)
	) name13222 (
		_w15113_,
		_w15116_,
		_w15119_,
		_w15122_,
		_w15123_
	);
	LUT3 #(
		.INIT('h80)
	) name13223 (
		\m0_addr_i[29]_pad ,
		_w8910_,
		_w8911_,
		_w15124_
	);
	LUT3 #(
		.INIT('h2a)
	) name13224 (
		\m7_addr_i[29]_pad ,
		_w8910_,
		_w8911_,
		_w15125_
	);
	LUT4 #(
		.INIT('h6e7f)
	) name13225 (
		_w8905_,
		_w8908_,
		_w15124_,
		_w15125_,
		_w15126_
	);
	LUT3 #(
		.INIT('h2a)
	) name13226 (
		\m1_addr_i[29]_pad ,
		_w8910_,
		_w8911_,
		_w15127_
	);
	LUT3 #(
		.INIT('h80)
	) name13227 (
		\m4_addr_i[29]_pad ,
		_w8910_,
		_w8911_,
		_w15128_
	);
	LUT4 #(
		.INIT('h5d7f)
	) name13228 (
		_w8905_,
		_w8908_,
		_w15127_,
		_w15128_,
		_w15129_
	);
	LUT3 #(
		.INIT('h80)
	) name13229 (
		\m2_addr_i[29]_pad ,
		_w8910_,
		_w8911_,
		_w15130_
	);
	LUT3 #(
		.INIT('h2a)
	) name13230 (
		\m3_addr_i[29]_pad ,
		_w8910_,
		_w8911_,
		_w15131_
	);
	LUT3 #(
		.INIT('h57)
	) name13231 (
		_w8909_,
		_w15130_,
		_w15131_,
		_w15132_
	);
	LUT3 #(
		.INIT('h2a)
	) name13232 (
		\m5_addr_i[29]_pad ,
		_w8910_,
		_w8911_,
		_w15133_
	);
	LUT3 #(
		.INIT('h80)
	) name13233 (
		\m6_addr_i[29]_pad ,
		_w8910_,
		_w8911_,
		_w15134_
	);
	LUT4 #(
		.INIT('hcedf)
	) name13234 (
		_w8905_,
		_w8908_,
		_w15133_,
		_w15134_,
		_w15135_
	);
	LUT4 #(
		.INIT('h7fff)
	) name13235 (
		_w15126_,
		_w15129_,
		_w15132_,
		_w15135_,
		_w15136_
	);
	LUT3 #(
		.INIT('h80)
	) name13236 (
		\m0_addr_i[2]_pad ,
		_w8910_,
		_w8911_,
		_w15137_
	);
	LUT3 #(
		.INIT('h2a)
	) name13237 (
		\m7_addr_i[2]_pad ,
		_w8910_,
		_w8911_,
		_w15138_
	);
	LUT4 #(
		.INIT('h6e7f)
	) name13238 (
		_w8905_,
		_w8908_,
		_w15137_,
		_w15138_,
		_w15139_
	);
	LUT3 #(
		.INIT('h80)
	) name13239 (
		\m6_addr_i[2]_pad ,
		_w8910_,
		_w8911_,
		_w15140_
	);
	LUT3 #(
		.INIT('h80)
	) name13240 (
		\m2_addr_i[2]_pad ,
		_w8910_,
		_w8911_,
		_w15141_
	);
	LUT4 #(
		.INIT('habef)
	) name13241 (
		_w8905_,
		_w8908_,
		_w15140_,
		_w15141_,
		_w15142_
	);
	LUT3 #(
		.INIT('h2a)
	) name13242 (
		\m5_addr_i[2]_pad ,
		_w8910_,
		_w8911_,
		_w15143_
	);
	LUT3 #(
		.INIT('h2a)
	) name13243 (
		\m1_addr_i[2]_pad ,
		_w8910_,
		_w8911_,
		_w15144_
	);
	LUT4 #(
		.INIT('h57df)
	) name13244 (
		_w8905_,
		_w8908_,
		_w15143_,
		_w15144_,
		_w15145_
	);
	LUT3 #(
		.INIT('h2a)
	) name13245 (
		\m3_addr_i[2]_pad ,
		_w8910_,
		_w8911_,
		_w15146_
	);
	LUT3 #(
		.INIT('h80)
	) name13246 (
		\m4_addr_i[2]_pad ,
		_w8910_,
		_w8911_,
		_w15147_
	);
	LUT4 #(
		.INIT('h9dbf)
	) name13247 (
		_w8905_,
		_w8908_,
		_w15146_,
		_w15147_,
		_w15148_
	);
	LUT4 #(
		.INIT('h7fff)
	) name13248 (
		_w15139_,
		_w15142_,
		_w15145_,
		_w15148_,
		_w15149_
	);
	LUT3 #(
		.INIT('h2a)
	) name13249 (
		\m1_addr_i[30]_pad ,
		_w8910_,
		_w8911_,
		_w15150_
	);
	LUT3 #(
		.INIT('h80)
	) name13250 (
		\m2_addr_i[30]_pad ,
		_w8910_,
		_w8911_,
		_w15151_
	);
	LUT4 #(
		.INIT('h3b7f)
	) name13251 (
		_w8905_,
		_w8908_,
		_w15150_,
		_w15151_,
		_w15152_
	);
	LUT3 #(
		.INIT('h2a)
	) name13252 (
		\m3_addr_i[30]_pad ,
		_w8910_,
		_w8911_,
		_w15153_
	);
	LUT3 #(
		.INIT('h80)
	) name13253 (
		\m6_addr_i[30]_pad ,
		_w8910_,
		_w8911_,
		_w15154_
	);
	LUT4 #(
		.INIT('haebf)
	) name13254 (
		_w8905_,
		_w8908_,
		_w15153_,
		_w15154_,
		_w15155_
	);
	LUT3 #(
		.INIT('h80)
	) name13255 (
		\m4_addr_i[30]_pad ,
		_w8910_,
		_w8911_,
		_w15156_
	);
	LUT3 #(
		.INIT('h2a)
	) name13256 (
		\m5_addr_i[30]_pad ,
		_w8910_,
		_w8911_,
		_w15157_
	);
	LUT3 #(
		.INIT('h57)
	) name13257 (
		_w8929_,
		_w15156_,
		_w15157_,
		_w15158_
	);
	LUT3 #(
		.INIT('h80)
	) name13258 (
		\m0_addr_i[30]_pad ,
		_w8910_,
		_w8911_,
		_w15159_
	);
	LUT3 #(
		.INIT('h2a)
	) name13259 (
		\m7_addr_i[30]_pad ,
		_w8910_,
		_w8911_,
		_w15160_
	);
	LUT4 #(
		.INIT('h6e7f)
	) name13260 (
		_w8905_,
		_w8908_,
		_w15159_,
		_w15160_,
		_w15161_
	);
	LUT4 #(
		.INIT('h7fff)
	) name13261 (
		_w15152_,
		_w15155_,
		_w15158_,
		_w15161_,
		_w15162_
	);
	LUT3 #(
		.INIT('h2a)
	) name13262 (
		\m5_addr_i[31]_pad ,
		_w8910_,
		_w8911_,
		_w15163_
	);
	LUT3 #(
		.INIT('h80)
	) name13263 (
		\m6_addr_i[31]_pad ,
		_w8910_,
		_w8911_,
		_w15164_
	);
	LUT4 #(
		.INIT('hcedf)
	) name13264 (
		_w8905_,
		_w8908_,
		_w15163_,
		_w15164_,
		_w15165_
	);
	LUT3 #(
		.INIT('h80)
	) name13265 (
		\m0_addr_i[31]_pad ,
		_w8910_,
		_w8911_,
		_w15166_
	);
	LUT3 #(
		.INIT('h80)
	) name13266 (
		\m4_addr_i[31]_pad ,
		_w8910_,
		_w8911_,
		_w15167_
	);
	LUT4 #(
		.INIT('h5d7f)
	) name13267 (
		_w8905_,
		_w8908_,
		_w15166_,
		_w15167_,
		_w15168_
	);
	LUT3 #(
		.INIT('h2a)
	) name13268 (
		\m7_addr_i[31]_pad ,
		_w8910_,
		_w8911_,
		_w15169_
	);
	LUT3 #(
		.INIT('h2a)
	) name13269 (
		\m3_addr_i[31]_pad ,
		_w8910_,
		_w8911_,
		_w15170_
	);
	LUT4 #(
		.INIT('habef)
	) name13270 (
		_w8905_,
		_w8908_,
		_w15169_,
		_w15170_,
		_w15171_
	);
	LUT3 #(
		.INIT('h2a)
	) name13271 (
		\m1_addr_i[31]_pad ,
		_w8910_,
		_w8911_,
		_w15172_
	);
	LUT3 #(
		.INIT('h80)
	) name13272 (
		\m2_addr_i[31]_pad ,
		_w8910_,
		_w8911_,
		_w15173_
	);
	LUT4 #(
		.INIT('h3b7f)
	) name13273 (
		_w8905_,
		_w8908_,
		_w15172_,
		_w15173_,
		_w15174_
	);
	LUT4 #(
		.INIT('h7fff)
	) name13274 (
		_w15165_,
		_w15168_,
		_w15171_,
		_w15174_,
		_w15175_
	);
	LUT3 #(
		.INIT('h80)
	) name13275 (
		\m6_addr_i[3]_pad ,
		_w8910_,
		_w8911_,
		_w15176_
	);
	LUT3 #(
		.INIT('h2a)
	) name13276 (
		\m5_addr_i[3]_pad ,
		_w8910_,
		_w8911_,
		_w15177_
	);
	LUT4 #(
		.INIT('hcdef)
	) name13277 (
		_w8905_,
		_w8908_,
		_w15176_,
		_w15177_,
		_w15178_
	);
	LUT3 #(
		.INIT('h80)
	) name13278 (
		\m0_addr_i[3]_pad ,
		_w8910_,
		_w8911_,
		_w15179_
	);
	LUT3 #(
		.INIT('h80)
	) name13279 (
		\m2_addr_i[3]_pad ,
		_w8910_,
		_w8911_,
		_w15180_
	);
	LUT4 #(
		.INIT('h3b7f)
	) name13280 (
		_w8905_,
		_w8908_,
		_w15179_,
		_w15180_,
		_w15181_
	);
	LUT3 #(
		.INIT('h2a)
	) name13281 (
		\m7_addr_i[3]_pad ,
		_w8910_,
		_w8911_,
		_w15182_
	);
	LUT3 #(
		.INIT('h2a)
	) name13282 (
		\m1_addr_i[3]_pad ,
		_w8910_,
		_w8911_,
		_w15183_
	);
	LUT4 #(
		.INIT('h67ef)
	) name13283 (
		_w8905_,
		_w8908_,
		_w15182_,
		_w15183_,
		_w15184_
	);
	LUT3 #(
		.INIT('h2a)
	) name13284 (
		\m3_addr_i[3]_pad ,
		_w8910_,
		_w8911_,
		_w15185_
	);
	LUT3 #(
		.INIT('h80)
	) name13285 (
		\m4_addr_i[3]_pad ,
		_w8910_,
		_w8911_,
		_w15186_
	);
	LUT4 #(
		.INIT('h9dbf)
	) name13286 (
		_w8905_,
		_w8908_,
		_w15185_,
		_w15186_,
		_w15187_
	);
	LUT4 #(
		.INIT('h7fff)
	) name13287 (
		_w15178_,
		_w15181_,
		_w15184_,
		_w15187_,
		_w15188_
	);
	LUT3 #(
		.INIT('h2a)
	) name13288 (
		\m1_addr_i[4]_pad ,
		_w8910_,
		_w8911_,
		_w15189_
	);
	LUT3 #(
		.INIT('h80)
	) name13289 (
		\m2_addr_i[4]_pad ,
		_w8910_,
		_w8911_,
		_w15190_
	);
	LUT4 #(
		.INIT('h3b7f)
	) name13290 (
		_w8905_,
		_w8908_,
		_w15189_,
		_w15190_,
		_w15191_
	);
	LUT3 #(
		.INIT('h80)
	) name13291 (
		\m0_addr_i[4]_pad ,
		_w8910_,
		_w8911_,
		_w15192_
	);
	LUT3 #(
		.INIT('h80)
	) name13292 (
		\m4_addr_i[4]_pad ,
		_w8910_,
		_w8911_,
		_w15193_
	);
	LUT4 #(
		.INIT('h5d7f)
	) name13293 (
		_w8905_,
		_w8908_,
		_w15192_,
		_w15193_,
		_w15194_
	);
	LUT3 #(
		.INIT('h2a)
	) name13294 (
		\m7_addr_i[4]_pad ,
		_w8910_,
		_w8911_,
		_w15195_
	);
	LUT3 #(
		.INIT('h2a)
	) name13295 (
		\m3_addr_i[4]_pad ,
		_w8910_,
		_w8911_,
		_w15196_
	);
	LUT4 #(
		.INIT('habef)
	) name13296 (
		_w8905_,
		_w8908_,
		_w15195_,
		_w15196_,
		_w15197_
	);
	LUT3 #(
		.INIT('h80)
	) name13297 (
		\m6_addr_i[4]_pad ,
		_w8910_,
		_w8911_,
		_w15198_
	);
	LUT3 #(
		.INIT('h2a)
	) name13298 (
		\m5_addr_i[4]_pad ,
		_w8910_,
		_w8911_,
		_w15199_
	);
	LUT4 #(
		.INIT('hcdef)
	) name13299 (
		_w8905_,
		_w8908_,
		_w15198_,
		_w15199_,
		_w15200_
	);
	LUT4 #(
		.INIT('h7fff)
	) name13300 (
		_w15191_,
		_w15194_,
		_w15197_,
		_w15200_,
		_w15201_
	);
	LUT3 #(
		.INIT('h2a)
	) name13301 (
		\m1_addr_i[5]_pad ,
		_w8910_,
		_w8911_,
		_w15202_
	);
	LUT3 #(
		.INIT('h80)
	) name13302 (
		\m2_addr_i[5]_pad ,
		_w8910_,
		_w8911_,
		_w15203_
	);
	LUT4 #(
		.INIT('h3b7f)
	) name13303 (
		_w8905_,
		_w8908_,
		_w15202_,
		_w15203_,
		_w15204_
	);
	LUT3 #(
		.INIT('h80)
	) name13304 (
		\m0_addr_i[5]_pad ,
		_w8910_,
		_w8911_,
		_w15205_
	);
	LUT3 #(
		.INIT('h80)
	) name13305 (
		\m4_addr_i[5]_pad ,
		_w8910_,
		_w8911_,
		_w15206_
	);
	LUT4 #(
		.INIT('h5d7f)
	) name13306 (
		_w8905_,
		_w8908_,
		_w15205_,
		_w15206_,
		_w15207_
	);
	LUT3 #(
		.INIT('h2a)
	) name13307 (
		\m7_addr_i[5]_pad ,
		_w8910_,
		_w8911_,
		_w15208_
	);
	LUT3 #(
		.INIT('h2a)
	) name13308 (
		\m3_addr_i[5]_pad ,
		_w8910_,
		_w8911_,
		_w15209_
	);
	LUT4 #(
		.INIT('habef)
	) name13309 (
		_w8905_,
		_w8908_,
		_w15208_,
		_w15209_,
		_w15210_
	);
	LUT3 #(
		.INIT('h80)
	) name13310 (
		\m6_addr_i[5]_pad ,
		_w8910_,
		_w8911_,
		_w15211_
	);
	LUT3 #(
		.INIT('h2a)
	) name13311 (
		\m5_addr_i[5]_pad ,
		_w8910_,
		_w8911_,
		_w15212_
	);
	LUT4 #(
		.INIT('hcdef)
	) name13312 (
		_w8905_,
		_w8908_,
		_w15211_,
		_w15212_,
		_w15213_
	);
	LUT4 #(
		.INIT('h7fff)
	) name13313 (
		_w15204_,
		_w15207_,
		_w15210_,
		_w15213_,
		_w15214_
	);
	LUT3 #(
		.INIT('h80)
	) name13314 (
		\m0_addr_i[6]_pad ,
		_w8910_,
		_w8911_,
		_w15215_
	);
	LUT3 #(
		.INIT('h2a)
	) name13315 (
		\m7_addr_i[6]_pad ,
		_w8910_,
		_w8911_,
		_w15216_
	);
	LUT4 #(
		.INIT('h6e7f)
	) name13316 (
		_w8905_,
		_w8908_,
		_w15215_,
		_w15216_,
		_w15217_
	);
	LUT3 #(
		.INIT('h2a)
	) name13317 (
		\m3_addr_i[6]_pad ,
		_w8910_,
		_w8911_,
		_w15218_
	);
	LUT3 #(
		.INIT('h80)
	) name13318 (
		\m2_addr_i[6]_pad ,
		_w8910_,
		_w8911_,
		_w15219_
	);
	LUT3 #(
		.INIT('h57)
	) name13319 (
		_w8909_,
		_w15218_,
		_w15219_,
		_w15220_
	);
	LUT3 #(
		.INIT('h80)
	) name13320 (
		\m4_addr_i[6]_pad ,
		_w8910_,
		_w8911_,
		_w15221_
	);
	LUT3 #(
		.INIT('h2a)
	) name13321 (
		\m1_addr_i[6]_pad ,
		_w8910_,
		_w8911_,
		_w15222_
	);
	LUT4 #(
		.INIT('h57df)
	) name13322 (
		_w8905_,
		_w8908_,
		_w15221_,
		_w15222_,
		_w15223_
	);
	LUT3 #(
		.INIT('h80)
	) name13323 (
		\m6_addr_i[6]_pad ,
		_w8910_,
		_w8911_,
		_w15224_
	);
	LUT3 #(
		.INIT('h2a)
	) name13324 (
		\m5_addr_i[6]_pad ,
		_w8910_,
		_w8911_,
		_w15225_
	);
	LUT4 #(
		.INIT('hcdef)
	) name13325 (
		_w8905_,
		_w8908_,
		_w15224_,
		_w15225_,
		_w15226_
	);
	LUT4 #(
		.INIT('h7fff)
	) name13326 (
		_w15217_,
		_w15220_,
		_w15223_,
		_w15226_,
		_w15227_
	);
	LUT3 #(
		.INIT('h80)
	) name13327 (
		\m0_addr_i[7]_pad ,
		_w8910_,
		_w8911_,
		_w15228_
	);
	LUT3 #(
		.INIT('h2a)
	) name13328 (
		\m7_addr_i[7]_pad ,
		_w8910_,
		_w8911_,
		_w15229_
	);
	LUT4 #(
		.INIT('h6e7f)
	) name13329 (
		_w8905_,
		_w8908_,
		_w15228_,
		_w15229_,
		_w15230_
	);
	LUT3 #(
		.INIT('h2a)
	) name13330 (
		\m1_addr_i[7]_pad ,
		_w8910_,
		_w8911_,
		_w15231_
	);
	LUT3 #(
		.INIT('h2a)
	) name13331 (
		\m5_addr_i[7]_pad ,
		_w8910_,
		_w8911_,
		_w15232_
	);
	LUT4 #(
		.INIT('h5d7f)
	) name13332 (
		_w8905_,
		_w8908_,
		_w15231_,
		_w15232_,
		_w15233_
	);
	LUT3 #(
		.INIT('h80)
	) name13333 (
		\m2_addr_i[7]_pad ,
		_w8910_,
		_w8911_,
		_w15234_
	);
	LUT3 #(
		.INIT('h80)
	) name13334 (
		\m6_addr_i[7]_pad ,
		_w8910_,
		_w8911_,
		_w15235_
	);
	LUT4 #(
		.INIT('haebf)
	) name13335 (
		_w8905_,
		_w8908_,
		_w15234_,
		_w15235_,
		_w15236_
	);
	LUT3 #(
		.INIT('h2a)
	) name13336 (
		\m3_addr_i[7]_pad ,
		_w8910_,
		_w8911_,
		_w15237_
	);
	LUT3 #(
		.INIT('h80)
	) name13337 (
		\m4_addr_i[7]_pad ,
		_w8910_,
		_w8911_,
		_w15238_
	);
	LUT4 #(
		.INIT('h9dbf)
	) name13338 (
		_w8905_,
		_w8908_,
		_w15237_,
		_w15238_,
		_w15239_
	);
	LUT4 #(
		.INIT('h7fff)
	) name13339 (
		_w15230_,
		_w15233_,
		_w15236_,
		_w15239_,
		_w15240_
	);
	LUT3 #(
		.INIT('h80)
	) name13340 (
		\m0_addr_i[8]_pad ,
		_w8910_,
		_w8911_,
		_w15241_
	);
	LUT3 #(
		.INIT('h2a)
	) name13341 (
		\m7_addr_i[8]_pad ,
		_w8910_,
		_w8911_,
		_w15242_
	);
	LUT4 #(
		.INIT('h6e7f)
	) name13342 (
		_w8905_,
		_w8908_,
		_w15241_,
		_w15242_,
		_w15243_
	);
	LUT3 #(
		.INIT('h80)
	) name13343 (
		\m6_addr_i[8]_pad ,
		_w8910_,
		_w8911_,
		_w15244_
	);
	LUT3 #(
		.INIT('h80)
	) name13344 (
		\m2_addr_i[8]_pad ,
		_w8910_,
		_w8911_,
		_w15245_
	);
	LUT4 #(
		.INIT('habef)
	) name13345 (
		_w8905_,
		_w8908_,
		_w15244_,
		_w15245_,
		_w15246_
	);
	LUT3 #(
		.INIT('h2a)
	) name13346 (
		\m5_addr_i[8]_pad ,
		_w8910_,
		_w8911_,
		_w15247_
	);
	LUT3 #(
		.INIT('h2a)
	) name13347 (
		\m1_addr_i[8]_pad ,
		_w8910_,
		_w8911_,
		_w15248_
	);
	LUT4 #(
		.INIT('h57df)
	) name13348 (
		_w8905_,
		_w8908_,
		_w15247_,
		_w15248_,
		_w15249_
	);
	LUT3 #(
		.INIT('h2a)
	) name13349 (
		\m3_addr_i[8]_pad ,
		_w8910_,
		_w8911_,
		_w15250_
	);
	LUT3 #(
		.INIT('h80)
	) name13350 (
		\m4_addr_i[8]_pad ,
		_w8910_,
		_w8911_,
		_w15251_
	);
	LUT4 #(
		.INIT('h9dbf)
	) name13351 (
		_w8905_,
		_w8908_,
		_w15250_,
		_w15251_,
		_w15252_
	);
	LUT4 #(
		.INIT('h7fff)
	) name13352 (
		_w15243_,
		_w15246_,
		_w15249_,
		_w15252_,
		_w15253_
	);
	LUT3 #(
		.INIT('h2a)
	) name13353 (
		\m1_addr_i[9]_pad ,
		_w8910_,
		_w8911_,
		_w15254_
	);
	LUT3 #(
		.INIT('h80)
	) name13354 (
		\m2_addr_i[9]_pad ,
		_w8910_,
		_w8911_,
		_w15255_
	);
	LUT4 #(
		.INIT('h3b7f)
	) name13355 (
		_w8905_,
		_w8908_,
		_w15254_,
		_w15255_,
		_w15256_
	);
	LUT3 #(
		.INIT('h80)
	) name13356 (
		\m6_addr_i[9]_pad ,
		_w8910_,
		_w8911_,
		_w15257_
	);
	LUT3 #(
		.INIT('h2a)
	) name13357 (
		\m7_addr_i[9]_pad ,
		_w8910_,
		_w8911_,
		_w15258_
	);
	LUT3 #(
		.INIT('h57)
	) name13358 (
		_w8917_,
		_w15257_,
		_w15258_,
		_w15259_
	);
	LUT3 #(
		.INIT('h2a)
	) name13359 (
		\m5_addr_i[9]_pad ,
		_w8910_,
		_w8911_,
		_w15260_
	);
	LUT3 #(
		.INIT('h80)
	) name13360 (
		\m0_addr_i[9]_pad ,
		_w8910_,
		_w8911_,
		_w15261_
	);
	LUT4 #(
		.INIT('h57df)
	) name13361 (
		_w8905_,
		_w8908_,
		_w15260_,
		_w15261_,
		_w15262_
	);
	LUT3 #(
		.INIT('h2a)
	) name13362 (
		\m3_addr_i[9]_pad ,
		_w8910_,
		_w8911_,
		_w15263_
	);
	LUT3 #(
		.INIT('h80)
	) name13363 (
		\m4_addr_i[9]_pad ,
		_w8910_,
		_w8911_,
		_w15264_
	);
	LUT4 #(
		.INIT('h9dbf)
	) name13364 (
		_w8905_,
		_w8908_,
		_w15263_,
		_w15264_,
		_w15265_
	);
	LUT4 #(
		.INIT('h7fff)
	) name13365 (
		_w15256_,
		_w15259_,
		_w15262_,
		_w15265_,
		_w15266_
	);
	LUT3 #(
		.INIT('h2a)
	) name13366 (
		\m3_data_i[0]_pad ,
		_w8910_,
		_w8911_,
		_w15267_
	);
	LUT3 #(
		.INIT('h80)
	) name13367 (
		\m4_data_i[0]_pad ,
		_w8910_,
		_w8911_,
		_w15268_
	);
	LUT4 #(
		.INIT('h9dbf)
	) name13368 (
		_w8905_,
		_w8908_,
		_w15267_,
		_w15268_,
		_w15269_
	);
	LUT3 #(
		.INIT('h2a)
	) name13369 (
		\m1_data_i[0]_pad ,
		_w8910_,
		_w8911_,
		_w15270_
	);
	LUT3 #(
		.INIT('h2a)
	) name13370 (
		\m5_data_i[0]_pad ,
		_w8910_,
		_w8911_,
		_w15271_
	);
	LUT4 #(
		.INIT('h5d7f)
	) name13371 (
		_w8905_,
		_w8908_,
		_w15270_,
		_w15271_,
		_w15272_
	);
	LUT3 #(
		.INIT('h80)
	) name13372 (
		\m2_data_i[0]_pad ,
		_w8910_,
		_w8911_,
		_w15273_
	);
	LUT3 #(
		.INIT('h80)
	) name13373 (
		\m6_data_i[0]_pad ,
		_w8910_,
		_w8911_,
		_w15274_
	);
	LUT4 #(
		.INIT('haebf)
	) name13374 (
		_w8905_,
		_w8908_,
		_w15273_,
		_w15274_,
		_w15275_
	);
	LUT3 #(
		.INIT('h80)
	) name13375 (
		\m0_data_i[0]_pad ,
		_w8910_,
		_w8911_,
		_w15276_
	);
	LUT3 #(
		.INIT('h2a)
	) name13376 (
		\m7_data_i[0]_pad ,
		_w8910_,
		_w8911_,
		_w15277_
	);
	LUT4 #(
		.INIT('h6e7f)
	) name13377 (
		_w8905_,
		_w8908_,
		_w15276_,
		_w15277_,
		_w15278_
	);
	LUT4 #(
		.INIT('h7fff)
	) name13378 (
		_w15269_,
		_w15272_,
		_w15275_,
		_w15278_,
		_w15279_
	);
	LUT3 #(
		.INIT('h80)
	) name13379 (
		\m0_data_i[10]_pad ,
		_w8910_,
		_w8911_,
		_w15280_
	);
	LUT3 #(
		.INIT('h2a)
	) name13380 (
		\m7_data_i[10]_pad ,
		_w8910_,
		_w8911_,
		_w15281_
	);
	LUT4 #(
		.INIT('h6e7f)
	) name13381 (
		_w8905_,
		_w8908_,
		_w15280_,
		_w15281_,
		_w15282_
	);
	LUT3 #(
		.INIT('h2a)
	) name13382 (
		\m1_data_i[10]_pad ,
		_w8910_,
		_w8911_,
		_w15283_
	);
	LUT3 #(
		.INIT('h80)
	) name13383 (
		\m4_data_i[10]_pad ,
		_w8910_,
		_w8911_,
		_w15284_
	);
	LUT4 #(
		.INIT('h5d7f)
	) name13384 (
		_w8905_,
		_w8908_,
		_w15283_,
		_w15284_,
		_w15285_
	);
	LUT3 #(
		.INIT('h80)
	) name13385 (
		\m2_data_i[10]_pad ,
		_w8910_,
		_w8911_,
		_w15286_
	);
	LUT3 #(
		.INIT('h2a)
	) name13386 (
		\m3_data_i[10]_pad ,
		_w8910_,
		_w8911_,
		_w15287_
	);
	LUT3 #(
		.INIT('h57)
	) name13387 (
		_w8909_,
		_w15286_,
		_w15287_,
		_w15288_
	);
	LUT3 #(
		.INIT('h80)
	) name13388 (
		\m6_data_i[10]_pad ,
		_w8910_,
		_w8911_,
		_w15289_
	);
	LUT3 #(
		.INIT('h2a)
	) name13389 (
		\m5_data_i[10]_pad ,
		_w8910_,
		_w8911_,
		_w15290_
	);
	LUT4 #(
		.INIT('hcdef)
	) name13390 (
		_w8905_,
		_w8908_,
		_w15289_,
		_w15290_,
		_w15291_
	);
	LUT4 #(
		.INIT('h7fff)
	) name13391 (
		_w15282_,
		_w15285_,
		_w15288_,
		_w15291_,
		_w15292_
	);
	LUT3 #(
		.INIT('h2a)
	) name13392 (
		\m1_data_i[11]_pad ,
		_w8910_,
		_w8911_,
		_w15293_
	);
	LUT3 #(
		.INIT('h80)
	) name13393 (
		\m2_data_i[11]_pad ,
		_w8910_,
		_w8911_,
		_w15294_
	);
	LUT4 #(
		.INIT('h3b7f)
	) name13394 (
		_w8905_,
		_w8908_,
		_w15293_,
		_w15294_,
		_w15295_
	);
	LUT3 #(
		.INIT('h80)
	) name13395 (
		\m0_data_i[11]_pad ,
		_w8910_,
		_w8911_,
		_w15296_
	);
	LUT3 #(
		.INIT('h80)
	) name13396 (
		\m4_data_i[11]_pad ,
		_w8910_,
		_w8911_,
		_w15297_
	);
	LUT4 #(
		.INIT('h5d7f)
	) name13397 (
		_w8905_,
		_w8908_,
		_w15296_,
		_w15297_,
		_w15298_
	);
	LUT3 #(
		.INIT('h2a)
	) name13398 (
		\m7_data_i[11]_pad ,
		_w8910_,
		_w8911_,
		_w15299_
	);
	LUT3 #(
		.INIT('h2a)
	) name13399 (
		\m3_data_i[11]_pad ,
		_w8910_,
		_w8911_,
		_w15300_
	);
	LUT4 #(
		.INIT('habef)
	) name13400 (
		_w8905_,
		_w8908_,
		_w15299_,
		_w15300_,
		_w15301_
	);
	LUT3 #(
		.INIT('h80)
	) name13401 (
		\m6_data_i[11]_pad ,
		_w8910_,
		_w8911_,
		_w15302_
	);
	LUT3 #(
		.INIT('h2a)
	) name13402 (
		\m5_data_i[11]_pad ,
		_w8910_,
		_w8911_,
		_w15303_
	);
	LUT4 #(
		.INIT('hcdef)
	) name13403 (
		_w8905_,
		_w8908_,
		_w15302_,
		_w15303_,
		_w15304_
	);
	LUT4 #(
		.INIT('h7fff)
	) name13404 (
		_w15295_,
		_w15298_,
		_w15301_,
		_w15304_,
		_w15305_
	);
	LUT3 #(
		.INIT('h2a)
	) name13405 (
		\m1_data_i[12]_pad ,
		_w8910_,
		_w8911_,
		_w15306_
	);
	LUT3 #(
		.INIT('h80)
	) name13406 (
		\m2_data_i[12]_pad ,
		_w8910_,
		_w8911_,
		_w15307_
	);
	LUT4 #(
		.INIT('h3b7f)
	) name13407 (
		_w8905_,
		_w8908_,
		_w15306_,
		_w15307_,
		_w15308_
	);
	LUT3 #(
		.INIT('h80)
	) name13408 (
		\m0_data_i[12]_pad ,
		_w8910_,
		_w8911_,
		_w15309_
	);
	LUT3 #(
		.INIT('h80)
	) name13409 (
		\m4_data_i[12]_pad ,
		_w8910_,
		_w8911_,
		_w15310_
	);
	LUT4 #(
		.INIT('h5d7f)
	) name13410 (
		_w8905_,
		_w8908_,
		_w15309_,
		_w15310_,
		_w15311_
	);
	LUT3 #(
		.INIT('h2a)
	) name13411 (
		\m7_data_i[12]_pad ,
		_w8910_,
		_w8911_,
		_w15312_
	);
	LUT3 #(
		.INIT('h2a)
	) name13412 (
		\m3_data_i[12]_pad ,
		_w8910_,
		_w8911_,
		_w15313_
	);
	LUT4 #(
		.INIT('habef)
	) name13413 (
		_w8905_,
		_w8908_,
		_w15312_,
		_w15313_,
		_w15314_
	);
	LUT3 #(
		.INIT('h80)
	) name13414 (
		\m6_data_i[12]_pad ,
		_w8910_,
		_w8911_,
		_w15315_
	);
	LUT3 #(
		.INIT('h2a)
	) name13415 (
		\m5_data_i[12]_pad ,
		_w8910_,
		_w8911_,
		_w15316_
	);
	LUT4 #(
		.INIT('hcdef)
	) name13416 (
		_w8905_,
		_w8908_,
		_w15315_,
		_w15316_,
		_w15317_
	);
	LUT4 #(
		.INIT('h7fff)
	) name13417 (
		_w15308_,
		_w15311_,
		_w15314_,
		_w15317_,
		_w15318_
	);
	LUT3 #(
		.INIT('h80)
	) name13418 (
		\m0_data_i[13]_pad ,
		_w8910_,
		_w8911_,
		_w15319_
	);
	LUT3 #(
		.INIT('h2a)
	) name13419 (
		\m7_data_i[13]_pad ,
		_w8910_,
		_w8911_,
		_w15320_
	);
	LUT4 #(
		.INIT('h6e7f)
	) name13420 (
		_w8905_,
		_w8908_,
		_w15319_,
		_w15320_,
		_w15321_
	);
	LUT3 #(
		.INIT('h80)
	) name13421 (
		\m6_data_i[13]_pad ,
		_w8910_,
		_w8911_,
		_w15322_
	);
	LUT3 #(
		.INIT('h80)
	) name13422 (
		\m2_data_i[13]_pad ,
		_w8910_,
		_w8911_,
		_w15323_
	);
	LUT4 #(
		.INIT('habef)
	) name13423 (
		_w8905_,
		_w8908_,
		_w15322_,
		_w15323_,
		_w15324_
	);
	LUT3 #(
		.INIT('h2a)
	) name13424 (
		\m5_data_i[13]_pad ,
		_w8910_,
		_w8911_,
		_w15325_
	);
	LUT3 #(
		.INIT('h2a)
	) name13425 (
		\m1_data_i[13]_pad ,
		_w8910_,
		_w8911_,
		_w15326_
	);
	LUT4 #(
		.INIT('h57df)
	) name13426 (
		_w8905_,
		_w8908_,
		_w15325_,
		_w15326_,
		_w15327_
	);
	LUT3 #(
		.INIT('h2a)
	) name13427 (
		\m3_data_i[13]_pad ,
		_w8910_,
		_w8911_,
		_w15328_
	);
	LUT3 #(
		.INIT('h80)
	) name13428 (
		\m4_data_i[13]_pad ,
		_w8910_,
		_w8911_,
		_w15329_
	);
	LUT4 #(
		.INIT('h9dbf)
	) name13429 (
		_w8905_,
		_w8908_,
		_w15328_,
		_w15329_,
		_w15330_
	);
	LUT4 #(
		.INIT('h7fff)
	) name13430 (
		_w15321_,
		_w15324_,
		_w15327_,
		_w15330_,
		_w15331_
	);
	LUT3 #(
		.INIT('h80)
	) name13431 (
		\m6_data_i[14]_pad ,
		_w8910_,
		_w8911_,
		_w15332_
	);
	LUT3 #(
		.INIT('h2a)
	) name13432 (
		\m5_data_i[14]_pad ,
		_w8910_,
		_w8911_,
		_w15333_
	);
	LUT4 #(
		.INIT('hcdef)
	) name13433 (
		_w8905_,
		_w8908_,
		_w15332_,
		_w15333_,
		_w15334_
	);
	LUT3 #(
		.INIT('h2a)
	) name13434 (
		\m3_data_i[14]_pad ,
		_w8910_,
		_w8911_,
		_w15335_
	);
	LUT3 #(
		.INIT('h80)
	) name13435 (
		\m2_data_i[14]_pad ,
		_w8910_,
		_w8911_,
		_w15336_
	);
	LUT3 #(
		.INIT('h57)
	) name13436 (
		_w8909_,
		_w15335_,
		_w15336_,
		_w15337_
	);
	LUT3 #(
		.INIT('h80)
	) name13437 (
		\m4_data_i[14]_pad ,
		_w8910_,
		_w8911_,
		_w15338_
	);
	LUT3 #(
		.INIT('h2a)
	) name13438 (
		\m1_data_i[14]_pad ,
		_w8910_,
		_w8911_,
		_w15339_
	);
	LUT4 #(
		.INIT('h57df)
	) name13439 (
		_w8905_,
		_w8908_,
		_w15338_,
		_w15339_,
		_w15340_
	);
	LUT3 #(
		.INIT('h80)
	) name13440 (
		\m0_data_i[14]_pad ,
		_w8910_,
		_w8911_,
		_w15341_
	);
	LUT3 #(
		.INIT('h2a)
	) name13441 (
		\m7_data_i[14]_pad ,
		_w8910_,
		_w8911_,
		_w15342_
	);
	LUT4 #(
		.INIT('h6e7f)
	) name13442 (
		_w8905_,
		_w8908_,
		_w15341_,
		_w15342_,
		_w15343_
	);
	LUT4 #(
		.INIT('h7fff)
	) name13443 (
		_w15334_,
		_w15337_,
		_w15340_,
		_w15343_,
		_w15344_
	);
	LUT3 #(
		.INIT('h2a)
	) name13444 (
		\m3_data_i[15]_pad ,
		_w8910_,
		_w8911_,
		_w15345_
	);
	LUT3 #(
		.INIT('h80)
	) name13445 (
		\m4_data_i[15]_pad ,
		_w8910_,
		_w8911_,
		_w15346_
	);
	LUT4 #(
		.INIT('h9dbf)
	) name13446 (
		_w8905_,
		_w8908_,
		_w15345_,
		_w15346_,
		_w15347_
	);
	LUT3 #(
		.INIT('h2a)
	) name13447 (
		\m1_data_i[15]_pad ,
		_w8910_,
		_w8911_,
		_w15348_
	);
	LUT3 #(
		.INIT('h2a)
	) name13448 (
		\m5_data_i[15]_pad ,
		_w8910_,
		_w8911_,
		_w15349_
	);
	LUT4 #(
		.INIT('h5d7f)
	) name13449 (
		_w8905_,
		_w8908_,
		_w15348_,
		_w15349_,
		_w15350_
	);
	LUT3 #(
		.INIT('h80)
	) name13450 (
		\m2_data_i[15]_pad ,
		_w8910_,
		_w8911_,
		_w15351_
	);
	LUT3 #(
		.INIT('h80)
	) name13451 (
		\m6_data_i[15]_pad ,
		_w8910_,
		_w8911_,
		_w15352_
	);
	LUT4 #(
		.INIT('haebf)
	) name13452 (
		_w8905_,
		_w8908_,
		_w15351_,
		_w15352_,
		_w15353_
	);
	LUT3 #(
		.INIT('h80)
	) name13453 (
		\m0_data_i[15]_pad ,
		_w8910_,
		_w8911_,
		_w15354_
	);
	LUT3 #(
		.INIT('h2a)
	) name13454 (
		\m7_data_i[15]_pad ,
		_w8910_,
		_w8911_,
		_w15355_
	);
	LUT4 #(
		.INIT('h6e7f)
	) name13455 (
		_w8905_,
		_w8908_,
		_w15354_,
		_w15355_,
		_w15356_
	);
	LUT4 #(
		.INIT('h7fff)
	) name13456 (
		_w15347_,
		_w15350_,
		_w15353_,
		_w15356_,
		_w15357_
	);
	LUT3 #(
		.INIT('h2a)
	) name13457 (
		\m3_data_i[16]_pad ,
		_w8910_,
		_w8911_,
		_w15358_
	);
	LUT3 #(
		.INIT('h80)
	) name13458 (
		\m4_data_i[16]_pad ,
		_w8910_,
		_w8911_,
		_w15359_
	);
	LUT4 #(
		.INIT('h9dbf)
	) name13459 (
		_w8905_,
		_w8908_,
		_w15358_,
		_w15359_,
		_w15360_
	);
	LUT3 #(
		.INIT('h2a)
	) name13460 (
		\m1_data_i[16]_pad ,
		_w8910_,
		_w8911_,
		_w15361_
	);
	LUT3 #(
		.INIT('h2a)
	) name13461 (
		\m5_data_i[16]_pad ,
		_w8910_,
		_w8911_,
		_w15362_
	);
	LUT4 #(
		.INIT('h5d7f)
	) name13462 (
		_w8905_,
		_w8908_,
		_w15361_,
		_w15362_,
		_w15363_
	);
	LUT3 #(
		.INIT('h80)
	) name13463 (
		\m2_data_i[16]_pad ,
		_w8910_,
		_w8911_,
		_w15364_
	);
	LUT3 #(
		.INIT('h80)
	) name13464 (
		\m6_data_i[16]_pad ,
		_w8910_,
		_w8911_,
		_w15365_
	);
	LUT4 #(
		.INIT('haebf)
	) name13465 (
		_w8905_,
		_w8908_,
		_w15364_,
		_w15365_,
		_w15366_
	);
	LUT3 #(
		.INIT('h80)
	) name13466 (
		\m0_data_i[16]_pad ,
		_w8910_,
		_w8911_,
		_w15367_
	);
	LUT3 #(
		.INIT('h2a)
	) name13467 (
		\m7_data_i[16]_pad ,
		_w8910_,
		_w8911_,
		_w15368_
	);
	LUT4 #(
		.INIT('h6e7f)
	) name13468 (
		_w8905_,
		_w8908_,
		_w15367_,
		_w15368_,
		_w15369_
	);
	LUT4 #(
		.INIT('h7fff)
	) name13469 (
		_w15360_,
		_w15363_,
		_w15366_,
		_w15369_,
		_w15370_
	);
	LUT3 #(
		.INIT('h80)
	) name13470 (
		\m6_data_i[17]_pad ,
		_w8910_,
		_w8911_,
		_w15371_
	);
	LUT3 #(
		.INIT('h2a)
	) name13471 (
		\m5_data_i[17]_pad ,
		_w8910_,
		_w8911_,
		_w15372_
	);
	LUT4 #(
		.INIT('hcdef)
	) name13472 (
		_w8905_,
		_w8908_,
		_w15371_,
		_w15372_,
		_w15373_
	);
	LUT3 #(
		.INIT('h2a)
	) name13473 (
		\m1_data_i[17]_pad ,
		_w8910_,
		_w8911_,
		_w15374_
	);
	LUT3 #(
		.INIT('h80)
	) name13474 (
		\m4_data_i[17]_pad ,
		_w8910_,
		_w8911_,
		_w15375_
	);
	LUT4 #(
		.INIT('h5d7f)
	) name13475 (
		_w8905_,
		_w8908_,
		_w15374_,
		_w15375_,
		_w15376_
	);
	LUT3 #(
		.INIT('h80)
	) name13476 (
		\m2_data_i[17]_pad ,
		_w8910_,
		_w8911_,
		_w15377_
	);
	LUT3 #(
		.INIT('h2a)
	) name13477 (
		\m3_data_i[17]_pad ,
		_w8910_,
		_w8911_,
		_w15378_
	);
	LUT3 #(
		.INIT('h57)
	) name13478 (
		_w8909_,
		_w15377_,
		_w15378_,
		_w15379_
	);
	LUT3 #(
		.INIT('h80)
	) name13479 (
		\m0_data_i[17]_pad ,
		_w8910_,
		_w8911_,
		_w15380_
	);
	LUT3 #(
		.INIT('h2a)
	) name13480 (
		\m7_data_i[17]_pad ,
		_w8910_,
		_w8911_,
		_w15381_
	);
	LUT4 #(
		.INIT('h6e7f)
	) name13481 (
		_w8905_,
		_w8908_,
		_w15380_,
		_w15381_,
		_w15382_
	);
	LUT4 #(
		.INIT('h7fff)
	) name13482 (
		_w15373_,
		_w15376_,
		_w15379_,
		_w15382_,
		_w15383_
	);
	LUT3 #(
		.INIT('h80)
	) name13483 (
		\m0_data_i[18]_pad ,
		_w8910_,
		_w8911_,
		_w15384_
	);
	LUT3 #(
		.INIT('h2a)
	) name13484 (
		\m7_data_i[18]_pad ,
		_w8910_,
		_w8911_,
		_w15385_
	);
	LUT4 #(
		.INIT('h6e7f)
	) name13485 (
		_w8905_,
		_w8908_,
		_w15384_,
		_w15385_,
		_w15386_
	);
	LUT3 #(
		.INIT('h2a)
	) name13486 (
		\m1_data_i[18]_pad ,
		_w8910_,
		_w8911_,
		_w15387_
	);
	LUT3 #(
		.INIT('h80)
	) name13487 (
		\m4_data_i[18]_pad ,
		_w8910_,
		_w8911_,
		_w15388_
	);
	LUT4 #(
		.INIT('h5d7f)
	) name13488 (
		_w8905_,
		_w8908_,
		_w15387_,
		_w15388_,
		_w15389_
	);
	LUT3 #(
		.INIT('h80)
	) name13489 (
		\m2_data_i[18]_pad ,
		_w8910_,
		_w8911_,
		_w15390_
	);
	LUT3 #(
		.INIT('h2a)
	) name13490 (
		\m3_data_i[18]_pad ,
		_w8910_,
		_w8911_,
		_w15391_
	);
	LUT3 #(
		.INIT('h57)
	) name13491 (
		_w8909_,
		_w15390_,
		_w15391_,
		_w15392_
	);
	LUT3 #(
		.INIT('h80)
	) name13492 (
		\m6_data_i[18]_pad ,
		_w8910_,
		_w8911_,
		_w15393_
	);
	LUT3 #(
		.INIT('h2a)
	) name13493 (
		\m5_data_i[18]_pad ,
		_w8910_,
		_w8911_,
		_w15394_
	);
	LUT4 #(
		.INIT('hcdef)
	) name13494 (
		_w8905_,
		_w8908_,
		_w15393_,
		_w15394_,
		_w15395_
	);
	LUT4 #(
		.INIT('h7fff)
	) name13495 (
		_w15386_,
		_w15389_,
		_w15392_,
		_w15395_,
		_w15396_
	);
	LUT3 #(
		.INIT('h2a)
	) name13496 (
		\m1_data_i[19]_pad ,
		_w8910_,
		_w8911_,
		_w15397_
	);
	LUT3 #(
		.INIT('h80)
	) name13497 (
		\m2_data_i[19]_pad ,
		_w8910_,
		_w8911_,
		_w15398_
	);
	LUT4 #(
		.INIT('h3b7f)
	) name13498 (
		_w8905_,
		_w8908_,
		_w15397_,
		_w15398_,
		_w15399_
	);
	LUT3 #(
		.INIT('h80)
	) name13499 (
		\m6_data_i[19]_pad ,
		_w8910_,
		_w8911_,
		_w15400_
	);
	LUT3 #(
		.INIT('h80)
	) name13500 (
		\m4_data_i[19]_pad ,
		_w8910_,
		_w8911_,
		_w15401_
	);
	LUT4 #(
		.INIT('hcdef)
	) name13501 (
		_w8905_,
		_w8908_,
		_w15400_,
		_w15401_,
		_w15402_
	);
	LUT3 #(
		.INIT('h2a)
	) name13502 (
		\m5_data_i[19]_pad ,
		_w8910_,
		_w8911_,
		_w15403_
	);
	LUT3 #(
		.INIT('h2a)
	) name13503 (
		\m3_data_i[19]_pad ,
		_w8910_,
		_w8911_,
		_w15404_
	);
	LUT4 #(
		.INIT('h9bdf)
	) name13504 (
		_w8905_,
		_w8908_,
		_w15403_,
		_w15404_,
		_w15405_
	);
	LUT3 #(
		.INIT('h80)
	) name13505 (
		\m0_data_i[19]_pad ,
		_w8910_,
		_w8911_,
		_w15406_
	);
	LUT3 #(
		.INIT('h2a)
	) name13506 (
		\m7_data_i[19]_pad ,
		_w8910_,
		_w8911_,
		_w15407_
	);
	LUT4 #(
		.INIT('h6e7f)
	) name13507 (
		_w8905_,
		_w8908_,
		_w15406_,
		_w15407_,
		_w15408_
	);
	LUT4 #(
		.INIT('h7fff)
	) name13508 (
		_w15399_,
		_w15402_,
		_w15405_,
		_w15408_,
		_w15409_
	);
	LUT3 #(
		.INIT('h2a)
	) name13509 (
		\m3_data_i[1]_pad ,
		_w8910_,
		_w8911_,
		_w15410_
	);
	LUT3 #(
		.INIT('h80)
	) name13510 (
		\m4_data_i[1]_pad ,
		_w8910_,
		_w8911_,
		_w15411_
	);
	LUT4 #(
		.INIT('h9dbf)
	) name13511 (
		_w8905_,
		_w8908_,
		_w15410_,
		_w15411_,
		_w15412_
	);
	LUT3 #(
		.INIT('h2a)
	) name13512 (
		\m1_data_i[1]_pad ,
		_w8910_,
		_w8911_,
		_w15413_
	);
	LUT3 #(
		.INIT('h2a)
	) name13513 (
		\m5_data_i[1]_pad ,
		_w8910_,
		_w8911_,
		_w15414_
	);
	LUT4 #(
		.INIT('h5d7f)
	) name13514 (
		_w8905_,
		_w8908_,
		_w15413_,
		_w15414_,
		_w15415_
	);
	LUT3 #(
		.INIT('h80)
	) name13515 (
		\m2_data_i[1]_pad ,
		_w8910_,
		_w8911_,
		_w15416_
	);
	LUT3 #(
		.INIT('h80)
	) name13516 (
		\m6_data_i[1]_pad ,
		_w8910_,
		_w8911_,
		_w15417_
	);
	LUT4 #(
		.INIT('haebf)
	) name13517 (
		_w8905_,
		_w8908_,
		_w15416_,
		_w15417_,
		_w15418_
	);
	LUT3 #(
		.INIT('h80)
	) name13518 (
		\m0_data_i[1]_pad ,
		_w8910_,
		_w8911_,
		_w15419_
	);
	LUT3 #(
		.INIT('h2a)
	) name13519 (
		\m7_data_i[1]_pad ,
		_w8910_,
		_w8911_,
		_w15420_
	);
	LUT4 #(
		.INIT('h6e7f)
	) name13520 (
		_w8905_,
		_w8908_,
		_w15419_,
		_w15420_,
		_w15421_
	);
	LUT4 #(
		.INIT('h7fff)
	) name13521 (
		_w15412_,
		_w15415_,
		_w15418_,
		_w15421_,
		_w15422_
	);
	LUT3 #(
		.INIT('h80)
	) name13522 (
		\m0_data_i[20]_pad ,
		_w8910_,
		_w8911_,
		_w15423_
	);
	LUT3 #(
		.INIT('h2a)
	) name13523 (
		\m7_data_i[20]_pad ,
		_w8910_,
		_w8911_,
		_w15424_
	);
	LUT4 #(
		.INIT('h6e7f)
	) name13524 (
		_w8905_,
		_w8908_,
		_w15423_,
		_w15424_,
		_w15425_
	);
	LUT3 #(
		.INIT('h2a)
	) name13525 (
		\m1_data_i[20]_pad ,
		_w8910_,
		_w8911_,
		_w15426_
	);
	LUT3 #(
		.INIT('h80)
	) name13526 (
		\m4_data_i[20]_pad ,
		_w8910_,
		_w8911_,
		_w15427_
	);
	LUT4 #(
		.INIT('h5d7f)
	) name13527 (
		_w8905_,
		_w8908_,
		_w15426_,
		_w15427_,
		_w15428_
	);
	LUT3 #(
		.INIT('h80)
	) name13528 (
		\m2_data_i[20]_pad ,
		_w8910_,
		_w8911_,
		_w15429_
	);
	LUT3 #(
		.INIT('h2a)
	) name13529 (
		\m3_data_i[20]_pad ,
		_w8910_,
		_w8911_,
		_w15430_
	);
	LUT3 #(
		.INIT('h57)
	) name13530 (
		_w8909_,
		_w15429_,
		_w15430_,
		_w15431_
	);
	LUT3 #(
		.INIT('h80)
	) name13531 (
		\m6_data_i[20]_pad ,
		_w8910_,
		_w8911_,
		_w15432_
	);
	LUT3 #(
		.INIT('h2a)
	) name13532 (
		\m5_data_i[20]_pad ,
		_w8910_,
		_w8911_,
		_w15433_
	);
	LUT4 #(
		.INIT('hcdef)
	) name13533 (
		_w8905_,
		_w8908_,
		_w15432_,
		_w15433_,
		_w15434_
	);
	LUT4 #(
		.INIT('h7fff)
	) name13534 (
		_w15425_,
		_w15428_,
		_w15431_,
		_w15434_,
		_w15435_
	);
	LUT3 #(
		.INIT('h2a)
	) name13535 (
		\m1_data_i[21]_pad ,
		_w8910_,
		_w8911_,
		_w15436_
	);
	LUT3 #(
		.INIT('h80)
	) name13536 (
		\m2_data_i[21]_pad ,
		_w8910_,
		_w8911_,
		_w15437_
	);
	LUT4 #(
		.INIT('h3b7f)
	) name13537 (
		_w8905_,
		_w8908_,
		_w15436_,
		_w15437_,
		_w15438_
	);
	LUT3 #(
		.INIT('h80)
	) name13538 (
		\m0_data_i[21]_pad ,
		_w8910_,
		_w8911_,
		_w15439_
	);
	LUT3 #(
		.INIT('h80)
	) name13539 (
		\m4_data_i[21]_pad ,
		_w8910_,
		_w8911_,
		_w15440_
	);
	LUT4 #(
		.INIT('h5d7f)
	) name13540 (
		_w8905_,
		_w8908_,
		_w15439_,
		_w15440_,
		_w15441_
	);
	LUT3 #(
		.INIT('h2a)
	) name13541 (
		\m7_data_i[21]_pad ,
		_w8910_,
		_w8911_,
		_w15442_
	);
	LUT3 #(
		.INIT('h2a)
	) name13542 (
		\m3_data_i[21]_pad ,
		_w8910_,
		_w8911_,
		_w15443_
	);
	LUT4 #(
		.INIT('habef)
	) name13543 (
		_w8905_,
		_w8908_,
		_w15442_,
		_w15443_,
		_w15444_
	);
	LUT3 #(
		.INIT('h80)
	) name13544 (
		\m6_data_i[21]_pad ,
		_w8910_,
		_w8911_,
		_w15445_
	);
	LUT3 #(
		.INIT('h2a)
	) name13545 (
		\m5_data_i[21]_pad ,
		_w8910_,
		_w8911_,
		_w15446_
	);
	LUT4 #(
		.INIT('hcdef)
	) name13546 (
		_w8905_,
		_w8908_,
		_w15445_,
		_w15446_,
		_w15447_
	);
	LUT4 #(
		.INIT('h7fff)
	) name13547 (
		_w15438_,
		_w15441_,
		_w15444_,
		_w15447_,
		_w15448_
	);
	LUT3 #(
		.INIT('h80)
	) name13548 (
		\m6_data_i[22]_pad ,
		_w8910_,
		_w8911_,
		_w15449_
	);
	LUT3 #(
		.INIT('h2a)
	) name13549 (
		\m5_data_i[22]_pad ,
		_w8910_,
		_w8911_,
		_w15450_
	);
	LUT4 #(
		.INIT('hcdef)
	) name13550 (
		_w8905_,
		_w8908_,
		_w15449_,
		_w15450_,
		_w15451_
	);
	LUT3 #(
		.INIT('h2a)
	) name13551 (
		\m3_data_i[22]_pad ,
		_w8910_,
		_w8911_,
		_w15452_
	);
	LUT3 #(
		.INIT('h2a)
	) name13552 (
		\m7_data_i[22]_pad ,
		_w8910_,
		_w8911_,
		_w15453_
	);
	LUT4 #(
		.INIT('haebf)
	) name13553 (
		_w8905_,
		_w8908_,
		_w15452_,
		_w15453_,
		_w15454_
	);
	LUT3 #(
		.INIT('h80)
	) name13554 (
		\m4_data_i[22]_pad ,
		_w8910_,
		_w8911_,
		_w15455_
	);
	LUT3 #(
		.INIT('h80)
	) name13555 (
		\m0_data_i[22]_pad ,
		_w8910_,
		_w8911_,
		_w15456_
	);
	LUT4 #(
		.INIT('h57df)
	) name13556 (
		_w8905_,
		_w8908_,
		_w15455_,
		_w15456_,
		_w15457_
	);
	LUT3 #(
		.INIT('h2a)
	) name13557 (
		\m1_data_i[22]_pad ,
		_w8910_,
		_w8911_,
		_w15458_
	);
	LUT3 #(
		.INIT('h80)
	) name13558 (
		\m2_data_i[22]_pad ,
		_w8910_,
		_w8911_,
		_w15459_
	);
	LUT4 #(
		.INIT('h3b7f)
	) name13559 (
		_w8905_,
		_w8908_,
		_w15458_,
		_w15459_,
		_w15460_
	);
	LUT4 #(
		.INIT('h7fff)
	) name13560 (
		_w15451_,
		_w15454_,
		_w15457_,
		_w15460_,
		_w15461_
	);
	LUT3 #(
		.INIT('h2a)
	) name13561 (
		\m1_data_i[23]_pad ,
		_w8910_,
		_w8911_,
		_w15462_
	);
	LUT3 #(
		.INIT('h80)
	) name13562 (
		\m2_data_i[23]_pad ,
		_w8910_,
		_w8911_,
		_w15463_
	);
	LUT4 #(
		.INIT('h3b7f)
	) name13563 (
		_w8905_,
		_w8908_,
		_w15462_,
		_w15463_,
		_w15464_
	);
	LUT3 #(
		.INIT('h80)
	) name13564 (
		\m0_data_i[23]_pad ,
		_w8910_,
		_w8911_,
		_w15465_
	);
	LUT3 #(
		.INIT('h80)
	) name13565 (
		\m4_data_i[23]_pad ,
		_w8910_,
		_w8911_,
		_w15466_
	);
	LUT4 #(
		.INIT('h5d7f)
	) name13566 (
		_w8905_,
		_w8908_,
		_w15465_,
		_w15466_,
		_w15467_
	);
	LUT3 #(
		.INIT('h2a)
	) name13567 (
		\m7_data_i[23]_pad ,
		_w8910_,
		_w8911_,
		_w15468_
	);
	LUT3 #(
		.INIT('h2a)
	) name13568 (
		\m3_data_i[23]_pad ,
		_w8910_,
		_w8911_,
		_w15469_
	);
	LUT4 #(
		.INIT('habef)
	) name13569 (
		_w8905_,
		_w8908_,
		_w15468_,
		_w15469_,
		_w15470_
	);
	LUT3 #(
		.INIT('h80)
	) name13570 (
		\m6_data_i[23]_pad ,
		_w8910_,
		_w8911_,
		_w15471_
	);
	LUT3 #(
		.INIT('h2a)
	) name13571 (
		\m5_data_i[23]_pad ,
		_w8910_,
		_w8911_,
		_w15472_
	);
	LUT4 #(
		.INIT('hcdef)
	) name13572 (
		_w8905_,
		_w8908_,
		_w15471_,
		_w15472_,
		_w15473_
	);
	LUT4 #(
		.INIT('h7fff)
	) name13573 (
		_w15464_,
		_w15467_,
		_w15470_,
		_w15473_,
		_w15474_
	);
	LUT3 #(
		.INIT('h2a)
	) name13574 (
		\m3_data_i[24]_pad ,
		_w8910_,
		_w8911_,
		_w15475_
	);
	LUT3 #(
		.INIT('h80)
	) name13575 (
		\m4_data_i[24]_pad ,
		_w8910_,
		_w8911_,
		_w15476_
	);
	LUT4 #(
		.INIT('h9dbf)
	) name13576 (
		_w8905_,
		_w8908_,
		_w15475_,
		_w15476_,
		_w15477_
	);
	LUT3 #(
		.INIT('h2a)
	) name13577 (
		\m1_data_i[24]_pad ,
		_w8910_,
		_w8911_,
		_w15478_
	);
	LUT3 #(
		.INIT('h2a)
	) name13578 (
		\m5_data_i[24]_pad ,
		_w8910_,
		_w8911_,
		_w15479_
	);
	LUT4 #(
		.INIT('h5d7f)
	) name13579 (
		_w8905_,
		_w8908_,
		_w15478_,
		_w15479_,
		_w15480_
	);
	LUT3 #(
		.INIT('h80)
	) name13580 (
		\m2_data_i[24]_pad ,
		_w8910_,
		_w8911_,
		_w15481_
	);
	LUT3 #(
		.INIT('h80)
	) name13581 (
		\m6_data_i[24]_pad ,
		_w8910_,
		_w8911_,
		_w15482_
	);
	LUT4 #(
		.INIT('haebf)
	) name13582 (
		_w8905_,
		_w8908_,
		_w15481_,
		_w15482_,
		_w15483_
	);
	LUT3 #(
		.INIT('h80)
	) name13583 (
		\m0_data_i[24]_pad ,
		_w8910_,
		_w8911_,
		_w15484_
	);
	LUT3 #(
		.INIT('h2a)
	) name13584 (
		\m7_data_i[24]_pad ,
		_w8910_,
		_w8911_,
		_w15485_
	);
	LUT4 #(
		.INIT('h6e7f)
	) name13585 (
		_w8905_,
		_w8908_,
		_w15484_,
		_w15485_,
		_w15486_
	);
	LUT4 #(
		.INIT('h7fff)
	) name13586 (
		_w15477_,
		_w15480_,
		_w15483_,
		_w15486_,
		_w15487_
	);
	LUT3 #(
		.INIT('h2a)
	) name13587 (
		\m3_data_i[25]_pad ,
		_w8910_,
		_w8911_,
		_w15488_
	);
	LUT3 #(
		.INIT('h80)
	) name13588 (
		\m4_data_i[25]_pad ,
		_w8910_,
		_w8911_,
		_w15489_
	);
	LUT4 #(
		.INIT('h9dbf)
	) name13589 (
		_w8905_,
		_w8908_,
		_w15488_,
		_w15489_,
		_w15490_
	);
	LUT3 #(
		.INIT('h80)
	) name13590 (
		\m0_data_i[25]_pad ,
		_w8910_,
		_w8911_,
		_w15491_
	);
	LUT3 #(
		.INIT('h80)
	) name13591 (
		\m2_data_i[25]_pad ,
		_w8910_,
		_w8911_,
		_w15492_
	);
	LUT4 #(
		.INIT('h3b7f)
	) name13592 (
		_w8905_,
		_w8908_,
		_w15491_,
		_w15492_,
		_w15493_
	);
	LUT3 #(
		.INIT('h2a)
	) name13593 (
		\m7_data_i[25]_pad ,
		_w8910_,
		_w8911_,
		_w15494_
	);
	LUT3 #(
		.INIT('h2a)
	) name13594 (
		\m1_data_i[25]_pad ,
		_w8910_,
		_w8911_,
		_w15495_
	);
	LUT4 #(
		.INIT('h67ef)
	) name13595 (
		_w8905_,
		_w8908_,
		_w15494_,
		_w15495_,
		_w15496_
	);
	LUT3 #(
		.INIT('h80)
	) name13596 (
		\m6_data_i[25]_pad ,
		_w8910_,
		_w8911_,
		_w15497_
	);
	LUT3 #(
		.INIT('h2a)
	) name13597 (
		\m5_data_i[25]_pad ,
		_w8910_,
		_w8911_,
		_w15498_
	);
	LUT4 #(
		.INIT('hcdef)
	) name13598 (
		_w8905_,
		_w8908_,
		_w15497_,
		_w15498_,
		_w15499_
	);
	LUT4 #(
		.INIT('h7fff)
	) name13599 (
		_w15490_,
		_w15493_,
		_w15496_,
		_w15499_,
		_w15500_
	);
	LUT3 #(
		.INIT('h2a)
	) name13600 (
		\m3_data_i[26]_pad ,
		_w8910_,
		_w8911_,
		_w15501_
	);
	LUT3 #(
		.INIT('h80)
	) name13601 (
		\m4_data_i[26]_pad ,
		_w8910_,
		_w8911_,
		_w15502_
	);
	LUT4 #(
		.INIT('h9dbf)
	) name13602 (
		_w8905_,
		_w8908_,
		_w15501_,
		_w15502_,
		_w15503_
	);
	LUT3 #(
		.INIT('h80)
	) name13603 (
		\m0_data_i[26]_pad ,
		_w8910_,
		_w8911_,
		_w15504_
	);
	LUT3 #(
		.INIT('h2a)
	) name13604 (
		\m5_data_i[26]_pad ,
		_w8910_,
		_w8911_,
		_w15505_
	);
	LUT4 #(
		.INIT('h5d7f)
	) name13605 (
		_w8905_,
		_w8908_,
		_w15504_,
		_w15505_,
		_w15506_
	);
	LUT3 #(
		.INIT('h2a)
	) name13606 (
		\m7_data_i[26]_pad ,
		_w8910_,
		_w8911_,
		_w15507_
	);
	LUT3 #(
		.INIT('h80)
	) name13607 (
		\m6_data_i[26]_pad ,
		_w8910_,
		_w8911_,
		_w15508_
	);
	LUT3 #(
		.INIT('h57)
	) name13608 (
		_w8917_,
		_w15507_,
		_w15508_,
		_w15509_
	);
	LUT3 #(
		.INIT('h2a)
	) name13609 (
		\m1_data_i[26]_pad ,
		_w8910_,
		_w8911_,
		_w15510_
	);
	LUT3 #(
		.INIT('h80)
	) name13610 (
		\m2_data_i[26]_pad ,
		_w8910_,
		_w8911_,
		_w15511_
	);
	LUT4 #(
		.INIT('h3b7f)
	) name13611 (
		_w8905_,
		_w8908_,
		_w15510_,
		_w15511_,
		_w15512_
	);
	LUT4 #(
		.INIT('h7fff)
	) name13612 (
		_w15503_,
		_w15506_,
		_w15509_,
		_w15512_,
		_w15513_
	);
	LUT3 #(
		.INIT('h2a)
	) name13613 (
		\m1_data_i[27]_pad ,
		_w8910_,
		_w8911_,
		_w15514_
	);
	LUT3 #(
		.INIT('h80)
	) name13614 (
		\m2_data_i[27]_pad ,
		_w8910_,
		_w8911_,
		_w15515_
	);
	LUT4 #(
		.INIT('h3b7f)
	) name13615 (
		_w8905_,
		_w8908_,
		_w15514_,
		_w15515_,
		_w15516_
	);
	LUT3 #(
		.INIT('h80)
	) name13616 (
		\m0_data_i[27]_pad ,
		_w8910_,
		_w8911_,
		_w15517_
	);
	LUT3 #(
		.INIT('h80)
	) name13617 (
		\m4_data_i[27]_pad ,
		_w8910_,
		_w8911_,
		_w15518_
	);
	LUT4 #(
		.INIT('h5d7f)
	) name13618 (
		_w8905_,
		_w8908_,
		_w15517_,
		_w15518_,
		_w15519_
	);
	LUT3 #(
		.INIT('h2a)
	) name13619 (
		\m7_data_i[27]_pad ,
		_w8910_,
		_w8911_,
		_w15520_
	);
	LUT3 #(
		.INIT('h2a)
	) name13620 (
		\m3_data_i[27]_pad ,
		_w8910_,
		_w8911_,
		_w15521_
	);
	LUT4 #(
		.INIT('habef)
	) name13621 (
		_w8905_,
		_w8908_,
		_w15520_,
		_w15521_,
		_w15522_
	);
	LUT3 #(
		.INIT('h80)
	) name13622 (
		\m6_data_i[27]_pad ,
		_w8910_,
		_w8911_,
		_w15523_
	);
	LUT3 #(
		.INIT('h2a)
	) name13623 (
		\m5_data_i[27]_pad ,
		_w8910_,
		_w8911_,
		_w15524_
	);
	LUT4 #(
		.INIT('hcdef)
	) name13624 (
		_w8905_,
		_w8908_,
		_w15523_,
		_w15524_,
		_w15525_
	);
	LUT4 #(
		.INIT('h7fff)
	) name13625 (
		_w15516_,
		_w15519_,
		_w15522_,
		_w15525_,
		_w15526_
	);
	LUT3 #(
		.INIT('h2a)
	) name13626 (
		\m3_data_i[28]_pad ,
		_w8910_,
		_w8911_,
		_w15527_
	);
	LUT3 #(
		.INIT('h80)
	) name13627 (
		\m4_data_i[28]_pad ,
		_w8910_,
		_w8911_,
		_w15528_
	);
	LUT4 #(
		.INIT('h9dbf)
	) name13628 (
		_w8905_,
		_w8908_,
		_w15527_,
		_w15528_,
		_w15529_
	);
	LUT3 #(
		.INIT('h80)
	) name13629 (
		\m6_data_i[28]_pad ,
		_w8910_,
		_w8911_,
		_w15530_
	);
	LUT3 #(
		.INIT('h2a)
	) name13630 (
		\m7_data_i[28]_pad ,
		_w8910_,
		_w8911_,
		_w15531_
	);
	LUT3 #(
		.INIT('h57)
	) name13631 (
		_w8917_,
		_w15530_,
		_w15531_,
		_w15532_
	);
	LUT3 #(
		.INIT('h2a)
	) name13632 (
		\m5_data_i[28]_pad ,
		_w8910_,
		_w8911_,
		_w15533_
	);
	LUT3 #(
		.INIT('h80)
	) name13633 (
		\m0_data_i[28]_pad ,
		_w8910_,
		_w8911_,
		_w15534_
	);
	LUT4 #(
		.INIT('h57df)
	) name13634 (
		_w8905_,
		_w8908_,
		_w15533_,
		_w15534_,
		_w15535_
	);
	LUT3 #(
		.INIT('h2a)
	) name13635 (
		\m1_data_i[28]_pad ,
		_w8910_,
		_w8911_,
		_w15536_
	);
	LUT3 #(
		.INIT('h80)
	) name13636 (
		\m2_data_i[28]_pad ,
		_w8910_,
		_w8911_,
		_w15537_
	);
	LUT4 #(
		.INIT('h3b7f)
	) name13637 (
		_w8905_,
		_w8908_,
		_w15536_,
		_w15537_,
		_w15538_
	);
	LUT4 #(
		.INIT('h7fff)
	) name13638 (
		_w15529_,
		_w15532_,
		_w15535_,
		_w15538_,
		_w15539_
	);
	LUT3 #(
		.INIT('h2a)
	) name13639 (
		\m1_data_i[29]_pad ,
		_w8910_,
		_w8911_,
		_w15540_
	);
	LUT3 #(
		.INIT('h80)
	) name13640 (
		\m2_data_i[29]_pad ,
		_w8910_,
		_w8911_,
		_w15541_
	);
	LUT4 #(
		.INIT('h3b7f)
	) name13641 (
		_w8905_,
		_w8908_,
		_w15540_,
		_w15541_,
		_w15542_
	);
	LUT3 #(
		.INIT('h80)
	) name13642 (
		\m0_data_i[29]_pad ,
		_w8910_,
		_w8911_,
		_w15543_
	);
	LUT3 #(
		.INIT('h80)
	) name13643 (
		\m4_data_i[29]_pad ,
		_w8910_,
		_w8911_,
		_w15544_
	);
	LUT4 #(
		.INIT('h5d7f)
	) name13644 (
		_w8905_,
		_w8908_,
		_w15543_,
		_w15544_,
		_w15545_
	);
	LUT3 #(
		.INIT('h2a)
	) name13645 (
		\m7_data_i[29]_pad ,
		_w8910_,
		_w8911_,
		_w15546_
	);
	LUT3 #(
		.INIT('h2a)
	) name13646 (
		\m3_data_i[29]_pad ,
		_w8910_,
		_w8911_,
		_w15547_
	);
	LUT4 #(
		.INIT('habef)
	) name13647 (
		_w8905_,
		_w8908_,
		_w15546_,
		_w15547_,
		_w15548_
	);
	LUT3 #(
		.INIT('h80)
	) name13648 (
		\m6_data_i[29]_pad ,
		_w8910_,
		_w8911_,
		_w15549_
	);
	LUT3 #(
		.INIT('h2a)
	) name13649 (
		\m5_data_i[29]_pad ,
		_w8910_,
		_w8911_,
		_w15550_
	);
	LUT4 #(
		.INIT('hcdef)
	) name13650 (
		_w8905_,
		_w8908_,
		_w15549_,
		_w15550_,
		_w15551_
	);
	LUT4 #(
		.INIT('h7fff)
	) name13651 (
		_w15542_,
		_w15545_,
		_w15548_,
		_w15551_,
		_w15552_
	);
	LUT3 #(
		.INIT('h2a)
	) name13652 (
		\m3_data_i[2]_pad ,
		_w8910_,
		_w8911_,
		_w15553_
	);
	LUT3 #(
		.INIT('h80)
	) name13653 (
		\m4_data_i[2]_pad ,
		_w8910_,
		_w8911_,
		_w15554_
	);
	LUT4 #(
		.INIT('h9dbf)
	) name13654 (
		_w8905_,
		_w8908_,
		_w15553_,
		_w15554_,
		_w15555_
	);
	LUT3 #(
		.INIT('h80)
	) name13655 (
		\m0_data_i[2]_pad ,
		_w8910_,
		_w8911_,
		_w15556_
	);
	LUT3 #(
		.INIT('h2a)
	) name13656 (
		\m5_data_i[2]_pad ,
		_w8910_,
		_w8911_,
		_w15557_
	);
	LUT4 #(
		.INIT('h5d7f)
	) name13657 (
		_w8905_,
		_w8908_,
		_w15556_,
		_w15557_,
		_w15558_
	);
	LUT3 #(
		.INIT('h2a)
	) name13658 (
		\m7_data_i[2]_pad ,
		_w8910_,
		_w8911_,
		_w15559_
	);
	LUT3 #(
		.INIT('h80)
	) name13659 (
		\m6_data_i[2]_pad ,
		_w8910_,
		_w8911_,
		_w15560_
	);
	LUT3 #(
		.INIT('h57)
	) name13660 (
		_w8917_,
		_w15559_,
		_w15560_,
		_w15561_
	);
	LUT3 #(
		.INIT('h2a)
	) name13661 (
		\m1_data_i[2]_pad ,
		_w8910_,
		_w8911_,
		_w15562_
	);
	LUT3 #(
		.INIT('h80)
	) name13662 (
		\m2_data_i[2]_pad ,
		_w8910_,
		_w8911_,
		_w15563_
	);
	LUT4 #(
		.INIT('h3b7f)
	) name13663 (
		_w8905_,
		_w8908_,
		_w15562_,
		_w15563_,
		_w15564_
	);
	LUT4 #(
		.INIT('h7fff)
	) name13664 (
		_w15555_,
		_w15558_,
		_w15561_,
		_w15564_,
		_w15565_
	);
	LUT3 #(
		.INIT('h2a)
	) name13665 (
		\m3_data_i[30]_pad ,
		_w8910_,
		_w8911_,
		_w15566_
	);
	LUT3 #(
		.INIT('h80)
	) name13666 (
		\m4_data_i[30]_pad ,
		_w8910_,
		_w8911_,
		_w15567_
	);
	LUT4 #(
		.INIT('h9dbf)
	) name13667 (
		_w8905_,
		_w8908_,
		_w15566_,
		_w15567_,
		_w15568_
	);
	LUT3 #(
		.INIT('h80)
	) name13668 (
		\m6_data_i[30]_pad ,
		_w8910_,
		_w8911_,
		_w15569_
	);
	LUT3 #(
		.INIT('h2a)
	) name13669 (
		\m7_data_i[30]_pad ,
		_w8910_,
		_w8911_,
		_w15570_
	);
	LUT3 #(
		.INIT('h57)
	) name13670 (
		_w8917_,
		_w15569_,
		_w15570_,
		_w15571_
	);
	LUT3 #(
		.INIT('h2a)
	) name13671 (
		\m5_data_i[30]_pad ,
		_w8910_,
		_w8911_,
		_w15572_
	);
	LUT3 #(
		.INIT('h80)
	) name13672 (
		\m0_data_i[30]_pad ,
		_w8910_,
		_w8911_,
		_w15573_
	);
	LUT4 #(
		.INIT('h57df)
	) name13673 (
		_w8905_,
		_w8908_,
		_w15572_,
		_w15573_,
		_w15574_
	);
	LUT3 #(
		.INIT('h2a)
	) name13674 (
		\m1_data_i[30]_pad ,
		_w8910_,
		_w8911_,
		_w15575_
	);
	LUT3 #(
		.INIT('h80)
	) name13675 (
		\m2_data_i[30]_pad ,
		_w8910_,
		_w8911_,
		_w15576_
	);
	LUT4 #(
		.INIT('h3b7f)
	) name13676 (
		_w8905_,
		_w8908_,
		_w15575_,
		_w15576_,
		_w15577_
	);
	LUT4 #(
		.INIT('h7fff)
	) name13677 (
		_w15568_,
		_w15571_,
		_w15574_,
		_w15577_,
		_w15578_
	);
	LUT3 #(
		.INIT('h2a)
	) name13678 (
		\m1_data_i[31]_pad ,
		_w8910_,
		_w8911_,
		_w15579_
	);
	LUT3 #(
		.INIT('h80)
	) name13679 (
		\m2_data_i[31]_pad ,
		_w8910_,
		_w8911_,
		_w15580_
	);
	LUT4 #(
		.INIT('h3b7f)
	) name13680 (
		_w8905_,
		_w8908_,
		_w15579_,
		_w15580_,
		_w15581_
	);
	LUT3 #(
		.INIT('h2a)
	) name13681 (
		\m3_data_i[31]_pad ,
		_w8910_,
		_w8911_,
		_w15582_
	);
	LUT3 #(
		.INIT('h2a)
	) name13682 (
		\m7_data_i[31]_pad ,
		_w8910_,
		_w8911_,
		_w15583_
	);
	LUT4 #(
		.INIT('haebf)
	) name13683 (
		_w8905_,
		_w8908_,
		_w15582_,
		_w15583_,
		_w15584_
	);
	LUT3 #(
		.INIT('h80)
	) name13684 (
		\m4_data_i[31]_pad ,
		_w8910_,
		_w8911_,
		_w15585_
	);
	LUT3 #(
		.INIT('h80)
	) name13685 (
		\m0_data_i[31]_pad ,
		_w8910_,
		_w8911_,
		_w15586_
	);
	LUT4 #(
		.INIT('h57df)
	) name13686 (
		_w8905_,
		_w8908_,
		_w15585_,
		_w15586_,
		_w15587_
	);
	LUT3 #(
		.INIT('h80)
	) name13687 (
		\m6_data_i[31]_pad ,
		_w8910_,
		_w8911_,
		_w15588_
	);
	LUT3 #(
		.INIT('h2a)
	) name13688 (
		\m5_data_i[31]_pad ,
		_w8910_,
		_w8911_,
		_w15589_
	);
	LUT4 #(
		.INIT('hcdef)
	) name13689 (
		_w8905_,
		_w8908_,
		_w15588_,
		_w15589_,
		_w15590_
	);
	LUT4 #(
		.INIT('h7fff)
	) name13690 (
		_w15581_,
		_w15584_,
		_w15587_,
		_w15590_,
		_w15591_
	);
	LUT3 #(
		.INIT('h80)
	) name13691 (
		\m0_data_i[3]_pad ,
		_w8910_,
		_w8911_,
		_w15592_
	);
	LUT3 #(
		.INIT('h2a)
	) name13692 (
		\m7_data_i[3]_pad ,
		_w8910_,
		_w8911_,
		_w15593_
	);
	LUT4 #(
		.INIT('h6e7f)
	) name13693 (
		_w8905_,
		_w8908_,
		_w15592_,
		_w15593_,
		_w15594_
	);
	LUT3 #(
		.INIT('h2a)
	) name13694 (
		\m1_data_i[3]_pad ,
		_w8910_,
		_w8911_,
		_w15595_
	);
	LUT3 #(
		.INIT('h2a)
	) name13695 (
		\m5_data_i[3]_pad ,
		_w8910_,
		_w8911_,
		_w15596_
	);
	LUT4 #(
		.INIT('h5d7f)
	) name13696 (
		_w8905_,
		_w8908_,
		_w15595_,
		_w15596_,
		_w15597_
	);
	LUT3 #(
		.INIT('h80)
	) name13697 (
		\m2_data_i[3]_pad ,
		_w8910_,
		_w8911_,
		_w15598_
	);
	LUT3 #(
		.INIT('h80)
	) name13698 (
		\m6_data_i[3]_pad ,
		_w8910_,
		_w8911_,
		_w15599_
	);
	LUT4 #(
		.INIT('haebf)
	) name13699 (
		_w8905_,
		_w8908_,
		_w15598_,
		_w15599_,
		_w15600_
	);
	LUT3 #(
		.INIT('h2a)
	) name13700 (
		\m3_data_i[3]_pad ,
		_w8910_,
		_w8911_,
		_w15601_
	);
	LUT3 #(
		.INIT('h80)
	) name13701 (
		\m4_data_i[3]_pad ,
		_w8910_,
		_w8911_,
		_w15602_
	);
	LUT4 #(
		.INIT('h9dbf)
	) name13702 (
		_w8905_,
		_w8908_,
		_w15601_,
		_w15602_,
		_w15603_
	);
	LUT4 #(
		.INIT('h7fff)
	) name13703 (
		_w15594_,
		_w15597_,
		_w15600_,
		_w15603_,
		_w15604_
	);
	LUT3 #(
		.INIT('h2a)
	) name13704 (
		\m1_data_i[4]_pad ,
		_w8910_,
		_w8911_,
		_w15605_
	);
	LUT3 #(
		.INIT('h80)
	) name13705 (
		\m2_data_i[4]_pad ,
		_w8910_,
		_w8911_,
		_w15606_
	);
	LUT4 #(
		.INIT('h3b7f)
	) name13706 (
		_w8905_,
		_w8908_,
		_w15605_,
		_w15606_,
		_w15607_
	);
	LUT3 #(
		.INIT('h80)
	) name13707 (
		\m0_data_i[4]_pad ,
		_w8910_,
		_w8911_,
		_w15608_
	);
	LUT3 #(
		.INIT('h2a)
	) name13708 (
		\m5_data_i[4]_pad ,
		_w8910_,
		_w8911_,
		_w15609_
	);
	LUT4 #(
		.INIT('h5d7f)
	) name13709 (
		_w8905_,
		_w8908_,
		_w15608_,
		_w15609_,
		_w15610_
	);
	LUT3 #(
		.INIT('h2a)
	) name13710 (
		\m7_data_i[4]_pad ,
		_w8910_,
		_w8911_,
		_w15611_
	);
	LUT3 #(
		.INIT('h80)
	) name13711 (
		\m6_data_i[4]_pad ,
		_w8910_,
		_w8911_,
		_w15612_
	);
	LUT3 #(
		.INIT('h57)
	) name13712 (
		_w8917_,
		_w15611_,
		_w15612_,
		_w15613_
	);
	LUT3 #(
		.INIT('h2a)
	) name13713 (
		\m3_data_i[4]_pad ,
		_w8910_,
		_w8911_,
		_w15614_
	);
	LUT3 #(
		.INIT('h80)
	) name13714 (
		\m4_data_i[4]_pad ,
		_w8910_,
		_w8911_,
		_w15615_
	);
	LUT4 #(
		.INIT('h9dbf)
	) name13715 (
		_w8905_,
		_w8908_,
		_w15614_,
		_w15615_,
		_w15616_
	);
	LUT4 #(
		.INIT('h7fff)
	) name13716 (
		_w15607_,
		_w15610_,
		_w15613_,
		_w15616_,
		_w15617_
	);
	LUT3 #(
		.INIT('h80)
	) name13717 (
		\m6_data_i[5]_pad ,
		_w8910_,
		_w8911_,
		_w15618_
	);
	LUT3 #(
		.INIT('h2a)
	) name13718 (
		\m5_data_i[5]_pad ,
		_w8910_,
		_w8911_,
		_w15619_
	);
	LUT4 #(
		.INIT('hcdef)
	) name13719 (
		_w8905_,
		_w8908_,
		_w15618_,
		_w15619_,
		_w15620_
	);
	LUT3 #(
		.INIT('h2a)
	) name13720 (
		\m1_data_i[5]_pad ,
		_w8910_,
		_w8911_,
		_w15621_
	);
	LUT3 #(
		.INIT('h2a)
	) name13721 (
		\m7_data_i[5]_pad ,
		_w8910_,
		_w8911_,
		_w15622_
	);
	LUT4 #(
		.INIT('h6e7f)
	) name13722 (
		_w8905_,
		_w8908_,
		_w15621_,
		_w15622_,
		_w15623_
	);
	LUT3 #(
		.INIT('h80)
	) name13723 (
		\m2_data_i[5]_pad ,
		_w8910_,
		_w8911_,
		_w15624_
	);
	LUT3 #(
		.INIT('h80)
	) name13724 (
		\m0_data_i[5]_pad ,
		_w8910_,
		_w8911_,
		_w15625_
	);
	LUT4 #(
		.INIT('h37bf)
	) name13725 (
		_w8905_,
		_w8908_,
		_w15624_,
		_w15625_,
		_w15626_
	);
	LUT3 #(
		.INIT('h2a)
	) name13726 (
		\m3_data_i[5]_pad ,
		_w8910_,
		_w8911_,
		_w15627_
	);
	LUT3 #(
		.INIT('h80)
	) name13727 (
		\m4_data_i[5]_pad ,
		_w8910_,
		_w8911_,
		_w15628_
	);
	LUT4 #(
		.INIT('h9dbf)
	) name13728 (
		_w8905_,
		_w8908_,
		_w15627_,
		_w15628_,
		_w15629_
	);
	LUT4 #(
		.INIT('h7fff)
	) name13729 (
		_w15620_,
		_w15623_,
		_w15626_,
		_w15629_,
		_w15630_
	);
	LUT3 #(
		.INIT('h2a)
	) name13730 (
		\m3_data_i[6]_pad ,
		_w8910_,
		_w8911_,
		_w15631_
	);
	LUT3 #(
		.INIT('h80)
	) name13731 (
		\m4_data_i[6]_pad ,
		_w8910_,
		_w8911_,
		_w15632_
	);
	LUT4 #(
		.INIT('h9dbf)
	) name13732 (
		_w8905_,
		_w8908_,
		_w15631_,
		_w15632_,
		_w15633_
	);
	LUT3 #(
		.INIT('h2a)
	) name13733 (
		\m1_data_i[6]_pad ,
		_w8910_,
		_w8911_,
		_w15634_
	);
	LUT3 #(
		.INIT('h2a)
	) name13734 (
		\m5_data_i[6]_pad ,
		_w8910_,
		_w8911_,
		_w15635_
	);
	LUT4 #(
		.INIT('h5d7f)
	) name13735 (
		_w8905_,
		_w8908_,
		_w15634_,
		_w15635_,
		_w15636_
	);
	LUT3 #(
		.INIT('h80)
	) name13736 (
		\m2_data_i[6]_pad ,
		_w8910_,
		_w8911_,
		_w15637_
	);
	LUT3 #(
		.INIT('h80)
	) name13737 (
		\m6_data_i[6]_pad ,
		_w8910_,
		_w8911_,
		_w15638_
	);
	LUT4 #(
		.INIT('haebf)
	) name13738 (
		_w8905_,
		_w8908_,
		_w15637_,
		_w15638_,
		_w15639_
	);
	LUT3 #(
		.INIT('h80)
	) name13739 (
		\m0_data_i[6]_pad ,
		_w8910_,
		_w8911_,
		_w15640_
	);
	LUT3 #(
		.INIT('h2a)
	) name13740 (
		\m7_data_i[6]_pad ,
		_w8910_,
		_w8911_,
		_w15641_
	);
	LUT4 #(
		.INIT('h6e7f)
	) name13741 (
		_w8905_,
		_w8908_,
		_w15640_,
		_w15641_,
		_w15642_
	);
	LUT4 #(
		.INIT('h7fff)
	) name13742 (
		_w15633_,
		_w15636_,
		_w15639_,
		_w15642_,
		_w15643_
	);
	LUT3 #(
		.INIT('h2a)
	) name13743 (
		\m1_data_i[7]_pad ,
		_w8910_,
		_w8911_,
		_w15644_
	);
	LUT3 #(
		.INIT('h80)
	) name13744 (
		\m2_data_i[7]_pad ,
		_w8910_,
		_w8911_,
		_w15645_
	);
	LUT4 #(
		.INIT('h3b7f)
	) name13745 (
		_w8905_,
		_w8908_,
		_w15644_,
		_w15645_,
		_w15646_
	);
	LUT3 #(
		.INIT('h80)
	) name13746 (
		\m0_data_i[7]_pad ,
		_w8910_,
		_w8911_,
		_w15647_
	);
	LUT3 #(
		.INIT('h2a)
	) name13747 (
		\m5_data_i[7]_pad ,
		_w8910_,
		_w8911_,
		_w15648_
	);
	LUT4 #(
		.INIT('h5d7f)
	) name13748 (
		_w8905_,
		_w8908_,
		_w15647_,
		_w15648_,
		_w15649_
	);
	LUT3 #(
		.INIT('h2a)
	) name13749 (
		\m7_data_i[7]_pad ,
		_w8910_,
		_w8911_,
		_w15650_
	);
	LUT3 #(
		.INIT('h80)
	) name13750 (
		\m6_data_i[7]_pad ,
		_w8910_,
		_w8911_,
		_w15651_
	);
	LUT3 #(
		.INIT('h57)
	) name13751 (
		_w8917_,
		_w15650_,
		_w15651_,
		_w15652_
	);
	LUT3 #(
		.INIT('h2a)
	) name13752 (
		\m3_data_i[7]_pad ,
		_w8910_,
		_w8911_,
		_w15653_
	);
	LUT3 #(
		.INIT('h80)
	) name13753 (
		\m4_data_i[7]_pad ,
		_w8910_,
		_w8911_,
		_w15654_
	);
	LUT4 #(
		.INIT('h9dbf)
	) name13754 (
		_w8905_,
		_w8908_,
		_w15653_,
		_w15654_,
		_w15655_
	);
	LUT4 #(
		.INIT('h7fff)
	) name13755 (
		_w15646_,
		_w15649_,
		_w15652_,
		_w15655_,
		_w15656_
	);
	LUT3 #(
		.INIT('h2a)
	) name13756 (
		\m1_data_i[8]_pad ,
		_w8910_,
		_w8911_,
		_w15657_
	);
	LUT3 #(
		.INIT('h80)
	) name13757 (
		\m2_data_i[8]_pad ,
		_w8910_,
		_w8911_,
		_w15658_
	);
	LUT4 #(
		.INIT('h3b7f)
	) name13758 (
		_w8905_,
		_w8908_,
		_w15657_,
		_w15658_,
		_w15659_
	);
	LUT3 #(
		.INIT('h80)
	) name13759 (
		\m0_data_i[8]_pad ,
		_w8910_,
		_w8911_,
		_w15660_
	);
	LUT3 #(
		.INIT('h80)
	) name13760 (
		\m4_data_i[8]_pad ,
		_w8910_,
		_w8911_,
		_w15661_
	);
	LUT4 #(
		.INIT('h5d7f)
	) name13761 (
		_w8905_,
		_w8908_,
		_w15660_,
		_w15661_,
		_w15662_
	);
	LUT3 #(
		.INIT('h2a)
	) name13762 (
		\m7_data_i[8]_pad ,
		_w8910_,
		_w8911_,
		_w15663_
	);
	LUT3 #(
		.INIT('h2a)
	) name13763 (
		\m3_data_i[8]_pad ,
		_w8910_,
		_w8911_,
		_w15664_
	);
	LUT4 #(
		.INIT('habef)
	) name13764 (
		_w8905_,
		_w8908_,
		_w15663_,
		_w15664_,
		_w15665_
	);
	LUT3 #(
		.INIT('h80)
	) name13765 (
		\m6_data_i[8]_pad ,
		_w8910_,
		_w8911_,
		_w15666_
	);
	LUT3 #(
		.INIT('h2a)
	) name13766 (
		\m5_data_i[8]_pad ,
		_w8910_,
		_w8911_,
		_w15667_
	);
	LUT4 #(
		.INIT('hcdef)
	) name13767 (
		_w8905_,
		_w8908_,
		_w15666_,
		_w15667_,
		_w15668_
	);
	LUT4 #(
		.INIT('h7fff)
	) name13768 (
		_w15659_,
		_w15662_,
		_w15665_,
		_w15668_,
		_w15669_
	);
	LUT3 #(
		.INIT('h80)
	) name13769 (
		\m0_data_i[9]_pad ,
		_w8910_,
		_w8911_,
		_w15670_
	);
	LUT3 #(
		.INIT('h2a)
	) name13770 (
		\m7_data_i[9]_pad ,
		_w8910_,
		_w8911_,
		_w15671_
	);
	LUT4 #(
		.INIT('h6e7f)
	) name13771 (
		_w8905_,
		_w8908_,
		_w15670_,
		_w15671_,
		_w15672_
	);
	LUT3 #(
		.INIT('h2a)
	) name13772 (
		\m1_data_i[9]_pad ,
		_w8910_,
		_w8911_,
		_w15673_
	);
	LUT3 #(
		.INIT('h2a)
	) name13773 (
		\m5_data_i[9]_pad ,
		_w8910_,
		_w8911_,
		_w15674_
	);
	LUT4 #(
		.INIT('h5d7f)
	) name13774 (
		_w8905_,
		_w8908_,
		_w15673_,
		_w15674_,
		_w15675_
	);
	LUT3 #(
		.INIT('h80)
	) name13775 (
		\m2_data_i[9]_pad ,
		_w8910_,
		_w8911_,
		_w15676_
	);
	LUT3 #(
		.INIT('h80)
	) name13776 (
		\m6_data_i[9]_pad ,
		_w8910_,
		_w8911_,
		_w15677_
	);
	LUT4 #(
		.INIT('haebf)
	) name13777 (
		_w8905_,
		_w8908_,
		_w15676_,
		_w15677_,
		_w15678_
	);
	LUT3 #(
		.INIT('h2a)
	) name13778 (
		\m3_data_i[9]_pad ,
		_w8910_,
		_w8911_,
		_w15679_
	);
	LUT3 #(
		.INIT('h80)
	) name13779 (
		\m4_data_i[9]_pad ,
		_w8910_,
		_w8911_,
		_w15680_
	);
	LUT4 #(
		.INIT('h9dbf)
	) name13780 (
		_w8905_,
		_w8908_,
		_w15679_,
		_w15680_,
		_w15681_
	);
	LUT4 #(
		.INIT('h7fff)
	) name13781 (
		_w15672_,
		_w15675_,
		_w15678_,
		_w15681_,
		_w15682_
	);
	LUT3 #(
		.INIT('h80)
	) name13782 (
		\m0_sel_i[0]_pad ,
		_w8910_,
		_w8911_,
		_w15683_
	);
	LUT3 #(
		.INIT('h2a)
	) name13783 (
		\m7_sel_i[0]_pad ,
		_w8910_,
		_w8911_,
		_w15684_
	);
	LUT4 #(
		.INIT('h6e7f)
	) name13784 (
		_w8905_,
		_w8908_,
		_w15683_,
		_w15684_,
		_w15685_
	);
	LUT3 #(
		.INIT('h2a)
	) name13785 (
		\m3_sel_i[0]_pad ,
		_w8910_,
		_w8911_,
		_w15686_
	);
	LUT3 #(
		.INIT('h80)
	) name13786 (
		\m2_sel_i[0]_pad ,
		_w8910_,
		_w8911_,
		_w15687_
	);
	LUT3 #(
		.INIT('h57)
	) name13787 (
		_w8909_,
		_w15686_,
		_w15687_,
		_w15688_
	);
	LUT3 #(
		.INIT('h80)
	) name13788 (
		\m4_sel_i[0]_pad ,
		_w8910_,
		_w8911_,
		_w15689_
	);
	LUT3 #(
		.INIT('h2a)
	) name13789 (
		\m1_sel_i[0]_pad ,
		_w8910_,
		_w8911_,
		_w15690_
	);
	LUT4 #(
		.INIT('h57df)
	) name13790 (
		_w8905_,
		_w8908_,
		_w15689_,
		_w15690_,
		_w15691_
	);
	LUT3 #(
		.INIT('h80)
	) name13791 (
		\m6_sel_i[0]_pad ,
		_w8910_,
		_w8911_,
		_w15692_
	);
	LUT3 #(
		.INIT('h2a)
	) name13792 (
		\m5_sel_i[0]_pad ,
		_w8910_,
		_w8911_,
		_w15693_
	);
	LUT4 #(
		.INIT('hcdef)
	) name13793 (
		_w8905_,
		_w8908_,
		_w15692_,
		_w15693_,
		_w15694_
	);
	LUT4 #(
		.INIT('h7fff)
	) name13794 (
		_w15685_,
		_w15688_,
		_w15691_,
		_w15694_,
		_w15695_
	);
	LUT3 #(
		.INIT('h80)
	) name13795 (
		\m0_sel_i[1]_pad ,
		_w8910_,
		_w8911_,
		_w15696_
	);
	LUT3 #(
		.INIT('h2a)
	) name13796 (
		\m7_sel_i[1]_pad ,
		_w8910_,
		_w8911_,
		_w15697_
	);
	LUT4 #(
		.INIT('h6e7f)
	) name13797 (
		_w8905_,
		_w8908_,
		_w15696_,
		_w15697_,
		_w15698_
	);
	LUT3 #(
		.INIT('h2a)
	) name13798 (
		\m1_sel_i[1]_pad ,
		_w8910_,
		_w8911_,
		_w15699_
	);
	LUT3 #(
		.INIT('h80)
	) name13799 (
		\m4_sel_i[1]_pad ,
		_w8910_,
		_w8911_,
		_w15700_
	);
	LUT4 #(
		.INIT('h5d7f)
	) name13800 (
		_w8905_,
		_w8908_,
		_w15699_,
		_w15700_,
		_w15701_
	);
	LUT3 #(
		.INIT('h80)
	) name13801 (
		\m2_sel_i[1]_pad ,
		_w8910_,
		_w8911_,
		_w15702_
	);
	LUT3 #(
		.INIT('h2a)
	) name13802 (
		\m3_sel_i[1]_pad ,
		_w8910_,
		_w8911_,
		_w15703_
	);
	LUT3 #(
		.INIT('h57)
	) name13803 (
		_w8909_,
		_w15702_,
		_w15703_,
		_w15704_
	);
	LUT3 #(
		.INIT('h80)
	) name13804 (
		\m6_sel_i[1]_pad ,
		_w8910_,
		_w8911_,
		_w15705_
	);
	LUT3 #(
		.INIT('h2a)
	) name13805 (
		\m5_sel_i[1]_pad ,
		_w8910_,
		_w8911_,
		_w15706_
	);
	LUT4 #(
		.INIT('hcdef)
	) name13806 (
		_w8905_,
		_w8908_,
		_w15705_,
		_w15706_,
		_w15707_
	);
	LUT4 #(
		.INIT('h7fff)
	) name13807 (
		_w15698_,
		_w15701_,
		_w15704_,
		_w15707_,
		_w15708_
	);
	LUT3 #(
		.INIT('h2a)
	) name13808 (
		\m1_sel_i[2]_pad ,
		_w8910_,
		_w8911_,
		_w15709_
	);
	LUT3 #(
		.INIT('h80)
	) name13809 (
		\m2_sel_i[2]_pad ,
		_w8910_,
		_w8911_,
		_w15710_
	);
	LUT4 #(
		.INIT('h3b7f)
	) name13810 (
		_w8905_,
		_w8908_,
		_w15709_,
		_w15710_,
		_w15711_
	);
	LUT3 #(
		.INIT('h80)
	) name13811 (
		\m0_sel_i[2]_pad ,
		_w8910_,
		_w8911_,
		_w15712_
	);
	LUT3 #(
		.INIT('h80)
	) name13812 (
		\m4_sel_i[2]_pad ,
		_w8910_,
		_w8911_,
		_w15713_
	);
	LUT4 #(
		.INIT('h5d7f)
	) name13813 (
		_w8905_,
		_w8908_,
		_w15712_,
		_w15713_,
		_w15714_
	);
	LUT3 #(
		.INIT('h2a)
	) name13814 (
		\m7_sel_i[2]_pad ,
		_w8910_,
		_w8911_,
		_w15715_
	);
	LUT3 #(
		.INIT('h2a)
	) name13815 (
		\m3_sel_i[2]_pad ,
		_w8910_,
		_w8911_,
		_w15716_
	);
	LUT4 #(
		.INIT('habef)
	) name13816 (
		_w8905_,
		_w8908_,
		_w15715_,
		_w15716_,
		_w15717_
	);
	LUT3 #(
		.INIT('h80)
	) name13817 (
		\m6_sel_i[2]_pad ,
		_w8910_,
		_w8911_,
		_w15718_
	);
	LUT3 #(
		.INIT('h2a)
	) name13818 (
		\m5_sel_i[2]_pad ,
		_w8910_,
		_w8911_,
		_w15719_
	);
	LUT4 #(
		.INIT('hcdef)
	) name13819 (
		_w8905_,
		_w8908_,
		_w15718_,
		_w15719_,
		_w15720_
	);
	LUT4 #(
		.INIT('h7fff)
	) name13820 (
		_w15711_,
		_w15714_,
		_w15717_,
		_w15720_,
		_w15721_
	);
	LUT3 #(
		.INIT('h2a)
	) name13821 (
		\m1_sel_i[3]_pad ,
		_w8910_,
		_w8911_,
		_w15722_
	);
	LUT3 #(
		.INIT('h80)
	) name13822 (
		\m2_sel_i[3]_pad ,
		_w8910_,
		_w8911_,
		_w15723_
	);
	LUT4 #(
		.INIT('h3b7f)
	) name13823 (
		_w8905_,
		_w8908_,
		_w15722_,
		_w15723_,
		_w15724_
	);
	LUT3 #(
		.INIT('h80)
	) name13824 (
		\m0_sel_i[3]_pad ,
		_w8910_,
		_w8911_,
		_w15725_
	);
	LUT3 #(
		.INIT('h80)
	) name13825 (
		\m4_sel_i[3]_pad ,
		_w8910_,
		_w8911_,
		_w15726_
	);
	LUT4 #(
		.INIT('h5d7f)
	) name13826 (
		_w8905_,
		_w8908_,
		_w15725_,
		_w15726_,
		_w15727_
	);
	LUT3 #(
		.INIT('h2a)
	) name13827 (
		\m7_sel_i[3]_pad ,
		_w8910_,
		_w8911_,
		_w15728_
	);
	LUT3 #(
		.INIT('h2a)
	) name13828 (
		\m3_sel_i[3]_pad ,
		_w8910_,
		_w8911_,
		_w15729_
	);
	LUT4 #(
		.INIT('habef)
	) name13829 (
		_w8905_,
		_w8908_,
		_w15728_,
		_w15729_,
		_w15730_
	);
	LUT3 #(
		.INIT('h80)
	) name13830 (
		\m6_sel_i[3]_pad ,
		_w8910_,
		_w8911_,
		_w15731_
	);
	LUT3 #(
		.INIT('h2a)
	) name13831 (
		\m5_sel_i[3]_pad ,
		_w8910_,
		_w8911_,
		_w15732_
	);
	LUT4 #(
		.INIT('hcdef)
	) name13832 (
		_w8905_,
		_w8908_,
		_w15731_,
		_w15732_,
		_w15733_
	);
	LUT4 #(
		.INIT('h7fff)
	) name13833 (
		_w15724_,
		_w15727_,
		_w15730_,
		_w15733_,
		_w15734_
	);
	LUT4 #(
		.INIT('h2a00)
	) name13834 (
		\m3_stb_i_pad ,
		_w8910_,
		_w8911_,
		_w9480_,
		_w15735_
	);
	LUT4 #(
		.INIT('h8000)
	) name13835 (
		\m2_stb_i_pad ,
		_w8910_,
		_w8911_,
		_w9451_,
		_w15736_
	);
	LUT3 #(
		.INIT('h57)
	) name13836 (
		_w8909_,
		_w15735_,
		_w15736_,
		_w15737_
	);
	LUT4 #(
		.INIT('h8000)
	) name13837 (
		\m6_stb_i_pad ,
		_w8910_,
		_w8911_,
		_w9559_,
		_w15738_
	);
	LUT4 #(
		.INIT('h2a00)
	) name13838 (
		\m1_stb_i_pad ,
		_w8910_,
		_w8911_,
		_w9413_,
		_w15739_
	);
	LUT4 #(
		.INIT('h67ef)
	) name13839 (
		_w8905_,
		_w8908_,
		_w15738_,
		_w15739_,
		_w15740_
	);
	LUT4 #(
		.INIT('h2a00)
	) name13840 (
		\m7_stb_i_pad ,
		_w8910_,
		_w8911_,
		_w9594_,
		_w15741_
	);
	LUT4 #(
		.INIT('h2a00)
	) name13841 (
		\m5_stb_i_pad ,
		_w8910_,
		_w8911_,
		_w9532_,
		_w15742_
	);
	LUT4 #(
		.INIT('hcdef)
	) name13842 (
		_w8905_,
		_w8908_,
		_w15741_,
		_w15742_,
		_w15743_
	);
	LUT4 #(
		.INIT('h8000)
	) name13843 (
		\m4_stb_i_pad ,
		_w8910_,
		_w8911_,
		_w9509_,
		_w15744_
	);
	LUT4 #(
		.INIT('h8000)
	) name13844 (
		\m0_stb_i_pad ,
		_w8910_,
		_w8911_,
		_w9381_,
		_w15745_
	);
	LUT4 #(
		.INIT('h57df)
	) name13845 (
		_w8905_,
		_w8908_,
		_w15744_,
		_w15745_,
		_w15746_
	);
	LUT4 #(
		.INIT('h7fff)
	) name13846 (
		_w15737_,
		_w15740_,
		_w15743_,
		_w15746_,
		_w15747_
	);
	LUT3 #(
		.INIT('h80)
	) name13847 (
		\m6_we_i_pad ,
		_w8910_,
		_w8911_,
		_w15748_
	);
	LUT3 #(
		.INIT('h2a)
	) name13848 (
		\m5_we_i_pad ,
		_w8910_,
		_w8911_,
		_w15749_
	);
	LUT4 #(
		.INIT('hcdef)
	) name13849 (
		_w8905_,
		_w8908_,
		_w15748_,
		_w15749_,
		_w15750_
	);
	LUT3 #(
		.INIT('h2a)
	) name13850 (
		\m3_we_i_pad ,
		_w8910_,
		_w8911_,
		_w15751_
	);
	LUT3 #(
		.INIT('h2a)
	) name13851 (
		\m7_we_i_pad ,
		_w8910_,
		_w8911_,
		_w15752_
	);
	LUT4 #(
		.INIT('haebf)
	) name13852 (
		_w8905_,
		_w8908_,
		_w15751_,
		_w15752_,
		_w15753_
	);
	LUT3 #(
		.INIT('h80)
	) name13853 (
		\m4_we_i_pad ,
		_w8910_,
		_w8911_,
		_w15754_
	);
	LUT3 #(
		.INIT('h80)
	) name13854 (
		\m0_we_i_pad ,
		_w8910_,
		_w8911_,
		_w15755_
	);
	LUT4 #(
		.INIT('h57df)
	) name13855 (
		_w8905_,
		_w8908_,
		_w15754_,
		_w15755_,
		_w15756_
	);
	LUT3 #(
		.INIT('h2a)
	) name13856 (
		\m1_we_i_pad ,
		_w8910_,
		_w8911_,
		_w15757_
	);
	LUT3 #(
		.INIT('h80)
	) name13857 (
		\m2_we_i_pad ,
		_w8910_,
		_w8911_,
		_w15758_
	);
	LUT4 #(
		.INIT('h3b7f)
	) name13858 (
		_w8905_,
		_w8908_,
		_w15757_,
		_w15758_,
		_w15759_
	);
	LUT4 #(
		.INIT('h7fff)
	) name13859 (
		_w15750_,
		_w15753_,
		_w15756_,
		_w15759_,
		_w15760_
	);
	LUT3 #(
		.INIT('h2a)
	) name13860 (
		\m1_addr_i[0]_pad ,
		_w8955_,
		_w8956_,
		_w15761_
	);
	LUT3 #(
		.INIT('h80)
	) name13861 (
		\m2_addr_i[0]_pad ,
		_w8955_,
		_w8956_,
		_w15762_
	);
	LUT4 #(
		.INIT('h3b7f)
	) name13862 (
		_w8950_,
		_w8953_,
		_w15761_,
		_w15762_,
		_w15763_
	);
	LUT3 #(
		.INIT('h80)
	) name13863 (
		\m0_addr_i[0]_pad ,
		_w8955_,
		_w8956_,
		_w15764_
	);
	LUT3 #(
		.INIT('h2a)
	) name13864 (
		\m5_addr_i[0]_pad ,
		_w8955_,
		_w8956_,
		_w15765_
	);
	LUT4 #(
		.INIT('h5d7f)
	) name13865 (
		_w8950_,
		_w8953_,
		_w15764_,
		_w15765_,
		_w15766_
	);
	LUT3 #(
		.INIT('h2a)
	) name13866 (
		\m7_addr_i[0]_pad ,
		_w8955_,
		_w8956_,
		_w15767_
	);
	LUT3 #(
		.INIT('h80)
	) name13867 (
		\m6_addr_i[0]_pad ,
		_w8955_,
		_w8956_,
		_w15768_
	);
	LUT3 #(
		.INIT('h57)
	) name13868 (
		_w8968_,
		_w15767_,
		_w15768_,
		_w15769_
	);
	LUT3 #(
		.INIT('h2a)
	) name13869 (
		\m3_addr_i[0]_pad ,
		_w8955_,
		_w8956_,
		_w15770_
	);
	LUT3 #(
		.INIT('h80)
	) name13870 (
		\m4_addr_i[0]_pad ,
		_w8955_,
		_w8956_,
		_w15771_
	);
	LUT4 #(
		.INIT('h9dbf)
	) name13871 (
		_w8950_,
		_w8953_,
		_w15770_,
		_w15771_,
		_w15772_
	);
	LUT4 #(
		.INIT('h7fff)
	) name13872 (
		_w15763_,
		_w15766_,
		_w15769_,
		_w15772_,
		_w15773_
	);
	LUT3 #(
		.INIT('h2a)
	) name13873 (
		\m1_addr_i[10]_pad ,
		_w8955_,
		_w8956_,
		_w15774_
	);
	LUT3 #(
		.INIT('h80)
	) name13874 (
		\m2_addr_i[10]_pad ,
		_w8955_,
		_w8956_,
		_w15775_
	);
	LUT4 #(
		.INIT('h3b7f)
	) name13875 (
		_w8950_,
		_w8953_,
		_w15774_,
		_w15775_,
		_w15776_
	);
	LUT3 #(
		.INIT('h80)
	) name13876 (
		\m6_addr_i[10]_pad ,
		_w8955_,
		_w8956_,
		_w15777_
	);
	LUT3 #(
		.INIT('h80)
	) name13877 (
		\m4_addr_i[10]_pad ,
		_w8955_,
		_w8956_,
		_w15778_
	);
	LUT4 #(
		.INIT('hcdef)
	) name13878 (
		_w8950_,
		_w8953_,
		_w15777_,
		_w15778_,
		_w15779_
	);
	LUT3 #(
		.INIT('h2a)
	) name13879 (
		\m5_addr_i[10]_pad ,
		_w8955_,
		_w8956_,
		_w15780_
	);
	LUT3 #(
		.INIT('h2a)
	) name13880 (
		\m3_addr_i[10]_pad ,
		_w8955_,
		_w8956_,
		_w15781_
	);
	LUT4 #(
		.INIT('h9bdf)
	) name13881 (
		_w8950_,
		_w8953_,
		_w15780_,
		_w15781_,
		_w15782_
	);
	LUT3 #(
		.INIT('h80)
	) name13882 (
		\m0_addr_i[10]_pad ,
		_w8955_,
		_w8956_,
		_w15783_
	);
	LUT3 #(
		.INIT('h2a)
	) name13883 (
		\m7_addr_i[10]_pad ,
		_w8955_,
		_w8956_,
		_w15784_
	);
	LUT4 #(
		.INIT('h6e7f)
	) name13884 (
		_w8950_,
		_w8953_,
		_w15783_,
		_w15784_,
		_w15785_
	);
	LUT4 #(
		.INIT('h7fff)
	) name13885 (
		_w15776_,
		_w15779_,
		_w15782_,
		_w15785_,
		_w15786_
	);
	LUT3 #(
		.INIT('h2a)
	) name13886 (
		\m1_addr_i[11]_pad ,
		_w8955_,
		_w8956_,
		_w15787_
	);
	LUT3 #(
		.INIT('h80)
	) name13887 (
		\m2_addr_i[11]_pad ,
		_w8955_,
		_w8956_,
		_w15788_
	);
	LUT4 #(
		.INIT('h3b7f)
	) name13888 (
		_w8950_,
		_w8953_,
		_w15787_,
		_w15788_,
		_w15789_
	);
	LUT3 #(
		.INIT('h2a)
	) name13889 (
		\m3_addr_i[11]_pad ,
		_w8955_,
		_w8956_,
		_w15790_
	);
	LUT3 #(
		.INIT('h2a)
	) name13890 (
		\m5_addr_i[11]_pad ,
		_w8955_,
		_w8956_,
		_w15791_
	);
	LUT4 #(
		.INIT('h9dbf)
	) name13891 (
		_w8950_,
		_w8953_,
		_w15790_,
		_w15791_,
		_w15792_
	);
	LUT3 #(
		.INIT('h80)
	) name13892 (
		\m4_addr_i[11]_pad ,
		_w8955_,
		_w8956_,
		_w15793_
	);
	LUT3 #(
		.INIT('h80)
	) name13893 (
		\m6_addr_i[11]_pad ,
		_w8955_,
		_w8956_,
		_w15794_
	);
	LUT4 #(
		.INIT('hcedf)
	) name13894 (
		_w8950_,
		_w8953_,
		_w15793_,
		_w15794_,
		_w15795_
	);
	LUT3 #(
		.INIT('h80)
	) name13895 (
		\m0_addr_i[11]_pad ,
		_w8955_,
		_w8956_,
		_w15796_
	);
	LUT3 #(
		.INIT('h2a)
	) name13896 (
		\m7_addr_i[11]_pad ,
		_w8955_,
		_w8956_,
		_w15797_
	);
	LUT4 #(
		.INIT('h6e7f)
	) name13897 (
		_w8950_,
		_w8953_,
		_w15796_,
		_w15797_,
		_w15798_
	);
	LUT4 #(
		.INIT('h7fff)
	) name13898 (
		_w15789_,
		_w15792_,
		_w15795_,
		_w15798_,
		_w15799_
	);
	LUT3 #(
		.INIT('h80)
	) name13899 (
		\m0_addr_i[12]_pad ,
		_w8955_,
		_w8956_,
		_w15800_
	);
	LUT3 #(
		.INIT('h2a)
	) name13900 (
		\m7_addr_i[12]_pad ,
		_w8955_,
		_w8956_,
		_w15801_
	);
	LUT4 #(
		.INIT('h6e7f)
	) name13901 (
		_w8950_,
		_w8953_,
		_w15800_,
		_w15801_,
		_w15802_
	);
	LUT3 #(
		.INIT('h80)
	) name13902 (
		\m6_addr_i[12]_pad ,
		_w8955_,
		_w8956_,
		_w15803_
	);
	LUT3 #(
		.INIT('h80)
	) name13903 (
		\m4_addr_i[12]_pad ,
		_w8955_,
		_w8956_,
		_w15804_
	);
	LUT4 #(
		.INIT('hcdef)
	) name13904 (
		_w8950_,
		_w8953_,
		_w15803_,
		_w15804_,
		_w15805_
	);
	LUT3 #(
		.INIT('h2a)
	) name13905 (
		\m5_addr_i[12]_pad ,
		_w8955_,
		_w8956_,
		_w15806_
	);
	LUT3 #(
		.INIT('h2a)
	) name13906 (
		\m3_addr_i[12]_pad ,
		_w8955_,
		_w8956_,
		_w15807_
	);
	LUT4 #(
		.INIT('h9bdf)
	) name13907 (
		_w8950_,
		_w8953_,
		_w15806_,
		_w15807_,
		_w15808_
	);
	LUT3 #(
		.INIT('h2a)
	) name13908 (
		\m1_addr_i[12]_pad ,
		_w8955_,
		_w8956_,
		_w15809_
	);
	LUT3 #(
		.INIT('h80)
	) name13909 (
		\m2_addr_i[12]_pad ,
		_w8955_,
		_w8956_,
		_w15810_
	);
	LUT4 #(
		.INIT('h3b7f)
	) name13910 (
		_w8950_,
		_w8953_,
		_w15809_,
		_w15810_,
		_w15811_
	);
	LUT4 #(
		.INIT('h7fff)
	) name13911 (
		_w15802_,
		_w15805_,
		_w15808_,
		_w15811_,
		_w15812_
	);
	LUT3 #(
		.INIT('h2a)
	) name13912 (
		\m3_addr_i[13]_pad ,
		_w8955_,
		_w8956_,
		_w15813_
	);
	LUT3 #(
		.INIT('h80)
	) name13913 (
		\m4_addr_i[13]_pad ,
		_w8955_,
		_w8956_,
		_w15814_
	);
	LUT4 #(
		.INIT('h9dbf)
	) name13914 (
		_w8950_,
		_w8953_,
		_w15813_,
		_w15814_,
		_w15815_
	);
	LUT3 #(
		.INIT('h2a)
	) name13915 (
		\m1_addr_i[13]_pad ,
		_w8955_,
		_w8956_,
		_w15816_
	);
	LUT3 #(
		.INIT('h2a)
	) name13916 (
		\m7_addr_i[13]_pad ,
		_w8955_,
		_w8956_,
		_w15817_
	);
	LUT4 #(
		.INIT('h6e7f)
	) name13917 (
		_w8950_,
		_w8953_,
		_w15816_,
		_w15817_,
		_w15818_
	);
	LUT3 #(
		.INIT('h80)
	) name13918 (
		\m2_addr_i[13]_pad ,
		_w8955_,
		_w8956_,
		_w15819_
	);
	LUT3 #(
		.INIT('h80)
	) name13919 (
		\m0_addr_i[13]_pad ,
		_w8955_,
		_w8956_,
		_w15820_
	);
	LUT4 #(
		.INIT('h37bf)
	) name13920 (
		_w8950_,
		_w8953_,
		_w15819_,
		_w15820_,
		_w15821_
	);
	LUT3 #(
		.INIT('h80)
	) name13921 (
		\m6_addr_i[13]_pad ,
		_w8955_,
		_w8956_,
		_w15822_
	);
	LUT3 #(
		.INIT('h2a)
	) name13922 (
		\m5_addr_i[13]_pad ,
		_w8955_,
		_w8956_,
		_w15823_
	);
	LUT4 #(
		.INIT('hcdef)
	) name13923 (
		_w8950_,
		_w8953_,
		_w15822_,
		_w15823_,
		_w15824_
	);
	LUT4 #(
		.INIT('h7fff)
	) name13924 (
		_w15815_,
		_w15818_,
		_w15821_,
		_w15824_,
		_w15825_
	);
	LUT3 #(
		.INIT('h2a)
	) name13925 (
		\m1_addr_i[14]_pad ,
		_w8955_,
		_w8956_,
		_w15826_
	);
	LUT3 #(
		.INIT('h80)
	) name13926 (
		\m2_addr_i[14]_pad ,
		_w8955_,
		_w8956_,
		_w15827_
	);
	LUT4 #(
		.INIT('h3b7f)
	) name13927 (
		_w8950_,
		_w8953_,
		_w15826_,
		_w15827_,
		_w15828_
	);
	LUT3 #(
		.INIT('h80)
	) name13928 (
		\m0_addr_i[14]_pad ,
		_w8955_,
		_w8956_,
		_w15829_
	);
	LUT3 #(
		.INIT('h80)
	) name13929 (
		\m4_addr_i[14]_pad ,
		_w8955_,
		_w8956_,
		_w15830_
	);
	LUT4 #(
		.INIT('h5d7f)
	) name13930 (
		_w8950_,
		_w8953_,
		_w15829_,
		_w15830_,
		_w15831_
	);
	LUT3 #(
		.INIT('h2a)
	) name13931 (
		\m7_addr_i[14]_pad ,
		_w8955_,
		_w8956_,
		_w15832_
	);
	LUT3 #(
		.INIT('h2a)
	) name13932 (
		\m3_addr_i[14]_pad ,
		_w8955_,
		_w8956_,
		_w15833_
	);
	LUT4 #(
		.INIT('habef)
	) name13933 (
		_w8950_,
		_w8953_,
		_w15832_,
		_w15833_,
		_w15834_
	);
	LUT3 #(
		.INIT('h80)
	) name13934 (
		\m6_addr_i[14]_pad ,
		_w8955_,
		_w8956_,
		_w15835_
	);
	LUT3 #(
		.INIT('h2a)
	) name13935 (
		\m5_addr_i[14]_pad ,
		_w8955_,
		_w8956_,
		_w15836_
	);
	LUT4 #(
		.INIT('hcdef)
	) name13936 (
		_w8950_,
		_w8953_,
		_w15835_,
		_w15836_,
		_w15837_
	);
	LUT4 #(
		.INIT('h7fff)
	) name13937 (
		_w15828_,
		_w15831_,
		_w15834_,
		_w15837_,
		_w15838_
	);
	LUT3 #(
		.INIT('h80)
	) name13938 (
		\m6_addr_i[15]_pad ,
		_w8955_,
		_w8956_,
		_w15839_
	);
	LUT3 #(
		.INIT('h2a)
	) name13939 (
		\m5_addr_i[15]_pad ,
		_w8955_,
		_w8956_,
		_w15840_
	);
	LUT4 #(
		.INIT('hcdef)
	) name13940 (
		_w8950_,
		_w8953_,
		_w15839_,
		_w15840_,
		_w15841_
	);
	LUT3 #(
		.INIT('h2a)
	) name13941 (
		\m3_addr_i[15]_pad ,
		_w8955_,
		_w8956_,
		_w15842_
	);
	LUT3 #(
		.INIT('h80)
	) name13942 (
		\m2_addr_i[15]_pad ,
		_w8955_,
		_w8956_,
		_w15843_
	);
	LUT3 #(
		.INIT('h57)
	) name13943 (
		_w8974_,
		_w15842_,
		_w15843_,
		_w15844_
	);
	LUT3 #(
		.INIT('h80)
	) name13944 (
		\m4_addr_i[15]_pad ,
		_w8955_,
		_w8956_,
		_w15845_
	);
	LUT3 #(
		.INIT('h2a)
	) name13945 (
		\m1_addr_i[15]_pad ,
		_w8955_,
		_w8956_,
		_w15846_
	);
	LUT4 #(
		.INIT('h57df)
	) name13946 (
		_w8950_,
		_w8953_,
		_w15845_,
		_w15846_,
		_w15847_
	);
	LUT3 #(
		.INIT('h80)
	) name13947 (
		\m0_addr_i[15]_pad ,
		_w8955_,
		_w8956_,
		_w15848_
	);
	LUT3 #(
		.INIT('h2a)
	) name13948 (
		\m7_addr_i[15]_pad ,
		_w8955_,
		_w8956_,
		_w15849_
	);
	LUT4 #(
		.INIT('h6e7f)
	) name13949 (
		_w8950_,
		_w8953_,
		_w15848_,
		_w15849_,
		_w15850_
	);
	LUT4 #(
		.INIT('h7fff)
	) name13950 (
		_w15841_,
		_w15844_,
		_w15847_,
		_w15850_,
		_w15851_
	);
	LUT3 #(
		.INIT('h80)
	) name13951 (
		\m0_addr_i[16]_pad ,
		_w8955_,
		_w8956_,
		_w15852_
	);
	LUT3 #(
		.INIT('h2a)
	) name13952 (
		\m7_addr_i[16]_pad ,
		_w8955_,
		_w8956_,
		_w15853_
	);
	LUT4 #(
		.INIT('h6e7f)
	) name13953 (
		_w8950_,
		_w8953_,
		_w15852_,
		_w15853_,
		_w15854_
	);
	LUT3 #(
		.INIT('h80)
	) name13954 (
		\m6_addr_i[16]_pad ,
		_w8955_,
		_w8956_,
		_w15855_
	);
	LUT3 #(
		.INIT('h80)
	) name13955 (
		\m4_addr_i[16]_pad ,
		_w8955_,
		_w8956_,
		_w15856_
	);
	LUT4 #(
		.INIT('hcdef)
	) name13956 (
		_w8950_,
		_w8953_,
		_w15855_,
		_w15856_,
		_w15857_
	);
	LUT3 #(
		.INIT('h2a)
	) name13957 (
		\m5_addr_i[16]_pad ,
		_w8955_,
		_w8956_,
		_w15858_
	);
	LUT3 #(
		.INIT('h2a)
	) name13958 (
		\m3_addr_i[16]_pad ,
		_w8955_,
		_w8956_,
		_w15859_
	);
	LUT4 #(
		.INIT('h9bdf)
	) name13959 (
		_w8950_,
		_w8953_,
		_w15858_,
		_w15859_,
		_w15860_
	);
	LUT3 #(
		.INIT('h2a)
	) name13960 (
		\m1_addr_i[16]_pad ,
		_w8955_,
		_w8956_,
		_w15861_
	);
	LUT3 #(
		.INIT('h80)
	) name13961 (
		\m2_addr_i[16]_pad ,
		_w8955_,
		_w8956_,
		_w15862_
	);
	LUT4 #(
		.INIT('h3b7f)
	) name13962 (
		_w8950_,
		_w8953_,
		_w15861_,
		_w15862_,
		_w15863_
	);
	LUT4 #(
		.INIT('h7fff)
	) name13963 (
		_w15854_,
		_w15857_,
		_w15860_,
		_w15863_,
		_w15864_
	);
	LUT3 #(
		.INIT('h80)
	) name13964 (
		\m6_addr_i[17]_pad ,
		_w8955_,
		_w8956_,
		_w15865_
	);
	LUT3 #(
		.INIT('h2a)
	) name13965 (
		\m5_addr_i[17]_pad ,
		_w8955_,
		_w8956_,
		_w15866_
	);
	LUT4 #(
		.INIT('hcdef)
	) name13966 (
		_w8950_,
		_w8953_,
		_w15865_,
		_w15866_,
		_w15867_
	);
	LUT3 #(
		.INIT('h80)
	) name13967 (
		\m0_addr_i[17]_pad ,
		_w8955_,
		_w8956_,
		_w15868_
	);
	LUT3 #(
		.INIT('h80)
	) name13968 (
		\m2_addr_i[17]_pad ,
		_w8955_,
		_w8956_,
		_w15869_
	);
	LUT4 #(
		.INIT('h3b7f)
	) name13969 (
		_w8950_,
		_w8953_,
		_w15868_,
		_w15869_,
		_w15870_
	);
	LUT3 #(
		.INIT('h2a)
	) name13970 (
		\m7_addr_i[17]_pad ,
		_w8955_,
		_w8956_,
		_w15871_
	);
	LUT3 #(
		.INIT('h2a)
	) name13971 (
		\m1_addr_i[17]_pad ,
		_w8955_,
		_w8956_,
		_w15872_
	);
	LUT4 #(
		.INIT('h67ef)
	) name13972 (
		_w8950_,
		_w8953_,
		_w15871_,
		_w15872_,
		_w15873_
	);
	LUT3 #(
		.INIT('h2a)
	) name13973 (
		\m3_addr_i[17]_pad ,
		_w8955_,
		_w8956_,
		_w15874_
	);
	LUT3 #(
		.INIT('h80)
	) name13974 (
		\m4_addr_i[17]_pad ,
		_w8955_,
		_w8956_,
		_w15875_
	);
	LUT4 #(
		.INIT('h9dbf)
	) name13975 (
		_w8950_,
		_w8953_,
		_w15874_,
		_w15875_,
		_w15876_
	);
	LUT4 #(
		.INIT('h7fff)
	) name13976 (
		_w15867_,
		_w15870_,
		_w15873_,
		_w15876_,
		_w15877_
	);
	LUT3 #(
		.INIT('h80)
	) name13977 (
		\m6_addr_i[18]_pad ,
		_w8955_,
		_w8956_,
		_w15878_
	);
	LUT3 #(
		.INIT('h2a)
	) name13978 (
		\m5_addr_i[18]_pad ,
		_w8955_,
		_w8956_,
		_w15879_
	);
	LUT4 #(
		.INIT('hcdef)
	) name13979 (
		_w8950_,
		_w8953_,
		_w15878_,
		_w15879_,
		_w15880_
	);
	LUT3 #(
		.INIT('h80)
	) name13980 (
		\m0_addr_i[18]_pad ,
		_w8955_,
		_w8956_,
		_w15881_
	);
	LUT3 #(
		.INIT('h80)
	) name13981 (
		\m4_addr_i[18]_pad ,
		_w8955_,
		_w8956_,
		_w15882_
	);
	LUT4 #(
		.INIT('h5d7f)
	) name13982 (
		_w8950_,
		_w8953_,
		_w15881_,
		_w15882_,
		_w15883_
	);
	LUT3 #(
		.INIT('h2a)
	) name13983 (
		\m7_addr_i[18]_pad ,
		_w8955_,
		_w8956_,
		_w15884_
	);
	LUT3 #(
		.INIT('h2a)
	) name13984 (
		\m3_addr_i[18]_pad ,
		_w8955_,
		_w8956_,
		_w15885_
	);
	LUT4 #(
		.INIT('habef)
	) name13985 (
		_w8950_,
		_w8953_,
		_w15884_,
		_w15885_,
		_w15886_
	);
	LUT3 #(
		.INIT('h2a)
	) name13986 (
		\m1_addr_i[18]_pad ,
		_w8955_,
		_w8956_,
		_w15887_
	);
	LUT3 #(
		.INIT('h80)
	) name13987 (
		\m2_addr_i[18]_pad ,
		_w8955_,
		_w8956_,
		_w15888_
	);
	LUT4 #(
		.INIT('h3b7f)
	) name13988 (
		_w8950_,
		_w8953_,
		_w15887_,
		_w15888_,
		_w15889_
	);
	LUT4 #(
		.INIT('h7fff)
	) name13989 (
		_w15880_,
		_w15883_,
		_w15886_,
		_w15889_,
		_w15890_
	);
	LUT3 #(
		.INIT('h80)
	) name13990 (
		\m6_addr_i[19]_pad ,
		_w8955_,
		_w8956_,
		_w15891_
	);
	LUT3 #(
		.INIT('h2a)
	) name13991 (
		\m5_addr_i[19]_pad ,
		_w8955_,
		_w8956_,
		_w15892_
	);
	LUT4 #(
		.INIT('hcdef)
	) name13992 (
		_w8950_,
		_w8953_,
		_w15891_,
		_w15892_,
		_w15893_
	);
	LUT3 #(
		.INIT('h80)
	) name13993 (
		\m0_addr_i[19]_pad ,
		_w8955_,
		_w8956_,
		_w15894_
	);
	LUT3 #(
		.INIT('h80)
	) name13994 (
		\m4_addr_i[19]_pad ,
		_w8955_,
		_w8956_,
		_w15895_
	);
	LUT4 #(
		.INIT('h5d7f)
	) name13995 (
		_w8950_,
		_w8953_,
		_w15894_,
		_w15895_,
		_w15896_
	);
	LUT3 #(
		.INIT('h2a)
	) name13996 (
		\m7_addr_i[19]_pad ,
		_w8955_,
		_w8956_,
		_w15897_
	);
	LUT3 #(
		.INIT('h2a)
	) name13997 (
		\m3_addr_i[19]_pad ,
		_w8955_,
		_w8956_,
		_w15898_
	);
	LUT4 #(
		.INIT('habef)
	) name13998 (
		_w8950_,
		_w8953_,
		_w15897_,
		_w15898_,
		_w15899_
	);
	LUT3 #(
		.INIT('h2a)
	) name13999 (
		\m1_addr_i[19]_pad ,
		_w8955_,
		_w8956_,
		_w15900_
	);
	LUT3 #(
		.INIT('h80)
	) name14000 (
		\m2_addr_i[19]_pad ,
		_w8955_,
		_w8956_,
		_w15901_
	);
	LUT4 #(
		.INIT('h3b7f)
	) name14001 (
		_w8950_,
		_w8953_,
		_w15900_,
		_w15901_,
		_w15902_
	);
	LUT4 #(
		.INIT('h7fff)
	) name14002 (
		_w15893_,
		_w15896_,
		_w15899_,
		_w15902_,
		_w15903_
	);
	LUT3 #(
		.INIT('h80)
	) name14003 (
		\m6_addr_i[1]_pad ,
		_w8955_,
		_w8956_,
		_w15904_
	);
	LUT3 #(
		.INIT('h2a)
	) name14004 (
		\m5_addr_i[1]_pad ,
		_w8955_,
		_w8956_,
		_w15905_
	);
	LUT4 #(
		.INIT('hcdef)
	) name14005 (
		_w8950_,
		_w8953_,
		_w15904_,
		_w15905_,
		_w15906_
	);
	LUT3 #(
		.INIT('h80)
	) name14006 (
		\m0_addr_i[1]_pad ,
		_w8955_,
		_w8956_,
		_w15907_
	);
	LUT3 #(
		.INIT('h80)
	) name14007 (
		\m4_addr_i[1]_pad ,
		_w8955_,
		_w8956_,
		_w15908_
	);
	LUT4 #(
		.INIT('h5d7f)
	) name14008 (
		_w8950_,
		_w8953_,
		_w15907_,
		_w15908_,
		_w15909_
	);
	LUT3 #(
		.INIT('h2a)
	) name14009 (
		\m7_addr_i[1]_pad ,
		_w8955_,
		_w8956_,
		_w15910_
	);
	LUT3 #(
		.INIT('h2a)
	) name14010 (
		\m3_addr_i[1]_pad ,
		_w8955_,
		_w8956_,
		_w15911_
	);
	LUT4 #(
		.INIT('habef)
	) name14011 (
		_w8950_,
		_w8953_,
		_w15910_,
		_w15911_,
		_w15912_
	);
	LUT3 #(
		.INIT('h2a)
	) name14012 (
		\m1_addr_i[1]_pad ,
		_w8955_,
		_w8956_,
		_w15913_
	);
	LUT3 #(
		.INIT('h80)
	) name14013 (
		\m2_addr_i[1]_pad ,
		_w8955_,
		_w8956_,
		_w15914_
	);
	LUT4 #(
		.INIT('h3b7f)
	) name14014 (
		_w8950_,
		_w8953_,
		_w15913_,
		_w15914_,
		_w15915_
	);
	LUT4 #(
		.INIT('h7fff)
	) name14015 (
		_w15906_,
		_w15909_,
		_w15912_,
		_w15915_,
		_w15916_
	);
	LUT3 #(
		.INIT('h2a)
	) name14016 (
		\m1_addr_i[20]_pad ,
		_w8955_,
		_w8956_,
		_w15917_
	);
	LUT3 #(
		.INIT('h80)
	) name14017 (
		\m2_addr_i[20]_pad ,
		_w8955_,
		_w8956_,
		_w15918_
	);
	LUT4 #(
		.INIT('h3b7f)
	) name14018 (
		_w8950_,
		_w8953_,
		_w15917_,
		_w15918_,
		_w15919_
	);
	LUT3 #(
		.INIT('h2a)
	) name14019 (
		\m3_addr_i[20]_pad ,
		_w8955_,
		_w8956_,
		_w15920_
	);
	LUT3 #(
		.INIT('h2a)
	) name14020 (
		\m7_addr_i[20]_pad ,
		_w8955_,
		_w8956_,
		_w15921_
	);
	LUT4 #(
		.INIT('haebf)
	) name14021 (
		_w8950_,
		_w8953_,
		_w15920_,
		_w15921_,
		_w15922_
	);
	LUT3 #(
		.INIT('h80)
	) name14022 (
		\m4_addr_i[20]_pad ,
		_w8955_,
		_w8956_,
		_w15923_
	);
	LUT3 #(
		.INIT('h80)
	) name14023 (
		\m0_addr_i[20]_pad ,
		_w8955_,
		_w8956_,
		_w15924_
	);
	LUT4 #(
		.INIT('h57df)
	) name14024 (
		_w8950_,
		_w8953_,
		_w15923_,
		_w15924_,
		_w15925_
	);
	LUT3 #(
		.INIT('h80)
	) name14025 (
		\m6_addr_i[20]_pad ,
		_w8955_,
		_w8956_,
		_w15926_
	);
	LUT3 #(
		.INIT('h2a)
	) name14026 (
		\m5_addr_i[20]_pad ,
		_w8955_,
		_w8956_,
		_w15927_
	);
	LUT4 #(
		.INIT('hcdef)
	) name14027 (
		_w8950_,
		_w8953_,
		_w15926_,
		_w15927_,
		_w15928_
	);
	LUT4 #(
		.INIT('h7fff)
	) name14028 (
		_w15919_,
		_w15922_,
		_w15925_,
		_w15928_,
		_w15929_
	);
	LUT3 #(
		.INIT('h2a)
	) name14029 (
		\m1_addr_i[21]_pad ,
		_w8955_,
		_w8956_,
		_w15930_
	);
	LUT3 #(
		.INIT('h80)
	) name14030 (
		\m2_addr_i[21]_pad ,
		_w8955_,
		_w8956_,
		_w15931_
	);
	LUT4 #(
		.INIT('h3b7f)
	) name14031 (
		_w8950_,
		_w8953_,
		_w15930_,
		_w15931_,
		_w15932_
	);
	LUT3 #(
		.INIT('h2a)
	) name14032 (
		\m3_addr_i[21]_pad ,
		_w8955_,
		_w8956_,
		_w15933_
	);
	LUT3 #(
		.INIT('h2a)
	) name14033 (
		\m5_addr_i[21]_pad ,
		_w8955_,
		_w8956_,
		_w15934_
	);
	LUT4 #(
		.INIT('h9dbf)
	) name14034 (
		_w8950_,
		_w8953_,
		_w15933_,
		_w15934_,
		_w15935_
	);
	LUT3 #(
		.INIT('h80)
	) name14035 (
		\m4_addr_i[21]_pad ,
		_w8955_,
		_w8956_,
		_w15936_
	);
	LUT3 #(
		.INIT('h80)
	) name14036 (
		\m6_addr_i[21]_pad ,
		_w8955_,
		_w8956_,
		_w15937_
	);
	LUT4 #(
		.INIT('hcedf)
	) name14037 (
		_w8950_,
		_w8953_,
		_w15936_,
		_w15937_,
		_w15938_
	);
	LUT3 #(
		.INIT('h80)
	) name14038 (
		\m0_addr_i[21]_pad ,
		_w8955_,
		_w8956_,
		_w15939_
	);
	LUT3 #(
		.INIT('h2a)
	) name14039 (
		\m7_addr_i[21]_pad ,
		_w8955_,
		_w8956_,
		_w15940_
	);
	LUT4 #(
		.INIT('h6e7f)
	) name14040 (
		_w8950_,
		_w8953_,
		_w15939_,
		_w15940_,
		_w15941_
	);
	LUT4 #(
		.INIT('h7fff)
	) name14041 (
		_w15932_,
		_w15935_,
		_w15938_,
		_w15941_,
		_w15942_
	);
	LUT3 #(
		.INIT('h80)
	) name14042 (
		\m0_addr_i[22]_pad ,
		_w8955_,
		_w8956_,
		_w15943_
	);
	LUT3 #(
		.INIT('h2a)
	) name14043 (
		\m7_addr_i[22]_pad ,
		_w8955_,
		_w8956_,
		_w15944_
	);
	LUT4 #(
		.INIT('h6e7f)
	) name14044 (
		_w8950_,
		_w8953_,
		_w15943_,
		_w15944_,
		_w15945_
	);
	LUT3 #(
		.INIT('h80)
	) name14045 (
		\m6_addr_i[22]_pad ,
		_w8955_,
		_w8956_,
		_w15946_
	);
	LUT3 #(
		.INIT('h80)
	) name14046 (
		\m2_addr_i[22]_pad ,
		_w8955_,
		_w8956_,
		_w15947_
	);
	LUT4 #(
		.INIT('habef)
	) name14047 (
		_w8950_,
		_w8953_,
		_w15946_,
		_w15947_,
		_w15948_
	);
	LUT3 #(
		.INIT('h2a)
	) name14048 (
		\m5_addr_i[22]_pad ,
		_w8955_,
		_w8956_,
		_w15949_
	);
	LUT3 #(
		.INIT('h2a)
	) name14049 (
		\m1_addr_i[22]_pad ,
		_w8955_,
		_w8956_,
		_w15950_
	);
	LUT4 #(
		.INIT('h57df)
	) name14050 (
		_w8950_,
		_w8953_,
		_w15949_,
		_w15950_,
		_w15951_
	);
	LUT3 #(
		.INIT('h2a)
	) name14051 (
		\m3_addr_i[22]_pad ,
		_w8955_,
		_w8956_,
		_w15952_
	);
	LUT3 #(
		.INIT('h80)
	) name14052 (
		\m4_addr_i[22]_pad ,
		_w8955_,
		_w8956_,
		_w15953_
	);
	LUT4 #(
		.INIT('h9dbf)
	) name14053 (
		_w8950_,
		_w8953_,
		_w15952_,
		_w15953_,
		_w15954_
	);
	LUT4 #(
		.INIT('h7fff)
	) name14054 (
		_w15945_,
		_w15948_,
		_w15951_,
		_w15954_,
		_w15955_
	);
	LUT3 #(
		.INIT('h2a)
	) name14055 (
		\m3_addr_i[23]_pad ,
		_w8955_,
		_w8956_,
		_w15956_
	);
	LUT3 #(
		.INIT('h80)
	) name14056 (
		\m4_addr_i[23]_pad ,
		_w8955_,
		_w8956_,
		_w15957_
	);
	LUT4 #(
		.INIT('h9dbf)
	) name14057 (
		_w8950_,
		_w8953_,
		_w15956_,
		_w15957_,
		_w15958_
	);
	LUT3 #(
		.INIT('h2a)
	) name14058 (
		\m1_addr_i[23]_pad ,
		_w8955_,
		_w8956_,
		_w15959_
	);
	LUT3 #(
		.INIT('h2a)
	) name14059 (
		\m5_addr_i[23]_pad ,
		_w8955_,
		_w8956_,
		_w15960_
	);
	LUT4 #(
		.INIT('h5d7f)
	) name14060 (
		_w8950_,
		_w8953_,
		_w15959_,
		_w15960_,
		_w15961_
	);
	LUT3 #(
		.INIT('h80)
	) name14061 (
		\m2_addr_i[23]_pad ,
		_w8955_,
		_w8956_,
		_w15962_
	);
	LUT3 #(
		.INIT('h80)
	) name14062 (
		\m6_addr_i[23]_pad ,
		_w8955_,
		_w8956_,
		_w15963_
	);
	LUT4 #(
		.INIT('haebf)
	) name14063 (
		_w8950_,
		_w8953_,
		_w15962_,
		_w15963_,
		_w15964_
	);
	LUT3 #(
		.INIT('h80)
	) name14064 (
		\m0_addr_i[23]_pad ,
		_w8955_,
		_w8956_,
		_w15965_
	);
	LUT3 #(
		.INIT('h2a)
	) name14065 (
		\m7_addr_i[23]_pad ,
		_w8955_,
		_w8956_,
		_w15966_
	);
	LUT4 #(
		.INIT('h6e7f)
	) name14066 (
		_w8950_,
		_w8953_,
		_w15965_,
		_w15966_,
		_w15967_
	);
	LUT4 #(
		.INIT('h7fff)
	) name14067 (
		_w15958_,
		_w15961_,
		_w15964_,
		_w15967_,
		_w15968_
	);
	LUT3 #(
		.INIT('h2a)
	) name14068 (
		\m1_addr_i[24]_pad ,
		_w8955_,
		_w8956_,
		_w15969_
	);
	LUT3 #(
		.INIT('h80)
	) name14069 (
		\m2_addr_i[24]_pad ,
		_w8955_,
		_w8956_,
		_w15970_
	);
	LUT4 #(
		.INIT('h3b7f)
	) name14070 (
		_w8950_,
		_w8953_,
		_w15969_,
		_w15970_,
		_w15971_
	);
	LUT3 #(
		.INIT('h80)
	) name14071 (
		\m0_addr_i[24]_pad ,
		_w8955_,
		_w8956_,
		_w15972_
	);
	LUT3 #(
		.INIT('h80)
	) name14072 (
		\m4_addr_i[24]_pad ,
		_w8955_,
		_w8956_,
		_w15973_
	);
	LUT4 #(
		.INIT('h5d7f)
	) name14073 (
		_w8950_,
		_w8953_,
		_w15972_,
		_w15973_,
		_w15974_
	);
	LUT3 #(
		.INIT('h2a)
	) name14074 (
		\m7_addr_i[24]_pad ,
		_w8955_,
		_w8956_,
		_w15975_
	);
	LUT3 #(
		.INIT('h2a)
	) name14075 (
		\m3_addr_i[24]_pad ,
		_w8955_,
		_w8956_,
		_w15976_
	);
	LUT4 #(
		.INIT('habef)
	) name14076 (
		_w8950_,
		_w8953_,
		_w15975_,
		_w15976_,
		_w15977_
	);
	LUT3 #(
		.INIT('h2a)
	) name14077 (
		\m5_addr_i[24]_pad ,
		_w8955_,
		_w8956_,
		_w15978_
	);
	LUT3 #(
		.INIT('h80)
	) name14078 (
		\m6_addr_i[24]_pad ,
		_w8955_,
		_w8956_,
		_w15979_
	);
	LUT4 #(
		.INIT('hcedf)
	) name14079 (
		_w8950_,
		_w8953_,
		_w15978_,
		_w15979_,
		_w15980_
	);
	LUT4 #(
		.INIT('h7fff)
	) name14080 (
		_w15971_,
		_w15974_,
		_w15977_,
		_w15980_,
		_w15981_
	);
	LUT3 #(
		.INIT('h80)
	) name14081 (
		\m0_addr_i[25]_pad ,
		_w8955_,
		_w8956_,
		_w15982_
	);
	LUT3 #(
		.INIT('h2a)
	) name14082 (
		\m7_addr_i[25]_pad ,
		_w8955_,
		_w8956_,
		_w15983_
	);
	LUT4 #(
		.INIT('h6e7f)
	) name14083 (
		_w8950_,
		_w8953_,
		_w15982_,
		_w15983_,
		_w15984_
	);
	LUT3 #(
		.INIT('h2a)
	) name14084 (
		\m1_addr_i[25]_pad ,
		_w8955_,
		_w8956_,
		_w15985_
	);
	LUT3 #(
		.INIT('h80)
	) name14085 (
		\m6_addr_i[25]_pad ,
		_w8955_,
		_w8956_,
		_w15986_
	);
	LUT4 #(
		.INIT('h6e7f)
	) name14086 (
		_w8950_,
		_w8953_,
		_w15985_,
		_w15986_,
		_w15987_
	);
	LUT3 #(
		.INIT('h80)
	) name14087 (
		\m2_addr_i[25]_pad ,
		_w8955_,
		_w8956_,
		_w15988_
	);
	LUT3 #(
		.INIT('h2a)
	) name14088 (
		\m5_addr_i[25]_pad ,
		_w8955_,
		_w8956_,
		_w15989_
	);
	LUT4 #(
		.INIT('h9dbf)
	) name14089 (
		_w8950_,
		_w8953_,
		_w15988_,
		_w15989_,
		_w15990_
	);
	LUT3 #(
		.INIT('h2a)
	) name14090 (
		\m3_addr_i[25]_pad ,
		_w8955_,
		_w8956_,
		_w15991_
	);
	LUT3 #(
		.INIT('h80)
	) name14091 (
		\m4_addr_i[25]_pad ,
		_w8955_,
		_w8956_,
		_w15992_
	);
	LUT4 #(
		.INIT('h9dbf)
	) name14092 (
		_w8950_,
		_w8953_,
		_w15991_,
		_w15992_,
		_w15993_
	);
	LUT4 #(
		.INIT('h7fff)
	) name14093 (
		_w15984_,
		_w15987_,
		_w15990_,
		_w15993_,
		_w15994_
	);
	LUT3 #(
		.INIT('h2a)
	) name14094 (
		\m3_addr_i[26]_pad ,
		_w8955_,
		_w8956_,
		_w15995_
	);
	LUT3 #(
		.INIT('h80)
	) name14095 (
		\m4_addr_i[26]_pad ,
		_w8955_,
		_w8956_,
		_w15996_
	);
	LUT4 #(
		.INIT('h9dbf)
	) name14096 (
		_w8950_,
		_w8953_,
		_w15995_,
		_w15996_,
		_w15997_
	);
	LUT3 #(
		.INIT('h2a)
	) name14097 (
		\m5_addr_i[26]_pad ,
		_w8955_,
		_w8956_,
		_w15998_
	);
	LUT3 #(
		.INIT('h80)
	) name14098 (
		\m2_addr_i[26]_pad ,
		_w8955_,
		_w8956_,
		_w15999_
	);
	LUT4 #(
		.INIT('h9bdf)
	) name14099 (
		_w8950_,
		_w8953_,
		_w15998_,
		_w15999_,
		_w16000_
	);
	LUT3 #(
		.INIT('h80)
	) name14100 (
		\m6_addr_i[26]_pad ,
		_w8955_,
		_w8956_,
		_w16001_
	);
	LUT3 #(
		.INIT('h2a)
	) name14101 (
		\m1_addr_i[26]_pad ,
		_w8955_,
		_w8956_,
		_w16002_
	);
	LUT4 #(
		.INIT('h67ef)
	) name14102 (
		_w8950_,
		_w8953_,
		_w16001_,
		_w16002_,
		_w16003_
	);
	LUT3 #(
		.INIT('h80)
	) name14103 (
		\m0_addr_i[26]_pad ,
		_w8955_,
		_w8956_,
		_w16004_
	);
	LUT3 #(
		.INIT('h2a)
	) name14104 (
		\m7_addr_i[26]_pad ,
		_w8955_,
		_w8956_,
		_w16005_
	);
	LUT4 #(
		.INIT('h6e7f)
	) name14105 (
		_w8950_,
		_w8953_,
		_w16004_,
		_w16005_,
		_w16006_
	);
	LUT4 #(
		.INIT('h7fff)
	) name14106 (
		_w15997_,
		_w16000_,
		_w16003_,
		_w16006_,
		_w16007_
	);
	LUT3 #(
		.INIT('h2a)
	) name14107 (
		\m3_addr_i[27]_pad ,
		_w8955_,
		_w8956_,
		_w16008_
	);
	LUT3 #(
		.INIT('h80)
	) name14108 (
		\m4_addr_i[27]_pad ,
		_w8955_,
		_w8956_,
		_w16009_
	);
	LUT4 #(
		.INIT('h9dbf)
	) name14109 (
		_w8950_,
		_w8953_,
		_w16008_,
		_w16009_,
		_w16010_
	);
	LUT3 #(
		.INIT('h2a)
	) name14110 (
		\m5_addr_i[27]_pad ,
		_w8955_,
		_w8956_,
		_w16011_
	);
	LUT3 #(
		.INIT('h2a)
	) name14111 (
		\m7_addr_i[27]_pad ,
		_w8955_,
		_w8956_,
		_w16012_
	);
	LUT4 #(
		.INIT('hcedf)
	) name14112 (
		_w8950_,
		_w8953_,
		_w16011_,
		_w16012_,
		_w16013_
	);
	LUT3 #(
		.INIT('h80)
	) name14113 (
		\m6_addr_i[27]_pad ,
		_w8955_,
		_w8956_,
		_w16014_
	);
	LUT3 #(
		.INIT('h80)
	) name14114 (
		\m0_addr_i[27]_pad ,
		_w8955_,
		_w8956_,
		_w16015_
	);
	LUT4 #(
		.INIT('h67ef)
	) name14115 (
		_w8950_,
		_w8953_,
		_w16014_,
		_w16015_,
		_w16016_
	);
	LUT3 #(
		.INIT('h2a)
	) name14116 (
		\m1_addr_i[27]_pad ,
		_w8955_,
		_w8956_,
		_w16017_
	);
	LUT3 #(
		.INIT('h80)
	) name14117 (
		\m2_addr_i[27]_pad ,
		_w8955_,
		_w8956_,
		_w16018_
	);
	LUT4 #(
		.INIT('h3b7f)
	) name14118 (
		_w8950_,
		_w8953_,
		_w16017_,
		_w16018_,
		_w16019_
	);
	LUT4 #(
		.INIT('h7fff)
	) name14119 (
		_w16010_,
		_w16013_,
		_w16016_,
		_w16019_,
		_w16020_
	);
	LUT3 #(
		.INIT('h2a)
	) name14120 (
		\m3_addr_i[28]_pad ,
		_w8955_,
		_w8956_,
		_w16021_
	);
	LUT3 #(
		.INIT('h80)
	) name14121 (
		\m4_addr_i[28]_pad ,
		_w8955_,
		_w8956_,
		_w16022_
	);
	LUT4 #(
		.INIT('h9dbf)
	) name14122 (
		_w8950_,
		_w8953_,
		_w16021_,
		_w16022_,
		_w16023_
	);
	LUT3 #(
		.INIT('h2a)
	) name14123 (
		\m5_addr_i[28]_pad ,
		_w8955_,
		_w8956_,
		_w16024_
	);
	LUT3 #(
		.INIT('h80)
	) name14124 (
		\m2_addr_i[28]_pad ,
		_w8955_,
		_w8956_,
		_w16025_
	);
	LUT4 #(
		.INIT('h9bdf)
	) name14125 (
		_w8950_,
		_w8953_,
		_w16024_,
		_w16025_,
		_w16026_
	);
	LUT3 #(
		.INIT('h80)
	) name14126 (
		\m6_addr_i[28]_pad ,
		_w8955_,
		_w8956_,
		_w16027_
	);
	LUT3 #(
		.INIT('h2a)
	) name14127 (
		\m1_addr_i[28]_pad ,
		_w8955_,
		_w8956_,
		_w16028_
	);
	LUT4 #(
		.INIT('h67ef)
	) name14128 (
		_w8950_,
		_w8953_,
		_w16027_,
		_w16028_,
		_w16029_
	);
	LUT3 #(
		.INIT('h80)
	) name14129 (
		\m0_addr_i[28]_pad ,
		_w8955_,
		_w8956_,
		_w16030_
	);
	LUT3 #(
		.INIT('h2a)
	) name14130 (
		\m7_addr_i[28]_pad ,
		_w8955_,
		_w8956_,
		_w16031_
	);
	LUT4 #(
		.INIT('h6e7f)
	) name14131 (
		_w8950_,
		_w8953_,
		_w16030_,
		_w16031_,
		_w16032_
	);
	LUT4 #(
		.INIT('h7fff)
	) name14132 (
		_w16023_,
		_w16026_,
		_w16029_,
		_w16032_,
		_w16033_
	);
	LUT3 #(
		.INIT('h2a)
	) name14133 (
		\m5_addr_i[29]_pad ,
		_w8955_,
		_w8956_,
		_w16034_
	);
	LUT3 #(
		.INIT('h80)
	) name14134 (
		\m6_addr_i[29]_pad ,
		_w8955_,
		_w8956_,
		_w16035_
	);
	LUT4 #(
		.INIT('hcedf)
	) name14135 (
		_w8950_,
		_w8953_,
		_w16034_,
		_w16035_,
		_w16036_
	);
	LUT3 #(
		.INIT('h2a)
	) name14136 (
		\m3_addr_i[29]_pad ,
		_w8955_,
		_w8956_,
		_w16037_
	);
	LUT3 #(
		.INIT('h80)
	) name14137 (
		\m2_addr_i[29]_pad ,
		_w8955_,
		_w8956_,
		_w16038_
	);
	LUT3 #(
		.INIT('h57)
	) name14138 (
		_w8974_,
		_w16037_,
		_w16038_,
		_w16039_
	);
	LUT3 #(
		.INIT('h80)
	) name14139 (
		\m4_addr_i[29]_pad ,
		_w8955_,
		_w8956_,
		_w16040_
	);
	LUT3 #(
		.INIT('h2a)
	) name14140 (
		\m1_addr_i[29]_pad ,
		_w8955_,
		_w8956_,
		_w16041_
	);
	LUT4 #(
		.INIT('h57df)
	) name14141 (
		_w8950_,
		_w8953_,
		_w16040_,
		_w16041_,
		_w16042_
	);
	LUT3 #(
		.INIT('h80)
	) name14142 (
		\m0_addr_i[29]_pad ,
		_w8955_,
		_w8956_,
		_w16043_
	);
	LUT3 #(
		.INIT('h2a)
	) name14143 (
		\m7_addr_i[29]_pad ,
		_w8955_,
		_w8956_,
		_w16044_
	);
	LUT4 #(
		.INIT('h6e7f)
	) name14144 (
		_w8950_,
		_w8953_,
		_w16043_,
		_w16044_,
		_w16045_
	);
	LUT4 #(
		.INIT('h7fff)
	) name14145 (
		_w16036_,
		_w16039_,
		_w16042_,
		_w16045_,
		_w16046_
	);
	LUT3 #(
		.INIT('h2a)
	) name14146 (
		\m3_addr_i[2]_pad ,
		_w8955_,
		_w8956_,
		_w16047_
	);
	LUT3 #(
		.INIT('h80)
	) name14147 (
		\m4_addr_i[2]_pad ,
		_w8955_,
		_w8956_,
		_w16048_
	);
	LUT4 #(
		.INIT('h9dbf)
	) name14148 (
		_w8950_,
		_w8953_,
		_w16047_,
		_w16048_,
		_w16049_
	);
	LUT3 #(
		.INIT('h80)
	) name14149 (
		\m0_addr_i[2]_pad ,
		_w8955_,
		_w8956_,
		_w16050_
	);
	LUT3 #(
		.INIT('h2a)
	) name14150 (
		\m5_addr_i[2]_pad ,
		_w8955_,
		_w8956_,
		_w16051_
	);
	LUT4 #(
		.INIT('h5d7f)
	) name14151 (
		_w8950_,
		_w8953_,
		_w16050_,
		_w16051_,
		_w16052_
	);
	LUT3 #(
		.INIT('h2a)
	) name14152 (
		\m7_addr_i[2]_pad ,
		_w8955_,
		_w8956_,
		_w16053_
	);
	LUT3 #(
		.INIT('h80)
	) name14153 (
		\m6_addr_i[2]_pad ,
		_w8955_,
		_w8956_,
		_w16054_
	);
	LUT3 #(
		.INIT('h57)
	) name14154 (
		_w8968_,
		_w16053_,
		_w16054_,
		_w16055_
	);
	LUT3 #(
		.INIT('h2a)
	) name14155 (
		\m1_addr_i[2]_pad ,
		_w8955_,
		_w8956_,
		_w16056_
	);
	LUT3 #(
		.INIT('h80)
	) name14156 (
		\m2_addr_i[2]_pad ,
		_w8955_,
		_w8956_,
		_w16057_
	);
	LUT4 #(
		.INIT('h3b7f)
	) name14157 (
		_w8950_,
		_w8953_,
		_w16056_,
		_w16057_,
		_w16058_
	);
	LUT4 #(
		.INIT('h7fff)
	) name14158 (
		_w16049_,
		_w16052_,
		_w16055_,
		_w16058_,
		_w16059_
	);
	LUT3 #(
		.INIT('h2a)
	) name14159 (
		\m1_addr_i[30]_pad ,
		_w8955_,
		_w8956_,
		_w16060_
	);
	LUT3 #(
		.INIT('h80)
	) name14160 (
		\m2_addr_i[30]_pad ,
		_w8955_,
		_w8956_,
		_w16061_
	);
	LUT4 #(
		.INIT('h3b7f)
	) name14161 (
		_w8950_,
		_w8953_,
		_w16060_,
		_w16061_,
		_w16062_
	);
	LUT3 #(
		.INIT('h80)
	) name14162 (
		\m0_addr_i[30]_pad ,
		_w8955_,
		_w8956_,
		_w16063_
	);
	LUT3 #(
		.INIT('h80)
	) name14163 (
		\m6_addr_i[30]_pad ,
		_w8955_,
		_w8956_,
		_w16064_
	);
	LUT4 #(
		.INIT('h6e7f)
	) name14164 (
		_w8950_,
		_w8953_,
		_w16063_,
		_w16064_,
		_w16065_
	);
	LUT3 #(
		.INIT('h2a)
	) name14165 (
		\m7_addr_i[30]_pad ,
		_w8955_,
		_w8956_,
		_w16066_
	);
	LUT3 #(
		.INIT('h2a)
	) name14166 (
		\m5_addr_i[30]_pad ,
		_w8955_,
		_w8956_,
		_w16067_
	);
	LUT4 #(
		.INIT('hcdef)
	) name14167 (
		_w8950_,
		_w8953_,
		_w16066_,
		_w16067_,
		_w16068_
	);
	LUT3 #(
		.INIT('h2a)
	) name14168 (
		\m3_addr_i[30]_pad ,
		_w8955_,
		_w8956_,
		_w16069_
	);
	LUT3 #(
		.INIT('h80)
	) name14169 (
		\m4_addr_i[30]_pad ,
		_w8955_,
		_w8956_,
		_w16070_
	);
	LUT4 #(
		.INIT('h9dbf)
	) name14170 (
		_w8950_,
		_w8953_,
		_w16069_,
		_w16070_,
		_w16071_
	);
	LUT4 #(
		.INIT('h7fff)
	) name14171 (
		_w16062_,
		_w16065_,
		_w16068_,
		_w16071_,
		_w16072_
	);
	LUT3 #(
		.INIT('h80)
	) name14172 (
		\m0_addr_i[31]_pad ,
		_w8955_,
		_w8956_,
		_w16073_
	);
	LUT3 #(
		.INIT('h2a)
	) name14173 (
		\m7_addr_i[31]_pad ,
		_w8955_,
		_w8956_,
		_w16074_
	);
	LUT4 #(
		.INIT('h6e7f)
	) name14174 (
		_w8950_,
		_w8953_,
		_w16073_,
		_w16074_,
		_w16075_
	);
	LUT3 #(
		.INIT('h2a)
	) name14175 (
		\m1_addr_i[31]_pad ,
		_w8955_,
		_w8956_,
		_w16076_
	);
	LUT3 #(
		.INIT('h80)
	) name14176 (
		\m6_addr_i[31]_pad ,
		_w8955_,
		_w8956_,
		_w16077_
	);
	LUT4 #(
		.INIT('h6e7f)
	) name14177 (
		_w8950_,
		_w8953_,
		_w16076_,
		_w16077_,
		_w16078_
	);
	LUT3 #(
		.INIT('h80)
	) name14178 (
		\m2_addr_i[31]_pad ,
		_w8955_,
		_w8956_,
		_w16079_
	);
	LUT3 #(
		.INIT('h2a)
	) name14179 (
		\m5_addr_i[31]_pad ,
		_w8955_,
		_w8956_,
		_w16080_
	);
	LUT4 #(
		.INIT('h9dbf)
	) name14180 (
		_w8950_,
		_w8953_,
		_w16079_,
		_w16080_,
		_w16081_
	);
	LUT3 #(
		.INIT('h2a)
	) name14181 (
		\m3_addr_i[31]_pad ,
		_w8955_,
		_w8956_,
		_w16082_
	);
	LUT3 #(
		.INIT('h80)
	) name14182 (
		\m4_addr_i[31]_pad ,
		_w8955_,
		_w8956_,
		_w16083_
	);
	LUT4 #(
		.INIT('h9dbf)
	) name14183 (
		_w8950_,
		_w8953_,
		_w16082_,
		_w16083_,
		_w16084_
	);
	LUT4 #(
		.INIT('h7fff)
	) name14184 (
		_w16075_,
		_w16078_,
		_w16081_,
		_w16084_,
		_w16085_
	);
	LUT3 #(
		.INIT('h80)
	) name14185 (
		\m0_addr_i[3]_pad ,
		_w8955_,
		_w8956_,
		_w16086_
	);
	LUT3 #(
		.INIT('h2a)
	) name14186 (
		\m7_addr_i[3]_pad ,
		_w8955_,
		_w8956_,
		_w16087_
	);
	LUT4 #(
		.INIT('h6e7f)
	) name14187 (
		_w8950_,
		_w8953_,
		_w16086_,
		_w16087_,
		_w16088_
	);
	LUT3 #(
		.INIT('h2a)
	) name14188 (
		\m1_addr_i[3]_pad ,
		_w8955_,
		_w8956_,
		_w16089_
	);
	LUT3 #(
		.INIT('h80)
	) name14189 (
		\m4_addr_i[3]_pad ,
		_w8955_,
		_w8956_,
		_w16090_
	);
	LUT4 #(
		.INIT('h5d7f)
	) name14190 (
		_w8950_,
		_w8953_,
		_w16089_,
		_w16090_,
		_w16091_
	);
	LUT3 #(
		.INIT('h80)
	) name14191 (
		\m2_addr_i[3]_pad ,
		_w8955_,
		_w8956_,
		_w16092_
	);
	LUT3 #(
		.INIT('h2a)
	) name14192 (
		\m3_addr_i[3]_pad ,
		_w8955_,
		_w8956_,
		_w16093_
	);
	LUT3 #(
		.INIT('h57)
	) name14193 (
		_w8974_,
		_w16092_,
		_w16093_,
		_w16094_
	);
	LUT3 #(
		.INIT('h80)
	) name14194 (
		\m6_addr_i[3]_pad ,
		_w8955_,
		_w8956_,
		_w16095_
	);
	LUT3 #(
		.INIT('h2a)
	) name14195 (
		\m5_addr_i[3]_pad ,
		_w8955_,
		_w8956_,
		_w16096_
	);
	LUT4 #(
		.INIT('hcdef)
	) name14196 (
		_w8950_,
		_w8953_,
		_w16095_,
		_w16096_,
		_w16097_
	);
	LUT4 #(
		.INIT('h7fff)
	) name14197 (
		_w16088_,
		_w16091_,
		_w16094_,
		_w16097_,
		_w16098_
	);
	LUT3 #(
		.INIT('h2a)
	) name14198 (
		\m1_addr_i[4]_pad ,
		_w8955_,
		_w8956_,
		_w16099_
	);
	LUT3 #(
		.INIT('h80)
	) name14199 (
		\m2_addr_i[4]_pad ,
		_w8955_,
		_w8956_,
		_w16100_
	);
	LUT4 #(
		.INIT('h3b7f)
	) name14200 (
		_w8950_,
		_w8953_,
		_w16099_,
		_w16100_,
		_w16101_
	);
	LUT3 #(
		.INIT('h80)
	) name14201 (
		\m6_addr_i[4]_pad ,
		_w8955_,
		_w8956_,
		_w16102_
	);
	LUT3 #(
		.INIT('h2a)
	) name14202 (
		\m7_addr_i[4]_pad ,
		_w8955_,
		_w8956_,
		_w16103_
	);
	LUT3 #(
		.INIT('h57)
	) name14203 (
		_w8968_,
		_w16102_,
		_w16103_,
		_w16104_
	);
	LUT3 #(
		.INIT('h2a)
	) name14204 (
		\m5_addr_i[4]_pad ,
		_w8955_,
		_w8956_,
		_w16105_
	);
	LUT3 #(
		.INIT('h80)
	) name14205 (
		\m0_addr_i[4]_pad ,
		_w8955_,
		_w8956_,
		_w16106_
	);
	LUT4 #(
		.INIT('h57df)
	) name14206 (
		_w8950_,
		_w8953_,
		_w16105_,
		_w16106_,
		_w16107_
	);
	LUT3 #(
		.INIT('h2a)
	) name14207 (
		\m3_addr_i[4]_pad ,
		_w8955_,
		_w8956_,
		_w16108_
	);
	LUT3 #(
		.INIT('h80)
	) name14208 (
		\m4_addr_i[4]_pad ,
		_w8955_,
		_w8956_,
		_w16109_
	);
	LUT4 #(
		.INIT('h9dbf)
	) name14209 (
		_w8950_,
		_w8953_,
		_w16108_,
		_w16109_,
		_w16110_
	);
	LUT4 #(
		.INIT('h7fff)
	) name14210 (
		_w16101_,
		_w16104_,
		_w16107_,
		_w16110_,
		_w16111_
	);
	LUT3 #(
		.INIT('h2a)
	) name14211 (
		\m3_addr_i[5]_pad ,
		_w8955_,
		_w8956_,
		_w16112_
	);
	LUT3 #(
		.INIT('h80)
	) name14212 (
		\m4_addr_i[5]_pad ,
		_w8955_,
		_w8956_,
		_w16113_
	);
	LUT4 #(
		.INIT('h9dbf)
	) name14213 (
		_w8950_,
		_w8953_,
		_w16112_,
		_w16113_,
		_w16114_
	);
	LUT3 #(
		.INIT('h80)
	) name14214 (
		\m0_addr_i[5]_pad ,
		_w8955_,
		_w8956_,
		_w16115_
	);
	LUT3 #(
		.INIT('h2a)
	) name14215 (
		\m5_addr_i[5]_pad ,
		_w8955_,
		_w8956_,
		_w16116_
	);
	LUT4 #(
		.INIT('h5d7f)
	) name14216 (
		_w8950_,
		_w8953_,
		_w16115_,
		_w16116_,
		_w16117_
	);
	LUT3 #(
		.INIT('h2a)
	) name14217 (
		\m7_addr_i[5]_pad ,
		_w8955_,
		_w8956_,
		_w16118_
	);
	LUT3 #(
		.INIT('h80)
	) name14218 (
		\m6_addr_i[5]_pad ,
		_w8955_,
		_w8956_,
		_w16119_
	);
	LUT3 #(
		.INIT('h57)
	) name14219 (
		_w8968_,
		_w16118_,
		_w16119_,
		_w16120_
	);
	LUT3 #(
		.INIT('h2a)
	) name14220 (
		\m1_addr_i[5]_pad ,
		_w8955_,
		_w8956_,
		_w16121_
	);
	LUT3 #(
		.INIT('h80)
	) name14221 (
		\m2_addr_i[5]_pad ,
		_w8955_,
		_w8956_,
		_w16122_
	);
	LUT4 #(
		.INIT('h3b7f)
	) name14222 (
		_w8950_,
		_w8953_,
		_w16121_,
		_w16122_,
		_w16123_
	);
	LUT4 #(
		.INIT('h7fff)
	) name14223 (
		_w16114_,
		_w16117_,
		_w16120_,
		_w16123_,
		_w16124_
	);
	LUT3 #(
		.INIT('h2a)
	) name14224 (
		\m3_addr_i[6]_pad ,
		_w8955_,
		_w8956_,
		_w16125_
	);
	LUT3 #(
		.INIT('h80)
	) name14225 (
		\m4_addr_i[6]_pad ,
		_w8955_,
		_w8956_,
		_w16126_
	);
	LUT4 #(
		.INIT('h9dbf)
	) name14226 (
		_w8950_,
		_w8953_,
		_w16125_,
		_w16126_,
		_w16127_
	);
	LUT3 #(
		.INIT('h2a)
	) name14227 (
		\m1_addr_i[6]_pad ,
		_w8955_,
		_w8956_,
		_w16128_
	);
	LUT3 #(
		.INIT('h2a)
	) name14228 (
		\m7_addr_i[6]_pad ,
		_w8955_,
		_w8956_,
		_w16129_
	);
	LUT4 #(
		.INIT('h6e7f)
	) name14229 (
		_w8950_,
		_w8953_,
		_w16128_,
		_w16129_,
		_w16130_
	);
	LUT3 #(
		.INIT('h80)
	) name14230 (
		\m2_addr_i[6]_pad ,
		_w8955_,
		_w8956_,
		_w16131_
	);
	LUT3 #(
		.INIT('h80)
	) name14231 (
		\m0_addr_i[6]_pad ,
		_w8955_,
		_w8956_,
		_w16132_
	);
	LUT4 #(
		.INIT('h37bf)
	) name14232 (
		_w8950_,
		_w8953_,
		_w16131_,
		_w16132_,
		_w16133_
	);
	LUT3 #(
		.INIT('h80)
	) name14233 (
		\m6_addr_i[6]_pad ,
		_w8955_,
		_w8956_,
		_w16134_
	);
	LUT3 #(
		.INIT('h2a)
	) name14234 (
		\m5_addr_i[6]_pad ,
		_w8955_,
		_w8956_,
		_w16135_
	);
	LUT4 #(
		.INIT('hcdef)
	) name14235 (
		_w8950_,
		_w8953_,
		_w16134_,
		_w16135_,
		_w16136_
	);
	LUT4 #(
		.INIT('h7fff)
	) name14236 (
		_w16127_,
		_w16130_,
		_w16133_,
		_w16136_,
		_w16137_
	);
	LUT3 #(
		.INIT('h2a)
	) name14237 (
		\m3_addr_i[7]_pad ,
		_w8955_,
		_w8956_,
		_w16138_
	);
	LUT3 #(
		.INIT('h80)
	) name14238 (
		\m4_addr_i[7]_pad ,
		_w8955_,
		_w8956_,
		_w16139_
	);
	LUT4 #(
		.INIT('h9dbf)
	) name14239 (
		_w8950_,
		_w8953_,
		_w16138_,
		_w16139_,
		_w16140_
	);
	LUT3 #(
		.INIT('h80)
	) name14240 (
		\m6_addr_i[7]_pad ,
		_w8955_,
		_w8956_,
		_w16141_
	);
	LUT3 #(
		.INIT('h80)
	) name14241 (
		\m2_addr_i[7]_pad ,
		_w8955_,
		_w8956_,
		_w16142_
	);
	LUT4 #(
		.INIT('habef)
	) name14242 (
		_w8950_,
		_w8953_,
		_w16141_,
		_w16142_,
		_w16143_
	);
	LUT3 #(
		.INIT('h2a)
	) name14243 (
		\m5_addr_i[7]_pad ,
		_w8955_,
		_w8956_,
		_w16144_
	);
	LUT3 #(
		.INIT('h2a)
	) name14244 (
		\m1_addr_i[7]_pad ,
		_w8955_,
		_w8956_,
		_w16145_
	);
	LUT4 #(
		.INIT('h57df)
	) name14245 (
		_w8950_,
		_w8953_,
		_w16144_,
		_w16145_,
		_w16146_
	);
	LUT3 #(
		.INIT('h80)
	) name14246 (
		\m0_addr_i[7]_pad ,
		_w8955_,
		_w8956_,
		_w16147_
	);
	LUT3 #(
		.INIT('h2a)
	) name14247 (
		\m7_addr_i[7]_pad ,
		_w8955_,
		_w8956_,
		_w16148_
	);
	LUT4 #(
		.INIT('h6e7f)
	) name14248 (
		_w8950_,
		_w8953_,
		_w16147_,
		_w16148_,
		_w16149_
	);
	LUT4 #(
		.INIT('h7fff)
	) name14249 (
		_w16140_,
		_w16143_,
		_w16146_,
		_w16149_,
		_w16150_
	);
	LUT3 #(
		.INIT('h80)
	) name14250 (
		\m6_addr_i[8]_pad ,
		_w8955_,
		_w8956_,
		_w16151_
	);
	LUT3 #(
		.INIT('h2a)
	) name14251 (
		\m5_addr_i[8]_pad ,
		_w8955_,
		_w8956_,
		_w16152_
	);
	LUT4 #(
		.INIT('hcdef)
	) name14252 (
		_w8950_,
		_w8953_,
		_w16151_,
		_w16152_,
		_w16153_
	);
	LUT3 #(
		.INIT('h80)
	) name14253 (
		\m0_addr_i[8]_pad ,
		_w8955_,
		_w8956_,
		_w16154_
	);
	LUT3 #(
		.INIT('h80)
	) name14254 (
		\m4_addr_i[8]_pad ,
		_w8955_,
		_w8956_,
		_w16155_
	);
	LUT4 #(
		.INIT('h5d7f)
	) name14255 (
		_w8950_,
		_w8953_,
		_w16154_,
		_w16155_,
		_w16156_
	);
	LUT3 #(
		.INIT('h2a)
	) name14256 (
		\m7_addr_i[8]_pad ,
		_w8955_,
		_w8956_,
		_w16157_
	);
	LUT3 #(
		.INIT('h2a)
	) name14257 (
		\m3_addr_i[8]_pad ,
		_w8955_,
		_w8956_,
		_w16158_
	);
	LUT4 #(
		.INIT('habef)
	) name14258 (
		_w8950_,
		_w8953_,
		_w16157_,
		_w16158_,
		_w16159_
	);
	LUT3 #(
		.INIT('h2a)
	) name14259 (
		\m1_addr_i[8]_pad ,
		_w8955_,
		_w8956_,
		_w16160_
	);
	LUT3 #(
		.INIT('h80)
	) name14260 (
		\m2_addr_i[8]_pad ,
		_w8955_,
		_w8956_,
		_w16161_
	);
	LUT4 #(
		.INIT('h3b7f)
	) name14261 (
		_w8950_,
		_w8953_,
		_w16160_,
		_w16161_,
		_w16162_
	);
	LUT4 #(
		.INIT('h7fff)
	) name14262 (
		_w16153_,
		_w16156_,
		_w16159_,
		_w16162_,
		_w16163_
	);
	LUT3 #(
		.INIT('h2a)
	) name14263 (
		\m1_addr_i[9]_pad ,
		_w8955_,
		_w8956_,
		_w16164_
	);
	LUT3 #(
		.INIT('h80)
	) name14264 (
		\m2_addr_i[9]_pad ,
		_w8955_,
		_w8956_,
		_w16165_
	);
	LUT4 #(
		.INIT('h3b7f)
	) name14265 (
		_w8950_,
		_w8953_,
		_w16164_,
		_w16165_,
		_w16166_
	);
	LUT3 #(
		.INIT('h2a)
	) name14266 (
		\m3_addr_i[9]_pad ,
		_w8955_,
		_w8956_,
		_w16167_
	);
	LUT3 #(
		.INIT('h2a)
	) name14267 (
		\m5_addr_i[9]_pad ,
		_w8955_,
		_w8956_,
		_w16168_
	);
	LUT4 #(
		.INIT('h9dbf)
	) name14268 (
		_w8950_,
		_w8953_,
		_w16167_,
		_w16168_,
		_w16169_
	);
	LUT3 #(
		.INIT('h80)
	) name14269 (
		\m4_addr_i[9]_pad ,
		_w8955_,
		_w8956_,
		_w16170_
	);
	LUT3 #(
		.INIT('h80)
	) name14270 (
		\m6_addr_i[9]_pad ,
		_w8955_,
		_w8956_,
		_w16171_
	);
	LUT4 #(
		.INIT('hcedf)
	) name14271 (
		_w8950_,
		_w8953_,
		_w16170_,
		_w16171_,
		_w16172_
	);
	LUT3 #(
		.INIT('h80)
	) name14272 (
		\m0_addr_i[9]_pad ,
		_w8955_,
		_w8956_,
		_w16173_
	);
	LUT3 #(
		.INIT('h2a)
	) name14273 (
		\m7_addr_i[9]_pad ,
		_w8955_,
		_w8956_,
		_w16174_
	);
	LUT4 #(
		.INIT('h6e7f)
	) name14274 (
		_w8950_,
		_w8953_,
		_w16173_,
		_w16174_,
		_w16175_
	);
	LUT4 #(
		.INIT('h7fff)
	) name14275 (
		_w16166_,
		_w16169_,
		_w16172_,
		_w16175_,
		_w16176_
	);
	LUT3 #(
		.INIT('h80)
	) name14276 (
		\m0_data_i[0]_pad ,
		_w8955_,
		_w8956_,
		_w16177_
	);
	LUT3 #(
		.INIT('h2a)
	) name14277 (
		\m7_data_i[0]_pad ,
		_w8955_,
		_w8956_,
		_w16178_
	);
	LUT4 #(
		.INIT('h6e7f)
	) name14278 (
		_w8950_,
		_w8953_,
		_w16177_,
		_w16178_,
		_w16179_
	);
	LUT3 #(
		.INIT('h80)
	) name14279 (
		\m6_data_i[0]_pad ,
		_w8955_,
		_w8956_,
		_w16180_
	);
	LUT3 #(
		.INIT('h80)
	) name14280 (
		\m2_data_i[0]_pad ,
		_w8955_,
		_w8956_,
		_w16181_
	);
	LUT4 #(
		.INIT('habef)
	) name14281 (
		_w8950_,
		_w8953_,
		_w16180_,
		_w16181_,
		_w16182_
	);
	LUT3 #(
		.INIT('h2a)
	) name14282 (
		\m5_data_i[0]_pad ,
		_w8955_,
		_w8956_,
		_w16183_
	);
	LUT3 #(
		.INIT('h2a)
	) name14283 (
		\m1_data_i[0]_pad ,
		_w8955_,
		_w8956_,
		_w16184_
	);
	LUT4 #(
		.INIT('h57df)
	) name14284 (
		_w8950_,
		_w8953_,
		_w16183_,
		_w16184_,
		_w16185_
	);
	LUT3 #(
		.INIT('h2a)
	) name14285 (
		\m3_data_i[0]_pad ,
		_w8955_,
		_w8956_,
		_w16186_
	);
	LUT3 #(
		.INIT('h80)
	) name14286 (
		\m4_data_i[0]_pad ,
		_w8955_,
		_w8956_,
		_w16187_
	);
	LUT4 #(
		.INIT('h9dbf)
	) name14287 (
		_w8950_,
		_w8953_,
		_w16186_,
		_w16187_,
		_w16188_
	);
	LUT4 #(
		.INIT('h7fff)
	) name14288 (
		_w16179_,
		_w16182_,
		_w16185_,
		_w16188_,
		_w16189_
	);
	LUT3 #(
		.INIT('h2a)
	) name14289 (
		\m1_data_i[10]_pad ,
		_w8955_,
		_w8956_,
		_w16190_
	);
	LUT3 #(
		.INIT('h80)
	) name14290 (
		\m2_data_i[10]_pad ,
		_w8955_,
		_w8956_,
		_w16191_
	);
	LUT4 #(
		.INIT('h3b7f)
	) name14291 (
		_w8950_,
		_w8953_,
		_w16190_,
		_w16191_,
		_w16192_
	);
	LUT3 #(
		.INIT('h80)
	) name14292 (
		\m0_data_i[10]_pad ,
		_w8955_,
		_w8956_,
		_w16193_
	);
	LUT3 #(
		.INIT('h80)
	) name14293 (
		\m4_data_i[10]_pad ,
		_w8955_,
		_w8956_,
		_w16194_
	);
	LUT4 #(
		.INIT('h5d7f)
	) name14294 (
		_w8950_,
		_w8953_,
		_w16193_,
		_w16194_,
		_w16195_
	);
	LUT3 #(
		.INIT('h2a)
	) name14295 (
		\m7_data_i[10]_pad ,
		_w8955_,
		_w8956_,
		_w16196_
	);
	LUT3 #(
		.INIT('h2a)
	) name14296 (
		\m3_data_i[10]_pad ,
		_w8955_,
		_w8956_,
		_w16197_
	);
	LUT4 #(
		.INIT('habef)
	) name14297 (
		_w8950_,
		_w8953_,
		_w16196_,
		_w16197_,
		_w16198_
	);
	LUT3 #(
		.INIT('h80)
	) name14298 (
		\m6_data_i[10]_pad ,
		_w8955_,
		_w8956_,
		_w16199_
	);
	LUT3 #(
		.INIT('h2a)
	) name14299 (
		\m5_data_i[10]_pad ,
		_w8955_,
		_w8956_,
		_w16200_
	);
	LUT4 #(
		.INIT('hcdef)
	) name14300 (
		_w8950_,
		_w8953_,
		_w16199_,
		_w16200_,
		_w16201_
	);
	LUT4 #(
		.INIT('h7fff)
	) name14301 (
		_w16192_,
		_w16195_,
		_w16198_,
		_w16201_,
		_w16202_
	);
	LUT3 #(
		.INIT('h2a)
	) name14302 (
		\m3_data_i[11]_pad ,
		_w8955_,
		_w8956_,
		_w16203_
	);
	LUT3 #(
		.INIT('h80)
	) name14303 (
		\m4_data_i[11]_pad ,
		_w8955_,
		_w8956_,
		_w16204_
	);
	LUT4 #(
		.INIT('h9dbf)
	) name14304 (
		_w8950_,
		_w8953_,
		_w16203_,
		_w16204_,
		_w16205_
	);
	LUT3 #(
		.INIT('h80)
	) name14305 (
		\m0_data_i[11]_pad ,
		_w8955_,
		_w8956_,
		_w16206_
	);
	LUT3 #(
		.INIT('h80)
	) name14306 (
		\m2_data_i[11]_pad ,
		_w8955_,
		_w8956_,
		_w16207_
	);
	LUT4 #(
		.INIT('h3b7f)
	) name14307 (
		_w8950_,
		_w8953_,
		_w16206_,
		_w16207_,
		_w16208_
	);
	LUT3 #(
		.INIT('h2a)
	) name14308 (
		\m7_data_i[11]_pad ,
		_w8955_,
		_w8956_,
		_w16209_
	);
	LUT3 #(
		.INIT('h2a)
	) name14309 (
		\m1_data_i[11]_pad ,
		_w8955_,
		_w8956_,
		_w16210_
	);
	LUT4 #(
		.INIT('h67ef)
	) name14310 (
		_w8950_,
		_w8953_,
		_w16209_,
		_w16210_,
		_w16211_
	);
	LUT3 #(
		.INIT('h80)
	) name14311 (
		\m6_data_i[11]_pad ,
		_w8955_,
		_w8956_,
		_w16212_
	);
	LUT3 #(
		.INIT('h2a)
	) name14312 (
		\m5_data_i[11]_pad ,
		_w8955_,
		_w8956_,
		_w16213_
	);
	LUT4 #(
		.INIT('hcdef)
	) name14313 (
		_w8950_,
		_w8953_,
		_w16212_,
		_w16213_,
		_w16214_
	);
	LUT4 #(
		.INIT('h7fff)
	) name14314 (
		_w16205_,
		_w16208_,
		_w16211_,
		_w16214_,
		_w16215_
	);
	LUT3 #(
		.INIT('h2a)
	) name14315 (
		\m1_data_i[12]_pad ,
		_w8955_,
		_w8956_,
		_w16216_
	);
	LUT3 #(
		.INIT('h80)
	) name14316 (
		\m2_data_i[12]_pad ,
		_w8955_,
		_w8956_,
		_w16217_
	);
	LUT4 #(
		.INIT('h3b7f)
	) name14317 (
		_w8950_,
		_w8953_,
		_w16216_,
		_w16217_,
		_w16218_
	);
	LUT3 #(
		.INIT('h80)
	) name14318 (
		\m0_data_i[12]_pad ,
		_w8955_,
		_w8956_,
		_w16219_
	);
	LUT3 #(
		.INIT('h80)
	) name14319 (
		\m4_data_i[12]_pad ,
		_w8955_,
		_w8956_,
		_w16220_
	);
	LUT4 #(
		.INIT('h5d7f)
	) name14320 (
		_w8950_,
		_w8953_,
		_w16219_,
		_w16220_,
		_w16221_
	);
	LUT3 #(
		.INIT('h2a)
	) name14321 (
		\m7_data_i[12]_pad ,
		_w8955_,
		_w8956_,
		_w16222_
	);
	LUT3 #(
		.INIT('h2a)
	) name14322 (
		\m3_data_i[12]_pad ,
		_w8955_,
		_w8956_,
		_w16223_
	);
	LUT4 #(
		.INIT('habef)
	) name14323 (
		_w8950_,
		_w8953_,
		_w16222_,
		_w16223_,
		_w16224_
	);
	LUT3 #(
		.INIT('h80)
	) name14324 (
		\m6_data_i[12]_pad ,
		_w8955_,
		_w8956_,
		_w16225_
	);
	LUT3 #(
		.INIT('h2a)
	) name14325 (
		\m5_data_i[12]_pad ,
		_w8955_,
		_w8956_,
		_w16226_
	);
	LUT4 #(
		.INIT('hcdef)
	) name14326 (
		_w8950_,
		_w8953_,
		_w16225_,
		_w16226_,
		_w16227_
	);
	LUT4 #(
		.INIT('h7fff)
	) name14327 (
		_w16218_,
		_w16221_,
		_w16224_,
		_w16227_,
		_w16228_
	);
	LUT3 #(
		.INIT('h2a)
	) name14328 (
		\m1_data_i[13]_pad ,
		_w8955_,
		_w8956_,
		_w16229_
	);
	LUT3 #(
		.INIT('h80)
	) name14329 (
		\m2_data_i[13]_pad ,
		_w8955_,
		_w8956_,
		_w16230_
	);
	LUT4 #(
		.INIT('h3b7f)
	) name14330 (
		_w8950_,
		_w8953_,
		_w16229_,
		_w16230_,
		_w16231_
	);
	LUT3 #(
		.INIT('h80)
	) name14331 (
		\m0_data_i[13]_pad ,
		_w8955_,
		_w8956_,
		_w16232_
	);
	LUT3 #(
		.INIT('h2a)
	) name14332 (
		\m5_data_i[13]_pad ,
		_w8955_,
		_w8956_,
		_w16233_
	);
	LUT4 #(
		.INIT('h5d7f)
	) name14333 (
		_w8950_,
		_w8953_,
		_w16232_,
		_w16233_,
		_w16234_
	);
	LUT3 #(
		.INIT('h2a)
	) name14334 (
		\m7_data_i[13]_pad ,
		_w8955_,
		_w8956_,
		_w16235_
	);
	LUT3 #(
		.INIT('h80)
	) name14335 (
		\m6_data_i[13]_pad ,
		_w8955_,
		_w8956_,
		_w16236_
	);
	LUT3 #(
		.INIT('h57)
	) name14336 (
		_w8968_,
		_w16235_,
		_w16236_,
		_w16237_
	);
	LUT3 #(
		.INIT('h2a)
	) name14337 (
		\m3_data_i[13]_pad ,
		_w8955_,
		_w8956_,
		_w16238_
	);
	LUT3 #(
		.INIT('h80)
	) name14338 (
		\m4_data_i[13]_pad ,
		_w8955_,
		_w8956_,
		_w16239_
	);
	LUT4 #(
		.INIT('h9dbf)
	) name14339 (
		_w8950_,
		_w8953_,
		_w16238_,
		_w16239_,
		_w16240_
	);
	LUT4 #(
		.INIT('h7fff)
	) name14340 (
		_w16231_,
		_w16234_,
		_w16237_,
		_w16240_,
		_w16241_
	);
	LUT3 #(
		.INIT('h2a)
	) name14341 (
		\m1_data_i[14]_pad ,
		_w8955_,
		_w8956_,
		_w16242_
	);
	LUT3 #(
		.INIT('h80)
	) name14342 (
		\m2_data_i[14]_pad ,
		_w8955_,
		_w8956_,
		_w16243_
	);
	LUT4 #(
		.INIT('h3b7f)
	) name14343 (
		_w8950_,
		_w8953_,
		_w16242_,
		_w16243_,
		_w16244_
	);
	LUT3 #(
		.INIT('h80)
	) name14344 (
		\m0_data_i[14]_pad ,
		_w8955_,
		_w8956_,
		_w16245_
	);
	LUT3 #(
		.INIT('h2a)
	) name14345 (
		\m5_data_i[14]_pad ,
		_w8955_,
		_w8956_,
		_w16246_
	);
	LUT4 #(
		.INIT('h5d7f)
	) name14346 (
		_w8950_,
		_w8953_,
		_w16245_,
		_w16246_,
		_w16247_
	);
	LUT3 #(
		.INIT('h2a)
	) name14347 (
		\m7_data_i[14]_pad ,
		_w8955_,
		_w8956_,
		_w16248_
	);
	LUT3 #(
		.INIT('h80)
	) name14348 (
		\m6_data_i[14]_pad ,
		_w8955_,
		_w8956_,
		_w16249_
	);
	LUT3 #(
		.INIT('h57)
	) name14349 (
		_w8968_,
		_w16248_,
		_w16249_,
		_w16250_
	);
	LUT3 #(
		.INIT('h2a)
	) name14350 (
		\m3_data_i[14]_pad ,
		_w8955_,
		_w8956_,
		_w16251_
	);
	LUT3 #(
		.INIT('h80)
	) name14351 (
		\m4_data_i[14]_pad ,
		_w8955_,
		_w8956_,
		_w16252_
	);
	LUT4 #(
		.INIT('h9dbf)
	) name14352 (
		_w8950_,
		_w8953_,
		_w16251_,
		_w16252_,
		_w16253_
	);
	LUT4 #(
		.INIT('h7fff)
	) name14353 (
		_w16244_,
		_w16247_,
		_w16250_,
		_w16253_,
		_w16254_
	);
	LUT3 #(
		.INIT('h2a)
	) name14354 (
		\m3_data_i[15]_pad ,
		_w8955_,
		_w8956_,
		_w16255_
	);
	LUT3 #(
		.INIT('h80)
	) name14355 (
		\m4_data_i[15]_pad ,
		_w8955_,
		_w8956_,
		_w16256_
	);
	LUT4 #(
		.INIT('h9dbf)
	) name14356 (
		_w8950_,
		_w8953_,
		_w16255_,
		_w16256_,
		_w16257_
	);
	LUT3 #(
		.INIT('h2a)
	) name14357 (
		\m1_data_i[15]_pad ,
		_w8955_,
		_w8956_,
		_w16258_
	);
	LUT3 #(
		.INIT('h2a)
	) name14358 (
		\m5_data_i[15]_pad ,
		_w8955_,
		_w8956_,
		_w16259_
	);
	LUT4 #(
		.INIT('h5d7f)
	) name14359 (
		_w8950_,
		_w8953_,
		_w16258_,
		_w16259_,
		_w16260_
	);
	LUT3 #(
		.INIT('h80)
	) name14360 (
		\m2_data_i[15]_pad ,
		_w8955_,
		_w8956_,
		_w16261_
	);
	LUT3 #(
		.INIT('h80)
	) name14361 (
		\m6_data_i[15]_pad ,
		_w8955_,
		_w8956_,
		_w16262_
	);
	LUT4 #(
		.INIT('haebf)
	) name14362 (
		_w8950_,
		_w8953_,
		_w16261_,
		_w16262_,
		_w16263_
	);
	LUT3 #(
		.INIT('h80)
	) name14363 (
		\m0_data_i[15]_pad ,
		_w8955_,
		_w8956_,
		_w16264_
	);
	LUT3 #(
		.INIT('h2a)
	) name14364 (
		\m7_data_i[15]_pad ,
		_w8955_,
		_w8956_,
		_w16265_
	);
	LUT4 #(
		.INIT('h6e7f)
	) name14365 (
		_w8950_,
		_w8953_,
		_w16264_,
		_w16265_,
		_w16266_
	);
	LUT4 #(
		.INIT('h7fff)
	) name14366 (
		_w16257_,
		_w16260_,
		_w16263_,
		_w16266_,
		_w16267_
	);
	LUT3 #(
		.INIT('h2a)
	) name14367 (
		\m1_data_i[16]_pad ,
		_w8955_,
		_w8956_,
		_w16268_
	);
	LUT3 #(
		.INIT('h80)
	) name14368 (
		\m2_data_i[16]_pad ,
		_w8955_,
		_w8956_,
		_w16269_
	);
	LUT4 #(
		.INIT('h3b7f)
	) name14369 (
		_w8950_,
		_w8953_,
		_w16268_,
		_w16269_,
		_w16270_
	);
	LUT3 #(
		.INIT('h80)
	) name14370 (
		\m0_data_i[16]_pad ,
		_w8955_,
		_w8956_,
		_w16271_
	);
	LUT3 #(
		.INIT('h80)
	) name14371 (
		\m4_data_i[16]_pad ,
		_w8955_,
		_w8956_,
		_w16272_
	);
	LUT4 #(
		.INIT('h5d7f)
	) name14372 (
		_w8950_,
		_w8953_,
		_w16271_,
		_w16272_,
		_w16273_
	);
	LUT3 #(
		.INIT('h2a)
	) name14373 (
		\m7_data_i[16]_pad ,
		_w8955_,
		_w8956_,
		_w16274_
	);
	LUT3 #(
		.INIT('h2a)
	) name14374 (
		\m3_data_i[16]_pad ,
		_w8955_,
		_w8956_,
		_w16275_
	);
	LUT4 #(
		.INIT('habef)
	) name14375 (
		_w8950_,
		_w8953_,
		_w16274_,
		_w16275_,
		_w16276_
	);
	LUT3 #(
		.INIT('h80)
	) name14376 (
		\m6_data_i[16]_pad ,
		_w8955_,
		_w8956_,
		_w16277_
	);
	LUT3 #(
		.INIT('h2a)
	) name14377 (
		\m5_data_i[16]_pad ,
		_w8955_,
		_w8956_,
		_w16278_
	);
	LUT4 #(
		.INIT('hcdef)
	) name14378 (
		_w8950_,
		_w8953_,
		_w16277_,
		_w16278_,
		_w16279_
	);
	LUT4 #(
		.INIT('h7fff)
	) name14379 (
		_w16270_,
		_w16273_,
		_w16276_,
		_w16279_,
		_w16280_
	);
	LUT3 #(
		.INIT('h80)
	) name14380 (
		\m0_data_i[17]_pad ,
		_w8955_,
		_w8956_,
		_w16281_
	);
	LUT3 #(
		.INIT('h2a)
	) name14381 (
		\m7_data_i[17]_pad ,
		_w8955_,
		_w8956_,
		_w16282_
	);
	LUT4 #(
		.INIT('h6e7f)
	) name14382 (
		_w8950_,
		_w8953_,
		_w16281_,
		_w16282_,
		_w16283_
	);
	LUT3 #(
		.INIT('h80)
	) name14383 (
		\m6_data_i[17]_pad ,
		_w8955_,
		_w8956_,
		_w16284_
	);
	LUT3 #(
		.INIT('h80)
	) name14384 (
		\m2_data_i[17]_pad ,
		_w8955_,
		_w8956_,
		_w16285_
	);
	LUT4 #(
		.INIT('habef)
	) name14385 (
		_w8950_,
		_w8953_,
		_w16284_,
		_w16285_,
		_w16286_
	);
	LUT3 #(
		.INIT('h2a)
	) name14386 (
		\m5_data_i[17]_pad ,
		_w8955_,
		_w8956_,
		_w16287_
	);
	LUT3 #(
		.INIT('h2a)
	) name14387 (
		\m1_data_i[17]_pad ,
		_w8955_,
		_w8956_,
		_w16288_
	);
	LUT4 #(
		.INIT('h57df)
	) name14388 (
		_w8950_,
		_w8953_,
		_w16287_,
		_w16288_,
		_w16289_
	);
	LUT3 #(
		.INIT('h2a)
	) name14389 (
		\m3_data_i[17]_pad ,
		_w8955_,
		_w8956_,
		_w16290_
	);
	LUT3 #(
		.INIT('h80)
	) name14390 (
		\m4_data_i[17]_pad ,
		_w8955_,
		_w8956_,
		_w16291_
	);
	LUT4 #(
		.INIT('h9dbf)
	) name14391 (
		_w8950_,
		_w8953_,
		_w16290_,
		_w16291_,
		_w16292_
	);
	LUT4 #(
		.INIT('h7fff)
	) name14392 (
		_w16283_,
		_w16286_,
		_w16289_,
		_w16292_,
		_w16293_
	);
	LUT3 #(
		.INIT('h2a)
	) name14393 (
		\m1_data_i[18]_pad ,
		_w8955_,
		_w8956_,
		_w16294_
	);
	LUT3 #(
		.INIT('h80)
	) name14394 (
		\m2_data_i[18]_pad ,
		_w8955_,
		_w8956_,
		_w16295_
	);
	LUT4 #(
		.INIT('h3b7f)
	) name14395 (
		_w8950_,
		_w8953_,
		_w16294_,
		_w16295_,
		_w16296_
	);
	LUT3 #(
		.INIT('h2a)
	) name14396 (
		\m3_data_i[18]_pad ,
		_w8955_,
		_w8956_,
		_w16297_
	);
	LUT3 #(
		.INIT('h2a)
	) name14397 (
		\m7_data_i[18]_pad ,
		_w8955_,
		_w8956_,
		_w16298_
	);
	LUT4 #(
		.INIT('haebf)
	) name14398 (
		_w8950_,
		_w8953_,
		_w16297_,
		_w16298_,
		_w16299_
	);
	LUT3 #(
		.INIT('h80)
	) name14399 (
		\m4_data_i[18]_pad ,
		_w8955_,
		_w8956_,
		_w16300_
	);
	LUT3 #(
		.INIT('h80)
	) name14400 (
		\m0_data_i[18]_pad ,
		_w8955_,
		_w8956_,
		_w16301_
	);
	LUT4 #(
		.INIT('h57df)
	) name14401 (
		_w8950_,
		_w8953_,
		_w16300_,
		_w16301_,
		_w16302_
	);
	LUT3 #(
		.INIT('h80)
	) name14402 (
		\m6_data_i[18]_pad ,
		_w8955_,
		_w8956_,
		_w16303_
	);
	LUT3 #(
		.INIT('h2a)
	) name14403 (
		\m5_data_i[18]_pad ,
		_w8955_,
		_w8956_,
		_w16304_
	);
	LUT4 #(
		.INIT('hcdef)
	) name14404 (
		_w8950_,
		_w8953_,
		_w16303_,
		_w16304_,
		_w16305_
	);
	LUT4 #(
		.INIT('h7fff)
	) name14405 (
		_w16296_,
		_w16299_,
		_w16302_,
		_w16305_,
		_w16306_
	);
	LUT3 #(
		.INIT('h2a)
	) name14406 (
		\m1_data_i[19]_pad ,
		_w8955_,
		_w8956_,
		_w16307_
	);
	LUT3 #(
		.INIT('h80)
	) name14407 (
		\m2_data_i[19]_pad ,
		_w8955_,
		_w8956_,
		_w16308_
	);
	LUT4 #(
		.INIT('h3b7f)
	) name14408 (
		_w8950_,
		_w8953_,
		_w16307_,
		_w16308_,
		_w16309_
	);
	LUT3 #(
		.INIT('h80)
	) name14409 (
		\m0_data_i[19]_pad ,
		_w8955_,
		_w8956_,
		_w16310_
	);
	LUT3 #(
		.INIT('h2a)
	) name14410 (
		\m5_data_i[19]_pad ,
		_w8955_,
		_w8956_,
		_w16311_
	);
	LUT4 #(
		.INIT('h5d7f)
	) name14411 (
		_w8950_,
		_w8953_,
		_w16310_,
		_w16311_,
		_w16312_
	);
	LUT3 #(
		.INIT('h2a)
	) name14412 (
		\m7_data_i[19]_pad ,
		_w8955_,
		_w8956_,
		_w16313_
	);
	LUT3 #(
		.INIT('h80)
	) name14413 (
		\m6_data_i[19]_pad ,
		_w8955_,
		_w8956_,
		_w16314_
	);
	LUT3 #(
		.INIT('h57)
	) name14414 (
		_w8968_,
		_w16313_,
		_w16314_,
		_w16315_
	);
	LUT3 #(
		.INIT('h2a)
	) name14415 (
		\m3_data_i[19]_pad ,
		_w8955_,
		_w8956_,
		_w16316_
	);
	LUT3 #(
		.INIT('h80)
	) name14416 (
		\m4_data_i[19]_pad ,
		_w8955_,
		_w8956_,
		_w16317_
	);
	LUT4 #(
		.INIT('h9dbf)
	) name14417 (
		_w8950_,
		_w8953_,
		_w16316_,
		_w16317_,
		_w16318_
	);
	LUT4 #(
		.INIT('h7fff)
	) name14418 (
		_w16309_,
		_w16312_,
		_w16315_,
		_w16318_,
		_w16319_
	);
	LUT3 #(
		.INIT('h2a)
	) name14419 (
		\m3_data_i[1]_pad ,
		_w8955_,
		_w8956_,
		_w16320_
	);
	LUT3 #(
		.INIT('h80)
	) name14420 (
		\m4_data_i[1]_pad ,
		_w8955_,
		_w8956_,
		_w16321_
	);
	LUT4 #(
		.INIT('h9dbf)
	) name14421 (
		_w8950_,
		_w8953_,
		_w16320_,
		_w16321_,
		_w16322_
	);
	LUT3 #(
		.INIT('h80)
	) name14422 (
		\m0_data_i[1]_pad ,
		_w8955_,
		_w8956_,
		_w16323_
	);
	LUT3 #(
		.INIT('h80)
	) name14423 (
		\m2_data_i[1]_pad ,
		_w8955_,
		_w8956_,
		_w16324_
	);
	LUT4 #(
		.INIT('h3b7f)
	) name14424 (
		_w8950_,
		_w8953_,
		_w16323_,
		_w16324_,
		_w16325_
	);
	LUT3 #(
		.INIT('h2a)
	) name14425 (
		\m7_data_i[1]_pad ,
		_w8955_,
		_w8956_,
		_w16326_
	);
	LUT3 #(
		.INIT('h2a)
	) name14426 (
		\m1_data_i[1]_pad ,
		_w8955_,
		_w8956_,
		_w16327_
	);
	LUT4 #(
		.INIT('h67ef)
	) name14427 (
		_w8950_,
		_w8953_,
		_w16326_,
		_w16327_,
		_w16328_
	);
	LUT3 #(
		.INIT('h80)
	) name14428 (
		\m6_data_i[1]_pad ,
		_w8955_,
		_w8956_,
		_w16329_
	);
	LUT3 #(
		.INIT('h2a)
	) name14429 (
		\m5_data_i[1]_pad ,
		_w8955_,
		_w8956_,
		_w16330_
	);
	LUT4 #(
		.INIT('hcdef)
	) name14430 (
		_w8950_,
		_w8953_,
		_w16329_,
		_w16330_,
		_w16331_
	);
	LUT4 #(
		.INIT('h7fff)
	) name14431 (
		_w16322_,
		_w16325_,
		_w16328_,
		_w16331_,
		_w16332_
	);
	LUT3 #(
		.INIT('h2a)
	) name14432 (
		\m1_data_i[20]_pad ,
		_w8955_,
		_w8956_,
		_w16333_
	);
	LUT3 #(
		.INIT('h80)
	) name14433 (
		\m2_data_i[20]_pad ,
		_w8955_,
		_w8956_,
		_w16334_
	);
	LUT4 #(
		.INIT('h3b7f)
	) name14434 (
		_w8950_,
		_w8953_,
		_w16333_,
		_w16334_,
		_w16335_
	);
	LUT3 #(
		.INIT('h80)
	) name14435 (
		\m0_data_i[20]_pad ,
		_w8955_,
		_w8956_,
		_w16336_
	);
	LUT3 #(
		.INIT('h80)
	) name14436 (
		\m4_data_i[20]_pad ,
		_w8955_,
		_w8956_,
		_w16337_
	);
	LUT4 #(
		.INIT('h5d7f)
	) name14437 (
		_w8950_,
		_w8953_,
		_w16336_,
		_w16337_,
		_w16338_
	);
	LUT3 #(
		.INIT('h2a)
	) name14438 (
		\m7_data_i[20]_pad ,
		_w8955_,
		_w8956_,
		_w16339_
	);
	LUT3 #(
		.INIT('h2a)
	) name14439 (
		\m3_data_i[20]_pad ,
		_w8955_,
		_w8956_,
		_w16340_
	);
	LUT4 #(
		.INIT('habef)
	) name14440 (
		_w8950_,
		_w8953_,
		_w16339_,
		_w16340_,
		_w16341_
	);
	LUT3 #(
		.INIT('h80)
	) name14441 (
		\m6_data_i[20]_pad ,
		_w8955_,
		_w8956_,
		_w16342_
	);
	LUT3 #(
		.INIT('h2a)
	) name14442 (
		\m5_data_i[20]_pad ,
		_w8955_,
		_w8956_,
		_w16343_
	);
	LUT4 #(
		.INIT('hcdef)
	) name14443 (
		_w8950_,
		_w8953_,
		_w16342_,
		_w16343_,
		_w16344_
	);
	LUT4 #(
		.INIT('h7fff)
	) name14444 (
		_w16335_,
		_w16338_,
		_w16341_,
		_w16344_,
		_w16345_
	);
	LUT3 #(
		.INIT('h2a)
	) name14445 (
		\m1_data_i[21]_pad ,
		_w8955_,
		_w8956_,
		_w16346_
	);
	LUT3 #(
		.INIT('h80)
	) name14446 (
		\m2_data_i[21]_pad ,
		_w8955_,
		_w8956_,
		_w16347_
	);
	LUT4 #(
		.INIT('h3b7f)
	) name14447 (
		_w8950_,
		_w8953_,
		_w16346_,
		_w16347_,
		_w16348_
	);
	LUT3 #(
		.INIT('h80)
	) name14448 (
		\m0_data_i[21]_pad ,
		_w8955_,
		_w8956_,
		_w16349_
	);
	LUT3 #(
		.INIT('h80)
	) name14449 (
		\m4_data_i[21]_pad ,
		_w8955_,
		_w8956_,
		_w16350_
	);
	LUT4 #(
		.INIT('h5d7f)
	) name14450 (
		_w8950_,
		_w8953_,
		_w16349_,
		_w16350_,
		_w16351_
	);
	LUT3 #(
		.INIT('h2a)
	) name14451 (
		\m7_data_i[21]_pad ,
		_w8955_,
		_w8956_,
		_w16352_
	);
	LUT3 #(
		.INIT('h2a)
	) name14452 (
		\m3_data_i[21]_pad ,
		_w8955_,
		_w8956_,
		_w16353_
	);
	LUT4 #(
		.INIT('habef)
	) name14453 (
		_w8950_,
		_w8953_,
		_w16352_,
		_w16353_,
		_w16354_
	);
	LUT3 #(
		.INIT('h80)
	) name14454 (
		\m6_data_i[21]_pad ,
		_w8955_,
		_w8956_,
		_w16355_
	);
	LUT3 #(
		.INIT('h2a)
	) name14455 (
		\m5_data_i[21]_pad ,
		_w8955_,
		_w8956_,
		_w16356_
	);
	LUT4 #(
		.INIT('hcdef)
	) name14456 (
		_w8950_,
		_w8953_,
		_w16355_,
		_w16356_,
		_w16357_
	);
	LUT4 #(
		.INIT('h7fff)
	) name14457 (
		_w16348_,
		_w16351_,
		_w16354_,
		_w16357_,
		_w16358_
	);
	LUT3 #(
		.INIT('h2a)
	) name14458 (
		\m1_data_i[22]_pad ,
		_w8955_,
		_w8956_,
		_w16359_
	);
	LUT3 #(
		.INIT('h80)
	) name14459 (
		\m2_data_i[22]_pad ,
		_w8955_,
		_w8956_,
		_w16360_
	);
	LUT4 #(
		.INIT('h3b7f)
	) name14460 (
		_w8950_,
		_w8953_,
		_w16359_,
		_w16360_,
		_w16361_
	);
	LUT3 #(
		.INIT('h80)
	) name14461 (
		\m0_data_i[22]_pad ,
		_w8955_,
		_w8956_,
		_w16362_
	);
	LUT3 #(
		.INIT('h80)
	) name14462 (
		\m4_data_i[22]_pad ,
		_w8955_,
		_w8956_,
		_w16363_
	);
	LUT4 #(
		.INIT('h5d7f)
	) name14463 (
		_w8950_,
		_w8953_,
		_w16362_,
		_w16363_,
		_w16364_
	);
	LUT3 #(
		.INIT('h2a)
	) name14464 (
		\m7_data_i[22]_pad ,
		_w8955_,
		_w8956_,
		_w16365_
	);
	LUT3 #(
		.INIT('h2a)
	) name14465 (
		\m3_data_i[22]_pad ,
		_w8955_,
		_w8956_,
		_w16366_
	);
	LUT4 #(
		.INIT('habef)
	) name14466 (
		_w8950_,
		_w8953_,
		_w16365_,
		_w16366_,
		_w16367_
	);
	LUT3 #(
		.INIT('h80)
	) name14467 (
		\m6_data_i[22]_pad ,
		_w8955_,
		_w8956_,
		_w16368_
	);
	LUT3 #(
		.INIT('h2a)
	) name14468 (
		\m5_data_i[22]_pad ,
		_w8955_,
		_w8956_,
		_w16369_
	);
	LUT4 #(
		.INIT('hcdef)
	) name14469 (
		_w8950_,
		_w8953_,
		_w16368_,
		_w16369_,
		_w16370_
	);
	LUT4 #(
		.INIT('h7fff)
	) name14470 (
		_w16361_,
		_w16364_,
		_w16367_,
		_w16370_,
		_w16371_
	);
	LUT3 #(
		.INIT('h2a)
	) name14471 (
		\m1_data_i[23]_pad ,
		_w8955_,
		_w8956_,
		_w16372_
	);
	LUT3 #(
		.INIT('h80)
	) name14472 (
		\m2_data_i[23]_pad ,
		_w8955_,
		_w8956_,
		_w16373_
	);
	LUT4 #(
		.INIT('h3b7f)
	) name14473 (
		_w8950_,
		_w8953_,
		_w16372_,
		_w16373_,
		_w16374_
	);
	LUT3 #(
		.INIT('h80)
	) name14474 (
		\m0_data_i[23]_pad ,
		_w8955_,
		_w8956_,
		_w16375_
	);
	LUT3 #(
		.INIT('h80)
	) name14475 (
		\m4_data_i[23]_pad ,
		_w8955_,
		_w8956_,
		_w16376_
	);
	LUT4 #(
		.INIT('h5d7f)
	) name14476 (
		_w8950_,
		_w8953_,
		_w16375_,
		_w16376_,
		_w16377_
	);
	LUT3 #(
		.INIT('h2a)
	) name14477 (
		\m7_data_i[23]_pad ,
		_w8955_,
		_w8956_,
		_w16378_
	);
	LUT3 #(
		.INIT('h2a)
	) name14478 (
		\m3_data_i[23]_pad ,
		_w8955_,
		_w8956_,
		_w16379_
	);
	LUT4 #(
		.INIT('habef)
	) name14479 (
		_w8950_,
		_w8953_,
		_w16378_,
		_w16379_,
		_w16380_
	);
	LUT3 #(
		.INIT('h80)
	) name14480 (
		\m6_data_i[23]_pad ,
		_w8955_,
		_w8956_,
		_w16381_
	);
	LUT3 #(
		.INIT('h2a)
	) name14481 (
		\m5_data_i[23]_pad ,
		_w8955_,
		_w8956_,
		_w16382_
	);
	LUT4 #(
		.INIT('hcdef)
	) name14482 (
		_w8950_,
		_w8953_,
		_w16381_,
		_w16382_,
		_w16383_
	);
	LUT4 #(
		.INIT('h7fff)
	) name14483 (
		_w16374_,
		_w16377_,
		_w16380_,
		_w16383_,
		_w16384_
	);
	LUT3 #(
		.INIT('h80)
	) name14484 (
		\m6_data_i[24]_pad ,
		_w8955_,
		_w8956_,
		_w16385_
	);
	LUT3 #(
		.INIT('h2a)
	) name14485 (
		\m5_data_i[24]_pad ,
		_w8955_,
		_w8956_,
		_w16386_
	);
	LUT4 #(
		.INIT('hcdef)
	) name14486 (
		_w8950_,
		_w8953_,
		_w16385_,
		_w16386_,
		_w16387_
	);
	LUT3 #(
		.INIT('h2a)
	) name14487 (
		\m1_data_i[24]_pad ,
		_w8955_,
		_w8956_,
		_w16388_
	);
	LUT3 #(
		.INIT('h80)
	) name14488 (
		\m4_data_i[24]_pad ,
		_w8955_,
		_w8956_,
		_w16389_
	);
	LUT4 #(
		.INIT('h5d7f)
	) name14489 (
		_w8950_,
		_w8953_,
		_w16388_,
		_w16389_,
		_w16390_
	);
	LUT3 #(
		.INIT('h80)
	) name14490 (
		\m2_data_i[24]_pad ,
		_w8955_,
		_w8956_,
		_w16391_
	);
	LUT3 #(
		.INIT('h2a)
	) name14491 (
		\m3_data_i[24]_pad ,
		_w8955_,
		_w8956_,
		_w16392_
	);
	LUT3 #(
		.INIT('h57)
	) name14492 (
		_w8974_,
		_w16391_,
		_w16392_,
		_w16393_
	);
	LUT3 #(
		.INIT('h80)
	) name14493 (
		\m0_data_i[24]_pad ,
		_w8955_,
		_w8956_,
		_w16394_
	);
	LUT3 #(
		.INIT('h2a)
	) name14494 (
		\m7_data_i[24]_pad ,
		_w8955_,
		_w8956_,
		_w16395_
	);
	LUT4 #(
		.INIT('h6e7f)
	) name14495 (
		_w8950_,
		_w8953_,
		_w16394_,
		_w16395_,
		_w16396_
	);
	LUT4 #(
		.INIT('h7fff)
	) name14496 (
		_w16387_,
		_w16390_,
		_w16393_,
		_w16396_,
		_w16397_
	);
	LUT3 #(
		.INIT('h2a)
	) name14497 (
		\m1_data_i[25]_pad ,
		_w8955_,
		_w8956_,
		_w16398_
	);
	LUT3 #(
		.INIT('h80)
	) name14498 (
		\m2_data_i[25]_pad ,
		_w8955_,
		_w8956_,
		_w16399_
	);
	LUT4 #(
		.INIT('h3b7f)
	) name14499 (
		_w8950_,
		_w8953_,
		_w16398_,
		_w16399_,
		_w16400_
	);
	LUT3 #(
		.INIT('h80)
	) name14500 (
		\m0_data_i[25]_pad ,
		_w8955_,
		_w8956_,
		_w16401_
	);
	LUT3 #(
		.INIT('h80)
	) name14501 (
		\m4_data_i[25]_pad ,
		_w8955_,
		_w8956_,
		_w16402_
	);
	LUT4 #(
		.INIT('h5d7f)
	) name14502 (
		_w8950_,
		_w8953_,
		_w16401_,
		_w16402_,
		_w16403_
	);
	LUT3 #(
		.INIT('h2a)
	) name14503 (
		\m7_data_i[25]_pad ,
		_w8955_,
		_w8956_,
		_w16404_
	);
	LUT3 #(
		.INIT('h2a)
	) name14504 (
		\m3_data_i[25]_pad ,
		_w8955_,
		_w8956_,
		_w16405_
	);
	LUT4 #(
		.INIT('habef)
	) name14505 (
		_w8950_,
		_w8953_,
		_w16404_,
		_w16405_,
		_w16406_
	);
	LUT3 #(
		.INIT('h80)
	) name14506 (
		\m6_data_i[25]_pad ,
		_w8955_,
		_w8956_,
		_w16407_
	);
	LUT3 #(
		.INIT('h2a)
	) name14507 (
		\m5_data_i[25]_pad ,
		_w8955_,
		_w8956_,
		_w16408_
	);
	LUT4 #(
		.INIT('hcdef)
	) name14508 (
		_w8950_,
		_w8953_,
		_w16407_,
		_w16408_,
		_w16409_
	);
	LUT4 #(
		.INIT('h7fff)
	) name14509 (
		_w16400_,
		_w16403_,
		_w16406_,
		_w16409_,
		_w16410_
	);
	LUT3 #(
		.INIT('h80)
	) name14510 (
		\m0_data_i[26]_pad ,
		_w8955_,
		_w8956_,
		_w16411_
	);
	LUT3 #(
		.INIT('h2a)
	) name14511 (
		\m7_data_i[26]_pad ,
		_w8955_,
		_w8956_,
		_w16412_
	);
	LUT4 #(
		.INIT('h6e7f)
	) name14512 (
		_w8950_,
		_w8953_,
		_w16411_,
		_w16412_,
		_w16413_
	);
	LUT3 #(
		.INIT('h2a)
	) name14513 (
		\m1_data_i[26]_pad ,
		_w8955_,
		_w8956_,
		_w16414_
	);
	LUT3 #(
		.INIT('h80)
	) name14514 (
		\m4_data_i[26]_pad ,
		_w8955_,
		_w8956_,
		_w16415_
	);
	LUT4 #(
		.INIT('h5d7f)
	) name14515 (
		_w8950_,
		_w8953_,
		_w16414_,
		_w16415_,
		_w16416_
	);
	LUT3 #(
		.INIT('h80)
	) name14516 (
		\m2_data_i[26]_pad ,
		_w8955_,
		_w8956_,
		_w16417_
	);
	LUT3 #(
		.INIT('h2a)
	) name14517 (
		\m3_data_i[26]_pad ,
		_w8955_,
		_w8956_,
		_w16418_
	);
	LUT3 #(
		.INIT('h57)
	) name14518 (
		_w8974_,
		_w16417_,
		_w16418_,
		_w16419_
	);
	LUT3 #(
		.INIT('h80)
	) name14519 (
		\m6_data_i[26]_pad ,
		_w8955_,
		_w8956_,
		_w16420_
	);
	LUT3 #(
		.INIT('h2a)
	) name14520 (
		\m5_data_i[26]_pad ,
		_w8955_,
		_w8956_,
		_w16421_
	);
	LUT4 #(
		.INIT('hcdef)
	) name14521 (
		_w8950_,
		_w8953_,
		_w16420_,
		_w16421_,
		_w16422_
	);
	LUT4 #(
		.INIT('h7fff)
	) name14522 (
		_w16413_,
		_w16416_,
		_w16419_,
		_w16422_,
		_w16423_
	);
	LUT3 #(
		.INIT('h80)
	) name14523 (
		\m0_data_i[27]_pad ,
		_w8955_,
		_w8956_,
		_w16424_
	);
	LUT3 #(
		.INIT('h2a)
	) name14524 (
		\m7_data_i[27]_pad ,
		_w8955_,
		_w8956_,
		_w16425_
	);
	LUT4 #(
		.INIT('h6e7f)
	) name14525 (
		_w8950_,
		_w8953_,
		_w16424_,
		_w16425_,
		_w16426_
	);
	LUT3 #(
		.INIT('h2a)
	) name14526 (
		\m1_data_i[27]_pad ,
		_w8955_,
		_w8956_,
		_w16427_
	);
	LUT3 #(
		.INIT('h80)
	) name14527 (
		\m4_data_i[27]_pad ,
		_w8955_,
		_w8956_,
		_w16428_
	);
	LUT4 #(
		.INIT('h5d7f)
	) name14528 (
		_w8950_,
		_w8953_,
		_w16427_,
		_w16428_,
		_w16429_
	);
	LUT3 #(
		.INIT('h80)
	) name14529 (
		\m2_data_i[27]_pad ,
		_w8955_,
		_w8956_,
		_w16430_
	);
	LUT3 #(
		.INIT('h2a)
	) name14530 (
		\m3_data_i[27]_pad ,
		_w8955_,
		_w8956_,
		_w16431_
	);
	LUT3 #(
		.INIT('h57)
	) name14531 (
		_w8974_,
		_w16430_,
		_w16431_,
		_w16432_
	);
	LUT3 #(
		.INIT('h80)
	) name14532 (
		\m6_data_i[27]_pad ,
		_w8955_,
		_w8956_,
		_w16433_
	);
	LUT3 #(
		.INIT('h2a)
	) name14533 (
		\m5_data_i[27]_pad ,
		_w8955_,
		_w8956_,
		_w16434_
	);
	LUT4 #(
		.INIT('hcdef)
	) name14534 (
		_w8950_,
		_w8953_,
		_w16433_,
		_w16434_,
		_w16435_
	);
	LUT4 #(
		.INIT('h7fff)
	) name14535 (
		_w16426_,
		_w16429_,
		_w16432_,
		_w16435_,
		_w16436_
	);
	LUT3 #(
		.INIT('h2a)
	) name14536 (
		\m1_data_i[28]_pad ,
		_w8955_,
		_w8956_,
		_w16437_
	);
	LUT3 #(
		.INIT('h80)
	) name14537 (
		\m2_data_i[28]_pad ,
		_w8955_,
		_w8956_,
		_w16438_
	);
	LUT4 #(
		.INIT('h3b7f)
	) name14538 (
		_w8950_,
		_w8953_,
		_w16437_,
		_w16438_,
		_w16439_
	);
	LUT3 #(
		.INIT('h80)
	) name14539 (
		\m0_data_i[28]_pad ,
		_w8955_,
		_w8956_,
		_w16440_
	);
	LUT3 #(
		.INIT('h80)
	) name14540 (
		\m4_data_i[28]_pad ,
		_w8955_,
		_w8956_,
		_w16441_
	);
	LUT4 #(
		.INIT('h5d7f)
	) name14541 (
		_w8950_,
		_w8953_,
		_w16440_,
		_w16441_,
		_w16442_
	);
	LUT3 #(
		.INIT('h2a)
	) name14542 (
		\m7_data_i[28]_pad ,
		_w8955_,
		_w8956_,
		_w16443_
	);
	LUT3 #(
		.INIT('h2a)
	) name14543 (
		\m3_data_i[28]_pad ,
		_w8955_,
		_w8956_,
		_w16444_
	);
	LUT4 #(
		.INIT('habef)
	) name14544 (
		_w8950_,
		_w8953_,
		_w16443_,
		_w16444_,
		_w16445_
	);
	LUT3 #(
		.INIT('h80)
	) name14545 (
		\m6_data_i[28]_pad ,
		_w8955_,
		_w8956_,
		_w16446_
	);
	LUT3 #(
		.INIT('h2a)
	) name14546 (
		\m5_data_i[28]_pad ,
		_w8955_,
		_w8956_,
		_w16447_
	);
	LUT4 #(
		.INIT('hcdef)
	) name14547 (
		_w8950_,
		_w8953_,
		_w16446_,
		_w16447_,
		_w16448_
	);
	LUT4 #(
		.INIT('h7fff)
	) name14548 (
		_w16439_,
		_w16442_,
		_w16445_,
		_w16448_,
		_w16449_
	);
	LUT3 #(
		.INIT('h2a)
	) name14549 (
		\m1_data_i[29]_pad ,
		_w8955_,
		_w8956_,
		_w16450_
	);
	LUT3 #(
		.INIT('h80)
	) name14550 (
		\m2_data_i[29]_pad ,
		_w8955_,
		_w8956_,
		_w16451_
	);
	LUT4 #(
		.INIT('h3b7f)
	) name14551 (
		_w8950_,
		_w8953_,
		_w16450_,
		_w16451_,
		_w16452_
	);
	LUT3 #(
		.INIT('h80)
	) name14552 (
		\m0_data_i[29]_pad ,
		_w8955_,
		_w8956_,
		_w16453_
	);
	LUT3 #(
		.INIT('h80)
	) name14553 (
		\m4_data_i[29]_pad ,
		_w8955_,
		_w8956_,
		_w16454_
	);
	LUT4 #(
		.INIT('h5d7f)
	) name14554 (
		_w8950_,
		_w8953_,
		_w16453_,
		_w16454_,
		_w16455_
	);
	LUT3 #(
		.INIT('h2a)
	) name14555 (
		\m7_data_i[29]_pad ,
		_w8955_,
		_w8956_,
		_w16456_
	);
	LUT3 #(
		.INIT('h2a)
	) name14556 (
		\m3_data_i[29]_pad ,
		_w8955_,
		_w8956_,
		_w16457_
	);
	LUT4 #(
		.INIT('habef)
	) name14557 (
		_w8950_,
		_w8953_,
		_w16456_,
		_w16457_,
		_w16458_
	);
	LUT3 #(
		.INIT('h80)
	) name14558 (
		\m6_data_i[29]_pad ,
		_w8955_,
		_w8956_,
		_w16459_
	);
	LUT3 #(
		.INIT('h2a)
	) name14559 (
		\m5_data_i[29]_pad ,
		_w8955_,
		_w8956_,
		_w16460_
	);
	LUT4 #(
		.INIT('hcdef)
	) name14560 (
		_w8950_,
		_w8953_,
		_w16459_,
		_w16460_,
		_w16461_
	);
	LUT4 #(
		.INIT('h7fff)
	) name14561 (
		_w16452_,
		_w16455_,
		_w16458_,
		_w16461_,
		_w16462_
	);
	LUT3 #(
		.INIT('h2a)
	) name14562 (
		\m1_data_i[2]_pad ,
		_w8955_,
		_w8956_,
		_w16463_
	);
	LUT3 #(
		.INIT('h80)
	) name14563 (
		\m2_data_i[2]_pad ,
		_w8955_,
		_w8956_,
		_w16464_
	);
	LUT4 #(
		.INIT('h3b7f)
	) name14564 (
		_w8950_,
		_w8953_,
		_w16463_,
		_w16464_,
		_w16465_
	);
	LUT3 #(
		.INIT('h80)
	) name14565 (
		\m0_data_i[2]_pad ,
		_w8955_,
		_w8956_,
		_w16466_
	);
	LUT3 #(
		.INIT('h2a)
	) name14566 (
		\m5_data_i[2]_pad ,
		_w8955_,
		_w8956_,
		_w16467_
	);
	LUT4 #(
		.INIT('h5d7f)
	) name14567 (
		_w8950_,
		_w8953_,
		_w16466_,
		_w16467_,
		_w16468_
	);
	LUT3 #(
		.INIT('h2a)
	) name14568 (
		\m7_data_i[2]_pad ,
		_w8955_,
		_w8956_,
		_w16469_
	);
	LUT3 #(
		.INIT('h80)
	) name14569 (
		\m6_data_i[2]_pad ,
		_w8955_,
		_w8956_,
		_w16470_
	);
	LUT3 #(
		.INIT('h57)
	) name14570 (
		_w8968_,
		_w16469_,
		_w16470_,
		_w16471_
	);
	LUT3 #(
		.INIT('h2a)
	) name14571 (
		\m3_data_i[2]_pad ,
		_w8955_,
		_w8956_,
		_w16472_
	);
	LUT3 #(
		.INIT('h80)
	) name14572 (
		\m4_data_i[2]_pad ,
		_w8955_,
		_w8956_,
		_w16473_
	);
	LUT4 #(
		.INIT('h9dbf)
	) name14573 (
		_w8950_,
		_w8953_,
		_w16472_,
		_w16473_,
		_w16474_
	);
	LUT4 #(
		.INIT('h7fff)
	) name14574 (
		_w16465_,
		_w16468_,
		_w16471_,
		_w16474_,
		_w16475_
	);
	LUT3 #(
		.INIT('h2a)
	) name14575 (
		\m1_data_i[30]_pad ,
		_w8955_,
		_w8956_,
		_w16476_
	);
	LUT3 #(
		.INIT('h80)
	) name14576 (
		\m2_data_i[30]_pad ,
		_w8955_,
		_w8956_,
		_w16477_
	);
	LUT4 #(
		.INIT('h3b7f)
	) name14577 (
		_w8950_,
		_w8953_,
		_w16476_,
		_w16477_,
		_w16478_
	);
	LUT3 #(
		.INIT('h80)
	) name14578 (
		\m0_data_i[30]_pad ,
		_w8955_,
		_w8956_,
		_w16479_
	);
	LUT3 #(
		.INIT('h80)
	) name14579 (
		\m4_data_i[30]_pad ,
		_w8955_,
		_w8956_,
		_w16480_
	);
	LUT4 #(
		.INIT('h5d7f)
	) name14580 (
		_w8950_,
		_w8953_,
		_w16479_,
		_w16480_,
		_w16481_
	);
	LUT3 #(
		.INIT('h2a)
	) name14581 (
		\m7_data_i[30]_pad ,
		_w8955_,
		_w8956_,
		_w16482_
	);
	LUT3 #(
		.INIT('h2a)
	) name14582 (
		\m3_data_i[30]_pad ,
		_w8955_,
		_w8956_,
		_w16483_
	);
	LUT4 #(
		.INIT('habef)
	) name14583 (
		_w8950_,
		_w8953_,
		_w16482_,
		_w16483_,
		_w16484_
	);
	LUT3 #(
		.INIT('h80)
	) name14584 (
		\m6_data_i[30]_pad ,
		_w8955_,
		_w8956_,
		_w16485_
	);
	LUT3 #(
		.INIT('h2a)
	) name14585 (
		\m5_data_i[30]_pad ,
		_w8955_,
		_w8956_,
		_w16486_
	);
	LUT4 #(
		.INIT('hcdef)
	) name14586 (
		_w8950_,
		_w8953_,
		_w16485_,
		_w16486_,
		_w16487_
	);
	LUT4 #(
		.INIT('h7fff)
	) name14587 (
		_w16478_,
		_w16481_,
		_w16484_,
		_w16487_,
		_w16488_
	);
	LUT3 #(
		.INIT('h2a)
	) name14588 (
		\m1_data_i[31]_pad ,
		_w8955_,
		_w8956_,
		_w16489_
	);
	LUT3 #(
		.INIT('h80)
	) name14589 (
		\m2_data_i[31]_pad ,
		_w8955_,
		_w8956_,
		_w16490_
	);
	LUT4 #(
		.INIT('h3b7f)
	) name14590 (
		_w8950_,
		_w8953_,
		_w16489_,
		_w16490_,
		_w16491_
	);
	LUT3 #(
		.INIT('h80)
	) name14591 (
		\m0_data_i[31]_pad ,
		_w8955_,
		_w8956_,
		_w16492_
	);
	LUT3 #(
		.INIT('h2a)
	) name14592 (
		\m5_data_i[31]_pad ,
		_w8955_,
		_w8956_,
		_w16493_
	);
	LUT4 #(
		.INIT('h5d7f)
	) name14593 (
		_w8950_,
		_w8953_,
		_w16492_,
		_w16493_,
		_w16494_
	);
	LUT3 #(
		.INIT('h2a)
	) name14594 (
		\m7_data_i[31]_pad ,
		_w8955_,
		_w8956_,
		_w16495_
	);
	LUT3 #(
		.INIT('h80)
	) name14595 (
		\m6_data_i[31]_pad ,
		_w8955_,
		_w8956_,
		_w16496_
	);
	LUT3 #(
		.INIT('h57)
	) name14596 (
		_w8968_,
		_w16495_,
		_w16496_,
		_w16497_
	);
	LUT3 #(
		.INIT('h2a)
	) name14597 (
		\m3_data_i[31]_pad ,
		_w8955_,
		_w8956_,
		_w16498_
	);
	LUT3 #(
		.INIT('h80)
	) name14598 (
		\m4_data_i[31]_pad ,
		_w8955_,
		_w8956_,
		_w16499_
	);
	LUT4 #(
		.INIT('h9dbf)
	) name14599 (
		_w8950_,
		_w8953_,
		_w16498_,
		_w16499_,
		_w16500_
	);
	LUT4 #(
		.INIT('h7fff)
	) name14600 (
		_w16491_,
		_w16494_,
		_w16497_,
		_w16500_,
		_w16501_
	);
	LUT3 #(
		.INIT('h80)
	) name14601 (
		\m0_data_i[3]_pad ,
		_w8955_,
		_w8956_,
		_w16502_
	);
	LUT3 #(
		.INIT('h2a)
	) name14602 (
		\m7_data_i[3]_pad ,
		_w8955_,
		_w8956_,
		_w16503_
	);
	LUT4 #(
		.INIT('h6e7f)
	) name14603 (
		_w8950_,
		_w8953_,
		_w16502_,
		_w16503_,
		_w16504_
	);
	LUT3 #(
		.INIT('h2a)
	) name14604 (
		\m1_data_i[3]_pad ,
		_w8955_,
		_w8956_,
		_w16505_
	);
	LUT3 #(
		.INIT('h2a)
	) name14605 (
		\m5_data_i[3]_pad ,
		_w8955_,
		_w8956_,
		_w16506_
	);
	LUT4 #(
		.INIT('h5d7f)
	) name14606 (
		_w8950_,
		_w8953_,
		_w16505_,
		_w16506_,
		_w16507_
	);
	LUT3 #(
		.INIT('h80)
	) name14607 (
		\m2_data_i[3]_pad ,
		_w8955_,
		_w8956_,
		_w16508_
	);
	LUT3 #(
		.INIT('h80)
	) name14608 (
		\m6_data_i[3]_pad ,
		_w8955_,
		_w8956_,
		_w16509_
	);
	LUT4 #(
		.INIT('haebf)
	) name14609 (
		_w8950_,
		_w8953_,
		_w16508_,
		_w16509_,
		_w16510_
	);
	LUT3 #(
		.INIT('h2a)
	) name14610 (
		\m3_data_i[3]_pad ,
		_w8955_,
		_w8956_,
		_w16511_
	);
	LUT3 #(
		.INIT('h80)
	) name14611 (
		\m4_data_i[3]_pad ,
		_w8955_,
		_w8956_,
		_w16512_
	);
	LUT4 #(
		.INIT('h9dbf)
	) name14612 (
		_w8950_,
		_w8953_,
		_w16511_,
		_w16512_,
		_w16513_
	);
	LUT4 #(
		.INIT('h7fff)
	) name14613 (
		_w16504_,
		_w16507_,
		_w16510_,
		_w16513_,
		_w16514_
	);
	LUT3 #(
		.INIT('h2a)
	) name14614 (
		\m1_data_i[4]_pad ,
		_w8955_,
		_w8956_,
		_w16515_
	);
	LUT3 #(
		.INIT('h80)
	) name14615 (
		\m2_data_i[4]_pad ,
		_w8955_,
		_w8956_,
		_w16516_
	);
	LUT4 #(
		.INIT('h3b7f)
	) name14616 (
		_w8950_,
		_w8953_,
		_w16515_,
		_w16516_,
		_w16517_
	);
	LUT3 #(
		.INIT('h80)
	) name14617 (
		\m0_data_i[4]_pad ,
		_w8955_,
		_w8956_,
		_w16518_
	);
	LUT3 #(
		.INIT('h80)
	) name14618 (
		\m4_data_i[4]_pad ,
		_w8955_,
		_w8956_,
		_w16519_
	);
	LUT4 #(
		.INIT('h5d7f)
	) name14619 (
		_w8950_,
		_w8953_,
		_w16518_,
		_w16519_,
		_w16520_
	);
	LUT3 #(
		.INIT('h2a)
	) name14620 (
		\m7_data_i[4]_pad ,
		_w8955_,
		_w8956_,
		_w16521_
	);
	LUT3 #(
		.INIT('h2a)
	) name14621 (
		\m3_data_i[4]_pad ,
		_w8955_,
		_w8956_,
		_w16522_
	);
	LUT4 #(
		.INIT('habef)
	) name14622 (
		_w8950_,
		_w8953_,
		_w16521_,
		_w16522_,
		_w16523_
	);
	LUT3 #(
		.INIT('h80)
	) name14623 (
		\m6_data_i[4]_pad ,
		_w8955_,
		_w8956_,
		_w16524_
	);
	LUT3 #(
		.INIT('h2a)
	) name14624 (
		\m5_data_i[4]_pad ,
		_w8955_,
		_w8956_,
		_w16525_
	);
	LUT4 #(
		.INIT('hcdef)
	) name14625 (
		_w8950_,
		_w8953_,
		_w16524_,
		_w16525_,
		_w16526_
	);
	LUT4 #(
		.INIT('h7fff)
	) name14626 (
		_w16517_,
		_w16520_,
		_w16523_,
		_w16526_,
		_w16527_
	);
	LUT3 #(
		.INIT('h2a)
	) name14627 (
		\m1_data_i[5]_pad ,
		_w8955_,
		_w8956_,
		_w16528_
	);
	LUT3 #(
		.INIT('h80)
	) name14628 (
		\m2_data_i[5]_pad ,
		_w8955_,
		_w8956_,
		_w16529_
	);
	LUT4 #(
		.INIT('h3b7f)
	) name14629 (
		_w8950_,
		_w8953_,
		_w16528_,
		_w16529_,
		_w16530_
	);
	LUT3 #(
		.INIT('h80)
	) name14630 (
		\m0_data_i[5]_pad ,
		_w8955_,
		_w8956_,
		_w16531_
	);
	LUT3 #(
		.INIT('h2a)
	) name14631 (
		\m5_data_i[5]_pad ,
		_w8955_,
		_w8956_,
		_w16532_
	);
	LUT4 #(
		.INIT('h5d7f)
	) name14632 (
		_w8950_,
		_w8953_,
		_w16531_,
		_w16532_,
		_w16533_
	);
	LUT3 #(
		.INIT('h2a)
	) name14633 (
		\m7_data_i[5]_pad ,
		_w8955_,
		_w8956_,
		_w16534_
	);
	LUT3 #(
		.INIT('h80)
	) name14634 (
		\m6_data_i[5]_pad ,
		_w8955_,
		_w8956_,
		_w16535_
	);
	LUT3 #(
		.INIT('h57)
	) name14635 (
		_w8968_,
		_w16534_,
		_w16535_,
		_w16536_
	);
	LUT3 #(
		.INIT('h2a)
	) name14636 (
		\m3_data_i[5]_pad ,
		_w8955_,
		_w8956_,
		_w16537_
	);
	LUT3 #(
		.INIT('h80)
	) name14637 (
		\m4_data_i[5]_pad ,
		_w8955_,
		_w8956_,
		_w16538_
	);
	LUT4 #(
		.INIT('h9dbf)
	) name14638 (
		_w8950_,
		_w8953_,
		_w16537_,
		_w16538_,
		_w16539_
	);
	LUT4 #(
		.INIT('h7fff)
	) name14639 (
		_w16530_,
		_w16533_,
		_w16536_,
		_w16539_,
		_w16540_
	);
	LUT3 #(
		.INIT('h2a)
	) name14640 (
		\m3_data_i[6]_pad ,
		_w8955_,
		_w8956_,
		_w16541_
	);
	LUT3 #(
		.INIT('h80)
	) name14641 (
		\m4_data_i[6]_pad ,
		_w8955_,
		_w8956_,
		_w16542_
	);
	LUT4 #(
		.INIT('h9dbf)
	) name14642 (
		_w8950_,
		_w8953_,
		_w16541_,
		_w16542_,
		_w16543_
	);
	LUT3 #(
		.INIT('h2a)
	) name14643 (
		\m1_data_i[6]_pad ,
		_w8955_,
		_w8956_,
		_w16544_
	);
	LUT3 #(
		.INIT('h2a)
	) name14644 (
		\m5_data_i[6]_pad ,
		_w8955_,
		_w8956_,
		_w16545_
	);
	LUT4 #(
		.INIT('h5d7f)
	) name14645 (
		_w8950_,
		_w8953_,
		_w16544_,
		_w16545_,
		_w16546_
	);
	LUT3 #(
		.INIT('h80)
	) name14646 (
		\m2_data_i[6]_pad ,
		_w8955_,
		_w8956_,
		_w16547_
	);
	LUT3 #(
		.INIT('h80)
	) name14647 (
		\m6_data_i[6]_pad ,
		_w8955_,
		_w8956_,
		_w16548_
	);
	LUT4 #(
		.INIT('haebf)
	) name14648 (
		_w8950_,
		_w8953_,
		_w16547_,
		_w16548_,
		_w16549_
	);
	LUT3 #(
		.INIT('h80)
	) name14649 (
		\m0_data_i[6]_pad ,
		_w8955_,
		_w8956_,
		_w16550_
	);
	LUT3 #(
		.INIT('h2a)
	) name14650 (
		\m7_data_i[6]_pad ,
		_w8955_,
		_w8956_,
		_w16551_
	);
	LUT4 #(
		.INIT('h6e7f)
	) name14651 (
		_w8950_,
		_w8953_,
		_w16550_,
		_w16551_,
		_w16552_
	);
	LUT4 #(
		.INIT('h7fff)
	) name14652 (
		_w16543_,
		_w16546_,
		_w16549_,
		_w16552_,
		_w16553_
	);
	LUT3 #(
		.INIT('h2a)
	) name14653 (
		\m3_data_i[7]_pad ,
		_w8955_,
		_w8956_,
		_w16554_
	);
	LUT3 #(
		.INIT('h80)
	) name14654 (
		\m4_data_i[7]_pad ,
		_w8955_,
		_w8956_,
		_w16555_
	);
	LUT4 #(
		.INIT('h9dbf)
	) name14655 (
		_w8950_,
		_w8953_,
		_w16554_,
		_w16555_,
		_w16556_
	);
	LUT3 #(
		.INIT('h80)
	) name14656 (
		\m0_data_i[7]_pad ,
		_w8955_,
		_w8956_,
		_w16557_
	);
	LUT3 #(
		.INIT('h80)
	) name14657 (
		\m2_data_i[7]_pad ,
		_w8955_,
		_w8956_,
		_w16558_
	);
	LUT4 #(
		.INIT('h3b7f)
	) name14658 (
		_w8950_,
		_w8953_,
		_w16557_,
		_w16558_,
		_w16559_
	);
	LUT3 #(
		.INIT('h2a)
	) name14659 (
		\m7_data_i[7]_pad ,
		_w8955_,
		_w8956_,
		_w16560_
	);
	LUT3 #(
		.INIT('h2a)
	) name14660 (
		\m1_data_i[7]_pad ,
		_w8955_,
		_w8956_,
		_w16561_
	);
	LUT4 #(
		.INIT('h67ef)
	) name14661 (
		_w8950_,
		_w8953_,
		_w16560_,
		_w16561_,
		_w16562_
	);
	LUT3 #(
		.INIT('h80)
	) name14662 (
		\m6_data_i[7]_pad ,
		_w8955_,
		_w8956_,
		_w16563_
	);
	LUT3 #(
		.INIT('h2a)
	) name14663 (
		\m5_data_i[7]_pad ,
		_w8955_,
		_w8956_,
		_w16564_
	);
	LUT4 #(
		.INIT('hcdef)
	) name14664 (
		_w8950_,
		_w8953_,
		_w16563_,
		_w16564_,
		_w16565_
	);
	LUT4 #(
		.INIT('h7fff)
	) name14665 (
		_w16556_,
		_w16559_,
		_w16562_,
		_w16565_,
		_w16566_
	);
	LUT3 #(
		.INIT('h2a)
	) name14666 (
		\m3_data_i[8]_pad ,
		_w8955_,
		_w8956_,
		_w16567_
	);
	LUT3 #(
		.INIT('h80)
	) name14667 (
		\m4_data_i[8]_pad ,
		_w8955_,
		_w8956_,
		_w16568_
	);
	LUT4 #(
		.INIT('h9dbf)
	) name14668 (
		_w8950_,
		_w8953_,
		_w16567_,
		_w16568_,
		_w16569_
	);
	LUT3 #(
		.INIT('h2a)
	) name14669 (
		\m1_data_i[8]_pad ,
		_w8955_,
		_w8956_,
		_w16570_
	);
	LUT3 #(
		.INIT('h2a)
	) name14670 (
		\m7_data_i[8]_pad ,
		_w8955_,
		_w8956_,
		_w16571_
	);
	LUT4 #(
		.INIT('h6e7f)
	) name14671 (
		_w8950_,
		_w8953_,
		_w16570_,
		_w16571_,
		_w16572_
	);
	LUT3 #(
		.INIT('h80)
	) name14672 (
		\m2_data_i[8]_pad ,
		_w8955_,
		_w8956_,
		_w16573_
	);
	LUT3 #(
		.INIT('h80)
	) name14673 (
		\m0_data_i[8]_pad ,
		_w8955_,
		_w8956_,
		_w16574_
	);
	LUT4 #(
		.INIT('h37bf)
	) name14674 (
		_w8950_,
		_w8953_,
		_w16573_,
		_w16574_,
		_w16575_
	);
	LUT3 #(
		.INIT('h80)
	) name14675 (
		\m6_data_i[8]_pad ,
		_w8955_,
		_w8956_,
		_w16576_
	);
	LUT3 #(
		.INIT('h2a)
	) name14676 (
		\m5_data_i[8]_pad ,
		_w8955_,
		_w8956_,
		_w16577_
	);
	LUT4 #(
		.INIT('hcdef)
	) name14677 (
		_w8950_,
		_w8953_,
		_w16576_,
		_w16577_,
		_w16578_
	);
	LUT4 #(
		.INIT('h7fff)
	) name14678 (
		_w16569_,
		_w16572_,
		_w16575_,
		_w16578_,
		_w16579_
	);
	LUT3 #(
		.INIT('h2a)
	) name14679 (
		\m1_data_i[9]_pad ,
		_w8955_,
		_w8956_,
		_w16580_
	);
	LUT3 #(
		.INIT('h80)
	) name14680 (
		\m2_data_i[9]_pad ,
		_w8955_,
		_w8956_,
		_w16581_
	);
	LUT4 #(
		.INIT('h3b7f)
	) name14681 (
		_w8950_,
		_w8953_,
		_w16580_,
		_w16581_,
		_w16582_
	);
	LUT3 #(
		.INIT('h80)
	) name14682 (
		\m0_data_i[9]_pad ,
		_w8955_,
		_w8956_,
		_w16583_
	);
	LUT3 #(
		.INIT('h2a)
	) name14683 (
		\m5_data_i[9]_pad ,
		_w8955_,
		_w8956_,
		_w16584_
	);
	LUT4 #(
		.INIT('h5d7f)
	) name14684 (
		_w8950_,
		_w8953_,
		_w16583_,
		_w16584_,
		_w16585_
	);
	LUT3 #(
		.INIT('h2a)
	) name14685 (
		\m7_data_i[9]_pad ,
		_w8955_,
		_w8956_,
		_w16586_
	);
	LUT3 #(
		.INIT('h80)
	) name14686 (
		\m6_data_i[9]_pad ,
		_w8955_,
		_w8956_,
		_w16587_
	);
	LUT3 #(
		.INIT('h57)
	) name14687 (
		_w8968_,
		_w16586_,
		_w16587_,
		_w16588_
	);
	LUT3 #(
		.INIT('h2a)
	) name14688 (
		\m3_data_i[9]_pad ,
		_w8955_,
		_w8956_,
		_w16589_
	);
	LUT3 #(
		.INIT('h80)
	) name14689 (
		\m4_data_i[9]_pad ,
		_w8955_,
		_w8956_,
		_w16590_
	);
	LUT4 #(
		.INIT('h9dbf)
	) name14690 (
		_w8950_,
		_w8953_,
		_w16589_,
		_w16590_,
		_w16591_
	);
	LUT4 #(
		.INIT('h7fff)
	) name14691 (
		_w16582_,
		_w16585_,
		_w16588_,
		_w16591_,
		_w16592_
	);
	LUT3 #(
		.INIT('h80)
	) name14692 (
		\m6_sel_i[0]_pad ,
		_w8955_,
		_w8956_,
		_w16593_
	);
	LUT3 #(
		.INIT('h2a)
	) name14693 (
		\m5_sel_i[0]_pad ,
		_w8955_,
		_w8956_,
		_w16594_
	);
	LUT4 #(
		.INIT('hcdef)
	) name14694 (
		_w8950_,
		_w8953_,
		_w16593_,
		_w16594_,
		_w16595_
	);
	LUT3 #(
		.INIT('h80)
	) name14695 (
		\m0_sel_i[0]_pad ,
		_w8955_,
		_w8956_,
		_w16596_
	);
	LUT3 #(
		.INIT('h80)
	) name14696 (
		\m4_sel_i[0]_pad ,
		_w8955_,
		_w8956_,
		_w16597_
	);
	LUT4 #(
		.INIT('h5d7f)
	) name14697 (
		_w8950_,
		_w8953_,
		_w16596_,
		_w16597_,
		_w16598_
	);
	LUT3 #(
		.INIT('h2a)
	) name14698 (
		\m7_sel_i[0]_pad ,
		_w8955_,
		_w8956_,
		_w16599_
	);
	LUT3 #(
		.INIT('h2a)
	) name14699 (
		\m3_sel_i[0]_pad ,
		_w8955_,
		_w8956_,
		_w16600_
	);
	LUT4 #(
		.INIT('habef)
	) name14700 (
		_w8950_,
		_w8953_,
		_w16599_,
		_w16600_,
		_w16601_
	);
	LUT3 #(
		.INIT('h2a)
	) name14701 (
		\m1_sel_i[0]_pad ,
		_w8955_,
		_w8956_,
		_w16602_
	);
	LUT3 #(
		.INIT('h80)
	) name14702 (
		\m2_sel_i[0]_pad ,
		_w8955_,
		_w8956_,
		_w16603_
	);
	LUT4 #(
		.INIT('h3b7f)
	) name14703 (
		_w8950_,
		_w8953_,
		_w16602_,
		_w16603_,
		_w16604_
	);
	LUT4 #(
		.INIT('h7fff)
	) name14704 (
		_w16595_,
		_w16598_,
		_w16601_,
		_w16604_,
		_w16605_
	);
	LUT3 #(
		.INIT('h80)
	) name14705 (
		\m0_sel_i[1]_pad ,
		_w8955_,
		_w8956_,
		_w16606_
	);
	LUT3 #(
		.INIT('h2a)
	) name14706 (
		\m7_sel_i[1]_pad ,
		_w8955_,
		_w8956_,
		_w16607_
	);
	LUT4 #(
		.INIT('h6e7f)
	) name14707 (
		_w8950_,
		_w8953_,
		_w16606_,
		_w16607_,
		_w16608_
	);
	LUT3 #(
		.INIT('h2a)
	) name14708 (
		\m1_sel_i[1]_pad ,
		_w8955_,
		_w8956_,
		_w16609_
	);
	LUT3 #(
		.INIT('h80)
	) name14709 (
		\m4_sel_i[1]_pad ,
		_w8955_,
		_w8956_,
		_w16610_
	);
	LUT4 #(
		.INIT('h5d7f)
	) name14710 (
		_w8950_,
		_w8953_,
		_w16609_,
		_w16610_,
		_w16611_
	);
	LUT3 #(
		.INIT('h80)
	) name14711 (
		\m2_sel_i[1]_pad ,
		_w8955_,
		_w8956_,
		_w16612_
	);
	LUT3 #(
		.INIT('h2a)
	) name14712 (
		\m3_sel_i[1]_pad ,
		_w8955_,
		_w8956_,
		_w16613_
	);
	LUT3 #(
		.INIT('h57)
	) name14713 (
		_w8974_,
		_w16612_,
		_w16613_,
		_w16614_
	);
	LUT3 #(
		.INIT('h80)
	) name14714 (
		\m6_sel_i[1]_pad ,
		_w8955_,
		_w8956_,
		_w16615_
	);
	LUT3 #(
		.INIT('h2a)
	) name14715 (
		\m5_sel_i[1]_pad ,
		_w8955_,
		_w8956_,
		_w16616_
	);
	LUT4 #(
		.INIT('hcdef)
	) name14716 (
		_w8950_,
		_w8953_,
		_w16615_,
		_w16616_,
		_w16617_
	);
	LUT4 #(
		.INIT('h7fff)
	) name14717 (
		_w16608_,
		_w16611_,
		_w16614_,
		_w16617_,
		_w16618_
	);
	LUT3 #(
		.INIT('h2a)
	) name14718 (
		\m3_sel_i[2]_pad ,
		_w8955_,
		_w8956_,
		_w16619_
	);
	LUT3 #(
		.INIT('h80)
	) name14719 (
		\m4_sel_i[2]_pad ,
		_w8955_,
		_w8956_,
		_w16620_
	);
	LUT4 #(
		.INIT('h9dbf)
	) name14720 (
		_w8950_,
		_w8953_,
		_w16619_,
		_w16620_,
		_w16621_
	);
	LUT3 #(
		.INIT('h80)
	) name14721 (
		\m0_sel_i[2]_pad ,
		_w8955_,
		_w8956_,
		_w16622_
	);
	LUT3 #(
		.INIT('h80)
	) name14722 (
		\m2_sel_i[2]_pad ,
		_w8955_,
		_w8956_,
		_w16623_
	);
	LUT4 #(
		.INIT('h3b7f)
	) name14723 (
		_w8950_,
		_w8953_,
		_w16622_,
		_w16623_,
		_w16624_
	);
	LUT3 #(
		.INIT('h2a)
	) name14724 (
		\m7_sel_i[2]_pad ,
		_w8955_,
		_w8956_,
		_w16625_
	);
	LUT3 #(
		.INIT('h2a)
	) name14725 (
		\m1_sel_i[2]_pad ,
		_w8955_,
		_w8956_,
		_w16626_
	);
	LUT4 #(
		.INIT('h67ef)
	) name14726 (
		_w8950_,
		_w8953_,
		_w16625_,
		_w16626_,
		_w16627_
	);
	LUT3 #(
		.INIT('h80)
	) name14727 (
		\m6_sel_i[2]_pad ,
		_w8955_,
		_w8956_,
		_w16628_
	);
	LUT3 #(
		.INIT('h2a)
	) name14728 (
		\m5_sel_i[2]_pad ,
		_w8955_,
		_w8956_,
		_w16629_
	);
	LUT4 #(
		.INIT('hcdef)
	) name14729 (
		_w8950_,
		_w8953_,
		_w16628_,
		_w16629_,
		_w16630_
	);
	LUT4 #(
		.INIT('h7fff)
	) name14730 (
		_w16621_,
		_w16624_,
		_w16627_,
		_w16630_,
		_w16631_
	);
	LUT3 #(
		.INIT('h2a)
	) name14731 (
		\m3_sel_i[3]_pad ,
		_w8955_,
		_w8956_,
		_w16632_
	);
	LUT3 #(
		.INIT('h80)
	) name14732 (
		\m4_sel_i[3]_pad ,
		_w8955_,
		_w8956_,
		_w16633_
	);
	LUT4 #(
		.INIT('h9dbf)
	) name14733 (
		_w8950_,
		_w8953_,
		_w16632_,
		_w16633_,
		_w16634_
	);
	LUT3 #(
		.INIT('h2a)
	) name14734 (
		\m1_sel_i[3]_pad ,
		_w8955_,
		_w8956_,
		_w16635_
	);
	LUT3 #(
		.INIT('h2a)
	) name14735 (
		\m5_sel_i[3]_pad ,
		_w8955_,
		_w8956_,
		_w16636_
	);
	LUT4 #(
		.INIT('h5d7f)
	) name14736 (
		_w8950_,
		_w8953_,
		_w16635_,
		_w16636_,
		_w16637_
	);
	LUT3 #(
		.INIT('h80)
	) name14737 (
		\m2_sel_i[3]_pad ,
		_w8955_,
		_w8956_,
		_w16638_
	);
	LUT3 #(
		.INIT('h80)
	) name14738 (
		\m6_sel_i[3]_pad ,
		_w8955_,
		_w8956_,
		_w16639_
	);
	LUT4 #(
		.INIT('haebf)
	) name14739 (
		_w8950_,
		_w8953_,
		_w16638_,
		_w16639_,
		_w16640_
	);
	LUT3 #(
		.INIT('h80)
	) name14740 (
		\m0_sel_i[3]_pad ,
		_w8955_,
		_w8956_,
		_w16641_
	);
	LUT3 #(
		.INIT('h2a)
	) name14741 (
		\m7_sel_i[3]_pad ,
		_w8955_,
		_w8956_,
		_w16642_
	);
	LUT4 #(
		.INIT('h6e7f)
	) name14742 (
		_w8950_,
		_w8953_,
		_w16641_,
		_w16642_,
		_w16643_
	);
	LUT4 #(
		.INIT('h7fff)
	) name14743 (
		_w16634_,
		_w16637_,
		_w16640_,
		_w16643_,
		_w16644_
	);
	LUT4 #(
		.INIT('h2a00)
	) name14744 (
		\m3_stb_i_pad ,
		_w8955_,
		_w8956_,
		_w9483_,
		_w16645_
	);
	LUT4 #(
		.INIT('h2a00)
	) name14745 (
		\m1_stb_i_pad ,
		_w8955_,
		_w8956_,
		_w9638_,
		_w16646_
	);
	LUT4 #(
		.INIT('h37bf)
	) name14746 (
		_w8950_,
		_w8953_,
		_w16645_,
		_w16646_,
		_w16647_
	);
	LUT4 #(
		.INIT('h8000)
	) name14747 (
		\m4_stb_i_pad ,
		_w8955_,
		_w8956_,
		_w9372_,
		_w16648_
	);
	LUT4 #(
		.INIT('h2a00)
	) name14748 (
		\m5_stb_i_pad ,
		_w8955_,
		_w8956_,
		_w9535_,
		_w16649_
	);
	LUT3 #(
		.INIT('h57)
	) name14749 (
		_w8954_,
		_w16648_,
		_w16649_,
		_w16650_
	);
	LUT4 #(
		.INIT('h8000)
	) name14750 (
		\m2_stb_i_pad ,
		_w8955_,
		_w8956_,
		_w9454_,
		_w16651_
	);
	LUT4 #(
		.INIT('h2a00)
	) name14751 (
		\m7_stb_i_pad ,
		_w8955_,
		_w8956_,
		_w9597_,
		_w16652_
	);
	LUT4 #(
		.INIT('haebf)
	) name14752 (
		_w8950_,
		_w8953_,
		_w16651_,
		_w16652_,
		_w16653_
	);
	LUT4 #(
		.INIT('h8000)
	) name14753 (
		\m6_stb_i_pad ,
		_w8955_,
		_w8956_,
		_w9562_,
		_w16654_
	);
	LUT4 #(
		.INIT('h8000)
	) name14754 (
		\m0_stb_i_pad ,
		_w8955_,
		_w8956_,
		_w9384_,
		_w16655_
	);
	LUT4 #(
		.INIT('h67ef)
	) name14755 (
		_w8950_,
		_w8953_,
		_w16654_,
		_w16655_,
		_w16656_
	);
	LUT4 #(
		.INIT('h7fff)
	) name14756 (
		_w16647_,
		_w16650_,
		_w16653_,
		_w16656_,
		_w16657_
	);
	LUT3 #(
		.INIT('h80)
	) name14757 (
		\m6_we_i_pad ,
		_w8955_,
		_w8956_,
		_w16658_
	);
	LUT3 #(
		.INIT('h2a)
	) name14758 (
		\m5_we_i_pad ,
		_w8955_,
		_w8956_,
		_w16659_
	);
	LUT4 #(
		.INIT('hcdef)
	) name14759 (
		_w8950_,
		_w8953_,
		_w16658_,
		_w16659_,
		_w16660_
	);
	LUT3 #(
		.INIT('h2a)
	) name14760 (
		\m3_we_i_pad ,
		_w8955_,
		_w8956_,
		_w16661_
	);
	LUT3 #(
		.INIT('h2a)
	) name14761 (
		\m7_we_i_pad ,
		_w8955_,
		_w8956_,
		_w16662_
	);
	LUT4 #(
		.INIT('haebf)
	) name14762 (
		_w8950_,
		_w8953_,
		_w16661_,
		_w16662_,
		_w16663_
	);
	LUT3 #(
		.INIT('h80)
	) name14763 (
		\m4_we_i_pad ,
		_w8955_,
		_w8956_,
		_w16664_
	);
	LUT3 #(
		.INIT('h80)
	) name14764 (
		\m0_we_i_pad ,
		_w8955_,
		_w8956_,
		_w16665_
	);
	LUT4 #(
		.INIT('h57df)
	) name14765 (
		_w8950_,
		_w8953_,
		_w16664_,
		_w16665_,
		_w16666_
	);
	LUT3 #(
		.INIT('h2a)
	) name14766 (
		\m1_we_i_pad ,
		_w8955_,
		_w8956_,
		_w16667_
	);
	LUT3 #(
		.INIT('h80)
	) name14767 (
		\m2_we_i_pad ,
		_w8955_,
		_w8956_,
		_w16668_
	);
	LUT4 #(
		.INIT('h3b7f)
	) name14768 (
		_w8950_,
		_w8953_,
		_w16667_,
		_w16668_,
		_w16669_
	);
	LUT4 #(
		.INIT('h7fff)
	) name14769 (
		_w16660_,
		_w16663_,
		_w16666_,
		_w16669_,
		_w16670_
	);
	LUT3 #(
		.INIT('h2a)
	) name14770 (
		\m3_addr_i[0]_pad ,
		_w9029_,
		_w9030_,
		_w16671_
	);
	LUT3 #(
		.INIT('h80)
	) name14771 (
		\m4_addr_i[0]_pad ,
		_w9029_,
		_w9030_,
		_w16672_
	);
	LUT4 #(
		.INIT('h9dbf)
	) name14772 (
		_w9024_,
		_w9027_,
		_w16671_,
		_w16672_,
		_w16673_
	);
	LUT3 #(
		.INIT('h80)
	) name14773 (
		\m6_addr_i[0]_pad ,
		_w9029_,
		_w9030_,
		_w16674_
	);
	LUT3 #(
		.INIT('h80)
	) name14774 (
		\m2_addr_i[0]_pad ,
		_w9029_,
		_w9030_,
		_w16675_
	);
	LUT4 #(
		.INIT('habef)
	) name14775 (
		_w9024_,
		_w9027_,
		_w16674_,
		_w16675_,
		_w16676_
	);
	LUT3 #(
		.INIT('h2a)
	) name14776 (
		\m5_addr_i[0]_pad ,
		_w9029_,
		_w9030_,
		_w16677_
	);
	LUT3 #(
		.INIT('h2a)
	) name14777 (
		\m1_addr_i[0]_pad ,
		_w9029_,
		_w9030_,
		_w16678_
	);
	LUT4 #(
		.INIT('h57df)
	) name14778 (
		_w9024_,
		_w9027_,
		_w16677_,
		_w16678_,
		_w16679_
	);
	LUT3 #(
		.INIT('h80)
	) name14779 (
		\m0_addr_i[0]_pad ,
		_w9029_,
		_w9030_,
		_w16680_
	);
	LUT3 #(
		.INIT('h2a)
	) name14780 (
		\m7_addr_i[0]_pad ,
		_w9029_,
		_w9030_,
		_w16681_
	);
	LUT4 #(
		.INIT('h6e7f)
	) name14781 (
		_w9024_,
		_w9027_,
		_w16680_,
		_w16681_,
		_w16682_
	);
	LUT4 #(
		.INIT('h7fff)
	) name14782 (
		_w16673_,
		_w16676_,
		_w16679_,
		_w16682_,
		_w16683_
	);
	LUT3 #(
		.INIT('h2a)
	) name14783 (
		\m3_addr_i[10]_pad ,
		_w9029_,
		_w9030_,
		_w16684_
	);
	LUT3 #(
		.INIT('h80)
	) name14784 (
		\m4_addr_i[10]_pad ,
		_w9029_,
		_w9030_,
		_w16685_
	);
	LUT4 #(
		.INIT('h9dbf)
	) name14785 (
		_w9024_,
		_w9027_,
		_w16684_,
		_w16685_,
		_w16686_
	);
	LUT3 #(
		.INIT('h2a)
	) name14786 (
		\m1_addr_i[10]_pad ,
		_w9029_,
		_w9030_,
		_w16687_
	);
	LUT3 #(
		.INIT('h2a)
	) name14787 (
		\m5_addr_i[10]_pad ,
		_w9029_,
		_w9030_,
		_w16688_
	);
	LUT4 #(
		.INIT('h5d7f)
	) name14788 (
		_w9024_,
		_w9027_,
		_w16687_,
		_w16688_,
		_w16689_
	);
	LUT3 #(
		.INIT('h80)
	) name14789 (
		\m2_addr_i[10]_pad ,
		_w9029_,
		_w9030_,
		_w16690_
	);
	LUT3 #(
		.INIT('h80)
	) name14790 (
		\m6_addr_i[10]_pad ,
		_w9029_,
		_w9030_,
		_w16691_
	);
	LUT4 #(
		.INIT('haebf)
	) name14791 (
		_w9024_,
		_w9027_,
		_w16690_,
		_w16691_,
		_w16692_
	);
	LUT3 #(
		.INIT('h80)
	) name14792 (
		\m0_addr_i[10]_pad ,
		_w9029_,
		_w9030_,
		_w16693_
	);
	LUT3 #(
		.INIT('h2a)
	) name14793 (
		\m7_addr_i[10]_pad ,
		_w9029_,
		_w9030_,
		_w16694_
	);
	LUT4 #(
		.INIT('h6e7f)
	) name14794 (
		_w9024_,
		_w9027_,
		_w16693_,
		_w16694_,
		_w16695_
	);
	LUT4 #(
		.INIT('h7fff)
	) name14795 (
		_w16686_,
		_w16689_,
		_w16692_,
		_w16695_,
		_w16696_
	);
	LUT3 #(
		.INIT('h2a)
	) name14796 (
		\m1_addr_i[11]_pad ,
		_w9029_,
		_w9030_,
		_w16697_
	);
	LUT3 #(
		.INIT('h80)
	) name14797 (
		\m2_addr_i[11]_pad ,
		_w9029_,
		_w9030_,
		_w16698_
	);
	LUT4 #(
		.INIT('h3b7f)
	) name14798 (
		_w9024_,
		_w9027_,
		_w16697_,
		_w16698_,
		_w16699_
	);
	LUT3 #(
		.INIT('h80)
	) name14799 (
		\m6_addr_i[11]_pad ,
		_w9029_,
		_w9030_,
		_w16700_
	);
	LUT3 #(
		.INIT('h2a)
	) name14800 (
		\m7_addr_i[11]_pad ,
		_w9029_,
		_w9030_,
		_w16701_
	);
	LUT3 #(
		.INIT('h57)
	) name14801 (
		_w9036_,
		_w16700_,
		_w16701_,
		_w16702_
	);
	LUT3 #(
		.INIT('h2a)
	) name14802 (
		\m5_addr_i[11]_pad ,
		_w9029_,
		_w9030_,
		_w16703_
	);
	LUT3 #(
		.INIT('h80)
	) name14803 (
		\m0_addr_i[11]_pad ,
		_w9029_,
		_w9030_,
		_w16704_
	);
	LUT4 #(
		.INIT('h57df)
	) name14804 (
		_w9024_,
		_w9027_,
		_w16703_,
		_w16704_,
		_w16705_
	);
	LUT3 #(
		.INIT('h2a)
	) name14805 (
		\m3_addr_i[11]_pad ,
		_w9029_,
		_w9030_,
		_w16706_
	);
	LUT3 #(
		.INIT('h80)
	) name14806 (
		\m4_addr_i[11]_pad ,
		_w9029_,
		_w9030_,
		_w16707_
	);
	LUT4 #(
		.INIT('h9dbf)
	) name14807 (
		_w9024_,
		_w9027_,
		_w16706_,
		_w16707_,
		_w16708_
	);
	LUT4 #(
		.INIT('h7fff)
	) name14808 (
		_w16699_,
		_w16702_,
		_w16705_,
		_w16708_,
		_w16709_
	);
	LUT3 #(
		.INIT('h80)
	) name14809 (
		\m0_addr_i[12]_pad ,
		_w9029_,
		_w9030_,
		_w16710_
	);
	LUT3 #(
		.INIT('h2a)
	) name14810 (
		\m7_addr_i[12]_pad ,
		_w9029_,
		_w9030_,
		_w16711_
	);
	LUT4 #(
		.INIT('h6e7f)
	) name14811 (
		_w9024_,
		_w9027_,
		_w16710_,
		_w16711_,
		_w16712_
	);
	LUT3 #(
		.INIT('h80)
	) name14812 (
		\m6_addr_i[12]_pad ,
		_w9029_,
		_w9030_,
		_w16713_
	);
	LUT3 #(
		.INIT('h80)
	) name14813 (
		\m2_addr_i[12]_pad ,
		_w9029_,
		_w9030_,
		_w16714_
	);
	LUT4 #(
		.INIT('habef)
	) name14814 (
		_w9024_,
		_w9027_,
		_w16713_,
		_w16714_,
		_w16715_
	);
	LUT3 #(
		.INIT('h2a)
	) name14815 (
		\m5_addr_i[12]_pad ,
		_w9029_,
		_w9030_,
		_w16716_
	);
	LUT3 #(
		.INIT('h2a)
	) name14816 (
		\m1_addr_i[12]_pad ,
		_w9029_,
		_w9030_,
		_w16717_
	);
	LUT4 #(
		.INIT('h57df)
	) name14817 (
		_w9024_,
		_w9027_,
		_w16716_,
		_w16717_,
		_w16718_
	);
	LUT3 #(
		.INIT('h2a)
	) name14818 (
		\m3_addr_i[12]_pad ,
		_w9029_,
		_w9030_,
		_w16719_
	);
	LUT3 #(
		.INIT('h80)
	) name14819 (
		\m4_addr_i[12]_pad ,
		_w9029_,
		_w9030_,
		_w16720_
	);
	LUT4 #(
		.INIT('h9dbf)
	) name14820 (
		_w9024_,
		_w9027_,
		_w16719_,
		_w16720_,
		_w16721_
	);
	LUT4 #(
		.INIT('h7fff)
	) name14821 (
		_w16712_,
		_w16715_,
		_w16718_,
		_w16721_,
		_w16722_
	);
	LUT3 #(
		.INIT('h2a)
	) name14822 (
		\m3_addr_i[13]_pad ,
		_w9029_,
		_w9030_,
		_w16723_
	);
	LUT3 #(
		.INIT('h80)
	) name14823 (
		\m4_addr_i[13]_pad ,
		_w9029_,
		_w9030_,
		_w16724_
	);
	LUT4 #(
		.INIT('h9dbf)
	) name14824 (
		_w9024_,
		_w9027_,
		_w16723_,
		_w16724_,
		_w16725_
	);
	LUT3 #(
		.INIT('h80)
	) name14825 (
		\m6_addr_i[13]_pad ,
		_w9029_,
		_w9030_,
		_w16726_
	);
	LUT3 #(
		.INIT('h80)
	) name14826 (
		\m2_addr_i[13]_pad ,
		_w9029_,
		_w9030_,
		_w16727_
	);
	LUT4 #(
		.INIT('habef)
	) name14827 (
		_w9024_,
		_w9027_,
		_w16726_,
		_w16727_,
		_w16728_
	);
	LUT3 #(
		.INIT('h2a)
	) name14828 (
		\m5_addr_i[13]_pad ,
		_w9029_,
		_w9030_,
		_w16729_
	);
	LUT3 #(
		.INIT('h2a)
	) name14829 (
		\m1_addr_i[13]_pad ,
		_w9029_,
		_w9030_,
		_w16730_
	);
	LUT4 #(
		.INIT('h57df)
	) name14830 (
		_w9024_,
		_w9027_,
		_w16729_,
		_w16730_,
		_w16731_
	);
	LUT3 #(
		.INIT('h80)
	) name14831 (
		\m0_addr_i[13]_pad ,
		_w9029_,
		_w9030_,
		_w16732_
	);
	LUT3 #(
		.INIT('h2a)
	) name14832 (
		\m7_addr_i[13]_pad ,
		_w9029_,
		_w9030_,
		_w16733_
	);
	LUT4 #(
		.INIT('h6e7f)
	) name14833 (
		_w9024_,
		_w9027_,
		_w16732_,
		_w16733_,
		_w16734_
	);
	LUT4 #(
		.INIT('h7fff)
	) name14834 (
		_w16725_,
		_w16728_,
		_w16731_,
		_w16734_,
		_w16735_
	);
	LUT3 #(
		.INIT('h2a)
	) name14835 (
		\m3_addr_i[14]_pad ,
		_w9029_,
		_w9030_,
		_w16736_
	);
	LUT3 #(
		.INIT('h80)
	) name14836 (
		\m4_addr_i[14]_pad ,
		_w9029_,
		_w9030_,
		_w16737_
	);
	LUT4 #(
		.INIT('h9dbf)
	) name14837 (
		_w9024_,
		_w9027_,
		_w16736_,
		_w16737_,
		_w16738_
	);
	LUT3 #(
		.INIT('h80)
	) name14838 (
		\m6_addr_i[14]_pad ,
		_w9029_,
		_w9030_,
		_w16739_
	);
	LUT3 #(
		.INIT('h80)
	) name14839 (
		\m2_addr_i[14]_pad ,
		_w9029_,
		_w9030_,
		_w16740_
	);
	LUT4 #(
		.INIT('habef)
	) name14840 (
		_w9024_,
		_w9027_,
		_w16739_,
		_w16740_,
		_w16741_
	);
	LUT3 #(
		.INIT('h2a)
	) name14841 (
		\m5_addr_i[14]_pad ,
		_w9029_,
		_w9030_,
		_w16742_
	);
	LUT3 #(
		.INIT('h2a)
	) name14842 (
		\m1_addr_i[14]_pad ,
		_w9029_,
		_w9030_,
		_w16743_
	);
	LUT4 #(
		.INIT('h57df)
	) name14843 (
		_w9024_,
		_w9027_,
		_w16742_,
		_w16743_,
		_w16744_
	);
	LUT3 #(
		.INIT('h80)
	) name14844 (
		\m0_addr_i[14]_pad ,
		_w9029_,
		_w9030_,
		_w16745_
	);
	LUT3 #(
		.INIT('h2a)
	) name14845 (
		\m7_addr_i[14]_pad ,
		_w9029_,
		_w9030_,
		_w16746_
	);
	LUT4 #(
		.INIT('h6e7f)
	) name14846 (
		_w9024_,
		_w9027_,
		_w16745_,
		_w16746_,
		_w16747_
	);
	LUT4 #(
		.INIT('h7fff)
	) name14847 (
		_w16738_,
		_w16741_,
		_w16744_,
		_w16747_,
		_w16748_
	);
	LUT3 #(
		.INIT('h2a)
	) name14848 (
		\m3_addr_i[15]_pad ,
		_w9029_,
		_w9030_,
		_w16749_
	);
	LUT3 #(
		.INIT('h80)
	) name14849 (
		\m4_addr_i[15]_pad ,
		_w9029_,
		_w9030_,
		_w16750_
	);
	LUT4 #(
		.INIT('h9dbf)
	) name14850 (
		_w9024_,
		_w9027_,
		_w16749_,
		_w16750_,
		_w16751_
	);
	LUT3 #(
		.INIT('h80)
	) name14851 (
		\m6_addr_i[15]_pad ,
		_w9029_,
		_w9030_,
		_w16752_
	);
	LUT3 #(
		.INIT('h80)
	) name14852 (
		\m2_addr_i[15]_pad ,
		_w9029_,
		_w9030_,
		_w16753_
	);
	LUT4 #(
		.INIT('habef)
	) name14853 (
		_w9024_,
		_w9027_,
		_w16752_,
		_w16753_,
		_w16754_
	);
	LUT3 #(
		.INIT('h2a)
	) name14854 (
		\m5_addr_i[15]_pad ,
		_w9029_,
		_w9030_,
		_w16755_
	);
	LUT3 #(
		.INIT('h2a)
	) name14855 (
		\m1_addr_i[15]_pad ,
		_w9029_,
		_w9030_,
		_w16756_
	);
	LUT4 #(
		.INIT('h57df)
	) name14856 (
		_w9024_,
		_w9027_,
		_w16755_,
		_w16756_,
		_w16757_
	);
	LUT3 #(
		.INIT('h80)
	) name14857 (
		\m0_addr_i[15]_pad ,
		_w9029_,
		_w9030_,
		_w16758_
	);
	LUT3 #(
		.INIT('h2a)
	) name14858 (
		\m7_addr_i[15]_pad ,
		_w9029_,
		_w9030_,
		_w16759_
	);
	LUT4 #(
		.INIT('h6e7f)
	) name14859 (
		_w9024_,
		_w9027_,
		_w16758_,
		_w16759_,
		_w16760_
	);
	LUT4 #(
		.INIT('h7fff)
	) name14860 (
		_w16751_,
		_w16754_,
		_w16757_,
		_w16760_,
		_w16761_
	);
	LUT3 #(
		.INIT('h2a)
	) name14861 (
		\m3_addr_i[16]_pad ,
		_w9029_,
		_w9030_,
		_w16762_
	);
	LUT3 #(
		.INIT('h80)
	) name14862 (
		\m4_addr_i[16]_pad ,
		_w9029_,
		_w9030_,
		_w16763_
	);
	LUT4 #(
		.INIT('h9dbf)
	) name14863 (
		_w9024_,
		_w9027_,
		_w16762_,
		_w16763_,
		_w16764_
	);
	LUT3 #(
		.INIT('h80)
	) name14864 (
		\m6_addr_i[16]_pad ,
		_w9029_,
		_w9030_,
		_w16765_
	);
	LUT3 #(
		.INIT('h80)
	) name14865 (
		\m2_addr_i[16]_pad ,
		_w9029_,
		_w9030_,
		_w16766_
	);
	LUT4 #(
		.INIT('habef)
	) name14866 (
		_w9024_,
		_w9027_,
		_w16765_,
		_w16766_,
		_w16767_
	);
	LUT3 #(
		.INIT('h2a)
	) name14867 (
		\m5_addr_i[16]_pad ,
		_w9029_,
		_w9030_,
		_w16768_
	);
	LUT3 #(
		.INIT('h2a)
	) name14868 (
		\m1_addr_i[16]_pad ,
		_w9029_,
		_w9030_,
		_w16769_
	);
	LUT4 #(
		.INIT('h57df)
	) name14869 (
		_w9024_,
		_w9027_,
		_w16768_,
		_w16769_,
		_w16770_
	);
	LUT3 #(
		.INIT('h80)
	) name14870 (
		\m0_addr_i[16]_pad ,
		_w9029_,
		_w9030_,
		_w16771_
	);
	LUT3 #(
		.INIT('h2a)
	) name14871 (
		\m7_addr_i[16]_pad ,
		_w9029_,
		_w9030_,
		_w16772_
	);
	LUT4 #(
		.INIT('h6e7f)
	) name14872 (
		_w9024_,
		_w9027_,
		_w16771_,
		_w16772_,
		_w16773_
	);
	LUT4 #(
		.INIT('h7fff)
	) name14873 (
		_w16764_,
		_w16767_,
		_w16770_,
		_w16773_,
		_w16774_
	);
	LUT3 #(
		.INIT('h2a)
	) name14874 (
		\m3_addr_i[17]_pad ,
		_w9029_,
		_w9030_,
		_w16775_
	);
	LUT3 #(
		.INIT('h80)
	) name14875 (
		\m4_addr_i[17]_pad ,
		_w9029_,
		_w9030_,
		_w16776_
	);
	LUT4 #(
		.INIT('h9dbf)
	) name14876 (
		_w9024_,
		_w9027_,
		_w16775_,
		_w16776_,
		_w16777_
	);
	LUT3 #(
		.INIT('h80)
	) name14877 (
		\m6_addr_i[17]_pad ,
		_w9029_,
		_w9030_,
		_w16778_
	);
	LUT3 #(
		.INIT('h80)
	) name14878 (
		\m2_addr_i[17]_pad ,
		_w9029_,
		_w9030_,
		_w16779_
	);
	LUT4 #(
		.INIT('habef)
	) name14879 (
		_w9024_,
		_w9027_,
		_w16778_,
		_w16779_,
		_w16780_
	);
	LUT3 #(
		.INIT('h2a)
	) name14880 (
		\m5_addr_i[17]_pad ,
		_w9029_,
		_w9030_,
		_w16781_
	);
	LUT3 #(
		.INIT('h2a)
	) name14881 (
		\m1_addr_i[17]_pad ,
		_w9029_,
		_w9030_,
		_w16782_
	);
	LUT4 #(
		.INIT('h57df)
	) name14882 (
		_w9024_,
		_w9027_,
		_w16781_,
		_w16782_,
		_w16783_
	);
	LUT3 #(
		.INIT('h80)
	) name14883 (
		\m0_addr_i[17]_pad ,
		_w9029_,
		_w9030_,
		_w16784_
	);
	LUT3 #(
		.INIT('h2a)
	) name14884 (
		\m7_addr_i[17]_pad ,
		_w9029_,
		_w9030_,
		_w16785_
	);
	LUT4 #(
		.INIT('h6e7f)
	) name14885 (
		_w9024_,
		_w9027_,
		_w16784_,
		_w16785_,
		_w16786_
	);
	LUT4 #(
		.INIT('h7fff)
	) name14886 (
		_w16777_,
		_w16780_,
		_w16783_,
		_w16786_,
		_w16787_
	);
	LUT3 #(
		.INIT('h2a)
	) name14887 (
		\m1_addr_i[18]_pad ,
		_w9029_,
		_w9030_,
		_w16788_
	);
	LUT3 #(
		.INIT('h80)
	) name14888 (
		\m2_addr_i[18]_pad ,
		_w9029_,
		_w9030_,
		_w16789_
	);
	LUT4 #(
		.INIT('h3b7f)
	) name14889 (
		_w9024_,
		_w9027_,
		_w16788_,
		_w16789_,
		_w16790_
	);
	LUT3 #(
		.INIT('h80)
	) name14890 (
		\m6_addr_i[18]_pad ,
		_w9029_,
		_w9030_,
		_w16791_
	);
	LUT3 #(
		.INIT('h2a)
	) name14891 (
		\m7_addr_i[18]_pad ,
		_w9029_,
		_w9030_,
		_w16792_
	);
	LUT3 #(
		.INIT('h57)
	) name14892 (
		_w9036_,
		_w16791_,
		_w16792_,
		_w16793_
	);
	LUT3 #(
		.INIT('h2a)
	) name14893 (
		\m5_addr_i[18]_pad ,
		_w9029_,
		_w9030_,
		_w16794_
	);
	LUT3 #(
		.INIT('h80)
	) name14894 (
		\m0_addr_i[18]_pad ,
		_w9029_,
		_w9030_,
		_w16795_
	);
	LUT4 #(
		.INIT('h57df)
	) name14895 (
		_w9024_,
		_w9027_,
		_w16794_,
		_w16795_,
		_w16796_
	);
	LUT3 #(
		.INIT('h2a)
	) name14896 (
		\m3_addr_i[18]_pad ,
		_w9029_,
		_w9030_,
		_w16797_
	);
	LUT3 #(
		.INIT('h80)
	) name14897 (
		\m4_addr_i[18]_pad ,
		_w9029_,
		_w9030_,
		_w16798_
	);
	LUT4 #(
		.INIT('h9dbf)
	) name14898 (
		_w9024_,
		_w9027_,
		_w16797_,
		_w16798_,
		_w16799_
	);
	LUT4 #(
		.INIT('h7fff)
	) name14899 (
		_w16790_,
		_w16793_,
		_w16796_,
		_w16799_,
		_w16800_
	);
	LUT3 #(
		.INIT('h80)
	) name14900 (
		\m0_addr_i[19]_pad ,
		_w9029_,
		_w9030_,
		_w16801_
	);
	LUT3 #(
		.INIT('h2a)
	) name14901 (
		\m7_addr_i[19]_pad ,
		_w9029_,
		_w9030_,
		_w16802_
	);
	LUT4 #(
		.INIT('h6e7f)
	) name14902 (
		_w9024_,
		_w9027_,
		_w16801_,
		_w16802_,
		_w16803_
	);
	LUT3 #(
		.INIT('h80)
	) name14903 (
		\m6_addr_i[19]_pad ,
		_w9029_,
		_w9030_,
		_w16804_
	);
	LUT3 #(
		.INIT('h80)
	) name14904 (
		\m4_addr_i[19]_pad ,
		_w9029_,
		_w9030_,
		_w16805_
	);
	LUT4 #(
		.INIT('hcdef)
	) name14905 (
		_w9024_,
		_w9027_,
		_w16804_,
		_w16805_,
		_w16806_
	);
	LUT3 #(
		.INIT('h2a)
	) name14906 (
		\m5_addr_i[19]_pad ,
		_w9029_,
		_w9030_,
		_w16807_
	);
	LUT3 #(
		.INIT('h2a)
	) name14907 (
		\m3_addr_i[19]_pad ,
		_w9029_,
		_w9030_,
		_w16808_
	);
	LUT4 #(
		.INIT('h9bdf)
	) name14908 (
		_w9024_,
		_w9027_,
		_w16807_,
		_w16808_,
		_w16809_
	);
	LUT3 #(
		.INIT('h2a)
	) name14909 (
		\m1_addr_i[19]_pad ,
		_w9029_,
		_w9030_,
		_w16810_
	);
	LUT3 #(
		.INIT('h80)
	) name14910 (
		\m2_addr_i[19]_pad ,
		_w9029_,
		_w9030_,
		_w16811_
	);
	LUT4 #(
		.INIT('h3b7f)
	) name14911 (
		_w9024_,
		_w9027_,
		_w16810_,
		_w16811_,
		_w16812_
	);
	LUT4 #(
		.INIT('h7fff)
	) name14912 (
		_w16803_,
		_w16806_,
		_w16809_,
		_w16812_,
		_w16813_
	);
	LUT3 #(
		.INIT('h2a)
	) name14913 (
		\m3_addr_i[1]_pad ,
		_w9029_,
		_w9030_,
		_w16814_
	);
	LUT3 #(
		.INIT('h80)
	) name14914 (
		\m4_addr_i[1]_pad ,
		_w9029_,
		_w9030_,
		_w16815_
	);
	LUT4 #(
		.INIT('h9dbf)
	) name14915 (
		_w9024_,
		_w9027_,
		_w16814_,
		_w16815_,
		_w16816_
	);
	LUT3 #(
		.INIT('h80)
	) name14916 (
		\m6_addr_i[1]_pad ,
		_w9029_,
		_w9030_,
		_w16817_
	);
	LUT3 #(
		.INIT('h80)
	) name14917 (
		\m2_addr_i[1]_pad ,
		_w9029_,
		_w9030_,
		_w16818_
	);
	LUT4 #(
		.INIT('habef)
	) name14918 (
		_w9024_,
		_w9027_,
		_w16817_,
		_w16818_,
		_w16819_
	);
	LUT3 #(
		.INIT('h2a)
	) name14919 (
		\m5_addr_i[1]_pad ,
		_w9029_,
		_w9030_,
		_w16820_
	);
	LUT3 #(
		.INIT('h2a)
	) name14920 (
		\m1_addr_i[1]_pad ,
		_w9029_,
		_w9030_,
		_w16821_
	);
	LUT4 #(
		.INIT('h57df)
	) name14921 (
		_w9024_,
		_w9027_,
		_w16820_,
		_w16821_,
		_w16822_
	);
	LUT3 #(
		.INIT('h80)
	) name14922 (
		\m0_addr_i[1]_pad ,
		_w9029_,
		_w9030_,
		_w16823_
	);
	LUT3 #(
		.INIT('h2a)
	) name14923 (
		\m7_addr_i[1]_pad ,
		_w9029_,
		_w9030_,
		_w16824_
	);
	LUT4 #(
		.INIT('h6e7f)
	) name14924 (
		_w9024_,
		_w9027_,
		_w16823_,
		_w16824_,
		_w16825_
	);
	LUT4 #(
		.INIT('h7fff)
	) name14925 (
		_w16816_,
		_w16819_,
		_w16822_,
		_w16825_,
		_w16826_
	);
	LUT3 #(
		.INIT('h80)
	) name14926 (
		\m6_addr_i[20]_pad ,
		_w9029_,
		_w9030_,
		_w16827_
	);
	LUT3 #(
		.INIT('h2a)
	) name14927 (
		\m5_addr_i[20]_pad ,
		_w9029_,
		_w9030_,
		_w16828_
	);
	LUT4 #(
		.INIT('hcdef)
	) name14928 (
		_w9024_,
		_w9027_,
		_w16827_,
		_w16828_,
		_w16829_
	);
	LUT3 #(
		.INIT('h2a)
	) name14929 (
		\m1_addr_i[20]_pad ,
		_w9029_,
		_w9030_,
		_w16830_
	);
	LUT3 #(
		.INIT('h80)
	) name14930 (
		\m4_addr_i[20]_pad ,
		_w9029_,
		_w9030_,
		_w16831_
	);
	LUT4 #(
		.INIT('h5d7f)
	) name14931 (
		_w9024_,
		_w9027_,
		_w16830_,
		_w16831_,
		_w16832_
	);
	LUT3 #(
		.INIT('h80)
	) name14932 (
		\m2_addr_i[20]_pad ,
		_w9029_,
		_w9030_,
		_w16833_
	);
	LUT3 #(
		.INIT('h2a)
	) name14933 (
		\m3_addr_i[20]_pad ,
		_w9029_,
		_w9030_,
		_w16834_
	);
	LUT3 #(
		.INIT('h57)
	) name14934 (
		_w9028_,
		_w16833_,
		_w16834_,
		_w16835_
	);
	LUT3 #(
		.INIT('h80)
	) name14935 (
		\m0_addr_i[20]_pad ,
		_w9029_,
		_w9030_,
		_w16836_
	);
	LUT3 #(
		.INIT('h2a)
	) name14936 (
		\m7_addr_i[20]_pad ,
		_w9029_,
		_w9030_,
		_w16837_
	);
	LUT4 #(
		.INIT('h6e7f)
	) name14937 (
		_w9024_,
		_w9027_,
		_w16836_,
		_w16837_,
		_w16838_
	);
	LUT4 #(
		.INIT('h7fff)
	) name14938 (
		_w16829_,
		_w16832_,
		_w16835_,
		_w16838_,
		_w16839_
	);
	LUT3 #(
		.INIT('h80)
	) name14939 (
		\m0_addr_i[21]_pad ,
		_w9029_,
		_w9030_,
		_w16840_
	);
	LUT3 #(
		.INIT('h2a)
	) name14940 (
		\m7_addr_i[21]_pad ,
		_w9029_,
		_w9030_,
		_w16841_
	);
	LUT4 #(
		.INIT('h6e7f)
	) name14941 (
		_w9024_,
		_w9027_,
		_w16840_,
		_w16841_,
		_w16842_
	);
	LUT3 #(
		.INIT('h2a)
	) name14942 (
		\m1_addr_i[21]_pad ,
		_w9029_,
		_w9030_,
		_w16843_
	);
	LUT3 #(
		.INIT('h80)
	) name14943 (
		\m4_addr_i[21]_pad ,
		_w9029_,
		_w9030_,
		_w16844_
	);
	LUT4 #(
		.INIT('h5d7f)
	) name14944 (
		_w9024_,
		_w9027_,
		_w16843_,
		_w16844_,
		_w16845_
	);
	LUT3 #(
		.INIT('h80)
	) name14945 (
		\m2_addr_i[21]_pad ,
		_w9029_,
		_w9030_,
		_w16846_
	);
	LUT3 #(
		.INIT('h2a)
	) name14946 (
		\m3_addr_i[21]_pad ,
		_w9029_,
		_w9030_,
		_w16847_
	);
	LUT3 #(
		.INIT('h57)
	) name14947 (
		_w9028_,
		_w16846_,
		_w16847_,
		_w16848_
	);
	LUT3 #(
		.INIT('h80)
	) name14948 (
		\m6_addr_i[21]_pad ,
		_w9029_,
		_w9030_,
		_w16849_
	);
	LUT3 #(
		.INIT('h2a)
	) name14949 (
		\m5_addr_i[21]_pad ,
		_w9029_,
		_w9030_,
		_w16850_
	);
	LUT4 #(
		.INIT('hcdef)
	) name14950 (
		_w9024_,
		_w9027_,
		_w16849_,
		_w16850_,
		_w16851_
	);
	LUT4 #(
		.INIT('h7fff)
	) name14951 (
		_w16842_,
		_w16845_,
		_w16848_,
		_w16851_,
		_w16852_
	);
	LUT3 #(
		.INIT('h80)
	) name14952 (
		\m0_addr_i[22]_pad ,
		_w9029_,
		_w9030_,
		_w16853_
	);
	LUT3 #(
		.INIT('h2a)
	) name14953 (
		\m7_addr_i[22]_pad ,
		_w9029_,
		_w9030_,
		_w16854_
	);
	LUT4 #(
		.INIT('h6e7f)
	) name14954 (
		_w9024_,
		_w9027_,
		_w16853_,
		_w16854_,
		_w16855_
	);
	LUT3 #(
		.INIT('h2a)
	) name14955 (
		\m3_addr_i[22]_pad ,
		_w9029_,
		_w9030_,
		_w16856_
	);
	LUT3 #(
		.INIT('h80)
	) name14956 (
		\m2_addr_i[22]_pad ,
		_w9029_,
		_w9030_,
		_w16857_
	);
	LUT3 #(
		.INIT('h57)
	) name14957 (
		_w9028_,
		_w16856_,
		_w16857_,
		_w16858_
	);
	LUT3 #(
		.INIT('h80)
	) name14958 (
		\m4_addr_i[22]_pad ,
		_w9029_,
		_w9030_,
		_w16859_
	);
	LUT3 #(
		.INIT('h2a)
	) name14959 (
		\m1_addr_i[22]_pad ,
		_w9029_,
		_w9030_,
		_w16860_
	);
	LUT4 #(
		.INIT('h57df)
	) name14960 (
		_w9024_,
		_w9027_,
		_w16859_,
		_w16860_,
		_w16861_
	);
	LUT3 #(
		.INIT('h80)
	) name14961 (
		\m6_addr_i[22]_pad ,
		_w9029_,
		_w9030_,
		_w16862_
	);
	LUT3 #(
		.INIT('h2a)
	) name14962 (
		\m5_addr_i[22]_pad ,
		_w9029_,
		_w9030_,
		_w16863_
	);
	LUT4 #(
		.INIT('hcdef)
	) name14963 (
		_w9024_,
		_w9027_,
		_w16862_,
		_w16863_,
		_w16864_
	);
	LUT4 #(
		.INIT('h7fff)
	) name14964 (
		_w16855_,
		_w16858_,
		_w16861_,
		_w16864_,
		_w16865_
	);
	LUT3 #(
		.INIT('h80)
	) name14965 (
		\m6_addr_i[23]_pad ,
		_w9029_,
		_w9030_,
		_w16866_
	);
	LUT3 #(
		.INIT('h2a)
	) name14966 (
		\m5_addr_i[23]_pad ,
		_w9029_,
		_w9030_,
		_w16867_
	);
	LUT4 #(
		.INIT('hcdef)
	) name14967 (
		_w9024_,
		_w9027_,
		_w16866_,
		_w16867_,
		_w16868_
	);
	LUT3 #(
		.INIT('h2a)
	) name14968 (
		\m3_addr_i[23]_pad ,
		_w9029_,
		_w9030_,
		_w16869_
	);
	LUT3 #(
		.INIT('h2a)
	) name14969 (
		\m7_addr_i[23]_pad ,
		_w9029_,
		_w9030_,
		_w16870_
	);
	LUT4 #(
		.INIT('haebf)
	) name14970 (
		_w9024_,
		_w9027_,
		_w16869_,
		_w16870_,
		_w16871_
	);
	LUT3 #(
		.INIT('h80)
	) name14971 (
		\m4_addr_i[23]_pad ,
		_w9029_,
		_w9030_,
		_w16872_
	);
	LUT3 #(
		.INIT('h80)
	) name14972 (
		\m0_addr_i[23]_pad ,
		_w9029_,
		_w9030_,
		_w16873_
	);
	LUT4 #(
		.INIT('h57df)
	) name14973 (
		_w9024_,
		_w9027_,
		_w16872_,
		_w16873_,
		_w16874_
	);
	LUT3 #(
		.INIT('h2a)
	) name14974 (
		\m1_addr_i[23]_pad ,
		_w9029_,
		_w9030_,
		_w16875_
	);
	LUT3 #(
		.INIT('h80)
	) name14975 (
		\m2_addr_i[23]_pad ,
		_w9029_,
		_w9030_,
		_w16876_
	);
	LUT4 #(
		.INIT('h3b7f)
	) name14976 (
		_w9024_,
		_w9027_,
		_w16875_,
		_w16876_,
		_w16877_
	);
	LUT4 #(
		.INIT('h7fff)
	) name14977 (
		_w16868_,
		_w16871_,
		_w16874_,
		_w16877_,
		_w16878_
	);
	LUT3 #(
		.INIT('h2a)
	) name14978 (
		\m3_addr_i[24]_pad ,
		_w9029_,
		_w9030_,
		_w16879_
	);
	LUT3 #(
		.INIT('h80)
	) name14979 (
		\m4_addr_i[24]_pad ,
		_w9029_,
		_w9030_,
		_w16880_
	);
	LUT4 #(
		.INIT('h9dbf)
	) name14980 (
		_w9024_,
		_w9027_,
		_w16879_,
		_w16880_,
		_w16881_
	);
	LUT3 #(
		.INIT('h2a)
	) name14981 (
		\m1_addr_i[24]_pad ,
		_w9029_,
		_w9030_,
		_w16882_
	);
	LUT3 #(
		.INIT('h80)
	) name14982 (
		\m6_addr_i[24]_pad ,
		_w9029_,
		_w9030_,
		_w16883_
	);
	LUT4 #(
		.INIT('h6e7f)
	) name14983 (
		_w9024_,
		_w9027_,
		_w16882_,
		_w16883_,
		_w16884_
	);
	LUT3 #(
		.INIT('h80)
	) name14984 (
		\m2_addr_i[24]_pad ,
		_w9029_,
		_w9030_,
		_w16885_
	);
	LUT3 #(
		.INIT('h2a)
	) name14985 (
		\m5_addr_i[24]_pad ,
		_w9029_,
		_w9030_,
		_w16886_
	);
	LUT4 #(
		.INIT('h9dbf)
	) name14986 (
		_w9024_,
		_w9027_,
		_w16885_,
		_w16886_,
		_w16887_
	);
	LUT3 #(
		.INIT('h80)
	) name14987 (
		\m0_addr_i[24]_pad ,
		_w9029_,
		_w9030_,
		_w16888_
	);
	LUT3 #(
		.INIT('h2a)
	) name14988 (
		\m7_addr_i[24]_pad ,
		_w9029_,
		_w9030_,
		_w16889_
	);
	LUT4 #(
		.INIT('h6e7f)
	) name14989 (
		_w9024_,
		_w9027_,
		_w16888_,
		_w16889_,
		_w16890_
	);
	LUT4 #(
		.INIT('h7fff)
	) name14990 (
		_w16881_,
		_w16884_,
		_w16887_,
		_w16890_,
		_w16891_
	);
	LUT3 #(
		.INIT('h80)
	) name14991 (
		\m0_addr_i[25]_pad ,
		_w9029_,
		_w9030_,
		_w16892_
	);
	LUT3 #(
		.INIT('h2a)
	) name14992 (
		\m7_addr_i[25]_pad ,
		_w9029_,
		_w9030_,
		_w16893_
	);
	LUT4 #(
		.INIT('h6e7f)
	) name14993 (
		_w9024_,
		_w9027_,
		_w16892_,
		_w16893_,
		_w16894_
	);
	LUT3 #(
		.INIT('h2a)
	) name14994 (
		\m3_addr_i[25]_pad ,
		_w9029_,
		_w9030_,
		_w16895_
	);
	LUT3 #(
		.INIT('h80)
	) name14995 (
		\m6_addr_i[25]_pad ,
		_w9029_,
		_w9030_,
		_w16896_
	);
	LUT4 #(
		.INIT('haebf)
	) name14996 (
		_w9024_,
		_w9027_,
		_w16895_,
		_w16896_,
		_w16897_
	);
	LUT3 #(
		.INIT('h80)
	) name14997 (
		\m4_addr_i[25]_pad ,
		_w9029_,
		_w9030_,
		_w16898_
	);
	LUT3 #(
		.INIT('h2a)
	) name14998 (
		\m5_addr_i[25]_pad ,
		_w9029_,
		_w9030_,
		_w16899_
	);
	LUT3 #(
		.INIT('h57)
	) name14999 (
		_w9042_,
		_w16898_,
		_w16899_,
		_w16900_
	);
	LUT3 #(
		.INIT('h2a)
	) name15000 (
		\m1_addr_i[25]_pad ,
		_w9029_,
		_w9030_,
		_w16901_
	);
	LUT3 #(
		.INIT('h80)
	) name15001 (
		\m2_addr_i[25]_pad ,
		_w9029_,
		_w9030_,
		_w16902_
	);
	LUT4 #(
		.INIT('h3b7f)
	) name15002 (
		_w9024_,
		_w9027_,
		_w16901_,
		_w16902_,
		_w16903_
	);
	LUT4 #(
		.INIT('h7fff)
	) name15003 (
		_w16894_,
		_w16897_,
		_w16900_,
		_w16903_,
		_w16904_
	);
	LUT3 #(
		.INIT('h2a)
	) name15004 (
		\m1_addr_i[26]_pad ,
		_w9029_,
		_w9030_,
		_w16905_
	);
	LUT3 #(
		.INIT('h80)
	) name15005 (
		\m2_addr_i[26]_pad ,
		_w9029_,
		_w9030_,
		_w16906_
	);
	LUT4 #(
		.INIT('h3b7f)
	) name15006 (
		_w9024_,
		_w9027_,
		_w16905_,
		_w16906_,
		_w16907_
	);
	LUT3 #(
		.INIT('h2a)
	) name15007 (
		\m3_addr_i[26]_pad ,
		_w9029_,
		_w9030_,
		_w16908_
	);
	LUT3 #(
		.INIT('h80)
	) name15008 (
		\m6_addr_i[26]_pad ,
		_w9029_,
		_w9030_,
		_w16909_
	);
	LUT4 #(
		.INIT('haebf)
	) name15009 (
		_w9024_,
		_w9027_,
		_w16908_,
		_w16909_,
		_w16910_
	);
	LUT3 #(
		.INIT('h80)
	) name15010 (
		\m4_addr_i[26]_pad ,
		_w9029_,
		_w9030_,
		_w16911_
	);
	LUT3 #(
		.INIT('h2a)
	) name15011 (
		\m5_addr_i[26]_pad ,
		_w9029_,
		_w9030_,
		_w16912_
	);
	LUT3 #(
		.INIT('h57)
	) name15012 (
		_w9042_,
		_w16911_,
		_w16912_,
		_w16913_
	);
	LUT3 #(
		.INIT('h80)
	) name15013 (
		\m0_addr_i[26]_pad ,
		_w9029_,
		_w9030_,
		_w16914_
	);
	LUT3 #(
		.INIT('h2a)
	) name15014 (
		\m7_addr_i[26]_pad ,
		_w9029_,
		_w9030_,
		_w16915_
	);
	LUT4 #(
		.INIT('h6e7f)
	) name15015 (
		_w9024_,
		_w9027_,
		_w16914_,
		_w16915_,
		_w16916_
	);
	LUT4 #(
		.INIT('h7fff)
	) name15016 (
		_w16907_,
		_w16910_,
		_w16913_,
		_w16916_,
		_w16917_
	);
	LUT3 #(
		.INIT('h2a)
	) name15017 (
		\m3_addr_i[27]_pad ,
		_w9029_,
		_w9030_,
		_w16918_
	);
	LUT3 #(
		.INIT('h80)
	) name15018 (
		\m4_addr_i[27]_pad ,
		_w9029_,
		_w9030_,
		_w16919_
	);
	LUT4 #(
		.INIT('h9dbf)
	) name15019 (
		_w9024_,
		_w9027_,
		_w16918_,
		_w16919_,
		_w16920_
	);
	LUT3 #(
		.INIT('h2a)
	) name15020 (
		\m5_addr_i[27]_pad ,
		_w9029_,
		_w9030_,
		_w16921_
	);
	LUT3 #(
		.INIT('h2a)
	) name15021 (
		\m7_addr_i[27]_pad ,
		_w9029_,
		_w9030_,
		_w16922_
	);
	LUT4 #(
		.INIT('hcedf)
	) name15022 (
		_w9024_,
		_w9027_,
		_w16921_,
		_w16922_,
		_w16923_
	);
	LUT3 #(
		.INIT('h80)
	) name15023 (
		\m6_addr_i[27]_pad ,
		_w9029_,
		_w9030_,
		_w16924_
	);
	LUT3 #(
		.INIT('h80)
	) name15024 (
		\m0_addr_i[27]_pad ,
		_w9029_,
		_w9030_,
		_w16925_
	);
	LUT4 #(
		.INIT('h67ef)
	) name15025 (
		_w9024_,
		_w9027_,
		_w16924_,
		_w16925_,
		_w16926_
	);
	LUT3 #(
		.INIT('h2a)
	) name15026 (
		\m1_addr_i[27]_pad ,
		_w9029_,
		_w9030_,
		_w16927_
	);
	LUT3 #(
		.INIT('h80)
	) name15027 (
		\m2_addr_i[27]_pad ,
		_w9029_,
		_w9030_,
		_w16928_
	);
	LUT4 #(
		.INIT('h3b7f)
	) name15028 (
		_w9024_,
		_w9027_,
		_w16927_,
		_w16928_,
		_w16929_
	);
	LUT4 #(
		.INIT('h7fff)
	) name15029 (
		_w16920_,
		_w16923_,
		_w16926_,
		_w16929_,
		_w16930_
	);
	LUT3 #(
		.INIT('h2a)
	) name15030 (
		\m1_addr_i[28]_pad ,
		_w9029_,
		_w9030_,
		_w16931_
	);
	LUT3 #(
		.INIT('h80)
	) name15031 (
		\m2_addr_i[28]_pad ,
		_w9029_,
		_w9030_,
		_w16932_
	);
	LUT4 #(
		.INIT('h3b7f)
	) name15032 (
		_w9024_,
		_w9027_,
		_w16931_,
		_w16932_,
		_w16933_
	);
	LUT3 #(
		.INIT('h2a)
	) name15033 (
		\m3_addr_i[28]_pad ,
		_w9029_,
		_w9030_,
		_w16934_
	);
	LUT3 #(
		.INIT('h2a)
	) name15034 (
		\m7_addr_i[28]_pad ,
		_w9029_,
		_w9030_,
		_w16935_
	);
	LUT4 #(
		.INIT('haebf)
	) name15035 (
		_w9024_,
		_w9027_,
		_w16934_,
		_w16935_,
		_w16936_
	);
	LUT3 #(
		.INIT('h80)
	) name15036 (
		\m4_addr_i[28]_pad ,
		_w9029_,
		_w9030_,
		_w16937_
	);
	LUT3 #(
		.INIT('h80)
	) name15037 (
		\m0_addr_i[28]_pad ,
		_w9029_,
		_w9030_,
		_w16938_
	);
	LUT4 #(
		.INIT('h57df)
	) name15038 (
		_w9024_,
		_w9027_,
		_w16937_,
		_w16938_,
		_w16939_
	);
	LUT3 #(
		.INIT('h2a)
	) name15039 (
		\m5_addr_i[28]_pad ,
		_w9029_,
		_w9030_,
		_w16940_
	);
	LUT3 #(
		.INIT('h80)
	) name15040 (
		\m6_addr_i[28]_pad ,
		_w9029_,
		_w9030_,
		_w16941_
	);
	LUT4 #(
		.INIT('hcedf)
	) name15041 (
		_w9024_,
		_w9027_,
		_w16940_,
		_w16941_,
		_w16942_
	);
	LUT4 #(
		.INIT('h7fff)
	) name15042 (
		_w16933_,
		_w16936_,
		_w16939_,
		_w16942_,
		_w16943_
	);
	LUT3 #(
		.INIT('h2a)
	) name15043 (
		\m3_addr_i[29]_pad ,
		_w9029_,
		_w9030_,
		_w16944_
	);
	LUT3 #(
		.INIT('h80)
	) name15044 (
		\m4_addr_i[29]_pad ,
		_w9029_,
		_w9030_,
		_w16945_
	);
	LUT4 #(
		.INIT('h9dbf)
	) name15045 (
		_w9024_,
		_w9027_,
		_w16944_,
		_w16945_,
		_w16946_
	);
	LUT3 #(
		.INIT('h2a)
	) name15046 (
		\m5_addr_i[29]_pad ,
		_w9029_,
		_w9030_,
		_w16947_
	);
	LUT3 #(
		.INIT('h80)
	) name15047 (
		\m2_addr_i[29]_pad ,
		_w9029_,
		_w9030_,
		_w16948_
	);
	LUT4 #(
		.INIT('h9bdf)
	) name15048 (
		_w9024_,
		_w9027_,
		_w16947_,
		_w16948_,
		_w16949_
	);
	LUT3 #(
		.INIT('h80)
	) name15049 (
		\m6_addr_i[29]_pad ,
		_w9029_,
		_w9030_,
		_w16950_
	);
	LUT3 #(
		.INIT('h2a)
	) name15050 (
		\m1_addr_i[29]_pad ,
		_w9029_,
		_w9030_,
		_w16951_
	);
	LUT4 #(
		.INIT('h67ef)
	) name15051 (
		_w9024_,
		_w9027_,
		_w16950_,
		_w16951_,
		_w16952_
	);
	LUT3 #(
		.INIT('h80)
	) name15052 (
		\m0_addr_i[29]_pad ,
		_w9029_,
		_w9030_,
		_w16953_
	);
	LUT3 #(
		.INIT('h2a)
	) name15053 (
		\m7_addr_i[29]_pad ,
		_w9029_,
		_w9030_,
		_w16954_
	);
	LUT4 #(
		.INIT('h6e7f)
	) name15054 (
		_w9024_,
		_w9027_,
		_w16953_,
		_w16954_,
		_w16955_
	);
	LUT4 #(
		.INIT('h7fff)
	) name15055 (
		_w16946_,
		_w16949_,
		_w16952_,
		_w16955_,
		_w16956_
	);
	LUT3 #(
		.INIT('h2a)
	) name15056 (
		\m3_addr_i[2]_pad ,
		_w9029_,
		_w9030_,
		_w16957_
	);
	LUT3 #(
		.INIT('h80)
	) name15057 (
		\m4_addr_i[2]_pad ,
		_w9029_,
		_w9030_,
		_w16958_
	);
	LUT4 #(
		.INIT('h9dbf)
	) name15058 (
		_w9024_,
		_w9027_,
		_w16957_,
		_w16958_,
		_w16959_
	);
	LUT3 #(
		.INIT('h80)
	) name15059 (
		\m6_addr_i[2]_pad ,
		_w9029_,
		_w9030_,
		_w16960_
	);
	LUT3 #(
		.INIT('h80)
	) name15060 (
		\m2_addr_i[2]_pad ,
		_w9029_,
		_w9030_,
		_w16961_
	);
	LUT4 #(
		.INIT('habef)
	) name15061 (
		_w9024_,
		_w9027_,
		_w16960_,
		_w16961_,
		_w16962_
	);
	LUT3 #(
		.INIT('h2a)
	) name15062 (
		\m5_addr_i[2]_pad ,
		_w9029_,
		_w9030_,
		_w16963_
	);
	LUT3 #(
		.INIT('h2a)
	) name15063 (
		\m1_addr_i[2]_pad ,
		_w9029_,
		_w9030_,
		_w16964_
	);
	LUT4 #(
		.INIT('h57df)
	) name15064 (
		_w9024_,
		_w9027_,
		_w16963_,
		_w16964_,
		_w16965_
	);
	LUT3 #(
		.INIT('h80)
	) name15065 (
		\m0_addr_i[2]_pad ,
		_w9029_,
		_w9030_,
		_w16966_
	);
	LUT3 #(
		.INIT('h2a)
	) name15066 (
		\m7_addr_i[2]_pad ,
		_w9029_,
		_w9030_,
		_w16967_
	);
	LUT4 #(
		.INIT('h6e7f)
	) name15067 (
		_w9024_,
		_w9027_,
		_w16966_,
		_w16967_,
		_w16968_
	);
	LUT4 #(
		.INIT('h7fff)
	) name15068 (
		_w16959_,
		_w16962_,
		_w16965_,
		_w16968_,
		_w16969_
	);
	LUT3 #(
		.INIT('h2a)
	) name15069 (
		\m1_addr_i[30]_pad ,
		_w9029_,
		_w9030_,
		_w16970_
	);
	LUT3 #(
		.INIT('h80)
	) name15070 (
		\m2_addr_i[30]_pad ,
		_w9029_,
		_w9030_,
		_w16971_
	);
	LUT4 #(
		.INIT('h3b7f)
	) name15071 (
		_w9024_,
		_w9027_,
		_w16970_,
		_w16971_,
		_w16972_
	);
	LUT3 #(
		.INIT('h2a)
	) name15072 (
		\m5_addr_i[30]_pad ,
		_w9029_,
		_w9030_,
		_w16973_
	);
	LUT3 #(
		.INIT('h80)
	) name15073 (
		\m4_addr_i[30]_pad ,
		_w9029_,
		_w9030_,
		_w16974_
	);
	LUT3 #(
		.INIT('h57)
	) name15074 (
		_w9042_,
		_w16973_,
		_w16974_,
		_w16975_
	);
	LUT3 #(
		.INIT('h80)
	) name15075 (
		\m6_addr_i[30]_pad ,
		_w9029_,
		_w9030_,
		_w16976_
	);
	LUT3 #(
		.INIT('h2a)
	) name15076 (
		\m3_addr_i[30]_pad ,
		_w9029_,
		_w9030_,
		_w16977_
	);
	LUT4 #(
		.INIT('habef)
	) name15077 (
		_w9024_,
		_w9027_,
		_w16976_,
		_w16977_,
		_w16978_
	);
	LUT3 #(
		.INIT('h80)
	) name15078 (
		\m0_addr_i[30]_pad ,
		_w9029_,
		_w9030_,
		_w16979_
	);
	LUT3 #(
		.INIT('h2a)
	) name15079 (
		\m7_addr_i[30]_pad ,
		_w9029_,
		_w9030_,
		_w16980_
	);
	LUT4 #(
		.INIT('h6e7f)
	) name15080 (
		_w9024_,
		_w9027_,
		_w16979_,
		_w16980_,
		_w16981_
	);
	LUT4 #(
		.INIT('h7fff)
	) name15081 (
		_w16972_,
		_w16975_,
		_w16978_,
		_w16981_,
		_w16982_
	);
	LUT3 #(
		.INIT('h80)
	) name15082 (
		\m0_addr_i[31]_pad ,
		_w9029_,
		_w9030_,
		_w16983_
	);
	LUT3 #(
		.INIT('h2a)
	) name15083 (
		\m7_addr_i[31]_pad ,
		_w9029_,
		_w9030_,
		_w16984_
	);
	LUT4 #(
		.INIT('h6e7f)
	) name15084 (
		_w9024_,
		_w9027_,
		_w16983_,
		_w16984_,
		_w16985_
	);
	LUT3 #(
		.INIT('h2a)
	) name15085 (
		\m1_addr_i[31]_pad ,
		_w9029_,
		_w9030_,
		_w16986_
	);
	LUT3 #(
		.INIT('h80)
	) name15086 (
		\m6_addr_i[31]_pad ,
		_w9029_,
		_w9030_,
		_w16987_
	);
	LUT4 #(
		.INIT('h6e7f)
	) name15087 (
		_w9024_,
		_w9027_,
		_w16986_,
		_w16987_,
		_w16988_
	);
	LUT3 #(
		.INIT('h80)
	) name15088 (
		\m2_addr_i[31]_pad ,
		_w9029_,
		_w9030_,
		_w16989_
	);
	LUT3 #(
		.INIT('h2a)
	) name15089 (
		\m5_addr_i[31]_pad ,
		_w9029_,
		_w9030_,
		_w16990_
	);
	LUT4 #(
		.INIT('h9dbf)
	) name15090 (
		_w9024_,
		_w9027_,
		_w16989_,
		_w16990_,
		_w16991_
	);
	LUT3 #(
		.INIT('h2a)
	) name15091 (
		\m3_addr_i[31]_pad ,
		_w9029_,
		_w9030_,
		_w16992_
	);
	LUT3 #(
		.INIT('h80)
	) name15092 (
		\m4_addr_i[31]_pad ,
		_w9029_,
		_w9030_,
		_w16993_
	);
	LUT4 #(
		.INIT('h9dbf)
	) name15093 (
		_w9024_,
		_w9027_,
		_w16992_,
		_w16993_,
		_w16994_
	);
	LUT4 #(
		.INIT('h7fff)
	) name15094 (
		_w16985_,
		_w16988_,
		_w16991_,
		_w16994_,
		_w16995_
	);
	LUT3 #(
		.INIT('h2a)
	) name15095 (
		\m3_addr_i[3]_pad ,
		_w9029_,
		_w9030_,
		_w16996_
	);
	LUT3 #(
		.INIT('h80)
	) name15096 (
		\m4_addr_i[3]_pad ,
		_w9029_,
		_w9030_,
		_w16997_
	);
	LUT4 #(
		.INIT('h9dbf)
	) name15097 (
		_w9024_,
		_w9027_,
		_w16996_,
		_w16997_,
		_w16998_
	);
	LUT3 #(
		.INIT('h80)
	) name15098 (
		\m6_addr_i[3]_pad ,
		_w9029_,
		_w9030_,
		_w16999_
	);
	LUT3 #(
		.INIT('h80)
	) name15099 (
		\m2_addr_i[3]_pad ,
		_w9029_,
		_w9030_,
		_w17000_
	);
	LUT4 #(
		.INIT('habef)
	) name15100 (
		_w9024_,
		_w9027_,
		_w16999_,
		_w17000_,
		_w17001_
	);
	LUT3 #(
		.INIT('h2a)
	) name15101 (
		\m5_addr_i[3]_pad ,
		_w9029_,
		_w9030_,
		_w17002_
	);
	LUT3 #(
		.INIT('h2a)
	) name15102 (
		\m1_addr_i[3]_pad ,
		_w9029_,
		_w9030_,
		_w17003_
	);
	LUT4 #(
		.INIT('h57df)
	) name15103 (
		_w9024_,
		_w9027_,
		_w17002_,
		_w17003_,
		_w17004_
	);
	LUT3 #(
		.INIT('h80)
	) name15104 (
		\m0_addr_i[3]_pad ,
		_w9029_,
		_w9030_,
		_w17005_
	);
	LUT3 #(
		.INIT('h2a)
	) name15105 (
		\m7_addr_i[3]_pad ,
		_w9029_,
		_w9030_,
		_w17006_
	);
	LUT4 #(
		.INIT('h6e7f)
	) name15106 (
		_w9024_,
		_w9027_,
		_w17005_,
		_w17006_,
		_w17007_
	);
	LUT4 #(
		.INIT('h7fff)
	) name15107 (
		_w16998_,
		_w17001_,
		_w17004_,
		_w17007_,
		_w17008_
	);
	LUT3 #(
		.INIT('h2a)
	) name15108 (
		\m3_addr_i[4]_pad ,
		_w9029_,
		_w9030_,
		_w17009_
	);
	LUT3 #(
		.INIT('h80)
	) name15109 (
		\m4_addr_i[4]_pad ,
		_w9029_,
		_w9030_,
		_w17010_
	);
	LUT4 #(
		.INIT('h9dbf)
	) name15110 (
		_w9024_,
		_w9027_,
		_w17009_,
		_w17010_,
		_w17011_
	);
	LUT3 #(
		.INIT('h80)
	) name15111 (
		\m6_addr_i[4]_pad ,
		_w9029_,
		_w9030_,
		_w17012_
	);
	LUT3 #(
		.INIT('h80)
	) name15112 (
		\m2_addr_i[4]_pad ,
		_w9029_,
		_w9030_,
		_w17013_
	);
	LUT4 #(
		.INIT('habef)
	) name15113 (
		_w9024_,
		_w9027_,
		_w17012_,
		_w17013_,
		_w17014_
	);
	LUT3 #(
		.INIT('h2a)
	) name15114 (
		\m5_addr_i[4]_pad ,
		_w9029_,
		_w9030_,
		_w17015_
	);
	LUT3 #(
		.INIT('h2a)
	) name15115 (
		\m1_addr_i[4]_pad ,
		_w9029_,
		_w9030_,
		_w17016_
	);
	LUT4 #(
		.INIT('h57df)
	) name15116 (
		_w9024_,
		_w9027_,
		_w17015_,
		_w17016_,
		_w17017_
	);
	LUT3 #(
		.INIT('h80)
	) name15117 (
		\m0_addr_i[4]_pad ,
		_w9029_,
		_w9030_,
		_w17018_
	);
	LUT3 #(
		.INIT('h2a)
	) name15118 (
		\m7_addr_i[4]_pad ,
		_w9029_,
		_w9030_,
		_w17019_
	);
	LUT4 #(
		.INIT('h6e7f)
	) name15119 (
		_w9024_,
		_w9027_,
		_w17018_,
		_w17019_,
		_w17020_
	);
	LUT4 #(
		.INIT('h7fff)
	) name15120 (
		_w17011_,
		_w17014_,
		_w17017_,
		_w17020_,
		_w17021_
	);
	LUT3 #(
		.INIT('h2a)
	) name15121 (
		\m3_addr_i[5]_pad ,
		_w9029_,
		_w9030_,
		_w17022_
	);
	LUT3 #(
		.INIT('h80)
	) name15122 (
		\m4_addr_i[5]_pad ,
		_w9029_,
		_w9030_,
		_w17023_
	);
	LUT4 #(
		.INIT('h9dbf)
	) name15123 (
		_w9024_,
		_w9027_,
		_w17022_,
		_w17023_,
		_w17024_
	);
	LUT3 #(
		.INIT('h80)
	) name15124 (
		\m6_addr_i[5]_pad ,
		_w9029_,
		_w9030_,
		_w17025_
	);
	LUT3 #(
		.INIT('h80)
	) name15125 (
		\m2_addr_i[5]_pad ,
		_w9029_,
		_w9030_,
		_w17026_
	);
	LUT4 #(
		.INIT('habef)
	) name15126 (
		_w9024_,
		_w9027_,
		_w17025_,
		_w17026_,
		_w17027_
	);
	LUT3 #(
		.INIT('h2a)
	) name15127 (
		\m5_addr_i[5]_pad ,
		_w9029_,
		_w9030_,
		_w17028_
	);
	LUT3 #(
		.INIT('h2a)
	) name15128 (
		\m1_addr_i[5]_pad ,
		_w9029_,
		_w9030_,
		_w17029_
	);
	LUT4 #(
		.INIT('h57df)
	) name15129 (
		_w9024_,
		_w9027_,
		_w17028_,
		_w17029_,
		_w17030_
	);
	LUT3 #(
		.INIT('h80)
	) name15130 (
		\m0_addr_i[5]_pad ,
		_w9029_,
		_w9030_,
		_w17031_
	);
	LUT3 #(
		.INIT('h2a)
	) name15131 (
		\m7_addr_i[5]_pad ,
		_w9029_,
		_w9030_,
		_w17032_
	);
	LUT4 #(
		.INIT('h6e7f)
	) name15132 (
		_w9024_,
		_w9027_,
		_w17031_,
		_w17032_,
		_w17033_
	);
	LUT4 #(
		.INIT('h7fff)
	) name15133 (
		_w17024_,
		_w17027_,
		_w17030_,
		_w17033_,
		_w17034_
	);
	LUT3 #(
		.INIT('h2a)
	) name15134 (
		\m3_addr_i[6]_pad ,
		_w9029_,
		_w9030_,
		_w17035_
	);
	LUT3 #(
		.INIT('h80)
	) name15135 (
		\m4_addr_i[6]_pad ,
		_w9029_,
		_w9030_,
		_w17036_
	);
	LUT4 #(
		.INIT('h9dbf)
	) name15136 (
		_w9024_,
		_w9027_,
		_w17035_,
		_w17036_,
		_w17037_
	);
	LUT3 #(
		.INIT('h80)
	) name15137 (
		\m6_addr_i[6]_pad ,
		_w9029_,
		_w9030_,
		_w17038_
	);
	LUT3 #(
		.INIT('h80)
	) name15138 (
		\m2_addr_i[6]_pad ,
		_w9029_,
		_w9030_,
		_w17039_
	);
	LUT4 #(
		.INIT('habef)
	) name15139 (
		_w9024_,
		_w9027_,
		_w17038_,
		_w17039_,
		_w17040_
	);
	LUT3 #(
		.INIT('h2a)
	) name15140 (
		\m5_addr_i[6]_pad ,
		_w9029_,
		_w9030_,
		_w17041_
	);
	LUT3 #(
		.INIT('h2a)
	) name15141 (
		\m1_addr_i[6]_pad ,
		_w9029_,
		_w9030_,
		_w17042_
	);
	LUT4 #(
		.INIT('h57df)
	) name15142 (
		_w9024_,
		_w9027_,
		_w17041_,
		_w17042_,
		_w17043_
	);
	LUT3 #(
		.INIT('h80)
	) name15143 (
		\m0_addr_i[6]_pad ,
		_w9029_,
		_w9030_,
		_w17044_
	);
	LUT3 #(
		.INIT('h2a)
	) name15144 (
		\m7_addr_i[6]_pad ,
		_w9029_,
		_w9030_,
		_w17045_
	);
	LUT4 #(
		.INIT('h6e7f)
	) name15145 (
		_w9024_,
		_w9027_,
		_w17044_,
		_w17045_,
		_w17046_
	);
	LUT4 #(
		.INIT('h7fff)
	) name15146 (
		_w17037_,
		_w17040_,
		_w17043_,
		_w17046_,
		_w17047_
	);
	LUT3 #(
		.INIT('h2a)
	) name15147 (
		\m1_addr_i[7]_pad ,
		_w9029_,
		_w9030_,
		_w17048_
	);
	LUT3 #(
		.INIT('h80)
	) name15148 (
		\m2_addr_i[7]_pad ,
		_w9029_,
		_w9030_,
		_w17049_
	);
	LUT4 #(
		.INIT('h3b7f)
	) name15149 (
		_w9024_,
		_w9027_,
		_w17048_,
		_w17049_,
		_w17050_
	);
	LUT3 #(
		.INIT('h80)
	) name15150 (
		\m6_addr_i[7]_pad ,
		_w9029_,
		_w9030_,
		_w17051_
	);
	LUT3 #(
		.INIT('h80)
	) name15151 (
		\m4_addr_i[7]_pad ,
		_w9029_,
		_w9030_,
		_w17052_
	);
	LUT4 #(
		.INIT('hcdef)
	) name15152 (
		_w9024_,
		_w9027_,
		_w17051_,
		_w17052_,
		_w17053_
	);
	LUT3 #(
		.INIT('h2a)
	) name15153 (
		\m5_addr_i[7]_pad ,
		_w9029_,
		_w9030_,
		_w17054_
	);
	LUT3 #(
		.INIT('h2a)
	) name15154 (
		\m3_addr_i[7]_pad ,
		_w9029_,
		_w9030_,
		_w17055_
	);
	LUT4 #(
		.INIT('h9bdf)
	) name15155 (
		_w9024_,
		_w9027_,
		_w17054_,
		_w17055_,
		_w17056_
	);
	LUT3 #(
		.INIT('h80)
	) name15156 (
		\m0_addr_i[7]_pad ,
		_w9029_,
		_w9030_,
		_w17057_
	);
	LUT3 #(
		.INIT('h2a)
	) name15157 (
		\m7_addr_i[7]_pad ,
		_w9029_,
		_w9030_,
		_w17058_
	);
	LUT4 #(
		.INIT('h6e7f)
	) name15158 (
		_w9024_,
		_w9027_,
		_w17057_,
		_w17058_,
		_w17059_
	);
	LUT4 #(
		.INIT('h7fff)
	) name15159 (
		_w17050_,
		_w17053_,
		_w17056_,
		_w17059_,
		_w17060_
	);
	LUT3 #(
		.INIT('h80)
	) name15160 (
		\m0_addr_i[8]_pad ,
		_w9029_,
		_w9030_,
		_w17061_
	);
	LUT3 #(
		.INIT('h2a)
	) name15161 (
		\m7_addr_i[8]_pad ,
		_w9029_,
		_w9030_,
		_w17062_
	);
	LUT4 #(
		.INIT('h6e7f)
	) name15162 (
		_w9024_,
		_w9027_,
		_w17061_,
		_w17062_,
		_w17063_
	);
	LUT3 #(
		.INIT('h80)
	) name15163 (
		\m6_addr_i[8]_pad ,
		_w9029_,
		_w9030_,
		_w17064_
	);
	LUT3 #(
		.INIT('h80)
	) name15164 (
		\m2_addr_i[8]_pad ,
		_w9029_,
		_w9030_,
		_w17065_
	);
	LUT4 #(
		.INIT('habef)
	) name15165 (
		_w9024_,
		_w9027_,
		_w17064_,
		_w17065_,
		_w17066_
	);
	LUT3 #(
		.INIT('h2a)
	) name15166 (
		\m5_addr_i[8]_pad ,
		_w9029_,
		_w9030_,
		_w17067_
	);
	LUT3 #(
		.INIT('h2a)
	) name15167 (
		\m1_addr_i[8]_pad ,
		_w9029_,
		_w9030_,
		_w17068_
	);
	LUT4 #(
		.INIT('h57df)
	) name15168 (
		_w9024_,
		_w9027_,
		_w17067_,
		_w17068_,
		_w17069_
	);
	LUT3 #(
		.INIT('h2a)
	) name15169 (
		\m3_addr_i[8]_pad ,
		_w9029_,
		_w9030_,
		_w17070_
	);
	LUT3 #(
		.INIT('h80)
	) name15170 (
		\m4_addr_i[8]_pad ,
		_w9029_,
		_w9030_,
		_w17071_
	);
	LUT4 #(
		.INIT('h9dbf)
	) name15171 (
		_w9024_,
		_w9027_,
		_w17070_,
		_w17071_,
		_w17072_
	);
	LUT4 #(
		.INIT('h7fff)
	) name15172 (
		_w17063_,
		_w17066_,
		_w17069_,
		_w17072_,
		_w17073_
	);
	LUT3 #(
		.INIT('h80)
	) name15173 (
		\m6_addr_i[9]_pad ,
		_w9029_,
		_w9030_,
		_w17074_
	);
	LUT3 #(
		.INIT('h2a)
	) name15174 (
		\m5_addr_i[9]_pad ,
		_w9029_,
		_w9030_,
		_w17075_
	);
	LUT4 #(
		.INIT('hcdef)
	) name15175 (
		_w9024_,
		_w9027_,
		_w17074_,
		_w17075_,
		_w17076_
	);
	LUT3 #(
		.INIT('h80)
	) name15176 (
		\m0_addr_i[9]_pad ,
		_w9029_,
		_w9030_,
		_w17077_
	);
	LUT3 #(
		.INIT('h80)
	) name15177 (
		\m4_addr_i[9]_pad ,
		_w9029_,
		_w9030_,
		_w17078_
	);
	LUT4 #(
		.INIT('h5d7f)
	) name15178 (
		_w9024_,
		_w9027_,
		_w17077_,
		_w17078_,
		_w17079_
	);
	LUT3 #(
		.INIT('h2a)
	) name15179 (
		\m7_addr_i[9]_pad ,
		_w9029_,
		_w9030_,
		_w17080_
	);
	LUT3 #(
		.INIT('h2a)
	) name15180 (
		\m3_addr_i[9]_pad ,
		_w9029_,
		_w9030_,
		_w17081_
	);
	LUT4 #(
		.INIT('habef)
	) name15181 (
		_w9024_,
		_w9027_,
		_w17080_,
		_w17081_,
		_w17082_
	);
	LUT3 #(
		.INIT('h2a)
	) name15182 (
		\m1_addr_i[9]_pad ,
		_w9029_,
		_w9030_,
		_w17083_
	);
	LUT3 #(
		.INIT('h80)
	) name15183 (
		\m2_addr_i[9]_pad ,
		_w9029_,
		_w9030_,
		_w17084_
	);
	LUT4 #(
		.INIT('h3b7f)
	) name15184 (
		_w9024_,
		_w9027_,
		_w17083_,
		_w17084_,
		_w17085_
	);
	LUT4 #(
		.INIT('h7fff)
	) name15185 (
		_w17076_,
		_w17079_,
		_w17082_,
		_w17085_,
		_w17086_
	);
	LUT3 #(
		.INIT('h2a)
	) name15186 (
		\m1_data_i[0]_pad ,
		_w9029_,
		_w9030_,
		_w17087_
	);
	LUT3 #(
		.INIT('h80)
	) name15187 (
		\m2_data_i[0]_pad ,
		_w9029_,
		_w9030_,
		_w17088_
	);
	LUT4 #(
		.INIT('h3b7f)
	) name15188 (
		_w9024_,
		_w9027_,
		_w17087_,
		_w17088_,
		_w17089_
	);
	LUT3 #(
		.INIT('h80)
	) name15189 (
		\m0_data_i[0]_pad ,
		_w9029_,
		_w9030_,
		_w17090_
	);
	LUT3 #(
		.INIT('h2a)
	) name15190 (
		\m5_data_i[0]_pad ,
		_w9029_,
		_w9030_,
		_w17091_
	);
	LUT4 #(
		.INIT('h5d7f)
	) name15191 (
		_w9024_,
		_w9027_,
		_w17090_,
		_w17091_,
		_w17092_
	);
	LUT3 #(
		.INIT('h2a)
	) name15192 (
		\m7_data_i[0]_pad ,
		_w9029_,
		_w9030_,
		_w17093_
	);
	LUT3 #(
		.INIT('h80)
	) name15193 (
		\m6_data_i[0]_pad ,
		_w9029_,
		_w9030_,
		_w17094_
	);
	LUT3 #(
		.INIT('h57)
	) name15194 (
		_w9036_,
		_w17093_,
		_w17094_,
		_w17095_
	);
	LUT3 #(
		.INIT('h2a)
	) name15195 (
		\m3_data_i[0]_pad ,
		_w9029_,
		_w9030_,
		_w17096_
	);
	LUT3 #(
		.INIT('h80)
	) name15196 (
		\m4_data_i[0]_pad ,
		_w9029_,
		_w9030_,
		_w17097_
	);
	LUT4 #(
		.INIT('h9dbf)
	) name15197 (
		_w9024_,
		_w9027_,
		_w17096_,
		_w17097_,
		_w17098_
	);
	LUT4 #(
		.INIT('h7fff)
	) name15198 (
		_w17089_,
		_w17092_,
		_w17095_,
		_w17098_,
		_w17099_
	);
	LUT3 #(
		.INIT('h80)
	) name15199 (
		\m0_data_i[10]_pad ,
		_w9029_,
		_w9030_,
		_w17100_
	);
	LUT3 #(
		.INIT('h2a)
	) name15200 (
		\m7_data_i[10]_pad ,
		_w9029_,
		_w9030_,
		_w17101_
	);
	LUT4 #(
		.INIT('h6e7f)
	) name15201 (
		_w9024_,
		_w9027_,
		_w17100_,
		_w17101_,
		_w17102_
	);
	LUT3 #(
		.INIT('h2a)
	) name15202 (
		\m1_data_i[10]_pad ,
		_w9029_,
		_w9030_,
		_w17103_
	);
	LUT3 #(
		.INIT('h80)
	) name15203 (
		\m4_data_i[10]_pad ,
		_w9029_,
		_w9030_,
		_w17104_
	);
	LUT4 #(
		.INIT('h5d7f)
	) name15204 (
		_w9024_,
		_w9027_,
		_w17103_,
		_w17104_,
		_w17105_
	);
	LUT3 #(
		.INIT('h80)
	) name15205 (
		\m2_data_i[10]_pad ,
		_w9029_,
		_w9030_,
		_w17106_
	);
	LUT3 #(
		.INIT('h2a)
	) name15206 (
		\m3_data_i[10]_pad ,
		_w9029_,
		_w9030_,
		_w17107_
	);
	LUT3 #(
		.INIT('h57)
	) name15207 (
		_w9028_,
		_w17106_,
		_w17107_,
		_w17108_
	);
	LUT3 #(
		.INIT('h80)
	) name15208 (
		\m6_data_i[10]_pad ,
		_w9029_,
		_w9030_,
		_w17109_
	);
	LUT3 #(
		.INIT('h2a)
	) name15209 (
		\m5_data_i[10]_pad ,
		_w9029_,
		_w9030_,
		_w17110_
	);
	LUT4 #(
		.INIT('hcdef)
	) name15210 (
		_w9024_,
		_w9027_,
		_w17109_,
		_w17110_,
		_w17111_
	);
	LUT4 #(
		.INIT('h7fff)
	) name15211 (
		_w17102_,
		_w17105_,
		_w17108_,
		_w17111_,
		_w17112_
	);
	LUT3 #(
		.INIT('h2a)
	) name15212 (
		\m1_data_i[11]_pad ,
		_w9029_,
		_w9030_,
		_w17113_
	);
	LUT3 #(
		.INIT('h80)
	) name15213 (
		\m2_data_i[11]_pad ,
		_w9029_,
		_w9030_,
		_w17114_
	);
	LUT4 #(
		.INIT('h3b7f)
	) name15214 (
		_w9024_,
		_w9027_,
		_w17113_,
		_w17114_,
		_w17115_
	);
	LUT3 #(
		.INIT('h80)
	) name15215 (
		\m0_data_i[11]_pad ,
		_w9029_,
		_w9030_,
		_w17116_
	);
	LUT3 #(
		.INIT('h2a)
	) name15216 (
		\m5_data_i[11]_pad ,
		_w9029_,
		_w9030_,
		_w17117_
	);
	LUT4 #(
		.INIT('h5d7f)
	) name15217 (
		_w9024_,
		_w9027_,
		_w17116_,
		_w17117_,
		_w17118_
	);
	LUT3 #(
		.INIT('h2a)
	) name15218 (
		\m7_data_i[11]_pad ,
		_w9029_,
		_w9030_,
		_w17119_
	);
	LUT3 #(
		.INIT('h80)
	) name15219 (
		\m6_data_i[11]_pad ,
		_w9029_,
		_w9030_,
		_w17120_
	);
	LUT3 #(
		.INIT('h57)
	) name15220 (
		_w9036_,
		_w17119_,
		_w17120_,
		_w17121_
	);
	LUT3 #(
		.INIT('h2a)
	) name15221 (
		\m3_data_i[11]_pad ,
		_w9029_,
		_w9030_,
		_w17122_
	);
	LUT3 #(
		.INIT('h80)
	) name15222 (
		\m4_data_i[11]_pad ,
		_w9029_,
		_w9030_,
		_w17123_
	);
	LUT4 #(
		.INIT('h9dbf)
	) name15223 (
		_w9024_,
		_w9027_,
		_w17122_,
		_w17123_,
		_w17124_
	);
	LUT4 #(
		.INIT('h7fff)
	) name15224 (
		_w17115_,
		_w17118_,
		_w17121_,
		_w17124_,
		_w17125_
	);
	LUT3 #(
		.INIT('h80)
	) name15225 (
		\m0_data_i[12]_pad ,
		_w9029_,
		_w9030_,
		_w17126_
	);
	LUT3 #(
		.INIT('h2a)
	) name15226 (
		\m7_data_i[12]_pad ,
		_w9029_,
		_w9030_,
		_w17127_
	);
	LUT4 #(
		.INIT('h6e7f)
	) name15227 (
		_w9024_,
		_w9027_,
		_w17126_,
		_w17127_,
		_w17128_
	);
	LUT3 #(
		.INIT('h2a)
	) name15228 (
		\m1_data_i[12]_pad ,
		_w9029_,
		_w9030_,
		_w17129_
	);
	LUT3 #(
		.INIT('h80)
	) name15229 (
		\m4_data_i[12]_pad ,
		_w9029_,
		_w9030_,
		_w17130_
	);
	LUT4 #(
		.INIT('h5d7f)
	) name15230 (
		_w9024_,
		_w9027_,
		_w17129_,
		_w17130_,
		_w17131_
	);
	LUT3 #(
		.INIT('h80)
	) name15231 (
		\m2_data_i[12]_pad ,
		_w9029_,
		_w9030_,
		_w17132_
	);
	LUT3 #(
		.INIT('h2a)
	) name15232 (
		\m3_data_i[12]_pad ,
		_w9029_,
		_w9030_,
		_w17133_
	);
	LUT3 #(
		.INIT('h57)
	) name15233 (
		_w9028_,
		_w17132_,
		_w17133_,
		_w17134_
	);
	LUT3 #(
		.INIT('h80)
	) name15234 (
		\m6_data_i[12]_pad ,
		_w9029_,
		_w9030_,
		_w17135_
	);
	LUT3 #(
		.INIT('h2a)
	) name15235 (
		\m5_data_i[12]_pad ,
		_w9029_,
		_w9030_,
		_w17136_
	);
	LUT4 #(
		.INIT('hcdef)
	) name15236 (
		_w9024_,
		_w9027_,
		_w17135_,
		_w17136_,
		_w17137_
	);
	LUT4 #(
		.INIT('h7fff)
	) name15237 (
		_w17128_,
		_w17131_,
		_w17134_,
		_w17137_,
		_w17138_
	);
	LUT3 #(
		.INIT('h2a)
	) name15238 (
		\m1_data_i[13]_pad ,
		_w9029_,
		_w9030_,
		_w17139_
	);
	LUT3 #(
		.INIT('h80)
	) name15239 (
		\m2_data_i[13]_pad ,
		_w9029_,
		_w9030_,
		_w17140_
	);
	LUT4 #(
		.INIT('h3b7f)
	) name15240 (
		_w9024_,
		_w9027_,
		_w17139_,
		_w17140_,
		_w17141_
	);
	LUT3 #(
		.INIT('h80)
	) name15241 (
		\m0_data_i[13]_pad ,
		_w9029_,
		_w9030_,
		_w17142_
	);
	LUT3 #(
		.INIT('h80)
	) name15242 (
		\m4_data_i[13]_pad ,
		_w9029_,
		_w9030_,
		_w17143_
	);
	LUT4 #(
		.INIT('h5d7f)
	) name15243 (
		_w9024_,
		_w9027_,
		_w17142_,
		_w17143_,
		_w17144_
	);
	LUT3 #(
		.INIT('h2a)
	) name15244 (
		\m7_data_i[13]_pad ,
		_w9029_,
		_w9030_,
		_w17145_
	);
	LUT3 #(
		.INIT('h2a)
	) name15245 (
		\m3_data_i[13]_pad ,
		_w9029_,
		_w9030_,
		_w17146_
	);
	LUT4 #(
		.INIT('habef)
	) name15246 (
		_w9024_,
		_w9027_,
		_w17145_,
		_w17146_,
		_w17147_
	);
	LUT3 #(
		.INIT('h80)
	) name15247 (
		\m6_data_i[13]_pad ,
		_w9029_,
		_w9030_,
		_w17148_
	);
	LUT3 #(
		.INIT('h2a)
	) name15248 (
		\m5_data_i[13]_pad ,
		_w9029_,
		_w9030_,
		_w17149_
	);
	LUT4 #(
		.INIT('hcdef)
	) name15249 (
		_w9024_,
		_w9027_,
		_w17148_,
		_w17149_,
		_w17150_
	);
	LUT4 #(
		.INIT('h7fff)
	) name15250 (
		_w17141_,
		_w17144_,
		_w17147_,
		_w17150_,
		_w17151_
	);
	LUT3 #(
		.INIT('h2a)
	) name15251 (
		\m3_data_i[14]_pad ,
		_w9029_,
		_w9030_,
		_w17152_
	);
	LUT3 #(
		.INIT('h80)
	) name15252 (
		\m4_data_i[14]_pad ,
		_w9029_,
		_w9030_,
		_w17153_
	);
	LUT4 #(
		.INIT('h9dbf)
	) name15253 (
		_w9024_,
		_w9027_,
		_w17152_,
		_w17153_,
		_w17154_
	);
	LUT3 #(
		.INIT('h80)
	) name15254 (
		\m6_data_i[14]_pad ,
		_w9029_,
		_w9030_,
		_w17155_
	);
	LUT3 #(
		.INIT('h80)
	) name15255 (
		\m2_data_i[14]_pad ,
		_w9029_,
		_w9030_,
		_w17156_
	);
	LUT4 #(
		.INIT('habef)
	) name15256 (
		_w9024_,
		_w9027_,
		_w17155_,
		_w17156_,
		_w17157_
	);
	LUT3 #(
		.INIT('h2a)
	) name15257 (
		\m5_data_i[14]_pad ,
		_w9029_,
		_w9030_,
		_w17158_
	);
	LUT3 #(
		.INIT('h2a)
	) name15258 (
		\m1_data_i[14]_pad ,
		_w9029_,
		_w9030_,
		_w17159_
	);
	LUT4 #(
		.INIT('h57df)
	) name15259 (
		_w9024_,
		_w9027_,
		_w17158_,
		_w17159_,
		_w17160_
	);
	LUT3 #(
		.INIT('h80)
	) name15260 (
		\m0_data_i[14]_pad ,
		_w9029_,
		_w9030_,
		_w17161_
	);
	LUT3 #(
		.INIT('h2a)
	) name15261 (
		\m7_data_i[14]_pad ,
		_w9029_,
		_w9030_,
		_w17162_
	);
	LUT4 #(
		.INIT('h6e7f)
	) name15262 (
		_w9024_,
		_w9027_,
		_w17161_,
		_w17162_,
		_w17163_
	);
	LUT4 #(
		.INIT('h7fff)
	) name15263 (
		_w17154_,
		_w17157_,
		_w17160_,
		_w17163_,
		_w17164_
	);
	LUT3 #(
		.INIT('h80)
	) name15264 (
		\m0_data_i[15]_pad ,
		_w9029_,
		_w9030_,
		_w17165_
	);
	LUT3 #(
		.INIT('h2a)
	) name15265 (
		\m7_data_i[15]_pad ,
		_w9029_,
		_w9030_,
		_w17166_
	);
	LUT4 #(
		.INIT('h6e7f)
	) name15266 (
		_w9024_,
		_w9027_,
		_w17165_,
		_w17166_,
		_w17167_
	);
	LUT3 #(
		.INIT('h80)
	) name15267 (
		\m6_data_i[15]_pad ,
		_w9029_,
		_w9030_,
		_w17168_
	);
	LUT3 #(
		.INIT('h80)
	) name15268 (
		\m4_data_i[15]_pad ,
		_w9029_,
		_w9030_,
		_w17169_
	);
	LUT4 #(
		.INIT('hcdef)
	) name15269 (
		_w9024_,
		_w9027_,
		_w17168_,
		_w17169_,
		_w17170_
	);
	LUT3 #(
		.INIT('h2a)
	) name15270 (
		\m5_data_i[15]_pad ,
		_w9029_,
		_w9030_,
		_w17171_
	);
	LUT3 #(
		.INIT('h2a)
	) name15271 (
		\m3_data_i[15]_pad ,
		_w9029_,
		_w9030_,
		_w17172_
	);
	LUT4 #(
		.INIT('h9bdf)
	) name15272 (
		_w9024_,
		_w9027_,
		_w17171_,
		_w17172_,
		_w17173_
	);
	LUT3 #(
		.INIT('h2a)
	) name15273 (
		\m1_data_i[15]_pad ,
		_w9029_,
		_w9030_,
		_w17174_
	);
	LUT3 #(
		.INIT('h80)
	) name15274 (
		\m2_data_i[15]_pad ,
		_w9029_,
		_w9030_,
		_w17175_
	);
	LUT4 #(
		.INIT('h3b7f)
	) name15275 (
		_w9024_,
		_w9027_,
		_w17174_,
		_w17175_,
		_w17176_
	);
	LUT4 #(
		.INIT('h7fff)
	) name15276 (
		_w17167_,
		_w17170_,
		_w17173_,
		_w17176_,
		_w17177_
	);
	LUT3 #(
		.INIT('h80)
	) name15277 (
		\m6_data_i[16]_pad ,
		_w9029_,
		_w9030_,
		_w17178_
	);
	LUT3 #(
		.INIT('h2a)
	) name15278 (
		\m5_data_i[16]_pad ,
		_w9029_,
		_w9030_,
		_w17179_
	);
	LUT4 #(
		.INIT('hcdef)
	) name15279 (
		_w9024_,
		_w9027_,
		_w17178_,
		_w17179_,
		_w17180_
	);
	LUT3 #(
		.INIT('h2a)
	) name15280 (
		\m3_data_i[16]_pad ,
		_w9029_,
		_w9030_,
		_w17181_
	);
	LUT3 #(
		.INIT('h2a)
	) name15281 (
		\m7_data_i[16]_pad ,
		_w9029_,
		_w9030_,
		_w17182_
	);
	LUT4 #(
		.INIT('haebf)
	) name15282 (
		_w9024_,
		_w9027_,
		_w17181_,
		_w17182_,
		_w17183_
	);
	LUT3 #(
		.INIT('h80)
	) name15283 (
		\m4_data_i[16]_pad ,
		_w9029_,
		_w9030_,
		_w17184_
	);
	LUT3 #(
		.INIT('h80)
	) name15284 (
		\m0_data_i[16]_pad ,
		_w9029_,
		_w9030_,
		_w17185_
	);
	LUT4 #(
		.INIT('h57df)
	) name15285 (
		_w9024_,
		_w9027_,
		_w17184_,
		_w17185_,
		_w17186_
	);
	LUT3 #(
		.INIT('h2a)
	) name15286 (
		\m1_data_i[16]_pad ,
		_w9029_,
		_w9030_,
		_w17187_
	);
	LUT3 #(
		.INIT('h80)
	) name15287 (
		\m2_data_i[16]_pad ,
		_w9029_,
		_w9030_,
		_w17188_
	);
	LUT4 #(
		.INIT('h3b7f)
	) name15288 (
		_w9024_,
		_w9027_,
		_w17187_,
		_w17188_,
		_w17189_
	);
	LUT4 #(
		.INIT('h7fff)
	) name15289 (
		_w17180_,
		_w17183_,
		_w17186_,
		_w17189_,
		_w17190_
	);
	LUT3 #(
		.INIT('h2a)
	) name15290 (
		\m1_data_i[17]_pad ,
		_w9029_,
		_w9030_,
		_w17191_
	);
	LUT3 #(
		.INIT('h80)
	) name15291 (
		\m2_data_i[17]_pad ,
		_w9029_,
		_w9030_,
		_w17192_
	);
	LUT4 #(
		.INIT('h3b7f)
	) name15292 (
		_w9024_,
		_w9027_,
		_w17191_,
		_w17192_,
		_w17193_
	);
	LUT3 #(
		.INIT('h80)
	) name15293 (
		\m0_data_i[17]_pad ,
		_w9029_,
		_w9030_,
		_w17194_
	);
	LUT3 #(
		.INIT('h2a)
	) name15294 (
		\m5_data_i[17]_pad ,
		_w9029_,
		_w9030_,
		_w17195_
	);
	LUT4 #(
		.INIT('h5d7f)
	) name15295 (
		_w9024_,
		_w9027_,
		_w17194_,
		_w17195_,
		_w17196_
	);
	LUT3 #(
		.INIT('h2a)
	) name15296 (
		\m7_data_i[17]_pad ,
		_w9029_,
		_w9030_,
		_w17197_
	);
	LUT3 #(
		.INIT('h80)
	) name15297 (
		\m6_data_i[17]_pad ,
		_w9029_,
		_w9030_,
		_w17198_
	);
	LUT3 #(
		.INIT('h57)
	) name15298 (
		_w9036_,
		_w17197_,
		_w17198_,
		_w17199_
	);
	LUT3 #(
		.INIT('h2a)
	) name15299 (
		\m3_data_i[17]_pad ,
		_w9029_,
		_w9030_,
		_w17200_
	);
	LUT3 #(
		.INIT('h80)
	) name15300 (
		\m4_data_i[17]_pad ,
		_w9029_,
		_w9030_,
		_w17201_
	);
	LUT4 #(
		.INIT('h9dbf)
	) name15301 (
		_w9024_,
		_w9027_,
		_w17200_,
		_w17201_,
		_w17202_
	);
	LUT4 #(
		.INIT('h7fff)
	) name15302 (
		_w17193_,
		_w17196_,
		_w17199_,
		_w17202_,
		_w17203_
	);
	LUT3 #(
		.INIT('h2a)
	) name15303 (
		\m1_data_i[18]_pad ,
		_w9029_,
		_w9030_,
		_w17204_
	);
	LUT3 #(
		.INIT('h80)
	) name15304 (
		\m2_data_i[18]_pad ,
		_w9029_,
		_w9030_,
		_w17205_
	);
	LUT4 #(
		.INIT('h3b7f)
	) name15305 (
		_w9024_,
		_w9027_,
		_w17204_,
		_w17205_,
		_w17206_
	);
	LUT3 #(
		.INIT('h80)
	) name15306 (
		\m0_data_i[18]_pad ,
		_w9029_,
		_w9030_,
		_w17207_
	);
	LUT3 #(
		.INIT('h2a)
	) name15307 (
		\m5_data_i[18]_pad ,
		_w9029_,
		_w9030_,
		_w17208_
	);
	LUT4 #(
		.INIT('h5d7f)
	) name15308 (
		_w9024_,
		_w9027_,
		_w17207_,
		_w17208_,
		_w17209_
	);
	LUT3 #(
		.INIT('h2a)
	) name15309 (
		\m7_data_i[18]_pad ,
		_w9029_,
		_w9030_,
		_w17210_
	);
	LUT3 #(
		.INIT('h80)
	) name15310 (
		\m6_data_i[18]_pad ,
		_w9029_,
		_w9030_,
		_w17211_
	);
	LUT3 #(
		.INIT('h57)
	) name15311 (
		_w9036_,
		_w17210_,
		_w17211_,
		_w17212_
	);
	LUT3 #(
		.INIT('h2a)
	) name15312 (
		\m3_data_i[18]_pad ,
		_w9029_,
		_w9030_,
		_w17213_
	);
	LUT3 #(
		.INIT('h80)
	) name15313 (
		\m4_data_i[18]_pad ,
		_w9029_,
		_w9030_,
		_w17214_
	);
	LUT4 #(
		.INIT('h9dbf)
	) name15314 (
		_w9024_,
		_w9027_,
		_w17213_,
		_w17214_,
		_w17215_
	);
	LUT4 #(
		.INIT('h7fff)
	) name15315 (
		_w17206_,
		_w17209_,
		_w17212_,
		_w17215_,
		_w17216_
	);
	LUT3 #(
		.INIT('h2a)
	) name15316 (
		\m1_data_i[19]_pad ,
		_w9029_,
		_w9030_,
		_w17217_
	);
	LUT3 #(
		.INIT('h80)
	) name15317 (
		\m2_data_i[19]_pad ,
		_w9029_,
		_w9030_,
		_w17218_
	);
	LUT4 #(
		.INIT('h3b7f)
	) name15318 (
		_w9024_,
		_w9027_,
		_w17217_,
		_w17218_,
		_w17219_
	);
	LUT3 #(
		.INIT('h80)
	) name15319 (
		\m0_data_i[19]_pad ,
		_w9029_,
		_w9030_,
		_w17220_
	);
	LUT3 #(
		.INIT('h80)
	) name15320 (
		\m4_data_i[19]_pad ,
		_w9029_,
		_w9030_,
		_w17221_
	);
	LUT4 #(
		.INIT('h5d7f)
	) name15321 (
		_w9024_,
		_w9027_,
		_w17220_,
		_w17221_,
		_w17222_
	);
	LUT3 #(
		.INIT('h2a)
	) name15322 (
		\m7_data_i[19]_pad ,
		_w9029_,
		_w9030_,
		_w17223_
	);
	LUT3 #(
		.INIT('h2a)
	) name15323 (
		\m3_data_i[19]_pad ,
		_w9029_,
		_w9030_,
		_w17224_
	);
	LUT4 #(
		.INIT('habef)
	) name15324 (
		_w9024_,
		_w9027_,
		_w17223_,
		_w17224_,
		_w17225_
	);
	LUT3 #(
		.INIT('h80)
	) name15325 (
		\m6_data_i[19]_pad ,
		_w9029_,
		_w9030_,
		_w17226_
	);
	LUT3 #(
		.INIT('h2a)
	) name15326 (
		\m5_data_i[19]_pad ,
		_w9029_,
		_w9030_,
		_w17227_
	);
	LUT4 #(
		.INIT('hcdef)
	) name15327 (
		_w9024_,
		_w9027_,
		_w17226_,
		_w17227_,
		_w17228_
	);
	LUT4 #(
		.INIT('h7fff)
	) name15328 (
		_w17219_,
		_w17222_,
		_w17225_,
		_w17228_,
		_w17229_
	);
	LUT3 #(
		.INIT('h2a)
	) name15329 (
		\m3_data_i[1]_pad ,
		_w9029_,
		_w9030_,
		_w17230_
	);
	LUT3 #(
		.INIT('h80)
	) name15330 (
		\m4_data_i[1]_pad ,
		_w9029_,
		_w9030_,
		_w17231_
	);
	LUT4 #(
		.INIT('h9dbf)
	) name15331 (
		_w9024_,
		_w9027_,
		_w17230_,
		_w17231_,
		_w17232_
	);
	LUT3 #(
		.INIT('h2a)
	) name15332 (
		\m1_data_i[1]_pad ,
		_w9029_,
		_w9030_,
		_w17233_
	);
	LUT3 #(
		.INIT('h2a)
	) name15333 (
		\m7_data_i[1]_pad ,
		_w9029_,
		_w9030_,
		_w17234_
	);
	LUT4 #(
		.INIT('h6e7f)
	) name15334 (
		_w9024_,
		_w9027_,
		_w17233_,
		_w17234_,
		_w17235_
	);
	LUT3 #(
		.INIT('h80)
	) name15335 (
		\m2_data_i[1]_pad ,
		_w9029_,
		_w9030_,
		_w17236_
	);
	LUT3 #(
		.INIT('h80)
	) name15336 (
		\m0_data_i[1]_pad ,
		_w9029_,
		_w9030_,
		_w17237_
	);
	LUT4 #(
		.INIT('h37bf)
	) name15337 (
		_w9024_,
		_w9027_,
		_w17236_,
		_w17237_,
		_w17238_
	);
	LUT3 #(
		.INIT('h80)
	) name15338 (
		\m6_data_i[1]_pad ,
		_w9029_,
		_w9030_,
		_w17239_
	);
	LUT3 #(
		.INIT('h2a)
	) name15339 (
		\m5_data_i[1]_pad ,
		_w9029_,
		_w9030_,
		_w17240_
	);
	LUT4 #(
		.INIT('hcdef)
	) name15340 (
		_w9024_,
		_w9027_,
		_w17239_,
		_w17240_,
		_w17241_
	);
	LUT4 #(
		.INIT('h7fff)
	) name15341 (
		_w17232_,
		_w17235_,
		_w17238_,
		_w17241_,
		_w17242_
	);
	LUT3 #(
		.INIT('h80)
	) name15342 (
		\m6_data_i[20]_pad ,
		_w9029_,
		_w9030_,
		_w17243_
	);
	LUT3 #(
		.INIT('h2a)
	) name15343 (
		\m5_data_i[20]_pad ,
		_w9029_,
		_w9030_,
		_w17244_
	);
	LUT4 #(
		.INIT('hcdef)
	) name15344 (
		_w9024_,
		_w9027_,
		_w17243_,
		_w17244_,
		_w17245_
	);
	LUT3 #(
		.INIT('h80)
	) name15345 (
		\m0_data_i[20]_pad ,
		_w9029_,
		_w9030_,
		_w17246_
	);
	LUT3 #(
		.INIT('h80)
	) name15346 (
		\m4_data_i[20]_pad ,
		_w9029_,
		_w9030_,
		_w17247_
	);
	LUT4 #(
		.INIT('h5d7f)
	) name15347 (
		_w9024_,
		_w9027_,
		_w17246_,
		_w17247_,
		_w17248_
	);
	LUT3 #(
		.INIT('h2a)
	) name15348 (
		\m7_data_i[20]_pad ,
		_w9029_,
		_w9030_,
		_w17249_
	);
	LUT3 #(
		.INIT('h2a)
	) name15349 (
		\m3_data_i[20]_pad ,
		_w9029_,
		_w9030_,
		_w17250_
	);
	LUT4 #(
		.INIT('habef)
	) name15350 (
		_w9024_,
		_w9027_,
		_w17249_,
		_w17250_,
		_w17251_
	);
	LUT3 #(
		.INIT('h2a)
	) name15351 (
		\m1_data_i[20]_pad ,
		_w9029_,
		_w9030_,
		_w17252_
	);
	LUT3 #(
		.INIT('h80)
	) name15352 (
		\m2_data_i[20]_pad ,
		_w9029_,
		_w9030_,
		_w17253_
	);
	LUT4 #(
		.INIT('h3b7f)
	) name15353 (
		_w9024_,
		_w9027_,
		_w17252_,
		_w17253_,
		_w17254_
	);
	LUT4 #(
		.INIT('h7fff)
	) name15354 (
		_w17245_,
		_w17248_,
		_w17251_,
		_w17254_,
		_w17255_
	);
	LUT3 #(
		.INIT('h2a)
	) name15355 (
		\m3_data_i[21]_pad ,
		_w9029_,
		_w9030_,
		_w17256_
	);
	LUT3 #(
		.INIT('h80)
	) name15356 (
		\m4_data_i[21]_pad ,
		_w9029_,
		_w9030_,
		_w17257_
	);
	LUT4 #(
		.INIT('h9dbf)
	) name15357 (
		_w9024_,
		_w9027_,
		_w17256_,
		_w17257_,
		_w17258_
	);
	LUT3 #(
		.INIT('h2a)
	) name15358 (
		\m1_data_i[21]_pad ,
		_w9029_,
		_w9030_,
		_w17259_
	);
	LUT3 #(
		.INIT('h2a)
	) name15359 (
		\m5_data_i[21]_pad ,
		_w9029_,
		_w9030_,
		_w17260_
	);
	LUT4 #(
		.INIT('h5d7f)
	) name15360 (
		_w9024_,
		_w9027_,
		_w17259_,
		_w17260_,
		_w17261_
	);
	LUT3 #(
		.INIT('h80)
	) name15361 (
		\m2_data_i[21]_pad ,
		_w9029_,
		_w9030_,
		_w17262_
	);
	LUT3 #(
		.INIT('h80)
	) name15362 (
		\m6_data_i[21]_pad ,
		_w9029_,
		_w9030_,
		_w17263_
	);
	LUT4 #(
		.INIT('haebf)
	) name15363 (
		_w9024_,
		_w9027_,
		_w17262_,
		_w17263_,
		_w17264_
	);
	LUT3 #(
		.INIT('h80)
	) name15364 (
		\m0_data_i[21]_pad ,
		_w9029_,
		_w9030_,
		_w17265_
	);
	LUT3 #(
		.INIT('h2a)
	) name15365 (
		\m7_data_i[21]_pad ,
		_w9029_,
		_w9030_,
		_w17266_
	);
	LUT4 #(
		.INIT('h6e7f)
	) name15366 (
		_w9024_,
		_w9027_,
		_w17265_,
		_w17266_,
		_w17267_
	);
	LUT4 #(
		.INIT('h7fff)
	) name15367 (
		_w17258_,
		_w17261_,
		_w17264_,
		_w17267_,
		_w17268_
	);
	LUT3 #(
		.INIT('h80)
	) name15368 (
		\m6_data_i[22]_pad ,
		_w9029_,
		_w9030_,
		_w17269_
	);
	LUT3 #(
		.INIT('h2a)
	) name15369 (
		\m5_data_i[22]_pad ,
		_w9029_,
		_w9030_,
		_w17270_
	);
	LUT4 #(
		.INIT('hcdef)
	) name15370 (
		_w9024_,
		_w9027_,
		_w17269_,
		_w17270_,
		_w17271_
	);
	LUT3 #(
		.INIT('h2a)
	) name15371 (
		\m3_data_i[22]_pad ,
		_w9029_,
		_w9030_,
		_w17272_
	);
	LUT3 #(
		.INIT('h80)
	) name15372 (
		\m2_data_i[22]_pad ,
		_w9029_,
		_w9030_,
		_w17273_
	);
	LUT3 #(
		.INIT('h57)
	) name15373 (
		_w9028_,
		_w17272_,
		_w17273_,
		_w17274_
	);
	LUT3 #(
		.INIT('h80)
	) name15374 (
		\m4_data_i[22]_pad ,
		_w9029_,
		_w9030_,
		_w17275_
	);
	LUT3 #(
		.INIT('h2a)
	) name15375 (
		\m1_data_i[22]_pad ,
		_w9029_,
		_w9030_,
		_w17276_
	);
	LUT4 #(
		.INIT('h57df)
	) name15376 (
		_w9024_,
		_w9027_,
		_w17275_,
		_w17276_,
		_w17277_
	);
	LUT3 #(
		.INIT('h80)
	) name15377 (
		\m0_data_i[22]_pad ,
		_w9029_,
		_w9030_,
		_w17278_
	);
	LUT3 #(
		.INIT('h2a)
	) name15378 (
		\m7_data_i[22]_pad ,
		_w9029_,
		_w9030_,
		_w17279_
	);
	LUT4 #(
		.INIT('h6e7f)
	) name15379 (
		_w9024_,
		_w9027_,
		_w17278_,
		_w17279_,
		_w17280_
	);
	LUT4 #(
		.INIT('h7fff)
	) name15380 (
		_w17271_,
		_w17274_,
		_w17277_,
		_w17280_,
		_w17281_
	);
	LUT3 #(
		.INIT('h80)
	) name15381 (
		\m6_data_i[23]_pad ,
		_w9029_,
		_w9030_,
		_w17282_
	);
	LUT3 #(
		.INIT('h2a)
	) name15382 (
		\m5_data_i[23]_pad ,
		_w9029_,
		_w9030_,
		_w17283_
	);
	LUT4 #(
		.INIT('hcdef)
	) name15383 (
		_w9024_,
		_w9027_,
		_w17282_,
		_w17283_,
		_w17284_
	);
	LUT3 #(
		.INIT('h80)
	) name15384 (
		\m0_data_i[23]_pad ,
		_w9029_,
		_w9030_,
		_w17285_
	);
	LUT3 #(
		.INIT('h80)
	) name15385 (
		\m2_data_i[23]_pad ,
		_w9029_,
		_w9030_,
		_w17286_
	);
	LUT4 #(
		.INIT('h3b7f)
	) name15386 (
		_w9024_,
		_w9027_,
		_w17285_,
		_w17286_,
		_w17287_
	);
	LUT3 #(
		.INIT('h2a)
	) name15387 (
		\m7_data_i[23]_pad ,
		_w9029_,
		_w9030_,
		_w17288_
	);
	LUT3 #(
		.INIT('h2a)
	) name15388 (
		\m1_data_i[23]_pad ,
		_w9029_,
		_w9030_,
		_w17289_
	);
	LUT4 #(
		.INIT('h67ef)
	) name15389 (
		_w9024_,
		_w9027_,
		_w17288_,
		_w17289_,
		_w17290_
	);
	LUT3 #(
		.INIT('h2a)
	) name15390 (
		\m3_data_i[23]_pad ,
		_w9029_,
		_w9030_,
		_w17291_
	);
	LUT3 #(
		.INIT('h80)
	) name15391 (
		\m4_data_i[23]_pad ,
		_w9029_,
		_w9030_,
		_w17292_
	);
	LUT4 #(
		.INIT('h9dbf)
	) name15392 (
		_w9024_,
		_w9027_,
		_w17291_,
		_w17292_,
		_w17293_
	);
	LUT4 #(
		.INIT('h7fff)
	) name15393 (
		_w17284_,
		_w17287_,
		_w17290_,
		_w17293_,
		_w17294_
	);
	LUT3 #(
		.INIT('h80)
	) name15394 (
		\m6_data_i[24]_pad ,
		_w9029_,
		_w9030_,
		_w17295_
	);
	LUT3 #(
		.INIT('h2a)
	) name15395 (
		\m5_data_i[24]_pad ,
		_w9029_,
		_w9030_,
		_w17296_
	);
	LUT4 #(
		.INIT('hcdef)
	) name15396 (
		_w9024_,
		_w9027_,
		_w17295_,
		_w17296_,
		_w17297_
	);
	LUT3 #(
		.INIT('h2a)
	) name15397 (
		\m1_data_i[24]_pad ,
		_w9029_,
		_w9030_,
		_w17298_
	);
	LUT3 #(
		.INIT('h2a)
	) name15398 (
		\m7_data_i[24]_pad ,
		_w9029_,
		_w9030_,
		_w17299_
	);
	LUT4 #(
		.INIT('h6e7f)
	) name15399 (
		_w9024_,
		_w9027_,
		_w17298_,
		_w17299_,
		_w17300_
	);
	LUT3 #(
		.INIT('h80)
	) name15400 (
		\m2_data_i[24]_pad ,
		_w9029_,
		_w9030_,
		_w17301_
	);
	LUT3 #(
		.INIT('h80)
	) name15401 (
		\m0_data_i[24]_pad ,
		_w9029_,
		_w9030_,
		_w17302_
	);
	LUT4 #(
		.INIT('h37bf)
	) name15402 (
		_w9024_,
		_w9027_,
		_w17301_,
		_w17302_,
		_w17303_
	);
	LUT3 #(
		.INIT('h2a)
	) name15403 (
		\m3_data_i[24]_pad ,
		_w9029_,
		_w9030_,
		_w17304_
	);
	LUT3 #(
		.INIT('h80)
	) name15404 (
		\m4_data_i[24]_pad ,
		_w9029_,
		_w9030_,
		_w17305_
	);
	LUT4 #(
		.INIT('h9dbf)
	) name15405 (
		_w9024_,
		_w9027_,
		_w17304_,
		_w17305_,
		_w17306_
	);
	LUT4 #(
		.INIT('h7fff)
	) name15406 (
		_w17297_,
		_w17300_,
		_w17303_,
		_w17306_,
		_w17307_
	);
	LUT3 #(
		.INIT('h2a)
	) name15407 (
		\m3_data_i[25]_pad ,
		_w9029_,
		_w9030_,
		_w17308_
	);
	LUT3 #(
		.INIT('h80)
	) name15408 (
		\m4_data_i[25]_pad ,
		_w9029_,
		_w9030_,
		_w17309_
	);
	LUT4 #(
		.INIT('h9dbf)
	) name15409 (
		_w9024_,
		_w9027_,
		_w17308_,
		_w17309_,
		_w17310_
	);
	LUT3 #(
		.INIT('h80)
	) name15410 (
		\m0_data_i[25]_pad ,
		_w9029_,
		_w9030_,
		_w17311_
	);
	LUT3 #(
		.INIT('h80)
	) name15411 (
		\m2_data_i[25]_pad ,
		_w9029_,
		_w9030_,
		_w17312_
	);
	LUT4 #(
		.INIT('h3b7f)
	) name15412 (
		_w9024_,
		_w9027_,
		_w17311_,
		_w17312_,
		_w17313_
	);
	LUT3 #(
		.INIT('h2a)
	) name15413 (
		\m7_data_i[25]_pad ,
		_w9029_,
		_w9030_,
		_w17314_
	);
	LUT3 #(
		.INIT('h2a)
	) name15414 (
		\m1_data_i[25]_pad ,
		_w9029_,
		_w9030_,
		_w17315_
	);
	LUT4 #(
		.INIT('h67ef)
	) name15415 (
		_w9024_,
		_w9027_,
		_w17314_,
		_w17315_,
		_w17316_
	);
	LUT3 #(
		.INIT('h80)
	) name15416 (
		\m6_data_i[25]_pad ,
		_w9029_,
		_w9030_,
		_w17317_
	);
	LUT3 #(
		.INIT('h2a)
	) name15417 (
		\m5_data_i[25]_pad ,
		_w9029_,
		_w9030_,
		_w17318_
	);
	LUT4 #(
		.INIT('hcdef)
	) name15418 (
		_w9024_,
		_w9027_,
		_w17317_,
		_w17318_,
		_w17319_
	);
	LUT4 #(
		.INIT('h7fff)
	) name15419 (
		_w17310_,
		_w17313_,
		_w17316_,
		_w17319_,
		_w17320_
	);
	LUT3 #(
		.INIT('h2a)
	) name15420 (
		\m1_data_i[26]_pad ,
		_w9029_,
		_w9030_,
		_w17321_
	);
	LUT3 #(
		.INIT('h80)
	) name15421 (
		\m2_data_i[26]_pad ,
		_w9029_,
		_w9030_,
		_w17322_
	);
	LUT4 #(
		.INIT('h3b7f)
	) name15422 (
		_w9024_,
		_w9027_,
		_w17321_,
		_w17322_,
		_w17323_
	);
	LUT3 #(
		.INIT('h80)
	) name15423 (
		\m0_data_i[26]_pad ,
		_w9029_,
		_w9030_,
		_w17324_
	);
	LUT3 #(
		.INIT('h2a)
	) name15424 (
		\m5_data_i[26]_pad ,
		_w9029_,
		_w9030_,
		_w17325_
	);
	LUT4 #(
		.INIT('h5d7f)
	) name15425 (
		_w9024_,
		_w9027_,
		_w17324_,
		_w17325_,
		_w17326_
	);
	LUT3 #(
		.INIT('h2a)
	) name15426 (
		\m7_data_i[26]_pad ,
		_w9029_,
		_w9030_,
		_w17327_
	);
	LUT3 #(
		.INIT('h80)
	) name15427 (
		\m6_data_i[26]_pad ,
		_w9029_,
		_w9030_,
		_w17328_
	);
	LUT3 #(
		.INIT('h57)
	) name15428 (
		_w9036_,
		_w17327_,
		_w17328_,
		_w17329_
	);
	LUT3 #(
		.INIT('h2a)
	) name15429 (
		\m3_data_i[26]_pad ,
		_w9029_,
		_w9030_,
		_w17330_
	);
	LUT3 #(
		.INIT('h80)
	) name15430 (
		\m4_data_i[26]_pad ,
		_w9029_,
		_w9030_,
		_w17331_
	);
	LUT4 #(
		.INIT('h9dbf)
	) name15431 (
		_w9024_,
		_w9027_,
		_w17330_,
		_w17331_,
		_w17332_
	);
	LUT4 #(
		.INIT('h7fff)
	) name15432 (
		_w17323_,
		_w17326_,
		_w17329_,
		_w17332_,
		_w17333_
	);
	LUT3 #(
		.INIT('h2a)
	) name15433 (
		\m1_data_i[27]_pad ,
		_w9029_,
		_w9030_,
		_w17334_
	);
	LUT3 #(
		.INIT('h80)
	) name15434 (
		\m2_data_i[27]_pad ,
		_w9029_,
		_w9030_,
		_w17335_
	);
	LUT4 #(
		.INIT('h3b7f)
	) name15435 (
		_w9024_,
		_w9027_,
		_w17334_,
		_w17335_,
		_w17336_
	);
	LUT3 #(
		.INIT('h2a)
	) name15436 (
		\m3_data_i[27]_pad ,
		_w9029_,
		_w9030_,
		_w17337_
	);
	LUT3 #(
		.INIT('h2a)
	) name15437 (
		\m7_data_i[27]_pad ,
		_w9029_,
		_w9030_,
		_w17338_
	);
	LUT4 #(
		.INIT('haebf)
	) name15438 (
		_w9024_,
		_w9027_,
		_w17337_,
		_w17338_,
		_w17339_
	);
	LUT3 #(
		.INIT('h80)
	) name15439 (
		\m4_data_i[27]_pad ,
		_w9029_,
		_w9030_,
		_w17340_
	);
	LUT3 #(
		.INIT('h80)
	) name15440 (
		\m0_data_i[27]_pad ,
		_w9029_,
		_w9030_,
		_w17341_
	);
	LUT4 #(
		.INIT('h57df)
	) name15441 (
		_w9024_,
		_w9027_,
		_w17340_,
		_w17341_,
		_w17342_
	);
	LUT3 #(
		.INIT('h80)
	) name15442 (
		\m6_data_i[27]_pad ,
		_w9029_,
		_w9030_,
		_w17343_
	);
	LUT3 #(
		.INIT('h2a)
	) name15443 (
		\m5_data_i[27]_pad ,
		_w9029_,
		_w9030_,
		_w17344_
	);
	LUT4 #(
		.INIT('hcdef)
	) name15444 (
		_w9024_,
		_w9027_,
		_w17343_,
		_w17344_,
		_w17345_
	);
	LUT4 #(
		.INIT('h7fff)
	) name15445 (
		_w17336_,
		_w17339_,
		_w17342_,
		_w17345_,
		_w17346_
	);
	LUT3 #(
		.INIT('h2a)
	) name15446 (
		\m3_data_i[28]_pad ,
		_w9029_,
		_w9030_,
		_w17347_
	);
	LUT3 #(
		.INIT('h80)
	) name15447 (
		\m4_data_i[28]_pad ,
		_w9029_,
		_w9030_,
		_w17348_
	);
	LUT4 #(
		.INIT('h9dbf)
	) name15448 (
		_w9024_,
		_w9027_,
		_w17347_,
		_w17348_,
		_w17349_
	);
	LUT3 #(
		.INIT('h80)
	) name15449 (
		\m6_data_i[28]_pad ,
		_w9029_,
		_w9030_,
		_w17350_
	);
	LUT3 #(
		.INIT('h80)
	) name15450 (
		\m2_data_i[28]_pad ,
		_w9029_,
		_w9030_,
		_w17351_
	);
	LUT4 #(
		.INIT('habef)
	) name15451 (
		_w9024_,
		_w9027_,
		_w17350_,
		_w17351_,
		_w17352_
	);
	LUT3 #(
		.INIT('h2a)
	) name15452 (
		\m5_data_i[28]_pad ,
		_w9029_,
		_w9030_,
		_w17353_
	);
	LUT3 #(
		.INIT('h2a)
	) name15453 (
		\m1_data_i[28]_pad ,
		_w9029_,
		_w9030_,
		_w17354_
	);
	LUT4 #(
		.INIT('h57df)
	) name15454 (
		_w9024_,
		_w9027_,
		_w17353_,
		_w17354_,
		_w17355_
	);
	LUT3 #(
		.INIT('h80)
	) name15455 (
		\m0_data_i[28]_pad ,
		_w9029_,
		_w9030_,
		_w17356_
	);
	LUT3 #(
		.INIT('h2a)
	) name15456 (
		\m7_data_i[28]_pad ,
		_w9029_,
		_w9030_,
		_w17357_
	);
	LUT4 #(
		.INIT('h6e7f)
	) name15457 (
		_w9024_,
		_w9027_,
		_w17356_,
		_w17357_,
		_w17358_
	);
	LUT4 #(
		.INIT('h7fff)
	) name15458 (
		_w17349_,
		_w17352_,
		_w17355_,
		_w17358_,
		_w17359_
	);
	LUT3 #(
		.INIT('h80)
	) name15459 (
		\m6_data_i[29]_pad ,
		_w9029_,
		_w9030_,
		_w17360_
	);
	LUT3 #(
		.INIT('h2a)
	) name15460 (
		\m5_data_i[29]_pad ,
		_w9029_,
		_w9030_,
		_w17361_
	);
	LUT4 #(
		.INIT('hcdef)
	) name15461 (
		_w9024_,
		_w9027_,
		_w17360_,
		_w17361_,
		_w17362_
	);
	LUT3 #(
		.INIT('h80)
	) name15462 (
		\m0_data_i[29]_pad ,
		_w9029_,
		_w9030_,
		_w17363_
	);
	LUT3 #(
		.INIT('h80)
	) name15463 (
		\m2_data_i[29]_pad ,
		_w9029_,
		_w9030_,
		_w17364_
	);
	LUT4 #(
		.INIT('h3b7f)
	) name15464 (
		_w9024_,
		_w9027_,
		_w17363_,
		_w17364_,
		_w17365_
	);
	LUT3 #(
		.INIT('h2a)
	) name15465 (
		\m7_data_i[29]_pad ,
		_w9029_,
		_w9030_,
		_w17366_
	);
	LUT3 #(
		.INIT('h2a)
	) name15466 (
		\m1_data_i[29]_pad ,
		_w9029_,
		_w9030_,
		_w17367_
	);
	LUT4 #(
		.INIT('h67ef)
	) name15467 (
		_w9024_,
		_w9027_,
		_w17366_,
		_w17367_,
		_w17368_
	);
	LUT3 #(
		.INIT('h2a)
	) name15468 (
		\m3_data_i[29]_pad ,
		_w9029_,
		_w9030_,
		_w17369_
	);
	LUT3 #(
		.INIT('h80)
	) name15469 (
		\m4_data_i[29]_pad ,
		_w9029_,
		_w9030_,
		_w17370_
	);
	LUT4 #(
		.INIT('h9dbf)
	) name15470 (
		_w9024_,
		_w9027_,
		_w17369_,
		_w17370_,
		_w17371_
	);
	LUT4 #(
		.INIT('h7fff)
	) name15471 (
		_w17362_,
		_w17365_,
		_w17368_,
		_w17371_,
		_w17372_
	);
	LUT3 #(
		.INIT('h2a)
	) name15472 (
		\m1_data_i[2]_pad ,
		_w9029_,
		_w9030_,
		_w17373_
	);
	LUT3 #(
		.INIT('h80)
	) name15473 (
		\m2_data_i[2]_pad ,
		_w9029_,
		_w9030_,
		_w17374_
	);
	LUT4 #(
		.INIT('h3b7f)
	) name15474 (
		_w9024_,
		_w9027_,
		_w17373_,
		_w17374_,
		_w17375_
	);
	LUT3 #(
		.INIT('h80)
	) name15475 (
		\m0_data_i[2]_pad ,
		_w9029_,
		_w9030_,
		_w17376_
	);
	LUT3 #(
		.INIT('h2a)
	) name15476 (
		\m5_data_i[2]_pad ,
		_w9029_,
		_w9030_,
		_w17377_
	);
	LUT4 #(
		.INIT('h5d7f)
	) name15477 (
		_w9024_,
		_w9027_,
		_w17376_,
		_w17377_,
		_w17378_
	);
	LUT3 #(
		.INIT('h2a)
	) name15478 (
		\m7_data_i[2]_pad ,
		_w9029_,
		_w9030_,
		_w17379_
	);
	LUT3 #(
		.INIT('h80)
	) name15479 (
		\m6_data_i[2]_pad ,
		_w9029_,
		_w9030_,
		_w17380_
	);
	LUT3 #(
		.INIT('h57)
	) name15480 (
		_w9036_,
		_w17379_,
		_w17380_,
		_w17381_
	);
	LUT3 #(
		.INIT('h2a)
	) name15481 (
		\m3_data_i[2]_pad ,
		_w9029_,
		_w9030_,
		_w17382_
	);
	LUT3 #(
		.INIT('h80)
	) name15482 (
		\m4_data_i[2]_pad ,
		_w9029_,
		_w9030_,
		_w17383_
	);
	LUT4 #(
		.INIT('h9dbf)
	) name15483 (
		_w9024_,
		_w9027_,
		_w17382_,
		_w17383_,
		_w17384_
	);
	LUT4 #(
		.INIT('h7fff)
	) name15484 (
		_w17375_,
		_w17378_,
		_w17381_,
		_w17384_,
		_w17385_
	);
	LUT3 #(
		.INIT('h2a)
	) name15485 (
		\m3_data_i[30]_pad ,
		_w9029_,
		_w9030_,
		_w17386_
	);
	LUT3 #(
		.INIT('h80)
	) name15486 (
		\m4_data_i[30]_pad ,
		_w9029_,
		_w9030_,
		_w17387_
	);
	LUT4 #(
		.INIT('h9dbf)
	) name15487 (
		_w9024_,
		_w9027_,
		_w17386_,
		_w17387_,
		_w17388_
	);
	LUT3 #(
		.INIT('h80)
	) name15488 (
		\m0_data_i[30]_pad ,
		_w9029_,
		_w9030_,
		_w17389_
	);
	LUT3 #(
		.INIT('h2a)
	) name15489 (
		\m5_data_i[30]_pad ,
		_w9029_,
		_w9030_,
		_w17390_
	);
	LUT4 #(
		.INIT('h5d7f)
	) name15490 (
		_w9024_,
		_w9027_,
		_w17389_,
		_w17390_,
		_w17391_
	);
	LUT3 #(
		.INIT('h2a)
	) name15491 (
		\m7_data_i[30]_pad ,
		_w9029_,
		_w9030_,
		_w17392_
	);
	LUT3 #(
		.INIT('h80)
	) name15492 (
		\m6_data_i[30]_pad ,
		_w9029_,
		_w9030_,
		_w17393_
	);
	LUT3 #(
		.INIT('h57)
	) name15493 (
		_w9036_,
		_w17392_,
		_w17393_,
		_w17394_
	);
	LUT3 #(
		.INIT('h2a)
	) name15494 (
		\m1_data_i[30]_pad ,
		_w9029_,
		_w9030_,
		_w17395_
	);
	LUT3 #(
		.INIT('h80)
	) name15495 (
		\m2_data_i[30]_pad ,
		_w9029_,
		_w9030_,
		_w17396_
	);
	LUT4 #(
		.INIT('h3b7f)
	) name15496 (
		_w9024_,
		_w9027_,
		_w17395_,
		_w17396_,
		_w17397_
	);
	LUT4 #(
		.INIT('h7fff)
	) name15497 (
		_w17388_,
		_w17391_,
		_w17394_,
		_w17397_,
		_w17398_
	);
	LUT3 #(
		.INIT('h2a)
	) name15498 (
		\m1_data_i[31]_pad ,
		_w9029_,
		_w9030_,
		_w17399_
	);
	LUT3 #(
		.INIT('h80)
	) name15499 (
		\m2_data_i[31]_pad ,
		_w9029_,
		_w9030_,
		_w17400_
	);
	LUT4 #(
		.INIT('h3b7f)
	) name15500 (
		_w9024_,
		_w9027_,
		_w17399_,
		_w17400_,
		_w17401_
	);
	LUT3 #(
		.INIT('h80)
	) name15501 (
		\m0_data_i[31]_pad ,
		_w9029_,
		_w9030_,
		_w17402_
	);
	LUT3 #(
		.INIT('h80)
	) name15502 (
		\m4_data_i[31]_pad ,
		_w9029_,
		_w9030_,
		_w17403_
	);
	LUT4 #(
		.INIT('h5d7f)
	) name15503 (
		_w9024_,
		_w9027_,
		_w17402_,
		_w17403_,
		_w17404_
	);
	LUT3 #(
		.INIT('h2a)
	) name15504 (
		\m7_data_i[31]_pad ,
		_w9029_,
		_w9030_,
		_w17405_
	);
	LUT3 #(
		.INIT('h2a)
	) name15505 (
		\m3_data_i[31]_pad ,
		_w9029_,
		_w9030_,
		_w17406_
	);
	LUT4 #(
		.INIT('habef)
	) name15506 (
		_w9024_,
		_w9027_,
		_w17405_,
		_w17406_,
		_w17407_
	);
	LUT3 #(
		.INIT('h80)
	) name15507 (
		\m6_data_i[31]_pad ,
		_w9029_,
		_w9030_,
		_w17408_
	);
	LUT3 #(
		.INIT('h2a)
	) name15508 (
		\m5_data_i[31]_pad ,
		_w9029_,
		_w9030_,
		_w17409_
	);
	LUT4 #(
		.INIT('hcdef)
	) name15509 (
		_w9024_,
		_w9027_,
		_w17408_,
		_w17409_,
		_w17410_
	);
	LUT4 #(
		.INIT('h7fff)
	) name15510 (
		_w17401_,
		_w17404_,
		_w17407_,
		_w17410_,
		_w17411_
	);
	LUT3 #(
		.INIT('h80)
	) name15511 (
		\m6_data_i[3]_pad ,
		_w9029_,
		_w9030_,
		_w17412_
	);
	LUT3 #(
		.INIT('h2a)
	) name15512 (
		\m5_data_i[3]_pad ,
		_w9029_,
		_w9030_,
		_w17413_
	);
	LUT4 #(
		.INIT('hcdef)
	) name15513 (
		_w9024_,
		_w9027_,
		_w17412_,
		_w17413_,
		_w17414_
	);
	LUT3 #(
		.INIT('h2a)
	) name15514 (
		\m1_data_i[3]_pad ,
		_w9029_,
		_w9030_,
		_w17415_
	);
	LUT3 #(
		.INIT('h80)
	) name15515 (
		\m4_data_i[3]_pad ,
		_w9029_,
		_w9030_,
		_w17416_
	);
	LUT4 #(
		.INIT('h5d7f)
	) name15516 (
		_w9024_,
		_w9027_,
		_w17415_,
		_w17416_,
		_w17417_
	);
	LUT3 #(
		.INIT('h80)
	) name15517 (
		\m2_data_i[3]_pad ,
		_w9029_,
		_w9030_,
		_w17418_
	);
	LUT3 #(
		.INIT('h2a)
	) name15518 (
		\m3_data_i[3]_pad ,
		_w9029_,
		_w9030_,
		_w17419_
	);
	LUT3 #(
		.INIT('h57)
	) name15519 (
		_w9028_,
		_w17418_,
		_w17419_,
		_w17420_
	);
	LUT3 #(
		.INIT('h80)
	) name15520 (
		\m0_data_i[3]_pad ,
		_w9029_,
		_w9030_,
		_w17421_
	);
	LUT3 #(
		.INIT('h2a)
	) name15521 (
		\m7_data_i[3]_pad ,
		_w9029_,
		_w9030_,
		_w17422_
	);
	LUT4 #(
		.INIT('h6e7f)
	) name15522 (
		_w9024_,
		_w9027_,
		_w17421_,
		_w17422_,
		_w17423_
	);
	LUT4 #(
		.INIT('h7fff)
	) name15523 (
		_w17414_,
		_w17417_,
		_w17420_,
		_w17423_,
		_w17424_
	);
	LUT3 #(
		.INIT('h2a)
	) name15524 (
		\m1_data_i[4]_pad ,
		_w9029_,
		_w9030_,
		_w17425_
	);
	LUT3 #(
		.INIT('h80)
	) name15525 (
		\m2_data_i[4]_pad ,
		_w9029_,
		_w9030_,
		_w17426_
	);
	LUT4 #(
		.INIT('h3b7f)
	) name15526 (
		_w9024_,
		_w9027_,
		_w17425_,
		_w17426_,
		_w17427_
	);
	LUT3 #(
		.INIT('h80)
	) name15527 (
		\m0_data_i[4]_pad ,
		_w9029_,
		_w9030_,
		_w17428_
	);
	LUT3 #(
		.INIT('h80)
	) name15528 (
		\m4_data_i[4]_pad ,
		_w9029_,
		_w9030_,
		_w17429_
	);
	LUT4 #(
		.INIT('h5d7f)
	) name15529 (
		_w9024_,
		_w9027_,
		_w17428_,
		_w17429_,
		_w17430_
	);
	LUT3 #(
		.INIT('h2a)
	) name15530 (
		\m7_data_i[4]_pad ,
		_w9029_,
		_w9030_,
		_w17431_
	);
	LUT3 #(
		.INIT('h2a)
	) name15531 (
		\m3_data_i[4]_pad ,
		_w9029_,
		_w9030_,
		_w17432_
	);
	LUT4 #(
		.INIT('habef)
	) name15532 (
		_w9024_,
		_w9027_,
		_w17431_,
		_w17432_,
		_w17433_
	);
	LUT3 #(
		.INIT('h80)
	) name15533 (
		\m6_data_i[4]_pad ,
		_w9029_,
		_w9030_,
		_w17434_
	);
	LUT3 #(
		.INIT('h2a)
	) name15534 (
		\m5_data_i[4]_pad ,
		_w9029_,
		_w9030_,
		_w17435_
	);
	LUT4 #(
		.INIT('hcdef)
	) name15535 (
		_w9024_,
		_w9027_,
		_w17434_,
		_w17435_,
		_w17436_
	);
	LUT4 #(
		.INIT('h7fff)
	) name15536 (
		_w17427_,
		_w17430_,
		_w17433_,
		_w17436_,
		_w17437_
	);
	LUT3 #(
		.INIT('h2a)
	) name15537 (
		\m3_data_i[5]_pad ,
		_w9029_,
		_w9030_,
		_w17438_
	);
	LUT3 #(
		.INIT('h80)
	) name15538 (
		\m4_data_i[5]_pad ,
		_w9029_,
		_w9030_,
		_w17439_
	);
	LUT4 #(
		.INIT('h9dbf)
	) name15539 (
		_w9024_,
		_w9027_,
		_w17438_,
		_w17439_,
		_w17440_
	);
	LUT3 #(
		.INIT('h80)
	) name15540 (
		\m0_data_i[5]_pad ,
		_w9029_,
		_w9030_,
		_w17441_
	);
	LUT3 #(
		.INIT('h80)
	) name15541 (
		\m2_data_i[5]_pad ,
		_w9029_,
		_w9030_,
		_w17442_
	);
	LUT4 #(
		.INIT('h3b7f)
	) name15542 (
		_w9024_,
		_w9027_,
		_w17441_,
		_w17442_,
		_w17443_
	);
	LUT3 #(
		.INIT('h2a)
	) name15543 (
		\m7_data_i[5]_pad ,
		_w9029_,
		_w9030_,
		_w17444_
	);
	LUT3 #(
		.INIT('h2a)
	) name15544 (
		\m1_data_i[5]_pad ,
		_w9029_,
		_w9030_,
		_w17445_
	);
	LUT4 #(
		.INIT('h67ef)
	) name15545 (
		_w9024_,
		_w9027_,
		_w17444_,
		_w17445_,
		_w17446_
	);
	LUT3 #(
		.INIT('h80)
	) name15546 (
		\m6_data_i[5]_pad ,
		_w9029_,
		_w9030_,
		_w17447_
	);
	LUT3 #(
		.INIT('h2a)
	) name15547 (
		\m5_data_i[5]_pad ,
		_w9029_,
		_w9030_,
		_w17448_
	);
	LUT4 #(
		.INIT('hcdef)
	) name15548 (
		_w9024_,
		_w9027_,
		_w17447_,
		_w17448_,
		_w17449_
	);
	LUT4 #(
		.INIT('h7fff)
	) name15549 (
		_w17440_,
		_w17443_,
		_w17446_,
		_w17449_,
		_w17450_
	);
	LUT3 #(
		.INIT('h2a)
	) name15550 (
		\m3_data_i[6]_pad ,
		_w9029_,
		_w9030_,
		_w17451_
	);
	LUT3 #(
		.INIT('h80)
	) name15551 (
		\m4_data_i[6]_pad ,
		_w9029_,
		_w9030_,
		_w17452_
	);
	LUT4 #(
		.INIT('h9dbf)
	) name15552 (
		_w9024_,
		_w9027_,
		_w17451_,
		_w17452_,
		_w17453_
	);
	LUT3 #(
		.INIT('h80)
	) name15553 (
		\m6_data_i[6]_pad ,
		_w9029_,
		_w9030_,
		_w17454_
	);
	LUT3 #(
		.INIT('h2a)
	) name15554 (
		\m7_data_i[6]_pad ,
		_w9029_,
		_w9030_,
		_w17455_
	);
	LUT3 #(
		.INIT('h57)
	) name15555 (
		_w9036_,
		_w17454_,
		_w17455_,
		_w17456_
	);
	LUT3 #(
		.INIT('h2a)
	) name15556 (
		\m5_data_i[6]_pad ,
		_w9029_,
		_w9030_,
		_w17457_
	);
	LUT3 #(
		.INIT('h80)
	) name15557 (
		\m0_data_i[6]_pad ,
		_w9029_,
		_w9030_,
		_w17458_
	);
	LUT4 #(
		.INIT('h57df)
	) name15558 (
		_w9024_,
		_w9027_,
		_w17457_,
		_w17458_,
		_w17459_
	);
	LUT3 #(
		.INIT('h2a)
	) name15559 (
		\m1_data_i[6]_pad ,
		_w9029_,
		_w9030_,
		_w17460_
	);
	LUT3 #(
		.INIT('h80)
	) name15560 (
		\m2_data_i[6]_pad ,
		_w9029_,
		_w9030_,
		_w17461_
	);
	LUT4 #(
		.INIT('h3b7f)
	) name15561 (
		_w9024_,
		_w9027_,
		_w17460_,
		_w17461_,
		_w17462_
	);
	LUT4 #(
		.INIT('h7fff)
	) name15562 (
		_w17453_,
		_w17456_,
		_w17459_,
		_w17462_,
		_w17463_
	);
	LUT3 #(
		.INIT('h2a)
	) name15563 (
		\m3_data_i[7]_pad ,
		_w9029_,
		_w9030_,
		_w17464_
	);
	LUT3 #(
		.INIT('h80)
	) name15564 (
		\m4_data_i[7]_pad ,
		_w9029_,
		_w9030_,
		_w17465_
	);
	LUT4 #(
		.INIT('h9dbf)
	) name15565 (
		_w9024_,
		_w9027_,
		_w17464_,
		_w17465_,
		_w17466_
	);
	LUT3 #(
		.INIT('h80)
	) name15566 (
		\m0_data_i[7]_pad ,
		_w9029_,
		_w9030_,
		_w17467_
	);
	LUT3 #(
		.INIT('h80)
	) name15567 (
		\m2_data_i[7]_pad ,
		_w9029_,
		_w9030_,
		_w17468_
	);
	LUT4 #(
		.INIT('h3b7f)
	) name15568 (
		_w9024_,
		_w9027_,
		_w17467_,
		_w17468_,
		_w17469_
	);
	LUT3 #(
		.INIT('h2a)
	) name15569 (
		\m7_data_i[7]_pad ,
		_w9029_,
		_w9030_,
		_w17470_
	);
	LUT3 #(
		.INIT('h2a)
	) name15570 (
		\m1_data_i[7]_pad ,
		_w9029_,
		_w9030_,
		_w17471_
	);
	LUT4 #(
		.INIT('h67ef)
	) name15571 (
		_w9024_,
		_w9027_,
		_w17470_,
		_w17471_,
		_w17472_
	);
	LUT3 #(
		.INIT('h80)
	) name15572 (
		\m6_data_i[7]_pad ,
		_w9029_,
		_w9030_,
		_w17473_
	);
	LUT3 #(
		.INIT('h2a)
	) name15573 (
		\m5_data_i[7]_pad ,
		_w9029_,
		_w9030_,
		_w17474_
	);
	LUT4 #(
		.INIT('hcdef)
	) name15574 (
		_w9024_,
		_w9027_,
		_w17473_,
		_w17474_,
		_w17475_
	);
	LUT4 #(
		.INIT('h7fff)
	) name15575 (
		_w17466_,
		_w17469_,
		_w17472_,
		_w17475_,
		_w17476_
	);
	LUT3 #(
		.INIT('h2a)
	) name15576 (
		\m1_data_i[8]_pad ,
		_w9029_,
		_w9030_,
		_w17477_
	);
	LUT3 #(
		.INIT('h80)
	) name15577 (
		\m2_data_i[8]_pad ,
		_w9029_,
		_w9030_,
		_w17478_
	);
	LUT4 #(
		.INIT('h3b7f)
	) name15578 (
		_w9024_,
		_w9027_,
		_w17477_,
		_w17478_,
		_w17479_
	);
	LUT3 #(
		.INIT('h80)
	) name15579 (
		\m0_data_i[8]_pad ,
		_w9029_,
		_w9030_,
		_w17480_
	);
	LUT3 #(
		.INIT('h80)
	) name15580 (
		\m4_data_i[8]_pad ,
		_w9029_,
		_w9030_,
		_w17481_
	);
	LUT4 #(
		.INIT('h5d7f)
	) name15581 (
		_w9024_,
		_w9027_,
		_w17480_,
		_w17481_,
		_w17482_
	);
	LUT3 #(
		.INIT('h2a)
	) name15582 (
		\m7_data_i[8]_pad ,
		_w9029_,
		_w9030_,
		_w17483_
	);
	LUT3 #(
		.INIT('h2a)
	) name15583 (
		\m3_data_i[8]_pad ,
		_w9029_,
		_w9030_,
		_w17484_
	);
	LUT4 #(
		.INIT('habef)
	) name15584 (
		_w9024_,
		_w9027_,
		_w17483_,
		_w17484_,
		_w17485_
	);
	LUT3 #(
		.INIT('h80)
	) name15585 (
		\m6_data_i[8]_pad ,
		_w9029_,
		_w9030_,
		_w17486_
	);
	LUT3 #(
		.INIT('h2a)
	) name15586 (
		\m5_data_i[8]_pad ,
		_w9029_,
		_w9030_,
		_w17487_
	);
	LUT4 #(
		.INIT('hcdef)
	) name15587 (
		_w9024_,
		_w9027_,
		_w17486_,
		_w17487_,
		_w17488_
	);
	LUT4 #(
		.INIT('h7fff)
	) name15588 (
		_w17479_,
		_w17482_,
		_w17485_,
		_w17488_,
		_w17489_
	);
	LUT3 #(
		.INIT('h2a)
	) name15589 (
		\m1_data_i[9]_pad ,
		_w9029_,
		_w9030_,
		_w17490_
	);
	LUT3 #(
		.INIT('h80)
	) name15590 (
		\m2_data_i[9]_pad ,
		_w9029_,
		_w9030_,
		_w17491_
	);
	LUT4 #(
		.INIT('h3b7f)
	) name15591 (
		_w9024_,
		_w9027_,
		_w17490_,
		_w17491_,
		_w17492_
	);
	LUT3 #(
		.INIT('h80)
	) name15592 (
		\m0_data_i[9]_pad ,
		_w9029_,
		_w9030_,
		_w17493_
	);
	LUT3 #(
		.INIT('h80)
	) name15593 (
		\m4_data_i[9]_pad ,
		_w9029_,
		_w9030_,
		_w17494_
	);
	LUT4 #(
		.INIT('h5d7f)
	) name15594 (
		_w9024_,
		_w9027_,
		_w17493_,
		_w17494_,
		_w17495_
	);
	LUT3 #(
		.INIT('h2a)
	) name15595 (
		\m7_data_i[9]_pad ,
		_w9029_,
		_w9030_,
		_w17496_
	);
	LUT3 #(
		.INIT('h2a)
	) name15596 (
		\m3_data_i[9]_pad ,
		_w9029_,
		_w9030_,
		_w17497_
	);
	LUT4 #(
		.INIT('habef)
	) name15597 (
		_w9024_,
		_w9027_,
		_w17496_,
		_w17497_,
		_w17498_
	);
	LUT3 #(
		.INIT('h80)
	) name15598 (
		\m6_data_i[9]_pad ,
		_w9029_,
		_w9030_,
		_w17499_
	);
	LUT3 #(
		.INIT('h2a)
	) name15599 (
		\m5_data_i[9]_pad ,
		_w9029_,
		_w9030_,
		_w17500_
	);
	LUT4 #(
		.INIT('hcdef)
	) name15600 (
		_w9024_,
		_w9027_,
		_w17499_,
		_w17500_,
		_w17501_
	);
	LUT4 #(
		.INIT('h7fff)
	) name15601 (
		_w17492_,
		_w17495_,
		_w17498_,
		_w17501_,
		_w17502_
	);
	LUT3 #(
		.INIT('h2a)
	) name15602 (
		\m3_sel_i[0]_pad ,
		_w9029_,
		_w9030_,
		_w17503_
	);
	LUT3 #(
		.INIT('h80)
	) name15603 (
		\m4_sel_i[0]_pad ,
		_w9029_,
		_w9030_,
		_w17504_
	);
	LUT4 #(
		.INIT('h9dbf)
	) name15604 (
		_w9024_,
		_w9027_,
		_w17503_,
		_w17504_,
		_w17505_
	);
	LUT3 #(
		.INIT('h80)
	) name15605 (
		\m6_sel_i[0]_pad ,
		_w9029_,
		_w9030_,
		_w17506_
	);
	LUT3 #(
		.INIT('h80)
	) name15606 (
		\m2_sel_i[0]_pad ,
		_w9029_,
		_w9030_,
		_w17507_
	);
	LUT4 #(
		.INIT('habef)
	) name15607 (
		_w9024_,
		_w9027_,
		_w17506_,
		_w17507_,
		_w17508_
	);
	LUT3 #(
		.INIT('h2a)
	) name15608 (
		\m5_sel_i[0]_pad ,
		_w9029_,
		_w9030_,
		_w17509_
	);
	LUT3 #(
		.INIT('h2a)
	) name15609 (
		\m1_sel_i[0]_pad ,
		_w9029_,
		_w9030_,
		_w17510_
	);
	LUT4 #(
		.INIT('h57df)
	) name15610 (
		_w9024_,
		_w9027_,
		_w17509_,
		_w17510_,
		_w17511_
	);
	LUT3 #(
		.INIT('h80)
	) name15611 (
		\m0_sel_i[0]_pad ,
		_w9029_,
		_w9030_,
		_w17512_
	);
	LUT3 #(
		.INIT('h2a)
	) name15612 (
		\m7_sel_i[0]_pad ,
		_w9029_,
		_w9030_,
		_w17513_
	);
	LUT4 #(
		.INIT('h6e7f)
	) name15613 (
		_w9024_,
		_w9027_,
		_w17512_,
		_w17513_,
		_w17514_
	);
	LUT4 #(
		.INIT('h7fff)
	) name15614 (
		_w17505_,
		_w17508_,
		_w17511_,
		_w17514_,
		_w17515_
	);
	LUT3 #(
		.INIT('h2a)
	) name15615 (
		\m3_sel_i[1]_pad ,
		_w9029_,
		_w9030_,
		_w17516_
	);
	LUT3 #(
		.INIT('h80)
	) name15616 (
		\m4_sel_i[1]_pad ,
		_w9029_,
		_w9030_,
		_w17517_
	);
	LUT4 #(
		.INIT('h9dbf)
	) name15617 (
		_w9024_,
		_w9027_,
		_w17516_,
		_w17517_,
		_w17518_
	);
	LUT3 #(
		.INIT('h80)
	) name15618 (
		\m6_sel_i[1]_pad ,
		_w9029_,
		_w9030_,
		_w17519_
	);
	LUT3 #(
		.INIT('h80)
	) name15619 (
		\m2_sel_i[1]_pad ,
		_w9029_,
		_w9030_,
		_w17520_
	);
	LUT4 #(
		.INIT('habef)
	) name15620 (
		_w9024_,
		_w9027_,
		_w17519_,
		_w17520_,
		_w17521_
	);
	LUT3 #(
		.INIT('h2a)
	) name15621 (
		\m5_sel_i[1]_pad ,
		_w9029_,
		_w9030_,
		_w17522_
	);
	LUT3 #(
		.INIT('h2a)
	) name15622 (
		\m1_sel_i[1]_pad ,
		_w9029_,
		_w9030_,
		_w17523_
	);
	LUT4 #(
		.INIT('h57df)
	) name15623 (
		_w9024_,
		_w9027_,
		_w17522_,
		_w17523_,
		_w17524_
	);
	LUT3 #(
		.INIT('h80)
	) name15624 (
		\m0_sel_i[1]_pad ,
		_w9029_,
		_w9030_,
		_w17525_
	);
	LUT3 #(
		.INIT('h2a)
	) name15625 (
		\m7_sel_i[1]_pad ,
		_w9029_,
		_w9030_,
		_w17526_
	);
	LUT4 #(
		.INIT('h6e7f)
	) name15626 (
		_w9024_,
		_w9027_,
		_w17525_,
		_w17526_,
		_w17527_
	);
	LUT4 #(
		.INIT('h7fff)
	) name15627 (
		_w17518_,
		_w17521_,
		_w17524_,
		_w17527_,
		_w17528_
	);
	LUT3 #(
		.INIT('h2a)
	) name15628 (
		\m3_sel_i[2]_pad ,
		_w9029_,
		_w9030_,
		_w17529_
	);
	LUT3 #(
		.INIT('h80)
	) name15629 (
		\m4_sel_i[2]_pad ,
		_w9029_,
		_w9030_,
		_w17530_
	);
	LUT4 #(
		.INIT('h9dbf)
	) name15630 (
		_w9024_,
		_w9027_,
		_w17529_,
		_w17530_,
		_w17531_
	);
	LUT3 #(
		.INIT('h80)
	) name15631 (
		\m6_sel_i[2]_pad ,
		_w9029_,
		_w9030_,
		_w17532_
	);
	LUT3 #(
		.INIT('h80)
	) name15632 (
		\m2_sel_i[2]_pad ,
		_w9029_,
		_w9030_,
		_w17533_
	);
	LUT4 #(
		.INIT('habef)
	) name15633 (
		_w9024_,
		_w9027_,
		_w17532_,
		_w17533_,
		_w17534_
	);
	LUT3 #(
		.INIT('h2a)
	) name15634 (
		\m5_sel_i[2]_pad ,
		_w9029_,
		_w9030_,
		_w17535_
	);
	LUT3 #(
		.INIT('h2a)
	) name15635 (
		\m1_sel_i[2]_pad ,
		_w9029_,
		_w9030_,
		_w17536_
	);
	LUT4 #(
		.INIT('h57df)
	) name15636 (
		_w9024_,
		_w9027_,
		_w17535_,
		_w17536_,
		_w17537_
	);
	LUT3 #(
		.INIT('h80)
	) name15637 (
		\m0_sel_i[2]_pad ,
		_w9029_,
		_w9030_,
		_w17538_
	);
	LUT3 #(
		.INIT('h2a)
	) name15638 (
		\m7_sel_i[2]_pad ,
		_w9029_,
		_w9030_,
		_w17539_
	);
	LUT4 #(
		.INIT('h6e7f)
	) name15639 (
		_w9024_,
		_w9027_,
		_w17538_,
		_w17539_,
		_w17540_
	);
	LUT4 #(
		.INIT('h7fff)
	) name15640 (
		_w17531_,
		_w17534_,
		_w17537_,
		_w17540_,
		_w17541_
	);
	LUT3 #(
		.INIT('h2a)
	) name15641 (
		\m3_sel_i[3]_pad ,
		_w9029_,
		_w9030_,
		_w17542_
	);
	LUT3 #(
		.INIT('h80)
	) name15642 (
		\m4_sel_i[3]_pad ,
		_w9029_,
		_w9030_,
		_w17543_
	);
	LUT4 #(
		.INIT('h9dbf)
	) name15643 (
		_w9024_,
		_w9027_,
		_w17542_,
		_w17543_,
		_w17544_
	);
	LUT3 #(
		.INIT('h80)
	) name15644 (
		\m6_sel_i[3]_pad ,
		_w9029_,
		_w9030_,
		_w17545_
	);
	LUT3 #(
		.INIT('h80)
	) name15645 (
		\m2_sel_i[3]_pad ,
		_w9029_,
		_w9030_,
		_w17546_
	);
	LUT4 #(
		.INIT('habef)
	) name15646 (
		_w9024_,
		_w9027_,
		_w17545_,
		_w17546_,
		_w17547_
	);
	LUT3 #(
		.INIT('h2a)
	) name15647 (
		\m5_sel_i[3]_pad ,
		_w9029_,
		_w9030_,
		_w17548_
	);
	LUT3 #(
		.INIT('h2a)
	) name15648 (
		\m1_sel_i[3]_pad ,
		_w9029_,
		_w9030_,
		_w17549_
	);
	LUT4 #(
		.INIT('h57df)
	) name15649 (
		_w9024_,
		_w9027_,
		_w17548_,
		_w17549_,
		_w17550_
	);
	LUT3 #(
		.INIT('h80)
	) name15650 (
		\m0_sel_i[3]_pad ,
		_w9029_,
		_w9030_,
		_w17551_
	);
	LUT3 #(
		.INIT('h2a)
	) name15651 (
		\m7_sel_i[3]_pad ,
		_w9029_,
		_w9030_,
		_w17552_
	);
	LUT4 #(
		.INIT('h6e7f)
	) name15652 (
		_w9024_,
		_w9027_,
		_w17551_,
		_w17552_,
		_w17553_
	);
	LUT4 #(
		.INIT('h7fff)
	) name15653 (
		_w17544_,
		_w17547_,
		_w17550_,
		_w17553_,
		_w17554_
	);
	LUT4 #(
		.INIT('h2a00)
	) name15654 (
		\m7_stb_i_pad ,
		_w9029_,
		_w9030_,
		_w9339_,
		_w17555_
	);
	LUT4 #(
		.INIT('h8000)
	) name15655 (
		\m6_stb_i_pad ,
		_w9029_,
		_w9030_,
		_w9565_,
		_w17556_
	);
	LUT3 #(
		.INIT('h57)
	) name15656 (
		_w9036_,
		_w17555_,
		_w17556_,
		_w17557_
	);
	LUT4 #(
		.INIT('h8000)
	) name15657 (
		\m4_stb_i_pad ,
		_w9029_,
		_w9030_,
		_w9512_,
		_w17558_
	);
	LUT4 #(
		.INIT('h2a00)
	) name15658 (
		\m1_stb_i_pad ,
		_w9029_,
		_w9030_,
		_w9635_,
		_w17559_
	);
	LUT4 #(
		.INIT('h57df)
	) name15659 (
		_w9024_,
		_w9027_,
		_w17558_,
		_w17559_,
		_w17560_
	);
	LUT4 #(
		.INIT('h2a00)
	) name15660 (
		\m5_stb_i_pad ,
		_w9029_,
		_w9030_,
		_w9354_,
		_w17561_
	);
	LUT4 #(
		.INIT('h2a00)
	) name15661 (
		\m3_stb_i_pad ,
		_w9029_,
		_w9030_,
		_w9486_,
		_w17562_
	);
	LUT4 #(
		.INIT('h9bdf)
	) name15662 (
		_w9024_,
		_w9027_,
		_w17561_,
		_w17562_,
		_w17563_
	);
	LUT4 #(
		.INIT('h8000)
	) name15663 (
		\m2_stb_i_pad ,
		_w9029_,
		_w9030_,
		_w9457_,
		_w17564_
	);
	LUT4 #(
		.INIT('h8000)
	) name15664 (
		\m0_stb_i_pad ,
		_w9029_,
		_w9030_,
		_w9650_,
		_w17565_
	);
	LUT4 #(
		.INIT('h37bf)
	) name15665 (
		_w9024_,
		_w9027_,
		_w17564_,
		_w17565_,
		_w17566_
	);
	LUT4 #(
		.INIT('h7fff)
	) name15666 (
		_w17557_,
		_w17560_,
		_w17563_,
		_w17566_,
		_w17567_
	);
	LUT3 #(
		.INIT('h2a)
	) name15667 (
		\m3_we_i_pad ,
		_w9029_,
		_w9030_,
		_w17568_
	);
	LUT3 #(
		.INIT('h80)
	) name15668 (
		\m4_we_i_pad ,
		_w9029_,
		_w9030_,
		_w17569_
	);
	LUT4 #(
		.INIT('h9dbf)
	) name15669 (
		_w9024_,
		_w9027_,
		_w17568_,
		_w17569_,
		_w17570_
	);
	LUT3 #(
		.INIT('h80)
	) name15670 (
		\m6_we_i_pad ,
		_w9029_,
		_w9030_,
		_w17571_
	);
	LUT3 #(
		.INIT('h80)
	) name15671 (
		\m2_we_i_pad ,
		_w9029_,
		_w9030_,
		_w17572_
	);
	LUT4 #(
		.INIT('habef)
	) name15672 (
		_w9024_,
		_w9027_,
		_w17571_,
		_w17572_,
		_w17573_
	);
	LUT3 #(
		.INIT('h2a)
	) name15673 (
		\m5_we_i_pad ,
		_w9029_,
		_w9030_,
		_w17574_
	);
	LUT3 #(
		.INIT('h2a)
	) name15674 (
		\m1_we_i_pad ,
		_w9029_,
		_w9030_,
		_w17575_
	);
	LUT4 #(
		.INIT('h57df)
	) name15675 (
		_w9024_,
		_w9027_,
		_w17574_,
		_w17575_,
		_w17576_
	);
	LUT3 #(
		.INIT('h80)
	) name15676 (
		\m0_we_i_pad ,
		_w9029_,
		_w9030_,
		_w17577_
	);
	LUT3 #(
		.INIT('h2a)
	) name15677 (
		\m7_we_i_pad ,
		_w9029_,
		_w9030_,
		_w17578_
	);
	LUT4 #(
		.INIT('h6e7f)
	) name15678 (
		_w9024_,
		_w9027_,
		_w17577_,
		_w17578_,
		_w17579_
	);
	LUT4 #(
		.INIT('h7fff)
	) name15679 (
		_w17570_,
		_w17573_,
		_w17576_,
		_w17579_,
		_w17580_
	);
	LUT3 #(
		.INIT('h80)
	) name15680 (
		\m6_addr_i[0]_pad ,
		_w9069_,
		_w9070_,
		_w17581_
	);
	LUT3 #(
		.INIT('h2a)
	) name15681 (
		\m5_addr_i[0]_pad ,
		_w9069_,
		_w9070_,
		_w17582_
	);
	LUT4 #(
		.INIT('hcdef)
	) name15682 (
		_w9064_,
		_w9067_,
		_w17581_,
		_w17582_,
		_w17583_
	);
	LUT3 #(
		.INIT('h80)
	) name15683 (
		\m0_addr_i[0]_pad ,
		_w9069_,
		_w9070_,
		_w17584_
	);
	LUT3 #(
		.INIT('h80)
	) name15684 (
		\m4_addr_i[0]_pad ,
		_w9069_,
		_w9070_,
		_w17585_
	);
	LUT4 #(
		.INIT('h5d7f)
	) name15685 (
		_w9064_,
		_w9067_,
		_w17584_,
		_w17585_,
		_w17586_
	);
	LUT3 #(
		.INIT('h2a)
	) name15686 (
		\m7_addr_i[0]_pad ,
		_w9069_,
		_w9070_,
		_w17587_
	);
	LUT3 #(
		.INIT('h2a)
	) name15687 (
		\m3_addr_i[0]_pad ,
		_w9069_,
		_w9070_,
		_w17588_
	);
	LUT4 #(
		.INIT('habef)
	) name15688 (
		_w9064_,
		_w9067_,
		_w17587_,
		_w17588_,
		_w17589_
	);
	LUT3 #(
		.INIT('h2a)
	) name15689 (
		\m1_addr_i[0]_pad ,
		_w9069_,
		_w9070_,
		_w17590_
	);
	LUT3 #(
		.INIT('h80)
	) name15690 (
		\m2_addr_i[0]_pad ,
		_w9069_,
		_w9070_,
		_w17591_
	);
	LUT4 #(
		.INIT('h3b7f)
	) name15691 (
		_w9064_,
		_w9067_,
		_w17590_,
		_w17591_,
		_w17592_
	);
	LUT4 #(
		.INIT('h7fff)
	) name15692 (
		_w17583_,
		_w17586_,
		_w17589_,
		_w17592_,
		_w17593_
	);
	LUT3 #(
		.INIT('h2a)
	) name15693 (
		\m3_addr_i[10]_pad ,
		_w9069_,
		_w9070_,
		_w17594_
	);
	LUT3 #(
		.INIT('h80)
	) name15694 (
		\m4_addr_i[10]_pad ,
		_w9069_,
		_w9070_,
		_w17595_
	);
	LUT4 #(
		.INIT('h9dbf)
	) name15695 (
		_w9064_,
		_w9067_,
		_w17594_,
		_w17595_,
		_w17596_
	);
	LUT3 #(
		.INIT('h80)
	) name15696 (
		\m6_addr_i[10]_pad ,
		_w9069_,
		_w9070_,
		_w17597_
	);
	LUT3 #(
		.INIT('h80)
	) name15697 (
		\m2_addr_i[10]_pad ,
		_w9069_,
		_w9070_,
		_w17598_
	);
	LUT4 #(
		.INIT('habef)
	) name15698 (
		_w9064_,
		_w9067_,
		_w17597_,
		_w17598_,
		_w17599_
	);
	LUT3 #(
		.INIT('h2a)
	) name15699 (
		\m5_addr_i[10]_pad ,
		_w9069_,
		_w9070_,
		_w17600_
	);
	LUT3 #(
		.INIT('h2a)
	) name15700 (
		\m1_addr_i[10]_pad ,
		_w9069_,
		_w9070_,
		_w17601_
	);
	LUT4 #(
		.INIT('h57df)
	) name15701 (
		_w9064_,
		_w9067_,
		_w17600_,
		_w17601_,
		_w17602_
	);
	LUT3 #(
		.INIT('h80)
	) name15702 (
		\m0_addr_i[10]_pad ,
		_w9069_,
		_w9070_,
		_w17603_
	);
	LUT3 #(
		.INIT('h2a)
	) name15703 (
		\m7_addr_i[10]_pad ,
		_w9069_,
		_w9070_,
		_w17604_
	);
	LUT4 #(
		.INIT('h6e7f)
	) name15704 (
		_w9064_,
		_w9067_,
		_w17603_,
		_w17604_,
		_w17605_
	);
	LUT4 #(
		.INIT('h7fff)
	) name15705 (
		_w17596_,
		_w17599_,
		_w17602_,
		_w17605_,
		_w17606_
	);
	LUT3 #(
		.INIT('h2a)
	) name15706 (
		\m3_addr_i[11]_pad ,
		_w9069_,
		_w9070_,
		_w17607_
	);
	LUT3 #(
		.INIT('h80)
	) name15707 (
		\m4_addr_i[11]_pad ,
		_w9069_,
		_w9070_,
		_w17608_
	);
	LUT4 #(
		.INIT('h9dbf)
	) name15708 (
		_w9064_,
		_w9067_,
		_w17607_,
		_w17608_,
		_w17609_
	);
	LUT3 #(
		.INIT('h80)
	) name15709 (
		\m6_addr_i[11]_pad ,
		_w9069_,
		_w9070_,
		_w17610_
	);
	LUT3 #(
		.INIT('h80)
	) name15710 (
		\m2_addr_i[11]_pad ,
		_w9069_,
		_w9070_,
		_w17611_
	);
	LUT4 #(
		.INIT('habef)
	) name15711 (
		_w9064_,
		_w9067_,
		_w17610_,
		_w17611_,
		_w17612_
	);
	LUT3 #(
		.INIT('h2a)
	) name15712 (
		\m5_addr_i[11]_pad ,
		_w9069_,
		_w9070_,
		_w17613_
	);
	LUT3 #(
		.INIT('h2a)
	) name15713 (
		\m1_addr_i[11]_pad ,
		_w9069_,
		_w9070_,
		_w17614_
	);
	LUT4 #(
		.INIT('h57df)
	) name15714 (
		_w9064_,
		_w9067_,
		_w17613_,
		_w17614_,
		_w17615_
	);
	LUT3 #(
		.INIT('h80)
	) name15715 (
		\m0_addr_i[11]_pad ,
		_w9069_,
		_w9070_,
		_w17616_
	);
	LUT3 #(
		.INIT('h2a)
	) name15716 (
		\m7_addr_i[11]_pad ,
		_w9069_,
		_w9070_,
		_w17617_
	);
	LUT4 #(
		.INIT('h6e7f)
	) name15717 (
		_w9064_,
		_w9067_,
		_w17616_,
		_w17617_,
		_w17618_
	);
	LUT4 #(
		.INIT('h7fff)
	) name15718 (
		_w17609_,
		_w17612_,
		_w17615_,
		_w17618_,
		_w17619_
	);
	LUT3 #(
		.INIT('h2a)
	) name15719 (
		\m3_addr_i[12]_pad ,
		_w9069_,
		_w9070_,
		_w17620_
	);
	LUT3 #(
		.INIT('h80)
	) name15720 (
		\m4_addr_i[12]_pad ,
		_w9069_,
		_w9070_,
		_w17621_
	);
	LUT4 #(
		.INIT('h9dbf)
	) name15721 (
		_w9064_,
		_w9067_,
		_w17620_,
		_w17621_,
		_w17622_
	);
	LUT3 #(
		.INIT('h80)
	) name15722 (
		\m6_addr_i[12]_pad ,
		_w9069_,
		_w9070_,
		_w17623_
	);
	LUT3 #(
		.INIT('h80)
	) name15723 (
		\m2_addr_i[12]_pad ,
		_w9069_,
		_w9070_,
		_w17624_
	);
	LUT4 #(
		.INIT('habef)
	) name15724 (
		_w9064_,
		_w9067_,
		_w17623_,
		_w17624_,
		_w17625_
	);
	LUT3 #(
		.INIT('h2a)
	) name15725 (
		\m5_addr_i[12]_pad ,
		_w9069_,
		_w9070_,
		_w17626_
	);
	LUT3 #(
		.INIT('h2a)
	) name15726 (
		\m1_addr_i[12]_pad ,
		_w9069_,
		_w9070_,
		_w17627_
	);
	LUT4 #(
		.INIT('h57df)
	) name15727 (
		_w9064_,
		_w9067_,
		_w17626_,
		_w17627_,
		_w17628_
	);
	LUT3 #(
		.INIT('h80)
	) name15728 (
		\m0_addr_i[12]_pad ,
		_w9069_,
		_w9070_,
		_w17629_
	);
	LUT3 #(
		.INIT('h2a)
	) name15729 (
		\m7_addr_i[12]_pad ,
		_w9069_,
		_w9070_,
		_w17630_
	);
	LUT4 #(
		.INIT('h6e7f)
	) name15730 (
		_w9064_,
		_w9067_,
		_w17629_,
		_w17630_,
		_w17631_
	);
	LUT4 #(
		.INIT('h7fff)
	) name15731 (
		_w17622_,
		_w17625_,
		_w17628_,
		_w17631_,
		_w17632_
	);
	LUT3 #(
		.INIT('h2a)
	) name15732 (
		\m3_addr_i[13]_pad ,
		_w9069_,
		_w9070_,
		_w17633_
	);
	LUT3 #(
		.INIT('h80)
	) name15733 (
		\m4_addr_i[13]_pad ,
		_w9069_,
		_w9070_,
		_w17634_
	);
	LUT4 #(
		.INIT('h9dbf)
	) name15734 (
		_w9064_,
		_w9067_,
		_w17633_,
		_w17634_,
		_w17635_
	);
	LUT3 #(
		.INIT('h80)
	) name15735 (
		\m6_addr_i[13]_pad ,
		_w9069_,
		_w9070_,
		_w17636_
	);
	LUT3 #(
		.INIT('h80)
	) name15736 (
		\m2_addr_i[13]_pad ,
		_w9069_,
		_w9070_,
		_w17637_
	);
	LUT4 #(
		.INIT('habef)
	) name15737 (
		_w9064_,
		_w9067_,
		_w17636_,
		_w17637_,
		_w17638_
	);
	LUT3 #(
		.INIT('h2a)
	) name15738 (
		\m5_addr_i[13]_pad ,
		_w9069_,
		_w9070_,
		_w17639_
	);
	LUT3 #(
		.INIT('h2a)
	) name15739 (
		\m1_addr_i[13]_pad ,
		_w9069_,
		_w9070_,
		_w17640_
	);
	LUT4 #(
		.INIT('h57df)
	) name15740 (
		_w9064_,
		_w9067_,
		_w17639_,
		_w17640_,
		_w17641_
	);
	LUT3 #(
		.INIT('h80)
	) name15741 (
		\m0_addr_i[13]_pad ,
		_w9069_,
		_w9070_,
		_w17642_
	);
	LUT3 #(
		.INIT('h2a)
	) name15742 (
		\m7_addr_i[13]_pad ,
		_w9069_,
		_w9070_,
		_w17643_
	);
	LUT4 #(
		.INIT('h6e7f)
	) name15743 (
		_w9064_,
		_w9067_,
		_w17642_,
		_w17643_,
		_w17644_
	);
	LUT4 #(
		.INIT('h7fff)
	) name15744 (
		_w17635_,
		_w17638_,
		_w17641_,
		_w17644_,
		_w17645_
	);
	LUT3 #(
		.INIT('h2a)
	) name15745 (
		\m3_addr_i[14]_pad ,
		_w9069_,
		_w9070_,
		_w17646_
	);
	LUT3 #(
		.INIT('h80)
	) name15746 (
		\m4_addr_i[14]_pad ,
		_w9069_,
		_w9070_,
		_w17647_
	);
	LUT4 #(
		.INIT('h9dbf)
	) name15747 (
		_w9064_,
		_w9067_,
		_w17646_,
		_w17647_,
		_w17648_
	);
	LUT3 #(
		.INIT('h80)
	) name15748 (
		\m6_addr_i[14]_pad ,
		_w9069_,
		_w9070_,
		_w17649_
	);
	LUT3 #(
		.INIT('h80)
	) name15749 (
		\m2_addr_i[14]_pad ,
		_w9069_,
		_w9070_,
		_w17650_
	);
	LUT4 #(
		.INIT('habef)
	) name15750 (
		_w9064_,
		_w9067_,
		_w17649_,
		_w17650_,
		_w17651_
	);
	LUT3 #(
		.INIT('h2a)
	) name15751 (
		\m5_addr_i[14]_pad ,
		_w9069_,
		_w9070_,
		_w17652_
	);
	LUT3 #(
		.INIT('h2a)
	) name15752 (
		\m1_addr_i[14]_pad ,
		_w9069_,
		_w9070_,
		_w17653_
	);
	LUT4 #(
		.INIT('h57df)
	) name15753 (
		_w9064_,
		_w9067_,
		_w17652_,
		_w17653_,
		_w17654_
	);
	LUT3 #(
		.INIT('h80)
	) name15754 (
		\m0_addr_i[14]_pad ,
		_w9069_,
		_w9070_,
		_w17655_
	);
	LUT3 #(
		.INIT('h2a)
	) name15755 (
		\m7_addr_i[14]_pad ,
		_w9069_,
		_w9070_,
		_w17656_
	);
	LUT4 #(
		.INIT('h6e7f)
	) name15756 (
		_w9064_,
		_w9067_,
		_w17655_,
		_w17656_,
		_w17657_
	);
	LUT4 #(
		.INIT('h7fff)
	) name15757 (
		_w17648_,
		_w17651_,
		_w17654_,
		_w17657_,
		_w17658_
	);
	LUT3 #(
		.INIT('h2a)
	) name15758 (
		\m3_addr_i[15]_pad ,
		_w9069_,
		_w9070_,
		_w17659_
	);
	LUT3 #(
		.INIT('h80)
	) name15759 (
		\m4_addr_i[15]_pad ,
		_w9069_,
		_w9070_,
		_w17660_
	);
	LUT4 #(
		.INIT('h9dbf)
	) name15760 (
		_w9064_,
		_w9067_,
		_w17659_,
		_w17660_,
		_w17661_
	);
	LUT3 #(
		.INIT('h80)
	) name15761 (
		\m6_addr_i[15]_pad ,
		_w9069_,
		_w9070_,
		_w17662_
	);
	LUT3 #(
		.INIT('h80)
	) name15762 (
		\m2_addr_i[15]_pad ,
		_w9069_,
		_w9070_,
		_w17663_
	);
	LUT4 #(
		.INIT('habef)
	) name15763 (
		_w9064_,
		_w9067_,
		_w17662_,
		_w17663_,
		_w17664_
	);
	LUT3 #(
		.INIT('h2a)
	) name15764 (
		\m5_addr_i[15]_pad ,
		_w9069_,
		_w9070_,
		_w17665_
	);
	LUT3 #(
		.INIT('h2a)
	) name15765 (
		\m1_addr_i[15]_pad ,
		_w9069_,
		_w9070_,
		_w17666_
	);
	LUT4 #(
		.INIT('h57df)
	) name15766 (
		_w9064_,
		_w9067_,
		_w17665_,
		_w17666_,
		_w17667_
	);
	LUT3 #(
		.INIT('h80)
	) name15767 (
		\m0_addr_i[15]_pad ,
		_w9069_,
		_w9070_,
		_w17668_
	);
	LUT3 #(
		.INIT('h2a)
	) name15768 (
		\m7_addr_i[15]_pad ,
		_w9069_,
		_w9070_,
		_w17669_
	);
	LUT4 #(
		.INIT('h6e7f)
	) name15769 (
		_w9064_,
		_w9067_,
		_w17668_,
		_w17669_,
		_w17670_
	);
	LUT4 #(
		.INIT('h7fff)
	) name15770 (
		_w17661_,
		_w17664_,
		_w17667_,
		_w17670_,
		_w17671_
	);
	LUT3 #(
		.INIT('h2a)
	) name15771 (
		\m3_addr_i[16]_pad ,
		_w9069_,
		_w9070_,
		_w17672_
	);
	LUT3 #(
		.INIT('h80)
	) name15772 (
		\m4_addr_i[16]_pad ,
		_w9069_,
		_w9070_,
		_w17673_
	);
	LUT4 #(
		.INIT('h9dbf)
	) name15773 (
		_w9064_,
		_w9067_,
		_w17672_,
		_w17673_,
		_w17674_
	);
	LUT3 #(
		.INIT('h80)
	) name15774 (
		\m6_addr_i[16]_pad ,
		_w9069_,
		_w9070_,
		_w17675_
	);
	LUT3 #(
		.INIT('h80)
	) name15775 (
		\m2_addr_i[16]_pad ,
		_w9069_,
		_w9070_,
		_w17676_
	);
	LUT4 #(
		.INIT('habef)
	) name15776 (
		_w9064_,
		_w9067_,
		_w17675_,
		_w17676_,
		_w17677_
	);
	LUT3 #(
		.INIT('h2a)
	) name15777 (
		\m5_addr_i[16]_pad ,
		_w9069_,
		_w9070_,
		_w17678_
	);
	LUT3 #(
		.INIT('h2a)
	) name15778 (
		\m1_addr_i[16]_pad ,
		_w9069_,
		_w9070_,
		_w17679_
	);
	LUT4 #(
		.INIT('h57df)
	) name15779 (
		_w9064_,
		_w9067_,
		_w17678_,
		_w17679_,
		_w17680_
	);
	LUT3 #(
		.INIT('h80)
	) name15780 (
		\m0_addr_i[16]_pad ,
		_w9069_,
		_w9070_,
		_w17681_
	);
	LUT3 #(
		.INIT('h2a)
	) name15781 (
		\m7_addr_i[16]_pad ,
		_w9069_,
		_w9070_,
		_w17682_
	);
	LUT4 #(
		.INIT('h6e7f)
	) name15782 (
		_w9064_,
		_w9067_,
		_w17681_,
		_w17682_,
		_w17683_
	);
	LUT4 #(
		.INIT('h7fff)
	) name15783 (
		_w17674_,
		_w17677_,
		_w17680_,
		_w17683_,
		_w17684_
	);
	LUT3 #(
		.INIT('h2a)
	) name15784 (
		\m3_addr_i[17]_pad ,
		_w9069_,
		_w9070_,
		_w17685_
	);
	LUT3 #(
		.INIT('h80)
	) name15785 (
		\m4_addr_i[17]_pad ,
		_w9069_,
		_w9070_,
		_w17686_
	);
	LUT4 #(
		.INIT('h9dbf)
	) name15786 (
		_w9064_,
		_w9067_,
		_w17685_,
		_w17686_,
		_w17687_
	);
	LUT3 #(
		.INIT('h80)
	) name15787 (
		\m6_addr_i[17]_pad ,
		_w9069_,
		_w9070_,
		_w17688_
	);
	LUT3 #(
		.INIT('h80)
	) name15788 (
		\m2_addr_i[17]_pad ,
		_w9069_,
		_w9070_,
		_w17689_
	);
	LUT4 #(
		.INIT('habef)
	) name15789 (
		_w9064_,
		_w9067_,
		_w17688_,
		_w17689_,
		_w17690_
	);
	LUT3 #(
		.INIT('h2a)
	) name15790 (
		\m5_addr_i[17]_pad ,
		_w9069_,
		_w9070_,
		_w17691_
	);
	LUT3 #(
		.INIT('h2a)
	) name15791 (
		\m1_addr_i[17]_pad ,
		_w9069_,
		_w9070_,
		_w17692_
	);
	LUT4 #(
		.INIT('h57df)
	) name15792 (
		_w9064_,
		_w9067_,
		_w17691_,
		_w17692_,
		_w17693_
	);
	LUT3 #(
		.INIT('h80)
	) name15793 (
		\m0_addr_i[17]_pad ,
		_w9069_,
		_w9070_,
		_w17694_
	);
	LUT3 #(
		.INIT('h2a)
	) name15794 (
		\m7_addr_i[17]_pad ,
		_w9069_,
		_w9070_,
		_w17695_
	);
	LUT4 #(
		.INIT('h6e7f)
	) name15795 (
		_w9064_,
		_w9067_,
		_w17694_,
		_w17695_,
		_w17696_
	);
	LUT4 #(
		.INIT('h7fff)
	) name15796 (
		_w17687_,
		_w17690_,
		_w17693_,
		_w17696_,
		_w17697_
	);
	LUT3 #(
		.INIT('h2a)
	) name15797 (
		\m3_addr_i[18]_pad ,
		_w9069_,
		_w9070_,
		_w17698_
	);
	LUT3 #(
		.INIT('h80)
	) name15798 (
		\m4_addr_i[18]_pad ,
		_w9069_,
		_w9070_,
		_w17699_
	);
	LUT4 #(
		.INIT('h9dbf)
	) name15799 (
		_w9064_,
		_w9067_,
		_w17698_,
		_w17699_,
		_w17700_
	);
	LUT3 #(
		.INIT('h80)
	) name15800 (
		\m6_addr_i[18]_pad ,
		_w9069_,
		_w9070_,
		_w17701_
	);
	LUT3 #(
		.INIT('h80)
	) name15801 (
		\m2_addr_i[18]_pad ,
		_w9069_,
		_w9070_,
		_w17702_
	);
	LUT4 #(
		.INIT('habef)
	) name15802 (
		_w9064_,
		_w9067_,
		_w17701_,
		_w17702_,
		_w17703_
	);
	LUT3 #(
		.INIT('h2a)
	) name15803 (
		\m5_addr_i[18]_pad ,
		_w9069_,
		_w9070_,
		_w17704_
	);
	LUT3 #(
		.INIT('h2a)
	) name15804 (
		\m1_addr_i[18]_pad ,
		_w9069_,
		_w9070_,
		_w17705_
	);
	LUT4 #(
		.INIT('h57df)
	) name15805 (
		_w9064_,
		_w9067_,
		_w17704_,
		_w17705_,
		_w17706_
	);
	LUT3 #(
		.INIT('h80)
	) name15806 (
		\m0_addr_i[18]_pad ,
		_w9069_,
		_w9070_,
		_w17707_
	);
	LUT3 #(
		.INIT('h2a)
	) name15807 (
		\m7_addr_i[18]_pad ,
		_w9069_,
		_w9070_,
		_w17708_
	);
	LUT4 #(
		.INIT('h6e7f)
	) name15808 (
		_w9064_,
		_w9067_,
		_w17707_,
		_w17708_,
		_w17709_
	);
	LUT4 #(
		.INIT('h7fff)
	) name15809 (
		_w17700_,
		_w17703_,
		_w17706_,
		_w17709_,
		_w17710_
	);
	LUT3 #(
		.INIT('h2a)
	) name15810 (
		\m3_addr_i[19]_pad ,
		_w9069_,
		_w9070_,
		_w17711_
	);
	LUT3 #(
		.INIT('h80)
	) name15811 (
		\m4_addr_i[19]_pad ,
		_w9069_,
		_w9070_,
		_w17712_
	);
	LUT4 #(
		.INIT('h9dbf)
	) name15812 (
		_w9064_,
		_w9067_,
		_w17711_,
		_w17712_,
		_w17713_
	);
	LUT3 #(
		.INIT('h80)
	) name15813 (
		\m6_addr_i[19]_pad ,
		_w9069_,
		_w9070_,
		_w17714_
	);
	LUT3 #(
		.INIT('h80)
	) name15814 (
		\m2_addr_i[19]_pad ,
		_w9069_,
		_w9070_,
		_w17715_
	);
	LUT4 #(
		.INIT('habef)
	) name15815 (
		_w9064_,
		_w9067_,
		_w17714_,
		_w17715_,
		_w17716_
	);
	LUT3 #(
		.INIT('h2a)
	) name15816 (
		\m5_addr_i[19]_pad ,
		_w9069_,
		_w9070_,
		_w17717_
	);
	LUT3 #(
		.INIT('h2a)
	) name15817 (
		\m1_addr_i[19]_pad ,
		_w9069_,
		_w9070_,
		_w17718_
	);
	LUT4 #(
		.INIT('h57df)
	) name15818 (
		_w9064_,
		_w9067_,
		_w17717_,
		_w17718_,
		_w17719_
	);
	LUT3 #(
		.INIT('h80)
	) name15819 (
		\m0_addr_i[19]_pad ,
		_w9069_,
		_w9070_,
		_w17720_
	);
	LUT3 #(
		.INIT('h2a)
	) name15820 (
		\m7_addr_i[19]_pad ,
		_w9069_,
		_w9070_,
		_w17721_
	);
	LUT4 #(
		.INIT('h6e7f)
	) name15821 (
		_w9064_,
		_w9067_,
		_w17720_,
		_w17721_,
		_w17722_
	);
	LUT4 #(
		.INIT('h7fff)
	) name15822 (
		_w17713_,
		_w17716_,
		_w17719_,
		_w17722_,
		_w17723_
	);
	LUT3 #(
		.INIT('h2a)
	) name15823 (
		\m3_addr_i[1]_pad ,
		_w9069_,
		_w9070_,
		_w17724_
	);
	LUT3 #(
		.INIT('h80)
	) name15824 (
		\m4_addr_i[1]_pad ,
		_w9069_,
		_w9070_,
		_w17725_
	);
	LUT4 #(
		.INIT('h9dbf)
	) name15825 (
		_w9064_,
		_w9067_,
		_w17724_,
		_w17725_,
		_w17726_
	);
	LUT3 #(
		.INIT('h80)
	) name15826 (
		\m6_addr_i[1]_pad ,
		_w9069_,
		_w9070_,
		_w17727_
	);
	LUT3 #(
		.INIT('h80)
	) name15827 (
		\m2_addr_i[1]_pad ,
		_w9069_,
		_w9070_,
		_w17728_
	);
	LUT4 #(
		.INIT('habef)
	) name15828 (
		_w9064_,
		_w9067_,
		_w17727_,
		_w17728_,
		_w17729_
	);
	LUT3 #(
		.INIT('h2a)
	) name15829 (
		\m5_addr_i[1]_pad ,
		_w9069_,
		_w9070_,
		_w17730_
	);
	LUT3 #(
		.INIT('h2a)
	) name15830 (
		\m1_addr_i[1]_pad ,
		_w9069_,
		_w9070_,
		_w17731_
	);
	LUT4 #(
		.INIT('h57df)
	) name15831 (
		_w9064_,
		_w9067_,
		_w17730_,
		_w17731_,
		_w17732_
	);
	LUT3 #(
		.INIT('h80)
	) name15832 (
		\m0_addr_i[1]_pad ,
		_w9069_,
		_w9070_,
		_w17733_
	);
	LUT3 #(
		.INIT('h2a)
	) name15833 (
		\m7_addr_i[1]_pad ,
		_w9069_,
		_w9070_,
		_w17734_
	);
	LUT4 #(
		.INIT('h6e7f)
	) name15834 (
		_w9064_,
		_w9067_,
		_w17733_,
		_w17734_,
		_w17735_
	);
	LUT4 #(
		.INIT('h7fff)
	) name15835 (
		_w17726_,
		_w17729_,
		_w17732_,
		_w17735_,
		_w17736_
	);
	LUT3 #(
		.INIT('h2a)
	) name15836 (
		\m3_addr_i[20]_pad ,
		_w9069_,
		_w9070_,
		_w17737_
	);
	LUT3 #(
		.INIT('h80)
	) name15837 (
		\m4_addr_i[20]_pad ,
		_w9069_,
		_w9070_,
		_w17738_
	);
	LUT4 #(
		.INIT('h9dbf)
	) name15838 (
		_w9064_,
		_w9067_,
		_w17737_,
		_w17738_,
		_w17739_
	);
	LUT3 #(
		.INIT('h80)
	) name15839 (
		\m6_addr_i[20]_pad ,
		_w9069_,
		_w9070_,
		_w17740_
	);
	LUT3 #(
		.INIT('h80)
	) name15840 (
		\m2_addr_i[20]_pad ,
		_w9069_,
		_w9070_,
		_w17741_
	);
	LUT4 #(
		.INIT('habef)
	) name15841 (
		_w9064_,
		_w9067_,
		_w17740_,
		_w17741_,
		_w17742_
	);
	LUT3 #(
		.INIT('h2a)
	) name15842 (
		\m5_addr_i[20]_pad ,
		_w9069_,
		_w9070_,
		_w17743_
	);
	LUT3 #(
		.INIT('h2a)
	) name15843 (
		\m1_addr_i[20]_pad ,
		_w9069_,
		_w9070_,
		_w17744_
	);
	LUT4 #(
		.INIT('h57df)
	) name15844 (
		_w9064_,
		_w9067_,
		_w17743_,
		_w17744_,
		_w17745_
	);
	LUT3 #(
		.INIT('h80)
	) name15845 (
		\m0_addr_i[20]_pad ,
		_w9069_,
		_w9070_,
		_w17746_
	);
	LUT3 #(
		.INIT('h2a)
	) name15846 (
		\m7_addr_i[20]_pad ,
		_w9069_,
		_w9070_,
		_w17747_
	);
	LUT4 #(
		.INIT('h6e7f)
	) name15847 (
		_w9064_,
		_w9067_,
		_w17746_,
		_w17747_,
		_w17748_
	);
	LUT4 #(
		.INIT('h7fff)
	) name15848 (
		_w17739_,
		_w17742_,
		_w17745_,
		_w17748_,
		_w17749_
	);
	LUT3 #(
		.INIT('h2a)
	) name15849 (
		\m3_addr_i[21]_pad ,
		_w9069_,
		_w9070_,
		_w17750_
	);
	LUT3 #(
		.INIT('h80)
	) name15850 (
		\m4_addr_i[21]_pad ,
		_w9069_,
		_w9070_,
		_w17751_
	);
	LUT4 #(
		.INIT('h9dbf)
	) name15851 (
		_w9064_,
		_w9067_,
		_w17750_,
		_w17751_,
		_w17752_
	);
	LUT3 #(
		.INIT('h80)
	) name15852 (
		\m6_addr_i[21]_pad ,
		_w9069_,
		_w9070_,
		_w17753_
	);
	LUT3 #(
		.INIT('h80)
	) name15853 (
		\m2_addr_i[21]_pad ,
		_w9069_,
		_w9070_,
		_w17754_
	);
	LUT4 #(
		.INIT('habef)
	) name15854 (
		_w9064_,
		_w9067_,
		_w17753_,
		_w17754_,
		_w17755_
	);
	LUT3 #(
		.INIT('h2a)
	) name15855 (
		\m5_addr_i[21]_pad ,
		_w9069_,
		_w9070_,
		_w17756_
	);
	LUT3 #(
		.INIT('h2a)
	) name15856 (
		\m1_addr_i[21]_pad ,
		_w9069_,
		_w9070_,
		_w17757_
	);
	LUT4 #(
		.INIT('h57df)
	) name15857 (
		_w9064_,
		_w9067_,
		_w17756_,
		_w17757_,
		_w17758_
	);
	LUT3 #(
		.INIT('h80)
	) name15858 (
		\m0_addr_i[21]_pad ,
		_w9069_,
		_w9070_,
		_w17759_
	);
	LUT3 #(
		.INIT('h2a)
	) name15859 (
		\m7_addr_i[21]_pad ,
		_w9069_,
		_w9070_,
		_w17760_
	);
	LUT4 #(
		.INIT('h6e7f)
	) name15860 (
		_w9064_,
		_w9067_,
		_w17759_,
		_w17760_,
		_w17761_
	);
	LUT4 #(
		.INIT('h7fff)
	) name15861 (
		_w17752_,
		_w17755_,
		_w17758_,
		_w17761_,
		_w17762_
	);
	LUT3 #(
		.INIT('h2a)
	) name15862 (
		\m3_addr_i[22]_pad ,
		_w9069_,
		_w9070_,
		_w17763_
	);
	LUT3 #(
		.INIT('h80)
	) name15863 (
		\m4_addr_i[22]_pad ,
		_w9069_,
		_w9070_,
		_w17764_
	);
	LUT4 #(
		.INIT('h9dbf)
	) name15864 (
		_w9064_,
		_w9067_,
		_w17763_,
		_w17764_,
		_w17765_
	);
	LUT3 #(
		.INIT('h80)
	) name15865 (
		\m6_addr_i[22]_pad ,
		_w9069_,
		_w9070_,
		_w17766_
	);
	LUT3 #(
		.INIT('h80)
	) name15866 (
		\m2_addr_i[22]_pad ,
		_w9069_,
		_w9070_,
		_w17767_
	);
	LUT4 #(
		.INIT('habef)
	) name15867 (
		_w9064_,
		_w9067_,
		_w17766_,
		_w17767_,
		_w17768_
	);
	LUT3 #(
		.INIT('h2a)
	) name15868 (
		\m5_addr_i[22]_pad ,
		_w9069_,
		_w9070_,
		_w17769_
	);
	LUT3 #(
		.INIT('h2a)
	) name15869 (
		\m1_addr_i[22]_pad ,
		_w9069_,
		_w9070_,
		_w17770_
	);
	LUT4 #(
		.INIT('h57df)
	) name15870 (
		_w9064_,
		_w9067_,
		_w17769_,
		_w17770_,
		_w17771_
	);
	LUT3 #(
		.INIT('h80)
	) name15871 (
		\m0_addr_i[22]_pad ,
		_w9069_,
		_w9070_,
		_w17772_
	);
	LUT3 #(
		.INIT('h2a)
	) name15872 (
		\m7_addr_i[22]_pad ,
		_w9069_,
		_w9070_,
		_w17773_
	);
	LUT4 #(
		.INIT('h6e7f)
	) name15873 (
		_w9064_,
		_w9067_,
		_w17772_,
		_w17773_,
		_w17774_
	);
	LUT4 #(
		.INIT('h7fff)
	) name15874 (
		_w17765_,
		_w17768_,
		_w17771_,
		_w17774_,
		_w17775_
	);
	LUT3 #(
		.INIT('h2a)
	) name15875 (
		\m3_addr_i[23]_pad ,
		_w9069_,
		_w9070_,
		_w17776_
	);
	LUT3 #(
		.INIT('h80)
	) name15876 (
		\m4_addr_i[23]_pad ,
		_w9069_,
		_w9070_,
		_w17777_
	);
	LUT4 #(
		.INIT('h9dbf)
	) name15877 (
		_w9064_,
		_w9067_,
		_w17776_,
		_w17777_,
		_w17778_
	);
	LUT3 #(
		.INIT('h80)
	) name15878 (
		\m6_addr_i[23]_pad ,
		_w9069_,
		_w9070_,
		_w17779_
	);
	LUT3 #(
		.INIT('h80)
	) name15879 (
		\m2_addr_i[23]_pad ,
		_w9069_,
		_w9070_,
		_w17780_
	);
	LUT4 #(
		.INIT('habef)
	) name15880 (
		_w9064_,
		_w9067_,
		_w17779_,
		_w17780_,
		_w17781_
	);
	LUT3 #(
		.INIT('h2a)
	) name15881 (
		\m5_addr_i[23]_pad ,
		_w9069_,
		_w9070_,
		_w17782_
	);
	LUT3 #(
		.INIT('h2a)
	) name15882 (
		\m1_addr_i[23]_pad ,
		_w9069_,
		_w9070_,
		_w17783_
	);
	LUT4 #(
		.INIT('h57df)
	) name15883 (
		_w9064_,
		_w9067_,
		_w17782_,
		_w17783_,
		_w17784_
	);
	LUT3 #(
		.INIT('h80)
	) name15884 (
		\m0_addr_i[23]_pad ,
		_w9069_,
		_w9070_,
		_w17785_
	);
	LUT3 #(
		.INIT('h2a)
	) name15885 (
		\m7_addr_i[23]_pad ,
		_w9069_,
		_w9070_,
		_w17786_
	);
	LUT4 #(
		.INIT('h6e7f)
	) name15886 (
		_w9064_,
		_w9067_,
		_w17785_,
		_w17786_,
		_w17787_
	);
	LUT4 #(
		.INIT('h7fff)
	) name15887 (
		_w17778_,
		_w17781_,
		_w17784_,
		_w17787_,
		_w17788_
	);
	LUT3 #(
		.INIT('h2a)
	) name15888 (
		\m3_addr_i[24]_pad ,
		_w9069_,
		_w9070_,
		_w17789_
	);
	LUT3 #(
		.INIT('h80)
	) name15889 (
		\m4_addr_i[24]_pad ,
		_w9069_,
		_w9070_,
		_w17790_
	);
	LUT4 #(
		.INIT('h9dbf)
	) name15890 (
		_w9064_,
		_w9067_,
		_w17789_,
		_w17790_,
		_w17791_
	);
	LUT3 #(
		.INIT('h2a)
	) name15891 (
		\m5_addr_i[24]_pad ,
		_w9069_,
		_w9070_,
		_w17792_
	);
	LUT3 #(
		.INIT('h80)
	) name15892 (
		\m2_addr_i[24]_pad ,
		_w9069_,
		_w9070_,
		_w17793_
	);
	LUT4 #(
		.INIT('h9bdf)
	) name15893 (
		_w9064_,
		_w9067_,
		_w17792_,
		_w17793_,
		_w17794_
	);
	LUT3 #(
		.INIT('h80)
	) name15894 (
		\m6_addr_i[24]_pad ,
		_w9069_,
		_w9070_,
		_w17795_
	);
	LUT3 #(
		.INIT('h2a)
	) name15895 (
		\m1_addr_i[24]_pad ,
		_w9069_,
		_w9070_,
		_w17796_
	);
	LUT4 #(
		.INIT('h67ef)
	) name15896 (
		_w9064_,
		_w9067_,
		_w17795_,
		_w17796_,
		_w17797_
	);
	LUT3 #(
		.INIT('h80)
	) name15897 (
		\m0_addr_i[24]_pad ,
		_w9069_,
		_w9070_,
		_w17798_
	);
	LUT3 #(
		.INIT('h2a)
	) name15898 (
		\m7_addr_i[24]_pad ,
		_w9069_,
		_w9070_,
		_w17799_
	);
	LUT4 #(
		.INIT('h6e7f)
	) name15899 (
		_w9064_,
		_w9067_,
		_w17798_,
		_w17799_,
		_w17800_
	);
	LUT4 #(
		.INIT('h7fff)
	) name15900 (
		_w17791_,
		_w17794_,
		_w17797_,
		_w17800_,
		_w17801_
	);
	LUT3 #(
		.INIT('h2a)
	) name15901 (
		\m3_addr_i[25]_pad ,
		_w9069_,
		_w9070_,
		_w17802_
	);
	LUT3 #(
		.INIT('h80)
	) name15902 (
		\m4_addr_i[25]_pad ,
		_w9069_,
		_w9070_,
		_w17803_
	);
	LUT4 #(
		.INIT('h9dbf)
	) name15903 (
		_w9064_,
		_w9067_,
		_w17802_,
		_w17803_,
		_w17804_
	);
	LUT3 #(
		.INIT('h2a)
	) name15904 (
		\m5_addr_i[25]_pad ,
		_w9069_,
		_w9070_,
		_w17805_
	);
	LUT3 #(
		.INIT('h80)
	) name15905 (
		\m2_addr_i[25]_pad ,
		_w9069_,
		_w9070_,
		_w17806_
	);
	LUT4 #(
		.INIT('h9bdf)
	) name15906 (
		_w9064_,
		_w9067_,
		_w17805_,
		_w17806_,
		_w17807_
	);
	LUT3 #(
		.INIT('h80)
	) name15907 (
		\m6_addr_i[25]_pad ,
		_w9069_,
		_w9070_,
		_w17808_
	);
	LUT3 #(
		.INIT('h2a)
	) name15908 (
		\m1_addr_i[25]_pad ,
		_w9069_,
		_w9070_,
		_w17809_
	);
	LUT4 #(
		.INIT('h67ef)
	) name15909 (
		_w9064_,
		_w9067_,
		_w17808_,
		_w17809_,
		_w17810_
	);
	LUT3 #(
		.INIT('h80)
	) name15910 (
		\m0_addr_i[25]_pad ,
		_w9069_,
		_w9070_,
		_w17811_
	);
	LUT3 #(
		.INIT('h2a)
	) name15911 (
		\m7_addr_i[25]_pad ,
		_w9069_,
		_w9070_,
		_w17812_
	);
	LUT4 #(
		.INIT('h6e7f)
	) name15912 (
		_w9064_,
		_w9067_,
		_w17811_,
		_w17812_,
		_w17813_
	);
	LUT4 #(
		.INIT('h7fff)
	) name15913 (
		_w17804_,
		_w17807_,
		_w17810_,
		_w17813_,
		_w17814_
	);
	LUT3 #(
		.INIT('h2a)
	) name15914 (
		\m3_addr_i[26]_pad ,
		_w9069_,
		_w9070_,
		_w17815_
	);
	LUT3 #(
		.INIT('h80)
	) name15915 (
		\m4_addr_i[26]_pad ,
		_w9069_,
		_w9070_,
		_w17816_
	);
	LUT4 #(
		.INIT('h9dbf)
	) name15916 (
		_w9064_,
		_w9067_,
		_w17815_,
		_w17816_,
		_w17817_
	);
	LUT3 #(
		.INIT('h2a)
	) name15917 (
		\m5_addr_i[26]_pad ,
		_w9069_,
		_w9070_,
		_w17818_
	);
	LUT3 #(
		.INIT('h80)
	) name15918 (
		\m2_addr_i[26]_pad ,
		_w9069_,
		_w9070_,
		_w17819_
	);
	LUT4 #(
		.INIT('h9bdf)
	) name15919 (
		_w9064_,
		_w9067_,
		_w17818_,
		_w17819_,
		_w17820_
	);
	LUT3 #(
		.INIT('h80)
	) name15920 (
		\m6_addr_i[26]_pad ,
		_w9069_,
		_w9070_,
		_w17821_
	);
	LUT3 #(
		.INIT('h2a)
	) name15921 (
		\m1_addr_i[26]_pad ,
		_w9069_,
		_w9070_,
		_w17822_
	);
	LUT4 #(
		.INIT('h67ef)
	) name15922 (
		_w9064_,
		_w9067_,
		_w17821_,
		_w17822_,
		_w17823_
	);
	LUT3 #(
		.INIT('h80)
	) name15923 (
		\m0_addr_i[26]_pad ,
		_w9069_,
		_w9070_,
		_w17824_
	);
	LUT3 #(
		.INIT('h2a)
	) name15924 (
		\m7_addr_i[26]_pad ,
		_w9069_,
		_w9070_,
		_w17825_
	);
	LUT4 #(
		.INIT('h6e7f)
	) name15925 (
		_w9064_,
		_w9067_,
		_w17824_,
		_w17825_,
		_w17826_
	);
	LUT4 #(
		.INIT('h7fff)
	) name15926 (
		_w17817_,
		_w17820_,
		_w17823_,
		_w17826_,
		_w17827_
	);
	LUT3 #(
		.INIT('h2a)
	) name15927 (
		\m3_addr_i[27]_pad ,
		_w9069_,
		_w9070_,
		_w17828_
	);
	LUT3 #(
		.INIT('h80)
	) name15928 (
		\m4_addr_i[27]_pad ,
		_w9069_,
		_w9070_,
		_w17829_
	);
	LUT4 #(
		.INIT('h9dbf)
	) name15929 (
		_w9064_,
		_w9067_,
		_w17828_,
		_w17829_,
		_w17830_
	);
	LUT3 #(
		.INIT('h2a)
	) name15930 (
		\m5_addr_i[27]_pad ,
		_w9069_,
		_w9070_,
		_w17831_
	);
	LUT3 #(
		.INIT('h80)
	) name15931 (
		\m2_addr_i[27]_pad ,
		_w9069_,
		_w9070_,
		_w17832_
	);
	LUT4 #(
		.INIT('h9bdf)
	) name15932 (
		_w9064_,
		_w9067_,
		_w17831_,
		_w17832_,
		_w17833_
	);
	LUT3 #(
		.INIT('h80)
	) name15933 (
		\m6_addr_i[27]_pad ,
		_w9069_,
		_w9070_,
		_w17834_
	);
	LUT3 #(
		.INIT('h2a)
	) name15934 (
		\m1_addr_i[27]_pad ,
		_w9069_,
		_w9070_,
		_w17835_
	);
	LUT4 #(
		.INIT('h67ef)
	) name15935 (
		_w9064_,
		_w9067_,
		_w17834_,
		_w17835_,
		_w17836_
	);
	LUT3 #(
		.INIT('h80)
	) name15936 (
		\m0_addr_i[27]_pad ,
		_w9069_,
		_w9070_,
		_w17837_
	);
	LUT3 #(
		.INIT('h2a)
	) name15937 (
		\m7_addr_i[27]_pad ,
		_w9069_,
		_w9070_,
		_w17838_
	);
	LUT4 #(
		.INIT('h6e7f)
	) name15938 (
		_w9064_,
		_w9067_,
		_w17837_,
		_w17838_,
		_w17839_
	);
	LUT4 #(
		.INIT('h7fff)
	) name15939 (
		_w17830_,
		_w17833_,
		_w17836_,
		_w17839_,
		_w17840_
	);
	LUT3 #(
		.INIT('h2a)
	) name15940 (
		\m3_addr_i[28]_pad ,
		_w9069_,
		_w9070_,
		_w17841_
	);
	LUT3 #(
		.INIT('h80)
	) name15941 (
		\m4_addr_i[28]_pad ,
		_w9069_,
		_w9070_,
		_w17842_
	);
	LUT4 #(
		.INIT('h9dbf)
	) name15942 (
		_w9064_,
		_w9067_,
		_w17841_,
		_w17842_,
		_w17843_
	);
	LUT3 #(
		.INIT('h2a)
	) name15943 (
		\m5_addr_i[28]_pad ,
		_w9069_,
		_w9070_,
		_w17844_
	);
	LUT3 #(
		.INIT('h80)
	) name15944 (
		\m2_addr_i[28]_pad ,
		_w9069_,
		_w9070_,
		_w17845_
	);
	LUT4 #(
		.INIT('h9bdf)
	) name15945 (
		_w9064_,
		_w9067_,
		_w17844_,
		_w17845_,
		_w17846_
	);
	LUT3 #(
		.INIT('h80)
	) name15946 (
		\m6_addr_i[28]_pad ,
		_w9069_,
		_w9070_,
		_w17847_
	);
	LUT3 #(
		.INIT('h2a)
	) name15947 (
		\m1_addr_i[28]_pad ,
		_w9069_,
		_w9070_,
		_w17848_
	);
	LUT4 #(
		.INIT('h67ef)
	) name15948 (
		_w9064_,
		_w9067_,
		_w17847_,
		_w17848_,
		_w17849_
	);
	LUT3 #(
		.INIT('h80)
	) name15949 (
		\m0_addr_i[28]_pad ,
		_w9069_,
		_w9070_,
		_w17850_
	);
	LUT3 #(
		.INIT('h2a)
	) name15950 (
		\m7_addr_i[28]_pad ,
		_w9069_,
		_w9070_,
		_w17851_
	);
	LUT4 #(
		.INIT('h6e7f)
	) name15951 (
		_w9064_,
		_w9067_,
		_w17850_,
		_w17851_,
		_w17852_
	);
	LUT4 #(
		.INIT('h7fff)
	) name15952 (
		_w17843_,
		_w17846_,
		_w17849_,
		_w17852_,
		_w17853_
	);
	LUT3 #(
		.INIT('h80)
	) name15953 (
		\m0_addr_i[29]_pad ,
		_w9069_,
		_w9070_,
		_w17854_
	);
	LUT3 #(
		.INIT('h2a)
	) name15954 (
		\m7_addr_i[29]_pad ,
		_w9069_,
		_w9070_,
		_w17855_
	);
	LUT4 #(
		.INIT('h6e7f)
	) name15955 (
		_w9064_,
		_w9067_,
		_w17854_,
		_w17855_,
		_w17856_
	);
	LUT3 #(
		.INIT('h2a)
	) name15956 (
		\m1_addr_i[29]_pad ,
		_w9069_,
		_w9070_,
		_w17857_
	);
	LUT3 #(
		.INIT('h80)
	) name15957 (
		\m4_addr_i[29]_pad ,
		_w9069_,
		_w9070_,
		_w17858_
	);
	LUT4 #(
		.INIT('h5d7f)
	) name15958 (
		_w9064_,
		_w9067_,
		_w17857_,
		_w17858_,
		_w17859_
	);
	LUT3 #(
		.INIT('h80)
	) name15959 (
		\m2_addr_i[29]_pad ,
		_w9069_,
		_w9070_,
		_w17860_
	);
	LUT3 #(
		.INIT('h2a)
	) name15960 (
		\m3_addr_i[29]_pad ,
		_w9069_,
		_w9070_,
		_w17861_
	);
	LUT3 #(
		.INIT('h57)
	) name15961 (
		_w9082_,
		_w17860_,
		_w17861_,
		_w17862_
	);
	LUT3 #(
		.INIT('h2a)
	) name15962 (
		\m5_addr_i[29]_pad ,
		_w9069_,
		_w9070_,
		_w17863_
	);
	LUT3 #(
		.INIT('h80)
	) name15963 (
		\m6_addr_i[29]_pad ,
		_w9069_,
		_w9070_,
		_w17864_
	);
	LUT4 #(
		.INIT('hcedf)
	) name15964 (
		_w9064_,
		_w9067_,
		_w17863_,
		_w17864_,
		_w17865_
	);
	LUT4 #(
		.INIT('h7fff)
	) name15965 (
		_w17856_,
		_w17859_,
		_w17862_,
		_w17865_,
		_w17866_
	);
	LUT3 #(
		.INIT('h2a)
	) name15966 (
		\m3_addr_i[2]_pad ,
		_w9069_,
		_w9070_,
		_w17867_
	);
	LUT3 #(
		.INIT('h80)
	) name15967 (
		\m4_addr_i[2]_pad ,
		_w9069_,
		_w9070_,
		_w17868_
	);
	LUT4 #(
		.INIT('h9dbf)
	) name15968 (
		_w9064_,
		_w9067_,
		_w17867_,
		_w17868_,
		_w17869_
	);
	LUT3 #(
		.INIT('h80)
	) name15969 (
		\m6_addr_i[2]_pad ,
		_w9069_,
		_w9070_,
		_w17870_
	);
	LUT3 #(
		.INIT('h80)
	) name15970 (
		\m2_addr_i[2]_pad ,
		_w9069_,
		_w9070_,
		_w17871_
	);
	LUT4 #(
		.INIT('habef)
	) name15971 (
		_w9064_,
		_w9067_,
		_w17870_,
		_w17871_,
		_w17872_
	);
	LUT3 #(
		.INIT('h2a)
	) name15972 (
		\m5_addr_i[2]_pad ,
		_w9069_,
		_w9070_,
		_w17873_
	);
	LUT3 #(
		.INIT('h2a)
	) name15973 (
		\m1_addr_i[2]_pad ,
		_w9069_,
		_w9070_,
		_w17874_
	);
	LUT4 #(
		.INIT('h57df)
	) name15974 (
		_w9064_,
		_w9067_,
		_w17873_,
		_w17874_,
		_w17875_
	);
	LUT3 #(
		.INIT('h80)
	) name15975 (
		\m0_addr_i[2]_pad ,
		_w9069_,
		_w9070_,
		_w17876_
	);
	LUT3 #(
		.INIT('h2a)
	) name15976 (
		\m7_addr_i[2]_pad ,
		_w9069_,
		_w9070_,
		_w17877_
	);
	LUT4 #(
		.INIT('h6e7f)
	) name15977 (
		_w9064_,
		_w9067_,
		_w17876_,
		_w17877_,
		_w17878_
	);
	LUT4 #(
		.INIT('h7fff)
	) name15978 (
		_w17869_,
		_w17872_,
		_w17875_,
		_w17878_,
		_w17879_
	);
	LUT3 #(
		.INIT('h2a)
	) name15979 (
		\m5_addr_i[30]_pad ,
		_w9069_,
		_w9070_,
		_w17880_
	);
	LUT3 #(
		.INIT('h80)
	) name15980 (
		\m6_addr_i[30]_pad ,
		_w9069_,
		_w9070_,
		_w17881_
	);
	LUT4 #(
		.INIT('hcedf)
	) name15981 (
		_w9064_,
		_w9067_,
		_w17880_,
		_w17881_,
		_w17882_
	);
	LUT3 #(
		.INIT('h80)
	) name15982 (
		\m0_addr_i[30]_pad ,
		_w9069_,
		_w9070_,
		_w17883_
	);
	LUT3 #(
		.INIT('h80)
	) name15983 (
		\m4_addr_i[30]_pad ,
		_w9069_,
		_w9070_,
		_w17884_
	);
	LUT4 #(
		.INIT('h5d7f)
	) name15984 (
		_w9064_,
		_w9067_,
		_w17883_,
		_w17884_,
		_w17885_
	);
	LUT3 #(
		.INIT('h2a)
	) name15985 (
		\m7_addr_i[30]_pad ,
		_w9069_,
		_w9070_,
		_w17886_
	);
	LUT3 #(
		.INIT('h2a)
	) name15986 (
		\m3_addr_i[30]_pad ,
		_w9069_,
		_w9070_,
		_w17887_
	);
	LUT4 #(
		.INIT('habef)
	) name15987 (
		_w9064_,
		_w9067_,
		_w17886_,
		_w17887_,
		_w17888_
	);
	LUT3 #(
		.INIT('h2a)
	) name15988 (
		\m1_addr_i[30]_pad ,
		_w9069_,
		_w9070_,
		_w17889_
	);
	LUT3 #(
		.INIT('h80)
	) name15989 (
		\m2_addr_i[30]_pad ,
		_w9069_,
		_w9070_,
		_w17890_
	);
	LUT4 #(
		.INIT('h3b7f)
	) name15990 (
		_w9064_,
		_w9067_,
		_w17889_,
		_w17890_,
		_w17891_
	);
	LUT4 #(
		.INIT('h7fff)
	) name15991 (
		_w17882_,
		_w17885_,
		_w17888_,
		_w17891_,
		_w17892_
	);
	LUT3 #(
		.INIT('h2a)
	) name15992 (
		\m5_addr_i[31]_pad ,
		_w9069_,
		_w9070_,
		_w17893_
	);
	LUT3 #(
		.INIT('h80)
	) name15993 (
		\m6_addr_i[31]_pad ,
		_w9069_,
		_w9070_,
		_w17894_
	);
	LUT4 #(
		.INIT('hcedf)
	) name15994 (
		_w9064_,
		_w9067_,
		_w17893_,
		_w17894_,
		_w17895_
	);
	LUT3 #(
		.INIT('h2a)
	) name15995 (
		\m3_addr_i[31]_pad ,
		_w9069_,
		_w9070_,
		_w17896_
	);
	LUT3 #(
		.INIT('h2a)
	) name15996 (
		\m7_addr_i[31]_pad ,
		_w9069_,
		_w9070_,
		_w17897_
	);
	LUT4 #(
		.INIT('haebf)
	) name15997 (
		_w9064_,
		_w9067_,
		_w17896_,
		_w17897_,
		_w17898_
	);
	LUT3 #(
		.INIT('h80)
	) name15998 (
		\m4_addr_i[31]_pad ,
		_w9069_,
		_w9070_,
		_w17899_
	);
	LUT3 #(
		.INIT('h80)
	) name15999 (
		\m0_addr_i[31]_pad ,
		_w9069_,
		_w9070_,
		_w17900_
	);
	LUT4 #(
		.INIT('h57df)
	) name16000 (
		_w9064_,
		_w9067_,
		_w17899_,
		_w17900_,
		_w17901_
	);
	LUT3 #(
		.INIT('h2a)
	) name16001 (
		\m1_addr_i[31]_pad ,
		_w9069_,
		_w9070_,
		_w17902_
	);
	LUT3 #(
		.INIT('h80)
	) name16002 (
		\m2_addr_i[31]_pad ,
		_w9069_,
		_w9070_,
		_w17903_
	);
	LUT4 #(
		.INIT('h3b7f)
	) name16003 (
		_w9064_,
		_w9067_,
		_w17902_,
		_w17903_,
		_w17904_
	);
	LUT4 #(
		.INIT('h7fff)
	) name16004 (
		_w17895_,
		_w17898_,
		_w17901_,
		_w17904_,
		_w17905_
	);
	LUT3 #(
		.INIT('h2a)
	) name16005 (
		\m3_addr_i[3]_pad ,
		_w9069_,
		_w9070_,
		_w17906_
	);
	LUT3 #(
		.INIT('h80)
	) name16006 (
		\m4_addr_i[3]_pad ,
		_w9069_,
		_w9070_,
		_w17907_
	);
	LUT4 #(
		.INIT('h9dbf)
	) name16007 (
		_w9064_,
		_w9067_,
		_w17906_,
		_w17907_,
		_w17908_
	);
	LUT3 #(
		.INIT('h80)
	) name16008 (
		\m6_addr_i[3]_pad ,
		_w9069_,
		_w9070_,
		_w17909_
	);
	LUT3 #(
		.INIT('h80)
	) name16009 (
		\m2_addr_i[3]_pad ,
		_w9069_,
		_w9070_,
		_w17910_
	);
	LUT4 #(
		.INIT('habef)
	) name16010 (
		_w9064_,
		_w9067_,
		_w17909_,
		_w17910_,
		_w17911_
	);
	LUT3 #(
		.INIT('h2a)
	) name16011 (
		\m5_addr_i[3]_pad ,
		_w9069_,
		_w9070_,
		_w17912_
	);
	LUT3 #(
		.INIT('h2a)
	) name16012 (
		\m1_addr_i[3]_pad ,
		_w9069_,
		_w9070_,
		_w17913_
	);
	LUT4 #(
		.INIT('h57df)
	) name16013 (
		_w9064_,
		_w9067_,
		_w17912_,
		_w17913_,
		_w17914_
	);
	LUT3 #(
		.INIT('h80)
	) name16014 (
		\m0_addr_i[3]_pad ,
		_w9069_,
		_w9070_,
		_w17915_
	);
	LUT3 #(
		.INIT('h2a)
	) name16015 (
		\m7_addr_i[3]_pad ,
		_w9069_,
		_w9070_,
		_w17916_
	);
	LUT4 #(
		.INIT('h6e7f)
	) name16016 (
		_w9064_,
		_w9067_,
		_w17915_,
		_w17916_,
		_w17917_
	);
	LUT4 #(
		.INIT('h7fff)
	) name16017 (
		_w17908_,
		_w17911_,
		_w17914_,
		_w17917_,
		_w17918_
	);
	LUT3 #(
		.INIT('h2a)
	) name16018 (
		\m3_addr_i[4]_pad ,
		_w9069_,
		_w9070_,
		_w17919_
	);
	LUT3 #(
		.INIT('h80)
	) name16019 (
		\m4_addr_i[4]_pad ,
		_w9069_,
		_w9070_,
		_w17920_
	);
	LUT4 #(
		.INIT('h9dbf)
	) name16020 (
		_w9064_,
		_w9067_,
		_w17919_,
		_w17920_,
		_w17921_
	);
	LUT3 #(
		.INIT('h80)
	) name16021 (
		\m6_addr_i[4]_pad ,
		_w9069_,
		_w9070_,
		_w17922_
	);
	LUT3 #(
		.INIT('h80)
	) name16022 (
		\m2_addr_i[4]_pad ,
		_w9069_,
		_w9070_,
		_w17923_
	);
	LUT4 #(
		.INIT('habef)
	) name16023 (
		_w9064_,
		_w9067_,
		_w17922_,
		_w17923_,
		_w17924_
	);
	LUT3 #(
		.INIT('h2a)
	) name16024 (
		\m5_addr_i[4]_pad ,
		_w9069_,
		_w9070_,
		_w17925_
	);
	LUT3 #(
		.INIT('h2a)
	) name16025 (
		\m1_addr_i[4]_pad ,
		_w9069_,
		_w9070_,
		_w17926_
	);
	LUT4 #(
		.INIT('h57df)
	) name16026 (
		_w9064_,
		_w9067_,
		_w17925_,
		_w17926_,
		_w17927_
	);
	LUT3 #(
		.INIT('h80)
	) name16027 (
		\m0_addr_i[4]_pad ,
		_w9069_,
		_w9070_,
		_w17928_
	);
	LUT3 #(
		.INIT('h2a)
	) name16028 (
		\m7_addr_i[4]_pad ,
		_w9069_,
		_w9070_,
		_w17929_
	);
	LUT4 #(
		.INIT('h6e7f)
	) name16029 (
		_w9064_,
		_w9067_,
		_w17928_,
		_w17929_,
		_w17930_
	);
	LUT4 #(
		.INIT('h7fff)
	) name16030 (
		_w17921_,
		_w17924_,
		_w17927_,
		_w17930_,
		_w17931_
	);
	LUT3 #(
		.INIT('h2a)
	) name16031 (
		\m3_addr_i[5]_pad ,
		_w9069_,
		_w9070_,
		_w17932_
	);
	LUT3 #(
		.INIT('h80)
	) name16032 (
		\m4_addr_i[5]_pad ,
		_w9069_,
		_w9070_,
		_w17933_
	);
	LUT4 #(
		.INIT('h9dbf)
	) name16033 (
		_w9064_,
		_w9067_,
		_w17932_,
		_w17933_,
		_w17934_
	);
	LUT3 #(
		.INIT('h80)
	) name16034 (
		\m6_addr_i[5]_pad ,
		_w9069_,
		_w9070_,
		_w17935_
	);
	LUT3 #(
		.INIT('h80)
	) name16035 (
		\m2_addr_i[5]_pad ,
		_w9069_,
		_w9070_,
		_w17936_
	);
	LUT4 #(
		.INIT('habef)
	) name16036 (
		_w9064_,
		_w9067_,
		_w17935_,
		_w17936_,
		_w17937_
	);
	LUT3 #(
		.INIT('h2a)
	) name16037 (
		\m5_addr_i[5]_pad ,
		_w9069_,
		_w9070_,
		_w17938_
	);
	LUT3 #(
		.INIT('h2a)
	) name16038 (
		\m1_addr_i[5]_pad ,
		_w9069_,
		_w9070_,
		_w17939_
	);
	LUT4 #(
		.INIT('h57df)
	) name16039 (
		_w9064_,
		_w9067_,
		_w17938_,
		_w17939_,
		_w17940_
	);
	LUT3 #(
		.INIT('h80)
	) name16040 (
		\m0_addr_i[5]_pad ,
		_w9069_,
		_w9070_,
		_w17941_
	);
	LUT3 #(
		.INIT('h2a)
	) name16041 (
		\m7_addr_i[5]_pad ,
		_w9069_,
		_w9070_,
		_w17942_
	);
	LUT4 #(
		.INIT('h6e7f)
	) name16042 (
		_w9064_,
		_w9067_,
		_w17941_,
		_w17942_,
		_w17943_
	);
	LUT4 #(
		.INIT('h7fff)
	) name16043 (
		_w17934_,
		_w17937_,
		_w17940_,
		_w17943_,
		_w17944_
	);
	LUT3 #(
		.INIT('h2a)
	) name16044 (
		\m1_addr_i[6]_pad ,
		_w9069_,
		_w9070_,
		_w17945_
	);
	LUT3 #(
		.INIT('h80)
	) name16045 (
		\m2_addr_i[6]_pad ,
		_w9069_,
		_w9070_,
		_w17946_
	);
	LUT4 #(
		.INIT('h3b7f)
	) name16046 (
		_w9064_,
		_w9067_,
		_w17945_,
		_w17946_,
		_w17947_
	);
	LUT3 #(
		.INIT('h80)
	) name16047 (
		\m6_addr_i[6]_pad ,
		_w9069_,
		_w9070_,
		_w17948_
	);
	LUT3 #(
		.INIT('h80)
	) name16048 (
		\m4_addr_i[6]_pad ,
		_w9069_,
		_w9070_,
		_w17949_
	);
	LUT4 #(
		.INIT('hcdef)
	) name16049 (
		_w9064_,
		_w9067_,
		_w17948_,
		_w17949_,
		_w17950_
	);
	LUT3 #(
		.INIT('h2a)
	) name16050 (
		\m5_addr_i[6]_pad ,
		_w9069_,
		_w9070_,
		_w17951_
	);
	LUT3 #(
		.INIT('h2a)
	) name16051 (
		\m3_addr_i[6]_pad ,
		_w9069_,
		_w9070_,
		_w17952_
	);
	LUT4 #(
		.INIT('h9bdf)
	) name16052 (
		_w9064_,
		_w9067_,
		_w17951_,
		_w17952_,
		_w17953_
	);
	LUT3 #(
		.INIT('h80)
	) name16053 (
		\m0_addr_i[6]_pad ,
		_w9069_,
		_w9070_,
		_w17954_
	);
	LUT3 #(
		.INIT('h2a)
	) name16054 (
		\m7_addr_i[6]_pad ,
		_w9069_,
		_w9070_,
		_w17955_
	);
	LUT4 #(
		.INIT('h6e7f)
	) name16055 (
		_w9064_,
		_w9067_,
		_w17954_,
		_w17955_,
		_w17956_
	);
	LUT4 #(
		.INIT('h7fff)
	) name16056 (
		_w17947_,
		_w17950_,
		_w17953_,
		_w17956_,
		_w17957_
	);
	LUT3 #(
		.INIT('h80)
	) name16057 (
		\m6_addr_i[7]_pad ,
		_w9069_,
		_w9070_,
		_w17958_
	);
	LUT3 #(
		.INIT('h2a)
	) name16058 (
		\m5_addr_i[7]_pad ,
		_w9069_,
		_w9070_,
		_w17959_
	);
	LUT4 #(
		.INIT('hcdef)
	) name16059 (
		_w9064_,
		_w9067_,
		_w17958_,
		_w17959_,
		_w17960_
	);
	LUT3 #(
		.INIT('h2a)
	) name16060 (
		\m3_addr_i[7]_pad ,
		_w9069_,
		_w9070_,
		_w17961_
	);
	LUT3 #(
		.INIT('h80)
	) name16061 (
		\m2_addr_i[7]_pad ,
		_w9069_,
		_w9070_,
		_w17962_
	);
	LUT3 #(
		.INIT('h57)
	) name16062 (
		_w9082_,
		_w17961_,
		_w17962_,
		_w17963_
	);
	LUT3 #(
		.INIT('h80)
	) name16063 (
		\m4_addr_i[7]_pad ,
		_w9069_,
		_w9070_,
		_w17964_
	);
	LUT3 #(
		.INIT('h2a)
	) name16064 (
		\m1_addr_i[7]_pad ,
		_w9069_,
		_w9070_,
		_w17965_
	);
	LUT4 #(
		.INIT('h57df)
	) name16065 (
		_w9064_,
		_w9067_,
		_w17964_,
		_w17965_,
		_w17966_
	);
	LUT3 #(
		.INIT('h80)
	) name16066 (
		\m0_addr_i[7]_pad ,
		_w9069_,
		_w9070_,
		_w17967_
	);
	LUT3 #(
		.INIT('h2a)
	) name16067 (
		\m7_addr_i[7]_pad ,
		_w9069_,
		_w9070_,
		_w17968_
	);
	LUT4 #(
		.INIT('h6e7f)
	) name16068 (
		_w9064_,
		_w9067_,
		_w17967_,
		_w17968_,
		_w17969_
	);
	LUT4 #(
		.INIT('h7fff)
	) name16069 (
		_w17960_,
		_w17963_,
		_w17966_,
		_w17969_,
		_w17970_
	);
	LUT3 #(
		.INIT('h80)
	) name16070 (
		\m6_addr_i[8]_pad ,
		_w9069_,
		_w9070_,
		_w17971_
	);
	LUT3 #(
		.INIT('h2a)
	) name16071 (
		\m5_addr_i[8]_pad ,
		_w9069_,
		_w9070_,
		_w17972_
	);
	LUT4 #(
		.INIT('hcdef)
	) name16072 (
		_w9064_,
		_w9067_,
		_w17971_,
		_w17972_,
		_w17973_
	);
	LUT3 #(
		.INIT('h80)
	) name16073 (
		\m0_addr_i[8]_pad ,
		_w9069_,
		_w9070_,
		_w17974_
	);
	LUT3 #(
		.INIT('h80)
	) name16074 (
		\m4_addr_i[8]_pad ,
		_w9069_,
		_w9070_,
		_w17975_
	);
	LUT4 #(
		.INIT('h5d7f)
	) name16075 (
		_w9064_,
		_w9067_,
		_w17974_,
		_w17975_,
		_w17976_
	);
	LUT3 #(
		.INIT('h2a)
	) name16076 (
		\m7_addr_i[8]_pad ,
		_w9069_,
		_w9070_,
		_w17977_
	);
	LUT3 #(
		.INIT('h2a)
	) name16077 (
		\m3_addr_i[8]_pad ,
		_w9069_,
		_w9070_,
		_w17978_
	);
	LUT4 #(
		.INIT('habef)
	) name16078 (
		_w9064_,
		_w9067_,
		_w17977_,
		_w17978_,
		_w17979_
	);
	LUT3 #(
		.INIT('h2a)
	) name16079 (
		\m1_addr_i[8]_pad ,
		_w9069_,
		_w9070_,
		_w17980_
	);
	LUT3 #(
		.INIT('h80)
	) name16080 (
		\m2_addr_i[8]_pad ,
		_w9069_,
		_w9070_,
		_w17981_
	);
	LUT4 #(
		.INIT('h3b7f)
	) name16081 (
		_w9064_,
		_w9067_,
		_w17980_,
		_w17981_,
		_w17982_
	);
	LUT4 #(
		.INIT('h7fff)
	) name16082 (
		_w17973_,
		_w17976_,
		_w17979_,
		_w17982_,
		_w17983_
	);
	LUT3 #(
		.INIT('h2a)
	) name16083 (
		\m3_addr_i[9]_pad ,
		_w9069_,
		_w9070_,
		_w17984_
	);
	LUT3 #(
		.INIT('h80)
	) name16084 (
		\m4_addr_i[9]_pad ,
		_w9069_,
		_w9070_,
		_w17985_
	);
	LUT4 #(
		.INIT('h9dbf)
	) name16085 (
		_w9064_,
		_w9067_,
		_w17984_,
		_w17985_,
		_w17986_
	);
	LUT3 #(
		.INIT('h80)
	) name16086 (
		\m6_addr_i[9]_pad ,
		_w9069_,
		_w9070_,
		_w17987_
	);
	LUT3 #(
		.INIT('h80)
	) name16087 (
		\m2_addr_i[9]_pad ,
		_w9069_,
		_w9070_,
		_w17988_
	);
	LUT4 #(
		.INIT('habef)
	) name16088 (
		_w9064_,
		_w9067_,
		_w17987_,
		_w17988_,
		_w17989_
	);
	LUT3 #(
		.INIT('h2a)
	) name16089 (
		\m5_addr_i[9]_pad ,
		_w9069_,
		_w9070_,
		_w17990_
	);
	LUT3 #(
		.INIT('h2a)
	) name16090 (
		\m1_addr_i[9]_pad ,
		_w9069_,
		_w9070_,
		_w17991_
	);
	LUT4 #(
		.INIT('h57df)
	) name16091 (
		_w9064_,
		_w9067_,
		_w17990_,
		_w17991_,
		_w17992_
	);
	LUT3 #(
		.INIT('h80)
	) name16092 (
		\m0_addr_i[9]_pad ,
		_w9069_,
		_w9070_,
		_w17993_
	);
	LUT3 #(
		.INIT('h2a)
	) name16093 (
		\m7_addr_i[9]_pad ,
		_w9069_,
		_w9070_,
		_w17994_
	);
	LUT4 #(
		.INIT('h6e7f)
	) name16094 (
		_w9064_,
		_w9067_,
		_w17993_,
		_w17994_,
		_w17995_
	);
	LUT4 #(
		.INIT('h7fff)
	) name16095 (
		_w17986_,
		_w17989_,
		_w17992_,
		_w17995_,
		_w17996_
	);
	LUT3 #(
		.INIT('h80)
	) name16096 (
		\m6_data_i[0]_pad ,
		_w9069_,
		_w9070_,
		_w17997_
	);
	LUT3 #(
		.INIT('h2a)
	) name16097 (
		\m5_data_i[0]_pad ,
		_w9069_,
		_w9070_,
		_w17998_
	);
	LUT4 #(
		.INIT('hcdef)
	) name16098 (
		_w9064_,
		_w9067_,
		_w17997_,
		_w17998_,
		_w17999_
	);
	LUT3 #(
		.INIT('h2a)
	) name16099 (
		\m3_data_i[0]_pad ,
		_w9069_,
		_w9070_,
		_w18000_
	);
	LUT3 #(
		.INIT('h80)
	) name16100 (
		\m2_data_i[0]_pad ,
		_w9069_,
		_w9070_,
		_w18001_
	);
	LUT3 #(
		.INIT('h57)
	) name16101 (
		_w9082_,
		_w18000_,
		_w18001_,
		_w18002_
	);
	LUT3 #(
		.INIT('h80)
	) name16102 (
		\m4_data_i[0]_pad ,
		_w9069_,
		_w9070_,
		_w18003_
	);
	LUT3 #(
		.INIT('h2a)
	) name16103 (
		\m1_data_i[0]_pad ,
		_w9069_,
		_w9070_,
		_w18004_
	);
	LUT4 #(
		.INIT('h57df)
	) name16104 (
		_w9064_,
		_w9067_,
		_w18003_,
		_w18004_,
		_w18005_
	);
	LUT3 #(
		.INIT('h80)
	) name16105 (
		\m0_data_i[0]_pad ,
		_w9069_,
		_w9070_,
		_w18006_
	);
	LUT3 #(
		.INIT('h2a)
	) name16106 (
		\m7_data_i[0]_pad ,
		_w9069_,
		_w9070_,
		_w18007_
	);
	LUT4 #(
		.INIT('h6e7f)
	) name16107 (
		_w9064_,
		_w9067_,
		_w18006_,
		_w18007_,
		_w18008_
	);
	LUT4 #(
		.INIT('h7fff)
	) name16108 (
		_w17999_,
		_w18002_,
		_w18005_,
		_w18008_,
		_w18009_
	);
	LUT3 #(
		.INIT('h80)
	) name16109 (
		\m0_data_i[10]_pad ,
		_w9069_,
		_w9070_,
		_w18010_
	);
	LUT3 #(
		.INIT('h2a)
	) name16110 (
		\m7_data_i[10]_pad ,
		_w9069_,
		_w9070_,
		_w18011_
	);
	LUT4 #(
		.INIT('h6e7f)
	) name16111 (
		_w9064_,
		_w9067_,
		_w18010_,
		_w18011_,
		_w18012_
	);
	LUT3 #(
		.INIT('h80)
	) name16112 (
		\m6_data_i[10]_pad ,
		_w9069_,
		_w9070_,
		_w18013_
	);
	LUT3 #(
		.INIT('h80)
	) name16113 (
		\m2_data_i[10]_pad ,
		_w9069_,
		_w9070_,
		_w18014_
	);
	LUT4 #(
		.INIT('habef)
	) name16114 (
		_w9064_,
		_w9067_,
		_w18013_,
		_w18014_,
		_w18015_
	);
	LUT3 #(
		.INIT('h2a)
	) name16115 (
		\m5_data_i[10]_pad ,
		_w9069_,
		_w9070_,
		_w18016_
	);
	LUT3 #(
		.INIT('h2a)
	) name16116 (
		\m1_data_i[10]_pad ,
		_w9069_,
		_w9070_,
		_w18017_
	);
	LUT4 #(
		.INIT('h57df)
	) name16117 (
		_w9064_,
		_w9067_,
		_w18016_,
		_w18017_,
		_w18018_
	);
	LUT3 #(
		.INIT('h2a)
	) name16118 (
		\m3_data_i[10]_pad ,
		_w9069_,
		_w9070_,
		_w18019_
	);
	LUT3 #(
		.INIT('h80)
	) name16119 (
		\m4_data_i[10]_pad ,
		_w9069_,
		_w9070_,
		_w18020_
	);
	LUT4 #(
		.INIT('h9dbf)
	) name16120 (
		_w9064_,
		_w9067_,
		_w18019_,
		_w18020_,
		_w18021_
	);
	LUT4 #(
		.INIT('h7fff)
	) name16121 (
		_w18012_,
		_w18015_,
		_w18018_,
		_w18021_,
		_w18022_
	);
	LUT3 #(
		.INIT('h80)
	) name16122 (
		\m0_data_i[11]_pad ,
		_w9069_,
		_w9070_,
		_w18023_
	);
	LUT3 #(
		.INIT('h2a)
	) name16123 (
		\m7_data_i[11]_pad ,
		_w9069_,
		_w9070_,
		_w18024_
	);
	LUT4 #(
		.INIT('h6e7f)
	) name16124 (
		_w9064_,
		_w9067_,
		_w18023_,
		_w18024_,
		_w18025_
	);
	LUT3 #(
		.INIT('h2a)
	) name16125 (
		\m1_data_i[11]_pad ,
		_w9069_,
		_w9070_,
		_w18026_
	);
	LUT3 #(
		.INIT('h80)
	) name16126 (
		\m4_data_i[11]_pad ,
		_w9069_,
		_w9070_,
		_w18027_
	);
	LUT4 #(
		.INIT('h5d7f)
	) name16127 (
		_w9064_,
		_w9067_,
		_w18026_,
		_w18027_,
		_w18028_
	);
	LUT3 #(
		.INIT('h80)
	) name16128 (
		\m2_data_i[11]_pad ,
		_w9069_,
		_w9070_,
		_w18029_
	);
	LUT3 #(
		.INIT('h2a)
	) name16129 (
		\m3_data_i[11]_pad ,
		_w9069_,
		_w9070_,
		_w18030_
	);
	LUT3 #(
		.INIT('h57)
	) name16130 (
		_w9082_,
		_w18029_,
		_w18030_,
		_w18031_
	);
	LUT3 #(
		.INIT('h80)
	) name16131 (
		\m6_data_i[11]_pad ,
		_w9069_,
		_w9070_,
		_w18032_
	);
	LUT3 #(
		.INIT('h2a)
	) name16132 (
		\m5_data_i[11]_pad ,
		_w9069_,
		_w9070_,
		_w18033_
	);
	LUT4 #(
		.INIT('hcdef)
	) name16133 (
		_w9064_,
		_w9067_,
		_w18032_,
		_w18033_,
		_w18034_
	);
	LUT4 #(
		.INIT('h7fff)
	) name16134 (
		_w18025_,
		_w18028_,
		_w18031_,
		_w18034_,
		_w18035_
	);
	LUT3 #(
		.INIT('h2a)
	) name16135 (
		\m3_data_i[12]_pad ,
		_w9069_,
		_w9070_,
		_w18036_
	);
	LUT3 #(
		.INIT('h80)
	) name16136 (
		\m4_data_i[12]_pad ,
		_w9069_,
		_w9070_,
		_w18037_
	);
	LUT4 #(
		.INIT('h9dbf)
	) name16137 (
		_w9064_,
		_w9067_,
		_w18036_,
		_w18037_,
		_w18038_
	);
	LUT3 #(
		.INIT('h80)
	) name16138 (
		\m0_data_i[12]_pad ,
		_w9069_,
		_w9070_,
		_w18039_
	);
	LUT3 #(
		.INIT('h2a)
	) name16139 (
		\m5_data_i[12]_pad ,
		_w9069_,
		_w9070_,
		_w18040_
	);
	LUT4 #(
		.INIT('h5d7f)
	) name16140 (
		_w9064_,
		_w9067_,
		_w18039_,
		_w18040_,
		_w18041_
	);
	LUT3 #(
		.INIT('h2a)
	) name16141 (
		\m7_data_i[12]_pad ,
		_w9069_,
		_w9070_,
		_w18042_
	);
	LUT3 #(
		.INIT('h80)
	) name16142 (
		\m6_data_i[12]_pad ,
		_w9069_,
		_w9070_,
		_w18043_
	);
	LUT3 #(
		.INIT('h57)
	) name16143 (
		_w9068_,
		_w18042_,
		_w18043_,
		_w18044_
	);
	LUT3 #(
		.INIT('h2a)
	) name16144 (
		\m1_data_i[12]_pad ,
		_w9069_,
		_w9070_,
		_w18045_
	);
	LUT3 #(
		.INIT('h80)
	) name16145 (
		\m2_data_i[12]_pad ,
		_w9069_,
		_w9070_,
		_w18046_
	);
	LUT4 #(
		.INIT('h3b7f)
	) name16146 (
		_w9064_,
		_w9067_,
		_w18045_,
		_w18046_,
		_w18047_
	);
	LUT4 #(
		.INIT('h7fff)
	) name16147 (
		_w18038_,
		_w18041_,
		_w18044_,
		_w18047_,
		_w18048_
	);
	LUT3 #(
		.INIT('h2a)
	) name16148 (
		\m3_data_i[13]_pad ,
		_w9069_,
		_w9070_,
		_w18049_
	);
	LUT3 #(
		.INIT('h80)
	) name16149 (
		\m4_data_i[13]_pad ,
		_w9069_,
		_w9070_,
		_w18050_
	);
	LUT4 #(
		.INIT('h9dbf)
	) name16150 (
		_w9064_,
		_w9067_,
		_w18049_,
		_w18050_,
		_w18051_
	);
	LUT3 #(
		.INIT('h80)
	) name16151 (
		\m0_data_i[13]_pad ,
		_w9069_,
		_w9070_,
		_w18052_
	);
	LUT3 #(
		.INIT('h80)
	) name16152 (
		\m2_data_i[13]_pad ,
		_w9069_,
		_w9070_,
		_w18053_
	);
	LUT4 #(
		.INIT('h3b7f)
	) name16153 (
		_w9064_,
		_w9067_,
		_w18052_,
		_w18053_,
		_w18054_
	);
	LUT3 #(
		.INIT('h2a)
	) name16154 (
		\m7_data_i[13]_pad ,
		_w9069_,
		_w9070_,
		_w18055_
	);
	LUT3 #(
		.INIT('h2a)
	) name16155 (
		\m1_data_i[13]_pad ,
		_w9069_,
		_w9070_,
		_w18056_
	);
	LUT4 #(
		.INIT('h67ef)
	) name16156 (
		_w9064_,
		_w9067_,
		_w18055_,
		_w18056_,
		_w18057_
	);
	LUT3 #(
		.INIT('h80)
	) name16157 (
		\m6_data_i[13]_pad ,
		_w9069_,
		_w9070_,
		_w18058_
	);
	LUT3 #(
		.INIT('h2a)
	) name16158 (
		\m5_data_i[13]_pad ,
		_w9069_,
		_w9070_,
		_w18059_
	);
	LUT4 #(
		.INIT('hcdef)
	) name16159 (
		_w9064_,
		_w9067_,
		_w18058_,
		_w18059_,
		_w18060_
	);
	LUT4 #(
		.INIT('h7fff)
	) name16160 (
		_w18051_,
		_w18054_,
		_w18057_,
		_w18060_,
		_w18061_
	);
	LUT3 #(
		.INIT('h2a)
	) name16161 (
		\m3_data_i[14]_pad ,
		_w9069_,
		_w9070_,
		_w18062_
	);
	LUT3 #(
		.INIT('h80)
	) name16162 (
		\m4_data_i[14]_pad ,
		_w9069_,
		_w9070_,
		_w18063_
	);
	LUT4 #(
		.INIT('h9dbf)
	) name16163 (
		_w9064_,
		_w9067_,
		_w18062_,
		_w18063_,
		_w18064_
	);
	LUT3 #(
		.INIT('h80)
	) name16164 (
		\m6_data_i[14]_pad ,
		_w9069_,
		_w9070_,
		_w18065_
	);
	LUT3 #(
		.INIT('h80)
	) name16165 (
		\m2_data_i[14]_pad ,
		_w9069_,
		_w9070_,
		_w18066_
	);
	LUT4 #(
		.INIT('habef)
	) name16166 (
		_w9064_,
		_w9067_,
		_w18065_,
		_w18066_,
		_w18067_
	);
	LUT3 #(
		.INIT('h2a)
	) name16167 (
		\m5_data_i[14]_pad ,
		_w9069_,
		_w9070_,
		_w18068_
	);
	LUT3 #(
		.INIT('h2a)
	) name16168 (
		\m1_data_i[14]_pad ,
		_w9069_,
		_w9070_,
		_w18069_
	);
	LUT4 #(
		.INIT('h57df)
	) name16169 (
		_w9064_,
		_w9067_,
		_w18068_,
		_w18069_,
		_w18070_
	);
	LUT3 #(
		.INIT('h80)
	) name16170 (
		\m0_data_i[14]_pad ,
		_w9069_,
		_w9070_,
		_w18071_
	);
	LUT3 #(
		.INIT('h2a)
	) name16171 (
		\m7_data_i[14]_pad ,
		_w9069_,
		_w9070_,
		_w18072_
	);
	LUT4 #(
		.INIT('h6e7f)
	) name16172 (
		_w9064_,
		_w9067_,
		_w18071_,
		_w18072_,
		_w18073_
	);
	LUT4 #(
		.INIT('h7fff)
	) name16173 (
		_w18064_,
		_w18067_,
		_w18070_,
		_w18073_,
		_w18074_
	);
	LUT3 #(
		.INIT('h2a)
	) name16174 (
		\m3_data_i[15]_pad ,
		_w9069_,
		_w9070_,
		_w18075_
	);
	LUT3 #(
		.INIT('h80)
	) name16175 (
		\m4_data_i[15]_pad ,
		_w9069_,
		_w9070_,
		_w18076_
	);
	LUT4 #(
		.INIT('h9dbf)
	) name16176 (
		_w9064_,
		_w9067_,
		_w18075_,
		_w18076_,
		_w18077_
	);
	LUT3 #(
		.INIT('h80)
	) name16177 (
		\m6_data_i[15]_pad ,
		_w9069_,
		_w9070_,
		_w18078_
	);
	LUT3 #(
		.INIT('h80)
	) name16178 (
		\m2_data_i[15]_pad ,
		_w9069_,
		_w9070_,
		_w18079_
	);
	LUT4 #(
		.INIT('habef)
	) name16179 (
		_w9064_,
		_w9067_,
		_w18078_,
		_w18079_,
		_w18080_
	);
	LUT3 #(
		.INIT('h2a)
	) name16180 (
		\m5_data_i[15]_pad ,
		_w9069_,
		_w9070_,
		_w18081_
	);
	LUT3 #(
		.INIT('h2a)
	) name16181 (
		\m1_data_i[15]_pad ,
		_w9069_,
		_w9070_,
		_w18082_
	);
	LUT4 #(
		.INIT('h57df)
	) name16182 (
		_w9064_,
		_w9067_,
		_w18081_,
		_w18082_,
		_w18083_
	);
	LUT3 #(
		.INIT('h80)
	) name16183 (
		\m0_data_i[15]_pad ,
		_w9069_,
		_w9070_,
		_w18084_
	);
	LUT3 #(
		.INIT('h2a)
	) name16184 (
		\m7_data_i[15]_pad ,
		_w9069_,
		_w9070_,
		_w18085_
	);
	LUT4 #(
		.INIT('h6e7f)
	) name16185 (
		_w9064_,
		_w9067_,
		_w18084_,
		_w18085_,
		_w18086_
	);
	LUT4 #(
		.INIT('h7fff)
	) name16186 (
		_w18077_,
		_w18080_,
		_w18083_,
		_w18086_,
		_w18087_
	);
	LUT3 #(
		.INIT('h2a)
	) name16187 (
		\m3_data_i[16]_pad ,
		_w9069_,
		_w9070_,
		_w18088_
	);
	LUT3 #(
		.INIT('h80)
	) name16188 (
		\m4_data_i[16]_pad ,
		_w9069_,
		_w9070_,
		_w18089_
	);
	LUT4 #(
		.INIT('h9dbf)
	) name16189 (
		_w9064_,
		_w9067_,
		_w18088_,
		_w18089_,
		_w18090_
	);
	LUT3 #(
		.INIT('h80)
	) name16190 (
		\m6_data_i[16]_pad ,
		_w9069_,
		_w9070_,
		_w18091_
	);
	LUT3 #(
		.INIT('h80)
	) name16191 (
		\m2_data_i[16]_pad ,
		_w9069_,
		_w9070_,
		_w18092_
	);
	LUT4 #(
		.INIT('habef)
	) name16192 (
		_w9064_,
		_w9067_,
		_w18091_,
		_w18092_,
		_w18093_
	);
	LUT3 #(
		.INIT('h2a)
	) name16193 (
		\m5_data_i[16]_pad ,
		_w9069_,
		_w9070_,
		_w18094_
	);
	LUT3 #(
		.INIT('h2a)
	) name16194 (
		\m1_data_i[16]_pad ,
		_w9069_,
		_w9070_,
		_w18095_
	);
	LUT4 #(
		.INIT('h57df)
	) name16195 (
		_w9064_,
		_w9067_,
		_w18094_,
		_w18095_,
		_w18096_
	);
	LUT3 #(
		.INIT('h80)
	) name16196 (
		\m0_data_i[16]_pad ,
		_w9069_,
		_w9070_,
		_w18097_
	);
	LUT3 #(
		.INIT('h2a)
	) name16197 (
		\m7_data_i[16]_pad ,
		_w9069_,
		_w9070_,
		_w18098_
	);
	LUT4 #(
		.INIT('h6e7f)
	) name16198 (
		_w9064_,
		_w9067_,
		_w18097_,
		_w18098_,
		_w18099_
	);
	LUT4 #(
		.INIT('h7fff)
	) name16199 (
		_w18090_,
		_w18093_,
		_w18096_,
		_w18099_,
		_w18100_
	);
	LUT3 #(
		.INIT('h2a)
	) name16200 (
		\m3_data_i[17]_pad ,
		_w9069_,
		_w9070_,
		_w18101_
	);
	LUT3 #(
		.INIT('h80)
	) name16201 (
		\m4_data_i[17]_pad ,
		_w9069_,
		_w9070_,
		_w18102_
	);
	LUT4 #(
		.INIT('h9dbf)
	) name16202 (
		_w9064_,
		_w9067_,
		_w18101_,
		_w18102_,
		_w18103_
	);
	LUT3 #(
		.INIT('h80)
	) name16203 (
		\m6_data_i[17]_pad ,
		_w9069_,
		_w9070_,
		_w18104_
	);
	LUT3 #(
		.INIT('h80)
	) name16204 (
		\m2_data_i[17]_pad ,
		_w9069_,
		_w9070_,
		_w18105_
	);
	LUT4 #(
		.INIT('habef)
	) name16205 (
		_w9064_,
		_w9067_,
		_w18104_,
		_w18105_,
		_w18106_
	);
	LUT3 #(
		.INIT('h2a)
	) name16206 (
		\m5_data_i[17]_pad ,
		_w9069_,
		_w9070_,
		_w18107_
	);
	LUT3 #(
		.INIT('h2a)
	) name16207 (
		\m1_data_i[17]_pad ,
		_w9069_,
		_w9070_,
		_w18108_
	);
	LUT4 #(
		.INIT('h57df)
	) name16208 (
		_w9064_,
		_w9067_,
		_w18107_,
		_w18108_,
		_w18109_
	);
	LUT3 #(
		.INIT('h80)
	) name16209 (
		\m0_data_i[17]_pad ,
		_w9069_,
		_w9070_,
		_w18110_
	);
	LUT3 #(
		.INIT('h2a)
	) name16210 (
		\m7_data_i[17]_pad ,
		_w9069_,
		_w9070_,
		_w18111_
	);
	LUT4 #(
		.INIT('h6e7f)
	) name16211 (
		_w9064_,
		_w9067_,
		_w18110_,
		_w18111_,
		_w18112_
	);
	LUT4 #(
		.INIT('h7fff)
	) name16212 (
		_w18103_,
		_w18106_,
		_w18109_,
		_w18112_,
		_w18113_
	);
	LUT3 #(
		.INIT('h2a)
	) name16213 (
		\m3_data_i[18]_pad ,
		_w9069_,
		_w9070_,
		_w18114_
	);
	LUT3 #(
		.INIT('h80)
	) name16214 (
		\m4_data_i[18]_pad ,
		_w9069_,
		_w9070_,
		_w18115_
	);
	LUT4 #(
		.INIT('h9dbf)
	) name16215 (
		_w9064_,
		_w9067_,
		_w18114_,
		_w18115_,
		_w18116_
	);
	LUT3 #(
		.INIT('h80)
	) name16216 (
		\m6_data_i[18]_pad ,
		_w9069_,
		_w9070_,
		_w18117_
	);
	LUT3 #(
		.INIT('h80)
	) name16217 (
		\m2_data_i[18]_pad ,
		_w9069_,
		_w9070_,
		_w18118_
	);
	LUT4 #(
		.INIT('habef)
	) name16218 (
		_w9064_,
		_w9067_,
		_w18117_,
		_w18118_,
		_w18119_
	);
	LUT3 #(
		.INIT('h2a)
	) name16219 (
		\m5_data_i[18]_pad ,
		_w9069_,
		_w9070_,
		_w18120_
	);
	LUT3 #(
		.INIT('h2a)
	) name16220 (
		\m1_data_i[18]_pad ,
		_w9069_,
		_w9070_,
		_w18121_
	);
	LUT4 #(
		.INIT('h57df)
	) name16221 (
		_w9064_,
		_w9067_,
		_w18120_,
		_w18121_,
		_w18122_
	);
	LUT3 #(
		.INIT('h80)
	) name16222 (
		\m0_data_i[18]_pad ,
		_w9069_,
		_w9070_,
		_w18123_
	);
	LUT3 #(
		.INIT('h2a)
	) name16223 (
		\m7_data_i[18]_pad ,
		_w9069_,
		_w9070_,
		_w18124_
	);
	LUT4 #(
		.INIT('h6e7f)
	) name16224 (
		_w9064_,
		_w9067_,
		_w18123_,
		_w18124_,
		_w18125_
	);
	LUT4 #(
		.INIT('h7fff)
	) name16225 (
		_w18116_,
		_w18119_,
		_w18122_,
		_w18125_,
		_w18126_
	);
	LUT3 #(
		.INIT('h2a)
	) name16226 (
		\m3_data_i[19]_pad ,
		_w9069_,
		_w9070_,
		_w18127_
	);
	LUT3 #(
		.INIT('h80)
	) name16227 (
		\m4_data_i[19]_pad ,
		_w9069_,
		_w9070_,
		_w18128_
	);
	LUT4 #(
		.INIT('h9dbf)
	) name16228 (
		_w9064_,
		_w9067_,
		_w18127_,
		_w18128_,
		_w18129_
	);
	LUT3 #(
		.INIT('h80)
	) name16229 (
		\m6_data_i[19]_pad ,
		_w9069_,
		_w9070_,
		_w18130_
	);
	LUT3 #(
		.INIT('h80)
	) name16230 (
		\m2_data_i[19]_pad ,
		_w9069_,
		_w9070_,
		_w18131_
	);
	LUT4 #(
		.INIT('habef)
	) name16231 (
		_w9064_,
		_w9067_,
		_w18130_,
		_w18131_,
		_w18132_
	);
	LUT3 #(
		.INIT('h2a)
	) name16232 (
		\m5_data_i[19]_pad ,
		_w9069_,
		_w9070_,
		_w18133_
	);
	LUT3 #(
		.INIT('h2a)
	) name16233 (
		\m1_data_i[19]_pad ,
		_w9069_,
		_w9070_,
		_w18134_
	);
	LUT4 #(
		.INIT('h57df)
	) name16234 (
		_w9064_,
		_w9067_,
		_w18133_,
		_w18134_,
		_w18135_
	);
	LUT3 #(
		.INIT('h80)
	) name16235 (
		\m0_data_i[19]_pad ,
		_w9069_,
		_w9070_,
		_w18136_
	);
	LUT3 #(
		.INIT('h2a)
	) name16236 (
		\m7_data_i[19]_pad ,
		_w9069_,
		_w9070_,
		_w18137_
	);
	LUT4 #(
		.INIT('h6e7f)
	) name16237 (
		_w9064_,
		_w9067_,
		_w18136_,
		_w18137_,
		_w18138_
	);
	LUT4 #(
		.INIT('h7fff)
	) name16238 (
		_w18129_,
		_w18132_,
		_w18135_,
		_w18138_,
		_w18139_
	);
	LUT3 #(
		.INIT('h2a)
	) name16239 (
		\m1_data_i[1]_pad ,
		_w9069_,
		_w9070_,
		_w18140_
	);
	LUT3 #(
		.INIT('h80)
	) name16240 (
		\m2_data_i[1]_pad ,
		_w9069_,
		_w9070_,
		_w18141_
	);
	LUT4 #(
		.INIT('h3b7f)
	) name16241 (
		_w9064_,
		_w9067_,
		_w18140_,
		_w18141_,
		_w18142_
	);
	LUT3 #(
		.INIT('h80)
	) name16242 (
		\m0_data_i[1]_pad ,
		_w9069_,
		_w9070_,
		_w18143_
	);
	LUT3 #(
		.INIT('h2a)
	) name16243 (
		\m5_data_i[1]_pad ,
		_w9069_,
		_w9070_,
		_w18144_
	);
	LUT4 #(
		.INIT('h5d7f)
	) name16244 (
		_w9064_,
		_w9067_,
		_w18143_,
		_w18144_,
		_w18145_
	);
	LUT3 #(
		.INIT('h2a)
	) name16245 (
		\m7_data_i[1]_pad ,
		_w9069_,
		_w9070_,
		_w18146_
	);
	LUT3 #(
		.INIT('h80)
	) name16246 (
		\m6_data_i[1]_pad ,
		_w9069_,
		_w9070_,
		_w18147_
	);
	LUT3 #(
		.INIT('h57)
	) name16247 (
		_w9068_,
		_w18146_,
		_w18147_,
		_w18148_
	);
	LUT3 #(
		.INIT('h2a)
	) name16248 (
		\m3_data_i[1]_pad ,
		_w9069_,
		_w9070_,
		_w18149_
	);
	LUT3 #(
		.INIT('h80)
	) name16249 (
		\m4_data_i[1]_pad ,
		_w9069_,
		_w9070_,
		_w18150_
	);
	LUT4 #(
		.INIT('h9dbf)
	) name16250 (
		_w9064_,
		_w9067_,
		_w18149_,
		_w18150_,
		_w18151_
	);
	LUT4 #(
		.INIT('h7fff)
	) name16251 (
		_w18142_,
		_w18145_,
		_w18148_,
		_w18151_,
		_w18152_
	);
	LUT3 #(
		.INIT('h2a)
	) name16252 (
		\m1_data_i[20]_pad ,
		_w9069_,
		_w9070_,
		_w18153_
	);
	LUT3 #(
		.INIT('h80)
	) name16253 (
		\m2_data_i[20]_pad ,
		_w9069_,
		_w9070_,
		_w18154_
	);
	LUT4 #(
		.INIT('h3b7f)
	) name16254 (
		_w9064_,
		_w9067_,
		_w18153_,
		_w18154_,
		_w18155_
	);
	LUT3 #(
		.INIT('h80)
	) name16255 (
		\m0_data_i[20]_pad ,
		_w9069_,
		_w9070_,
		_w18156_
	);
	LUT3 #(
		.INIT('h80)
	) name16256 (
		\m4_data_i[20]_pad ,
		_w9069_,
		_w9070_,
		_w18157_
	);
	LUT4 #(
		.INIT('h5d7f)
	) name16257 (
		_w9064_,
		_w9067_,
		_w18156_,
		_w18157_,
		_w18158_
	);
	LUT3 #(
		.INIT('h2a)
	) name16258 (
		\m7_data_i[20]_pad ,
		_w9069_,
		_w9070_,
		_w18159_
	);
	LUT3 #(
		.INIT('h2a)
	) name16259 (
		\m3_data_i[20]_pad ,
		_w9069_,
		_w9070_,
		_w18160_
	);
	LUT4 #(
		.INIT('habef)
	) name16260 (
		_w9064_,
		_w9067_,
		_w18159_,
		_w18160_,
		_w18161_
	);
	LUT3 #(
		.INIT('h80)
	) name16261 (
		\m6_data_i[20]_pad ,
		_w9069_,
		_w9070_,
		_w18162_
	);
	LUT3 #(
		.INIT('h2a)
	) name16262 (
		\m5_data_i[20]_pad ,
		_w9069_,
		_w9070_,
		_w18163_
	);
	LUT4 #(
		.INIT('hcdef)
	) name16263 (
		_w9064_,
		_w9067_,
		_w18162_,
		_w18163_,
		_w18164_
	);
	LUT4 #(
		.INIT('h7fff)
	) name16264 (
		_w18155_,
		_w18158_,
		_w18161_,
		_w18164_,
		_w18165_
	);
	LUT3 #(
		.INIT('h2a)
	) name16265 (
		\m1_data_i[21]_pad ,
		_w9069_,
		_w9070_,
		_w18166_
	);
	LUT3 #(
		.INIT('h80)
	) name16266 (
		\m2_data_i[21]_pad ,
		_w9069_,
		_w9070_,
		_w18167_
	);
	LUT4 #(
		.INIT('h3b7f)
	) name16267 (
		_w9064_,
		_w9067_,
		_w18166_,
		_w18167_,
		_w18168_
	);
	LUT3 #(
		.INIT('h80)
	) name16268 (
		\m0_data_i[21]_pad ,
		_w9069_,
		_w9070_,
		_w18169_
	);
	LUT3 #(
		.INIT('h80)
	) name16269 (
		\m4_data_i[21]_pad ,
		_w9069_,
		_w9070_,
		_w18170_
	);
	LUT4 #(
		.INIT('h5d7f)
	) name16270 (
		_w9064_,
		_w9067_,
		_w18169_,
		_w18170_,
		_w18171_
	);
	LUT3 #(
		.INIT('h2a)
	) name16271 (
		\m7_data_i[21]_pad ,
		_w9069_,
		_w9070_,
		_w18172_
	);
	LUT3 #(
		.INIT('h2a)
	) name16272 (
		\m3_data_i[21]_pad ,
		_w9069_,
		_w9070_,
		_w18173_
	);
	LUT4 #(
		.INIT('habef)
	) name16273 (
		_w9064_,
		_w9067_,
		_w18172_,
		_w18173_,
		_w18174_
	);
	LUT3 #(
		.INIT('h80)
	) name16274 (
		\m6_data_i[21]_pad ,
		_w9069_,
		_w9070_,
		_w18175_
	);
	LUT3 #(
		.INIT('h2a)
	) name16275 (
		\m5_data_i[21]_pad ,
		_w9069_,
		_w9070_,
		_w18176_
	);
	LUT4 #(
		.INIT('hcdef)
	) name16276 (
		_w9064_,
		_w9067_,
		_w18175_,
		_w18176_,
		_w18177_
	);
	LUT4 #(
		.INIT('h7fff)
	) name16277 (
		_w18168_,
		_w18171_,
		_w18174_,
		_w18177_,
		_w18178_
	);
	LUT3 #(
		.INIT('h2a)
	) name16278 (
		\m1_data_i[22]_pad ,
		_w9069_,
		_w9070_,
		_w18179_
	);
	LUT3 #(
		.INIT('h80)
	) name16279 (
		\m2_data_i[22]_pad ,
		_w9069_,
		_w9070_,
		_w18180_
	);
	LUT4 #(
		.INIT('h3b7f)
	) name16280 (
		_w9064_,
		_w9067_,
		_w18179_,
		_w18180_,
		_w18181_
	);
	LUT3 #(
		.INIT('h80)
	) name16281 (
		\m0_data_i[22]_pad ,
		_w9069_,
		_w9070_,
		_w18182_
	);
	LUT3 #(
		.INIT('h2a)
	) name16282 (
		\m5_data_i[22]_pad ,
		_w9069_,
		_w9070_,
		_w18183_
	);
	LUT4 #(
		.INIT('h5d7f)
	) name16283 (
		_w9064_,
		_w9067_,
		_w18182_,
		_w18183_,
		_w18184_
	);
	LUT3 #(
		.INIT('h2a)
	) name16284 (
		\m7_data_i[22]_pad ,
		_w9069_,
		_w9070_,
		_w18185_
	);
	LUT3 #(
		.INIT('h80)
	) name16285 (
		\m6_data_i[22]_pad ,
		_w9069_,
		_w9070_,
		_w18186_
	);
	LUT3 #(
		.INIT('h57)
	) name16286 (
		_w9068_,
		_w18185_,
		_w18186_,
		_w18187_
	);
	LUT3 #(
		.INIT('h2a)
	) name16287 (
		\m3_data_i[22]_pad ,
		_w9069_,
		_w9070_,
		_w18188_
	);
	LUT3 #(
		.INIT('h80)
	) name16288 (
		\m4_data_i[22]_pad ,
		_w9069_,
		_w9070_,
		_w18189_
	);
	LUT4 #(
		.INIT('h9dbf)
	) name16289 (
		_w9064_,
		_w9067_,
		_w18188_,
		_w18189_,
		_w18190_
	);
	LUT4 #(
		.INIT('h7fff)
	) name16290 (
		_w18181_,
		_w18184_,
		_w18187_,
		_w18190_,
		_w18191_
	);
	LUT3 #(
		.INIT('h2a)
	) name16291 (
		\m1_data_i[23]_pad ,
		_w9069_,
		_w9070_,
		_w18192_
	);
	LUT3 #(
		.INIT('h80)
	) name16292 (
		\m2_data_i[23]_pad ,
		_w9069_,
		_w9070_,
		_w18193_
	);
	LUT4 #(
		.INIT('h3b7f)
	) name16293 (
		_w9064_,
		_w9067_,
		_w18192_,
		_w18193_,
		_w18194_
	);
	LUT3 #(
		.INIT('h80)
	) name16294 (
		\m0_data_i[23]_pad ,
		_w9069_,
		_w9070_,
		_w18195_
	);
	LUT3 #(
		.INIT('h80)
	) name16295 (
		\m4_data_i[23]_pad ,
		_w9069_,
		_w9070_,
		_w18196_
	);
	LUT4 #(
		.INIT('h5d7f)
	) name16296 (
		_w9064_,
		_w9067_,
		_w18195_,
		_w18196_,
		_w18197_
	);
	LUT3 #(
		.INIT('h2a)
	) name16297 (
		\m7_data_i[23]_pad ,
		_w9069_,
		_w9070_,
		_w18198_
	);
	LUT3 #(
		.INIT('h2a)
	) name16298 (
		\m3_data_i[23]_pad ,
		_w9069_,
		_w9070_,
		_w18199_
	);
	LUT4 #(
		.INIT('habef)
	) name16299 (
		_w9064_,
		_w9067_,
		_w18198_,
		_w18199_,
		_w18200_
	);
	LUT3 #(
		.INIT('h80)
	) name16300 (
		\m6_data_i[23]_pad ,
		_w9069_,
		_w9070_,
		_w18201_
	);
	LUT3 #(
		.INIT('h2a)
	) name16301 (
		\m5_data_i[23]_pad ,
		_w9069_,
		_w9070_,
		_w18202_
	);
	LUT4 #(
		.INIT('hcdef)
	) name16302 (
		_w9064_,
		_w9067_,
		_w18201_,
		_w18202_,
		_w18203_
	);
	LUT4 #(
		.INIT('h7fff)
	) name16303 (
		_w18194_,
		_w18197_,
		_w18200_,
		_w18203_,
		_w18204_
	);
	LUT3 #(
		.INIT('h2a)
	) name16304 (
		\m3_data_i[24]_pad ,
		_w9069_,
		_w9070_,
		_w18205_
	);
	LUT3 #(
		.INIT('h80)
	) name16305 (
		\m4_data_i[24]_pad ,
		_w9069_,
		_w9070_,
		_w18206_
	);
	LUT4 #(
		.INIT('h9dbf)
	) name16306 (
		_w9064_,
		_w9067_,
		_w18205_,
		_w18206_,
		_w18207_
	);
	LUT3 #(
		.INIT('h80)
	) name16307 (
		\m6_data_i[24]_pad ,
		_w9069_,
		_w9070_,
		_w18208_
	);
	LUT3 #(
		.INIT('h80)
	) name16308 (
		\m2_data_i[24]_pad ,
		_w9069_,
		_w9070_,
		_w18209_
	);
	LUT4 #(
		.INIT('habef)
	) name16309 (
		_w9064_,
		_w9067_,
		_w18208_,
		_w18209_,
		_w18210_
	);
	LUT3 #(
		.INIT('h2a)
	) name16310 (
		\m5_data_i[24]_pad ,
		_w9069_,
		_w9070_,
		_w18211_
	);
	LUT3 #(
		.INIT('h2a)
	) name16311 (
		\m1_data_i[24]_pad ,
		_w9069_,
		_w9070_,
		_w18212_
	);
	LUT4 #(
		.INIT('h57df)
	) name16312 (
		_w9064_,
		_w9067_,
		_w18211_,
		_w18212_,
		_w18213_
	);
	LUT3 #(
		.INIT('h80)
	) name16313 (
		\m0_data_i[24]_pad ,
		_w9069_,
		_w9070_,
		_w18214_
	);
	LUT3 #(
		.INIT('h2a)
	) name16314 (
		\m7_data_i[24]_pad ,
		_w9069_,
		_w9070_,
		_w18215_
	);
	LUT4 #(
		.INIT('h6e7f)
	) name16315 (
		_w9064_,
		_w9067_,
		_w18214_,
		_w18215_,
		_w18216_
	);
	LUT4 #(
		.INIT('h7fff)
	) name16316 (
		_w18207_,
		_w18210_,
		_w18213_,
		_w18216_,
		_w18217_
	);
	LUT3 #(
		.INIT('h2a)
	) name16317 (
		\m3_data_i[25]_pad ,
		_w9069_,
		_w9070_,
		_w18218_
	);
	LUT3 #(
		.INIT('h80)
	) name16318 (
		\m4_data_i[25]_pad ,
		_w9069_,
		_w9070_,
		_w18219_
	);
	LUT4 #(
		.INIT('h9dbf)
	) name16319 (
		_w9064_,
		_w9067_,
		_w18218_,
		_w18219_,
		_w18220_
	);
	LUT3 #(
		.INIT('h80)
	) name16320 (
		\m6_data_i[25]_pad ,
		_w9069_,
		_w9070_,
		_w18221_
	);
	LUT3 #(
		.INIT('h80)
	) name16321 (
		\m2_data_i[25]_pad ,
		_w9069_,
		_w9070_,
		_w18222_
	);
	LUT4 #(
		.INIT('habef)
	) name16322 (
		_w9064_,
		_w9067_,
		_w18221_,
		_w18222_,
		_w18223_
	);
	LUT3 #(
		.INIT('h2a)
	) name16323 (
		\m5_data_i[25]_pad ,
		_w9069_,
		_w9070_,
		_w18224_
	);
	LUT3 #(
		.INIT('h2a)
	) name16324 (
		\m1_data_i[25]_pad ,
		_w9069_,
		_w9070_,
		_w18225_
	);
	LUT4 #(
		.INIT('h57df)
	) name16325 (
		_w9064_,
		_w9067_,
		_w18224_,
		_w18225_,
		_w18226_
	);
	LUT3 #(
		.INIT('h80)
	) name16326 (
		\m0_data_i[25]_pad ,
		_w9069_,
		_w9070_,
		_w18227_
	);
	LUT3 #(
		.INIT('h2a)
	) name16327 (
		\m7_data_i[25]_pad ,
		_w9069_,
		_w9070_,
		_w18228_
	);
	LUT4 #(
		.INIT('h6e7f)
	) name16328 (
		_w9064_,
		_w9067_,
		_w18227_,
		_w18228_,
		_w18229_
	);
	LUT4 #(
		.INIT('h7fff)
	) name16329 (
		_w18220_,
		_w18223_,
		_w18226_,
		_w18229_,
		_w18230_
	);
	LUT3 #(
		.INIT('h2a)
	) name16330 (
		\m3_data_i[26]_pad ,
		_w9069_,
		_w9070_,
		_w18231_
	);
	LUT3 #(
		.INIT('h80)
	) name16331 (
		\m4_data_i[26]_pad ,
		_w9069_,
		_w9070_,
		_w18232_
	);
	LUT4 #(
		.INIT('h9dbf)
	) name16332 (
		_w9064_,
		_w9067_,
		_w18231_,
		_w18232_,
		_w18233_
	);
	LUT3 #(
		.INIT('h80)
	) name16333 (
		\m6_data_i[26]_pad ,
		_w9069_,
		_w9070_,
		_w18234_
	);
	LUT3 #(
		.INIT('h80)
	) name16334 (
		\m2_data_i[26]_pad ,
		_w9069_,
		_w9070_,
		_w18235_
	);
	LUT4 #(
		.INIT('habef)
	) name16335 (
		_w9064_,
		_w9067_,
		_w18234_,
		_w18235_,
		_w18236_
	);
	LUT3 #(
		.INIT('h2a)
	) name16336 (
		\m5_data_i[26]_pad ,
		_w9069_,
		_w9070_,
		_w18237_
	);
	LUT3 #(
		.INIT('h2a)
	) name16337 (
		\m1_data_i[26]_pad ,
		_w9069_,
		_w9070_,
		_w18238_
	);
	LUT4 #(
		.INIT('h57df)
	) name16338 (
		_w9064_,
		_w9067_,
		_w18237_,
		_w18238_,
		_w18239_
	);
	LUT3 #(
		.INIT('h80)
	) name16339 (
		\m0_data_i[26]_pad ,
		_w9069_,
		_w9070_,
		_w18240_
	);
	LUT3 #(
		.INIT('h2a)
	) name16340 (
		\m7_data_i[26]_pad ,
		_w9069_,
		_w9070_,
		_w18241_
	);
	LUT4 #(
		.INIT('h6e7f)
	) name16341 (
		_w9064_,
		_w9067_,
		_w18240_,
		_w18241_,
		_w18242_
	);
	LUT4 #(
		.INIT('h7fff)
	) name16342 (
		_w18233_,
		_w18236_,
		_w18239_,
		_w18242_,
		_w18243_
	);
	LUT3 #(
		.INIT('h2a)
	) name16343 (
		\m3_data_i[27]_pad ,
		_w9069_,
		_w9070_,
		_w18244_
	);
	LUT3 #(
		.INIT('h80)
	) name16344 (
		\m4_data_i[27]_pad ,
		_w9069_,
		_w9070_,
		_w18245_
	);
	LUT4 #(
		.INIT('h9dbf)
	) name16345 (
		_w9064_,
		_w9067_,
		_w18244_,
		_w18245_,
		_w18246_
	);
	LUT3 #(
		.INIT('h80)
	) name16346 (
		\m6_data_i[27]_pad ,
		_w9069_,
		_w9070_,
		_w18247_
	);
	LUT3 #(
		.INIT('h80)
	) name16347 (
		\m2_data_i[27]_pad ,
		_w9069_,
		_w9070_,
		_w18248_
	);
	LUT4 #(
		.INIT('habef)
	) name16348 (
		_w9064_,
		_w9067_,
		_w18247_,
		_w18248_,
		_w18249_
	);
	LUT3 #(
		.INIT('h2a)
	) name16349 (
		\m5_data_i[27]_pad ,
		_w9069_,
		_w9070_,
		_w18250_
	);
	LUT3 #(
		.INIT('h2a)
	) name16350 (
		\m1_data_i[27]_pad ,
		_w9069_,
		_w9070_,
		_w18251_
	);
	LUT4 #(
		.INIT('h57df)
	) name16351 (
		_w9064_,
		_w9067_,
		_w18250_,
		_w18251_,
		_w18252_
	);
	LUT3 #(
		.INIT('h80)
	) name16352 (
		\m0_data_i[27]_pad ,
		_w9069_,
		_w9070_,
		_w18253_
	);
	LUT3 #(
		.INIT('h2a)
	) name16353 (
		\m7_data_i[27]_pad ,
		_w9069_,
		_w9070_,
		_w18254_
	);
	LUT4 #(
		.INIT('h6e7f)
	) name16354 (
		_w9064_,
		_w9067_,
		_w18253_,
		_w18254_,
		_w18255_
	);
	LUT4 #(
		.INIT('h7fff)
	) name16355 (
		_w18246_,
		_w18249_,
		_w18252_,
		_w18255_,
		_w18256_
	);
	LUT3 #(
		.INIT('h2a)
	) name16356 (
		\m3_data_i[28]_pad ,
		_w9069_,
		_w9070_,
		_w18257_
	);
	LUT3 #(
		.INIT('h80)
	) name16357 (
		\m4_data_i[28]_pad ,
		_w9069_,
		_w9070_,
		_w18258_
	);
	LUT4 #(
		.INIT('h9dbf)
	) name16358 (
		_w9064_,
		_w9067_,
		_w18257_,
		_w18258_,
		_w18259_
	);
	LUT3 #(
		.INIT('h80)
	) name16359 (
		\m6_data_i[28]_pad ,
		_w9069_,
		_w9070_,
		_w18260_
	);
	LUT3 #(
		.INIT('h80)
	) name16360 (
		\m2_data_i[28]_pad ,
		_w9069_,
		_w9070_,
		_w18261_
	);
	LUT4 #(
		.INIT('habef)
	) name16361 (
		_w9064_,
		_w9067_,
		_w18260_,
		_w18261_,
		_w18262_
	);
	LUT3 #(
		.INIT('h2a)
	) name16362 (
		\m5_data_i[28]_pad ,
		_w9069_,
		_w9070_,
		_w18263_
	);
	LUT3 #(
		.INIT('h2a)
	) name16363 (
		\m1_data_i[28]_pad ,
		_w9069_,
		_w9070_,
		_w18264_
	);
	LUT4 #(
		.INIT('h57df)
	) name16364 (
		_w9064_,
		_w9067_,
		_w18263_,
		_w18264_,
		_w18265_
	);
	LUT3 #(
		.INIT('h80)
	) name16365 (
		\m0_data_i[28]_pad ,
		_w9069_,
		_w9070_,
		_w18266_
	);
	LUT3 #(
		.INIT('h2a)
	) name16366 (
		\m7_data_i[28]_pad ,
		_w9069_,
		_w9070_,
		_w18267_
	);
	LUT4 #(
		.INIT('h6e7f)
	) name16367 (
		_w9064_,
		_w9067_,
		_w18266_,
		_w18267_,
		_w18268_
	);
	LUT4 #(
		.INIT('h7fff)
	) name16368 (
		_w18259_,
		_w18262_,
		_w18265_,
		_w18268_,
		_w18269_
	);
	LUT3 #(
		.INIT('h2a)
	) name16369 (
		\m3_data_i[29]_pad ,
		_w9069_,
		_w9070_,
		_w18270_
	);
	LUT3 #(
		.INIT('h80)
	) name16370 (
		\m4_data_i[29]_pad ,
		_w9069_,
		_w9070_,
		_w18271_
	);
	LUT4 #(
		.INIT('h9dbf)
	) name16371 (
		_w9064_,
		_w9067_,
		_w18270_,
		_w18271_,
		_w18272_
	);
	LUT3 #(
		.INIT('h80)
	) name16372 (
		\m6_data_i[29]_pad ,
		_w9069_,
		_w9070_,
		_w18273_
	);
	LUT3 #(
		.INIT('h80)
	) name16373 (
		\m2_data_i[29]_pad ,
		_w9069_,
		_w9070_,
		_w18274_
	);
	LUT4 #(
		.INIT('habef)
	) name16374 (
		_w9064_,
		_w9067_,
		_w18273_,
		_w18274_,
		_w18275_
	);
	LUT3 #(
		.INIT('h2a)
	) name16375 (
		\m5_data_i[29]_pad ,
		_w9069_,
		_w9070_,
		_w18276_
	);
	LUT3 #(
		.INIT('h2a)
	) name16376 (
		\m1_data_i[29]_pad ,
		_w9069_,
		_w9070_,
		_w18277_
	);
	LUT4 #(
		.INIT('h57df)
	) name16377 (
		_w9064_,
		_w9067_,
		_w18276_,
		_w18277_,
		_w18278_
	);
	LUT3 #(
		.INIT('h80)
	) name16378 (
		\m0_data_i[29]_pad ,
		_w9069_,
		_w9070_,
		_w18279_
	);
	LUT3 #(
		.INIT('h2a)
	) name16379 (
		\m7_data_i[29]_pad ,
		_w9069_,
		_w9070_,
		_w18280_
	);
	LUT4 #(
		.INIT('h6e7f)
	) name16380 (
		_w9064_,
		_w9067_,
		_w18279_,
		_w18280_,
		_w18281_
	);
	LUT4 #(
		.INIT('h7fff)
	) name16381 (
		_w18272_,
		_w18275_,
		_w18278_,
		_w18281_,
		_w18282_
	);
	LUT3 #(
		.INIT('h80)
	) name16382 (
		\m0_data_i[2]_pad ,
		_w9069_,
		_w9070_,
		_w18283_
	);
	LUT3 #(
		.INIT('h2a)
	) name16383 (
		\m7_data_i[2]_pad ,
		_w9069_,
		_w9070_,
		_w18284_
	);
	LUT4 #(
		.INIT('h6e7f)
	) name16384 (
		_w9064_,
		_w9067_,
		_w18283_,
		_w18284_,
		_w18285_
	);
	LUT3 #(
		.INIT('h2a)
	) name16385 (
		\m1_data_i[2]_pad ,
		_w9069_,
		_w9070_,
		_w18286_
	);
	LUT3 #(
		.INIT('h2a)
	) name16386 (
		\m5_data_i[2]_pad ,
		_w9069_,
		_w9070_,
		_w18287_
	);
	LUT4 #(
		.INIT('h5d7f)
	) name16387 (
		_w9064_,
		_w9067_,
		_w18286_,
		_w18287_,
		_w18288_
	);
	LUT3 #(
		.INIT('h80)
	) name16388 (
		\m2_data_i[2]_pad ,
		_w9069_,
		_w9070_,
		_w18289_
	);
	LUT3 #(
		.INIT('h80)
	) name16389 (
		\m6_data_i[2]_pad ,
		_w9069_,
		_w9070_,
		_w18290_
	);
	LUT4 #(
		.INIT('haebf)
	) name16390 (
		_w9064_,
		_w9067_,
		_w18289_,
		_w18290_,
		_w18291_
	);
	LUT3 #(
		.INIT('h2a)
	) name16391 (
		\m3_data_i[2]_pad ,
		_w9069_,
		_w9070_,
		_w18292_
	);
	LUT3 #(
		.INIT('h80)
	) name16392 (
		\m4_data_i[2]_pad ,
		_w9069_,
		_w9070_,
		_w18293_
	);
	LUT4 #(
		.INIT('h9dbf)
	) name16393 (
		_w9064_,
		_w9067_,
		_w18292_,
		_w18293_,
		_w18294_
	);
	LUT4 #(
		.INIT('h7fff)
	) name16394 (
		_w18285_,
		_w18288_,
		_w18291_,
		_w18294_,
		_w18295_
	);
	LUT3 #(
		.INIT('h2a)
	) name16395 (
		\m3_data_i[30]_pad ,
		_w9069_,
		_w9070_,
		_w18296_
	);
	LUT3 #(
		.INIT('h80)
	) name16396 (
		\m4_data_i[30]_pad ,
		_w9069_,
		_w9070_,
		_w18297_
	);
	LUT4 #(
		.INIT('h9dbf)
	) name16397 (
		_w9064_,
		_w9067_,
		_w18296_,
		_w18297_,
		_w18298_
	);
	LUT3 #(
		.INIT('h80)
	) name16398 (
		\m6_data_i[30]_pad ,
		_w9069_,
		_w9070_,
		_w18299_
	);
	LUT3 #(
		.INIT('h80)
	) name16399 (
		\m2_data_i[30]_pad ,
		_w9069_,
		_w9070_,
		_w18300_
	);
	LUT4 #(
		.INIT('habef)
	) name16400 (
		_w9064_,
		_w9067_,
		_w18299_,
		_w18300_,
		_w18301_
	);
	LUT3 #(
		.INIT('h2a)
	) name16401 (
		\m5_data_i[30]_pad ,
		_w9069_,
		_w9070_,
		_w18302_
	);
	LUT3 #(
		.INIT('h2a)
	) name16402 (
		\m1_data_i[30]_pad ,
		_w9069_,
		_w9070_,
		_w18303_
	);
	LUT4 #(
		.INIT('h57df)
	) name16403 (
		_w9064_,
		_w9067_,
		_w18302_,
		_w18303_,
		_w18304_
	);
	LUT3 #(
		.INIT('h80)
	) name16404 (
		\m0_data_i[30]_pad ,
		_w9069_,
		_w9070_,
		_w18305_
	);
	LUT3 #(
		.INIT('h2a)
	) name16405 (
		\m7_data_i[30]_pad ,
		_w9069_,
		_w9070_,
		_w18306_
	);
	LUT4 #(
		.INIT('h6e7f)
	) name16406 (
		_w9064_,
		_w9067_,
		_w18305_,
		_w18306_,
		_w18307_
	);
	LUT4 #(
		.INIT('h7fff)
	) name16407 (
		_w18298_,
		_w18301_,
		_w18304_,
		_w18307_,
		_w18308_
	);
	LUT3 #(
		.INIT('h2a)
	) name16408 (
		\m3_data_i[31]_pad ,
		_w9069_,
		_w9070_,
		_w18309_
	);
	LUT3 #(
		.INIT('h80)
	) name16409 (
		\m4_data_i[31]_pad ,
		_w9069_,
		_w9070_,
		_w18310_
	);
	LUT4 #(
		.INIT('h9dbf)
	) name16410 (
		_w9064_,
		_w9067_,
		_w18309_,
		_w18310_,
		_w18311_
	);
	LUT3 #(
		.INIT('h80)
	) name16411 (
		\m6_data_i[31]_pad ,
		_w9069_,
		_w9070_,
		_w18312_
	);
	LUT3 #(
		.INIT('h80)
	) name16412 (
		\m2_data_i[31]_pad ,
		_w9069_,
		_w9070_,
		_w18313_
	);
	LUT4 #(
		.INIT('habef)
	) name16413 (
		_w9064_,
		_w9067_,
		_w18312_,
		_w18313_,
		_w18314_
	);
	LUT3 #(
		.INIT('h2a)
	) name16414 (
		\m5_data_i[31]_pad ,
		_w9069_,
		_w9070_,
		_w18315_
	);
	LUT3 #(
		.INIT('h2a)
	) name16415 (
		\m1_data_i[31]_pad ,
		_w9069_,
		_w9070_,
		_w18316_
	);
	LUT4 #(
		.INIT('h57df)
	) name16416 (
		_w9064_,
		_w9067_,
		_w18315_,
		_w18316_,
		_w18317_
	);
	LUT3 #(
		.INIT('h80)
	) name16417 (
		\m0_data_i[31]_pad ,
		_w9069_,
		_w9070_,
		_w18318_
	);
	LUT3 #(
		.INIT('h2a)
	) name16418 (
		\m7_data_i[31]_pad ,
		_w9069_,
		_w9070_,
		_w18319_
	);
	LUT4 #(
		.INIT('h6e7f)
	) name16419 (
		_w9064_,
		_w9067_,
		_w18318_,
		_w18319_,
		_w18320_
	);
	LUT4 #(
		.INIT('h7fff)
	) name16420 (
		_w18311_,
		_w18314_,
		_w18317_,
		_w18320_,
		_w18321_
	);
	LUT3 #(
		.INIT('h2a)
	) name16421 (
		\m3_data_i[3]_pad ,
		_w9069_,
		_w9070_,
		_w18322_
	);
	LUT3 #(
		.INIT('h80)
	) name16422 (
		\m4_data_i[3]_pad ,
		_w9069_,
		_w9070_,
		_w18323_
	);
	LUT4 #(
		.INIT('h9dbf)
	) name16423 (
		_w9064_,
		_w9067_,
		_w18322_,
		_w18323_,
		_w18324_
	);
	LUT3 #(
		.INIT('h80)
	) name16424 (
		\m6_data_i[3]_pad ,
		_w9069_,
		_w9070_,
		_w18325_
	);
	LUT3 #(
		.INIT('h2a)
	) name16425 (
		\m7_data_i[3]_pad ,
		_w9069_,
		_w9070_,
		_w18326_
	);
	LUT3 #(
		.INIT('h57)
	) name16426 (
		_w9068_,
		_w18325_,
		_w18326_,
		_w18327_
	);
	LUT3 #(
		.INIT('h2a)
	) name16427 (
		\m5_data_i[3]_pad ,
		_w9069_,
		_w9070_,
		_w18328_
	);
	LUT3 #(
		.INIT('h80)
	) name16428 (
		\m0_data_i[3]_pad ,
		_w9069_,
		_w9070_,
		_w18329_
	);
	LUT4 #(
		.INIT('h57df)
	) name16429 (
		_w9064_,
		_w9067_,
		_w18328_,
		_w18329_,
		_w18330_
	);
	LUT3 #(
		.INIT('h2a)
	) name16430 (
		\m1_data_i[3]_pad ,
		_w9069_,
		_w9070_,
		_w18331_
	);
	LUT3 #(
		.INIT('h80)
	) name16431 (
		\m2_data_i[3]_pad ,
		_w9069_,
		_w9070_,
		_w18332_
	);
	LUT4 #(
		.INIT('h3b7f)
	) name16432 (
		_w9064_,
		_w9067_,
		_w18331_,
		_w18332_,
		_w18333_
	);
	LUT4 #(
		.INIT('h7fff)
	) name16433 (
		_w18324_,
		_w18327_,
		_w18330_,
		_w18333_,
		_w18334_
	);
	LUT3 #(
		.INIT('h80)
	) name16434 (
		\m6_data_i[4]_pad ,
		_w9069_,
		_w9070_,
		_w18335_
	);
	LUT3 #(
		.INIT('h2a)
	) name16435 (
		\m5_data_i[4]_pad ,
		_w9069_,
		_w9070_,
		_w18336_
	);
	LUT4 #(
		.INIT('hcdef)
	) name16436 (
		_w9064_,
		_w9067_,
		_w18335_,
		_w18336_,
		_w18337_
	);
	LUT3 #(
		.INIT('h2a)
	) name16437 (
		\m1_data_i[4]_pad ,
		_w9069_,
		_w9070_,
		_w18338_
	);
	LUT3 #(
		.INIT('h80)
	) name16438 (
		\m4_data_i[4]_pad ,
		_w9069_,
		_w9070_,
		_w18339_
	);
	LUT4 #(
		.INIT('h5d7f)
	) name16439 (
		_w9064_,
		_w9067_,
		_w18338_,
		_w18339_,
		_w18340_
	);
	LUT3 #(
		.INIT('h80)
	) name16440 (
		\m2_data_i[4]_pad ,
		_w9069_,
		_w9070_,
		_w18341_
	);
	LUT3 #(
		.INIT('h2a)
	) name16441 (
		\m3_data_i[4]_pad ,
		_w9069_,
		_w9070_,
		_w18342_
	);
	LUT3 #(
		.INIT('h57)
	) name16442 (
		_w9082_,
		_w18341_,
		_w18342_,
		_w18343_
	);
	LUT3 #(
		.INIT('h80)
	) name16443 (
		\m0_data_i[4]_pad ,
		_w9069_,
		_w9070_,
		_w18344_
	);
	LUT3 #(
		.INIT('h2a)
	) name16444 (
		\m7_data_i[4]_pad ,
		_w9069_,
		_w9070_,
		_w18345_
	);
	LUT4 #(
		.INIT('h6e7f)
	) name16445 (
		_w9064_,
		_w9067_,
		_w18344_,
		_w18345_,
		_w18346_
	);
	LUT4 #(
		.INIT('h7fff)
	) name16446 (
		_w18337_,
		_w18340_,
		_w18343_,
		_w18346_,
		_w18347_
	);
	LUT3 #(
		.INIT('h2a)
	) name16447 (
		\m1_data_i[5]_pad ,
		_w9069_,
		_w9070_,
		_w18348_
	);
	LUT3 #(
		.INIT('h80)
	) name16448 (
		\m2_data_i[5]_pad ,
		_w9069_,
		_w9070_,
		_w18349_
	);
	LUT4 #(
		.INIT('h3b7f)
	) name16449 (
		_w9064_,
		_w9067_,
		_w18348_,
		_w18349_,
		_w18350_
	);
	LUT3 #(
		.INIT('h2a)
	) name16450 (
		\m3_data_i[5]_pad ,
		_w9069_,
		_w9070_,
		_w18351_
	);
	LUT3 #(
		.INIT('h2a)
	) name16451 (
		\m7_data_i[5]_pad ,
		_w9069_,
		_w9070_,
		_w18352_
	);
	LUT4 #(
		.INIT('haebf)
	) name16452 (
		_w9064_,
		_w9067_,
		_w18351_,
		_w18352_,
		_w18353_
	);
	LUT3 #(
		.INIT('h80)
	) name16453 (
		\m4_data_i[5]_pad ,
		_w9069_,
		_w9070_,
		_w18354_
	);
	LUT3 #(
		.INIT('h80)
	) name16454 (
		\m0_data_i[5]_pad ,
		_w9069_,
		_w9070_,
		_w18355_
	);
	LUT4 #(
		.INIT('h57df)
	) name16455 (
		_w9064_,
		_w9067_,
		_w18354_,
		_w18355_,
		_w18356_
	);
	LUT3 #(
		.INIT('h80)
	) name16456 (
		\m6_data_i[5]_pad ,
		_w9069_,
		_w9070_,
		_w18357_
	);
	LUT3 #(
		.INIT('h2a)
	) name16457 (
		\m5_data_i[5]_pad ,
		_w9069_,
		_w9070_,
		_w18358_
	);
	LUT4 #(
		.INIT('hcdef)
	) name16458 (
		_w9064_,
		_w9067_,
		_w18357_,
		_w18358_,
		_w18359_
	);
	LUT4 #(
		.INIT('h7fff)
	) name16459 (
		_w18350_,
		_w18353_,
		_w18356_,
		_w18359_,
		_w18360_
	);
	LUT3 #(
		.INIT('h2a)
	) name16460 (
		\m3_data_i[6]_pad ,
		_w9069_,
		_w9070_,
		_w18361_
	);
	LUT3 #(
		.INIT('h80)
	) name16461 (
		\m4_data_i[6]_pad ,
		_w9069_,
		_w9070_,
		_w18362_
	);
	LUT4 #(
		.INIT('h9dbf)
	) name16462 (
		_w9064_,
		_w9067_,
		_w18361_,
		_w18362_,
		_w18363_
	);
	LUT3 #(
		.INIT('h80)
	) name16463 (
		\m0_data_i[6]_pad ,
		_w9069_,
		_w9070_,
		_w18364_
	);
	LUT3 #(
		.INIT('h2a)
	) name16464 (
		\m5_data_i[6]_pad ,
		_w9069_,
		_w9070_,
		_w18365_
	);
	LUT4 #(
		.INIT('h5d7f)
	) name16465 (
		_w9064_,
		_w9067_,
		_w18364_,
		_w18365_,
		_w18366_
	);
	LUT3 #(
		.INIT('h2a)
	) name16466 (
		\m7_data_i[6]_pad ,
		_w9069_,
		_w9070_,
		_w18367_
	);
	LUT3 #(
		.INIT('h80)
	) name16467 (
		\m6_data_i[6]_pad ,
		_w9069_,
		_w9070_,
		_w18368_
	);
	LUT3 #(
		.INIT('h57)
	) name16468 (
		_w9068_,
		_w18367_,
		_w18368_,
		_w18369_
	);
	LUT3 #(
		.INIT('h2a)
	) name16469 (
		\m1_data_i[6]_pad ,
		_w9069_,
		_w9070_,
		_w18370_
	);
	LUT3 #(
		.INIT('h80)
	) name16470 (
		\m2_data_i[6]_pad ,
		_w9069_,
		_w9070_,
		_w18371_
	);
	LUT4 #(
		.INIT('h3b7f)
	) name16471 (
		_w9064_,
		_w9067_,
		_w18370_,
		_w18371_,
		_w18372_
	);
	LUT4 #(
		.INIT('h7fff)
	) name16472 (
		_w18363_,
		_w18366_,
		_w18369_,
		_w18372_,
		_w18373_
	);
	LUT3 #(
		.INIT('h2a)
	) name16473 (
		\m3_data_i[7]_pad ,
		_w9069_,
		_w9070_,
		_w18374_
	);
	LUT3 #(
		.INIT('h80)
	) name16474 (
		\m4_data_i[7]_pad ,
		_w9069_,
		_w9070_,
		_w18375_
	);
	LUT4 #(
		.INIT('h9dbf)
	) name16475 (
		_w9064_,
		_w9067_,
		_w18374_,
		_w18375_,
		_w18376_
	);
	LUT3 #(
		.INIT('h80)
	) name16476 (
		\m6_data_i[7]_pad ,
		_w9069_,
		_w9070_,
		_w18377_
	);
	LUT3 #(
		.INIT('h80)
	) name16477 (
		\m2_data_i[7]_pad ,
		_w9069_,
		_w9070_,
		_w18378_
	);
	LUT4 #(
		.INIT('habef)
	) name16478 (
		_w9064_,
		_w9067_,
		_w18377_,
		_w18378_,
		_w18379_
	);
	LUT3 #(
		.INIT('h2a)
	) name16479 (
		\m5_data_i[7]_pad ,
		_w9069_,
		_w9070_,
		_w18380_
	);
	LUT3 #(
		.INIT('h2a)
	) name16480 (
		\m1_data_i[7]_pad ,
		_w9069_,
		_w9070_,
		_w18381_
	);
	LUT4 #(
		.INIT('h57df)
	) name16481 (
		_w9064_,
		_w9067_,
		_w18380_,
		_w18381_,
		_w18382_
	);
	LUT3 #(
		.INIT('h80)
	) name16482 (
		\m0_data_i[7]_pad ,
		_w9069_,
		_w9070_,
		_w18383_
	);
	LUT3 #(
		.INIT('h2a)
	) name16483 (
		\m7_data_i[7]_pad ,
		_w9069_,
		_w9070_,
		_w18384_
	);
	LUT4 #(
		.INIT('h6e7f)
	) name16484 (
		_w9064_,
		_w9067_,
		_w18383_,
		_w18384_,
		_w18385_
	);
	LUT4 #(
		.INIT('h7fff)
	) name16485 (
		_w18376_,
		_w18379_,
		_w18382_,
		_w18385_,
		_w18386_
	);
	LUT3 #(
		.INIT('h80)
	) name16486 (
		\m0_data_i[8]_pad ,
		_w9069_,
		_w9070_,
		_w18387_
	);
	LUT3 #(
		.INIT('h2a)
	) name16487 (
		\m7_data_i[8]_pad ,
		_w9069_,
		_w9070_,
		_w18388_
	);
	LUT4 #(
		.INIT('h6e7f)
	) name16488 (
		_w9064_,
		_w9067_,
		_w18387_,
		_w18388_,
		_w18389_
	);
	LUT3 #(
		.INIT('h2a)
	) name16489 (
		\m1_data_i[8]_pad ,
		_w9069_,
		_w9070_,
		_w18390_
	);
	LUT3 #(
		.INIT('h80)
	) name16490 (
		\m4_data_i[8]_pad ,
		_w9069_,
		_w9070_,
		_w18391_
	);
	LUT4 #(
		.INIT('h5d7f)
	) name16491 (
		_w9064_,
		_w9067_,
		_w18390_,
		_w18391_,
		_w18392_
	);
	LUT3 #(
		.INIT('h80)
	) name16492 (
		\m2_data_i[8]_pad ,
		_w9069_,
		_w9070_,
		_w18393_
	);
	LUT3 #(
		.INIT('h2a)
	) name16493 (
		\m3_data_i[8]_pad ,
		_w9069_,
		_w9070_,
		_w18394_
	);
	LUT3 #(
		.INIT('h57)
	) name16494 (
		_w9082_,
		_w18393_,
		_w18394_,
		_w18395_
	);
	LUT3 #(
		.INIT('h80)
	) name16495 (
		\m6_data_i[8]_pad ,
		_w9069_,
		_w9070_,
		_w18396_
	);
	LUT3 #(
		.INIT('h2a)
	) name16496 (
		\m5_data_i[8]_pad ,
		_w9069_,
		_w9070_,
		_w18397_
	);
	LUT4 #(
		.INIT('hcdef)
	) name16497 (
		_w9064_,
		_w9067_,
		_w18396_,
		_w18397_,
		_w18398_
	);
	LUT4 #(
		.INIT('h7fff)
	) name16498 (
		_w18389_,
		_w18392_,
		_w18395_,
		_w18398_,
		_w18399_
	);
	LUT3 #(
		.INIT('h80)
	) name16499 (
		\m6_data_i[9]_pad ,
		_w9069_,
		_w9070_,
		_w18400_
	);
	LUT3 #(
		.INIT('h2a)
	) name16500 (
		\m5_data_i[9]_pad ,
		_w9069_,
		_w9070_,
		_w18401_
	);
	LUT4 #(
		.INIT('hcdef)
	) name16501 (
		_w9064_,
		_w9067_,
		_w18400_,
		_w18401_,
		_w18402_
	);
	LUT3 #(
		.INIT('h2a)
	) name16502 (
		\m3_data_i[9]_pad ,
		_w9069_,
		_w9070_,
		_w18403_
	);
	LUT3 #(
		.INIT('h2a)
	) name16503 (
		\m7_data_i[9]_pad ,
		_w9069_,
		_w9070_,
		_w18404_
	);
	LUT4 #(
		.INIT('haebf)
	) name16504 (
		_w9064_,
		_w9067_,
		_w18403_,
		_w18404_,
		_w18405_
	);
	LUT3 #(
		.INIT('h80)
	) name16505 (
		\m4_data_i[9]_pad ,
		_w9069_,
		_w9070_,
		_w18406_
	);
	LUT3 #(
		.INIT('h80)
	) name16506 (
		\m0_data_i[9]_pad ,
		_w9069_,
		_w9070_,
		_w18407_
	);
	LUT4 #(
		.INIT('h57df)
	) name16507 (
		_w9064_,
		_w9067_,
		_w18406_,
		_w18407_,
		_w18408_
	);
	LUT3 #(
		.INIT('h2a)
	) name16508 (
		\m1_data_i[9]_pad ,
		_w9069_,
		_w9070_,
		_w18409_
	);
	LUT3 #(
		.INIT('h80)
	) name16509 (
		\m2_data_i[9]_pad ,
		_w9069_,
		_w9070_,
		_w18410_
	);
	LUT4 #(
		.INIT('h3b7f)
	) name16510 (
		_w9064_,
		_w9067_,
		_w18409_,
		_w18410_,
		_w18411_
	);
	LUT4 #(
		.INIT('h7fff)
	) name16511 (
		_w18402_,
		_w18405_,
		_w18408_,
		_w18411_,
		_w18412_
	);
	LUT3 #(
		.INIT('h2a)
	) name16512 (
		\m3_sel_i[0]_pad ,
		_w9069_,
		_w9070_,
		_w18413_
	);
	LUT3 #(
		.INIT('h80)
	) name16513 (
		\m4_sel_i[0]_pad ,
		_w9069_,
		_w9070_,
		_w18414_
	);
	LUT4 #(
		.INIT('h9dbf)
	) name16514 (
		_w9064_,
		_w9067_,
		_w18413_,
		_w18414_,
		_w18415_
	);
	LUT3 #(
		.INIT('h80)
	) name16515 (
		\m6_sel_i[0]_pad ,
		_w9069_,
		_w9070_,
		_w18416_
	);
	LUT3 #(
		.INIT('h80)
	) name16516 (
		\m2_sel_i[0]_pad ,
		_w9069_,
		_w9070_,
		_w18417_
	);
	LUT4 #(
		.INIT('habef)
	) name16517 (
		_w9064_,
		_w9067_,
		_w18416_,
		_w18417_,
		_w18418_
	);
	LUT3 #(
		.INIT('h2a)
	) name16518 (
		\m5_sel_i[0]_pad ,
		_w9069_,
		_w9070_,
		_w18419_
	);
	LUT3 #(
		.INIT('h2a)
	) name16519 (
		\m1_sel_i[0]_pad ,
		_w9069_,
		_w9070_,
		_w18420_
	);
	LUT4 #(
		.INIT('h57df)
	) name16520 (
		_w9064_,
		_w9067_,
		_w18419_,
		_w18420_,
		_w18421_
	);
	LUT3 #(
		.INIT('h80)
	) name16521 (
		\m0_sel_i[0]_pad ,
		_w9069_,
		_w9070_,
		_w18422_
	);
	LUT3 #(
		.INIT('h2a)
	) name16522 (
		\m7_sel_i[0]_pad ,
		_w9069_,
		_w9070_,
		_w18423_
	);
	LUT4 #(
		.INIT('h6e7f)
	) name16523 (
		_w9064_,
		_w9067_,
		_w18422_,
		_w18423_,
		_w18424_
	);
	LUT4 #(
		.INIT('h7fff)
	) name16524 (
		_w18415_,
		_w18418_,
		_w18421_,
		_w18424_,
		_w18425_
	);
	LUT3 #(
		.INIT('h2a)
	) name16525 (
		\m3_sel_i[1]_pad ,
		_w9069_,
		_w9070_,
		_w18426_
	);
	LUT3 #(
		.INIT('h80)
	) name16526 (
		\m4_sel_i[1]_pad ,
		_w9069_,
		_w9070_,
		_w18427_
	);
	LUT4 #(
		.INIT('h9dbf)
	) name16527 (
		_w9064_,
		_w9067_,
		_w18426_,
		_w18427_,
		_w18428_
	);
	LUT3 #(
		.INIT('h80)
	) name16528 (
		\m6_sel_i[1]_pad ,
		_w9069_,
		_w9070_,
		_w18429_
	);
	LUT3 #(
		.INIT('h80)
	) name16529 (
		\m2_sel_i[1]_pad ,
		_w9069_,
		_w9070_,
		_w18430_
	);
	LUT4 #(
		.INIT('habef)
	) name16530 (
		_w9064_,
		_w9067_,
		_w18429_,
		_w18430_,
		_w18431_
	);
	LUT3 #(
		.INIT('h2a)
	) name16531 (
		\m5_sel_i[1]_pad ,
		_w9069_,
		_w9070_,
		_w18432_
	);
	LUT3 #(
		.INIT('h2a)
	) name16532 (
		\m1_sel_i[1]_pad ,
		_w9069_,
		_w9070_,
		_w18433_
	);
	LUT4 #(
		.INIT('h57df)
	) name16533 (
		_w9064_,
		_w9067_,
		_w18432_,
		_w18433_,
		_w18434_
	);
	LUT3 #(
		.INIT('h80)
	) name16534 (
		\m0_sel_i[1]_pad ,
		_w9069_,
		_w9070_,
		_w18435_
	);
	LUT3 #(
		.INIT('h2a)
	) name16535 (
		\m7_sel_i[1]_pad ,
		_w9069_,
		_w9070_,
		_w18436_
	);
	LUT4 #(
		.INIT('h6e7f)
	) name16536 (
		_w9064_,
		_w9067_,
		_w18435_,
		_w18436_,
		_w18437_
	);
	LUT4 #(
		.INIT('h7fff)
	) name16537 (
		_w18428_,
		_w18431_,
		_w18434_,
		_w18437_,
		_w18438_
	);
	LUT3 #(
		.INIT('h80)
	) name16538 (
		\m6_sel_i[2]_pad ,
		_w9069_,
		_w9070_,
		_w18439_
	);
	LUT3 #(
		.INIT('h2a)
	) name16539 (
		\m5_sel_i[2]_pad ,
		_w9069_,
		_w9070_,
		_w18440_
	);
	LUT4 #(
		.INIT('hcdef)
	) name16540 (
		_w9064_,
		_w9067_,
		_w18439_,
		_w18440_,
		_w18441_
	);
	LUT3 #(
		.INIT('h80)
	) name16541 (
		\m0_sel_i[2]_pad ,
		_w9069_,
		_w9070_,
		_w18442_
	);
	LUT3 #(
		.INIT('h80)
	) name16542 (
		\m4_sel_i[2]_pad ,
		_w9069_,
		_w9070_,
		_w18443_
	);
	LUT4 #(
		.INIT('h5d7f)
	) name16543 (
		_w9064_,
		_w9067_,
		_w18442_,
		_w18443_,
		_w18444_
	);
	LUT3 #(
		.INIT('h2a)
	) name16544 (
		\m7_sel_i[2]_pad ,
		_w9069_,
		_w9070_,
		_w18445_
	);
	LUT3 #(
		.INIT('h2a)
	) name16545 (
		\m3_sel_i[2]_pad ,
		_w9069_,
		_w9070_,
		_w18446_
	);
	LUT4 #(
		.INIT('habef)
	) name16546 (
		_w9064_,
		_w9067_,
		_w18445_,
		_w18446_,
		_w18447_
	);
	LUT3 #(
		.INIT('h2a)
	) name16547 (
		\m1_sel_i[2]_pad ,
		_w9069_,
		_w9070_,
		_w18448_
	);
	LUT3 #(
		.INIT('h80)
	) name16548 (
		\m2_sel_i[2]_pad ,
		_w9069_,
		_w9070_,
		_w18449_
	);
	LUT4 #(
		.INIT('h3b7f)
	) name16549 (
		_w9064_,
		_w9067_,
		_w18448_,
		_w18449_,
		_w18450_
	);
	LUT4 #(
		.INIT('h7fff)
	) name16550 (
		_w18441_,
		_w18444_,
		_w18447_,
		_w18450_,
		_w18451_
	);
	LUT3 #(
		.INIT('h80)
	) name16551 (
		\m6_sel_i[3]_pad ,
		_w9069_,
		_w9070_,
		_w18452_
	);
	LUT3 #(
		.INIT('h2a)
	) name16552 (
		\m5_sel_i[3]_pad ,
		_w9069_,
		_w9070_,
		_w18453_
	);
	LUT4 #(
		.INIT('hcdef)
	) name16553 (
		_w9064_,
		_w9067_,
		_w18452_,
		_w18453_,
		_w18454_
	);
	LUT3 #(
		.INIT('h80)
	) name16554 (
		\m0_sel_i[3]_pad ,
		_w9069_,
		_w9070_,
		_w18455_
	);
	LUT3 #(
		.INIT('h80)
	) name16555 (
		\m4_sel_i[3]_pad ,
		_w9069_,
		_w9070_,
		_w18456_
	);
	LUT4 #(
		.INIT('h5d7f)
	) name16556 (
		_w9064_,
		_w9067_,
		_w18455_,
		_w18456_,
		_w18457_
	);
	LUT3 #(
		.INIT('h2a)
	) name16557 (
		\m7_sel_i[3]_pad ,
		_w9069_,
		_w9070_,
		_w18458_
	);
	LUT3 #(
		.INIT('h2a)
	) name16558 (
		\m3_sel_i[3]_pad ,
		_w9069_,
		_w9070_,
		_w18459_
	);
	LUT4 #(
		.INIT('habef)
	) name16559 (
		_w9064_,
		_w9067_,
		_w18458_,
		_w18459_,
		_w18460_
	);
	LUT3 #(
		.INIT('h2a)
	) name16560 (
		\m1_sel_i[3]_pad ,
		_w9069_,
		_w9070_,
		_w18461_
	);
	LUT3 #(
		.INIT('h80)
	) name16561 (
		\m2_sel_i[3]_pad ,
		_w9069_,
		_w9070_,
		_w18462_
	);
	LUT4 #(
		.INIT('h3b7f)
	) name16562 (
		_w9064_,
		_w9067_,
		_w18461_,
		_w18462_,
		_w18463_
	);
	LUT4 #(
		.INIT('h7fff)
	) name16563 (
		_w18454_,
		_w18457_,
		_w18460_,
		_w18463_,
		_w18464_
	);
	LUT4 #(
		.INIT('h2a00)
	) name16564 (
		\m3_stb_i_pad ,
		_w9069_,
		_w9070_,
		_w9489_,
		_w18465_
	);
	LUT4 #(
		.INIT('h8000)
	) name16565 (
		\m2_stb_i_pad ,
		_w9069_,
		_w9070_,
		_w9629_,
		_w18466_
	);
	LUT3 #(
		.INIT('h57)
	) name16566 (
		_w9082_,
		_w18465_,
		_w18466_,
		_w18467_
	);
	LUT4 #(
		.INIT('h8000)
	) name16567 (
		\m6_stb_i_pad ,
		_w9069_,
		_w9070_,
		_w9568_,
		_w18468_
	);
	LUT4 #(
		.INIT('h2a00)
	) name16568 (
		\m7_stb_i_pad ,
		_w9069_,
		_w9070_,
		_w9600_,
		_w18469_
	);
	LUT3 #(
		.INIT('h57)
	) name16569 (
		_w9068_,
		_w18468_,
		_w18469_,
		_w18470_
	);
	LUT4 #(
		.INIT('h2a00)
	) name16570 (
		\m1_stb_i_pad ,
		_w9069_,
		_w9070_,
		_w9419_,
		_w18471_
	);
	LUT4 #(
		.INIT('h2a00)
	) name16571 (
		\m5_stb_i_pad ,
		_w9069_,
		_w9070_,
		_w9538_,
		_w18472_
	);
	LUT4 #(
		.INIT('h5d7f)
	) name16572 (
		_w9064_,
		_w9067_,
		_w18471_,
		_w18472_,
		_w18473_
	);
	LUT4 #(
		.INIT('h8000)
	) name16573 (
		\m4_stb_i_pad ,
		_w9069_,
		_w9070_,
		_w9369_,
		_w18474_
	);
	LUT4 #(
		.INIT('h8000)
	) name16574 (
		\m0_stb_i_pad ,
		_w9069_,
		_w9070_,
		_w9647_,
		_w18475_
	);
	LUT4 #(
		.INIT('h57df)
	) name16575 (
		_w9064_,
		_w9067_,
		_w18474_,
		_w18475_,
		_w18476_
	);
	LUT4 #(
		.INIT('h7fff)
	) name16576 (
		_w18467_,
		_w18470_,
		_w18473_,
		_w18476_,
		_w18477_
	);
	LUT3 #(
		.INIT('h2a)
	) name16577 (
		\m3_we_i_pad ,
		_w9069_,
		_w9070_,
		_w18478_
	);
	LUT3 #(
		.INIT('h80)
	) name16578 (
		\m4_we_i_pad ,
		_w9069_,
		_w9070_,
		_w18479_
	);
	LUT4 #(
		.INIT('h9dbf)
	) name16579 (
		_w9064_,
		_w9067_,
		_w18478_,
		_w18479_,
		_w18480_
	);
	LUT3 #(
		.INIT('h80)
	) name16580 (
		\m6_we_i_pad ,
		_w9069_,
		_w9070_,
		_w18481_
	);
	LUT3 #(
		.INIT('h80)
	) name16581 (
		\m2_we_i_pad ,
		_w9069_,
		_w9070_,
		_w18482_
	);
	LUT4 #(
		.INIT('habef)
	) name16582 (
		_w9064_,
		_w9067_,
		_w18481_,
		_w18482_,
		_w18483_
	);
	LUT3 #(
		.INIT('h2a)
	) name16583 (
		\m5_we_i_pad ,
		_w9069_,
		_w9070_,
		_w18484_
	);
	LUT3 #(
		.INIT('h2a)
	) name16584 (
		\m1_we_i_pad ,
		_w9069_,
		_w9070_,
		_w18485_
	);
	LUT4 #(
		.INIT('h57df)
	) name16585 (
		_w9064_,
		_w9067_,
		_w18484_,
		_w18485_,
		_w18486_
	);
	LUT3 #(
		.INIT('h80)
	) name16586 (
		\m0_we_i_pad ,
		_w9069_,
		_w9070_,
		_w18487_
	);
	LUT3 #(
		.INIT('h2a)
	) name16587 (
		\m7_we_i_pad ,
		_w9069_,
		_w9070_,
		_w18488_
	);
	LUT4 #(
		.INIT('h6e7f)
	) name16588 (
		_w9064_,
		_w9067_,
		_w18487_,
		_w18488_,
		_w18489_
	);
	LUT4 #(
		.INIT('h7fff)
	) name16589 (
		_w18480_,
		_w18483_,
		_w18486_,
		_w18489_,
		_w18490_
	);
	LUT3 #(
		.INIT('h2a)
	) name16590 (
		\m3_addr_i[0]_pad ,
		_w9137_,
		_w9138_,
		_w18491_
	);
	LUT3 #(
		.INIT('h80)
	) name16591 (
		\m4_addr_i[0]_pad ,
		_w9137_,
		_w9138_,
		_w18492_
	);
	LUT4 #(
		.INIT('h9bdf)
	) name16592 (
		_w9132_,
		_w9135_,
		_w18491_,
		_w18492_,
		_w18493_
	);
	LUT3 #(
		.INIT('h80)
	) name16593 (
		\m6_addr_i[0]_pad ,
		_w9137_,
		_w9138_,
		_w18494_
	);
	LUT3 #(
		.INIT('h80)
	) name16594 (
		\m2_addr_i[0]_pad ,
		_w9137_,
		_w9138_,
		_w18495_
	);
	LUT4 #(
		.INIT('hcdef)
	) name16595 (
		_w9132_,
		_w9135_,
		_w18494_,
		_w18495_,
		_w18496_
	);
	LUT3 #(
		.INIT('h2a)
	) name16596 (
		\m5_addr_i[0]_pad ,
		_w9137_,
		_w9138_,
		_w18497_
	);
	LUT3 #(
		.INIT('h2a)
	) name16597 (
		\m1_addr_i[0]_pad ,
		_w9137_,
		_w9138_,
		_w18498_
	);
	LUT4 #(
		.INIT('h37bf)
	) name16598 (
		_w9132_,
		_w9135_,
		_w18497_,
		_w18498_,
		_w18499_
	);
	LUT3 #(
		.INIT('h80)
	) name16599 (
		\m0_addr_i[0]_pad ,
		_w9137_,
		_w9138_,
		_w18500_
	);
	LUT3 #(
		.INIT('h2a)
	) name16600 (
		\m7_addr_i[0]_pad ,
		_w9137_,
		_w9138_,
		_w18501_
	);
	LUT4 #(
		.INIT('h6e7f)
	) name16601 (
		_w9132_,
		_w9135_,
		_w18500_,
		_w18501_,
		_w18502_
	);
	LUT4 #(
		.INIT('h7fff)
	) name16602 (
		_w18493_,
		_w18496_,
		_w18499_,
		_w18502_,
		_w18503_
	);
	LUT3 #(
		.INIT('h2a)
	) name16603 (
		\m1_addr_i[10]_pad ,
		_w9137_,
		_w9138_,
		_w18504_
	);
	LUT3 #(
		.INIT('h80)
	) name16604 (
		\m2_addr_i[10]_pad ,
		_w9137_,
		_w9138_,
		_w18505_
	);
	LUT4 #(
		.INIT('h5d7f)
	) name16605 (
		_w9132_,
		_w9135_,
		_w18504_,
		_w18505_,
		_w18506_
	);
	LUT3 #(
		.INIT('h80)
	) name16606 (
		\m6_addr_i[10]_pad ,
		_w9137_,
		_w9138_,
		_w18507_
	);
	LUT3 #(
		.INIT('h2a)
	) name16607 (
		\m7_addr_i[10]_pad ,
		_w9137_,
		_w9138_,
		_w18508_
	);
	LUT3 #(
		.INIT('h57)
	) name16608 (
		_w9150_,
		_w18507_,
		_w18508_,
		_w18509_
	);
	LUT3 #(
		.INIT('h2a)
	) name16609 (
		\m5_addr_i[10]_pad ,
		_w9137_,
		_w9138_,
		_w18510_
	);
	LUT3 #(
		.INIT('h80)
	) name16610 (
		\m0_addr_i[10]_pad ,
		_w9137_,
		_w9138_,
		_w18511_
	);
	LUT4 #(
		.INIT('h37bf)
	) name16611 (
		_w9132_,
		_w9135_,
		_w18510_,
		_w18511_,
		_w18512_
	);
	LUT3 #(
		.INIT('h2a)
	) name16612 (
		\m3_addr_i[10]_pad ,
		_w9137_,
		_w9138_,
		_w18513_
	);
	LUT3 #(
		.INIT('h80)
	) name16613 (
		\m4_addr_i[10]_pad ,
		_w9137_,
		_w9138_,
		_w18514_
	);
	LUT4 #(
		.INIT('h9bdf)
	) name16614 (
		_w9132_,
		_w9135_,
		_w18513_,
		_w18514_,
		_w18515_
	);
	LUT4 #(
		.INIT('h7fff)
	) name16615 (
		_w18506_,
		_w18509_,
		_w18512_,
		_w18515_,
		_w18516_
	);
	LUT3 #(
		.INIT('h2a)
	) name16616 (
		\m3_addr_i[11]_pad ,
		_w9137_,
		_w9138_,
		_w18517_
	);
	LUT3 #(
		.INIT('h80)
	) name16617 (
		\m4_addr_i[11]_pad ,
		_w9137_,
		_w9138_,
		_w18518_
	);
	LUT4 #(
		.INIT('h9bdf)
	) name16618 (
		_w9132_,
		_w9135_,
		_w18517_,
		_w18518_,
		_w18519_
	);
	LUT3 #(
		.INIT('h80)
	) name16619 (
		\m6_addr_i[11]_pad ,
		_w9137_,
		_w9138_,
		_w18520_
	);
	LUT3 #(
		.INIT('h80)
	) name16620 (
		\m2_addr_i[11]_pad ,
		_w9137_,
		_w9138_,
		_w18521_
	);
	LUT4 #(
		.INIT('hcdef)
	) name16621 (
		_w9132_,
		_w9135_,
		_w18520_,
		_w18521_,
		_w18522_
	);
	LUT3 #(
		.INIT('h2a)
	) name16622 (
		\m5_addr_i[11]_pad ,
		_w9137_,
		_w9138_,
		_w18523_
	);
	LUT3 #(
		.INIT('h2a)
	) name16623 (
		\m1_addr_i[11]_pad ,
		_w9137_,
		_w9138_,
		_w18524_
	);
	LUT4 #(
		.INIT('h37bf)
	) name16624 (
		_w9132_,
		_w9135_,
		_w18523_,
		_w18524_,
		_w18525_
	);
	LUT3 #(
		.INIT('h80)
	) name16625 (
		\m0_addr_i[11]_pad ,
		_w9137_,
		_w9138_,
		_w18526_
	);
	LUT3 #(
		.INIT('h2a)
	) name16626 (
		\m7_addr_i[11]_pad ,
		_w9137_,
		_w9138_,
		_w18527_
	);
	LUT4 #(
		.INIT('h6e7f)
	) name16627 (
		_w9132_,
		_w9135_,
		_w18526_,
		_w18527_,
		_w18528_
	);
	LUT4 #(
		.INIT('h7fff)
	) name16628 (
		_w18519_,
		_w18522_,
		_w18525_,
		_w18528_,
		_w18529_
	);
	LUT3 #(
		.INIT('h2a)
	) name16629 (
		\m3_addr_i[12]_pad ,
		_w9137_,
		_w9138_,
		_w18530_
	);
	LUT3 #(
		.INIT('h80)
	) name16630 (
		\m4_addr_i[12]_pad ,
		_w9137_,
		_w9138_,
		_w18531_
	);
	LUT4 #(
		.INIT('h9bdf)
	) name16631 (
		_w9132_,
		_w9135_,
		_w18530_,
		_w18531_,
		_w18532_
	);
	LUT3 #(
		.INIT('h80)
	) name16632 (
		\m6_addr_i[12]_pad ,
		_w9137_,
		_w9138_,
		_w18533_
	);
	LUT3 #(
		.INIT('h80)
	) name16633 (
		\m2_addr_i[12]_pad ,
		_w9137_,
		_w9138_,
		_w18534_
	);
	LUT4 #(
		.INIT('hcdef)
	) name16634 (
		_w9132_,
		_w9135_,
		_w18533_,
		_w18534_,
		_w18535_
	);
	LUT3 #(
		.INIT('h2a)
	) name16635 (
		\m5_addr_i[12]_pad ,
		_w9137_,
		_w9138_,
		_w18536_
	);
	LUT3 #(
		.INIT('h2a)
	) name16636 (
		\m1_addr_i[12]_pad ,
		_w9137_,
		_w9138_,
		_w18537_
	);
	LUT4 #(
		.INIT('h37bf)
	) name16637 (
		_w9132_,
		_w9135_,
		_w18536_,
		_w18537_,
		_w18538_
	);
	LUT3 #(
		.INIT('h80)
	) name16638 (
		\m0_addr_i[12]_pad ,
		_w9137_,
		_w9138_,
		_w18539_
	);
	LUT3 #(
		.INIT('h2a)
	) name16639 (
		\m7_addr_i[12]_pad ,
		_w9137_,
		_w9138_,
		_w18540_
	);
	LUT4 #(
		.INIT('h6e7f)
	) name16640 (
		_w9132_,
		_w9135_,
		_w18539_,
		_w18540_,
		_w18541_
	);
	LUT4 #(
		.INIT('h7fff)
	) name16641 (
		_w18532_,
		_w18535_,
		_w18538_,
		_w18541_,
		_w18542_
	);
	LUT3 #(
		.INIT('h2a)
	) name16642 (
		\m3_addr_i[13]_pad ,
		_w9137_,
		_w9138_,
		_w18543_
	);
	LUT3 #(
		.INIT('h80)
	) name16643 (
		\m4_addr_i[13]_pad ,
		_w9137_,
		_w9138_,
		_w18544_
	);
	LUT4 #(
		.INIT('h9bdf)
	) name16644 (
		_w9132_,
		_w9135_,
		_w18543_,
		_w18544_,
		_w18545_
	);
	LUT3 #(
		.INIT('h80)
	) name16645 (
		\m6_addr_i[13]_pad ,
		_w9137_,
		_w9138_,
		_w18546_
	);
	LUT3 #(
		.INIT('h80)
	) name16646 (
		\m2_addr_i[13]_pad ,
		_w9137_,
		_w9138_,
		_w18547_
	);
	LUT4 #(
		.INIT('hcdef)
	) name16647 (
		_w9132_,
		_w9135_,
		_w18546_,
		_w18547_,
		_w18548_
	);
	LUT3 #(
		.INIT('h2a)
	) name16648 (
		\m5_addr_i[13]_pad ,
		_w9137_,
		_w9138_,
		_w18549_
	);
	LUT3 #(
		.INIT('h2a)
	) name16649 (
		\m1_addr_i[13]_pad ,
		_w9137_,
		_w9138_,
		_w18550_
	);
	LUT4 #(
		.INIT('h37bf)
	) name16650 (
		_w9132_,
		_w9135_,
		_w18549_,
		_w18550_,
		_w18551_
	);
	LUT3 #(
		.INIT('h80)
	) name16651 (
		\m0_addr_i[13]_pad ,
		_w9137_,
		_w9138_,
		_w18552_
	);
	LUT3 #(
		.INIT('h2a)
	) name16652 (
		\m7_addr_i[13]_pad ,
		_w9137_,
		_w9138_,
		_w18553_
	);
	LUT4 #(
		.INIT('h6e7f)
	) name16653 (
		_w9132_,
		_w9135_,
		_w18552_,
		_w18553_,
		_w18554_
	);
	LUT4 #(
		.INIT('h7fff)
	) name16654 (
		_w18545_,
		_w18548_,
		_w18551_,
		_w18554_,
		_w18555_
	);
	LUT3 #(
		.INIT('h2a)
	) name16655 (
		\m1_addr_i[14]_pad ,
		_w9137_,
		_w9138_,
		_w18556_
	);
	LUT3 #(
		.INIT('h80)
	) name16656 (
		\m2_addr_i[14]_pad ,
		_w9137_,
		_w9138_,
		_w18557_
	);
	LUT4 #(
		.INIT('h5d7f)
	) name16657 (
		_w9132_,
		_w9135_,
		_w18556_,
		_w18557_,
		_w18558_
	);
	LUT3 #(
		.INIT('h80)
	) name16658 (
		\m6_addr_i[14]_pad ,
		_w9137_,
		_w9138_,
		_w18559_
	);
	LUT3 #(
		.INIT('h2a)
	) name16659 (
		\m7_addr_i[14]_pad ,
		_w9137_,
		_w9138_,
		_w18560_
	);
	LUT3 #(
		.INIT('h57)
	) name16660 (
		_w9150_,
		_w18559_,
		_w18560_,
		_w18561_
	);
	LUT3 #(
		.INIT('h2a)
	) name16661 (
		\m5_addr_i[14]_pad ,
		_w9137_,
		_w9138_,
		_w18562_
	);
	LUT3 #(
		.INIT('h80)
	) name16662 (
		\m0_addr_i[14]_pad ,
		_w9137_,
		_w9138_,
		_w18563_
	);
	LUT4 #(
		.INIT('h37bf)
	) name16663 (
		_w9132_,
		_w9135_,
		_w18562_,
		_w18563_,
		_w18564_
	);
	LUT3 #(
		.INIT('h2a)
	) name16664 (
		\m3_addr_i[14]_pad ,
		_w9137_,
		_w9138_,
		_w18565_
	);
	LUT3 #(
		.INIT('h80)
	) name16665 (
		\m4_addr_i[14]_pad ,
		_w9137_,
		_w9138_,
		_w18566_
	);
	LUT4 #(
		.INIT('h9bdf)
	) name16666 (
		_w9132_,
		_w9135_,
		_w18565_,
		_w18566_,
		_w18567_
	);
	LUT4 #(
		.INIT('h7fff)
	) name16667 (
		_w18558_,
		_w18561_,
		_w18564_,
		_w18567_,
		_w18568_
	);
	LUT3 #(
		.INIT('h80)
	) name16668 (
		\m6_addr_i[15]_pad ,
		_w9137_,
		_w9138_,
		_w18569_
	);
	LUT3 #(
		.INIT('h2a)
	) name16669 (
		\m5_addr_i[15]_pad ,
		_w9137_,
		_w9138_,
		_w18570_
	);
	LUT4 #(
		.INIT('habef)
	) name16670 (
		_w9132_,
		_w9135_,
		_w18569_,
		_w18570_,
		_w18571_
	);
	LUT3 #(
		.INIT('h80)
	) name16671 (
		\m0_addr_i[15]_pad ,
		_w9137_,
		_w9138_,
		_w18572_
	);
	LUT3 #(
		.INIT('h80)
	) name16672 (
		\m4_addr_i[15]_pad ,
		_w9137_,
		_w9138_,
		_w18573_
	);
	LUT4 #(
		.INIT('h3b7f)
	) name16673 (
		_w9132_,
		_w9135_,
		_w18572_,
		_w18573_,
		_w18574_
	);
	LUT3 #(
		.INIT('h2a)
	) name16674 (
		\m7_addr_i[15]_pad ,
		_w9137_,
		_w9138_,
		_w18575_
	);
	LUT3 #(
		.INIT('h2a)
	) name16675 (
		\m3_addr_i[15]_pad ,
		_w9137_,
		_w9138_,
		_w18576_
	);
	LUT4 #(
		.INIT('hcdef)
	) name16676 (
		_w9132_,
		_w9135_,
		_w18575_,
		_w18576_,
		_w18577_
	);
	LUT3 #(
		.INIT('h2a)
	) name16677 (
		\m1_addr_i[15]_pad ,
		_w9137_,
		_w9138_,
		_w18578_
	);
	LUT3 #(
		.INIT('h80)
	) name16678 (
		\m2_addr_i[15]_pad ,
		_w9137_,
		_w9138_,
		_w18579_
	);
	LUT4 #(
		.INIT('h5d7f)
	) name16679 (
		_w9132_,
		_w9135_,
		_w18578_,
		_w18579_,
		_w18580_
	);
	LUT4 #(
		.INIT('h7fff)
	) name16680 (
		_w18571_,
		_w18574_,
		_w18577_,
		_w18580_,
		_w18581_
	);
	LUT3 #(
		.INIT('h2a)
	) name16681 (
		\m3_addr_i[16]_pad ,
		_w9137_,
		_w9138_,
		_w18582_
	);
	LUT3 #(
		.INIT('h80)
	) name16682 (
		\m4_addr_i[16]_pad ,
		_w9137_,
		_w9138_,
		_w18583_
	);
	LUT4 #(
		.INIT('h9bdf)
	) name16683 (
		_w9132_,
		_w9135_,
		_w18582_,
		_w18583_,
		_w18584_
	);
	LUT3 #(
		.INIT('h80)
	) name16684 (
		\m6_addr_i[16]_pad ,
		_w9137_,
		_w9138_,
		_w18585_
	);
	LUT3 #(
		.INIT('h2a)
	) name16685 (
		\m7_addr_i[16]_pad ,
		_w9137_,
		_w9138_,
		_w18586_
	);
	LUT3 #(
		.INIT('h57)
	) name16686 (
		_w9150_,
		_w18585_,
		_w18586_,
		_w18587_
	);
	LUT3 #(
		.INIT('h2a)
	) name16687 (
		\m5_addr_i[16]_pad ,
		_w9137_,
		_w9138_,
		_w18588_
	);
	LUT3 #(
		.INIT('h80)
	) name16688 (
		\m0_addr_i[16]_pad ,
		_w9137_,
		_w9138_,
		_w18589_
	);
	LUT4 #(
		.INIT('h37bf)
	) name16689 (
		_w9132_,
		_w9135_,
		_w18588_,
		_w18589_,
		_w18590_
	);
	LUT3 #(
		.INIT('h2a)
	) name16690 (
		\m1_addr_i[16]_pad ,
		_w9137_,
		_w9138_,
		_w18591_
	);
	LUT3 #(
		.INIT('h80)
	) name16691 (
		\m2_addr_i[16]_pad ,
		_w9137_,
		_w9138_,
		_w18592_
	);
	LUT4 #(
		.INIT('h5d7f)
	) name16692 (
		_w9132_,
		_w9135_,
		_w18591_,
		_w18592_,
		_w18593_
	);
	LUT4 #(
		.INIT('h7fff)
	) name16693 (
		_w18584_,
		_w18587_,
		_w18590_,
		_w18593_,
		_w18594_
	);
	LUT3 #(
		.INIT('h2a)
	) name16694 (
		\m3_addr_i[17]_pad ,
		_w9137_,
		_w9138_,
		_w18595_
	);
	LUT3 #(
		.INIT('h80)
	) name16695 (
		\m4_addr_i[17]_pad ,
		_w9137_,
		_w9138_,
		_w18596_
	);
	LUT4 #(
		.INIT('h9bdf)
	) name16696 (
		_w9132_,
		_w9135_,
		_w18595_,
		_w18596_,
		_w18597_
	);
	LUT3 #(
		.INIT('h80)
	) name16697 (
		\m6_addr_i[17]_pad ,
		_w9137_,
		_w9138_,
		_w18598_
	);
	LUT3 #(
		.INIT('h80)
	) name16698 (
		\m2_addr_i[17]_pad ,
		_w9137_,
		_w9138_,
		_w18599_
	);
	LUT4 #(
		.INIT('hcdef)
	) name16699 (
		_w9132_,
		_w9135_,
		_w18598_,
		_w18599_,
		_w18600_
	);
	LUT3 #(
		.INIT('h2a)
	) name16700 (
		\m5_addr_i[17]_pad ,
		_w9137_,
		_w9138_,
		_w18601_
	);
	LUT3 #(
		.INIT('h2a)
	) name16701 (
		\m1_addr_i[17]_pad ,
		_w9137_,
		_w9138_,
		_w18602_
	);
	LUT4 #(
		.INIT('h37bf)
	) name16702 (
		_w9132_,
		_w9135_,
		_w18601_,
		_w18602_,
		_w18603_
	);
	LUT3 #(
		.INIT('h80)
	) name16703 (
		\m0_addr_i[17]_pad ,
		_w9137_,
		_w9138_,
		_w18604_
	);
	LUT3 #(
		.INIT('h2a)
	) name16704 (
		\m7_addr_i[17]_pad ,
		_w9137_,
		_w9138_,
		_w18605_
	);
	LUT4 #(
		.INIT('h6e7f)
	) name16705 (
		_w9132_,
		_w9135_,
		_w18604_,
		_w18605_,
		_w18606_
	);
	LUT4 #(
		.INIT('h7fff)
	) name16706 (
		_w18597_,
		_w18600_,
		_w18603_,
		_w18606_,
		_w18607_
	);
	LUT3 #(
		.INIT('h2a)
	) name16707 (
		\m3_addr_i[18]_pad ,
		_w9137_,
		_w9138_,
		_w18608_
	);
	LUT3 #(
		.INIT('h80)
	) name16708 (
		\m4_addr_i[18]_pad ,
		_w9137_,
		_w9138_,
		_w18609_
	);
	LUT4 #(
		.INIT('h9bdf)
	) name16709 (
		_w9132_,
		_w9135_,
		_w18608_,
		_w18609_,
		_w18610_
	);
	LUT3 #(
		.INIT('h80)
	) name16710 (
		\m6_addr_i[18]_pad ,
		_w9137_,
		_w9138_,
		_w18611_
	);
	LUT3 #(
		.INIT('h2a)
	) name16711 (
		\m7_addr_i[18]_pad ,
		_w9137_,
		_w9138_,
		_w18612_
	);
	LUT3 #(
		.INIT('h57)
	) name16712 (
		_w9150_,
		_w18611_,
		_w18612_,
		_w18613_
	);
	LUT3 #(
		.INIT('h2a)
	) name16713 (
		\m5_addr_i[18]_pad ,
		_w9137_,
		_w9138_,
		_w18614_
	);
	LUT3 #(
		.INIT('h80)
	) name16714 (
		\m0_addr_i[18]_pad ,
		_w9137_,
		_w9138_,
		_w18615_
	);
	LUT4 #(
		.INIT('h37bf)
	) name16715 (
		_w9132_,
		_w9135_,
		_w18614_,
		_w18615_,
		_w18616_
	);
	LUT3 #(
		.INIT('h2a)
	) name16716 (
		\m1_addr_i[18]_pad ,
		_w9137_,
		_w9138_,
		_w18617_
	);
	LUT3 #(
		.INIT('h80)
	) name16717 (
		\m2_addr_i[18]_pad ,
		_w9137_,
		_w9138_,
		_w18618_
	);
	LUT4 #(
		.INIT('h5d7f)
	) name16718 (
		_w9132_,
		_w9135_,
		_w18617_,
		_w18618_,
		_w18619_
	);
	LUT4 #(
		.INIT('h7fff)
	) name16719 (
		_w18610_,
		_w18613_,
		_w18616_,
		_w18619_,
		_w18620_
	);
	LUT3 #(
		.INIT('h2a)
	) name16720 (
		\m3_addr_i[19]_pad ,
		_w9137_,
		_w9138_,
		_w18621_
	);
	LUT3 #(
		.INIT('h80)
	) name16721 (
		\m4_addr_i[19]_pad ,
		_w9137_,
		_w9138_,
		_w18622_
	);
	LUT4 #(
		.INIT('h9bdf)
	) name16722 (
		_w9132_,
		_w9135_,
		_w18621_,
		_w18622_,
		_w18623_
	);
	LUT3 #(
		.INIT('h80)
	) name16723 (
		\m6_addr_i[19]_pad ,
		_w9137_,
		_w9138_,
		_w18624_
	);
	LUT3 #(
		.INIT('h80)
	) name16724 (
		\m2_addr_i[19]_pad ,
		_w9137_,
		_w9138_,
		_w18625_
	);
	LUT4 #(
		.INIT('hcdef)
	) name16725 (
		_w9132_,
		_w9135_,
		_w18624_,
		_w18625_,
		_w18626_
	);
	LUT3 #(
		.INIT('h2a)
	) name16726 (
		\m5_addr_i[19]_pad ,
		_w9137_,
		_w9138_,
		_w18627_
	);
	LUT3 #(
		.INIT('h2a)
	) name16727 (
		\m1_addr_i[19]_pad ,
		_w9137_,
		_w9138_,
		_w18628_
	);
	LUT4 #(
		.INIT('h37bf)
	) name16728 (
		_w9132_,
		_w9135_,
		_w18627_,
		_w18628_,
		_w18629_
	);
	LUT3 #(
		.INIT('h80)
	) name16729 (
		\m0_addr_i[19]_pad ,
		_w9137_,
		_w9138_,
		_w18630_
	);
	LUT3 #(
		.INIT('h2a)
	) name16730 (
		\m7_addr_i[19]_pad ,
		_w9137_,
		_w9138_,
		_w18631_
	);
	LUT4 #(
		.INIT('h6e7f)
	) name16731 (
		_w9132_,
		_w9135_,
		_w18630_,
		_w18631_,
		_w18632_
	);
	LUT4 #(
		.INIT('h7fff)
	) name16732 (
		_w18623_,
		_w18626_,
		_w18629_,
		_w18632_,
		_w18633_
	);
	LUT3 #(
		.INIT('h2a)
	) name16733 (
		\m3_addr_i[1]_pad ,
		_w9137_,
		_w9138_,
		_w18634_
	);
	LUT3 #(
		.INIT('h80)
	) name16734 (
		\m4_addr_i[1]_pad ,
		_w9137_,
		_w9138_,
		_w18635_
	);
	LUT4 #(
		.INIT('h9bdf)
	) name16735 (
		_w9132_,
		_w9135_,
		_w18634_,
		_w18635_,
		_w18636_
	);
	LUT3 #(
		.INIT('h80)
	) name16736 (
		\m6_addr_i[1]_pad ,
		_w9137_,
		_w9138_,
		_w18637_
	);
	LUT3 #(
		.INIT('h80)
	) name16737 (
		\m2_addr_i[1]_pad ,
		_w9137_,
		_w9138_,
		_w18638_
	);
	LUT4 #(
		.INIT('hcdef)
	) name16738 (
		_w9132_,
		_w9135_,
		_w18637_,
		_w18638_,
		_w18639_
	);
	LUT3 #(
		.INIT('h2a)
	) name16739 (
		\m5_addr_i[1]_pad ,
		_w9137_,
		_w9138_,
		_w18640_
	);
	LUT3 #(
		.INIT('h2a)
	) name16740 (
		\m1_addr_i[1]_pad ,
		_w9137_,
		_w9138_,
		_w18641_
	);
	LUT4 #(
		.INIT('h37bf)
	) name16741 (
		_w9132_,
		_w9135_,
		_w18640_,
		_w18641_,
		_w18642_
	);
	LUT3 #(
		.INIT('h80)
	) name16742 (
		\m0_addr_i[1]_pad ,
		_w9137_,
		_w9138_,
		_w18643_
	);
	LUT3 #(
		.INIT('h2a)
	) name16743 (
		\m7_addr_i[1]_pad ,
		_w9137_,
		_w9138_,
		_w18644_
	);
	LUT4 #(
		.INIT('h6e7f)
	) name16744 (
		_w9132_,
		_w9135_,
		_w18643_,
		_w18644_,
		_w18645_
	);
	LUT4 #(
		.INIT('h7fff)
	) name16745 (
		_w18636_,
		_w18639_,
		_w18642_,
		_w18645_,
		_w18646_
	);
	LUT3 #(
		.INIT('h2a)
	) name16746 (
		\m3_addr_i[20]_pad ,
		_w9137_,
		_w9138_,
		_w18647_
	);
	LUT3 #(
		.INIT('h80)
	) name16747 (
		\m4_addr_i[20]_pad ,
		_w9137_,
		_w9138_,
		_w18648_
	);
	LUT4 #(
		.INIT('h9bdf)
	) name16748 (
		_w9132_,
		_w9135_,
		_w18647_,
		_w18648_,
		_w18649_
	);
	LUT3 #(
		.INIT('h80)
	) name16749 (
		\m6_addr_i[20]_pad ,
		_w9137_,
		_w9138_,
		_w18650_
	);
	LUT3 #(
		.INIT('h80)
	) name16750 (
		\m2_addr_i[20]_pad ,
		_w9137_,
		_w9138_,
		_w18651_
	);
	LUT4 #(
		.INIT('hcdef)
	) name16751 (
		_w9132_,
		_w9135_,
		_w18650_,
		_w18651_,
		_w18652_
	);
	LUT3 #(
		.INIT('h2a)
	) name16752 (
		\m5_addr_i[20]_pad ,
		_w9137_,
		_w9138_,
		_w18653_
	);
	LUT3 #(
		.INIT('h2a)
	) name16753 (
		\m1_addr_i[20]_pad ,
		_w9137_,
		_w9138_,
		_w18654_
	);
	LUT4 #(
		.INIT('h37bf)
	) name16754 (
		_w9132_,
		_w9135_,
		_w18653_,
		_w18654_,
		_w18655_
	);
	LUT3 #(
		.INIT('h80)
	) name16755 (
		\m0_addr_i[20]_pad ,
		_w9137_,
		_w9138_,
		_w18656_
	);
	LUT3 #(
		.INIT('h2a)
	) name16756 (
		\m7_addr_i[20]_pad ,
		_w9137_,
		_w9138_,
		_w18657_
	);
	LUT4 #(
		.INIT('h6e7f)
	) name16757 (
		_w9132_,
		_w9135_,
		_w18656_,
		_w18657_,
		_w18658_
	);
	LUT4 #(
		.INIT('h7fff)
	) name16758 (
		_w18649_,
		_w18652_,
		_w18655_,
		_w18658_,
		_w18659_
	);
	LUT3 #(
		.INIT('h2a)
	) name16759 (
		\m3_addr_i[21]_pad ,
		_w9137_,
		_w9138_,
		_w18660_
	);
	LUT3 #(
		.INIT('h80)
	) name16760 (
		\m4_addr_i[21]_pad ,
		_w9137_,
		_w9138_,
		_w18661_
	);
	LUT4 #(
		.INIT('h9bdf)
	) name16761 (
		_w9132_,
		_w9135_,
		_w18660_,
		_w18661_,
		_w18662_
	);
	LUT3 #(
		.INIT('h80)
	) name16762 (
		\m6_addr_i[21]_pad ,
		_w9137_,
		_w9138_,
		_w18663_
	);
	LUT3 #(
		.INIT('h80)
	) name16763 (
		\m2_addr_i[21]_pad ,
		_w9137_,
		_w9138_,
		_w18664_
	);
	LUT4 #(
		.INIT('hcdef)
	) name16764 (
		_w9132_,
		_w9135_,
		_w18663_,
		_w18664_,
		_w18665_
	);
	LUT3 #(
		.INIT('h2a)
	) name16765 (
		\m5_addr_i[21]_pad ,
		_w9137_,
		_w9138_,
		_w18666_
	);
	LUT3 #(
		.INIT('h2a)
	) name16766 (
		\m1_addr_i[21]_pad ,
		_w9137_,
		_w9138_,
		_w18667_
	);
	LUT4 #(
		.INIT('h37bf)
	) name16767 (
		_w9132_,
		_w9135_,
		_w18666_,
		_w18667_,
		_w18668_
	);
	LUT3 #(
		.INIT('h80)
	) name16768 (
		\m0_addr_i[21]_pad ,
		_w9137_,
		_w9138_,
		_w18669_
	);
	LUT3 #(
		.INIT('h2a)
	) name16769 (
		\m7_addr_i[21]_pad ,
		_w9137_,
		_w9138_,
		_w18670_
	);
	LUT4 #(
		.INIT('h6e7f)
	) name16770 (
		_w9132_,
		_w9135_,
		_w18669_,
		_w18670_,
		_w18671_
	);
	LUT4 #(
		.INIT('h7fff)
	) name16771 (
		_w18662_,
		_w18665_,
		_w18668_,
		_w18671_,
		_w18672_
	);
	LUT3 #(
		.INIT('h2a)
	) name16772 (
		\m3_addr_i[22]_pad ,
		_w9137_,
		_w9138_,
		_w18673_
	);
	LUT3 #(
		.INIT('h80)
	) name16773 (
		\m4_addr_i[22]_pad ,
		_w9137_,
		_w9138_,
		_w18674_
	);
	LUT4 #(
		.INIT('h9bdf)
	) name16774 (
		_w9132_,
		_w9135_,
		_w18673_,
		_w18674_,
		_w18675_
	);
	LUT3 #(
		.INIT('h80)
	) name16775 (
		\m6_addr_i[22]_pad ,
		_w9137_,
		_w9138_,
		_w18676_
	);
	LUT3 #(
		.INIT('h80)
	) name16776 (
		\m2_addr_i[22]_pad ,
		_w9137_,
		_w9138_,
		_w18677_
	);
	LUT4 #(
		.INIT('hcdef)
	) name16777 (
		_w9132_,
		_w9135_,
		_w18676_,
		_w18677_,
		_w18678_
	);
	LUT3 #(
		.INIT('h2a)
	) name16778 (
		\m5_addr_i[22]_pad ,
		_w9137_,
		_w9138_,
		_w18679_
	);
	LUT3 #(
		.INIT('h2a)
	) name16779 (
		\m1_addr_i[22]_pad ,
		_w9137_,
		_w9138_,
		_w18680_
	);
	LUT4 #(
		.INIT('h37bf)
	) name16780 (
		_w9132_,
		_w9135_,
		_w18679_,
		_w18680_,
		_w18681_
	);
	LUT3 #(
		.INIT('h80)
	) name16781 (
		\m0_addr_i[22]_pad ,
		_w9137_,
		_w9138_,
		_w18682_
	);
	LUT3 #(
		.INIT('h2a)
	) name16782 (
		\m7_addr_i[22]_pad ,
		_w9137_,
		_w9138_,
		_w18683_
	);
	LUT4 #(
		.INIT('h6e7f)
	) name16783 (
		_w9132_,
		_w9135_,
		_w18682_,
		_w18683_,
		_w18684_
	);
	LUT4 #(
		.INIT('h7fff)
	) name16784 (
		_w18675_,
		_w18678_,
		_w18681_,
		_w18684_,
		_w18685_
	);
	LUT3 #(
		.INIT('h2a)
	) name16785 (
		\m3_addr_i[23]_pad ,
		_w9137_,
		_w9138_,
		_w18686_
	);
	LUT3 #(
		.INIT('h80)
	) name16786 (
		\m4_addr_i[23]_pad ,
		_w9137_,
		_w9138_,
		_w18687_
	);
	LUT4 #(
		.INIT('h9bdf)
	) name16787 (
		_w9132_,
		_w9135_,
		_w18686_,
		_w18687_,
		_w18688_
	);
	LUT3 #(
		.INIT('h80)
	) name16788 (
		\m6_addr_i[23]_pad ,
		_w9137_,
		_w9138_,
		_w18689_
	);
	LUT3 #(
		.INIT('h80)
	) name16789 (
		\m2_addr_i[23]_pad ,
		_w9137_,
		_w9138_,
		_w18690_
	);
	LUT4 #(
		.INIT('hcdef)
	) name16790 (
		_w9132_,
		_w9135_,
		_w18689_,
		_w18690_,
		_w18691_
	);
	LUT3 #(
		.INIT('h2a)
	) name16791 (
		\m5_addr_i[23]_pad ,
		_w9137_,
		_w9138_,
		_w18692_
	);
	LUT3 #(
		.INIT('h2a)
	) name16792 (
		\m1_addr_i[23]_pad ,
		_w9137_,
		_w9138_,
		_w18693_
	);
	LUT4 #(
		.INIT('h37bf)
	) name16793 (
		_w9132_,
		_w9135_,
		_w18692_,
		_w18693_,
		_w18694_
	);
	LUT3 #(
		.INIT('h80)
	) name16794 (
		\m0_addr_i[23]_pad ,
		_w9137_,
		_w9138_,
		_w18695_
	);
	LUT3 #(
		.INIT('h2a)
	) name16795 (
		\m7_addr_i[23]_pad ,
		_w9137_,
		_w9138_,
		_w18696_
	);
	LUT4 #(
		.INIT('h6e7f)
	) name16796 (
		_w9132_,
		_w9135_,
		_w18695_,
		_w18696_,
		_w18697_
	);
	LUT4 #(
		.INIT('h7fff)
	) name16797 (
		_w18688_,
		_w18691_,
		_w18694_,
		_w18697_,
		_w18698_
	);
	LUT3 #(
		.INIT('h2a)
	) name16798 (
		\m3_addr_i[24]_pad ,
		_w9137_,
		_w9138_,
		_w18699_
	);
	LUT3 #(
		.INIT('h80)
	) name16799 (
		\m4_addr_i[24]_pad ,
		_w9137_,
		_w9138_,
		_w18700_
	);
	LUT4 #(
		.INIT('h9bdf)
	) name16800 (
		_w9132_,
		_w9135_,
		_w18699_,
		_w18700_,
		_w18701_
	);
	LUT3 #(
		.INIT('h2a)
	) name16801 (
		\m5_addr_i[24]_pad ,
		_w9137_,
		_w9138_,
		_w18702_
	);
	LUT3 #(
		.INIT('h80)
	) name16802 (
		\m2_addr_i[24]_pad ,
		_w9137_,
		_w9138_,
		_w18703_
	);
	LUT4 #(
		.INIT('h9dbf)
	) name16803 (
		_w9132_,
		_w9135_,
		_w18702_,
		_w18703_,
		_w18704_
	);
	LUT3 #(
		.INIT('h80)
	) name16804 (
		\m6_addr_i[24]_pad ,
		_w9137_,
		_w9138_,
		_w18705_
	);
	LUT3 #(
		.INIT('h2a)
	) name16805 (
		\m1_addr_i[24]_pad ,
		_w9137_,
		_w9138_,
		_w18706_
	);
	LUT4 #(
		.INIT('h67ef)
	) name16806 (
		_w9132_,
		_w9135_,
		_w18705_,
		_w18706_,
		_w18707_
	);
	LUT3 #(
		.INIT('h80)
	) name16807 (
		\m0_addr_i[24]_pad ,
		_w9137_,
		_w9138_,
		_w18708_
	);
	LUT3 #(
		.INIT('h2a)
	) name16808 (
		\m7_addr_i[24]_pad ,
		_w9137_,
		_w9138_,
		_w18709_
	);
	LUT4 #(
		.INIT('h6e7f)
	) name16809 (
		_w9132_,
		_w9135_,
		_w18708_,
		_w18709_,
		_w18710_
	);
	LUT4 #(
		.INIT('h7fff)
	) name16810 (
		_w18701_,
		_w18704_,
		_w18707_,
		_w18710_,
		_w18711_
	);
	LUT3 #(
		.INIT('h2a)
	) name16811 (
		\m3_addr_i[25]_pad ,
		_w9137_,
		_w9138_,
		_w18712_
	);
	LUT3 #(
		.INIT('h80)
	) name16812 (
		\m4_addr_i[25]_pad ,
		_w9137_,
		_w9138_,
		_w18713_
	);
	LUT4 #(
		.INIT('h9bdf)
	) name16813 (
		_w9132_,
		_w9135_,
		_w18712_,
		_w18713_,
		_w18714_
	);
	LUT3 #(
		.INIT('h2a)
	) name16814 (
		\m5_addr_i[25]_pad ,
		_w9137_,
		_w9138_,
		_w18715_
	);
	LUT3 #(
		.INIT('h80)
	) name16815 (
		\m2_addr_i[25]_pad ,
		_w9137_,
		_w9138_,
		_w18716_
	);
	LUT4 #(
		.INIT('h9dbf)
	) name16816 (
		_w9132_,
		_w9135_,
		_w18715_,
		_w18716_,
		_w18717_
	);
	LUT3 #(
		.INIT('h80)
	) name16817 (
		\m6_addr_i[25]_pad ,
		_w9137_,
		_w9138_,
		_w18718_
	);
	LUT3 #(
		.INIT('h2a)
	) name16818 (
		\m1_addr_i[25]_pad ,
		_w9137_,
		_w9138_,
		_w18719_
	);
	LUT4 #(
		.INIT('h67ef)
	) name16819 (
		_w9132_,
		_w9135_,
		_w18718_,
		_w18719_,
		_w18720_
	);
	LUT3 #(
		.INIT('h80)
	) name16820 (
		\m0_addr_i[25]_pad ,
		_w9137_,
		_w9138_,
		_w18721_
	);
	LUT3 #(
		.INIT('h2a)
	) name16821 (
		\m7_addr_i[25]_pad ,
		_w9137_,
		_w9138_,
		_w18722_
	);
	LUT4 #(
		.INIT('h6e7f)
	) name16822 (
		_w9132_,
		_w9135_,
		_w18721_,
		_w18722_,
		_w18723_
	);
	LUT4 #(
		.INIT('h7fff)
	) name16823 (
		_w18714_,
		_w18717_,
		_w18720_,
		_w18723_,
		_w18724_
	);
	LUT3 #(
		.INIT('h2a)
	) name16824 (
		\m3_addr_i[26]_pad ,
		_w9137_,
		_w9138_,
		_w18725_
	);
	LUT3 #(
		.INIT('h80)
	) name16825 (
		\m4_addr_i[26]_pad ,
		_w9137_,
		_w9138_,
		_w18726_
	);
	LUT4 #(
		.INIT('h9bdf)
	) name16826 (
		_w9132_,
		_w9135_,
		_w18725_,
		_w18726_,
		_w18727_
	);
	LUT3 #(
		.INIT('h2a)
	) name16827 (
		\m5_addr_i[26]_pad ,
		_w9137_,
		_w9138_,
		_w18728_
	);
	LUT3 #(
		.INIT('h80)
	) name16828 (
		\m2_addr_i[26]_pad ,
		_w9137_,
		_w9138_,
		_w18729_
	);
	LUT4 #(
		.INIT('h9dbf)
	) name16829 (
		_w9132_,
		_w9135_,
		_w18728_,
		_w18729_,
		_w18730_
	);
	LUT3 #(
		.INIT('h80)
	) name16830 (
		\m6_addr_i[26]_pad ,
		_w9137_,
		_w9138_,
		_w18731_
	);
	LUT3 #(
		.INIT('h2a)
	) name16831 (
		\m1_addr_i[26]_pad ,
		_w9137_,
		_w9138_,
		_w18732_
	);
	LUT4 #(
		.INIT('h67ef)
	) name16832 (
		_w9132_,
		_w9135_,
		_w18731_,
		_w18732_,
		_w18733_
	);
	LUT3 #(
		.INIT('h80)
	) name16833 (
		\m0_addr_i[26]_pad ,
		_w9137_,
		_w9138_,
		_w18734_
	);
	LUT3 #(
		.INIT('h2a)
	) name16834 (
		\m7_addr_i[26]_pad ,
		_w9137_,
		_w9138_,
		_w18735_
	);
	LUT4 #(
		.INIT('h6e7f)
	) name16835 (
		_w9132_,
		_w9135_,
		_w18734_,
		_w18735_,
		_w18736_
	);
	LUT4 #(
		.INIT('h7fff)
	) name16836 (
		_w18727_,
		_w18730_,
		_w18733_,
		_w18736_,
		_w18737_
	);
	LUT3 #(
		.INIT('h2a)
	) name16837 (
		\m3_addr_i[27]_pad ,
		_w9137_,
		_w9138_,
		_w18738_
	);
	LUT3 #(
		.INIT('h80)
	) name16838 (
		\m4_addr_i[27]_pad ,
		_w9137_,
		_w9138_,
		_w18739_
	);
	LUT4 #(
		.INIT('h9bdf)
	) name16839 (
		_w9132_,
		_w9135_,
		_w18738_,
		_w18739_,
		_w18740_
	);
	LUT3 #(
		.INIT('h2a)
	) name16840 (
		\m5_addr_i[27]_pad ,
		_w9137_,
		_w9138_,
		_w18741_
	);
	LUT3 #(
		.INIT('h80)
	) name16841 (
		\m2_addr_i[27]_pad ,
		_w9137_,
		_w9138_,
		_w18742_
	);
	LUT4 #(
		.INIT('h9dbf)
	) name16842 (
		_w9132_,
		_w9135_,
		_w18741_,
		_w18742_,
		_w18743_
	);
	LUT3 #(
		.INIT('h80)
	) name16843 (
		\m6_addr_i[27]_pad ,
		_w9137_,
		_w9138_,
		_w18744_
	);
	LUT3 #(
		.INIT('h2a)
	) name16844 (
		\m1_addr_i[27]_pad ,
		_w9137_,
		_w9138_,
		_w18745_
	);
	LUT4 #(
		.INIT('h67ef)
	) name16845 (
		_w9132_,
		_w9135_,
		_w18744_,
		_w18745_,
		_w18746_
	);
	LUT3 #(
		.INIT('h80)
	) name16846 (
		\m0_addr_i[27]_pad ,
		_w9137_,
		_w9138_,
		_w18747_
	);
	LUT3 #(
		.INIT('h2a)
	) name16847 (
		\m7_addr_i[27]_pad ,
		_w9137_,
		_w9138_,
		_w18748_
	);
	LUT4 #(
		.INIT('h6e7f)
	) name16848 (
		_w9132_,
		_w9135_,
		_w18747_,
		_w18748_,
		_w18749_
	);
	LUT4 #(
		.INIT('h7fff)
	) name16849 (
		_w18740_,
		_w18743_,
		_w18746_,
		_w18749_,
		_w18750_
	);
	LUT3 #(
		.INIT('h2a)
	) name16850 (
		\m3_addr_i[28]_pad ,
		_w9137_,
		_w9138_,
		_w18751_
	);
	LUT3 #(
		.INIT('h80)
	) name16851 (
		\m4_addr_i[28]_pad ,
		_w9137_,
		_w9138_,
		_w18752_
	);
	LUT4 #(
		.INIT('h9bdf)
	) name16852 (
		_w9132_,
		_w9135_,
		_w18751_,
		_w18752_,
		_w18753_
	);
	LUT3 #(
		.INIT('h2a)
	) name16853 (
		\m5_addr_i[28]_pad ,
		_w9137_,
		_w9138_,
		_w18754_
	);
	LUT3 #(
		.INIT('h80)
	) name16854 (
		\m2_addr_i[28]_pad ,
		_w9137_,
		_w9138_,
		_w18755_
	);
	LUT4 #(
		.INIT('h9dbf)
	) name16855 (
		_w9132_,
		_w9135_,
		_w18754_,
		_w18755_,
		_w18756_
	);
	LUT3 #(
		.INIT('h80)
	) name16856 (
		\m6_addr_i[28]_pad ,
		_w9137_,
		_w9138_,
		_w18757_
	);
	LUT3 #(
		.INIT('h2a)
	) name16857 (
		\m1_addr_i[28]_pad ,
		_w9137_,
		_w9138_,
		_w18758_
	);
	LUT4 #(
		.INIT('h67ef)
	) name16858 (
		_w9132_,
		_w9135_,
		_w18757_,
		_w18758_,
		_w18759_
	);
	LUT3 #(
		.INIT('h80)
	) name16859 (
		\m0_addr_i[28]_pad ,
		_w9137_,
		_w9138_,
		_w18760_
	);
	LUT3 #(
		.INIT('h2a)
	) name16860 (
		\m7_addr_i[28]_pad ,
		_w9137_,
		_w9138_,
		_w18761_
	);
	LUT4 #(
		.INIT('h6e7f)
	) name16861 (
		_w9132_,
		_w9135_,
		_w18760_,
		_w18761_,
		_w18762_
	);
	LUT4 #(
		.INIT('h7fff)
	) name16862 (
		_w18753_,
		_w18756_,
		_w18759_,
		_w18762_,
		_w18763_
	);
	LUT3 #(
		.INIT('h2a)
	) name16863 (
		\m3_addr_i[29]_pad ,
		_w9137_,
		_w9138_,
		_w18764_
	);
	LUT3 #(
		.INIT('h80)
	) name16864 (
		\m4_addr_i[29]_pad ,
		_w9137_,
		_w9138_,
		_w18765_
	);
	LUT4 #(
		.INIT('h9bdf)
	) name16865 (
		_w9132_,
		_w9135_,
		_w18764_,
		_w18765_,
		_w18766_
	);
	LUT3 #(
		.INIT('h2a)
	) name16866 (
		\m5_addr_i[29]_pad ,
		_w9137_,
		_w9138_,
		_w18767_
	);
	LUT3 #(
		.INIT('h80)
	) name16867 (
		\m2_addr_i[29]_pad ,
		_w9137_,
		_w9138_,
		_w18768_
	);
	LUT4 #(
		.INIT('h9dbf)
	) name16868 (
		_w9132_,
		_w9135_,
		_w18767_,
		_w18768_,
		_w18769_
	);
	LUT3 #(
		.INIT('h80)
	) name16869 (
		\m6_addr_i[29]_pad ,
		_w9137_,
		_w9138_,
		_w18770_
	);
	LUT3 #(
		.INIT('h2a)
	) name16870 (
		\m1_addr_i[29]_pad ,
		_w9137_,
		_w9138_,
		_w18771_
	);
	LUT4 #(
		.INIT('h67ef)
	) name16871 (
		_w9132_,
		_w9135_,
		_w18770_,
		_w18771_,
		_w18772_
	);
	LUT3 #(
		.INIT('h80)
	) name16872 (
		\m0_addr_i[29]_pad ,
		_w9137_,
		_w9138_,
		_w18773_
	);
	LUT3 #(
		.INIT('h2a)
	) name16873 (
		\m7_addr_i[29]_pad ,
		_w9137_,
		_w9138_,
		_w18774_
	);
	LUT4 #(
		.INIT('h6e7f)
	) name16874 (
		_w9132_,
		_w9135_,
		_w18773_,
		_w18774_,
		_w18775_
	);
	LUT4 #(
		.INIT('h7fff)
	) name16875 (
		_w18766_,
		_w18769_,
		_w18772_,
		_w18775_,
		_w18776_
	);
	LUT3 #(
		.INIT('h80)
	) name16876 (
		\m6_addr_i[2]_pad ,
		_w9137_,
		_w9138_,
		_w18777_
	);
	LUT3 #(
		.INIT('h2a)
	) name16877 (
		\m5_addr_i[2]_pad ,
		_w9137_,
		_w9138_,
		_w18778_
	);
	LUT4 #(
		.INIT('habef)
	) name16878 (
		_w9132_,
		_w9135_,
		_w18777_,
		_w18778_,
		_w18779_
	);
	LUT3 #(
		.INIT('h80)
	) name16879 (
		\m0_addr_i[2]_pad ,
		_w9137_,
		_w9138_,
		_w18780_
	);
	LUT3 #(
		.INIT('h80)
	) name16880 (
		\m4_addr_i[2]_pad ,
		_w9137_,
		_w9138_,
		_w18781_
	);
	LUT4 #(
		.INIT('h3b7f)
	) name16881 (
		_w9132_,
		_w9135_,
		_w18780_,
		_w18781_,
		_w18782_
	);
	LUT3 #(
		.INIT('h2a)
	) name16882 (
		\m7_addr_i[2]_pad ,
		_w9137_,
		_w9138_,
		_w18783_
	);
	LUT3 #(
		.INIT('h2a)
	) name16883 (
		\m3_addr_i[2]_pad ,
		_w9137_,
		_w9138_,
		_w18784_
	);
	LUT4 #(
		.INIT('hcdef)
	) name16884 (
		_w9132_,
		_w9135_,
		_w18783_,
		_w18784_,
		_w18785_
	);
	LUT3 #(
		.INIT('h2a)
	) name16885 (
		\m1_addr_i[2]_pad ,
		_w9137_,
		_w9138_,
		_w18786_
	);
	LUT3 #(
		.INIT('h80)
	) name16886 (
		\m2_addr_i[2]_pad ,
		_w9137_,
		_w9138_,
		_w18787_
	);
	LUT4 #(
		.INIT('h5d7f)
	) name16887 (
		_w9132_,
		_w9135_,
		_w18786_,
		_w18787_,
		_w18788_
	);
	LUT4 #(
		.INIT('h7fff)
	) name16888 (
		_w18779_,
		_w18782_,
		_w18785_,
		_w18788_,
		_w18789_
	);
	LUT3 #(
		.INIT('h2a)
	) name16889 (
		\m3_addr_i[30]_pad ,
		_w9137_,
		_w9138_,
		_w18790_
	);
	LUT3 #(
		.INIT('h80)
	) name16890 (
		\m4_addr_i[30]_pad ,
		_w9137_,
		_w9138_,
		_w18791_
	);
	LUT4 #(
		.INIT('h9bdf)
	) name16891 (
		_w9132_,
		_w9135_,
		_w18790_,
		_w18791_,
		_w18792_
	);
	LUT3 #(
		.INIT('h2a)
	) name16892 (
		\m5_addr_i[30]_pad ,
		_w9137_,
		_w9138_,
		_w18793_
	);
	LUT3 #(
		.INIT('h80)
	) name16893 (
		\m2_addr_i[30]_pad ,
		_w9137_,
		_w9138_,
		_w18794_
	);
	LUT4 #(
		.INIT('h9dbf)
	) name16894 (
		_w9132_,
		_w9135_,
		_w18793_,
		_w18794_,
		_w18795_
	);
	LUT3 #(
		.INIT('h80)
	) name16895 (
		\m6_addr_i[30]_pad ,
		_w9137_,
		_w9138_,
		_w18796_
	);
	LUT3 #(
		.INIT('h2a)
	) name16896 (
		\m1_addr_i[30]_pad ,
		_w9137_,
		_w9138_,
		_w18797_
	);
	LUT4 #(
		.INIT('h67ef)
	) name16897 (
		_w9132_,
		_w9135_,
		_w18796_,
		_w18797_,
		_w18798_
	);
	LUT3 #(
		.INIT('h80)
	) name16898 (
		\m0_addr_i[30]_pad ,
		_w9137_,
		_w9138_,
		_w18799_
	);
	LUT3 #(
		.INIT('h2a)
	) name16899 (
		\m7_addr_i[30]_pad ,
		_w9137_,
		_w9138_,
		_w18800_
	);
	LUT4 #(
		.INIT('h6e7f)
	) name16900 (
		_w9132_,
		_w9135_,
		_w18799_,
		_w18800_,
		_w18801_
	);
	LUT4 #(
		.INIT('h7fff)
	) name16901 (
		_w18792_,
		_w18795_,
		_w18798_,
		_w18801_,
		_w18802_
	);
	LUT3 #(
		.INIT('h2a)
	) name16902 (
		\m3_addr_i[31]_pad ,
		_w9137_,
		_w9138_,
		_w18803_
	);
	LUT3 #(
		.INIT('h80)
	) name16903 (
		\m4_addr_i[31]_pad ,
		_w9137_,
		_w9138_,
		_w18804_
	);
	LUT4 #(
		.INIT('h9bdf)
	) name16904 (
		_w9132_,
		_w9135_,
		_w18803_,
		_w18804_,
		_w18805_
	);
	LUT3 #(
		.INIT('h2a)
	) name16905 (
		\m5_addr_i[31]_pad ,
		_w9137_,
		_w9138_,
		_w18806_
	);
	LUT3 #(
		.INIT('h80)
	) name16906 (
		\m2_addr_i[31]_pad ,
		_w9137_,
		_w9138_,
		_w18807_
	);
	LUT4 #(
		.INIT('h9dbf)
	) name16907 (
		_w9132_,
		_w9135_,
		_w18806_,
		_w18807_,
		_w18808_
	);
	LUT3 #(
		.INIT('h80)
	) name16908 (
		\m6_addr_i[31]_pad ,
		_w9137_,
		_w9138_,
		_w18809_
	);
	LUT3 #(
		.INIT('h2a)
	) name16909 (
		\m1_addr_i[31]_pad ,
		_w9137_,
		_w9138_,
		_w18810_
	);
	LUT4 #(
		.INIT('h67ef)
	) name16910 (
		_w9132_,
		_w9135_,
		_w18809_,
		_w18810_,
		_w18811_
	);
	LUT3 #(
		.INIT('h80)
	) name16911 (
		\m0_addr_i[31]_pad ,
		_w9137_,
		_w9138_,
		_w18812_
	);
	LUT3 #(
		.INIT('h2a)
	) name16912 (
		\m7_addr_i[31]_pad ,
		_w9137_,
		_w9138_,
		_w18813_
	);
	LUT4 #(
		.INIT('h6e7f)
	) name16913 (
		_w9132_,
		_w9135_,
		_w18812_,
		_w18813_,
		_w18814_
	);
	LUT4 #(
		.INIT('h7fff)
	) name16914 (
		_w18805_,
		_w18808_,
		_w18811_,
		_w18814_,
		_w18815_
	);
	LUT3 #(
		.INIT('h2a)
	) name16915 (
		\m3_addr_i[3]_pad ,
		_w9137_,
		_w9138_,
		_w18816_
	);
	LUT3 #(
		.INIT('h80)
	) name16916 (
		\m4_addr_i[3]_pad ,
		_w9137_,
		_w9138_,
		_w18817_
	);
	LUT4 #(
		.INIT('h9bdf)
	) name16917 (
		_w9132_,
		_w9135_,
		_w18816_,
		_w18817_,
		_w18818_
	);
	LUT3 #(
		.INIT('h80)
	) name16918 (
		\m6_addr_i[3]_pad ,
		_w9137_,
		_w9138_,
		_w18819_
	);
	LUT3 #(
		.INIT('h80)
	) name16919 (
		\m2_addr_i[3]_pad ,
		_w9137_,
		_w9138_,
		_w18820_
	);
	LUT4 #(
		.INIT('hcdef)
	) name16920 (
		_w9132_,
		_w9135_,
		_w18819_,
		_w18820_,
		_w18821_
	);
	LUT3 #(
		.INIT('h2a)
	) name16921 (
		\m5_addr_i[3]_pad ,
		_w9137_,
		_w9138_,
		_w18822_
	);
	LUT3 #(
		.INIT('h2a)
	) name16922 (
		\m1_addr_i[3]_pad ,
		_w9137_,
		_w9138_,
		_w18823_
	);
	LUT4 #(
		.INIT('h37bf)
	) name16923 (
		_w9132_,
		_w9135_,
		_w18822_,
		_w18823_,
		_w18824_
	);
	LUT3 #(
		.INIT('h80)
	) name16924 (
		\m0_addr_i[3]_pad ,
		_w9137_,
		_w9138_,
		_w18825_
	);
	LUT3 #(
		.INIT('h2a)
	) name16925 (
		\m7_addr_i[3]_pad ,
		_w9137_,
		_w9138_,
		_w18826_
	);
	LUT4 #(
		.INIT('h6e7f)
	) name16926 (
		_w9132_,
		_w9135_,
		_w18825_,
		_w18826_,
		_w18827_
	);
	LUT4 #(
		.INIT('h7fff)
	) name16927 (
		_w18818_,
		_w18821_,
		_w18824_,
		_w18827_,
		_w18828_
	);
	LUT3 #(
		.INIT('h80)
	) name16928 (
		\m6_addr_i[4]_pad ,
		_w9137_,
		_w9138_,
		_w18829_
	);
	LUT3 #(
		.INIT('h2a)
	) name16929 (
		\m5_addr_i[4]_pad ,
		_w9137_,
		_w9138_,
		_w18830_
	);
	LUT4 #(
		.INIT('habef)
	) name16930 (
		_w9132_,
		_w9135_,
		_w18829_,
		_w18830_,
		_w18831_
	);
	LUT3 #(
		.INIT('h80)
	) name16931 (
		\m0_addr_i[4]_pad ,
		_w9137_,
		_w9138_,
		_w18832_
	);
	LUT3 #(
		.INIT('h80)
	) name16932 (
		\m4_addr_i[4]_pad ,
		_w9137_,
		_w9138_,
		_w18833_
	);
	LUT4 #(
		.INIT('h3b7f)
	) name16933 (
		_w9132_,
		_w9135_,
		_w18832_,
		_w18833_,
		_w18834_
	);
	LUT3 #(
		.INIT('h2a)
	) name16934 (
		\m7_addr_i[4]_pad ,
		_w9137_,
		_w9138_,
		_w18835_
	);
	LUT3 #(
		.INIT('h2a)
	) name16935 (
		\m3_addr_i[4]_pad ,
		_w9137_,
		_w9138_,
		_w18836_
	);
	LUT4 #(
		.INIT('hcdef)
	) name16936 (
		_w9132_,
		_w9135_,
		_w18835_,
		_w18836_,
		_w18837_
	);
	LUT3 #(
		.INIT('h2a)
	) name16937 (
		\m1_addr_i[4]_pad ,
		_w9137_,
		_w9138_,
		_w18838_
	);
	LUT3 #(
		.INIT('h80)
	) name16938 (
		\m2_addr_i[4]_pad ,
		_w9137_,
		_w9138_,
		_w18839_
	);
	LUT4 #(
		.INIT('h5d7f)
	) name16939 (
		_w9132_,
		_w9135_,
		_w18838_,
		_w18839_,
		_w18840_
	);
	LUT4 #(
		.INIT('h7fff)
	) name16940 (
		_w18831_,
		_w18834_,
		_w18837_,
		_w18840_,
		_w18841_
	);
	LUT3 #(
		.INIT('h2a)
	) name16941 (
		\m3_addr_i[5]_pad ,
		_w9137_,
		_w9138_,
		_w18842_
	);
	LUT3 #(
		.INIT('h80)
	) name16942 (
		\m4_addr_i[5]_pad ,
		_w9137_,
		_w9138_,
		_w18843_
	);
	LUT4 #(
		.INIT('h9bdf)
	) name16943 (
		_w9132_,
		_w9135_,
		_w18842_,
		_w18843_,
		_w18844_
	);
	LUT3 #(
		.INIT('h80)
	) name16944 (
		\m6_addr_i[5]_pad ,
		_w9137_,
		_w9138_,
		_w18845_
	);
	LUT3 #(
		.INIT('h80)
	) name16945 (
		\m2_addr_i[5]_pad ,
		_w9137_,
		_w9138_,
		_w18846_
	);
	LUT4 #(
		.INIT('hcdef)
	) name16946 (
		_w9132_,
		_w9135_,
		_w18845_,
		_w18846_,
		_w18847_
	);
	LUT3 #(
		.INIT('h2a)
	) name16947 (
		\m5_addr_i[5]_pad ,
		_w9137_,
		_w9138_,
		_w18848_
	);
	LUT3 #(
		.INIT('h2a)
	) name16948 (
		\m1_addr_i[5]_pad ,
		_w9137_,
		_w9138_,
		_w18849_
	);
	LUT4 #(
		.INIT('h37bf)
	) name16949 (
		_w9132_,
		_w9135_,
		_w18848_,
		_w18849_,
		_w18850_
	);
	LUT3 #(
		.INIT('h80)
	) name16950 (
		\m0_addr_i[5]_pad ,
		_w9137_,
		_w9138_,
		_w18851_
	);
	LUT3 #(
		.INIT('h2a)
	) name16951 (
		\m7_addr_i[5]_pad ,
		_w9137_,
		_w9138_,
		_w18852_
	);
	LUT4 #(
		.INIT('h6e7f)
	) name16952 (
		_w9132_,
		_w9135_,
		_w18851_,
		_w18852_,
		_w18853_
	);
	LUT4 #(
		.INIT('h7fff)
	) name16953 (
		_w18844_,
		_w18847_,
		_w18850_,
		_w18853_,
		_w18854_
	);
	LUT3 #(
		.INIT('h2a)
	) name16954 (
		\m3_addr_i[6]_pad ,
		_w9137_,
		_w9138_,
		_w18855_
	);
	LUT3 #(
		.INIT('h80)
	) name16955 (
		\m4_addr_i[6]_pad ,
		_w9137_,
		_w9138_,
		_w18856_
	);
	LUT4 #(
		.INIT('h9bdf)
	) name16956 (
		_w9132_,
		_w9135_,
		_w18855_,
		_w18856_,
		_w18857_
	);
	LUT3 #(
		.INIT('h80)
	) name16957 (
		\m6_addr_i[6]_pad ,
		_w9137_,
		_w9138_,
		_w18858_
	);
	LUT3 #(
		.INIT('h80)
	) name16958 (
		\m2_addr_i[6]_pad ,
		_w9137_,
		_w9138_,
		_w18859_
	);
	LUT4 #(
		.INIT('hcdef)
	) name16959 (
		_w9132_,
		_w9135_,
		_w18858_,
		_w18859_,
		_w18860_
	);
	LUT3 #(
		.INIT('h2a)
	) name16960 (
		\m5_addr_i[6]_pad ,
		_w9137_,
		_w9138_,
		_w18861_
	);
	LUT3 #(
		.INIT('h2a)
	) name16961 (
		\m1_addr_i[6]_pad ,
		_w9137_,
		_w9138_,
		_w18862_
	);
	LUT4 #(
		.INIT('h37bf)
	) name16962 (
		_w9132_,
		_w9135_,
		_w18861_,
		_w18862_,
		_w18863_
	);
	LUT3 #(
		.INIT('h80)
	) name16963 (
		\m0_addr_i[6]_pad ,
		_w9137_,
		_w9138_,
		_w18864_
	);
	LUT3 #(
		.INIT('h2a)
	) name16964 (
		\m7_addr_i[6]_pad ,
		_w9137_,
		_w9138_,
		_w18865_
	);
	LUT4 #(
		.INIT('h6e7f)
	) name16965 (
		_w9132_,
		_w9135_,
		_w18864_,
		_w18865_,
		_w18866_
	);
	LUT4 #(
		.INIT('h7fff)
	) name16966 (
		_w18857_,
		_w18860_,
		_w18863_,
		_w18866_,
		_w18867_
	);
	LUT3 #(
		.INIT('h2a)
	) name16967 (
		\m3_addr_i[7]_pad ,
		_w9137_,
		_w9138_,
		_w18868_
	);
	LUT3 #(
		.INIT('h80)
	) name16968 (
		\m4_addr_i[7]_pad ,
		_w9137_,
		_w9138_,
		_w18869_
	);
	LUT4 #(
		.INIT('h9bdf)
	) name16969 (
		_w9132_,
		_w9135_,
		_w18868_,
		_w18869_,
		_w18870_
	);
	LUT3 #(
		.INIT('h80)
	) name16970 (
		\m6_addr_i[7]_pad ,
		_w9137_,
		_w9138_,
		_w18871_
	);
	LUT3 #(
		.INIT('h80)
	) name16971 (
		\m2_addr_i[7]_pad ,
		_w9137_,
		_w9138_,
		_w18872_
	);
	LUT4 #(
		.INIT('hcdef)
	) name16972 (
		_w9132_,
		_w9135_,
		_w18871_,
		_w18872_,
		_w18873_
	);
	LUT3 #(
		.INIT('h2a)
	) name16973 (
		\m5_addr_i[7]_pad ,
		_w9137_,
		_w9138_,
		_w18874_
	);
	LUT3 #(
		.INIT('h2a)
	) name16974 (
		\m1_addr_i[7]_pad ,
		_w9137_,
		_w9138_,
		_w18875_
	);
	LUT4 #(
		.INIT('h37bf)
	) name16975 (
		_w9132_,
		_w9135_,
		_w18874_,
		_w18875_,
		_w18876_
	);
	LUT3 #(
		.INIT('h80)
	) name16976 (
		\m0_addr_i[7]_pad ,
		_w9137_,
		_w9138_,
		_w18877_
	);
	LUT3 #(
		.INIT('h2a)
	) name16977 (
		\m7_addr_i[7]_pad ,
		_w9137_,
		_w9138_,
		_w18878_
	);
	LUT4 #(
		.INIT('h6e7f)
	) name16978 (
		_w9132_,
		_w9135_,
		_w18877_,
		_w18878_,
		_w18879_
	);
	LUT4 #(
		.INIT('h7fff)
	) name16979 (
		_w18870_,
		_w18873_,
		_w18876_,
		_w18879_,
		_w18880_
	);
	LUT3 #(
		.INIT('h2a)
	) name16980 (
		\m3_addr_i[8]_pad ,
		_w9137_,
		_w9138_,
		_w18881_
	);
	LUT3 #(
		.INIT('h80)
	) name16981 (
		\m4_addr_i[8]_pad ,
		_w9137_,
		_w9138_,
		_w18882_
	);
	LUT4 #(
		.INIT('h9bdf)
	) name16982 (
		_w9132_,
		_w9135_,
		_w18881_,
		_w18882_,
		_w18883_
	);
	LUT3 #(
		.INIT('h80)
	) name16983 (
		\m6_addr_i[8]_pad ,
		_w9137_,
		_w9138_,
		_w18884_
	);
	LUT3 #(
		.INIT('h80)
	) name16984 (
		\m2_addr_i[8]_pad ,
		_w9137_,
		_w9138_,
		_w18885_
	);
	LUT4 #(
		.INIT('hcdef)
	) name16985 (
		_w9132_,
		_w9135_,
		_w18884_,
		_w18885_,
		_w18886_
	);
	LUT3 #(
		.INIT('h2a)
	) name16986 (
		\m5_addr_i[8]_pad ,
		_w9137_,
		_w9138_,
		_w18887_
	);
	LUT3 #(
		.INIT('h2a)
	) name16987 (
		\m1_addr_i[8]_pad ,
		_w9137_,
		_w9138_,
		_w18888_
	);
	LUT4 #(
		.INIT('h37bf)
	) name16988 (
		_w9132_,
		_w9135_,
		_w18887_,
		_w18888_,
		_w18889_
	);
	LUT3 #(
		.INIT('h80)
	) name16989 (
		\m0_addr_i[8]_pad ,
		_w9137_,
		_w9138_,
		_w18890_
	);
	LUT3 #(
		.INIT('h2a)
	) name16990 (
		\m7_addr_i[8]_pad ,
		_w9137_,
		_w9138_,
		_w18891_
	);
	LUT4 #(
		.INIT('h6e7f)
	) name16991 (
		_w9132_,
		_w9135_,
		_w18890_,
		_w18891_,
		_w18892_
	);
	LUT4 #(
		.INIT('h7fff)
	) name16992 (
		_w18883_,
		_w18886_,
		_w18889_,
		_w18892_,
		_w18893_
	);
	LUT3 #(
		.INIT('h2a)
	) name16993 (
		\m3_addr_i[9]_pad ,
		_w9137_,
		_w9138_,
		_w18894_
	);
	LUT3 #(
		.INIT('h80)
	) name16994 (
		\m4_addr_i[9]_pad ,
		_w9137_,
		_w9138_,
		_w18895_
	);
	LUT4 #(
		.INIT('h9bdf)
	) name16995 (
		_w9132_,
		_w9135_,
		_w18894_,
		_w18895_,
		_w18896_
	);
	LUT3 #(
		.INIT('h80)
	) name16996 (
		\m6_addr_i[9]_pad ,
		_w9137_,
		_w9138_,
		_w18897_
	);
	LUT3 #(
		.INIT('h80)
	) name16997 (
		\m2_addr_i[9]_pad ,
		_w9137_,
		_w9138_,
		_w18898_
	);
	LUT4 #(
		.INIT('hcdef)
	) name16998 (
		_w9132_,
		_w9135_,
		_w18897_,
		_w18898_,
		_w18899_
	);
	LUT3 #(
		.INIT('h2a)
	) name16999 (
		\m5_addr_i[9]_pad ,
		_w9137_,
		_w9138_,
		_w18900_
	);
	LUT3 #(
		.INIT('h2a)
	) name17000 (
		\m1_addr_i[9]_pad ,
		_w9137_,
		_w9138_,
		_w18901_
	);
	LUT4 #(
		.INIT('h37bf)
	) name17001 (
		_w9132_,
		_w9135_,
		_w18900_,
		_w18901_,
		_w18902_
	);
	LUT3 #(
		.INIT('h80)
	) name17002 (
		\m0_addr_i[9]_pad ,
		_w9137_,
		_w9138_,
		_w18903_
	);
	LUT3 #(
		.INIT('h2a)
	) name17003 (
		\m7_addr_i[9]_pad ,
		_w9137_,
		_w9138_,
		_w18904_
	);
	LUT4 #(
		.INIT('h6e7f)
	) name17004 (
		_w9132_,
		_w9135_,
		_w18903_,
		_w18904_,
		_w18905_
	);
	LUT4 #(
		.INIT('h7fff)
	) name17005 (
		_w18896_,
		_w18899_,
		_w18902_,
		_w18905_,
		_w18906_
	);
	LUT3 #(
		.INIT('h2a)
	) name17006 (
		\m3_data_i[0]_pad ,
		_w9137_,
		_w9138_,
		_w18907_
	);
	LUT3 #(
		.INIT('h80)
	) name17007 (
		\m4_data_i[0]_pad ,
		_w9137_,
		_w9138_,
		_w18908_
	);
	LUT4 #(
		.INIT('h9bdf)
	) name17008 (
		_w9132_,
		_w9135_,
		_w18907_,
		_w18908_,
		_w18909_
	);
	LUT3 #(
		.INIT('h80)
	) name17009 (
		\m6_data_i[0]_pad ,
		_w9137_,
		_w9138_,
		_w18910_
	);
	LUT3 #(
		.INIT('h80)
	) name17010 (
		\m2_data_i[0]_pad ,
		_w9137_,
		_w9138_,
		_w18911_
	);
	LUT4 #(
		.INIT('hcdef)
	) name17011 (
		_w9132_,
		_w9135_,
		_w18910_,
		_w18911_,
		_w18912_
	);
	LUT3 #(
		.INIT('h2a)
	) name17012 (
		\m5_data_i[0]_pad ,
		_w9137_,
		_w9138_,
		_w18913_
	);
	LUT3 #(
		.INIT('h2a)
	) name17013 (
		\m1_data_i[0]_pad ,
		_w9137_,
		_w9138_,
		_w18914_
	);
	LUT4 #(
		.INIT('h37bf)
	) name17014 (
		_w9132_,
		_w9135_,
		_w18913_,
		_w18914_,
		_w18915_
	);
	LUT3 #(
		.INIT('h80)
	) name17015 (
		\m0_data_i[0]_pad ,
		_w9137_,
		_w9138_,
		_w18916_
	);
	LUT3 #(
		.INIT('h2a)
	) name17016 (
		\m7_data_i[0]_pad ,
		_w9137_,
		_w9138_,
		_w18917_
	);
	LUT4 #(
		.INIT('h6e7f)
	) name17017 (
		_w9132_,
		_w9135_,
		_w18916_,
		_w18917_,
		_w18918_
	);
	LUT4 #(
		.INIT('h7fff)
	) name17018 (
		_w18909_,
		_w18912_,
		_w18915_,
		_w18918_,
		_w18919_
	);
	LUT3 #(
		.INIT('h2a)
	) name17019 (
		\m3_data_i[10]_pad ,
		_w9137_,
		_w9138_,
		_w18920_
	);
	LUT3 #(
		.INIT('h80)
	) name17020 (
		\m4_data_i[10]_pad ,
		_w9137_,
		_w9138_,
		_w18921_
	);
	LUT4 #(
		.INIT('h9bdf)
	) name17021 (
		_w9132_,
		_w9135_,
		_w18920_,
		_w18921_,
		_w18922_
	);
	LUT3 #(
		.INIT('h80)
	) name17022 (
		\m6_data_i[10]_pad ,
		_w9137_,
		_w9138_,
		_w18923_
	);
	LUT3 #(
		.INIT('h2a)
	) name17023 (
		\m7_data_i[10]_pad ,
		_w9137_,
		_w9138_,
		_w18924_
	);
	LUT3 #(
		.INIT('h57)
	) name17024 (
		_w9150_,
		_w18923_,
		_w18924_,
		_w18925_
	);
	LUT3 #(
		.INIT('h2a)
	) name17025 (
		\m5_data_i[10]_pad ,
		_w9137_,
		_w9138_,
		_w18926_
	);
	LUT3 #(
		.INIT('h80)
	) name17026 (
		\m0_data_i[10]_pad ,
		_w9137_,
		_w9138_,
		_w18927_
	);
	LUT4 #(
		.INIT('h37bf)
	) name17027 (
		_w9132_,
		_w9135_,
		_w18926_,
		_w18927_,
		_w18928_
	);
	LUT3 #(
		.INIT('h2a)
	) name17028 (
		\m1_data_i[10]_pad ,
		_w9137_,
		_w9138_,
		_w18929_
	);
	LUT3 #(
		.INIT('h80)
	) name17029 (
		\m2_data_i[10]_pad ,
		_w9137_,
		_w9138_,
		_w18930_
	);
	LUT4 #(
		.INIT('h5d7f)
	) name17030 (
		_w9132_,
		_w9135_,
		_w18929_,
		_w18930_,
		_w18931_
	);
	LUT4 #(
		.INIT('h7fff)
	) name17031 (
		_w18922_,
		_w18925_,
		_w18928_,
		_w18931_,
		_w18932_
	);
	LUT3 #(
		.INIT('h2a)
	) name17032 (
		\m3_data_i[11]_pad ,
		_w9137_,
		_w9138_,
		_w18933_
	);
	LUT3 #(
		.INIT('h80)
	) name17033 (
		\m4_data_i[11]_pad ,
		_w9137_,
		_w9138_,
		_w18934_
	);
	LUT4 #(
		.INIT('h9bdf)
	) name17034 (
		_w9132_,
		_w9135_,
		_w18933_,
		_w18934_,
		_w18935_
	);
	LUT3 #(
		.INIT('h80)
	) name17035 (
		\m6_data_i[11]_pad ,
		_w9137_,
		_w9138_,
		_w18936_
	);
	LUT3 #(
		.INIT('h80)
	) name17036 (
		\m2_data_i[11]_pad ,
		_w9137_,
		_w9138_,
		_w18937_
	);
	LUT4 #(
		.INIT('hcdef)
	) name17037 (
		_w9132_,
		_w9135_,
		_w18936_,
		_w18937_,
		_w18938_
	);
	LUT3 #(
		.INIT('h2a)
	) name17038 (
		\m5_data_i[11]_pad ,
		_w9137_,
		_w9138_,
		_w18939_
	);
	LUT3 #(
		.INIT('h2a)
	) name17039 (
		\m1_data_i[11]_pad ,
		_w9137_,
		_w9138_,
		_w18940_
	);
	LUT4 #(
		.INIT('h37bf)
	) name17040 (
		_w9132_,
		_w9135_,
		_w18939_,
		_w18940_,
		_w18941_
	);
	LUT3 #(
		.INIT('h80)
	) name17041 (
		\m0_data_i[11]_pad ,
		_w9137_,
		_w9138_,
		_w18942_
	);
	LUT3 #(
		.INIT('h2a)
	) name17042 (
		\m7_data_i[11]_pad ,
		_w9137_,
		_w9138_,
		_w18943_
	);
	LUT4 #(
		.INIT('h6e7f)
	) name17043 (
		_w9132_,
		_w9135_,
		_w18942_,
		_w18943_,
		_w18944_
	);
	LUT4 #(
		.INIT('h7fff)
	) name17044 (
		_w18935_,
		_w18938_,
		_w18941_,
		_w18944_,
		_w18945_
	);
	LUT3 #(
		.INIT('h2a)
	) name17045 (
		\m3_data_i[12]_pad ,
		_w9137_,
		_w9138_,
		_w18946_
	);
	LUT3 #(
		.INIT('h80)
	) name17046 (
		\m4_data_i[12]_pad ,
		_w9137_,
		_w9138_,
		_w18947_
	);
	LUT4 #(
		.INIT('h9bdf)
	) name17047 (
		_w9132_,
		_w9135_,
		_w18946_,
		_w18947_,
		_w18948_
	);
	LUT3 #(
		.INIT('h80)
	) name17048 (
		\m6_data_i[12]_pad ,
		_w9137_,
		_w9138_,
		_w18949_
	);
	LUT3 #(
		.INIT('h80)
	) name17049 (
		\m2_data_i[12]_pad ,
		_w9137_,
		_w9138_,
		_w18950_
	);
	LUT4 #(
		.INIT('hcdef)
	) name17050 (
		_w9132_,
		_w9135_,
		_w18949_,
		_w18950_,
		_w18951_
	);
	LUT3 #(
		.INIT('h2a)
	) name17051 (
		\m5_data_i[12]_pad ,
		_w9137_,
		_w9138_,
		_w18952_
	);
	LUT3 #(
		.INIT('h2a)
	) name17052 (
		\m1_data_i[12]_pad ,
		_w9137_,
		_w9138_,
		_w18953_
	);
	LUT4 #(
		.INIT('h37bf)
	) name17053 (
		_w9132_,
		_w9135_,
		_w18952_,
		_w18953_,
		_w18954_
	);
	LUT3 #(
		.INIT('h80)
	) name17054 (
		\m0_data_i[12]_pad ,
		_w9137_,
		_w9138_,
		_w18955_
	);
	LUT3 #(
		.INIT('h2a)
	) name17055 (
		\m7_data_i[12]_pad ,
		_w9137_,
		_w9138_,
		_w18956_
	);
	LUT4 #(
		.INIT('h6e7f)
	) name17056 (
		_w9132_,
		_w9135_,
		_w18955_,
		_w18956_,
		_w18957_
	);
	LUT4 #(
		.INIT('h7fff)
	) name17057 (
		_w18948_,
		_w18951_,
		_w18954_,
		_w18957_,
		_w18958_
	);
	LUT3 #(
		.INIT('h2a)
	) name17058 (
		\m3_data_i[13]_pad ,
		_w9137_,
		_w9138_,
		_w18959_
	);
	LUT3 #(
		.INIT('h80)
	) name17059 (
		\m4_data_i[13]_pad ,
		_w9137_,
		_w9138_,
		_w18960_
	);
	LUT4 #(
		.INIT('h9bdf)
	) name17060 (
		_w9132_,
		_w9135_,
		_w18959_,
		_w18960_,
		_w18961_
	);
	LUT3 #(
		.INIT('h80)
	) name17061 (
		\m6_data_i[13]_pad ,
		_w9137_,
		_w9138_,
		_w18962_
	);
	LUT3 #(
		.INIT('h80)
	) name17062 (
		\m2_data_i[13]_pad ,
		_w9137_,
		_w9138_,
		_w18963_
	);
	LUT4 #(
		.INIT('hcdef)
	) name17063 (
		_w9132_,
		_w9135_,
		_w18962_,
		_w18963_,
		_w18964_
	);
	LUT3 #(
		.INIT('h2a)
	) name17064 (
		\m5_data_i[13]_pad ,
		_w9137_,
		_w9138_,
		_w18965_
	);
	LUT3 #(
		.INIT('h2a)
	) name17065 (
		\m1_data_i[13]_pad ,
		_w9137_,
		_w9138_,
		_w18966_
	);
	LUT4 #(
		.INIT('h37bf)
	) name17066 (
		_w9132_,
		_w9135_,
		_w18965_,
		_w18966_,
		_w18967_
	);
	LUT3 #(
		.INIT('h80)
	) name17067 (
		\m0_data_i[13]_pad ,
		_w9137_,
		_w9138_,
		_w18968_
	);
	LUT3 #(
		.INIT('h2a)
	) name17068 (
		\m7_data_i[13]_pad ,
		_w9137_,
		_w9138_,
		_w18969_
	);
	LUT4 #(
		.INIT('h6e7f)
	) name17069 (
		_w9132_,
		_w9135_,
		_w18968_,
		_w18969_,
		_w18970_
	);
	LUT4 #(
		.INIT('h7fff)
	) name17070 (
		_w18961_,
		_w18964_,
		_w18967_,
		_w18970_,
		_w18971_
	);
	LUT3 #(
		.INIT('h2a)
	) name17071 (
		\m3_data_i[14]_pad ,
		_w9137_,
		_w9138_,
		_w18972_
	);
	LUT3 #(
		.INIT('h80)
	) name17072 (
		\m4_data_i[14]_pad ,
		_w9137_,
		_w9138_,
		_w18973_
	);
	LUT4 #(
		.INIT('h9bdf)
	) name17073 (
		_w9132_,
		_w9135_,
		_w18972_,
		_w18973_,
		_w18974_
	);
	LUT3 #(
		.INIT('h80)
	) name17074 (
		\m6_data_i[14]_pad ,
		_w9137_,
		_w9138_,
		_w18975_
	);
	LUT3 #(
		.INIT('h80)
	) name17075 (
		\m2_data_i[14]_pad ,
		_w9137_,
		_w9138_,
		_w18976_
	);
	LUT4 #(
		.INIT('hcdef)
	) name17076 (
		_w9132_,
		_w9135_,
		_w18975_,
		_w18976_,
		_w18977_
	);
	LUT3 #(
		.INIT('h2a)
	) name17077 (
		\m5_data_i[14]_pad ,
		_w9137_,
		_w9138_,
		_w18978_
	);
	LUT3 #(
		.INIT('h2a)
	) name17078 (
		\m1_data_i[14]_pad ,
		_w9137_,
		_w9138_,
		_w18979_
	);
	LUT4 #(
		.INIT('h37bf)
	) name17079 (
		_w9132_,
		_w9135_,
		_w18978_,
		_w18979_,
		_w18980_
	);
	LUT3 #(
		.INIT('h80)
	) name17080 (
		\m0_data_i[14]_pad ,
		_w9137_,
		_w9138_,
		_w18981_
	);
	LUT3 #(
		.INIT('h2a)
	) name17081 (
		\m7_data_i[14]_pad ,
		_w9137_,
		_w9138_,
		_w18982_
	);
	LUT4 #(
		.INIT('h6e7f)
	) name17082 (
		_w9132_,
		_w9135_,
		_w18981_,
		_w18982_,
		_w18983_
	);
	LUT4 #(
		.INIT('h7fff)
	) name17083 (
		_w18974_,
		_w18977_,
		_w18980_,
		_w18983_,
		_w18984_
	);
	LUT3 #(
		.INIT('h2a)
	) name17084 (
		\m3_data_i[15]_pad ,
		_w9137_,
		_w9138_,
		_w18985_
	);
	LUT3 #(
		.INIT('h80)
	) name17085 (
		\m4_data_i[15]_pad ,
		_w9137_,
		_w9138_,
		_w18986_
	);
	LUT4 #(
		.INIT('h9bdf)
	) name17086 (
		_w9132_,
		_w9135_,
		_w18985_,
		_w18986_,
		_w18987_
	);
	LUT3 #(
		.INIT('h80)
	) name17087 (
		\m6_data_i[15]_pad ,
		_w9137_,
		_w9138_,
		_w18988_
	);
	LUT3 #(
		.INIT('h80)
	) name17088 (
		\m2_data_i[15]_pad ,
		_w9137_,
		_w9138_,
		_w18989_
	);
	LUT4 #(
		.INIT('hcdef)
	) name17089 (
		_w9132_,
		_w9135_,
		_w18988_,
		_w18989_,
		_w18990_
	);
	LUT3 #(
		.INIT('h2a)
	) name17090 (
		\m5_data_i[15]_pad ,
		_w9137_,
		_w9138_,
		_w18991_
	);
	LUT3 #(
		.INIT('h2a)
	) name17091 (
		\m1_data_i[15]_pad ,
		_w9137_,
		_w9138_,
		_w18992_
	);
	LUT4 #(
		.INIT('h37bf)
	) name17092 (
		_w9132_,
		_w9135_,
		_w18991_,
		_w18992_,
		_w18993_
	);
	LUT3 #(
		.INIT('h80)
	) name17093 (
		\m0_data_i[15]_pad ,
		_w9137_,
		_w9138_,
		_w18994_
	);
	LUT3 #(
		.INIT('h2a)
	) name17094 (
		\m7_data_i[15]_pad ,
		_w9137_,
		_w9138_,
		_w18995_
	);
	LUT4 #(
		.INIT('h6e7f)
	) name17095 (
		_w9132_,
		_w9135_,
		_w18994_,
		_w18995_,
		_w18996_
	);
	LUT4 #(
		.INIT('h7fff)
	) name17096 (
		_w18987_,
		_w18990_,
		_w18993_,
		_w18996_,
		_w18997_
	);
	LUT3 #(
		.INIT('h2a)
	) name17097 (
		\m3_data_i[16]_pad ,
		_w9137_,
		_w9138_,
		_w18998_
	);
	LUT3 #(
		.INIT('h80)
	) name17098 (
		\m4_data_i[16]_pad ,
		_w9137_,
		_w9138_,
		_w18999_
	);
	LUT4 #(
		.INIT('h9bdf)
	) name17099 (
		_w9132_,
		_w9135_,
		_w18998_,
		_w18999_,
		_w19000_
	);
	LUT3 #(
		.INIT('h80)
	) name17100 (
		\m6_data_i[16]_pad ,
		_w9137_,
		_w9138_,
		_w19001_
	);
	LUT3 #(
		.INIT('h80)
	) name17101 (
		\m2_data_i[16]_pad ,
		_w9137_,
		_w9138_,
		_w19002_
	);
	LUT4 #(
		.INIT('hcdef)
	) name17102 (
		_w9132_,
		_w9135_,
		_w19001_,
		_w19002_,
		_w19003_
	);
	LUT3 #(
		.INIT('h2a)
	) name17103 (
		\m5_data_i[16]_pad ,
		_w9137_,
		_w9138_,
		_w19004_
	);
	LUT3 #(
		.INIT('h2a)
	) name17104 (
		\m1_data_i[16]_pad ,
		_w9137_,
		_w9138_,
		_w19005_
	);
	LUT4 #(
		.INIT('h37bf)
	) name17105 (
		_w9132_,
		_w9135_,
		_w19004_,
		_w19005_,
		_w19006_
	);
	LUT3 #(
		.INIT('h80)
	) name17106 (
		\m0_data_i[16]_pad ,
		_w9137_,
		_w9138_,
		_w19007_
	);
	LUT3 #(
		.INIT('h2a)
	) name17107 (
		\m7_data_i[16]_pad ,
		_w9137_,
		_w9138_,
		_w19008_
	);
	LUT4 #(
		.INIT('h6e7f)
	) name17108 (
		_w9132_,
		_w9135_,
		_w19007_,
		_w19008_,
		_w19009_
	);
	LUT4 #(
		.INIT('h7fff)
	) name17109 (
		_w19000_,
		_w19003_,
		_w19006_,
		_w19009_,
		_w19010_
	);
	LUT3 #(
		.INIT('h2a)
	) name17110 (
		\m3_data_i[17]_pad ,
		_w9137_,
		_w9138_,
		_w19011_
	);
	LUT3 #(
		.INIT('h80)
	) name17111 (
		\m4_data_i[17]_pad ,
		_w9137_,
		_w9138_,
		_w19012_
	);
	LUT4 #(
		.INIT('h9bdf)
	) name17112 (
		_w9132_,
		_w9135_,
		_w19011_,
		_w19012_,
		_w19013_
	);
	LUT3 #(
		.INIT('h80)
	) name17113 (
		\m6_data_i[17]_pad ,
		_w9137_,
		_w9138_,
		_w19014_
	);
	LUT3 #(
		.INIT('h80)
	) name17114 (
		\m2_data_i[17]_pad ,
		_w9137_,
		_w9138_,
		_w19015_
	);
	LUT4 #(
		.INIT('hcdef)
	) name17115 (
		_w9132_,
		_w9135_,
		_w19014_,
		_w19015_,
		_w19016_
	);
	LUT3 #(
		.INIT('h2a)
	) name17116 (
		\m5_data_i[17]_pad ,
		_w9137_,
		_w9138_,
		_w19017_
	);
	LUT3 #(
		.INIT('h2a)
	) name17117 (
		\m1_data_i[17]_pad ,
		_w9137_,
		_w9138_,
		_w19018_
	);
	LUT4 #(
		.INIT('h37bf)
	) name17118 (
		_w9132_,
		_w9135_,
		_w19017_,
		_w19018_,
		_w19019_
	);
	LUT3 #(
		.INIT('h80)
	) name17119 (
		\m0_data_i[17]_pad ,
		_w9137_,
		_w9138_,
		_w19020_
	);
	LUT3 #(
		.INIT('h2a)
	) name17120 (
		\m7_data_i[17]_pad ,
		_w9137_,
		_w9138_,
		_w19021_
	);
	LUT4 #(
		.INIT('h6e7f)
	) name17121 (
		_w9132_,
		_w9135_,
		_w19020_,
		_w19021_,
		_w19022_
	);
	LUT4 #(
		.INIT('h7fff)
	) name17122 (
		_w19013_,
		_w19016_,
		_w19019_,
		_w19022_,
		_w19023_
	);
	LUT3 #(
		.INIT('h2a)
	) name17123 (
		\m3_data_i[18]_pad ,
		_w9137_,
		_w9138_,
		_w19024_
	);
	LUT3 #(
		.INIT('h80)
	) name17124 (
		\m4_data_i[18]_pad ,
		_w9137_,
		_w9138_,
		_w19025_
	);
	LUT4 #(
		.INIT('h9bdf)
	) name17125 (
		_w9132_,
		_w9135_,
		_w19024_,
		_w19025_,
		_w19026_
	);
	LUT3 #(
		.INIT('h80)
	) name17126 (
		\m6_data_i[18]_pad ,
		_w9137_,
		_w9138_,
		_w19027_
	);
	LUT3 #(
		.INIT('h80)
	) name17127 (
		\m2_data_i[18]_pad ,
		_w9137_,
		_w9138_,
		_w19028_
	);
	LUT4 #(
		.INIT('hcdef)
	) name17128 (
		_w9132_,
		_w9135_,
		_w19027_,
		_w19028_,
		_w19029_
	);
	LUT3 #(
		.INIT('h2a)
	) name17129 (
		\m5_data_i[18]_pad ,
		_w9137_,
		_w9138_,
		_w19030_
	);
	LUT3 #(
		.INIT('h2a)
	) name17130 (
		\m1_data_i[18]_pad ,
		_w9137_,
		_w9138_,
		_w19031_
	);
	LUT4 #(
		.INIT('h37bf)
	) name17131 (
		_w9132_,
		_w9135_,
		_w19030_,
		_w19031_,
		_w19032_
	);
	LUT3 #(
		.INIT('h80)
	) name17132 (
		\m0_data_i[18]_pad ,
		_w9137_,
		_w9138_,
		_w19033_
	);
	LUT3 #(
		.INIT('h2a)
	) name17133 (
		\m7_data_i[18]_pad ,
		_w9137_,
		_w9138_,
		_w19034_
	);
	LUT4 #(
		.INIT('h6e7f)
	) name17134 (
		_w9132_,
		_w9135_,
		_w19033_,
		_w19034_,
		_w19035_
	);
	LUT4 #(
		.INIT('h7fff)
	) name17135 (
		_w19026_,
		_w19029_,
		_w19032_,
		_w19035_,
		_w19036_
	);
	LUT3 #(
		.INIT('h80)
	) name17136 (
		\m6_data_i[19]_pad ,
		_w9137_,
		_w9138_,
		_w19037_
	);
	LUT3 #(
		.INIT('h2a)
	) name17137 (
		\m5_data_i[19]_pad ,
		_w9137_,
		_w9138_,
		_w19038_
	);
	LUT4 #(
		.INIT('habef)
	) name17138 (
		_w9132_,
		_w9135_,
		_w19037_,
		_w19038_,
		_w19039_
	);
	LUT3 #(
		.INIT('h80)
	) name17139 (
		\m0_data_i[19]_pad ,
		_w9137_,
		_w9138_,
		_w19040_
	);
	LUT3 #(
		.INIT('h80)
	) name17140 (
		\m4_data_i[19]_pad ,
		_w9137_,
		_w9138_,
		_w19041_
	);
	LUT4 #(
		.INIT('h3b7f)
	) name17141 (
		_w9132_,
		_w9135_,
		_w19040_,
		_w19041_,
		_w19042_
	);
	LUT3 #(
		.INIT('h2a)
	) name17142 (
		\m7_data_i[19]_pad ,
		_w9137_,
		_w9138_,
		_w19043_
	);
	LUT3 #(
		.INIT('h2a)
	) name17143 (
		\m3_data_i[19]_pad ,
		_w9137_,
		_w9138_,
		_w19044_
	);
	LUT4 #(
		.INIT('hcdef)
	) name17144 (
		_w9132_,
		_w9135_,
		_w19043_,
		_w19044_,
		_w19045_
	);
	LUT3 #(
		.INIT('h2a)
	) name17145 (
		\m1_data_i[19]_pad ,
		_w9137_,
		_w9138_,
		_w19046_
	);
	LUT3 #(
		.INIT('h80)
	) name17146 (
		\m2_data_i[19]_pad ,
		_w9137_,
		_w9138_,
		_w19047_
	);
	LUT4 #(
		.INIT('h5d7f)
	) name17147 (
		_w9132_,
		_w9135_,
		_w19046_,
		_w19047_,
		_w19048_
	);
	LUT4 #(
		.INIT('h7fff)
	) name17148 (
		_w19039_,
		_w19042_,
		_w19045_,
		_w19048_,
		_w19049_
	);
	LUT3 #(
		.INIT('h2a)
	) name17149 (
		\m3_data_i[1]_pad ,
		_w9137_,
		_w9138_,
		_w19050_
	);
	LUT3 #(
		.INIT('h80)
	) name17150 (
		\m4_data_i[1]_pad ,
		_w9137_,
		_w9138_,
		_w19051_
	);
	LUT4 #(
		.INIT('h9bdf)
	) name17151 (
		_w9132_,
		_w9135_,
		_w19050_,
		_w19051_,
		_w19052_
	);
	LUT3 #(
		.INIT('h80)
	) name17152 (
		\m6_data_i[1]_pad ,
		_w9137_,
		_w9138_,
		_w19053_
	);
	LUT3 #(
		.INIT('h80)
	) name17153 (
		\m2_data_i[1]_pad ,
		_w9137_,
		_w9138_,
		_w19054_
	);
	LUT4 #(
		.INIT('hcdef)
	) name17154 (
		_w9132_,
		_w9135_,
		_w19053_,
		_w19054_,
		_w19055_
	);
	LUT3 #(
		.INIT('h2a)
	) name17155 (
		\m5_data_i[1]_pad ,
		_w9137_,
		_w9138_,
		_w19056_
	);
	LUT3 #(
		.INIT('h2a)
	) name17156 (
		\m1_data_i[1]_pad ,
		_w9137_,
		_w9138_,
		_w19057_
	);
	LUT4 #(
		.INIT('h37bf)
	) name17157 (
		_w9132_,
		_w9135_,
		_w19056_,
		_w19057_,
		_w19058_
	);
	LUT3 #(
		.INIT('h80)
	) name17158 (
		\m0_data_i[1]_pad ,
		_w9137_,
		_w9138_,
		_w19059_
	);
	LUT3 #(
		.INIT('h2a)
	) name17159 (
		\m7_data_i[1]_pad ,
		_w9137_,
		_w9138_,
		_w19060_
	);
	LUT4 #(
		.INIT('h6e7f)
	) name17160 (
		_w9132_,
		_w9135_,
		_w19059_,
		_w19060_,
		_w19061_
	);
	LUT4 #(
		.INIT('h7fff)
	) name17161 (
		_w19052_,
		_w19055_,
		_w19058_,
		_w19061_,
		_w19062_
	);
	LUT3 #(
		.INIT('h2a)
	) name17162 (
		\m3_data_i[20]_pad ,
		_w9137_,
		_w9138_,
		_w19063_
	);
	LUT3 #(
		.INIT('h80)
	) name17163 (
		\m4_data_i[20]_pad ,
		_w9137_,
		_w9138_,
		_w19064_
	);
	LUT4 #(
		.INIT('h9bdf)
	) name17164 (
		_w9132_,
		_w9135_,
		_w19063_,
		_w19064_,
		_w19065_
	);
	LUT3 #(
		.INIT('h80)
	) name17165 (
		\m6_data_i[20]_pad ,
		_w9137_,
		_w9138_,
		_w19066_
	);
	LUT3 #(
		.INIT('h80)
	) name17166 (
		\m2_data_i[20]_pad ,
		_w9137_,
		_w9138_,
		_w19067_
	);
	LUT4 #(
		.INIT('hcdef)
	) name17167 (
		_w9132_,
		_w9135_,
		_w19066_,
		_w19067_,
		_w19068_
	);
	LUT3 #(
		.INIT('h2a)
	) name17168 (
		\m5_data_i[20]_pad ,
		_w9137_,
		_w9138_,
		_w19069_
	);
	LUT3 #(
		.INIT('h2a)
	) name17169 (
		\m1_data_i[20]_pad ,
		_w9137_,
		_w9138_,
		_w19070_
	);
	LUT4 #(
		.INIT('h37bf)
	) name17170 (
		_w9132_,
		_w9135_,
		_w19069_,
		_w19070_,
		_w19071_
	);
	LUT3 #(
		.INIT('h80)
	) name17171 (
		\m0_data_i[20]_pad ,
		_w9137_,
		_w9138_,
		_w19072_
	);
	LUT3 #(
		.INIT('h2a)
	) name17172 (
		\m7_data_i[20]_pad ,
		_w9137_,
		_w9138_,
		_w19073_
	);
	LUT4 #(
		.INIT('h6e7f)
	) name17173 (
		_w9132_,
		_w9135_,
		_w19072_,
		_w19073_,
		_w19074_
	);
	LUT4 #(
		.INIT('h7fff)
	) name17174 (
		_w19065_,
		_w19068_,
		_w19071_,
		_w19074_,
		_w19075_
	);
	LUT3 #(
		.INIT('h2a)
	) name17175 (
		\m1_data_i[21]_pad ,
		_w9137_,
		_w9138_,
		_w19076_
	);
	LUT3 #(
		.INIT('h80)
	) name17176 (
		\m2_data_i[21]_pad ,
		_w9137_,
		_w9138_,
		_w19077_
	);
	LUT4 #(
		.INIT('h5d7f)
	) name17177 (
		_w9132_,
		_w9135_,
		_w19076_,
		_w19077_,
		_w19078_
	);
	LUT3 #(
		.INIT('h80)
	) name17178 (
		\m6_data_i[21]_pad ,
		_w9137_,
		_w9138_,
		_w19079_
	);
	LUT3 #(
		.INIT('h2a)
	) name17179 (
		\m7_data_i[21]_pad ,
		_w9137_,
		_w9138_,
		_w19080_
	);
	LUT3 #(
		.INIT('h57)
	) name17180 (
		_w9150_,
		_w19079_,
		_w19080_,
		_w19081_
	);
	LUT3 #(
		.INIT('h2a)
	) name17181 (
		\m5_data_i[21]_pad ,
		_w9137_,
		_w9138_,
		_w19082_
	);
	LUT3 #(
		.INIT('h80)
	) name17182 (
		\m0_data_i[21]_pad ,
		_w9137_,
		_w9138_,
		_w19083_
	);
	LUT4 #(
		.INIT('h37bf)
	) name17183 (
		_w9132_,
		_w9135_,
		_w19082_,
		_w19083_,
		_w19084_
	);
	LUT3 #(
		.INIT('h2a)
	) name17184 (
		\m3_data_i[21]_pad ,
		_w9137_,
		_w9138_,
		_w19085_
	);
	LUT3 #(
		.INIT('h80)
	) name17185 (
		\m4_data_i[21]_pad ,
		_w9137_,
		_w9138_,
		_w19086_
	);
	LUT4 #(
		.INIT('h9bdf)
	) name17186 (
		_w9132_,
		_w9135_,
		_w19085_,
		_w19086_,
		_w19087_
	);
	LUT4 #(
		.INIT('h7fff)
	) name17187 (
		_w19078_,
		_w19081_,
		_w19084_,
		_w19087_,
		_w19088_
	);
	LUT3 #(
		.INIT('h2a)
	) name17188 (
		\m3_data_i[22]_pad ,
		_w9137_,
		_w9138_,
		_w19089_
	);
	LUT3 #(
		.INIT('h80)
	) name17189 (
		\m4_data_i[22]_pad ,
		_w9137_,
		_w9138_,
		_w19090_
	);
	LUT4 #(
		.INIT('h9bdf)
	) name17190 (
		_w9132_,
		_w9135_,
		_w19089_,
		_w19090_,
		_w19091_
	);
	LUT3 #(
		.INIT('h80)
	) name17191 (
		\m6_data_i[22]_pad ,
		_w9137_,
		_w9138_,
		_w19092_
	);
	LUT3 #(
		.INIT('h80)
	) name17192 (
		\m2_data_i[22]_pad ,
		_w9137_,
		_w9138_,
		_w19093_
	);
	LUT4 #(
		.INIT('hcdef)
	) name17193 (
		_w9132_,
		_w9135_,
		_w19092_,
		_w19093_,
		_w19094_
	);
	LUT3 #(
		.INIT('h2a)
	) name17194 (
		\m5_data_i[22]_pad ,
		_w9137_,
		_w9138_,
		_w19095_
	);
	LUT3 #(
		.INIT('h2a)
	) name17195 (
		\m1_data_i[22]_pad ,
		_w9137_,
		_w9138_,
		_w19096_
	);
	LUT4 #(
		.INIT('h37bf)
	) name17196 (
		_w9132_,
		_w9135_,
		_w19095_,
		_w19096_,
		_w19097_
	);
	LUT3 #(
		.INIT('h80)
	) name17197 (
		\m0_data_i[22]_pad ,
		_w9137_,
		_w9138_,
		_w19098_
	);
	LUT3 #(
		.INIT('h2a)
	) name17198 (
		\m7_data_i[22]_pad ,
		_w9137_,
		_w9138_,
		_w19099_
	);
	LUT4 #(
		.INIT('h6e7f)
	) name17199 (
		_w9132_,
		_w9135_,
		_w19098_,
		_w19099_,
		_w19100_
	);
	LUT4 #(
		.INIT('h7fff)
	) name17200 (
		_w19091_,
		_w19094_,
		_w19097_,
		_w19100_,
		_w19101_
	);
	LUT3 #(
		.INIT('h2a)
	) name17201 (
		\m3_data_i[23]_pad ,
		_w9137_,
		_w9138_,
		_w19102_
	);
	LUT3 #(
		.INIT('h80)
	) name17202 (
		\m4_data_i[23]_pad ,
		_w9137_,
		_w9138_,
		_w19103_
	);
	LUT4 #(
		.INIT('h9bdf)
	) name17203 (
		_w9132_,
		_w9135_,
		_w19102_,
		_w19103_,
		_w19104_
	);
	LUT3 #(
		.INIT('h80)
	) name17204 (
		\m6_data_i[23]_pad ,
		_w9137_,
		_w9138_,
		_w19105_
	);
	LUT3 #(
		.INIT('h80)
	) name17205 (
		\m2_data_i[23]_pad ,
		_w9137_,
		_w9138_,
		_w19106_
	);
	LUT4 #(
		.INIT('hcdef)
	) name17206 (
		_w9132_,
		_w9135_,
		_w19105_,
		_w19106_,
		_w19107_
	);
	LUT3 #(
		.INIT('h2a)
	) name17207 (
		\m5_data_i[23]_pad ,
		_w9137_,
		_w9138_,
		_w19108_
	);
	LUT3 #(
		.INIT('h2a)
	) name17208 (
		\m1_data_i[23]_pad ,
		_w9137_,
		_w9138_,
		_w19109_
	);
	LUT4 #(
		.INIT('h37bf)
	) name17209 (
		_w9132_,
		_w9135_,
		_w19108_,
		_w19109_,
		_w19110_
	);
	LUT3 #(
		.INIT('h80)
	) name17210 (
		\m0_data_i[23]_pad ,
		_w9137_,
		_w9138_,
		_w19111_
	);
	LUT3 #(
		.INIT('h2a)
	) name17211 (
		\m7_data_i[23]_pad ,
		_w9137_,
		_w9138_,
		_w19112_
	);
	LUT4 #(
		.INIT('h6e7f)
	) name17212 (
		_w9132_,
		_w9135_,
		_w19111_,
		_w19112_,
		_w19113_
	);
	LUT4 #(
		.INIT('h7fff)
	) name17213 (
		_w19104_,
		_w19107_,
		_w19110_,
		_w19113_,
		_w19114_
	);
	LUT3 #(
		.INIT('h2a)
	) name17214 (
		\m3_data_i[24]_pad ,
		_w9137_,
		_w9138_,
		_w19115_
	);
	LUT3 #(
		.INIT('h80)
	) name17215 (
		\m4_data_i[24]_pad ,
		_w9137_,
		_w9138_,
		_w19116_
	);
	LUT4 #(
		.INIT('h9bdf)
	) name17216 (
		_w9132_,
		_w9135_,
		_w19115_,
		_w19116_,
		_w19117_
	);
	LUT3 #(
		.INIT('h80)
	) name17217 (
		\m6_data_i[24]_pad ,
		_w9137_,
		_w9138_,
		_w19118_
	);
	LUT3 #(
		.INIT('h80)
	) name17218 (
		\m2_data_i[24]_pad ,
		_w9137_,
		_w9138_,
		_w19119_
	);
	LUT4 #(
		.INIT('hcdef)
	) name17219 (
		_w9132_,
		_w9135_,
		_w19118_,
		_w19119_,
		_w19120_
	);
	LUT3 #(
		.INIT('h2a)
	) name17220 (
		\m5_data_i[24]_pad ,
		_w9137_,
		_w9138_,
		_w19121_
	);
	LUT3 #(
		.INIT('h2a)
	) name17221 (
		\m1_data_i[24]_pad ,
		_w9137_,
		_w9138_,
		_w19122_
	);
	LUT4 #(
		.INIT('h37bf)
	) name17222 (
		_w9132_,
		_w9135_,
		_w19121_,
		_w19122_,
		_w19123_
	);
	LUT3 #(
		.INIT('h80)
	) name17223 (
		\m0_data_i[24]_pad ,
		_w9137_,
		_w9138_,
		_w19124_
	);
	LUT3 #(
		.INIT('h2a)
	) name17224 (
		\m7_data_i[24]_pad ,
		_w9137_,
		_w9138_,
		_w19125_
	);
	LUT4 #(
		.INIT('h6e7f)
	) name17225 (
		_w9132_,
		_w9135_,
		_w19124_,
		_w19125_,
		_w19126_
	);
	LUT4 #(
		.INIT('h7fff)
	) name17226 (
		_w19117_,
		_w19120_,
		_w19123_,
		_w19126_,
		_w19127_
	);
	LUT3 #(
		.INIT('h2a)
	) name17227 (
		\m3_data_i[25]_pad ,
		_w9137_,
		_w9138_,
		_w19128_
	);
	LUT3 #(
		.INIT('h80)
	) name17228 (
		\m4_data_i[25]_pad ,
		_w9137_,
		_w9138_,
		_w19129_
	);
	LUT4 #(
		.INIT('h9bdf)
	) name17229 (
		_w9132_,
		_w9135_,
		_w19128_,
		_w19129_,
		_w19130_
	);
	LUT3 #(
		.INIT('h80)
	) name17230 (
		\m6_data_i[25]_pad ,
		_w9137_,
		_w9138_,
		_w19131_
	);
	LUT3 #(
		.INIT('h80)
	) name17231 (
		\m2_data_i[25]_pad ,
		_w9137_,
		_w9138_,
		_w19132_
	);
	LUT4 #(
		.INIT('hcdef)
	) name17232 (
		_w9132_,
		_w9135_,
		_w19131_,
		_w19132_,
		_w19133_
	);
	LUT3 #(
		.INIT('h2a)
	) name17233 (
		\m5_data_i[25]_pad ,
		_w9137_,
		_w9138_,
		_w19134_
	);
	LUT3 #(
		.INIT('h2a)
	) name17234 (
		\m1_data_i[25]_pad ,
		_w9137_,
		_w9138_,
		_w19135_
	);
	LUT4 #(
		.INIT('h37bf)
	) name17235 (
		_w9132_,
		_w9135_,
		_w19134_,
		_w19135_,
		_w19136_
	);
	LUT3 #(
		.INIT('h80)
	) name17236 (
		\m0_data_i[25]_pad ,
		_w9137_,
		_w9138_,
		_w19137_
	);
	LUT3 #(
		.INIT('h2a)
	) name17237 (
		\m7_data_i[25]_pad ,
		_w9137_,
		_w9138_,
		_w19138_
	);
	LUT4 #(
		.INIT('h6e7f)
	) name17238 (
		_w9132_,
		_w9135_,
		_w19137_,
		_w19138_,
		_w19139_
	);
	LUT4 #(
		.INIT('h7fff)
	) name17239 (
		_w19130_,
		_w19133_,
		_w19136_,
		_w19139_,
		_w19140_
	);
	LUT3 #(
		.INIT('h2a)
	) name17240 (
		\m3_data_i[26]_pad ,
		_w9137_,
		_w9138_,
		_w19141_
	);
	LUT3 #(
		.INIT('h80)
	) name17241 (
		\m4_data_i[26]_pad ,
		_w9137_,
		_w9138_,
		_w19142_
	);
	LUT4 #(
		.INIT('h9bdf)
	) name17242 (
		_w9132_,
		_w9135_,
		_w19141_,
		_w19142_,
		_w19143_
	);
	LUT3 #(
		.INIT('h80)
	) name17243 (
		\m6_data_i[26]_pad ,
		_w9137_,
		_w9138_,
		_w19144_
	);
	LUT3 #(
		.INIT('h80)
	) name17244 (
		\m2_data_i[26]_pad ,
		_w9137_,
		_w9138_,
		_w19145_
	);
	LUT4 #(
		.INIT('hcdef)
	) name17245 (
		_w9132_,
		_w9135_,
		_w19144_,
		_w19145_,
		_w19146_
	);
	LUT3 #(
		.INIT('h2a)
	) name17246 (
		\m5_data_i[26]_pad ,
		_w9137_,
		_w9138_,
		_w19147_
	);
	LUT3 #(
		.INIT('h2a)
	) name17247 (
		\m1_data_i[26]_pad ,
		_w9137_,
		_w9138_,
		_w19148_
	);
	LUT4 #(
		.INIT('h37bf)
	) name17248 (
		_w9132_,
		_w9135_,
		_w19147_,
		_w19148_,
		_w19149_
	);
	LUT3 #(
		.INIT('h80)
	) name17249 (
		\m0_data_i[26]_pad ,
		_w9137_,
		_w9138_,
		_w19150_
	);
	LUT3 #(
		.INIT('h2a)
	) name17250 (
		\m7_data_i[26]_pad ,
		_w9137_,
		_w9138_,
		_w19151_
	);
	LUT4 #(
		.INIT('h6e7f)
	) name17251 (
		_w9132_,
		_w9135_,
		_w19150_,
		_w19151_,
		_w19152_
	);
	LUT4 #(
		.INIT('h7fff)
	) name17252 (
		_w19143_,
		_w19146_,
		_w19149_,
		_w19152_,
		_w19153_
	);
	LUT3 #(
		.INIT('h2a)
	) name17253 (
		\m3_data_i[27]_pad ,
		_w9137_,
		_w9138_,
		_w19154_
	);
	LUT3 #(
		.INIT('h80)
	) name17254 (
		\m4_data_i[27]_pad ,
		_w9137_,
		_w9138_,
		_w19155_
	);
	LUT4 #(
		.INIT('h9bdf)
	) name17255 (
		_w9132_,
		_w9135_,
		_w19154_,
		_w19155_,
		_w19156_
	);
	LUT3 #(
		.INIT('h80)
	) name17256 (
		\m6_data_i[27]_pad ,
		_w9137_,
		_w9138_,
		_w19157_
	);
	LUT3 #(
		.INIT('h80)
	) name17257 (
		\m2_data_i[27]_pad ,
		_w9137_,
		_w9138_,
		_w19158_
	);
	LUT4 #(
		.INIT('hcdef)
	) name17258 (
		_w9132_,
		_w9135_,
		_w19157_,
		_w19158_,
		_w19159_
	);
	LUT3 #(
		.INIT('h2a)
	) name17259 (
		\m5_data_i[27]_pad ,
		_w9137_,
		_w9138_,
		_w19160_
	);
	LUT3 #(
		.INIT('h2a)
	) name17260 (
		\m1_data_i[27]_pad ,
		_w9137_,
		_w9138_,
		_w19161_
	);
	LUT4 #(
		.INIT('h37bf)
	) name17261 (
		_w9132_,
		_w9135_,
		_w19160_,
		_w19161_,
		_w19162_
	);
	LUT3 #(
		.INIT('h80)
	) name17262 (
		\m0_data_i[27]_pad ,
		_w9137_,
		_w9138_,
		_w19163_
	);
	LUT3 #(
		.INIT('h2a)
	) name17263 (
		\m7_data_i[27]_pad ,
		_w9137_,
		_w9138_,
		_w19164_
	);
	LUT4 #(
		.INIT('h6e7f)
	) name17264 (
		_w9132_,
		_w9135_,
		_w19163_,
		_w19164_,
		_w19165_
	);
	LUT4 #(
		.INIT('h7fff)
	) name17265 (
		_w19156_,
		_w19159_,
		_w19162_,
		_w19165_,
		_w19166_
	);
	LUT3 #(
		.INIT('h2a)
	) name17266 (
		\m3_data_i[28]_pad ,
		_w9137_,
		_w9138_,
		_w19167_
	);
	LUT3 #(
		.INIT('h80)
	) name17267 (
		\m4_data_i[28]_pad ,
		_w9137_,
		_w9138_,
		_w19168_
	);
	LUT4 #(
		.INIT('h9bdf)
	) name17268 (
		_w9132_,
		_w9135_,
		_w19167_,
		_w19168_,
		_w19169_
	);
	LUT3 #(
		.INIT('h80)
	) name17269 (
		\m6_data_i[28]_pad ,
		_w9137_,
		_w9138_,
		_w19170_
	);
	LUT3 #(
		.INIT('h80)
	) name17270 (
		\m2_data_i[28]_pad ,
		_w9137_,
		_w9138_,
		_w19171_
	);
	LUT4 #(
		.INIT('hcdef)
	) name17271 (
		_w9132_,
		_w9135_,
		_w19170_,
		_w19171_,
		_w19172_
	);
	LUT3 #(
		.INIT('h2a)
	) name17272 (
		\m5_data_i[28]_pad ,
		_w9137_,
		_w9138_,
		_w19173_
	);
	LUT3 #(
		.INIT('h2a)
	) name17273 (
		\m1_data_i[28]_pad ,
		_w9137_,
		_w9138_,
		_w19174_
	);
	LUT4 #(
		.INIT('h37bf)
	) name17274 (
		_w9132_,
		_w9135_,
		_w19173_,
		_w19174_,
		_w19175_
	);
	LUT3 #(
		.INIT('h80)
	) name17275 (
		\m0_data_i[28]_pad ,
		_w9137_,
		_w9138_,
		_w19176_
	);
	LUT3 #(
		.INIT('h2a)
	) name17276 (
		\m7_data_i[28]_pad ,
		_w9137_,
		_w9138_,
		_w19177_
	);
	LUT4 #(
		.INIT('h6e7f)
	) name17277 (
		_w9132_,
		_w9135_,
		_w19176_,
		_w19177_,
		_w19178_
	);
	LUT4 #(
		.INIT('h7fff)
	) name17278 (
		_w19169_,
		_w19172_,
		_w19175_,
		_w19178_,
		_w19179_
	);
	LUT3 #(
		.INIT('h2a)
	) name17279 (
		\m3_data_i[29]_pad ,
		_w9137_,
		_w9138_,
		_w19180_
	);
	LUT3 #(
		.INIT('h80)
	) name17280 (
		\m4_data_i[29]_pad ,
		_w9137_,
		_w9138_,
		_w19181_
	);
	LUT4 #(
		.INIT('h9bdf)
	) name17281 (
		_w9132_,
		_w9135_,
		_w19180_,
		_w19181_,
		_w19182_
	);
	LUT3 #(
		.INIT('h80)
	) name17282 (
		\m0_data_i[29]_pad ,
		_w9137_,
		_w9138_,
		_w19183_
	);
	LUT3 #(
		.INIT('h2a)
	) name17283 (
		\m5_data_i[29]_pad ,
		_w9137_,
		_w9138_,
		_w19184_
	);
	LUT4 #(
		.INIT('h3b7f)
	) name17284 (
		_w9132_,
		_w9135_,
		_w19183_,
		_w19184_,
		_w19185_
	);
	LUT3 #(
		.INIT('h2a)
	) name17285 (
		\m7_data_i[29]_pad ,
		_w9137_,
		_w9138_,
		_w19186_
	);
	LUT3 #(
		.INIT('h80)
	) name17286 (
		\m6_data_i[29]_pad ,
		_w9137_,
		_w9138_,
		_w19187_
	);
	LUT3 #(
		.INIT('h57)
	) name17287 (
		_w9150_,
		_w19186_,
		_w19187_,
		_w19188_
	);
	LUT3 #(
		.INIT('h2a)
	) name17288 (
		\m1_data_i[29]_pad ,
		_w9137_,
		_w9138_,
		_w19189_
	);
	LUT3 #(
		.INIT('h80)
	) name17289 (
		\m2_data_i[29]_pad ,
		_w9137_,
		_w9138_,
		_w19190_
	);
	LUT4 #(
		.INIT('h5d7f)
	) name17290 (
		_w9132_,
		_w9135_,
		_w19189_,
		_w19190_,
		_w19191_
	);
	LUT4 #(
		.INIT('h7fff)
	) name17291 (
		_w19182_,
		_w19185_,
		_w19188_,
		_w19191_,
		_w19192_
	);
	LUT3 #(
		.INIT('h2a)
	) name17292 (
		\m3_data_i[2]_pad ,
		_w9137_,
		_w9138_,
		_w19193_
	);
	LUT3 #(
		.INIT('h80)
	) name17293 (
		\m4_data_i[2]_pad ,
		_w9137_,
		_w9138_,
		_w19194_
	);
	LUT4 #(
		.INIT('h9bdf)
	) name17294 (
		_w9132_,
		_w9135_,
		_w19193_,
		_w19194_,
		_w19195_
	);
	LUT3 #(
		.INIT('h80)
	) name17295 (
		\m6_data_i[2]_pad ,
		_w9137_,
		_w9138_,
		_w19196_
	);
	LUT3 #(
		.INIT('h80)
	) name17296 (
		\m2_data_i[2]_pad ,
		_w9137_,
		_w9138_,
		_w19197_
	);
	LUT4 #(
		.INIT('hcdef)
	) name17297 (
		_w9132_,
		_w9135_,
		_w19196_,
		_w19197_,
		_w19198_
	);
	LUT3 #(
		.INIT('h2a)
	) name17298 (
		\m5_data_i[2]_pad ,
		_w9137_,
		_w9138_,
		_w19199_
	);
	LUT3 #(
		.INIT('h2a)
	) name17299 (
		\m1_data_i[2]_pad ,
		_w9137_,
		_w9138_,
		_w19200_
	);
	LUT4 #(
		.INIT('h37bf)
	) name17300 (
		_w9132_,
		_w9135_,
		_w19199_,
		_w19200_,
		_w19201_
	);
	LUT3 #(
		.INIT('h80)
	) name17301 (
		\m0_data_i[2]_pad ,
		_w9137_,
		_w9138_,
		_w19202_
	);
	LUT3 #(
		.INIT('h2a)
	) name17302 (
		\m7_data_i[2]_pad ,
		_w9137_,
		_w9138_,
		_w19203_
	);
	LUT4 #(
		.INIT('h6e7f)
	) name17303 (
		_w9132_,
		_w9135_,
		_w19202_,
		_w19203_,
		_w19204_
	);
	LUT4 #(
		.INIT('h7fff)
	) name17304 (
		_w19195_,
		_w19198_,
		_w19201_,
		_w19204_,
		_w19205_
	);
	LUT3 #(
		.INIT('h2a)
	) name17305 (
		\m3_data_i[30]_pad ,
		_w9137_,
		_w9138_,
		_w19206_
	);
	LUT3 #(
		.INIT('h80)
	) name17306 (
		\m4_data_i[30]_pad ,
		_w9137_,
		_w9138_,
		_w19207_
	);
	LUT4 #(
		.INIT('h9bdf)
	) name17307 (
		_w9132_,
		_w9135_,
		_w19206_,
		_w19207_,
		_w19208_
	);
	LUT3 #(
		.INIT('h80)
	) name17308 (
		\m0_data_i[30]_pad ,
		_w9137_,
		_w9138_,
		_w19209_
	);
	LUT3 #(
		.INIT('h2a)
	) name17309 (
		\m5_data_i[30]_pad ,
		_w9137_,
		_w9138_,
		_w19210_
	);
	LUT4 #(
		.INIT('h3b7f)
	) name17310 (
		_w9132_,
		_w9135_,
		_w19209_,
		_w19210_,
		_w19211_
	);
	LUT3 #(
		.INIT('h2a)
	) name17311 (
		\m7_data_i[30]_pad ,
		_w9137_,
		_w9138_,
		_w19212_
	);
	LUT3 #(
		.INIT('h80)
	) name17312 (
		\m6_data_i[30]_pad ,
		_w9137_,
		_w9138_,
		_w19213_
	);
	LUT3 #(
		.INIT('h57)
	) name17313 (
		_w9150_,
		_w19212_,
		_w19213_,
		_w19214_
	);
	LUT3 #(
		.INIT('h2a)
	) name17314 (
		\m1_data_i[30]_pad ,
		_w9137_,
		_w9138_,
		_w19215_
	);
	LUT3 #(
		.INIT('h80)
	) name17315 (
		\m2_data_i[30]_pad ,
		_w9137_,
		_w9138_,
		_w19216_
	);
	LUT4 #(
		.INIT('h5d7f)
	) name17316 (
		_w9132_,
		_w9135_,
		_w19215_,
		_w19216_,
		_w19217_
	);
	LUT4 #(
		.INIT('h7fff)
	) name17317 (
		_w19208_,
		_w19211_,
		_w19214_,
		_w19217_,
		_w19218_
	);
	LUT3 #(
		.INIT('h2a)
	) name17318 (
		\m1_data_i[31]_pad ,
		_w9137_,
		_w9138_,
		_w19219_
	);
	LUT3 #(
		.INIT('h80)
	) name17319 (
		\m2_data_i[31]_pad ,
		_w9137_,
		_w9138_,
		_w19220_
	);
	LUT4 #(
		.INIT('h5d7f)
	) name17320 (
		_w9132_,
		_w9135_,
		_w19219_,
		_w19220_,
		_w19221_
	);
	LUT3 #(
		.INIT('h80)
	) name17321 (
		\m6_data_i[31]_pad ,
		_w9137_,
		_w9138_,
		_w19222_
	);
	LUT3 #(
		.INIT('h2a)
	) name17322 (
		\m7_data_i[31]_pad ,
		_w9137_,
		_w9138_,
		_w19223_
	);
	LUT3 #(
		.INIT('h57)
	) name17323 (
		_w9150_,
		_w19222_,
		_w19223_,
		_w19224_
	);
	LUT3 #(
		.INIT('h2a)
	) name17324 (
		\m5_data_i[31]_pad ,
		_w9137_,
		_w9138_,
		_w19225_
	);
	LUT3 #(
		.INIT('h80)
	) name17325 (
		\m0_data_i[31]_pad ,
		_w9137_,
		_w9138_,
		_w19226_
	);
	LUT4 #(
		.INIT('h37bf)
	) name17326 (
		_w9132_,
		_w9135_,
		_w19225_,
		_w19226_,
		_w19227_
	);
	LUT3 #(
		.INIT('h2a)
	) name17327 (
		\m3_data_i[31]_pad ,
		_w9137_,
		_w9138_,
		_w19228_
	);
	LUT3 #(
		.INIT('h80)
	) name17328 (
		\m4_data_i[31]_pad ,
		_w9137_,
		_w9138_,
		_w19229_
	);
	LUT4 #(
		.INIT('h9bdf)
	) name17329 (
		_w9132_,
		_w9135_,
		_w19228_,
		_w19229_,
		_w19230_
	);
	LUT4 #(
		.INIT('h7fff)
	) name17330 (
		_w19221_,
		_w19224_,
		_w19227_,
		_w19230_,
		_w19231_
	);
	LUT3 #(
		.INIT('h2a)
	) name17331 (
		\m3_data_i[3]_pad ,
		_w9137_,
		_w9138_,
		_w19232_
	);
	LUT3 #(
		.INIT('h80)
	) name17332 (
		\m4_data_i[3]_pad ,
		_w9137_,
		_w9138_,
		_w19233_
	);
	LUT4 #(
		.INIT('h9bdf)
	) name17333 (
		_w9132_,
		_w9135_,
		_w19232_,
		_w19233_,
		_w19234_
	);
	LUT3 #(
		.INIT('h80)
	) name17334 (
		\m6_data_i[3]_pad ,
		_w9137_,
		_w9138_,
		_w19235_
	);
	LUT3 #(
		.INIT('h80)
	) name17335 (
		\m2_data_i[3]_pad ,
		_w9137_,
		_w9138_,
		_w19236_
	);
	LUT4 #(
		.INIT('hcdef)
	) name17336 (
		_w9132_,
		_w9135_,
		_w19235_,
		_w19236_,
		_w19237_
	);
	LUT3 #(
		.INIT('h2a)
	) name17337 (
		\m5_data_i[3]_pad ,
		_w9137_,
		_w9138_,
		_w19238_
	);
	LUT3 #(
		.INIT('h2a)
	) name17338 (
		\m1_data_i[3]_pad ,
		_w9137_,
		_w9138_,
		_w19239_
	);
	LUT4 #(
		.INIT('h37bf)
	) name17339 (
		_w9132_,
		_w9135_,
		_w19238_,
		_w19239_,
		_w19240_
	);
	LUT3 #(
		.INIT('h80)
	) name17340 (
		\m0_data_i[3]_pad ,
		_w9137_,
		_w9138_,
		_w19241_
	);
	LUT3 #(
		.INIT('h2a)
	) name17341 (
		\m7_data_i[3]_pad ,
		_w9137_,
		_w9138_,
		_w19242_
	);
	LUT4 #(
		.INIT('h6e7f)
	) name17342 (
		_w9132_,
		_w9135_,
		_w19241_,
		_w19242_,
		_w19243_
	);
	LUT4 #(
		.INIT('h7fff)
	) name17343 (
		_w19234_,
		_w19237_,
		_w19240_,
		_w19243_,
		_w19244_
	);
	LUT3 #(
		.INIT('h80)
	) name17344 (
		\m6_data_i[4]_pad ,
		_w9137_,
		_w9138_,
		_w19245_
	);
	LUT3 #(
		.INIT('h2a)
	) name17345 (
		\m5_data_i[4]_pad ,
		_w9137_,
		_w9138_,
		_w19246_
	);
	LUT4 #(
		.INIT('habef)
	) name17346 (
		_w9132_,
		_w9135_,
		_w19245_,
		_w19246_,
		_w19247_
	);
	LUT3 #(
		.INIT('h2a)
	) name17347 (
		\m3_data_i[4]_pad ,
		_w9137_,
		_w9138_,
		_w19248_
	);
	LUT3 #(
		.INIT('h80)
	) name17348 (
		\m2_data_i[4]_pad ,
		_w9137_,
		_w9138_,
		_w19249_
	);
	LUT3 #(
		.INIT('h57)
	) name17349 (
		_w9144_,
		_w19248_,
		_w19249_,
		_w19250_
	);
	LUT3 #(
		.INIT('h80)
	) name17350 (
		\m4_data_i[4]_pad ,
		_w9137_,
		_w9138_,
		_w19251_
	);
	LUT3 #(
		.INIT('h2a)
	) name17351 (
		\m1_data_i[4]_pad ,
		_w9137_,
		_w9138_,
		_w19252_
	);
	LUT4 #(
		.INIT('h37bf)
	) name17352 (
		_w9132_,
		_w9135_,
		_w19251_,
		_w19252_,
		_w19253_
	);
	LUT3 #(
		.INIT('h80)
	) name17353 (
		\m0_data_i[4]_pad ,
		_w9137_,
		_w9138_,
		_w19254_
	);
	LUT3 #(
		.INIT('h2a)
	) name17354 (
		\m7_data_i[4]_pad ,
		_w9137_,
		_w9138_,
		_w19255_
	);
	LUT4 #(
		.INIT('h6e7f)
	) name17355 (
		_w9132_,
		_w9135_,
		_w19254_,
		_w19255_,
		_w19256_
	);
	LUT4 #(
		.INIT('h7fff)
	) name17356 (
		_w19247_,
		_w19250_,
		_w19253_,
		_w19256_,
		_w19257_
	);
	LUT3 #(
		.INIT('h2a)
	) name17357 (
		\m3_data_i[5]_pad ,
		_w9137_,
		_w9138_,
		_w19258_
	);
	LUT3 #(
		.INIT('h80)
	) name17358 (
		\m4_data_i[5]_pad ,
		_w9137_,
		_w9138_,
		_w19259_
	);
	LUT4 #(
		.INIT('h9bdf)
	) name17359 (
		_w9132_,
		_w9135_,
		_w19258_,
		_w19259_,
		_w19260_
	);
	LUT3 #(
		.INIT('h80)
	) name17360 (
		\m6_data_i[5]_pad ,
		_w9137_,
		_w9138_,
		_w19261_
	);
	LUT3 #(
		.INIT('h80)
	) name17361 (
		\m2_data_i[5]_pad ,
		_w9137_,
		_w9138_,
		_w19262_
	);
	LUT4 #(
		.INIT('hcdef)
	) name17362 (
		_w9132_,
		_w9135_,
		_w19261_,
		_w19262_,
		_w19263_
	);
	LUT3 #(
		.INIT('h2a)
	) name17363 (
		\m5_data_i[5]_pad ,
		_w9137_,
		_w9138_,
		_w19264_
	);
	LUT3 #(
		.INIT('h2a)
	) name17364 (
		\m1_data_i[5]_pad ,
		_w9137_,
		_w9138_,
		_w19265_
	);
	LUT4 #(
		.INIT('h37bf)
	) name17365 (
		_w9132_,
		_w9135_,
		_w19264_,
		_w19265_,
		_w19266_
	);
	LUT3 #(
		.INIT('h80)
	) name17366 (
		\m0_data_i[5]_pad ,
		_w9137_,
		_w9138_,
		_w19267_
	);
	LUT3 #(
		.INIT('h2a)
	) name17367 (
		\m7_data_i[5]_pad ,
		_w9137_,
		_w9138_,
		_w19268_
	);
	LUT4 #(
		.INIT('h6e7f)
	) name17368 (
		_w9132_,
		_w9135_,
		_w19267_,
		_w19268_,
		_w19269_
	);
	LUT4 #(
		.INIT('h7fff)
	) name17369 (
		_w19260_,
		_w19263_,
		_w19266_,
		_w19269_,
		_w19270_
	);
	LUT3 #(
		.INIT('h2a)
	) name17370 (
		\m3_data_i[6]_pad ,
		_w9137_,
		_w9138_,
		_w19271_
	);
	LUT3 #(
		.INIT('h80)
	) name17371 (
		\m4_data_i[6]_pad ,
		_w9137_,
		_w9138_,
		_w19272_
	);
	LUT4 #(
		.INIT('h9bdf)
	) name17372 (
		_w9132_,
		_w9135_,
		_w19271_,
		_w19272_,
		_w19273_
	);
	LUT3 #(
		.INIT('h80)
	) name17373 (
		\m6_data_i[6]_pad ,
		_w9137_,
		_w9138_,
		_w19274_
	);
	LUT3 #(
		.INIT('h80)
	) name17374 (
		\m2_data_i[6]_pad ,
		_w9137_,
		_w9138_,
		_w19275_
	);
	LUT4 #(
		.INIT('hcdef)
	) name17375 (
		_w9132_,
		_w9135_,
		_w19274_,
		_w19275_,
		_w19276_
	);
	LUT3 #(
		.INIT('h2a)
	) name17376 (
		\m5_data_i[6]_pad ,
		_w9137_,
		_w9138_,
		_w19277_
	);
	LUT3 #(
		.INIT('h2a)
	) name17377 (
		\m1_data_i[6]_pad ,
		_w9137_,
		_w9138_,
		_w19278_
	);
	LUT4 #(
		.INIT('h37bf)
	) name17378 (
		_w9132_,
		_w9135_,
		_w19277_,
		_w19278_,
		_w19279_
	);
	LUT3 #(
		.INIT('h80)
	) name17379 (
		\m0_data_i[6]_pad ,
		_w9137_,
		_w9138_,
		_w19280_
	);
	LUT3 #(
		.INIT('h2a)
	) name17380 (
		\m7_data_i[6]_pad ,
		_w9137_,
		_w9138_,
		_w19281_
	);
	LUT4 #(
		.INIT('h6e7f)
	) name17381 (
		_w9132_,
		_w9135_,
		_w19280_,
		_w19281_,
		_w19282_
	);
	LUT4 #(
		.INIT('h7fff)
	) name17382 (
		_w19273_,
		_w19276_,
		_w19279_,
		_w19282_,
		_w19283_
	);
	LUT3 #(
		.INIT('h80)
	) name17383 (
		\m6_data_i[7]_pad ,
		_w9137_,
		_w9138_,
		_w19284_
	);
	LUT3 #(
		.INIT('h2a)
	) name17384 (
		\m5_data_i[7]_pad ,
		_w9137_,
		_w9138_,
		_w19285_
	);
	LUT4 #(
		.INIT('habef)
	) name17385 (
		_w9132_,
		_w9135_,
		_w19284_,
		_w19285_,
		_w19286_
	);
	LUT3 #(
		.INIT('h80)
	) name17386 (
		\m0_data_i[7]_pad ,
		_w9137_,
		_w9138_,
		_w19287_
	);
	LUT3 #(
		.INIT('h80)
	) name17387 (
		\m4_data_i[7]_pad ,
		_w9137_,
		_w9138_,
		_w19288_
	);
	LUT4 #(
		.INIT('h3b7f)
	) name17388 (
		_w9132_,
		_w9135_,
		_w19287_,
		_w19288_,
		_w19289_
	);
	LUT3 #(
		.INIT('h2a)
	) name17389 (
		\m7_data_i[7]_pad ,
		_w9137_,
		_w9138_,
		_w19290_
	);
	LUT3 #(
		.INIT('h2a)
	) name17390 (
		\m3_data_i[7]_pad ,
		_w9137_,
		_w9138_,
		_w19291_
	);
	LUT4 #(
		.INIT('hcdef)
	) name17391 (
		_w9132_,
		_w9135_,
		_w19290_,
		_w19291_,
		_w19292_
	);
	LUT3 #(
		.INIT('h2a)
	) name17392 (
		\m1_data_i[7]_pad ,
		_w9137_,
		_w9138_,
		_w19293_
	);
	LUT3 #(
		.INIT('h80)
	) name17393 (
		\m2_data_i[7]_pad ,
		_w9137_,
		_w9138_,
		_w19294_
	);
	LUT4 #(
		.INIT('h5d7f)
	) name17394 (
		_w9132_,
		_w9135_,
		_w19293_,
		_w19294_,
		_w19295_
	);
	LUT4 #(
		.INIT('h7fff)
	) name17395 (
		_w19286_,
		_w19289_,
		_w19292_,
		_w19295_,
		_w19296_
	);
	LUT3 #(
		.INIT('h2a)
	) name17396 (
		\m3_data_i[8]_pad ,
		_w9137_,
		_w9138_,
		_w19297_
	);
	LUT3 #(
		.INIT('h80)
	) name17397 (
		\m4_data_i[8]_pad ,
		_w9137_,
		_w9138_,
		_w19298_
	);
	LUT4 #(
		.INIT('h9bdf)
	) name17398 (
		_w9132_,
		_w9135_,
		_w19297_,
		_w19298_,
		_w19299_
	);
	LUT3 #(
		.INIT('h80)
	) name17399 (
		\m6_data_i[8]_pad ,
		_w9137_,
		_w9138_,
		_w19300_
	);
	LUT3 #(
		.INIT('h80)
	) name17400 (
		\m2_data_i[8]_pad ,
		_w9137_,
		_w9138_,
		_w19301_
	);
	LUT4 #(
		.INIT('hcdef)
	) name17401 (
		_w9132_,
		_w9135_,
		_w19300_,
		_w19301_,
		_w19302_
	);
	LUT3 #(
		.INIT('h2a)
	) name17402 (
		\m5_data_i[8]_pad ,
		_w9137_,
		_w9138_,
		_w19303_
	);
	LUT3 #(
		.INIT('h2a)
	) name17403 (
		\m1_data_i[8]_pad ,
		_w9137_,
		_w9138_,
		_w19304_
	);
	LUT4 #(
		.INIT('h37bf)
	) name17404 (
		_w9132_,
		_w9135_,
		_w19303_,
		_w19304_,
		_w19305_
	);
	LUT3 #(
		.INIT('h80)
	) name17405 (
		\m0_data_i[8]_pad ,
		_w9137_,
		_w9138_,
		_w19306_
	);
	LUT3 #(
		.INIT('h2a)
	) name17406 (
		\m7_data_i[8]_pad ,
		_w9137_,
		_w9138_,
		_w19307_
	);
	LUT4 #(
		.INIT('h6e7f)
	) name17407 (
		_w9132_,
		_w9135_,
		_w19306_,
		_w19307_,
		_w19308_
	);
	LUT4 #(
		.INIT('h7fff)
	) name17408 (
		_w19299_,
		_w19302_,
		_w19305_,
		_w19308_,
		_w19309_
	);
	LUT3 #(
		.INIT('h2a)
	) name17409 (
		\m3_data_i[9]_pad ,
		_w9137_,
		_w9138_,
		_w19310_
	);
	LUT3 #(
		.INIT('h80)
	) name17410 (
		\m4_data_i[9]_pad ,
		_w9137_,
		_w9138_,
		_w19311_
	);
	LUT4 #(
		.INIT('h9bdf)
	) name17411 (
		_w9132_,
		_w9135_,
		_w19310_,
		_w19311_,
		_w19312_
	);
	LUT3 #(
		.INIT('h80)
	) name17412 (
		\m6_data_i[9]_pad ,
		_w9137_,
		_w9138_,
		_w19313_
	);
	LUT3 #(
		.INIT('h80)
	) name17413 (
		\m2_data_i[9]_pad ,
		_w9137_,
		_w9138_,
		_w19314_
	);
	LUT4 #(
		.INIT('hcdef)
	) name17414 (
		_w9132_,
		_w9135_,
		_w19313_,
		_w19314_,
		_w19315_
	);
	LUT3 #(
		.INIT('h2a)
	) name17415 (
		\m5_data_i[9]_pad ,
		_w9137_,
		_w9138_,
		_w19316_
	);
	LUT3 #(
		.INIT('h2a)
	) name17416 (
		\m1_data_i[9]_pad ,
		_w9137_,
		_w9138_,
		_w19317_
	);
	LUT4 #(
		.INIT('h37bf)
	) name17417 (
		_w9132_,
		_w9135_,
		_w19316_,
		_w19317_,
		_w19318_
	);
	LUT3 #(
		.INIT('h80)
	) name17418 (
		\m0_data_i[9]_pad ,
		_w9137_,
		_w9138_,
		_w19319_
	);
	LUT3 #(
		.INIT('h2a)
	) name17419 (
		\m7_data_i[9]_pad ,
		_w9137_,
		_w9138_,
		_w19320_
	);
	LUT4 #(
		.INIT('h6e7f)
	) name17420 (
		_w9132_,
		_w9135_,
		_w19319_,
		_w19320_,
		_w19321_
	);
	LUT4 #(
		.INIT('h7fff)
	) name17421 (
		_w19312_,
		_w19315_,
		_w19318_,
		_w19321_,
		_w19322_
	);
	LUT3 #(
		.INIT('h2a)
	) name17422 (
		\m3_sel_i[0]_pad ,
		_w9137_,
		_w9138_,
		_w19323_
	);
	LUT3 #(
		.INIT('h80)
	) name17423 (
		\m4_sel_i[0]_pad ,
		_w9137_,
		_w9138_,
		_w19324_
	);
	LUT4 #(
		.INIT('h9bdf)
	) name17424 (
		_w9132_,
		_w9135_,
		_w19323_,
		_w19324_,
		_w19325_
	);
	LUT3 #(
		.INIT('h80)
	) name17425 (
		\m6_sel_i[0]_pad ,
		_w9137_,
		_w9138_,
		_w19326_
	);
	LUT3 #(
		.INIT('h80)
	) name17426 (
		\m2_sel_i[0]_pad ,
		_w9137_,
		_w9138_,
		_w19327_
	);
	LUT4 #(
		.INIT('hcdef)
	) name17427 (
		_w9132_,
		_w9135_,
		_w19326_,
		_w19327_,
		_w19328_
	);
	LUT3 #(
		.INIT('h2a)
	) name17428 (
		\m5_sel_i[0]_pad ,
		_w9137_,
		_w9138_,
		_w19329_
	);
	LUT3 #(
		.INIT('h2a)
	) name17429 (
		\m1_sel_i[0]_pad ,
		_w9137_,
		_w9138_,
		_w19330_
	);
	LUT4 #(
		.INIT('h37bf)
	) name17430 (
		_w9132_,
		_w9135_,
		_w19329_,
		_w19330_,
		_w19331_
	);
	LUT3 #(
		.INIT('h80)
	) name17431 (
		\m0_sel_i[0]_pad ,
		_w9137_,
		_w9138_,
		_w19332_
	);
	LUT3 #(
		.INIT('h2a)
	) name17432 (
		\m7_sel_i[0]_pad ,
		_w9137_,
		_w9138_,
		_w19333_
	);
	LUT4 #(
		.INIT('h6e7f)
	) name17433 (
		_w9132_,
		_w9135_,
		_w19332_,
		_w19333_,
		_w19334_
	);
	LUT4 #(
		.INIT('h7fff)
	) name17434 (
		_w19325_,
		_w19328_,
		_w19331_,
		_w19334_,
		_w19335_
	);
	LUT3 #(
		.INIT('h2a)
	) name17435 (
		\m3_sel_i[1]_pad ,
		_w9137_,
		_w9138_,
		_w19336_
	);
	LUT3 #(
		.INIT('h80)
	) name17436 (
		\m4_sel_i[1]_pad ,
		_w9137_,
		_w9138_,
		_w19337_
	);
	LUT4 #(
		.INIT('h9bdf)
	) name17437 (
		_w9132_,
		_w9135_,
		_w19336_,
		_w19337_,
		_w19338_
	);
	LUT3 #(
		.INIT('h80)
	) name17438 (
		\m6_sel_i[1]_pad ,
		_w9137_,
		_w9138_,
		_w19339_
	);
	LUT3 #(
		.INIT('h80)
	) name17439 (
		\m2_sel_i[1]_pad ,
		_w9137_,
		_w9138_,
		_w19340_
	);
	LUT4 #(
		.INIT('hcdef)
	) name17440 (
		_w9132_,
		_w9135_,
		_w19339_,
		_w19340_,
		_w19341_
	);
	LUT3 #(
		.INIT('h2a)
	) name17441 (
		\m5_sel_i[1]_pad ,
		_w9137_,
		_w9138_,
		_w19342_
	);
	LUT3 #(
		.INIT('h2a)
	) name17442 (
		\m1_sel_i[1]_pad ,
		_w9137_,
		_w9138_,
		_w19343_
	);
	LUT4 #(
		.INIT('h37bf)
	) name17443 (
		_w9132_,
		_w9135_,
		_w19342_,
		_w19343_,
		_w19344_
	);
	LUT3 #(
		.INIT('h80)
	) name17444 (
		\m0_sel_i[1]_pad ,
		_w9137_,
		_w9138_,
		_w19345_
	);
	LUT3 #(
		.INIT('h2a)
	) name17445 (
		\m7_sel_i[1]_pad ,
		_w9137_,
		_w9138_,
		_w19346_
	);
	LUT4 #(
		.INIT('h6e7f)
	) name17446 (
		_w9132_,
		_w9135_,
		_w19345_,
		_w19346_,
		_w19347_
	);
	LUT4 #(
		.INIT('h7fff)
	) name17447 (
		_w19338_,
		_w19341_,
		_w19344_,
		_w19347_,
		_w19348_
	);
	LUT3 #(
		.INIT('h80)
	) name17448 (
		\m6_sel_i[2]_pad ,
		_w9137_,
		_w9138_,
		_w19349_
	);
	LUT3 #(
		.INIT('h2a)
	) name17449 (
		\m5_sel_i[2]_pad ,
		_w9137_,
		_w9138_,
		_w19350_
	);
	LUT4 #(
		.INIT('habef)
	) name17450 (
		_w9132_,
		_w9135_,
		_w19349_,
		_w19350_,
		_w19351_
	);
	LUT3 #(
		.INIT('h2a)
	) name17451 (
		\m3_sel_i[2]_pad ,
		_w9137_,
		_w9138_,
		_w19352_
	);
	LUT3 #(
		.INIT('h80)
	) name17452 (
		\m2_sel_i[2]_pad ,
		_w9137_,
		_w9138_,
		_w19353_
	);
	LUT3 #(
		.INIT('h57)
	) name17453 (
		_w9144_,
		_w19352_,
		_w19353_,
		_w19354_
	);
	LUT3 #(
		.INIT('h80)
	) name17454 (
		\m4_sel_i[2]_pad ,
		_w9137_,
		_w9138_,
		_w19355_
	);
	LUT3 #(
		.INIT('h2a)
	) name17455 (
		\m1_sel_i[2]_pad ,
		_w9137_,
		_w9138_,
		_w19356_
	);
	LUT4 #(
		.INIT('h37bf)
	) name17456 (
		_w9132_,
		_w9135_,
		_w19355_,
		_w19356_,
		_w19357_
	);
	LUT3 #(
		.INIT('h80)
	) name17457 (
		\m0_sel_i[2]_pad ,
		_w9137_,
		_w9138_,
		_w19358_
	);
	LUT3 #(
		.INIT('h2a)
	) name17458 (
		\m7_sel_i[2]_pad ,
		_w9137_,
		_w9138_,
		_w19359_
	);
	LUT4 #(
		.INIT('h6e7f)
	) name17459 (
		_w9132_,
		_w9135_,
		_w19358_,
		_w19359_,
		_w19360_
	);
	LUT4 #(
		.INIT('h7fff)
	) name17460 (
		_w19351_,
		_w19354_,
		_w19357_,
		_w19360_,
		_w19361_
	);
	LUT3 #(
		.INIT('h2a)
	) name17461 (
		\m1_sel_i[3]_pad ,
		_w9137_,
		_w9138_,
		_w19362_
	);
	LUT3 #(
		.INIT('h80)
	) name17462 (
		\m2_sel_i[3]_pad ,
		_w9137_,
		_w9138_,
		_w19363_
	);
	LUT4 #(
		.INIT('h5d7f)
	) name17463 (
		_w9132_,
		_w9135_,
		_w19362_,
		_w19363_,
		_w19364_
	);
	LUT3 #(
		.INIT('h80)
	) name17464 (
		\m6_sel_i[3]_pad ,
		_w9137_,
		_w9138_,
		_w19365_
	);
	LUT3 #(
		.INIT('h80)
	) name17465 (
		\m4_sel_i[3]_pad ,
		_w9137_,
		_w9138_,
		_w19366_
	);
	LUT4 #(
		.INIT('habef)
	) name17466 (
		_w9132_,
		_w9135_,
		_w19365_,
		_w19366_,
		_w19367_
	);
	LUT3 #(
		.INIT('h2a)
	) name17467 (
		\m5_sel_i[3]_pad ,
		_w9137_,
		_w9138_,
		_w19368_
	);
	LUT3 #(
		.INIT('h2a)
	) name17468 (
		\m3_sel_i[3]_pad ,
		_w9137_,
		_w9138_,
		_w19369_
	);
	LUT4 #(
		.INIT('h9dbf)
	) name17469 (
		_w9132_,
		_w9135_,
		_w19368_,
		_w19369_,
		_w19370_
	);
	LUT3 #(
		.INIT('h80)
	) name17470 (
		\m0_sel_i[3]_pad ,
		_w9137_,
		_w9138_,
		_w19371_
	);
	LUT3 #(
		.INIT('h2a)
	) name17471 (
		\m7_sel_i[3]_pad ,
		_w9137_,
		_w9138_,
		_w19372_
	);
	LUT4 #(
		.INIT('h6e7f)
	) name17472 (
		_w9132_,
		_w9135_,
		_w19371_,
		_w19372_,
		_w19373_
	);
	LUT4 #(
		.INIT('h7fff)
	) name17473 (
		_w19364_,
		_w19367_,
		_w19370_,
		_w19373_,
		_w19374_
	);
	LUT4 #(
		.INIT('h2a00)
	) name17474 (
		\m3_stb_i_pad ,
		_w9137_,
		_w9138_,
		_w9497_,
		_w19375_
	);
	LUT4 #(
		.INIT('h8000)
	) name17475 (
		\m2_stb_i_pad ,
		_w9137_,
		_w9138_,
		_w9632_,
		_w19376_
	);
	LUT3 #(
		.INIT('h57)
	) name17476 (
		_w9144_,
		_w19375_,
		_w19376_,
		_w19377_
	);
	LUT4 #(
		.INIT('h8000)
	) name17477 (
		\m4_stb_i_pad ,
		_w9137_,
		_w9138_,
		_w9515_,
		_w19378_
	);
	LUT4 #(
		.INIT('h8000)
	) name17478 (
		\m6_stb_i_pad ,
		_w9137_,
		_w9138_,
		_w9571_,
		_w19379_
	);
	LUT4 #(
		.INIT('haebf)
	) name17479 (
		_w9132_,
		_w9135_,
		_w19378_,
		_w19379_,
		_w19380_
	);
	LUT4 #(
		.INIT('h2a00)
	) name17480 (
		\m5_stb_i_pad ,
		_w9137_,
		_w9138_,
		_w9348_,
		_w19381_
	);
	LUT4 #(
		.INIT('h2a00)
	) name17481 (
		\m7_stb_i_pad ,
		_w9137_,
		_w9138_,
		_w9603_,
		_w19382_
	);
	LUT4 #(
		.INIT('haebf)
	) name17482 (
		_w9132_,
		_w9135_,
		_w19381_,
		_w19382_,
		_w19383_
	);
	LUT4 #(
		.INIT('h2a00)
	) name17483 (
		\m1_stb_i_pad ,
		_w9137_,
		_w9138_,
		_w9422_,
		_w19384_
	);
	LUT4 #(
		.INIT('h8000)
	) name17484 (
		\m0_stb_i_pad ,
		_w9137_,
		_w9138_,
		_w9390_,
		_w19385_
	);
	LUT3 #(
		.INIT('h57)
	) name17485 (
		_w9136_,
		_w19384_,
		_w19385_,
		_w19386_
	);
	LUT4 #(
		.INIT('h7fff)
	) name17486 (
		_w19377_,
		_w19380_,
		_w19383_,
		_w19386_,
		_w19387_
	);
	LUT3 #(
		.INIT('h2a)
	) name17487 (
		\m3_we_i_pad ,
		_w9137_,
		_w9138_,
		_w19388_
	);
	LUT3 #(
		.INIT('h80)
	) name17488 (
		\m4_we_i_pad ,
		_w9137_,
		_w9138_,
		_w19389_
	);
	LUT4 #(
		.INIT('h9bdf)
	) name17489 (
		_w9132_,
		_w9135_,
		_w19388_,
		_w19389_,
		_w19390_
	);
	LUT3 #(
		.INIT('h80)
	) name17490 (
		\m6_we_i_pad ,
		_w9137_,
		_w9138_,
		_w19391_
	);
	LUT3 #(
		.INIT('h80)
	) name17491 (
		\m2_we_i_pad ,
		_w9137_,
		_w9138_,
		_w19392_
	);
	LUT4 #(
		.INIT('hcdef)
	) name17492 (
		_w9132_,
		_w9135_,
		_w19391_,
		_w19392_,
		_w19393_
	);
	LUT3 #(
		.INIT('h2a)
	) name17493 (
		\m5_we_i_pad ,
		_w9137_,
		_w9138_,
		_w19394_
	);
	LUT3 #(
		.INIT('h2a)
	) name17494 (
		\m1_we_i_pad ,
		_w9137_,
		_w9138_,
		_w19395_
	);
	LUT4 #(
		.INIT('h37bf)
	) name17495 (
		_w9132_,
		_w9135_,
		_w19394_,
		_w19395_,
		_w19396_
	);
	LUT3 #(
		.INIT('h80)
	) name17496 (
		\m0_we_i_pad ,
		_w9137_,
		_w9138_,
		_w19397_
	);
	LUT3 #(
		.INIT('h2a)
	) name17497 (
		\m7_we_i_pad ,
		_w9137_,
		_w9138_,
		_w19398_
	);
	LUT4 #(
		.INIT('h6e7f)
	) name17498 (
		_w9132_,
		_w9135_,
		_w19397_,
		_w19398_,
		_w19399_
	);
	LUT4 #(
		.INIT('h7fff)
	) name17499 (
		_w19390_,
		_w19393_,
		_w19396_,
		_w19399_,
		_w19400_
	);
	LUT3 #(
		.INIT('h2a)
	) name17500 (
		\m7_addr_i[0]_pad ,
		_w1901_,
		_w1902_,
		_w19401_
	);
	LUT3 #(
		.INIT('h2a)
	) name17501 (
		\m6_addr_i[0]_pad ,
		_w1908_,
		_w1909_,
		_w19402_
	);
	LUT4 #(
		.INIT('h153f)
	) name17502 (
		_w1907_,
		_w1918_,
		_w19401_,
		_w19402_,
		_w19403_
	);
	LUT3 #(
		.INIT('h2a)
	) name17503 (
		\m5_addr_i[0]_pad ,
		_w1901_,
		_w1902_,
		_w19404_
	);
	LUT3 #(
		.INIT('h2a)
	) name17504 (
		\m2_addr_i[0]_pad ,
		_w1908_,
		_w1909_,
		_w19405_
	);
	LUT4 #(
		.INIT('h153f)
	) name17505 (
		_w1914_,
		_w1920_,
		_w19404_,
		_w19405_,
		_w19406_
	);
	LUT3 #(
		.INIT('h80)
	) name17506 (
		\m4_addr_i[0]_pad ,
		_w1908_,
		_w1909_,
		_w19407_
	);
	LUT3 #(
		.INIT('h80)
	) name17507 (
		\m3_addr_i[0]_pad ,
		_w1901_,
		_w1902_,
		_w19408_
	);
	LUT4 #(
		.INIT('h135f)
	) name17508 (
		_w1907_,
		_w1918_,
		_w19407_,
		_w19408_,
		_w19409_
	);
	LUT3 #(
		.INIT('h80)
	) name17509 (
		\m1_addr_i[0]_pad ,
		_w1901_,
		_w1902_,
		_w19410_
	);
	LUT3 #(
		.INIT('h80)
	) name17510 (
		\m0_addr_i[0]_pad ,
		_w1908_,
		_w1909_,
		_w19411_
	);
	LUT4 #(
		.INIT('h153f)
	) name17511 (
		_w1914_,
		_w1920_,
		_w19410_,
		_w19411_,
		_w19412_
	);
	LUT4 #(
		.INIT('h7fff)
	) name17512 (
		_w19403_,
		_w19406_,
		_w19409_,
		_w19412_,
		_w19413_
	);
	LUT3 #(
		.INIT('h2a)
	) name17513 (
		\m7_addr_i[10]_pad ,
		_w1901_,
		_w1902_,
		_w19414_
	);
	LUT3 #(
		.INIT('h2a)
	) name17514 (
		\m6_addr_i[10]_pad ,
		_w1908_,
		_w1909_,
		_w19415_
	);
	LUT4 #(
		.INIT('h153f)
	) name17515 (
		_w1907_,
		_w1918_,
		_w19414_,
		_w19415_,
		_w19416_
	);
	LUT3 #(
		.INIT('h2a)
	) name17516 (
		\m5_addr_i[10]_pad ,
		_w1901_,
		_w1902_,
		_w19417_
	);
	LUT3 #(
		.INIT('h2a)
	) name17517 (
		\m2_addr_i[10]_pad ,
		_w1908_,
		_w1909_,
		_w19418_
	);
	LUT4 #(
		.INIT('h153f)
	) name17518 (
		_w1914_,
		_w1920_,
		_w19417_,
		_w19418_,
		_w19419_
	);
	LUT3 #(
		.INIT('h80)
	) name17519 (
		\m4_addr_i[10]_pad ,
		_w1908_,
		_w1909_,
		_w19420_
	);
	LUT3 #(
		.INIT('h80)
	) name17520 (
		\m3_addr_i[10]_pad ,
		_w1901_,
		_w1902_,
		_w19421_
	);
	LUT4 #(
		.INIT('h135f)
	) name17521 (
		_w1907_,
		_w1918_,
		_w19420_,
		_w19421_,
		_w19422_
	);
	LUT3 #(
		.INIT('h80)
	) name17522 (
		\m1_addr_i[10]_pad ,
		_w1901_,
		_w1902_,
		_w19423_
	);
	LUT3 #(
		.INIT('h80)
	) name17523 (
		\m0_addr_i[10]_pad ,
		_w1908_,
		_w1909_,
		_w19424_
	);
	LUT4 #(
		.INIT('h153f)
	) name17524 (
		_w1914_,
		_w1920_,
		_w19423_,
		_w19424_,
		_w19425_
	);
	LUT4 #(
		.INIT('h7fff)
	) name17525 (
		_w19416_,
		_w19419_,
		_w19422_,
		_w19425_,
		_w19426_
	);
	LUT3 #(
		.INIT('h2a)
	) name17526 (
		\m7_addr_i[11]_pad ,
		_w1901_,
		_w1902_,
		_w19427_
	);
	LUT3 #(
		.INIT('h2a)
	) name17527 (
		\m6_addr_i[11]_pad ,
		_w1908_,
		_w1909_,
		_w19428_
	);
	LUT4 #(
		.INIT('h153f)
	) name17528 (
		_w1907_,
		_w1918_,
		_w19427_,
		_w19428_,
		_w19429_
	);
	LUT3 #(
		.INIT('h2a)
	) name17529 (
		\m5_addr_i[11]_pad ,
		_w1901_,
		_w1902_,
		_w19430_
	);
	LUT3 #(
		.INIT('h2a)
	) name17530 (
		\m2_addr_i[11]_pad ,
		_w1908_,
		_w1909_,
		_w19431_
	);
	LUT4 #(
		.INIT('h153f)
	) name17531 (
		_w1914_,
		_w1920_,
		_w19430_,
		_w19431_,
		_w19432_
	);
	LUT3 #(
		.INIT('h80)
	) name17532 (
		\m4_addr_i[11]_pad ,
		_w1908_,
		_w1909_,
		_w19433_
	);
	LUT3 #(
		.INIT('h80)
	) name17533 (
		\m3_addr_i[11]_pad ,
		_w1901_,
		_w1902_,
		_w19434_
	);
	LUT4 #(
		.INIT('h135f)
	) name17534 (
		_w1907_,
		_w1918_,
		_w19433_,
		_w19434_,
		_w19435_
	);
	LUT3 #(
		.INIT('h80)
	) name17535 (
		\m1_addr_i[11]_pad ,
		_w1901_,
		_w1902_,
		_w19436_
	);
	LUT3 #(
		.INIT('h80)
	) name17536 (
		\m0_addr_i[11]_pad ,
		_w1908_,
		_w1909_,
		_w19437_
	);
	LUT4 #(
		.INIT('h153f)
	) name17537 (
		_w1914_,
		_w1920_,
		_w19436_,
		_w19437_,
		_w19438_
	);
	LUT4 #(
		.INIT('h7fff)
	) name17538 (
		_w19429_,
		_w19432_,
		_w19435_,
		_w19438_,
		_w19439_
	);
	LUT3 #(
		.INIT('h2a)
	) name17539 (
		\m7_addr_i[12]_pad ,
		_w1901_,
		_w1902_,
		_w19440_
	);
	LUT3 #(
		.INIT('h2a)
	) name17540 (
		\m6_addr_i[12]_pad ,
		_w1908_,
		_w1909_,
		_w19441_
	);
	LUT4 #(
		.INIT('h153f)
	) name17541 (
		_w1907_,
		_w1918_,
		_w19440_,
		_w19441_,
		_w19442_
	);
	LUT3 #(
		.INIT('h2a)
	) name17542 (
		\m5_addr_i[12]_pad ,
		_w1901_,
		_w1902_,
		_w19443_
	);
	LUT3 #(
		.INIT('h2a)
	) name17543 (
		\m2_addr_i[12]_pad ,
		_w1908_,
		_w1909_,
		_w19444_
	);
	LUT4 #(
		.INIT('h153f)
	) name17544 (
		_w1914_,
		_w1920_,
		_w19443_,
		_w19444_,
		_w19445_
	);
	LUT3 #(
		.INIT('h80)
	) name17545 (
		\m4_addr_i[12]_pad ,
		_w1908_,
		_w1909_,
		_w19446_
	);
	LUT3 #(
		.INIT('h80)
	) name17546 (
		\m3_addr_i[12]_pad ,
		_w1901_,
		_w1902_,
		_w19447_
	);
	LUT4 #(
		.INIT('h135f)
	) name17547 (
		_w1907_,
		_w1918_,
		_w19446_,
		_w19447_,
		_w19448_
	);
	LUT3 #(
		.INIT('h80)
	) name17548 (
		\m1_addr_i[12]_pad ,
		_w1901_,
		_w1902_,
		_w19449_
	);
	LUT3 #(
		.INIT('h80)
	) name17549 (
		\m0_addr_i[12]_pad ,
		_w1908_,
		_w1909_,
		_w19450_
	);
	LUT4 #(
		.INIT('h153f)
	) name17550 (
		_w1914_,
		_w1920_,
		_w19449_,
		_w19450_,
		_w19451_
	);
	LUT4 #(
		.INIT('h7fff)
	) name17551 (
		_w19442_,
		_w19445_,
		_w19448_,
		_w19451_,
		_w19452_
	);
	LUT3 #(
		.INIT('h2a)
	) name17552 (
		\m7_addr_i[13]_pad ,
		_w1901_,
		_w1902_,
		_w19453_
	);
	LUT3 #(
		.INIT('h2a)
	) name17553 (
		\m6_addr_i[13]_pad ,
		_w1908_,
		_w1909_,
		_w19454_
	);
	LUT4 #(
		.INIT('h153f)
	) name17554 (
		_w1907_,
		_w1918_,
		_w19453_,
		_w19454_,
		_w19455_
	);
	LUT3 #(
		.INIT('h2a)
	) name17555 (
		\m5_addr_i[13]_pad ,
		_w1901_,
		_w1902_,
		_w19456_
	);
	LUT3 #(
		.INIT('h2a)
	) name17556 (
		\m2_addr_i[13]_pad ,
		_w1908_,
		_w1909_,
		_w19457_
	);
	LUT4 #(
		.INIT('h153f)
	) name17557 (
		_w1914_,
		_w1920_,
		_w19456_,
		_w19457_,
		_w19458_
	);
	LUT3 #(
		.INIT('h80)
	) name17558 (
		\m4_addr_i[13]_pad ,
		_w1908_,
		_w1909_,
		_w19459_
	);
	LUT3 #(
		.INIT('h80)
	) name17559 (
		\m3_addr_i[13]_pad ,
		_w1901_,
		_w1902_,
		_w19460_
	);
	LUT4 #(
		.INIT('h135f)
	) name17560 (
		_w1907_,
		_w1918_,
		_w19459_,
		_w19460_,
		_w19461_
	);
	LUT3 #(
		.INIT('h80)
	) name17561 (
		\m1_addr_i[13]_pad ,
		_w1901_,
		_w1902_,
		_w19462_
	);
	LUT3 #(
		.INIT('h80)
	) name17562 (
		\m0_addr_i[13]_pad ,
		_w1908_,
		_w1909_,
		_w19463_
	);
	LUT4 #(
		.INIT('h153f)
	) name17563 (
		_w1914_,
		_w1920_,
		_w19462_,
		_w19463_,
		_w19464_
	);
	LUT4 #(
		.INIT('h7fff)
	) name17564 (
		_w19455_,
		_w19458_,
		_w19461_,
		_w19464_,
		_w19465_
	);
	LUT3 #(
		.INIT('h2a)
	) name17565 (
		\m7_addr_i[14]_pad ,
		_w1901_,
		_w1902_,
		_w19466_
	);
	LUT3 #(
		.INIT('h2a)
	) name17566 (
		\m6_addr_i[14]_pad ,
		_w1908_,
		_w1909_,
		_w19467_
	);
	LUT4 #(
		.INIT('h153f)
	) name17567 (
		_w1907_,
		_w1918_,
		_w19466_,
		_w19467_,
		_w19468_
	);
	LUT3 #(
		.INIT('h2a)
	) name17568 (
		\m5_addr_i[14]_pad ,
		_w1901_,
		_w1902_,
		_w19469_
	);
	LUT3 #(
		.INIT('h2a)
	) name17569 (
		\m2_addr_i[14]_pad ,
		_w1908_,
		_w1909_,
		_w19470_
	);
	LUT4 #(
		.INIT('h153f)
	) name17570 (
		_w1914_,
		_w1920_,
		_w19469_,
		_w19470_,
		_w19471_
	);
	LUT3 #(
		.INIT('h80)
	) name17571 (
		\m4_addr_i[14]_pad ,
		_w1908_,
		_w1909_,
		_w19472_
	);
	LUT3 #(
		.INIT('h80)
	) name17572 (
		\m3_addr_i[14]_pad ,
		_w1901_,
		_w1902_,
		_w19473_
	);
	LUT4 #(
		.INIT('h135f)
	) name17573 (
		_w1907_,
		_w1918_,
		_w19472_,
		_w19473_,
		_w19474_
	);
	LUT3 #(
		.INIT('h80)
	) name17574 (
		\m1_addr_i[14]_pad ,
		_w1901_,
		_w1902_,
		_w19475_
	);
	LUT3 #(
		.INIT('h80)
	) name17575 (
		\m0_addr_i[14]_pad ,
		_w1908_,
		_w1909_,
		_w19476_
	);
	LUT4 #(
		.INIT('h153f)
	) name17576 (
		_w1914_,
		_w1920_,
		_w19475_,
		_w19476_,
		_w19477_
	);
	LUT4 #(
		.INIT('h7fff)
	) name17577 (
		_w19468_,
		_w19471_,
		_w19474_,
		_w19477_,
		_w19478_
	);
	LUT3 #(
		.INIT('h80)
	) name17578 (
		\m3_addr_i[15]_pad ,
		_w1901_,
		_w1902_,
		_w19479_
	);
	LUT3 #(
		.INIT('h2a)
	) name17579 (
		\m2_addr_i[15]_pad ,
		_w1908_,
		_w1909_,
		_w19480_
	);
	LUT4 #(
		.INIT('h153f)
	) name17580 (
		_w1914_,
		_w1918_,
		_w19479_,
		_w19480_,
		_w19481_
	);
	LUT3 #(
		.INIT('h2a)
	) name17581 (
		\m5_addr_i[15]_pad ,
		_w1901_,
		_w1902_,
		_w19482_
	);
	LUT3 #(
		.INIT('h80)
	) name17582 (
		\m0_addr_i[15]_pad ,
		_w1908_,
		_w1909_,
		_w19483_
	);
	LUT4 #(
		.INIT('h153f)
	) name17583 (
		_w1914_,
		_w1920_,
		_w19482_,
		_w19483_,
		_w19484_
	);
	LUT3 #(
		.INIT('h80)
	) name17584 (
		\m4_addr_i[15]_pad ,
		_w1908_,
		_w1909_,
		_w19485_
	);
	LUT3 #(
		.INIT('h80)
	) name17585 (
		\m1_addr_i[15]_pad ,
		_w1901_,
		_w1902_,
		_w19486_
	);
	LUT4 #(
		.INIT('h135f)
	) name17586 (
		_w1907_,
		_w1920_,
		_w19485_,
		_w19486_,
		_w19487_
	);
	LUT3 #(
		.INIT('h2a)
	) name17587 (
		\m7_addr_i[15]_pad ,
		_w1901_,
		_w1902_,
		_w19488_
	);
	LUT3 #(
		.INIT('h2a)
	) name17588 (
		\m6_addr_i[15]_pad ,
		_w1908_,
		_w1909_,
		_w19489_
	);
	LUT4 #(
		.INIT('h153f)
	) name17589 (
		_w1907_,
		_w1918_,
		_w19488_,
		_w19489_,
		_w19490_
	);
	LUT4 #(
		.INIT('h7fff)
	) name17590 (
		_w19481_,
		_w19484_,
		_w19487_,
		_w19490_,
		_w19491_
	);
	LUT3 #(
		.INIT('h2a)
	) name17591 (
		\m7_addr_i[16]_pad ,
		_w1901_,
		_w1902_,
		_w19492_
	);
	LUT3 #(
		.INIT('h2a)
	) name17592 (
		\m6_addr_i[16]_pad ,
		_w1908_,
		_w1909_,
		_w19493_
	);
	LUT4 #(
		.INIT('h153f)
	) name17593 (
		_w1907_,
		_w1918_,
		_w19492_,
		_w19493_,
		_w19494_
	);
	LUT3 #(
		.INIT('h2a)
	) name17594 (
		\m5_addr_i[16]_pad ,
		_w1901_,
		_w1902_,
		_w19495_
	);
	LUT3 #(
		.INIT('h2a)
	) name17595 (
		\m2_addr_i[16]_pad ,
		_w1908_,
		_w1909_,
		_w19496_
	);
	LUT4 #(
		.INIT('h153f)
	) name17596 (
		_w1914_,
		_w1920_,
		_w19495_,
		_w19496_,
		_w19497_
	);
	LUT3 #(
		.INIT('h80)
	) name17597 (
		\m4_addr_i[16]_pad ,
		_w1908_,
		_w1909_,
		_w19498_
	);
	LUT3 #(
		.INIT('h80)
	) name17598 (
		\m3_addr_i[16]_pad ,
		_w1901_,
		_w1902_,
		_w19499_
	);
	LUT4 #(
		.INIT('h135f)
	) name17599 (
		_w1907_,
		_w1918_,
		_w19498_,
		_w19499_,
		_w19500_
	);
	LUT3 #(
		.INIT('h80)
	) name17600 (
		\m1_addr_i[16]_pad ,
		_w1901_,
		_w1902_,
		_w19501_
	);
	LUT3 #(
		.INIT('h80)
	) name17601 (
		\m0_addr_i[16]_pad ,
		_w1908_,
		_w1909_,
		_w19502_
	);
	LUT4 #(
		.INIT('h153f)
	) name17602 (
		_w1914_,
		_w1920_,
		_w19501_,
		_w19502_,
		_w19503_
	);
	LUT4 #(
		.INIT('h7fff)
	) name17603 (
		_w19494_,
		_w19497_,
		_w19500_,
		_w19503_,
		_w19504_
	);
	LUT3 #(
		.INIT('h2a)
	) name17604 (
		\m5_addr_i[17]_pad ,
		_w1901_,
		_w1902_,
		_w19505_
	);
	LUT3 #(
		.INIT('h80)
	) name17605 (
		\m4_addr_i[17]_pad ,
		_w1908_,
		_w1909_,
		_w19506_
	);
	LUT4 #(
		.INIT('h153f)
	) name17606 (
		_w1907_,
		_w1920_,
		_w19505_,
		_w19506_,
		_w19507_
	);
	LUT3 #(
		.INIT('h2a)
	) name17607 (
		\m7_addr_i[17]_pad ,
		_w1901_,
		_w1902_,
		_w19508_
	);
	LUT3 #(
		.INIT('h2a)
	) name17608 (
		\m2_addr_i[17]_pad ,
		_w1908_,
		_w1909_,
		_w19509_
	);
	LUT4 #(
		.INIT('h153f)
	) name17609 (
		_w1914_,
		_w1918_,
		_w19508_,
		_w19509_,
		_w19510_
	);
	LUT3 #(
		.INIT('h2a)
	) name17610 (
		\m6_addr_i[17]_pad ,
		_w1908_,
		_w1909_,
		_w19511_
	);
	LUT3 #(
		.INIT('h80)
	) name17611 (
		\m3_addr_i[17]_pad ,
		_w1901_,
		_w1902_,
		_w19512_
	);
	LUT4 #(
		.INIT('h135f)
	) name17612 (
		_w1907_,
		_w1918_,
		_w19511_,
		_w19512_,
		_w19513_
	);
	LUT3 #(
		.INIT('h80)
	) name17613 (
		\m1_addr_i[17]_pad ,
		_w1901_,
		_w1902_,
		_w19514_
	);
	LUT3 #(
		.INIT('h80)
	) name17614 (
		\m0_addr_i[17]_pad ,
		_w1908_,
		_w1909_,
		_w19515_
	);
	LUT4 #(
		.INIT('h153f)
	) name17615 (
		_w1914_,
		_w1920_,
		_w19514_,
		_w19515_,
		_w19516_
	);
	LUT4 #(
		.INIT('h7fff)
	) name17616 (
		_w19507_,
		_w19510_,
		_w19513_,
		_w19516_,
		_w19517_
	);
	LUT3 #(
		.INIT('h2a)
	) name17617 (
		\m7_addr_i[18]_pad ,
		_w1901_,
		_w1902_,
		_w19518_
	);
	LUT3 #(
		.INIT('h2a)
	) name17618 (
		\m6_addr_i[18]_pad ,
		_w1908_,
		_w1909_,
		_w19519_
	);
	LUT4 #(
		.INIT('h153f)
	) name17619 (
		_w1907_,
		_w1918_,
		_w19518_,
		_w19519_,
		_w19520_
	);
	LUT3 #(
		.INIT('h2a)
	) name17620 (
		\m5_addr_i[18]_pad ,
		_w1901_,
		_w1902_,
		_w19521_
	);
	LUT3 #(
		.INIT('h2a)
	) name17621 (
		\m2_addr_i[18]_pad ,
		_w1908_,
		_w1909_,
		_w19522_
	);
	LUT4 #(
		.INIT('h153f)
	) name17622 (
		_w1914_,
		_w1920_,
		_w19521_,
		_w19522_,
		_w19523_
	);
	LUT3 #(
		.INIT('h80)
	) name17623 (
		\m4_addr_i[18]_pad ,
		_w1908_,
		_w1909_,
		_w19524_
	);
	LUT3 #(
		.INIT('h80)
	) name17624 (
		\m3_addr_i[18]_pad ,
		_w1901_,
		_w1902_,
		_w19525_
	);
	LUT4 #(
		.INIT('h135f)
	) name17625 (
		_w1907_,
		_w1918_,
		_w19524_,
		_w19525_,
		_w19526_
	);
	LUT3 #(
		.INIT('h80)
	) name17626 (
		\m1_addr_i[18]_pad ,
		_w1901_,
		_w1902_,
		_w19527_
	);
	LUT3 #(
		.INIT('h80)
	) name17627 (
		\m0_addr_i[18]_pad ,
		_w1908_,
		_w1909_,
		_w19528_
	);
	LUT4 #(
		.INIT('h153f)
	) name17628 (
		_w1914_,
		_w1920_,
		_w19527_,
		_w19528_,
		_w19529_
	);
	LUT4 #(
		.INIT('h7fff)
	) name17629 (
		_w19520_,
		_w19523_,
		_w19526_,
		_w19529_,
		_w19530_
	);
	LUT3 #(
		.INIT('h2a)
	) name17630 (
		\m7_addr_i[19]_pad ,
		_w1901_,
		_w1902_,
		_w19531_
	);
	LUT3 #(
		.INIT('h2a)
	) name17631 (
		\m6_addr_i[19]_pad ,
		_w1908_,
		_w1909_,
		_w19532_
	);
	LUT4 #(
		.INIT('h153f)
	) name17632 (
		_w1907_,
		_w1918_,
		_w19531_,
		_w19532_,
		_w19533_
	);
	LUT3 #(
		.INIT('h2a)
	) name17633 (
		\m5_addr_i[19]_pad ,
		_w1901_,
		_w1902_,
		_w19534_
	);
	LUT3 #(
		.INIT('h2a)
	) name17634 (
		\m2_addr_i[19]_pad ,
		_w1908_,
		_w1909_,
		_w19535_
	);
	LUT4 #(
		.INIT('h153f)
	) name17635 (
		_w1914_,
		_w1920_,
		_w19534_,
		_w19535_,
		_w19536_
	);
	LUT3 #(
		.INIT('h80)
	) name17636 (
		\m4_addr_i[19]_pad ,
		_w1908_,
		_w1909_,
		_w19537_
	);
	LUT3 #(
		.INIT('h80)
	) name17637 (
		\m3_addr_i[19]_pad ,
		_w1901_,
		_w1902_,
		_w19538_
	);
	LUT4 #(
		.INIT('h135f)
	) name17638 (
		_w1907_,
		_w1918_,
		_w19537_,
		_w19538_,
		_w19539_
	);
	LUT3 #(
		.INIT('h80)
	) name17639 (
		\m1_addr_i[19]_pad ,
		_w1901_,
		_w1902_,
		_w19540_
	);
	LUT3 #(
		.INIT('h80)
	) name17640 (
		\m0_addr_i[19]_pad ,
		_w1908_,
		_w1909_,
		_w19541_
	);
	LUT4 #(
		.INIT('h153f)
	) name17641 (
		_w1914_,
		_w1920_,
		_w19540_,
		_w19541_,
		_w19542_
	);
	LUT4 #(
		.INIT('h7fff)
	) name17642 (
		_w19533_,
		_w19536_,
		_w19539_,
		_w19542_,
		_w19543_
	);
	LUT3 #(
		.INIT('h2a)
	) name17643 (
		\m7_addr_i[1]_pad ,
		_w1901_,
		_w1902_,
		_w19544_
	);
	LUT3 #(
		.INIT('h2a)
	) name17644 (
		\m6_addr_i[1]_pad ,
		_w1908_,
		_w1909_,
		_w19545_
	);
	LUT4 #(
		.INIT('h153f)
	) name17645 (
		_w1907_,
		_w1918_,
		_w19544_,
		_w19545_,
		_w19546_
	);
	LUT3 #(
		.INIT('h2a)
	) name17646 (
		\m5_addr_i[1]_pad ,
		_w1901_,
		_w1902_,
		_w19547_
	);
	LUT3 #(
		.INIT('h2a)
	) name17647 (
		\m2_addr_i[1]_pad ,
		_w1908_,
		_w1909_,
		_w19548_
	);
	LUT4 #(
		.INIT('h153f)
	) name17648 (
		_w1914_,
		_w1920_,
		_w19547_,
		_w19548_,
		_w19549_
	);
	LUT3 #(
		.INIT('h80)
	) name17649 (
		\m4_addr_i[1]_pad ,
		_w1908_,
		_w1909_,
		_w19550_
	);
	LUT3 #(
		.INIT('h80)
	) name17650 (
		\m3_addr_i[1]_pad ,
		_w1901_,
		_w1902_,
		_w19551_
	);
	LUT4 #(
		.INIT('h135f)
	) name17651 (
		_w1907_,
		_w1918_,
		_w19550_,
		_w19551_,
		_w19552_
	);
	LUT3 #(
		.INIT('h80)
	) name17652 (
		\m1_addr_i[1]_pad ,
		_w1901_,
		_w1902_,
		_w19553_
	);
	LUT3 #(
		.INIT('h80)
	) name17653 (
		\m0_addr_i[1]_pad ,
		_w1908_,
		_w1909_,
		_w19554_
	);
	LUT4 #(
		.INIT('h153f)
	) name17654 (
		_w1914_,
		_w1920_,
		_w19553_,
		_w19554_,
		_w19555_
	);
	LUT4 #(
		.INIT('h7fff)
	) name17655 (
		_w19546_,
		_w19549_,
		_w19552_,
		_w19555_,
		_w19556_
	);
	LUT3 #(
		.INIT('h2a)
	) name17656 (
		\m7_addr_i[20]_pad ,
		_w1901_,
		_w1902_,
		_w19557_
	);
	LUT3 #(
		.INIT('h2a)
	) name17657 (
		\m6_addr_i[20]_pad ,
		_w1908_,
		_w1909_,
		_w19558_
	);
	LUT4 #(
		.INIT('h153f)
	) name17658 (
		_w1907_,
		_w1918_,
		_w19557_,
		_w19558_,
		_w19559_
	);
	LUT3 #(
		.INIT('h2a)
	) name17659 (
		\m5_addr_i[20]_pad ,
		_w1901_,
		_w1902_,
		_w19560_
	);
	LUT3 #(
		.INIT('h2a)
	) name17660 (
		\m2_addr_i[20]_pad ,
		_w1908_,
		_w1909_,
		_w19561_
	);
	LUT4 #(
		.INIT('h153f)
	) name17661 (
		_w1914_,
		_w1920_,
		_w19560_,
		_w19561_,
		_w19562_
	);
	LUT3 #(
		.INIT('h80)
	) name17662 (
		\m4_addr_i[20]_pad ,
		_w1908_,
		_w1909_,
		_w19563_
	);
	LUT3 #(
		.INIT('h80)
	) name17663 (
		\m3_addr_i[20]_pad ,
		_w1901_,
		_w1902_,
		_w19564_
	);
	LUT4 #(
		.INIT('h135f)
	) name17664 (
		_w1907_,
		_w1918_,
		_w19563_,
		_w19564_,
		_w19565_
	);
	LUT3 #(
		.INIT('h80)
	) name17665 (
		\m1_addr_i[20]_pad ,
		_w1901_,
		_w1902_,
		_w19566_
	);
	LUT3 #(
		.INIT('h80)
	) name17666 (
		\m0_addr_i[20]_pad ,
		_w1908_,
		_w1909_,
		_w19567_
	);
	LUT4 #(
		.INIT('h153f)
	) name17667 (
		_w1914_,
		_w1920_,
		_w19566_,
		_w19567_,
		_w19568_
	);
	LUT4 #(
		.INIT('h7fff)
	) name17668 (
		_w19559_,
		_w19562_,
		_w19565_,
		_w19568_,
		_w19569_
	);
	LUT3 #(
		.INIT('h80)
	) name17669 (
		\m3_addr_i[21]_pad ,
		_w1901_,
		_w1902_,
		_w19570_
	);
	LUT3 #(
		.INIT('h2a)
	) name17670 (
		\m2_addr_i[21]_pad ,
		_w1908_,
		_w1909_,
		_w19571_
	);
	LUT4 #(
		.INIT('h153f)
	) name17671 (
		_w1914_,
		_w1918_,
		_w19570_,
		_w19571_,
		_w19572_
	);
	LUT3 #(
		.INIT('h2a)
	) name17672 (
		\m5_addr_i[21]_pad ,
		_w1901_,
		_w1902_,
		_w19573_
	);
	LUT3 #(
		.INIT('h80)
	) name17673 (
		\m0_addr_i[21]_pad ,
		_w1908_,
		_w1909_,
		_w19574_
	);
	LUT4 #(
		.INIT('h153f)
	) name17674 (
		_w1914_,
		_w1920_,
		_w19573_,
		_w19574_,
		_w19575_
	);
	LUT3 #(
		.INIT('h80)
	) name17675 (
		\m4_addr_i[21]_pad ,
		_w1908_,
		_w1909_,
		_w19576_
	);
	LUT3 #(
		.INIT('h80)
	) name17676 (
		\m1_addr_i[21]_pad ,
		_w1901_,
		_w1902_,
		_w19577_
	);
	LUT4 #(
		.INIT('h135f)
	) name17677 (
		_w1907_,
		_w1920_,
		_w19576_,
		_w19577_,
		_w19578_
	);
	LUT3 #(
		.INIT('h2a)
	) name17678 (
		\m7_addr_i[21]_pad ,
		_w1901_,
		_w1902_,
		_w19579_
	);
	LUT3 #(
		.INIT('h2a)
	) name17679 (
		\m6_addr_i[21]_pad ,
		_w1908_,
		_w1909_,
		_w19580_
	);
	LUT4 #(
		.INIT('h153f)
	) name17680 (
		_w1907_,
		_w1918_,
		_w19579_,
		_w19580_,
		_w19581_
	);
	LUT4 #(
		.INIT('h7fff)
	) name17681 (
		_w19572_,
		_w19575_,
		_w19578_,
		_w19581_,
		_w19582_
	);
	LUT3 #(
		.INIT('h2a)
	) name17682 (
		\m7_addr_i[22]_pad ,
		_w1901_,
		_w1902_,
		_w19583_
	);
	LUT3 #(
		.INIT('h2a)
	) name17683 (
		\m6_addr_i[22]_pad ,
		_w1908_,
		_w1909_,
		_w19584_
	);
	LUT4 #(
		.INIT('h153f)
	) name17684 (
		_w1907_,
		_w1918_,
		_w19583_,
		_w19584_,
		_w19585_
	);
	LUT3 #(
		.INIT('h2a)
	) name17685 (
		\m5_addr_i[22]_pad ,
		_w1901_,
		_w1902_,
		_w19586_
	);
	LUT3 #(
		.INIT('h2a)
	) name17686 (
		\m2_addr_i[22]_pad ,
		_w1908_,
		_w1909_,
		_w19587_
	);
	LUT4 #(
		.INIT('h153f)
	) name17687 (
		_w1914_,
		_w1920_,
		_w19586_,
		_w19587_,
		_w19588_
	);
	LUT3 #(
		.INIT('h80)
	) name17688 (
		\m4_addr_i[22]_pad ,
		_w1908_,
		_w1909_,
		_w19589_
	);
	LUT3 #(
		.INIT('h80)
	) name17689 (
		\m3_addr_i[22]_pad ,
		_w1901_,
		_w1902_,
		_w19590_
	);
	LUT4 #(
		.INIT('h135f)
	) name17690 (
		_w1907_,
		_w1918_,
		_w19589_,
		_w19590_,
		_w19591_
	);
	LUT3 #(
		.INIT('h80)
	) name17691 (
		\m1_addr_i[22]_pad ,
		_w1901_,
		_w1902_,
		_w19592_
	);
	LUT3 #(
		.INIT('h80)
	) name17692 (
		\m0_addr_i[22]_pad ,
		_w1908_,
		_w1909_,
		_w19593_
	);
	LUT4 #(
		.INIT('h153f)
	) name17693 (
		_w1914_,
		_w1920_,
		_w19592_,
		_w19593_,
		_w19594_
	);
	LUT4 #(
		.INIT('h7fff)
	) name17694 (
		_w19585_,
		_w19588_,
		_w19591_,
		_w19594_,
		_w19595_
	);
	LUT3 #(
		.INIT('h2a)
	) name17695 (
		\m7_addr_i[23]_pad ,
		_w1901_,
		_w1902_,
		_w19596_
	);
	LUT3 #(
		.INIT('h2a)
	) name17696 (
		\m6_addr_i[23]_pad ,
		_w1908_,
		_w1909_,
		_w19597_
	);
	LUT4 #(
		.INIT('h153f)
	) name17697 (
		_w1907_,
		_w1918_,
		_w19596_,
		_w19597_,
		_w19598_
	);
	LUT3 #(
		.INIT('h2a)
	) name17698 (
		\m5_addr_i[23]_pad ,
		_w1901_,
		_w1902_,
		_w19599_
	);
	LUT3 #(
		.INIT('h2a)
	) name17699 (
		\m2_addr_i[23]_pad ,
		_w1908_,
		_w1909_,
		_w19600_
	);
	LUT4 #(
		.INIT('h153f)
	) name17700 (
		_w1914_,
		_w1920_,
		_w19599_,
		_w19600_,
		_w19601_
	);
	LUT3 #(
		.INIT('h80)
	) name17701 (
		\m4_addr_i[23]_pad ,
		_w1908_,
		_w1909_,
		_w19602_
	);
	LUT3 #(
		.INIT('h80)
	) name17702 (
		\m3_addr_i[23]_pad ,
		_w1901_,
		_w1902_,
		_w19603_
	);
	LUT4 #(
		.INIT('h135f)
	) name17703 (
		_w1907_,
		_w1918_,
		_w19602_,
		_w19603_,
		_w19604_
	);
	LUT3 #(
		.INIT('h80)
	) name17704 (
		\m1_addr_i[23]_pad ,
		_w1901_,
		_w1902_,
		_w19605_
	);
	LUT3 #(
		.INIT('h80)
	) name17705 (
		\m0_addr_i[23]_pad ,
		_w1908_,
		_w1909_,
		_w19606_
	);
	LUT4 #(
		.INIT('h153f)
	) name17706 (
		_w1914_,
		_w1920_,
		_w19605_,
		_w19606_,
		_w19607_
	);
	LUT4 #(
		.INIT('h7fff)
	) name17707 (
		_w19598_,
		_w19601_,
		_w19604_,
		_w19607_,
		_w19608_
	);
	LUT3 #(
		.INIT('h80)
	) name17708 (
		\m4_addr_i[28]_pad ,
		_w1908_,
		_w1909_,
		_w19609_
	);
	LUT3 #(
		.INIT('h80)
	) name17709 (
		\m3_addr_i[28]_pad ,
		_w1901_,
		_w1902_,
		_w19610_
	);
	LUT4 #(
		.INIT('h135f)
	) name17710 (
		_w1907_,
		_w1918_,
		_w19609_,
		_w19610_,
		_w19611_
	);
	LUT3 #(
		.INIT('h80)
	) name17711 (
		\m1_addr_i[28]_pad ,
		_w1901_,
		_w1902_,
		_w19612_
	);
	LUT3 #(
		.INIT('h2a)
	) name17712 (
		\m6_addr_i[28]_pad ,
		_w1908_,
		_w1909_,
		_w19613_
	);
	LUT4 #(
		.INIT('h153f)
	) name17713 (
		_w1907_,
		_w1920_,
		_w19612_,
		_w19613_,
		_w19614_
	);
	LUT3 #(
		.INIT('h2a)
	) name17714 (
		\m2_addr_i[28]_pad ,
		_w1908_,
		_w1909_,
		_w19615_
	);
	LUT3 #(
		.INIT('h2a)
	) name17715 (
		\m5_addr_i[28]_pad ,
		_w1901_,
		_w1902_,
		_w19616_
	);
	LUT4 #(
		.INIT('h135f)
	) name17716 (
		_w1914_,
		_w1920_,
		_w19615_,
		_w19616_,
		_w19617_
	);
	LUT3 #(
		.INIT('h80)
	) name17717 (
		\m0_addr_i[28]_pad ,
		_w1908_,
		_w1909_,
		_w19618_
	);
	LUT3 #(
		.INIT('h2a)
	) name17718 (
		\m7_addr_i[28]_pad ,
		_w1901_,
		_w1902_,
		_w19619_
	);
	LUT4 #(
		.INIT('h135f)
	) name17719 (
		_w1914_,
		_w1918_,
		_w19618_,
		_w19619_,
		_w19620_
	);
	LUT4 #(
		.INIT('h7fff)
	) name17720 (
		_w19611_,
		_w19614_,
		_w19617_,
		_w19620_,
		_w19621_
	);
	LUT3 #(
		.INIT('h80)
	) name17721 (
		\m1_addr_i[29]_pad ,
		_w1901_,
		_w1902_,
		_w19622_
	);
	LUT3 #(
		.INIT('h2a)
	) name17722 (
		\m2_addr_i[29]_pad ,
		_w1908_,
		_w1909_,
		_w19623_
	);
	LUT4 #(
		.INIT('h153f)
	) name17723 (
		_w1914_,
		_w1920_,
		_w19622_,
		_w19623_,
		_w19624_
	);
	LUT3 #(
		.INIT('h80)
	) name17724 (
		\m0_addr_i[29]_pad ,
		_w1908_,
		_w1909_,
		_w19625_
	);
	LUT3 #(
		.INIT('h80)
	) name17725 (
		\m3_addr_i[29]_pad ,
		_w1901_,
		_w1902_,
		_w19626_
	);
	LUT4 #(
		.INIT('h135f)
	) name17726 (
		_w1914_,
		_w1918_,
		_w19625_,
		_w19626_,
		_w19627_
	);
	LUT3 #(
		.INIT('h2a)
	) name17727 (
		\m7_addr_i[29]_pad ,
		_w1901_,
		_w1902_,
		_w19628_
	);
	LUT3 #(
		.INIT('h80)
	) name17728 (
		\m4_addr_i[29]_pad ,
		_w1908_,
		_w1909_,
		_w19629_
	);
	LUT4 #(
		.INIT('h153f)
	) name17729 (
		_w1907_,
		_w1918_,
		_w19628_,
		_w19629_,
		_w19630_
	);
	LUT3 #(
		.INIT('h2a)
	) name17730 (
		\m5_addr_i[29]_pad ,
		_w1901_,
		_w1902_,
		_w19631_
	);
	LUT3 #(
		.INIT('h2a)
	) name17731 (
		\m6_addr_i[29]_pad ,
		_w1908_,
		_w1909_,
		_w19632_
	);
	LUT4 #(
		.INIT('h153f)
	) name17732 (
		_w1907_,
		_w1920_,
		_w19631_,
		_w19632_,
		_w19633_
	);
	LUT4 #(
		.INIT('h7fff)
	) name17733 (
		_w19624_,
		_w19627_,
		_w19630_,
		_w19633_,
		_w19634_
	);
	LUT3 #(
		.INIT('h80)
	) name17734 (
		\m4_addr_i[30]_pad ,
		_w1908_,
		_w1909_,
		_w19635_
	);
	LUT3 #(
		.INIT('h80)
	) name17735 (
		\m3_addr_i[30]_pad ,
		_w1901_,
		_w1902_,
		_w19636_
	);
	LUT4 #(
		.INIT('h135f)
	) name17736 (
		_w1907_,
		_w1918_,
		_w19635_,
		_w19636_,
		_w19637_
	);
	LUT3 #(
		.INIT('h80)
	) name17737 (
		\m1_addr_i[30]_pad ,
		_w1901_,
		_w1902_,
		_w19638_
	);
	LUT3 #(
		.INIT('h2a)
	) name17738 (
		\m6_addr_i[30]_pad ,
		_w1908_,
		_w1909_,
		_w19639_
	);
	LUT4 #(
		.INIT('h153f)
	) name17739 (
		_w1907_,
		_w1920_,
		_w19638_,
		_w19639_,
		_w19640_
	);
	LUT3 #(
		.INIT('h2a)
	) name17740 (
		\m2_addr_i[30]_pad ,
		_w1908_,
		_w1909_,
		_w19641_
	);
	LUT3 #(
		.INIT('h2a)
	) name17741 (
		\m5_addr_i[30]_pad ,
		_w1901_,
		_w1902_,
		_w19642_
	);
	LUT4 #(
		.INIT('h135f)
	) name17742 (
		_w1914_,
		_w1920_,
		_w19641_,
		_w19642_,
		_w19643_
	);
	LUT3 #(
		.INIT('h80)
	) name17743 (
		\m0_addr_i[30]_pad ,
		_w1908_,
		_w1909_,
		_w19644_
	);
	LUT3 #(
		.INIT('h2a)
	) name17744 (
		\m7_addr_i[30]_pad ,
		_w1901_,
		_w1902_,
		_w19645_
	);
	LUT4 #(
		.INIT('h135f)
	) name17745 (
		_w1914_,
		_w1918_,
		_w19644_,
		_w19645_,
		_w19646_
	);
	LUT4 #(
		.INIT('h7fff)
	) name17746 (
		_w19637_,
		_w19640_,
		_w19643_,
		_w19646_,
		_w19647_
	);
	LUT3 #(
		.INIT('h80)
	) name17747 (
		\m4_addr_i[31]_pad ,
		_w1908_,
		_w1909_,
		_w19648_
	);
	LUT3 #(
		.INIT('h80)
	) name17748 (
		\m3_addr_i[31]_pad ,
		_w1901_,
		_w1902_,
		_w19649_
	);
	LUT4 #(
		.INIT('h135f)
	) name17749 (
		_w1907_,
		_w1918_,
		_w19648_,
		_w19649_,
		_w19650_
	);
	LUT3 #(
		.INIT('h80)
	) name17750 (
		\m1_addr_i[31]_pad ,
		_w1901_,
		_w1902_,
		_w19651_
	);
	LUT3 #(
		.INIT('h2a)
	) name17751 (
		\m6_addr_i[31]_pad ,
		_w1908_,
		_w1909_,
		_w19652_
	);
	LUT4 #(
		.INIT('h153f)
	) name17752 (
		_w1907_,
		_w1920_,
		_w19651_,
		_w19652_,
		_w19653_
	);
	LUT3 #(
		.INIT('h2a)
	) name17753 (
		\m2_addr_i[31]_pad ,
		_w1908_,
		_w1909_,
		_w19654_
	);
	LUT3 #(
		.INIT('h2a)
	) name17754 (
		\m5_addr_i[31]_pad ,
		_w1901_,
		_w1902_,
		_w19655_
	);
	LUT4 #(
		.INIT('h135f)
	) name17755 (
		_w1914_,
		_w1920_,
		_w19654_,
		_w19655_,
		_w19656_
	);
	LUT3 #(
		.INIT('h80)
	) name17756 (
		\m0_addr_i[31]_pad ,
		_w1908_,
		_w1909_,
		_w19657_
	);
	LUT3 #(
		.INIT('h2a)
	) name17757 (
		\m7_addr_i[31]_pad ,
		_w1901_,
		_w1902_,
		_w19658_
	);
	LUT4 #(
		.INIT('h135f)
	) name17758 (
		_w1914_,
		_w1918_,
		_w19657_,
		_w19658_,
		_w19659_
	);
	LUT4 #(
		.INIT('h7fff)
	) name17759 (
		_w19650_,
		_w19653_,
		_w19656_,
		_w19659_,
		_w19660_
	);
	LUT3 #(
		.INIT('h2a)
	) name17760 (
		\m7_addr_i[6]_pad ,
		_w1901_,
		_w1902_,
		_w19661_
	);
	LUT3 #(
		.INIT('h2a)
	) name17761 (
		\m6_addr_i[6]_pad ,
		_w1908_,
		_w1909_,
		_w19662_
	);
	LUT4 #(
		.INIT('h153f)
	) name17762 (
		_w1907_,
		_w1918_,
		_w19661_,
		_w19662_,
		_w19663_
	);
	LUT3 #(
		.INIT('h2a)
	) name17763 (
		\m5_addr_i[6]_pad ,
		_w1901_,
		_w1902_,
		_w19664_
	);
	LUT3 #(
		.INIT('h2a)
	) name17764 (
		\m2_addr_i[6]_pad ,
		_w1908_,
		_w1909_,
		_w19665_
	);
	LUT4 #(
		.INIT('h153f)
	) name17765 (
		_w1914_,
		_w1920_,
		_w19664_,
		_w19665_,
		_w19666_
	);
	LUT3 #(
		.INIT('h80)
	) name17766 (
		\m4_addr_i[6]_pad ,
		_w1908_,
		_w1909_,
		_w19667_
	);
	LUT3 #(
		.INIT('h80)
	) name17767 (
		\m3_addr_i[6]_pad ,
		_w1901_,
		_w1902_,
		_w19668_
	);
	LUT4 #(
		.INIT('h135f)
	) name17768 (
		_w1907_,
		_w1918_,
		_w19667_,
		_w19668_,
		_w19669_
	);
	LUT3 #(
		.INIT('h80)
	) name17769 (
		\m1_addr_i[6]_pad ,
		_w1901_,
		_w1902_,
		_w19670_
	);
	LUT3 #(
		.INIT('h80)
	) name17770 (
		\m0_addr_i[6]_pad ,
		_w1908_,
		_w1909_,
		_w19671_
	);
	LUT4 #(
		.INIT('h153f)
	) name17771 (
		_w1914_,
		_w1920_,
		_w19670_,
		_w19671_,
		_w19672_
	);
	LUT4 #(
		.INIT('h7fff)
	) name17772 (
		_w19663_,
		_w19666_,
		_w19669_,
		_w19672_,
		_w19673_
	);
	LUT3 #(
		.INIT('h2a)
	) name17773 (
		\m7_addr_i[7]_pad ,
		_w1901_,
		_w1902_,
		_w19674_
	);
	LUT3 #(
		.INIT('h2a)
	) name17774 (
		\m6_addr_i[7]_pad ,
		_w1908_,
		_w1909_,
		_w19675_
	);
	LUT4 #(
		.INIT('h153f)
	) name17775 (
		_w1907_,
		_w1918_,
		_w19674_,
		_w19675_,
		_w19676_
	);
	LUT3 #(
		.INIT('h2a)
	) name17776 (
		\m5_addr_i[7]_pad ,
		_w1901_,
		_w1902_,
		_w19677_
	);
	LUT3 #(
		.INIT('h2a)
	) name17777 (
		\m2_addr_i[7]_pad ,
		_w1908_,
		_w1909_,
		_w19678_
	);
	LUT4 #(
		.INIT('h153f)
	) name17778 (
		_w1914_,
		_w1920_,
		_w19677_,
		_w19678_,
		_w19679_
	);
	LUT3 #(
		.INIT('h80)
	) name17779 (
		\m4_addr_i[7]_pad ,
		_w1908_,
		_w1909_,
		_w19680_
	);
	LUT3 #(
		.INIT('h80)
	) name17780 (
		\m3_addr_i[7]_pad ,
		_w1901_,
		_w1902_,
		_w19681_
	);
	LUT4 #(
		.INIT('h135f)
	) name17781 (
		_w1907_,
		_w1918_,
		_w19680_,
		_w19681_,
		_w19682_
	);
	LUT3 #(
		.INIT('h80)
	) name17782 (
		\m1_addr_i[7]_pad ,
		_w1901_,
		_w1902_,
		_w19683_
	);
	LUT3 #(
		.INIT('h80)
	) name17783 (
		\m0_addr_i[7]_pad ,
		_w1908_,
		_w1909_,
		_w19684_
	);
	LUT4 #(
		.INIT('h153f)
	) name17784 (
		_w1914_,
		_w1920_,
		_w19683_,
		_w19684_,
		_w19685_
	);
	LUT4 #(
		.INIT('h7fff)
	) name17785 (
		_w19676_,
		_w19679_,
		_w19682_,
		_w19685_,
		_w19686_
	);
	LUT3 #(
		.INIT('h2a)
	) name17786 (
		\m7_addr_i[8]_pad ,
		_w1901_,
		_w1902_,
		_w19687_
	);
	LUT3 #(
		.INIT('h2a)
	) name17787 (
		\m6_addr_i[8]_pad ,
		_w1908_,
		_w1909_,
		_w19688_
	);
	LUT4 #(
		.INIT('h153f)
	) name17788 (
		_w1907_,
		_w1918_,
		_w19687_,
		_w19688_,
		_w19689_
	);
	LUT3 #(
		.INIT('h2a)
	) name17789 (
		\m5_addr_i[8]_pad ,
		_w1901_,
		_w1902_,
		_w19690_
	);
	LUT3 #(
		.INIT('h2a)
	) name17790 (
		\m2_addr_i[8]_pad ,
		_w1908_,
		_w1909_,
		_w19691_
	);
	LUT4 #(
		.INIT('h153f)
	) name17791 (
		_w1914_,
		_w1920_,
		_w19690_,
		_w19691_,
		_w19692_
	);
	LUT3 #(
		.INIT('h80)
	) name17792 (
		\m4_addr_i[8]_pad ,
		_w1908_,
		_w1909_,
		_w19693_
	);
	LUT3 #(
		.INIT('h80)
	) name17793 (
		\m3_addr_i[8]_pad ,
		_w1901_,
		_w1902_,
		_w19694_
	);
	LUT4 #(
		.INIT('h135f)
	) name17794 (
		_w1907_,
		_w1918_,
		_w19693_,
		_w19694_,
		_w19695_
	);
	LUT3 #(
		.INIT('h80)
	) name17795 (
		\m1_addr_i[8]_pad ,
		_w1901_,
		_w1902_,
		_w19696_
	);
	LUT3 #(
		.INIT('h80)
	) name17796 (
		\m0_addr_i[8]_pad ,
		_w1908_,
		_w1909_,
		_w19697_
	);
	LUT4 #(
		.INIT('h153f)
	) name17797 (
		_w1914_,
		_w1920_,
		_w19696_,
		_w19697_,
		_w19698_
	);
	LUT4 #(
		.INIT('h7fff)
	) name17798 (
		_w19689_,
		_w19692_,
		_w19695_,
		_w19698_,
		_w19699_
	);
	LUT3 #(
		.INIT('h80)
	) name17799 (
		\m3_addr_i[9]_pad ,
		_w1901_,
		_w1902_,
		_w19700_
	);
	LUT3 #(
		.INIT('h2a)
	) name17800 (
		\m2_addr_i[9]_pad ,
		_w1908_,
		_w1909_,
		_w19701_
	);
	LUT4 #(
		.INIT('h153f)
	) name17801 (
		_w1914_,
		_w1918_,
		_w19700_,
		_w19701_,
		_w19702_
	);
	LUT3 #(
		.INIT('h2a)
	) name17802 (
		\m5_addr_i[9]_pad ,
		_w1901_,
		_w1902_,
		_w19703_
	);
	LUT3 #(
		.INIT('h80)
	) name17803 (
		\m0_addr_i[9]_pad ,
		_w1908_,
		_w1909_,
		_w19704_
	);
	LUT4 #(
		.INIT('h153f)
	) name17804 (
		_w1914_,
		_w1920_,
		_w19703_,
		_w19704_,
		_w19705_
	);
	LUT3 #(
		.INIT('h80)
	) name17805 (
		\m4_addr_i[9]_pad ,
		_w1908_,
		_w1909_,
		_w19706_
	);
	LUT3 #(
		.INIT('h80)
	) name17806 (
		\m1_addr_i[9]_pad ,
		_w1901_,
		_w1902_,
		_w19707_
	);
	LUT4 #(
		.INIT('h135f)
	) name17807 (
		_w1907_,
		_w1920_,
		_w19706_,
		_w19707_,
		_w19708_
	);
	LUT3 #(
		.INIT('h2a)
	) name17808 (
		\m7_addr_i[9]_pad ,
		_w1901_,
		_w1902_,
		_w19709_
	);
	LUT3 #(
		.INIT('h2a)
	) name17809 (
		\m6_addr_i[9]_pad ,
		_w1908_,
		_w1909_,
		_w19710_
	);
	LUT4 #(
		.INIT('h153f)
	) name17810 (
		_w1907_,
		_w1918_,
		_w19709_,
		_w19710_,
		_w19711_
	);
	LUT4 #(
		.INIT('h7fff)
	) name17811 (
		_w19702_,
		_w19705_,
		_w19708_,
		_w19711_,
		_w19712_
	);
	LUT3 #(
		.INIT('h15)
	) name17812 (
		_w2016_,
		_w2045_,
		_w2097_,
		_w19713_
	);
	LUT3 #(
		.INIT('h2a)
	) name17813 (
		\m7_data_i[16]_pad ,
		_w1901_,
		_w1902_,
		_w19714_
	);
	LUT3 #(
		.INIT('h2a)
	) name17814 (
		\m6_data_i[16]_pad ,
		_w1908_,
		_w1909_,
		_w19715_
	);
	LUT4 #(
		.INIT('h153f)
	) name17815 (
		_w1907_,
		_w1918_,
		_w19714_,
		_w19715_,
		_w19716_
	);
	LUT3 #(
		.INIT('h2a)
	) name17816 (
		\m5_data_i[16]_pad ,
		_w1901_,
		_w1902_,
		_w19717_
	);
	LUT3 #(
		.INIT('h2a)
	) name17817 (
		\m2_data_i[16]_pad ,
		_w1908_,
		_w1909_,
		_w19718_
	);
	LUT4 #(
		.INIT('h153f)
	) name17818 (
		_w1914_,
		_w1920_,
		_w19717_,
		_w19718_,
		_w19719_
	);
	LUT3 #(
		.INIT('h80)
	) name17819 (
		\m4_data_i[16]_pad ,
		_w1908_,
		_w1909_,
		_w19720_
	);
	LUT3 #(
		.INIT('h80)
	) name17820 (
		\m3_data_i[16]_pad ,
		_w1901_,
		_w1902_,
		_w19721_
	);
	LUT4 #(
		.INIT('h135f)
	) name17821 (
		_w1907_,
		_w1918_,
		_w19720_,
		_w19721_,
		_w19722_
	);
	LUT3 #(
		.INIT('h80)
	) name17822 (
		\m1_data_i[16]_pad ,
		_w1901_,
		_w1902_,
		_w19723_
	);
	LUT3 #(
		.INIT('h80)
	) name17823 (
		\m0_data_i[16]_pad ,
		_w1908_,
		_w1909_,
		_w19724_
	);
	LUT4 #(
		.INIT('h153f)
	) name17824 (
		_w1914_,
		_w1920_,
		_w19723_,
		_w19724_,
		_w19725_
	);
	LUT4 #(
		.INIT('h7fff)
	) name17825 (
		_w19716_,
		_w19719_,
		_w19722_,
		_w19725_,
		_w19726_
	);
	LUT3 #(
		.INIT('h2a)
	) name17826 (
		\m7_data_i[17]_pad ,
		_w1901_,
		_w1902_,
		_w19727_
	);
	LUT3 #(
		.INIT('h2a)
	) name17827 (
		\m6_data_i[17]_pad ,
		_w1908_,
		_w1909_,
		_w19728_
	);
	LUT4 #(
		.INIT('h153f)
	) name17828 (
		_w1907_,
		_w1918_,
		_w19727_,
		_w19728_,
		_w19729_
	);
	LUT3 #(
		.INIT('h2a)
	) name17829 (
		\m5_data_i[17]_pad ,
		_w1901_,
		_w1902_,
		_w19730_
	);
	LUT3 #(
		.INIT('h80)
	) name17830 (
		\m0_data_i[17]_pad ,
		_w1908_,
		_w1909_,
		_w19731_
	);
	LUT4 #(
		.INIT('h153f)
	) name17831 (
		_w1914_,
		_w1920_,
		_w19730_,
		_w19731_,
		_w19732_
	);
	LUT3 #(
		.INIT('h80)
	) name17832 (
		\m4_data_i[17]_pad ,
		_w1908_,
		_w1909_,
		_w19733_
	);
	LUT3 #(
		.INIT('h80)
	) name17833 (
		\m1_data_i[17]_pad ,
		_w1901_,
		_w1902_,
		_w19734_
	);
	LUT4 #(
		.INIT('h135f)
	) name17834 (
		_w1907_,
		_w1920_,
		_w19733_,
		_w19734_,
		_w19735_
	);
	LUT3 #(
		.INIT('h80)
	) name17835 (
		\m3_data_i[17]_pad ,
		_w1901_,
		_w1902_,
		_w19736_
	);
	LUT3 #(
		.INIT('h2a)
	) name17836 (
		\m2_data_i[17]_pad ,
		_w1908_,
		_w1909_,
		_w19737_
	);
	LUT4 #(
		.INIT('h153f)
	) name17837 (
		_w1914_,
		_w1918_,
		_w19736_,
		_w19737_,
		_w19738_
	);
	LUT4 #(
		.INIT('h7fff)
	) name17838 (
		_w19729_,
		_w19732_,
		_w19735_,
		_w19738_,
		_w19739_
	);
	LUT3 #(
		.INIT('h2a)
	) name17839 (
		\m7_data_i[18]_pad ,
		_w1901_,
		_w1902_,
		_w19740_
	);
	LUT3 #(
		.INIT('h2a)
	) name17840 (
		\m6_data_i[18]_pad ,
		_w1908_,
		_w1909_,
		_w19741_
	);
	LUT4 #(
		.INIT('h153f)
	) name17841 (
		_w1907_,
		_w1918_,
		_w19740_,
		_w19741_,
		_w19742_
	);
	LUT3 #(
		.INIT('h2a)
	) name17842 (
		\m5_data_i[18]_pad ,
		_w1901_,
		_w1902_,
		_w19743_
	);
	LUT3 #(
		.INIT('h2a)
	) name17843 (
		\m2_data_i[18]_pad ,
		_w1908_,
		_w1909_,
		_w19744_
	);
	LUT4 #(
		.INIT('h153f)
	) name17844 (
		_w1914_,
		_w1920_,
		_w19743_,
		_w19744_,
		_w19745_
	);
	LUT3 #(
		.INIT('h80)
	) name17845 (
		\m4_data_i[18]_pad ,
		_w1908_,
		_w1909_,
		_w19746_
	);
	LUT3 #(
		.INIT('h80)
	) name17846 (
		\m3_data_i[18]_pad ,
		_w1901_,
		_w1902_,
		_w19747_
	);
	LUT4 #(
		.INIT('h135f)
	) name17847 (
		_w1907_,
		_w1918_,
		_w19746_,
		_w19747_,
		_w19748_
	);
	LUT3 #(
		.INIT('h80)
	) name17848 (
		\m1_data_i[18]_pad ,
		_w1901_,
		_w1902_,
		_w19749_
	);
	LUT3 #(
		.INIT('h80)
	) name17849 (
		\m0_data_i[18]_pad ,
		_w1908_,
		_w1909_,
		_w19750_
	);
	LUT4 #(
		.INIT('h153f)
	) name17850 (
		_w1914_,
		_w1920_,
		_w19749_,
		_w19750_,
		_w19751_
	);
	LUT4 #(
		.INIT('h7fff)
	) name17851 (
		_w19742_,
		_w19745_,
		_w19748_,
		_w19751_,
		_w19752_
	);
	LUT3 #(
		.INIT('h2a)
	) name17852 (
		\m5_data_i[19]_pad ,
		_w1901_,
		_w1902_,
		_w19753_
	);
	LUT3 #(
		.INIT('h80)
	) name17853 (
		\m4_data_i[19]_pad ,
		_w1908_,
		_w1909_,
		_w19754_
	);
	LUT4 #(
		.INIT('h153f)
	) name17854 (
		_w1907_,
		_w1920_,
		_w19753_,
		_w19754_,
		_w19755_
	);
	LUT3 #(
		.INIT('h2a)
	) name17855 (
		\m7_data_i[19]_pad ,
		_w1901_,
		_w1902_,
		_w19756_
	);
	LUT3 #(
		.INIT('h2a)
	) name17856 (
		\m2_data_i[19]_pad ,
		_w1908_,
		_w1909_,
		_w19757_
	);
	LUT4 #(
		.INIT('h153f)
	) name17857 (
		_w1914_,
		_w1918_,
		_w19756_,
		_w19757_,
		_w19758_
	);
	LUT3 #(
		.INIT('h2a)
	) name17858 (
		\m6_data_i[19]_pad ,
		_w1908_,
		_w1909_,
		_w19759_
	);
	LUT3 #(
		.INIT('h80)
	) name17859 (
		\m3_data_i[19]_pad ,
		_w1901_,
		_w1902_,
		_w19760_
	);
	LUT4 #(
		.INIT('h135f)
	) name17860 (
		_w1907_,
		_w1918_,
		_w19759_,
		_w19760_,
		_w19761_
	);
	LUT3 #(
		.INIT('h80)
	) name17861 (
		\m1_data_i[19]_pad ,
		_w1901_,
		_w1902_,
		_w19762_
	);
	LUT3 #(
		.INIT('h80)
	) name17862 (
		\m0_data_i[19]_pad ,
		_w1908_,
		_w1909_,
		_w19763_
	);
	LUT4 #(
		.INIT('h153f)
	) name17863 (
		_w1914_,
		_w1920_,
		_w19762_,
		_w19763_,
		_w19764_
	);
	LUT4 #(
		.INIT('h7fff)
	) name17864 (
		_w19755_,
		_w19758_,
		_w19761_,
		_w19764_,
		_w19765_
	);
	LUT3 #(
		.INIT('h2a)
	) name17865 (
		\m7_data_i[20]_pad ,
		_w1901_,
		_w1902_,
		_w19766_
	);
	LUT3 #(
		.INIT('h2a)
	) name17866 (
		\m6_data_i[20]_pad ,
		_w1908_,
		_w1909_,
		_w19767_
	);
	LUT4 #(
		.INIT('h153f)
	) name17867 (
		_w1907_,
		_w1918_,
		_w19766_,
		_w19767_,
		_w19768_
	);
	LUT3 #(
		.INIT('h2a)
	) name17868 (
		\m5_data_i[20]_pad ,
		_w1901_,
		_w1902_,
		_w19769_
	);
	LUT3 #(
		.INIT('h2a)
	) name17869 (
		\m2_data_i[20]_pad ,
		_w1908_,
		_w1909_,
		_w19770_
	);
	LUT4 #(
		.INIT('h153f)
	) name17870 (
		_w1914_,
		_w1920_,
		_w19769_,
		_w19770_,
		_w19771_
	);
	LUT3 #(
		.INIT('h80)
	) name17871 (
		\m4_data_i[20]_pad ,
		_w1908_,
		_w1909_,
		_w19772_
	);
	LUT3 #(
		.INIT('h80)
	) name17872 (
		\m3_data_i[20]_pad ,
		_w1901_,
		_w1902_,
		_w19773_
	);
	LUT4 #(
		.INIT('h135f)
	) name17873 (
		_w1907_,
		_w1918_,
		_w19772_,
		_w19773_,
		_w19774_
	);
	LUT3 #(
		.INIT('h80)
	) name17874 (
		\m1_data_i[20]_pad ,
		_w1901_,
		_w1902_,
		_w19775_
	);
	LUT3 #(
		.INIT('h80)
	) name17875 (
		\m0_data_i[20]_pad ,
		_w1908_,
		_w1909_,
		_w19776_
	);
	LUT4 #(
		.INIT('h153f)
	) name17876 (
		_w1914_,
		_w1920_,
		_w19775_,
		_w19776_,
		_w19777_
	);
	LUT4 #(
		.INIT('h7fff)
	) name17877 (
		_w19768_,
		_w19771_,
		_w19774_,
		_w19777_,
		_w19778_
	);
	LUT3 #(
		.INIT('h2a)
	) name17878 (
		\m5_data_i[21]_pad ,
		_w1901_,
		_w1902_,
		_w19779_
	);
	LUT3 #(
		.INIT('h80)
	) name17879 (
		\m4_data_i[21]_pad ,
		_w1908_,
		_w1909_,
		_w19780_
	);
	LUT4 #(
		.INIT('h153f)
	) name17880 (
		_w1907_,
		_w1920_,
		_w19779_,
		_w19780_,
		_w19781_
	);
	LUT3 #(
		.INIT('h2a)
	) name17881 (
		\m7_data_i[21]_pad ,
		_w1901_,
		_w1902_,
		_w19782_
	);
	LUT3 #(
		.INIT('h2a)
	) name17882 (
		\m2_data_i[21]_pad ,
		_w1908_,
		_w1909_,
		_w19783_
	);
	LUT4 #(
		.INIT('h153f)
	) name17883 (
		_w1914_,
		_w1918_,
		_w19782_,
		_w19783_,
		_w19784_
	);
	LUT3 #(
		.INIT('h2a)
	) name17884 (
		\m6_data_i[21]_pad ,
		_w1908_,
		_w1909_,
		_w19785_
	);
	LUT3 #(
		.INIT('h80)
	) name17885 (
		\m3_data_i[21]_pad ,
		_w1901_,
		_w1902_,
		_w19786_
	);
	LUT4 #(
		.INIT('h135f)
	) name17886 (
		_w1907_,
		_w1918_,
		_w19785_,
		_w19786_,
		_w19787_
	);
	LUT3 #(
		.INIT('h80)
	) name17887 (
		\m1_data_i[21]_pad ,
		_w1901_,
		_w1902_,
		_w19788_
	);
	LUT3 #(
		.INIT('h80)
	) name17888 (
		\m0_data_i[21]_pad ,
		_w1908_,
		_w1909_,
		_w19789_
	);
	LUT4 #(
		.INIT('h153f)
	) name17889 (
		_w1914_,
		_w1920_,
		_w19788_,
		_w19789_,
		_w19790_
	);
	LUT4 #(
		.INIT('h7fff)
	) name17890 (
		_w19781_,
		_w19784_,
		_w19787_,
		_w19790_,
		_w19791_
	);
	LUT3 #(
		.INIT('h2a)
	) name17891 (
		\m7_data_i[22]_pad ,
		_w1901_,
		_w1902_,
		_w19792_
	);
	LUT3 #(
		.INIT('h2a)
	) name17892 (
		\m6_data_i[22]_pad ,
		_w1908_,
		_w1909_,
		_w19793_
	);
	LUT4 #(
		.INIT('h153f)
	) name17893 (
		_w1907_,
		_w1918_,
		_w19792_,
		_w19793_,
		_w19794_
	);
	LUT3 #(
		.INIT('h2a)
	) name17894 (
		\m5_data_i[22]_pad ,
		_w1901_,
		_w1902_,
		_w19795_
	);
	LUT3 #(
		.INIT('h2a)
	) name17895 (
		\m2_data_i[22]_pad ,
		_w1908_,
		_w1909_,
		_w19796_
	);
	LUT4 #(
		.INIT('h153f)
	) name17896 (
		_w1914_,
		_w1920_,
		_w19795_,
		_w19796_,
		_w19797_
	);
	LUT3 #(
		.INIT('h80)
	) name17897 (
		\m4_data_i[22]_pad ,
		_w1908_,
		_w1909_,
		_w19798_
	);
	LUT3 #(
		.INIT('h80)
	) name17898 (
		\m3_data_i[22]_pad ,
		_w1901_,
		_w1902_,
		_w19799_
	);
	LUT4 #(
		.INIT('h135f)
	) name17899 (
		_w1907_,
		_w1918_,
		_w19798_,
		_w19799_,
		_w19800_
	);
	LUT3 #(
		.INIT('h80)
	) name17900 (
		\m1_data_i[22]_pad ,
		_w1901_,
		_w1902_,
		_w19801_
	);
	LUT3 #(
		.INIT('h80)
	) name17901 (
		\m0_data_i[22]_pad ,
		_w1908_,
		_w1909_,
		_w19802_
	);
	LUT4 #(
		.INIT('h153f)
	) name17902 (
		_w1914_,
		_w1920_,
		_w19801_,
		_w19802_,
		_w19803_
	);
	LUT4 #(
		.INIT('h7fff)
	) name17903 (
		_w19794_,
		_w19797_,
		_w19800_,
		_w19803_,
		_w19804_
	);
	LUT3 #(
		.INIT('h2a)
	) name17904 (
		\m7_data_i[23]_pad ,
		_w1901_,
		_w1902_,
		_w19805_
	);
	LUT3 #(
		.INIT('h2a)
	) name17905 (
		\m6_data_i[23]_pad ,
		_w1908_,
		_w1909_,
		_w19806_
	);
	LUT4 #(
		.INIT('h153f)
	) name17906 (
		_w1907_,
		_w1918_,
		_w19805_,
		_w19806_,
		_w19807_
	);
	LUT3 #(
		.INIT('h2a)
	) name17907 (
		\m5_data_i[23]_pad ,
		_w1901_,
		_w1902_,
		_w19808_
	);
	LUT3 #(
		.INIT('h2a)
	) name17908 (
		\m2_data_i[23]_pad ,
		_w1908_,
		_w1909_,
		_w19809_
	);
	LUT4 #(
		.INIT('h153f)
	) name17909 (
		_w1914_,
		_w1920_,
		_w19808_,
		_w19809_,
		_w19810_
	);
	LUT3 #(
		.INIT('h80)
	) name17910 (
		\m4_data_i[23]_pad ,
		_w1908_,
		_w1909_,
		_w19811_
	);
	LUT3 #(
		.INIT('h80)
	) name17911 (
		\m3_data_i[23]_pad ,
		_w1901_,
		_w1902_,
		_w19812_
	);
	LUT4 #(
		.INIT('h135f)
	) name17912 (
		_w1907_,
		_w1918_,
		_w19811_,
		_w19812_,
		_w19813_
	);
	LUT3 #(
		.INIT('h80)
	) name17913 (
		\m1_data_i[23]_pad ,
		_w1901_,
		_w1902_,
		_w19814_
	);
	LUT3 #(
		.INIT('h80)
	) name17914 (
		\m0_data_i[23]_pad ,
		_w1908_,
		_w1909_,
		_w19815_
	);
	LUT4 #(
		.INIT('h153f)
	) name17915 (
		_w1914_,
		_w1920_,
		_w19814_,
		_w19815_,
		_w19816_
	);
	LUT4 #(
		.INIT('h7fff)
	) name17916 (
		_w19807_,
		_w19810_,
		_w19813_,
		_w19816_,
		_w19817_
	);
	LUT3 #(
		.INIT('h2a)
	) name17917 (
		\m7_data_i[24]_pad ,
		_w1901_,
		_w1902_,
		_w19818_
	);
	LUT3 #(
		.INIT('h2a)
	) name17918 (
		\m6_data_i[24]_pad ,
		_w1908_,
		_w1909_,
		_w19819_
	);
	LUT4 #(
		.INIT('h153f)
	) name17919 (
		_w1907_,
		_w1918_,
		_w19818_,
		_w19819_,
		_w19820_
	);
	LUT3 #(
		.INIT('h2a)
	) name17920 (
		\m5_data_i[24]_pad ,
		_w1901_,
		_w1902_,
		_w19821_
	);
	LUT3 #(
		.INIT('h2a)
	) name17921 (
		\m2_data_i[24]_pad ,
		_w1908_,
		_w1909_,
		_w19822_
	);
	LUT4 #(
		.INIT('h153f)
	) name17922 (
		_w1914_,
		_w1920_,
		_w19821_,
		_w19822_,
		_w19823_
	);
	LUT3 #(
		.INIT('h80)
	) name17923 (
		\m4_data_i[24]_pad ,
		_w1908_,
		_w1909_,
		_w19824_
	);
	LUT3 #(
		.INIT('h80)
	) name17924 (
		\m3_data_i[24]_pad ,
		_w1901_,
		_w1902_,
		_w19825_
	);
	LUT4 #(
		.INIT('h135f)
	) name17925 (
		_w1907_,
		_w1918_,
		_w19824_,
		_w19825_,
		_w19826_
	);
	LUT3 #(
		.INIT('h80)
	) name17926 (
		\m1_data_i[24]_pad ,
		_w1901_,
		_w1902_,
		_w19827_
	);
	LUT3 #(
		.INIT('h80)
	) name17927 (
		\m0_data_i[24]_pad ,
		_w1908_,
		_w1909_,
		_w19828_
	);
	LUT4 #(
		.INIT('h153f)
	) name17928 (
		_w1914_,
		_w1920_,
		_w19827_,
		_w19828_,
		_w19829_
	);
	LUT4 #(
		.INIT('h7fff)
	) name17929 (
		_w19820_,
		_w19823_,
		_w19826_,
		_w19829_,
		_w19830_
	);
	LUT3 #(
		.INIT('h2a)
	) name17930 (
		\m7_data_i[25]_pad ,
		_w1901_,
		_w1902_,
		_w19831_
	);
	LUT3 #(
		.INIT('h2a)
	) name17931 (
		\m6_data_i[25]_pad ,
		_w1908_,
		_w1909_,
		_w19832_
	);
	LUT4 #(
		.INIT('h153f)
	) name17932 (
		_w1907_,
		_w1918_,
		_w19831_,
		_w19832_,
		_w19833_
	);
	LUT3 #(
		.INIT('h2a)
	) name17933 (
		\m5_data_i[25]_pad ,
		_w1901_,
		_w1902_,
		_w19834_
	);
	LUT3 #(
		.INIT('h2a)
	) name17934 (
		\m2_data_i[25]_pad ,
		_w1908_,
		_w1909_,
		_w19835_
	);
	LUT4 #(
		.INIT('h153f)
	) name17935 (
		_w1914_,
		_w1920_,
		_w19834_,
		_w19835_,
		_w19836_
	);
	LUT3 #(
		.INIT('h80)
	) name17936 (
		\m4_data_i[25]_pad ,
		_w1908_,
		_w1909_,
		_w19837_
	);
	LUT3 #(
		.INIT('h80)
	) name17937 (
		\m3_data_i[25]_pad ,
		_w1901_,
		_w1902_,
		_w19838_
	);
	LUT4 #(
		.INIT('h135f)
	) name17938 (
		_w1907_,
		_w1918_,
		_w19837_,
		_w19838_,
		_w19839_
	);
	LUT3 #(
		.INIT('h80)
	) name17939 (
		\m1_data_i[25]_pad ,
		_w1901_,
		_w1902_,
		_w19840_
	);
	LUT3 #(
		.INIT('h80)
	) name17940 (
		\m0_data_i[25]_pad ,
		_w1908_,
		_w1909_,
		_w19841_
	);
	LUT4 #(
		.INIT('h153f)
	) name17941 (
		_w1914_,
		_w1920_,
		_w19840_,
		_w19841_,
		_w19842_
	);
	LUT4 #(
		.INIT('h7fff)
	) name17942 (
		_w19833_,
		_w19836_,
		_w19839_,
		_w19842_,
		_w19843_
	);
	LUT3 #(
		.INIT('h2a)
	) name17943 (
		\m7_data_i[26]_pad ,
		_w1901_,
		_w1902_,
		_w19844_
	);
	LUT3 #(
		.INIT('h2a)
	) name17944 (
		\m6_data_i[26]_pad ,
		_w1908_,
		_w1909_,
		_w19845_
	);
	LUT4 #(
		.INIT('h153f)
	) name17945 (
		_w1907_,
		_w1918_,
		_w19844_,
		_w19845_,
		_w19846_
	);
	LUT3 #(
		.INIT('h2a)
	) name17946 (
		\m5_data_i[26]_pad ,
		_w1901_,
		_w1902_,
		_w19847_
	);
	LUT3 #(
		.INIT('h2a)
	) name17947 (
		\m2_data_i[26]_pad ,
		_w1908_,
		_w1909_,
		_w19848_
	);
	LUT4 #(
		.INIT('h153f)
	) name17948 (
		_w1914_,
		_w1920_,
		_w19847_,
		_w19848_,
		_w19849_
	);
	LUT3 #(
		.INIT('h80)
	) name17949 (
		\m4_data_i[26]_pad ,
		_w1908_,
		_w1909_,
		_w19850_
	);
	LUT3 #(
		.INIT('h80)
	) name17950 (
		\m3_data_i[26]_pad ,
		_w1901_,
		_w1902_,
		_w19851_
	);
	LUT4 #(
		.INIT('h135f)
	) name17951 (
		_w1907_,
		_w1918_,
		_w19850_,
		_w19851_,
		_w19852_
	);
	LUT3 #(
		.INIT('h80)
	) name17952 (
		\m1_data_i[26]_pad ,
		_w1901_,
		_w1902_,
		_w19853_
	);
	LUT3 #(
		.INIT('h80)
	) name17953 (
		\m0_data_i[26]_pad ,
		_w1908_,
		_w1909_,
		_w19854_
	);
	LUT4 #(
		.INIT('h153f)
	) name17954 (
		_w1914_,
		_w1920_,
		_w19853_,
		_w19854_,
		_w19855_
	);
	LUT4 #(
		.INIT('h7fff)
	) name17955 (
		_w19846_,
		_w19849_,
		_w19852_,
		_w19855_,
		_w19856_
	);
	LUT3 #(
		.INIT('h2a)
	) name17956 (
		\m7_data_i[27]_pad ,
		_w1901_,
		_w1902_,
		_w19857_
	);
	LUT3 #(
		.INIT('h2a)
	) name17957 (
		\m6_data_i[27]_pad ,
		_w1908_,
		_w1909_,
		_w19858_
	);
	LUT4 #(
		.INIT('h153f)
	) name17958 (
		_w1907_,
		_w1918_,
		_w19857_,
		_w19858_,
		_w19859_
	);
	LUT3 #(
		.INIT('h2a)
	) name17959 (
		\m5_data_i[27]_pad ,
		_w1901_,
		_w1902_,
		_w19860_
	);
	LUT3 #(
		.INIT('h2a)
	) name17960 (
		\m2_data_i[27]_pad ,
		_w1908_,
		_w1909_,
		_w19861_
	);
	LUT4 #(
		.INIT('h153f)
	) name17961 (
		_w1914_,
		_w1920_,
		_w19860_,
		_w19861_,
		_w19862_
	);
	LUT3 #(
		.INIT('h80)
	) name17962 (
		\m4_data_i[27]_pad ,
		_w1908_,
		_w1909_,
		_w19863_
	);
	LUT3 #(
		.INIT('h80)
	) name17963 (
		\m3_data_i[27]_pad ,
		_w1901_,
		_w1902_,
		_w19864_
	);
	LUT4 #(
		.INIT('h135f)
	) name17964 (
		_w1907_,
		_w1918_,
		_w19863_,
		_w19864_,
		_w19865_
	);
	LUT3 #(
		.INIT('h80)
	) name17965 (
		\m1_data_i[27]_pad ,
		_w1901_,
		_w1902_,
		_w19866_
	);
	LUT3 #(
		.INIT('h80)
	) name17966 (
		\m0_data_i[27]_pad ,
		_w1908_,
		_w1909_,
		_w19867_
	);
	LUT4 #(
		.INIT('h153f)
	) name17967 (
		_w1914_,
		_w1920_,
		_w19866_,
		_w19867_,
		_w19868_
	);
	LUT4 #(
		.INIT('h7fff)
	) name17968 (
		_w19859_,
		_w19862_,
		_w19865_,
		_w19868_,
		_w19869_
	);
	LUT3 #(
		.INIT('h2a)
	) name17969 (
		\m7_data_i[28]_pad ,
		_w1901_,
		_w1902_,
		_w19870_
	);
	LUT3 #(
		.INIT('h2a)
	) name17970 (
		\m6_data_i[28]_pad ,
		_w1908_,
		_w1909_,
		_w19871_
	);
	LUT4 #(
		.INIT('h153f)
	) name17971 (
		_w1907_,
		_w1918_,
		_w19870_,
		_w19871_,
		_w19872_
	);
	LUT3 #(
		.INIT('h2a)
	) name17972 (
		\m5_data_i[28]_pad ,
		_w1901_,
		_w1902_,
		_w19873_
	);
	LUT3 #(
		.INIT('h2a)
	) name17973 (
		\m2_data_i[28]_pad ,
		_w1908_,
		_w1909_,
		_w19874_
	);
	LUT4 #(
		.INIT('h153f)
	) name17974 (
		_w1914_,
		_w1920_,
		_w19873_,
		_w19874_,
		_w19875_
	);
	LUT3 #(
		.INIT('h80)
	) name17975 (
		\m4_data_i[28]_pad ,
		_w1908_,
		_w1909_,
		_w19876_
	);
	LUT3 #(
		.INIT('h80)
	) name17976 (
		\m3_data_i[28]_pad ,
		_w1901_,
		_w1902_,
		_w19877_
	);
	LUT4 #(
		.INIT('h135f)
	) name17977 (
		_w1907_,
		_w1918_,
		_w19876_,
		_w19877_,
		_w19878_
	);
	LUT3 #(
		.INIT('h80)
	) name17978 (
		\m1_data_i[28]_pad ,
		_w1901_,
		_w1902_,
		_w19879_
	);
	LUT3 #(
		.INIT('h80)
	) name17979 (
		\m0_data_i[28]_pad ,
		_w1908_,
		_w1909_,
		_w19880_
	);
	LUT4 #(
		.INIT('h153f)
	) name17980 (
		_w1914_,
		_w1920_,
		_w19879_,
		_w19880_,
		_w19881_
	);
	LUT4 #(
		.INIT('h7fff)
	) name17981 (
		_w19872_,
		_w19875_,
		_w19878_,
		_w19881_,
		_w19882_
	);
	LUT3 #(
		.INIT('h2a)
	) name17982 (
		\m5_data_i[29]_pad ,
		_w1901_,
		_w1902_,
		_w19883_
	);
	LUT3 #(
		.INIT('h80)
	) name17983 (
		\m4_data_i[29]_pad ,
		_w1908_,
		_w1909_,
		_w19884_
	);
	LUT4 #(
		.INIT('h153f)
	) name17984 (
		_w1907_,
		_w1920_,
		_w19883_,
		_w19884_,
		_w19885_
	);
	LUT3 #(
		.INIT('h80)
	) name17985 (
		\m3_data_i[29]_pad ,
		_w1901_,
		_w1902_,
		_w19886_
	);
	LUT3 #(
		.INIT('h80)
	) name17986 (
		\m0_data_i[29]_pad ,
		_w1908_,
		_w1909_,
		_w19887_
	);
	LUT4 #(
		.INIT('h153f)
	) name17987 (
		_w1914_,
		_w1918_,
		_w19886_,
		_w19887_,
		_w19888_
	);
	LUT3 #(
		.INIT('h2a)
	) name17988 (
		\m2_data_i[29]_pad ,
		_w1908_,
		_w1909_,
		_w19889_
	);
	LUT3 #(
		.INIT('h80)
	) name17989 (
		\m1_data_i[29]_pad ,
		_w1901_,
		_w1902_,
		_w19890_
	);
	LUT4 #(
		.INIT('h135f)
	) name17990 (
		_w1914_,
		_w1920_,
		_w19889_,
		_w19890_,
		_w19891_
	);
	LUT3 #(
		.INIT('h2a)
	) name17991 (
		\m7_data_i[29]_pad ,
		_w1901_,
		_w1902_,
		_w19892_
	);
	LUT3 #(
		.INIT('h2a)
	) name17992 (
		\m6_data_i[29]_pad ,
		_w1908_,
		_w1909_,
		_w19893_
	);
	LUT4 #(
		.INIT('h153f)
	) name17993 (
		_w1907_,
		_w1918_,
		_w19892_,
		_w19893_,
		_w19894_
	);
	LUT4 #(
		.INIT('h7fff)
	) name17994 (
		_w19885_,
		_w19888_,
		_w19891_,
		_w19894_,
		_w19895_
	);
	LUT3 #(
		.INIT('h80)
	) name17995 (
		\m3_data_i[30]_pad ,
		_w1901_,
		_w1902_,
		_w19896_
	);
	LUT3 #(
		.INIT('h2a)
	) name17996 (
		\m2_data_i[30]_pad ,
		_w1908_,
		_w1909_,
		_w19897_
	);
	LUT4 #(
		.INIT('h153f)
	) name17997 (
		_w1914_,
		_w1918_,
		_w19896_,
		_w19897_,
		_w19898_
	);
	LUT3 #(
		.INIT('h2a)
	) name17998 (
		\m5_data_i[30]_pad ,
		_w1901_,
		_w1902_,
		_w19899_
	);
	LUT3 #(
		.INIT('h2a)
	) name17999 (
		\m6_data_i[30]_pad ,
		_w1908_,
		_w1909_,
		_w19900_
	);
	LUT4 #(
		.INIT('h153f)
	) name18000 (
		_w1907_,
		_w1920_,
		_w19899_,
		_w19900_,
		_w19901_
	);
	LUT3 #(
		.INIT('h80)
	) name18001 (
		\m4_data_i[30]_pad ,
		_w1908_,
		_w1909_,
		_w19902_
	);
	LUT3 #(
		.INIT('h2a)
	) name18002 (
		\m7_data_i[30]_pad ,
		_w1901_,
		_w1902_,
		_w19903_
	);
	LUT4 #(
		.INIT('h135f)
	) name18003 (
		_w1907_,
		_w1918_,
		_w19902_,
		_w19903_,
		_w19904_
	);
	LUT3 #(
		.INIT('h80)
	) name18004 (
		\m1_data_i[30]_pad ,
		_w1901_,
		_w1902_,
		_w19905_
	);
	LUT3 #(
		.INIT('h80)
	) name18005 (
		\m0_data_i[30]_pad ,
		_w1908_,
		_w1909_,
		_w19906_
	);
	LUT4 #(
		.INIT('h153f)
	) name18006 (
		_w1914_,
		_w1920_,
		_w19905_,
		_w19906_,
		_w19907_
	);
	LUT4 #(
		.INIT('h7fff)
	) name18007 (
		_w19898_,
		_w19901_,
		_w19904_,
		_w19907_,
		_w19908_
	);
	LUT3 #(
		.INIT('h2a)
	) name18008 (
		\m7_data_i[31]_pad ,
		_w1901_,
		_w1902_,
		_w19909_
	);
	LUT3 #(
		.INIT('h2a)
	) name18009 (
		\m6_data_i[31]_pad ,
		_w1908_,
		_w1909_,
		_w19910_
	);
	LUT4 #(
		.INIT('h153f)
	) name18010 (
		_w1907_,
		_w1918_,
		_w19909_,
		_w19910_,
		_w19911_
	);
	LUT3 #(
		.INIT('h2a)
	) name18011 (
		\m5_data_i[31]_pad ,
		_w1901_,
		_w1902_,
		_w19912_
	);
	LUT3 #(
		.INIT('h2a)
	) name18012 (
		\m2_data_i[31]_pad ,
		_w1908_,
		_w1909_,
		_w19913_
	);
	LUT4 #(
		.INIT('h153f)
	) name18013 (
		_w1914_,
		_w1920_,
		_w19912_,
		_w19913_,
		_w19914_
	);
	LUT3 #(
		.INIT('h80)
	) name18014 (
		\m4_data_i[31]_pad ,
		_w1908_,
		_w1909_,
		_w19915_
	);
	LUT3 #(
		.INIT('h80)
	) name18015 (
		\m3_data_i[31]_pad ,
		_w1901_,
		_w1902_,
		_w19916_
	);
	LUT4 #(
		.INIT('h135f)
	) name18016 (
		_w1907_,
		_w1918_,
		_w19915_,
		_w19916_,
		_w19917_
	);
	LUT3 #(
		.INIT('h80)
	) name18017 (
		\m1_data_i[31]_pad ,
		_w1901_,
		_w1902_,
		_w19918_
	);
	LUT3 #(
		.INIT('h80)
	) name18018 (
		\m0_data_i[31]_pad ,
		_w1908_,
		_w1909_,
		_w19919_
	);
	LUT4 #(
		.INIT('h153f)
	) name18019 (
		_w1914_,
		_w1920_,
		_w19918_,
		_w19919_,
		_w19920_
	);
	LUT4 #(
		.INIT('h7fff)
	) name18020 (
		_w19911_,
		_w19914_,
		_w19917_,
		_w19920_,
		_w19921_
	);
	LUT3 #(
		.INIT('h2a)
	) name18021 (
		\m7_sel_i[0]_pad ,
		_w1901_,
		_w1902_,
		_w19922_
	);
	LUT3 #(
		.INIT('h2a)
	) name18022 (
		\m6_sel_i[0]_pad ,
		_w1908_,
		_w1909_,
		_w19923_
	);
	LUT4 #(
		.INIT('h153f)
	) name18023 (
		_w1907_,
		_w1918_,
		_w19922_,
		_w19923_,
		_w19924_
	);
	LUT3 #(
		.INIT('h2a)
	) name18024 (
		\m5_sel_i[0]_pad ,
		_w1901_,
		_w1902_,
		_w19925_
	);
	LUT3 #(
		.INIT('h2a)
	) name18025 (
		\m2_sel_i[0]_pad ,
		_w1908_,
		_w1909_,
		_w19926_
	);
	LUT4 #(
		.INIT('h153f)
	) name18026 (
		_w1914_,
		_w1920_,
		_w19925_,
		_w19926_,
		_w19927_
	);
	LUT3 #(
		.INIT('h80)
	) name18027 (
		\m4_sel_i[0]_pad ,
		_w1908_,
		_w1909_,
		_w19928_
	);
	LUT3 #(
		.INIT('h80)
	) name18028 (
		\m3_sel_i[0]_pad ,
		_w1901_,
		_w1902_,
		_w19929_
	);
	LUT4 #(
		.INIT('h135f)
	) name18029 (
		_w1907_,
		_w1918_,
		_w19928_,
		_w19929_,
		_w19930_
	);
	LUT3 #(
		.INIT('h80)
	) name18030 (
		\m1_sel_i[0]_pad ,
		_w1901_,
		_w1902_,
		_w19931_
	);
	LUT3 #(
		.INIT('h80)
	) name18031 (
		\m0_sel_i[0]_pad ,
		_w1908_,
		_w1909_,
		_w19932_
	);
	LUT4 #(
		.INIT('h153f)
	) name18032 (
		_w1914_,
		_w1920_,
		_w19931_,
		_w19932_,
		_w19933_
	);
	LUT4 #(
		.INIT('h7fff)
	) name18033 (
		_w19924_,
		_w19927_,
		_w19930_,
		_w19933_,
		_w19934_
	);
	LUT3 #(
		.INIT('h2a)
	) name18034 (
		\m7_sel_i[1]_pad ,
		_w1901_,
		_w1902_,
		_w19935_
	);
	LUT3 #(
		.INIT('h2a)
	) name18035 (
		\m6_sel_i[1]_pad ,
		_w1908_,
		_w1909_,
		_w19936_
	);
	LUT4 #(
		.INIT('h153f)
	) name18036 (
		_w1907_,
		_w1918_,
		_w19935_,
		_w19936_,
		_w19937_
	);
	LUT3 #(
		.INIT('h2a)
	) name18037 (
		\m5_sel_i[1]_pad ,
		_w1901_,
		_w1902_,
		_w19938_
	);
	LUT3 #(
		.INIT('h2a)
	) name18038 (
		\m2_sel_i[1]_pad ,
		_w1908_,
		_w1909_,
		_w19939_
	);
	LUT4 #(
		.INIT('h153f)
	) name18039 (
		_w1914_,
		_w1920_,
		_w19938_,
		_w19939_,
		_w19940_
	);
	LUT3 #(
		.INIT('h80)
	) name18040 (
		\m4_sel_i[1]_pad ,
		_w1908_,
		_w1909_,
		_w19941_
	);
	LUT3 #(
		.INIT('h80)
	) name18041 (
		\m3_sel_i[1]_pad ,
		_w1901_,
		_w1902_,
		_w19942_
	);
	LUT4 #(
		.INIT('h135f)
	) name18042 (
		_w1907_,
		_w1918_,
		_w19941_,
		_w19942_,
		_w19943_
	);
	LUT3 #(
		.INIT('h80)
	) name18043 (
		\m1_sel_i[1]_pad ,
		_w1901_,
		_w1902_,
		_w19944_
	);
	LUT3 #(
		.INIT('h80)
	) name18044 (
		\m0_sel_i[1]_pad ,
		_w1908_,
		_w1909_,
		_w19945_
	);
	LUT4 #(
		.INIT('h153f)
	) name18045 (
		_w1914_,
		_w1920_,
		_w19944_,
		_w19945_,
		_w19946_
	);
	LUT4 #(
		.INIT('h7fff)
	) name18046 (
		_w19937_,
		_w19940_,
		_w19943_,
		_w19946_,
		_w19947_
	);
	LUT3 #(
		.INIT('h2a)
	) name18047 (
		\m7_sel_i[2]_pad ,
		_w1901_,
		_w1902_,
		_w19948_
	);
	LUT3 #(
		.INIT('h2a)
	) name18048 (
		\m6_sel_i[2]_pad ,
		_w1908_,
		_w1909_,
		_w19949_
	);
	LUT4 #(
		.INIT('h153f)
	) name18049 (
		_w1907_,
		_w1918_,
		_w19948_,
		_w19949_,
		_w19950_
	);
	LUT3 #(
		.INIT('h2a)
	) name18050 (
		\m5_sel_i[2]_pad ,
		_w1901_,
		_w1902_,
		_w19951_
	);
	LUT3 #(
		.INIT('h2a)
	) name18051 (
		\m2_sel_i[2]_pad ,
		_w1908_,
		_w1909_,
		_w19952_
	);
	LUT4 #(
		.INIT('h153f)
	) name18052 (
		_w1914_,
		_w1920_,
		_w19951_,
		_w19952_,
		_w19953_
	);
	LUT3 #(
		.INIT('h80)
	) name18053 (
		\m4_sel_i[2]_pad ,
		_w1908_,
		_w1909_,
		_w19954_
	);
	LUT3 #(
		.INIT('h80)
	) name18054 (
		\m3_sel_i[2]_pad ,
		_w1901_,
		_w1902_,
		_w19955_
	);
	LUT4 #(
		.INIT('h135f)
	) name18055 (
		_w1907_,
		_w1918_,
		_w19954_,
		_w19955_,
		_w19956_
	);
	LUT3 #(
		.INIT('h80)
	) name18056 (
		\m1_sel_i[2]_pad ,
		_w1901_,
		_w1902_,
		_w19957_
	);
	LUT3 #(
		.INIT('h80)
	) name18057 (
		\m0_sel_i[2]_pad ,
		_w1908_,
		_w1909_,
		_w19958_
	);
	LUT4 #(
		.INIT('h153f)
	) name18058 (
		_w1914_,
		_w1920_,
		_w19957_,
		_w19958_,
		_w19959_
	);
	LUT4 #(
		.INIT('h7fff)
	) name18059 (
		_w19950_,
		_w19953_,
		_w19956_,
		_w19959_,
		_w19960_
	);
	LUT3 #(
		.INIT('h80)
	) name18060 (
		\m3_sel_i[3]_pad ,
		_w1901_,
		_w1902_,
		_w19961_
	);
	LUT3 #(
		.INIT('h2a)
	) name18061 (
		\m2_sel_i[3]_pad ,
		_w1908_,
		_w1909_,
		_w19962_
	);
	LUT4 #(
		.INIT('h153f)
	) name18062 (
		_w1914_,
		_w1918_,
		_w19961_,
		_w19962_,
		_w19963_
	);
	LUT3 #(
		.INIT('h2a)
	) name18063 (
		\m5_sel_i[3]_pad ,
		_w1901_,
		_w1902_,
		_w19964_
	);
	LUT3 #(
		.INIT('h80)
	) name18064 (
		\m0_sel_i[3]_pad ,
		_w1908_,
		_w1909_,
		_w19965_
	);
	LUT4 #(
		.INIT('h153f)
	) name18065 (
		_w1914_,
		_w1920_,
		_w19964_,
		_w19965_,
		_w19966_
	);
	LUT3 #(
		.INIT('h80)
	) name18066 (
		\m4_sel_i[3]_pad ,
		_w1908_,
		_w1909_,
		_w19967_
	);
	LUT3 #(
		.INIT('h80)
	) name18067 (
		\m1_sel_i[3]_pad ,
		_w1901_,
		_w1902_,
		_w19968_
	);
	LUT4 #(
		.INIT('h135f)
	) name18068 (
		_w1907_,
		_w1920_,
		_w19967_,
		_w19968_,
		_w19969_
	);
	LUT3 #(
		.INIT('h2a)
	) name18069 (
		\m7_sel_i[3]_pad ,
		_w1901_,
		_w1902_,
		_w19970_
	);
	LUT3 #(
		.INIT('h2a)
	) name18070 (
		\m6_sel_i[3]_pad ,
		_w1908_,
		_w1909_,
		_w19971_
	);
	LUT4 #(
		.INIT('h153f)
	) name18071 (
		_w1907_,
		_w1918_,
		_w19970_,
		_w19971_,
		_w19972_
	);
	LUT4 #(
		.INIT('h7fff)
	) name18072 (
		_w19963_,
		_w19966_,
		_w19969_,
		_w19972_,
		_w19973_
	);
	LUT3 #(
		.INIT('h2a)
	) name18073 (
		\m3_addr_i[0]_pad ,
		_w9103_,
		_w9104_,
		_w19974_
	);
	LUT3 #(
		.INIT('h80)
	) name18074 (
		\m4_addr_i[0]_pad ,
		_w9103_,
		_w9104_,
		_w19975_
	);
	LUT4 #(
		.INIT('h9dbf)
	) name18075 (
		_w9098_,
		_w9101_,
		_w19974_,
		_w19975_,
		_w19976_
	);
	LUT3 #(
		.INIT('h80)
	) name18076 (
		\m6_addr_i[0]_pad ,
		_w9103_,
		_w9104_,
		_w19977_
	);
	LUT3 #(
		.INIT('h80)
	) name18077 (
		\m2_addr_i[0]_pad ,
		_w9103_,
		_w9104_,
		_w19978_
	);
	LUT4 #(
		.INIT('habef)
	) name18078 (
		_w9098_,
		_w9101_,
		_w19977_,
		_w19978_,
		_w19979_
	);
	LUT3 #(
		.INIT('h2a)
	) name18079 (
		\m5_addr_i[0]_pad ,
		_w9103_,
		_w9104_,
		_w19980_
	);
	LUT3 #(
		.INIT('h2a)
	) name18080 (
		\m1_addr_i[0]_pad ,
		_w9103_,
		_w9104_,
		_w19981_
	);
	LUT4 #(
		.INIT('h57df)
	) name18081 (
		_w9098_,
		_w9101_,
		_w19980_,
		_w19981_,
		_w19982_
	);
	LUT3 #(
		.INIT('h80)
	) name18082 (
		\m0_addr_i[0]_pad ,
		_w9103_,
		_w9104_,
		_w19983_
	);
	LUT3 #(
		.INIT('h2a)
	) name18083 (
		\m7_addr_i[0]_pad ,
		_w9103_,
		_w9104_,
		_w19984_
	);
	LUT4 #(
		.INIT('h6e7f)
	) name18084 (
		_w9098_,
		_w9101_,
		_w19983_,
		_w19984_,
		_w19985_
	);
	LUT4 #(
		.INIT('h7fff)
	) name18085 (
		_w19976_,
		_w19979_,
		_w19982_,
		_w19985_,
		_w19986_
	);
	LUT3 #(
		.INIT('h2a)
	) name18086 (
		\m3_addr_i[10]_pad ,
		_w9103_,
		_w9104_,
		_w19987_
	);
	LUT3 #(
		.INIT('h80)
	) name18087 (
		\m4_addr_i[10]_pad ,
		_w9103_,
		_w9104_,
		_w19988_
	);
	LUT4 #(
		.INIT('h9dbf)
	) name18088 (
		_w9098_,
		_w9101_,
		_w19987_,
		_w19988_,
		_w19989_
	);
	LUT3 #(
		.INIT('h80)
	) name18089 (
		\m6_addr_i[10]_pad ,
		_w9103_,
		_w9104_,
		_w19990_
	);
	LUT3 #(
		.INIT('h80)
	) name18090 (
		\m2_addr_i[10]_pad ,
		_w9103_,
		_w9104_,
		_w19991_
	);
	LUT4 #(
		.INIT('habef)
	) name18091 (
		_w9098_,
		_w9101_,
		_w19990_,
		_w19991_,
		_w19992_
	);
	LUT3 #(
		.INIT('h2a)
	) name18092 (
		\m5_addr_i[10]_pad ,
		_w9103_,
		_w9104_,
		_w19993_
	);
	LUT3 #(
		.INIT('h2a)
	) name18093 (
		\m1_addr_i[10]_pad ,
		_w9103_,
		_w9104_,
		_w19994_
	);
	LUT4 #(
		.INIT('h57df)
	) name18094 (
		_w9098_,
		_w9101_,
		_w19993_,
		_w19994_,
		_w19995_
	);
	LUT3 #(
		.INIT('h80)
	) name18095 (
		\m0_addr_i[10]_pad ,
		_w9103_,
		_w9104_,
		_w19996_
	);
	LUT3 #(
		.INIT('h2a)
	) name18096 (
		\m7_addr_i[10]_pad ,
		_w9103_,
		_w9104_,
		_w19997_
	);
	LUT4 #(
		.INIT('h6e7f)
	) name18097 (
		_w9098_,
		_w9101_,
		_w19996_,
		_w19997_,
		_w19998_
	);
	LUT4 #(
		.INIT('h7fff)
	) name18098 (
		_w19989_,
		_w19992_,
		_w19995_,
		_w19998_,
		_w19999_
	);
	LUT3 #(
		.INIT('h80)
	) name18099 (
		\m0_addr_i[11]_pad ,
		_w9103_,
		_w9104_,
		_w20000_
	);
	LUT3 #(
		.INIT('h2a)
	) name18100 (
		\m7_addr_i[11]_pad ,
		_w9103_,
		_w9104_,
		_w20001_
	);
	LUT4 #(
		.INIT('h6e7f)
	) name18101 (
		_w9098_,
		_w9101_,
		_w20000_,
		_w20001_,
		_w20002_
	);
	LUT3 #(
		.INIT('h80)
	) name18102 (
		\m6_addr_i[11]_pad ,
		_w9103_,
		_w9104_,
		_w20003_
	);
	LUT3 #(
		.INIT('h80)
	) name18103 (
		\m2_addr_i[11]_pad ,
		_w9103_,
		_w9104_,
		_w20004_
	);
	LUT4 #(
		.INIT('habef)
	) name18104 (
		_w9098_,
		_w9101_,
		_w20003_,
		_w20004_,
		_w20005_
	);
	LUT3 #(
		.INIT('h2a)
	) name18105 (
		\m5_addr_i[11]_pad ,
		_w9103_,
		_w9104_,
		_w20006_
	);
	LUT3 #(
		.INIT('h2a)
	) name18106 (
		\m1_addr_i[11]_pad ,
		_w9103_,
		_w9104_,
		_w20007_
	);
	LUT4 #(
		.INIT('h57df)
	) name18107 (
		_w9098_,
		_w9101_,
		_w20006_,
		_w20007_,
		_w20008_
	);
	LUT3 #(
		.INIT('h2a)
	) name18108 (
		\m3_addr_i[11]_pad ,
		_w9103_,
		_w9104_,
		_w20009_
	);
	LUT3 #(
		.INIT('h80)
	) name18109 (
		\m4_addr_i[11]_pad ,
		_w9103_,
		_w9104_,
		_w20010_
	);
	LUT4 #(
		.INIT('h9dbf)
	) name18110 (
		_w9098_,
		_w9101_,
		_w20009_,
		_w20010_,
		_w20011_
	);
	LUT4 #(
		.INIT('h7fff)
	) name18111 (
		_w20002_,
		_w20005_,
		_w20008_,
		_w20011_,
		_w20012_
	);
	LUT3 #(
		.INIT('h2a)
	) name18112 (
		\m1_addr_i[12]_pad ,
		_w9103_,
		_w9104_,
		_w20013_
	);
	LUT3 #(
		.INIT('h80)
	) name18113 (
		\m2_addr_i[12]_pad ,
		_w9103_,
		_w9104_,
		_w20014_
	);
	LUT4 #(
		.INIT('h3b7f)
	) name18114 (
		_w9098_,
		_w9101_,
		_w20013_,
		_w20014_,
		_w20015_
	);
	LUT3 #(
		.INIT('h80)
	) name18115 (
		\m0_addr_i[12]_pad ,
		_w9103_,
		_w9104_,
		_w20016_
	);
	LUT3 #(
		.INIT('h80)
	) name18116 (
		\m4_addr_i[12]_pad ,
		_w9103_,
		_w9104_,
		_w20017_
	);
	LUT4 #(
		.INIT('h5d7f)
	) name18117 (
		_w9098_,
		_w9101_,
		_w20016_,
		_w20017_,
		_w20018_
	);
	LUT3 #(
		.INIT('h2a)
	) name18118 (
		\m7_addr_i[12]_pad ,
		_w9103_,
		_w9104_,
		_w20019_
	);
	LUT3 #(
		.INIT('h2a)
	) name18119 (
		\m3_addr_i[12]_pad ,
		_w9103_,
		_w9104_,
		_w20020_
	);
	LUT4 #(
		.INIT('habef)
	) name18120 (
		_w9098_,
		_w9101_,
		_w20019_,
		_w20020_,
		_w20021_
	);
	LUT3 #(
		.INIT('h80)
	) name18121 (
		\m6_addr_i[12]_pad ,
		_w9103_,
		_w9104_,
		_w20022_
	);
	LUT3 #(
		.INIT('h2a)
	) name18122 (
		\m5_addr_i[12]_pad ,
		_w9103_,
		_w9104_,
		_w20023_
	);
	LUT4 #(
		.INIT('hcdef)
	) name18123 (
		_w9098_,
		_w9101_,
		_w20022_,
		_w20023_,
		_w20024_
	);
	LUT4 #(
		.INIT('h7fff)
	) name18124 (
		_w20015_,
		_w20018_,
		_w20021_,
		_w20024_,
		_w20025_
	);
	LUT3 #(
		.INIT('h2a)
	) name18125 (
		\m3_addr_i[13]_pad ,
		_w9103_,
		_w9104_,
		_w20026_
	);
	LUT3 #(
		.INIT('h80)
	) name18126 (
		\m4_addr_i[13]_pad ,
		_w9103_,
		_w9104_,
		_w20027_
	);
	LUT4 #(
		.INIT('h9dbf)
	) name18127 (
		_w9098_,
		_w9101_,
		_w20026_,
		_w20027_,
		_w20028_
	);
	LUT3 #(
		.INIT('h80)
	) name18128 (
		\m6_addr_i[13]_pad ,
		_w9103_,
		_w9104_,
		_w20029_
	);
	LUT3 #(
		.INIT('h2a)
	) name18129 (
		\m7_addr_i[13]_pad ,
		_w9103_,
		_w9104_,
		_w20030_
	);
	LUT3 #(
		.INIT('h57)
	) name18130 (
		_w9102_,
		_w20029_,
		_w20030_,
		_w20031_
	);
	LUT3 #(
		.INIT('h2a)
	) name18131 (
		\m5_addr_i[13]_pad ,
		_w9103_,
		_w9104_,
		_w20032_
	);
	LUT3 #(
		.INIT('h80)
	) name18132 (
		\m0_addr_i[13]_pad ,
		_w9103_,
		_w9104_,
		_w20033_
	);
	LUT4 #(
		.INIT('h57df)
	) name18133 (
		_w9098_,
		_w9101_,
		_w20032_,
		_w20033_,
		_w20034_
	);
	LUT3 #(
		.INIT('h2a)
	) name18134 (
		\m1_addr_i[13]_pad ,
		_w9103_,
		_w9104_,
		_w20035_
	);
	LUT3 #(
		.INIT('h80)
	) name18135 (
		\m2_addr_i[13]_pad ,
		_w9103_,
		_w9104_,
		_w20036_
	);
	LUT4 #(
		.INIT('h3b7f)
	) name18136 (
		_w9098_,
		_w9101_,
		_w20035_,
		_w20036_,
		_w20037_
	);
	LUT4 #(
		.INIT('h7fff)
	) name18137 (
		_w20028_,
		_w20031_,
		_w20034_,
		_w20037_,
		_w20038_
	);
	LUT3 #(
		.INIT('h2a)
	) name18138 (
		\m3_addr_i[14]_pad ,
		_w9103_,
		_w9104_,
		_w20039_
	);
	LUT3 #(
		.INIT('h80)
	) name18139 (
		\m4_addr_i[14]_pad ,
		_w9103_,
		_w9104_,
		_w20040_
	);
	LUT4 #(
		.INIT('h9dbf)
	) name18140 (
		_w9098_,
		_w9101_,
		_w20039_,
		_w20040_,
		_w20041_
	);
	LUT3 #(
		.INIT('h80)
	) name18141 (
		\m6_addr_i[14]_pad ,
		_w9103_,
		_w9104_,
		_w20042_
	);
	LUT3 #(
		.INIT('h80)
	) name18142 (
		\m2_addr_i[14]_pad ,
		_w9103_,
		_w9104_,
		_w20043_
	);
	LUT4 #(
		.INIT('habef)
	) name18143 (
		_w9098_,
		_w9101_,
		_w20042_,
		_w20043_,
		_w20044_
	);
	LUT3 #(
		.INIT('h2a)
	) name18144 (
		\m5_addr_i[14]_pad ,
		_w9103_,
		_w9104_,
		_w20045_
	);
	LUT3 #(
		.INIT('h2a)
	) name18145 (
		\m1_addr_i[14]_pad ,
		_w9103_,
		_w9104_,
		_w20046_
	);
	LUT4 #(
		.INIT('h57df)
	) name18146 (
		_w9098_,
		_w9101_,
		_w20045_,
		_w20046_,
		_w20047_
	);
	LUT3 #(
		.INIT('h80)
	) name18147 (
		\m0_addr_i[14]_pad ,
		_w9103_,
		_w9104_,
		_w20048_
	);
	LUT3 #(
		.INIT('h2a)
	) name18148 (
		\m7_addr_i[14]_pad ,
		_w9103_,
		_w9104_,
		_w20049_
	);
	LUT4 #(
		.INIT('h6e7f)
	) name18149 (
		_w9098_,
		_w9101_,
		_w20048_,
		_w20049_,
		_w20050_
	);
	LUT4 #(
		.INIT('h7fff)
	) name18150 (
		_w20041_,
		_w20044_,
		_w20047_,
		_w20050_,
		_w20051_
	);
	LUT3 #(
		.INIT('h2a)
	) name18151 (
		\m3_addr_i[15]_pad ,
		_w9103_,
		_w9104_,
		_w20052_
	);
	LUT3 #(
		.INIT('h80)
	) name18152 (
		\m4_addr_i[15]_pad ,
		_w9103_,
		_w9104_,
		_w20053_
	);
	LUT4 #(
		.INIT('h9dbf)
	) name18153 (
		_w9098_,
		_w9101_,
		_w20052_,
		_w20053_,
		_w20054_
	);
	LUT3 #(
		.INIT('h80)
	) name18154 (
		\m6_addr_i[15]_pad ,
		_w9103_,
		_w9104_,
		_w20055_
	);
	LUT3 #(
		.INIT('h80)
	) name18155 (
		\m2_addr_i[15]_pad ,
		_w9103_,
		_w9104_,
		_w20056_
	);
	LUT4 #(
		.INIT('habef)
	) name18156 (
		_w9098_,
		_w9101_,
		_w20055_,
		_w20056_,
		_w20057_
	);
	LUT3 #(
		.INIT('h2a)
	) name18157 (
		\m5_addr_i[15]_pad ,
		_w9103_,
		_w9104_,
		_w20058_
	);
	LUT3 #(
		.INIT('h2a)
	) name18158 (
		\m1_addr_i[15]_pad ,
		_w9103_,
		_w9104_,
		_w20059_
	);
	LUT4 #(
		.INIT('h57df)
	) name18159 (
		_w9098_,
		_w9101_,
		_w20058_,
		_w20059_,
		_w20060_
	);
	LUT3 #(
		.INIT('h80)
	) name18160 (
		\m0_addr_i[15]_pad ,
		_w9103_,
		_w9104_,
		_w20061_
	);
	LUT3 #(
		.INIT('h2a)
	) name18161 (
		\m7_addr_i[15]_pad ,
		_w9103_,
		_w9104_,
		_w20062_
	);
	LUT4 #(
		.INIT('h6e7f)
	) name18162 (
		_w9098_,
		_w9101_,
		_w20061_,
		_w20062_,
		_w20063_
	);
	LUT4 #(
		.INIT('h7fff)
	) name18163 (
		_w20054_,
		_w20057_,
		_w20060_,
		_w20063_,
		_w20064_
	);
	LUT3 #(
		.INIT('h2a)
	) name18164 (
		\m1_addr_i[16]_pad ,
		_w9103_,
		_w9104_,
		_w20065_
	);
	LUT3 #(
		.INIT('h80)
	) name18165 (
		\m2_addr_i[16]_pad ,
		_w9103_,
		_w9104_,
		_w20066_
	);
	LUT4 #(
		.INIT('h3b7f)
	) name18166 (
		_w9098_,
		_w9101_,
		_w20065_,
		_w20066_,
		_w20067_
	);
	LUT3 #(
		.INIT('h80)
	) name18167 (
		\m6_addr_i[16]_pad ,
		_w9103_,
		_w9104_,
		_w20068_
	);
	LUT3 #(
		.INIT('h2a)
	) name18168 (
		\m7_addr_i[16]_pad ,
		_w9103_,
		_w9104_,
		_w20069_
	);
	LUT3 #(
		.INIT('h57)
	) name18169 (
		_w9102_,
		_w20068_,
		_w20069_,
		_w20070_
	);
	LUT3 #(
		.INIT('h2a)
	) name18170 (
		\m5_addr_i[16]_pad ,
		_w9103_,
		_w9104_,
		_w20071_
	);
	LUT3 #(
		.INIT('h80)
	) name18171 (
		\m0_addr_i[16]_pad ,
		_w9103_,
		_w9104_,
		_w20072_
	);
	LUT4 #(
		.INIT('h57df)
	) name18172 (
		_w9098_,
		_w9101_,
		_w20071_,
		_w20072_,
		_w20073_
	);
	LUT3 #(
		.INIT('h2a)
	) name18173 (
		\m3_addr_i[16]_pad ,
		_w9103_,
		_w9104_,
		_w20074_
	);
	LUT3 #(
		.INIT('h80)
	) name18174 (
		\m4_addr_i[16]_pad ,
		_w9103_,
		_w9104_,
		_w20075_
	);
	LUT4 #(
		.INIT('h9dbf)
	) name18175 (
		_w9098_,
		_w9101_,
		_w20074_,
		_w20075_,
		_w20076_
	);
	LUT4 #(
		.INIT('h7fff)
	) name18176 (
		_w20067_,
		_w20070_,
		_w20073_,
		_w20076_,
		_w20077_
	);
	LUT3 #(
		.INIT('h80)
	) name18177 (
		\m6_addr_i[17]_pad ,
		_w9103_,
		_w9104_,
		_w20078_
	);
	LUT3 #(
		.INIT('h2a)
	) name18178 (
		\m5_addr_i[17]_pad ,
		_w9103_,
		_w9104_,
		_w20079_
	);
	LUT4 #(
		.INIT('hcdef)
	) name18179 (
		_w9098_,
		_w9101_,
		_w20078_,
		_w20079_,
		_w20080_
	);
	LUT3 #(
		.INIT('h80)
	) name18180 (
		\m0_addr_i[17]_pad ,
		_w9103_,
		_w9104_,
		_w20081_
	);
	LUT3 #(
		.INIT('h80)
	) name18181 (
		\m4_addr_i[17]_pad ,
		_w9103_,
		_w9104_,
		_w20082_
	);
	LUT4 #(
		.INIT('h5d7f)
	) name18182 (
		_w9098_,
		_w9101_,
		_w20081_,
		_w20082_,
		_w20083_
	);
	LUT3 #(
		.INIT('h2a)
	) name18183 (
		\m7_addr_i[17]_pad ,
		_w9103_,
		_w9104_,
		_w20084_
	);
	LUT3 #(
		.INIT('h2a)
	) name18184 (
		\m3_addr_i[17]_pad ,
		_w9103_,
		_w9104_,
		_w20085_
	);
	LUT4 #(
		.INIT('habef)
	) name18185 (
		_w9098_,
		_w9101_,
		_w20084_,
		_w20085_,
		_w20086_
	);
	LUT3 #(
		.INIT('h2a)
	) name18186 (
		\m1_addr_i[17]_pad ,
		_w9103_,
		_w9104_,
		_w20087_
	);
	LUT3 #(
		.INIT('h80)
	) name18187 (
		\m2_addr_i[17]_pad ,
		_w9103_,
		_w9104_,
		_w20088_
	);
	LUT4 #(
		.INIT('h3b7f)
	) name18188 (
		_w9098_,
		_w9101_,
		_w20087_,
		_w20088_,
		_w20089_
	);
	LUT4 #(
		.INIT('h7fff)
	) name18189 (
		_w20080_,
		_w20083_,
		_w20086_,
		_w20089_,
		_w20090_
	);
	LUT3 #(
		.INIT('h2a)
	) name18190 (
		\m3_addr_i[18]_pad ,
		_w9103_,
		_w9104_,
		_w20091_
	);
	LUT3 #(
		.INIT('h80)
	) name18191 (
		\m4_addr_i[18]_pad ,
		_w9103_,
		_w9104_,
		_w20092_
	);
	LUT4 #(
		.INIT('h9dbf)
	) name18192 (
		_w9098_,
		_w9101_,
		_w20091_,
		_w20092_,
		_w20093_
	);
	LUT3 #(
		.INIT('h80)
	) name18193 (
		\m6_addr_i[18]_pad ,
		_w9103_,
		_w9104_,
		_w20094_
	);
	LUT3 #(
		.INIT('h80)
	) name18194 (
		\m2_addr_i[18]_pad ,
		_w9103_,
		_w9104_,
		_w20095_
	);
	LUT4 #(
		.INIT('habef)
	) name18195 (
		_w9098_,
		_w9101_,
		_w20094_,
		_w20095_,
		_w20096_
	);
	LUT3 #(
		.INIT('h2a)
	) name18196 (
		\m5_addr_i[18]_pad ,
		_w9103_,
		_w9104_,
		_w20097_
	);
	LUT3 #(
		.INIT('h2a)
	) name18197 (
		\m1_addr_i[18]_pad ,
		_w9103_,
		_w9104_,
		_w20098_
	);
	LUT4 #(
		.INIT('h57df)
	) name18198 (
		_w9098_,
		_w9101_,
		_w20097_,
		_w20098_,
		_w20099_
	);
	LUT3 #(
		.INIT('h80)
	) name18199 (
		\m0_addr_i[18]_pad ,
		_w9103_,
		_w9104_,
		_w20100_
	);
	LUT3 #(
		.INIT('h2a)
	) name18200 (
		\m7_addr_i[18]_pad ,
		_w9103_,
		_w9104_,
		_w20101_
	);
	LUT4 #(
		.INIT('h6e7f)
	) name18201 (
		_w9098_,
		_w9101_,
		_w20100_,
		_w20101_,
		_w20102_
	);
	LUT4 #(
		.INIT('h7fff)
	) name18202 (
		_w20093_,
		_w20096_,
		_w20099_,
		_w20102_,
		_w20103_
	);
	LUT3 #(
		.INIT('h2a)
	) name18203 (
		\m3_addr_i[19]_pad ,
		_w9103_,
		_w9104_,
		_w20104_
	);
	LUT3 #(
		.INIT('h80)
	) name18204 (
		\m4_addr_i[19]_pad ,
		_w9103_,
		_w9104_,
		_w20105_
	);
	LUT4 #(
		.INIT('h9dbf)
	) name18205 (
		_w9098_,
		_w9101_,
		_w20104_,
		_w20105_,
		_w20106_
	);
	LUT3 #(
		.INIT('h80)
	) name18206 (
		\m6_addr_i[19]_pad ,
		_w9103_,
		_w9104_,
		_w20107_
	);
	LUT3 #(
		.INIT('h80)
	) name18207 (
		\m2_addr_i[19]_pad ,
		_w9103_,
		_w9104_,
		_w20108_
	);
	LUT4 #(
		.INIT('habef)
	) name18208 (
		_w9098_,
		_w9101_,
		_w20107_,
		_w20108_,
		_w20109_
	);
	LUT3 #(
		.INIT('h2a)
	) name18209 (
		\m5_addr_i[19]_pad ,
		_w9103_,
		_w9104_,
		_w20110_
	);
	LUT3 #(
		.INIT('h2a)
	) name18210 (
		\m1_addr_i[19]_pad ,
		_w9103_,
		_w9104_,
		_w20111_
	);
	LUT4 #(
		.INIT('h57df)
	) name18211 (
		_w9098_,
		_w9101_,
		_w20110_,
		_w20111_,
		_w20112_
	);
	LUT3 #(
		.INIT('h80)
	) name18212 (
		\m0_addr_i[19]_pad ,
		_w9103_,
		_w9104_,
		_w20113_
	);
	LUT3 #(
		.INIT('h2a)
	) name18213 (
		\m7_addr_i[19]_pad ,
		_w9103_,
		_w9104_,
		_w20114_
	);
	LUT4 #(
		.INIT('h6e7f)
	) name18214 (
		_w9098_,
		_w9101_,
		_w20113_,
		_w20114_,
		_w20115_
	);
	LUT4 #(
		.INIT('h7fff)
	) name18215 (
		_w20106_,
		_w20109_,
		_w20112_,
		_w20115_,
		_w20116_
	);
	LUT3 #(
		.INIT('h2a)
	) name18216 (
		\m3_addr_i[1]_pad ,
		_w9103_,
		_w9104_,
		_w20117_
	);
	LUT3 #(
		.INIT('h80)
	) name18217 (
		\m4_addr_i[1]_pad ,
		_w9103_,
		_w9104_,
		_w20118_
	);
	LUT4 #(
		.INIT('h9dbf)
	) name18218 (
		_w9098_,
		_w9101_,
		_w20117_,
		_w20118_,
		_w20119_
	);
	LUT3 #(
		.INIT('h80)
	) name18219 (
		\m6_addr_i[1]_pad ,
		_w9103_,
		_w9104_,
		_w20120_
	);
	LUT3 #(
		.INIT('h80)
	) name18220 (
		\m2_addr_i[1]_pad ,
		_w9103_,
		_w9104_,
		_w20121_
	);
	LUT4 #(
		.INIT('habef)
	) name18221 (
		_w9098_,
		_w9101_,
		_w20120_,
		_w20121_,
		_w20122_
	);
	LUT3 #(
		.INIT('h2a)
	) name18222 (
		\m5_addr_i[1]_pad ,
		_w9103_,
		_w9104_,
		_w20123_
	);
	LUT3 #(
		.INIT('h2a)
	) name18223 (
		\m1_addr_i[1]_pad ,
		_w9103_,
		_w9104_,
		_w20124_
	);
	LUT4 #(
		.INIT('h57df)
	) name18224 (
		_w9098_,
		_w9101_,
		_w20123_,
		_w20124_,
		_w20125_
	);
	LUT3 #(
		.INIT('h80)
	) name18225 (
		\m0_addr_i[1]_pad ,
		_w9103_,
		_w9104_,
		_w20126_
	);
	LUT3 #(
		.INIT('h2a)
	) name18226 (
		\m7_addr_i[1]_pad ,
		_w9103_,
		_w9104_,
		_w20127_
	);
	LUT4 #(
		.INIT('h6e7f)
	) name18227 (
		_w9098_,
		_w9101_,
		_w20126_,
		_w20127_,
		_w20128_
	);
	LUT4 #(
		.INIT('h7fff)
	) name18228 (
		_w20119_,
		_w20122_,
		_w20125_,
		_w20128_,
		_w20129_
	);
	LUT3 #(
		.INIT('h2a)
	) name18229 (
		\m1_addr_i[20]_pad ,
		_w9103_,
		_w9104_,
		_w20130_
	);
	LUT3 #(
		.INIT('h80)
	) name18230 (
		\m2_addr_i[20]_pad ,
		_w9103_,
		_w9104_,
		_w20131_
	);
	LUT4 #(
		.INIT('h3b7f)
	) name18231 (
		_w9098_,
		_w9101_,
		_w20130_,
		_w20131_,
		_w20132_
	);
	LUT3 #(
		.INIT('h2a)
	) name18232 (
		\m3_addr_i[20]_pad ,
		_w9103_,
		_w9104_,
		_w20133_
	);
	LUT3 #(
		.INIT('h2a)
	) name18233 (
		\m7_addr_i[20]_pad ,
		_w9103_,
		_w9104_,
		_w20134_
	);
	LUT4 #(
		.INIT('haebf)
	) name18234 (
		_w9098_,
		_w9101_,
		_w20133_,
		_w20134_,
		_w20135_
	);
	LUT3 #(
		.INIT('h80)
	) name18235 (
		\m4_addr_i[20]_pad ,
		_w9103_,
		_w9104_,
		_w20136_
	);
	LUT3 #(
		.INIT('h80)
	) name18236 (
		\m0_addr_i[20]_pad ,
		_w9103_,
		_w9104_,
		_w20137_
	);
	LUT4 #(
		.INIT('h57df)
	) name18237 (
		_w9098_,
		_w9101_,
		_w20136_,
		_w20137_,
		_w20138_
	);
	LUT3 #(
		.INIT('h80)
	) name18238 (
		\m6_addr_i[20]_pad ,
		_w9103_,
		_w9104_,
		_w20139_
	);
	LUT3 #(
		.INIT('h2a)
	) name18239 (
		\m5_addr_i[20]_pad ,
		_w9103_,
		_w9104_,
		_w20140_
	);
	LUT4 #(
		.INIT('hcdef)
	) name18240 (
		_w9098_,
		_w9101_,
		_w20139_,
		_w20140_,
		_w20141_
	);
	LUT4 #(
		.INIT('h7fff)
	) name18241 (
		_w20132_,
		_w20135_,
		_w20138_,
		_w20141_,
		_w20142_
	);
	LUT3 #(
		.INIT('h80)
	) name18242 (
		\m0_addr_i[21]_pad ,
		_w9103_,
		_w9104_,
		_w20143_
	);
	LUT3 #(
		.INIT('h2a)
	) name18243 (
		\m7_addr_i[21]_pad ,
		_w9103_,
		_w9104_,
		_w20144_
	);
	LUT4 #(
		.INIT('h6e7f)
	) name18244 (
		_w9098_,
		_w9101_,
		_w20143_,
		_w20144_,
		_w20145_
	);
	LUT3 #(
		.INIT('h2a)
	) name18245 (
		\m1_addr_i[21]_pad ,
		_w9103_,
		_w9104_,
		_w20146_
	);
	LUT3 #(
		.INIT('h2a)
	) name18246 (
		\m5_addr_i[21]_pad ,
		_w9103_,
		_w9104_,
		_w20147_
	);
	LUT4 #(
		.INIT('h5d7f)
	) name18247 (
		_w9098_,
		_w9101_,
		_w20146_,
		_w20147_,
		_w20148_
	);
	LUT3 #(
		.INIT('h80)
	) name18248 (
		\m2_addr_i[21]_pad ,
		_w9103_,
		_w9104_,
		_w20149_
	);
	LUT3 #(
		.INIT('h80)
	) name18249 (
		\m6_addr_i[21]_pad ,
		_w9103_,
		_w9104_,
		_w20150_
	);
	LUT4 #(
		.INIT('haebf)
	) name18250 (
		_w9098_,
		_w9101_,
		_w20149_,
		_w20150_,
		_w20151_
	);
	LUT3 #(
		.INIT('h2a)
	) name18251 (
		\m3_addr_i[21]_pad ,
		_w9103_,
		_w9104_,
		_w20152_
	);
	LUT3 #(
		.INIT('h80)
	) name18252 (
		\m4_addr_i[21]_pad ,
		_w9103_,
		_w9104_,
		_w20153_
	);
	LUT4 #(
		.INIT('h9dbf)
	) name18253 (
		_w9098_,
		_w9101_,
		_w20152_,
		_w20153_,
		_w20154_
	);
	LUT4 #(
		.INIT('h7fff)
	) name18254 (
		_w20145_,
		_w20148_,
		_w20151_,
		_w20154_,
		_w20155_
	);
	LUT3 #(
		.INIT('h2a)
	) name18255 (
		\m1_addr_i[22]_pad ,
		_w9103_,
		_w9104_,
		_w20156_
	);
	LUT3 #(
		.INIT('h80)
	) name18256 (
		\m2_addr_i[22]_pad ,
		_w9103_,
		_w9104_,
		_w20157_
	);
	LUT4 #(
		.INIT('h3b7f)
	) name18257 (
		_w9098_,
		_w9101_,
		_w20156_,
		_w20157_,
		_w20158_
	);
	LUT3 #(
		.INIT('h2a)
	) name18258 (
		\m3_addr_i[22]_pad ,
		_w9103_,
		_w9104_,
		_w20159_
	);
	LUT3 #(
		.INIT('h2a)
	) name18259 (
		\m7_addr_i[22]_pad ,
		_w9103_,
		_w9104_,
		_w20160_
	);
	LUT4 #(
		.INIT('haebf)
	) name18260 (
		_w9098_,
		_w9101_,
		_w20159_,
		_w20160_,
		_w20161_
	);
	LUT3 #(
		.INIT('h80)
	) name18261 (
		\m4_addr_i[22]_pad ,
		_w9103_,
		_w9104_,
		_w20162_
	);
	LUT3 #(
		.INIT('h80)
	) name18262 (
		\m0_addr_i[22]_pad ,
		_w9103_,
		_w9104_,
		_w20163_
	);
	LUT4 #(
		.INIT('h57df)
	) name18263 (
		_w9098_,
		_w9101_,
		_w20162_,
		_w20163_,
		_w20164_
	);
	LUT3 #(
		.INIT('h80)
	) name18264 (
		\m6_addr_i[22]_pad ,
		_w9103_,
		_w9104_,
		_w20165_
	);
	LUT3 #(
		.INIT('h2a)
	) name18265 (
		\m5_addr_i[22]_pad ,
		_w9103_,
		_w9104_,
		_w20166_
	);
	LUT4 #(
		.INIT('hcdef)
	) name18266 (
		_w9098_,
		_w9101_,
		_w20165_,
		_w20166_,
		_w20167_
	);
	LUT4 #(
		.INIT('h7fff)
	) name18267 (
		_w20158_,
		_w20161_,
		_w20164_,
		_w20167_,
		_w20168_
	);
	LUT3 #(
		.INIT('h2a)
	) name18268 (
		\m1_addr_i[23]_pad ,
		_w9103_,
		_w9104_,
		_w20169_
	);
	LUT3 #(
		.INIT('h80)
	) name18269 (
		\m2_addr_i[23]_pad ,
		_w9103_,
		_w9104_,
		_w20170_
	);
	LUT4 #(
		.INIT('h3b7f)
	) name18270 (
		_w9098_,
		_w9101_,
		_w20169_,
		_w20170_,
		_w20171_
	);
	LUT3 #(
		.INIT('h80)
	) name18271 (
		\m0_addr_i[23]_pad ,
		_w9103_,
		_w9104_,
		_w20172_
	);
	LUT3 #(
		.INIT('h2a)
	) name18272 (
		\m5_addr_i[23]_pad ,
		_w9103_,
		_w9104_,
		_w20173_
	);
	LUT4 #(
		.INIT('h5d7f)
	) name18273 (
		_w9098_,
		_w9101_,
		_w20172_,
		_w20173_,
		_w20174_
	);
	LUT3 #(
		.INIT('h2a)
	) name18274 (
		\m7_addr_i[23]_pad ,
		_w9103_,
		_w9104_,
		_w20175_
	);
	LUT3 #(
		.INIT('h80)
	) name18275 (
		\m6_addr_i[23]_pad ,
		_w9103_,
		_w9104_,
		_w20176_
	);
	LUT3 #(
		.INIT('h57)
	) name18276 (
		_w9102_,
		_w20175_,
		_w20176_,
		_w20177_
	);
	LUT3 #(
		.INIT('h2a)
	) name18277 (
		\m3_addr_i[23]_pad ,
		_w9103_,
		_w9104_,
		_w20178_
	);
	LUT3 #(
		.INIT('h80)
	) name18278 (
		\m4_addr_i[23]_pad ,
		_w9103_,
		_w9104_,
		_w20179_
	);
	LUT4 #(
		.INIT('h9dbf)
	) name18279 (
		_w9098_,
		_w9101_,
		_w20178_,
		_w20179_,
		_w20180_
	);
	LUT4 #(
		.INIT('h7fff)
	) name18280 (
		_w20171_,
		_w20174_,
		_w20177_,
		_w20180_,
		_w20181_
	);
	LUT3 #(
		.INIT('h2a)
	) name18281 (
		\m5_addr_i[24]_pad ,
		_w9103_,
		_w9104_,
		_w20182_
	);
	LUT3 #(
		.INIT('h80)
	) name18282 (
		\m6_addr_i[24]_pad ,
		_w9103_,
		_w9104_,
		_w20183_
	);
	LUT4 #(
		.INIT('hcedf)
	) name18283 (
		_w9098_,
		_w9101_,
		_w20182_,
		_w20183_,
		_w20184_
	);
	LUT3 #(
		.INIT('h2a)
	) name18284 (
		\m1_addr_i[24]_pad ,
		_w9103_,
		_w9104_,
		_w20185_
	);
	LUT3 #(
		.INIT('h2a)
	) name18285 (
		\m7_addr_i[24]_pad ,
		_w9103_,
		_w9104_,
		_w20186_
	);
	LUT4 #(
		.INIT('h6e7f)
	) name18286 (
		_w9098_,
		_w9101_,
		_w20185_,
		_w20186_,
		_w20187_
	);
	LUT3 #(
		.INIT('h80)
	) name18287 (
		\m2_addr_i[24]_pad ,
		_w9103_,
		_w9104_,
		_w20188_
	);
	LUT3 #(
		.INIT('h80)
	) name18288 (
		\m0_addr_i[24]_pad ,
		_w9103_,
		_w9104_,
		_w20189_
	);
	LUT4 #(
		.INIT('h37bf)
	) name18289 (
		_w9098_,
		_w9101_,
		_w20188_,
		_w20189_,
		_w20190_
	);
	LUT3 #(
		.INIT('h2a)
	) name18290 (
		\m3_addr_i[24]_pad ,
		_w9103_,
		_w9104_,
		_w20191_
	);
	LUT3 #(
		.INIT('h80)
	) name18291 (
		\m4_addr_i[24]_pad ,
		_w9103_,
		_w9104_,
		_w20192_
	);
	LUT4 #(
		.INIT('h9dbf)
	) name18292 (
		_w9098_,
		_w9101_,
		_w20191_,
		_w20192_,
		_w20193_
	);
	LUT4 #(
		.INIT('h7fff)
	) name18293 (
		_w20184_,
		_w20187_,
		_w20190_,
		_w20193_,
		_w20194_
	);
	LUT3 #(
		.INIT('h2a)
	) name18294 (
		\m1_addr_i[25]_pad ,
		_w9103_,
		_w9104_,
		_w20195_
	);
	LUT3 #(
		.INIT('h80)
	) name18295 (
		\m2_addr_i[25]_pad ,
		_w9103_,
		_w9104_,
		_w20196_
	);
	LUT4 #(
		.INIT('h3b7f)
	) name18296 (
		_w9098_,
		_w9101_,
		_w20195_,
		_w20196_,
		_w20197_
	);
	LUT3 #(
		.INIT('h80)
	) name18297 (
		\m0_addr_i[25]_pad ,
		_w9103_,
		_w9104_,
		_w20198_
	);
	LUT3 #(
		.INIT('h80)
	) name18298 (
		\m4_addr_i[25]_pad ,
		_w9103_,
		_w9104_,
		_w20199_
	);
	LUT4 #(
		.INIT('h5d7f)
	) name18299 (
		_w9098_,
		_w9101_,
		_w20198_,
		_w20199_,
		_w20200_
	);
	LUT3 #(
		.INIT('h2a)
	) name18300 (
		\m7_addr_i[25]_pad ,
		_w9103_,
		_w9104_,
		_w20201_
	);
	LUT3 #(
		.INIT('h2a)
	) name18301 (
		\m3_addr_i[25]_pad ,
		_w9103_,
		_w9104_,
		_w20202_
	);
	LUT4 #(
		.INIT('habef)
	) name18302 (
		_w9098_,
		_w9101_,
		_w20201_,
		_w20202_,
		_w20203_
	);
	LUT3 #(
		.INIT('h2a)
	) name18303 (
		\m5_addr_i[25]_pad ,
		_w9103_,
		_w9104_,
		_w20204_
	);
	LUT3 #(
		.INIT('h80)
	) name18304 (
		\m6_addr_i[25]_pad ,
		_w9103_,
		_w9104_,
		_w20205_
	);
	LUT4 #(
		.INIT('hcedf)
	) name18305 (
		_w9098_,
		_w9101_,
		_w20204_,
		_w20205_,
		_w20206_
	);
	LUT4 #(
		.INIT('h7fff)
	) name18306 (
		_w20197_,
		_w20200_,
		_w20203_,
		_w20206_,
		_w20207_
	);
	LUT3 #(
		.INIT('h2a)
	) name18307 (
		\m3_addr_i[26]_pad ,
		_w9103_,
		_w9104_,
		_w20208_
	);
	LUT3 #(
		.INIT('h80)
	) name18308 (
		\m4_addr_i[26]_pad ,
		_w9103_,
		_w9104_,
		_w20209_
	);
	LUT4 #(
		.INIT('h9dbf)
	) name18309 (
		_w9098_,
		_w9101_,
		_w20208_,
		_w20209_,
		_w20210_
	);
	LUT3 #(
		.INIT('h2a)
	) name18310 (
		\m1_addr_i[26]_pad ,
		_w9103_,
		_w9104_,
		_w20211_
	);
	LUT3 #(
		.INIT('h2a)
	) name18311 (
		\m7_addr_i[26]_pad ,
		_w9103_,
		_w9104_,
		_w20212_
	);
	LUT4 #(
		.INIT('h6e7f)
	) name18312 (
		_w9098_,
		_w9101_,
		_w20211_,
		_w20212_,
		_w20213_
	);
	LUT3 #(
		.INIT('h80)
	) name18313 (
		\m2_addr_i[26]_pad ,
		_w9103_,
		_w9104_,
		_w20214_
	);
	LUT3 #(
		.INIT('h80)
	) name18314 (
		\m0_addr_i[26]_pad ,
		_w9103_,
		_w9104_,
		_w20215_
	);
	LUT4 #(
		.INIT('h37bf)
	) name18315 (
		_w9098_,
		_w9101_,
		_w20214_,
		_w20215_,
		_w20216_
	);
	LUT3 #(
		.INIT('h2a)
	) name18316 (
		\m5_addr_i[26]_pad ,
		_w9103_,
		_w9104_,
		_w20217_
	);
	LUT3 #(
		.INIT('h80)
	) name18317 (
		\m6_addr_i[26]_pad ,
		_w9103_,
		_w9104_,
		_w20218_
	);
	LUT4 #(
		.INIT('hcedf)
	) name18318 (
		_w9098_,
		_w9101_,
		_w20217_,
		_w20218_,
		_w20219_
	);
	LUT4 #(
		.INIT('h7fff)
	) name18319 (
		_w20210_,
		_w20213_,
		_w20216_,
		_w20219_,
		_w20220_
	);
	LUT3 #(
		.INIT('h2a)
	) name18320 (
		\m1_addr_i[27]_pad ,
		_w9103_,
		_w9104_,
		_w20221_
	);
	LUT3 #(
		.INIT('h80)
	) name18321 (
		\m2_addr_i[27]_pad ,
		_w9103_,
		_w9104_,
		_w20222_
	);
	LUT4 #(
		.INIT('h3b7f)
	) name18322 (
		_w9098_,
		_w9101_,
		_w20221_,
		_w20222_,
		_w20223_
	);
	LUT3 #(
		.INIT('h80)
	) name18323 (
		\m0_addr_i[27]_pad ,
		_w9103_,
		_w9104_,
		_w20224_
	);
	LUT3 #(
		.INIT('h80)
	) name18324 (
		\m6_addr_i[27]_pad ,
		_w9103_,
		_w9104_,
		_w20225_
	);
	LUT4 #(
		.INIT('h6e7f)
	) name18325 (
		_w9098_,
		_w9101_,
		_w20224_,
		_w20225_,
		_w20226_
	);
	LUT3 #(
		.INIT('h2a)
	) name18326 (
		\m7_addr_i[27]_pad ,
		_w9103_,
		_w9104_,
		_w20227_
	);
	LUT3 #(
		.INIT('h2a)
	) name18327 (
		\m5_addr_i[27]_pad ,
		_w9103_,
		_w9104_,
		_w20228_
	);
	LUT4 #(
		.INIT('hcdef)
	) name18328 (
		_w9098_,
		_w9101_,
		_w20227_,
		_w20228_,
		_w20229_
	);
	LUT3 #(
		.INIT('h2a)
	) name18329 (
		\m3_addr_i[27]_pad ,
		_w9103_,
		_w9104_,
		_w20230_
	);
	LUT3 #(
		.INIT('h80)
	) name18330 (
		\m4_addr_i[27]_pad ,
		_w9103_,
		_w9104_,
		_w20231_
	);
	LUT4 #(
		.INIT('h9dbf)
	) name18331 (
		_w9098_,
		_w9101_,
		_w20230_,
		_w20231_,
		_w20232_
	);
	LUT4 #(
		.INIT('h7fff)
	) name18332 (
		_w20223_,
		_w20226_,
		_w20229_,
		_w20232_,
		_w20233_
	);
	LUT3 #(
		.INIT('h2a)
	) name18333 (
		\m1_addr_i[28]_pad ,
		_w9103_,
		_w9104_,
		_w20234_
	);
	LUT3 #(
		.INIT('h80)
	) name18334 (
		\m2_addr_i[28]_pad ,
		_w9103_,
		_w9104_,
		_w20235_
	);
	LUT4 #(
		.INIT('h3b7f)
	) name18335 (
		_w9098_,
		_w9101_,
		_w20234_,
		_w20235_,
		_w20236_
	);
	LUT3 #(
		.INIT('h80)
	) name18336 (
		\m0_addr_i[28]_pad ,
		_w9103_,
		_w9104_,
		_w20237_
	);
	LUT3 #(
		.INIT('h80)
	) name18337 (
		\m4_addr_i[28]_pad ,
		_w9103_,
		_w9104_,
		_w20238_
	);
	LUT4 #(
		.INIT('h5d7f)
	) name18338 (
		_w9098_,
		_w9101_,
		_w20237_,
		_w20238_,
		_w20239_
	);
	LUT3 #(
		.INIT('h2a)
	) name18339 (
		\m7_addr_i[28]_pad ,
		_w9103_,
		_w9104_,
		_w20240_
	);
	LUT3 #(
		.INIT('h2a)
	) name18340 (
		\m3_addr_i[28]_pad ,
		_w9103_,
		_w9104_,
		_w20241_
	);
	LUT4 #(
		.INIT('habef)
	) name18341 (
		_w9098_,
		_w9101_,
		_w20240_,
		_w20241_,
		_w20242_
	);
	LUT3 #(
		.INIT('h2a)
	) name18342 (
		\m5_addr_i[28]_pad ,
		_w9103_,
		_w9104_,
		_w20243_
	);
	LUT3 #(
		.INIT('h80)
	) name18343 (
		\m6_addr_i[28]_pad ,
		_w9103_,
		_w9104_,
		_w20244_
	);
	LUT4 #(
		.INIT('hcedf)
	) name18344 (
		_w9098_,
		_w9101_,
		_w20243_,
		_w20244_,
		_w20245_
	);
	LUT4 #(
		.INIT('h7fff)
	) name18345 (
		_w20236_,
		_w20239_,
		_w20242_,
		_w20245_,
		_w20246_
	);
	LUT3 #(
		.INIT('h80)
	) name18346 (
		\m0_addr_i[29]_pad ,
		_w9103_,
		_w9104_,
		_w20247_
	);
	LUT3 #(
		.INIT('h2a)
	) name18347 (
		\m7_addr_i[29]_pad ,
		_w9103_,
		_w9104_,
		_w20248_
	);
	LUT4 #(
		.INIT('h6e7f)
	) name18348 (
		_w9098_,
		_w9101_,
		_w20247_,
		_w20248_,
		_w20249_
	);
	LUT3 #(
		.INIT('h2a)
	) name18349 (
		\m5_addr_i[29]_pad ,
		_w9103_,
		_w9104_,
		_w20250_
	);
	LUT3 #(
		.INIT('h80)
	) name18350 (
		\m4_addr_i[29]_pad ,
		_w9103_,
		_w9104_,
		_w20251_
	);
	LUT3 #(
		.INIT('h57)
	) name18351 (
		_w9116_,
		_w20250_,
		_w20251_,
		_w20252_
	);
	LUT3 #(
		.INIT('h80)
	) name18352 (
		\m6_addr_i[29]_pad ,
		_w9103_,
		_w9104_,
		_w20253_
	);
	LUT3 #(
		.INIT('h2a)
	) name18353 (
		\m3_addr_i[29]_pad ,
		_w9103_,
		_w9104_,
		_w20254_
	);
	LUT4 #(
		.INIT('habef)
	) name18354 (
		_w9098_,
		_w9101_,
		_w20253_,
		_w20254_,
		_w20255_
	);
	LUT3 #(
		.INIT('h2a)
	) name18355 (
		\m1_addr_i[29]_pad ,
		_w9103_,
		_w9104_,
		_w20256_
	);
	LUT3 #(
		.INIT('h80)
	) name18356 (
		\m2_addr_i[29]_pad ,
		_w9103_,
		_w9104_,
		_w20257_
	);
	LUT4 #(
		.INIT('h3b7f)
	) name18357 (
		_w9098_,
		_w9101_,
		_w20256_,
		_w20257_,
		_w20258_
	);
	LUT4 #(
		.INIT('h7fff)
	) name18358 (
		_w20249_,
		_w20252_,
		_w20255_,
		_w20258_,
		_w20259_
	);
	LUT3 #(
		.INIT('h2a)
	) name18359 (
		\m3_addr_i[2]_pad ,
		_w9103_,
		_w9104_,
		_w20260_
	);
	LUT3 #(
		.INIT('h80)
	) name18360 (
		\m4_addr_i[2]_pad ,
		_w9103_,
		_w9104_,
		_w20261_
	);
	LUT4 #(
		.INIT('h9dbf)
	) name18361 (
		_w9098_,
		_w9101_,
		_w20260_,
		_w20261_,
		_w20262_
	);
	LUT3 #(
		.INIT('h80)
	) name18362 (
		\m6_addr_i[2]_pad ,
		_w9103_,
		_w9104_,
		_w20263_
	);
	LUT3 #(
		.INIT('h80)
	) name18363 (
		\m2_addr_i[2]_pad ,
		_w9103_,
		_w9104_,
		_w20264_
	);
	LUT4 #(
		.INIT('habef)
	) name18364 (
		_w9098_,
		_w9101_,
		_w20263_,
		_w20264_,
		_w20265_
	);
	LUT3 #(
		.INIT('h2a)
	) name18365 (
		\m5_addr_i[2]_pad ,
		_w9103_,
		_w9104_,
		_w20266_
	);
	LUT3 #(
		.INIT('h2a)
	) name18366 (
		\m1_addr_i[2]_pad ,
		_w9103_,
		_w9104_,
		_w20267_
	);
	LUT4 #(
		.INIT('h57df)
	) name18367 (
		_w9098_,
		_w9101_,
		_w20266_,
		_w20267_,
		_w20268_
	);
	LUT3 #(
		.INIT('h80)
	) name18368 (
		\m0_addr_i[2]_pad ,
		_w9103_,
		_w9104_,
		_w20269_
	);
	LUT3 #(
		.INIT('h2a)
	) name18369 (
		\m7_addr_i[2]_pad ,
		_w9103_,
		_w9104_,
		_w20270_
	);
	LUT4 #(
		.INIT('h6e7f)
	) name18370 (
		_w9098_,
		_w9101_,
		_w20269_,
		_w20270_,
		_w20271_
	);
	LUT4 #(
		.INIT('h7fff)
	) name18371 (
		_w20262_,
		_w20265_,
		_w20268_,
		_w20271_,
		_w20272_
	);
	LUT3 #(
		.INIT('h2a)
	) name18372 (
		\m3_addr_i[30]_pad ,
		_w9103_,
		_w9104_,
		_w20273_
	);
	LUT3 #(
		.INIT('h80)
	) name18373 (
		\m4_addr_i[30]_pad ,
		_w9103_,
		_w9104_,
		_w20274_
	);
	LUT4 #(
		.INIT('h9dbf)
	) name18374 (
		_w9098_,
		_w9101_,
		_w20273_,
		_w20274_,
		_w20275_
	);
	LUT3 #(
		.INIT('h80)
	) name18375 (
		\m0_addr_i[30]_pad ,
		_w9103_,
		_w9104_,
		_w20276_
	);
	LUT3 #(
		.INIT('h80)
	) name18376 (
		\m6_addr_i[30]_pad ,
		_w9103_,
		_w9104_,
		_w20277_
	);
	LUT4 #(
		.INIT('h6e7f)
	) name18377 (
		_w9098_,
		_w9101_,
		_w20276_,
		_w20277_,
		_w20278_
	);
	LUT3 #(
		.INIT('h2a)
	) name18378 (
		\m7_addr_i[30]_pad ,
		_w9103_,
		_w9104_,
		_w20279_
	);
	LUT3 #(
		.INIT('h2a)
	) name18379 (
		\m5_addr_i[30]_pad ,
		_w9103_,
		_w9104_,
		_w20280_
	);
	LUT4 #(
		.INIT('hcdef)
	) name18380 (
		_w9098_,
		_w9101_,
		_w20279_,
		_w20280_,
		_w20281_
	);
	LUT3 #(
		.INIT('h2a)
	) name18381 (
		\m1_addr_i[30]_pad ,
		_w9103_,
		_w9104_,
		_w20282_
	);
	LUT3 #(
		.INIT('h80)
	) name18382 (
		\m2_addr_i[30]_pad ,
		_w9103_,
		_w9104_,
		_w20283_
	);
	LUT4 #(
		.INIT('h3b7f)
	) name18383 (
		_w9098_,
		_w9101_,
		_w20282_,
		_w20283_,
		_w20284_
	);
	LUT4 #(
		.INIT('h7fff)
	) name18384 (
		_w20275_,
		_w20278_,
		_w20281_,
		_w20284_,
		_w20285_
	);
	LUT3 #(
		.INIT('h2a)
	) name18385 (
		\m5_addr_i[31]_pad ,
		_w9103_,
		_w9104_,
		_w20286_
	);
	LUT3 #(
		.INIT('h80)
	) name18386 (
		\m6_addr_i[31]_pad ,
		_w9103_,
		_w9104_,
		_w20287_
	);
	LUT4 #(
		.INIT('hcedf)
	) name18387 (
		_w9098_,
		_w9101_,
		_w20286_,
		_w20287_,
		_w20288_
	);
	LUT3 #(
		.INIT('h2a)
	) name18388 (
		\m1_addr_i[31]_pad ,
		_w9103_,
		_w9104_,
		_w20289_
	);
	LUT3 #(
		.INIT('h80)
	) name18389 (
		\m4_addr_i[31]_pad ,
		_w9103_,
		_w9104_,
		_w20290_
	);
	LUT4 #(
		.INIT('h5d7f)
	) name18390 (
		_w9098_,
		_w9101_,
		_w20289_,
		_w20290_,
		_w20291_
	);
	LUT3 #(
		.INIT('h80)
	) name18391 (
		\m2_addr_i[31]_pad ,
		_w9103_,
		_w9104_,
		_w20292_
	);
	LUT3 #(
		.INIT('h2a)
	) name18392 (
		\m3_addr_i[31]_pad ,
		_w9103_,
		_w9104_,
		_w20293_
	);
	LUT3 #(
		.INIT('h57)
	) name18393 (
		_w9110_,
		_w20292_,
		_w20293_,
		_w20294_
	);
	LUT3 #(
		.INIT('h80)
	) name18394 (
		\m0_addr_i[31]_pad ,
		_w9103_,
		_w9104_,
		_w20295_
	);
	LUT3 #(
		.INIT('h2a)
	) name18395 (
		\m7_addr_i[31]_pad ,
		_w9103_,
		_w9104_,
		_w20296_
	);
	LUT4 #(
		.INIT('h6e7f)
	) name18396 (
		_w9098_,
		_w9101_,
		_w20295_,
		_w20296_,
		_w20297_
	);
	LUT4 #(
		.INIT('h7fff)
	) name18397 (
		_w20288_,
		_w20291_,
		_w20294_,
		_w20297_,
		_w20298_
	);
	LUT3 #(
		.INIT('h2a)
	) name18398 (
		\m3_addr_i[3]_pad ,
		_w9103_,
		_w9104_,
		_w20299_
	);
	LUT3 #(
		.INIT('h80)
	) name18399 (
		\m4_addr_i[3]_pad ,
		_w9103_,
		_w9104_,
		_w20300_
	);
	LUT4 #(
		.INIT('h9dbf)
	) name18400 (
		_w9098_,
		_w9101_,
		_w20299_,
		_w20300_,
		_w20301_
	);
	LUT3 #(
		.INIT('h80)
	) name18401 (
		\m6_addr_i[3]_pad ,
		_w9103_,
		_w9104_,
		_w20302_
	);
	LUT3 #(
		.INIT('h80)
	) name18402 (
		\m2_addr_i[3]_pad ,
		_w9103_,
		_w9104_,
		_w20303_
	);
	LUT4 #(
		.INIT('habef)
	) name18403 (
		_w9098_,
		_w9101_,
		_w20302_,
		_w20303_,
		_w20304_
	);
	LUT3 #(
		.INIT('h2a)
	) name18404 (
		\m5_addr_i[3]_pad ,
		_w9103_,
		_w9104_,
		_w20305_
	);
	LUT3 #(
		.INIT('h2a)
	) name18405 (
		\m1_addr_i[3]_pad ,
		_w9103_,
		_w9104_,
		_w20306_
	);
	LUT4 #(
		.INIT('h57df)
	) name18406 (
		_w9098_,
		_w9101_,
		_w20305_,
		_w20306_,
		_w20307_
	);
	LUT3 #(
		.INIT('h80)
	) name18407 (
		\m0_addr_i[3]_pad ,
		_w9103_,
		_w9104_,
		_w20308_
	);
	LUT3 #(
		.INIT('h2a)
	) name18408 (
		\m7_addr_i[3]_pad ,
		_w9103_,
		_w9104_,
		_w20309_
	);
	LUT4 #(
		.INIT('h6e7f)
	) name18409 (
		_w9098_,
		_w9101_,
		_w20308_,
		_w20309_,
		_w20310_
	);
	LUT4 #(
		.INIT('h7fff)
	) name18410 (
		_w20301_,
		_w20304_,
		_w20307_,
		_w20310_,
		_w20311_
	);
	LUT3 #(
		.INIT('h2a)
	) name18411 (
		\m3_addr_i[4]_pad ,
		_w9103_,
		_w9104_,
		_w20312_
	);
	LUT3 #(
		.INIT('h80)
	) name18412 (
		\m4_addr_i[4]_pad ,
		_w9103_,
		_w9104_,
		_w20313_
	);
	LUT4 #(
		.INIT('h9dbf)
	) name18413 (
		_w9098_,
		_w9101_,
		_w20312_,
		_w20313_,
		_w20314_
	);
	LUT3 #(
		.INIT('h80)
	) name18414 (
		\m6_addr_i[4]_pad ,
		_w9103_,
		_w9104_,
		_w20315_
	);
	LUT3 #(
		.INIT('h80)
	) name18415 (
		\m2_addr_i[4]_pad ,
		_w9103_,
		_w9104_,
		_w20316_
	);
	LUT4 #(
		.INIT('habef)
	) name18416 (
		_w9098_,
		_w9101_,
		_w20315_,
		_w20316_,
		_w20317_
	);
	LUT3 #(
		.INIT('h2a)
	) name18417 (
		\m5_addr_i[4]_pad ,
		_w9103_,
		_w9104_,
		_w20318_
	);
	LUT3 #(
		.INIT('h2a)
	) name18418 (
		\m1_addr_i[4]_pad ,
		_w9103_,
		_w9104_,
		_w20319_
	);
	LUT4 #(
		.INIT('h57df)
	) name18419 (
		_w9098_,
		_w9101_,
		_w20318_,
		_w20319_,
		_w20320_
	);
	LUT3 #(
		.INIT('h80)
	) name18420 (
		\m0_addr_i[4]_pad ,
		_w9103_,
		_w9104_,
		_w20321_
	);
	LUT3 #(
		.INIT('h2a)
	) name18421 (
		\m7_addr_i[4]_pad ,
		_w9103_,
		_w9104_,
		_w20322_
	);
	LUT4 #(
		.INIT('h6e7f)
	) name18422 (
		_w9098_,
		_w9101_,
		_w20321_,
		_w20322_,
		_w20323_
	);
	LUT4 #(
		.INIT('h7fff)
	) name18423 (
		_w20314_,
		_w20317_,
		_w20320_,
		_w20323_,
		_w20324_
	);
	LUT3 #(
		.INIT('h2a)
	) name18424 (
		\m3_addr_i[5]_pad ,
		_w9103_,
		_w9104_,
		_w20325_
	);
	LUT3 #(
		.INIT('h80)
	) name18425 (
		\m4_addr_i[5]_pad ,
		_w9103_,
		_w9104_,
		_w20326_
	);
	LUT4 #(
		.INIT('h9dbf)
	) name18426 (
		_w9098_,
		_w9101_,
		_w20325_,
		_w20326_,
		_w20327_
	);
	LUT3 #(
		.INIT('h80)
	) name18427 (
		\m6_addr_i[5]_pad ,
		_w9103_,
		_w9104_,
		_w20328_
	);
	LUT3 #(
		.INIT('h80)
	) name18428 (
		\m2_addr_i[5]_pad ,
		_w9103_,
		_w9104_,
		_w20329_
	);
	LUT4 #(
		.INIT('habef)
	) name18429 (
		_w9098_,
		_w9101_,
		_w20328_,
		_w20329_,
		_w20330_
	);
	LUT3 #(
		.INIT('h2a)
	) name18430 (
		\m5_addr_i[5]_pad ,
		_w9103_,
		_w9104_,
		_w20331_
	);
	LUT3 #(
		.INIT('h2a)
	) name18431 (
		\m1_addr_i[5]_pad ,
		_w9103_,
		_w9104_,
		_w20332_
	);
	LUT4 #(
		.INIT('h57df)
	) name18432 (
		_w9098_,
		_w9101_,
		_w20331_,
		_w20332_,
		_w20333_
	);
	LUT3 #(
		.INIT('h80)
	) name18433 (
		\m0_addr_i[5]_pad ,
		_w9103_,
		_w9104_,
		_w20334_
	);
	LUT3 #(
		.INIT('h2a)
	) name18434 (
		\m7_addr_i[5]_pad ,
		_w9103_,
		_w9104_,
		_w20335_
	);
	LUT4 #(
		.INIT('h6e7f)
	) name18435 (
		_w9098_,
		_w9101_,
		_w20334_,
		_w20335_,
		_w20336_
	);
	LUT4 #(
		.INIT('h7fff)
	) name18436 (
		_w20327_,
		_w20330_,
		_w20333_,
		_w20336_,
		_w20337_
	);
	LUT3 #(
		.INIT('h2a)
	) name18437 (
		\m3_addr_i[6]_pad ,
		_w9103_,
		_w9104_,
		_w20338_
	);
	LUT3 #(
		.INIT('h80)
	) name18438 (
		\m4_addr_i[6]_pad ,
		_w9103_,
		_w9104_,
		_w20339_
	);
	LUT4 #(
		.INIT('h9dbf)
	) name18439 (
		_w9098_,
		_w9101_,
		_w20338_,
		_w20339_,
		_w20340_
	);
	LUT3 #(
		.INIT('h80)
	) name18440 (
		\m6_addr_i[6]_pad ,
		_w9103_,
		_w9104_,
		_w20341_
	);
	LUT3 #(
		.INIT('h80)
	) name18441 (
		\m2_addr_i[6]_pad ,
		_w9103_,
		_w9104_,
		_w20342_
	);
	LUT4 #(
		.INIT('habef)
	) name18442 (
		_w9098_,
		_w9101_,
		_w20341_,
		_w20342_,
		_w20343_
	);
	LUT3 #(
		.INIT('h2a)
	) name18443 (
		\m5_addr_i[6]_pad ,
		_w9103_,
		_w9104_,
		_w20344_
	);
	LUT3 #(
		.INIT('h2a)
	) name18444 (
		\m1_addr_i[6]_pad ,
		_w9103_,
		_w9104_,
		_w20345_
	);
	LUT4 #(
		.INIT('h57df)
	) name18445 (
		_w9098_,
		_w9101_,
		_w20344_,
		_w20345_,
		_w20346_
	);
	LUT3 #(
		.INIT('h80)
	) name18446 (
		\m0_addr_i[6]_pad ,
		_w9103_,
		_w9104_,
		_w20347_
	);
	LUT3 #(
		.INIT('h2a)
	) name18447 (
		\m7_addr_i[6]_pad ,
		_w9103_,
		_w9104_,
		_w20348_
	);
	LUT4 #(
		.INIT('h6e7f)
	) name18448 (
		_w9098_,
		_w9101_,
		_w20347_,
		_w20348_,
		_w20349_
	);
	LUT4 #(
		.INIT('h7fff)
	) name18449 (
		_w20340_,
		_w20343_,
		_w20346_,
		_w20349_,
		_w20350_
	);
	LUT3 #(
		.INIT('h2a)
	) name18450 (
		\m3_addr_i[7]_pad ,
		_w9103_,
		_w9104_,
		_w20351_
	);
	LUT3 #(
		.INIT('h80)
	) name18451 (
		\m4_addr_i[7]_pad ,
		_w9103_,
		_w9104_,
		_w20352_
	);
	LUT4 #(
		.INIT('h9dbf)
	) name18452 (
		_w9098_,
		_w9101_,
		_w20351_,
		_w20352_,
		_w20353_
	);
	LUT3 #(
		.INIT('h80)
	) name18453 (
		\m6_addr_i[7]_pad ,
		_w9103_,
		_w9104_,
		_w20354_
	);
	LUT3 #(
		.INIT('h80)
	) name18454 (
		\m2_addr_i[7]_pad ,
		_w9103_,
		_w9104_,
		_w20355_
	);
	LUT4 #(
		.INIT('habef)
	) name18455 (
		_w9098_,
		_w9101_,
		_w20354_,
		_w20355_,
		_w20356_
	);
	LUT3 #(
		.INIT('h2a)
	) name18456 (
		\m5_addr_i[7]_pad ,
		_w9103_,
		_w9104_,
		_w20357_
	);
	LUT3 #(
		.INIT('h2a)
	) name18457 (
		\m1_addr_i[7]_pad ,
		_w9103_,
		_w9104_,
		_w20358_
	);
	LUT4 #(
		.INIT('h57df)
	) name18458 (
		_w9098_,
		_w9101_,
		_w20357_,
		_w20358_,
		_w20359_
	);
	LUT3 #(
		.INIT('h80)
	) name18459 (
		\m0_addr_i[7]_pad ,
		_w9103_,
		_w9104_,
		_w20360_
	);
	LUT3 #(
		.INIT('h2a)
	) name18460 (
		\m7_addr_i[7]_pad ,
		_w9103_,
		_w9104_,
		_w20361_
	);
	LUT4 #(
		.INIT('h6e7f)
	) name18461 (
		_w9098_,
		_w9101_,
		_w20360_,
		_w20361_,
		_w20362_
	);
	LUT4 #(
		.INIT('h7fff)
	) name18462 (
		_w20353_,
		_w20356_,
		_w20359_,
		_w20362_,
		_w20363_
	);
	LUT3 #(
		.INIT('h2a)
	) name18463 (
		\m3_addr_i[8]_pad ,
		_w9103_,
		_w9104_,
		_w20364_
	);
	LUT3 #(
		.INIT('h80)
	) name18464 (
		\m4_addr_i[8]_pad ,
		_w9103_,
		_w9104_,
		_w20365_
	);
	LUT4 #(
		.INIT('h9dbf)
	) name18465 (
		_w9098_,
		_w9101_,
		_w20364_,
		_w20365_,
		_w20366_
	);
	LUT3 #(
		.INIT('h80)
	) name18466 (
		\m6_addr_i[8]_pad ,
		_w9103_,
		_w9104_,
		_w20367_
	);
	LUT3 #(
		.INIT('h80)
	) name18467 (
		\m2_addr_i[8]_pad ,
		_w9103_,
		_w9104_,
		_w20368_
	);
	LUT4 #(
		.INIT('habef)
	) name18468 (
		_w9098_,
		_w9101_,
		_w20367_,
		_w20368_,
		_w20369_
	);
	LUT3 #(
		.INIT('h2a)
	) name18469 (
		\m5_addr_i[8]_pad ,
		_w9103_,
		_w9104_,
		_w20370_
	);
	LUT3 #(
		.INIT('h2a)
	) name18470 (
		\m1_addr_i[8]_pad ,
		_w9103_,
		_w9104_,
		_w20371_
	);
	LUT4 #(
		.INIT('h57df)
	) name18471 (
		_w9098_,
		_w9101_,
		_w20370_,
		_w20371_,
		_w20372_
	);
	LUT3 #(
		.INIT('h80)
	) name18472 (
		\m0_addr_i[8]_pad ,
		_w9103_,
		_w9104_,
		_w20373_
	);
	LUT3 #(
		.INIT('h2a)
	) name18473 (
		\m7_addr_i[8]_pad ,
		_w9103_,
		_w9104_,
		_w20374_
	);
	LUT4 #(
		.INIT('h6e7f)
	) name18474 (
		_w9098_,
		_w9101_,
		_w20373_,
		_w20374_,
		_w20375_
	);
	LUT4 #(
		.INIT('h7fff)
	) name18475 (
		_w20366_,
		_w20369_,
		_w20372_,
		_w20375_,
		_w20376_
	);
	LUT3 #(
		.INIT('h2a)
	) name18476 (
		\m3_addr_i[9]_pad ,
		_w9103_,
		_w9104_,
		_w20377_
	);
	LUT3 #(
		.INIT('h80)
	) name18477 (
		\m4_addr_i[9]_pad ,
		_w9103_,
		_w9104_,
		_w20378_
	);
	LUT4 #(
		.INIT('h9dbf)
	) name18478 (
		_w9098_,
		_w9101_,
		_w20377_,
		_w20378_,
		_w20379_
	);
	LUT3 #(
		.INIT('h80)
	) name18479 (
		\m6_addr_i[9]_pad ,
		_w9103_,
		_w9104_,
		_w20380_
	);
	LUT3 #(
		.INIT('h80)
	) name18480 (
		\m2_addr_i[9]_pad ,
		_w9103_,
		_w9104_,
		_w20381_
	);
	LUT4 #(
		.INIT('habef)
	) name18481 (
		_w9098_,
		_w9101_,
		_w20380_,
		_w20381_,
		_w20382_
	);
	LUT3 #(
		.INIT('h2a)
	) name18482 (
		\m5_addr_i[9]_pad ,
		_w9103_,
		_w9104_,
		_w20383_
	);
	LUT3 #(
		.INIT('h2a)
	) name18483 (
		\m1_addr_i[9]_pad ,
		_w9103_,
		_w9104_,
		_w20384_
	);
	LUT4 #(
		.INIT('h57df)
	) name18484 (
		_w9098_,
		_w9101_,
		_w20383_,
		_w20384_,
		_w20385_
	);
	LUT3 #(
		.INIT('h80)
	) name18485 (
		\m0_addr_i[9]_pad ,
		_w9103_,
		_w9104_,
		_w20386_
	);
	LUT3 #(
		.INIT('h2a)
	) name18486 (
		\m7_addr_i[9]_pad ,
		_w9103_,
		_w9104_,
		_w20387_
	);
	LUT4 #(
		.INIT('h6e7f)
	) name18487 (
		_w9098_,
		_w9101_,
		_w20386_,
		_w20387_,
		_w20388_
	);
	LUT4 #(
		.INIT('h7fff)
	) name18488 (
		_w20379_,
		_w20382_,
		_w20385_,
		_w20388_,
		_w20389_
	);
	LUT3 #(
		.INIT('h2a)
	) name18489 (
		\m1_data_i[0]_pad ,
		_w9103_,
		_w9104_,
		_w20390_
	);
	LUT3 #(
		.INIT('h80)
	) name18490 (
		\m2_data_i[0]_pad ,
		_w9103_,
		_w9104_,
		_w20391_
	);
	LUT4 #(
		.INIT('h3b7f)
	) name18491 (
		_w9098_,
		_w9101_,
		_w20390_,
		_w20391_,
		_w20392_
	);
	LUT3 #(
		.INIT('h80)
	) name18492 (
		\m0_data_i[0]_pad ,
		_w9103_,
		_w9104_,
		_w20393_
	);
	LUT3 #(
		.INIT('h80)
	) name18493 (
		\m4_data_i[0]_pad ,
		_w9103_,
		_w9104_,
		_w20394_
	);
	LUT4 #(
		.INIT('h5d7f)
	) name18494 (
		_w9098_,
		_w9101_,
		_w20393_,
		_w20394_,
		_w20395_
	);
	LUT3 #(
		.INIT('h2a)
	) name18495 (
		\m7_data_i[0]_pad ,
		_w9103_,
		_w9104_,
		_w20396_
	);
	LUT3 #(
		.INIT('h2a)
	) name18496 (
		\m3_data_i[0]_pad ,
		_w9103_,
		_w9104_,
		_w20397_
	);
	LUT4 #(
		.INIT('habef)
	) name18497 (
		_w9098_,
		_w9101_,
		_w20396_,
		_w20397_,
		_w20398_
	);
	LUT3 #(
		.INIT('h80)
	) name18498 (
		\m6_data_i[0]_pad ,
		_w9103_,
		_w9104_,
		_w20399_
	);
	LUT3 #(
		.INIT('h2a)
	) name18499 (
		\m5_data_i[0]_pad ,
		_w9103_,
		_w9104_,
		_w20400_
	);
	LUT4 #(
		.INIT('hcdef)
	) name18500 (
		_w9098_,
		_w9101_,
		_w20399_,
		_w20400_,
		_w20401_
	);
	LUT4 #(
		.INIT('h7fff)
	) name18501 (
		_w20392_,
		_w20395_,
		_w20398_,
		_w20401_,
		_w20402_
	);
	LUT3 #(
		.INIT('h80)
	) name18502 (
		\m6_data_i[10]_pad ,
		_w9103_,
		_w9104_,
		_w20403_
	);
	LUT3 #(
		.INIT('h2a)
	) name18503 (
		\m5_data_i[10]_pad ,
		_w9103_,
		_w9104_,
		_w20404_
	);
	LUT4 #(
		.INIT('hcdef)
	) name18504 (
		_w9098_,
		_w9101_,
		_w20403_,
		_w20404_,
		_w20405_
	);
	LUT3 #(
		.INIT('h2a)
	) name18505 (
		\m1_data_i[10]_pad ,
		_w9103_,
		_w9104_,
		_w20406_
	);
	LUT3 #(
		.INIT('h80)
	) name18506 (
		\m4_data_i[10]_pad ,
		_w9103_,
		_w9104_,
		_w20407_
	);
	LUT4 #(
		.INIT('h5d7f)
	) name18507 (
		_w9098_,
		_w9101_,
		_w20406_,
		_w20407_,
		_w20408_
	);
	LUT3 #(
		.INIT('h80)
	) name18508 (
		\m2_data_i[10]_pad ,
		_w9103_,
		_w9104_,
		_w20409_
	);
	LUT3 #(
		.INIT('h2a)
	) name18509 (
		\m3_data_i[10]_pad ,
		_w9103_,
		_w9104_,
		_w20410_
	);
	LUT3 #(
		.INIT('h57)
	) name18510 (
		_w9110_,
		_w20409_,
		_w20410_,
		_w20411_
	);
	LUT3 #(
		.INIT('h80)
	) name18511 (
		\m0_data_i[10]_pad ,
		_w9103_,
		_w9104_,
		_w20412_
	);
	LUT3 #(
		.INIT('h2a)
	) name18512 (
		\m7_data_i[10]_pad ,
		_w9103_,
		_w9104_,
		_w20413_
	);
	LUT4 #(
		.INIT('h6e7f)
	) name18513 (
		_w9098_,
		_w9101_,
		_w20412_,
		_w20413_,
		_w20414_
	);
	LUT4 #(
		.INIT('h7fff)
	) name18514 (
		_w20405_,
		_w20408_,
		_w20411_,
		_w20414_,
		_w20415_
	);
	LUT3 #(
		.INIT('h80)
	) name18515 (
		\m6_data_i[11]_pad ,
		_w9103_,
		_w9104_,
		_w20416_
	);
	LUT3 #(
		.INIT('h2a)
	) name18516 (
		\m5_data_i[11]_pad ,
		_w9103_,
		_w9104_,
		_w20417_
	);
	LUT4 #(
		.INIT('hcdef)
	) name18517 (
		_w9098_,
		_w9101_,
		_w20416_,
		_w20417_,
		_w20418_
	);
	LUT3 #(
		.INIT('h2a)
	) name18518 (
		\m3_data_i[11]_pad ,
		_w9103_,
		_w9104_,
		_w20419_
	);
	LUT3 #(
		.INIT('h80)
	) name18519 (
		\m2_data_i[11]_pad ,
		_w9103_,
		_w9104_,
		_w20420_
	);
	LUT3 #(
		.INIT('h57)
	) name18520 (
		_w9110_,
		_w20419_,
		_w20420_,
		_w20421_
	);
	LUT3 #(
		.INIT('h80)
	) name18521 (
		\m4_data_i[11]_pad ,
		_w9103_,
		_w9104_,
		_w20422_
	);
	LUT3 #(
		.INIT('h2a)
	) name18522 (
		\m1_data_i[11]_pad ,
		_w9103_,
		_w9104_,
		_w20423_
	);
	LUT4 #(
		.INIT('h57df)
	) name18523 (
		_w9098_,
		_w9101_,
		_w20422_,
		_w20423_,
		_w20424_
	);
	LUT3 #(
		.INIT('h80)
	) name18524 (
		\m0_data_i[11]_pad ,
		_w9103_,
		_w9104_,
		_w20425_
	);
	LUT3 #(
		.INIT('h2a)
	) name18525 (
		\m7_data_i[11]_pad ,
		_w9103_,
		_w9104_,
		_w20426_
	);
	LUT4 #(
		.INIT('h6e7f)
	) name18526 (
		_w9098_,
		_w9101_,
		_w20425_,
		_w20426_,
		_w20427_
	);
	LUT4 #(
		.INIT('h7fff)
	) name18527 (
		_w20418_,
		_w20421_,
		_w20424_,
		_w20427_,
		_w20428_
	);
	LUT3 #(
		.INIT('h80)
	) name18528 (
		\m0_data_i[12]_pad ,
		_w9103_,
		_w9104_,
		_w20429_
	);
	LUT3 #(
		.INIT('h2a)
	) name18529 (
		\m7_data_i[12]_pad ,
		_w9103_,
		_w9104_,
		_w20430_
	);
	LUT4 #(
		.INIT('h6e7f)
	) name18530 (
		_w9098_,
		_w9101_,
		_w20429_,
		_w20430_,
		_w20431_
	);
	LUT3 #(
		.INIT('h80)
	) name18531 (
		\m6_data_i[12]_pad ,
		_w9103_,
		_w9104_,
		_w20432_
	);
	LUT3 #(
		.INIT('h80)
	) name18532 (
		\m4_data_i[12]_pad ,
		_w9103_,
		_w9104_,
		_w20433_
	);
	LUT4 #(
		.INIT('hcdef)
	) name18533 (
		_w9098_,
		_w9101_,
		_w20432_,
		_w20433_,
		_w20434_
	);
	LUT3 #(
		.INIT('h2a)
	) name18534 (
		\m5_data_i[12]_pad ,
		_w9103_,
		_w9104_,
		_w20435_
	);
	LUT3 #(
		.INIT('h2a)
	) name18535 (
		\m3_data_i[12]_pad ,
		_w9103_,
		_w9104_,
		_w20436_
	);
	LUT4 #(
		.INIT('h9bdf)
	) name18536 (
		_w9098_,
		_w9101_,
		_w20435_,
		_w20436_,
		_w20437_
	);
	LUT3 #(
		.INIT('h2a)
	) name18537 (
		\m1_data_i[12]_pad ,
		_w9103_,
		_w9104_,
		_w20438_
	);
	LUT3 #(
		.INIT('h80)
	) name18538 (
		\m2_data_i[12]_pad ,
		_w9103_,
		_w9104_,
		_w20439_
	);
	LUT4 #(
		.INIT('h3b7f)
	) name18539 (
		_w9098_,
		_w9101_,
		_w20438_,
		_w20439_,
		_w20440_
	);
	LUT4 #(
		.INIT('h7fff)
	) name18540 (
		_w20431_,
		_w20434_,
		_w20437_,
		_w20440_,
		_w20441_
	);
	LUT3 #(
		.INIT('h2a)
	) name18541 (
		\m3_data_i[13]_pad ,
		_w9103_,
		_w9104_,
		_w20442_
	);
	LUT3 #(
		.INIT('h80)
	) name18542 (
		\m4_data_i[13]_pad ,
		_w9103_,
		_w9104_,
		_w20443_
	);
	LUT4 #(
		.INIT('h9dbf)
	) name18543 (
		_w9098_,
		_w9101_,
		_w20442_,
		_w20443_,
		_w20444_
	);
	LUT3 #(
		.INIT('h80)
	) name18544 (
		\m0_data_i[13]_pad ,
		_w9103_,
		_w9104_,
		_w20445_
	);
	LUT3 #(
		.INIT('h2a)
	) name18545 (
		\m5_data_i[13]_pad ,
		_w9103_,
		_w9104_,
		_w20446_
	);
	LUT4 #(
		.INIT('h5d7f)
	) name18546 (
		_w9098_,
		_w9101_,
		_w20445_,
		_w20446_,
		_w20447_
	);
	LUT3 #(
		.INIT('h2a)
	) name18547 (
		\m7_data_i[13]_pad ,
		_w9103_,
		_w9104_,
		_w20448_
	);
	LUT3 #(
		.INIT('h80)
	) name18548 (
		\m6_data_i[13]_pad ,
		_w9103_,
		_w9104_,
		_w20449_
	);
	LUT3 #(
		.INIT('h57)
	) name18549 (
		_w9102_,
		_w20448_,
		_w20449_,
		_w20450_
	);
	LUT3 #(
		.INIT('h2a)
	) name18550 (
		\m1_data_i[13]_pad ,
		_w9103_,
		_w9104_,
		_w20451_
	);
	LUT3 #(
		.INIT('h80)
	) name18551 (
		\m2_data_i[13]_pad ,
		_w9103_,
		_w9104_,
		_w20452_
	);
	LUT4 #(
		.INIT('h3b7f)
	) name18552 (
		_w9098_,
		_w9101_,
		_w20451_,
		_w20452_,
		_w20453_
	);
	LUT4 #(
		.INIT('h7fff)
	) name18553 (
		_w20444_,
		_w20447_,
		_w20450_,
		_w20453_,
		_w20454_
	);
	LUT3 #(
		.INIT('h80)
	) name18554 (
		\m6_data_i[14]_pad ,
		_w9103_,
		_w9104_,
		_w20455_
	);
	LUT3 #(
		.INIT('h2a)
	) name18555 (
		\m5_data_i[14]_pad ,
		_w9103_,
		_w9104_,
		_w20456_
	);
	LUT4 #(
		.INIT('hcdef)
	) name18556 (
		_w9098_,
		_w9101_,
		_w20455_,
		_w20456_,
		_w20457_
	);
	LUT3 #(
		.INIT('h2a)
	) name18557 (
		\m1_data_i[14]_pad ,
		_w9103_,
		_w9104_,
		_w20458_
	);
	LUT3 #(
		.INIT('h80)
	) name18558 (
		\m4_data_i[14]_pad ,
		_w9103_,
		_w9104_,
		_w20459_
	);
	LUT4 #(
		.INIT('h5d7f)
	) name18559 (
		_w9098_,
		_w9101_,
		_w20458_,
		_w20459_,
		_w20460_
	);
	LUT3 #(
		.INIT('h80)
	) name18560 (
		\m2_data_i[14]_pad ,
		_w9103_,
		_w9104_,
		_w20461_
	);
	LUT3 #(
		.INIT('h2a)
	) name18561 (
		\m3_data_i[14]_pad ,
		_w9103_,
		_w9104_,
		_w20462_
	);
	LUT3 #(
		.INIT('h57)
	) name18562 (
		_w9110_,
		_w20461_,
		_w20462_,
		_w20463_
	);
	LUT3 #(
		.INIT('h80)
	) name18563 (
		\m0_data_i[14]_pad ,
		_w9103_,
		_w9104_,
		_w20464_
	);
	LUT3 #(
		.INIT('h2a)
	) name18564 (
		\m7_data_i[14]_pad ,
		_w9103_,
		_w9104_,
		_w20465_
	);
	LUT4 #(
		.INIT('h6e7f)
	) name18565 (
		_w9098_,
		_w9101_,
		_w20464_,
		_w20465_,
		_w20466_
	);
	LUT4 #(
		.INIT('h7fff)
	) name18566 (
		_w20457_,
		_w20460_,
		_w20463_,
		_w20466_,
		_w20467_
	);
	LUT3 #(
		.INIT('h2a)
	) name18567 (
		\m3_data_i[15]_pad ,
		_w9103_,
		_w9104_,
		_w20468_
	);
	LUT3 #(
		.INIT('h80)
	) name18568 (
		\m4_data_i[15]_pad ,
		_w9103_,
		_w9104_,
		_w20469_
	);
	LUT4 #(
		.INIT('h9dbf)
	) name18569 (
		_w9098_,
		_w9101_,
		_w20468_,
		_w20469_,
		_w20470_
	);
	LUT3 #(
		.INIT('h80)
	) name18570 (
		\m0_data_i[15]_pad ,
		_w9103_,
		_w9104_,
		_w20471_
	);
	LUT3 #(
		.INIT('h80)
	) name18571 (
		\m2_data_i[15]_pad ,
		_w9103_,
		_w9104_,
		_w20472_
	);
	LUT4 #(
		.INIT('h3b7f)
	) name18572 (
		_w9098_,
		_w9101_,
		_w20471_,
		_w20472_,
		_w20473_
	);
	LUT3 #(
		.INIT('h2a)
	) name18573 (
		\m7_data_i[15]_pad ,
		_w9103_,
		_w9104_,
		_w20474_
	);
	LUT3 #(
		.INIT('h2a)
	) name18574 (
		\m1_data_i[15]_pad ,
		_w9103_,
		_w9104_,
		_w20475_
	);
	LUT4 #(
		.INIT('h67ef)
	) name18575 (
		_w9098_,
		_w9101_,
		_w20474_,
		_w20475_,
		_w20476_
	);
	LUT3 #(
		.INIT('h80)
	) name18576 (
		\m6_data_i[15]_pad ,
		_w9103_,
		_w9104_,
		_w20477_
	);
	LUT3 #(
		.INIT('h2a)
	) name18577 (
		\m5_data_i[15]_pad ,
		_w9103_,
		_w9104_,
		_w20478_
	);
	LUT4 #(
		.INIT('hcdef)
	) name18578 (
		_w9098_,
		_w9101_,
		_w20477_,
		_w20478_,
		_w20479_
	);
	LUT4 #(
		.INIT('h7fff)
	) name18579 (
		_w20470_,
		_w20473_,
		_w20476_,
		_w20479_,
		_w20480_
	);
	LUT3 #(
		.INIT('h2a)
	) name18580 (
		\m1_data_i[16]_pad ,
		_w9103_,
		_w9104_,
		_w20481_
	);
	LUT3 #(
		.INIT('h80)
	) name18581 (
		\m2_data_i[16]_pad ,
		_w9103_,
		_w9104_,
		_w20482_
	);
	LUT4 #(
		.INIT('h3b7f)
	) name18582 (
		_w9098_,
		_w9101_,
		_w20481_,
		_w20482_,
		_w20483_
	);
	LUT3 #(
		.INIT('h80)
	) name18583 (
		\m0_data_i[16]_pad ,
		_w9103_,
		_w9104_,
		_w20484_
	);
	LUT3 #(
		.INIT('h2a)
	) name18584 (
		\m5_data_i[16]_pad ,
		_w9103_,
		_w9104_,
		_w20485_
	);
	LUT4 #(
		.INIT('h5d7f)
	) name18585 (
		_w9098_,
		_w9101_,
		_w20484_,
		_w20485_,
		_w20486_
	);
	LUT3 #(
		.INIT('h2a)
	) name18586 (
		\m7_data_i[16]_pad ,
		_w9103_,
		_w9104_,
		_w20487_
	);
	LUT3 #(
		.INIT('h80)
	) name18587 (
		\m6_data_i[16]_pad ,
		_w9103_,
		_w9104_,
		_w20488_
	);
	LUT3 #(
		.INIT('h57)
	) name18588 (
		_w9102_,
		_w20487_,
		_w20488_,
		_w20489_
	);
	LUT3 #(
		.INIT('h2a)
	) name18589 (
		\m3_data_i[16]_pad ,
		_w9103_,
		_w9104_,
		_w20490_
	);
	LUT3 #(
		.INIT('h80)
	) name18590 (
		\m4_data_i[16]_pad ,
		_w9103_,
		_w9104_,
		_w20491_
	);
	LUT4 #(
		.INIT('h9dbf)
	) name18591 (
		_w9098_,
		_w9101_,
		_w20490_,
		_w20491_,
		_w20492_
	);
	LUT4 #(
		.INIT('h7fff)
	) name18592 (
		_w20483_,
		_w20486_,
		_w20489_,
		_w20492_,
		_w20493_
	);
	LUT3 #(
		.INIT('h2a)
	) name18593 (
		\m3_data_i[17]_pad ,
		_w9103_,
		_w9104_,
		_w20494_
	);
	LUT3 #(
		.INIT('h80)
	) name18594 (
		\m4_data_i[17]_pad ,
		_w9103_,
		_w9104_,
		_w20495_
	);
	LUT4 #(
		.INIT('h9dbf)
	) name18595 (
		_w9098_,
		_w9101_,
		_w20494_,
		_w20495_,
		_w20496_
	);
	LUT3 #(
		.INIT('h80)
	) name18596 (
		\m0_data_i[17]_pad ,
		_w9103_,
		_w9104_,
		_w20497_
	);
	LUT3 #(
		.INIT('h80)
	) name18597 (
		\m2_data_i[17]_pad ,
		_w9103_,
		_w9104_,
		_w20498_
	);
	LUT4 #(
		.INIT('h3b7f)
	) name18598 (
		_w9098_,
		_w9101_,
		_w20497_,
		_w20498_,
		_w20499_
	);
	LUT3 #(
		.INIT('h2a)
	) name18599 (
		\m7_data_i[17]_pad ,
		_w9103_,
		_w9104_,
		_w20500_
	);
	LUT3 #(
		.INIT('h2a)
	) name18600 (
		\m1_data_i[17]_pad ,
		_w9103_,
		_w9104_,
		_w20501_
	);
	LUT4 #(
		.INIT('h67ef)
	) name18601 (
		_w9098_,
		_w9101_,
		_w20500_,
		_w20501_,
		_w20502_
	);
	LUT3 #(
		.INIT('h80)
	) name18602 (
		\m6_data_i[17]_pad ,
		_w9103_,
		_w9104_,
		_w20503_
	);
	LUT3 #(
		.INIT('h2a)
	) name18603 (
		\m5_data_i[17]_pad ,
		_w9103_,
		_w9104_,
		_w20504_
	);
	LUT4 #(
		.INIT('hcdef)
	) name18604 (
		_w9098_,
		_w9101_,
		_w20503_,
		_w20504_,
		_w20505_
	);
	LUT4 #(
		.INIT('h7fff)
	) name18605 (
		_w20496_,
		_w20499_,
		_w20502_,
		_w20505_,
		_w20506_
	);
	LUT3 #(
		.INIT('h2a)
	) name18606 (
		\m3_data_i[18]_pad ,
		_w9103_,
		_w9104_,
		_w20507_
	);
	LUT3 #(
		.INIT('h80)
	) name18607 (
		\m4_data_i[18]_pad ,
		_w9103_,
		_w9104_,
		_w20508_
	);
	LUT4 #(
		.INIT('h9dbf)
	) name18608 (
		_w9098_,
		_w9101_,
		_w20507_,
		_w20508_,
		_w20509_
	);
	LUT3 #(
		.INIT('h80)
	) name18609 (
		\m0_data_i[18]_pad ,
		_w9103_,
		_w9104_,
		_w20510_
	);
	LUT3 #(
		.INIT('h80)
	) name18610 (
		\m2_data_i[18]_pad ,
		_w9103_,
		_w9104_,
		_w20511_
	);
	LUT4 #(
		.INIT('h3b7f)
	) name18611 (
		_w9098_,
		_w9101_,
		_w20510_,
		_w20511_,
		_w20512_
	);
	LUT3 #(
		.INIT('h2a)
	) name18612 (
		\m7_data_i[18]_pad ,
		_w9103_,
		_w9104_,
		_w20513_
	);
	LUT3 #(
		.INIT('h2a)
	) name18613 (
		\m1_data_i[18]_pad ,
		_w9103_,
		_w9104_,
		_w20514_
	);
	LUT4 #(
		.INIT('h67ef)
	) name18614 (
		_w9098_,
		_w9101_,
		_w20513_,
		_w20514_,
		_w20515_
	);
	LUT3 #(
		.INIT('h80)
	) name18615 (
		\m6_data_i[18]_pad ,
		_w9103_,
		_w9104_,
		_w20516_
	);
	LUT3 #(
		.INIT('h2a)
	) name18616 (
		\m5_data_i[18]_pad ,
		_w9103_,
		_w9104_,
		_w20517_
	);
	LUT4 #(
		.INIT('hcdef)
	) name18617 (
		_w9098_,
		_w9101_,
		_w20516_,
		_w20517_,
		_w20518_
	);
	LUT4 #(
		.INIT('h7fff)
	) name18618 (
		_w20509_,
		_w20512_,
		_w20515_,
		_w20518_,
		_w20519_
	);
	LUT3 #(
		.INIT('h2a)
	) name18619 (
		\m3_data_i[19]_pad ,
		_w9103_,
		_w9104_,
		_w20520_
	);
	LUT3 #(
		.INIT('h80)
	) name18620 (
		\m4_data_i[19]_pad ,
		_w9103_,
		_w9104_,
		_w20521_
	);
	LUT4 #(
		.INIT('h9dbf)
	) name18621 (
		_w9098_,
		_w9101_,
		_w20520_,
		_w20521_,
		_w20522_
	);
	LUT3 #(
		.INIT('h80)
	) name18622 (
		\m6_data_i[19]_pad ,
		_w9103_,
		_w9104_,
		_w20523_
	);
	LUT3 #(
		.INIT('h80)
	) name18623 (
		\m2_data_i[19]_pad ,
		_w9103_,
		_w9104_,
		_w20524_
	);
	LUT4 #(
		.INIT('habef)
	) name18624 (
		_w9098_,
		_w9101_,
		_w20523_,
		_w20524_,
		_w20525_
	);
	LUT3 #(
		.INIT('h2a)
	) name18625 (
		\m5_data_i[19]_pad ,
		_w9103_,
		_w9104_,
		_w20526_
	);
	LUT3 #(
		.INIT('h2a)
	) name18626 (
		\m1_data_i[19]_pad ,
		_w9103_,
		_w9104_,
		_w20527_
	);
	LUT4 #(
		.INIT('h57df)
	) name18627 (
		_w9098_,
		_w9101_,
		_w20526_,
		_w20527_,
		_w20528_
	);
	LUT3 #(
		.INIT('h80)
	) name18628 (
		\m0_data_i[19]_pad ,
		_w9103_,
		_w9104_,
		_w20529_
	);
	LUT3 #(
		.INIT('h2a)
	) name18629 (
		\m7_data_i[19]_pad ,
		_w9103_,
		_w9104_,
		_w20530_
	);
	LUT4 #(
		.INIT('h6e7f)
	) name18630 (
		_w9098_,
		_w9101_,
		_w20529_,
		_w20530_,
		_w20531_
	);
	LUT4 #(
		.INIT('h7fff)
	) name18631 (
		_w20522_,
		_w20525_,
		_w20528_,
		_w20531_,
		_w20532_
	);
	LUT3 #(
		.INIT('h2a)
	) name18632 (
		\m3_data_i[1]_pad ,
		_w9103_,
		_w9104_,
		_w20533_
	);
	LUT3 #(
		.INIT('h80)
	) name18633 (
		\m4_data_i[1]_pad ,
		_w9103_,
		_w9104_,
		_w20534_
	);
	LUT4 #(
		.INIT('h9dbf)
	) name18634 (
		_w9098_,
		_w9101_,
		_w20533_,
		_w20534_,
		_w20535_
	);
	LUT3 #(
		.INIT('h2a)
	) name18635 (
		\m1_data_i[1]_pad ,
		_w9103_,
		_w9104_,
		_w20536_
	);
	LUT3 #(
		.INIT('h2a)
	) name18636 (
		\m5_data_i[1]_pad ,
		_w9103_,
		_w9104_,
		_w20537_
	);
	LUT4 #(
		.INIT('h5d7f)
	) name18637 (
		_w9098_,
		_w9101_,
		_w20536_,
		_w20537_,
		_w20538_
	);
	LUT3 #(
		.INIT('h80)
	) name18638 (
		\m2_data_i[1]_pad ,
		_w9103_,
		_w9104_,
		_w20539_
	);
	LUT3 #(
		.INIT('h80)
	) name18639 (
		\m6_data_i[1]_pad ,
		_w9103_,
		_w9104_,
		_w20540_
	);
	LUT4 #(
		.INIT('haebf)
	) name18640 (
		_w9098_,
		_w9101_,
		_w20539_,
		_w20540_,
		_w20541_
	);
	LUT3 #(
		.INIT('h80)
	) name18641 (
		\m0_data_i[1]_pad ,
		_w9103_,
		_w9104_,
		_w20542_
	);
	LUT3 #(
		.INIT('h2a)
	) name18642 (
		\m7_data_i[1]_pad ,
		_w9103_,
		_w9104_,
		_w20543_
	);
	LUT4 #(
		.INIT('h6e7f)
	) name18643 (
		_w9098_,
		_w9101_,
		_w20542_,
		_w20543_,
		_w20544_
	);
	LUT4 #(
		.INIT('h7fff)
	) name18644 (
		_w20535_,
		_w20538_,
		_w20541_,
		_w20544_,
		_w20545_
	);
	LUT3 #(
		.INIT('h2a)
	) name18645 (
		\m3_data_i[20]_pad ,
		_w9103_,
		_w9104_,
		_w20546_
	);
	LUT3 #(
		.INIT('h80)
	) name18646 (
		\m4_data_i[20]_pad ,
		_w9103_,
		_w9104_,
		_w20547_
	);
	LUT4 #(
		.INIT('h9dbf)
	) name18647 (
		_w9098_,
		_w9101_,
		_w20546_,
		_w20547_,
		_w20548_
	);
	LUT3 #(
		.INIT('h2a)
	) name18648 (
		\m1_data_i[20]_pad ,
		_w9103_,
		_w9104_,
		_w20549_
	);
	LUT3 #(
		.INIT('h2a)
	) name18649 (
		\m5_data_i[20]_pad ,
		_w9103_,
		_w9104_,
		_w20550_
	);
	LUT4 #(
		.INIT('h5d7f)
	) name18650 (
		_w9098_,
		_w9101_,
		_w20549_,
		_w20550_,
		_w20551_
	);
	LUT3 #(
		.INIT('h80)
	) name18651 (
		\m2_data_i[20]_pad ,
		_w9103_,
		_w9104_,
		_w20552_
	);
	LUT3 #(
		.INIT('h80)
	) name18652 (
		\m6_data_i[20]_pad ,
		_w9103_,
		_w9104_,
		_w20553_
	);
	LUT4 #(
		.INIT('haebf)
	) name18653 (
		_w9098_,
		_w9101_,
		_w20552_,
		_w20553_,
		_w20554_
	);
	LUT3 #(
		.INIT('h80)
	) name18654 (
		\m0_data_i[20]_pad ,
		_w9103_,
		_w9104_,
		_w20555_
	);
	LUT3 #(
		.INIT('h2a)
	) name18655 (
		\m7_data_i[20]_pad ,
		_w9103_,
		_w9104_,
		_w20556_
	);
	LUT4 #(
		.INIT('h6e7f)
	) name18656 (
		_w9098_,
		_w9101_,
		_w20555_,
		_w20556_,
		_w20557_
	);
	LUT4 #(
		.INIT('h7fff)
	) name18657 (
		_w20548_,
		_w20551_,
		_w20554_,
		_w20557_,
		_w20558_
	);
	LUT3 #(
		.INIT('h80)
	) name18658 (
		\m6_data_i[21]_pad ,
		_w9103_,
		_w9104_,
		_w20559_
	);
	LUT3 #(
		.INIT('h2a)
	) name18659 (
		\m5_data_i[21]_pad ,
		_w9103_,
		_w9104_,
		_w20560_
	);
	LUT4 #(
		.INIT('hcdef)
	) name18660 (
		_w9098_,
		_w9101_,
		_w20559_,
		_w20560_,
		_w20561_
	);
	LUT3 #(
		.INIT('h80)
	) name18661 (
		\m0_data_i[21]_pad ,
		_w9103_,
		_w9104_,
		_w20562_
	);
	LUT3 #(
		.INIT('h80)
	) name18662 (
		\m4_data_i[21]_pad ,
		_w9103_,
		_w9104_,
		_w20563_
	);
	LUT4 #(
		.INIT('h5d7f)
	) name18663 (
		_w9098_,
		_w9101_,
		_w20562_,
		_w20563_,
		_w20564_
	);
	LUT3 #(
		.INIT('h2a)
	) name18664 (
		\m7_data_i[21]_pad ,
		_w9103_,
		_w9104_,
		_w20565_
	);
	LUT3 #(
		.INIT('h2a)
	) name18665 (
		\m3_data_i[21]_pad ,
		_w9103_,
		_w9104_,
		_w20566_
	);
	LUT4 #(
		.INIT('habef)
	) name18666 (
		_w9098_,
		_w9101_,
		_w20565_,
		_w20566_,
		_w20567_
	);
	LUT3 #(
		.INIT('h2a)
	) name18667 (
		\m1_data_i[21]_pad ,
		_w9103_,
		_w9104_,
		_w20568_
	);
	LUT3 #(
		.INIT('h80)
	) name18668 (
		\m2_data_i[21]_pad ,
		_w9103_,
		_w9104_,
		_w20569_
	);
	LUT4 #(
		.INIT('h3b7f)
	) name18669 (
		_w9098_,
		_w9101_,
		_w20568_,
		_w20569_,
		_w20570_
	);
	LUT4 #(
		.INIT('h7fff)
	) name18670 (
		_w20561_,
		_w20564_,
		_w20567_,
		_w20570_,
		_w20571_
	);
	LUT3 #(
		.INIT('h2a)
	) name18671 (
		\m3_data_i[22]_pad ,
		_w9103_,
		_w9104_,
		_w20572_
	);
	LUT3 #(
		.INIT('h80)
	) name18672 (
		\m4_data_i[22]_pad ,
		_w9103_,
		_w9104_,
		_w20573_
	);
	LUT4 #(
		.INIT('h9dbf)
	) name18673 (
		_w9098_,
		_w9101_,
		_w20572_,
		_w20573_,
		_w20574_
	);
	LUT3 #(
		.INIT('h80)
	) name18674 (
		\m6_data_i[22]_pad ,
		_w9103_,
		_w9104_,
		_w20575_
	);
	LUT3 #(
		.INIT('h80)
	) name18675 (
		\m2_data_i[22]_pad ,
		_w9103_,
		_w9104_,
		_w20576_
	);
	LUT4 #(
		.INIT('habef)
	) name18676 (
		_w9098_,
		_w9101_,
		_w20575_,
		_w20576_,
		_w20577_
	);
	LUT3 #(
		.INIT('h2a)
	) name18677 (
		\m5_data_i[22]_pad ,
		_w9103_,
		_w9104_,
		_w20578_
	);
	LUT3 #(
		.INIT('h2a)
	) name18678 (
		\m1_data_i[22]_pad ,
		_w9103_,
		_w9104_,
		_w20579_
	);
	LUT4 #(
		.INIT('h57df)
	) name18679 (
		_w9098_,
		_w9101_,
		_w20578_,
		_w20579_,
		_w20580_
	);
	LUT3 #(
		.INIT('h80)
	) name18680 (
		\m0_data_i[22]_pad ,
		_w9103_,
		_w9104_,
		_w20581_
	);
	LUT3 #(
		.INIT('h2a)
	) name18681 (
		\m7_data_i[22]_pad ,
		_w9103_,
		_w9104_,
		_w20582_
	);
	LUT4 #(
		.INIT('h6e7f)
	) name18682 (
		_w9098_,
		_w9101_,
		_w20581_,
		_w20582_,
		_w20583_
	);
	LUT4 #(
		.INIT('h7fff)
	) name18683 (
		_w20574_,
		_w20577_,
		_w20580_,
		_w20583_,
		_w20584_
	);
	LUT3 #(
		.INIT('h80)
	) name18684 (
		\m0_data_i[23]_pad ,
		_w9103_,
		_w9104_,
		_w20585_
	);
	LUT3 #(
		.INIT('h2a)
	) name18685 (
		\m7_data_i[23]_pad ,
		_w9103_,
		_w9104_,
		_w20586_
	);
	LUT4 #(
		.INIT('h6e7f)
	) name18686 (
		_w9098_,
		_w9101_,
		_w20585_,
		_w20586_,
		_w20587_
	);
	LUT3 #(
		.INIT('h2a)
	) name18687 (
		\m1_data_i[23]_pad ,
		_w9103_,
		_w9104_,
		_w20588_
	);
	LUT3 #(
		.INIT('h2a)
	) name18688 (
		\m5_data_i[23]_pad ,
		_w9103_,
		_w9104_,
		_w20589_
	);
	LUT4 #(
		.INIT('h5d7f)
	) name18689 (
		_w9098_,
		_w9101_,
		_w20588_,
		_w20589_,
		_w20590_
	);
	LUT3 #(
		.INIT('h80)
	) name18690 (
		\m2_data_i[23]_pad ,
		_w9103_,
		_w9104_,
		_w20591_
	);
	LUT3 #(
		.INIT('h80)
	) name18691 (
		\m6_data_i[23]_pad ,
		_w9103_,
		_w9104_,
		_w20592_
	);
	LUT4 #(
		.INIT('haebf)
	) name18692 (
		_w9098_,
		_w9101_,
		_w20591_,
		_w20592_,
		_w20593_
	);
	LUT3 #(
		.INIT('h2a)
	) name18693 (
		\m3_data_i[23]_pad ,
		_w9103_,
		_w9104_,
		_w20594_
	);
	LUT3 #(
		.INIT('h80)
	) name18694 (
		\m4_data_i[23]_pad ,
		_w9103_,
		_w9104_,
		_w20595_
	);
	LUT4 #(
		.INIT('h9dbf)
	) name18695 (
		_w9098_,
		_w9101_,
		_w20594_,
		_w20595_,
		_w20596_
	);
	LUT4 #(
		.INIT('h7fff)
	) name18696 (
		_w20587_,
		_w20590_,
		_w20593_,
		_w20596_,
		_w20597_
	);
	LUT3 #(
		.INIT('h2a)
	) name18697 (
		\m1_data_i[24]_pad ,
		_w9103_,
		_w9104_,
		_w20598_
	);
	LUT3 #(
		.INIT('h80)
	) name18698 (
		\m2_data_i[24]_pad ,
		_w9103_,
		_w9104_,
		_w20599_
	);
	LUT4 #(
		.INIT('h3b7f)
	) name18699 (
		_w9098_,
		_w9101_,
		_w20598_,
		_w20599_,
		_w20600_
	);
	LUT3 #(
		.INIT('h80)
	) name18700 (
		\m6_data_i[24]_pad ,
		_w9103_,
		_w9104_,
		_w20601_
	);
	LUT3 #(
		.INIT('h80)
	) name18701 (
		\m4_data_i[24]_pad ,
		_w9103_,
		_w9104_,
		_w20602_
	);
	LUT4 #(
		.INIT('hcdef)
	) name18702 (
		_w9098_,
		_w9101_,
		_w20601_,
		_w20602_,
		_w20603_
	);
	LUT3 #(
		.INIT('h2a)
	) name18703 (
		\m5_data_i[24]_pad ,
		_w9103_,
		_w9104_,
		_w20604_
	);
	LUT3 #(
		.INIT('h2a)
	) name18704 (
		\m3_data_i[24]_pad ,
		_w9103_,
		_w9104_,
		_w20605_
	);
	LUT4 #(
		.INIT('h9bdf)
	) name18705 (
		_w9098_,
		_w9101_,
		_w20604_,
		_w20605_,
		_w20606_
	);
	LUT3 #(
		.INIT('h80)
	) name18706 (
		\m0_data_i[24]_pad ,
		_w9103_,
		_w9104_,
		_w20607_
	);
	LUT3 #(
		.INIT('h2a)
	) name18707 (
		\m7_data_i[24]_pad ,
		_w9103_,
		_w9104_,
		_w20608_
	);
	LUT4 #(
		.INIT('h6e7f)
	) name18708 (
		_w9098_,
		_w9101_,
		_w20607_,
		_w20608_,
		_w20609_
	);
	LUT4 #(
		.INIT('h7fff)
	) name18709 (
		_w20600_,
		_w20603_,
		_w20606_,
		_w20609_,
		_w20610_
	);
	LUT3 #(
		.INIT('h80)
	) name18710 (
		\m6_data_i[25]_pad ,
		_w9103_,
		_w9104_,
		_w20611_
	);
	LUT3 #(
		.INIT('h2a)
	) name18711 (
		\m5_data_i[25]_pad ,
		_w9103_,
		_w9104_,
		_w20612_
	);
	LUT4 #(
		.INIT('hcdef)
	) name18712 (
		_w9098_,
		_w9101_,
		_w20611_,
		_w20612_,
		_w20613_
	);
	LUT3 #(
		.INIT('h80)
	) name18713 (
		\m0_data_i[25]_pad ,
		_w9103_,
		_w9104_,
		_w20614_
	);
	LUT3 #(
		.INIT('h80)
	) name18714 (
		\m4_data_i[25]_pad ,
		_w9103_,
		_w9104_,
		_w20615_
	);
	LUT4 #(
		.INIT('h5d7f)
	) name18715 (
		_w9098_,
		_w9101_,
		_w20614_,
		_w20615_,
		_w20616_
	);
	LUT3 #(
		.INIT('h2a)
	) name18716 (
		\m7_data_i[25]_pad ,
		_w9103_,
		_w9104_,
		_w20617_
	);
	LUT3 #(
		.INIT('h2a)
	) name18717 (
		\m3_data_i[25]_pad ,
		_w9103_,
		_w9104_,
		_w20618_
	);
	LUT4 #(
		.INIT('habef)
	) name18718 (
		_w9098_,
		_w9101_,
		_w20617_,
		_w20618_,
		_w20619_
	);
	LUT3 #(
		.INIT('h2a)
	) name18719 (
		\m1_data_i[25]_pad ,
		_w9103_,
		_w9104_,
		_w20620_
	);
	LUT3 #(
		.INIT('h80)
	) name18720 (
		\m2_data_i[25]_pad ,
		_w9103_,
		_w9104_,
		_w20621_
	);
	LUT4 #(
		.INIT('h3b7f)
	) name18721 (
		_w9098_,
		_w9101_,
		_w20620_,
		_w20621_,
		_w20622_
	);
	LUT4 #(
		.INIT('h7fff)
	) name18722 (
		_w20613_,
		_w20616_,
		_w20619_,
		_w20622_,
		_w20623_
	);
	LUT3 #(
		.INIT('h2a)
	) name18723 (
		\m1_data_i[26]_pad ,
		_w9103_,
		_w9104_,
		_w20624_
	);
	LUT3 #(
		.INIT('h80)
	) name18724 (
		\m2_data_i[26]_pad ,
		_w9103_,
		_w9104_,
		_w20625_
	);
	LUT4 #(
		.INIT('h3b7f)
	) name18725 (
		_w9098_,
		_w9101_,
		_w20624_,
		_w20625_,
		_w20626_
	);
	LUT3 #(
		.INIT('h2a)
	) name18726 (
		\m3_data_i[26]_pad ,
		_w9103_,
		_w9104_,
		_w20627_
	);
	LUT3 #(
		.INIT('h2a)
	) name18727 (
		\m5_data_i[26]_pad ,
		_w9103_,
		_w9104_,
		_w20628_
	);
	LUT4 #(
		.INIT('h9dbf)
	) name18728 (
		_w9098_,
		_w9101_,
		_w20627_,
		_w20628_,
		_w20629_
	);
	LUT3 #(
		.INIT('h80)
	) name18729 (
		\m4_data_i[26]_pad ,
		_w9103_,
		_w9104_,
		_w20630_
	);
	LUT3 #(
		.INIT('h80)
	) name18730 (
		\m6_data_i[26]_pad ,
		_w9103_,
		_w9104_,
		_w20631_
	);
	LUT4 #(
		.INIT('hcedf)
	) name18731 (
		_w9098_,
		_w9101_,
		_w20630_,
		_w20631_,
		_w20632_
	);
	LUT3 #(
		.INIT('h80)
	) name18732 (
		\m0_data_i[26]_pad ,
		_w9103_,
		_w9104_,
		_w20633_
	);
	LUT3 #(
		.INIT('h2a)
	) name18733 (
		\m7_data_i[26]_pad ,
		_w9103_,
		_w9104_,
		_w20634_
	);
	LUT4 #(
		.INIT('h6e7f)
	) name18734 (
		_w9098_,
		_w9101_,
		_w20633_,
		_w20634_,
		_w20635_
	);
	LUT4 #(
		.INIT('h7fff)
	) name18735 (
		_w20626_,
		_w20629_,
		_w20632_,
		_w20635_,
		_w20636_
	);
	LUT3 #(
		.INIT('h80)
	) name18736 (
		\m0_data_i[27]_pad ,
		_w9103_,
		_w9104_,
		_w20637_
	);
	LUT3 #(
		.INIT('h2a)
	) name18737 (
		\m7_data_i[27]_pad ,
		_w9103_,
		_w9104_,
		_w20638_
	);
	LUT4 #(
		.INIT('h6e7f)
	) name18738 (
		_w9098_,
		_w9101_,
		_w20637_,
		_w20638_,
		_w20639_
	);
	LUT3 #(
		.INIT('h2a)
	) name18739 (
		\m3_data_i[27]_pad ,
		_w9103_,
		_w9104_,
		_w20640_
	);
	LUT3 #(
		.INIT('h80)
	) name18740 (
		\m2_data_i[27]_pad ,
		_w9103_,
		_w9104_,
		_w20641_
	);
	LUT3 #(
		.INIT('h57)
	) name18741 (
		_w9110_,
		_w20640_,
		_w20641_,
		_w20642_
	);
	LUT3 #(
		.INIT('h80)
	) name18742 (
		\m4_data_i[27]_pad ,
		_w9103_,
		_w9104_,
		_w20643_
	);
	LUT3 #(
		.INIT('h2a)
	) name18743 (
		\m1_data_i[27]_pad ,
		_w9103_,
		_w9104_,
		_w20644_
	);
	LUT4 #(
		.INIT('h57df)
	) name18744 (
		_w9098_,
		_w9101_,
		_w20643_,
		_w20644_,
		_w20645_
	);
	LUT3 #(
		.INIT('h80)
	) name18745 (
		\m6_data_i[27]_pad ,
		_w9103_,
		_w9104_,
		_w20646_
	);
	LUT3 #(
		.INIT('h2a)
	) name18746 (
		\m5_data_i[27]_pad ,
		_w9103_,
		_w9104_,
		_w20647_
	);
	LUT4 #(
		.INIT('hcdef)
	) name18747 (
		_w9098_,
		_w9101_,
		_w20646_,
		_w20647_,
		_w20648_
	);
	LUT4 #(
		.INIT('h7fff)
	) name18748 (
		_w20639_,
		_w20642_,
		_w20645_,
		_w20648_,
		_w20649_
	);
	LUT3 #(
		.INIT('h2a)
	) name18749 (
		\m1_data_i[28]_pad ,
		_w9103_,
		_w9104_,
		_w20650_
	);
	LUT3 #(
		.INIT('h80)
	) name18750 (
		\m2_data_i[28]_pad ,
		_w9103_,
		_w9104_,
		_w20651_
	);
	LUT4 #(
		.INIT('h3b7f)
	) name18751 (
		_w9098_,
		_w9101_,
		_w20650_,
		_w20651_,
		_w20652_
	);
	LUT3 #(
		.INIT('h80)
	) name18752 (
		\m0_data_i[28]_pad ,
		_w9103_,
		_w9104_,
		_w20653_
	);
	LUT3 #(
		.INIT('h2a)
	) name18753 (
		\m5_data_i[28]_pad ,
		_w9103_,
		_w9104_,
		_w20654_
	);
	LUT4 #(
		.INIT('h5d7f)
	) name18754 (
		_w9098_,
		_w9101_,
		_w20653_,
		_w20654_,
		_w20655_
	);
	LUT3 #(
		.INIT('h2a)
	) name18755 (
		\m7_data_i[28]_pad ,
		_w9103_,
		_w9104_,
		_w20656_
	);
	LUT3 #(
		.INIT('h80)
	) name18756 (
		\m6_data_i[28]_pad ,
		_w9103_,
		_w9104_,
		_w20657_
	);
	LUT3 #(
		.INIT('h57)
	) name18757 (
		_w9102_,
		_w20656_,
		_w20657_,
		_w20658_
	);
	LUT3 #(
		.INIT('h2a)
	) name18758 (
		\m3_data_i[28]_pad ,
		_w9103_,
		_w9104_,
		_w20659_
	);
	LUT3 #(
		.INIT('h80)
	) name18759 (
		\m4_data_i[28]_pad ,
		_w9103_,
		_w9104_,
		_w20660_
	);
	LUT4 #(
		.INIT('h9dbf)
	) name18760 (
		_w9098_,
		_w9101_,
		_w20659_,
		_w20660_,
		_w20661_
	);
	LUT4 #(
		.INIT('h7fff)
	) name18761 (
		_w20652_,
		_w20655_,
		_w20658_,
		_w20661_,
		_w20662_
	);
	LUT3 #(
		.INIT('h2a)
	) name18762 (
		\m1_data_i[29]_pad ,
		_w9103_,
		_w9104_,
		_w20663_
	);
	LUT3 #(
		.INIT('h80)
	) name18763 (
		\m2_data_i[29]_pad ,
		_w9103_,
		_w9104_,
		_w20664_
	);
	LUT4 #(
		.INIT('h3b7f)
	) name18764 (
		_w9098_,
		_w9101_,
		_w20663_,
		_w20664_,
		_w20665_
	);
	LUT3 #(
		.INIT('h80)
	) name18765 (
		\m0_data_i[29]_pad ,
		_w9103_,
		_w9104_,
		_w20666_
	);
	LUT3 #(
		.INIT('h80)
	) name18766 (
		\m4_data_i[29]_pad ,
		_w9103_,
		_w9104_,
		_w20667_
	);
	LUT4 #(
		.INIT('h5d7f)
	) name18767 (
		_w9098_,
		_w9101_,
		_w20666_,
		_w20667_,
		_w20668_
	);
	LUT3 #(
		.INIT('h2a)
	) name18768 (
		\m7_data_i[29]_pad ,
		_w9103_,
		_w9104_,
		_w20669_
	);
	LUT3 #(
		.INIT('h2a)
	) name18769 (
		\m3_data_i[29]_pad ,
		_w9103_,
		_w9104_,
		_w20670_
	);
	LUT4 #(
		.INIT('habef)
	) name18770 (
		_w9098_,
		_w9101_,
		_w20669_,
		_w20670_,
		_w20671_
	);
	LUT3 #(
		.INIT('h80)
	) name18771 (
		\m6_data_i[29]_pad ,
		_w9103_,
		_w9104_,
		_w20672_
	);
	LUT3 #(
		.INIT('h2a)
	) name18772 (
		\m5_data_i[29]_pad ,
		_w9103_,
		_w9104_,
		_w20673_
	);
	LUT4 #(
		.INIT('hcdef)
	) name18773 (
		_w9098_,
		_w9101_,
		_w20672_,
		_w20673_,
		_w20674_
	);
	LUT4 #(
		.INIT('h7fff)
	) name18774 (
		_w20665_,
		_w20668_,
		_w20671_,
		_w20674_,
		_w20675_
	);
	LUT3 #(
		.INIT('h80)
	) name18775 (
		\m6_data_i[2]_pad ,
		_w9103_,
		_w9104_,
		_w20676_
	);
	LUT3 #(
		.INIT('h2a)
	) name18776 (
		\m5_data_i[2]_pad ,
		_w9103_,
		_w9104_,
		_w20677_
	);
	LUT4 #(
		.INIT('hcdef)
	) name18777 (
		_w9098_,
		_w9101_,
		_w20676_,
		_w20677_,
		_w20678_
	);
	LUT3 #(
		.INIT('h2a)
	) name18778 (
		\m3_data_i[2]_pad ,
		_w9103_,
		_w9104_,
		_w20679_
	);
	LUT3 #(
		.INIT('h2a)
	) name18779 (
		\m7_data_i[2]_pad ,
		_w9103_,
		_w9104_,
		_w20680_
	);
	LUT4 #(
		.INIT('haebf)
	) name18780 (
		_w9098_,
		_w9101_,
		_w20679_,
		_w20680_,
		_w20681_
	);
	LUT3 #(
		.INIT('h80)
	) name18781 (
		\m4_data_i[2]_pad ,
		_w9103_,
		_w9104_,
		_w20682_
	);
	LUT3 #(
		.INIT('h80)
	) name18782 (
		\m0_data_i[2]_pad ,
		_w9103_,
		_w9104_,
		_w20683_
	);
	LUT4 #(
		.INIT('h57df)
	) name18783 (
		_w9098_,
		_w9101_,
		_w20682_,
		_w20683_,
		_w20684_
	);
	LUT3 #(
		.INIT('h2a)
	) name18784 (
		\m1_data_i[2]_pad ,
		_w9103_,
		_w9104_,
		_w20685_
	);
	LUT3 #(
		.INIT('h80)
	) name18785 (
		\m2_data_i[2]_pad ,
		_w9103_,
		_w9104_,
		_w20686_
	);
	LUT4 #(
		.INIT('h3b7f)
	) name18786 (
		_w9098_,
		_w9101_,
		_w20685_,
		_w20686_,
		_w20687_
	);
	LUT4 #(
		.INIT('h7fff)
	) name18787 (
		_w20678_,
		_w20681_,
		_w20684_,
		_w20687_,
		_w20688_
	);
	LUT3 #(
		.INIT('h2a)
	) name18788 (
		\m1_data_i[30]_pad ,
		_w9103_,
		_w9104_,
		_w20689_
	);
	LUT3 #(
		.INIT('h80)
	) name18789 (
		\m2_data_i[30]_pad ,
		_w9103_,
		_w9104_,
		_w20690_
	);
	LUT4 #(
		.INIT('h3b7f)
	) name18790 (
		_w9098_,
		_w9101_,
		_w20689_,
		_w20690_,
		_w20691_
	);
	LUT3 #(
		.INIT('h80)
	) name18791 (
		\m0_data_i[30]_pad ,
		_w9103_,
		_w9104_,
		_w20692_
	);
	LUT3 #(
		.INIT('h80)
	) name18792 (
		\m4_data_i[30]_pad ,
		_w9103_,
		_w9104_,
		_w20693_
	);
	LUT4 #(
		.INIT('h5d7f)
	) name18793 (
		_w9098_,
		_w9101_,
		_w20692_,
		_w20693_,
		_w20694_
	);
	LUT3 #(
		.INIT('h2a)
	) name18794 (
		\m7_data_i[30]_pad ,
		_w9103_,
		_w9104_,
		_w20695_
	);
	LUT3 #(
		.INIT('h2a)
	) name18795 (
		\m3_data_i[30]_pad ,
		_w9103_,
		_w9104_,
		_w20696_
	);
	LUT4 #(
		.INIT('habef)
	) name18796 (
		_w9098_,
		_w9101_,
		_w20695_,
		_w20696_,
		_w20697_
	);
	LUT3 #(
		.INIT('h80)
	) name18797 (
		\m6_data_i[30]_pad ,
		_w9103_,
		_w9104_,
		_w20698_
	);
	LUT3 #(
		.INIT('h2a)
	) name18798 (
		\m5_data_i[30]_pad ,
		_w9103_,
		_w9104_,
		_w20699_
	);
	LUT4 #(
		.INIT('hcdef)
	) name18799 (
		_w9098_,
		_w9101_,
		_w20698_,
		_w20699_,
		_w20700_
	);
	LUT4 #(
		.INIT('h7fff)
	) name18800 (
		_w20691_,
		_w20694_,
		_w20697_,
		_w20700_,
		_w20701_
	);
	LUT3 #(
		.INIT('h80)
	) name18801 (
		\m0_data_i[31]_pad ,
		_w9103_,
		_w9104_,
		_w20702_
	);
	LUT3 #(
		.INIT('h2a)
	) name18802 (
		\m7_data_i[31]_pad ,
		_w9103_,
		_w9104_,
		_w20703_
	);
	LUT4 #(
		.INIT('h6e7f)
	) name18803 (
		_w9098_,
		_w9101_,
		_w20702_,
		_w20703_,
		_w20704_
	);
	LUT3 #(
		.INIT('h2a)
	) name18804 (
		\m1_data_i[31]_pad ,
		_w9103_,
		_w9104_,
		_w20705_
	);
	LUT3 #(
		.INIT('h80)
	) name18805 (
		\m4_data_i[31]_pad ,
		_w9103_,
		_w9104_,
		_w20706_
	);
	LUT4 #(
		.INIT('h5d7f)
	) name18806 (
		_w9098_,
		_w9101_,
		_w20705_,
		_w20706_,
		_w20707_
	);
	LUT3 #(
		.INIT('h80)
	) name18807 (
		\m2_data_i[31]_pad ,
		_w9103_,
		_w9104_,
		_w20708_
	);
	LUT3 #(
		.INIT('h2a)
	) name18808 (
		\m3_data_i[31]_pad ,
		_w9103_,
		_w9104_,
		_w20709_
	);
	LUT3 #(
		.INIT('h57)
	) name18809 (
		_w9110_,
		_w20708_,
		_w20709_,
		_w20710_
	);
	LUT3 #(
		.INIT('h80)
	) name18810 (
		\m6_data_i[31]_pad ,
		_w9103_,
		_w9104_,
		_w20711_
	);
	LUT3 #(
		.INIT('h2a)
	) name18811 (
		\m5_data_i[31]_pad ,
		_w9103_,
		_w9104_,
		_w20712_
	);
	LUT4 #(
		.INIT('hcdef)
	) name18812 (
		_w9098_,
		_w9101_,
		_w20711_,
		_w20712_,
		_w20713_
	);
	LUT4 #(
		.INIT('h7fff)
	) name18813 (
		_w20704_,
		_w20707_,
		_w20710_,
		_w20713_,
		_w20714_
	);
	LUT3 #(
		.INIT('h2a)
	) name18814 (
		\m1_data_i[3]_pad ,
		_w9103_,
		_w9104_,
		_w20715_
	);
	LUT3 #(
		.INIT('h80)
	) name18815 (
		\m2_data_i[3]_pad ,
		_w9103_,
		_w9104_,
		_w20716_
	);
	LUT4 #(
		.INIT('h3b7f)
	) name18816 (
		_w9098_,
		_w9101_,
		_w20715_,
		_w20716_,
		_w20717_
	);
	LUT3 #(
		.INIT('h80)
	) name18817 (
		\m0_data_i[3]_pad ,
		_w9103_,
		_w9104_,
		_w20718_
	);
	LUT3 #(
		.INIT('h2a)
	) name18818 (
		\m5_data_i[3]_pad ,
		_w9103_,
		_w9104_,
		_w20719_
	);
	LUT4 #(
		.INIT('h5d7f)
	) name18819 (
		_w9098_,
		_w9101_,
		_w20718_,
		_w20719_,
		_w20720_
	);
	LUT3 #(
		.INIT('h2a)
	) name18820 (
		\m7_data_i[3]_pad ,
		_w9103_,
		_w9104_,
		_w20721_
	);
	LUT3 #(
		.INIT('h80)
	) name18821 (
		\m6_data_i[3]_pad ,
		_w9103_,
		_w9104_,
		_w20722_
	);
	LUT3 #(
		.INIT('h57)
	) name18822 (
		_w9102_,
		_w20721_,
		_w20722_,
		_w20723_
	);
	LUT3 #(
		.INIT('h2a)
	) name18823 (
		\m3_data_i[3]_pad ,
		_w9103_,
		_w9104_,
		_w20724_
	);
	LUT3 #(
		.INIT('h80)
	) name18824 (
		\m4_data_i[3]_pad ,
		_w9103_,
		_w9104_,
		_w20725_
	);
	LUT4 #(
		.INIT('h9dbf)
	) name18825 (
		_w9098_,
		_w9101_,
		_w20724_,
		_w20725_,
		_w20726_
	);
	LUT4 #(
		.INIT('h7fff)
	) name18826 (
		_w20717_,
		_w20720_,
		_w20723_,
		_w20726_,
		_w20727_
	);
	LUT3 #(
		.INIT('h2a)
	) name18827 (
		\m3_data_i[4]_pad ,
		_w9103_,
		_w9104_,
		_w20728_
	);
	LUT3 #(
		.INIT('h80)
	) name18828 (
		\m4_data_i[4]_pad ,
		_w9103_,
		_w9104_,
		_w20729_
	);
	LUT4 #(
		.INIT('h9dbf)
	) name18829 (
		_w9098_,
		_w9101_,
		_w20728_,
		_w20729_,
		_w20730_
	);
	LUT3 #(
		.INIT('h2a)
	) name18830 (
		\m1_data_i[4]_pad ,
		_w9103_,
		_w9104_,
		_w20731_
	);
	LUT3 #(
		.INIT('h2a)
	) name18831 (
		\m5_data_i[4]_pad ,
		_w9103_,
		_w9104_,
		_w20732_
	);
	LUT4 #(
		.INIT('h5d7f)
	) name18832 (
		_w9098_,
		_w9101_,
		_w20731_,
		_w20732_,
		_w20733_
	);
	LUT3 #(
		.INIT('h80)
	) name18833 (
		\m2_data_i[4]_pad ,
		_w9103_,
		_w9104_,
		_w20734_
	);
	LUT3 #(
		.INIT('h80)
	) name18834 (
		\m6_data_i[4]_pad ,
		_w9103_,
		_w9104_,
		_w20735_
	);
	LUT4 #(
		.INIT('haebf)
	) name18835 (
		_w9098_,
		_w9101_,
		_w20734_,
		_w20735_,
		_w20736_
	);
	LUT3 #(
		.INIT('h80)
	) name18836 (
		\m0_data_i[4]_pad ,
		_w9103_,
		_w9104_,
		_w20737_
	);
	LUT3 #(
		.INIT('h2a)
	) name18837 (
		\m7_data_i[4]_pad ,
		_w9103_,
		_w9104_,
		_w20738_
	);
	LUT4 #(
		.INIT('h6e7f)
	) name18838 (
		_w9098_,
		_w9101_,
		_w20737_,
		_w20738_,
		_w20739_
	);
	LUT4 #(
		.INIT('h7fff)
	) name18839 (
		_w20730_,
		_w20733_,
		_w20736_,
		_w20739_,
		_w20740_
	);
	LUT3 #(
		.INIT('h80)
	) name18840 (
		\m6_data_i[5]_pad ,
		_w9103_,
		_w9104_,
		_w20741_
	);
	LUT3 #(
		.INIT('h2a)
	) name18841 (
		\m5_data_i[5]_pad ,
		_w9103_,
		_w9104_,
		_w20742_
	);
	LUT4 #(
		.INIT('hcdef)
	) name18842 (
		_w9098_,
		_w9101_,
		_w20741_,
		_w20742_,
		_w20743_
	);
	LUT3 #(
		.INIT('h80)
	) name18843 (
		\m0_data_i[5]_pad ,
		_w9103_,
		_w9104_,
		_w20744_
	);
	LUT3 #(
		.INIT('h80)
	) name18844 (
		\m4_data_i[5]_pad ,
		_w9103_,
		_w9104_,
		_w20745_
	);
	LUT4 #(
		.INIT('h5d7f)
	) name18845 (
		_w9098_,
		_w9101_,
		_w20744_,
		_w20745_,
		_w20746_
	);
	LUT3 #(
		.INIT('h2a)
	) name18846 (
		\m7_data_i[5]_pad ,
		_w9103_,
		_w9104_,
		_w20747_
	);
	LUT3 #(
		.INIT('h2a)
	) name18847 (
		\m3_data_i[5]_pad ,
		_w9103_,
		_w9104_,
		_w20748_
	);
	LUT4 #(
		.INIT('habef)
	) name18848 (
		_w9098_,
		_w9101_,
		_w20747_,
		_w20748_,
		_w20749_
	);
	LUT3 #(
		.INIT('h2a)
	) name18849 (
		\m1_data_i[5]_pad ,
		_w9103_,
		_w9104_,
		_w20750_
	);
	LUT3 #(
		.INIT('h80)
	) name18850 (
		\m2_data_i[5]_pad ,
		_w9103_,
		_w9104_,
		_w20751_
	);
	LUT4 #(
		.INIT('h3b7f)
	) name18851 (
		_w9098_,
		_w9101_,
		_w20750_,
		_w20751_,
		_w20752_
	);
	LUT4 #(
		.INIT('h7fff)
	) name18852 (
		_w20743_,
		_w20746_,
		_w20749_,
		_w20752_,
		_w20753_
	);
	LUT3 #(
		.INIT('h2a)
	) name18853 (
		\m1_data_i[6]_pad ,
		_w9103_,
		_w9104_,
		_w20754_
	);
	LUT3 #(
		.INIT('h80)
	) name18854 (
		\m2_data_i[6]_pad ,
		_w9103_,
		_w9104_,
		_w20755_
	);
	LUT4 #(
		.INIT('h3b7f)
	) name18855 (
		_w9098_,
		_w9101_,
		_w20754_,
		_w20755_,
		_w20756_
	);
	LUT3 #(
		.INIT('h2a)
	) name18856 (
		\m3_data_i[6]_pad ,
		_w9103_,
		_w9104_,
		_w20757_
	);
	LUT3 #(
		.INIT('h2a)
	) name18857 (
		\m5_data_i[6]_pad ,
		_w9103_,
		_w9104_,
		_w20758_
	);
	LUT4 #(
		.INIT('h9dbf)
	) name18858 (
		_w9098_,
		_w9101_,
		_w20757_,
		_w20758_,
		_w20759_
	);
	LUT3 #(
		.INIT('h80)
	) name18859 (
		\m4_data_i[6]_pad ,
		_w9103_,
		_w9104_,
		_w20760_
	);
	LUT3 #(
		.INIT('h80)
	) name18860 (
		\m6_data_i[6]_pad ,
		_w9103_,
		_w9104_,
		_w20761_
	);
	LUT4 #(
		.INIT('hcedf)
	) name18861 (
		_w9098_,
		_w9101_,
		_w20760_,
		_w20761_,
		_w20762_
	);
	LUT3 #(
		.INIT('h80)
	) name18862 (
		\m0_data_i[6]_pad ,
		_w9103_,
		_w9104_,
		_w20763_
	);
	LUT3 #(
		.INIT('h2a)
	) name18863 (
		\m7_data_i[6]_pad ,
		_w9103_,
		_w9104_,
		_w20764_
	);
	LUT4 #(
		.INIT('h6e7f)
	) name18864 (
		_w9098_,
		_w9101_,
		_w20763_,
		_w20764_,
		_w20765_
	);
	LUT4 #(
		.INIT('h7fff)
	) name18865 (
		_w20756_,
		_w20759_,
		_w20762_,
		_w20765_,
		_w20766_
	);
	LUT3 #(
		.INIT('h80)
	) name18866 (
		\m6_data_i[7]_pad ,
		_w9103_,
		_w9104_,
		_w20767_
	);
	LUT3 #(
		.INIT('h2a)
	) name18867 (
		\m5_data_i[7]_pad ,
		_w9103_,
		_w9104_,
		_w20768_
	);
	LUT4 #(
		.INIT('hcdef)
	) name18868 (
		_w9098_,
		_w9101_,
		_w20767_,
		_w20768_,
		_w20769_
	);
	LUT3 #(
		.INIT('h2a)
	) name18869 (
		\m3_data_i[7]_pad ,
		_w9103_,
		_w9104_,
		_w20770_
	);
	LUT3 #(
		.INIT('h80)
	) name18870 (
		\m2_data_i[7]_pad ,
		_w9103_,
		_w9104_,
		_w20771_
	);
	LUT3 #(
		.INIT('h57)
	) name18871 (
		_w9110_,
		_w20770_,
		_w20771_,
		_w20772_
	);
	LUT3 #(
		.INIT('h80)
	) name18872 (
		\m4_data_i[7]_pad ,
		_w9103_,
		_w9104_,
		_w20773_
	);
	LUT3 #(
		.INIT('h2a)
	) name18873 (
		\m1_data_i[7]_pad ,
		_w9103_,
		_w9104_,
		_w20774_
	);
	LUT4 #(
		.INIT('h57df)
	) name18874 (
		_w9098_,
		_w9101_,
		_w20773_,
		_w20774_,
		_w20775_
	);
	LUT3 #(
		.INIT('h80)
	) name18875 (
		\m0_data_i[7]_pad ,
		_w9103_,
		_w9104_,
		_w20776_
	);
	LUT3 #(
		.INIT('h2a)
	) name18876 (
		\m7_data_i[7]_pad ,
		_w9103_,
		_w9104_,
		_w20777_
	);
	LUT4 #(
		.INIT('h6e7f)
	) name18877 (
		_w9098_,
		_w9101_,
		_w20776_,
		_w20777_,
		_w20778_
	);
	LUT4 #(
		.INIT('h7fff)
	) name18878 (
		_w20769_,
		_w20772_,
		_w20775_,
		_w20778_,
		_w20779_
	);
	LUT3 #(
		.INIT('h80)
	) name18879 (
		\m6_data_i[8]_pad ,
		_w9103_,
		_w9104_,
		_w20780_
	);
	LUT3 #(
		.INIT('h2a)
	) name18880 (
		\m5_data_i[8]_pad ,
		_w9103_,
		_w9104_,
		_w20781_
	);
	LUT4 #(
		.INIT('hcdef)
	) name18881 (
		_w9098_,
		_w9101_,
		_w20780_,
		_w20781_,
		_w20782_
	);
	LUT3 #(
		.INIT('h2a)
	) name18882 (
		\m3_data_i[8]_pad ,
		_w9103_,
		_w9104_,
		_w20783_
	);
	LUT3 #(
		.INIT('h2a)
	) name18883 (
		\m7_data_i[8]_pad ,
		_w9103_,
		_w9104_,
		_w20784_
	);
	LUT4 #(
		.INIT('haebf)
	) name18884 (
		_w9098_,
		_w9101_,
		_w20783_,
		_w20784_,
		_w20785_
	);
	LUT3 #(
		.INIT('h80)
	) name18885 (
		\m4_data_i[8]_pad ,
		_w9103_,
		_w9104_,
		_w20786_
	);
	LUT3 #(
		.INIT('h80)
	) name18886 (
		\m0_data_i[8]_pad ,
		_w9103_,
		_w9104_,
		_w20787_
	);
	LUT4 #(
		.INIT('h57df)
	) name18887 (
		_w9098_,
		_w9101_,
		_w20786_,
		_w20787_,
		_w20788_
	);
	LUT3 #(
		.INIT('h2a)
	) name18888 (
		\m1_data_i[8]_pad ,
		_w9103_,
		_w9104_,
		_w20789_
	);
	LUT3 #(
		.INIT('h80)
	) name18889 (
		\m2_data_i[8]_pad ,
		_w9103_,
		_w9104_,
		_w20790_
	);
	LUT4 #(
		.INIT('h3b7f)
	) name18890 (
		_w9098_,
		_w9101_,
		_w20789_,
		_w20790_,
		_w20791_
	);
	LUT4 #(
		.INIT('h7fff)
	) name18891 (
		_w20782_,
		_w20785_,
		_w20788_,
		_w20791_,
		_w20792_
	);
	LUT3 #(
		.INIT('h80)
	) name18892 (
		\m6_data_i[9]_pad ,
		_w9103_,
		_w9104_,
		_w20793_
	);
	LUT3 #(
		.INIT('h2a)
	) name18893 (
		\m5_data_i[9]_pad ,
		_w9103_,
		_w9104_,
		_w20794_
	);
	LUT4 #(
		.INIT('hcdef)
	) name18894 (
		_w9098_,
		_w9101_,
		_w20793_,
		_w20794_,
		_w20795_
	);
	LUT3 #(
		.INIT('h2a)
	) name18895 (
		\m1_data_i[9]_pad ,
		_w9103_,
		_w9104_,
		_w20796_
	);
	LUT3 #(
		.INIT('h2a)
	) name18896 (
		\m7_data_i[9]_pad ,
		_w9103_,
		_w9104_,
		_w20797_
	);
	LUT4 #(
		.INIT('h6e7f)
	) name18897 (
		_w9098_,
		_w9101_,
		_w20796_,
		_w20797_,
		_w20798_
	);
	LUT3 #(
		.INIT('h80)
	) name18898 (
		\m2_data_i[9]_pad ,
		_w9103_,
		_w9104_,
		_w20799_
	);
	LUT3 #(
		.INIT('h80)
	) name18899 (
		\m0_data_i[9]_pad ,
		_w9103_,
		_w9104_,
		_w20800_
	);
	LUT4 #(
		.INIT('h37bf)
	) name18900 (
		_w9098_,
		_w9101_,
		_w20799_,
		_w20800_,
		_w20801_
	);
	LUT3 #(
		.INIT('h2a)
	) name18901 (
		\m3_data_i[9]_pad ,
		_w9103_,
		_w9104_,
		_w20802_
	);
	LUT3 #(
		.INIT('h80)
	) name18902 (
		\m4_data_i[9]_pad ,
		_w9103_,
		_w9104_,
		_w20803_
	);
	LUT4 #(
		.INIT('h9dbf)
	) name18903 (
		_w9098_,
		_w9101_,
		_w20802_,
		_w20803_,
		_w20804_
	);
	LUT4 #(
		.INIT('h7fff)
	) name18904 (
		_w20795_,
		_w20798_,
		_w20801_,
		_w20804_,
		_w20805_
	);
	LUT3 #(
		.INIT('h2a)
	) name18905 (
		\m3_sel_i[0]_pad ,
		_w9103_,
		_w9104_,
		_w20806_
	);
	LUT3 #(
		.INIT('h80)
	) name18906 (
		\m4_sel_i[0]_pad ,
		_w9103_,
		_w9104_,
		_w20807_
	);
	LUT4 #(
		.INIT('h9dbf)
	) name18907 (
		_w9098_,
		_w9101_,
		_w20806_,
		_w20807_,
		_w20808_
	);
	LUT3 #(
		.INIT('h80)
	) name18908 (
		\m6_sel_i[0]_pad ,
		_w9103_,
		_w9104_,
		_w20809_
	);
	LUT3 #(
		.INIT('h80)
	) name18909 (
		\m2_sel_i[0]_pad ,
		_w9103_,
		_w9104_,
		_w20810_
	);
	LUT4 #(
		.INIT('habef)
	) name18910 (
		_w9098_,
		_w9101_,
		_w20809_,
		_w20810_,
		_w20811_
	);
	LUT3 #(
		.INIT('h2a)
	) name18911 (
		\m5_sel_i[0]_pad ,
		_w9103_,
		_w9104_,
		_w20812_
	);
	LUT3 #(
		.INIT('h2a)
	) name18912 (
		\m1_sel_i[0]_pad ,
		_w9103_,
		_w9104_,
		_w20813_
	);
	LUT4 #(
		.INIT('h57df)
	) name18913 (
		_w9098_,
		_w9101_,
		_w20812_,
		_w20813_,
		_w20814_
	);
	LUT3 #(
		.INIT('h80)
	) name18914 (
		\m0_sel_i[0]_pad ,
		_w9103_,
		_w9104_,
		_w20815_
	);
	LUT3 #(
		.INIT('h2a)
	) name18915 (
		\m7_sel_i[0]_pad ,
		_w9103_,
		_w9104_,
		_w20816_
	);
	LUT4 #(
		.INIT('h6e7f)
	) name18916 (
		_w9098_,
		_w9101_,
		_w20815_,
		_w20816_,
		_w20817_
	);
	LUT4 #(
		.INIT('h7fff)
	) name18917 (
		_w20808_,
		_w20811_,
		_w20814_,
		_w20817_,
		_w20818_
	);
	LUT3 #(
		.INIT('h80)
	) name18918 (
		\m0_sel_i[1]_pad ,
		_w9103_,
		_w9104_,
		_w20819_
	);
	LUT3 #(
		.INIT('h2a)
	) name18919 (
		\m7_sel_i[1]_pad ,
		_w9103_,
		_w9104_,
		_w20820_
	);
	LUT4 #(
		.INIT('h6e7f)
	) name18920 (
		_w9098_,
		_w9101_,
		_w20819_,
		_w20820_,
		_w20821_
	);
	LUT3 #(
		.INIT('h80)
	) name18921 (
		\m6_sel_i[1]_pad ,
		_w9103_,
		_w9104_,
		_w20822_
	);
	LUT3 #(
		.INIT('h80)
	) name18922 (
		\m2_sel_i[1]_pad ,
		_w9103_,
		_w9104_,
		_w20823_
	);
	LUT4 #(
		.INIT('habef)
	) name18923 (
		_w9098_,
		_w9101_,
		_w20822_,
		_w20823_,
		_w20824_
	);
	LUT3 #(
		.INIT('h2a)
	) name18924 (
		\m5_sel_i[1]_pad ,
		_w9103_,
		_w9104_,
		_w20825_
	);
	LUT3 #(
		.INIT('h2a)
	) name18925 (
		\m1_sel_i[1]_pad ,
		_w9103_,
		_w9104_,
		_w20826_
	);
	LUT4 #(
		.INIT('h57df)
	) name18926 (
		_w9098_,
		_w9101_,
		_w20825_,
		_w20826_,
		_w20827_
	);
	LUT3 #(
		.INIT('h2a)
	) name18927 (
		\m3_sel_i[1]_pad ,
		_w9103_,
		_w9104_,
		_w20828_
	);
	LUT3 #(
		.INIT('h80)
	) name18928 (
		\m4_sel_i[1]_pad ,
		_w9103_,
		_w9104_,
		_w20829_
	);
	LUT4 #(
		.INIT('h9dbf)
	) name18929 (
		_w9098_,
		_w9101_,
		_w20828_,
		_w20829_,
		_w20830_
	);
	LUT4 #(
		.INIT('h7fff)
	) name18930 (
		_w20821_,
		_w20824_,
		_w20827_,
		_w20830_,
		_w20831_
	);
	LUT3 #(
		.INIT('h2a)
	) name18931 (
		\m1_sel_i[2]_pad ,
		_w9103_,
		_w9104_,
		_w20832_
	);
	LUT3 #(
		.INIT('h80)
	) name18932 (
		\m2_sel_i[2]_pad ,
		_w9103_,
		_w9104_,
		_w20833_
	);
	LUT4 #(
		.INIT('h3b7f)
	) name18933 (
		_w9098_,
		_w9101_,
		_w20832_,
		_w20833_,
		_w20834_
	);
	LUT3 #(
		.INIT('h2a)
	) name18934 (
		\m3_sel_i[2]_pad ,
		_w9103_,
		_w9104_,
		_w20835_
	);
	LUT3 #(
		.INIT('h2a)
	) name18935 (
		\m7_sel_i[2]_pad ,
		_w9103_,
		_w9104_,
		_w20836_
	);
	LUT4 #(
		.INIT('haebf)
	) name18936 (
		_w9098_,
		_w9101_,
		_w20835_,
		_w20836_,
		_w20837_
	);
	LUT3 #(
		.INIT('h80)
	) name18937 (
		\m4_sel_i[2]_pad ,
		_w9103_,
		_w9104_,
		_w20838_
	);
	LUT3 #(
		.INIT('h80)
	) name18938 (
		\m0_sel_i[2]_pad ,
		_w9103_,
		_w9104_,
		_w20839_
	);
	LUT4 #(
		.INIT('h57df)
	) name18939 (
		_w9098_,
		_w9101_,
		_w20838_,
		_w20839_,
		_w20840_
	);
	LUT3 #(
		.INIT('h80)
	) name18940 (
		\m6_sel_i[2]_pad ,
		_w9103_,
		_w9104_,
		_w20841_
	);
	LUT3 #(
		.INIT('h2a)
	) name18941 (
		\m5_sel_i[2]_pad ,
		_w9103_,
		_w9104_,
		_w20842_
	);
	LUT4 #(
		.INIT('hcdef)
	) name18942 (
		_w9098_,
		_w9101_,
		_w20841_,
		_w20842_,
		_w20843_
	);
	LUT4 #(
		.INIT('h7fff)
	) name18943 (
		_w20834_,
		_w20837_,
		_w20840_,
		_w20843_,
		_w20844_
	);
	LUT3 #(
		.INIT('h2a)
	) name18944 (
		\m3_sel_i[3]_pad ,
		_w9103_,
		_w9104_,
		_w20845_
	);
	LUT3 #(
		.INIT('h80)
	) name18945 (
		\m4_sel_i[3]_pad ,
		_w9103_,
		_w9104_,
		_w20846_
	);
	LUT4 #(
		.INIT('h9dbf)
	) name18946 (
		_w9098_,
		_w9101_,
		_w20845_,
		_w20846_,
		_w20847_
	);
	LUT3 #(
		.INIT('h80)
	) name18947 (
		\m6_sel_i[3]_pad ,
		_w9103_,
		_w9104_,
		_w20848_
	);
	LUT3 #(
		.INIT('h80)
	) name18948 (
		\m2_sel_i[3]_pad ,
		_w9103_,
		_w9104_,
		_w20849_
	);
	LUT4 #(
		.INIT('habef)
	) name18949 (
		_w9098_,
		_w9101_,
		_w20848_,
		_w20849_,
		_w20850_
	);
	LUT3 #(
		.INIT('h2a)
	) name18950 (
		\m5_sel_i[3]_pad ,
		_w9103_,
		_w9104_,
		_w20851_
	);
	LUT3 #(
		.INIT('h2a)
	) name18951 (
		\m1_sel_i[3]_pad ,
		_w9103_,
		_w9104_,
		_w20852_
	);
	LUT4 #(
		.INIT('h57df)
	) name18952 (
		_w9098_,
		_w9101_,
		_w20851_,
		_w20852_,
		_w20853_
	);
	LUT3 #(
		.INIT('h80)
	) name18953 (
		\m0_sel_i[3]_pad ,
		_w9103_,
		_w9104_,
		_w20854_
	);
	LUT3 #(
		.INIT('h2a)
	) name18954 (
		\m7_sel_i[3]_pad ,
		_w9103_,
		_w9104_,
		_w20855_
	);
	LUT4 #(
		.INIT('h6e7f)
	) name18955 (
		_w9098_,
		_w9101_,
		_w20854_,
		_w20855_,
		_w20856_
	);
	LUT4 #(
		.INIT('h7fff)
	) name18956 (
		_w20847_,
		_w20850_,
		_w20853_,
		_w20856_,
		_w20857_
	);
	LUT4 #(
		.INIT('h2a00)
	) name18957 (
		\m1_stb_i_pad ,
		_w9103_,
		_w9104_,
		_w9322_,
		_w20858_
	);
	LUT4 #(
		.INIT('h8000)
	) name18958 (
		\m6_stb_i_pad ,
		_w9103_,
		_w9104_,
		_w9312_,
		_w20859_
	);
	LUT4 #(
		.INIT('h6e7f)
	) name18959 (
		_w9098_,
		_w9101_,
		_w20858_,
		_w20859_,
		_w20860_
	);
	LUT4 #(
		.INIT('h8000)
	) name18960 (
		\m2_stb_i_pad ,
		_w9103_,
		_w9104_,
		_w9288_,
		_w20861_
	);
	LUT4 #(
		.INIT('h2a00)
	) name18961 (
		\m3_stb_i_pad ,
		_w9103_,
		_w9104_,
		_w9295_,
		_w20862_
	);
	LUT3 #(
		.INIT('h57)
	) name18962 (
		_w9110_,
		_w20861_,
		_w20862_,
		_w20863_
	);
	LUT4 #(
		.INIT('h8000)
	) name18963 (
		\m0_stb_i_pad ,
		_w9103_,
		_w9104_,
		_w9277_,
		_w20864_
	);
	LUT4 #(
		.INIT('h2a00)
	) name18964 (
		\m5_stb_i_pad ,
		_w9103_,
		_w9104_,
		_w9269_,
		_w20865_
	);
	LUT4 #(
		.INIT('h5d7f)
	) name18965 (
		_w9098_,
		_w9101_,
		_w20864_,
		_w20865_,
		_w20866_
	);
	LUT4 #(
		.INIT('h8000)
	) name18966 (
		\m4_stb_i_pad ,
		_w9103_,
		_w9104_,
		_w9302_,
		_w20867_
	);
	LUT4 #(
		.INIT('h2a00)
	) name18967 (
		\m7_stb_i_pad ,
		_w9103_,
		_w9104_,
		_w9319_,
		_w20868_
	);
	LUT4 #(
		.INIT('hcedf)
	) name18968 (
		_w9098_,
		_w9101_,
		_w20867_,
		_w20868_,
		_w20869_
	);
	LUT4 #(
		.INIT('h7fff)
	) name18969 (
		_w20860_,
		_w20863_,
		_w20866_,
		_w20869_,
		_w20870_
	);
	LUT3 #(
		.INIT('h2a)
	) name18970 (
		\m3_we_i_pad ,
		_w9103_,
		_w9104_,
		_w20871_
	);
	LUT3 #(
		.INIT('h80)
	) name18971 (
		\m4_we_i_pad ,
		_w9103_,
		_w9104_,
		_w20872_
	);
	LUT4 #(
		.INIT('h9dbf)
	) name18972 (
		_w9098_,
		_w9101_,
		_w20871_,
		_w20872_,
		_w20873_
	);
	LUT3 #(
		.INIT('h80)
	) name18973 (
		\m6_we_i_pad ,
		_w9103_,
		_w9104_,
		_w20874_
	);
	LUT3 #(
		.INIT('h80)
	) name18974 (
		\m2_we_i_pad ,
		_w9103_,
		_w9104_,
		_w20875_
	);
	LUT4 #(
		.INIT('habef)
	) name18975 (
		_w9098_,
		_w9101_,
		_w20874_,
		_w20875_,
		_w20876_
	);
	LUT3 #(
		.INIT('h2a)
	) name18976 (
		\m5_we_i_pad ,
		_w9103_,
		_w9104_,
		_w20877_
	);
	LUT3 #(
		.INIT('h2a)
	) name18977 (
		\m1_we_i_pad ,
		_w9103_,
		_w9104_,
		_w20878_
	);
	LUT4 #(
		.INIT('h57df)
	) name18978 (
		_w9098_,
		_w9101_,
		_w20877_,
		_w20878_,
		_w20879_
	);
	LUT3 #(
		.INIT('h80)
	) name18979 (
		\m0_we_i_pad ,
		_w9103_,
		_w9104_,
		_w20880_
	);
	LUT3 #(
		.INIT('h2a)
	) name18980 (
		\m7_we_i_pad ,
		_w9103_,
		_w9104_,
		_w20881_
	);
	LUT4 #(
		.INIT('h6e7f)
	) name18981 (
		_w9098_,
		_w9101_,
		_w20880_,
		_w20881_,
		_w20882_
	);
	LUT4 #(
		.INIT('h7fff)
	) name18982 (
		_w20873_,
		_w20876_,
		_w20879_,
		_w20882_,
		_w20883_
	);
	LUT3 #(
		.INIT('h2a)
	) name18983 (
		\m3_addr_i[0]_pad ,
		_w9171_,
		_w9172_,
		_w20884_
	);
	LUT3 #(
		.INIT('h80)
	) name18984 (
		\m4_addr_i[0]_pad ,
		_w9171_,
		_w9172_,
		_w20885_
	);
	LUT4 #(
		.INIT('h9dbf)
	) name18985 (
		_w9166_,
		_w9169_,
		_w20884_,
		_w20885_,
		_w20886_
	);
	LUT3 #(
		.INIT('h80)
	) name18986 (
		\m6_addr_i[0]_pad ,
		_w9171_,
		_w9172_,
		_w20887_
	);
	LUT3 #(
		.INIT('h80)
	) name18987 (
		\m2_addr_i[0]_pad ,
		_w9171_,
		_w9172_,
		_w20888_
	);
	LUT4 #(
		.INIT('habef)
	) name18988 (
		_w9166_,
		_w9169_,
		_w20887_,
		_w20888_,
		_w20889_
	);
	LUT3 #(
		.INIT('h2a)
	) name18989 (
		\m5_addr_i[0]_pad ,
		_w9171_,
		_w9172_,
		_w20890_
	);
	LUT3 #(
		.INIT('h2a)
	) name18990 (
		\m1_addr_i[0]_pad ,
		_w9171_,
		_w9172_,
		_w20891_
	);
	LUT4 #(
		.INIT('h57df)
	) name18991 (
		_w9166_,
		_w9169_,
		_w20890_,
		_w20891_,
		_w20892_
	);
	LUT3 #(
		.INIT('h80)
	) name18992 (
		\m0_addr_i[0]_pad ,
		_w9171_,
		_w9172_,
		_w20893_
	);
	LUT3 #(
		.INIT('h2a)
	) name18993 (
		\m7_addr_i[0]_pad ,
		_w9171_,
		_w9172_,
		_w20894_
	);
	LUT4 #(
		.INIT('h6e7f)
	) name18994 (
		_w9166_,
		_w9169_,
		_w20893_,
		_w20894_,
		_w20895_
	);
	LUT4 #(
		.INIT('h7fff)
	) name18995 (
		_w20886_,
		_w20889_,
		_w20892_,
		_w20895_,
		_w20896_
	);
	LUT3 #(
		.INIT('h2a)
	) name18996 (
		\m3_addr_i[10]_pad ,
		_w9171_,
		_w9172_,
		_w20897_
	);
	LUT3 #(
		.INIT('h80)
	) name18997 (
		\m4_addr_i[10]_pad ,
		_w9171_,
		_w9172_,
		_w20898_
	);
	LUT4 #(
		.INIT('h9dbf)
	) name18998 (
		_w9166_,
		_w9169_,
		_w20897_,
		_w20898_,
		_w20899_
	);
	LUT3 #(
		.INIT('h80)
	) name18999 (
		\m6_addr_i[10]_pad ,
		_w9171_,
		_w9172_,
		_w20900_
	);
	LUT3 #(
		.INIT('h80)
	) name19000 (
		\m2_addr_i[10]_pad ,
		_w9171_,
		_w9172_,
		_w20901_
	);
	LUT4 #(
		.INIT('habef)
	) name19001 (
		_w9166_,
		_w9169_,
		_w20900_,
		_w20901_,
		_w20902_
	);
	LUT3 #(
		.INIT('h2a)
	) name19002 (
		\m5_addr_i[10]_pad ,
		_w9171_,
		_w9172_,
		_w20903_
	);
	LUT3 #(
		.INIT('h2a)
	) name19003 (
		\m1_addr_i[10]_pad ,
		_w9171_,
		_w9172_,
		_w20904_
	);
	LUT4 #(
		.INIT('h57df)
	) name19004 (
		_w9166_,
		_w9169_,
		_w20903_,
		_w20904_,
		_w20905_
	);
	LUT3 #(
		.INIT('h80)
	) name19005 (
		\m0_addr_i[10]_pad ,
		_w9171_,
		_w9172_,
		_w20906_
	);
	LUT3 #(
		.INIT('h2a)
	) name19006 (
		\m7_addr_i[10]_pad ,
		_w9171_,
		_w9172_,
		_w20907_
	);
	LUT4 #(
		.INIT('h6e7f)
	) name19007 (
		_w9166_,
		_w9169_,
		_w20906_,
		_w20907_,
		_w20908_
	);
	LUT4 #(
		.INIT('h7fff)
	) name19008 (
		_w20899_,
		_w20902_,
		_w20905_,
		_w20908_,
		_w20909_
	);
	LUT3 #(
		.INIT('h2a)
	) name19009 (
		\m3_addr_i[11]_pad ,
		_w9171_,
		_w9172_,
		_w20910_
	);
	LUT3 #(
		.INIT('h80)
	) name19010 (
		\m4_addr_i[11]_pad ,
		_w9171_,
		_w9172_,
		_w20911_
	);
	LUT4 #(
		.INIT('h9dbf)
	) name19011 (
		_w9166_,
		_w9169_,
		_w20910_,
		_w20911_,
		_w20912_
	);
	LUT3 #(
		.INIT('h80)
	) name19012 (
		\m6_addr_i[11]_pad ,
		_w9171_,
		_w9172_,
		_w20913_
	);
	LUT3 #(
		.INIT('h80)
	) name19013 (
		\m2_addr_i[11]_pad ,
		_w9171_,
		_w9172_,
		_w20914_
	);
	LUT4 #(
		.INIT('habef)
	) name19014 (
		_w9166_,
		_w9169_,
		_w20913_,
		_w20914_,
		_w20915_
	);
	LUT3 #(
		.INIT('h2a)
	) name19015 (
		\m5_addr_i[11]_pad ,
		_w9171_,
		_w9172_,
		_w20916_
	);
	LUT3 #(
		.INIT('h2a)
	) name19016 (
		\m1_addr_i[11]_pad ,
		_w9171_,
		_w9172_,
		_w20917_
	);
	LUT4 #(
		.INIT('h57df)
	) name19017 (
		_w9166_,
		_w9169_,
		_w20916_,
		_w20917_,
		_w20918_
	);
	LUT3 #(
		.INIT('h80)
	) name19018 (
		\m0_addr_i[11]_pad ,
		_w9171_,
		_w9172_,
		_w20919_
	);
	LUT3 #(
		.INIT('h2a)
	) name19019 (
		\m7_addr_i[11]_pad ,
		_w9171_,
		_w9172_,
		_w20920_
	);
	LUT4 #(
		.INIT('h6e7f)
	) name19020 (
		_w9166_,
		_w9169_,
		_w20919_,
		_w20920_,
		_w20921_
	);
	LUT4 #(
		.INIT('h7fff)
	) name19021 (
		_w20912_,
		_w20915_,
		_w20918_,
		_w20921_,
		_w20922_
	);
	LUT3 #(
		.INIT('h2a)
	) name19022 (
		\m3_addr_i[12]_pad ,
		_w9171_,
		_w9172_,
		_w20923_
	);
	LUT3 #(
		.INIT('h80)
	) name19023 (
		\m4_addr_i[12]_pad ,
		_w9171_,
		_w9172_,
		_w20924_
	);
	LUT4 #(
		.INIT('h9dbf)
	) name19024 (
		_w9166_,
		_w9169_,
		_w20923_,
		_w20924_,
		_w20925_
	);
	LUT3 #(
		.INIT('h80)
	) name19025 (
		\m6_addr_i[12]_pad ,
		_w9171_,
		_w9172_,
		_w20926_
	);
	LUT3 #(
		.INIT('h80)
	) name19026 (
		\m2_addr_i[12]_pad ,
		_w9171_,
		_w9172_,
		_w20927_
	);
	LUT4 #(
		.INIT('habef)
	) name19027 (
		_w9166_,
		_w9169_,
		_w20926_,
		_w20927_,
		_w20928_
	);
	LUT3 #(
		.INIT('h2a)
	) name19028 (
		\m5_addr_i[12]_pad ,
		_w9171_,
		_w9172_,
		_w20929_
	);
	LUT3 #(
		.INIT('h2a)
	) name19029 (
		\m1_addr_i[12]_pad ,
		_w9171_,
		_w9172_,
		_w20930_
	);
	LUT4 #(
		.INIT('h57df)
	) name19030 (
		_w9166_,
		_w9169_,
		_w20929_,
		_w20930_,
		_w20931_
	);
	LUT3 #(
		.INIT('h80)
	) name19031 (
		\m0_addr_i[12]_pad ,
		_w9171_,
		_w9172_,
		_w20932_
	);
	LUT3 #(
		.INIT('h2a)
	) name19032 (
		\m7_addr_i[12]_pad ,
		_w9171_,
		_w9172_,
		_w20933_
	);
	LUT4 #(
		.INIT('h6e7f)
	) name19033 (
		_w9166_,
		_w9169_,
		_w20932_,
		_w20933_,
		_w20934_
	);
	LUT4 #(
		.INIT('h7fff)
	) name19034 (
		_w20925_,
		_w20928_,
		_w20931_,
		_w20934_,
		_w20935_
	);
	LUT3 #(
		.INIT('h2a)
	) name19035 (
		\m3_addr_i[13]_pad ,
		_w9171_,
		_w9172_,
		_w20936_
	);
	LUT3 #(
		.INIT('h80)
	) name19036 (
		\m4_addr_i[13]_pad ,
		_w9171_,
		_w9172_,
		_w20937_
	);
	LUT4 #(
		.INIT('h9dbf)
	) name19037 (
		_w9166_,
		_w9169_,
		_w20936_,
		_w20937_,
		_w20938_
	);
	LUT3 #(
		.INIT('h80)
	) name19038 (
		\m6_addr_i[13]_pad ,
		_w9171_,
		_w9172_,
		_w20939_
	);
	LUT3 #(
		.INIT('h80)
	) name19039 (
		\m2_addr_i[13]_pad ,
		_w9171_,
		_w9172_,
		_w20940_
	);
	LUT4 #(
		.INIT('habef)
	) name19040 (
		_w9166_,
		_w9169_,
		_w20939_,
		_w20940_,
		_w20941_
	);
	LUT3 #(
		.INIT('h2a)
	) name19041 (
		\m5_addr_i[13]_pad ,
		_w9171_,
		_w9172_,
		_w20942_
	);
	LUT3 #(
		.INIT('h2a)
	) name19042 (
		\m1_addr_i[13]_pad ,
		_w9171_,
		_w9172_,
		_w20943_
	);
	LUT4 #(
		.INIT('h57df)
	) name19043 (
		_w9166_,
		_w9169_,
		_w20942_,
		_w20943_,
		_w20944_
	);
	LUT3 #(
		.INIT('h80)
	) name19044 (
		\m0_addr_i[13]_pad ,
		_w9171_,
		_w9172_,
		_w20945_
	);
	LUT3 #(
		.INIT('h2a)
	) name19045 (
		\m7_addr_i[13]_pad ,
		_w9171_,
		_w9172_,
		_w20946_
	);
	LUT4 #(
		.INIT('h6e7f)
	) name19046 (
		_w9166_,
		_w9169_,
		_w20945_,
		_w20946_,
		_w20947_
	);
	LUT4 #(
		.INIT('h7fff)
	) name19047 (
		_w20938_,
		_w20941_,
		_w20944_,
		_w20947_,
		_w20948_
	);
	LUT3 #(
		.INIT('h2a)
	) name19048 (
		\m3_addr_i[14]_pad ,
		_w9171_,
		_w9172_,
		_w20949_
	);
	LUT3 #(
		.INIT('h80)
	) name19049 (
		\m4_addr_i[14]_pad ,
		_w9171_,
		_w9172_,
		_w20950_
	);
	LUT4 #(
		.INIT('h9dbf)
	) name19050 (
		_w9166_,
		_w9169_,
		_w20949_,
		_w20950_,
		_w20951_
	);
	LUT3 #(
		.INIT('h80)
	) name19051 (
		\m6_addr_i[14]_pad ,
		_w9171_,
		_w9172_,
		_w20952_
	);
	LUT3 #(
		.INIT('h80)
	) name19052 (
		\m2_addr_i[14]_pad ,
		_w9171_,
		_w9172_,
		_w20953_
	);
	LUT4 #(
		.INIT('habef)
	) name19053 (
		_w9166_,
		_w9169_,
		_w20952_,
		_w20953_,
		_w20954_
	);
	LUT3 #(
		.INIT('h2a)
	) name19054 (
		\m5_addr_i[14]_pad ,
		_w9171_,
		_w9172_,
		_w20955_
	);
	LUT3 #(
		.INIT('h2a)
	) name19055 (
		\m1_addr_i[14]_pad ,
		_w9171_,
		_w9172_,
		_w20956_
	);
	LUT4 #(
		.INIT('h57df)
	) name19056 (
		_w9166_,
		_w9169_,
		_w20955_,
		_w20956_,
		_w20957_
	);
	LUT3 #(
		.INIT('h80)
	) name19057 (
		\m0_addr_i[14]_pad ,
		_w9171_,
		_w9172_,
		_w20958_
	);
	LUT3 #(
		.INIT('h2a)
	) name19058 (
		\m7_addr_i[14]_pad ,
		_w9171_,
		_w9172_,
		_w20959_
	);
	LUT4 #(
		.INIT('h6e7f)
	) name19059 (
		_w9166_,
		_w9169_,
		_w20958_,
		_w20959_,
		_w20960_
	);
	LUT4 #(
		.INIT('h7fff)
	) name19060 (
		_w20951_,
		_w20954_,
		_w20957_,
		_w20960_,
		_w20961_
	);
	LUT3 #(
		.INIT('h2a)
	) name19061 (
		\m3_addr_i[15]_pad ,
		_w9171_,
		_w9172_,
		_w20962_
	);
	LUT3 #(
		.INIT('h80)
	) name19062 (
		\m4_addr_i[15]_pad ,
		_w9171_,
		_w9172_,
		_w20963_
	);
	LUT4 #(
		.INIT('h9dbf)
	) name19063 (
		_w9166_,
		_w9169_,
		_w20962_,
		_w20963_,
		_w20964_
	);
	LUT3 #(
		.INIT('h80)
	) name19064 (
		\m6_addr_i[15]_pad ,
		_w9171_,
		_w9172_,
		_w20965_
	);
	LUT3 #(
		.INIT('h80)
	) name19065 (
		\m2_addr_i[15]_pad ,
		_w9171_,
		_w9172_,
		_w20966_
	);
	LUT4 #(
		.INIT('habef)
	) name19066 (
		_w9166_,
		_w9169_,
		_w20965_,
		_w20966_,
		_w20967_
	);
	LUT3 #(
		.INIT('h2a)
	) name19067 (
		\m5_addr_i[15]_pad ,
		_w9171_,
		_w9172_,
		_w20968_
	);
	LUT3 #(
		.INIT('h2a)
	) name19068 (
		\m1_addr_i[15]_pad ,
		_w9171_,
		_w9172_,
		_w20969_
	);
	LUT4 #(
		.INIT('h57df)
	) name19069 (
		_w9166_,
		_w9169_,
		_w20968_,
		_w20969_,
		_w20970_
	);
	LUT3 #(
		.INIT('h80)
	) name19070 (
		\m0_addr_i[15]_pad ,
		_w9171_,
		_w9172_,
		_w20971_
	);
	LUT3 #(
		.INIT('h2a)
	) name19071 (
		\m7_addr_i[15]_pad ,
		_w9171_,
		_w9172_,
		_w20972_
	);
	LUT4 #(
		.INIT('h6e7f)
	) name19072 (
		_w9166_,
		_w9169_,
		_w20971_,
		_w20972_,
		_w20973_
	);
	LUT4 #(
		.INIT('h7fff)
	) name19073 (
		_w20964_,
		_w20967_,
		_w20970_,
		_w20973_,
		_w20974_
	);
	LUT3 #(
		.INIT('h2a)
	) name19074 (
		\m3_addr_i[16]_pad ,
		_w9171_,
		_w9172_,
		_w20975_
	);
	LUT3 #(
		.INIT('h80)
	) name19075 (
		\m4_addr_i[16]_pad ,
		_w9171_,
		_w9172_,
		_w20976_
	);
	LUT4 #(
		.INIT('h9dbf)
	) name19076 (
		_w9166_,
		_w9169_,
		_w20975_,
		_w20976_,
		_w20977_
	);
	LUT3 #(
		.INIT('h80)
	) name19077 (
		\m6_addr_i[16]_pad ,
		_w9171_,
		_w9172_,
		_w20978_
	);
	LUT3 #(
		.INIT('h80)
	) name19078 (
		\m2_addr_i[16]_pad ,
		_w9171_,
		_w9172_,
		_w20979_
	);
	LUT4 #(
		.INIT('habef)
	) name19079 (
		_w9166_,
		_w9169_,
		_w20978_,
		_w20979_,
		_w20980_
	);
	LUT3 #(
		.INIT('h2a)
	) name19080 (
		\m5_addr_i[16]_pad ,
		_w9171_,
		_w9172_,
		_w20981_
	);
	LUT3 #(
		.INIT('h2a)
	) name19081 (
		\m1_addr_i[16]_pad ,
		_w9171_,
		_w9172_,
		_w20982_
	);
	LUT4 #(
		.INIT('h57df)
	) name19082 (
		_w9166_,
		_w9169_,
		_w20981_,
		_w20982_,
		_w20983_
	);
	LUT3 #(
		.INIT('h80)
	) name19083 (
		\m0_addr_i[16]_pad ,
		_w9171_,
		_w9172_,
		_w20984_
	);
	LUT3 #(
		.INIT('h2a)
	) name19084 (
		\m7_addr_i[16]_pad ,
		_w9171_,
		_w9172_,
		_w20985_
	);
	LUT4 #(
		.INIT('h6e7f)
	) name19085 (
		_w9166_,
		_w9169_,
		_w20984_,
		_w20985_,
		_w20986_
	);
	LUT4 #(
		.INIT('h7fff)
	) name19086 (
		_w20977_,
		_w20980_,
		_w20983_,
		_w20986_,
		_w20987_
	);
	LUT3 #(
		.INIT('h2a)
	) name19087 (
		\m3_addr_i[17]_pad ,
		_w9171_,
		_w9172_,
		_w20988_
	);
	LUT3 #(
		.INIT('h80)
	) name19088 (
		\m4_addr_i[17]_pad ,
		_w9171_,
		_w9172_,
		_w20989_
	);
	LUT4 #(
		.INIT('h9dbf)
	) name19089 (
		_w9166_,
		_w9169_,
		_w20988_,
		_w20989_,
		_w20990_
	);
	LUT3 #(
		.INIT('h80)
	) name19090 (
		\m6_addr_i[17]_pad ,
		_w9171_,
		_w9172_,
		_w20991_
	);
	LUT3 #(
		.INIT('h80)
	) name19091 (
		\m2_addr_i[17]_pad ,
		_w9171_,
		_w9172_,
		_w20992_
	);
	LUT4 #(
		.INIT('habef)
	) name19092 (
		_w9166_,
		_w9169_,
		_w20991_,
		_w20992_,
		_w20993_
	);
	LUT3 #(
		.INIT('h2a)
	) name19093 (
		\m5_addr_i[17]_pad ,
		_w9171_,
		_w9172_,
		_w20994_
	);
	LUT3 #(
		.INIT('h2a)
	) name19094 (
		\m1_addr_i[17]_pad ,
		_w9171_,
		_w9172_,
		_w20995_
	);
	LUT4 #(
		.INIT('h57df)
	) name19095 (
		_w9166_,
		_w9169_,
		_w20994_,
		_w20995_,
		_w20996_
	);
	LUT3 #(
		.INIT('h80)
	) name19096 (
		\m0_addr_i[17]_pad ,
		_w9171_,
		_w9172_,
		_w20997_
	);
	LUT3 #(
		.INIT('h2a)
	) name19097 (
		\m7_addr_i[17]_pad ,
		_w9171_,
		_w9172_,
		_w20998_
	);
	LUT4 #(
		.INIT('h6e7f)
	) name19098 (
		_w9166_,
		_w9169_,
		_w20997_,
		_w20998_,
		_w20999_
	);
	LUT4 #(
		.INIT('h7fff)
	) name19099 (
		_w20990_,
		_w20993_,
		_w20996_,
		_w20999_,
		_w21000_
	);
	LUT3 #(
		.INIT('h2a)
	) name19100 (
		\m3_addr_i[18]_pad ,
		_w9171_,
		_w9172_,
		_w21001_
	);
	LUT3 #(
		.INIT('h80)
	) name19101 (
		\m4_addr_i[18]_pad ,
		_w9171_,
		_w9172_,
		_w21002_
	);
	LUT4 #(
		.INIT('h9dbf)
	) name19102 (
		_w9166_,
		_w9169_,
		_w21001_,
		_w21002_,
		_w21003_
	);
	LUT3 #(
		.INIT('h80)
	) name19103 (
		\m6_addr_i[18]_pad ,
		_w9171_,
		_w9172_,
		_w21004_
	);
	LUT3 #(
		.INIT('h80)
	) name19104 (
		\m2_addr_i[18]_pad ,
		_w9171_,
		_w9172_,
		_w21005_
	);
	LUT4 #(
		.INIT('habef)
	) name19105 (
		_w9166_,
		_w9169_,
		_w21004_,
		_w21005_,
		_w21006_
	);
	LUT3 #(
		.INIT('h2a)
	) name19106 (
		\m5_addr_i[18]_pad ,
		_w9171_,
		_w9172_,
		_w21007_
	);
	LUT3 #(
		.INIT('h2a)
	) name19107 (
		\m1_addr_i[18]_pad ,
		_w9171_,
		_w9172_,
		_w21008_
	);
	LUT4 #(
		.INIT('h57df)
	) name19108 (
		_w9166_,
		_w9169_,
		_w21007_,
		_w21008_,
		_w21009_
	);
	LUT3 #(
		.INIT('h80)
	) name19109 (
		\m0_addr_i[18]_pad ,
		_w9171_,
		_w9172_,
		_w21010_
	);
	LUT3 #(
		.INIT('h2a)
	) name19110 (
		\m7_addr_i[18]_pad ,
		_w9171_,
		_w9172_,
		_w21011_
	);
	LUT4 #(
		.INIT('h6e7f)
	) name19111 (
		_w9166_,
		_w9169_,
		_w21010_,
		_w21011_,
		_w21012_
	);
	LUT4 #(
		.INIT('h7fff)
	) name19112 (
		_w21003_,
		_w21006_,
		_w21009_,
		_w21012_,
		_w21013_
	);
	LUT3 #(
		.INIT('h2a)
	) name19113 (
		\m3_addr_i[19]_pad ,
		_w9171_,
		_w9172_,
		_w21014_
	);
	LUT3 #(
		.INIT('h80)
	) name19114 (
		\m4_addr_i[19]_pad ,
		_w9171_,
		_w9172_,
		_w21015_
	);
	LUT4 #(
		.INIT('h9dbf)
	) name19115 (
		_w9166_,
		_w9169_,
		_w21014_,
		_w21015_,
		_w21016_
	);
	LUT3 #(
		.INIT('h80)
	) name19116 (
		\m6_addr_i[19]_pad ,
		_w9171_,
		_w9172_,
		_w21017_
	);
	LUT3 #(
		.INIT('h80)
	) name19117 (
		\m2_addr_i[19]_pad ,
		_w9171_,
		_w9172_,
		_w21018_
	);
	LUT4 #(
		.INIT('habef)
	) name19118 (
		_w9166_,
		_w9169_,
		_w21017_,
		_w21018_,
		_w21019_
	);
	LUT3 #(
		.INIT('h2a)
	) name19119 (
		\m5_addr_i[19]_pad ,
		_w9171_,
		_w9172_,
		_w21020_
	);
	LUT3 #(
		.INIT('h2a)
	) name19120 (
		\m1_addr_i[19]_pad ,
		_w9171_,
		_w9172_,
		_w21021_
	);
	LUT4 #(
		.INIT('h57df)
	) name19121 (
		_w9166_,
		_w9169_,
		_w21020_,
		_w21021_,
		_w21022_
	);
	LUT3 #(
		.INIT('h80)
	) name19122 (
		\m0_addr_i[19]_pad ,
		_w9171_,
		_w9172_,
		_w21023_
	);
	LUT3 #(
		.INIT('h2a)
	) name19123 (
		\m7_addr_i[19]_pad ,
		_w9171_,
		_w9172_,
		_w21024_
	);
	LUT4 #(
		.INIT('h6e7f)
	) name19124 (
		_w9166_,
		_w9169_,
		_w21023_,
		_w21024_,
		_w21025_
	);
	LUT4 #(
		.INIT('h7fff)
	) name19125 (
		_w21016_,
		_w21019_,
		_w21022_,
		_w21025_,
		_w21026_
	);
	LUT3 #(
		.INIT('h2a)
	) name19126 (
		\m3_addr_i[1]_pad ,
		_w9171_,
		_w9172_,
		_w21027_
	);
	LUT3 #(
		.INIT('h80)
	) name19127 (
		\m4_addr_i[1]_pad ,
		_w9171_,
		_w9172_,
		_w21028_
	);
	LUT4 #(
		.INIT('h9dbf)
	) name19128 (
		_w9166_,
		_w9169_,
		_w21027_,
		_w21028_,
		_w21029_
	);
	LUT3 #(
		.INIT('h80)
	) name19129 (
		\m6_addr_i[1]_pad ,
		_w9171_,
		_w9172_,
		_w21030_
	);
	LUT3 #(
		.INIT('h80)
	) name19130 (
		\m2_addr_i[1]_pad ,
		_w9171_,
		_w9172_,
		_w21031_
	);
	LUT4 #(
		.INIT('habef)
	) name19131 (
		_w9166_,
		_w9169_,
		_w21030_,
		_w21031_,
		_w21032_
	);
	LUT3 #(
		.INIT('h2a)
	) name19132 (
		\m5_addr_i[1]_pad ,
		_w9171_,
		_w9172_,
		_w21033_
	);
	LUT3 #(
		.INIT('h2a)
	) name19133 (
		\m1_addr_i[1]_pad ,
		_w9171_,
		_w9172_,
		_w21034_
	);
	LUT4 #(
		.INIT('h57df)
	) name19134 (
		_w9166_,
		_w9169_,
		_w21033_,
		_w21034_,
		_w21035_
	);
	LUT3 #(
		.INIT('h80)
	) name19135 (
		\m0_addr_i[1]_pad ,
		_w9171_,
		_w9172_,
		_w21036_
	);
	LUT3 #(
		.INIT('h2a)
	) name19136 (
		\m7_addr_i[1]_pad ,
		_w9171_,
		_w9172_,
		_w21037_
	);
	LUT4 #(
		.INIT('h6e7f)
	) name19137 (
		_w9166_,
		_w9169_,
		_w21036_,
		_w21037_,
		_w21038_
	);
	LUT4 #(
		.INIT('h7fff)
	) name19138 (
		_w21029_,
		_w21032_,
		_w21035_,
		_w21038_,
		_w21039_
	);
	LUT3 #(
		.INIT('h2a)
	) name19139 (
		\m3_addr_i[20]_pad ,
		_w9171_,
		_w9172_,
		_w21040_
	);
	LUT3 #(
		.INIT('h80)
	) name19140 (
		\m4_addr_i[20]_pad ,
		_w9171_,
		_w9172_,
		_w21041_
	);
	LUT4 #(
		.INIT('h9dbf)
	) name19141 (
		_w9166_,
		_w9169_,
		_w21040_,
		_w21041_,
		_w21042_
	);
	LUT3 #(
		.INIT('h80)
	) name19142 (
		\m6_addr_i[20]_pad ,
		_w9171_,
		_w9172_,
		_w21043_
	);
	LUT3 #(
		.INIT('h80)
	) name19143 (
		\m2_addr_i[20]_pad ,
		_w9171_,
		_w9172_,
		_w21044_
	);
	LUT4 #(
		.INIT('habef)
	) name19144 (
		_w9166_,
		_w9169_,
		_w21043_,
		_w21044_,
		_w21045_
	);
	LUT3 #(
		.INIT('h2a)
	) name19145 (
		\m5_addr_i[20]_pad ,
		_w9171_,
		_w9172_,
		_w21046_
	);
	LUT3 #(
		.INIT('h2a)
	) name19146 (
		\m1_addr_i[20]_pad ,
		_w9171_,
		_w9172_,
		_w21047_
	);
	LUT4 #(
		.INIT('h57df)
	) name19147 (
		_w9166_,
		_w9169_,
		_w21046_,
		_w21047_,
		_w21048_
	);
	LUT3 #(
		.INIT('h80)
	) name19148 (
		\m0_addr_i[20]_pad ,
		_w9171_,
		_w9172_,
		_w21049_
	);
	LUT3 #(
		.INIT('h2a)
	) name19149 (
		\m7_addr_i[20]_pad ,
		_w9171_,
		_w9172_,
		_w21050_
	);
	LUT4 #(
		.INIT('h6e7f)
	) name19150 (
		_w9166_,
		_w9169_,
		_w21049_,
		_w21050_,
		_w21051_
	);
	LUT4 #(
		.INIT('h7fff)
	) name19151 (
		_w21042_,
		_w21045_,
		_w21048_,
		_w21051_,
		_w21052_
	);
	LUT3 #(
		.INIT('h2a)
	) name19152 (
		\m3_addr_i[21]_pad ,
		_w9171_,
		_w9172_,
		_w21053_
	);
	LUT3 #(
		.INIT('h80)
	) name19153 (
		\m4_addr_i[21]_pad ,
		_w9171_,
		_w9172_,
		_w21054_
	);
	LUT4 #(
		.INIT('h9dbf)
	) name19154 (
		_w9166_,
		_w9169_,
		_w21053_,
		_w21054_,
		_w21055_
	);
	LUT3 #(
		.INIT('h80)
	) name19155 (
		\m6_addr_i[21]_pad ,
		_w9171_,
		_w9172_,
		_w21056_
	);
	LUT3 #(
		.INIT('h80)
	) name19156 (
		\m2_addr_i[21]_pad ,
		_w9171_,
		_w9172_,
		_w21057_
	);
	LUT4 #(
		.INIT('habef)
	) name19157 (
		_w9166_,
		_w9169_,
		_w21056_,
		_w21057_,
		_w21058_
	);
	LUT3 #(
		.INIT('h2a)
	) name19158 (
		\m5_addr_i[21]_pad ,
		_w9171_,
		_w9172_,
		_w21059_
	);
	LUT3 #(
		.INIT('h2a)
	) name19159 (
		\m1_addr_i[21]_pad ,
		_w9171_,
		_w9172_,
		_w21060_
	);
	LUT4 #(
		.INIT('h57df)
	) name19160 (
		_w9166_,
		_w9169_,
		_w21059_,
		_w21060_,
		_w21061_
	);
	LUT3 #(
		.INIT('h80)
	) name19161 (
		\m0_addr_i[21]_pad ,
		_w9171_,
		_w9172_,
		_w21062_
	);
	LUT3 #(
		.INIT('h2a)
	) name19162 (
		\m7_addr_i[21]_pad ,
		_w9171_,
		_w9172_,
		_w21063_
	);
	LUT4 #(
		.INIT('h6e7f)
	) name19163 (
		_w9166_,
		_w9169_,
		_w21062_,
		_w21063_,
		_w21064_
	);
	LUT4 #(
		.INIT('h7fff)
	) name19164 (
		_w21055_,
		_w21058_,
		_w21061_,
		_w21064_,
		_w21065_
	);
	LUT3 #(
		.INIT('h2a)
	) name19165 (
		\m3_addr_i[22]_pad ,
		_w9171_,
		_w9172_,
		_w21066_
	);
	LUT3 #(
		.INIT('h80)
	) name19166 (
		\m4_addr_i[22]_pad ,
		_w9171_,
		_w9172_,
		_w21067_
	);
	LUT4 #(
		.INIT('h9dbf)
	) name19167 (
		_w9166_,
		_w9169_,
		_w21066_,
		_w21067_,
		_w21068_
	);
	LUT3 #(
		.INIT('h80)
	) name19168 (
		\m6_addr_i[22]_pad ,
		_w9171_,
		_w9172_,
		_w21069_
	);
	LUT3 #(
		.INIT('h80)
	) name19169 (
		\m2_addr_i[22]_pad ,
		_w9171_,
		_w9172_,
		_w21070_
	);
	LUT4 #(
		.INIT('habef)
	) name19170 (
		_w9166_,
		_w9169_,
		_w21069_,
		_w21070_,
		_w21071_
	);
	LUT3 #(
		.INIT('h2a)
	) name19171 (
		\m5_addr_i[22]_pad ,
		_w9171_,
		_w9172_,
		_w21072_
	);
	LUT3 #(
		.INIT('h2a)
	) name19172 (
		\m1_addr_i[22]_pad ,
		_w9171_,
		_w9172_,
		_w21073_
	);
	LUT4 #(
		.INIT('h57df)
	) name19173 (
		_w9166_,
		_w9169_,
		_w21072_,
		_w21073_,
		_w21074_
	);
	LUT3 #(
		.INIT('h80)
	) name19174 (
		\m0_addr_i[22]_pad ,
		_w9171_,
		_w9172_,
		_w21075_
	);
	LUT3 #(
		.INIT('h2a)
	) name19175 (
		\m7_addr_i[22]_pad ,
		_w9171_,
		_w9172_,
		_w21076_
	);
	LUT4 #(
		.INIT('h6e7f)
	) name19176 (
		_w9166_,
		_w9169_,
		_w21075_,
		_w21076_,
		_w21077_
	);
	LUT4 #(
		.INIT('h7fff)
	) name19177 (
		_w21068_,
		_w21071_,
		_w21074_,
		_w21077_,
		_w21078_
	);
	LUT3 #(
		.INIT('h2a)
	) name19178 (
		\m3_addr_i[23]_pad ,
		_w9171_,
		_w9172_,
		_w21079_
	);
	LUT3 #(
		.INIT('h80)
	) name19179 (
		\m4_addr_i[23]_pad ,
		_w9171_,
		_w9172_,
		_w21080_
	);
	LUT4 #(
		.INIT('h9dbf)
	) name19180 (
		_w9166_,
		_w9169_,
		_w21079_,
		_w21080_,
		_w21081_
	);
	LUT3 #(
		.INIT('h80)
	) name19181 (
		\m6_addr_i[23]_pad ,
		_w9171_,
		_w9172_,
		_w21082_
	);
	LUT3 #(
		.INIT('h80)
	) name19182 (
		\m2_addr_i[23]_pad ,
		_w9171_,
		_w9172_,
		_w21083_
	);
	LUT4 #(
		.INIT('habef)
	) name19183 (
		_w9166_,
		_w9169_,
		_w21082_,
		_w21083_,
		_w21084_
	);
	LUT3 #(
		.INIT('h2a)
	) name19184 (
		\m5_addr_i[23]_pad ,
		_w9171_,
		_w9172_,
		_w21085_
	);
	LUT3 #(
		.INIT('h2a)
	) name19185 (
		\m1_addr_i[23]_pad ,
		_w9171_,
		_w9172_,
		_w21086_
	);
	LUT4 #(
		.INIT('h57df)
	) name19186 (
		_w9166_,
		_w9169_,
		_w21085_,
		_w21086_,
		_w21087_
	);
	LUT3 #(
		.INIT('h80)
	) name19187 (
		\m0_addr_i[23]_pad ,
		_w9171_,
		_w9172_,
		_w21088_
	);
	LUT3 #(
		.INIT('h2a)
	) name19188 (
		\m7_addr_i[23]_pad ,
		_w9171_,
		_w9172_,
		_w21089_
	);
	LUT4 #(
		.INIT('h6e7f)
	) name19189 (
		_w9166_,
		_w9169_,
		_w21088_,
		_w21089_,
		_w21090_
	);
	LUT4 #(
		.INIT('h7fff)
	) name19190 (
		_w21081_,
		_w21084_,
		_w21087_,
		_w21090_,
		_w21091_
	);
	LUT3 #(
		.INIT('h2a)
	) name19191 (
		\m3_addr_i[24]_pad ,
		_w9171_,
		_w9172_,
		_w21092_
	);
	LUT3 #(
		.INIT('h80)
	) name19192 (
		\m4_addr_i[24]_pad ,
		_w9171_,
		_w9172_,
		_w21093_
	);
	LUT4 #(
		.INIT('h9dbf)
	) name19193 (
		_w9166_,
		_w9169_,
		_w21092_,
		_w21093_,
		_w21094_
	);
	LUT3 #(
		.INIT('h2a)
	) name19194 (
		\m5_addr_i[24]_pad ,
		_w9171_,
		_w9172_,
		_w21095_
	);
	LUT3 #(
		.INIT('h80)
	) name19195 (
		\m2_addr_i[24]_pad ,
		_w9171_,
		_w9172_,
		_w21096_
	);
	LUT4 #(
		.INIT('h9bdf)
	) name19196 (
		_w9166_,
		_w9169_,
		_w21095_,
		_w21096_,
		_w21097_
	);
	LUT3 #(
		.INIT('h80)
	) name19197 (
		\m6_addr_i[24]_pad ,
		_w9171_,
		_w9172_,
		_w21098_
	);
	LUT3 #(
		.INIT('h2a)
	) name19198 (
		\m1_addr_i[24]_pad ,
		_w9171_,
		_w9172_,
		_w21099_
	);
	LUT4 #(
		.INIT('h67ef)
	) name19199 (
		_w9166_,
		_w9169_,
		_w21098_,
		_w21099_,
		_w21100_
	);
	LUT3 #(
		.INIT('h80)
	) name19200 (
		\m0_addr_i[24]_pad ,
		_w9171_,
		_w9172_,
		_w21101_
	);
	LUT3 #(
		.INIT('h2a)
	) name19201 (
		\m7_addr_i[24]_pad ,
		_w9171_,
		_w9172_,
		_w21102_
	);
	LUT4 #(
		.INIT('h6e7f)
	) name19202 (
		_w9166_,
		_w9169_,
		_w21101_,
		_w21102_,
		_w21103_
	);
	LUT4 #(
		.INIT('h7fff)
	) name19203 (
		_w21094_,
		_w21097_,
		_w21100_,
		_w21103_,
		_w21104_
	);
	LUT3 #(
		.INIT('h2a)
	) name19204 (
		\m3_addr_i[25]_pad ,
		_w9171_,
		_w9172_,
		_w21105_
	);
	LUT3 #(
		.INIT('h80)
	) name19205 (
		\m4_addr_i[25]_pad ,
		_w9171_,
		_w9172_,
		_w21106_
	);
	LUT4 #(
		.INIT('h9dbf)
	) name19206 (
		_w9166_,
		_w9169_,
		_w21105_,
		_w21106_,
		_w21107_
	);
	LUT3 #(
		.INIT('h2a)
	) name19207 (
		\m5_addr_i[25]_pad ,
		_w9171_,
		_w9172_,
		_w21108_
	);
	LUT3 #(
		.INIT('h80)
	) name19208 (
		\m2_addr_i[25]_pad ,
		_w9171_,
		_w9172_,
		_w21109_
	);
	LUT4 #(
		.INIT('h9bdf)
	) name19209 (
		_w9166_,
		_w9169_,
		_w21108_,
		_w21109_,
		_w21110_
	);
	LUT3 #(
		.INIT('h80)
	) name19210 (
		\m6_addr_i[25]_pad ,
		_w9171_,
		_w9172_,
		_w21111_
	);
	LUT3 #(
		.INIT('h2a)
	) name19211 (
		\m1_addr_i[25]_pad ,
		_w9171_,
		_w9172_,
		_w21112_
	);
	LUT4 #(
		.INIT('h67ef)
	) name19212 (
		_w9166_,
		_w9169_,
		_w21111_,
		_w21112_,
		_w21113_
	);
	LUT3 #(
		.INIT('h80)
	) name19213 (
		\m0_addr_i[25]_pad ,
		_w9171_,
		_w9172_,
		_w21114_
	);
	LUT3 #(
		.INIT('h2a)
	) name19214 (
		\m7_addr_i[25]_pad ,
		_w9171_,
		_w9172_,
		_w21115_
	);
	LUT4 #(
		.INIT('h6e7f)
	) name19215 (
		_w9166_,
		_w9169_,
		_w21114_,
		_w21115_,
		_w21116_
	);
	LUT4 #(
		.INIT('h7fff)
	) name19216 (
		_w21107_,
		_w21110_,
		_w21113_,
		_w21116_,
		_w21117_
	);
	LUT3 #(
		.INIT('h2a)
	) name19217 (
		\m3_addr_i[26]_pad ,
		_w9171_,
		_w9172_,
		_w21118_
	);
	LUT3 #(
		.INIT('h80)
	) name19218 (
		\m4_addr_i[26]_pad ,
		_w9171_,
		_w9172_,
		_w21119_
	);
	LUT4 #(
		.INIT('h9dbf)
	) name19219 (
		_w9166_,
		_w9169_,
		_w21118_,
		_w21119_,
		_w21120_
	);
	LUT3 #(
		.INIT('h2a)
	) name19220 (
		\m5_addr_i[26]_pad ,
		_w9171_,
		_w9172_,
		_w21121_
	);
	LUT3 #(
		.INIT('h80)
	) name19221 (
		\m2_addr_i[26]_pad ,
		_w9171_,
		_w9172_,
		_w21122_
	);
	LUT4 #(
		.INIT('h9bdf)
	) name19222 (
		_w9166_,
		_w9169_,
		_w21121_,
		_w21122_,
		_w21123_
	);
	LUT3 #(
		.INIT('h80)
	) name19223 (
		\m6_addr_i[26]_pad ,
		_w9171_,
		_w9172_,
		_w21124_
	);
	LUT3 #(
		.INIT('h2a)
	) name19224 (
		\m1_addr_i[26]_pad ,
		_w9171_,
		_w9172_,
		_w21125_
	);
	LUT4 #(
		.INIT('h67ef)
	) name19225 (
		_w9166_,
		_w9169_,
		_w21124_,
		_w21125_,
		_w21126_
	);
	LUT3 #(
		.INIT('h80)
	) name19226 (
		\m0_addr_i[26]_pad ,
		_w9171_,
		_w9172_,
		_w21127_
	);
	LUT3 #(
		.INIT('h2a)
	) name19227 (
		\m7_addr_i[26]_pad ,
		_w9171_,
		_w9172_,
		_w21128_
	);
	LUT4 #(
		.INIT('h6e7f)
	) name19228 (
		_w9166_,
		_w9169_,
		_w21127_,
		_w21128_,
		_w21129_
	);
	LUT4 #(
		.INIT('h7fff)
	) name19229 (
		_w21120_,
		_w21123_,
		_w21126_,
		_w21129_,
		_w21130_
	);
	LUT3 #(
		.INIT('h2a)
	) name19230 (
		\m3_addr_i[27]_pad ,
		_w9171_,
		_w9172_,
		_w21131_
	);
	LUT3 #(
		.INIT('h80)
	) name19231 (
		\m4_addr_i[27]_pad ,
		_w9171_,
		_w9172_,
		_w21132_
	);
	LUT4 #(
		.INIT('h9dbf)
	) name19232 (
		_w9166_,
		_w9169_,
		_w21131_,
		_w21132_,
		_w21133_
	);
	LUT3 #(
		.INIT('h2a)
	) name19233 (
		\m5_addr_i[27]_pad ,
		_w9171_,
		_w9172_,
		_w21134_
	);
	LUT3 #(
		.INIT('h80)
	) name19234 (
		\m2_addr_i[27]_pad ,
		_w9171_,
		_w9172_,
		_w21135_
	);
	LUT4 #(
		.INIT('h9bdf)
	) name19235 (
		_w9166_,
		_w9169_,
		_w21134_,
		_w21135_,
		_w21136_
	);
	LUT3 #(
		.INIT('h80)
	) name19236 (
		\m6_addr_i[27]_pad ,
		_w9171_,
		_w9172_,
		_w21137_
	);
	LUT3 #(
		.INIT('h2a)
	) name19237 (
		\m1_addr_i[27]_pad ,
		_w9171_,
		_w9172_,
		_w21138_
	);
	LUT4 #(
		.INIT('h67ef)
	) name19238 (
		_w9166_,
		_w9169_,
		_w21137_,
		_w21138_,
		_w21139_
	);
	LUT3 #(
		.INIT('h80)
	) name19239 (
		\m0_addr_i[27]_pad ,
		_w9171_,
		_w9172_,
		_w21140_
	);
	LUT3 #(
		.INIT('h2a)
	) name19240 (
		\m7_addr_i[27]_pad ,
		_w9171_,
		_w9172_,
		_w21141_
	);
	LUT4 #(
		.INIT('h6e7f)
	) name19241 (
		_w9166_,
		_w9169_,
		_w21140_,
		_w21141_,
		_w21142_
	);
	LUT4 #(
		.INIT('h7fff)
	) name19242 (
		_w21133_,
		_w21136_,
		_w21139_,
		_w21142_,
		_w21143_
	);
	LUT3 #(
		.INIT('h2a)
	) name19243 (
		\m3_addr_i[28]_pad ,
		_w9171_,
		_w9172_,
		_w21144_
	);
	LUT3 #(
		.INIT('h80)
	) name19244 (
		\m4_addr_i[28]_pad ,
		_w9171_,
		_w9172_,
		_w21145_
	);
	LUT4 #(
		.INIT('h9dbf)
	) name19245 (
		_w9166_,
		_w9169_,
		_w21144_,
		_w21145_,
		_w21146_
	);
	LUT3 #(
		.INIT('h2a)
	) name19246 (
		\m5_addr_i[28]_pad ,
		_w9171_,
		_w9172_,
		_w21147_
	);
	LUT3 #(
		.INIT('h80)
	) name19247 (
		\m2_addr_i[28]_pad ,
		_w9171_,
		_w9172_,
		_w21148_
	);
	LUT4 #(
		.INIT('h9bdf)
	) name19248 (
		_w9166_,
		_w9169_,
		_w21147_,
		_w21148_,
		_w21149_
	);
	LUT3 #(
		.INIT('h80)
	) name19249 (
		\m6_addr_i[28]_pad ,
		_w9171_,
		_w9172_,
		_w21150_
	);
	LUT3 #(
		.INIT('h2a)
	) name19250 (
		\m1_addr_i[28]_pad ,
		_w9171_,
		_w9172_,
		_w21151_
	);
	LUT4 #(
		.INIT('h67ef)
	) name19251 (
		_w9166_,
		_w9169_,
		_w21150_,
		_w21151_,
		_w21152_
	);
	LUT3 #(
		.INIT('h80)
	) name19252 (
		\m0_addr_i[28]_pad ,
		_w9171_,
		_w9172_,
		_w21153_
	);
	LUT3 #(
		.INIT('h2a)
	) name19253 (
		\m7_addr_i[28]_pad ,
		_w9171_,
		_w9172_,
		_w21154_
	);
	LUT4 #(
		.INIT('h6e7f)
	) name19254 (
		_w9166_,
		_w9169_,
		_w21153_,
		_w21154_,
		_w21155_
	);
	LUT4 #(
		.INIT('h7fff)
	) name19255 (
		_w21146_,
		_w21149_,
		_w21152_,
		_w21155_,
		_w21156_
	);
	LUT3 #(
		.INIT('h2a)
	) name19256 (
		\m3_addr_i[29]_pad ,
		_w9171_,
		_w9172_,
		_w21157_
	);
	LUT3 #(
		.INIT('h80)
	) name19257 (
		\m4_addr_i[29]_pad ,
		_w9171_,
		_w9172_,
		_w21158_
	);
	LUT4 #(
		.INIT('h9dbf)
	) name19258 (
		_w9166_,
		_w9169_,
		_w21157_,
		_w21158_,
		_w21159_
	);
	LUT3 #(
		.INIT('h2a)
	) name19259 (
		\m5_addr_i[29]_pad ,
		_w9171_,
		_w9172_,
		_w21160_
	);
	LUT3 #(
		.INIT('h80)
	) name19260 (
		\m2_addr_i[29]_pad ,
		_w9171_,
		_w9172_,
		_w21161_
	);
	LUT4 #(
		.INIT('h9bdf)
	) name19261 (
		_w9166_,
		_w9169_,
		_w21160_,
		_w21161_,
		_w21162_
	);
	LUT3 #(
		.INIT('h80)
	) name19262 (
		\m6_addr_i[29]_pad ,
		_w9171_,
		_w9172_,
		_w21163_
	);
	LUT3 #(
		.INIT('h2a)
	) name19263 (
		\m1_addr_i[29]_pad ,
		_w9171_,
		_w9172_,
		_w21164_
	);
	LUT4 #(
		.INIT('h67ef)
	) name19264 (
		_w9166_,
		_w9169_,
		_w21163_,
		_w21164_,
		_w21165_
	);
	LUT3 #(
		.INIT('h80)
	) name19265 (
		\m0_addr_i[29]_pad ,
		_w9171_,
		_w9172_,
		_w21166_
	);
	LUT3 #(
		.INIT('h2a)
	) name19266 (
		\m7_addr_i[29]_pad ,
		_w9171_,
		_w9172_,
		_w21167_
	);
	LUT4 #(
		.INIT('h6e7f)
	) name19267 (
		_w9166_,
		_w9169_,
		_w21166_,
		_w21167_,
		_w21168_
	);
	LUT4 #(
		.INIT('h7fff)
	) name19268 (
		_w21159_,
		_w21162_,
		_w21165_,
		_w21168_,
		_w21169_
	);
	LUT3 #(
		.INIT('h2a)
	) name19269 (
		\m3_addr_i[2]_pad ,
		_w9171_,
		_w9172_,
		_w21170_
	);
	LUT3 #(
		.INIT('h80)
	) name19270 (
		\m4_addr_i[2]_pad ,
		_w9171_,
		_w9172_,
		_w21171_
	);
	LUT4 #(
		.INIT('h9dbf)
	) name19271 (
		_w9166_,
		_w9169_,
		_w21170_,
		_w21171_,
		_w21172_
	);
	LUT3 #(
		.INIT('h80)
	) name19272 (
		\m6_addr_i[2]_pad ,
		_w9171_,
		_w9172_,
		_w21173_
	);
	LUT3 #(
		.INIT('h80)
	) name19273 (
		\m2_addr_i[2]_pad ,
		_w9171_,
		_w9172_,
		_w21174_
	);
	LUT4 #(
		.INIT('habef)
	) name19274 (
		_w9166_,
		_w9169_,
		_w21173_,
		_w21174_,
		_w21175_
	);
	LUT3 #(
		.INIT('h2a)
	) name19275 (
		\m5_addr_i[2]_pad ,
		_w9171_,
		_w9172_,
		_w21176_
	);
	LUT3 #(
		.INIT('h2a)
	) name19276 (
		\m1_addr_i[2]_pad ,
		_w9171_,
		_w9172_,
		_w21177_
	);
	LUT4 #(
		.INIT('h57df)
	) name19277 (
		_w9166_,
		_w9169_,
		_w21176_,
		_w21177_,
		_w21178_
	);
	LUT3 #(
		.INIT('h80)
	) name19278 (
		\m0_addr_i[2]_pad ,
		_w9171_,
		_w9172_,
		_w21179_
	);
	LUT3 #(
		.INIT('h2a)
	) name19279 (
		\m7_addr_i[2]_pad ,
		_w9171_,
		_w9172_,
		_w21180_
	);
	LUT4 #(
		.INIT('h6e7f)
	) name19280 (
		_w9166_,
		_w9169_,
		_w21179_,
		_w21180_,
		_w21181_
	);
	LUT4 #(
		.INIT('h7fff)
	) name19281 (
		_w21172_,
		_w21175_,
		_w21178_,
		_w21181_,
		_w21182_
	);
	LUT3 #(
		.INIT('h2a)
	) name19282 (
		\m3_addr_i[30]_pad ,
		_w9171_,
		_w9172_,
		_w21183_
	);
	LUT3 #(
		.INIT('h80)
	) name19283 (
		\m4_addr_i[30]_pad ,
		_w9171_,
		_w9172_,
		_w21184_
	);
	LUT4 #(
		.INIT('h9dbf)
	) name19284 (
		_w9166_,
		_w9169_,
		_w21183_,
		_w21184_,
		_w21185_
	);
	LUT3 #(
		.INIT('h2a)
	) name19285 (
		\m5_addr_i[30]_pad ,
		_w9171_,
		_w9172_,
		_w21186_
	);
	LUT3 #(
		.INIT('h80)
	) name19286 (
		\m2_addr_i[30]_pad ,
		_w9171_,
		_w9172_,
		_w21187_
	);
	LUT4 #(
		.INIT('h9bdf)
	) name19287 (
		_w9166_,
		_w9169_,
		_w21186_,
		_w21187_,
		_w21188_
	);
	LUT3 #(
		.INIT('h80)
	) name19288 (
		\m6_addr_i[30]_pad ,
		_w9171_,
		_w9172_,
		_w21189_
	);
	LUT3 #(
		.INIT('h2a)
	) name19289 (
		\m1_addr_i[30]_pad ,
		_w9171_,
		_w9172_,
		_w21190_
	);
	LUT4 #(
		.INIT('h67ef)
	) name19290 (
		_w9166_,
		_w9169_,
		_w21189_,
		_w21190_,
		_w21191_
	);
	LUT3 #(
		.INIT('h80)
	) name19291 (
		\m0_addr_i[30]_pad ,
		_w9171_,
		_w9172_,
		_w21192_
	);
	LUT3 #(
		.INIT('h2a)
	) name19292 (
		\m7_addr_i[30]_pad ,
		_w9171_,
		_w9172_,
		_w21193_
	);
	LUT4 #(
		.INIT('h6e7f)
	) name19293 (
		_w9166_,
		_w9169_,
		_w21192_,
		_w21193_,
		_w21194_
	);
	LUT4 #(
		.INIT('h7fff)
	) name19294 (
		_w21185_,
		_w21188_,
		_w21191_,
		_w21194_,
		_w21195_
	);
	LUT3 #(
		.INIT('h2a)
	) name19295 (
		\m3_addr_i[31]_pad ,
		_w9171_,
		_w9172_,
		_w21196_
	);
	LUT3 #(
		.INIT('h80)
	) name19296 (
		\m4_addr_i[31]_pad ,
		_w9171_,
		_w9172_,
		_w21197_
	);
	LUT4 #(
		.INIT('h9dbf)
	) name19297 (
		_w9166_,
		_w9169_,
		_w21196_,
		_w21197_,
		_w21198_
	);
	LUT3 #(
		.INIT('h2a)
	) name19298 (
		\m5_addr_i[31]_pad ,
		_w9171_,
		_w9172_,
		_w21199_
	);
	LUT3 #(
		.INIT('h80)
	) name19299 (
		\m2_addr_i[31]_pad ,
		_w9171_,
		_w9172_,
		_w21200_
	);
	LUT4 #(
		.INIT('h9bdf)
	) name19300 (
		_w9166_,
		_w9169_,
		_w21199_,
		_w21200_,
		_w21201_
	);
	LUT3 #(
		.INIT('h80)
	) name19301 (
		\m6_addr_i[31]_pad ,
		_w9171_,
		_w9172_,
		_w21202_
	);
	LUT3 #(
		.INIT('h2a)
	) name19302 (
		\m1_addr_i[31]_pad ,
		_w9171_,
		_w9172_,
		_w21203_
	);
	LUT4 #(
		.INIT('h67ef)
	) name19303 (
		_w9166_,
		_w9169_,
		_w21202_,
		_w21203_,
		_w21204_
	);
	LUT3 #(
		.INIT('h80)
	) name19304 (
		\m0_addr_i[31]_pad ,
		_w9171_,
		_w9172_,
		_w21205_
	);
	LUT3 #(
		.INIT('h2a)
	) name19305 (
		\m7_addr_i[31]_pad ,
		_w9171_,
		_w9172_,
		_w21206_
	);
	LUT4 #(
		.INIT('h6e7f)
	) name19306 (
		_w9166_,
		_w9169_,
		_w21205_,
		_w21206_,
		_w21207_
	);
	LUT4 #(
		.INIT('h7fff)
	) name19307 (
		_w21198_,
		_w21201_,
		_w21204_,
		_w21207_,
		_w21208_
	);
	LUT3 #(
		.INIT('h2a)
	) name19308 (
		\m3_addr_i[3]_pad ,
		_w9171_,
		_w9172_,
		_w21209_
	);
	LUT3 #(
		.INIT('h80)
	) name19309 (
		\m4_addr_i[3]_pad ,
		_w9171_,
		_w9172_,
		_w21210_
	);
	LUT4 #(
		.INIT('h9dbf)
	) name19310 (
		_w9166_,
		_w9169_,
		_w21209_,
		_w21210_,
		_w21211_
	);
	LUT3 #(
		.INIT('h80)
	) name19311 (
		\m6_addr_i[3]_pad ,
		_w9171_,
		_w9172_,
		_w21212_
	);
	LUT3 #(
		.INIT('h80)
	) name19312 (
		\m2_addr_i[3]_pad ,
		_w9171_,
		_w9172_,
		_w21213_
	);
	LUT4 #(
		.INIT('habef)
	) name19313 (
		_w9166_,
		_w9169_,
		_w21212_,
		_w21213_,
		_w21214_
	);
	LUT3 #(
		.INIT('h2a)
	) name19314 (
		\m5_addr_i[3]_pad ,
		_w9171_,
		_w9172_,
		_w21215_
	);
	LUT3 #(
		.INIT('h2a)
	) name19315 (
		\m1_addr_i[3]_pad ,
		_w9171_,
		_w9172_,
		_w21216_
	);
	LUT4 #(
		.INIT('h57df)
	) name19316 (
		_w9166_,
		_w9169_,
		_w21215_,
		_w21216_,
		_w21217_
	);
	LUT3 #(
		.INIT('h80)
	) name19317 (
		\m0_addr_i[3]_pad ,
		_w9171_,
		_w9172_,
		_w21218_
	);
	LUT3 #(
		.INIT('h2a)
	) name19318 (
		\m7_addr_i[3]_pad ,
		_w9171_,
		_w9172_,
		_w21219_
	);
	LUT4 #(
		.INIT('h6e7f)
	) name19319 (
		_w9166_,
		_w9169_,
		_w21218_,
		_w21219_,
		_w21220_
	);
	LUT4 #(
		.INIT('h7fff)
	) name19320 (
		_w21211_,
		_w21214_,
		_w21217_,
		_w21220_,
		_w21221_
	);
	LUT3 #(
		.INIT('h2a)
	) name19321 (
		\m3_addr_i[4]_pad ,
		_w9171_,
		_w9172_,
		_w21222_
	);
	LUT3 #(
		.INIT('h80)
	) name19322 (
		\m4_addr_i[4]_pad ,
		_w9171_,
		_w9172_,
		_w21223_
	);
	LUT4 #(
		.INIT('h9dbf)
	) name19323 (
		_w9166_,
		_w9169_,
		_w21222_,
		_w21223_,
		_w21224_
	);
	LUT3 #(
		.INIT('h80)
	) name19324 (
		\m6_addr_i[4]_pad ,
		_w9171_,
		_w9172_,
		_w21225_
	);
	LUT3 #(
		.INIT('h80)
	) name19325 (
		\m2_addr_i[4]_pad ,
		_w9171_,
		_w9172_,
		_w21226_
	);
	LUT4 #(
		.INIT('habef)
	) name19326 (
		_w9166_,
		_w9169_,
		_w21225_,
		_w21226_,
		_w21227_
	);
	LUT3 #(
		.INIT('h2a)
	) name19327 (
		\m5_addr_i[4]_pad ,
		_w9171_,
		_w9172_,
		_w21228_
	);
	LUT3 #(
		.INIT('h2a)
	) name19328 (
		\m1_addr_i[4]_pad ,
		_w9171_,
		_w9172_,
		_w21229_
	);
	LUT4 #(
		.INIT('h57df)
	) name19329 (
		_w9166_,
		_w9169_,
		_w21228_,
		_w21229_,
		_w21230_
	);
	LUT3 #(
		.INIT('h80)
	) name19330 (
		\m0_addr_i[4]_pad ,
		_w9171_,
		_w9172_,
		_w21231_
	);
	LUT3 #(
		.INIT('h2a)
	) name19331 (
		\m7_addr_i[4]_pad ,
		_w9171_,
		_w9172_,
		_w21232_
	);
	LUT4 #(
		.INIT('h6e7f)
	) name19332 (
		_w9166_,
		_w9169_,
		_w21231_,
		_w21232_,
		_w21233_
	);
	LUT4 #(
		.INIT('h7fff)
	) name19333 (
		_w21224_,
		_w21227_,
		_w21230_,
		_w21233_,
		_w21234_
	);
	LUT3 #(
		.INIT('h2a)
	) name19334 (
		\m3_addr_i[5]_pad ,
		_w9171_,
		_w9172_,
		_w21235_
	);
	LUT3 #(
		.INIT('h80)
	) name19335 (
		\m4_addr_i[5]_pad ,
		_w9171_,
		_w9172_,
		_w21236_
	);
	LUT4 #(
		.INIT('h9dbf)
	) name19336 (
		_w9166_,
		_w9169_,
		_w21235_,
		_w21236_,
		_w21237_
	);
	LUT3 #(
		.INIT('h80)
	) name19337 (
		\m6_addr_i[5]_pad ,
		_w9171_,
		_w9172_,
		_w21238_
	);
	LUT3 #(
		.INIT('h80)
	) name19338 (
		\m2_addr_i[5]_pad ,
		_w9171_,
		_w9172_,
		_w21239_
	);
	LUT4 #(
		.INIT('habef)
	) name19339 (
		_w9166_,
		_w9169_,
		_w21238_,
		_w21239_,
		_w21240_
	);
	LUT3 #(
		.INIT('h2a)
	) name19340 (
		\m5_addr_i[5]_pad ,
		_w9171_,
		_w9172_,
		_w21241_
	);
	LUT3 #(
		.INIT('h2a)
	) name19341 (
		\m1_addr_i[5]_pad ,
		_w9171_,
		_w9172_,
		_w21242_
	);
	LUT4 #(
		.INIT('h57df)
	) name19342 (
		_w9166_,
		_w9169_,
		_w21241_,
		_w21242_,
		_w21243_
	);
	LUT3 #(
		.INIT('h80)
	) name19343 (
		\m0_addr_i[5]_pad ,
		_w9171_,
		_w9172_,
		_w21244_
	);
	LUT3 #(
		.INIT('h2a)
	) name19344 (
		\m7_addr_i[5]_pad ,
		_w9171_,
		_w9172_,
		_w21245_
	);
	LUT4 #(
		.INIT('h6e7f)
	) name19345 (
		_w9166_,
		_w9169_,
		_w21244_,
		_w21245_,
		_w21246_
	);
	LUT4 #(
		.INIT('h7fff)
	) name19346 (
		_w21237_,
		_w21240_,
		_w21243_,
		_w21246_,
		_w21247_
	);
	LUT3 #(
		.INIT('h2a)
	) name19347 (
		\m3_addr_i[6]_pad ,
		_w9171_,
		_w9172_,
		_w21248_
	);
	LUT3 #(
		.INIT('h80)
	) name19348 (
		\m4_addr_i[6]_pad ,
		_w9171_,
		_w9172_,
		_w21249_
	);
	LUT4 #(
		.INIT('h9dbf)
	) name19349 (
		_w9166_,
		_w9169_,
		_w21248_,
		_w21249_,
		_w21250_
	);
	LUT3 #(
		.INIT('h80)
	) name19350 (
		\m6_addr_i[6]_pad ,
		_w9171_,
		_w9172_,
		_w21251_
	);
	LUT3 #(
		.INIT('h80)
	) name19351 (
		\m2_addr_i[6]_pad ,
		_w9171_,
		_w9172_,
		_w21252_
	);
	LUT4 #(
		.INIT('habef)
	) name19352 (
		_w9166_,
		_w9169_,
		_w21251_,
		_w21252_,
		_w21253_
	);
	LUT3 #(
		.INIT('h2a)
	) name19353 (
		\m5_addr_i[6]_pad ,
		_w9171_,
		_w9172_,
		_w21254_
	);
	LUT3 #(
		.INIT('h2a)
	) name19354 (
		\m1_addr_i[6]_pad ,
		_w9171_,
		_w9172_,
		_w21255_
	);
	LUT4 #(
		.INIT('h57df)
	) name19355 (
		_w9166_,
		_w9169_,
		_w21254_,
		_w21255_,
		_w21256_
	);
	LUT3 #(
		.INIT('h80)
	) name19356 (
		\m0_addr_i[6]_pad ,
		_w9171_,
		_w9172_,
		_w21257_
	);
	LUT3 #(
		.INIT('h2a)
	) name19357 (
		\m7_addr_i[6]_pad ,
		_w9171_,
		_w9172_,
		_w21258_
	);
	LUT4 #(
		.INIT('h6e7f)
	) name19358 (
		_w9166_,
		_w9169_,
		_w21257_,
		_w21258_,
		_w21259_
	);
	LUT4 #(
		.INIT('h7fff)
	) name19359 (
		_w21250_,
		_w21253_,
		_w21256_,
		_w21259_,
		_w21260_
	);
	LUT3 #(
		.INIT('h2a)
	) name19360 (
		\m3_addr_i[7]_pad ,
		_w9171_,
		_w9172_,
		_w21261_
	);
	LUT3 #(
		.INIT('h80)
	) name19361 (
		\m4_addr_i[7]_pad ,
		_w9171_,
		_w9172_,
		_w21262_
	);
	LUT4 #(
		.INIT('h9dbf)
	) name19362 (
		_w9166_,
		_w9169_,
		_w21261_,
		_w21262_,
		_w21263_
	);
	LUT3 #(
		.INIT('h80)
	) name19363 (
		\m6_addr_i[7]_pad ,
		_w9171_,
		_w9172_,
		_w21264_
	);
	LUT3 #(
		.INIT('h80)
	) name19364 (
		\m2_addr_i[7]_pad ,
		_w9171_,
		_w9172_,
		_w21265_
	);
	LUT4 #(
		.INIT('habef)
	) name19365 (
		_w9166_,
		_w9169_,
		_w21264_,
		_w21265_,
		_w21266_
	);
	LUT3 #(
		.INIT('h2a)
	) name19366 (
		\m5_addr_i[7]_pad ,
		_w9171_,
		_w9172_,
		_w21267_
	);
	LUT3 #(
		.INIT('h2a)
	) name19367 (
		\m1_addr_i[7]_pad ,
		_w9171_,
		_w9172_,
		_w21268_
	);
	LUT4 #(
		.INIT('h57df)
	) name19368 (
		_w9166_,
		_w9169_,
		_w21267_,
		_w21268_,
		_w21269_
	);
	LUT3 #(
		.INIT('h80)
	) name19369 (
		\m0_addr_i[7]_pad ,
		_w9171_,
		_w9172_,
		_w21270_
	);
	LUT3 #(
		.INIT('h2a)
	) name19370 (
		\m7_addr_i[7]_pad ,
		_w9171_,
		_w9172_,
		_w21271_
	);
	LUT4 #(
		.INIT('h6e7f)
	) name19371 (
		_w9166_,
		_w9169_,
		_w21270_,
		_w21271_,
		_w21272_
	);
	LUT4 #(
		.INIT('h7fff)
	) name19372 (
		_w21263_,
		_w21266_,
		_w21269_,
		_w21272_,
		_w21273_
	);
	LUT3 #(
		.INIT('h2a)
	) name19373 (
		\m3_addr_i[8]_pad ,
		_w9171_,
		_w9172_,
		_w21274_
	);
	LUT3 #(
		.INIT('h80)
	) name19374 (
		\m4_addr_i[8]_pad ,
		_w9171_,
		_w9172_,
		_w21275_
	);
	LUT4 #(
		.INIT('h9dbf)
	) name19375 (
		_w9166_,
		_w9169_,
		_w21274_,
		_w21275_,
		_w21276_
	);
	LUT3 #(
		.INIT('h80)
	) name19376 (
		\m6_addr_i[8]_pad ,
		_w9171_,
		_w9172_,
		_w21277_
	);
	LUT3 #(
		.INIT('h80)
	) name19377 (
		\m2_addr_i[8]_pad ,
		_w9171_,
		_w9172_,
		_w21278_
	);
	LUT4 #(
		.INIT('habef)
	) name19378 (
		_w9166_,
		_w9169_,
		_w21277_,
		_w21278_,
		_w21279_
	);
	LUT3 #(
		.INIT('h2a)
	) name19379 (
		\m5_addr_i[8]_pad ,
		_w9171_,
		_w9172_,
		_w21280_
	);
	LUT3 #(
		.INIT('h2a)
	) name19380 (
		\m1_addr_i[8]_pad ,
		_w9171_,
		_w9172_,
		_w21281_
	);
	LUT4 #(
		.INIT('h57df)
	) name19381 (
		_w9166_,
		_w9169_,
		_w21280_,
		_w21281_,
		_w21282_
	);
	LUT3 #(
		.INIT('h80)
	) name19382 (
		\m0_addr_i[8]_pad ,
		_w9171_,
		_w9172_,
		_w21283_
	);
	LUT3 #(
		.INIT('h2a)
	) name19383 (
		\m7_addr_i[8]_pad ,
		_w9171_,
		_w9172_,
		_w21284_
	);
	LUT4 #(
		.INIT('h6e7f)
	) name19384 (
		_w9166_,
		_w9169_,
		_w21283_,
		_w21284_,
		_w21285_
	);
	LUT4 #(
		.INIT('h7fff)
	) name19385 (
		_w21276_,
		_w21279_,
		_w21282_,
		_w21285_,
		_w21286_
	);
	LUT3 #(
		.INIT('h2a)
	) name19386 (
		\m3_addr_i[9]_pad ,
		_w9171_,
		_w9172_,
		_w21287_
	);
	LUT3 #(
		.INIT('h80)
	) name19387 (
		\m4_addr_i[9]_pad ,
		_w9171_,
		_w9172_,
		_w21288_
	);
	LUT4 #(
		.INIT('h9dbf)
	) name19388 (
		_w9166_,
		_w9169_,
		_w21287_,
		_w21288_,
		_w21289_
	);
	LUT3 #(
		.INIT('h80)
	) name19389 (
		\m6_addr_i[9]_pad ,
		_w9171_,
		_w9172_,
		_w21290_
	);
	LUT3 #(
		.INIT('h80)
	) name19390 (
		\m2_addr_i[9]_pad ,
		_w9171_,
		_w9172_,
		_w21291_
	);
	LUT4 #(
		.INIT('habef)
	) name19391 (
		_w9166_,
		_w9169_,
		_w21290_,
		_w21291_,
		_w21292_
	);
	LUT3 #(
		.INIT('h2a)
	) name19392 (
		\m5_addr_i[9]_pad ,
		_w9171_,
		_w9172_,
		_w21293_
	);
	LUT3 #(
		.INIT('h2a)
	) name19393 (
		\m1_addr_i[9]_pad ,
		_w9171_,
		_w9172_,
		_w21294_
	);
	LUT4 #(
		.INIT('h57df)
	) name19394 (
		_w9166_,
		_w9169_,
		_w21293_,
		_w21294_,
		_w21295_
	);
	LUT3 #(
		.INIT('h80)
	) name19395 (
		\m0_addr_i[9]_pad ,
		_w9171_,
		_w9172_,
		_w21296_
	);
	LUT3 #(
		.INIT('h2a)
	) name19396 (
		\m7_addr_i[9]_pad ,
		_w9171_,
		_w9172_,
		_w21297_
	);
	LUT4 #(
		.INIT('h6e7f)
	) name19397 (
		_w9166_,
		_w9169_,
		_w21296_,
		_w21297_,
		_w21298_
	);
	LUT4 #(
		.INIT('h7fff)
	) name19398 (
		_w21289_,
		_w21292_,
		_w21295_,
		_w21298_,
		_w21299_
	);
	LUT3 #(
		.INIT('h2a)
	) name19399 (
		\m3_data_i[0]_pad ,
		_w9171_,
		_w9172_,
		_w21300_
	);
	LUT3 #(
		.INIT('h80)
	) name19400 (
		\m4_data_i[0]_pad ,
		_w9171_,
		_w9172_,
		_w21301_
	);
	LUT4 #(
		.INIT('h9dbf)
	) name19401 (
		_w9166_,
		_w9169_,
		_w21300_,
		_w21301_,
		_w21302_
	);
	LUT3 #(
		.INIT('h80)
	) name19402 (
		\m6_data_i[0]_pad ,
		_w9171_,
		_w9172_,
		_w21303_
	);
	LUT3 #(
		.INIT('h80)
	) name19403 (
		\m2_data_i[0]_pad ,
		_w9171_,
		_w9172_,
		_w21304_
	);
	LUT4 #(
		.INIT('habef)
	) name19404 (
		_w9166_,
		_w9169_,
		_w21303_,
		_w21304_,
		_w21305_
	);
	LUT3 #(
		.INIT('h2a)
	) name19405 (
		\m5_data_i[0]_pad ,
		_w9171_,
		_w9172_,
		_w21306_
	);
	LUT3 #(
		.INIT('h2a)
	) name19406 (
		\m1_data_i[0]_pad ,
		_w9171_,
		_w9172_,
		_w21307_
	);
	LUT4 #(
		.INIT('h57df)
	) name19407 (
		_w9166_,
		_w9169_,
		_w21306_,
		_w21307_,
		_w21308_
	);
	LUT3 #(
		.INIT('h80)
	) name19408 (
		\m0_data_i[0]_pad ,
		_w9171_,
		_w9172_,
		_w21309_
	);
	LUT3 #(
		.INIT('h2a)
	) name19409 (
		\m7_data_i[0]_pad ,
		_w9171_,
		_w9172_,
		_w21310_
	);
	LUT4 #(
		.INIT('h6e7f)
	) name19410 (
		_w9166_,
		_w9169_,
		_w21309_,
		_w21310_,
		_w21311_
	);
	LUT4 #(
		.INIT('h7fff)
	) name19411 (
		_w21302_,
		_w21305_,
		_w21308_,
		_w21311_,
		_w21312_
	);
	LUT3 #(
		.INIT('h2a)
	) name19412 (
		\m3_data_i[10]_pad ,
		_w9171_,
		_w9172_,
		_w21313_
	);
	LUT3 #(
		.INIT('h80)
	) name19413 (
		\m4_data_i[10]_pad ,
		_w9171_,
		_w9172_,
		_w21314_
	);
	LUT4 #(
		.INIT('h9dbf)
	) name19414 (
		_w9166_,
		_w9169_,
		_w21313_,
		_w21314_,
		_w21315_
	);
	LUT3 #(
		.INIT('h80)
	) name19415 (
		\m6_data_i[10]_pad ,
		_w9171_,
		_w9172_,
		_w21316_
	);
	LUT3 #(
		.INIT('h80)
	) name19416 (
		\m2_data_i[10]_pad ,
		_w9171_,
		_w9172_,
		_w21317_
	);
	LUT4 #(
		.INIT('habef)
	) name19417 (
		_w9166_,
		_w9169_,
		_w21316_,
		_w21317_,
		_w21318_
	);
	LUT3 #(
		.INIT('h2a)
	) name19418 (
		\m5_data_i[10]_pad ,
		_w9171_,
		_w9172_,
		_w21319_
	);
	LUT3 #(
		.INIT('h2a)
	) name19419 (
		\m1_data_i[10]_pad ,
		_w9171_,
		_w9172_,
		_w21320_
	);
	LUT4 #(
		.INIT('h57df)
	) name19420 (
		_w9166_,
		_w9169_,
		_w21319_,
		_w21320_,
		_w21321_
	);
	LUT3 #(
		.INIT('h80)
	) name19421 (
		\m0_data_i[10]_pad ,
		_w9171_,
		_w9172_,
		_w21322_
	);
	LUT3 #(
		.INIT('h2a)
	) name19422 (
		\m7_data_i[10]_pad ,
		_w9171_,
		_w9172_,
		_w21323_
	);
	LUT4 #(
		.INIT('h6e7f)
	) name19423 (
		_w9166_,
		_w9169_,
		_w21322_,
		_w21323_,
		_w21324_
	);
	LUT4 #(
		.INIT('h7fff)
	) name19424 (
		_w21315_,
		_w21318_,
		_w21321_,
		_w21324_,
		_w21325_
	);
	LUT3 #(
		.INIT('h2a)
	) name19425 (
		\m3_data_i[11]_pad ,
		_w9171_,
		_w9172_,
		_w21326_
	);
	LUT3 #(
		.INIT('h80)
	) name19426 (
		\m4_data_i[11]_pad ,
		_w9171_,
		_w9172_,
		_w21327_
	);
	LUT4 #(
		.INIT('h9dbf)
	) name19427 (
		_w9166_,
		_w9169_,
		_w21326_,
		_w21327_,
		_w21328_
	);
	LUT3 #(
		.INIT('h80)
	) name19428 (
		\m6_data_i[11]_pad ,
		_w9171_,
		_w9172_,
		_w21329_
	);
	LUT3 #(
		.INIT('h80)
	) name19429 (
		\m2_data_i[11]_pad ,
		_w9171_,
		_w9172_,
		_w21330_
	);
	LUT4 #(
		.INIT('habef)
	) name19430 (
		_w9166_,
		_w9169_,
		_w21329_,
		_w21330_,
		_w21331_
	);
	LUT3 #(
		.INIT('h2a)
	) name19431 (
		\m5_data_i[11]_pad ,
		_w9171_,
		_w9172_,
		_w21332_
	);
	LUT3 #(
		.INIT('h2a)
	) name19432 (
		\m1_data_i[11]_pad ,
		_w9171_,
		_w9172_,
		_w21333_
	);
	LUT4 #(
		.INIT('h57df)
	) name19433 (
		_w9166_,
		_w9169_,
		_w21332_,
		_w21333_,
		_w21334_
	);
	LUT3 #(
		.INIT('h80)
	) name19434 (
		\m0_data_i[11]_pad ,
		_w9171_,
		_w9172_,
		_w21335_
	);
	LUT3 #(
		.INIT('h2a)
	) name19435 (
		\m7_data_i[11]_pad ,
		_w9171_,
		_w9172_,
		_w21336_
	);
	LUT4 #(
		.INIT('h6e7f)
	) name19436 (
		_w9166_,
		_w9169_,
		_w21335_,
		_w21336_,
		_w21337_
	);
	LUT4 #(
		.INIT('h7fff)
	) name19437 (
		_w21328_,
		_w21331_,
		_w21334_,
		_w21337_,
		_w21338_
	);
	LUT3 #(
		.INIT('h2a)
	) name19438 (
		\m3_data_i[12]_pad ,
		_w9171_,
		_w9172_,
		_w21339_
	);
	LUT3 #(
		.INIT('h80)
	) name19439 (
		\m4_data_i[12]_pad ,
		_w9171_,
		_w9172_,
		_w21340_
	);
	LUT4 #(
		.INIT('h9dbf)
	) name19440 (
		_w9166_,
		_w9169_,
		_w21339_,
		_w21340_,
		_w21341_
	);
	LUT3 #(
		.INIT('h80)
	) name19441 (
		\m6_data_i[12]_pad ,
		_w9171_,
		_w9172_,
		_w21342_
	);
	LUT3 #(
		.INIT('h80)
	) name19442 (
		\m2_data_i[12]_pad ,
		_w9171_,
		_w9172_,
		_w21343_
	);
	LUT4 #(
		.INIT('habef)
	) name19443 (
		_w9166_,
		_w9169_,
		_w21342_,
		_w21343_,
		_w21344_
	);
	LUT3 #(
		.INIT('h2a)
	) name19444 (
		\m5_data_i[12]_pad ,
		_w9171_,
		_w9172_,
		_w21345_
	);
	LUT3 #(
		.INIT('h2a)
	) name19445 (
		\m1_data_i[12]_pad ,
		_w9171_,
		_w9172_,
		_w21346_
	);
	LUT4 #(
		.INIT('h57df)
	) name19446 (
		_w9166_,
		_w9169_,
		_w21345_,
		_w21346_,
		_w21347_
	);
	LUT3 #(
		.INIT('h80)
	) name19447 (
		\m0_data_i[12]_pad ,
		_w9171_,
		_w9172_,
		_w21348_
	);
	LUT3 #(
		.INIT('h2a)
	) name19448 (
		\m7_data_i[12]_pad ,
		_w9171_,
		_w9172_,
		_w21349_
	);
	LUT4 #(
		.INIT('h6e7f)
	) name19449 (
		_w9166_,
		_w9169_,
		_w21348_,
		_w21349_,
		_w21350_
	);
	LUT4 #(
		.INIT('h7fff)
	) name19450 (
		_w21341_,
		_w21344_,
		_w21347_,
		_w21350_,
		_w21351_
	);
	LUT3 #(
		.INIT('h2a)
	) name19451 (
		\m3_data_i[13]_pad ,
		_w9171_,
		_w9172_,
		_w21352_
	);
	LUT3 #(
		.INIT('h80)
	) name19452 (
		\m4_data_i[13]_pad ,
		_w9171_,
		_w9172_,
		_w21353_
	);
	LUT4 #(
		.INIT('h9dbf)
	) name19453 (
		_w9166_,
		_w9169_,
		_w21352_,
		_w21353_,
		_w21354_
	);
	LUT3 #(
		.INIT('h80)
	) name19454 (
		\m6_data_i[13]_pad ,
		_w9171_,
		_w9172_,
		_w21355_
	);
	LUT3 #(
		.INIT('h80)
	) name19455 (
		\m2_data_i[13]_pad ,
		_w9171_,
		_w9172_,
		_w21356_
	);
	LUT4 #(
		.INIT('habef)
	) name19456 (
		_w9166_,
		_w9169_,
		_w21355_,
		_w21356_,
		_w21357_
	);
	LUT3 #(
		.INIT('h2a)
	) name19457 (
		\m5_data_i[13]_pad ,
		_w9171_,
		_w9172_,
		_w21358_
	);
	LUT3 #(
		.INIT('h2a)
	) name19458 (
		\m1_data_i[13]_pad ,
		_w9171_,
		_w9172_,
		_w21359_
	);
	LUT4 #(
		.INIT('h57df)
	) name19459 (
		_w9166_,
		_w9169_,
		_w21358_,
		_w21359_,
		_w21360_
	);
	LUT3 #(
		.INIT('h80)
	) name19460 (
		\m0_data_i[13]_pad ,
		_w9171_,
		_w9172_,
		_w21361_
	);
	LUT3 #(
		.INIT('h2a)
	) name19461 (
		\m7_data_i[13]_pad ,
		_w9171_,
		_w9172_,
		_w21362_
	);
	LUT4 #(
		.INIT('h6e7f)
	) name19462 (
		_w9166_,
		_w9169_,
		_w21361_,
		_w21362_,
		_w21363_
	);
	LUT4 #(
		.INIT('h7fff)
	) name19463 (
		_w21354_,
		_w21357_,
		_w21360_,
		_w21363_,
		_w21364_
	);
	LUT3 #(
		.INIT('h2a)
	) name19464 (
		\m3_data_i[14]_pad ,
		_w9171_,
		_w9172_,
		_w21365_
	);
	LUT3 #(
		.INIT('h80)
	) name19465 (
		\m4_data_i[14]_pad ,
		_w9171_,
		_w9172_,
		_w21366_
	);
	LUT4 #(
		.INIT('h9dbf)
	) name19466 (
		_w9166_,
		_w9169_,
		_w21365_,
		_w21366_,
		_w21367_
	);
	LUT3 #(
		.INIT('h80)
	) name19467 (
		\m6_data_i[14]_pad ,
		_w9171_,
		_w9172_,
		_w21368_
	);
	LUT3 #(
		.INIT('h80)
	) name19468 (
		\m2_data_i[14]_pad ,
		_w9171_,
		_w9172_,
		_w21369_
	);
	LUT4 #(
		.INIT('habef)
	) name19469 (
		_w9166_,
		_w9169_,
		_w21368_,
		_w21369_,
		_w21370_
	);
	LUT3 #(
		.INIT('h2a)
	) name19470 (
		\m5_data_i[14]_pad ,
		_w9171_,
		_w9172_,
		_w21371_
	);
	LUT3 #(
		.INIT('h2a)
	) name19471 (
		\m1_data_i[14]_pad ,
		_w9171_,
		_w9172_,
		_w21372_
	);
	LUT4 #(
		.INIT('h57df)
	) name19472 (
		_w9166_,
		_w9169_,
		_w21371_,
		_w21372_,
		_w21373_
	);
	LUT3 #(
		.INIT('h80)
	) name19473 (
		\m0_data_i[14]_pad ,
		_w9171_,
		_w9172_,
		_w21374_
	);
	LUT3 #(
		.INIT('h2a)
	) name19474 (
		\m7_data_i[14]_pad ,
		_w9171_,
		_w9172_,
		_w21375_
	);
	LUT4 #(
		.INIT('h6e7f)
	) name19475 (
		_w9166_,
		_w9169_,
		_w21374_,
		_w21375_,
		_w21376_
	);
	LUT4 #(
		.INIT('h7fff)
	) name19476 (
		_w21367_,
		_w21370_,
		_w21373_,
		_w21376_,
		_w21377_
	);
	LUT3 #(
		.INIT('h2a)
	) name19477 (
		\m3_data_i[15]_pad ,
		_w9171_,
		_w9172_,
		_w21378_
	);
	LUT3 #(
		.INIT('h80)
	) name19478 (
		\m4_data_i[15]_pad ,
		_w9171_,
		_w9172_,
		_w21379_
	);
	LUT4 #(
		.INIT('h9dbf)
	) name19479 (
		_w9166_,
		_w9169_,
		_w21378_,
		_w21379_,
		_w21380_
	);
	LUT3 #(
		.INIT('h80)
	) name19480 (
		\m6_data_i[15]_pad ,
		_w9171_,
		_w9172_,
		_w21381_
	);
	LUT3 #(
		.INIT('h80)
	) name19481 (
		\m2_data_i[15]_pad ,
		_w9171_,
		_w9172_,
		_w21382_
	);
	LUT4 #(
		.INIT('habef)
	) name19482 (
		_w9166_,
		_w9169_,
		_w21381_,
		_w21382_,
		_w21383_
	);
	LUT3 #(
		.INIT('h2a)
	) name19483 (
		\m5_data_i[15]_pad ,
		_w9171_,
		_w9172_,
		_w21384_
	);
	LUT3 #(
		.INIT('h2a)
	) name19484 (
		\m1_data_i[15]_pad ,
		_w9171_,
		_w9172_,
		_w21385_
	);
	LUT4 #(
		.INIT('h57df)
	) name19485 (
		_w9166_,
		_w9169_,
		_w21384_,
		_w21385_,
		_w21386_
	);
	LUT3 #(
		.INIT('h80)
	) name19486 (
		\m0_data_i[15]_pad ,
		_w9171_,
		_w9172_,
		_w21387_
	);
	LUT3 #(
		.INIT('h2a)
	) name19487 (
		\m7_data_i[15]_pad ,
		_w9171_,
		_w9172_,
		_w21388_
	);
	LUT4 #(
		.INIT('h6e7f)
	) name19488 (
		_w9166_,
		_w9169_,
		_w21387_,
		_w21388_,
		_w21389_
	);
	LUT4 #(
		.INIT('h7fff)
	) name19489 (
		_w21380_,
		_w21383_,
		_w21386_,
		_w21389_,
		_w21390_
	);
	LUT3 #(
		.INIT('h2a)
	) name19490 (
		\m3_data_i[16]_pad ,
		_w9171_,
		_w9172_,
		_w21391_
	);
	LUT3 #(
		.INIT('h80)
	) name19491 (
		\m4_data_i[16]_pad ,
		_w9171_,
		_w9172_,
		_w21392_
	);
	LUT4 #(
		.INIT('h9dbf)
	) name19492 (
		_w9166_,
		_w9169_,
		_w21391_,
		_w21392_,
		_w21393_
	);
	LUT3 #(
		.INIT('h80)
	) name19493 (
		\m6_data_i[16]_pad ,
		_w9171_,
		_w9172_,
		_w21394_
	);
	LUT3 #(
		.INIT('h80)
	) name19494 (
		\m2_data_i[16]_pad ,
		_w9171_,
		_w9172_,
		_w21395_
	);
	LUT4 #(
		.INIT('habef)
	) name19495 (
		_w9166_,
		_w9169_,
		_w21394_,
		_w21395_,
		_w21396_
	);
	LUT3 #(
		.INIT('h2a)
	) name19496 (
		\m5_data_i[16]_pad ,
		_w9171_,
		_w9172_,
		_w21397_
	);
	LUT3 #(
		.INIT('h2a)
	) name19497 (
		\m1_data_i[16]_pad ,
		_w9171_,
		_w9172_,
		_w21398_
	);
	LUT4 #(
		.INIT('h57df)
	) name19498 (
		_w9166_,
		_w9169_,
		_w21397_,
		_w21398_,
		_w21399_
	);
	LUT3 #(
		.INIT('h80)
	) name19499 (
		\m0_data_i[16]_pad ,
		_w9171_,
		_w9172_,
		_w21400_
	);
	LUT3 #(
		.INIT('h2a)
	) name19500 (
		\m7_data_i[16]_pad ,
		_w9171_,
		_w9172_,
		_w21401_
	);
	LUT4 #(
		.INIT('h6e7f)
	) name19501 (
		_w9166_,
		_w9169_,
		_w21400_,
		_w21401_,
		_w21402_
	);
	LUT4 #(
		.INIT('h7fff)
	) name19502 (
		_w21393_,
		_w21396_,
		_w21399_,
		_w21402_,
		_w21403_
	);
	LUT3 #(
		.INIT('h2a)
	) name19503 (
		\m3_data_i[17]_pad ,
		_w9171_,
		_w9172_,
		_w21404_
	);
	LUT3 #(
		.INIT('h80)
	) name19504 (
		\m4_data_i[17]_pad ,
		_w9171_,
		_w9172_,
		_w21405_
	);
	LUT4 #(
		.INIT('h9dbf)
	) name19505 (
		_w9166_,
		_w9169_,
		_w21404_,
		_w21405_,
		_w21406_
	);
	LUT3 #(
		.INIT('h80)
	) name19506 (
		\m6_data_i[17]_pad ,
		_w9171_,
		_w9172_,
		_w21407_
	);
	LUT3 #(
		.INIT('h80)
	) name19507 (
		\m2_data_i[17]_pad ,
		_w9171_,
		_w9172_,
		_w21408_
	);
	LUT4 #(
		.INIT('habef)
	) name19508 (
		_w9166_,
		_w9169_,
		_w21407_,
		_w21408_,
		_w21409_
	);
	LUT3 #(
		.INIT('h2a)
	) name19509 (
		\m5_data_i[17]_pad ,
		_w9171_,
		_w9172_,
		_w21410_
	);
	LUT3 #(
		.INIT('h2a)
	) name19510 (
		\m1_data_i[17]_pad ,
		_w9171_,
		_w9172_,
		_w21411_
	);
	LUT4 #(
		.INIT('h57df)
	) name19511 (
		_w9166_,
		_w9169_,
		_w21410_,
		_w21411_,
		_w21412_
	);
	LUT3 #(
		.INIT('h80)
	) name19512 (
		\m0_data_i[17]_pad ,
		_w9171_,
		_w9172_,
		_w21413_
	);
	LUT3 #(
		.INIT('h2a)
	) name19513 (
		\m7_data_i[17]_pad ,
		_w9171_,
		_w9172_,
		_w21414_
	);
	LUT4 #(
		.INIT('h6e7f)
	) name19514 (
		_w9166_,
		_w9169_,
		_w21413_,
		_w21414_,
		_w21415_
	);
	LUT4 #(
		.INIT('h7fff)
	) name19515 (
		_w21406_,
		_w21409_,
		_w21412_,
		_w21415_,
		_w21416_
	);
	LUT3 #(
		.INIT('h2a)
	) name19516 (
		\m3_data_i[18]_pad ,
		_w9171_,
		_w9172_,
		_w21417_
	);
	LUT3 #(
		.INIT('h80)
	) name19517 (
		\m4_data_i[18]_pad ,
		_w9171_,
		_w9172_,
		_w21418_
	);
	LUT4 #(
		.INIT('h9dbf)
	) name19518 (
		_w9166_,
		_w9169_,
		_w21417_,
		_w21418_,
		_w21419_
	);
	LUT3 #(
		.INIT('h80)
	) name19519 (
		\m6_data_i[18]_pad ,
		_w9171_,
		_w9172_,
		_w21420_
	);
	LUT3 #(
		.INIT('h80)
	) name19520 (
		\m2_data_i[18]_pad ,
		_w9171_,
		_w9172_,
		_w21421_
	);
	LUT4 #(
		.INIT('habef)
	) name19521 (
		_w9166_,
		_w9169_,
		_w21420_,
		_w21421_,
		_w21422_
	);
	LUT3 #(
		.INIT('h2a)
	) name19522 (
		\m5_data_i[18]_pad ,
		_w9171_,
		_w9172_,
		_w21423_
	);
	LUT3 #(
		.INIT('h2a)
	) name19523 (
		\m1_data_i[18]_pad ,
		_w9171_,
		_w9172_,
		_w21424_
	);
	LUT4 #(
		.INIT('h57df)
	) name19524 (
		_w9166_,
		_w9169_,
		_w21423_,
		_w21424_,
		_w21425_
	);
	LUT3 #(
		.INIT('h80)
	) name19525 (
		\m0_data_i[18]_pad ,
		_w9171_,
		_w9172_,
		_w21426_
	);
	LUT3 #(
		.INIT('h2a)
	) name19526 (
		\m7_data_i[18]_pad ,
		_w9171_,
		_w9172_,
		_w21427_
	);
	LUT4 #(
		.INIT('h6e7f)
	) name19527 (
		_w9166_,
		_w9169_,
		_w21426_,
		_w21427_,
		_w21428_
	);
	LUT4 #(
		.INIT('h7fff)
	) name19528 (
		_w21419_,
		_w21422_,
		_w21425_,
		_w21428_,
		_w21429_
	);
	LUT3 #(
		.INIT('h2a)
	) name19529 (
		\m3_data_i[19]_pad ,
		_w9171_,
		_w9172_,
		_w21430_
	);
	LUT3 #(
		.INIT('h80)
	) name19530 (
		\m4_data_i[19]_pad ,
		_w9171_,
		_w9172_,
		_w21431_
	);
	LUT4 #(
		.INIT('h9dbf)
	) name19531 (
		_w9166_,
		_w9169_,
		_w21430_,
		_w21431_,
		_w21432_
	);
	LUT3 #(
		.INIT('h80)
	) name19532 (
		\m6_data_i[19]_pad ,
		_w9171_,
		_w9172_,
		_w21433_
	);
	LUT3 #(
		.INIT('h80)
	) name19533 (
		\m2_data_i[19]_pad ,
		_w9171_,
		_w9172_,
		_w21434_
	);
	LUT4 #(
		.INIT('habef)
	) name19534 (
		_w9166_,
		_w9169_,
		_w21433_,
		_w21434_,
		_w21435_
	);
	LUT3 #(
		.INIT('h2a)
	) name19535 (
		\m5_data_i[19]_pad ,
		_w9171_,
		_w9172_,
		_w21436_
	);
	LUT3 #(
		.INIT('h2a)
	) name19536 (
		\m1_data_i[19]_pad ,
		_w9171_,
		_w9172_,
		_w21437_
	);
	LUT4 #(
		.INIT('h57df)
	) name19537 (
		_w9166_,
		_w9169_,
		_w21436_,
		_w21437_,
		_w21438_
	);
	LUT3 #(
		.INIT('h80)
	) name19538 (
		\m0_data_i[19]_pad ,
		_w9171_,
		_w9172_,
		_w21439_
	);
	LUT3 #(
		.INIT('h2a)
	) name19539 (
		\m7_data_i[19]_pad ,
		_w9171_,
		_w9172_,
		_w21440_
	);
	LUT4 #(
		.INIT('h6e7f)
	) name19540 (
		_w9166_,
		_w9169_,
		_w21439_,
		_w21440_,
		_w21441_
	);
	LUT4 #(
		.INIT('h7fff)
	) name19541 (
		_w21432_,
		_w21435_,
		_w21438_,
		_w21441_,
		_w21442_
	);
	LUT3 #(
		.INIT('h2a)
	) name19542 (
		\m3_data_i[1]_pad ,
		_w9171_,
		_w9172_,
		_w21443_
	);
	LUT3 #(
		.INIT('h80)
	) name19543 (
		\m4_data_i[1]_pad ,
		_w9171_,
		_w9172_,
		_w21444_
	);
	LUT4 #(
		.INIT('h9dbf)
	) name19544 (
		_w9166_,
		_w9169_,
		_w21443_,
		_w21444_,
		_w21445_
	);
	LUT3 #(
		.INIT('h80)
	) name19545 (
		\m6_data_i[1]_pad ,
		_w9171_,
		_w9172_,
		_w21446_
	);
	LUT3 #(
		.INIT('h80)
	) name19546 (
		\m2_data_i[1]_pad ,
		_w9171_,
		_w9172_,
		_w21447_
	);
	LUT4 #(
		.INIT('habef)
	) name19547 (
		_w9166_,
		_w9169_,
		_w21446_,
		_w21447_,
		_w21448_
	);
	LUT3 #(
		.INIT('h2a)
	) name19548 (
		\m5_data_i[1]_pad ,
		_w9171_,
		_w9172_,
		_w21449_
	);
	LUT3 #(
		.INIT('h2a)
	) name19549 (
		\m1_data_i[1]_pad ,
		_w9171_,
		_w9172_,
		_w21450_
	);
	LUT4 #(
		.INIT('h57df)
	) name19550 (
		_w9166_,
		_w9169_,
		_w21449_,
		_w21450_,
		_w21451_
	);
	LUT3 #(
		.INIT('h80)
	) name19551 (
		\m0_data_i[1]_pad ,
		_w9171_,
		_w9172_,
		_w21452_
	);
	LUT3 #(
		.INIT('h2a)
	) name19552 (
		\m7_data_i[1]_pad ,
		_w9171_,
		_w9172_,
		_w21453_
	);
	LUT4 #(
		.INIT('h6e7f)
	) name19553 (
		_w9166_,
		_w9169_,
		_w21452_,
		_w21453_,
		_w21454_
	);
	LUT4 #(
		.INIT('h7fff)
	) name19554 (
		_w21445_,
		_w21448_,
		_w21451_,
		_w21454_,
		_w21455_
	);
	LUT3 #(
		.INIT('h2a)
	) name19555 (
		\m3_data_i[20]_pad ,
		_w9171_,
		_w9172_,
		_w21456_
	);
	LUT3 #(
		.INIT('h80)
	) name19556 (
		\m4_data_i[20]_pad ,
		_w9171_,
		_w9172_,
		_w21457_
	);
	LUT4 #(
		.INIT('h9dbf)
	) name19557 (
		_w9166_,
		_w9169_,
		_w21456_,
		_w21457_,
		_w21458_
	);
	LUT3 #(
		.INIT('h80)
	) name19558 (
		\m6_data_i[20]_pad ,
		_w9171_,
		_w9172_,
		_w21459_
	);
	LUT3 #(
		.INIT('h80)
	) name19559 (
		\m2_data_i[20]_pad ,
		_w9171_,
		_w9172_,
		_w21460_
	);
	LUT4 #(
		.INIT('habef)
	) name19560 (
		_w9166_,
		_w9169_,
		_w21459_,
		_w21460_,
		_w21461_
	);
	LUT3 #(
		.INIT('h2a)
	) name19561 (
		\m5_data_i[20]_pad ,
		_w9171_,
		_w9172_,
		_w21462_
	);
	LUT3 #(
		.INIT('h2a)
	) name19562 (
		\m1_data_i[20]_pad ,
		_w9171_,
		_w9172_,
		_w21463_
	);
	LUT4 #(
		.INIT('h57df)
	) name19563 (
		_w9166_,
		_w9169_,
		_w21462_,
		_w21463_,
		_w21464_
	);
	LUT3 #(
		.INIT('h80)
	) name19564 (
		\m0_data_i[20]_pad ,
		_w9171_,
		_w9172_,
		_w21465_
	);
	LUT3 #(
		.INIT('h2a)
	) name19565 (
		\m7_data_i[20]_pad ,
		_w9171_,
		_w9172_,
		_w21466_
	);
	LUT4 #(
		.INIT('h6e7f)
	) name19566 (
		_w9166_,
		_w9169_,
		_w21465_,
		_w21466_,
		_w21467_
	);
	LUT4 #(
		.INIT('h7fff)
	) name19567 (
		_w21458_,
		_w21461_,
		_w21464_,
		_w21467_,
		_w21468_
	);
	LUT3 #(
		.INIT('h2a)
	) name19568 (
		\m3_data_i[21]_pad ,
		_w9171_,
		_w9172_,
		_w21469_
	);
	LUT3 #(
		.INIT('h80)
	) name19569 (
		\m4_data_i[21]_pad ,
		_w9171_,
		_w9172_,
		_w21470_
	);
	LUT4 #(
		.INIT('h9dbf)
	) name19570 (
		_w9166_,
		_w9169_,
		_w21469_,
		_w21470_,
		_w21471_
	);
	LUT3 #(
		.INIT('h80)
	) name19571 (
		\m6_data_i[21]_pad ,
		_w9171_,
		_w9172_,
		_w21472_
	);
	LUT3 #(
		.INIT('h80)
	) name19572 (
		\m2_data_i[21]_pad ,
		_w9171_,
		_w9172_,
		_w21473_
	);
	LUT4 #(
		.INIT('habef)
	) name19573 (
		_w9166_,
		_w9169_,
		_w21472_,
		_w21473_,
		_w21474_
	);
	LUT3 #(
		.INIT('h2a)
	) name19574 (
		\m5_data_i[21]_pad ,
		_w9171_,
		_w9172_,
		_w21475_
	);
	LUT3 #(
		.INIT('h2a)
	) name19575 (
		\m1_data_i[21]_pad ,
		_w9171_,
		_w9172_,
		_w21476_
	);
	LUT4 #(
		.INIT('h57df)
	) name19576 (
		_w9166_,
		_w9169_,
		_w21475_,
		_w21476_,
		_w21477_
	);
	LUT3 #(
		.INIT('h80)
	) name19577 (
		\m0_data_i[21]_pad ,
		_w9171_,
		_w9172_,
		_w21478_
	);
	LUT3 #(
		.INIT('h2a)
	) name19578 (
		\m7_data_i[21]_pad ,
		_w9171_,
		_w9172_,
		_w21479_
	);
	LUT4 #(
		.INIT('h6e7f)
	) name19579 (
		_w9166_,
		_w9169_,
		_w21478_,
		_w21479_,
		_w21480_
	);
	LUT4 #(
		.INIT('h7fff)
	) name19580 (
		_w21471_,
		_w21474_,
		_w21477_,
		_w21480_,
		_w21481_
	);
	LUT3 #(
		.INIT('h2a)
	) name19581 (
		\m3_data_i[22]_pad ,
		_w9171_,
		_w9172_,
		_w21482_
	);
	LUT3 #(
		.INIT('h80)
	) name19582 (
		\m4_data_i[22]_pad ,
		_w9171_,
		_w9172_,
		_w21483_
	);
	LUT4 #(
		.INIT('h9dbf)
	) name19583 (
		_w9166_,
		_w9169_,
		_w21482_,
		_w21483_,
		_w21484_
	);
	LUT3 #(
		.INIT('h80)
	) name19584 (
		\m6_data_i[22]_pad ,
		_w9171_,
		_w9172_,
		_w21485_
	);
	LUT3 #(
		.INIT('h80)
	) name19585 (
		\m2_data_i[22]_pad ,
		_w9171_,
		_w9172_,
		_w21486_
	);
	LUT4 #(
		.INIT('habef)
	) name19586 (
		_w9166_,
		_w9169_,
		_w21485_,
		_w21486_,
		_w21487_
	);
	LUT3 #(
		.INIT('h2a)
	) name19587 (
		\m5_data_i[22]_pad ,
		_w9171_,
		_w9172_,
		_w21488_
	);
	LUT3 #(
		.INIT('h2a)
	) name19588 (
		\m1_data_i[22]_pad ,
		_w9171_,
		_w9172_,
		_w21489_
	);
	LUT4 #(
		.INIT('h57df)
	) name19589 (
		_w9166_,
		_w9169_,
		_w21488_,
		_w21489_,
		_w21490_
	);
	LUT3 #(
		.INIT('h80)
	) name19590 (
		\m0_data_i[22]_pad ,
		_w9171_,
		_w9172_,
		_w21491_
	);
	LUT3 #(
		.INIT('h2a)
	) name19591 (
		\m7_data_i[22]_pad ,
		_w9171_,
		_w9172_,
		_w21492_
	);
	LUT4 #(
		.INIT('h6e7f)
	) name19592 (
		_w9166_,
		_w9169_,
		_w21491_,
		_w21492_,
		_w21493_
	);
	LUT4 #(
		.INIT('h7fff)
	) name19593 (
		_w21484_,
		_w21487_,
		_w21490_,
		_w21493_,
		_w21494_
	);
	LUT3 #(
		.INIT('h2a)
	) name19594 (
		\m3_data_i[23]_pad ,
		_w9171_,
		_w9172_,
		_w21495_
	);
	LUT3 #(
		.INIT('h80)
	) name19595 (
		\m4_data_i[23]_pad ,
		_w9171_,
		_w9172_,
		_w21496_
	);
	LUT4 #(
		.INIT('h9dbf)
	) name19596 (
		_w9166_,
		_w9169_,
		_w21495_,
		_w21496_,
		_w21497_
	);
	LUT3 #(
		.INIT('h80)
	) name19597 (
		\m6_data_i[23]_pad ,
		_w9171_,
		_w9172_,
		_w21498_
	);
	LUT3 #(
		.INIT('h80)
	) name19598 (
		\m2_data_i[23]_pad ,
		_w9171_,
		_w9172_,
		_w21499_
	);
	LUT4 #(
		.INIT('habef)
	) name19599 (
		_w9166_,
		_w9169_,
		_w21498_,
		_w21499_,
		_w21500_
	);
	LUT3 #(
		.INIT('h2a)
	) name19600 (
		\m5_data_i[23]_pad ,
		_w9171_,
		_w9172_,
		_w21501_
	);
	LUT3 #(
		.INIT('h2a)
	) name19601 (
		\m1_data_i[23]_pad ,
		_w9171_,
		_w9172_,
		_w21502_
	);
	LUT4 #(
		.INIT('h57df)
	) name19602 (
		_w9166_,
		_w9169_,
		_w21501_,
		_w21502_,
		_w21503_
	);
	LUT3 #(
		.INIT('h80)
	) name19603 (
		\m0_data_i[23]_pad ,
		_w9171_,
		_w9172_,
		_w21504_
	);
	LUT3 #(
		.INIT('h2a)
	) name19604 (
		\m7_data_i[23]_pad ,
		_w9171_,
		_w9172_,
		_w21505_
	);
	LUT4 #(
		.INIT('h6e7f)
	) name19605 (
		_w9166_,
		_w9169_,
		_w21504_,
		_w21505_,
		_w21506_
	);
	LUT4 #(
		.INIT('h7fff)
	) name19606 (
		_w21497_,
		_w21500_,
		_w21503_,
		_w21506_,
		_w21507_
	);
	LUT3 #(
		.INIT('h2a)
	) name19607 (
		\m3_data_i[24]_pad ,
		_w9171_,
		_w9172_,
		_w21508_
	);
	LUT3 #(
		.INIT('h80)
	) name19608 (
		\m4_data_i[24]_pad ,
		_w9171_,
		_w9172_,
		_w21509_
	);
	LUT4 #(
		.INIT('h9dbf)
	) name19609 (
		_w9166_,
		_w9169_,
		_w21508_,
		_w21509_,
		_w21510_
	);
	LUT3 #(
		.INIT('h80)
	) name19610 (
		\m6_data_i[24]_pad ,
		_w9171_,
		_w9172_,
		_w21511_
	);
	LUT3 #(
		.INIT('h80)
	) name19611 (
		\m2_data_i[24]_pad ,
		_w9171_,
		_w9172_,
		_w21512_
	);
	LUT4 #(
		.INIT('habef)
	) name19612 (
		_w9166_,
		_w9169_,
		_w21511_,
		_w21512_,
		_w21513_
	);
	LUT3 #(
		.INIT('h2a)
	) name19613 (
		\m5_data_i[24]_pad ,
		_w9171_,
		_w9172_,
		_w21514_
	);
	LUT3 #(
		.INIT('h2a)
	) name19614 (
		\m1_data_i[24]_pad ,
		_w9171_,
		_w9172_,
		_w21515_
	);
	LUT4 #(
		.INIT('h57df)
	) name19615 (
		_w9166_,
		_w9169_,
		_w21514_,
		_w21515_,
		_w21516_
	);
	LUT3 #(
		.INIT('h80)
	) name19616 (
		\m0_data_i[24]_pad ,
		_w9171_,
		_w9172_,
		_w21517_
	);
	LUT3 #(
		.INIT('h2a)
	) name19617 (
		\m7_data_i[24]_pad ,
		_w9171_,
		_w9172_,
		_w21518_
	);
	LUT4 #(
		.INIT('h6e7f)
	) name19618 (
		_w9166_,
		_w9169_,
		_w21517_,
		_w21518_,
		_w21519_
	);
	LUT4 #(
		.INIT('h7fff)
	) name19619 (
		_w21510_,
		_w21513_,
		_w21516_,
		_w21519_,
		_w21520_
	);
	LUT3 #(
		.INIT('h2a)
	) name19620 (
		\m3_data_i[25]_pad ,
		_w9171_,
		_w9172_,
		_w21521_
	);
	LUT3 #(
		.INIT('h80)
	) name19621 (
		\m4_data_i[25]_pad ,
		_w9171_,
		_w9172_,
		_w21522_
	);
	LUT4 #(
		.INIT('h9dbf)
	) name19622 (
		_w9166_,
		_w9169_,
		_w21521_,
		_w21522_,
		_w21523_
	);
	LUT3 #(
		.INIT('h80)
	) name19623 (
		\m6_data_i[25]_pad ,
		_w9171_,
		_w9172_,
		_w21524_
	);
	LUT3 #(
		.INIT('h80)
	) name19624 (
		\m2_data_i[25]_pad ,
		_w9171_,
		_w9172_,
		_w21525_
	);
	LUT4 #(
		.INIT('habef)
	) name19625 (
		_w9166_,
		_w9169_,
		_w21524_,
		_w21525_,
		_w21526_
	);
	LUT3 #(
		.INIT('h2a)
	) name19626 (
		\m5_data_i[25]_pad ,
		_w9171_,
		_w9172_,
		_w21527_
	);
	LUT3 #(
		.INIT('h2a)
	) name19627 (
		\m1_data_i[25]_pad ,
		_w9171_,
		_w9172_,
		_w21528_
	);
	LUT4 #(
		.INIT('h57df)
	) name19628 (
		_w9166_,
		_w9169_,
		_w21527_,
		_w21528_,
		_w21529_
	);
	LUT3 #(
		.INIT('h80)
	) name19629 (
		\m0_data_i[25]_pad ,
		_w9171_,
		_w9172_,
		_w21530_
	);
	LUT3 #(
		.INIT('h2a)
	) name19630 (
		\m7_data_i[25]_pad ,
		_w9171_,
		_w9172_,
		_w21531_
	);
	LUT4 #(
		.INIT('h6e7f)
	) name19631 (
		_w9166_,
		_w9169_,
		_w21530_,
		_w21531_,
		_w21532_
	);
	LUT4 #(
		.INIT('h7fff)
	) name19632 (
		_w21523_,
		_w21526_,
		_w21529_,
		_w21532_,
		_w21533_
	);
	LUT3 #(
		.INIT('h80)
	) name19633 (
		\m0_data_i[26]_pad ,
		_w9171_,
		_w9172_,
		_w21534_
	);
	LUT3 #(
		.INIT('h2a)
	) name19634 (
		\m7_data_i[26]_pad ,
		_w9171_,
		_w9172_,
		_w21535_
	);
	LUT4 #(
		.INIT('h6e7f)
	) name19635 (
		_w9166_,
		_w9169_,
		_w21534_,
		_w21535_,
		_w21536_
	);
	LUT3 #(
		.INIT('h2a)
	) name19636 (
		\m1_data_i[26]_pad ,
		_w9171_,
		_w9172_,
		_w21537_
	);
	LUT3 #(
		.INIT('h80)
	) name19637 (
		\m4_data_i[26]_pad ,
		_w9171_,
		_w9172_,
		_w21538_
	);
	LUT4 #(
		.INIT('h5d7f)
	) name19638 (
		_w9166_,
		_w9169_,
		_w21537_,
		_w21538_,
		_w21539_
	);
	LUT3 #(
		.INIT('h80)
	) name19639 (
		\m2_data_i[26]_pad ,
		_w9171_,
		_w9172_,
		_w21540_
	);
	LUT3 #(
		.INIT('h2a)
	) name19640 (
		\m3_data_i[26]_pad ,
		_w9171_,
		_w9172_,
		_w21541_
	);
	LUT3 #(
		.INIT('h57)
	) name19641 (
		_w9190_,
		_w21540_,
		_w21541_,
		_w21542_
	);
	LUT3 #(
		.INIT('h80)
	) name19642 (
		\m6_data_i[26]_pad ,
		_w9171_,
		_w9172_,
		_w21543_
	);
	LUT3 #(
		.INIT('h2a)
	) name19643 (
		\m5_data_i[26]_pad ,
		_w9171_,
		_w9172_,
		_w21544_
	);
	LUT4 #(
		.INIT('hcdef)
	) name19644 (
		_w9166_,
		_w9169_,
		_w21543_,
		_w21544_,
		_w21545_
	);
	LUT4 #(
		.INIT('h7fff)
	) name19645 (
		_w21536_,
		_w21539_,
		_w21542_,
		_w21545_,
		_w21546_
	);
	LUT3 #(
		.INIT('h2a)
	) name19646 (
		\m1_data_i[27]_pad ,
		_w9171_,
		_w9172_,
		_w21547_
	);
	LUT3 #(
		.INIT('h80)
	) name19647 (
		\m2_data_i[27]_pad ,
		_w9171_,
		_w9172_,
		_w21548_
	);
	LUT4 #(
		.INIT('h3b7f)
	) name19648 (
		_w9166_,
		_w9169_,
		_w21547_,
		_w21548_,
		_w21549_
	);
	LUT3 #(
		.INIT('h80)
	) name19649 (
		\m6_data_i[27]_pad ,
		_w9171_,
		_w9172_,
		_w21550_
	);
	LUT3 #(
		.INIT('h2a)
	) name19650 (
		\m7_data_i[27]_pad ,
		_w9171_,
		_w9172_,
		_w21551_
	);
	LUT3 #(
		.INIT('h57)
	) name19651 (
		_w9184_,
		_w21550_,
		_w21551_,
		_w21552_
	);
	LUT3 #(
		.INIT('h2a)
	) name19652 (
		\m5_data_i[27]_pad ,
		_w9171_,
		_w9172_,
		_w21553_
	);
	LUT3 #(
		.INIT('h80)
	) name19653 (
		\m0_data_i[27]_pad ,
		_w9171_,
		_w9172_,
		_w21554_
	);
	LUT4 #(
		.INIT('h57df)
	) name19654 (
		_w9166_,
		_w9169_,
		_w21553_,
		_w21554_,
		_w21555_
	);
	LUT3 #(
		.INIT('h2a)
	) name19655 (
		\m3_data_i[27]_pad ,
		_w9171_,
		_w9172_,
		_w21556_
	);
	LUT3 #(
		.INIT('h80)
	) name19656 (
		\m4_data_i[27]_pad ,
		_w9171_,
		_w9172_,
		_w21557_
	);
	LUT4 #(
		.INIT('h9dbf)
	) name19657 (
		_w9166_,
		_w9169_,
		_w21556_,
		_w21557_,
		_w21558_
	);
	LUT4 #(
		.INIT('h7fff)
	) name19658 (
		_w21549_,
		_w21552_,
		_w21555_,
		_w21558_,
		_w21559_
	);
	LUT3 #(
		.INIT('h2a)
	) name19659 (
		\m1_data_i[28]_pad ,
		_w9171_,
		_w9172_,
		_w21560_
	);
	LUT3 #(
		.INIT('h80)
	) name19660 (
		\m2_data_i[28]_pad ,
		_w9171_,
		_w9172_,
		_w21561_
	);
	LUT4 #(
		.INIT('h3b7f)
	) name19661 (
		_w9166_,
		_w9169_,
		_w21560_,
		_w21561_,
		_w21562_
	);
	LUT3 #(
		.INIT('h80)
	) name19662 (
		\m0_data_i[28]_pad ,
		_w9171_,
		_w9172_,
		_w21563_
	);
	LUT3 #(
		.INIT('h80)
	) name19663 (
		\m4_data_i[28]_pad ,
		_w9171_,
		_w9172_,
		_w21564_
	);
	LUT4 #(
		.INIT('h5d7f)
	) name19664 (
		_w9166_,
		_w9169_,
		_w21563_,
		_w21564_,
		_w21565_
	);
	LUT3 #(
		.INIT('h2a)
	) name19665 (
		\m7_data_i[28]_pad ,
		_w9171_,
		_w9172_,
		_w21566_
	);
	LUT3 #(
		.INIT('h2a)
	) name19666 (
		\m3_data_i[28]_pad ,
		_w9171_,
		_w9172_,
		_w21567_
	);
	LUT4 #(
		.INIT('habef)
	) name19667 (
		_w9166_,
		_w9169_,
		_w21566_,
		_w21567_,
		_w21568_
	);
	LUT3 #(
		.INIT('h80)
	) name19668 (
		\m6_data_i[28]_pad ,
		_w9171_,
		_w9172_,
		_w21569_
	);
	LUT3 #(
		.INIT('h2a)
	) name19669 (
		\m5_data_i[28]_pad ,
		_w9171_,
		_w9172_,
		_w21570_
	);
	LUT4 #(
		.INIT('hcdef)
	) name19670 (
		_w9166_,
		_w9169_,
		_w21569_,
		_w21570_,
		_w21571_
	);
	LUT4 #(
		.INIT('h7fff)
	) name19671 (
		_w21562_,
		_w21565_,
		_w21568_,
		_w21571_,
		_w21572_
	);
	LUT3 #(
		.INIT('h2a)
	) name19672 (
		\m3_data_i[29]_pad ,
		_w9171_,
		_w9172_,
		_w21573_
	);
	LUT3 #(
		.INIT('h80)
	) name19673 (
		\m4_data_i[29]_pad ,
		_w9171_,
		_w9172_,
		_w21574_
	);
	LUT4 #(
		.INIT('h9dbf)
	) name19674 (
		_w9166_,
		_w9169_,
		_w21573_,
		_w21574_,
		_w21575_
	);
	LUT3 #(
		.INIT('h80)
	) name19675 (
		\m6_data_i[29]_pad ,
		_w9171_,
		_w9172_,
		_w21576_
	);
	LUT3 #(
		.INIT('h2a)
	) name19676 (
		\m7_data_i[29]_pad ,
		_w9171_,
		_w9172_,
		_w21577_
	);
	LUT3 #(
		.INIT('h57)
	) name19677 (
		_w9184_,
		_w21576_,
		_w21577_,
		_w21578_
	);
	LUT3 #(
		.INIT('h2a)
	) name19678 (
		\m5_data_i[29]_pad ,
		_w9171_,
		_w9172_,
		_w21579_
	);
	LUT3 #(
		.INIT('h80)
	) name19679 (
		\m0_data_i[29]_pad ,
		_w9171_,
		_w9172_,
		_w21580_
	);
	LUT4 #(
		.INIT('h57df)
	) name19680 (
		_w9166_,
		_w9169_,
		_w21579_,
		_w21580_,
		_w21581_
	);
	LUT3 #(
		.INIT('h2a)
	) name19681 (
		\m1_data_i[29]_pad ,
		_w9171_,
		_w9172_,
		_w21582_
	);
	LUT3 #(
		.INIT('h80)
	) name19682 (
		\m2_data_i[29]_pad ,
		_w9171_,
		_w9172_,
		_w21583_
	);
	LUT4 #(
		.INIT('h3b7f)
	) name19683 (
		_w9166_,
		_w9169_,
		_w21582_,
		_w21583_,
		_w21584_
	);
	LUT4 #(
		.INIT('h7fff)
	) name19684 (
		_w21575_,
		_w21578_,
		_w21581_,
		_w21584_,
		_w21585_
	);
	LUT3 #(
		.INIT('h2a)
	) name19685 (
		\m3_data_i[2]_pad ,
		_w9171_,
		_w9172_,
		_w21586_
	);
	LUT3 #(
		.INIT('h80)
	) name19686 (
		\m4_data_i[2]_pad ,
		_w9171_,
		_w9172_,
		_w21587_
	);
	LUT4 #(
		.INIT('h9dbf)
	) name19687 (
		_w9166_,
		_w9169_,
		_w21586_,
		_w21587_,
		_w21588_
	);
	LUT3 #(
		.INIT('h80)
	) name19688 (
		\m6_data_i[2]_pad ,
		_w9171_,
		_w9172_,
		_w21589_
	);
	LUT3 #(
		.INIT('h80)
	) name19689 (
		\m2_data_i[2]_pad ,
		_w9171_,
		_w9172_,
		_w21590_
	);
	LUT4 #(
		.INIT('habef)
	) name19690 (
		_w9166_,
		_w9169_,
		_w21589_,
		_w21590_,
		_w21591_
	);
	LUT3 #(
		.INIT('h2a)
	) name19691 (
		\m5_data_i[2]_pad ,
		_w9171_,
		_w9172_,
		_w21592_
	);
	LUT3 #(
		.INIT('h2a)
	) name19692 (
		\m1_data_i[2]_pad ,
		_w9171_,
		_w9172_,
		_w21593_
	);
	LUT4 #(
		.INIT('h57df)
	) name19693 (
		_w9166_,
		_w9169_,
		_w21592_,
		_w21593_,
		_w21594_
	);
	LUT3 #(
		.INIT('h80)
	) name19694 (
		\m0_data_i[2]_pad ,
		_w9171_,
		_w9172_,
		_w21595_
	);
	LUT3 #(
		.INIT('h2a)
	) name19695 (
		\m7_data_i[2]_pad ,
		_w9171_,
		_w9172_,
		_w21596_
	);
	LUT4 #(
		.INIT('h6e7f)
	) name19696 (
		_w9166_,
		_w9169_,
		_w21595_,
		_w21596_,
		_w21597_
	);
	LUT4 #(
		.INIT('h7fff)
	) name19697 (
		_w21588_,
		_w21591_,
		_w21594_,
		_w21597_,
		_w21598_
	);
	LUT3 #(
		.INIT('h2a)
	) name19698 (
		\m1_data_i[30]_pad ,
		_w9171_,
		_w9172_,
		_w21599_
	);
	LUT3 #(
		.INIT('h80)
	) name19699 (
		\m2_data_i[30]_pad ,
		_w9171_,
		_w9172_,
		_w21600_
	);
	LUT4 #(
		.INIT('h3b7f)
	) name19700 (
		_w9166_,
		_w9169_,
		_w21599_,
		_w21600_,
		_w21601_
	);
	LUT3 #(
		.INIT('h2a)
	) name19701 (
		\m3_data_i[30]_pad ,
		_w9171_,
		_w9172_,
		_w21602_
	);
	LUT3 #(
		.INIT('h2a)
	) name19702 (
		\m7_data_i[30]_pad ,
		_w9171_,
		_w9172_,
		_w21603_
	);
	LUT4 #(
		.INIT('haebf)
	) name19703 (
		_w9166_,
		_w9169_,
		_w21602_,
		_w21603_,
		_w21604_
	);
	LUT3 #(
		.INIT('h80)
	) name19704 (
		\m4_data_i[30]_pad ,
		_w9171_,
		_w9172_,
		_w21605_
	);
	LUT3 #(
		.INIT('h80)
	) name19705 (
		\m0_data_i[30]_pad ,
		_w9171_,
		_w9172_,
		_w21606_
	);
	LUT4 #(
		.INIT('h57df)
	) name19706 (
		_w9166_,
		_w9169_,
		_w21605_,
		_w21606_,
		_w21607_
	);
	LUT3 #(
		.INIT('h80)
	) name19707 (
		\m6_data_i[30]_pad ,
		_w9171_,
		_w9172_,
		_w21608_
	);
	LUT3 #(
		.INIT('h2a)
	) name19708 (
		\m5_data_i[30]_pad ,
		_w9171_,
		_w9172_,
		_w21609_
	);
	LUT4 #(
		.INIT('hcdef)
	) name19709 (
		_w9166_,
		_w9169_,
		_w21608_,
		_w21609_,
		_w21610_
	);
	LUT4 #(
		.INIT('h7fff)
	) name19710 (
		_w21601_,
		_w21604_,
		_w21607_,
		_w21610_,
		_w21611_
	);
	LUT3 #(
		.INIT('h2a)
	) name19711 (
		\m1_data_i[31]_pad ,
		_w9171_,
		_w9172_,
		_w21612_
	);
	LUT3 #(
		.INIT('h80)
	) name19712 (
		\m2_data_i[31]_pad ,
		_w9171_,
		_w9172_,
		_w21613_
	);
	LUT4 #(
		.INIT('h3b7f)
	) name19713 (
		_w9166_,
		_w9169_,
		_w21612_,
		_w21613_,
		_w21614_
	);
	LUT3 #(
		.INIT('h80)
	) name19714 (
		\m6_data_i[31]_pad ,
		_w9171_,
		_w9172_,
		_w21615_
	);
	LUT3 #(
		.INIT('h80)
	) name19715 (
		\m4_data_i[31]_pad ,
		_w9171_,
		_w9172_,
		_w21616_
	);
	LUT4 #(
		.INIT('hcdef)
	) name19716 (
		_w9166_,
		_w9169_,
		_w21615_,
		_w21616_,
		_w21617_
	);
	LUT3 #(
		.INIT('h2a)
	) name19717 (
		\m5_data_i[31]_pad ,
		_w9171_,
		_w9172_,
		_w21618_
	);
	LUT3 #(
		.INIT('h2a)
	) name19718 (
		\m3_data_i[31]_pad ,
		_w9171_,
		_w9172_,
		_w21619_
	);
	LUT4 #(
		.INIT('h9bdf)
	) name19719 (
		_w9166_,
		_w9169_,
		_w21618_,
		_w21619_,
		_w21620_
	);
	LUT3 #(
		.INIT('h80)
	) name19720 (
		\m0_data_i[31]_pad ,
		_w9171_,
		_w9172_,
		_w21621_
	);
	LUT3 #(
		.INIT('h2a)
	) name19721 (
		\m7_data_i[31]_pad ,
		_w9171_,
		_w9172_,
		_w21622_
	);
	LUT4 #(
		.INIT('h6e7f)
	) name19722 (
		_w9166_,
		_w9169_,
		_w21621_,
		_w21622_,
		_w21623_
	);
	LUT4 #(
		.INIT('h7fff)
	) name19723 (
		_w21614_,
		_w21617_,
		_w21620_,
		_w21623_,
		_w21624_
	);
	LUT3 #(
		.INIT('h2a)
	) name19724 (
		\m3_data_i[3]_pad ,
		_w9171_,
		_w9172_,
		_w21625_
	);
	LUT3 #(
		.INIT('h80)
	) name19725 (
		\m4_data_i[3]_pad ,
		_w9171_,
		_w9172_,
		_w21626_
	);
	LUT4 #(
		.INIT('h9dbf)
	) name19726 (
		_w9166_,
		_w9169_,
		_w21625_,
		_w21626_,
		_w21627_
	);
	LUT3 #(
		.INIT('h80)
	) name19727 (
		\m6_data_i[3]_pad ,
		_w9171_,
		_w9172_,
		_w21628_
	);
	LUT3 #(
		.INIT('h80)
	) name19728 (
		\m2_data_i[3]_pad ,
		_w9171_,
		_w9172_,
		_w21629_
	);
	LUT4 #(
		.INIT('habef)
	) name19729 (
		_w9166_,
		_w9169_,
		_w21628_,
		_w21629_,
		_w21630_
	);
	LUT3 #(
		.INIT('h2a)
	) name19730 (
		\m5_data_i[3]_pad ,
		_w9171_,
		_w9172_,
		_w21631_
	);
	LUT3 #(
		.INIT('h2a)
	) name19731 (
		\m1_data_i[3]_pad ,
		_w9171_,
		_w9172_,
		_w21632_
	);
	LUT4 #(
		.INIT('h57df)
	) name19732 (
		_w9166_,
		_w9169_,
		_w21631_,
		_w21632_,
		_w21633_
	);
	LUT3 #(
		.INIT('h80)
	) name19733 (
		\m0_data_i[3]_pad ,
		_w9171_,
		_w9172_,
		_w21634_
	);
	LUT3 #(
		.INIT('h2a)
	) name19734 (
		\m7_data_i[3]_pad ,
		_w9171_,
		_w9172_,
		_w21635_
	);
	LUT4 #(
		.INIT('h6e7f)
	) name19735 (
		_w9166_,
		_w9169_,
		_w21634_,
		_w21635_,
		_w21636_
	);
	LUT4 #(
		.INIT('h7fff)
	) name19736 (
		_w21627_,
		_w21630_,
		_w21633_,
		_w21636_,
		_w21637_
	);
	LUT3 #(
		.INIT('h2a)
	) name19737 (
		\m3_data_i[4]_pad ,
		_w9171_,
		_w9172_,
		_w21638_
	);
	LUT3 #(
		.INIT('h80)
	) name19738 (
		\m4_data_i[4]_pad ,
		_w9171_,
		_w9172_,
		_w21639_
	);
	LUT4 #(
		.INIT('h9dbf)
	) name19739 (
		_w9166_,
		_w9169_,
		_w21638_,
		_w21639_,
		_w21640_
	);
	LUT3 #(
		.INIT('h80)
	) name19740 (
		\m6_data_i[4]_pad ,
		_w9171_,
		_w9172_,
		_w21641_
	);
	LUT3 #(
		.INIT('h80)
	) name19741 (
		\m2_data_i[4]_pad ,
		_w9171_,
		_w9172_,
		_w21642_
	);
	LUT4 #(
		.INIT('habef)
	) name19742 (
		_w9166_,
		_w9169_,
		_w21641_,
		_w21642_,
		_w21643_
	);
	LUT3 #(
		.INIT('h2a)
	) name19743 (
		\m5_data_i[4]_pad ,
		_w9171_,
		_w9172_,
		_w21644_
	);
	LUT3 #(
		.INIT('h2a)
	) name19744 (
		\m1_data_i[4]_pad ,
		_w9171_,
		_w9172_,
		_w21645_
	);
	LUT4 #(
		.INIT('h57df)
	) name19745 (
		_w9166_,
		_w9169_,
		_w21644_,
		_w21645_,
		_w21646_
	);
	LUT3 #(
		.INIT('h80)
	) name19746 (
		\m0_data_i[4]_pad ,
		_w9171_,
		_w9172_,
		_w21647_
	);
	LUT3 #(
		.INIT('h2a)
	) name19747 (
		\m7_data_i[4]_pad ,
		_w9171_,
		_w9172_,
		_w21648_
	);
	LUT4 #(
		.INIT('h6e7f)
	) name19748 (
		_w9166_,
		_w9169_,
		_w21647_,
		_w21648_,
		_w21649_
	);
	LUT4 #(
		.INIT('h7fff)
	) name19749 (
		_w21640_,
		_w21643_,
		_w21646_,
		_w21649_,
		_w21650_
	);
	LUT3 #(
		.INIT('h2a)
	) name19750 (
		\m3_data_i[5]_pad ,
		_w9171_,
		_w9172_,
		_w21651_
	);
	LUT3 #(
		.INIT('h80)
	) name19751 (
		\m4_data_i[5]_pad ,
		_w9171_,
		_w9172_,
		_w21652_
	);
	LUT4 #(
		.INIT('h9dbf)
	) name19752 (
		_w9166_,
		_w9169_,
		_w21651_,
		_w21652_,
		_w21653_
	);
	LUT3 #(
		.INIT('h80)
	) name19753 (
		\m6_data_i[5]_pad ,
		_w9171_,
		_w9172_,
		_w21654_
	);
	LUT3 #(
		.INIT('h80)
	) name19754 (
		\m2_data_i[5]_pad ,
		_w9171_,
		_w9172_,
		_w21655_
	);
	LUT4 #(
		.INIT('habef)
	) name19755 (
		_w9166_,
		_w9169_,
		_w21654_,
		_w21655_,
		_w21656_
	);
	LUT3 #(
		.INIT('h2a)
	) name19756 (
		\m5_data_i[5]_pad ,
		_w9171_,
		_w9172_,
		_w21657_
	);
	LUT3 #(
		.INIT('h2a)
	) name19757 (
		\m1_data_i[5]_pad ,
		_w9171_,
		_w9172_,
		_w21658_
	);
	LUT4 #(
		.INIT('h57df)
	) name19758 (
		_w9166_,
		_w9169_,
		_w21657_,
		_w21658_,
		_w21659_
	);
	LUT3 #(
		.INIT('h80)
	) name19759 (
		\m0_data_i[5]_pad ,
		_w9171_,
		_w9172_,
		_w21660_
	);
	LUT3 #(
		.INIT('h2a)
	) name19760 (
		\m7_data_i[5]_pad ,
		_w9171_,
		_w9172_,
		_w21661_
	);
	LUT4 #(
		.INIT('h6e7f)
	) name19761 (
		_w9166_,
		_w9169_,
		_w21660_,
		_w21661_,
		_w21662_
	);
	LUT4 #(
		.INIT('h7fff)
	) name19762 (
		_w21653_,
		_w21656_,
		_w21659_,
		_w21662_,
		_w21663_
	);
	LUT3 #(
		.INIT('h2a)
	) name19763 (
		\m3_data_i[6]_pad ,
		_w9171_,
		_w9172_,
		_w21664_
	);
	LUT3 #(
		.INIT('h80)
	) name19764 (
		\m4_data_i[6]_pad ,
		_w9171_,
		_w9172_,
		_w21665_
	);
	LUT4 #(
		.INIT('h9dbf)
	) name19765 (
		_w9166_,
		_w9169_,
		_w21664_,
		_w21665_,
		_w21666_
	);
	LUT3 #(
		.INIT('h80)
	) name19766 (
		\m6_data_i[6]_pad ,
		_w9171_,
		_w9172_,
		_w21667_
	);
	LUT3 #(
		.INIT('h80)
	) name19767 (
		\m2_data_i[6]_pad ,
		_w9171_,
		_w9172_,
		_w21668_
	);
	LUT4 #(
		.INIT('habef)
	) name19768 (
		_w9166_,
		_w9169_,
		_w21667_,
		_w21668_,
		_w21669_
	);
	LUT3 #(
		.INIT('h2a)
	) name19769 (
		\m5_data_i[6]_pad ,
		_w9171_,
		_w9172_,
		_w21670_
	);
	LUT3 #(
		.INIT('h2a)
	) name19770 (
		\m1_data_i[6]_pad ,
		_w9171_,
		_w9172_,
		_w21671_
	);
	LUT4 #(
		.INIT('h57df)
	) name19771 (
		_w9166_,
		_w9169_,
		_w21670_,
		_w21671_,
		_w21672_
	);
	LUT3 #(
		.INIT('h80)
	) name19772 (
		\m0_data_i[6]_pad ,
		_w9171_,
		_w9172_,
		_w21673_
	);
	LUT3 #(
		.INIT('h2a)
	) name19773 (
		\m7_data_i[6]_pad ,
		_w9171_,
		_w9172_,
		_w21674_
	);
	LUT4 #(
		.INIT('h6e7f)
	) name19774 (
		_w9166_,
		_w9169_,
		_w21673_,
		_w21674_,
		_w21675_
	);
	LUT4 #(
		.INIT('h7fff)
	) name19775 (
		_w21666_,
		_w21669_,
		_w21672_,
		_w21675_,
		_w21676_
	);
	LUT3 #(
		.INIT('h2a)
	) name19776 (
		\m3_data_i[7]_pad ,
		_w9171_,
		_w9172_,
		_w21677_
	);
	LUT3 #(
		.INIT('h80)
	) name19777 (
		\m4_data_i[7]_pad ,
		_w9171_,
		_w9172_,
		_w21678_
	);
	LUT4 #(
		.INIT('h9dbf)
	) name19778 (
		_w9166_,
		_w9169_,
		_w21677_,
		_w21678_,
		_w21679_
	);
	LUT3 #(
		.INIT('h80)
	) name19779 (
		\m6_data_i[7]_pad ,
		_w9171_,
		_w9172_,
		_w21680_
	);
	LUT3 #(
		.INIT('h80)
	) name19780 (
		\m2_data_i[7]_pad ,
		_w9171_,
		_w9172_,
		_w21681_
	);
	LUT4 #(
		.INIT('habef)
	) name19781 (
		_w9166_,
		_w9169_,
		_w21680_,
		_w21681_,
		_w21682_
	);
	LUT3 #(
		.INIT('h2a)
	) name19782 (
		\m5_data_i[7]_pad ,
		_w9171_,
		_w9172_,
		_w21683_
	);
	LUT3 #(
		.INIT('h2a)
	) name19783 (
		\m1_data_i[7]_pad ,
		_w9171_,
		_w9172_,
		_w21684_
	);
	LUT4 #(
		.INIT('h57df)
	) name19784 (
		_w9166_,
		_w9169_,
		_w21683_,
		_w21684_,
		_w21685_
	);
	LUT3 #(
		.INIT('h80)
	) name19785 (
		\m0_data_i[7]_pad ,
		_w9171_,
		_w9172_,
		_w21686_
	);
	LUT3 #(
		.INIT('h2a)
	) name19786 (
		\m7_data_i[7]_pad ,
		_w9171_,
		_w9172_,
		_w21687_
	);
	LUT4 #(
		.INIT('h6e7f)
	) name19787 (
		_w9166_,
		_w9169_,
		_w21686_,
		_w21687_,
		_w21688_
	);
	LUT4 #(
		.INIT('h7fff)
	) name19788 (
		_w21679_,
		_w21682_,
		_w21685_,
		_w21688_,
		_w21689_
	);
	LUT3 #(
		.INIT('h2a)
	) name19789 (
		\m3_data_i[8]_pad ,
		_w9171_,
		_w9172_,
		_w21690_
	);
	LUT3 #(
		.INIT('h80)
	) name19790 (
		\m4_data_i[8]_pad ,
		_w9171_,
		_w9172_,
		_w21691_
	);
	LUT4 #(
		.INIT('h9dbf)
	) name19791 (
		_w9166_,
		_w9169_,
		_w21690_,
		_w21691_,
		_w21692_
	);
	LUT3 #(
		.INIT('h80)
	) name19792 (
		\m6_data_i[8]_pad ,
		_w9171_,
		_w9172_,
		_w21693_
	);
	LUT3 #(
		.INIT('h80)
	) name19793 (
		\m2_data_i[8]_pad ,
		_w9171_,
		_w9172_,
		_w21694_
	);
	LUT4 #(
		.INIT('habef)
	) name19794 (
		_w9166_,
		_w9169_,
		_w21693_,
		_w21694_,
		_w21695_
	);
	LUT3 #(
		.INIT('h2a)
	) name19795 (
		\m5_data_i[8]_pad ,
		_w9171_,
		_w9172_,
		_w21696_
	);
	LUT3 #(
		.INIT('h2a)
	) name19796 (
		\m1_data_i[8]_pad ,
		_w9171_,
		_w9172_,
		_w21697_
	);
	LUT4 #(
		.INIT('h57df)
	) name19797 (
		_w9166_,
		_w9169_,
		_w21696_,
		_w21697_,
		_w21698_
	);
	LUT3 #(
		.INIT('h80)
	) name19798 (
		\m0_data_i[8]_pad ,
		_w9171_,
		_w9172_,
		_w21699_
	);
	LUT3 #(
		.INIT('h2a)
	) name19799 (
		\m7_data_i[8]_pad ,
		_w9171_,
		_w9172_,
		_w21700_
	);
	LUT4 #(
		.INIT('h6e7f)
	) name19800 (
		_w9166_,
		_w9169_,
		_w21699_,
		_w21700_,
		_w21701_
	);
	LUT4 #(
		.INIT('h7fff)
	) name19801 (
		_w21692_,
		_w21695_,
		_w21698_,
		_w21701_,
		_w21702_
	);
	LUT3 #(
		.INIT('h2a)
	) name19802 (
		\m3_data_i[9]_pad ,
		_w9171_,
		_w9172_,
		_w21703_
	);
	LUT3 #(
		.INIT('h80)
	) name19803 (
		\m4_data_i[9]_pad ,
		_w9171_,
		_w9172_,
		_w21704_
	);
	LUT4 #(
		.INIT('h9dbf)
	) name19804 (
		_w9166_,
		_w9169_,
		_w21703_,
		_w21704_,
		_w21705_
	);
	LUT3 #(
		.INIT('h80)
	) name19805 (
		\m6_data_i[9]_pad ,
		_w9171_,
		_w9172_,
		_w21706_
	);
	LUT3 #(
		.INIT('h80)
	) name19806 (
		\m2_data_i[9]_pad ,
		_w9171_,
		_w9172_,
		_w21707_
	);
	LUT4 #(
		.INIT('habef)
	) name19807 (
		_w9166_,
		_w9169_,
		_w21706_,
		_w21707_,
		_w21708_
	);
	LUT3 #(
		.INIT('h2a)
	) name19808 (
		\m5_data_i[9]_pad ,
		_w9171_,
		_w9172_,
		_w21709_
	);
	LUT3 #(
		.INIT('h2a)
	) name19809 (
		\m1_data_i[9]_pad ,
		_w9171_,
		_w9172_,
		_w21710_
	);
	LUT4 #(
		.INIT('h57df)
	) name19810 (
		_w9166_,
		_w9169_,
		_w21709_,
		_w21710_,
		_w21711_
	);
	LUT3 #(
		.INIT('h80)
	) name19811 (
		\m0_data_i[9]_pad ,
		_w9171_,
		_w9172_,
		_w21712_
	);
	LUT3 #(
		.INIT('h2a)
	) name19812 (
		\m7_data_i[9]_pad ,
		_w9171_,
		_w9172_,
		_w21713_
	);
	LUT4 #(
		.INIT('h6e7f)
	) name19813 (
		_w9166_,
		_w9169_,
		_w21712_,
		_w21713_,
		_w21714_
	);
	LUT4 #(
		.INIT('h7fff)
	) name19814 (
		_w21705_,
		_w21708_,
		_w21711_,
		_w21714_,
		_w21715_
	);
	LUT3 #(
		.INIT('h2a)
	) name19815 (
		\m3_sel_i[0]_pad ,
		_w9171_,
		_w9172_,
		_w21716_
	);
	LUT3 #(
		.INIT('h80)
	) name19816 (
		\m4_sel_i[0]_pad ,
		_w9171_,
		_w9172_,
		_w21717_
	);
	LUT4 #(
		.INIT('h9dbf)
	) name19817 (
		_w9166_,
		_w9169_,
		_w21716_,
		_w21717_,
		_w21718_
	);
	LUT3 #(
		.INIT('h80)
	) name19818 (
		\m6_sel_i[0]_pad ,
		_w9171_,
		_w9172_,
		_w21719_
	);
	LUT3 #(
		.INIT('h80)
	) name19819 (
		\m2_sel_i[0]_pad ,
		_w9171_,
		_w9172_,
		_w21720_
	);
	LUT4 #(
		.INIT('habef)
	) name19820 (
		_w9166_,
		_w9169_,
		_w21719_,
		_w21720_,
		_w21721_
	);
	LUT3 #(
		.INIT('h2a)
	) name19821 (
		\m5_sel_i[0]_pad ,
		_w9171_,
		_w9172_,
		_w21722_
	);
	LUT3 #(
		.INIT('h2a)
	) name19822 (
		\m1_sel_i[0]_pad ,
		_w9171_,
		_w9172_,
		_w21723_
	);
	LUT4 #(
		.INIT('h57df)
	) name19823 (
		_w9166_,
		_w9169_,
		_w21722_,
		_w21723_,
		_w21724_
	);
	LUT3 #(
		.INIT('h80)
	) name19824 (
		\m0_sel_i[0]_pad ,
		_w9171_,
		_w9172_,
		_w21725_
	);
	LUT3 #(
		.INIT('h2a)
	) name19825 (
		\m7_sel_i[0]_pad ,
		_w9171_,
		_w9172_,
		_w21726_
	);
	LUT4 #(
		.INIT('h6e7f)
	) name19826 (
		_w9166_,
		_w9169_,
		_w21725_,
		_w21726_,
		_w21727_
	);
	LUT4 #(
		.INIT('h7fff)
	) name19827 (
		_w21718_,
		_w21721_,
		_w21724_,
		_w21727_,
		_w21728_
	);
	LUT3 #(
		.INIT('h2a)
	) name19828 (
		\m3_sel_i[1]_pad ,
		_w9171_,
		_w9172_,
		_w21729_
	);
	LUT3 #(
		.INIT('h80)
	) name19829 (
		\m4_sel_i[1]_pad ,
		_w9171_,
		_w9172_,
		_w21730_
	);
	LUT4 #(
		.INIT('h9dbf)
	) name19830 (
		_w9166_,
		_w9169_,
		_w21729_,
		_w21730_,
		_w21731_
	);
	LUT3 #(
		.INIT('h80)
	) name19831 (
		\m6_sel_i[1]_pad ,
		_w9171_,
		_w9172_,
		_w21732_
	);
	LUT3 #(
		.INIT('h80)
	) name19832 (
		\m2_sel_i[1]_pad ,
		_w9171_,
		_w9172_,
		_w21733_
	);
	LUT4 #(
		.INIT('habef)
	) name19833 (
		_w9166_,
		_w9169_,
		_w21732_,
		_w21733_,
		_w21734_
	);
	LUT3 #(
		.INIT('h2a)
	) name19834 (
		\m5_sel_i[1]_pad ,
		_w9171_,
		_w9172_,
		_w21735_
	);
	LUT3 #(
		.INIT('h2a)
	) name19835 (
		\m1_sel_i[1]_pad ,
		_w9171_,
		_w9172_,
		_w21736_
	);
	LUT4 #(
		.INIT('h57df)
	) name19836 (
		_w9166_,
		_w9169_,
		_w21735_,
		_w21736_,
		_w21737_
	);
	LUT3 #(
		.INIT('h80)
	) name19837 (
		\m0_sel_i[1]_pad ,
		_w9171_,
		_w9172_,
		_w21738_
	);
	LUT3 #(
		.INIT('h2a)
	) name19838 (
		\m7_sel_i[1]_pad ,
		_w9171_,
		_w9172_,
		_w21739_
	);
	LUT4 #(
		.INIT('h6e7f)
	) name19839 (
		_w9166_,
		_w9169_,
		_w21738_,
		_w21739_,
		_w21740_
	);
	LUT4 #(
		.INIT('h7fff)
	) name19840 (
		_w21731_,
		_w21734_,
		_w21737_,
		_w21740_,
		_w21741_
	);
	LUT3 #(
		.INIT('h2a)
	) name19841 (
		\m3_sel_i[2]_pad ,
		_w9171_,
		_w9172_,
		_w21742_
	);
	LUT3 #(
		.INIT('h80)
	) name19842 (
		\m4_sel_i[2]_pad ,
		_w9171_,
		_w9172_,
		_w21743_
	);
	LUT4 #(
		.INIT('h9dbf)
	) name19843 (
		_w9166_,
		_w9169_,
		_w21742_,
		_w21743_,
		_w21744_
	);
	LUT3 #(
		.INIT('h80)
	) name19844 (
		\m6_sel_i[2]_pad ,
		_w9171_,
		_w9172_,
		_w21745_
	);
	LUT3 #(
		.INIT('h80)
	) name19845 (
		\m2_sel_i[2]_pad ,
		_w9171_,
		_w9172_,
		_w21746_
	);
	LUT4 #(
		.INIT('habef)
	) name19846 (
		_w9166_,
		_w9169_,
		_w21745_,
		_w21746_,
		_w21747_
	);
	LUT3 #(
		.INIT('h2a)
	) name19847 (
		\m5_sel_i[2]_pad ,
		_w9171_,
		_w9172_,
		_w21748_
	);
	LUT3 #(
		.INIT('h2a)
	) name19848 (
		\m1_sel_i[2]_pad ,
		_w9171_,
		_w9172_,
		_w21749_
	);
	LUT4 #(
		.INIT('h57df)
	) name19849 (
		_w9166_,
		_w9169_,
		_w21748_,
		_w21749_,
		_w21750_
	);
	LUT3 #(
		.INIT('h80)
	) name19850 (
		\m0_sel_i[2]_pad ,
		_w9171_,
		_w9172_,
		_w21751_
	);
	LUT3 #(
		.INIT('h2a)
	) name19851 (
		\m7_sel_i[2]_pad ,
		_w9171_,
		_w9172_,
		_w21752_
	);
	LUT4 #(
		.INIT('h6e7f)
	) name19852 (
		_w9166_,
		_w9169_,
		_w21751_,
		_w21752_,
		_w21753_
	);
	LUT4 #(
		.INIT('h7fff)
	) name19853 (
		_w21744_,
		_w21747_,
		_w21750_,
		_w21753_,
		_w21754_
	);
	LUT3 #(
		.INIT('h2a)
	) name19854 (
		\m3_sel_i[3]_pad ,
		_w9171_,
		_w9172_,
		_w21755_
	);
	LUT3 #(
		.INIT('h80)
	) name19855 (
		\m4_sel_i[3]_pad ,
		_w9171_,
		_w9172_,
		_w21756_
	);
	LUT4 #(
		.INIT('h9dbf)
	) name19856 (
		_w9166_,
		_w9169_,
		_w21755_,
		_w21756_,
		_w21757_
	);
	LUT3 #(
		.INIT('h80)
	) name19857 (
		\m6_sel_i[3]_pad ,
		_w9171_,
		_w9172_,
		_w21758_
	);
	LUT3 #(
		.INIT('h80)
	) name19858 (
		\m2_sel_i[3]_pad ,
		_w9171_,
		_w9172_,
		_w21759_
	);
	LUT4 #(
		.INIT('habef)
	) name19859 (
		_w9166_,
		_w9169_,
		_w21758_,
		_w21759_,
		_w21760_
	);
	LUT3 #(
		.INIT('h2a)
	) name19860 (
		\m5_sel_i[3]_pad ,
		_w9171_,
		_w9172_,
		_w21761_
	);
	LUT3 #(
		.INIT('h2a)
	) name19861 (
		\m1_sel_i[3]_pad ,
		_w9171_,
		_w9172_,
		_w21762_
	);
	LUT4 #(
		.INIT('h57df)
	) name19862 (
		_w9166_,
		_w9169_,
		_w21761_,
		_w21762_,
		_w21763_
	);
	LUT3 #(
		.INIT('h80)
	) name19863 (
		\m0_sel_i[3]_pad ,
		_w9171_,
		_w9172_,
		_w21764_
	);
	LUT3 #(
		.INIT('h2a)
	) name19864 (
		\m7_sel_i[3]_pad ,
		_w9171_,
		_w9172_,
		_w21765_
	);
	LUT4 #(
		.INIT('h6e7f)
	) name19865 (
		_w9166_,
		_w9169_,
		_w21764_,
		_w21765_,
		_w21766_
	);
	LUT4 #(
		.INIT('h7fff)
	) name19866 (
		_w21757_,
		_w21760_,
		_w21763_,
		_w21766_,
		_w21767_
	);
	LUT4 #(
		.INIT('h2a00)
	) name19867 (
		\m5_stb_i_pad ,
		_w9171_,
		_w9172_,
		_w9541_,
		_w21768_
	);
	LUT4 #(
		.INIT('h8000)
	) name19868 (
		\m4_stb_i_pad ,
		_w9171_,
		_w9172_,
		_w9520_,
		_w21769_
	);
	LUT3 #(
		.INIT('h57)
	) name19869 (
		_w9170_,
		_w21768_,
		_w21769_,
		_w21770_
	);
	LUT4 #(
		.INIT('h8000)
	) name19870 (
		\m2_stb_i_pad ,
		_w9171_,
		_w9172_,
		_w9462_,
		_w21771_
	);
	LUT4 #(
		.INIT('h2a00)
	) name19871 (
		\m1_stb_i_pad ,
		_w9171_,
		_w9172_,
		_w9427_,
		_w21772_
	);
	LUT4 #(
		.INIT('h37bf)
	) name19872 (
		_w9166_,
		_w9169_,
		_w21771_,
		_w21772_,
		_w21773_
	);
	LUT4 #(
		.INIT('h2a00)
	) name19873 (
		\m3_stb_i_pad ,
		_w9171_,
		_w9172_,
		_w9494_,
		_w21774_
	);
	LUT4 #(
		.INIT('h2a00)
	) name19874 (
		\m7_stb_i_pad ,
		_w9171_,
		_w9172_,
		_w9608_,
		_w21775_
	);
	LUT4 #(
		.INIT('haebf)
	) name19875 (
		_w9166_,
		_w9169_,
		_w21774_,
		_w21775_,
		_w21776_
	);
	LUT4 #(
		.INIT('h8000)
	) name19876 (
		\m6_stb_i_pad ,
		_w9171_,
		_w9172_,
		_w9576_,
		_w21777_
	);
	LUT4 #(
		.INIT('h8000)
	) name19877 (
		\m0_stb_i_pad ,
		_w9171_,
		_w9172_,
		_w9395_,
		_w21778_
	);
	LUT4 #(
		.INIT('h67ef)
	) name19878 (
		_w9166_,
		_w9169_,
		_w21777_,
		_w21778_,
		_w21779_
	);
	LUT4 #(
		.INIT('h7fff)
	) name19879 (
		_w21770_,
		_w21773_,
		_w21776_,
		_w21779_,
		_w21780_
	);
	LUT3 #(
		.INIT('h2a)
	) name19880 (
		\m3_we_i_pad ,
		_w9171_,
		_w9172_,
		_w21781_
	);
	LUT3 #(
		.INIT('h80)
	) name19881 (
		\m4_we_i_pad ,
		_w9171_,
		_w9172_,
		_w21782_
	);
	LUT4 #(
		.INIT('h9dbf)
	) name19882 (
		_w9166_,
		_w9169_,
		_w21781_,
		_w21782_,
		_w21783_
	);
	LUT3 #(
		.INIT('h80)
	) name19883 (
		\m6_we_i_pad ,
		_w9171_,
		_w9172_,
		_w21784_
	);
	LUT3 #(
		.INIT('h80)
	) name19884 (
		\m2_we_i_pad ,
		_w9171_,
		_w9172_,
		_w21785_
	);
	LUT4 #(
		.INIT('habef)
	) name19885 (
		_w9166_,
		_w9169_,
		_w21784_,
		_w21785_,
		_w21786_
	);
	LUT3 #(
		.INIT('h2a)
	) name19886 (
		\m5_we_i_pad ,
		_w9171_,
		_w9172_,
		_w21787_
	);
	LUT3 #(
		.INIT('h2a)
	) name19887 (
		\m1_we_i_pad ,
		_w9171_,
		_w9172_,
		_w21788_
	);
	LUT4 #(
		.INIT('h57df)
	) name19888 (
		_w9166_,
		_w9169_,
		_w21787_,
		_w21788_,
		_w21789_
	);
	LUT3 #(
		.INIT('h80)
	) name19889 (
		\m0_we_i_pad ,
		_w9171_,
		_w9172_,
		_w21790_
	);
	LUT3 #(
		.INIT('h2a)
	) name19890 (
		\m7_we_i_pad ,
		_w9171_,
		_w9172_,
		_w21791_
	);
	LUT4 #(
		.INIT('h6e7f)
	) name19891 (
		_w9166_,
		_w9169_,
		_w21790_,
		_w21791_,
		_w21792_
	);
	LUT4 #(
		.INIT('h7fff)
	) name19892 (
		_w21783_,
		_w21786_,
		_w21789_,
		_w21792_,
		_w21793_
	);
	LUT3 #(
		.INIT('h2a)
	) name19893 (
		\m1_addr_i[0]_pad ,
		_w9205_,
		_w9206_,
		_w21794_
	);
	LUT3 #(
		.INIT('h80)
	) name19894 (
		\m2_addr_i[0]_pad ,
		_w9205_,
		_w9206_,
		_w21795_
	);
	LUT4 #(
		.INIT('h3b7f)
	) name19895 (
		_w9200_,
		_w9203_,
		_w21794_,
		_w21795_,
		_w21796_
	);
	LUT3 #(
		.INIT('h80)
	) name19896 (
		\m6_addr_i[0]_pad ,
		_w9205_,
		_w9206_,
		_w21797_
	);
	LUT3 #(
		.INIT('h2a)
	) name19897 (
		\m7_addr_i[0]_pad ,
		_w9205_,
		_w9206_,
		_w21798_
	);
	LUT3 #(
		.INIT('h57)
	) name19898 (
		_w9218_,
		_w21797_,
		_w21798_,
		_w21799_
	);
	LUT3 #(
		.INIT('h2a)
	) name19899 (
		\m5_addr_i[0]_pad ,
		_w9205_,
		_w9206_,
		_w21800_
	);
	LUT3 #(
		.INIT('h80)
	) name19900 (
		\m0_addr_i[0]_pad ,
		_w9205_,
		_w9206_,
		_w21801_
	);
	LUT4 #(
		.INIT('h57df)
	) name19901 (
		_w9200_,
		_w9203_,
		_w21800_,
		_w21801_,
		_w21802_
	);
	LUT3 #(
		.INIT('h2a)
	) name19902 (
		\m3_addr_i[0]_pad ,
		_w9205_,
		_w9206_,
		_w21803_
	);
	LUT3 #(
		.INIT('h80)
	) name19903 (
		\m4_addr_i[0]_pad ,
		_w9205_,
		_w9206_,
		_w21804_
	);
	LUT4 #(
		.INIT('h9dbf)
	) name19904 (
		_w9200_,
		_w9203_,
		_w21803_,
		_w21804_,
		_w21805_
	);
	LUT4 #(
		.INIT('h7fff)
	) name19905 (
		_w21796_,
		_w21799_,
		_w21802_,
		_w21805_,
		_w21806_
	);
	LUT3 #(
		.INIT('h2a)
	) name19906 (
		\m3_addr_i[10]_pad ,
		_w9205_,
		_w9206_,
		_w21807_
	);
	LUT3 #(
		.INIT('h80)
	) name19907 (
		\m4_addr_i[10]_pad ,
		_w9205_,
		_w9206_,
		_w21808_
	);
	LUT4 #(
		.INIT('h9dbf)
	) name19908 (
		_w9200_,
		_w9203_,
		_w21807_,
		_w21808_,
		_w21809_
	);
	LUT3 #(
		.INIT('h80)
	) name19909 (
		\m6_addr_i[10]_pad ,
		_w9205_,
		_w9206_,
		_w21810_
	);
	LUT3 #(
		.INIT('h80)
	) name19910 (
		\m2_addr_i[10]_pad ,
		_w9205_,
		_w9206_,
		_w21811_
	);
	LUT4 #(
		.INIT('habef)
	) name19911 (
		_w9200_,
		_w9203_,
		_w21810_,
		_w21811_,
		_w21812_
	);
	LUT3 #(
		.INIT('h2a)
	) name19912 (
		\m5_addr_i[10]_pad ,
		_w9205_,
		_w9206_,
		_w21813_
	);
	LUT3 #(
		.INIT('h2a)
	) name19913 (
		\m1_addr_i[10]_pad ,
		_w9205_,
		_w9206_,
		_w21814_
	);
	LUT4 #(
		.INIT('h57df)
	) name19914 (
		_w9200_,
		_w9203_,
		_w21813_,
		_w21814_,
		_w21815_
	);
	LUT3 #(
		.INIT('h80)
	) name19915 (
		\m0_addr_i[10]_pad ,
		_w9205_,
		_w9206_,
		_w21816_
	);
	LUT3 #(
		.INIT('h2a)
	) name19916 (
		\m7_addr_i[10]_pad ,
		_w9205_,
		_w9206_,
		_w21817_
	);
	LUT4 #(
		.INIT('h6e7f)
	) name19917 (
		_w9200_,
		_w9203_,
		_w21816_,
		_w21817_,
		_w21818_
	);
	LUT4 #(
		.INIT('h7fff)
	) name19918 (
		_w21809_,
		_w21812_,
		_w21815_,
		_w21818_,
		_w21819_
	);
	LUT3 #(
		.INIT('h2a)
	) name19919 (
		\m3_addr_i[11]_pad ,
		_w9205_,
		_w9206_,
		_w21820_
	);
	LUT3 #(
		.INIT('h80)
	) name19920 (
		\m4_addr_i[11]_pad ,
		_w9205_,
		_w9206_,
		_w21821_
	);
	LUT4 #(
		.INIT('h9dbf)
	) name19921 (
		_w9200_,
		_w9203_,
		_w21820_,
		_w21821_,
		_w21822_
	);
	LUT3 #(
		.INIT('h80)
	) name19922 (
		\m6_addr_i[11]_pad ,
		_w9205_,
		_w9206_,
		_w21823_
	);
	LUT3 #(
		.INIT('h80)
	) name19923 (
		\m2_addr_i[11]_pad ,
		_w9205_,
		_w9206_,
		_w21824_
	);
	LUT4 #(
		.INIT('habef)
	) name19924 (
		_w9200_,
		_w9203_,
		_w21823_,
		_w21824_,
		_w21825_
	);
	LUT3 #(
		.INIT('h2a)
	) name19925 (
		\m5_addr_i[11]_pad ,
		_w9205_,
		_w9206_,
		_w21826_
	);
	LUT3 #(
		.INIT('h2a)
	) name19926 (
		\m1_addr_i[11]_pad ,
		_w9205_,
		_w9206_,
		_w21827_
	);
	LUT4 #(
		.INIT('h57df)
	) name19927 (
		_w9200_,
		_w9203_,
		_w21826_,
		_w21827_,
		_w21828_
	);
	LUT3 #(
		.INIT('h80)
	) name19928 (
		\m0_addr_i[11]_pad ,
		_w9205_,
		_w9206_,
		_w21829_
	);
	LUT3 #(
		.INIT('h2a)
	) name19929 (
		\m7_addr_i[11]_pad ,
		_w9205_,
		_w9206_,
		_w21830_
	);
	LUT4 #(
		.INIT('h6e7f)
	) name19930 (
		_w9200_,
		_w9203_,
		_w21829_,
		_w21830_,
		_w21831_
	);
	LUT4 #(
		.INIT('h7fff)
	) name19931 (
		_w21822_,
		_w21825_,
		_w21828_,
		_w21831_,
		_w21832_
	);
	LUT3 #(
		.INIT('h2a)
	) name19932 (
		\m3_addr_i[12]_pad ,
		_w9205_,
		_w9206_,
		_w21833_
	);
	LUT3 #(
		.INIT('h80)
	) name19933 (
		\m4_addr_i[12]_pad ,
		_w9205_,
		_w9206_,
		_w21834_
	);
	LUT4 #(
		.INIT('h9dbf)
	) name19934 (
		_w9200_,
		_w9203_,
		_w21833_,
		_w21834_,
		_w21835_
	);
	LUT3 #(
		.INIT('h80)
	) name19935 (
		\m6_addr_i[12]_pad ,
		_w9205_,
		_w9206_,
		_w21836_
	);
	LUT3 #(
		.INIT('h80)
	) name19936 (
		\m2_addr_i[12]_pad ,
		_w9205_,
		_w9206_,
		_w21837_
	);
	LUT4 #(
		.INIT('habef)
	) name19937 (
		_w9200_,
		_w9203_,
		_w21836_,
		_w21837_,
		_w21838_
	);
	LUT3 #(
		.INIT('h2a)
	) name19938 (
		\m5_addr_i[12]_pad ,
		_w9205_,
		_w9206_,
		_w21839_
	);
	LUT3 #(
		.INIT('h2a)
	) name19939 (
		\m1_addr_i[12]_pad ,
		_w9205_,
		_w9206_,
		_w21840_
	);
	LUT4 #(
		.INIT('h57df)
	) name19940 (
		_w9200_,
		_w9203_,
		_w21839_,
		_w21840_,
		_w21841_
	);
	LUT3 #(
		.INIT('h80)
	) name19941 (
		\m0_addr_i[12]_pad ,
		_w9205_,
		_w9206_,
		_w21842_
	);
	LUT3 #(
		.INIT('h2a)
	) name19942 (
		\m7_addr_i[12]_pad ,
		_w9205_,
		_w9206_,
		_w21843_
	);
	LUT4 #(
		.INIT('h6e7f)
	) name19943 (
		_w9200_,
		_w9203_,
		_w21842_,
		_w21843_,
		_w21844_
	);
	LUT4 #(
		.INIT('h7fff)
	) name19944 (
		_w21835_,
		_w21838_,
		_w21841_,
		_w21844_,
		_w21845_
	);
	LUT3 #(
		.INIT('h2a)
	) name19945 (
		\m3_addr_i[13]_pad ,
		_w9205_,
		_w9206_,
		_w21846_
	);
	LUT3 #(
		.INIT('h80)
	) name19946 (
		\m4_addr_i[13]_pad ,
		_w9205_,
		_w9206_,
		_w21847_
	);
	LUT4 #(
		.INIT('h9dbf)
	) name19947 (
		_w9200_,
		_w9203_,
		_w21846_,
		_w21847_,
		_w21848_
	);
	LUT3 #(
		.INIT('h80)
	) name19948 (
		\m6_addr_i[13]_pad ,
		_w9205_,
		_w9206_,
		_w21849_
	);
	LUT3 #(
		.INIT('h80)
	) name19949 (
		\m2_addr_i[13]_pad ,
		_w9205_,
		_w9206_,
		_w21850_
	);
	LUT4 #(
		.INIT('habef)
	) name19950 (
		_w9200_,
		_w9203_,
		_w21849_,
		_w21850_,
		_w21851_
	);
	LUT3 #(
		.INIT('h2a)
	) name19951 (
		\m5_addr_i[13]_pad ,
		_w9205_,
		_w9206_,
		_w21852_
	);
	LUT3 #(
		.INIT('h2a)
	) name19952 (
		\m1_addr_i[13]_pad ,
		_w9205_,
		_w9206_,
		_w21853_
	);
	LUT4 #(
		.INIT('h57df)
	) name19953 (
		_w9200_,
		_w9203_,
		_w21852_,
		_w21853_,
		_w21854_
	);
	LUT3 #(
		.INIT('h80)
	) name19954 (
		\m0_addr_i[13]_pad ,
		_w9205_,
		_w9206_,
		_w21855_
	);
	LUT3 #(
		.INIT('h2a)
	) name19955 (
		\m7_addr_i[13]_pad ,
		_w9205_,
		_w9206_,
		_w21856_
	);
	LUT4 #(
		.INIT('h6e7f)
	) name19956 (
		_w9200_,
		_w9203_,
		_w21855_,
		_w21856_,
		_w21857_
	);
	LUT4 #(
		.INIT('h7fff)
	) name19957 (
		_w21848_,
		_w21851_,
		_w21854_,
		_w21857_,
		_w21858_
	);
	LUT3 #(
		.INIT('h2a)
	) name19958 (
		\m3_addr_i[14]_pad ,
		_w9205_,
		_w9206_,
		_w21859_
	);
	LUT3 #(
		.INIT('h80)
	) name19959 (
		\m4_addr_i[14]_pad ,
		_w9205_,
		_w9206_,
		_w21860_
	);
	LUT4 #(
		.INIT('h9dbf)
	) name19960 (
		_w9200_,
		_w9203_,
		_w21859_,
		_w21860_,
		_w21861_
	);
	LUT3 #(
		.INIT('h80)
	) name19961 (
		\m6_addr_i[14]_pad ,
		_w9205_,
		_w9206_,
		_w21862_
	);
	LUT3 #(
		.INIT('h80)
	) name19962 (
		\m2_addr_i[14]_pad ,
		_w9205_,
		_w9206_,
		_w21863_
	);
	LUT4 #(
		.INIT('habef)
	) name19963 (
		_w9200_,
		_w9203_,
		_w21862_,
		_w21863_,
		_w21864_
	);
	LUT3 #(
		.INIT('h2a)
	) name19964 (
		\m5_addr_i[14]_pad ,
		_w9205_,
		_w9206_,
		_w21865_
	);
	LUT3 #(
		.INIT('h2a)
	) name19965 (
		\m1_addr_i[14]_pad ,
		_w9205_,
		_w9206_,
		_w21866_
	);
	LUT4 #(
		.INIT('h57df)
	) name19966 (
		_w9200_,
		_w9203_,
		_w21865_,
		_w21866_,
		_w21867_
	);
	LUT3 #(
		.INIT('h80)
	) name19967 (
		\m0_addr_i[14]_pad ,
		_w9205_,
		_w9206_,
		_w21868_
	);
	LUT3 #(
		.INIT('h2a)
	) name19968 (
		\m7_addr_i[14]_pad ,
		_w9205_,
		_w9206_,
		_w21869_
	);
	LUT4 #(
		.INIT('h6e7f)
	) name19969 (
		_w9200_,
		_w9203_,
		_w21868_,
		_w21869_,
		_w21870_
	);
	LUT4 #(
		.INIT('h7fff)
	) name19970 (
		_w21861_,
		_w21864_,
		_w21867_,
		_w21870_,
		_w21871_
	);
	LUT3 #(
		.INIT('h2a)
	) name19971 (
		\m3_addr_i[15]_pad ,
		_w9205_,
		_w9206_,
		_w21872_
	);
	LUT3 #(
		.INIT('h80)
	) name19972 (
		\m4_addr_i[15]_pad ,
		_w9205_,
		_w9206_,
		_w21873_
	);
	LUT4 #(
		.INIT('h9dbf)
	) name19973 (
		_w9200_,
		_w9203_,
		_w21872_,
		_w21873_,
		_w21874_
	);
	LUT3 #(
		.INIT('h80)
	) name19974 (
		\m6_addr_i[15]_pad ,
		_w9205_,
		_w9206_,
		_w21875_
	);
	LUT3 #(
		.INIT('h80)
	) name19975 (
		\m2_addr_i[15]_pad ,
		_w9205_,
		_w9206_,
		_w21876_
	);
	LUT4 #(
		.INIT('habef)
	) name19976 (
		_w9200_,
		_w9203_,
		_w21875_,
		_w21876_,
		_w21877_
	);
	LUT3 #(
		.INIT('h2a)
	) name19977 (
		\m5_addr_i[15]_pad ,
		_w9205_,
		_w9206_,
		_w21878_
	);
	LUT3 #(
		.INIT('h2a)
	) name19978 (
		\m1_addr_i[15]_pad ,
		_w9205_,
		_w9206_,
		_w21879_
	);
	LUT4 #(
		.INIT('h57df)
	) name19979 (
		_w9200_,
		_w9203_,
		_w21878_,
		_w21879_,
		_w21880_
	);
	LUT3 #(
		.INIT('h80)
	) name19980 (
		\m0_addr_i[15]_pad ,
		_w9205_,
		_w9206_,
		_w21881_
	);
	LUT3 #(
		.INIT('h2a)
	) name19981 (
		\m7_addr_i[15]_pad ,
		_w9205_,
		_w9206_,
		_w21882_
	);
	LUT4 #(
		.INIT('h6e7f)
	) name19982 (
		_w9200_,
		_w9203_,
		_w21881_,
		_w21882_,
		_w21883_
	);
	LUT4 #(
		.INIT('h7fff)
	) name19983 (
		_w21874_,
		_w21877_,
		_w21880_,
		_w21883_,
		_w21884_
	);
	LUT3 #(
		.INIT('h2a)
	) name19984 (
		\m3_addr_i[16]_pad ,
		_w9205_,
		_w9206_,
		_w21885_
	);
	LUT3 #(
		.INIT('h80)
	) name19985 (
		\m4_addr_i[16]_pad ,
		_w9205_,
		_w9206_,
		_w21886_
	);
	LUT4 #(
		.INIT('h9dbf)
	) name19986 (
		_w9200_,
		_w9203_,
		_w21885_,
		_w21886_,
		_w21887_
	);
	LUT3 #(
		.INIT('h80)
	) name19987 (
		\m6_addr_i[16]_pad ,
		_w9205_,
		_w9206_,
		_w21888_
	);
	LUT3 #(
		.INIT('h80)
	) name19988 (
		\m2_addr_i[16]_pad ,
		_w9205_,
		_w9206_,
		_w21889_
	);
	LUT4 #(
		.INIT('habef)
	) name19989 (
		_w9200_,
		_w9203_,
		_w21888_,
		_w21889_,
		_w21890_
	);
	LUT3 #(
		.INIT('h2a)
	) name19990 (
		\m5_addr_i[16]_pad ,
		_w9205_,
		_w9206_,
		_w21891_
	);
	LUT3 #(
		.INIT('h2a)
	) name19991 (
		\m1_addr_i[16]_pad ,
		_w9205_,
		_w9206_,
		_w21892_
	);
	LUT4 #(
		.INIT('h57df)
	) name19992 (
		_w9200_,
		_w9203_,
		_w21891_,
		_w21892_,
		_w21893_
	);
	LUT3 #(
		.INIT('h80)
	) name19993 (
		\m0_addr_i[16]_pad ,
		_w9205_,
		_w9206_,
		_w21894_
	);
	LUT3 #(
		.INIT('h2a)
	) name19994 (
		\m7_addr_i[16]_pad ,
		_w9205_,
		_w9206_,
		_w21895_
	);
	LUT4 #(
		.INIT('h6e7f)
	) name19995 (
		_w9200_,
		_w9203_,
		_w21894_,
		_w21895_,
		_w21896_
	);
	LUT4 #(
		.INIT('h7fff)
	) name19996 (
		_w21887_,
		_w21890_,
		_w21893_,
		_w21896_,
		_w21897_
	);
	LUT3 #(
		.INIT('h2a)
	) name19997 (
		\m3_addr_i[17]_pad ,
		_w9205_,
		_w9206_,
		_w21898_
	);
	LUT3 #(
		.INIT('h80)
	) name19998 (
		\m4_addr_i[17]_pad ,
		_w9205_,
		_w9206_,
		_w21899_
	);
	LUT4 #(
		.INIT('h9dbf)
	) name19999 (
		_w9200_,
		_w9203_,
		_w21898_,
		_w21899_,
		_w21900_
	);
	LUT3 #(
		.INIT('h80)
	) name20000 (
		\m6_addr_i[17]_pad ,
		_w9205_,
		_w9206_,
		_w21901_
	);
	LUT3 #(
		.INIT('h80)
	) name20001 (
		\m2_addr_i[17]_pad ,
		_w9205_,
		_w9206_,
		_w21902_
	);
	LUT4 #(
		.INIT('habef)
	) name20002 (
		_w9200_,
		_w9203_,
		_w21901_,
		_w21902_,
		_w21903_
	);
	LUT3 #(
		.INIT('h2a)
	) name20003 (
		\m5_addr_i[17]_pad ,
		_w9205_,
		_w9206_,
		_w21904_
	);
	LUT3 #(
		.INIT('h2a)
	) name20004 (
		\m1_addr_i[17]_pad ,
		_w9205_,
		_w9206_,
		_w21905_
	);
	LUT4 #(
		.INIT('h57df)
	) name20005 (
		_w9200_,
		_w9203_,
		_w21904_,
		_w21905_,
		_w21906_
	);
	LUT3 #(
		.INIT('h80)
	) name20006 (
		\m0_addr_i[17]_pad ,
		_w9205_,
		_w9206_,
		_w21907_
	);
	LUT3 #(
		.INIT('h2a)
	) name20007 (
		\m7_addr_i[17]_pad ,
		_w9205_,
		_w9206_,
		_w21908_
	);
	LUT4 #(
		.INIT('h6e7f)
	) name20008 (
		_w9200_,
		_w9203_,
		_w21907_,
		_w21908_,
		_w21909_
	);
	LUT4 #(
		.INIT('h7fff)
	) name20009 (
		_w21900_,
		_w21903_,
		_w21906_,
		_w21909_,
		_w21910_
	);
	LUT3 #(
		.INIT('h2a)
	) name20010 (
		\m3_addr_i[18]_pad ,
		_w9205_,
		_w9206_,
		_w21911_
	);
	LUT3 #(
		.INIT('h80)
	) name20011 (
		\m4_addr_i[18]_pad ,
		_w9205_,
		_w9206_,
		_w21912_
	);
	LUT4 #(
		.INIT('h9dbf)
	) name20012 (
		_w9200_,
		_w9203_,
		_w21911_,
		_w21912_,
		_w21913_
	);
	LUT3 #(
		.INIT('h80)
	) name20013 (
		\m6_addr_i[18]_pad ,
		_w9205_,
		_w9206_,
		_w21914_
	);
	LUT3 #(
		.INIT('h80)
	) name20014 (
		\m2_addr_i[18]_pad ,
		_w9205_,
		_w9206_,
		_w21915_
	);
	LUT4 #(
		.INIT('habef)
	) name20015 (
		_w9200_,
		_w9203_,
		_w21914_,
		_w21915_,
		_w21916_
	);
	LUT3 #(
		.INIT('h2a)
	) name20016 (
		\m5_addr_i[18]_pad ,
		_w9205_,
		_w9206_,
		_w21917_
	);
	LUT3 #(
		.INIT('h2a)
	) name20017 (
		\m1_addr_i[18]_pad ,
		_w9205_,
		_w9206_,
		_w21918_
	);
	LUT4 #(
		.INIT('h57df)
	) name20018 (
		_w9200_,
		_w9203_,
		_w21917_,
		_w21918_,
		_w21919_
	);
	LUT3 #(
		.INIT('h80)
	) name20019 (
		\m0_addr_i[18]_pad ,
		_w9205_,
		_w9206_,
		_w21920_
	);
	LUT3 #(
		.INIT('h2a)
	) name20020 (
		\m7_addr_i[18]_pad ,
		_w9205_,
		_w9206_,
		_w21921_
	);
	LUT4 #(
		.INIT('h6e7f)
	) name20021 (
		_w9200_,
		_w9203_,
		_w21920_,
		_w21921_,
		_w21922_
	);
	LUT4 #(
		.INIT('h7fff)
	) name20022 (
		_w21913_,
		_w21916_,
		_w21919_,
		_w21922_,
		_w21923_
	);
	LUT3 #(
		.INIT('h2a)
	) name20023 (
		\m3_addr_i[19]_pad ,
		_w9205_,
		_w9206_,
		_w21924_
	);
	LUT3 #(
		.INIT('h80)
	) name20024 (
		\m4_addr_i[19]_pad ,
		_w9205_,
		_w9206_,
		_w21925_
	);
	LUT4 #(
		.INIT('h9dbf)
	) name20025 (
		_w9200_,
		_w9203_,
		_w21924_,
		_w21925_,
		_w21926_
	);
	LUT3 #(
		.INIT('h80)
	) name20026 (
		\m6_addr_i[19]_pad ,
		_w9205_,
		_w9206_,
		_w21927_
	);
	LUT3 #(
		.INIT('h80)
	) name20027 (
		\m2_addr_i[19]_pad ,
		_w9205_,
		_w9206_,
		_w21928_
	);
	LUT4 #(
		.INIT('habef)
	) name20028 (
		_w9200_,
		_w9203_,
		_w21927_,
		_w21928_,
		_w21929_
	);
	LUT3 #(
		.INIT('h2a)
	) name20029 (
		\m5_addr_i[19]_pad ,
		_w9205_,
		_w9206_,
		_w21930_
	);
	LUT3 #(
		.INIT('h2a)
	) name20030 (
		\m1_addr_i[19]_pad ,
		_w9205_,
		_w9206_,
		_w21931_
	);
	LUT4 #(
		.INIT('h57df)
	) name20031 (
		_w9200_,
		_w9203_,
		_w21930_,
		_w21931_,
		_w21932_
	);
	LUT3 #(
		.INIT('h80)
	) name20032 (
		\m0_addr_i[19]_pad ,
		_w9205_,
		_w9206_,
		_w21933_
	);
	LUT3 #(
		.INIT('h2a)
	) name20033 (
		\m7_addr_i[19]_pad ,
		_w9205_,
		_w9206_,
		_w21934_
	);
	LUT4 #(
		.INIT('h6e7f)
	) name20034 (
		_w9200_,
		_w9203_,
		_w21933_,
		_w21934_,
		_w21935_
	);
	LUT4 #(
		.INIT('h7fff)
	) name20035 (
		_w21926_,
		_w21929_,
		_w21932_,
		_w21935_,
		_w21936_
	);
	LUT3 #(
		.INIT('h2a)
	) name20036 (
		\m3_addr_i[1]_pad ,
		_w9205_,
		_w9206_,
		_w21937_
	);
	LUT3 #(
		.INIT('h80)
	) name20037 (
		\m4_addr_i[1]_pad ,
		_w9205_,
		_w9206_,
		_w21938_
	);
	LUT4 #(
		.INIT('h9dbf)
	) name20038 (
		_w9200_,
		_w9203_,
		_w21937_,
		_w21938_,
		_w21939_
	);
	LUT3 #(
		.INIT('h80)
	) name20039 (
		\m6_addr_i[1]_pad ,
		_w9205_,
		_w9206_,
		_w21940_
	);
	LUT3 #(
		.INIT('h80)
	) name20040 (
		\m2_addr_i[1]_pad ,
		_w9205_,
		_w9206_,
		_w21941_
	);
	LUT4 #(
		.INIT('habef)
	) name20041 (
		_w9200_,
		_w9203_,
		_w21940_,
		_w21941_,
		_w21942_
	);
	LUT3 #(
		.INIT('h2a)
	) name20042 (
		\m5_addr_i[1]_pad ,
		_w9205_,
		_w9206_,
		_w21943_
	);
	LUT3 #(
		.INIT('h2a)
	) name20043 (
		\m1_addr_i[1]_pad ,
		_w9205_,
		_w9206_,
		_w21944_
	);
	LUT4 #(
		.INIT('h57df)
	) name20044 (
		_w9200_,
		_w9203_,
		_w21943_,
		_w21944_,
		_w21945_
	);
	LUT3 #(
		.INIT('h80)
	) name20045 (
		\m0_addr_i[1]_pad ,
		_w9205_,
		_w9206_,
		_w21946_
	);
	LUT3 #(
		.INIT('h2a)
	) name20046 (
		\m7_addr_i[1]_pad ,
		_w9205_,
		_w9206_,
		_w21947_
	);
	LUT4 #(
		.INIT('h6e7f)
	) name20047 (
		_w9200_,
		_w9203_,
		_w21946_,
		_w21947_,
		_w21948_
	);
	LUT4 #(
		.INIT('h7fff)
	) name20048 (
		_w21939_,
		_w21942_,
		_w21945_,
		_w21948_,
		_w21949_
	);
	LUT3 #(
		.INIT('h2a)
	) name20049 (
		\m3_addr_i[20]_pad ,
		_w9205_,
		_w9206_,
		_w21950_
	);
	LUT3 #(
		.INIT('h80)
	) name20050 (
		\m4_addr_i[20]_pad ,
		_w9205_,
		_w9206_,
		_w21951_
	);
	LUT4 #(
		.INIT('h9dbf)
	) name20051 (
		_w9200_,
		_w9203_,
		_w21950_,
		_w21951_,
		_w21952_
	);
	LUT3 #(
		.INIT('h80)
	) name20052 (
		\m6_addr_i[20]_pad ,
		_w9205_,
		_w9206_,
		_w21953_
	);
	LUT3 #(
		.INIT('h80)
	) name20053 (
		\m2_addr_i[20]_pad ,
		_w9205_,
		_w9206_,
		_w21954_
	);
	LUT4 #(
		.INIT('habef)
	) name20054 (
		_w9200_,
		_w9203_,
		_w21953_,
		_w21954_,
		_w21955_
	);
	LUT3 #(
		.INIT('h2a)
	) name20055 (
		\m5_addr_i[20]_pad ,
		_w9205_,
		_w9206_,
		_w21956_
	);
	LUT3 #(
		.INIT('h2a)
	) name20056 (
		\m1_addr_i[20]_pad ,
		_w9205_,
		_w9206_,
		_w21957_
	);
	LUT4 #(
		.INIT('h57df)
	) name20057 (
		_w9200_,
		_w9203_,
		_w21956_,
		_w21957_,
		_w21958_
	);
	LUT3 #(
		.INIT('h80)
	) name20058 (
		\m0_addr_i[20]_pad ,
		_w9205_,
		_w9206_,
		_w21959_
	);
	LUT3 #(
		.INIT('h2a)
	) name20059 (
		\m7_addr_i[20]_pad ,
		_w9205_,
		_w9206_,
		_w21960_
	);
	LUT4 #(
		.INIT('h6e7f)
	) name20060 (
		_w9200_,
		_w9203_,
		_w21959_,
		_w21960_,
		_w21961_
	);
	LUT4 #(
		.INIT('h7fff)
	) name20061 (
		_w21952_,
		_w21955_,
		_w21958_,
		_w21961_,
		_w21962_
	);
	LUT3 #(
		.INIT('h2a)
	) name20062 (
		\m3_addr_i[21]_pad ,
		_w9205_,
		_w9206_,
		_w21963_
	);
	LUT3 #(
		.INIT('h80)
	) name20063 (
		\m4_addr_i[21]_pad ,
		_w9205_,
		_w9206_,
		_w21964_
	);
	LUT4 #(
		.INIT('h9dbf)
	) name20064 (
		_w9200_,
		_w9203_,
		_w21963_,
		_w21964_,
		_w21965_
	);
	LUT3 #(
		.INIT('h80)
	) name20065 (
		\m6_addr_i[21]_pad ,
		_w9205_,
		_w9206_,
		_w21966_
	);
	LUT3 #(
		.INIT('h80)
	) name20066 (
		\m2_addr_i[21]_pad ,
		_w9205_,
		_w9206_,
		_w21967_
	);
	LUT4 #(
		.INIT('habef)
	) name20067 (
		_w9200_,
		_w9203_,
		_w21966_,
		_w21967_,
		_w21968_
	);
	LUT3 #(
		.INIT('h2a)
	) name20068 (
		\m5_addr_i[21]_pad ,
		_w9205_,
		_w9206_,
		_w21969_
	);
	LUT3 #(
		.INIT('h2a)
	) name20069 (
		\m1_addr_i[21]_pad ,
		_w9205_,
		_w9206_,
		_w21970_
	);
	LUT4 #(
		.INIT('h57df)
	) name20070 (
		_w9200_,
		_w9203_,
		_w21969_,
		_w21970_,
		_w21971_
	);
	LUT3 #(
		.INIT('h80)
	) name20071 (
		\m0_addr_i[21]_pad ,
		_w9205_,
		_w9206_,
		_w21972_
	);
	LUT3 #(
		.INIT('h2a)
	) name20072 (
		\m7_addr_i[21]_pad ,
		_w9205_,
		_w9206_,
		_w21973_
	);
	LUT4 #(
		.INIT('h6e7f)
	) name20073 (
		_w9200_,
		_w9203_,
		_w21972_,
		_w21973_,
		_w21974_
	);
	LUT4 #(
		.INIT('h7fff)
	) name20074 (
		_w21965_,
		_w21968_,
		_w21971_,
		_w21974_,
		_w21975_
	);
	LUT3 #(
		.INIT('h2a)
	) name20075 (
		\m3_addr_i[22]_pad ,
		_w9205_,
		_w9206_,
		_w21976_
	);
	LUT3 #(
		.INIT('h80)
	) name20076 (
		\m4_addr_i[22]_pad ,
		_w9205_,
		_w9206_,
		_w21977_
	);
	LUT4 #(
		.INIT('h9dbf)
	) name20077 (
		_w9200_,
		_w9203_,
		_w21976_,
		_w21977_,
		_w21978_
	);
	LUT3 #(
		.INIT('h80)
	) name20078 (
		\m6_addr_i[22]_pad ,
		_w9205_,
		_w9206_,
		_w21979_
	);
	LUT3 #(
		.INIT('h80)
	) name20079 (
		\m2_addr_i[22]_pad ,
		_w9205_,
		_w9206_,
		_w21980_
	);
	LUT4 #(
		.INIT('habef)
	) name20080 (
		_w9200_,
		_w9203_,
		_w21979_,
		_w21980_,
		_w21981_
	);
	LUT3 #(
		.INIT('h2a)
	) name20081 (
		\m5_addr_i[22]_pad ,
		_w9205_,
		_w9206_,
		_w21982_
	);
	LUT3 #(
		.INIT('h2a)
	) name20082 (
		\m1_addr_i[22]_pad ,
		_w9205_,
		_w9206_,
		_w21983_
	);
	LUT4 #(
		.INIT('h57df)
	) name20083 (
		_w9200_,
		_w9203_,
		_w21982_,
		_w21983_,
		_w21984_
	);
	LUT3 #(
		.INIT('h80)
	) name20084 (
		\m0_addr_i[22]_pad ,
		_w9205_,
		_w9206_,
		_w21985_
	);
	LUT3 #(
		.INIT('h2a)
	) name20085 (
		\m7_addr_i[22]_pad ,
		_w9205_,
		_w9206_,
		_w21986_
	);
	LUT4 #(
		.INIT('h6e7f)
	) name20086 (
		_w9200_,
		_w9203_,
		_w21985_,
		_w21986_,
		_w21987_
	);
	LUT4 #(
		.INIT('h7fff)
	) name20087 (
		_w21978_,
		_w21981_,
		_w21984_,
		_w21987_,
		_w21988_
	);
	LUT3 #(
		.INIT('h2a)
	) name20088 (
		\m3_addr_i[23]_pad ,
		_w9205_,
		_w9206_,
		_w21989_
	);
	LUT3 #(
		.INIT('h80)
	) name20089 (
		\m4_addr_i[23]_pad ,
		_w9205_,
		_w9206_,
		_w21990_
	);
	LUT4 #(
		.INIT('h9dbf)
	) name20090 (
		_w9200_,
		_w9203_,
		_w21989_,
		_w21990_,
		_w21991_
	);
	LUT3 #(
		.INIT('h80)
	) name20091 (
		\m6_addr_i[23]_pad ,
		_w9205_,
		_w9206_,
		_w21992_
	);
	LUT3 #(
		.INIT('h80)
	) name20092 (
		\m2_addr_i[23]_pad ,
		_w9205_,
		_w9206_,
		_w21993_
	);
	LUT4 #(
		.INIT('habef)
	) name20093 (
		_w9200_,
		_w9203_,
		_w21992_,
		_w21993_,
		_w21994_
	);
	LUT3 #(
		.INIT('h2a)
	) name20094 (
		\m5_addr_i[23]_pad ,
		_w9205_,
		_w9206_,
		_w21995_
	);
	LUT3 #(
		.INIT('h2a)
	) name20095 (
		\m1_addr_i[23]_pad ,
		_w9205_,
		_w9206_,
		_w21996_
	);
	LUT4 #(
		.INIT('h57df)
	) name20096 (
		_w9200_,
		_w9203_,
		_w21995_,
		_w21996_,
		_w21997_
	);
	LUT3 #(
		.INIT('h80)
	) name20097 (
		\m0_addr_i[23]_pad ,
		_w9205_,
		_w9206_,
		_w21998_
	);
	LUT3 #(
		.INIT('h2a)
	) name20098 (
		\m7_addr_i[23]_pad ,
		_w9205_,
		_w9206_,
		_w21999_
	);
	LUT4 #(
		.INIT('h6e7f)
	) name20099 (
		_w9200_,
		_w9203_,
		_w21998_,
		_w21999_,
		_w22000_
	);
	LUT4 #(
		.INIT('h7fff)
	) name20100 (
		_w21991_,
		_w21994_,
		_w21997_,
		_w22000_,
		_w22001_
	);
	LUT3 #(
		.INIT('h2a)
	) name20101 (
		\m3_addr_i[24]_pad ,
		_w9205_,
		_w9206_,
		_w22002_
	);
	LUT3 #(
		.INIT('h80)
	) name20102 (
		\m4_addr_i[24]_pad ,
		_w9205_,
		_w9206_,
		_w22003_
	);
	LUT4 #(
		.INIT('h9dbf)
	) name20103 (
		_w9200_,
		_w9203_,
		_w22002_,
		_w22003_,
		_w22004_
	);
	LUT3 #(
		.INIT('h2a)
	) name20104 (
		\m5_addr_i[24]_pad ,
		_w9205_,
		_w9206_,
		_w22005_
	);
	LUT3 #(
		.INIT('h80)
	) name20105 (
		\m2_addr_i[24]_pad ,
		_w9205_,
		_w9206_,
		_w22006_
	);
	LUT4 #(
		.INIT('h9bdf)
	) name20106 (
		_w9200_,
		_w9203_,
		_w22005_,
		_w22006_,
		_w22007_
	);
	LUT3 #(
		.INIT('h80)
	) name20107 (
		\m6_addr_i[24]_pad ,
		_w9205_,
		_w9206_,
		_w22008_
	);
	LUT3 #(
		.INIT('h2a)
	) name20108 (
		\m1_addr_i[24]_pad ,
		_w9205_,
		_w9206_,
		_w22009_
	);
	LUT4 #(
		.INIT('h67ef)
	) name20109 (
		_w9200_,
		_w9203_,
		_w22008_,
		_w22009_,
		_w22010_
	);
	LUT3 #(
		.INIT('h80)
	) name20110 (
		\m0_addr_i[24]_pad ,
		_w9205_,
		_w9206_,
		_w22011_
	);
	LUT3 #(
		.INIT('h2a)
	) name20111 (
		\m7_addr_i[24]_pad ,
		_w9205_,
		_w9206_,
		_w22012_
	);
	LUT4 #(
		.INIT('h6e7f)
	) name20112 (
		_w9200_,
		_w9203_,
		_w22011_,
		_w22012_,
		_w22013_
	);
	LUT4 #(
		.INIT('h7fff)
	) name20113 (
		_w22004_,
		_w22007_,
		_w22010_,
		_w22013_,
		_w22014_
	);
	LUT3 #(
		.INIT('h2a)
	) name20114 (
		\m3_addr_i[25]_pad ,
		_w9205_,
		_w9206_,
		_w22015_
	);
	LUT3 #(
		.INIT('h80)
	) name20115 (
		\m4_addr_i[25]_pad ,
		_w9205_,
		_w9206_,
		_w22016_
	);
	LUT4 #(
		.INIT('h9dbf)
	) name20116 (
		_w9200_,
		_w9203_,
		_w22015_,
		_w22016_,
		_w22017_
	);
	LUT3 #(
		.INIT('h2a)
	) name20117 (
		\m5_addr_i[25]_pad ,
		_w9205_,
		_w9206_,
		_w22018_
	);
	LUT3 #(
		.INIT('h80)
	) name20118 (
		\m2_addr_i[25]_pad ,
		_w9205_,
		_w9206_,
		_w22019_
	);
	LUT4 #(
		.INIT('h9bdf)
	) name20119 (
		_w9200_,
		_w9203_,
		_w22018_,
		_w22019_,
		_w22020_
	);
	LUT3 #(
		.INIT('h80)
	) name20120 (
		\m6_addr_i[25]_pad ,
		_w9205_,
		_w9206_,
		_w22021_
	);
	LUT3 #(
		.INIT('h2a)
	) name20121 (
		\m1_addr_i[25]_pad ,
		_w9205_,
		_w9206_,
		_w22022_
	);
	LUT4 #(
		.INIT('h67ef)
	) name20122 (
		_w9200_,
		_w9203_,
		_w22021_,
		_w22022_,
		_w22023_
	);
	LUT3 #(
		.INIT('h80)
	) name20123 (
		\m0_addr_i[25]_pad ,
		_w9205_,
		_w9206_,
		_w22024_
	);
	LUT3 #(
		.INIT('h2a)
	) name20124 (
		\m7_addr_i[25]_pad ,
		_w9205_,
		_w9206_,
		_w22025_
	);
	LUT4 #(
		.INIT('h6e7f)
	) name20125 (
		_w9200_,
		_w9203_,
		_w22024_,
		_w22025_,
		_w22026_
	);
	LUT4 #(
		.INIT('h7fff)
	) name20126 (
		_w22017_,
		_w22020_,
		_w22023_,
		_w22026_,
		_w22027_
	);
	LUT3 #(
		.INIT('h2a)
	) name20127 (
		\m3_addr_i[26]_pad ,
		_w9205_,
		_w9206_,
		_w22028_
	);
	LUT3 #(
		.INIT('h80)
	) name20128 (
		\m4_addr_i[26]_pad ,
		_w9205_,
		_w9206_,
		_w22029_
	);
	LUT4 #(
		.INIT('h9dbf)
	) name20129 (
		_w9200_,
		_w9203_,
		_w22028_,
		_w22029_,
		_w22030_
	);
	LUT3 #(
		.INIT('h2a)
	) name20130 (
		\m5_addr_i[26]_pad ,
		_w9205_,
		_w9206_,
		_w22031_
	);
	LUT3 #(
		.INIT('h80)
	) name20131 (
		\m2_addr_i[26]_pad ,
		_w9205_,
		_w9206_,
		_w22032_
	);
	LUT4 #(
		.INIT('h9bdf)
	) name20132 (
		_w9200_,
		_w9203_,
		_w22031_,
		_w22032_,
		_w22033_
	);
	LUT3 #(
		.INIT('h80)
	) name20133 (
		\m6_addr_i[26]_pad ,
		_w9205_,
		_w9206_,
		_w22034_
	);
	LUT3 #(
		.INIT('h2a)
	) name20134 (
		\m1_addr_i[26]_pad ,
		_w9205_,
		_w9206_,
		_w22035_
	);
	LUT4 #(
		.INIT('h67ef)
	) name20135 (
		_w9200_,
		_w9203_,
		_w22034_,
		_w22035_,
		_w22036_
	);
	LUT3 #(
		.INIT('h80)
	) name20136 (
		\m0_addr_i[26]_pad ,
		_w9205_,
		_w9206_,
		_w22037_
	);
	LUT3 #(
		.INIT('h2a)
	) name20137 (
		\m7_addr_i[26]_pad ,
		_w9205_,
		_w9206_,
		_w22038_
	);
	LUT4 #(
		.INIT('h6e7f)
	) name20138 (
		_w9200_,
		_w9203_,
		_w22037_,
		_w22038_,
		_w22039_
	);
	LUT4 #(
		.INIT('h7fff)
	) name20139 (
		_w22030_,
		_w22033_,
		_w22036_,
		_w22039_,
		_w22040_
	);
	LUT3 #(
		.INIT('h2a)
	) name20140 (
		\m3_addr_i[27]_pad ,
		_w9205_,
		_w9206_,
		_w22041_
	);
	LUT3 #(
		.INIT('h80)
	) name20141 (
		\m4_addr_i[27]_pad ,
		_w9205_,
		_w9206_,
		_w22042_
	);
	LUT4 #(
		.INIT('h9dbf)
	) name20142 (
		_w9200_,
		_w9203_,
		_w22041_,
		_w22042_,
		_w22043_
	);
	LUT3 #(
		.INIT('h2a)
	) name20143 (
		\m5_addr_i[27]_pad ,
		_w9205_,
		_w9206_,
		_w22044_
	);
	LUT3 #(
		.INIT('h80)
	) name20144 (
		\m2_addr_i[27]_pad ,
		_w9205_,
		_w9206_,
		_w22045_
	);
	LUT4 #(
		.INIT('h9bdf)
	) name20145 (
		_w9200_,
		_w9203_,
		_w22044_,
		_w22045_,
		_w22046_
	);
	LUT3 #(
		.INIT('h80)
	) name20146 (
		\m6_addr_i[27]_pad ,
		_w9205_,
		_w9206_,
		_w22047_
	);
	LUT3 #(
		.INIT('h2a)
	) name20147 (
		\m1_addr_i[27]_pad ,
		_w9205_,
		_w9206_,
		_w22048_
	);
	LUT4 #(
		.INIT('h67ef)
	) name20148 (
		_w9200_,
		_w9203_,
		_w22047_,
		_w22048_,
		_w22049_
	);
	LUT3 #(
		.INIT('h80)
	) name20149 (
		\m0_addr_i[27]_pad ,
		_w9205_,
		_w9206_,
		_w22050_
	);
	LUT3 #(
		.INIT('h2a)
	) name20150 (
		\m7_addr_i[27]_pad ,
		_w9205_,
		_w9206_,
		_w22051_
	);
	LUT4 #(
		.INIT('h6e7f)
	) name20151 (
		_w9200_,
		_w9203_,
		_w22050_,
		_w22051_,
		_w22052_
	);
	LUT4 #(
		.INIT('h7fff)
	) name20152 (
		_w22043_,
		_w22046_,
		_w22049_,
		_w22052_,
		_w22053_
	);
	LUT3 #(
		.INIT('h2a)
	) name20153 (
		\m3_addr_i[28]_pad ,
		_w9205_,
		_w9206_,
		_w22054_
	);
	LUT3 #(
		.INIT('h80)
	) name20154 (
		\m4_addr_i[28]_pad ,
		_w9205_,
		_w9206_,
		_w22055_
	);
	LUT4 #(
		.INIT('h9dbf)
	) name20155 (
		_w9200_,
		_w9203_,
		_w22054_,
		_w22055_,
		_w22056_
	);
	LUT3 #(
		.INIT('h2a)
	) name20156 (
		\m5_addr_i[28]_pad ,
		_w9205_,
		_w9206_,
		_w22057_
	);
	LUT3 #(
		.INIT('h80)
	) name20157 (
		\m2_addr_i[28]_pad ,
		_w9205_,
		_w9206_,
		_w22058_
	);
	LUT4 #(
		.INIT('h9bdf)
	) name20158 (
		_w9200_,
		_w9203_,
		_w22057_,
		_w22058_,
		_w22059_
	);
	LUT3 #(
		.INIT('h80)
	) name20159 (
		\m6_addr_i[28]_pad ,
		_w9205_,
		_w9206_,
		_w22060_
	);
	LUT3 #(
		.INIT('h2a)
	) name20160 (
		\m1_addr_i[28]_pad ,
		_w9205_,
		_w9206_,
		_w22061_
	);
	LUT4 #(
		.INIT('h67ef)
	) name20161 (
		_w9200_,
		_w9203_,
		_w22060_,
		_w22061_,
		_w22062_
	);
	LUT3 #(
		.INIT('h80)
	) name20162 (
		\m0_addr_i[28]_pad ,
		_w9205_,
		_w9206_,
		_w22063_
	);
	LUT3 #(
		.INIT('h2a)
	) name20163 (
		\m7_addr_i[28]_pad ,
		_w9205_,
		_w9206_,
		_w22064_
	);
	LUT4 #(
		.INIT('h6e7f)
	) name20164 (
		_w9200_,
		_w9203_,
		_w22063_,
		_w22064_,
		_w22065_
	);
	LUT4 #(
		.INIT('h7fff)
	) name20165 (
		_w22056_,
		_w22059_,
		_w22062_,
		_w22065_,
		_w22066_
	);
	LUT3 #(
		.INIT('h2a)
	) name20166 (
		\m3_addr_i[29]_pad ,
		_w9205_,
		_w9206_,
		_w22067_
	);
	LUT3 #(
		.INIT('h80)
	) name20167 (
		\m4_addr_i[29]_pad ,
		_w9205_,
		_w9206_,
		_w22068_
	);
	LUT4 #(
		.INIT('h9dbf)
	) name20168 (
		_w9200_,
		_w9203_,
		_w22067_,
		_w22068_,
		_w22069_
	);
	LUT3 #(
		.INIT('h2a)
	) name20169 (
		\m5_addr_i[29]_pad ,
		_w9205_,
		_w9206_,
		_w22070_
	);
	LUT3 #(
		.INIT('h80)
	) name20170 (
		\m2_addr_i[29]_pad ,
		_w9205_,
		_w9206_,
		_w22071_
	);
	LUT4 #(
		.INIT('h9bdf)
	) name20171 (
		_w9200_,
		_w9203_,
		_w22070_,
		_w22071_,
		_w22072_
	);
	LUT3 #(
		.INIT('h80)
	) name20172 (
		\m6_addr_i[29]_pad ,
		_w9205_,
		_w9206_,
		_w22073_
	);
	LUT3 #(
		.INIT('h2a)
	) name20173 (
		\m1_addr_i[29]_pad ,
		_w9205_,
		_w9206_,
		_w22074_
	);
	LUT4 #(
		.INIT('h67ef)
	) name20174 (
		_w9200_,
		_w9203_,
		_w22073_,
		_w22074_,
		_w22075_
	);
	LUT3 #(
		.INIT('h80)
	) name20175 (
		\m0_addr_i[29]_pad ,
		_w9205_,
		_w9206_,
		_w22076_
	);
	LUT3 #(
		.INIT('h2a)
	) name20176 (
		\m7_addr_i[29]_pad ,
		_w9205_,
		_w9206_,
		_w22077_
	);
	LUT4 #(
		.INIT('h6e7f)
	) name20177 (
		_w9200_,
		_w9203_,
		_w22076_,
		_w22077_,
		_w22078_
	);
	LUT4 #(
		.INIT('h7fff)
	) name20178 (
		_w22069_,
		_w22072_,
		_w22075_,
		_w22078_,
		_w22079_
	);
	LUT3 #(
		.INIT('h2a)
	) name20179 (
		\m3_addr_i[2]_pad ,
		_w9205_,
		_w9206_,
		_w22080_
	);
	LUT3 #(
		.INIT('h80)
	) name20180 (
		\m4_addr_i[2]_pad ,
		_w9205_,
		_w9206_,
		_w22081_
	);
	LUT4 #(
		.INIT('h9dbf)
	) name20181 (
		_w9200_,
		_w9203_,
		_w22080_,
		_w22081_,
		_w22082_
	);
	LUT3 #(
		.INIT('h80)
	) name20182 (
		\m6_addr_i[2]_pad ,
		_w9205_,
		_w9206_,
		_w22083_
	);
	LUT3 #(
		.INIT('h80)
	) name20183 (
		\m2_addr_i[2]_pad ,
		_w9205_,
		_w9206_,
		_w22084_
	);
	LUT4 #(
		.INIT('habef)
	) name20184 (
		_w9200_,
		_w9203_,
		_w22083_,
		_w22084_,
		_w22085_
	);
	LUT3 #(
		.INIT('h2a)
	) name20185 (
		\m5_addr_i[2]_pad ,
		_w9205_,
		_w9206_,
		_w22086_
	);
	LUT3 #(
		.INIT('h2a)
	) name20186 (
		\m1_addr_i[2]_pad ,
		_w9205_,
		_w9206_,
		_w22087_
	);
	LUT4 #(
		.INIT('h57df)
	) name20187 (
		_w9200_,
		_w9203_,
		_w22086_,
		_w22087_,
		_w22088_
	);
	LUT3 #(
		.INIT('h80)
	) name20188 (
		\m0_addr_i[2]_pad ,
		_w9205_,
		_w9206_,
		_w22089_
	);
	LUT3 #(
		.INIT('h2a)
	) name20189 (
		\m7_addr_i[2]_pad ,
		_w9205_,
		_w9206_,
		_w22090_
	);
	LUT4 #(
		.INIT('h6e7f)
	) name20190 (
		_w9200_,
		_w9203_,
		_w22089_,
		_w22090_,
		_w22091_
	);
	LUT4 #(
		.INIT('h7fff)
	) name20191 (
		_w22082_,
		_w22085_,
		_w22088_,
		_w22091_,
		_w22092_
	);
	LUT3 #(
		.INIT('h2a)
	) name20192 (
		\m3_addr_i[30]_pad ,
		_w9205_,
		_w9206_,
		_w22093_
	);
	LUT3 #(
		.INIT('h80)
	) name20193 (
		\m4_addr_i[30]_pad ,
		_w9205_,
		_w9206_,
		_w22094_
	);
	LUT4 #(
		.INIT('h9dbf)
	) name20194 (
		_w9200_,
		_w9203_,
		_w22093_,
		_w22094_,
		_w22095_
	);
	LUT3 #(
		.INIT('h2a)
	) name20195 (
		\m5_addr_i[30]_pad ,
		_w9205_,
		_w9206_,
		_w22096_
	);
	LUT3 #(
		.INIT('h80)
	) name20196 (
		\m2_addr_i[30]_pad ,
		_w9205_,
		_w9206_,
		_w22097_
	);
	LUT4 #(
		.INIT('h9bdf)
	) name20197 (
		_w9200_,
		_w9203_,
		_w22096_,
		_w22097_,
		_w22098_
	);
	LUT3 #(
		.INIT('h80)
	) name20198 (
		\m6_addr_i[30]_pad ,
		_w9205_,
		_w9206_,
		_w22099_
	);
	LUT3 #(
		.INIT('h2a)
	) name20199 (
		\m1_addr_i[30]_pad ,
		_w9205_,
		_w9206_,
		_w22100_
	);
	LUT4 #(
		.INIT('h67ef)
	) name20200 (
		_w9200_,
		_w9203_,
		_w22099_,
		_w22100_,
		_w22101_
	);
	LUT3 #(
		.INIT('h80)
	) name20201 (
		\m0_addr_i[30]_pad ,
		_w9205_,
		_w9206_,
		_w22102_
	);
	LUT3 #(
		.INIT('h2a)
	) name20202 (
		\m7_addr_i[30]_pad ,
		_w9205_,
		_w9206_,
		_w22103_
	);
	LUT4 #(
		.INIT('h6e7f)
	) name20203 (
		_w9200_,
		_w9203_,
		_w22102_,
		_w22103_,
		_w22104_
	);
	LUT4 #(
		.INIT('h7fff)
	) name20204 (
		_w22095_,
		_w22098_,
		_w22101_,
		_w22104_,
		_w22105_
	);
	LUT3 #(
		.INIT('h2a)
	) name20205 (
		\m3_addr_i[31]_pad ,
		_w9205_,
		_w9206_,
		_w22106_
	);
	LUT3 #(
		.INIT('h80)
	) name20206 (
		\m4_addr_i[31]_pad ,
		_w9205_,
		_w9206_,
		_w22107_
	);
	LUT4 #(
		.INIT('h9dbf)
	) name20207 (
		_w9200_,
		_w9203_,
		_w22106_,
		_w22107_,
		_w22108_
	);
	LUT3 #(
		.INIT('h2a)
	) name20208 (
		\m5_addr_i[31]_pad ,
		_w9205_,
		_w9206_,
		_w22109_
	);
	LUT3 #(
		.INIT('h80)
	) name20209 (
		\m2_addr_i[31]_pad ,
		_w9205_,
		_w9206_,
		_w22110_
	);
	LUT4 #(
		.INIT('h9bdf)
	) name20210 (
		_w9200_,
		_w9203_,
		_w22109_,
		_w22110_,
		_w22111_
	);
	LUT3 #(
		.INIT('h80)
	) name20211 (
		\m6_addr_i[31]_pad ,
		_w9205_,
		_w9206_,
		_w22112_
	);
	LUT3 #(
		.INIT('h2a)
	) name20212 (
		\m1_addr_i[31]_pad ,
		_w9205_,
		_w9206_,
		_w22113_
	);
	LUT4 #(
		.INIT('h67ef)
	) name20213 (
		_w9200_,
		_w9203_,
		_w22112_,
		_w22113_,
		_w22114_
	);
	LUT3 #(
		.INIT('h80)
	) name20214 (
		\m0_addr_i[31]_pad ,
		_w9205_,
		_w9206_,
		_w22115_
	);
	LUT3 #(
		.INIT('h2a)
	) name20215 (
		\m7_addr_i[31]_pad ,
		_w9205_,
		_w9206_,
		_w22116_
	);
	LUT4 #(
		.INIT('h6e7f)
	) name20216 (
		_w9200_,
		_w9203_,
		_w22115_,
		_w22116_,
		_w22117_
	);
	LUT4 #(
		.INIT('h7fff)
	) name20217 (
		_w22108_,
		_w22111_,
		_w22114_,
		_w22117_,
		_w22118_
	);
	LUT3 #(
		.INIT('h2a)
	) name20218 (
		\m3_addr_i[3]_pad ,
		_w9205_,
		_w9206_,
		_w22119_
	);
	LUT3 #(
		.INIT('h80)
	) name20219 (
		\m4_addr_i[3]_pad ,
		_w9205_,
		_w9206_,
		_w22120_
	);
	LUT4 #(
		.INIT('h9dbf)
	) name20220 (
		_w9200_,
		_w9203_,
		_w22119_,
		_w22120_,
		_w22121_
	);
	LUT3 #(
		.INIT('h80)
	) name20221 (
		\m6_addr_i[3]_pad ,
		_w9205_,
		_w9206_,
		_w22122_
	);
	LUT3 #(
		.INIT('h80)
	) name20222 (
		\m2_addr_i[3]_pad ,
		_w9205_,
		_w9206_,
		_w22123_
	);
	LUT4 #(
		.INIT('habef)
	) name20223 (
		_w9200_,
		_w9203_,
		_w22122_,
		_w22123_,
		_w22124_
	);
	LUT3 #(
		.INIT('h2a)
	) name20224 (
		\m5_addr_i[3]_pad ,
		_w9205_,
		_w9206_,
		_w22125_
	);
	LUT3 #(
		.INIT('h2a)
	) name20225 (
		\m1_addr_i[3]_pad ,
		_w9205_,
		_w9206_,
		_w22126_
	);
	LUT4 #(
		.INIT('h57df)
	) name20226 (
		_w9200_,
		_w9203_,
		_w22125_,
		_w22126_,
		_w22127_
	);
	LUT3 #(
		.INIT('h80)
	) name20227 (
		\m0_addr_i[3]_pad ,
		_w9205_,
		_w9206_,
		_w22128_
	);
	LUT3 #(
		.INIT('h2a)
	) name20228 (
		\m7_addr_i[3]_pad ,
		_w9205_,
		_w9206_,
		_w22129_
	);
	LUT4 #(
		.INIT('h6e7f)
	) name20229 (
		_w9200_,
		_w9203_,
		_w22128_,
		_w22129_,
		_w22130_
	);
	LUT4 #(
		.INIT('h7fff)
	) name20230 (
		_w22121_,
		_w22124_,
		_w22127_,
		_w22130_,
		_w22131_
	);
	LUT3 #(
		.INIT('h2a)
	) name20231 (
		\m3_addr_i[4]_pad ,
		_w9205_,
		_w9206_,
		_w22132_
	);
	LUT3 #(
		.INIT('h80)
	) name20232 (
		\m4_addr_i[4]_pad ,
		_w9205_,
		_w9206_,
		_w22133_
	);
	LUT4 #(
		.INIT('h9dbf)
	) name20233 (
		_w9200_,
		_w9203_,
		_w22132_,
		_w22133_,
		_w22134_
	);
	LUT3 #(
		.INIT('h80)
	) name20234 (
		\m6_addr_i[4]_pad ,
		_w9205_,
		_w9206_,
		_w22135_
	);
	LUT3 #(
		.INIT('h80)
	) name20235 (
		\m2_addr_i[4]_pad ,
		_w9205_,
		_w9206_,
		_w22136_
	);
	LUT4 #(
		.INIT('habef)
	) name20236 (
		_w9200_,
		_w9203_,
		_w22135_,
		_w22136_,
		_w22137_
	);
	LUT3 #(
		.INIT('h2a)
	) name20237 (
		\m5_addr_i[4]_pad ,
		_w9205_,
		_w9206_,
		_w22138_
	);
	LUT3 #(
		.INIT('h2a)
	) name20238 (
		\m1_addr_i[4]_pad ,
		_w9205_,
		_w9206_,
		_w22139_
	);
	LUT4 #(
		.INIT('h57df)
	) name20239 (
		_w9200_,
		_w9203_,
		_w22138_,
		_w22139_,
		_w22140_
	);
	LUT3 #(
		.INIT('h80)
	) name20240 (
		\m0_addr_i[4]_pad ,
		_w9205_,
		_w9206_,
		_w22141_
	);
	LUT3 #(
		.INIT('h2a)
	) name20241 (
		\m7_addr_i[4]_pad ,
		_w9205_,
		_w9206_,
		_w22142_
	);
	LUT4 #(
		.INIT('h6e7f)
	) name20242 (
		_w9200_,
		_w9203_,
		_w22141_,
		_w22142_,
		_w22143_
	);
	LUT4 #(
		.INIT('h7fff)
	) name20243 (
		_w22134_,
		_w22137_,
		_w22140_,
		_w22143_,
		_w22144_
	);
	LUT3 #(
		.INIT('h2a)
	) name20244 (
		\m3_addr_i[5]_pad ,
		_w9205_,
		_w9206_,
		_w22145_
	);
	LUT3 #(
		.INIT('h80)
	) name20245 (
		\m4_addr_i[5]_pad ,
		_w9205_,
		_w9206_,
		_w22146_
	);
	LUT4 #(
		.INIT('h9dbf)
	) name20246 (
		_w9200_,
		_w9203_,
		_w22145_,
		_w22146_,
		_w22147_
	);
	LUT3 #(
		.INIT('h80)
	) name20247 (
		\m6_addr_i[5]_pad ,
		_w9205_,
		_w9206_,
		_w22148_
	);
	LUT3 #(
		.INIT('h80)
	) name20248 (
		\m2_addr_i[5]_pad ,
		_w9205_,
		_w9206_,
		_w22149_
	);
	LUT4 #(
		.INIT('habef)
	) name20249 (
		_w9200_,
		_w9203_,
		_w22148_,
		_w22149_,
		_w22150_
	);
	LUT3 #(
		.INIT('h2a)
	) name20250 (
		\m5_addr_i[5]_pad ,
		_w9205_,
		_w9206_,
		_w22151_
	);
	LUT3 #(
		.INIT('h2a)
	) name20251 (
		\m1_addr_i[5]_pad ,
		_w9205_,
		_w9206_,
		_w22152_
	);
	LUT4 #(
		.INIT('h57df)
	) name20252 (
		_w9200_,
		_w9203_,
		_w22151_,
		_w22152_,
		_w22153_
	);
	LUT3 #(
		.INIT('h80)
	) name20253 (
		\m0_addr_i[5]_pad ,
		_w9205_,
		_w9206_,
		_w22154_
	);
	LUT3 #(
		.INIT('h2a)
	) name20254 (
		\m7_addr_i[5]_pad ,
		_w9205_,
		_w9206_,
		_w22155_
	);
	LUT4 #(
		.INIT('h6e7f)
	) name20255 (
		_w9200_,
		_w9203_,
		_w22154_,
		_w22155_,
		_w22156_
	);
	LUT4 #(
		.INIT('h7fff)
	) name20256 (
		_w22147_,
		_w22150_,
		_w22153_,
		_w22156_,
		_w22157_
	);
	LUT3 #(
		.INIT('h2a)
	) name20257 (
		\m3_addr_i[6]_pad ,
		_w9205_,
		_w9206_,
		_w22158_
	);
	LUT3 #(
		.INIT('h80)
	) name20258 (
		\m4_addr_i[6]_pad ,
		_w9205_,
		_w9206_,
		_w22159_
	);
	LUT4 #(
		.INIT('h9dbf)
	) name20259 (
		_w9200_,
		_w9203_,
		_w22158_,
		_w22159_,
		_w22160_
	);
	LUT3 #(
		.INIT('h80)
	) name20260 (
		\m6_addr_i[6]_pad ,
		_w9205_,
		_w9206_,
		_w22161_
	);
	LUT3 #(
		.INIT('h80)
	) name20261 (
		\m2_addr_i[6]_pad ,
		_w9205_,
		_w9206_,
		_w22162_
	);
	LUT4 #(
		.INIT('habef)
	) name20262 (
		_w9200_,
		_w9203_,
		_w22161_,
		_w22162_,
		_w22163_
	);
	LUT3 #(
		.INIT('h2a)
	) name20263 (
		\m5_addr_i[6]_pad ,
		_w9205_,
		_w9206_,
		_w22164_
	);
	LUT3 #(
		.INIT('h2a)
	) name20264 (
		\m1_addr_i[6]_pad ,
		_w9205_,
		_w9206_,
		_w22165_
	);
	LUT4 #(
		.INIT('h57df)
	) name20265 (
		_w9200_,
		_w9203_,
		_w22164_,
		_w22165_,
		_w22166_
	);
	LUT3 #(
		.INIT('h80)
	) name20266 (
		\m0_addr_i[6]_pad ,
		_w9205_,
		_w9206_,
		_w22167_
	);
	LUT3 #(
		.INIT('h2a)
	) name20267 (
		\m7_addr_i[6]_pad ,
		_w9205_,
		_w9206_,
		_w22168_
	);
	LUT4 #(
		.INIT('h6e7f)
	) name20268 (
		_w9200_,
		_w9203_,
		_w22167_,
		_w22168_,
		_w22169_
	);
	LUT4 #(
		.INIT('h7fff)
	) name20269 (
		_w22160_,
		_w22163_,
		_w22166_,
		_w22169_,
		_w22170_
	);
	LUT3 #(
		.INIT('h2a)
	) name20270 (
		\m3_addr_i[7]_pad ,
		_w9205_,
		_w9206_,
		_w22171_
	);
	LUT3 #(
		.INIT('h80)
	) name20271 (
		\m4_addr_i[7]_pad ,
		_w9205_,
		_w9206_,
		_w22172_
	);
	LUT4 #(
		.INIT('h9dbf)
	) name20272 (
		_w9200_,
		_w9203_,
		_w22171_,
		_w22172_,
		_w22173_
	);
	LUT3 #(
		.INIT('h80)
	) name20273 (
		\m6_addr_i[7]_pad ,
		_w9205_,
		_w9206_,
		_w22174_
	);
	LUT3 #(
		.INIT('h80)
	) name20274 (
		\m2_addr_i[7]_pad ,
		_w9205_,
		_w9206_,
		_w22175_
	);
	LUT4 #(
		.INIT('habef)
	) name20275 (
		_w9200_,
		_w9203_,
		_w22174_,
		_w22175_,
		_w22176_
	);
	LUT3 #(
		.INIT('h2a)
	) name20276 (
		\m5_addr_i[7]_pad ,
		_w9205_,
		_w9206_,
		_w22177_
	);
	LUT3 #(
		.INIT('h2a)
	) name20277 (
		\m1_addr_i[7]_pad ,
		_w9205_,
		_w9206_,
		_w22178_
	);
	LUT4 #(
		.INIT('h57df)
	) name20278 (
		_w9200_,
		_w9203_,
		_w22177_,
		_w22178_,
		_w22179_
	);
	LUT3 #(
		.INIT('h80)
	) name20279 (
		\m0_addr_i[7]_pad ,
		_w9205_,
		_w9206_,
		_w22180_
	);
	LUT3 #(
		.INIT('h2a)
	) name20280 (
		\m7_addr_i[7]_pad ,
		_w9205_,
		_w9206_,
		_w22181_
	);
	LUT4 #(
		.INIT('h6e7f)
	) name20281 (
		_w9200_,
		_w9203_,
		_w22180_,
		_w22181_,
		_w22182_
	);
	LUT4 #(
		.INIT('h7fff)
	) name20282 (
		_w22173_,
		_w22176_,
		_w22179_,
		_w22182_,
		_w22183_
	);
	LUT3 #(
		.INIT('h2a)
	) name20283 (
		\m3_addr_i[8]_pad ,
		_w9205_,
		_w9206_,
		_w22184_
	);
	LUT3 #(
		.INIT('h80)
	) name20284 (
		\m4_addr_i[8]_pad ,
		_w9205_,
		_w9206_,
		_w22185_
	);
	LUT4 #(
		.INIT('h9dbf)
	) name20285 (
		_w9200_,
		_w9203_,
		_w22184_,
		_w22185_,
		_w22186_
	);
	LUT3 #(
		.INIT('h80)
	) name20286 (
		\m6_addr_i[8]_pad ,
		_w9205_,
		_w9206_,
		_w22187_
	);
	LUT3 #(
		.INIT('h80)
	) name20287 (
		\m2_addr_i[8]_pad ,
		_w9205_,
		_w9206_,
		_w22188_
	);
	LUT4 #(
		.INIT('habef)
	) name20288 (
		_w9200_,
		_w9203_,
		_w22187_,
		_w22188_,
		_w22189_
	);
	LUT3 #(
		.INIT('h2a)
	) name20289 (
		\m5_addr_i[8]_pad ,
		_w9205_,
		_w9206_,
		_w22190_
	);
	LUT3 #(
		.INIT('h2a)
	) name20290 (
		\m1_addr_i[8]_pad ,
		_w9205_,
		_w9206_,
		_w22191_
	);
	LUT4 #(
		.INIT('h57df)
	) name20291 (
		_w9200_,
		_w9203_,
		_w22190_,
		_w22191_,
		_w22192_
	);
	LUT3 #(
		.INIT('h80)
	) name20292 (
		\m0_addr_i[8]_pad ,
		_w9205_,
		_w9206_,
		_w22193_
	);
	LUT3 #(
		.INIT('h2a)
	) name20293 (
		\m7_addr_i[8]_pad ,
		_w9205_,
		_w9206_,
		_w22194_
	);
	LUT4 #(
		.INIT('h6e7f)
	) name20294 (
		_w9200_,
		_w9203_,
		_w22193_,
		_w22194_,
		_w22195_
	);
	LUT4 #(
		.INIT('h7fff)
	) name20295 (
		_w22186_,
		_w22189_,
		_w22192_,
		_w22195_,
		_w22196_
	);
	LUT3 #(
		.INIT('h2a)
	) name20296 (
		\m3_addr_i[9]_pad ,
		_w9205_,
		_w9206_,
		_w22197_
	);
	LUT3 #(
		.INIT('h80)
	) name20297 (
		\m4_addr_i[9]_pad ,
		_w9205_,
		_w9206_,
		_w22198_
	);
	LUT4 #(
		.INIT('h9dbf)
	) name20298 (
		_w9200_,
		_w9203_,
		_w22197_,
		_w22198_,
		_w22199_
	);
	LUT3 #(
		.INIT('h80)
	) name20299 (
		\m6_addr_i[9]_pad ,
		_w9205_,
		_w9206_,
		_w22200_
	);
	LUT3 #(
		.INIT('h80)
	) name20300 (
		\m2_addr_i[9]_pad ,
		_w9205_,
		_w9206_,
		_w22201_
	);
	LUT4 #(
		.INIT('habef)
	) name20301 (
		_w9200_,
		_w9203_,
		_w22200_,
		_w22201_,
		_w22202_
	);
	LUT3 #(
		.INIT('h2a)
	) name20302 (
		\m5_addr_i[9]_pad ,
		_w9205_,
		_w9206_,
		_w22203_
	);
	LUT3 #(
		.INIT('h2a)
	) name20303 (
		\m1_addr_i[9]_pad ,
		_w9205_,
		_w9206_,
		_w22204_
	);
	LUT4 #(
		.INIT('h57df)
	) name20304 (
		_w9200_,
		_w9203_,
		_w22203_,
		_w22204_,
		_w22205_
	);
	LUT3 #(
		.INIT('h80)
	) name20305 (
		\m0_addr_i[9]_pad ,
		_w9205_,
		_w9206_,
		_w22206_
	);
	LUT3 #(
		.INIT('h2a)
	) name20306 (
		\m7_addr_i[9]_pad ,
		_w9205_,
		_w9206_,
		_w22207_
	);
	LUT4 #(
		.INIT('h6e7f)
	) name20307 (
		_w9200_,
		_w9203_,
		_w22206_,
		_w22207_,
		_w22208_
	);
	LUT4 #(
		.INIT('h7fff)
	) name20308 (
		_w22199_,
		_w22202_,
		_w22205_,
		_w22208_,
		_w22209_
	);
	LUT3 #(
		.INIT('h2a)
	) name20309 (
		\m3_data_i[0]_pad ,
		_w9205_,
		_w9206_,
		_w22210_
	);
	LUT3 #(
		.INIT('h80)
	) name20310 (
		\m4_data_i[0]_pad ,
		_w9205_,
		_w9206_,
		_w22211_
	);
	LUT4 #(
		.INIT('h9dbf)
	) name20311 (
		_w9200_,
		_w9203_,
		_w22210_,
		_w22211_,
		_w22212_
	);
	LUT3 #(
		.INIT('h80)
	) name20312 (
		\m6_data_i[0]_pad ,
		_w9205_,
		_w9206_,
		_w22213_
	);
	LUT3 #(
		.INIT('h80)
	) name20313 (
		\m2_data_i[0]_pad ,
		_w9205_,
		_w9206_,
		_w22214_
	);
	LUT4 #(
		.INIT('habef)
	) name20314 (
		_w9200_,
		_w9203_,
		_w22213_,
		_w22214_,
		_w22215_
	);
	LUT3 #(
		.INIT('h2a)
	) name20315 (
		\m5_data_i[0]_pad ,
		_w9205_,
		_w9206_,
		_w22216_
	);
	LUT3 #(
		.INIT('h2a)
	) name20316 (
		\m1_data_i[0]_pad ,
		_w9205_,
		_w9206_,
		_w22217_
	);
	LUT4 #(
		.INIT('h57df)
	) name20317 (
		_w9200_,
		_w9203_,
		_w22216_,
		_w22217_,
		_w22218_
	);
	LUT3 #(
		.INIT('h80)
	) name20318 (
		\m0_data_i[0]_pad ,
		_w9205_,
		_w9206_,
		_w22219_
	);
	LUT3 #(
		.INIT('h2a)
	) name20319 (
		\m7_data_i[0]_pad ,
		_w9205_,
		_w9206_,
		_w22220_
	);
	LUT4 #(
		.INIT('h6e7f)
	) name20320 (
		_w9200_,
		_w9203_,
		_w22219_,
		_w22220_,
		_w22221_
	);
	LUT4 #(
		.INIT('h7fff)
	) name20321 (
		_w22212_,
		_w22215_,
		_w22218_,
		_w22221_,
		_w22222_
	);
	LUT3 #(
		.INIT('h2a)
	) name20322 (
		\m3_data_i[10]_pad ,
		_w9205_,
		_w9206_,
		_w22223_
	);
	LUT3 #(
		.INIT('h80)
	) name20323 (
		\m4_data_i[10]_pad ,
		_w9205_,
		_w9206_,
		_w22224_
	);
	LUT4 #(
		.INIT('h9dbf)
	) name20324 (
		_w9200_,
		_w9203_,
		_w22223_,
		_w22224_,
		_w22225_
	);
	LUT3 #(
		.INIT('h80)
	) name20325 (
		\m6_data_i[10]_pad ,
		_w9205_,
		_w9206_,
		_w22226_
	);
	LUT3 #(
		.INIT('h80)
	) name20326 (
		\m2_data_i[10]_pad ,
		_w9205_,
		_w9206_,
		_w22227_
	);
	LUT4 #(
		.INIT('habef)
	) name20327 (
		_w9200_,
		_w9203_,
		_w22226_,
		_w22227_,
		_w22228_
	);
	LUT3 #(
		.INIT('h2a)
	) name20328 (
		\m5_data_i[10]_pad ,
		_w9205_,
		_w9206_,
		_w22229_
	);
	LUT3 #(
		.INIT('h2a)
	) name20329 (
		\m1_data_i[10]_pad ,
		_w9205_,
		_w9206_,
		_w22230_
	);
	LUT4 #(
		.INIT('h57df)
	) name20330 (
		_w9200_,
		_w9203_,
		_w22229_,
		_w22230_,
		_w22231_
	);
	LUT3 #(
		.INIT('h80)
	) name20331 (
		\m0_data_i[10]_pad ,
		_w9205_,
		_w9206_,
		_w22232_
	);
	LUT3 #(
		.INIT('h2a)
	) name20332 (
		\m7_data_i[10]_pad ,
		_w9205_,
		_w9206_,
		_w22233_
	);
	LUT4 #(
		.INIT('h6e7f)
	) name20333 (
		_w9200_,
		_w9203_,
		_w22232_,
		_w22233_,
		_w22234_
	);
	LUT4 #(
		.INIT('h7fff)
	) name20334 (
		_w22225_,
		_w22228_,
		_w22231_,
		_w22234_,
		_w22235_
	);
	LUT3 #(
		.INIT('h2a)
	) name20335 (
		\m3_data_i[11]_pad ,
		_w9205_,
		_w9206_,
		_w22236_
	);
	LUT3 #(
		.INIT('h80)
	) name20336 (
		\m4_data_i[11]_pad ,
		_w9205_,
		_w9206_,
		_w22237_
	);
	LUT4 #(
		.INIT('h9dbf)
	) name20337 (
		_w9200_,
		_w9203_,
		_w22236_,
		_w22237_,
		_w22238_
	);
	LUT3 #(
		.INIT('h80)
	) name20338 (
		\m6_data_i[11]_pad ,
		_w9205_,
		_w9206_,
		_w22239_
	);
	LUT3 #(
		.INIT('h80)
	) name20339 (
		\m2_data_i[11]_pad ,
		_w9205_,
		_w9206_,
		_w22240_
	);
	LUT4 #(
		.INIT('habef)
	) name20340 (
		_w9200_,
		_w9203_,
		_w22239_,
		_w22240_,
		_w22241_
	);
	LUT3 #(
		.INIT('h2a)
	) name20341 (
		\m5_data_i[11]_pad ,
		_w9205_,
		_w9206_,
		_w22242_
	);
	LUT3 #(
		.INIT('h2a)
	) name20342 (
		\m1_data_i[11]_pad ,
		_w9205_,
		_w9206_,
		_w22243_
	);
	LUT4 #(
		.INIT('h57df)
	) name20343 (
		_w9200_,
		_w9203_,
		_w22242_,
		_w22243_,
		_w22244_
	);
	LUT3 #(
		.INIT('h80)
	) name20344 (
		\m0_data_i[11]_pad ,
		_w9205_,
		_w9206_,
		_w22245_
	);
	LUT3 #(
		.INIT('h2a)
	) name20345 (
		\m7_data_i[11]_pad ,
		_w9205_,
		_w9206_,
		_w22246_
	);
	LUT4 #(
		.INIT('h6e7f)
	) name20346 (
		_w9200_,
		_w9203_,
		_w22245_,
		_w22246_,
		_w22247_
	);
	LUT4 #(
		.INIT('h7fff)
	) name20347 (
		_w22238_,
		_w22241_,
		_w22244_,
		_w22247_,
		_w22248_
	);
	LUT3 #(
		.INIT('h2a)
	) name20348 (
		\m3_data_i[12]_pad ,
		_w9205_,
		_w9206_,
		_w22249_
	);
	LUT3 #(
		.INIT('h80)
	) name20349 (
		\m4_data_i[12]_pad ,
		_w9205_,
		_w9206_,
		_w22250_
	);
	LUT4 #(
		.INIT('h9dbf)
	) name20350 (
		_w9200_,
		_w9203_,
		_w22249_,
		_w22250_,
		_w22251_
	);
	LUT3 #(
		.INIT('h80)
	) name20351 (
		\m6_data_i[12]_pad ,
		_w9205_,
		_w9206_,
		_w22252_
	);
	LUT3 #(
		.INIT('h80)
	) name20352 (
		\m2_data_i[12]_pad ,
		_w9205_,
		_w9206_,
		_w22253_
	);
	LUT4 #(
		.INIT('habef)
	) name20353 (
		_w9200_,
		_w9203_,
		_w22252_,
		_w22253_,
		_w22254_
	);
	LUT3 #(
		.INIT('h2a)
	) name20354 (
		\m5_data_i[12]_pad ,
		_w9205_,
		_w9206_,
		_w22255_
	);
	LUT3 #(
		.INIT('h2a)
	) name20355 (
		\m1_data_i[12]_pad ,
		_w9205_,
		_w9206_,
		_w22256_
	);
	LUT4 #(
		.INIT('h57df)
	) name20356 (
		_w9200_,
		_w9203_,
		_w22255_,
		_w22256_,
		_w22257_
	);
	LUT3 #(
		.INIT('h80)
	) name20357 (
		\m0_data_i[12]_pad ,
		_w9205_,
		_w9206_,
		_w22258_
	);
	LUT3 #(
		.INIT('h2a)
	) name20358 (
		\m7_data_i[12]_pad ,
		_w9205_,
		_w9206_,
		_w22259_
	);
	LUT4 #(
		.INIT('h6e7f)
	) name20359 (
		_w9200_,
		_w9203_,
		_w22258_,
		_w22259_,
		_w22260_
	);
	LUT4 #(
		.INIT('h7fff)
	) name20360 (
		_w22251_,
		_w22254_,
		_w22257_,
		_w22260_,
		_w22261_
	);
	LUT3 #(
		.INIT('h2a)
	) name20361 (
		\m3_data_i[13]_pad ,
		_w9205_,
		_w9206_,
		_w22262_
	);
	LUT3 #(
		.INIT('h80)
	) name20362 (
		\m4_data_i[13]_pad ,
		_w9205_,
		_w9206_,
		_w22263_
	);
	LUT4 #(
		.INIT('h9dbf)
	) name20363 (
		_w9200_,
		_w9203_,
		_w22262_,
		_w22263_,
		_w22264_
	);
	LUT3 #(
		.INIT('h80)
	) name20364 (
		\m6_data_i[13]_pad ,
		_w9205_,
		_w9206_,
		_w22265_
	);
	LUT3 #(
		.INIT('h80)
	) name20365 (
		\m2_data_i[13]_pad ,
		_w9205_,
		_w9206_,
		_w22266_
	);
	LUT4 #(
		.INIT('habef)
	) name20366 (
		_w9200_,
		_w9203_,
		_w22265_,
		_w22266_,
		_w22267_
	);
	LUT3 #(
		.INIT('h2a)
	) name20367 (
		\m5_data_i[13]_pad ,
		_w9205_,
		_w9206_,
		_w22268_
	);
	LUT3 #(
		.INIT('h2a)
	) name20368 (
		\m1_data_i[13]_pad ,
		_w9205_,
		_w9206_,
		_w22269_
	);
	LUT4 #(
		.INIT('h57df)
	) name20369 (
		_w9200_,
		_w9203_,
		_w22268_,
		_w22269_,
		_w22270_
	);
	LUT3 #(
		.INIT('h80)
	) name20370 (
		\m0_data_i[13]_pad ,
		_w9205_,
		_w9206_,
		_w22271_
	);
	LUT3 #(
		.INIT('h2a)
	) name20371 (
		\m7_data_i[13]_pad ,
		_w9205_,
		_w9206_,
		_w22272_
	);
	LUT4 #(
		.INIT('h6e7f)
	) name20372 (
		_w9200_,
		_w9203_,
		_w22271_,
		_w22272_,
		_w22273_
	);
	LUT4 #(
		.INIT('h7fff)
	) name20373 (
		_w22264_,
		_w22267_,
		_w22270_,
		_w22273_,
		_w22274_
	);
	LUT3 #(
		.INIT('h2a)
	) name20374 (
		\m3_data_i[14]_pad ,
		_w9205_,
		_w9206_,
		_w22275_
	);
	LUT3 #(
		.INIT('h80)
	) name20375 (
		\m4_data_i[14]_pad ,
		_w9205_,
		_w9206_,
		_w22276_
	);
	LUT4 #(
		.INIT('h9dbf)
	) name20376 (
		_w9200_,
		_w9203_,
		_w22275_,
		_w22276_,
		_w22277_
	);
	LUT3 #(
		.INIT('h80)
	) name20377 (
		\m6_data_i[14]_pad ,
		_w9205_,
		_w9206_,
		_w22278_
	);
	LUT3 #(
		.INIT('h80)
	) name20378 (
		\m2_data_i[14]_pad ,
		_w9205_,
		_w9206_,
		_w22279_
	);
	LUT4 #(
		.INIT('habef)
	) name20379 (
		_w9200_,
		_w9203_,
		_w22278_,
		_w22279_,
		_w22280_
	);
	LUT3 #(
		.INIT('h2a)
	) name20380 (
		\m5_data_i[14]_pad ,
		_w9205_,
		_w9206_,
		_w22281_
	);
	LUT3 #(
		.INIT('h2a)
	) name20381 (
		\m1_data_i[14]_pad ,
		_w9205_,
		_w9206_,
		_w22282_
	);
	LUT4 #(
		.INIT('h57df)
	) name20382 (
		_w9200_,
		_w9203_,
		_w22281_,
		_w22282_,
		_w22283_
	);
	LUT3 #(
		.INIT('h80)
	) name20383 (
		\m0_data_i[14]_pad ,
		_w9205_,
		_w9206_,
		_w22284_
	);
	LUT3 #(
		.INIT('h2a)
	) name20384 (
		\m7_data_i[14]_pad ,
		_w9205_,
		_w9206_,
		_w22285_
	);
	LUT4 #(
		.INIT('h6e7f)
	) name20385 (
		_w9200_,
		_w9203_,
		_w22284_,
		_w22285_,
		_w22286_
	);
	LUT4 #(
		.INIT('h7fff)
	) name20386 (
		_w22277_,
		_w22280_,
		_w22283_,
		_w22286_,
		_w22287_
	);
	LUT3 #(
		.INIT('h2a)
	) name20387 (
		\m3_data_i[15]_pad ,
		_w9205_,
		_w9206_,
		_w22288_
	);
	LUT3 #(
		.INIT('h80)
	) name20388 (
		\m4_data_i[15]_pad ,
		_w9205_,
		_w9206_,
		_w22289_
	);
	LUT4 #(
		.INIT('h9dbf)
	) name20389 (
		_w9200_,
		_w9203_,
		_w22288_,
		_w22289_,
		_w22290_
	);
	LUT3 #(
		.INIT('h80)
	) name20390 (
		\m6_data_i[15]_pad ,
		_w9205_,
		_w9206_,
		_w22291_
	);
	LUT3 #(
		.INIT('h80)
	) name20391 (
		\m2_data_i[15]_pad ,
		_w9205_,
		_w9206_,
		_w22292_
	);
	LUT4 #(
		.INIT('habef)
	) name20392 (
		_w9200_,
		_w9203_,
		_w22291_,
		_w22292_,
		_w22293_
	);
	LUT3 #(
		.INIT('h2a)
	) name20393 (
		\m5_data_i[15]_pad ,
		_w9205_,
		_w9206_,
		_w22294_
	);
	LUT3 #(
		.INIT('h2a)
	) name20394 (
		\m1_data_i[15]_pad ,
		_w9205_,
		_w9206_,
		_w22295_
	);
	LUT4 #(
		.INIT('h57df)
	) name20395 (
		_w9200_,
		_w9203_,
		_w22294_,
		_w22295_,
		_w22296_
	);
	LUT3 #(
		.INIT('h80)
	) name20396 (
		\m0_data_i[15]_pad ,
		_w9205_,
		_w9206_,
		_w22297_
	);
	LUT3 #(
		.INIT('h2a)
	) name20397 (
		\m7_data_i[15]_pad ,
		_w9205_,
		_w9206_,
		_w22298_
	);
	LUT4 #(
		.INIT('h6e7f)
	) name20398 (
		_w9200_,
		_w9203_,
		_w22297_,
		_w22298_,
		_w22299_
	);
	LUT4 #(
		.INIT('h7fff)
	) name20399 (
		_w22290_,
		_w22293_,
		_w22296_,
		_w22299_,
		_w22300_
	);
	LUT3 #(
		.INIT('h2a)
	) name20400 (
		\m3_data_i[16]_pad ,
		_w9205_,
		_w9206_,
		_w22301_
	);
	LUT3 #(
		.INIT('h80)
	) name20401 (
		\m4_data_i[16]_pad ,
		_w9205_,
		_w9206_,
		_w22302_
	);
	LUT4 #(
		.INIT('h9dbf)
	) name20402 (
		_w9200_,
		_w9203_,
		_w22301_,
		_w22302_,
		_w22303_
	);
	LUT3 #(
		.INIT('h80)
	) name20403 (
		\m6_data_i[16]_pad ,
		_w9205_,
		_w9206_,
		_w22304_
	);
	LUT3 #(
		.INIT('h80)
	) name20404 (
		\m2_data_i[16]_pad ,
		_w9205_,
		_w9206_,
		_w22305_
	);
	LUT4 #(
		.INIT('habef)
	) name20405 (
		_w9200_,
		_w9203_,
		_w22304_,
		_w22305_,
		_w22306_
	);
	LUT3 #(
		.INIT('h2a)
	) name20406 (
		\m5_data_i[16]_pad ,
		_w9205_,
		_w9206_,
		_w22307_
	);
	LUT3 #(
		.INIT('h2a)
	) name20407 (
		\m1_data_i[16]_pad ,
		_w9205_,
		_w9206_,
		_w22308_
	);
	LUT4 #(
		.INIT('h57df)
	) name20408 (
		_w9200_,
		_w9203_,
		_w22307_,
		_w22308_,
		_w22309_
	);
	LUT3 #(
		.INIT('h80)
	) name20409 (
		\m0_data_i[16]_pad ,
		_w9205_,
		_w9206_,
		_w22310_
	);
	LUT3 #(
		.INIT('h2a)
	) name20410 (
		\m7_data_i[16]_pad ,
		_w9205_,
		_w9206_,
		_w22311_
	);
	LUT4 #(
		.INIT('h6e7f)
	) name20411 (
		_w9200_,
		_w9203_,
		_w22310_,
		_w22311_,
		_w22312_
	);
	LUT4 #(
		.INIT('h7fff)
	) name20412 (
		_w22303_,
		_w22306_,
		_w22309_,
		_w22312_,
		_w22313_
	);
	LUT3 #(
		.INIT('h2a)
	) name20413 (
		\m3_data_i[17]_pad ,
		_w9205_,
		_w9206_,
		_w22314_
	);
	LUT3 #(
		.INIT('h80)
	) name20414 (
		\m4_data_i[17]_pad ,
		_w9205_,
		_w9206_,
		_w22315_
	);
	LUT4 #(
		.INIT('h9dbf)
	) name20415 (
		_w9200_,
		_w9203_,
		_w22314_,
		_w22315_,
		_w22316_
	);
	LUT3 #(
		.INIT('h80)
	) name20416 (
		\m6_data_i[17]_pad ,
		_w9205_,
		_w9206_,
		_w22317_
	);
	LUT3 #(
		.INIT('h80)
	) name20417 (
		\m2_data_i[17]_pad ,
		_w9205_,
		_w9206_,
		_w22318_
	);
	LUT4 #(
		.INIT('habef)
	) name20418 (
		_w9200_,
		_w9203_,
		_w22317_,
		_w22318_,
		_w22319_
	);
	LUT3 #(
		.INIT('h2a)
	) name20419 (
		\m5_data_i[17]_pad ,
		_w9205_,
		_w9206_,
		_w22320_
	);
	LUT3 #(
		.INIT('h2a)
	) name20420 (
		\m1_data_i[17]_pad ,
		_w9205_,
		_w9206_,
		_w22321_
	);
	LUT4 #(
		.INIT('h57df)
	) name20421 (
		_w9200_,
		_w9203_,
		_w22320_,
		_w22321_,
		_w22322_
	);
	LUT3 #(
		.INIT('h80)
	) name20422 (
		\m0_data_i[17]_pad ,
		_w9205_,
		_w9206_,
		_w22323_
	);
	LUT3 #(
		.INIT('h2a)
	) name20423 (
		\m7_data_i[17]_pad ,
		_w9205_,
		_w9206_,
		_w22324_
	);
	LUT4 #(
		.INIT('h6e7f)
	) name20424 (
		_w9200_,
		_w9203_,
		_w22323_,
		_w22324_,
		_w22325_
	);
	LUT4 #(
		.INIT('h7fff)
	) name20425 (
		_w22316_,
		_w22319_,
		_w22322_,
		_w22325_,
		_w22326_
	);
	LUT3 #(
		.INIT('h2a)
	) name20426 (
		\m3_data_i[18]_pad ,
		_w9205_,
		_w9206_,
		_w22327_
	);
	LUT3 #(
		.INIT('h80)
	) name20427 (
		\m4_data_i[18]_pad ,
		_w9205_,
		_w9206_,
		_w22328_
	);
	LUT4 #(
		.INIT('h9dbf)
	) name20428 (
		_w9200_,
		_w9203_,
		_w22327_,
		_w22328_,
		_w22329_
	);
	LUT3 #(
		.INIT('h80)
	) name20429 (
		\m6_data_i[18]_pad ,
		_w9205_,
		_w9206_,
		_w22330_
	);
	LUT3 #(
		.INIT('h80)
	) name20430 (
		\m2_data_i[18]_pad ,
		_w9205_,
		_w9206_,
		_w22331_
	);
	LUT4 #(
		.INIT('habef)
	) name20431 (
		_w9200_,
		_w9203_,
		_w22330_,
		_w22331_,
		_w22332_
	);
	LUT3 #(
		.INIT('h2a)
	) name20432 (
		\m5_data_i[18]_pad ,
		_w9205_,
		_w9206_,
		_w22333_
	);
	LUT3 #(
		.INIT('h2a)
	) name20433 (
		\m1_data_i[18]_pad ,
		_w9205_,
		_w9206_,
		_w22334_
	);
	LUT4 #(
		.INIT('h57df)
	) name20434 (
		_w9200_,
		_w9203_,
		_w22333_,
		_w22334_,
		_w22335_
	);
	LUT3 #(
		.INIT('h80)
	) name20435 (
		\m0_data_i[18]_pad ,
		_w9205_,
		_w9206_,
		_w22336_
	);
	LUT3 #(
		.INIT('h2a)
	) name20436 (
		\m7_data_i[18]_pad ,
		_w9205_,
		_w9206_,
		_w22337_
	);
	LUT4 #(
		.INIT('h6e7f)
	) name20437 (
		_w9200_,
		_w9203_,
		_w22336_,
		_w22337_,
		_w22338_
	);
	LUT4 #(
		.INIT('h7fff)
	) name20438 (
		_w22329_,
		_w22332_,
		_w22335_,
		_w22338_,
		_w22339_
	);
	LUT3 #(
		.INIT('h2a)
	) name20439 (
		\m3_data_i[19]_pad ,
		_w9205_,
		_w9206_,
		_w22340_
	);
	LUT3 #(
		.INIT('h80)
	) name20440 (
		\m4_data_i[19]_pad ,
		_w9205_,
		_w9206_,
		_w22341_
	);
	LUT4 #(
		.INIT('h9dbf)
	) name20441 (
		_w9200_,
		_w9203_,
		_w22340_,
		_w22341_,
		_w22342_
	);
	LUT3 #(
		.INIT('h80)
	) name20442 (
		\m6_data_i[19]_pad ,
		_w9205_,
		_w9206_,
		_w22343_
	);
	LUT3 #(
		.INIT('h80)
	) name20443 (
		\m2_data_i[19]_pad ,
		_w9205_,
		_w9206_,
		_w22344_
	);
	LUT4 #(
		.INIT('habef)
	) name20444 (
		_w9200_,
		_w9203_,
		_w22343_,
		_w22344_,
		_w22345_
	);
	LUT3 #(
		.INIT('h2a)
	) name20445 (
		\m5_data_i[19]_pad ,
		_w9205_,
		_w9206_,
		_w22346_
	);
	LUT3 #(
		.INIT('h2a)
	) name20446 (
		\m1_data_i[19]_pad ,
		_w9205_,
		_w9206_,
		_w22347_
	);
	LUT4 #(
		.INIT('h57df)
	) name20447 (
		_w9200_,
		_w9203_,
		_w22346_,
		_w22347_,
		_w22348_
	);
	LUT3 #(
		.INIT('h80)
	) name20448 (
		\m0_data_i[19]_pad ,
		_w9205_,
		_w9206_,
		_w22349_
	);
	LUT3 #(
		.INIT('h2a)
	) name20449 (
		\m7_data_i[19]_pad ,
		_w9205_,
		_w9206_,
		_w22350_
	);
	LUT4 #(
		.INIT('h6e7f)
	) name20450 (
		_w9200_,
		_w9203_,
		_w22349_,
		_w22350_,
		_w22351_
	);
	LUT4 #(
		.INIT('h7fff)
	) name20451 (
		_w22342_,
		_w22345_,
		_w22348_,
		_w22351_,
		_w22352_
	);
	LUT3 #(
		.INIT('h2a)
	) name20452 (
		\m3_data_i[1]_pad ,
		_w9205_,
		_w9206_,
		_w22353_
	);
	LUT3 #(
		.INIT('h80)
	) name20453 (
		\m4_data_i[1]_pad ,
		_w9205_,
		_w9206_,
		_w22354_
	);
	LUT4 #(
		.INIT('h9dbf)
	) name20454 (
		_w9200_,
		_w9203_,
		_w22353_,
		_w22354_,
		_w22355_
	);
	LUT3 #(
		.INIT('h80)
	) name20455 (
		\m6_data_i[1]_pad ,
		_w9205_,
		_w9206_,
		_w22356_
	);
	LUT3 #(
		.INIT('h80)
	) name20456 (
		\m2_data_i[1]_pad ,
		_w9205_,
		_w9206_,
		_w22357_
	);
	LUT4 #(
		.INIT('habef)
	) name20457 (
		_w9200_,
		_w9203_,
		_w22356_,
		_w22357_,
		_w22358_
	);
	LUT3 #(
		.INIT('h2a)
	) name20458 (
		\m5_data_i[1]_pad ,
		_w9205_,
		_w9206_,
		_w22359_
	);
	LUT3 #(
		.INIT('h2a)
	) name20459 (
		\m1_data_i[1]_pad ,
		_w9205_,
		_w9206_,
		_w22360_
	);
	LUT4 #(
		.INIT('h57df)
	) name20460 (
		_w9200_,
		_w9203_,
		_w22359_,
		_w22360_,
		_w22361_
	);
	LUT3 #(
		.INIT('h80)
	) name20461 (
		\m0_data_i[1]_pad ,
		_w9205_,
		_w9206_,
		_w22362_
	);
	LUT3 #(
		.INIT('h2a)
	) name20462 (
		\m7_data_i[1]_pad ,
		_w9205_,
		_w9206_,
		_w22363_
	);
	LUT4 #(
		.INIT('h6e7f)
	) name20463 (
		_w9200_,
		_w9203_,
		_w22362_,
		_w22363_,
		_w22364_
	);
	LUT4 #(
		.INIT('h7fff)
	) name20464 (
		_w22355_,
		_w22358_,
		_w22361_,
		_w22364_,
		_w22365_
	);
	LUT3 #(
		.INIT('h2a)
	) name20465 (
		\m3_data_i[20]_pad ,
		_w9205_,
		_w9206_,
		_w22366_
	);
	LUT3 #(
		.INIT('h80)
	) name20466 (
		\m4_data_i[20]_pad ,
		_w9205_,
		_w9206_,
		_w22367_
	);
	LUT4 #(
		.INIT('h9dbf)
	) name20467 (
		_w9200_,
		_w9203_,
		_w22366_,
		_w22367_,
		_w22368_
	);
	LUT3 #(
		.INIT('h80)
	) name20468 (
		\m6_data_i[20]_pad ,
		_w9205_,
		_w9206_,
		_w22369_
	);
	LUT3 #(
		.INIT('h80)
	) name20469 (
		\m2_data_i[20]_pad ,
		_w9205_,
		_w9206_,
		_w22370_
	);
	LUT4 #(
		.INIT('habef)
	) name20470 (
		_w9200_,
		_w9203_,
		_w22369_,
		_w22370_,
		_w22371_
	);
	LUT3 #(
		.INIT('h2a)
	) name20471 (
		\m5_data_i[20]_pad ,
		_w9205_,
		_w9206_,
		_w22372_
	);
	LUT3 #(
		.INIT('h2a)
	) name20472 (
		\m1_data_i[20]_pad ,
		_w9205_,
		_w9206_,
		_w22373_
	);
	LUT4 #(
		.INIT('h57df)
	) name20473 (
		_w9200_,
		_w9203_,
		_w22372_,
		_w22373_,
		_w22374_
	);
	LUT3 #(
		.INIT('h80)
	) name20474 (
		\m0_data_i[20]_pad ,
		_w9205_,
		_w9206_,
		_w22375_
	);
	LUT3 #(
		.INIT('h2a)
	) name20475 (
		\m7_data_i[20]_pad ,
		_w9205_,
		_w9206_,
		_w22376_
	);
	LUT4 #(
		.INIT('h6e7f)
	) name20476 (
		_w9200_,
		_w9203_,
		_w22375_,
		_w22376_,
		_w22377_
	);
	LUT4 #(
		.INIT('h7fff)
	) name20477 (
		_w22368_,
		_w22371_,
		_w22374_,
		_w22377_,
		_w22378_
	);
	LUT3 #(
		.INIT('h2a)
	) name20478 (
		\m3_data_i[21]_pad ,
		_w9205_,
		_w9206_,
		_w22379_
	);
	LUT3 #(
		.INIT('h80)
	) name20479 (
		\m4_data_i[21]_pad ,
		_w9205_,
		_w9206_,
		_w22380_
	);
	LUT4 #(
		.INIT('h9dbf)
	) name20480 (
		_w9200_,
		_w9203_,
		_w22379_,
		_w22380_,
		_w22381_
	);
	LUT3 #(
		.INIT('h80)
	) name20481 (
		\m6_data_i[21]_pad ,
		_w9205_,
		_w9206_,
		_w22382_
	);
	LUT3 #(
		.INIT('h80)
	) name20482 (
		\m2_data_i[21]_pad ,
		_w9205_,
		_w9206_,
		_w22383_
	);
	LUT4 #(
		.INIT('habef)
	) name20483 (
		_w9200_,
		_w9203_,
		_w22382_,
		_w22383_,
		_w22384_
	);
	LUT3 #(
		.INIT('h2a)
	) name20484 (
		\m5_data_i[21]_pad ,
		_w9205_,
		_w9206_,
		_w22385_
	);
	LUT3 #(
		.INIT('h2a)
	) name20485 (
		\m1_data_i[21]_pad ,
		_w9205_,
		_w9206_,
		_w22386_
	);
	LUT4 #(
		.INIT('h57df)
	) name20486 (
		_w9200_,
		_w9203_,
		_w22385_,
		_w22386_,
		_w22387_
	);
	LUT3 #(
		.INIT('h80)
	) name20487 (
		\m0_data_i[21]_pad ,
		_w9205_,
		_w9206_,
		_w22388_
	);
	LUT3 #(
		.INIT('h2a)
	) name20488 (
		\m7_data_i[21]_pad ,
		_w9205_,
		_w9206_,
		_w22389_
	);
	LUT4 #(
		.INIT('h6e7f)
	) name20489 (
		_w9200_,
		_w9203_,
		_w22388_,
		_w22389_,
		_w22390_
	);
	LUT4 #(
		.INIT('h7fff)
	) name20490 (
		_w22381_,
		_w22384_,
		_w22387_,
		_w22390_,
		_w22391_
	);
	LUT3 #(
		.INIT('h2a)
	) name20491 (
		\m3_data_i[22]_pad ,
		_w9205_,
		_w9206_,
		_w22392_
	);
	LUT3 #(
		.INIT('h80)
	) name20492 (
		\m4_data_i[22]_pad ,
		_w9205_,
		_w9206_,
		_w22393_
	);
	LUT4 #(
		.INIT('h9dbf)
	) name20493 (
		_w9200_,
		_w9203_,
		_w22392_,
		_w22393_,
		_w22394_
	);
	LUT3 #(
		.INIT('h80)
	) name20494 (
		\m6_data_i[22]_pad ,
		_w9205_,
		_w9206_,
		_w22395_
	);
	LUT3 #(
		.INIT('h80)
	) name20495 (
		\m2_data_i[22]_pad ,
		_w9205_,
		_w9206_,
		_w22396_
	);
	LUT4 #(
		.INIT('habef)
	) name20496 (
		_w9200_,
		_w9203_,
		_w22395_,
		_w22396_,
		_w22397_
	);
	LUT3 #(
		.INIT('h2a)
	) name20497 (
		\m5_data_i[22]_pad ,
		_w9205_,
		_w9206_,
		_w22398_
	);
	LUT3 #(
		.INIT('h2a)
	) name20498 (
		\m1_data_i[22]_pad ,
		_w9205_,
		_w9206_,
		_w22399_
	);
	LUT4 #(
		.INIT('h57df)
	) name20499 (
		_w9200_,
		_w9203_,
		_w22398_,
		_w22399_,
		_w22400_
	);
	LUT3 #(
		.INIT('h80)
	) name20500 (
		\m0_data_i[22]_pad ,
		_w9205_,
		_w9206_,
		_w22401_
	);
	LUT3 #(
		.INIT('h2a)
	) name20501 (
		\m7_data_i[22]_pad ,
		_w9205_,
		_w9206_,
		_w22402_
	);
	LUT4 #(
		.INIT('h6e7f)
	) name20502 (
		_w9200_,
		_w9203_,
		_w22401_,
		_w22402_,
		_w22403_
	);
	LUT4 #(
		.INIT('h7fff)
	) name20503 (
		_w22394_,
		_w22397_,
		_w22400_,
		_w22403_,
		_w22404_
	);
	LUT3 #(
		.INIT('h2a)
	) name20504 (
		\m3_data_i[23]_pad ,
		_w9205_,
		_w9206_,
		_w22405_
	);
	LUT3 #(
		.INIT('h80)
	) name20505 (
		\m4_data_i[23]_pad ,
		_w9205_,
		_w9206_,
		_w22406_
	);
	LUT4 #(
		.INIT('h9dbf)
	) name20506 (
		_w9200_,
		_w9203_,
		_w22405_,
		_w22406_,
		_w22407_
	);
	LUT3 #(
		.INIT('h80)
	) name20507 (
		\m6_data_i[23]_pad ,
		_w9205_,
		_w9206_,
		_w22408_
	);
	LUT3 #(
		.INIT('h80)
	) name20508 (
		\m2_data_i[23]_pad ,
		_w9205_,
		_w9206_,
		_w22409_
	);
	LUT4 #(
		.INIT('habef)
	) name20509 (
		_w9200_,
		_w9203_,
		_w22408_,
		_w22409_,
		_w22410_
	);
	LUT3 #(
		.INIT('h2a)
	) name20510 (
		\m5_data_i[23]_pad ,
		_w9205_,
		_w9206_,
		_w22411_
	);
	LUT3 #(
		.INIT('h2a)
	) name20511 (
		\m1_data_i[23]_pad ,
		_w9205_,
		_w9206_,
		_w22412_
	);
	LUT4 #(
		.INIT('h57df)
	) name20512 (
		_w9200_,
		_w9203_,
		_w22411_,
		_w22412_,
		_w22413_
	);
	LUT3 #(
		.INIT('h80)
	) name20513 (
		\m0_data_i[23]_pad ,
		_w9205_,
		_w9206_,
		_w22414_
	);
	LUT3 #(
		.INIT('h2a)
	) name20514 (
		\m7_data_i[23]_pad ,
		_w9205_,
		_w9206_,
		_w22415_
	);
	LUT4 #(
		.INIT('h6e7f)
	) name20515 (
		_w9200_,
		_w9203_,
		_w22414_,
		_w22415_,
		_w22416_
	);
	LUT4 #(
		.INIT('h7fff)
	) name20516 (
		_w22407_,
		_w22410_,
		_w22413_,
		_w22416_,
		_w22417_
	);
	LUT3 #(
		.INIT('h2a)
	) name20517 (
		\m3_data_i[24]_pad ,
		_w9205_,
		_w9206_,
		_w22418_
	);
	LUT3 #(
		.INIT('h80)
	) name20518 (
		\m4_data_i[24]_pad ,
		_w9205_,
		_w9206_,
		_w22419_
	);
	LUT4 #(
		.INIT('h9dbf)
	) name20519 (
		_w9200_,
		_w9203_,
		_w22418_,
		_w22419_,
		_w22420_
	);
	LUT3 #(
		.INIT('h80)
	) name20520 (
		\m6_data_i[24]_pad ,
		_w9205_,
		_w9206_,
		_w22421_
	);
	LUT3 #(
		.INIT('h80)
	) name20521 (
		\m2_data_i[24]_pad ,
		_w9205_,
		_w9206_,
		_w22422_
	);
	LUT4 #(
		.INIT('habef)
	) name20522 (
		_w9200_,
		_w9203_,
		_w22421_,
		_w22422_,
		_w22423_
	);
	LUT3 #(
		.INIT('h2a)
	) name20523 (
		\m5_data_i[24]_pad ,
		_w9205_,
		_w9206_,
		_w22424_
	);
	LUT3 #(
		.INIT('h2a)
	) name20524 (
		\m1_data_i[24]_pad ,
		_w9205_,
		_w9206_,
		_w22425_
	);
	LUT4 #(
		.INIT('h57df)
	) name20525 (
		_w9200_,
		_w9203_,
		_w22424_,
		_w22425_,
		_w22426_
	);
	LUT3 #(
		.INIT('h80)
	) name20526 (
		\m0_data_i[24]_pad ,
		_w9205_,
		_w9206_,
		_w22427_
	);
	LUT3 #(
		.INIT('h2a)
	) name20527 (
		\m7_data_i[24]_pad ,
		_w9205_,
		_w9206_,
		_w22428_
	);
	LUT4 #(
		.INIT('h6e7f)
	) name20528 (
		_w9200_,
		_w9203_,
		_w22427_,
		_w22428_,
		_w22429_
	);
	LUT4 #(
		.INIT('h7fff)
	) name20529 (
		_w22420_,
		_w22423_,
		_w22426_,
		_w22429_,
		_w22430_
	);
	LUT3 #(
		.INIT('h2a)
	) name20530 (
		\m3_data_i[25]_pad ,
		_w9205_,
		_w9206_,
		_w22431_
	);
	LUT3 #(
		.INIT('h80)
	) name20531 (
		\m4_data_i[25]_pad ,
		_w9205_,
		_w9206_,
		_w22432_
	);
	LUT4 #(
		.INIT('h9dbf)
	) name20532 (
		_w9200_,
		_w9203_,
		_w22431_,
		_w22432_,
		_w22433_
	);
	LUT3 #(
		.INIT('h80)
	) name20533 (
		\m6_data_i[25]_pad ,
		_w9205_,
		_w9206_,
		_w22434_
	);
	LUT3 #(
		.INIT('h80)
	) name20534 (
		\m2_data_i[25]_pad ,
		_w9205_,
		_w9206_,
		_w22435_
	);
	LUT4 #(
		.INIT('habef)
	) name20535 (
		_w9200_,
		_w9203_,
		_w22434_,
		_w22435_,
		_w22436_
	);
	LUT3 #(
		.INIT('h2a)
	) name20536 (
		\m5_data_i[25]_pad ,
		_w9205_,
		_w9206_,
		_w22437_
	);
	LUT3 #(
		.INIT('h2a)
	) name20537 (
		\m1_data_i[25]_pad ,
		_w9205_,
		_w9206_,
		_w22438_
	);
	LUT4 #(
		.INIT('h57df)
	) name20538 (
		_w9200_,
		_w9203_,
		_w22437_,
		_w22438_,
		_w22439_
	);
	LUT3 #(
		.INIT('h80)
	) name20539 (
		\m0_data_i[25]_pad ,
		_w9205_,
		_w9206_,
		_w22440_
	);
	LUT3 #(
		.INIT('h2a)
	) name20540 (
		\m7_data_i[25]_pad ,
		_w9205_,
		_w9206_,
		_w22441_
	);
	LUT4 #(
		.INIT('h6e7f)
	) name20541 (
		_w9200_,
		_w9203_,
		_w22440_,
		_w22441_,
		_w22442_
	);
	LUT4 #(
		.INIT('h7fff)
	) name20542 (
		_w22433_,
		_w22436_,
		_w22439_,
		_w22442_,
		_w22443_
	);
	LUT3 #(
		.INIT('h2a)
	) name20543 (
		\m3_data_i[26]_pad ,
		_w9205_,
		_w9206_,
		_w22444_
	);
	LUT3 #(
		.INIT('h80)
	) name20544 (
		\m4_data_i[26]_pad ,
		_w9205_,
		_w9206_,
		_w22445_
	);
	LUT4 #(
		.INIT('h9dbf)
	) name20545 (
		_w9200_,
		_w9203_,
		_w22444_,
		_w22445_,
		_w22446_
	);
	LUT3 #(
		.INIT('h80)
	) name20546 (
		\m6_data_i[26]_pad ,
		_w9205_,
		_w9206_,
		_w22447_
	);
	LUT3 #(
		.INIT('h80)
	) name20547 (
		\m2_data_i[26]_pad ,
		_w9205_,
		_w9206_,
		_w22448_
	);
	LUT4 #(
		.INIT('habef)
	) name20548 (
		_w9200_,
		_w9203_,
		_w22447_,
		_w22448_,
		_w22449_
	);
	LUT3 #(
		.INIT('h2a)
	) name20549 (
		\m5_data_i[26]_pad ,
		_w9205_,
		_w9206_,
		_w22450_
	);
	LUT3 #(
		.INIT('h2a)
	) name20550 (
		\m1_data_i[26]_pad ,
		_w9205_,
		_w9206_,
		_w22451_
	);
	LUT4 #(
		.INIT('h57df)
	) name20551 (
		_w9200_,
		_w9203_,
		_w22450_,
		_w22451_,
		_w22452_
	);
	LUT3 #(
		.INIT('h80)
	) name20552 (
		\m0_data_i[26]_pad ,
		_w9205_,
		_w9206_,
		_w22453_
	);
	LUT3 #(
		.INIT('h2a)
	) name20553 (
		\m7_data_i[26]_pad ,
		_w9205_,
		_w9206_,
		_w22454_
	);
	LUT4 #(
		.INIT('h6e7f)
	) name20554 (
		_w9200_,
		_w9203_,
		_w22453_,
		_w22454_,
		_w22455_
	);
	LUT4 #(
		.INIT('h7fff)
	) name20555 (
		_w22446_,
		_w22449_,
		_w22452_,
		_w22455_,
		_w22456_
	);
	LUT3 #(
		.INIT('h2a)
	) name20556 (
		\m3_data_i[27]_pad ,
		_w9205_,
		_w9206_,
		_w22457_
	);
	LUT3 #(
		.INIT('h80)
	) name20557 (
		\m4_data_i[27]_pad ,
		_w9205_,
		_w9206_,
		_w22458_
	);
	LUT4 #(
		.INIT('h9dbf)
	) name20558 (
		_w9200_,
		_w9203_,
		_w22457_,
		_w22458_,
		_w22459_
	);
	LUT3 #(
		.INIT('h80)
	) name20559 (
		\m6_data_i[27]_pad ,
		_w9205_,
		_w9206_,
		_w22460_
	);
	LUT3 #(
		.INIT('h80)
	) name20560 (
		\m2_data_i[27]_pad ,
		_w9205_,
		_w9206_,
		_w22461_
	);
	LUT4 #(
		.INIT('habef)
	) name20561 (
		_w9200_,
		_w9203_,
		_w22460_,
		_w22461_,
		_w22462_
	);
	LUT3 #(
		.INIT('h2a)
	) name20562 (
		\m5_data_i[27]_pad ,
		_w9205_,
		_w9206_,
		_w22463_
	);
	LUT3 #(
		.INIT('h2a)
	) name20563 (
		\m1_data_i[27]_pad ,
		_w9205_,
		_w9206_,
		_w22464_
	);
	LUT4 #(
		.INIT('h57df)
	) name20564 (
		_w9200_,
		_w9203_,
		_w22463_,
		_w22464_,
		_w22465_
	);
	LUT3 #(
		.INIT('h80)
	) name20565 (
		\m0_data_i[27]_pad ,
		_w9205_,
		_w9206_,
		_w22466_
	);
	LUT3 #(
		.INIT('h2a)
	) name20566 (
		\m7_data_i[27]_pad ,
		_w9205_,
		_w9206_,
		_w22467_
	);
	LUT4 #(
		.INIT('h6e7f)
	) name20567 (
		_w9200_,
		_w9203_,
		_w22466_,
		_w22467_,
		_w22468_
	);
	LUT4 #(
		.INIT('h7fff)
	) name20568 (
		_w22459_,
		_w22462_,
		_w22465_,
		_w22468_,
		_w22469_
	);
	LUT3 #(
		.INIT('h2a)
	) name20569 (
		\m3_data_i[28]_pad ,
		_w9205_,
		_w9206_,
		_w22470_
	);
	LUT3 #(
		.INIT('h80)
	) name20570 (
		\m4_data_i[28]_pad ,
		_w9205_,
		_w9206_,
		_w22471_
	);
	LUT4 #(
		.INIT('h9dbf)
	) name20571 (
		_w9200_,
		_w9203_,
		_w22470_,
		_w22471_,
		_w22472_
	);
	LUT3 #(
		.INIT('h80)
	) name20572 (
		\m6_data_i[28]_pad ,
		_w9205_,
		_w9206_,
		_w22473_
	);
	LUT3 #(
		.INIT('h80)
	) name20573 (
		\m2_data_i[28]_pad ,
		_w9205_,
		_w9206_,
		_w22474_
	);
	LUT4 #(
		.INIT('habef)
	) name20574 (
		_w9200_,
		_w9203_,
		_w22473_,
		_w22474_,
		_w22475_
	);
	LUT3 #(
		.INIT('h2a)
	) name20575 (
		\m5_data_i[28]_pad ,
		_w9205_,
		_w9206_,
		_w22476_
	);
	LUT3 #(
		.INIT('h2a)
	) name20576 (
		\m1_data_i[28]_pad ,
		_w9205_,
		_w9206_,
		_w22477_
	);
	LUT4 #(
		.INIT('h57df)
	) name20577 (
		_w9200_,
		_w9203_,
		_w22476_,
		_w22477_,
		_w22478_
	);
	LUT3 #(
		.INIT('h80)
	) name20578 (
		\m0_data_i[28]_pad ,
		_w9205_,
		_w9206_,
		_w22479_
	);
	LUT3 #(
		.INIT('h2a)
	) name20579 (
		\m7_data_i[28]_pad ,
		_w9205_,
		_w9206_,
		_w22480_
	);
	LUT4 #(
		.INIT('h6e7f)
	) name20580 (
		_w9200_,
		_w9203_,
		_w22479_,
		_w22480_,
		_w22481_
	);
	LUT4 #(
		.INIT('h7fff)
	) name20581 (
		_w22472_,
		_w22475_,
		_w22478_,
		_w22481_,
		_w22482_
	);
	LUT3 #(
		.INIT('h2a)
	) name20582 (
		\m3_data_i[29]_pad ,
		_w9205_,
		_w9206_,
		_w22483_
	);
	LUT3 #(
		.INIT('h80)
	) name20583 (
		\m4_data_i[29]_pad ,
		_w9205_,
		_w9206_,
		_w22484_
	);
	LUT4 #(
		.INIT('h9dbf)
	) name20584 (
		_w9200_,
		_w9203_,
		_w22483_,
		_w22484_,
		_w22485_
	);
	LUT3 #(
		.INIT('h80)
	) name20585 (
		\m6_data_i[29]_pad ,
		_w9205_,
		_w9206_,
		_w22486_
	);
	LUT3 #(
		.INIT('h80)
	) name20586 (
		\m2_data_i[29]_pad ,
		_w9205_,
		_w9206_,
		_w22487_
	);
	LUT4 #(
		.INIT('habef)
	) name20587 (
		_w9200_,
		_w9203_,
		_w22486_,
		_w22487_,
		_w22488_
	);
	LUT3 #(
		.INIT('h2a)
	) name20588 (
		\m5_data_i[29]_pad ,
		_w9205_,
		_w9206_,
		_w22489_
	);
	LUT3 #(
		.INIT('h2a)
	) name20589 (
		\m1_data_i[29]_pad ,
		_w9205_,
		_w9206_,
		_w22490_
	);
	LUT4 #(
		.INIT('h57df)
	) name20590 (
		_w9200_,
		_w9203_,
		_w22489_,
		_w22490_,
		_w22491_
	);
	LUT3 #(
		.INIT('h80)
	) name20591 (
		\m0_data_i[29]_pad ,
		_w9205_,
		_w9206_,
		_w22492_
	);
	LUT3 #(
		.INIT('h2a)
	) name20592 (
		\m7_data_i[29]_pad ,
		_w9205_,
		_w9206_,
		_w22493_
	);
	LUT4 #(
		.INIT('h6e7f)
	) name20593 (
		_w9200_,
		_w9203_,
		_w22492_,
		_w22493_,
		_w22494_
	);
	LUT4 #(
		.INIT('h7fff)
	) name20594 (
		_w22485_,
		_w22488_,
		_w22491_,
		_w22494_,
		_w22495_
	);
	LUT3 #(
		.INIT('h2a)
	) name20595 (
		\m3_data_i[2]_pad ,
		_w9205_,
		_w9206_,
		_w22496_
	);
	LUT3 #(
		.INIT('h80)
	) name20596 (
		\m4_data_i[2]_pad ,
		_w9205_,
		_w9206_,
		_w22497_
	);
	LUT4 #(
		.INIT('h9dbf)
	) name20597 (
		_w9200_,
		_w9203_,
		_w22496_,
		_w22497_,
		_w22498_
	);
	LUT3 #(
		.INIT('h80)
	) name20598 (
		\m6_data_i[2]_pad ,
		_w9205_,
		_w9206_,
		_w22499_
	);
	LUT3 #(
		.INIT('h80)
	) name20599 (
		\m2_data_i[2]_pad ,
		_w9205_,
		_w9206_,
		_w22500_
	);
	LUT4 #(
		.INIT('habef)
	) name20600 (
		_w9200_,
		_w9203_,
		_w22499_,
		_w22500_,
		_w22501_
	);
	LUT3 #(
		.INIT('h2a)
	) name20601 (
		\m5_data_i[2]_pad ,
		_w9205_,
		_w9206_,
		_w22502_
	);
	LUT3 #(
		.INIT('h2a)
	) name20602 (
		\m1_data_i[2]_pad ,
		_w9205_,
		_w9206_,
		_w22503_
	);
	LUT4 #(
		.INIT('h57df)
	) name20603 (
		_w9200_,
		_w9203_,
		_w22502_,
		_w22503_,
		_w22504_
	);
	LUT3 #(
		.INIT('h80)
	) name20604 (
		\m0_data_i[2]_pad ,
		_w9205_,
		_w9206_,
		_w22505_
	);
	LUT3 #(
		.INIT('h2a)
	) name20605 (
		\m7_data_i[2]_pad ,
		_w9205_,
		_w9206_,
		_w22506_
	);
	LUT4 #(
		.INIT('h6e7f)
	) name20606 (
		_w9200_,
		_w9203_,
		_w22505_,
		_w22506_,
		_w22507_
	);
	LUT4 #(
		.INIT('h7fff)
	) name20607 (
		_w22498_,
		_w22501_,
		_w22504_,
		_w22507_,
		_w22508_
	);
	LUT3 #(
		.INIT('h2a)
	) name20608 (
		\m3_data_i[30]_pad ,
		_w9205_,
		_w9206_,
		_w22509_
	);
	LUT3 #(
		.INIT('h80)
	) name20609 (
		\m4_data_i[30]_pad ,
		_w9205_,
		_w9206_,
		_w22510_
	);
	LUT4 #(
		.INIT('h9dbf)
	) name20610 (
		_w9200_,
		_w9203_,
		_w22509_,
		_w22510_,
		_w22511_
	);
	LUT3 #(
		.INIT('h80)
	) name20611 (
		\m6_data_i[30]_pad ,
		_w9205_,
		_w9206_,
		_w22512_
	);
	LUT3 #(
		.INIT('h80)
	) name20612 (
		\m2_data_i[30]_pad ,
		_w9205_,
		_w9206_,
		_w22513_
	);
	LUT4 #(
		.INIT('habef)
	) name20613 (
		_w9200_,
		_w9203_,
		_w22512_,
		_w22513_,
		_w22514_
	);
	LUT3 #(
		.INIT('h2a)
	) name20614 (
		\m5_data_i[30]_pad ,
		_w9205_,
		_w9206_,
		_w22515_
	);
	LUT3 #(
		.INIT('h2a)
	) name20615 (
		\m1_data_i[30]_pad ,
		_w9205_,
		_w9206_,
		_w22516_
	);
	LUT4 #(
		.INIT('h57df)
	) name20616 (
		_w9200_,
		_w9203_,
		_w22515_,
		_w22516_,
		_w22517_
	);
	LUT3 #(
		.INIT('h80)
	) name20617 (
		\m0_data_i[30]_pad ,
		_w9205_,
		_w9206_,
		_w22518_
	);
	LUT3 #(
		.INIT('h2a)
	) name20618 (
		\m7_data_i[30]_pad ,
		_w9205_,
		_w9206_,
		_w22519_
	);
	LUT4 #(
		.INIT('h6e7f)
	) name20619 (
		_w9200_,
		_w9203_,
		_w22518_,
		_w22519_,
		_w22520_
	);
	LUT4 #(
		.INIT('h7fff)
	) name20620 (
		_w22511_,
		_w22514_,
		_w22517_,
		_w22520_,
		_w22521_
	);
	LUT3 #(
		.INIT('h2a)
	) name20621 (
		\m3_data_i[31]_pad ,
		_w9205_,
		_w9206_,
		_w22522_
	);
	LUT3 #(
		.INIT('h80)
	) name20622 (
		\m4_data_i[31]_pad ,
		_w9205_,
		_w9206_,
		_w22523_
	);
	LUT4 #(
		.INIT('h9dbf)
	) name20623 (
		_w9200_,
		_w9203_,
		_w22522_,
		_w22523_,
		_w22524_
	);
	LUT3 #(
		.INIT('h80)
	) name20624 (
		\m6_data_i[31]_pad ,
		_w9205_,
		_w9206_,
		_w22525_
	);
	LUT3 #(
		.INIT('h80)
	) name20625 (
		\m2_data_i[31]_pad ,
		_w9205_,
		_w9206_,
		_w22526_
	);
	LUT4 #(
		.INIT('habef)
	) name20626 (
		_w9200_,
		_w9203_,
		_w22525_,
		_w22526_,
		_w22527_
	);
	LUT3 #(
		.INIT('h2a)
	) name20627 (
		\m5_data_i[31]_pad ,
		_w9205_,
		_w9206_,
		_w22528_
	);
	LUT3 #(
		.INIT('h2a)
	) name20628 (
		\m1_data_i[31]_pad ,
		_w9205_,
		_w9206_,
		_w22529_
	);
	LUT4 #(
		.INIT('h57df)
	) name20629 (
		_w9200_,
		_w9203_,
		_w22528_,
		_w22529_,
		_w22530_
	);
	LUT3 #(
		.INIT('h80)
	) name20630 (
		\m0_data_i[31]_pad ,
		_w9205_,
		_w9206_,
		_w22531_
	);
	LUT3 #(
		.INIT('h2a)
	) name20631 (
		\m7_data_i[31]_pad ,
		_w9205_,
		_w9206_,
		_w22532_
	);
	LUT4 #(
		.INIT('h6e7f)
	) name20632 (
		_w9200_,
		_w9203_,
		_w22531_,
		_w22532_,
		_w22533_
	);
	LUT4 #(
		.INIT('h7fff)
	) name20633 (
		_w22524_,
		_w22527_,
		_w22530_,
		_w22533_,
		_w22534_
	);
	LUT3 #(
		.INIT('h2a)
	) name20634 (
		\m3_data_i[3]_pad ,
		_w9205_,
		_w9206_,
		_w22535_
	);
	LUT3 #(
		.INIT('h80)
	) name20635 (
		\m4_data_i[3]_pad ,
		_w9205_,
		_w9206_,
		_w22536_
	);
	LUT4 #(
		.INIT('h9dbf)
	) name20636 (
		_w9200_,
		_w9203_,
		_w22535_,
		_w22536_,
		_w22537_
	);
	LUT3 #(
		.INIT('h80)
	) name20637 (
		\m6_data_i[3]_pad ,
		_w9205_,
		_w9206_,
		_w22538_
	);
	LUT3 #(
		.INIT('h80)
	) name20638 (
		\m2_data_i[3]_pad ,
		_w9205_,
		_w9206_,
		_w22539_
	);
	LUT4 #(
		.INIT('habef)
	) name20639 (
		_w9200_,
		_w9203_,
		_w22538_,
		_w22539_,
		_w22540_
	);
	LUT3 #(
		.INIT('h2a)
	) name20640 (
		\m5_data_i[3]_pad ,
		_w9205_,
		_w9206_,
		_w22541_
	);
	LUT3 #(
		.INIT('h2a)
	) name20641 (
		\m1_data_i[3]_pad ,
		_w9205_,
		_w9206_,
		_w22542_
	);
	LUT4 #(
		.INIT('h57df)
	) name20642 (
		_w9200_,
		_w9203_,
		_w22541_,
		_w22542_,
		_w22543_
	);
	LUT3 #(
		.INIT('h80)
	) name20643 (
		\m0_data_i[3]_pad ,
		_w9205_,
		_w9206_,
		_w22544_
	);
	LUT3 #(
		.INIT('h2a)
	) name20644 (
		\m7_data_i[3]_pad ,
		_w9205_,
		_w9206_,
		_w22545_
	);
	LUT4 #(
		.INIT('h6e7f)
	) name20645 (
		_w9200_,
		_w9203_,
		_w22544_,
		_w22545_,
		_w22546_
	);
	LUT4 #(
		.INIT('h7fff)
	) name20646 (
		_w22537_,
		_w22540_,
		_w22543_,
		_w22546_,
		_w22547_
	);
	LUT3 #(
		.INIT('h2a)
	) name20647 (
		\m3_data_i[4]_pad ,
		_w9205_,
		_w9206_,
		_w22548_
	);
	LUT3 #(
		.INIT('h80)
	) name20648 (
		\m4_data_i[4]_pad ,
		_w9205_,
		_w9206_,
		_w22549_
	);
	LUT4 #(
		.INIT('h9dbf)
	) name20649 (
		_w9200_,
		_w9203_,
		_w22548_,
		_w22549_,
		_w22550_
	);
	LUT3 #(
		.INIT('h80)
	) name20650 (
		\m6_data_i[4]_pad ,
		_w9205_,
		_w9206_,
		_w22551_
	);
	LUT3 #(
		.INIT('h80)
	) name20651 (
		\m2_data_i[4]_pad ,
		_w9205_,
		_w9206_,
		_w22552_
	);
	LUT4 #(
		.INIT('habef)
	) name20652 (
		_w9200_,
		_w9203_,
		_w22551_,
		_w22552_,
		_w22553_
	);
	LUT3 #(
		.INIT('h2a)
	) name20653 (
		\m5_data_i[4]_pad ,
		_w9205_,
		_w9206_,
		_w22554_
	);
	LUT3 #(
		.INIT('h2a)
	) name20654 (
		\m1_data_i[4]_pad ,
		_w9205_,
		_w9206_,
		_w22555_
	);
	LUT4 #(
		.INIT('h57df)
	) name20655 (
		_w9200_,
		_w9203_,
		_w22554_,
		_w22555_,
		_w22556_
	);
	LUT3 #(
		.INIT('h80)
	) name20656 (
		\m0_data_i[4]_pad ,
		_w9205_,
		_w9206_,
		_w22557_
	);
	LUT3 #(
		.INIT('h2a)
	) name20657 (
		\m7_data_i[4]_pad ,
		_w9205_,
		_w9206_,
		_w22558_
	);
	LUT4 #(
		.INIT('h6e7f)
	) name20658 (
		_w9200_,
		_w9203_,
		_w22557_,
		_w22558_,
		_w22559_
	);
	LUT4 #(
		.INIT('h7fff)
	) name20659 (
		_w22550_,
		_w22553_,
		_w22556_,
		_w22559_,
		_w22560_
	);
	LUT3 #(
		.INIT('h2a)
	) name20660 (
		\m3_data_i[5]_pad ,
		_w9205_,
		_w9206_,
		_w22561_
	);
	LUT3 #(
		.INIT('h80)
	) name20661 (
		\m4_data_i[5]_pad ,
		_w9205_,
		_w9206_,
		_w22562_
	);
	LUT4 #(
		.INIT('h9dbf)
	) name20662 (
		_w9200_,
		_w9203_,
		_w22561_,
		_w22562_,
		_w22563_
	);
	LUT3 #(
		.INIT('h80)
	) name20663 (
		\m6_data_i[5]_pad ,
		_w9205_,
		_w9206_,
		_w22564_
	);
	LUT3 #(
		.INIT('h80)
	) name20664 (
		\m2_data_i[5]_pad ,
		_w9205_,
		_w9206_,
		_w22565_
	);
	LUT4 #(
		.INIT('habef)
	) name20665 (
		_w9200_,
		_w9203_,
		_w22564_,
		_w22565_,
		_w22566_
	);
	LUT3 #(
		.INIT('h2a)
	) name20666 (
		\m5_data_i[5]_pad ,
		_w9205_,
		_w9206_,
		_w22567_
	);
	LUT3 #(
		.INIT('h2a)
	) name20667 (
		\m1_data_i[5]_pad ,
		_w9205_,
		_w9206_,
		_w22568_
	);
	LUT4 #(
		.INIT('h57df)
	) name20668 (
		_w9200_,
		_w9203_,
		_w22567_,
		_w22568_,
		_w22569_
	);
	LUT3 #(
		.INIT('h80)
	) name20669 (
		\m0_data_i[5]_pad ,
		_w9205_,
		_w9206_,
		_w22570_
	);
	LUT3 #(
		.INIT('h2a)
	) name20670 (
		\m7_data_i[5]_pad ,
		_w9205_,
		_w9206_,
		_w22571_
	);
	LUT4 #(
		.INIT('h6e7f)
	) name20671 (
		_w9200_,
		_w9203_,
		_w22570_,
		_w22571_,
		_w22572_
	);
	LUT4 #(
		.INIT('h7fff)
	) name20672 (
		_w22563_,
		_w22566_,
		_w22569_,
		_w22572_,
		_w22573_
	);
	LUT3 #(
		.INIT('h2a)
	) name20673 (
		\m3_data_i[6]_pad ,
		_w9205_,
		_w9206_,
		_w22574_
	);
	LUT3 #(
		.INIT('h80)
	) name20674 (
		\m4_data_i[6]_pad ,
		_w9205_,
		_w9206_,
		_w22575_
	);
	LUT4 #(
		.INIT('h9dbf)
	) name20675 (
		_w9200_,
		_w9203_,
		_w22574_,
		_w22575_,
		_w22576_
	);
	LUT3 #(
		.INIT('h80)
	) name20676 (
		\m6_data_i[6]_pad ,
		_w9205_,
		_w9206_,
		_w22577_
	);
	LUT3 #(
		.INIT('h80)
	) name20677 (
		\m2_data_i[6]_pad ,
		_w9205_,
		_w9206_,
		_w22578_
	);
	LUT4 #(
		.INIT('habef)
	) name20678 (
		_w9200_,
		_w9203_,
		_w22577_,
		_w22578_,
		_w22579_
	);
	LUT3 #(
		.INIT('h2a)
	) name20679 (
		\m5_data_i[6]_pad ,
		_w9205_,
		_w9206_,
		_w22580_
	);
	LUT3 #(
		.INIT('h2a)
	) name20680 (
		\m1_data_i[6]_pad ,
		_w9205_,
		_w9206_,
		_w22581_
	);
	LUT4 #(
		.INIT('h57df)
	) name20681 (
		_w9200_,
		_w9203_,
		_w22580_,
		_w22581_,
		_w22582_
	);
	LUT3 #(
		.INIT('h80)
	) name20682 (
		\m0_data_i[6]_pad ,
		_w9205_,
		_w9206_,
		_w22583_
	);
	LUT3 #(
		.INIT('h2a)
	) name20683 (
		\m7_data_i[6]_pad ,
		_w9205_,
		_w9206_,
		_w22584_
	);
	LUT4 #(
		.INIT('h6e7f)
	) name20684 (
		_w9200_,
		_w9203_,
		_w22583_,
		_w22584_,
		_w22585_
	);
	LUT4 #(
		.INIT('h7fff)
	) name20685 (
		_w22576_,
		_w22579_,
		_w22582_,
		_w22585_,
		_w22586_
	);
	LUT3 #(
		.INIT('h2a)
	) name20686 (
		\m3_data_i[7]_pad ,
		_w9205_,
		_w9206_,
		_w22587_
	);
	LUT3 #(
		.INIT('h80)
	) name20687 (
		\m4_data_i[7]_pad ,
		_w9205_,
		_w9206_,
		_w22588_
	);
	LUT4 #(
		.INIT('h9dbf)
	) name20688 (
		_w9200_,
		_w9203_,
		_w22587_,
		_w22588_,
		_w22589_
	);
	LUT3 #(
		.INIT('h80)
	) name20689 (
		\m6_data_i[7]_pad ,
		_w9205_,
		_w9206_,
		_w22590_
	);
	LUT3 #(
		.INIT('h80)
	) name20690 (
		\m2_data_i[7]_pad ,
		_w9205_,
		_w9206_,
		_w22591_
	);
	LUT4 #(
		.INIT('habef)
	) name20691 (
		_w9200_,
		_w9203_,
		_w22590_,
		_w22591_,
		_w22592_
	);
	LUT3 #(
		.INIT('h2a)
	) name20692 (
		\m5_data_i[7]_pad ,
		_w9205_,
		_w9206_,
		_w22593_
	);
	LUT3 #(
		.INIT('h2a)
	) name20693 (
		\m1_data_i[7]_pad ,
		_w9205_,
		_w9206_,
		_w22594_
	);
	LUT4 #(
		.INIT('h57df)
	) name20694 (
		_w9200_,
		_w9203_,
		_w22593_,
		_w22594_,
		_w22595_
	);
	LUT3 #(
		.INIT('h80)
	) name20695 (
		\m0_data_i[7]_pad ,
		_w9205_,
		_w9206_,
		_w22596_
	);
	LUT3 #(
		.INIT('h2a)
	) name20696 (
		\m7_data_i[7]_pad ,
		_w9205_,
		_w9206_,
		_w22597_
	);
	LUT4 #(
		.INIT('h6e7f)
	) name20697 (
		_w9200_,
		_w9203_,
		_w22596_,
		_w22597_,
		_w22598_
	);
	LUT4 #(
		.INIT('h7fff)
	) name20698 (
		_w22589_,
		_w22592_,
		_w22595_,
		_w22598_,
		_w22599_
	);
	LUT3 #(
		.INIT('h2a)
	) name20699 (
		\m3_data_i[8]_pad ,
		_w9205_,
		_w9206_,
		_w22600_
	);
	LUT3 #(
		.INIT('h80)
	) name20700 (
		\m4_data_i[8]_pad ,
		_w9205_,
		_w9206_,
		_w22601_
	);
	LUT4 #(
		.INIT('h9dbf)
	) name20701 (
		_w9200_,
		_w9203_,
		_w22600_,
		_w22601_,
		_w22602_
	);
	LUT3 #(
		.INIT('h80)
	) name20702 (
		\m6_data_i[8]_pad ,
		_w9205_,
		_w9206_,
		_w22603_
	);
	LUT3 #(
		.INIT('h80)
	) name20703 (
		\m2_data_i[8]_pad ,
		_w9205_,
		_w9206_,
		_w22604_
	);
	LUT4 #(
		.INIT('habef)
	) name20704 (
		_w9200_,
		_w9203_,
		_w22603_,
		_w22604_,
		_w22605_
	);
	LUT3 #(
		.INIT('h2a)
	) name20705 (
		\m5_data_i[8]_pad ,
		_w9205_,
		_w9206_,
		_w22606_
	);
	LUT3 #(
		.INIT('h2a)
	) name20706 (
		\m1_data_i[8]_pad ,
		_w9205_,
		_w9206_,
		_w22607_
	);
	LUT4 #(
		.INIT('h57df)
	) name20707 (
		_w9200_,
		_w9203_,
		_w22606_,
		_w22607_,
		_w22608_
	);
	LUT3 #(
		.INIT('h80)
	) name20708 (
		\m0_data_i[8]_pad ,
		_w9205_,
		_w9206_,
		_w22609_
	);
	LUT3 #(
		.INIT('h2a)
	) name20709 (
		\m7_data_i[8]_pad ,
		_w9205_,
		_w9206_,
		_w22610_
	);
	LUT4 #(
		.INIT('h6e7f)
	) name20710 (
		_w9200_,
		_w9203_,
		_w22609_,
		_w22610_,
		_w22611_
	);
	LUT4 #(
		.INIT('h7fff)
	) name20711 (
		_w22602_,
		_w22605_,
		_w22608_,
		_w22611_,
		_w22612_
	);
	LUT3 #(
		.INIT('h2a)
	) name20712 (
		\m3_data_i[9]_pad ,
		_w9205_,
		_w9206_,
		_w22613_
	);
	LUT3 #(
		.INIT('h80)
	) name20713 (
		\m4_data_i[9]_pad ,
		_w9205_,
		_w9206_,
		_w22614_
	);
	LUT4 #(
		.INIT('h9dbf)
	) name20714 (
		_w9200_,
		_w9203_,
		_w22613_,
		_w22614_,
		_w22615_
	);
	LUT3 #(
		.INIT('h80)
	) name20715 (
		\m6_data_i[9]_pad ,
		_w9205_,
		_w9206_,
		_w22616_
	);
	LUT3 #(
		.INIT('h80)
	) name20716 (
		\m2_data_i[9]_pad ,
		_w9205_,
		_w9206_,
		_w22617_
	);
	LUT4 #(
		.INIT('habef)
	) name20717 (
		_w9200_,
		_w9203_,
		_w22616_,
		_w22617_,
		_w22618_
	);
	LUT3 #(
		.INIT('h2a)
	) name20718 (
		\m5_data_i[9]_pad ,
		_w9205_,
		_w9206_,
		_w22619_
	);
	LUT3 #(
		.INIT('h2a)
	) name20719 (
		\m1_data_i[9]_pad ,
		_w9205_,
		_w9206_,
		_w22620_
	);
	LUT4 #(
		.INIT('h57df)
	) name20720 (
		_w9200_,
		_w9203_,
		_w22619_,
		_w22620_,
		_w22621_
	);
	LUT3 #(
		.INIT('h80)
	) name20721 (
		\m0_data_i[9]_pad ,
		_w9205_,
		_w9206_,
		_w22622_
	);
	LUT3 #(
		.INIT('h2a)
	) name20722 (
		\m7_data_i[9]_pad ,
		_w9205_,
		_w9206_,
		_w22623_
	);
	LUT4 #(
		.INIT('h6e7f)
	) name20723 (
		_w9200_,
		_w9203_,
		_w22622_,
		_w22623_,
		_w22624_
	);
	LUT4 #(
		.INIT('h7fff)
	) name20724 (
		_w22615_,
		_w22618_,
		_w22621_,
		_w22624_,
		_w22625_
	);
	LUT3 #(
		.INIT('h2a)
	) name20725 (
		\m3_sel_i[0]_pad ,
		_w9205_,
		_w9206_,
		_w22626_
	);
	LUT3 #(
		.INIT('h80)
	) name20726 (
		\m4_sel_i[0]_pad ,
		_w9205_,
		_w9206_,
		_w22627_
	);
	LUT4 #(
		.INIT('h9dbf)
	) name20727 (
		_w9200_,
		_w9203_,
		_w22626_,
		_w22627_,
		_w22628_
	);
	LUT3 #(
		.INIT('h80)
	) name20728 (
		\m6_sel_i[0]_pad ,
		_w9205_,
		_w9206_,
		_w22629_
	);
	LUT3 #(
		.INIT('h80)
	) name20729 (
		\m2_sel_i[0]_pad ,
		_w9205_,
		_w9206_,
		_w22630_
	);
	LUT4 #(
		.INIT('habef)
	) name20730 (
		_w9200_,
		_w9203_,
		_w22629_,
		_w22630_,
		_w22631_
	);
	LUT3 #(
		.INIT('h2a)
	) name20731 (
		\m5_sel_i[0]_pad ,
		_w9205_,
		_w9206_,
		_w22632_
	);
	LUT3 #(
		.INIT('h2a)
	) name20732 (
		\m1_sel_i[0]_pad ,
		_w9205_,
		_w9206_,
		_w22633_
	);
	LUT4 #(
		.INIT('h57df)
	) name20733 (
		_w9200_,
		_w9203_,
		_w22632_,
		_w22633_,
		_w22634_
	);
	LUT3 #(
		.INIT('h80)
	) name20734 (
		\m0_sel_i[0]_pad ,
		_w9205_,
		_w9206_,
		_w22635_
	);
	LUT3 #(
		.INIT('h2a)
	) name20735 (
		\m7_sel_i[0]_pad ,
		_w9205_,
		_w9206_,
		_w22636_
	);
	LUT4 #(
		.INIT('h6e7f)
	) name20736 (
		_w9200_,
		_w9203_,
		_w22635_,
		_w22636_,
		_w22637_
	);
	LUT4 #(
		.INIT('h7fff)
	) name20737 (
		_w22628_,
		_w22631_,
		_w22634_,
		_w22637_,
		_w22638_
	);
	LUT3 #(
		.INIT('h2a)
	) name20738 (
		\m3_sel_i[1]_pad ,
		_w9205_,
		_w9206_,
		_w22639_
	);
	LUT3 #(
		.INIT('h80)
	) name20739 (
		\m4_sel_i[1]_pad ,
		_w9205_,
		_w9206_,
		_w22640_
	);
	LUT4 #(
		.INIT('h9dbf)
	) name20740 (
		_w9200_,
		_w9203_,
		_w22639_,
		_w22640_,
		_w22641_
	);
	LUT3 #(
		.INIT('h80)
	) name20741 (
		\m6_sel_i[1]_pad ,
		_w9205_,
		_w9206_,
		_w22642_
	);
	LUT3 #(
		.INIT('h80)
	) name20742 (
		\m2_sel_i[1]_pad ,
		_w9205_,
		_w9206_,
		_w22643_
	);
	LUT4 #(
		.INIT('habef)
	) name20743 (
		_w9200_,
		_w9203_,
		_w22642_,
		_w22643_,
		_w22644_
	);
	LUT3 #(
		.INIT('h2a)
	) name20744 (
		\m5_sel_i[1]_pad ,
		_w9205_,
		_w9206_,
		_w22645_
	);
	LUT3 #(
		.INIT('h2a)
	) name20745 (
		\m1_sel_i[1]_pad ,
		_w9205_,
		_w9206_,
		_w22646_
	);
	LUT4 #(
		.INIT('h57df)
	) name20746 (
		_w9200_,
		_w9203_,
		_w22645_,
		_w22646_,
		_w22647_
	);
	LUT3 #(
		.INIT('h80)
	) name20747 (
		\m0_sel_i[1]_pad ,
		_w9205_,
		_w9206_,
		_w22648_
	);
	LUT3 #(
		.INIT('h2a)
	) name20748 (
		\m7_sel_i[1]_pad ,
		_w9205_,
		_w9206_,
		_w22649_
	);
	LUT4 #(
		.INIT('h6e7f)
	) name20749 (
		_w9200_,
		_w9203_,
		_w22648_,
		_w22649_,
		_w22650_
	);
	LUT4 #(
		.INIT('h7fff)
	) name20750 (
		_w22641_,
		_w22644_,
		_w22647_,
		_w22650_,
		_w22651_
	);
	LUT3 #(
		.INIT('h2a)
	) name20751 (
		\m3_sel_i[2]_pad ,
		_w9205_,
		_w9206_,
		_w22652_
	);
	LUT3 #(
		.INIT('h80)
	) name20752 (
		\m4_sel_i[2]_pad ,
		_w9205_,
		_w9206_,
		_w22653_
	);
	LUT4 #(
		.INIT('h9dbf)
	) name20753 (
		_w9200_,
		_w9203_,
		_w22652_,
		_w22653_,
		_w22654_
	);
	LUT3 #(
		.INIT('h80)
	) name20754 (
		\m6_sel_i[2]_pad ,
		_w9205_,
		_w9206_,
		_w22655_
	);
	LUT3 #(
		.INIT('h80)
	) name20755 (
		\m2_sel_i[2]_pad ,
		_w9205_,
		_w9206_,
		_w22656_
	);
	LUT4 #(
		.INIT('habef)
	) name20756 (
		_w9200_,
		_w9203_,
		_w22655_,
		_w22656_,
		_w22657_
	);
	LUT3 #(
		.INIT('h2a)
	) name20757 (
		\m5_sel_i[2]_pad ,
		_w9205_,
		_w9206_,
		_w22658_
	);
	LUT3 #(
		.INIT('h2a)
	) name20758 (
		\m1_sel_i[2]_pad ,
		_w9205_,
		_w9206_,
		_w22659_
	);
	LUT4 #(
		.INIT('h57df)
	) name20759 (
		_w9200_,
		_w9203_,
		_w22658_,
		_w22659_,
		_w22660_
	);
	LUT3 #(
		.INIT('h80)
	) name20760 (
		\m0_sel_i[2]_pad ,
		_w9205_,
		_w9206_,
		_w22661_
	);
	LUT3 #(
		.INIT('h2a)
	) name20761 (
		\m7_sel_i[2]_pad ,
		_w9205_,
		_w9206_,
		_w22662_
	);
	LUT4 #(
		.INIT('h6e7f)
	) name20762 (
		_w9200_,
		_w9203_,
		_w22661_,
		_w22662_,
		_w22663_
	);
	LUT4 #(
		.INIT('h7fff)
	) name20763 (
		_w22654_,
		_w22657_,
		_w22660_,
		_w22663_,
		_w22664_
	);
	LUT3 #(
		.INIT('h2a)
	) name20764 (
		\m3_sel_i[3]_pad ,
		_w9205_,
		_w9206_,
		_w22665_
	);
	LUT3 #(
		.INIT('h80)
	) name20765 (
		\m4_sel_i[3]_pad ,
		_w9205_,
		_w9206_,
		_w22666_
	);
	LUT4 #(
		.INIT('h9dbf)
	) name20766 (
		_w9200_,
		_w9203_,
		_w22665_,
		_w22666_,
		_w22667_
	);
	LUT3 #(
		.INIT('h80)
	) name20767 (
		\m6_sel_i[3]_pad ,
		_w9205_,
		_w9206_,
		_w22668_
	);
	LUT3 #(
		.INIT('h80)
	) name20768 (
		\m2_sel_i[3]_pad ,
		_w9205_,
		_w9206_,
		_w22669_
	);
	LUT4 #(
		.INIT('habef)
	) name20769 (
		_w9200_,
		_w9203_,
		_w22668_,
		_w22669_,
		_w22670_
	);
	LUT3 #(
		.INIT('h2a)
	) name20770 (
		\m5_sel_i[3]_pad ,
		_w9205_,
		_w9206_,
		_w22671_
	);
	LUT3 #(
		.INIT('h2a)
	) name20771 (
		\m1_sel_i[3]_pad ,
		_w9205_,
		_w9206_,
		_w22672_
	);
	LUT4 #(
		.INIT('h57df)
	) name20772 (
		_w9200_,
		_w9203_,
		_w22671_,
		_w22672_,
		_w22673_
	);
	LUT3 #(
		.INIT('h80)
	) name20773 (
		\m0_sel_i[3]_pad ,
		_w9205_,
		_w9206_,
		_w22674_
	);
	LUT3 #(
		.INIT('h2a)
	) name20774 (
		\m7_sel_i[3]_pad ,
		_w9205_,
		_w9206_,
		_w22675_
	);
	LUT4 #(
		.INIT('h6e7f)
	) name20775 (
		_w9200_,
		_w9203_,
		_w22674_,
		_w22675_,
		_w22676_
	);
	LUT4 #(
		.INIT('h7fff)
	) name20776 (
		_w22667_,
		_w22670_,
		_w22673_,
		_w22676_,
		_w22677_
	);
	LUT4 #(
		.INIT('h2a00)
	) name20777 (
		\m7_stb_i_pad ,
		_w9205_,
		_w9206_,
		_w9611_,
		_w22678_
	);
	LUT4 #(
		.INIT('h8000)
	) name20778 (
		\m6_stb_i_pad ,
		_w9205_,
		_w9206_,
		_w9579_,
		_w22679_
	);
	LUT3 #(
		.INIT('h57)
	) name20779 (
		_w9218_,
		_w22678_,
		_w22679_,
		_w22680_
	);
	LUT4 #(
		.INIT('h8000)
	) name20780 (
		\m2_stb_i_pad ,
		_w9205_,
		_w9206_,
		_w9465_,
		_w22681_
	);
	LUT4 #(
		.INIT('h2a00)
	) name20781 (
		\m3_stb_i_pad ,
		_w9205_,
		_w9206_,
		_w9416_,
		_w22682_
	);
	LUT3 #(
		.INIT('h57)
	) name20782 (
		_w9212_,
		_w22681_,
		_w22682_,
		_w22683_
	);
	LUT4 #(
		.INIT('h2a00)
	) name20783 (
		\m1_stb_i_pad ,
		_w9205_,
		_w9206_,
		_w9430_,
		_w22684_
	);
	LUT4 #(
		.INIT('h2a00)
	) name20784 (
		\m5_stb_i_pad ,
		_w9205_,
		_w9206_,
		_w9351_,
		_w22685_
	);
	LUT4 #(
		.INIT('h5d7f)
	) name20785 (
		_w9200_,
		_w9203_,
		_w22684_,
		_w22685_,
		_w22686_
	);
	LUT4 #(
		.INIT('h8000)
	) name20786 (
		\m4_stb_i_pad ,
		_w9205_,
		_w9206_,
		_w9523_,
		_w22687_
	);
	LUT4 #(
		.INIT('h8000)
	) name20787 (
		\m0_stb_i_pad ,
		_w9205_,
		_w9206_,
		_w9398_,
		_w22688_
	);
	LUT4 #(
		.INIT('h57df)
	) name20788 (
		_w9200_,
		_w9203_,
		_w22687_,
		_w22688_,
		_w22689_
	);
	LUT4 #(
		.INIT('h7fff)
	) name20789 (
		_w22680_,
		_w22683_,
		_w22686_,
		_w22689_,
		_w22690_
	);
	LUT3 #(
		.INIT('h2a)
	) name20790 (
		\m3_we_i_pad ,
		_w9205_,
		_w9206_,
		_w22691_
	);
	LUT3 #(
		.INIT('h80)
	) name20791 (
		\m4_we_i_pad ,
		_w9205_,
		_w9206_,
		_w22692_
	);
	LUT4 #(
		.INIT('h9dbf)
	) name20792 (
		_w9200_,
		_w9203_,
		_w22691_,
		_w22692_,
		_w22693_
	);
	LUT3 #(
		.INIT('h80)
	) name20793 (
		\m6_we_i_pad ,
		_w9205_,
		_w9206_,
		_w22694_
	);
	LUT3 #(
		.INIT('h80)
	) name20794 (
		\m2_we_i_pad ,
		_w9205_,
		_w9206_,
		_w22695_
	);
	LUT4 #(
		.INIT('habef)
	) name20795 (
		_w9200_,
		_w9203_,
		_w22694_,
		_w22695_,
		_w22696_
	);
	LUT3 #(
		.INIT('h2a)
	) name20796 (
		\m5_we_i_pad ,
		_w9205_,
		_w9206_,
		_w22697_
	);
	LUT3 #(
		.INIT('h2a)
	) name20797 (
		\m1_we_i_pad ,
		_w9205_,
		_w9206_,
		_w22698_
	);
	LUT4 #(
		.INIT('h57df)
	) name20798 (
		_w9200_,
		_w9203_,
		_w22697_,
		_w22698_,
		_w22699_
	);
	LUT3 #(
		.INIT('h80)
	) name20799 (
		\m0_we_i_pad ,
		_w9205_,
		_w9206_,
		_w22700_
	);
	LUT3 #(
		.INIT('h2a)
	) name20800 (
		\m7_we_i_pad ,
		_w9205_,
		_w9206_,
		_w22701_
	);
	LUT4 #(
		.INIT('h6e7f)
	) name20801 (
		_w9200_,
		_w9203_,
		_w22700_,
		_w22701_,
		_w22702_
	);
	LUT4 #(
		.INIT('h7fff)
	) name20802 (
		_w22693_,
		_w22696_,
		_w22699_,
		_w22702_,
		_w22703_
	);
	LUT3 #(
		.INIT('h2a)
	) name20803 (
		\m3_addr_i[0]_pad ,
		_w8655_,
		_w8656_,
		_w22704_
	);
	LUT3 #(
		.INIT('h80)
	) name20804 (
		\m4_addr_i[0]_pad ,
		_w8655_,
		_w8656_,
		_w22705_
	);
	LUT4 #(
		.INIT('h9dbf)
	) name20805 (
		_w8650_,
		_w8653_,
		_w22704_,
		_w22705_,
		_w22706_
	);
	LUT3 #(
		.INIT('h80)
	) name20806 (
		\m6_addr_i[0]_pad ,
		_w8655_,
		_w8656_,
		_w22707_
	);
	LUT3 #(
		.INIT('h80)
	) name20807 (
		\m2_addr_i[0]_pad ,
		_w8655_,
		_w8656_,
		_w22708_
	);
	LUT4 #(
		.INIT('habef)
	) name20808 (
		_w8650_,
		_w8653_,
		_w22707_,
		_w22708_,
		_w22709_
	);
	LUT3 #(
		.INIT('h2a)
	) name20809 (
		\m5_addr_i[0]_pad ,
		_w8655_,
		_w8656_,
		_w22710_
	);
	LUT3 #(
		.INIT('h2a)
	) name20810 (
		\m1_addr_i[0]_pad ,
		_w8655_,
		_w8656_,
		_w22711_
	);
	LUT4 #(
		.INIT('h57df)
	) name20811 (
		_w8650_,
		_w8653_,
		_w22710_,
		_w22711_,
		_w22712_
	);
	LUT3 #(
		.INIT('h80)
	) name20812 (
		\m0_addr_i[0]_pad ,
		_w8655_,
		_w8656_,
		_w22713_
	);
	LUT3 #(
		.INIT('h2a)
	) name20813 (
		\m7_addr_i[0]_pad ,
		_w8655_,
		_w8656_,
		_w22714_
	);
	LUT4 #(
		.INIT('h6e7f)
	) name20814 (
		_w8650_,
		_w8653_,
		_w22713_,
		_w22714_,
		_w22715_
	);
	LUT4 #(
		.INIT('h7fff)
	) name20815 (
		_w22706_,
		_w22709_,
		_w22712_,
		_w22715_,
		_w22716_
	);
	LUT3 #(
		.INIT('h2a)
	) name20816 (
		\m3_addr_i[10]_pad ,
		_w8655_,
		_w8656_,
		_w22717_
	);
	LUT3 #(
		.INIT('h80)
	) name20817 (
		\m4_addr_i[10]_pad ,
		_w8655_,
		_w8656_,
		_w22718_
	);
	LUT4 #(
		.INIT('h9dbf)
	) name20818 (
		_w8650_,
		_w8653_,
		_w22717_,
		_w22718_,
		_w22719_
	);
	LUT3 #(
		.INIT('h80)
	) name20819 (
		\m6_addr_i[10]_pad ,
		_w8655_,
		_w8656_,
		_w22720_
	);
	LUT3 #(
		.INIT('h80)
	) name20820 (
		\m2_addr_i[10]_pad ,
		_w8655_,
		_w8656_,
		_w22721_
	);
	LUT4 #(
		.INIT('habef)
	) name20821 (
		_w8650_,
		_w8653_,
		_w22720_,
		_w22721_,
		_w22722_
	);
	LUT3 #(
		.INIT('h2a)
	) name20822 (
		\m5_addr_i[10]_pad ,
		_w8655_,
		_w8656_,
		_w22723_
	);
	LUT3 #(
		.INIT('h2a)
	) name20823 (
		\m1_addr_i[10]_pad ,
		_w8655_,
		_w8656_,
		_w22724_
	);
	LUT4 #(
		.INIT('h57df)
	) name20824 (
		_w8650_,
		_w8653_,
		_w22723_,
		_w22724_,
		_w22725_
	);
	LUT3 #(
		.INIT('h80)
	) name20825 (
		\m0_addr_i[10]_pad ,
		_w8655_,
		_w8656_,
		_w22726_
	);
	LUT3 #(
		.INIT('h2a)
	) name20826 (
		\m7_addr_i[10]_pad ,
		_w8655_,
		_w8656_,
		_w22727_
	);
	LUT4 #(
		.INIT('h6e7f)
	) name20827 (
		_w8650_,
		_w8653_,
		_w22726_,
		_w22727_,
		_w22728_
	);
	LUT4 #(
		.INIT('h7fff)
	) name20828 (
		_w22719_,
		_w22722_,
		_w22725_,
		_w22728_,
		_w22729_
	);
	LUT3 #(
		.INIT('h2a)
	) name20829 (
		\m3_addr_i[11]_pad ,
		_w8655_,
		_w8656_,
		_w22730_
	);
	LUT3 #(
		.INIT('h80)
	) name20830 (
		\m4_addr_i[11]_pad ,
		_w8655_,
		_w8656_,
		_w22731_
	);
	LUT4 #(
		.INIT('h9dbf)
	) name20831 (
		_w8650_,
		_w8653_,
		_w22730_,
		_w22731_,
		_w22732_
	);
	LUT3 #(
		.INIT('h80)
	) name20832 (
		\m6_addr_i[11]_pad ,
		_w8655_,
		_w8656_,
		_w22733_
	);
	LUT3 #(
		.INIT('h80)
	) name20833 (
		\m2_addr_i[11]_pad ,
		_w8655_,
		_w8656_,
		_w22734_
	);
	LUT4 #(
		.INIT('habef)
	) name20834 (
		_w8650_,
		_w8653_,
		_w22733_,
		_w22734_,
		_w22735_
	);
	LUT3 #(
		.INIT('h2a)
	) name20835 (
		\m5_addr_i[11]_pad ,
		_w8655_,
		_w8656_,
		_w22736_
	);
	LUT3 #(
		.INIT('h2a)
	) name20836 (
		\m1_addr_i[11]_pad ,
		_w8655_,
		_w8656_,
		_w22737_
	);
	LUT4 #(
		.INIT('h57df)
	) name20837 (
		_w8650_,
		_w8653_,
		_w22736_,
		_w22737_,
		_w22738_
	);
	LUT3 #(
		.INIT('h80)
	) name20838 (
		\m0_addr_i[11]_pad ,
		_w8655_,
		_w8656_,
		_w22739_
	);
	LUT3 #(
		.INIT('h2a)
	) name20839 (
		\m7_addr_i[11]_pad ,
		_w8655_,
		_w8656_,
		_w22740_
	);
	LUT4 #(
		.INIT('h6e7f)
	) name20840 (
		_w8650_,
		_w8653_,
		_w22739_,
		_w22740_,
		_w22741_
	);
	LUT4 #(
		.INIT('h7fff)
	) name20841 (
		_w22732_,
		_w22735_,
		_w22738_,
		_w22741_,
		_w22742_
	);
	LUT3 #(
		.INIT('h2a)
	) name20842 (
		\m3_addr_i[12]_pad ,
		_w8655_,
		_w8656_,
		_w22743_
	);
	LUT3 #(
		.INIT('h80)
	) name20843 (
		\m4_addr_i[12]_pad ,
		_w8655_,
		_w8656_,
		_w22744_
	);
	LUT4 #(
		.INIT('h9dbf)
	) name20844 (
		_w8650_,
		_w8653_,
		_w22743_,
		_w22744_,
		_w22745_
	);
	LUT3 #(
		.INIT('h80)
	) name20845 (
		\m6_addr_i[12]_pad ,
		_w8655_,
		_w8656_,
		_w22746_
	);
	LUT3 #(
		.INIT('h80)
	) name20846 (
		\m2_addr_i[12]_pad ,
		_w8655_,
		_w8656_,
		_w22747_
	);
	LUT4 #(
		.INIT('habef)
	) name20847 (
		_w8650_,
		_w8653_,
		_w22746_,
		_w22747_,
		_w22748_
	);
	LUT3 #(
		.INIT('h2a)
	) name20848 (
		\m5_addr_i[12]_pad ,
		_w8655_,
		_w8656_,
		_w22749_
	);
	LUT3 #(
		.INIT('h2a)
	) name20849 (
		\m1_addr_i[12]_pad ,
		_w8655_,
		_w8656_,
		_w22750_
	);
	LUT4 #(
		.INIT('h57df)
	) name20850 (
		_w8650_,
		_w8653_,
		_w22749_,
		_w22750_,
		_w22751_
	);
	LUT3 #(
		.INIT('h80)
	) name20851 (
		\m0_addr_i[12]_pad ,
		_w8655_,
		_w8656_,
		_w22752_
	);
	LUT3 #(
		.INIT('h2a)
	) name20852 (
		\m7_addr_i[12]_pad ,
		_w8655_,
		_w8656_,
		_w22753_
	);
	LUT4 #(
		.INIT('h6e7f)
	) name20853 (
		_w8650_,
		_w8653_,
		_w22752_,
		_w22753_,
		_w22754_
	);
	LUT4 #(
		.INIT('h7fff)
	) name20854 (
		_w22745_,
		_w22748_,
		_w22751_,
		_w22754_,
		_w22755_
	);
	LUT3 #(
		.INIT('h2a)
	) name20855 (
		\m3_addr_i[13]_pad ,
		_w8655_,
		_w8656_,
		_w22756_
	);
	LUT3 #(
		.INIT('h80)
	) name20856 (
		\m4_addr_i[13]_pad ,
		_w8655_,
		_w8656_,
		_w22757_
	);
	LUT4 #(
		.INIT('h9dbf)
	) name20857 (
		_w8650_,
		_w8653_,
		_w22756_,
		_w22757_,
		_w22758_
	);
	LUT3 #(
		.INIT('h80)
	) name20858 (
		\m6_addr_i[13]_pad ,
		_w8655_,
		_w8656_,
		_w22759_
	);
	LUT3 #(
		.INIT('h80)
	) name20859 (
		\m2_addr_i[13]_pad ,
		_w8655_,
		_w8656_,
		_w22760_
	);
	LUT4 #(
		.INIT('habef)
	) name20860 (
		_w8650_,
		_w8653_,
		_w22759_,
		_w22760_,
		_w22761_
	);
	LUT3 #(
		.INIT('h2a)
	) name20861 (
		\m5_addr_i[13]_pad ,
		_w8655_,
		_w8656_,
		_w22762_
	);
	LUT3 #(
		.INIT('h2a)
	) name20862 (
		\m1_addr_i[13]_pad ,
		_w8655_,
		_w8656_,
		_w22763_
	);
	LUT4 #(
		.INIT('h57df)
	) name20863 (
		_w8650_,
		_w8653_,
		_w22762_,
		_w22763_,
		_w22764_
	);
	LUT3 #(
		.INIT('h80)
	) name20864 (
		\m0_addr_i[13]_pad ,
		_w8655_,
		_w8656_,
		_w22765_
	);
	LUT3 #(
		.INIT('h2a)
	) name20865 (
		\m7_addr_i[13]_pad ,
		_w8655_,
		_w8656_,
		_w22766_
	);
	LUT4 #(
		.INIT('h6e7f)
	) name20866 (
		_w8650_,
		_w8653_,
		_w22765_,
		_w22766_,
		_w22767_
	);
	LUT4 #(
		.INIT('h7fff)
	) name20867 (
		_w22758_,
		_w22761_,
		_w22764_,
		_w22767_,
		_w22768_
	);
	LUT3 #(
		.INIT('h2a)
	) name20868 (
		\m3_addr_i[14]_pad ,
		_w8655_,
		_w8656_,
		_w22769_
	);
	LUT3 #(
		.INIT('h80)
	) name20869 (
		\m4_addr_i[14]_pad ,
		_w8655_,
		_w8656_,
		_w22770_
	);
	LUT4 #(
		.INIT('h9dbf)
	) name20870 (
		_w8650_,
		_w8653_,
		_w22769_,
		_w22770_,
		_w22771_
	);
	LUT3 #(
		.INIT('h80)
	) name20871 (
		\m6_addr_i[14]_pad ,
		_w8655_,
		_w8656_,
		_w22772_
	);
	LUT3 #(
		.INIT('h80)
	) name20872 (
		\m2_addr_i[14]_pad ,
		_w8655_,
		_w8656_,
		_w22773_
	);
	LUT4 #(
		.INIT('habef)
	) name20873 (
		_w8650_,
		_w8653_,
		_w22772_,
		_w22773_,
		_w22774_
	);
	LUT3 #(
		.INIT('h2a)
	) name20874 (
		\m5_addr_i[14]_pad ,
		_w8655_,
		_w8656_,
		_w22775_
	);
	LUT3 #(
		.INIT('h2a)
	) name20875 (
		\m1_addr_i[14]_pad ,
		_w8655_,
		_w8656_,
		_w22776_
	);
	LUT4 #(
		.INIT('h57df)
	) name20876 (
		_w8650_,
		_w8653_,
		_w22775_,
		_w22776_,
		_w22777_
	);
	LUT3 #(
		.INIT('h80)
	) name20877 (
		\m0_addr_i[14]_pad ,
		_w8655_,
		_w8656_,
		_w22778_
	);
	LUT3 #(
		.INIT('h2a)
	) name20878 (
		\m7_addr_i[14]_pad ,
		_w8655_,
		_w8656_,
		_w22779_
	);
	LUT4 #(
		.INIT('h6e7f)
	) name20879 (
		_w8650_,
		_w8653_,
		_w22778_,
		_w22779_,
		_w22780_
	);
	LUT4 #(
		.INIT('h7fff)
	) name20880 (
		_w22771_,
		_w22774_,
		_w22777_,
		_w22780_,
		_w22781_
	);
	LUT3 #(
		.INIT('h2a)
	) name20881 (
		\m3_addr_i[15]_pad ,
		_w8655_,
		_w8656_,
		_w22782_
	);
	LUT3 #(
		.INIT('h80)
	) name20882 (
		\m4_addr_i[15]_pad ,
		_w8655_,
		_w8656_,
		_w22783_
	);
	LUT4 #(
		.INIT('h9dbf)
	) name20883 (
		_w8650_,
		_w8653_,
		_w22782_,
		_w22783_,
		_w22784_
	);
	LUT3 #(
		.INIT('h80)
	) name20884 (
		\m6_addr_i[15]_pad ,
		_w8655_,
		_w8656_,
		_w22785_
	);
	LUT3 #(
		.INIT('h80)
	) name20885 (
		\m2_addr_i[15]_pad ,
		_w8655_,
		_w8656_,
		_w22786_
	);
	LUT4 #(
		.INIT('habef)
	) name20886 (
		_w8650_,
		_w8653_,
		_w22785_,
		_w22786_,
		_w22787_
	);
	LUT3 #(
		.INIT('h2a)
	) name20887 (
		\m5_addr_i[15]_pad ,
		_w8655_,
		_w8656_,
		_w22788_
	);
	LUT3 #(
		.INIT('h2a)
	) name20888 (
		\m1_addr_i[15]_pad ,
		_w8655_,
		_w8656_,
		_w22789_
	);
	LUT4 #(
		.INIT('h57df)
	) name20889 (
		_w8650_,
		_w8653_,
		_w22788_,
		_w22789_,
		_w22790_
	);
	LUT3 #(
		.INIT('h80)
	) name20890 (
		\m0_addr_i[15]_pad ,
		_w8655_,
		_w8656_,
		_w22791_
	);
	LUT3 #(
		.INIT('h2a)
	) name20891 (
		\m7_addr_i[15]_pad ,
		_w8655_,
		_w8656_,
		_w22792_
	);
	LUT4 #(
		.INIT('h6e7f)
	) name20892 (
		_w8650_,
		_w8653_,
		_w22791_,
		_w22792_,
		_w22793_
	);
	LUT4 #(
		.INIT('h7fff)
	) name20893 (
		_w22784_,
		_w22787_,
		_w22790_,
		_w22793_,
		_w22794_
	);
	LUT3 #(
		.INIT('h2a)
	) name20894 (
		\m3_addr_i[16]_pad ,
		_w8655_,
		_w8656_,
		_w22795_
	);
	LUT3 #(
		.INIT('h80)
	) name20895 (
		\m4_addr_i[16]_pad ,
		_w8655_,
		_w8656_,
		_w22796_
	);
	LUT4 #(
		.INIT('h9dbf)
	) name20896 (
		_w8650_,
		_w8653_,
		_w22795_,
		_w22796_,
		_w22797_
	);
	LUT3 #(
		.INIT('h80)
	) name20897 (
		\m6_addr_i[16]_pad ,
		_w8655_,
		_w8656_,
		_w22798_
	);
	LUT3 #(
		.INIT('h80)
	) name20898 (
		\m2_addr_i[16]_pad ,
		_w8655_,
		_w8656_,
		_w22799_
	);
	LUT4 #(
		.INIT('habef)
	) name20899 (
		_w8650_,
		_w8653_,
		_w22798_,
		_w22799_,
		_w22800_
	);
	LUT3 #(
		.INIT('h2a)
	) name20900 (
		\m5_addr_i[16]_pad ,
		_w8655_,
		_w8656_,
		_w22801_
	);
	LUT3 #(
		.INIT('h2a)
	) name20901 (
		\m1_addr_i[16]_pad ,
		_w8655_,
		_w8656_,
		_w22802_
	);
	LUT4 #(
		.INIT('h57df)
	) name20902 (
		_w8650_,
		_w8653_,
		_w22801_,
		_w22802_,
		_w22803_
	);
	LUT3 #(
		.INIT('h80)
	) name20903 (
		\m0_addr_i[16]_pad ,
		_w8655_,
		_w8656_,
		_w22804_
	);
	LUT3 #(
		.INIT('h2a)
	) name20904 (
		\m7_addr_i[16]_pad ,
		_w8655_,
		_w8656_,
		_w22805_
	);
	LUT4 #(
		.INIT('h6e7f)
	) name20905 (
		_w8650_,
		_w8653_,
		_w22804_,
		_w22805_,
		_w22806_
	);
	LUT4 #(
		.INIT('h7fff)
	) name20906 (
		_w22797_,
		_w22800_,
		_w22803_,
		_w22806_,
		_w22807_
	);
	LUT3 #(
		.INIT('h2a)
	) name20907 (
		\m3_addr_i[17]_pad ,
		_w8655_,
		_w8656_,
		_w22808_
	);
	LUT3 #(
		.INIT('h80)
	) name20908 (
		\m4_addr_i[17]_pad ,
		_w8655_,
		_w8656_,
		_w22809_
	);
	LUT4 #(
		.INIT('h9dbf)
	) name20909 (
		_w8650_,
		_w8653_,
		_w22808_,
		_w22809_,
		_w22810_
	);
	LUT3 #(
		.INIT('h80)
	) name20910 (
		\m6_addr_i[17]_pad ,
		_w8655_,
		_w8656_,
		_w22811_
	);
	LUT3 #(
		.INIT('h80)
	) name20911 (
		\m2_addr_i[17]_pad ,
		_w8655_,
		_w8656_,
		_w22812_
	);
	LUT4 #(
		.INIT('habef)
	) name20912 (
		_w8650_,
		_w8653_,
		_w22811_,
		_w22812_,
		_w22813_
	);
	LUT3 #(
		.INIT('h2a)
	) name20913 (
		\m5_addr_i[17]_pad ,
		_w8655_,
		_w8656_,
		_w22814_
	);
	LUT3 #(
		.INIT('h2a)
	) name20914 (
		\m1_addr_i[17]_pad ,
		_w8655_,
		_w8656_,
		_w22815_
	);
	LUT4 #(
		.INIT('h57df)
	) name20915 (
		_w8650_,
		_w8653_,
		_w22814_,
		_w22815_,
		_w22816_
	);
	LUT3 #(
		.INIT('h80)
	) name20916 (
		\m0_addr_i[17]_pad ,
		_w8655_,
		_w8656_,
		_w22817_
	);
	LUT3 #(
		.INIT('h2a)
	) name20917 (
		\m7_addr_i[17]_pad ,
		_w8655_,
		_w8656_,
		_w22818_
	);
	LUT4 #(
		.INIT('h6e7f)
	) name20918 (
		_w8650_,
		_w8653_,
		_w22817_,
		_w22818_,
		_w22819_
	);
	LUT4 #(
		.INIT('h7fff)
	) name20919 (
		_w22810_,
		_w22813_,
		_w22816_,
		_w22819_,
		_w22820_
	);
	LUT3 #(
		.INIT('h2a)
	) name20920 (
		\m3_addr_i[18]_pad ,
		_w8655_,
		_w8656_,
		_w22821_
	);
	LUT3 #(
		.INIT('h80)
	) name20921 (
		\m4_addr_i[18]_pad ,
		_w8655_,
		_w8656_,
		_w22822_
	);
	LUT4 #(
		.INIT('h9dbf)
	) name20922 (
		_w8650_,
		_w8653_,
		_w22821_,
		_w22822_,
		_w22823_
	);
	LUT3 #(
		.INIT('h80)
	) name20923 (
		\m6_addr_i[18]_pad ,
		_w8655_,
		_w8656_,
		_w22824_
	);
	LUT3 #(
		.INIT('h80)
	) name20924 (
		\m2_addr_i[18]_pad ,
		_w8655_,
		_w8656_,
		_w22825_
	);
	LUT4 #(
		.INIT('habef)
	) name20925 (
		_w8650_,
		_w8653_,
		_w22824_,
		_w22825_,
		_w22826_
	);
	LUT3 #(
		.INIT('h2a)
	) name20926 (
		\m5_addr_i[18]_pad ,
		_w8655_,
		_w8656_,
		_w22827_
	);
	LUT3 #(
		.INIT('h2a)
	) name20927 (
		\m1_addr_i[18]_pad ,
		_w8655_,
		_w8656_,
		_w22828_
	);
	LUT4 #(
		.INIT('h57df)
	) name20928 (
		_w8650_,
		_w8653_,
		_w22827_,
		_w22828_,
		_w22829_
	);
	LUT3 #(
		.INIT('h80)
	) name20929 (
		\m0_addr_i[18]_pad ,
		_w8655_,
		_w8656_,
		_w22830_
	);
	LUT3 #(
		.INIT('h2a)
	) name20930 (
		\m7_addr_i[18]_pad ,
		_w8655_,
		_w8656_,
		_w22831_
	);
	LUT4 #(
		.INIT('h6e7f)
	) name20931 (
		_w8650_,
		_w8653_,
		_w22830_,
		_w22831_,
		_w22832_
	);
	LUT4 #(
		.INIT('h7fff)
	) name20932 (
		_w22823_,
		_w22826_,
		_w22829_,
		_w22832_,
		_w22833_
	);
	LUT3 #(
		.INIT('h2a)
	) name20933 (
		\m3_addr_i[19]_pad ,
		_w8655_,
		_w8656_,
		_w22834_
	);
	LUT3 #(
		.INIT('h80)
	) name20934 (
		\m4_addr_i[19]_pad ,
		_w8655_,
		_w8656_,
		_w22835_
	);
	LUT4 #(
		.INIT('h9dbf)
	) name20935 (
		_w8650_,
		_w8653_,
		_w22834_,
		_w22835_,
		_w22836_
	);
	LUT3 #(
		.INIT('h80)
	) name20936 (
		\m6_addr_i[19]_pad ,
		_w8655_,
		_w8656_,
		_w22837_
	);
	LUT3 #(
		.INIT('h80)
	) name20937 (
		\m2_addr_i[19]_pad ,
		_w8655_,
		_w8656_,
		_w22838_
	);
	LUT4 #(
		.INIT('habef)
	) name20938 (
		_w8650_,
		_w8653_,
		_w22837_,
		_w22838_,
		_w22839_
	);
	LUT3 #(
		.INIT('h2a)
	) name20939 (
		\m5_addr_i[19]_pad ,
		_w8655_,
		_w8656_,
		_w22840_
	);
	LUT3 #(
		.INIT('h2a)
	) name20940 (
		\m1_addr_i[19]_pad ,
		_w8655_,
		_w8656_,
		_w22841_
	);
	LUT4 #(
		.INIT('h57df)
	) name20941 (
		_w8650_,
		_w8653_,
		_w22840_,
		_w22841_,
		_w22842_
	);
	LUT3 #(
		.INIT('h80)
	) name20942 (
		\m0_addr_i[19]_pad ,
		_w8655_,
		_w8656_,
		_w22843_
	);
	LUT3 #(
		.INIT('h2a)
	) name20943 (
		\m7_addr_i[19]_pad ,
		_w8655_,
		_w8656_,
		_w22844_
	);
	LUT4 #(
		.INIT('h6e7f)
	) name20944 (
		_w8650_,
		_w8653_,
		_w22843_,
		_w22844_,
		_w22845_
	);
	LUT4 #(
		.INIT('h7fff)
	) name20945 (
		_w22836_,
		_w22839_,
		_w22842_,
		_w22845_,
		_w22846_
	);
	LUT3 #(
		.INIT('h2a)
	) name20946 (
		\m3_addr_i[1]_pad ,
		_w8655_,
		_w8656_,
		_w22847_
	);
	LUT3 #(
		.INIT('h80)
	) name20947 (
		\m4_addr_i[1]_pad ,
		_w8655_,
		_w8656_,
		_w22848_
	);
	LUT4 #(
		.INIT('h9dbf)
	) name20948 (
		_w8650_,
		_w8653_,
		_w22847_,
		_w22848_,
		_w22849_
	);
	LUT3 #(
		.INIT('h80)
	) name20949 (
		\m6_addr_i[1]_pad ,
		_w8655_,
		_w8656_,
		_w22850_
	);
	LUT3 #(
		.INIT('h80)
	) name20950 (
		\m2_addr_i[1]_pad ,
		_w8655_,
		_w8656_,
		_w22851_
	);
	LUT4 #(
		.INIT('habef)
	) name20951 (
		_w8650_,
		_w8653_,
		_w22850_,
		_w22851_,
		_w22852_
	);
	LUT3 #(
		.INIT('h2a)
	) name20952 (
		\m5_addr_i[1]_pad ,
		_w8655_,
		_w8656_,
		_w22853_
	);
	LUT3 #(
		.INIT('h2a)
	) name20953 (
		\m1_addr_i[1]_pad ,
		_w8655_,
		_w8656_,
		_w22854_
	);
	LUT4 #(
		.INIT('h57df)
	) name20954 (
		_w8650_,
		_w8653_,
		_w22853_,
		_w22854_,
		_w22855_
	);
	LUT3 #(
		.INIT('h80)
	) name20955 (
		\m0_addr_i[1]_pad ,
		_w8655_,
		_w8656_,
		_w22856_
	);
	LUT3 #(
		.INIT('h2a)
	) name20956 (
		\m7_addr_i[1]_pad ,
		_w8655_,
		_w8656_,
		_w22857_
	);
	LUT4 #(
		.INIT('h6e7f)
	) name20957 (
		_w8650_,
		_w8653_,
		_w22856_,
		_w22857_,
		_w22858_
	);
	LUT4 #(
		.INIT('h7fff)
	) name20958 (
		_w22849_,
		_w22852_,
		_w22855_,
		_w22858_,
		_w22859_
	);
	LUT3 #(
		.INIT('h2a)
	) name20959 (
		\m3_addr_i[20]_pad ,
		_w8655_,
		_w8656_,
		_w22860_
	);
	LUT3 #(
		.INIT('h80)
	) name20960 (
		\m4_addr_i[20]_pad ,
		_w8655_,
		_w8656_,
		_w22861_
	);
	LUT4 #(
		.INIT('h9dbf)
	) name20961 (
		_w8650_,
		_w8653_,
		_w22860_,
		_w22861_,
		_w22862_
	);
	LUT3 #(
		.INIT('h80)
	) name20962 (
		\m6_addr_i[20]_pad ,
		_w8655_,
		_w8656_,
		_w22863_
	);
	LUT3 #(
		.INIT('h80)
	) name20963 (
		\m2_addr_i[20]_pad ,
		_w8655_,
		_w8656_,
		_w22864_
	);
	LUT4 #(
		.INIT('habef)
	) name20964 (
		_w8650_,
		_w8653_,
		_w22863_,
		_w22864_,
		_w22865_
	);
	LUT3 #(
		.INIT('h2a)
	) name20965 (
		\m5_addr_i[20]_pad ,
		_w8655_,
		_w8656_,
		_w22866_
	);
	LUT3 #(
		.INIT('h2a)
	) name20966 (
		\m1_addr_i[20]_pad ,
		_w8655_,
		_w8656_,
		_w22867_
	);
	LUT4 #(
		.INIT('h57df)
	) name20967 (
		_w8650_,
		_w8653_,
		_w22866_,
		_w22867_,
		_w22868_
	);
	LUT3 #(
		.INIT('h80)
	) name20968 (
		\m0_addr_i[20]_pad ,
		_w8655_,
		_w8656_,
		_w22869_
	);
	LUT3 #(
		.INIT('h2a)
	) name20969 (
		\m7_addr_i[20]_pad ,
		_w8655_,
		_w8656_,
		_w22870_
	);
	LUT4 #(
		.INIT('h6e7f)
	) name20970 (
		_w8650_,
		_w8653_,
		_w22869_,
		_w22870_,
		_w22871_
	);
	LUT4 #(
		.INIT('h7fff)
	) name20971 (
		_w22862_,
		_w22865_,
		_w22868_,
		_w22871_,
		_w22872_
	);
	LUT3 #(
		.INIT('h2a)
	) name20972 (
		\m3_addr_i[21]_pad ,
		_w8655_,
		_w8656_,
		_w22873_
	);
	LUT3 #(
		.INIT('h80)
	) name20973 (
		\m4_addr_i[21]_pad ,
		_w8655_,
		_w8656_,
		_w22874_
	);
	LUT4 #(
		.INIT('h9dbf)
	) name20974 (
		_w8650_,
		_w8653_,
		_w22873_,
		_w22874_,
		_w22875_
	);
	LUT3 #(
		.INIT('h80)
	) name20975 (
		\m6_addr_i[21]_pad ,
		_w8655_,
		_w8656_,
		_w22876_
	);
	LUT3 #(
		.INIT('h80)
	) name20976 (
		\m2_addr_i[21]_pad ,
		_w8655_,
		_w8656_,
		_w22877_
	);
	LUT4 #(
		.INIT('habef)
	) name20977 (
		_w8650_,
		_w8653_,
		_w22876_,
		_w22877_,
		_w22878_
	);
	LUT3 #(
		.INIT('h2a)
	) name20978 (
		\m5_addr_i[21]_pad ,
		_w8655_,
		_w8656_,
		_w22879_
	);
	LUT3 #(
		.INIT('h2a)
	) name20979 (
		\m1_addr_i[21]_pad ,
		_w8655_,
		_w8656_,
		_w22880_
	);
	LUT4 #(
		.INIT('h57df)
	) name20980 (
		_w8650_,
		_w8653_,
		_w22879_,
		_w22880_,
		_w22881_
	);
	LUT3 #(
		.INIT('h80)
	) name20981 (
		\m0_addr_i[21]_pad ,
		_w8655_,
		_w8656_,
		_w22882_
	);
	LUT3 #(
		.INIT('h2a)
	) name20982 (
		\m7_addr_i[21]_pad ,
		_w8655_,
		_w8656_,
		_w22883_
	);
	LUT4 #(
		.INIT('h6e7f)
	) name20983 (
		_w8650_,
		_w8653_,
		_w22882_,
		_w22883_,
		_w22884_
	);
	LUT4 #(
		.INIT('h7fff)
	) name20984 (
		_w22875_,
		_w22878_,
		_w22881_,
		_w22884_,
		_w22885_
	);
	LUT3 #(
		.INIT('h2a)
	) name20985 (
		\m3_addr_i[22]_pad ,
		_w8655_,
		_w8656_,
		_w22886_
	);
	LUT3 #(
		.INIT('h80)
	) name20986 (
		\m4_addr_i[22]_pad ,
		_w8655_,
		_w8656_,
		_w22887_
	);
	LUT4 #(
		.INIT('h9dbf)
	) name20987 (
		_w8650_,
		_w8653_,
		_w22886_,
		_w22887_,
		_w22888_
	);
	LUT3 #(
		.INIT('h80)
	) name20988 (
		\m6_addr_i[22]_pad ,
		_w8655_,
		_w8656_,
		_w22889_
	);
	LUT3 #(
		.INIT('h80)
	) name20989 (
		\m2_addr_i[22]_pad ,
		_w8655_,
		_w8656_,
		_w22890_
	);
	LUT4 #(
		.INIT('habef)
	) name20990 (
		_w8650_,
		_w8653_,
		_w22889_,
		_w22890_,
		_w22891_
	);
	LUT3 #(
		.INIT('h2a)
	) name20991 (
		\m5_addr_i[22]_pad ,
		_w8655_,
		_w8656_,
		_w22892_
	);
	LUT3 #(
		.INIT('h2a)
	) name20992 (
		\m1_addr_i[22]_pad ,
		_w8655_,
		_w8656_,
		_w22893_
	);
	LUT4 #(
		.INIT('h57df)
	) name20993 (
		_w8650_,
		_w8653_,
		_w22892_,
		_w22893_,
		_w22894_
	);
	LUT3 #(
		.INIT('h80)
	) name20994 (
		\m0_addr_i[22]_pad ,
		_w8655_,
		_w8656_,
		_w22895_
	);
	LUT3 #(
		.INIT('h2a)
	) name20995 (
		\m7_addr_i[22]_pad ,
		_w8655_,
		_w8656_,
		_w22896_
	);
	LUT4 #(
		.INIT('h6e7f)
	) name20996 (
		_w8650_,
		_w8653_,
		_w22895_,
		_w22896_,
		_w22897_
	);
	LUT4 #(
		.INIT('h7fff)
	) name20997 (
		_w22888_,
		_w22891_,
		_w22894_,
		_w22897_,
		_w22898_
	);
	LUT3 #(
		.INIT('h2a)
	) name20998 (
		\m3_addr_i[23]_pad ,
		_w8655_,
		_w8656_,
		_w22899_
	);
	LUT3 #(
		.INIT('h80)
	) name20999 (
		\m4_addr_i[23]_pad ,
		_w8655_,
		_w8656_,
		_w22900_
	);
	LUT4 #(
		.INIT('h9dbf)
	) name21000 (
		_w8650_,
		_w8653_,
		_w22899_,
		_w22900_,
		_w22901_
	);
	LUT3 #(
		.INIT('h80)
	) name21001 (
		\m6_addr_i[23]_pad ,
		_w8655_,
		_w8656_,
		_w22902_
	);
	LUT3 #(
		.INIT('h80)
	) name21002 (
		\m2_addr_i[23]_pad ,
		_w8655_,
		_w8656_,
		_w22903_
	);
	LUT4 #(
		.INIT('habef)
	) name21003 (
		_w8650_,
		_w8653_,
		_w22902_,
		_w22903_,
		_w22904_
	);
	LUT3 #(
		.INIT('h2a)
	) name21004 (
		\m5_addr_i[23]_pad ,
		_w8655_,
		_w8656_,
		_w22905_
	);
	LUT3 #(
		.INIT('h2a)
	) name21005 (
		\m1_addr_i[23]_pad ,
		_w8655_,
		_w8656_,
		_w22906_
	);
	LUT4 #(
		.INIT('h57df)
	) name21006 (
		_w8650_,
		_w8653_,
		_w22905_,
		_w22906_,
		_w22907_
	);
	LUT3 #(
		.INIT('h80)
	) name21007 (
		\m0_addr_i[23]_pad ,
		_w8655_,
		_w8656_,
		_w22908_
	);
	LUT3 #(
		.INIT('h2a)
	) name21008 (
		\m7_addr_i[23]_pad ,
		_w8655_,
		_w8656_,
		_w22909_
	);
	LUT4 #(
		.INIT('h6e7f)
	) name21009 (
		_w8650_,
		_w8653_,
		_w22908_,
		_w22909_,
		_w22910_
	);
	LUT4 #(
		.INIT('h7fff)
	) name21010 (
		_w22901_,
		_w22904_,
		_w22907_,
		_w22910_,
		_w22911_
	);
	LUT3 #(
		.INIT('h2a)
	) name21011 (
		\m3_addr_i[24]_pad ,
		_w8655_,
		_w8656_,
		_w22912_
	);
	LUT3 #(
		.INIT('h80)
	) name21012 (
		\m4_addr_i[24]_pad ,
		_w8655_,
		_w8656_,
		_w22913_
	);
	LUT4 #(
		.INIT('h9dbf)
	) name21013 (
		_w8650_,
		_w8653_,
		_w22912_,
		_w22913_,
		_w22914_
	);
	LUT3 #(
		.INIT('h2a)
	) name21014 (
		\m5_addr_i[24]_pad ,
		_w8655_,
		_w8656_,
		_w22915_
	);
	LUT3 #(
		.INIT('h80)
	) name21015 (
		\m2_addr_i[24]_pad ,
		_w8655_,
		_w8656_,
		_w22916_
	);
	LUT4 #(
		.INIT('h9bdf)
	) name21016 (
		_w8650_,
		_w8653_,
		_w22915_,
		_w22916_,
		_w22917_
	);
	LUT3 #(
		.INIT('h80)
	) name21017 (
		\m6_addr_i[24]_pad ,
		_w8655_,
		_w8656_,
		_w22918_
	);
	LUT3 #(
		.INIT('h2a)
	) name21018 (
		\m1_addr_i[24]_pad ,
		_w8655_,
		_w8656_,
		_w22919_
	);
	LUT4 #(
		.INIT('h67ef)
	) name21019 (
		_w8650_,
		_w8653_,
		_w22918_,
		_w22919_,
		_w22920_
	);
	LUT3 #(
		.INIT('h80)
	) name21020 (
		\m0_addr_i[24]_pad ,
		_w8655_,
		_w8656_,
		_w22921_
	);
	LUT3 #(
		.INIT('h2a)
	) name21021 (
		\m7_addr_i[24]_pad ,
		_w8655_,
		_w8656_,
		_w22922_
	);
	LUT4 #(
		.INIT('h6e7f)
	) name21022 (
		_w8650_,
		_w8653_,
		_w22921_,
		_w22922_,
		_w22923_
	);
	LUT4 #(
		.INIT('h7fff)
	) name21023 (
		_w22914_,
		_w22917_,
		_w22920_,
		_w22923_,
		_w22924_
	);
	LUT3 #(
		.INIT('h2a)
	) name21024 (
		\m3_addr_i[25]_pad ,
		_w8655_,
		_w8656_,
		_w22925_
	);
	LUT3 #(
		.INIT('h80)
	) name21025 (
		\m4_addr_i[25]_pad ,
		_w8655_,
		_w8656_,
		_w22926_
	);
	LUT4 #(
		.INIT('h9dbf)
	) name21026 (
		_w8650_,
		_w8653_,
		_w22925_,
		_w22926_,
		_w22927_
	);
	LUT3 #(
		.INIT('h2a)
	) name21027 (
		\m5_addr_i[25]_pad ,
		_w8655_,
		_w8656_,
		_w22928_
	);
	LUT3 #(
		.INIT('h80)
	) name21028 (
		\m2_addr_i[25]_pad ,
		_w8655_,
		_w8656_,
		_w22929_
	);
	LUT4 #(
		.INIT('h9bdf)
	) name21029 (
		_w8650_,
		_w8653_,
		_w22928_,
		_w22929_,
		_w22930_
	);
	LUT3 #(
		.INIT('h80)
	) name21030 (
		\m6_addr_i[25]_pad ,
		_w8655_,
		_w8656_,
		_w22931_
	);
	LUT3 #(
		.INIT('h2a)
	) name21031 (
		\m1_addr_i[25]_pad ,
		_w8655_,
		_w8656_,
		_w22932_
	);
	LUT4 #(
		.INIT('h67ef)
	) name21032 (
		_w8650_,
		_w8653_,
		_w22931_,
		_w22932_,
		_w22933_
	);
	LUT3 #(
		.INIT('h80)
	) name21033 (
		\m0_addr_i[25]_pad ,
		_w8655_,
		_w8656_,
		_w22934_
	);
	LUT3 #(
		.INIT('h2a)
	) name21034 (
		\m7_addr_i[25]_pad ,
		_w8655_,
		_w8656_,
		_w22935_
	);
	LUT4 #(
		.INIT('h6e7f)
	) name21035 (
		_w8650_,
		_w8653_,
		_w22934_,
		_w22935_,
		_w22936_
	);
	LUT4 #(
		.INIT('h7fff)
	) name21036 (
		_w22927_,
		_w22930_,
		_w22933_,
		_w22936_,
		_w22937_
	);
	LUT3 #(
		.INIT('h2a)
	) name21037 (
		\m3_addr_i[26]_pad ,
		_w8655_,
		_w8656_,
		_w22938_
	);
	LUT3 #(
		.INIT('h80)
	) name21038 (
		\m4_addr_i[26]_pad ,
		_w8655_,
		_w8656_,
		_w22939_
	);
	LUT4 #(
		.INIT('h9dbf)
	) name21039 (
		_w8650_,
		_w8653_,
		_w22938_,
		_w22939_,
		_w22940_
	);
	LUT3 #(
		.INIT('h2a)
	) name21040 (
		\m5_addr_i[26]_pad ,
		_w8655_,
		_w8656_,
		_w22941_
	);
	LUT3 #(
		.INIT('h80)
	) name21041 (
		\m2_addr_i[26]_pad ,
		_w8655_,
		_w8656_,
		_w22942_
	);
	LUT4 #(
		.INIT('h9bdf)
	) name21042 (
		_w8650_,
		_w8653_,
		_w22941_,
		_w22942_,
		_w22943_
	);
	LUT3 #(
		.INIT('h80)
	) name21043 (
		\m6_addr_i[26]_pad ,
		_w8655_,
		_w8656_,
		_w22944_
	);
	LUT3 #(
		.INIT('h2a)
	) name21044 (
		\m1_addr_i[26]_pad ,
		_w8655_,
		_w8656_,
		_w22945_
	);
	LUT4 #(
		.INIT('h67ef)
	) name21045 (
		_w8650_,
		_w8653_,
		_w22944_,
		_w22945_,
		_w22946_
	);
	LUT3 #(
		.INIT('h80)
	) name21046 (
		\m0_addr_i[26]_pad ,
		_w8655_,
		_w8656_,
		_w22947_
	);
	LUT3 #(
		.INIT('h2a)
	) name21047 (
		\m7_addr_i[26]_pad ,
		_w8655_,
		_w8656_,
		_w22948_
	);
	LUT4 #(
		.INIT('h6e7f)
	) name21048 (
		_w8650_,
		_w8653_,
		_w22947_,
		_w22948_,
		_w22949_
	);
	LUT4 #(
		.INIT('h7fff)
	) name21049 (
		_w22940_,
		_w22943_,
		_w22946_,
		_w22949_,
		_w22950_
	);
	LUT3 #(
		.INIT('h2a)
	) name21050 (
		\m3_addr_i[27]_pad ,
		_w8655_,
		_w8656_,
		_w22951_
	);
	LUT3 #(
		.INIT('h80)
	) name21051 (
		\m4_addr_i[27]_pad ,
		_w8655_,
		_w8656_,
		_w22952_
	);
	LUT4 #(
		.INIT('h9dbf)
	) name21052 (
		_w8650_,
		_w8653_,
		_w22951_,
		_w22952_,
		_w22953_
	);
	LUT3 #(
		.INIT('h2a)
	) name21053 (
		\m5_addr_i[27]_pad ,
		_w8655_,
		_w8656_,
		_w22954_
	);
	LUT3 #(
		.INIT('h80)
	) name21054 (
		\m2_addr_i[27]_pad ,
		_w8655_,
		_w8656_,
		_w22955_
	);
	LUT4 #(
		.INIT('h9bdf)
	) name21055 (
		_w8650_,
		_w8653_,
		_w22954_,
		_w22955_,
		_w22956_
	);
	LUT3 #(
		.INIT('h80)
	) name21056 (
		\m6_addr_i[27]_pad ,
		_w8655_,
		_w8656_,
		_w22957_
	);
	LUT3 #(
		.INIT('h2a)
	) name21057 (
		\m1_addr_i[27]_pad ,
		_w8655_,
		_w8656_,
		_w22958_
	);
	LUT4 #(
		.INIT('h67ef)
	) name21058 (
		_w8650_,
		_w8653_,
		_w22957_,
		_w22958_,
		_w22959_
	);
	LUT3 #(
		.INIT('h80)
	) name21059 (
		\m0_addr_i[27]_pad ,
		_w8655_,
		_w8656_,
		_w22960_
	);
	LUT3 #(
		.INIT('h2a)
	) name21060 (
		\m7_addr_i[27]_pad ,
		_w8655_,
		_w8656_,
		_w22961_
	);
	LUT4 #(
		.INIT('h6e7f)
	) name21061 (
		_w8650_,
		_w8653_,
		_w22960_,
		_w22961_,
		_w22962_
	);
	LUT4 #(
		.INIT('h7fff)
	) name21062 (
		_w22953_,
		_w22956_,
		_w22959_,
		_w22962_,
		_w22963_
	);
	LUT3 #(
		.INIT('h2a)
	) name21063 (
		\m3_addr_i[28]_pad ,
		_w8655_,
		_w8656_,
		_w22964_
	);
	LUT3 #(
		.INIT('h80)
	) name21064 (
		\m4_addr_i[28]_pad ,
		_w8655_,
		_w8656_,
		_w22965_
	);
	LUT4 #(
		.INIT('h9dbf)
	) name21065 (
		_w8650_,
		_w8653_,
		_w22964_,
		_w22965_,
		_w22966_
	);
	LUT3 #(
		.INIT('h2a)
	) name21066 (
		\m5_addr_i[28]_pad ,
		_w8655_,
		_w8656_,
		_w22967_
	);
	LUT3 #(
		.INIT('h80)
	) name21067 (
		\m2_addr_i[28]_pad ,
		_w8655_,
		_w8656_,
		_w22968_
	);
	LUT4 #(
		.INIT('h9bdf)
	) name21068 (
		_w8650_,
		_w8653_,
		_w22967_,
		_w22968_,
		_w22969_
	);
	LUT3 #(
		.INIT('h80)
	) name21069 (
		\m6_addr_i[28]_pad ,
		_w8655_,
		_w8656_,
		_w22970_
	);
	LUT3 #(
		.INIT('h2a)
	) name21070 (
		\m1_addr_i[28]_pad ,
		_w8655_,
		_w8656_,
		_w22971_
	);
	LUT4 #(
		.INIT('h67ef)
	) name21071 (
		_w8650_,
		_w8653_,
		_w22970_,
		_w22971_,
		_w22972_
	);
	LUT3 #(
		.INIT('h80)
	) name21072 (
		\m0_addr_i[28]_pad ,
		_w8655_,
		_w8656_,
		_w22973_
	);
	LUT3 #(
		.INIT('h2a)
	) name21073 (
		\m7_addr_i[28]_pad ,
		_w8655_,
		_w8656_,
		_w22974_
	);
	LUT4 #(
		.INIT('h6e7f)
	) name21074 (
		_w8650_,
		_w8653_,
		_w22973_,
		_w22974_,
		_w22975_
	);
	LUT4 #(
		.INIT('h7fff)
	) name21075 (
		_w22966_,
		_w22969_,
		_w22972_,
		_w22975_,
		_w22976_
	);
	LUT3 #(
		.INIT('h2a)
	) name21076 (
		\m3_addr_i[29]_pad ,
		_w8655_,
		_w8656_,
		_w22977_
	);
	LUT3 #(
		.INIT('h80)
	) name21077 (
		\m4_addr_i[29]_pad ,
		_w8655_,
		_w8656_,
		_w22978_
	);
	LUT4 #(
		.INIT('h9dbf)
	) name21078 (
		_w8650_,
		_w8653_,
		_w22977_,
		_w22978_,
		_w22979_
	);
	LUT3 #(
		.INIT('h2a)
	) name21079 (
		\m5_addr_i[29]_pad ,
		_w8655_,
		_w8656_,
		_w22980_
	);
	LUT3 #(
		.INIT('h80)
	) name21080 (
		\m2_addr_i[29]_pad ,
		_w8655_,
		_w8656_,
		_w22981_
	);
	LUT4 #(
		.INIT('h9bdf)
	) name21081 (
		_w8650_,
		_w8653_,
		_w22980_,
		_w22981_,
		_w22982_
	);
	LUT3 #(
		.INIT('h80)
	) name21082 (
		\m6_addr_i[29]_pad ,
		_w8655_,
		_w8656_,
		_w22983_
	);
	LUT3 #(
		.INIT('h2a)
	) name21083 (
		\m1_addr_i[29]_pad ,
		_w8655_,
		_w8656_,
		_w22984_
	);
	LUT4 #(
		.INIT('h67ef)
	) name21084 (
		_w8650_,
		_w8653_,
		_w22983_,
		_w22984_,
		_w22985_
	);
	LUT3 #(
		.INIT('h80)
	) name21085 (
		\m0_addr_i[29]_pad ,
		_w8655_,
		_w8656_,
		_w22986_
	);
	LUT3 #(
		.INIT('h2a)
	) name21086 (
		\m7_addr_i[29]_pad ,
		_w8655_,
		_w8656_,
		_w22987_
	);
	LUT4 #(
		.INIT('h6e7f)
	) name21087 (
		_w8650_,
		_w8653_,
		_w22986_,
		_w22987_,
		_w22988_
	);
	LUT4 #(
		.INIT('h7fff)
	) name21088 (
		_w22979_,
		_w22982_,
		_w22985_,
		_w22988_,
		_w22989_
	);
	LUT3 #(
		.INIT('h2a)
	) name21089 (
		\m3_addr_i[2]_pad ,
		_w8655_,
		_w8656_,
		_w22990_
	);
	LUT3 #(
		.INIT('h80)
	) name21090 (
		\m4_addr_i[2]_pad ,
		_w8655_,
		_w8656_,
		_w22991_
	);
	LUT4 #(
		.INIT('h9dbf)
	) name21091 (
		_w8650_,
		_w8653_,
		_w22990_,
		_w22991_,
		_w22992_
	);
	LUT3 #(
		.INIT('h80)
	) name21092 (
		\m6_addr_i[2]_pad ,
		_w8655_,
		_w8656_,
		_w22993_
	);
	LUT3 #(
		.INIT('h80)
	) name21093 (
		\m2_addr_i[2]_pad ,
		_w8655_,
		_w8656_,
		_w22994_
	);
	LUT4 #(
		.INIT('habef)
	) name21094 (
		_w8650_,
		_w8653_,
		_w22993_,
		_w22994_,
		_w22995_
	);
	LUT3 #(
		.INIT('h2a)
	) name21095 (
		\m5_addr_i[2]_pad ,
		_w8655_,
		_w8656_,
		_w22996_
	);
	LUT3 #(
		.INIT('h2a)
	) name21096 (
		\m1_addr_i[2]_pad ,
		_w8655_,
		_w8656_,
		_w22997_
	);
	LUT4 #(
		.INIT('h57df)
	) name21097 (
		_w8650_,
		_w8653_,
		_w22996_,
		_w22997_,
		_w22998_
	);
	LUT3 #(
		.INIT('h80)
	) name21098 (
		\m0_addr_i[2]_pad ,
		_w8655_,
		_w8656_,
		_w22999_
	);
	LUT3 #(
		.INIT('h2a)
	) name21099 (
		\m7_addr_i[2]_pad ,
		_w8655_,
		_w8656_,
		_w23000_
	);
	LUT4 #(
		.INIT('h6e7f)
	) name21100 (
		_w8650_,
		_w8653_,
		_w22999_,
		_w23000_,
		_w23001_
	);
	LUT4 #(
		.INIT('h7fff)
	) name21101 (
		_w22992_,
		_w22995_,
		_w22998_,
		_w23001_,
		_w23002_
	);
	LUT3 #(
		.INIT('h2a)
	) name21102 (
		\m3_addr_i[30]_pad ,
		_w8655_,
		_w8656_,
		_w23003_
	);
	LUT3 #(
		.INIT('h80)
	) name21103 (
		\m4_addr_i[30]_pad ,
		_w8655_,
		_w8656_,
		_w23004_
	);
	LUT4 #(
		.INIT('h9dbf)
	) name21104 (
		_w8650_,
		_w8653_,
		_w23003_,
		_w23004_,
		_w23005_
	);
	LUT3 #(
		.INIT('h2a)
	) name21105 (
		\m5_addr_i[30]_pad ,
		_w8655_,
		_w8656_,
		_w23006_
	);
	LUT3 #(
		.INIT('h80)
	) name21106 (
		\m2_addr_i[30]_pad ,
		_w8655_,
		_w8656_,
		_w23007_
	);
	LUT4 #(
		.INIT('h9bdf)
	) name21107 (
		_w8650_,
		_w8653_,
		_w23006_,
		_w23007_,
		_w23008_
	);
	LUT3 #(
		.INIT('h80)
	) name21108 (
		\m6_addr_i[30]_pad ,
		_w8655_,
		_w8656_,
		_w23009_
	);
	LUT3 #(
		.INIT('h2a)
	) name21109 (
		\m1_addr_i[30]_pad ,
		_w8655_,
		_w8656_,
		_w23010_
	);
	LUT4 #(
		.INIT('h67ef)
	) name21110 (
		_w8650_,
		_w8653_,
		_w23009_,
		_w23010_,
		_w23011_
	);
	LUT3 #(
		.INIT('h80)
	) name21111 (
		\m0_addr_i[30]_pad ,
		_w8655_,
		_w8656_,
		_w23012_
	);
	LUT3 #(
		.INIT('h2a)
	) name21112 (
		\m7_addr_i[30]_pad ,
		_w8655_,
		_w8656_,
		_w23013_
	);
	LUT4 #(
		.INIT('h6e7f)
	) name21113 (
		_w8650_,
		_w8653_,
		_w23012_,
		_w23013_,
		_w23014_
	);
	LUT4 #(
		.INIT('h7fff)
	) name21114 (
		_w23005_,
		_w23008_,
		_w23011_,
		_w23014_,
		_w23015_
	);
	LUT3 #(
		.INIT('h2a)
	) name21115 (
		\m3_addr_i[31]_pad ,
		_w8655_,
		_w8656_,
		_w23016_
	);
	LUT3 #(
		.INIT('h80)
	) name21116 (
		\m4_addr_i[31]_pad ,
		_w8655_,
		_w8656_,
		_w23017_
	);
	LUT4 #(
		.INIT('h9dbf)
	) name21117 (
		_w8650_,
		_w8653_,
		_w23016_,
		_w23017_,
		_w23018_
	);
	LUT3 #(
		.INIT('h2a)
	) name21118 (
		\m5_addr_i[31]_pad ,
		_w8655_,
		_w8656_,
		_w23019_
	);
	LUT3 #(
		.INIT('h80)
	) name21119 (
		\m2_addr_i[31]_pad ,
		_w8655_,
		_w8656_,
		_w23020_
	);
	LUT4 #(
		.INIT('h9bdf)
	) name21120 (
		_w8650_,
		_w8653_,
		_w23019_,
		_w23020_,
		_w23021_
	);
	LUT3 #(
		.INIT('h80)
	) name21121 (
		\m6_addr_i[31]_pad ,
		_w8655_,
		_w8656_,
		_w23022_
	);
	LUT3 #(
		.INIT('h2a)
	) name21122 (
		\m1_addr_i[31]_pad ,
		_w8655_,
		_w8656_,
		_w23023_
	);
	LUT4 #(
		.INIT('h67ef)
	) name21123 (
		_w8650_,
		_w8653_,
		_w23022_,
		_w23023_,
		_w23024_
	);
	LUT3 #(
		.INIT('h80)
	) name21124 (
		\m0_addr_i[31]_pad ,
		_w8655_,
		_w8656_,
		_w23025_
	);
	LUT3 #(
		.INIT('h2a)
	) name21125 (
		\m7_addr_i[31]_pad ,
		_w8655_,
		_w8656_,
		_w23026_
	);
	LUT4 #(
		.INIT('h6e7f)
	) name21126 (
		_w8650_,
		_w8653_,
		_w23025_,
		_w23026_,
		_w23027_
	);
	LUT4 #(
		.INIT('h7fff)
	) name21127 (
		_w23018_,
		_w23021_,
		_w23024_,
		_w23027_,
		_w23028_
	);
	LUT3 #(
		.INIT('h2a)
	) name21128 (
		\m3_addr_i[3]_pad ,
		_w8655_,
		_w8656_,
		_w23029_
	);
	LUT3 #(
		.INIT('h80)
	) name21129 (
		\m4_addr_i[3]_pad ,
		_w8655_,
		_w8656_,
		_w23030_
	);
	LUT4 #(
		.INIT('h9dbf)
	) name21130 (
		_w8650_,
		_w8653_,
		_w23029_,
		_w23030_,
		_w23031_
	);
	LUT3 #(
		.INIT('h80)
	) name21131 (
		\m6_addr_i[3]_pad ,
		_w8655_,
		_w8656_,
		_w23032_
	);
	LUT3 #(
		.INIT('h80)
	) name21132 (
		\m2_addr_i[3]_pad ,
		_w8655_,
		_w8656_,
		_w23033_
	);
	LUT4 #(
		.INIT('habef)
	) name21133 (
		_w8650_,
		_w8653_,
		_w23032_,
		_w23033_,
		_w23034_
	);
	LUT3 #(
		.INIT('h2a)
	) name21134 (
		\m5_addr_i[3]_pad ,
		_w8655_,
		_w8656_,
		_w23035_
	);
	LUT3 #(
		.INIT('h2a)
	) name21135 (
		\m1_addr_i[3]_pad ,
		_w8655_,
		_w8656_,
		_w23036_
	);
	LUT4 #(
		.INIT('h57df)
	) name21136 (
		_w8650_,
		_w8653_,
		_w23035_,
		_w23036_,
		_w23037_
	);
	LUT3 #(
		.INIT('h80)
	) name21137 (
		\m0_addr_i[3]_pad ,
		_w8655_,
		_w8656_,
		_w23038_
	);
	LUT3 #(
		.INIT('h2a)
	) name21138 (
		\m7_addr_i[3]_pad ,
		_w8655_,
		_w8656_,
		_w23039_
	);
	LUT4 #(
		.INIT('h6e7f)
	) name21139 (
		_w8650_,
		_w8653_,
		_w23038_,
		_w23039_,
		_w23040_
	);
	LUT4 #(
		.INIT('h7fff)
	) name21140 (
		_w23031_,
		_w23034_,
		_w23037_,
		_w23040_,
		_w23041_
	);
	LUT3 #(
		.INIT('h2a)
	) name21141 (
		\m3_addr_i[4]_pad ,
		_w8655_,
		_w8656_,
		_w23042_
	);
	LUT3 #(
		.INIT('h80)
	) name21142 (
		\m4_addr_i[4]_pad ,
		_w8655_,
		_w8656_,
		_w23043_
	);
	LUT4 #(
		.INIT('h9dbf)
	) name21143 (
		_w8650_,
		_w8653_,
		_w23042_,
		_w23043_,
		_w23044_
	);
	LUT3 #(
		.INIT('h80)
	) name21144 (
		\m6_addr_i[4]_pad ,
		_w8655_,
		_w8656_,
		_w23045_
	);
	LUT3 #(
		.INIT('h80)
	) name21145 (
		\m2_addr_i[4]_pad ,
		_w8655_,
		_w8656_,
		_w23046_
	);
	LUT4 #(
		.INIT('habef)
	) name21146 (
		_w8650_,
		_w8653_,
		_w23045_,
		_w23046_,
		_w23047_
	);
	LUT3 #(
		.INIT('h2a)
	) name21147 (
		\m5_addr_i[4]_pad ,
		_w8655_,
		_w8656_,
		_w23048_
	);
	LUT3 #(
		.INIT('h2a)
	) name21148 (
		\m1_addr_i[4]_pad ,
		_w8655_,
		_w8656_,
		_w23049_
	);
	LUT4 #(
		.INIT('h57df)
	) name21149 (
		_w8650_,
		_w8653_,
		_w23048_,
		_w23049_,
		_w23050_
	);
	LUT3 #(
		.INIT('h80)
	) name21150 (
		\m0_addr_i[4]_pad ,
		_w8655_,
		_w8656_,
		_w23051_
	);
	LUT3 #(
		.INIT('h2a)
	) name21151 (
		\m7_addr_i[4]_pad ,
		_w8655_,
		_w8656_,
		_w23052_
	);
	LUT4 #(
		.INIT('h6e7f)
	) name21152 (
		_w8650_,
		_w8653_,
		_w23051_,
		_w23052_,
		_w23053_
	);
	LUT4 #(
		.INIT('h7fff)
	) name21153 (
		_w23044_,
		_w23047_,
		_w23050_,
		_w23053_,
		_w23054_
	);
	LUT3 #(
		.INIT('h2a)
	) name21154 (
		\m3_addr_i[5]_pad ,
		_w8655_,
		_w8656_,
		_w23055_
	);
	LUT3 #(
		.INIT('h80)
	) name21155 (
		\m4_addr_i[5]_pad ,
		_w8655_,
		_w8656_,
		_w23056_
	);
	LUT4 #(
		.INIT('h9dbf)
	) name21156 (
		_w8650_,
		_w8653_,
		_w23055_,
		_w23056_,
		_w23057_
	);
	LUT3 #(
		.INIT('h80)
	) name21157 (
		\m6_addr_i[5]_pad ,
		_w8655_,
		_w8656_,
		_w23058_
	);
	LUT3 #(
		.INIT('h80)
	) name21158 (
		\m2_addr_i[5]_pad ,
		_w8655_,
		_w8656_,
		_w23059_
	);
	LUT4 #(
		.INIT('habef)
	) name21159 (
		_w8650_,
		_w8653_,
		_w23058_,
		_w23059_,
		_w23060_
	);
	LUT3 #(
		.INIT('h2a)
	) name21160 (
		\m5_addr_i[5]_pad ,
		_w8655_,
		_w8656_,
		_w23061_
	);
	LUT3 #(
		.INIT('h2a)
	) name21161 (
		\m1_addr_i[5]_pad ,
		_w8655_,
		_w8656_,
		_w23062_
	);
	LUT4 #(
		.INIT('h57df)
	) name21162 (
		_w8650_,
		_w8653_,
		_w23061_,
		_w23062_,
		_w23063_
	);
	LUT3 #(
		.INIT('h80)
	) name21163 (
		\m0_addr_i[5]_pad ,
		_w8655_,
		_w8656_,
		_w23064_
	);
	LUT3 #(
		.INIT('h2a)
	) name21164 (
		\m7_addr_i[5]_pad ,
		_w8655_,
		_w8656_,
		_w23065_
	);
	LUT4 #(
		.INIT('h6e7f)
	) name21165 (
		_w8650_,
		_w8653_,
		_w23064_,
		_w23065_,
		_w23066_
	);
	LUT4 #(
		.INIT('h7fff)
	) name21166 (
		_w23057_,
		_w23060_,
		_w23063_,
		_w23066_,
		_w23067_
	);
	LUT3 #(
		.INIT('h2a)
	) name21167 (
		\m3_addr_i[6]_pad ,
		_w8655_,
		_w8656_,
		_w23068_
	);
	LUT3 #(
		.INIT('h80)
	) name21168 (
		\m4_addr_i[6]_pad ,
		_w8655_,
		_w8656_,
		_w23069_
	);
	LUT4 #(
		.INIT('h9dbf)
	) name21169 (
		_w8650_,
		_w8653_,
		_w23068_,
		_w23069_,
		_w23070_
	);
	LUT3 #(
		.INIT('h80)
	) name21170 (
		\m6_addr_i[6]_pad ,
		_w8655_,
		_w8656_,
		_w23071_
	);
	LUT3 #(
		.INIT('h80)
	) name21171 (
		\m2_addr_i[6]_pad ,
		_w8655_,
		_w8656_,
		_w23072_
	);
	LUT4 #(
		.INIT('habef)
	) name21172 (
		_w8650_,
		_w8653_,
		_w23071_,
		_w23072_,
		_w23073_
	);
	LUT3 #(
		.INIT('h2a)
	) name21173 (
		\m5_addr_i[6]_pad ,
		_w8655_,
		_w8656_,
		_w23074_
	);
	LUT3 #(
		.INIT('h2a)
	) name21174 (
		\m1_addr_i[6]_pad ,
		_w8655_,
		_w8656_,
		_w23075_
	);
	LUT4 #(
		.INIT('h57df)
	) name21175 (
		_w8650_,
		_w8653_,
		_w23074_,
		_w23075_,
		_w23076_
	);
	LUT3 #(
		.INIT('h80)
	) name21176 (
		\m0_addr_i[6]_pad ,
		_w8655_,
		_w8656_,
		_w23077_
	);
	LUT3 #(
		.INIT('h2a)
	) name21177 (
		\m7_addr_i[6]_pad ,
		_w8655_,
		_w8656_,
		_w23078_
	);
	LUT4 #(
		.INIT('h6e7f)
	) name21178 (
		_w8650_,
		_w8653_,
		_w23077_,
		_w23078_,
		_w23079_
	);
	LUT4 #(
		.INIT('h7fff)
	) name21179 (
		_w23070_,
		_w23073_,
		_w23076_,
		_w23079_,
		_w23080_
	);
	LUT3 #(
		.INIT('h2a)
	) name21180 (
		\m3_addr_i[7]_pad ,
		_w8655_,
		_w8656_,
		_w23081_
	);
	LUT3 #(
		.INIT('h80)
	) name21181 (
		\m4_addr_i[7]_pad ,
		_w8655_,
		_w8656_,
		_w23082_
	);
	LUT4 #(
		.INIT('h9dbf)
	) name21182 (
		_w8650_,
		_w8653_,
		_w23081_,
		_w23082_,
		_w23083_
	);
	LUT3 #(
		.INIT('h80)
	) name21183 (
		\m6_addr_i[7]_pad ,
		_w8655_,
		_w8656_,
		_w23084_
	);
	LUT3 #(
		.INIT('h80)
	) name21184 (
		\m2_addr_i[7]_pad ,
		_w8655_,
		_w8656_,
		_w23085_
	);
	LUT4 #(
		.INIT('habef)
	) name21185 (
		_w8650_,
		_w8653_,
		_w23084_,
		_w23085_,
		_w23086_
	);
	LUT3 #(
		.INIT('h2a)
	) name21186 (
		\m5_addr_i[7]_pad ,
		_w8655_,
		_w8656_,
		_w23087_
	);
	LUT3 #(
		.INIT('h2a)
	) name21187 (
		\m1_addr_i[7]_pad ,
		_w8655_,
		_w8656_,
		_w23088_
	);
	LUT4 #(
		.INIT('h57df)
	) name21188 (
		_w8650_,
		_w8653_,
		_w23087_,
		_w23088_,
		_w23089_
	);
	LUT3 #(
		.INIT('h80)
	) name21189 (
		\m0_addr_i[7]_pad ,
		_w8655_,
		_w8656_,
		_w23090_
	);
	LUT3 #(
		.INIT('h2a)
	) name21190 (
		\m7_addr_i[7]_pad ,
		_w8655_,
		_w8656_,
		_w23091_
	);
	LUT4 #(
		.INIT('h6e7f)
	) name21191 (
		_w8650_,
		_w8653_,
		_w23090_,
		_w23091_,
		_w23092_
	);
	LUT4 #(
		.INIT('h7fff)
	) name21192 (
		_w23083_,
		_w23086_,
		_w23089_,
		_w23092_,
		_w23093_
	);
	LUT3 #(
		.INIT('h2a)
	) name21193 (
		\m3_addr_i[8]_pad ,
		_w8655_,
		_w8656_,
		_w23094_
	);
	LUT3 #(
		.INIT('h80)
	) name21194 (
		\m4_addr_i[8]_pad ,
		_w8655_,
		_w8656_,
		_w23095_
	);
	LUT4 #(
		.INIT('h9dbf)
	) name21195 (
		_w8650_,
		_w8653_,
		_w23094_,
		_w23095_,
		_w23096_
	);
	LUT3 #(
		.INIT('h80)
	) name21196 (
		\m6_addr_i[8]_pad ,
		_w8655_,
		_w8656_,
		_w23097_
	);
	LUT3 #(
		.INIT('h80)
	) name21197 (
		\m2_addr_i[8]_pad ,
		_w8655_,
		_w8656_,
		_w23098_
	);
	LUT4 #(
		.INIT('habef)
	) name21198 (
		_w8650_,
		_w8653_,
		_w23097_,
		_w23098_,
		_w23099_
	);
	LUT3 #(
		.INIT('h2a)
	) name21199 (
		\m5_addr_i[8]_pad ,
		_w8655_,
		_w8656_,
		_w23100_
	);
	LUT3 #(
		.INIT('h2a)
	) name21200 (
		\m1_addr_i[8]_pad ,
		_w8655_,
		_w8656_,
		_w23101_
	);
	LUT4 #(
		.INIT('h57df)
	) name21201 (
		_w8650_,
		_w8653_,
		_w23100_,
		_w23101_,
		_w23102_
	);
	LUT3 #(
		.INIT('h80)
	) name21202 (
		\m0_addr_i[8]_pad ,
		_w8655_,
		_w8656_,
		_w23103_
	);
	LUT3 #(
		.INIT('h2a)
	) name21203 (
		\m7_addr_i[8]_pad ,
		_w8655_,
		_w8656_,
		_w23104_
	);
	LUT4 #(
		.INIT('h6e7f)
	) name21204 (
		_w8650_,
		_w8653_,
		_w23103_,
		_w23104_,
		_w23105_
	);
	LUT4 #(
		.INIT('h7fff)
	) name21205 (
		_w23096_,
		_w23099_,
		_w23102_,
		_w23105_,
		_w23106_
	);
	LUT3 #(
		.INIT('h2a)
	) name21206 (
		\m3_addr_i[9]_pad ,
		_w8655_,
		_w8656_,
		_w23107_
	);
	LUT3 #(
		.INIT('h80)
	) name21207 (
		\m4_addr_i[9]_pad ,
		_w8655_,
		_w8656_,
		_w23108_
	);
	LUT4 #(
		.INIT('h9dbf)
	) name21208 (
		_w8650_,
		_w8653_,
		_w23107_,
		_w23108_,
		_w23109_
	);
	LUT3 #(
		.INIT('h80)
	) name21209 (
		\m6_addr_i[9]_pad ,
		_w8655_,
		_w8656_,
		_w23110_
	);
	LUT3 #(
		.INIT('h80)
	) name21210 (
		\m2_addr_i[9]_pad ,
		_w8655_,
		_w8656_,
		_w23111_
	);
	LUT4 #(
		.INIT('habef)
	) name21211 (
		_w8650_,
		_w8653_,
		_w23110_,
		_w23111_,
		_w23112_
	);
	LUT3 #(
		.INIT('h2a)
	) name21212 (
		\m5_addr_i[9]_pad ,
		_w8655_,
		_w8656_,
		_w23113_
	);
	LUT3 #(
		.INIT('h2a)
	) name21213 (
		\m1_addr_i[9]_pad ,
		_w8655_,
		_w8656_,
		_w23114_
	);
	LUT4 #(
		.INIT('h57df)
	) name21214 (
		_w8650_,
		_w8653_,
		_w23113_,
		_w23114_,
		_w23115_
	);
	LUT3 #(
		.INIT('h80)
	) name21215 (
		\m0_addr_i[9]_pad ,
		_w8655_,
		_w8656_,
		_w23116_
	);
	LUT3 #(
		.INIT('h2a)
	) name21216 (
		\m7_addr_i[9]_pad ,
		_w8655_,
		_w8656_,
		_w23117_
	);
	LUT4 #(
		.INIT('h6e7f)
	) name21217 (
		_w8650_,
		_w8653_,
		_w23116_,
		_w23117_,
		_w23118_
	);
	LUT4 #(
		.INIT('h7fff)
	) name21218 (
		_w23109_,
		_w23112_,
		_w23115_,
		_w23118_,
		_w23119_
	);
	LUT3 #(
		.INIT('h2a)
	) name21219 (
		\m3_data_i[0]_pad ,
		_w8655_,
		_w8656_,
		_w23120_
	);
	LUT3 #(
		.INIT('h80)
	) name21220 (
		\m4_data_i[0]_pad ,
		_w8655_,
		_w8656_,
		_w23121_
	);
	LUT4 #(
		.INIT('h9dbf)
	) name21221 (
		_w8650_,
		_w8653_,
		_w23120_,
		_w23121_,
		_w23122_
	);
	LUT3 #(
		.INIT('h80)
	) name21222 (
		\m6_data_i[0]_pad ,
		_w8655_,
		_w8656_,
		_w23123_
	);
	LUT3 #(
		.INIT('h80)
	) name21223 (
		\m2_data_i[0]_pad ,
		_w8655_,
		_w8656_,
		_w23124_
	);
	LUT4 #(
		.INIT('habef)
	) name21224 (
		_w8650_,
		_w8653_,
		_w23123_,
		_w23124_,
		_w23125_
	);
	LUT3 #(
		.INIT('h2a)
	) name21225 (
		\m5_data_i[0]_pad ,
		_w8655_,
		_w8656_,
		_w23126_
	);
	LUT3 #(
		.INIT('h2a)
	) name21226 (
		\m1_data_i[0]_pad ,
		_w8655_,
		_w8656_,
		_w23127_
	);
	LUT4 #(
		.INIT('h57df)
	) name21227 (
		_w8650_,
		_w8653_,
		_w23126_,
		_w23127_,
		_w23128_
	);
	LUT3 #(
		.INIT('h80)
	) name21228 (
		\m0_data_i[0]_pad ,
		_w8655_,
		_w8656_,
		_w23129_
	);
	LUT3 #(
		.INIT('h2a)
	) name21229 (
		\m7_data_i[0]_pad ,
		_w8655_,
		_w8656_,
		_w23130_
	);
	LUT4 #(
		.INIT('h6e7f)
	) name21230 (
		_w8650_,
		_w8653_,
		_w23129_,
		_w23130_,
		_w23131_
	);
	LUT4 #(
		.INIT('h7fff)
	) name21231 (
		_w23122_,
		_w23125_,
		_w23128_,
		_w23131_,
		_w23132_
	);
	LUT3 #(
		.INIT('h2a)
	) name21232 (
		\m3_data_i[10]_pad ,
		_w8655_,
		_w8656_,
		_w23133_
	);
	LUT3 #(
		.INIT('h80)
	) name21233 (
		\m4_data_i[10]_pad ,
		_w8655_,
		_w8656_,
		_w23134_
	);
	LUT4 #(
		.INIT('h9dbf)
	) name21234 (
		_w8650_,
		_w8653_,
		_w23133_,
		_w23134_,
		_w23135_
	);
	LUT3 #(
		.INIT('h80)
	) name21235 (
		\m6_data_i[10]_pad ,
		_w8655_,
		_w8656_,
		_w23136_
	);
	LUT3 #(
		.INIT('h80)
	) name21236 (
		\m2_data_i[10]_pad ,
		_w8655_,
		_w8656_,
		_w23137_
	);
	LUT4 #(
		.INIT('habef)
	) name21237 (
		_w8650_,
		_w8653_,
		_w23136_,
		_w23137_,
		_w23138_
	);
	LUT3 #(
		.INIT('h2a)
	) name21238 (
		\m5_data_i[10]_pad ,
		_w8655_,
		_w8656_,
		_w23139_
	);
	LUT3 #(
		.INIT('h2a)
	) name21239 (
		\m1_data_i[10]_pad ,
		_w8655_,
		_w8656_,
		_w23140_
	);
	LUT4 #(
		.INIT('h57df)
	) name21240 (
		_w8650_,
		_w8653_,
		_w23139_,
		_w23140_,
		_w23141_
	);
	LUT3 #(
		.INIT('h80)
	) name21241 (
		\m0_data_i[10]_pad ,
		_w8655_,
		_w8656_,
		_w23142_
	);
	LUT3 #(
		.INIT('h2a)
	) name21242 (
		\m7_data_i[10]_pad ,
		_w8655_,
		_w8656_,
		_w23143_
	);
	LUT4 #(
		.INIT('h6e7f)
	) name21243 (
		_w8650_,
		_w8653_,
		_w23142_,
		_w23143_,
		_w23144_
	);
	LUT4 #(
		.INIT('h7fff)
	) name21244 (
		_w23135_,
		_w23138_,
		_w23141_,
		_w23144_,
		_w23145_
	);
	LUT3 #(
		.INIT('h2a)
	) name21245 (
		\m3_data_i[11]_pad ,
		_w8655_,
		_w8656_,
		_w23146_
	);
	LUT3 #(
		.INIT('h80)
	) name21246 (
		\m4_data_i[11]_pad ,
		_w8655_,
		_w8656_,
		_w23147_
	);
	LUT4 #(
		.INIT('h9dbf)
	) name21247 (
		_w8650_,
		_w8653_,
		_w23146_,
		_w23147_,
		_w23148_
	);
	LUT3 #(
		.INIT('h80)
	) name21248 (
		\m6_data_i[11]_pad ,
		_w8655_,
		_w8656_,
		_w23149_
	);
	LUT3 #(
		.INIT('h80)
	) name21249 (
		\m2_data_i[11]_pad ,
		_w8655_,
		_w8656_,
		_w23150_
	);
	LUT4 #(
		.INIT('habef)
	) name21250 (
		_w8650_,
		_w8653_,
		_w23149_,
		_w23150_,
		_w23151_
	);
	LUT3 #(
		.INIT('h2a)
	) name21251 (
		\m5_data_i[11]_pad ,
		_w8655_,
		_w8656_,
		_w23152_
	);
	LUT3 #(
		.INIT('h2a)
	) name21252 (
		\m1_data_i[11]_pad ,
		_w8655_,
		_w8656_,
		_w23153_
	);
	LUT4 #(
		.INIT('h57df)
	) name21253 (
		_w8650_,
		_w8653_,
		_w23152_,
		_w23153_,
		_w23154_
	);
	LUT3 #(
		.INIT('h80)
	) name21254 (
		\m0_data_i[11]_pad ,
		_w8655_,
		_w8656_,
		_w23155_
	);
	LUT3 #(
		.INIT('h2a)
	) name21255 (
		\m7_data_i[11]_pad ,
		_w8655_,
		_w8656_,
		_w23156_
	);
	LUT4 #(
		.INIT('h6e7f)
	) name21256 (
		_w8650_,
		_w8653_,
		_w23155_,
		_w23156_,
		_w23157_
	);
	LUT4 #(
		.INIT('h7fff)
	) name21257 (
		_w23148_,
		_w23151_,
		_w23154_,
		_w23157_,
		_w23158_
	);
	LUT3 #(
		.INIT('h2a)
	) name21258 (
		\m3_data_i[12]_pad ,
		_w8655_,
		_w8656_,
		_w23159_
	);
	LUT3 #(
		.INIT('h80)
	) name21259 (
		\m4_data_i[12]_pad ,
		_w8655_,
		_w8656_,
		_w23160_
	);
	LUT4 #(
		.INIT('h9dbf)
	) name21260 (
		_w8650_,
		_w8653_,
		_w23159_,
		_w23160_,
		_w23161_
	);
	LUT3 #(
		.INIT('h80)
	) name21261 (
		\m6_data_i[12]_pad ,
		_w8655_,
		_w8656_,
		_w23162_
	);
	LUT3 #(
		.INIT('h80)
	) name21262 (
		\m2_data_i[12]_pad ,
		_w8655_,
		_w8656_,
		_w23163_
	);
	LUT4 #(
		.INIT('habef)
	) name21263 (
		_w8650_,
		_w8653_,
		_w23162_,
		_w23163_,
		_w23164_
	);
	LUT3 #(
		.INIT('h2a)
	) name21264 (
		\m5_data_i[12]_pad ,
		_w8655_,
		_w8656_,
		_w23165_
	);
	LUT3 #(
		.INIT('h2a)
	) name21265 (
		\m1_data_i[12]_pad ,
		_w8655_,
		_w8656_,
		_w23166_
	);
	LUT4 #(
		.INIT('h57df)
	) name21266 (
		_w8650_,
		_w8653_,
		_w23165_,
		_w23166_,
		_w23167_
	);
	LUT3 #(
		.INIT('h80)
	) name21267 (
		\m0_data_i[12]_pad ,
		_w8655_,
		_w8656_,
		_w23168_
	);
	LUT3 #(
		.INIT('h2a)
	) name21268 (
		\m7_data_i[12]_pad ,
		_w8655_,
		_w8656_,
		_w23169_
	);
	LUT4 #(
		.INIT('h6e7f)
	) name21269 (
		_w8650_,
		_w8653_,
		_w23168_,
		_w23169_,
		_w23170_
	);
	LUT4 #(
		.INIT('h7fff)
	) name21270 (
		_w23161_,
		_w23164_,
		_w23167_,
		_w23170_,
		_w23171_
	);
	LUT3 #(
		.INIT('h2a)
	) name21271 (
		\m3_data_i[13]_pad ,
		_w8655_,
		_w8656_,
		_w23172_
	);
	LUT3 #(
		.INIT('h80)
	) name21272 (
		\m4_data_i[13]_pad ,
		_w8655_,
		_w8656_,
		_w23173_
	);
	LUT4 #(
		.INIT('h9dbf)
	) name21273 (
		_w8650_,
		_w8653_,
		_w23172_,
		_w23173_,
		_w23174_
	);
	LUT3 #(
		.INIT('h80)
	) name21274 (
		\m6_data_i[13]_pad ,
		_w8655_,
		_w8656_,
		_w23175_
	);
	LUT3 #(
		.INIT('h80)
	) name21275 (
		\m2_data_i[13]_pad ,
		_w8655_,
		_w8656_,
		_w23176_
	);
	LUT4 #(
		.INIT('habef)
	) name21276 (
		_w8650_,
		_w8653_,
		_w23175_,
		_w23176_,
		_w23177_
	);
	LUT3 #(
		.INIT('h2a)
	) name21277 (
		\m5_data_i[13]_pad ,
		_w8655_,
		_w8656_,
		_w23178_
	);
	LUT3 #(
		.INIT('h2a)
	) name21278 (
		\m1_data_i[13]_pad ,
		_w8655_,
		_w8656_,
		_w23179_
	);
	LUT4 #(
		.INIT('h57df)
	) name21279 (
		_w8650_,
		_w8653_,
		_w23178_,
		_w23179_,
		_w23180_
	);
	LUT3 #(
		.INIT('h80)
	) name21280 (
		\m0_data_i[13]_pad ,
		_w8655_,
		_w8656_,
		_w23181_
	);
	LUT3 #(
		.INIT('h2a)
	) name21281 (
		\m7_data_i[13]_pad ,
		_w8655_,
		_w8656_,
		_w23182_
	);
	LUT4 #(
		.INIT('h6e7f)
	) name21282 (
		_w8650_,
		_w8653_,
		_w23181_,
		_w23182_,
		_w23183_
	);
	LUT4 #(
		.INIT('h7fff)
	) name21283 (
		_w23174_,
		_w23177_,
		_w23180_,
		_w23183_,
		_w23184_
	);
	LUT3 #(
		.INIT('h2a)
	) name21284 (
		\m3_data_i[14]_pad ,
		_w8655_,
		_w8656_,
		_w23185_
	);
	LUT3 #(
		.INIT('h80)
	) name21285 (
		\m4_data_i[14]_pad ,
		_w8655_,
		_w8656_,
		_w23186_
	);
	LUT4 #(
		.INIT('h9dbf)
	) name21286 (
		_w8650_,
		_w8653_,
		_w23185_,
		_w23186_,
		_w23187_
	);
	LUT3 #(
		.INIT('h80)
	) name21287 (
		\m6_data_i[14]_pad ,
		_w8655_,
		_w8656_,
		_w23188_
	);
	LUT3 #(
		.INIT('h80)
	) name21288 (
		\m2_data_i[14]_pad ,
		_w8655_,
		_w8656_,
		_w23189_
	);
	LUT4 #(
		.INIT('habef)
	) name21289 (
		_w8650_,
		_w8653_,
		_w23188_,
		_w23189_,
		_w23190_
	);
	LUT3 #(
		.INIT('h2a)
	) name21290 (
		\m5_data_i[14]_pad ,
		_w8655_,
		_w8656_,
		_w23191_
	);
	LUT3 #(
		.INIT('h2a)
	) name21291 (
		\m1_data_i[14]_pad ,
		_w8655_,
		_w8656_,
		_w23192_
	);
	LUT4 #(
		.INIT('h57df)
	) name21292 (
		_w8650_,
		_w8653_,
		_w23191_,
		_w23192_,
		_w23193_
	);
	LUT3 #(
		.INIT('h80)
	) name21293 (
		\m0_data_i[14]_pad ,
		_w8655_,
		_w8656_,
		_w23194_
	);
	LUT3 #(
		.INIT('h2a)
	) name21294 (
		\m7_data_i[14]_pad ,
		_w8655_,
		_w8656_,
		_w23195_
	);
	LUT4 #(
		.INIT('h6e7f)
	) name21295 (
		_w8650_,
		_w8653_,
		_w23194_,
		_w23195_,
		_w23196_
	);
	LUT4 #(
		.INIT('h7fff)
	) name21296 (
		_w23187_,
		_w23190_,
		_w23193_,
		_w23196_,
		_w23197_
	);
	LUT3 #(
		.INIT('h2a)
	) name21297 (
		\m3_data_i[15]_pad ,
		_w8655_,
		_w8656_,
		_w23198_
	);
	LUT3 #(
		.INIT('h80)
	) name21298 (
		\m4_data_i[15]_pad ,
		_w8655_,
		_w8656_,
		_w23199_
	);
	LUT4 #(
		.INIT('h9dbf)
	) name21299 (
		_w8650_,
		_w8653_,
		_w23198_,
		_w23199_,
		_w23200_
	);
	LUT3 #(
		.INIT('h80)
	) name21300 (
		\m6_data_i[15]_pad ,
		_w8655_,
		_w8656_,
		_w23201_
	);
	LUT3 #(
		.INIT('h80)
	) name21301 (
		\m2_data_i[15]_pad ,
		_w8655_,
		_w8656_,
		_w23202_
	);
	LUT4 #(
		.INIT('habef)
	) name21302 (
		_w8650_,
		_w8653_,
		_w23201_,
		_w23202_,
		_w23203_
	);
	LUT3 #(
		.INIT('h2a)
	) name21303 (
		\m5_data_i[15]_pad ,
		_w8655_,
		_w8656_,
		_w23204_
	);
	LUT3 #(
		.INIT('h2a)
	) name21304 (
		\m1_data_i[15]_pad ,
		_w8655_,
		_w8656_,
		_w23205_
	);
	LUT4 #(
		.INIT('h57df)
	) name21305 (
		_w8650_,
		_w8653_,
		_w23204_,
		_w23205_,
		_w23206_
	);
	LUT3 #(
		.INIT('h80)
	) name21306 (
		\m0_data_i[15]_pad ,
		_w8655_,
		_w8656_,
		_w23207_
	);
	LUT3 #(
		.INIT('h2a)
	) name21307 (
		\m7_data_i[15]_pad ,
		_w8655_,
		_w8656_,
		_w23208_
	);
	LUT4 #(
		.INIT('h6e7f)
	) name21308 (
		_w8650_,
		_w8653_,
		_w23207_,
		_w23208_,
		_w23209_
	);
	LUT4 #(
		.INIT('h7fff)
	) name21309 (
		_w23200_,
		_w23203_,
		_w23206_,
		_w23209_,
		_w23210_
	);
	LUT3 #(
		.INIT('h2a)
	) name21310 (
		\m3_data_i[16]_pad ,
		_w8655_,
		_w8656_,
		_w23211_
	);
	LUT3 #(
		.INIT('h80)
	) name21311 (
		\m4_data_i[16]_pad ,
		_w8655_,
		_w8656_,
		_w23212_
	);
	LUT4 #(
		.INIT('h9dbf)
	) name21312 (
		_w8650_,
		_w8653_,
		_w23211_,
		_w23212_,
		_w23213_
	);
	LUT3 #(
		.INIT('h80)
	) name21313 (
		\m6_data_i[16]_pad ,
		_w8655_,
		_w8656_,
		_w23214_
	);
	LUT3 #(
		.INIT('h80)
	) name21314 (
		\m2_data_i[16]_pad ,
		_w8655_,
		_w8656_,
		_w23215_
	);
	LUT4 #(
		.INIT('habef)
	) name21315 (
		_w8650_,
		_w8653_,
		_w23214_,
		_w23215_,
		_w23216_
	);
	LUT3 #(
		.INIT('h2a)
	) name21316 (
		\m5_data_i[16]_pad ,
		_w8655_,
		_w8656_,
		_w23217_
	);
	LUT3 #(
		.INIT('h2a)
	) name21317 (
		\m1_data_i[16]_pad ,
		_w8655_,
		_w8656_,
		_w23218_
	);
	LUT4 #(
		.INIT('h57df)
	) name21318 (
		_w8650_,
		_w8653_,
		_w23217_,
		_w23218_,
		_w23219_
	);
	LUT3 #(
		.INIT('h80)
	) name21319 (
		\m0_data_i[16]_pad ,
		_w8655_,
		_w8656_,
		_w23220_
	);
	LUT3 #(
		.INIT('h2a)
	) name21320 (
		\m7_data_i[16]_pad ,
		_w8655_,
		_w8656_,
		_w23221_
	);
	LUT4 #(
		.INIT('h6e7f)
	) name21321 (
		_w8650_,
		_w8653_,
		_w23220_,
		_w23221_,
		_w23222_
	);
	LUT4 #(
		.INIT('h7fff)
	) name21322 (
		_w23213_,
		_w23216_,
		_w23219_,
		_w23222_,
		_w23223_
	);
	LUT3 #(
		.INIT('h2a)
	) name21323 (
		\m3_data_i[17]_pad ,
		_w8655_,
		_w8656_,
		_w23224_
	);
	LUT3 #(
		.INIT('h80)
	) name21324 (
		\m4_data_i[17]_pad ,
		_w8655_,
		_w8656_,
		_w23225_
	);
	LUT4 #(
		.INIT('h9dbf)
	) name21325 (
		_w8650_,
		_w8653_,
		_w23224_,
		_w23225_,
		_w23226_
	);
	LUT3 #(
		.INIT('h80)
	) name21326 (
		\m6_data_i[17]_pad ,
		_w8655_,
		_w8656_,
		_w23227_
	);
	LUT3 #(
		.INIT('h80)
	) name21327 (
		\m2_data_i[17]_pad ,
		_w8655_,
		_w8656_,
		_w23228_
	);
	LUT4 #(
		.INIT('habef)
	) name21328 (
		_w8650_,
		_w8653_,
		_w23227_,
		_w23228_,
		_w23229_
	);
	LUT3 #(
		.INIT('h2a)
	) name21329 (
		\m5_data_i[17]_pad ,
		_w8655_,
		_w8656_,
		_w23230_
	);
	LUT3 #(
		.INIT('h2a)
	) name21330 (
		\m1_data_i[17]_pad ,
		_w8655_,
		_w8656_,
		_w23231_
	);
	LUT4 #(
		.INIT('h57df)
	) name21331 (
		_w8650_,
		_w8653_,
		_w23230_,
		_w23231_,
		_w23232_
	);
	LUT3 #(
		.INIT('h80)
	) name21332 (
		\m0_data_i[17]_pad ,
		_w8655_,
		_w8656_,
		_w23233_
	);
	LUT3 #(
		.INIT('h2a)
	) name21333 (
		\m7_data_i[17]_pad ,
		_w8655_,
		_w8656_,
		_w23234_
	);
	LUT4 #(
		.INIT('h6e7f)
	) name21334 (
		_w8650_,
		_w8653_,
		_w23233_,
		_w23234_,
		_w23235_
	);
	LUT4 #(
		.INIT('h7fff)
	) name21335 (
		_w23226_,
		_w23229_,
		_w23232_,
		_w23235_,
		_w23236_
	);
	LUT3 #(
		.INIT('h2a)
	) name21336 (
		\m3_data_i[18]_pad ,
		_w8655_,
		_w8656_,
		_w23237_
	);
	LUT3 #(
		.INIT('h80)
	) name21337 (
		\m4_data_i[18]_pad ,
		_w8655_,
		_w8656_,
		_w23238_
	);
	LUT4 #(
		.INIT('h9dbf)
	) name21338 (
		_w8650_,
		_w8653_,
		_w23237_,
		_w23238_,
		_w23239_
	);
	LUT3 #(
		.INIT('h80)
	) name21339 (
		\m6_data_i[18]_pad ,
		_w8655_,
		_w8656_,
		_w23240_
	);
	LUT3 #(
		.INIT('h80)
	) name21340 (
		\m2_data_i[18]_pad ,
		_w8655_,
		_w8656_,
		_w23241_
	);
	LUT4 #(
		.INIT('habef)
	) name21341 (
		_w8650_,
		_w8653_,
		_w23240_,
		_w23241_,
		_w23242_
	);
	LUT3 #(
		.INIT('h2a)
	) name21342 (
		\m5_data_i[18]_pad ,
		_w8655_,
		_w8656_,
		_w23243_
	);
	LUT3 #(
		.INIT('h2a)
	) name21343 (
		\m1_data_i[18]_pad ,
		_w8655_,
		_w8656_,
		_w23244_
	);
	LUT4 #(
		.INIT('h57df)
	) name21344 (
		_w8650_,
		_w8653_,
		_w23243_,
		_w23244_,
		_w23245_
	);
	LUT3 #(
		.INIT('h80)
	) name21345 (
		\m0_data_i[18]_pad ,
		_w8655_,
		_w8656_,
		_w23246_
	);
	LUT3 #(
		.INIT('h2a)
	) name21346 (
		\m7_data_i[18]_pad ,
		_w8655_,
		_w8656_,
		_w23247_
	);
	LUT4 #(
		.INIT('h6e7f)
	) name21347 (
		_w8650_,
		_w8653_,
		_w23246_,
		_w23247_,
		_w23248_
	);
	LUT4 #(
		.INIT('h7fff)
	) name21348 (
		_w23239_,
		_w23242_,
		_w23245_,
		_w23248_,
		_w23249_
	);
	LUT3 #(
		.INIT('h2a)
	) name21349 (
		\m3_data_i[19]_pad ,
		_w8655_,
		_w8656_,
		_w23250_
	);
	LUT3 #(
		.INIT('h80)
	) name21350 (
		\m4_data_i[19]_pad ,
		_w8655_,
		_w8656_,
		_w23251_
	);
	LUT4 #(
		.INIT('h9dbf)
	) name21351 (
		_w8650_,
		_w8653_,
		_w23250_,
		_w23251_,
		_w23252_
	);
	LUT3 #(
		.INIT('h80)
	) name21352 (
		\m6_data_i[19]_pad ,
		_w8655_,
		_w8656_,
		_w23253_
	);
	LUT3 #(
		.INIT('h80)
	) name21353 (
		\m2_data_i[19]_pad ,
		_w8655_,
		_w8656_,
		_w23254_
	);
	LUT4 #(
		.INIT('habef)
	) name21354 (
		_w8650_,
		_w8653_,
		_w23253_,
		_w23254_,
		_w23255_
	);
	LUT3 #(
		.INIT('h2a)
	) name21355 (
		\m5_data_i[19]_pad ,
		_w8655_,
		_w8656_,
		_w23256_
	);
	LUT3 #(
		.INIT('h2a)
	) name21356 (
		\m1_data_i[19]_pad ,
		_w8655_,
		_w8656_,
		_w23257_
	);
	LUT4 #(
		.INIT('h57df)
	) name21357 (
		_w8650_,
		_w8653_,
		_w23256_,
		_w23257_,
		_w23258_
	);
	LUT3 #(
		.INIT('h80)
	) name21358 (
		\m0_data_i[19]_pad ,
		_w8655_,
		_w8656_,
		_w23259_
	);
	LUT3 #(
		.INIT('h2a)
	) name21359 (
		\m7_data_i[19]_pad ,
		_w8655_,
		_w8656_,
		_w23260_
	);
	LUT4 #(
		.INIT('h6e7f)
	) name21360 (
		_w8650_,
		_w8653_,
		_w23259_,
		_w23260_,
		_w23261_
	);
	LUT4 #(
		.INIT('h7fff)
	) name21361 (
		_w23252_,
		_w23255_,
		_w23258_,
		_w23261_,
		_w23262_
	);
	LUT3 #(
		.INIT('h2a)
	) name21362 (
		\m3_data_i[1]_pad ,
		_w8655_,
		_w8656_,
		_w23263_
	);
	LUT3 #(
		.INIT('h80)
	) name21363 (
		\m4_data_i[1]_pad ,
		_w8655_,
		_w8656_,
		_w23264_
	);
	LUT4 #(
		.INIT('h9dbf)
	) name21364 (
		_w8650_,
		_w8653_,
		_w23263_,
		_w23264_,
		_w23265_
	);
	LUT3 #(
		.INIT('h80)
	) name21365 (
		\m6_data_i[1]_pad ,
		_w8655_,
		_w8656_,
		_w23266_
	);
	LUT3 #(
		.INIT('h80)
	) name21366 (
		\m2_data_i[1]_pad ,
		_w8655_,
		_w8656_,
		_w23267_
	);
	LUT4 #(
		.INIT('habef)
	) name21367 (
		_w8650_,
		_w8653_,
		_w23266_,
		_w23267_,
		_w23268_
	);
	LUT3 #(
		.INIT('h2a)
	) name21368 (
		\m5_data_i[1]_pad ,
		_w8655_,
		_w8656_,
		_w23269_
	);
	LUT3 #(
		.INIT('h2a)
	) name21369 (
		\m1_data_i[1]_pad ,
		_w8655_,
		_w8656_,
		_w23270_
	);
	LUT4 #(
		.INIT('h57df)
	) name21370 (
		_w8650_,
		_w8653_,
		_w23269_,
		_w23270_,
		_w23271_
	);
	LUT3 #(
		.INIT('h80)
	) name21371 (
		\m0_data_i[1]_pad ,
		_w8655_,
		_w8656_,
		_w23272_
	);
	LUT3 #(
		.INIT('h2a)
	) name21372 (
		\m7_data_i[1]_pad ,
		_w8655_,
		_w8656_,
		_w23273_
	);
	LUT4 #(
		.INIT('h6e7f)
	) name21373 (
		_w8650_,
		_w8653_,
		_w23272_,
		_w23273_,
		_w23274_
	);
	LUT4 #(
		.INIT('h7fff)
	) name21374 (
		_w23265_,
		_w23268_,
		_w23271_,
		_w23274_,
		_w23275_
	);
	LUT3 #(
		.INIT('h2a)
	) name21375 (
		\m3_data_i[20]_pad ,
		_w8655_,
		_w8656_,
		_w23276_
	);
	LUT3 #(
		.INIT('h80)
	) name21376 (
		\m4_data_i[20]_pad ,
		_w8655_,
		_w8656_,
		_w23277_
	);
	LUT4 #(
		.INIT('h9dbf)
	) name21377 (
		_w8650_,
		_w8653_,
		_w23276_,
		_w23277_,
		_w23278_
	);
	LUT3 #(
		.INIT('h80)
	) name21378 (
		\m6_data_i[20]_pad ,
		_w8655_,
		_w8656_,
		_w23279_
	);
	LUT3 #(
		.INIT('h80)
	) name21379 (
		\m2_data_i[20]_pad ,
		_w8655_,
		_w8656_,
		_w23280_
	);
	LUT4 #(
		.INIT('habef)
	) name21380 (
		_w8650_,
		_w8653_,
		_w23279_,
		_w23280_,
		_w23281_
	);
	LUT3 #(
		.INIT('h2a)
	) name21381 (
		\m5_data_i[20]_pad ,
		_w8655_,
		_w8656_,
		_w23282_
	);
	LUT3 #(
		.INIT('h2a)
	) name21382 (
		\m1_data_i[20]_pad ,
		_w8655_,
		_w8656_,
		_w23283_
	);
	LUT4 #(
		.INIT('h57df)
	) name21383 (
		_w8650_,
		_w8653_,
		_w23282_,
		_w23283_,
		_w23284_
	);
	LUT3 #(
		.INIT('h80)
	) name21384 (
		\m0_data_i[20]_pad ,
		_w8655_,
		_w8656_,
		_w23285_
	);
	LUT3 #(
		.INIT('h2a)
	) name21385 (
		\m7_data_i[20]_pad ,
		_w8655_,
		_w8656_,
		_w23286_
	);
	LUT4 #(
		.INIT('h6e7f)
	) name21386 (
		_w8650_,
		_w8653_,
		_w23285_,
		_w23286_,
		_w23287_
	);
	LUT4 #(
		.INIT('h7fff)
	) name21387 (
		_w23278_,
		_w23281_,
		_w23284_,
		_w23287_,
		_w23288_
	);
	LUT3 #(
		.INIT('h2a)
	) name21388 (
		\m3_data_i[21]_pad ,
		_w8655_,
		_w8656_,
		_w23289_
	);
	LUT3 #(
		.INIT('h80)
	) name21389 (
		\m4_data_i[21]_pad ,
		_w8655_,
		_w8656_,
		_w23290_
	);
	LUT4 #(
		.INIT('h9dbf)
	) name21390 (
		_w8650_,
		_w8653_,
		_w23289_,
		_w23290_,
		_w23291_
	);
	LUT3 #(
		.INIT('h80)
	) name21391 (
		\m6_data_i[21]_pad ,
		_w8655_,
		_w8656_,
		_w23292_
	);
	LUT3 #(
		.INIT('h80)
	) name21392 (
		\m2_data_i[21]_pad ,
		_w8655_,
		_w8656_,
		_w23293_
	);
	LUT4 #(
		.INIT('habef)
	) name21393 (
		_w8650_,
		_w8653_,
		_w23292_,
		_w23293_,
		_w23294_
	);
	LUT3 #(
		.INIT('h2a)
	) name21394 (
		\m5_data_i[21]_pad ,
		_w8655_,
		_w8656_,
		_w23295_
	);
	LUT3 #(
		.INIT('h2a)
	) name21395 (
		\m1_data_i[21]_pad ,
		_w8655_,
		_w8656_,
		_w23296_
	);
	LUT4 #(
		.INIT('h57df)
	) name21396 (
		_w8650_,
		_w8653_,
		_w23295_,
		_w23296_,
		_w23297_
	);
	LUT3 #(
		.INIT('h80)
	) name21397 (
		\m0_data_i[21]_pad ,
		_w8655_,
		_w8656_,
		_w23298_
	);
	LUT3 #(
		.INIT('h2a)
	) name21398 (
		\m7_data_i[21]_pad ,
		_w8655_,
		_w8656_,
		_w23299_
	);
	LUT4 #(
		.INIT('h6e7f)
	) name21399 (
		_w8650_,
		_w8653_,
		_w23298_,
		_w23299_,
		_w23300_
	);
	LUT4 #(
		.INIT('h7fff)
	) name21400 (
		_w23291_,
		_w23294_,
		_w23297_,
		_w23300_,
		_w23301_
	);
	LUT3 #(
		.INIT('h2a)
	) name21401 (
		\m3_data_i[22]_pad ,
		_w8655_,
		_w8656_,
		_w23302_
	);
	LUT3 #(
		.INIT('h80)
	) name21402 (
		\m4_data_i[22]_pad ,
		_w8655_,
		_w8656_,
		_w23303_
	);
	LUT4 #(
		.INIT('h9dbf)
	) name21403 (
		_w8650_,
		_w8653_,
		_w23302_,
		_w23303_,
		_w23304_
	);
	LUT3 #(
		.INIT('h80)
	) name21404 (
		\m6_data_i[22]_pad ,
		_w8655_,
		_w8656_,
		_w23305_
	);
	LUT3 #(
		.INIT('h80)
	) name21405 (
		\m2_data_i[22]_pad ,
		_w8655_,
		_w8656_,
		_w23306_
	);
	LUT4 #(
		.INIT('habef)
	) name21406 (
		_w8650_,
		_w8653_,
		_w23305_,
		_w23306_,
		_w23307_
	);
	LUT3 #(
		.INIT('h2a)
	) name21407 (
		\m5_data_i[22]_pad ,
		_w8655_,
		_w8656_,
		_w23308_
	);
	LUT3 #(
		.INIT('h2a)
	) name21408 (
		\m1_data_i[22]_pad ,
		_w8655_,
		_w8656_,
		_w23309_
	);
	LUT4 #(
		.INIT('h57df)
	) name21409 (
		_w8650_,
		_w8653_,
		_w23308_,
		_w23309_,
		_w23310_
	);
	LUT3 #(
		.INIT('h80)
	) name21410 (
		\m0_data_i[22]_pad ,
		_w8655_,
		_w8656_,
		_w23311_
	);
	LUT3 #(
		.INIT('h2a)
	) name21411 (
		\m7_data_i[22]_pad ,
		_w8655_,
		_w8656_,
		_w23312_
	);
	LUT4 #(
		.INIT('h6e7f)
	) name21412 (
		_w8650_,
		_w8653_,
		_w23311_,
		_w23312_,
		_w23313_
	);
	LUT4 #(
		.INIT('h7fff)
	) name21413 (
		_w23304_,
		_w23307_,
		_w23310_,
		_w23313_,
		_w23314_
	);
	LUT3 #(
		.INIT('h2a)
	) name21414 (
		\m3_data_i[23]_pad ,
		_w8655_,
		_w8656_,
		_w23315_
	);
	LUT3 #(
		.INIT('h80)
	) name21415 (
		\m4_data_i[23]_pad ,
		_w8655_,
		_w8656_,
		_w23316_
	);
	LUT4 #(
		.INIT('h9dbf)
	) name21416 (
		_w8650_,
		_w8653_,
		_w23315_,
		_w23316_,
		_w23317_
	);
	LUT3 #(
		.INIT('h80)
	) name21417 (
		\m6_data_i[23]_pad ,
		_w8655_,
		_w8656_,
		_w23318_
	);
	LUT3 #(
		.INIT('h80)
	) name21418 (
		\m2_data_i[23]_pad ,
		_w8655_,
		_w8656_,
		_w23319_
	);
	LUT4 #(
		.INIT('habef)
	) name21419 (
		_w8650_,
		_w8653_,
		_w23318_,
		_w23319_,
		_w23320_
	);
	LUT3 #(
		.INIT('h2a)
	) name21420 (
		\m5_data_i[23]_pad ,
		_w8655_,
		_w8656_,
		_w23321_
	);
	LUT3 #(
		.INIT('h2a)
	) name21421 (
		\m1_data_i[23]_pad ,
		_w8655_,
		_w8656_,
		_w23322_
	);
	LUT4 #(
		.INIT('h57df)
	) name21422 (
		_w8650_,
		_w8653_,
		_w23321_,
		_w23322_,
		_w23323_
	);
	LUT3 #(
		.INIT('h80)
	) name21423 (
		\m0_data_i[23]_pad ,
		_w8655_,
		_w8656_,
		_w23324_
	);
	LUT3 #(
		.INIT('h2a)
	) name21424 (
		\m7_data_i[23]_pad ,
		_w8655_,
		_w8656_,
		_w23325_
	);
	LUT4 #(
		.INIT('h6e7f)
	) name21425 (
		_w8650_,
		_w8653_,
		_w23324_,
		_w23325_,
		_w23326_
	);
	LUT4 #(
		.INIT('h7fff)
	) name21426 (
		_w23317_,
		_w23320_,
		_w23323_,
		_w23326_,
		_w23327_
	);
	LUT3 #(
		.INIT('h2a)
	) name21427 (
		\m3_data_i[24]_pad ,
		_w8655_,
		_w8656_,
		_w23328_
	);
	LUT3 #(
		.INIT('h80)
	) name21428 (
		\m4_data_i[24]_pad ,
		_w8655_,
		_w8656_,
		_w23329_
	);
	LUT4 #(
		.INIT('h9dbf)
	) name21429 (
		_w8650_,
		_w8653_,
		_w23328_,
		_w23329_,
		_w23330_
	);
	LUT3 #(
		.INIT('h80)
	) name21430 (
		\m6_data_i[24]_pad ,
		_w8655_,
		_w8656_,
		_w23331_
	);
	LUT3 #(
		.INIT('h80)
	) name21431 (
		\m2_data_i[24]_pad ,
		_w8655_,
		_w8656_,
		_w23332_
	);
	LUT4 #(
		.INIT('habef)
	) name21432 (
		_w8650_,
		_w8653_,
		_w23331_,
		_w23332_,
		_w23333_
	);
	LUT3 #(
		.INIT('h2a)
	) name21433 (
		\m5_data_i[24]_pad ,
		_w8655_,
		_w8656_,
		_w23334_
	);
	LUT3 #(
		.INIT('h2a)
	) name21434 (
		\m1_data_i[24]_pad ,
		_w8655_,
		_w8656_,
		_w23335_
	);
	LUT4 #(
		.INIT('h57df)
	) name21435 (
		_w8650_,
		_w8653_,
		_w23334_,
		_w23335_,
		_w23336_
	);
	LUT3 #(
		.INIT('h80)
	) name21436 (
		\m0_data_i[24]_pad ,
		_w8655_,
		_w8656_,
		_w23337_
	);
	LUT3 #(
		.INIT('h2a)
	) name21437 (
		\m7_data_i[24]_pad ,
		_w8655_,
		_w8656_,
		_w23338_
	);
	LUT4 #(
		.INIT('h6e7f)
	) name21438 (
		_w8650_,
		_w8653_,
		_w23337_,
		_w23338_,
		_w23339_
	);
	LUT4 #(
		.INIT('h7fff)
	) name21439 (
		_w23330_,
		_w23333_,
		_w23336_,
		_w23339_,
		_w23340_
	);
	LUT3 #(
		.INIT('h2a)
	) name21440 (
		\m3_data_i[25]_pad ,
		_w8655_,
		_w8656_,
		_w23341_
	);
	LUT3 #(
		.INIT('h80)
	) name21441 (
		\m4_data_i[25]_pad ,
		_w8655_,
		_w8656_,
		_w23342_
	);
	LUT4 #(
		.INIT('h9dbf)
	) name21442 (
		_w8650_,
		_w8653_,
		_w23341_,
		_w23342_,
		_w23343_
	);
	LUT3 #(
		.INIT('h80)
	) name21443 (
		\m6_data_i[25]_pad ,
		_w8655_,
		_w8656_,
		_w23344_
	);
	LUT3 #(
		.INIT('h80)
	) name21444 (
		\m2_data_i[25]_pad ,
		_w8655_,
		_w8656_,
		_w23345_
	);
	LUT4 #(
		.INIT('habef)
	) name21445 (
		_w8650_,
		_w8653_,
		_w23344_,
		_w23345_,
		_w23346_
	);
	LUT3 #(
		.INIT('h2a)
	) name21446 (
		\m5_data_i[25]_pad ,
		_w8655_,
		_w8656_,
		_w23347_
	);
	LUT3 #(
		.INIT('h2a)
	) name21447 (
		\m1_data_i[25]_pad ,
		_w8655_,
		_w8656_,
		_w23348_
	);
	LUT4 #(
		.INIT('h57df)
	) name21448 (
		_w8650_,
		_w8653_,
		_w23347_,
		_w23348_,
		_w23349_
	);
	LUT3 #(
		.INIT('h80)
	) name21449 (
		\m0_data_i[25]_pad ,
		_w8655_,
		_w8656_,
		_w23350_
	);
	LUT3 #(
		.INIT('h2a)
	) name21450 (
		\m7_data_i[25]_pad ,
		_w8655_,
		_w8656_,
		_w23351_
	);
	LUT4 #(
		.INIT('h6e7f)
	) name21451 (
		_w8650_,
		_w8653_,
		_w23350_,
		_w23351_,
		_w23352_
	);
	LUT4 #(
		.INIT('h7fff)
	) name21452 (
		_w23343_,
		_w23346_,
		_w23349_,
		_w23352_,
		_w23353_
	);
	LUT3 #(
		.INIT('h2a)
	) name21453 (
		\m3_data_i[26]_pad ,
		_w8655_,
		_w8656_,
		_w23354_
	);
	LUT3 #(
		.INIT('h80)
	) name21454 (
		\m4_data_i[26]_pad ,
		_w8655_,
		_w8656_,
		_w23355_
	);
	LUT4 #(
		.INIT('h9dbf)
	) name21455 (
		_w8650_,
		_w8653_,
		_w23354_,
		_w23355_,
		_w23356_
	);
	LUT3 #(
		.INIT('h80)
	) name21456 (
		\m6_data_i[26]_pad ,
		_w8655_,
		_w8656_,
		_w23357_
	);
	LUT3 #(
		.INIT('h80)
	) name21457 (
		\m2_data_i[26]_pad ,
		_w8655_,
		_w8656_,
		_w23358_
	);
	LUT4 #(
		.INIT('habef)
	) name21458 (
		_w8650_,
		_w8653_,
		_w23357_,
		_w23358_,
		_w23359_
	);
	LUT3 #(
		.INIT('h2a)
	) name21459 (
		\m5_data_i[26]_pad ,
		_w8655_,
		_w8656_,
		_w23360_
	);
	LUT3 #(
		.INIT('h2a)
	) name21460 (
		\m1_data_i[26]_pad ,
		_w8655_,
		_w8656_,
		_w23361_
	);
	LUT4 #(
		.INIT('h57df)
	) name21461 (
		_w8650_,
		_w8653_,
		_w23360_,
		_w23361_,
		_w23362_
	);
	LUT3 #(
		.INIT('h80)
	) name21462 (
		\m0_data_i[26]_pad ,
		_w8655_,
		_w8656_,
		_w23363_
	);
	LUT3 #(
		.INIT('h2a)
	) name21463 (
		\m7_data_i[26]_pad ,
		_w8655_,
		_w8656_,
		_w23364_
	);
	LUT4 #(
		.INIT('h6e7f)
	) name21464 (
		_w8650_,
		_w8653_,
		_w23363_,
		_w23364_,
		_w23365_
	);
	LUT4 #(
		.INIT('h7fff)
	) name21465 (
		_w23356_,
		_w23359_,
		_w23362_,
		_w23365_,
		_w23366_
	);
	LUT3 #(
		.INIT('h2a)
	) name21466 (
		\m3_data_i[27]_pad ,
		_w8655_,
		_w8656_,
		_w23367_
	);
	LUT3 #(
		.INIT('h80)
	) name21467 (
		\m4_data_i[27]_pad ,
		_w8655_,
		_w8656_,
		_w23368_
	);
	LUT4 #(
		.INIT('h9dbf)
	) name21468 (
		_w8650_,
		_w8653_,
		_w23367_,
		_w23368_,
		_w23369_
	);
	LUT3 #(
		.INIT('h80)
	) name21469 (
		\m6_data_i[27]_pad ,
		_w8655_,
		_w8656_,
		_w23370_
	);
	LUT3 #(
		.INIT('h80)
	) name21470 (
		\m2_data_i[27]_pad ,
		_w8655_,
		_w8656_,
		_w23371_
	);
	LUT4 #(
		.INIT('habef)
	) name21471 (
		_w8650_,
		_w8653_,
		_w23370_,
		_w23371_,
		_w23372_
	);
	LUT3 #(
		.INIT('h2a)
	) name21472 (
		\m5_data_i[27]_pad ,
		_w8655_,
		_w8656_,
		_w23373_
	);
	LUT3 #(
		.INIT('h2a)
	) name21473 (
		\m1_data_i[27]_pad ,
		_w8655_,
		_w8656_,
		_w23374_
	);
	LUT4 #(
		.INIT('h57df)
	) name21474 (
		_w8650_,
		_w8653_,
		_w23373_,
		_w23374_,
		_w23375_
	);
	LUT3 #(
		.INIT('h80)
	) name21475 (
		\m0_data_i[27]_pad ,
		_w8655_,
		_w8656_,
		_w23376_
	);
	LUT3 #(
		.INIT('h2a)
	) name21476 (
		\m7_data_i[27]_pad ,
		_w8655_,
		_w8656_,
		_w23377_
	);
	LUT4 #(
		.INIT('h6e7f)
	) name21477 (
		_w8650_,
		_w8653_,
		_w23376_,
		_w23377_,
		_w23378_
	);
	LUT4 #(
		.INIT('h7fff)
	) name21478 (
		_w23369_,
		_w23372_,
		_w23375_,
		_w23378_,
		_w23379_
	);
	LUT3 #(
		.INIT('h2a)
	) name21479 (
		\m3_data_i[28]_pad ,
		_w8655_,
		_w8656_,
		_w23380_
	);
	LUT3 #(
		.INIT('h80)
	) name21480 (
		\m4_data_i[28]_pad ,
		_w8655_,
		_w8656_,
		_w23381_
	);
	LUT4 #(
		.INIT('h9dbf)
	) name21481 (
		_w8650_,
		_w8653_,
		_w23380_,
		_w23381_,
		_w23382_
	);
	LUT3 #(
		.INIT('h80)
	) name21482 (
		\m6_data_i[28]_pad ,
		_w8655_,
		_w8656_,
		_w23383_
	);
	LUT3 #(
		.INIT('h80)
	) name21483 (
		\m2_data_i[28]_pad ,
		_w8655_,
		_w8656_,
		_w23384_
	);
	LUT4 #(
		.INIT('habef)
	) name21484 (
		_w8650_,
		_w8653_,
		_w23383_,
		_w23384_,
		_w23385_
	);
	LUT3 #(
		.INIT('h2a)
	) name21485 (
		\m5_data_i[28]_pad ,
		_w8655_,
		_w8656_,
		_w23386_
	);
	LUT3 #(
		.INIT('h2a)
	) name21486 (
		\m1_data_i[28]_pad ,
		_w8655_,
		_w8656_,
		_w23387_
	);
	LUT4 #(
		.INIT('h57df)
	) name21487 (
		_w8650_,
		_w8653_,
		_w23386_,
		_w23387_,
		_w23388_
	);
	LUT3 #(
		.INIT('h80)
	) name21488 (
		\m0_data_i[28]_pad ,
		_w8655_,
		_w8656_,
		_w23389_
	);
	LUT3 #(
		.INIT('h2a)
	) name21489 (
		\m7_data_i[28]_pad ,
		_w8655_,
		_w8656_,
		_w23390_
	);
	LUT4 #(
		.INIT('h6e7f)
	) name21490 (
		_w8650_,
		_w8653_,
		_w23389_,
		_w23390_,
		_w23391_
	);
	LUT4 #(
		.INIT('h7fff)
	) name21491 (
		_w23382_,
		_w23385_,
		_w23388_,
		_w23391_,
		_w23392_
	);
	LUT3 #(
		.INIT('h2a)
	) name21492 (
		\m3_data_i[29]_pad ,
		_w8655_,
		_w8656_,
		_w23393_
	);
	LUT3 #(
		.INIT('h80)
	) name21493 (
		\m4_data_i[29]_pad ,
		_w8655_,
		_w8656_,
		_w23394_
	);
	LUT4 #(
		.INIT('h9dbf)
	) name21494 (
		_w8650_,
		_w8653_,
		_w23393_,
		_w23394_,
		_w23395_
	);
	LUT3 #(
		.INIT('h80)
	) name21495 (
		\m6_data_i[29]_pad ,
		_w8655_,
		_w8656_,
		_w23396_
	);
	LUT3 #(
		.INIT('h80)
	) name21496 (
		\m2_data_i[29]_pad ,
		_w8655_,
		_w8656_,
		_w23397_
	);
	LUT4 #(
		.INIT('habef)
	) name21497 (
		_w8650_,
		_w8653_,
		_w23396_,
		_w23397_,
		_w23398_
	);
	LUT3 #(
		.INIT('h2a)
	) name21498 (
		\m5_data_i[29]_pad ,
		_w8655_,
		_w8656_,
		_w23399_
	);
	LUT3 #(
		.INIT('h2a)
	) name21499 (
		\m1_data_i[29]_pad ,
		_w8655_,
		_w8656_,
		_w23400_
	);
	LUT4 #(
		.INIT('h57df)
	) name21500 (
		_w8650_,
		_w8653_,
		_w23399_,
		_w23400_,
		_w23401_
	);
	LUT3 #(
		.INIT('h80)
	) name21501 (
		\m0_data_i[29]_pad ,
		_w8655_,
		_w8656_,
		_w23402_
	);
	LUT3 #(
		.INIT('h2a)
	) name21502 (
		\m7_data_i[29]_pad ,
		_w8655_,
		_w8656_,
		_w23403_
	);
	LUT4 #(
		.INIT('h6e7f)
	) name21503 (
		_w8650_,
		_w8653_,
		_w23402_,
		_w23403_,
		_w23404_
	);
	LUT4 #(
		.INIT('h7fff)
	) name21504 (
		_w23395_,
		_w23398_,
		_w23401_,
		_w23404_,
		_w23405_
	);
	LUT3 #(
		.INIT('h2a)
	) name21505 (
		\m3_data_i[2]_pad ,
		_w8655_,
		_w8656_,
		_w23406_
	);
	LUT3 #(
		.INIT('h80)
	) name21506 (
		\m4_data_i[2]_pad ,
		_w8655_,
		_w8656_,
		_w23407_
	);
	LUT4 #(
		.INIT('h9dbf)
	) name21507 (
		_w8650_,
		_w8653_,
		_w23406_,
		_w23407_,
		_w23408_
	);
	LUT3 #(
		.INIT('h80)
	) name21508 (
		\m6_data_i[2]_pad ,
		_w8655_,
		_w8656_,
		_w23409_
	);
	LUT3 #(
		.INIT('h80)
	) name21509 (
		\m2_data_i[2]_pad ,
		_w8655_,
		_w8656_,
		_w23410_
	);
	LUT4 #(
		.INIT('habef)
	) name21510 (
		_w8650_,
		_w8653_,
		_w23409_,
		_w23410_,
		_w23411_
	);
	LUT3 #(
		.INIT('h2a)
	) name21511 (
		\m5_data_i[2]_pad ,
		_w8655_,
		_w8656_,
		_w23412_
	);
	LUT3 #(
		.INIT('h2a)
	) name21512 (
		\m1_data_i[2]_pad ,
		_w8655_,
		_w8656_,
		_w23413_
	);
	LUT4 #(
		.INIT('h57df)
	) name21513 (
		_w8650_,
		_w8653_,
		_w23412_,
		_w23413_,
		_w23414_
	);
	LUT3 #(
		.INIT('h80)
	) name21514 (
		\m0_data_i[2]_pad ,
		_w8655_,
		_w8656_,
		_w23415_
	);
	LUT3 #(
		.INIT('h2a)
	) name21515 (
		\m7_data_i[2]_pad ,
		_w8655_,
		_w8656_,
		_w23416_
	);
	LUT4 #(
		.INIT('h6e7f)
	) name21516 (
		_w8650_,
		_w8653_,
		_w23415_,
		_w23416_,
		_w23417_
	);
	LUT4 #(
		.INIT('h7fff)
	) name21517 (
		_w23408_,
		_w23411_,
		_w23414_,
		_w23417_,
		_w23418_
	);
	LUT3 #(
		.INIT('h2a)
	) name21518 (
		\m3_data_i[30]_pad ,
		_w8655_,
		_w8656_,
		_w23419_
	);
	LUT3 #(
		.INIT('h80)
	) name21519 (
		\m4_data_i[30]_pad ,
		_w8655_,
		_w8656_,
		_w23420_
	);
	LUT4 #(
		.INIT('h9dbf)
	) name21520 (
		_w8650_,
		_w8653_,
		_w23419_,
		_w23420_,
		_w23421_
	);
	LUT3 #(
		.INIT('h80)
	) name21521 (
		\m6_data_i[30]_pad ,
		_w8655_,
		_w8656_,
		_w23422_
	);
	LUT3 #(
		.INIT('h80)
	) name21522 (
		\m2_data_i[30]_pad ,
		_w8655_,
		_w8656_,
		_w23423_
	);
	LUT4 #(
		.INIT('habef)
	) name21523 (
		_w8650_,
		_w8653_,
		_w23422_,
		_w23423_,
		_w23424_
	);
	LUT3 #(
		.INIT('h2a)
	) name21524 (
		\m5_data_i[30]_pad ,
		_w8655_,
		_w8656_,
		_w23425_
	);
	LUT3 #(
		.INIT('h2a)
	) name21525 (
		\m1_data_i[30]_pad ,
		_w8655_,
		_w8656_,
		_w23426_
	);
	LUT4 #(
		.INIT('h57df)
	) name21526 (
		_w8650_,
		_w8653_,
		_w23425_,
		_w23426_,
		_w23427_
	);
	LUT3 #(
		.INIT('h80)
	) name21527 (
		\m0_data_i[30]_pad ,
		_w8655_,
		_w8656_,
		_w23428_
	);
	LUT3 #(
		.INIT('h2a)
	) name21528 (
		\m7_data_i[30]_pad ,
		_w8655_,
		_w8656_,
		_w23429_
	);
	LUT4 #(
		.INIT('h6e7f)
	) name21529 (
		_w8650_,
		_w8653_,
		_w23428_,
		_w23429_,
		_w23430_
	);
	LUT4 #(
		.INIT('h7fff)
	) name21530 (
		_w23421_,
		_w23424_,
		_w23427_,
		_w23430_,
		_w23431_
	);
	LUT3 #(
		.INIT('h2a)
	) name21531 (
		\m3_data_i[31]_pad ,
		_w8655_,
		_w8656_,
		_w23432_
	);
	LUT3 #(
		.INIT('h80)
	) name21532 (
		\m4_data_i[31]_pad ,
		_w8655_,
		_w8656_,
		_w23433_
	);
	LUT4 #(
		.INIT('h9dbf)
	) name21533 (
		_w8650_,
		_w8653_,
		_w23432_,
		_w23433_,
		_w23434_
	);
	LUT3 #(
		.INIT('h80)
	) name21534 (
		\m6_data_i[31]_pad ,
		_w8655_,
		_w8656_,
		_w23435_
	);
	LUT3 #(
		.INIT('h80)
	) name21535 (
		\m2_data_i[31]_pad ,
		_w8655_,
		_w8656_,
		_w23436_
	);
	LUT4 #(
		.INIT('habef)
	) name21536 (
		_w8650_,
		_w8653_,
		_w23435_,
		_w23436_,
		_w23437_
	);
	LUT3 #(
		.INIT('h2a)
	) name21537 (
		\m5_data_i[31]_pad ,
		_w8655_,
		_w8656_,
		_w23438_
	);
	LUT3 #(
		.INIT('h2a)
	) name21538 (
		\m1_data_i[31]_pad ,
		_w8655_,
		_w8656_,
		_w23439_
	);
	LUT4 #(
		.INIT('h57df)
	) name21539 (
		_w8650_,
		_w8653_,
		_w23438_,
		_w23439_,
		_w23440_
	);
	LUT3 #(
		.INIT('h80)
	) name21540 (
		\m0_data_i[31]_pad ,
		_w8655_,
		_w8656_,
		_w23441_
	);
	LUT3 #(
		.INIT('h2a)
	) name21541 (
		\m7_data_i[31]_pad ,
		_w8655_,
		_w8656_,
		_w23442_
	);
	LUT4 #(
		.INIT('h6e7f)
	) name21542 (
		_w8650_,
		_w8653_,
		_w23441_,
		_w23442_,
		_w23443_
	);
	LUT4 #(
		.INIT('h7fff)
	) name21543 (
		_w23434_,
		_w23437_,
		_w23440_,
		_w23443_,
		_w23444_
	);
	LUT3 #(
		.INIT('h2a)
	) name21544 (
		\m3_data_i[3]_pad ,
		_w8655_,
		_w8656_,
		_w23445_
	);
	LUT3 #(
		.INIT('h80)
	) name21545 (
		\m4_data_i[3]_pad ,
		_w8655_,
		_w8656_,
		_w23446_
	);
	LUT4 #(
		.INIT('h9dbf)
	) name21546 (
		_w8650_,
		_w8653_,
		_w23445_,
		_w23446_,
		_w23447_
	);
	LUT3 #(
		.INIT('h80)
	) name21547 (
		\m6_data_i[3]_pad ,
		_w8655_,
		_w8656_,
		_w23448_
	);
	LUT3 #(
		.INIT('h80)
	) name21548 (
		\m2_data_i[3]_pad ,
		_w8655_,
		_w8656_,
		_w23449_
	);
	LUT4 #(
		.INIT('habef)
	) name21549 (
		_w8650_,
		_w8653_,
		_w23448_,
		_w23449_,
		_w23450_
	);
	LUT3 #(
		.INIT('h2a)
	) name21550 (
		\m5_data_i[3]_pad ,
		_w8655_,
		_w8656_,
		_w23451_
	);
	LUT3 #(
		.INIT('h2a)
	) name21551 (
		\m1_data_i[3]_pad ,
		_w8655_,
		_w8656_,
		_w23452_
	);
	LUT4 #(
		.INIT('h57df)
	) name21552 (
		_w8650_,
		_w8653_,
		_w23451_,
		_w23452_,
		_w23453_
	);
	LUT3 #(
		.INIT('h80)
	) name21553 (
		\m0_data_i[3]_pad ,
		_w8655_,
		_w8656_,
		_w23454_
	);
	LUT3 #(
		.INIT('h2a)
	) name21554 (
		\m7_data_i[3]_pad ,
		_w8655_,
		_w8656_,
		_w23455_
	);
	LUT4 #(
		.INIT('h6e7f)
	) name21555 (
		_w8650_,
		_w8653_,
		_w23454_,
		_w23455_,
		_w23456_
	);
	LUT4 #(
		.INIT('h7fff)
	) name21556 (
		_w23447_,
		_w23450_,
		_w23453_,
		_w23456_,
		_w23457_
	);
	LUT3 #(
		.INIT('h2a)
	) name21557 (
		\m3_data_i[4]_pad ,
		_w8655_,
		_w8656_,
		_w23458_
	);
	LUT3 #(
		.INIT('h80)
	) name21558 (
		\m4_data_i[4]_pad ,
		_w8655_,
		_w8656_,
		_w23459_
	);
	LUT4 #(
		.INIT('h9dbf)
	) name21559 (
		_w8650_,
		_w8653_,
		_w23458_,
		_w23459_,
		_w23460_
	);
	LUT3 #(
		.INIT('h80)
	) name21560 (
		\m6_data_i[4]_pad ,
		_w8655_,
		_w8656_,
		_w23461_
	);
	LUT3 #(
		.INIT('h80)
	) name21561 (
		\m2_data_i[4]_pad ,
		_w8655_,
		_w8656_,
		_w23462_
	);
	LUT4 #(
		.INIT('habef)
	) name21562 (
		_w8650_,
		_w8653_,
		_w23461_,
		_w23462_,
		_w23463_
	);
	LUT3 #(
		.INIT('h2a)
	) name21563 (
		\m5_data_i[4]_pad ,
		_w8655_,
		_w8656_,
		_w23464_
	);
	LUT3 #(
		.INIT('h2a)
	) name21564 (
		\m1_data_i[4]_pad ,
		_w8655_,
		_w8656_,
		_w23465_
	);
	LUT4 #(
		.INIT('h57df)
	) name21565 (
		_w8650_,
		_w8653_,
		_w23464_,
		_w23465_,
		_w23466_
	);
	LUT3 #(
		.INIT('h80)
	) name21566 (
		\m0_data_i[4]_pad ,
		_w8655_,
		_w8656_,
		_w23467_
	);
	LUT3 #(
		.INIT('h2a)
	) name21567 (
		\m7_data_i[4]_pad ,
		_w8655_,
		_w8656_,
		_w23468_
	);
	LUT4 #(
		.INIT('h6e7f)
	) name21568 (
		_w8650_,
		_w8653_,
		_w23467_,
		_w23468_,
		_w23469_
	);
	LUT4 #(
		.INIT('h7fff)
	) name21569 (
		_w23460_,
		_w23463_,
		_w23466_,
		_w23469_,
		_w23470_
	);
	LUT3 #(
		.INIT('h2a)
	) name21570 (
		\m3_data_i[5]_pad ,
		_w8655_,
		_w8656_,
		_w23471_
	);
	LUT3 #(
		.INIT('h80)
	) name21571 (
		\m4_data_i[5]_pad ,
		_w8655_,
		_w8656_,
		_w23472_
	);
	LUT4 #(
		.INIT('h9dbf)
	) name21572 (
		_w8650_,
		_w8653_,
		_w23471_,
		_w23472_,
		_w23473_
	);
	LUT3 #(
		.INIT('h80)
	) name21573 (
		\m6_data_i[5]_pad ,
		_w8655_,
		_w8656_,
		_w23474_
	);
	LUT3 #(
		.INIT('h80)
	) name21574 (
		\m2_data_i[5]_pad ,
		_w8655_,
		_w8656_,
		_w23475_
	);
	LUT4 #(
		.INIT('habef)
	) name21575 (
		_w8650_,
		_w8653_,
		_w23474_,
		_w23475_,
		_w23476_
	);
	LUT3 #(
		.INIT('h2a)
	) name21576 (
		\m5_data_i[5]_pad ,
		_w8655_,
		_w8656_,
		_w23477_
	);
	LUT3 #(
		.INIT('h2a)
	) name21577 (
		\m1_data_i[5]_pad ,
		_w8655_,
		_w8656_,
		_w23478_
	);
	LUT4 #(
		.INIT('h57df)
	) name21578 (
		_w8650_,
		_w8653_,
		_w23477_,
		_w23478_,
		_w23479_
	);
	LUT3 #(
		.INIT('h80)
	) name21579 (
		\m0_data_i[5]_pad ,
		_w8655_,
		_w8656_,
		_w23480_
	);
	LUT3 #(
		.INIT('h2a)
	) name21580 (
		\m7_data_i[5]_pad ,
		_w8655_,
		_w8656_,
		_w23481_
	);
	LUT4 #(
		.INIT('h6e7f)
	) name21581 (
		_w8650_,
		_w8653_,
		_w23480_,
		_w23481_,
		_w23482_
	);
	LUT4 #(
		.INIT('h7fff)
	) name21582 (
		_w23473_,
		_w23476_,
		_w23479_,
		_w23482_,
		_w23483_
	);
	LUT3 #(
		.INIT('h2a)
	) name21583 (
		\m3_data_i[6]_pad ,
		_w8655_,
		_w8656_,
		_w23484_
	);
	LUT3 #(
		.INIT('h80)
	) name21584 (
		\m4_data_i[6]_pad ,
		_w8655_,
		_w8656_,
		_w23485_
	);
	LUT4 #(
		.INIT('h9dbf)
	) name21585 (
		_w8650_,
		_w8653_,
		_w23484_,
		_w23485_,
		_w23486_
	);
	LUT3 #(
		.INIT('h80)
	) name21586 (
		\m6_data_i[6]_pad ,
		_w8655_,
		_w8656_,
		_w23487_
	);
	LUT3 #(
		.INIT('h80)
	) name21587 (
		\m2_data_i[6]_pad ,
		_w8655_,
		_w8656_,
		_w23488_
	);
	LUT4 #(
		.INIT('habef)
	) name21588 (
		_w8650_,
		_w8653_,
		_w23487_,
		_w23488_,
		_w23489_
	);
	LUT3 #(
		.INIT('h2a)
	) name21589 (
		\m5_data_i[6]_pad ,
		_w8655_,
		_w8656_,
		_w23490_
	);
	LUT3 #(
		.INIT('h2a)
	) name21590 (
		\m1_data_i[6]_pad ,
		_w8655_,
		_w8656_,
		_w23491_
	);
	LUT4 #(
		.INIT('h57df)
	) name21591 (
		_w8650_,
		_w8653_,
		_w23490_,
		_w23491_,
		_w23492_
	);
	LUT3 #(
		.INIT('h80)
	) name21592 (
		\m0_data_i[6]_pad ,
		_w8655_,
		_w8656_,
		_w23493_
	);
	LUT3 #(
		.INIT('h2a)
	) name21593 (
		\m7_data_i[6]_pad ,
		_w8655_,
		_w8656_,
		_w23494_
	);
	LUT4 #(
		.INIT('h6e7f)
	) name21594 (
		_w8650_,
		_w8653_,
		_w23493_,
		_w23494_,
		_w23495_
	);
	LUT4 #(
		.INIT('h7fff)
	) name21595 (
		_w23486_,
		_w23489_,
		_w23492_,
		_w23495_,
		_w23496_
	);
	LUT3 #(
		.INIT('h2a)
	) name21596 (
		\m3_data_i[7]_pad ,
		_w8655_,
		_w8656_,
		_w23497_
	);
	LUT3 #(
		.INIT('h80)
	) name21597 (
		\m4_data_i[7]_pad ,
		_w8655_,
		_w8656_,
		_w23498_
	);
	LUT4 #(
		.INIT('h9dbf)
	) name21598 (
		_w8650_,
		_w8653_,
		_w23497_,
		_w23498_,
		_w23499_
	);
	LUT3 #(
		.INIT('h80)
	) name21599 (
		\m6_data_i[7]_pad ,
		_w8655_,
		_w8656_,
		_w23500_
	);
	LUT3 #(
		.INIT('h80)
	) name21600 (
		\m2_data_i[7]_pad ,
		_w8655_,
		_w8656_,
		_w23501_
	);
	LUT4 #(
		.INIT('habef)
	) name21601 (
		_w8650_,
		_w8653_,
		_w23500_,
		_w23501_,
		_w23502_
	);
	LUT3 #(
		.INIT('h2a)
	) name21602 (
		\m5_data_i[7]_pad ,
		_w8655_,
		_w8656_,
		_w23503_
	);
	LUT3 #(
		.INIT('h2a)
	) name21603 (
		\m1_data_i[7]_pad ,
		_w8655_,
		_w8656_,
		_w23504_
	);
	LUT4 #(
		.INIT('h57df)
	) name21604 (
		_w8650_,
		_w8653_,
		_w23503_,
		_w23504_,
		_w23505_
	);
	LUT3 #(
		.INIT('h80)
	) name21605 (
		\m0_data_i[7]_pad ,
		_w8655_,
		_w8656_,
		_w23506_
	);
	LUT3 #(
		.INIT('h2a)
	) name21606 (
		\m7_data_i[7]_pad ,
		_w8655_,
		_w8656_,
		_w23507_
	);
	LUT4 #(
		.INIT('h6e7f)
	) name21607 (
		_w8650_,
		_w8653_,
		_w23506_,
		_w23507_,
		_w23508_
	);
	LUT4 #(
		.INIT('h7fff)
	) name21608 (
		_w23499_,
		_w23502_,
		_w23505_,
		_w23508_,
		_w23509_
	);
	LUT3 #(
		.INIT('h2a)
	) name21609 (
		\m3_data_i[8]_pad ,
		_w8655_,
		_w8656_,
		_w23510_
	);
	LUT3 #(
		.INIT('h80)
	) name21610 (
		\m4_data_i[8]_pad ,
		_w8655_,
		_w8656_,
		_w23511_
	);
	LUT4 #(
		.INIT('h9dbf)
	) name21611 (
		_w8650_,
		_w8653_,
		_w23510_,
		_w23511_,
		_w23512_
	);
	LUT3 #(
		.INIT('h80)
	) name21612 (
		\m6_data_i[8]_pad ,
		_w8655_,
		_w8656_,
		_w23513_
	);
	LUT3 #(
		.INIT('h80)
	) name21613 (
		\m2_data_i[8]_pad ,
		_w8655_,
		_w8656_,
		_w23514_
	);
	LUT4 #(
		.INIT('habef)
	) name21614 (
		_w8650_,
		_w8653_,
		_w23513_,
		_w23514_,
		_w23515_
	);
	LUT3 #(
		.INIT('h2a)
	) name21615 (
		\m5_data_i[8]_pad ,
		_w8655_,
		_w8656_,
		_w23516_
	);
	LUT3 #(
		.INIT('h2a)
	) name21616 (
		\m1_data_i[8]_pad ,
		_w8655_,
		_w8656_,
		_w23517_
	);
	LUT4 #(
		.INIT('h57df)
	) name21617 (
		_w8650_,
		_w8653_,
		_w23516_,
		_w23517_,
		_w23518_
	);
	LUT3 #(
		.INIT('h80)
	) name21618 (
		\m0_data_i[8]_pad ,
		_w8655_,
		_w8656_,
		_w23519_
	);
	LUT3 #(
		.INIT('h2a)
	) name21619 (
		\m7_data_i[8]_pad ,
		_w8655_,
		_w8656_,
		_w23520_
	);
	LUT4 #(
		.INIT('h6e7f)
	) name21620 (
		_w8650_,
		_w8653_,
		_w23519_,
		_w23520_,
		_w23521_
	);
	LUT4 #(
		.INIT('h7fff)
	) name21621 (
		_w23512_,
		_w23515_,
		_w23518_,
		_w23521_,
		_w23522_
	);
	LUT3 #(
		.INIT('h2a)
	) name21622 (
		\m3_data_i[9]_pad ,
		_w8655_,
		_w8656_,
		_w23523_
	);
	LUT3 #(
		.INIT('h80)
	) name21623 (
		\m4_data_i[9]_pad ,
		_w8655_,
		_w8656_,
		_w23524_
	);
	LUT4 #(
		.INIT('h9dbf)
	) name21624 (
		_w8650_,
		_w8653_,
		_w23523_,
		_w23524_,
		_w23525_
	);
	LUT3 #(
		.INIT('h80)
	) name21625 (
		\m6_data_i[9]_pad ,
		_w8655_,
		_w8656_,
		_w23526_
	);
	LUT3 #(
		.INIT('h80)
	) name21626 (
		\m2_data_i[9]_pad ,
		_w8655_,
		_w8656_,
		_w23527_
	);
	LUT4 #(
		.INIT('habef)
	) name21627 (
		_w8650_,
		_w8653_,
		_w23526_,
		_w23527_,
		_w23528_
	);
	LUT3 #(
		.INIT('h2a)
	) name21628 (
		\m5_data_i[9]_pad ,
		_w8655_,
		_w8656_,
		_w23529_
	);
	LUT3 #(
		.INIT('h2a)
	) name21629 (
		\m1_data_i[9]_pad ,
		_w8655_,
		_w8656_,
		_w23530_
	);
	LUT4 #(
		.INIT('h57df)
	) name21630 (
		_w8650_,
		_w8653_,
		_w23529_,
		_w23530_,
		_w23531_
	);
	LUT3 #(
		.INIT('h80)
	) name21631 (
		\m0_data_i[9]_pad ,
		_w8655_,
		_w8656_,
		_w23532_
	);
	LUT3 #(
		.INIT('h2a)
	) name21632 (
		\m7_data_i[9]_pad ,
		_w8655_,
		_w8656_,
		_w23533_
	);
	LUT4 #(
		.INIT('h6e7f)
	) name21633 (
		_w8650_,
		_w8653_,
		_w23532_,
		_w23533_,
		_w23534_
	);
	LUT4 #(
		.INIT('h7fff)
	) name21634 (
		_w23525_,
		_w23528_,
		_w23531_,
		_w23534_,
		_w23535_
	);
	LUT3 #(
		.INIT('h2a)
	) name21635 (
		\m3_sel_i[0]_pad ,
		_w8655_,
		_w8656_,
		_w23536_
	);
	LUT3 #(
		.INIT('h80)
	) name21636 (
		\m4_sel_i[0]_pad ,
		_w8655_,
		_w8656_,
		_w23537_
	);
	LUT4 #(
		.INIT('h9dbf)
	) name21637 (
		_w8650_,
		_w8653_,
		_w23536_,
		_w23537_,
		_w23538_
	);
	LUT3 #(
		.INIT('h80)
	) name21638 (
		\m6_sel_i[0]_pad ,
		_w8655_,
		_w8656_,
		_w23539_
	);
	LUT3 #(
		.INIT('h80)
	) name21639 (
		\m2_sel_i[0]_pad ,
		_w8655_,
		_w8656_,
		_w23540_
	);
	LUT4 #(
		.INIT('habef)
	) name21640 (
		_w8650_,
		_w8653_,
		_w23539_,
		_w23540_,
		_w23541_
	);
	LUT3 #(
		.INIT('h2a)
	) name21641 (
		\m5_sel_i[0]_pad ,
		_w8655_,
		_w8656_,
		_w23542_
	);
	LUT3 #(
		.INIT('h2a)
	) name21642 (
		\m1_sel_i[0]_pad ,
		_w8655_,
		_w8656_,
		_w23543_
	);
	LUT4 #(
		.INIT('h57df)
	) name21643 (
		_w8650_,
		_w8653_,
		_w23542_,
		_w23543_,
		_w23544_
	);
	LUT3 #(
		.INIT('h80)
	) name21644 (
		\m0_sel_i[0]_pad ,
		_w8655_,
		_w8656_,
		_w23545_
	);
	LUT3 #(
		.INIT('h2a)
	) name21645 (
		\m7_sel_i[0]_pad ,
		_w8655_,
		_w8656_,
		_w23546_
	);
	LUT4 #(
		.INIT('h6e7f)
	) name21646 (
		_w8650_,
		_w8653_,
		_w23545_,
		_w23546_,
		_w23547_
	);
	LUT4 #(
		.INIT('h7fff)
	) name21647 (
		_w23538_,
		_w23541_,
		_w23544_,
		_w23547_,
		_w23548_
	);
	LUT3 #(
		.INIT('h2a)
	) name21648 (
		\m3_sel_i[1]_pad ,
		_w8655_,
		_w8656_,
		_w23549_
	);
	LUT3 #(
		.INIT('h80)
	) name21649 (
		\m4_sel_i[1]_pad ,
		_w8655_,
		_w8656_,
		_w23550_
	);
	LUT4 #(
		.INIT('h9dbf)
	) name21650 (
		_w8650_,
		_w8653_,
		_w23549_,
		_w23550_,
		_w23551_
	);
	LUT3 #(
		.INIT('h80)
	) name21651 (
		\m6_sel_i[1]_pad ,
		_w8655_,
		_w8656_,
		_w23552_
	);
	LUT3 #(
		.INIT('h80)
	) name21652 (
		\m2_sel_i[1]_pad ,
		_w8655_,
		_w8656_,
		_w23553_
	);
	LUT4 #(
		.INIT('habef)
	) name21653 (
		_w8650_,
		_w8653_,
		_w23552_,
		_w23553_,
		_w23554_
	);
	LUT3 #(
		.INIT('h2a)
	) name21654 (
		\m5_sel_i[1]_pad ,
		_w8655_,
		_w8656_,
		_w23555_
	);
	LUT3 #(
		.INIT('h2a)
	) name21655 (
		\m1_sel_i[1]_pad ,
		_w8655_,
		_w8656_,
		_w23556_
	);
	LUT4 #(
		.INIT('h57df)
	) name21656 (
		_w8650_,
		_w8653_,
		_w23555_,
		_w23556_,
		_w23557_
	);
	LUT3 #(
		.INIT('h80)
	) name21657 (
		\m0_sel_i[1]_pad ,
		_w8655_,
		_w8656_,
		_w23558_
	);
	LUT3 #(
		.INIT('h2a)
	) name21658 (
		\m7_sel_i[1]_pad ,
		_w8655_,
		_w8656_,
		_w23559_
	);
	LUT4 #(
		.INIT('h6e7f)
	) name21659 (
		_w8650_,
		_w8653_,
		_w23558_,
		_w23559_,
		_w23560_
	);
	LUT4 #(
		.INIT('h7fff)
	) name21660 (
		_w23551_,
		_w23554_,
		_w23557_,
		_w23560_,
		_w23561_
	);
	LUT3 #(
		.INIT('h2a)
	) name21661 (
		\m3_sel_i[2]_pad ,
		_w8655_,
		_w8656_,
		_w23562_
	);
	LUT3 #(
		.INIT('h80)
	) name21662 (
		\m4_sel_i[2]_pad ,
		_w8655_,
		_w8656_,
		_w23563_
	);
	LUT4 #(
		.INIT('h9dbf)
	) name21663 (
		_w8650_,
		_w8653_,
		_w23562_,
		_w23563_,
		_w23564_
	);
	LUT3 #(
		.INIT('h80)
	) name21664 (
		\m6_sel_i[2]_pad ,
		_w8655_,
		_w8656_,
		_w23565_
	);
	LUT3 #(
		.INIT('h80)
	) name21665 (
		\m2_sel_i[2]_pad ,
		_w8655_,
		_w8656_,
		_w23566_
	);
	LUT4 #(
		.INIT('habef)
	) name21666 (
		_w8650_,
		_w8653_,
		_w23565_,
		_w23566_,
		_w23567_
	);
	LUT3 #(
		.INIT('h2a)
	) name21667 (
		\m5_sel_i[2]_pad ,
		_w8655_,
		_w8656_,
		_w23568_
	);
	LUT3 #(
		.INIT('h2a)
	) name21668 (
		\m1_sel_i[2]_pad ,
		_w8655_,
		_w8656_,
		_w23569_
	);
	LUT4 #(
		.INIT('h57df)
	) name21669 (
		_w8650_,
		_w8653_,
		_w23568_,
		_w23569_,
		_w23570_
	);
	LUT3 #(
		.INIT('h80)
	) name21670 (
		\m0_sel_i[2]_pad ,
		_w8655_,
		_w8656_,
		_w23571_
	);
	LUT3 #(
		.INIT('h2a)
	) name21671 (
		\m7_sel_i[2]_pad ,
		_w8655_,
		_w8656_,
		_w23572_
	);
	LUT4 #(
		.INIT('h6e7f)
	) name21672 (
		_w8650_,
		_w8653_,
		_w23571_,
		_w23572_,
		_w23573_
	);
	LUT4 #(
		.INIT('h7fff)
	) name21673 (
		_w23564_,
		_w23567_,
		_w23570_,
		_w23573_,
		_w23574_
	);
	LUT3 #(
		.INIT('h2a)
	) name21674 (
		\m3_sel_i[3]_pad ,
		_w8655_,
		_w8656_,
		_w23575_
	);
	LUT3 #(
		.INIT('h80)
	) name21675 (
		\m4_sel_i[3]_pad ,
		_w8655_,
		_w8656_,
		_w23576_
	);
	LUT4 #(
		.INIT('h9dbf)
	) name21676 (
		_w8650_,
		_w8653_,
		_w23575_,
		_w23576_,
		_w23577_
	);
	LUT3 #(
		.INIT('h80)
	) name21677 (
		\m6_sel_i[3]_pad ,
		_w8655_,
		_w8656_,
		_w23578_
	);
	LUT3 #(
		.INIT('h80)
	) name21678 (
		\m2_sel_i[3]_pad ,
		_w8655_,
		_w8656_,
		_w23579_
	);
	LUT4 #(
		.INIT('habef)
	) name21679 (
		_w8650_,
		_w8653_,
		_w23578_,
		_w23579_,
		_w23580_
	);
	LUT3 #(
		.INIT('h2a)
	) name21680 (
		\m5_sel_i[3]_pad ,
		_w8655_,
		_w8656_,
		_w23581_
	);
	LUT3 #(
		.INIT('h2a)
	) name21681 (
		\m1_sel_i[3]_pad ,
		_w8655_,
		_w8656_,
		_w23582_
	);
	LUT4 #(
		.INIT('h57df)
	) name21682 (
		_w8650_,
		_w8653_,
		_w23581_,
		_w23582_,
		_w23583_
	);
	LUT3 #(
		.INIT('h80)
	) name21683 (
		\m0_sel_i[3]_pad ,
		_w8655_,
		_w8656_,
		_w23584_
	);
	LUT3 #(
		.INIT('h2a)
	) name21684 (
		\m7_sel_i[3]_pad ,
		_w8655_,
		_w8656_,
		_w23585_
	);
	LUT4 #(
		.INIT('h6e7f)
	) name21685 (
		_w8650_,
		_w8653_,
		_w23584_,
		_w23585_,
		_w23586_
	);
	LUT4 #(
		.INIT('h7fff)
	) name21686 (
		_w23577_,
		_w23580_,
		_w23583_,
		_w23586_,
		_w23587_
	);
	LUT4 #(
		.INIT('h2a00)
	) name21687 (
		\m3_stb_i_pad ,
		_w8655_,
		_w8656_,
		_w9500_,
		_w23588_
	);
	LUT4 #(
		.INIT('h8000)
	) name21688 (
		\m2_stb_i_pad ,
		_w8655_,
		_w8656_,
		_w9468_,
		_w23589_
	);
	LUT3 #(
		.INIT('h57)
	) name21689 (
		_w8668_,
		_w23588_,
		_w23589_,
		_w23590_
	);
	LUT4 #(
		.INIT('h8000)
	) name21690 (
		\m4_stb_i_pad ,
		_w8655_,
		_w8656_,
		_w9366_,
		_w23591_
	);
	LUT4 #(
		.INIT('h2a00)
	) name21691 (
		\m1_stb_i_pad ,
		_w8655_,
		_w8656_,
		_w9433_,
		_w23592_
	);
	LUT4 #(
		.INIT('h57df)
	) name21692 (
		_w8650_,
		_w8653_,
		_w23591_,
		_w23592_,
		_w23593_
	);
	LUT4 #(
		.INIT('h2a00)
	) name21693 (
		\m5_stb_i_pad ,
		_w8655_,
		_w8656_,
		_w9544_,
		_w23594_
	);
	LUT4 #(
		.INIT('h2a00)
	) name21694 (
		\m7_stb_i_pad ,
		_w8655_,
		_w8656_,
		_w9614_,
		_w23595_
	);
	LUT4 #(
		.INIT('hcedf)
	) name21695 (
		_w8650_,
		_w8653_,
		_w23594_,
		_w23595_,
		_w23596_
	);
	LUT4 #(
		.INIT('h8000)
	) name21696 (
		\m6_stb_i_pad ,
		_w8655_,
		_w8656_,
		_w9582_,
		_w23597_
	);
	LUT4 #(
		.INIT('h8000)
	) name21697 (
		\m0_stb_i_pad ,
		_w8655_,
		_w8656_,
		_w9644_,
		_w23598_
	);
	LUT4 #(
		.INIT('h67ef)
	) name21698 (
		_w8650_,
		_w8653_,
		_w23597_,
		_w23598_,
		_w23599_
	);
	LUT4 #(
		.INIT('h7fff)
	) name21699 (
		_w23590_,
		_w23593_,
		_w23596_,
		_w23599_,
		_w23600_
	);
	LUT3 #(
		.INIT('h2a)
	) name21700 (
		\m3_we_i_pad ,
		_w8655_,
		_w8656_,
		_w23601_
	);
	LUT3 #(
		.INIT('h80)
	) name21701 (
		\m4_we_i_pad ,
		_w8655_,
		_w8656_,
		_w23602_
	);
	LUT4 #(
		.INIT('h9dbf)
	) name21702 (
		_w8650_,
		_w8653_,
		_w23601_,
		_w23602_,
		_w23603_
	);
	LUT3 #(
		.INIT('h80)
	) name21703 (
		\m6_we_i_pad ,
		_w8655_,
		_w8656_,
		_w23604_
	);
	LUT3 #(
		.INIT('h80)
	) name21704 (
		\m2_we_i_pad ,
		_w8655_,
		_w8656_,
		_w23605_
	);
	LUT4 #(
		.INIT('habef)
	) name21705 (
		_w8650_,
		_w8653_,
		_w23604_,
		_w23605_,
		_w23606_
	);
	LUT3 #(
		.INIT('h2a)
	) name21706 (
		\m5_we_i_pad ,
		_w8655_,
		_w8656_,
		_w23607_
	);
	LUT3 #(
		.INIT('h2a)
	) name21707 (
		\m1_we_i_pad ,
		_w8655_,
		_w8656_,
		_w23608_
	);
	LUT4 #(
		.INIT('h57df)
	) name21708 (
		_w8650_,
		_w8653_,
		_w23607_,
		_w23608_,
		_w23609_
	);
	LUT3 #(
		.INIT('h80)
	) name21709 (
		\m0_we_i_pad ,
		_w8655_,
		_w8656_,
		_w23610_
	);
	LUT3 #(
		.INIT('h2a)
	) name21710 (
		\m7_we_i_pad ,
		_w8655_,
		_w8656_,
		_w23611_
	);
	LUT4 #(
		.INIT('h6e7f)
	) name21711 (
		_w8650_,
		_w8653_,
		_w23610_,
		_w23611_,
		_w23612_
	);
	LUT4 #(
		.INIT('h7fff)
	) name21712 (
		_w23603_,
		_w23606_,
		_w23609_,
		_w23612_,
		_w23613_
	);
	LUT3 #(
		.INIT('h2a)
	) name21713 (
		\m3_addr_i[0]_pad ,
		_w8699_,
		_w8700_,
		_w23614_
	);
	LUT3 #(
		.INIT('h80)
	) name21714 (
		\m4_addr_i[0]_pad ,
		_w8699_,
		_w8700_,
		_w23615_
	);
	LUT4 #(
		.INIT('h9dbf)
	) name21715 (
		_w8694_,
		_w8697_,
		_w23614_,
		_w23615_,
		_w23616_
	);
	LUT3 #(
		.INIT('h80)
	) name21716 (
		\m6_addr_i[0]_pad ,
		_w8699_,
		_w8700_,
		_w23617_
	);
	LUT3 #(
		.INIT('h2a)
	) name21717 (
		\m7_addr_i[0]_pad ,
		_w8699_,
		_w8700_,
		_w23618_
	);
	LUT3 #(
		.INIT('h57)
	) name21718 (
		_w8712_,
		_w23617_,
		_w23618_,
		_w23619_
	);
	LUT3 #(
		.INIT('h2a)
	) name21719 (
		\m5_addr_i[0]_pad ,
		_w8699_,
		_w8700_,
		_w23620_
	);
	LUT3 #(
		.INIT('h80)
	) name21720 (
		\m0_addr_i[0]_pad ,
		_w8699_,
		_w8700_,
		_w23621_
	);
	LUT4 #(
		.INIT('h57df)
	) name21721 (
		_w8694_,
		_w8697_,
		_w23620_,
		_w23621_,
		_w23622_
	);
	LUT3 #(
		.INIT('h2a)
	) name21722 (
		\m1_addr_i[0]_pad ,
		_w8699_,
		_w8700_,
		_w23623_
	);
	LUT3 #(
		.INIT('h80)
	) name21723 (
		\m2_addr_i[0]_pad ,
		_w8699_,
		_w8700_,
		_w23624_
	);
	LUT4 #(
		.INIT('h3b7f)
	) name21724 (
		_w8694_,
		_w8697_,
		_w23623_,
		_w23624_,
		_w23625_
	);
	LUT4 #(
		.INIT('h7fff)
	) name21725 (
		_w23616_,
		_w23619_,
		_w23622_,
		_w23625_,
		_w23626_
	);
	LUT3 #(
		.INIT('h2a)
	) name21726 (
		\m3_addr_i[10]_pad ,
		_w8699_,
		_w8700_,
		_w23627_
	);
	LUT3 #(
		.INIT('h80)
	) name21727 (
		\m4_addr_i[10]_pad ,
		_w8699_,
		_w8700_,
		_w23628_
	);
	LUT4 #(
		.INIT('h9dbf)
	) name21728 (
		_w8694_,
		_w8697_,
		_w23627_,
		_w23628_,
		_w23629_
	);
	LUT3 #(
		.INIT('h80)
	) name21729 (
		\m6_addr_i[10]_pad ,
		_w8699_,
		_w8700_,
		_w23630_
	);
	LUT3 #(
		.INIT('h80)
	) name21730 (
		\m2_addr_i[10]_pad ,
		_w8699_,
		_w8700_,
		_w23631_
	);
	LUT4 #(
		.INIT('habef)
	) name21731 (
		_w8694_,
		_w8697_,
		_w23630_,
		_w23631_,
		_w23632_
	);
	LUT3 #(
		.INIT('h2a)
	) name21732 (
		\m5_addr_i[10]_pad ,
		_w8699_,
		_w8700_,
		_w23633_
	);
	LUT3 #(
		.INIT('h2a)
	) name21733 (
		\m1_addr_i[10]_pad ,
		_w8699_,
		_w8700_,
		_w23634_
	);
	LUT4 #(
		.INIT('h57df)
	) name21734 (
		_w8694_,
		_w8697_,
		_w23633_,
		_w23634_,
		_w23635_
	);
	LUT3 #(
		.INIT('h80)
	) name21735 (
		\m0_addr_i[10]_pad ,
		_w8699_,
		_w8700_,
		_w23636_
	);
	LUT3 #(
		.INIT('h2a)
	) name21736 (
		\m7_addr_i[10]_pad ,
		_w8699_,
		_w8700_,
		_w23637_
	);
	LUT4 #(
		.INIT('h6e7f)
	) name21737 (
		_w8694_,
		_w8697_,
		_w23636_,
		_w23637_,
		_w23638_
	);
	LUT4 #(
		.INIT('h7fff)
	) name21738 (
		_w23629_,
		_w23632_,
		_w23635_,
		_w23638_,
		_w23639_
	);
	LUT3 #(
		.INIT('h2a)
	) name21739 (
		\m3_addr_i[11]_pad ,
		_w8699_,
		_w8700_,
		_w23640_
	);
	LUT3 #(
		.INIT('h80)
	) name21740 (
		\m4_addr_i[11]_pad ,
		_w8699_,
		_w8700_,
		_w23641_
	);
	LUT4 #(
		.INIT('h9dbf)
	) name21741 (
		_w8694_,
		_w8697_,
		_w23640_,
		_w23641_,
		_w23642_
	);
	LUT3 #(
		.INIT('h80)
	) name21742 (
		\m6_addr_i[11]_pad ,
		_w8699_,
		_w8700_,
		_w23643_
	);
	LUT3 #(
		.INIT('h80)
	) name21743 (
		\m2_addr_i[11]_pad ,
		_w8699_,
		_w8700_,
		_w23644_
	);
	LUT4 #(
		.INIT('habef)
	) name21744 (
		_w8694_,
		_w8697_,
		_w23643_,
		_w23644_,
		_w23645_
	);
	LUT3 #(
		.INIT('h2a)
	) name21745 (
		\m5_addr_i[11]_pad ,
		_w8699_,
		_w8700_,
		_w23646_
	);
	LUT3 #(
		.INIT('h2a)
	) name21746 (
		\m1_addr_i[11]_pad ,
		_w8699_,
		_w8700_,
		_w23647_
	);
	LUT4 #(
		.INIT('h57df)
	) name21747 (
		_w8694_,
		_w8697_,
		_w23646_,
		_w23647_,
		_w23648_
	);
	LUT3 #(
		.INIT('h80)
	) name21748 (
		\m0_addr_i[11]_pad ,
		_w8699_,
		_w8700_,
		_w23649_
	);
	LUT3 #(
		.INIT('h2a)
	) name21749 (
		\m7_addr_i[11]_pad ,
		_w8699_,
		_w8700_,
		_w23650_
	);
	LUT4 #(
		.INIT('h6e7f)
	) name21750 (
		_w8694_,
		_w8697_,
		_w23649_,
		_w23650_,
		_w23651_
	);
	LUT4 #(
		.INIT('h7fff)
	) name21751 (
		_w23642_,
		_w23645_,
		_w23648_,
		_w23651_,
		_w23652_
	);
	LUT3 #(
		.INIT('h80)
	) name21752 (
		\m6_addr_i[12]_pad ,
		_w8699_,
		_w8700_,
		_w23653_
	);
	LUT3 #(
		.INIT('h2a)
	) name21753 (
		\m5_addr_i[12]_pad ,
		_w8699_,
		_w8700_,
		_w23654_
	);
	LUT4 #(
		.INIT('hcdef)
	) name21754 (
		_w8694_,
		_w8697_,
		_w23653_,
		_w23654_,
		_w23655_
	);
	LUT3 #(
		.INIT('h2a)
	) name21755 (
		\m1_addr_i[12]_pad ,
		_w8699_,
		_w8700_,
		_w23656_
	);
	LUT3 #(
		.INIT('h80)
	) name21756 (
		\m4_addr_i[12]_pad ,
		_w8699_,
		_w8700_,
		_w23657_
	);
	LUT4 #(
		.INIT('h5d7f)
	) name21757 (
		_w8694_,
		_w8697_,
		_w23656_,
		_w23657_,
		_w23658_
	);
	LUT3 #(
		.INIT('h80)
	) name21758 (
		\m2_addr_i[12]_pad ,
		_w8699_,
		_w8700_,
		_w23659_
	);
	LUT3 #(
		.INIT('h2a)
	) name21759 (
		\m3_addr_i[12]_pad ,
		_w8699_,
		_w8700_,
		_w23660_
	);
	LUT3 #(
		.INIT('h57)
	) name21760 (
		_w8698_,
		_w23659_,
		_w23660_,
		_w23661_
	);
	LUT3 #(
		.INIT('h80)
	) name21761 (
		\m0_addr_i[12]_pad ,
		_w8699_,
		_w8700_,
		_w23662_
	);
	LUT3 #(
		.INIT('h2a)
	) name21762 (
		\m7_addr_i[12]_pad ,
		_w8699_,
		_w8700_,
		_w23663_
	);
	LUT4 #(
		.INIT('h6e7f)
	) name21763 (
		_w8694_,
		_w8697_,
		_w23662_,
		_w23663_,
		_w23664_
	);
	LUT4 #(
		.INIT('h7fff)
	) name21764 (
		_w23655_,
		_w23658_,
		_w23661_,
		_w23664_,
		_w23665_
	);
	LUT3 #(
		.INIT('h80)
	) name21765 (
		\m6_addr_i[13]_pad ,
		_w8699_,
		_w8700_,
		_w23666_
	);
	LUT3 #(
		.INIT('h2a)
	) name21766 (
		\m5_addr_i[13]_pad ,
		_w8699_,
		_w8700_,
		_w23667_
	);
	LUT4 #(
		.INIT('hcdef)
	) name21767 (
		_w8694_,
		_w8697_,
		_w23666_,
		_w23667_,
		_w23668_
	);
	LUT3 #(
		.INIT('h80)
	) name21768 (
		\m0_addr_i[13]_pad ,
		_w8699_,
		_w8700_,
		_w23669_
	);
	LUT3 #(
		.INIT('h80)
	) name21769 (
		\m4_addr_i[13]_pad ,
		_w8699_,
		_w8700_,
		_w23670_
	);
	LUT4 #(
		.INIT('h5d7f)
	) name21770 (
		_w8694_,
		_w8697_,
		_w23669_,
		_w23670_,
		_w23671_
	);
	LUT3 #(
		.INIT('h2a)
	) name21771 (
		\m7_addr_i[13]_pad ,
		_w8699_,
		_w8700_,
		_w23672_
	);
	LUT3 #(
		.INIT('h2a)
	) name21772 (
		\m3_addr_i[13]_pad ,
		_w8699_,
		_w8700_,
		_w23673_
	);
	LUT4 #(
		.INIT('habef)
	) name21773 (
		_w8694_,
		_w8697_,
		_w23672_,
		_w23673_,
		_w23674_
	);
	LUT3 #(
		.INIT('h2a)
	) name21774 (
		\m1_addr_i[13]_pad ,
		_w8699_,
		_w8700_,
		_w23675_
	);
	LUT3 #(
		.INIT('h80)
	) name21775 (
		\m2_addr_i[13]_pad ,
		_w8699_,
		_w8700_,
		_w23676_
	);
	LUT4 #(
		.INIT('h3b7f)
	) name21776 (
		_w8694_,
		_w8697_,
		_w23675_,
		_w23676_,
		_w23677_
	);
	LUT4 #(
		.INIT('h7fff)
	) name21777 (
		_w23668_,
		_w23671_,
		_w23674_,
		_w23677_,
		_w23678_
	);
	LUT3 #(
		.INIT('h2a)
	) name21778 (
		\m3_addr_i[14]_pad ,
		_w8699_,
		_w8700_,
		_w23679_
	);
	LUT3 #(
		.INIT('h80)
	) name21779 (
		\m4_addr_i[14]_pad ,
		_w8699_,
		_w8700_,
		_w23680_
	);
	LUT4 #(
		.INIT('h9dbf)
	) name21780 (
		_w8694_,
		_w8697_,
		_w23679_,
		_w23680_,
		_w23681_
	);
	LUT3 #(
		.INIT('h80)
	) name21781 (
		\m6_addr_i[14]_pad ,
		_w8699_,
		_w8700_,
		_w23682_
	);
	LUT3 #(
		.INIT('h80)
	) name21782 (
		\m2_addr_i[14]_pad ,
		_w8699_,
		_w8700_,
		_w23683_
	);
	LUT4 #(
		.INIT('habef)
	) name21783 (
		_w8694_,
		_w8697_,
		_w23682_,
		_w23683_,
		_w23684_
	);
	LUT3 #(
		.INIT('h2a)
	) name21784 (
		\m5_addr_i[14]_pad ,
		_w8699_,
		_w8700_,
		_w23685_
	);
	LUT3 #(
		.INIT('h2a)
	) name21785 (
		\m1_addr_i[14]_pad ,
		_w8699_,
		_w8700_,
		_w23686_
	);
	LUT4 #(
		.INIT('h57df)
	) name21786 (
		_w8694_,
		_w8697_,
		_w23685_,
		_w23686_,
		_w23687_
	);
	LUT3 #(
		.INIT('h80)
	) name21787 (
		\m0_addr_i[14]_pad ,
		_w8699_,
		_w8700_,
		_w23688_
	);
	LUT3 #(
		.INIT('h2a)
	) name21788 (
		\m7_addr_i[14]_pad ,
		_w8699_,
		_w8700_,
		_w23689_
	);
	LUT4 #(
		.INIT('h6e7f)
	) name21789 (
		_w8694_,
		_w8697_,
		_w23688_,
		_w23689_,
		_w23690_
	);
	LUT4 #(
		.INIT('h7fff)
	) name21790 (
		_w23681_,
		_w23684_,
		_w23687_,
		_w23690_,
		_w23691_
	);
	LUT3 #(
		.INIT('h80)
	) name21791 (
		\m6_addr_i[15]_pad ,
		_w8699_,
		_w8700_,
		_w23692_
	);
	LUT3 #(
		.INIT('h2a)
	) name21792 (
		\m5_addr_i[15]_pad ,
		_w8699_,
		_w8700_,
		_w23693_
	);
	LUT4 #(
		.INIT('hcdef)
	) name21793 (
		_w8694_,
		_w8697_,
		_w23692_,
		_w23693_,
		_w23694_
	);
	LUT3 #(
		.INIT('h2a)
	) name21794 (
		\m3_addr_i[15]_pad ,
		_w8699_,
		_w8700_,
		_w23695_
	);
	LUT3 #(
		.INIT('h80)
	) name21795 (
		\m2_addr_i[15]_pad ,
		_w8699_,
		_w8700_,
		_w23696_
	);
	LUT3 #(
		.INIT('h57)
	) name21796 (
		_w8698_,
		_w23695_,
		_w23696_,
		_w23697_
	);
	LUT3 #(
		.INIT('h80)
	) name21797 (
		\m4_addr_i[15]_pad ,
		_w8699_,
		_w8700_,
		_w23698_
	);
	LUT3 #(
		.INIT('h2a)
	) name21798 (
		\m1_addr_i[15]_pad ,
		_w8699_,
		_w8700_,
		_w23699_
	);
	LUT4 #(
		.INIT('h57df)
	) name21799 (
		_w8694_,
		_w8697_,
		_w23698_,
		_w23699_,
		_w23700_
	);
	LUT3 #(
		.INIT('h80)
	) name21800 (
		\m0_addr_i[15]_pad ,
		_w8699_,
		_w8700_,
		_w23701_
	);
	LUT3 #(
		.INIT('h2a)
	) name21801 (
		\m7_addr_i[15]_pad ,
		_w8699_,
		_w8700_,
		_w23702_
	);
	LUT4 #(
		.INIT('h6e7f)
	) name21802 (
		_w8694_,
		_w8697_,
		_w23701_,
		_w23702_,
		_w23703_
	);
	LUT4 #(
		.INIT('h7fff)
	) name21803 (
		_w23694_,
		_w23697_,
		_w23700_,
		_w23703_,
		_w23704_
	);
	LUT3 #(
		.INIT('h2a)
	) name21804 (
		\m3_addr_i[16]_pad ,
		_w8699_,
		_w8700_,
		_w23705_
	);
	LUT3 #(
		.INIT('h80)
	) name21805 (
		\m4_addr_i[16]_pad ,
		_w8699_,
		_w8700_,
		_w23706_
	);
	LUT4 #(
		.INIT('h9dbf)
	) name21806 (
		_w8694_,
		_w8697_,
		_w23705_,
		_w23706_,
		_w23707_
	);
	LUT3 #(
		.INIT('h80)
	) name21807 (
		\m6_addr_i[16]_pad ,
		_w8699_,
		_w8700_,
		_w23708_
	);
	LUT3 #(
		.INIT('h80)
	) name21808 (
		\m2_addr_i[16]_pad ,
		_w8699_,
		_w8700_,
		_w23709_
	);
	LUT4 #(
		.INIT('habef)
	) name21809 (
		_w8694_,
		_w8697_,
		_w23708_,
		_w23709_,
		_w23710_
	);
	LUT3 #(
		.INIT('h2a)
	) name21810 (
		\m5_addr_i[16]_pad ,
		_w8699_,
		_w8700_,
		_w23711_
	);
	LUT3 #(
		.INIT('h2a)
	) name21811 (
		\m1_addr_i[16]_pad ,
		_w8699_,
		_w8700_,
		_w23712_
	);
	LUT4 #(
		.INIT('h57df)
	) name21812 (
		_w8694_,
		_w8697_,
		_w23711_,
		_w23712_,
		_w23713_
	);
	LUT3 #(
		.INIT('h80)
	) name21813 (
		\m0_addr_i[16]_pad ,
		_w8699_,
		_w8700_,
		_w23714_
	);
	LUT3 #(
		.INIT('h2a)
	) name21814 (
		\m7_addr_i[16]_pad ,
		_w8699_,
		_w8700_,
		_w23715_
	);
	LUT4 #(
		.INIT('h6e7f)
	) name21815 (
		_w8694_,
		_w8697_,
		_w23714_,
		_w23715_,
		_w23716_
	);
	LUT4 #(
		.INIT('h7fff)
	) name21816 (
		_w23707_,
		_w23710_,
		_w23713_,
		_w23716_,
		_w23717_
	);
	LUT3 #(
		.INIT('h80)
	) name21817 (
		\m6_addr_i[17]_pad ,
		_w8699_,
		_w8700_,
		_w23718_
	);
	LUT3 #(
		.INIT('h2a)
	) name21818 (
		\m5_addr_i[17]_pad ,
		_w8699_,
		_w8700_,
		_w23719_
	);
	LUT4 #(
		.INIT('hcdef)
	) name21819 (
		_w8694_,
		_w8697_,
		_w23718_,
		_w23719_,
		_w23720_
	);
	LUT3 #(
		.INIT('h2a)
	) name21820 (
		\m1_addr_i[17]_pad ,
		_w8699_,
		_w8700_,
		_w23721_
	);
	LUT3 #(
		.INIT('h80)
	) name21821 (
		\m4_addr_i[17]_pad ,
		_w8699_,
		_w8700_,
		_w23722_
	);
	LUT4 #(
		.INIT('h5d7f)
	) name21822 (
		_w8694_,
		_w8697_,
		_w23721_,
		_w23722_,
		_w23723_
	);
	LUT3 #(
		.INIT('h80)
	) name21823 (
		\m2_addr_i[17]_pad ,
		_w8699_,
		_w8700_,
		_w23724_
	);
	LUT3 #(
		.INIT('h2a)
	) name21824 (
		\m3_addr_i[17]_pad ,
		_w8699_,
		_w8700_,
		_w23725_
	);
	LUT3 #(
		.INIT('h57)
	) name21825 (
		_w8698_,
		_w23724_,
		_w23725_,
		_w23726_
	);
	LUT3 #(
		.INIT('h80)
	) name21826 (
		\m0_addr_i[17]_pad ,
		_w8699_,
		_w8700_,
		_w23727_
	);
	LUT3 #(
		.INIT('h2a)
	) name21827 (
		\m7_addr_i[17]_pad ,
		_w8699_,
		_w8700_,
		_w23728_
	);
	LUT4 #(
		.INIT('h6e7f)
	) name21828 (
		_w8694_,
		_w8697_,
		_w23727_,
		_w23728_,
		_w23729_
	);
	LUT4 #(
		.INIT('h7fff)
	) name21829 (
		_w23720_,
		_w23723_,
		_w23726_,
		_w23729_,
		_w23730_
	);
	LUT3 #(
		.INIT('h2a)
	) name21830 (
		\m3_addr_i[18]_pad ,
		_w8699_,
		_w8700_,
		_w23731_
	);
	LUT3 #(
		.INIT('h80)
	) name21831 (
		\m4_addr_i[18]_pad ,
		_w8699_,
		_w8700_,
		_w23732_
	);
	LUT4 #(
		.INIT('h9dbf)
	) name21832 (
		_w8694_,
		_w8697_,
		_w23731_,
		_w23732_,
		_w23733_
	);
	LUT3 #(
		.INIT('h80)
	) name21833 (
		\m6_addr_i[18]_pad ,
		_w8699_,
		_w8700_,
		_w23734_
	);
	LUT3 #(
		.INIT('h80)
	) name21834 (
		\m2_addr_i[18]_pad ,
		_w8699_,
		_w8700_,
		_w23735_
	);
	LUT4 #(
		.INIT('habef)
	) name21835 (
		_w8694_,
		_w8697_,
		_w23734_,
		_w23735_,
		_w23736_
	);
	LUT3 #(
		.INIT('h2a)
	) name21836 (
		\m5_addr_i[18]_pad ,
		_w8699_,
		_w8700_,
		_w23737_
	);
	LUT3 #(
		.INIT('h2a)
	) name21837 (
		\m1_addr_i[18]_pad ,
		_w8699_,
		_w8700_,
		_w23738_
	);
	LUT4 #(
		.INIT('h57df)
	) name21838 (
		_w8694_,
		_w8697_,
		_w23737_,
		_w23738_,
		_w23739_
	);
	LUT3 #(
		.INIT('h80)
	) name21839 (
		\m0_addr_i[18]_pad ,
		_w8699_,
		_w8700_,
		_w23740_
	);
	LUT3 #(
		.INIT('h2a)
	) name21840 (
		\m7_addr_i[18]_pad ,
		_w8699_,
		_w8700_,
		_w23741_
	);
	LUT4 #(
		.INIT('h6e7f)
	) name21841 (
		_w8694_,
		_w8697_,
		_w23740_,
		_w23741_,
		_w23742_
	);
	LUT4 #(
		.INIT('h7fff)
	) name21842 (
		_w23733_,
		_w23736_,
		_w23739_,
		_w23742_,
		_w23743_
	);
	LUT3 #(
		.INIT('h2a)
	) name21843 (
		\m3_addr_i[19]_pad ,
		_w8699_,
		_w8700_,
		_w23744_
	);
	LUT3 #(
		.INIT('h80)
	) name21844 (
		\m4_addr_i[19]_pad ,
		_w8699_,
		_w8700_,
		_w23745_
	);
	LUT4 #(
		.INIT('h9dbf)
	) name21845 (
		_w8694_,
		_w8697_,
		_w23744_,
		_w23745_,
		_w23746_
	);
	LUT3 #(
		.INIT('h80)
	) name21846 (
		\m6_addr_i[19]_pad ,
		_w8699_,
		_w8700_,
		_w23747_
	);
	LUT3 #(
		.INIT('h80)
	) name21847 (
		\m2_addr_i[19]_pad ,
		_w8699_,
		_w8700_,
		_w23748_
	);
	LUT4 #(
		.INIT('habef)
	) name21848 (
		_w8694_,
		_w8697_,
		_w23747_,
		_w23748_,
		_w23749_
	);
	LUT3 #(
		.INIT('h2a)
	) name21849 (
		\m5_addr_i[19]_pad ,
		_w8699_,
		_w8700_,
		_w23750_
	);
	LUT3 #(
		.INIT('h2a)
	) name21850 (
		\m1_addr_i[19]_pad ,
		_w8699_,
		_w8700_,
		_w23751_
	);
	LUT4 #(
		.INIT('h57df)
	) name21851 (
		_w8694_,
		_w8697_,
		_w23750_,
		_w23751_,
		_w23752_
	);
	LUT3 #(
		.INIT('h80)
	) name21852 (
		\m0_addr_i[19]_pad ,
		_w8699_,
		_w8700_,
		_w23753_
	);
	LUT3 #(
		.INIT('h2a)
	) name21853 (
		\m7_addr_i[19]_pad ,
		_w8699_,
		_w8700_,
		_w23754_
	);
	LUT4 #(
		.INIT('h6e7f)
	) name21854 (
		_w8694_,
		_w8697_,
		_w23753_,
		_w23754_,
		_w23755_
	);
	LUT4 #(
		.INIT('h7fff)
	) name21855 (
		_w23746_,
		_w23749_,
		_w23752_,
		_w23755_,
		_w23756_
	);
	LUT3 #(
		.INIT('h2a)
	) name21856 (
		\m3_addr_i[1]_pad ,
		_w8699_,
		_w8700_,
		_w23757_
	);
	LUT3 #(
		.INIT('h80)
	) name21857 (
		\m4_addr_i[1]_pad ,
		_w8699_,
		_w8700_,
		_w23758_
	);
	LUT4 #(
		.INIT('h9dbf)
	) name21858 (
		_w8694_,
		_w8697_,
		_w23757_,
		_w23758_,
		_w23759_
	);
	LUT3 #(
		.INIT('h80)
	) name21859 (
		\m6_addr_i[1]_pad ,
		_w8699_,
		_w8700_,
		_w23760_
	);
	LUT3 #(
		.INIT('h80)
	) name21860 (
		\m2_addr_i[1]_pad ,
		_w8699_,
		_w8700_,
		_w23761_
	);
	LUT4 #(
		.INIT('habef)
	) name21861 (
		_w8694_,
		_w8697_,
		_w23760_,
		_w23761_,
		_w23762_
	);
	LUT3 #(
		.INIT('h2a)
	) name21862 (
		\m5_addr_i[1]_pad ,
		_w8699_,
		_w8700_,
		_w23763_
	);
	LUT3 #(
		.INIT('h2a)
	) name21863 (
		\m1_addr_i[1]_pad ,
		_w8699_,
		_w8700_,
		_w23764_
	);
	LUT4 #(
		.INIT('h57df)
	) name21864 (
		_w8694_,
		_w8697_,
		_w23763_,
		_w23764_,
		_w23765_
	);
	LUT3 #(
		.INIT('h80)
	) name21865 (
		\m0_addr_i[1]_pad ,
		_w8699_,
		_w8700_,
		_w23766_
	);
	LUT3 #(
		.INIT('h2a)
	) name21866 (
		\m7_addr_i[1]_pad ,
		_w8699_,
		_w8700_,
		_w23767_
	);
	LUT4 #(
		.INIT('h6e7f)
	) name21867 (
		_w8694_,
		_w8697_,
		_w23766_,
		_w23767_,
		_w23768_
	);
	LUT4 #(
		.INIT('h7fff)
	) name21868 (
		_w23759_,
		_w23762_,
		_w23765_,
		_w23768_,
		_w23769_
	);
	LUT3 #(
		.INIT('h2a)
	) name21869 (
		\m3_addr_i[20]_pad ,
		_w8699_,
		_w8700_,
		_w23770_
	);
	LUT3 #(
		.INIT('h80)
	) name21870 (
		\m4_addr_i[20]_pad ,
		_w8699_,
		_w8700_,
		_w23771_
	);
	LUT4 #(
		.INIT('h9dbf)
	) name21871 (
		_w8694_,
		_w8697_,
		_w23770_,
		_w23771_,
		_w23772_
	);
	LUT3 #(
		.INIT('h80)
	) name21872 (
		\m6_addr_i[20]_pad ,
		_w8699_,
		_w8700_,
		_w23773_
	);
	LUT3 #(
		.INIT('h80)
	) name21873 (
		\m2_addr_i[20]_pad ,
		_w8699_,
		_w8700_,
		_w23774_
	);
	LUT4 #(
		.INIT('habef)
	) name21874 (
		_w8694_,
		_w8697_,
		_w23773_,
		_w23774_,
		_w23775_
	);
	LUT3 #(
		.INIT('h2a)
	) name21875 (
		\m5_addr_i[20]_pad ,
		_w8699_,
		_w8700_,
		_w23776_
	);
	LUT3 #(
		.INIT('h2a)
	) name21876 (
		\m1_addr_i[20]_pad ,
		_w8699_,
		_w8700_,
		_w23777_
	);
	LUT4 #(
		.INIT('h57df)
	) name21877 (
		_w8694_,
		_w8697_,
		_w23776_,
		_w23777_,
		_w23778_
	);
	LUT3 #(
		.INIT('h80)
	) name21878 (
		\m0_addr_i[20]_pad ,
		_w8699_,
		_w8700_,
		_w23779_
	);
	LUT3 #(
		.INIT('h2a)
	) name21879 (
		\m7_addr_i[20]_pad ,
		_w8699_,
		_w8700_,
		_w23780_
	);
	LUT4 #(
		.INIT('h6e7f)
	) name21880 (
		_w8694_,
		_w8697_,
		_w23779_,
		_w23780_,
		_w23781_
	);
	LUT4 #(
		.INIT('h7fff)
	) name21881 (
		_w23772_,
		_w23775_,
		_w23778_,
		_w23781_,
		_w23782_
	);
	LUT3 #(
		.INIT('h2a)
	) name21882 (
		\m3_addr_i[21]_pad ,
		_w8699_,
		_w8700_,
		_w23783_
	);
	LUT3 #(
		.INIT('h80)
	) name21883 (
		\m4_addr_i[21]_pad ,
		_w8699_,
		_w8700_,
		_w23784_
	);
	LUT4 #(
		.INIT('h9dbf)
	) name21884 (
		_w8694_,
		_w8697_,
		_w23783_,
		_w23784_,
		_w23785_
	);
	LUT3 #(
		.INIT('h80)
	) name21885 (
		\m6_addr_i[21]_pad ,
		_w8699_,
		_w8700_,
		_w23786_
	);
	LUT3 #(
		.INIT('h80)
	) name21886 (
		\m2_addr_i[21]_pad ,
		_w8699_,
		_w8700_,
		_w23787_
	);
	LUT4 #(
		.INIT('habef)
	) name21887 (
		_w8694_,
		_w8697_,
		_w23786_,
		_w23787_,
		_w23788_
	);
	LUT3 #(
		.INIT('h2a)
	) name21888 (
		\m5_addr_i[21]_pad ,
		_w8699_,
		_w8700_,
		_w23789_
	);
	LUT3 #(
		.INIT('h2a)
	) name21889 (
		\m1_addr_i[21]_pad ,
		_w8699_,
		_w8700_,
		_w23790_
	);
	LUT4 #(
		.INIT('h57df)
	) name21890 (
		_w8694_,
		_w8697_,
		_w23789_,
		_w23790_,
		_w23791_
	);
	LUT3 #(
		.INIT('h80)
	) name21891 (
		\m0_addr_i[21]_pad ,
		_w8699_,
		_w8700_,
		_w23792_
	);
	LUT3 #(
		.INIT('h2a)
	) name21892 (
		\m7_addr_i[21]_pad ,
		_w8699_,
		_w8700_,
		_w23793_
	);
	LUT4 #(
		.INIT('h6e7f)
	) name21893 (
		_w8694_,
		_w8697_,
		_w23792_,
		_w23793_,
		_w23794_
	);
	LUT4 #(
		.INIT('h7fff)
	) name21894 (
		_w23785_,
		_w23788_,
		_w23791_,
		_w23794_,
		_w23795_
	);
	LUT3 #(
		.INIT('h80)
	) name21895 (
		\m0_addr_i[22]_pad ,
		_w8699_,
		_w8700_,
		_w23796_
	);
	LUT3 #(
		.INIT('h2a)
	) name21896 (
		\m7_addr_i[22]_pad ,
		_w8699_,
		_w8700_,
		_w23797_
	);
	LUT4 #(
		.INIT('h6e7f)
	) name21897 (
		_w8694_,
		_w8697_,
		_w23796_,
		_w23797_,
		_w23798_
	);
	LUT3 #(
		.INIT('h80)
	) name21898 (
		\m6_addr_i[22]_pad ,
		_w8699_,
		_w8700_,
		_w23799_
	);
	LUT3 #(
		.INIT('h80)
	) name21899 (
		\m2_addr_i[22]_pad ,
		_w8699_,
		_w8700_,
		_w23800_
	);
	LUT4 #(
		.INIT('habef)
	) name21900 (
		_w8694_,
		_w8697_,
		_w23799_,
		_w23800_,
		_w23801_
	);
	LUT3 #(
		.INIT('h2a)
	) name21901 (
		\m5_addr_i[22]_pad ,
		_w8699_,
		_w8700_,
		_w23802_
	);
	LUT3 #(
		.INIT('h2a)
	) name21902 (
		\m1_addr_i[22]_pad ,
		_w8699_,
		_w8700_,
		_w23803_
	);
	LUT4 #(
		.INIT('h57df)
	) name21903 (
		_w8694_,
		_w8697_,
		_w23802_,
		_w23803_,
		_w23804_
	);
	LUT3 #(
		.INIT('h2a)
	) name21904 (
		\m3_addr_i[22]_pad ,
		_w8699_,
		_w8700_,
		_w23805_
	);
	LUT3 #(
		.INIT('h80)
	) name21905 (
		\m4_addr_i[22]_pad ,
		_w8699_,
		_w8700_,
		_w23806_
	);
	LUT4 #(
		.INIT('h9dbf)
	) name21906 (
		_w8694_,
		_w8697_,
		_w23805_,
		_w23806_,
		_w23807_
	);
	LUT4 #(
		.INIT('h7fff)
	) name21907 (
		_w23798_,
		_w23801_,
		_w23804_,
		_w23807_,
		_w23808_
	);
	LUT3 #(
		.INIT('h2a)
	) name21908 (
		\m3_addr_i[23]_pad ,
		_w8699_,
		_w8700_,
		_w23809_
	);
	LUT3 #(
		.INIT('h80)
	) name21909 (
		\m4_addr_i[23]_pad ,
		_w8699_,
		_w8700_,
		_w23810_
	);
	LUT4 #(
		.INIT('h9dbf)
	) name21910 (
		_w8694_,
		_w8697_,
		_w23809_,
		_w23810_,
		_w23811_
	);
	LUT3 #(
		.INIT('h80)
	) name21911 (
		\m6_addr_i[23]_pad ,
		_w8699_,
		_w8700_,
		_w23812_
	);
	LUT3 #(
		.INIT('h80)
	) name21912 (
		\m2_addr_i[23]_pad ,
		_w8699_,
		_w8700_,
		_w23813_
	);
	LUT4 #(
		.INIT('habef)
	) name21913 (
		_w8694_,
		_w8697_,
		_w23812_,
		_w23813_,
		_w23814_
	);
	LUT3 #(
		.INIT('h2a)
	) name21914 (
		\m5_addr_i[23]_pad ,
		_w8699_,
		_w8700_,
		_w23815_
	);
	LUT3 #(
		.INIT('h2a)
	) name21915 (
		\m1_addr_i[23]_pad ,
		_w8699_,
		_w8700_,
		_w23816_
	);
	LUT4 #(
		.INIT('h57df)
	) name21916 (
		_w8694_,
		_w8697_,
		_w23815_,
		_w23816_,
		_w23817_
	);
	LUT3 #(
		.INIT('h80)
	) name21917 (
		\m0_addr_i[23]_pad ,
		_w8699_,
		_w8700_,
		_w23818_
	);
	LUT3 #(
		.INIT('h2a)
	) name21918 (
		\m7_addr_i[23]_pad ,
		_w8699_,
		_w8700_,
		_w23819_
	);
	LUT4 #(
		.INIT('h6e7f)
	) name21919 (
		_w8694_,
		_w8697_,
		_w23818_,
		_w23819_,
		_w23820_
	);
	LUT4 #(
		.INIT('h7fff)
	) name21920 (
		_w23811_,
		_w23814_,
		_w23817_,
		_w23820_,
		_w23821_
	);
	LUT3 #(
		.INIT('h2a)
	) name21921 (
		\m3_addr_i[24]_pad ,
		_w8699_,
		_w8700_,
		_w23822_
	);
	LUT3 #(
		.INIT('h80)
	) name21922 (
		\m4_addr_i[24]_pad ,
		_w8699_,
		_w8700_,
		_w23823_
	);
	LUT4 #(
		.INIT('h9dbf)
	) name21923 (
		_w8694_,
		_w8697_,
		_w23822_,
		_w23823_,
		_w23824_
	);
	LUT3 #(
		.INIT('h2a)
	) name21924 (
		\m5_addr_i[24]_pad ,
		_w8699_,
		_w8700_,
		_w23825_
	);
	LUT3 #(
		.INIT('h80)
	) name21925 (
		\m2_addr_i[24]_pad ,
		_w8699_,
		_w8700_,
		_w23826_
	);
	LUT4 #(
		.INIT('h9bdf)
	) name21926 (
		_w8694_,
		_w8697_,
		_w23825_,
		_w23826_,
		_w23827_
	);
	LUT3 #(
		.INIT('h80)
	) name21927 (
		\m6_addr_i[24]_pad ,
		_w8699_,
		_w8700_,
		_w23828_
	);
	LUT3 #(
		.INIT('h2a)
	) name21928 (
		\m1_addr_i[24]_pad ,
		_w8699_,
		_w8700_,
		_w23829_
	);
	LUT4 #(
		.INIT('h67ef)
	) name21929 (
		_w8694_,
		_w8697_,
		_w23828_,
		_w23829_,
		_w23830_
	);
	LUT3 #(
		.INIT('h80)
	) name21930 (
		\m0_addr_i[24]_pad ,
		_w8699_,
		_w8700_,
		_w23831_
	);
	LUT3 #(
		.INIT('h2a)
	) name21931 (
		\m7_addr_i[24]_pad ,
		_w8699_,
		_w8700_,
		_w23832_
	);
	LUT4 #(
		.INIT('h6e7f)
	) name21932 (
		_w8694_,
		_w8697_,
		_w23831_,
		_w23832_,
		_w23833_
	);
	LUT4 #(
		.INIT('h7fff)
	) name21933 (
		_w23824_,
		_w23827_,
		_w23830_,
		_w23833_,
		_w23834_
	);
	LUT3 #(
		.INIT('h2a)
	) name21934 (
		\m5_addr_i[25]_pad ,
		_w8699_,
		_w8700_,
		_w23835_
	);
	LUT3 #(
		.INIT('h80)
	) name21935 (
		\m6_addr_i[25]_pad ,
		_w8699_,
		_w8700_,
		_w23836_
	);
	LUT4 #(
		.INIT('hcedf)
	) name21936 (
		_w8694_,
		_w8697_,
		_w23835_,
		_w23836_,
		_w23837_
	);
	LUT3 #(
		.INIT('h80)
	) name21937 (
		\m0_addr_i[25]_pad ,
		_w8699_,
		_w8700_,
		_w23838_
	);
	LUT3 #(
		.INIT('h80)
	) name21938 (
		\m4_addr_i[25]_pad ,
		_w8699_,
		_w8700_,
		_w23839_
	);
	LUT4 #(
		.INIT('h5d7f)
	) name21939 (
		_w8694_,
		_w8697_,
		_w23838_,
		_w23839_,
		_w23840_
	);
	LUT3 #(
		.INIT('h2a)
	) name21940 (
		\m7_addr_i[25]_pad ,
		_w8699_,
		_w8700_,
		_w23841_
	);
	LUT3 #(
		.INIT('h2a)
	) name21941 (
		\m3_addr_i[25]_pad ,
		_w8699_,
		_w8700_,
		_w23842_
	);
	LUT4 #(
		.INIT('habef)
	) name21942 (
		_w8694_,
		_w8697_,
		_w23841_,
		_w23842_,
		_w23843_
	);
	LUT3 #(
		.INIT('h2a)
	) name21943 (
		\m1_addr_i[25]_pad ,
		_w8699_,
		_w8700_,
		_w23844_
	);
	LUT3 #(
		.INIT('h80)
	) name21944 (
		\m2_addr_i[25]_pad ,
		_w8699_,
		_w8700_,
		_w23845_
	);
	LUT4 #(
		.INIT('h3b7f)
	) name21945 (
		_w8694_,
		_w8697_,
		_w23844_,
		_w23845_,
		_w23846_
	);
	LUT4 #(
		.INIT('h7fff)
	) name21946 (
		_w23837_,
		_w23840_,
		_w23843_,
		_w23846_,
		_w23847_
	);
	LUT3 #(
		.INIT('h2a)
	) name21947 (
		\m5_addr_i[26]_pad ,
		_w8699_,
		_w8700_,
		_w23848_
	);
	LUT3 #(
		.INIT('h80)
	) name21948 (
		\m6_addr_i[26]_pad ,
		_w8699_,
		_w8700_,
		_w23849_
	);
	LUT4 #(
		.INIT('hcedf)
	) name21949 (
		_w8694_,
		_w8697_,
		_w23848_,
		_w23849_,
		_w23850_
	);
	LUT3 #(
		.INIT('h2a)
	) name21950 (
		\m1_addr_i[26]_pad ,
		_w8699_,
		_w8700_,
		_w23851_
	);
	LUT3 #(
		.INIT('h80)
	) name21951 (
		\m4_addr_i[26]_pad ,
		_w8699_,
		_w8700_,
		_w23852_
	);
	LUT4 #(
		.INIT('h5d7f)
	) name21952 (
		_w8694_,
		_w8697_,
		_w23851_,
		_w23852_,
		_w23853_
	);
	LUT3 #(
		.INIT('h80)
	) name21953 (
		\m2_addr_i[26]_pad ,
		_w8699_,
		_w8700_,
		_w23854_
	);
	LUT3 #(
		.INIT('h2a)
	) name21954 (
		\m3_addr_i[26]_pad ,
		_w8699_,
		_w8700_,
		_w23855_
	);
	LUT3 #(
		.INIT('h57)
	) name21955 (
		_w8698_,
		_w23854_,
		_w23855_,
		_w23856_
	);
	LUT3 #(
		.INIT('h80)
	) name21956 (
		\m0_addr_i[26]_pad ,
		_w8699_,
		_w8700_,
		_w23857_
	);
	LUT3 #(
		.INIT('h2a)
	) name21957 (
		\m7_addr_i[26]_pad ,
		_w8699_,
		_w8700_,
		_w23858_
	);
	LUT4 #(
		.INIT('h6e7f)
	) name21958 (
		_w8694_,
		_w8697_,
		_w23857_,
		_w23858_,
		_w23859_
	);
	LUT4 #(
		.INIT('h7fff)
	) name21959 (
		_w23850_,
		_w23853_,
		_w23856_,
		_w23859_,
		_w23860_
	);
	LUT3 #(
		.INIT('h2a)
	) name21960 (
		\m3_addr_i[27]_pad ,
		_w8699_,
		_w8700_,
		_w23861_
	);
	LUT3 #(
		.INIT('h80)
	) name21961 (
		\m4_addr_i[27]_pad ,
		_w8699_,
		_w8700_,
		_w23862_
	);
	LUT4 #(
		.INIT('h9dbf)
	) name21962 (
		_w8694_,
		_w8697_,
		_w23861_,
		_w23862_,
		_w23863_
	);
	LUT3 #(
		.INIT('h80)
	) name21963 (
		\m0_addr_i[27]_pad ,
		_w8699_,
		_w8700_,
		_w23864_
	);
	LUT3 #(
		.INIT('h80)
	) name21964 (
		\m6_addr_i[27]_pad ,
		_w8699_,
		_w8700_,
		_w23865_
	);
	LUT4 #(
		.INIT('h6e7f)
	) name21965 (
		_w8694_,
		_w8697_,
		_w23864_,
		_w23865_,
		_w23866_
	);
	LUT3 #(
		.INIT('h2a)
	) name21966 (
		\m7_addr_i[27]_pad ,
		_w8699_,
		_w8700_,
		_w23867_
	);
	LUT3 #(
		.INIT('h2a)
	) name21967 (
		\m5_addr_i[27]_pad ,
		_w8699_,
		_w8700_,
		_w23868_
	);
	LUT4 #(
		.INIT('hcdef)
	) name21968 (
		_w8694_,
		_w8697_,
		_w23867_,
		_w23868_,
		_w23869_
	);
	LUT3 #(
		.INIT('h2a)
	) name21969 (
		\m1_addr_i[27]_pad ,
		_w8699_,
		_w8700_,
		_w23870_
	);
	LUT3 #(
		.INIT('h80)
	) name21970 (
		\m2_addr_i[27]_pad ,
		_w8699_,
		_w8700_,
		_w23871_
	);
	LUT4 #(
		.INIT('h3b7f)
	) name21971 (
		_w8694_,
		_w8697_,
		_w23870_,
		_w23871_,
		_w23872_
	);
	LUT4 #(
		.INIT('h7fff)
	) name21972 (
		_w23863_,
		_w23866_,
		_w23869_,
		_w23872_,
		_w23873_
	);
	LUT3 #(
		.INIT('h2a)
	) name21973 (
		\m3_addr_i[28]_pad ,
		_w8699_,
		_w8700_,
		_w23874_
	);
	LUT3 #(
		.INIT('h80)
	) name21974 (
		\m4_addr_i[28]_pad ,
		_w8699_,
		_w8700_,
		_w23875_
	);
	LUT4 #(
		.INIT('h9dbf)
	) name21975 (
		_w8694_,
		_w8697_,
		_w23874_,
		_w23875_,
		_w23876_
	);
	LUT3 #(
		.INIT('h2a)
	) name21976 (
		\m1_addr_i[28]_pad ,
		_w8699_,
		_w8700_,
		_w23877_
	);
	LUT3 #(
		.INIT('h2a)
	) name21977 (
		\m7_addr_i[28]_pad ,
		_w8699_,
		_w8700_,
		_w23878_
	);
	LUT4 #(
		.INIT('h6e7f)
	) name21978 (
		_w8694_,
		_w8697_,
		_w23877_,
		_w23878_,
		_w23879_
	);
	LUT3 #(
		.INIT('h80)
	) name21979 (
		\m2_addr_i[28]_pad ,
		_w8699_,
		_w8700_,
		_w23880_
	);
	LUT3 #(
		.INIT('h80)
	) name21980 (
		\m0_addr_i[28]_pad ,
		_w8699_,
		_w8700_,
		_w23881_
	);
	LUT4 #(
		.INIT('h37bf)
	) name21981 (
		_w8694_,
		_w8697_,
		_w23880_,
		_w23881_,
		_w23882_
	);
	LUT3 #(
		.INIT('h2a)
	) name21982 (
		\m5_addr_i[28]_pad ,
		_w8699_,
		_w8700_,
		_w23883_
	);
	LUT3 #(
		.INIT('h80)
	) name21983 (
		\m6_addr_i[28]_pad ,
		_w8699_,
		_w8700_,
		_w23884_
	);
	LUT4 #(
		.INIT('hcedf)
	) name21984 (
		_w8694_,
		_w8697_,
		_w23883_,
		_w23884_,
		_w23885_
	);
	LUT4 #(
		.INIT('h7fff)
	) name21985 (
		_w23876_,
		_w23879_,
		_w23882_,
		_w23885_,
		_w23886_
	);
	LUT3 #(
		.INIT('h2a)
	) name21986 (
		\m5_addr_i[29]_pad ,
		_w8699_,
		_w8700_,
		_w23887_
	);
	LUT3 #(
		.INIT('h80)
	) name21987 (
		\m6_addr_i[29]_pad ,
		_w8699_,
		_w8700_,
		_w23888_
	);
	LUT4 #(
		.INIT('hcedf)
	) name21988 (
		_w8694_,
		_w8697_,
		_w23887_,
		_w23888_,
		_w23889_
	);
	LUT3 #(
		.INIT('h80)
	) name21989 (
		\m0_addr_i[29]_pad ,
		_w8699_,
		_w8700_,
		_w23890_
	);
	LUT3 #(
		.INIT('h80)
	) name21990 (
		\m4_addr_i[29]_pad ,
		_w8699_,
		_w8700_,
		_w23891_
	);
	LUT4 #(
		.INIT('h5d7f)
	) name21991 (
		_w8694_,
		_w8697_,
		_w23890_,
		_w23891_,
		_w23892_
	);
	LUT3 #(
		.INIT('h2a)
	) name21992 (
		\m7_addr_i[29]_pad ,
		_w8699_,
		_w8700_,
		_w23893_
	);
	LUT3 #(
		.INIT('h2a)
	) name21993 (
		\m3_addr_i[29]_pad ,
		_w8699_,
		_w8700_,
		_w23894_
	);
	LUT4 #(
		.INIT('habef)
	) name21994 (
		_w8694_,
		_w8697_,
		_w23893_,
		_w23894_,
		_w23895_
	);
	LUT3 #(
		.INIT('h2a)
	) name21995 (
		\m1_addr_i[29]_pad ,
		_w8699_,
		_w8700_,
		_w23896_
	);
	LUT3 #(
		.INIT('h80)
	) name21996 (
		\m2_addr_i[29]_pad ,
		_w8699_,
		_w8700_,
		_w23897_
	);
	LUT4 #(
		.INIT('h3b7f)
	) name21997 (
		_w8694_,
		_w8697_,
		_w23896_,
		_w23897_,
		_w23898_
	);
	LUT4 #(
		.INIT('h7fff)
	) name21998 (
		_w23889_,
		_w23892_,
		_w23895_,
		_w23898_,
		_w23899_
	);
	LUT3 #(
		.INIT('h80)
	) name21999 (
		\m0_addr_i[2]_pad ,
		_w8699_,
		_w8700_,
		_w23900_
	);
	LUT3 #(
		.INIT('h2a)
	) name22000 (
		\m7_addr_i[2]_pad ,
		_w8699_,
		_w8700_,
		_w23901_
	);
	LUT4 #(
		.INIT('h6e7f)
	) name22001 (
		_w8694_,
		_w8697_,
		_w23900_,
		_w23901_,
		_w23902_
	);
	LUT3 #(
		.INIT('h2a)
	) name22002 (
		\m1_addr_i[2]_pad ,
		_w8699_,
		_w8700_,
		_w23903_
	);
	LUT3 #(
		.INIT('h2a)
	) name22003 (
		\m5_addr_i[2]_pad ,
		_w8699_,
		_w8700_,
		_w23904_
	);
	LUT4 #(
		.INIT('h5d7f)
	) name22004 (
		_w8694_,
		_w8697_,
		_w23903_,
		_w23904_,
		_w23905_
	);
	LUT3 #(
		.INIT('h80)
	) name22005 (
		\m2_addr_i[2]_pad ,
		_w8699_,
		_w8700_,
		_w23906_
	);
	LUT3 #(
		.INIT('h80)
	) name22006 (
		\m6_addr_i[2]_pad ,
		_w8699_,
		_w8700_,
		_w23907_
	);
	LUT4 #(
		.INIT('haebf)
	) name22007 (
		_w8694_,
		_w8697_,
		_w23906_,
		_w23907_,
		_w23908_
	);
	LUT3 #(
		.INIT('h2a)
	) name22008 (
		\m3_addr_i[2]_pad ,
		_w8699_,
		_w8700_,
		_w23909_
	);
	LUT3 #(
		.INIT('h80)
	) name22009 (
		\m4_addr_i[2]_pad ,
		_w8699_,
		_w8700_,
		_w23910_
	);
	LUT4 #(
		.INIT('h9dbf)
	) name22010 (
		_w8694_,
		_w8697_,
		_w23909_,
		_w23910_,
		_w23911_
	);
	LUT4 #(
		.INIT('h7fff)
	) name22011 (
		_w23902_,
		_w23905_,
		_w23908_,
		_w23911_,
		_w23912_
	);
	LUT3 #(
		.INIT('h2a)
	) name22012 (
		\m5_addr_i[30]_pad ,
		_w8699_,
		_w8700_,
		_w23913_
	);
	LUT3 #(
		.INIT('h80)
	) name22013 (
		\m6_addr_i[30]_pad ,
		_w8699_,
		_w8700_,
		_w23914_
	);
	LUT4 #(
		.INIT('hcedf)
	) name22014 (
		_w8694_,
		_w8697_,
		_w23913_,
		_w23914_,
		_w23915_
	);
	LUT3 #(
		.INIT('h80)
	) name22015 (
		\m0_addr_i[30]_pad ,
		_w8699_,
		_w8700_,
		_w23916_
	);
	LUT3 #(
		.INIT('h80)
	) name22016 (
		\m4_addr_i[30]_pad ,
		_w8699_,
		_w8700_,
		_w23917_
	);
	LUT4 #(
		.INIT('h5d7f)
	) name22017 (
		_w8694_,
		_w8697_,
		_w23916_,
		_w23917_,
		_w23918_
	);
	LUT3 #(
		.INIT('h2a)
	) name22018 (
		\m7_addr_i[30]_pad ,
		_w8699_,
		_w8700_,
		_w23919_
	);
	LUT3 #(
		.INIT('h2a)
	) name22019 (
		\m3_addr_i[30]_pad ,
		_w8699_,
		_w8700_,
		_w23920_
	);
	LUT4 #(
		.INIT('habef)
	) name22020 (
		_w8694_,
		_w8697_,
		_w23919_,
		_w23920_,
		_w23921_
	);
	LUT3 #(
		.INIT('h2a)
	) name22021 (
		\m1_addr_i[30]_pad ,
		_w8699_,
		_w8700_,
		_w23922_
	);
	LUT3 #(
		.INIT('h80)
	) name22022 (
		\m2_addr_i[30]_pad ,
		_w8699_,
		_w8700_,
		_w23923_
	);
	LUT4 #(
		.INIT('h3b7f)
	) name22023 (
		_w8694_,
		_w8697_,
		_w23922_,
		_w23923_,
		_w23924_
	);
	LUT4 #(
		.INIT('h7fff)
	) name22024 (
		_w23915_,
		_w23918_,
		_w23921_,
		_w23924_,
		_w23925_
	);
	LUT3 #(
		.INIT('h2a)
	) name22025 (
		\m5_addr_i[31]_pad ,
		_w8699_,
		_w8700_,
		_w23926_
	);
	LUT3 #(
		.INIT('h80)
	) name22026 (
		\m6_addr_i[31]_pad ,
		_w8699_,
		_w8700_,
		_w23927_
	);
	LUT4 #(
		.INIT('hcedf)
	) name22027 (
		_w8694_,
		_w8697_,
		_w23926_,
		_w23927_,
		_w23928_
	);
	LUT3 #(
		.INIT('h2a)
	) name22028 (
		\m3_addr_i[31]_pad ,
		_w8699_,
		_w8700_,
		_w23929_
	);
	LUT3 #(
		.INIT('h80)
	) name22029 (
		\m2_addr_i[31]_pad ,
		_w8699_,
		_w8700_,
		_w23930_
	);
	LUT3 #(
		.INIT('h57)
	) name22030 (
		_w8698_,
		_w23929_,
		_w23930_,
		_w23931_
	);
	LUT3 #(
		.INIT('h80)
	) name22031 (
		\m4_addr_i[31]_pad ,
		_w8699_,
		_w8700_,
		_w23932_
	);
	LUT3 #(
		.INIT('h2a)
	) name22032 (
		\m1_addr_i[31]_pad ,
		_w8699_,
		_w8700_,
		_w23933_
	);
	LUT4 #(
		.INIT('h57df)
	) name22033 (
		_w8694_,
		_w8697_,
		_w23932_,
		_w23933_,
		_w23934_
	);
	LUT3 #(
		.INIT('h80)
	) name22034 (
		\m0_addr_i[31]_pad ,
		_w8699_,
		_w8700_,
		_w23935_
	);
	LUT3 #(
		.INIT('h2a)
	) name22035 (
		\m7_addr_i[31]_pad ,
		_w8699_,
		_w8700_,
		_w23936_
	);
	LUT4 #(
		.INIT('h6e7f)
	) name22036 (
		_w8694_,
		_w8697_,
		_w23935_,
		_w23936_,
		_w23937_
	);
	LUT4 #(
		.INIT('h7fff)
	) name22037 (
		_w23928_,
		_w23931_,
		_w23934_,
		_w23937_,
		_w23938_
	);
	LUT3 #(
		.INIT('h2a)
	) name22038 (
		\m1_addr_i[3]_pad ,
		_w8699_,
		_w8700_,
		_w23939_
	);
	LUT3 #(
		.INIT('h80)
	) name22039 (
		\m2_addr_i[3]_pad ,
		_w8699_,
		_w8700_,
		_w23940_
	);
	LUT4 #(
		.INIT('h3b7f)
	) name22040 (
		_w8694_,
		_w8697_,
		_w23939_,
		_w23940_,
		_w23941_
	);
	LUT3 #(
		.INIT('h80)
	) name22041 (
		\m0_addr_i[3]_pad ,
		_w8699_,
		_w8700_,
		_w23942_
	);
	LUT3 #(
		.INIT('h80)
	) name22042 (
		\m4_addr_i[3]_pad ,
		_w8699_,
		_w8700_,
		_w23943_
	);
	LUT4 #(
		.INIT('h5d7f)
	) name22043 (
		_w8694_,
		_w8697_,
		_w23942_,
		_w23943_,
		_w23944_
	);
	LUT3 #(
		.INIT('h2a)
	) name22044 (
		\m7_addr_i[3]_pad ,
		_w8699_,
		_w8700_,
		_w23945_
	);
	LUT3 #(
		.INIT('h2a)
	) name22045 (
		\m3_addr_i[3]_pad ,
		_w8699_,
		_w8700_,
		_w23946_
	);
	LUT4 #(
		.INIT('habef)
	) name22046 (
		_w8694_,
		_w8697_,
		_w23945_,
		_w23946_,
		_w23947_
	);
	LUT3 #(
		.INIT('h80)
	) name22047 (
		\m6_addr_i[3]_pad ,
		_w8699_,
		_w8700_,
		_w23948_
	);
	LUT3 #(
		.INIT('h2a)
	) name22048 (
		\m5_addr_i[3]_pad ,
		_w8699_,
		_w8700_,
		_w23949_
	);
	LUT4 #(
		.INIT('hcdef)
	) name22049 (
		_w8694_,
		_w8697_,
		_w23948_,
		_w23949_,
		_w23950_
	);
	LUT4 #(
		.INIT('h7fff)
	) name22050 (
		_w23941_,
		_w23944_,
		_w23947_,
		_w23950_,
		_w23951_
	);
	LUT3 #(
		.INIT('h80)
	) name22051 (
		\m6_addr_i[4]_pad ,
		_w8699_,
		_w8700_,
		_w23952_
	);
	LUT3 #(
		.INIT('h2a)
	) name22052 (
		\m5_addr_i[4]_pad ,
		_w8699_,
		_w8700_,
		_w23953_
	);
	LUT4 #(
		.INIT('hcdef)
	) name22053 (
		_w8694_,
		_w8697_,
		_w23952_,
		_w23953_,
		_w23954_
	);
	LUT3 #(
		.INIT('h80)
	) name22054 (
		\m0_addr_i[4]_pad ,
		_w8699_,
		_w8700_,
		_w23955_
	);
	LUT3 #(
		.INIT('h80)
	) name22055 (
		\m4_addr_i[4]_pad ,
		_w8699_,
		_w8700_,
		_w23956_
	);
	LUT4 #(
		.INIT('h5d7f)
	) name22056 (
		_w8694_,
		_w8697_,
		_w23955_,
		_w23956_,
		_w23957_
	);
	LUT3 #(
		.INIT('h2a)
	) name22057 (
		\m7_addr_i[4]_pad ,
		_w8699_,
		_w8700_,
		_w23958_
	);
	LUT3 #(
		.INIT('h2a)
	) name22058 (
		\m3_addr_i[4]_pad ,
		_w8699_,
		_w8700_,
		_w23959_
	);
	LUT4 #(
		.INIT('habef)
	) name22059 (
		_w8694_,
		_w8697_,
		_w23958_,
		_w23959_,
		_w23960_
	);
	LUT3 #(
		.INIT('h2a)
	) name22060 (
		\m1_addr_i[4]_pad ,
		_w8699_,
		_w8700_,
		_w23961_
	);
	LUT3 #(
		.INIT('h80)
	) name22061 (
		\m2_addr_i[4]_pad ,
		_w8699_,
		_w8700_,
		_w23962_
	);
	LUT4 #(
		.INIT('h3b7f)
	) name22062 (
		_w8694_,
		_w8697_,
		_w23961_,
		_w23962_,
		_w23963_
	);
	LUT4 #(
		.INIT('h7fff)
	) name22063 (
		_w23954_,
		_w23957_,
		_w23960_,
		_w23963_,
		_w23964_
	);
	LUT3 #(
		.INIT('h80)
	) name22064 (
		\m6_addr_i[5]_pad ,
		_w8699_,
		_w8700_,
		_w23965_
	);
	LUT3 #(
		.INIT('h2a)
	) name22065 (
		\m5_addr_i[5]_pad ,
		_w8699_,
		_w8700_,
		_w23966_
	);
	LUT4 #(
		.INIT('hcdef)
	) name22066 (
		_w8694_,
		_w8697_,
		_w23965_,
		_w23966_,
		_w23967_
	);
	LUT3 #(
		.INIT('h2a)
	) name22067 (
		\m1_addr_i[5]_pad ,
		_w8699_,
		_w8700_,
		_w23968_
	);
	LUT3 #(
		.INIT('h80)
	) name22068 (
		\m4_addr_i[5]_pad ,
		_w8699_,
		_w8700_,
		_w23969_
	);
	LUT4 #(
		.INIT('h5d7f)
	) name22069 (
		_w8694_,
		_w8697_,
		_w23968_,
		_w23969_,
		_w23970_
	);
	LUT3 #(
		.INIT('h80)
	) name22070 (
		\m2_addr_i[5]_pad ,
		_w8699_,
		_w8700_,
		_w23971_
	);
	LUT3 #(
		.INIT('h2a)
	) name22071 (
		\m3_addr_i[5]_pad ,
		_w8699_,
		_w8700_,
		_w23972_
	);
	LUT3 #(
		.INIT('h57)
	) name22072 (
		_w8698_,
		_w23971_,
		_w23972_,
		_w23973_
	);
	LUT3 #(
		.INIT('h80)
	) name22073 (
		\m0_addr_i[5]_pad ,
		_w8699_,
		_w8700_,
		_w23974_
	);
	LUT3 #(
		.INIT('h2a)
	) name22074 (
		\m7_addr_i[5]_pad ,
		_w8699_,
		_w8700_,
		_w23975_
	);
	LUT4 #(
		.INIT('h6e7f)
	) name22075 (
		_w8694_,
		_w8697_,
		_w23974_,
		_w23975_,
		_w23976_
	);
	LUT4 #(
		.INIT('h7fff)
	) name22076 (
		_w23967_,
		_w23970_,
		_w23973_,
		_w23976_,
		_w23977_
	);
	LUT3 #(
		.INIT('h80)
	) name22077 (
		\m6_addr_i[6]_pad ,
		_w8699_,
		_w8700_,
		_w23978_
	);
	LUT3 #(
		.INIT('h2a)
	) name22078 (
		\m5_addr_i[6]_pad ,
		_w8699_,
		_w8700_,
		_w23979_
	);
	LUT4 #(
		.INIT('hcdef)
	) name22079 (
		_w8694_,
		_w8697_,
		_w23978_,
		_w23979_,
		_w23980_
	);
	LUT3 #(
		.INIT('h80)
	) name22080 (
		\m0_addr_i[6]_pad ,
		_w8699_,
		_w8700_,
		_w23981_
	);
	LUT3 #(
		.INIT('h80)
	) name22081 (
		\m4_addr_i[6]_pad ,
		_w8699_,
		_w8700_,
		_w23982_
	);
	LUT4 #(
		.INIT('h5d7f)
	) name22082 (
		_w8694_,
		_w8697_,
		_w23981_,
		_w23982_,
		_w23983_
	);
	LUT3 #(
		.INIT('h2a)
	) name22083 (
		\m7_addr_i[6]_pad ,
		_w8699_,
		_w8700_,
		_w23984_
	);
	LUT3 #(
		.INIT('h2a)
	) name22084 (
		\m3_addr_i[6]_pad ,
		_w8699_,
		_w8700_,
		_w23985_
	);
	LUT4 #(
		.INIT('habef)
	) name22085 (
		_w8694_,
		_w8697_,
		_w23984_,
		_w23985_,
		_w23986_
	);
	LUT3 #(
		.INIT('h2a)
	) name22086 (
		\m1_addr_i[6]_pad ,
		_w8699_,
		_w8700_,
		_w23987_
	);
	LUT3 #(
		.INIT('h80)
	) name22087 (
		\m2_addr_i[6]_pad ,
		_w8699_,
		_w8700_,
		_w23988_
	);
	LUT4 #(
		.INIT('h3b7f)
	) name22088 (
		_w8694_,
		_w8697_,
		_w23987_,
		_w23988_,
		_w23989_
	);
	LUT4 #(
		.INIT('h7fff)
	) name22089 (
		_w23980_,
		_w23983_,
		_w23986_,
		_w23989_,
		_w23990_
	);
	LUT3 #(
		.INIT('h2a)
	) name22090 (
		\m3_addr_i[7]_pad ,
		_w8699_,
		_w8700_,
		_w23991_
	);
	LUT3 #(
		.INIT('h80)
	) name22091 (
		\m4_addr_i[7]_pad ,
		_w8699_,
		_w8700_,
		_w23992_
	);
	LUT4 #(
		.INIT('h9dbf)
	) name22092 (
		_w8694_,
		_w8697_,
		_w23991_,
		_w23992_,
		_w23993_
	);
	LUT3 #(
		.INIT('h2a)
	) name22093 (
		\m1_addr_i[7]_pad ,
		_w8699_,
		_w8700_,
		_w23994_
	);
	LUT3 #(
		.INIT('h2a)
	) name22094 (
		\m5_addr_i[7]_pad ,
		_w8699_,
		_w8700_,
		_w23995_
	);
	LUT4 #(
		.INIT('h5d7f)
	) name22095 (
		_w8694_,
		_w8697_,
		_w23994_,
		_w23995_,
		_w23996_
	);
	LUT3 #(
		.INIT('h80)
	) name22096 (
		\m2_addr_i[7]_pad ,
		_w8699_,
		_w8700_,
		_w23997_
	);
	LUT3 #(
		.INIT('h80)
	) name22097 (
		\m6_addr_i[7]_pad ,
		_w8699_,
		_w8700_,
		_w23998_
	);
	LUT4 #(
		.INIT('haebf)
	) name22098 (
		_w8694_,
		_w8697_,
		_w23997_,
		_w23998_,
		_w23999_
	);
	LUT3 #(
		.INIT('h80)
	) name22099 (
		\m0_addr_i[7]_pad ,
		_w8699_,
		_w8700_,
		_w24000_
	);
	LUT3 #(
		.INIT('h2a)
	) name22100 (
		\m7_addr_i[7]_pad ,
		_w8699_,
		_w8700_,
		_w24001_
	);
	LUT4 #(
		.INIT('h6e7f)
	) name22101 (
		_w8694_,
		_w8697_,
		_w24000_,
		_w24001_,
		_w24002_
	);
	LUT4 #(
		.INIT('h7fff)
	) name22102 (
		_w23993_,
		_w23996_,
		_w23999_,
		_w24002_,
		_w24003_
	);
	LUT3 #(
		.INIT('h80)
	) name22103 (
		\m0_addr_i[8]_pad ,
		_w8699_,
		_w8700_,
		_w24004_
	);
	LUT3 #(
		.INIT('h2a)
	) name22104 (
		\m7_addr_i[8]_pad ,
		_w8699_,
		_w8700_,
		_w24005_
	);
	LUT4 #(
		.INIT('h6e7f)
	) name22105 (
		_w8694_,
		_w8697_,
		_w24004_,
		_w24005_,
		_w24006_
	);
	LUT3 #(
		.INIT('h2a)
	) name22106 (
		\m3_addr_i[8]_pad ,
		_w8699_,
		_w8700_,
		_w24007_
	);
	LUT3 #(
		.INIT('h2a)
	) name22107 (
		\m5_addr_i[8]_pad ,
		_w8699_,
		_w8700_,
		_w24008_
	);
	LUT4 #(
		.INIT('h9dbf)
	) name22108 (
		_w8694_,
		_w8697_,
		_w24007_,
		_w24008_,
		_w24009_
	);
	LUT3 #(
		.INIT('h80)
	) name22109 (
		\m4_addr_i[8]_pad ,
		_w8699_,
		_w8700_,
		_w24010_
	);
	LUT3 #(
		.INIT('h80)
	) name22110 (
		\m6_addr_i[8]_pad ,
		_w8699_,
		_w8700_,
		_w24011_
	);
	LUT4 #(
		.INIT('hcedf)
	) name22111 (
		_w8694_,
		_w8697_,
		_w24010_,
		_w24011_,
		_w24012_
	);
	LUT3 #(
		.INIT('h2a)
	) name22112 (
		\m1_addr_i[8]_pad ,
		_w8699_,
		_w8700_,
		_w24013_
	);
	LUT3 #(
		.INIT('h80)
	) name22113 (
		\m2_addr_i[8]_pad ,
		_w8699_,
		_w8700_,
		_w24014_
	);
	LUT4 #(
		.INIT('h3b7f)
	) name22114 (
		_w8694_,
		_w8697_,
		_w24013_,
		_w24014_,
		_w24015_
	);
	LUT4 #(
		.INIT('h7fff)
	) name22115 (
		_w24006_,
		_w24009_,
		_w24012_,
		_w24015_,
		_w24016_
	);
	LUT3 #(
		.INIT('h80)
	) name22116 (
		\m6_addr_i[9]_pad ,
		_w8699_,
		_w8700_,
		_w24017_
	);
	LUT3 #(
		.INIT('h2a)
	) name22117 (
		\m5_addr_i[9]_pad ,
		_w8699_,
		_w8700_,
		_w24018_
	);
	LUT4 #(
		.INIT('hcdef)
	) name22118 (
		_w8694_,
		_w8697_,
		_w24017_,
		_w24018_,
		_w24019_
	);
	LUT3 #(
		.INIT('h80)
	) name22119 (
		\m0_addr_i[9]_pad ,
		_w8699_,
		_w8700_,
		_w24020_
	);
	LUT3 #(
		.INIT('h80)
	) name22120 (
		\m4_addr_i[9]_pad ,
		_w8699_,
		_w8700_,
		_w24021_
	);
	LUT4 #(
		.INIT('h5d7f)
	) name22121 (
		_w8694_,
		_w8697_,
		_w24020_,
		_w24021_,
		_w24022_
	);
	LUT3 #(
		.INIT('h2a)
	) name22122 (
		\m7_addr_i[9]_pad ,
		_w8699_,
		_w8700_,
		_w24023_
	);
	LUT3 #(
		.INIT('h2a)
	) name22123 (
		\m3_addr_i[9]_pad ,
		_w8699_,
		_w8700_,
		_w24024_
	);
	LUT4 #(
		.INIT('habef)
	) name22124 (
		_w8694_,
		_w8697_,
		_w24023_,
		_w24024_,
		_w24025_
	);
	LUT3 #(
		.INIT('h2a)
	) name22125 (
		\m1_addr_i[9]_pad ,
		_w8699_,
		_w8700_,
		_w24026_
	);
	LUT3 #(
		.INIT('h80)
	) name22126 (
		\m2_addr_i[9]_pad ,
		_w8699_,
		_w8700_,
		_w24027_
	);
	LUT4 #(
		.INIT('h3b7f)
	) name22127 (
		_w8694_,
		_w8697_,
		_w24026_,
		_w24027_,
		_w24028_
	);
	LUT4 #(
		.INIT('h7fff)
	) name22128 (
		_w24019_,
		_w24022_,
		_w24025_,
		_w24028_,
		_w24029_
	);
	LUT3 #(
		.INIT('h2a)
	) name22129 (
		\m3_data_i[0]_pad ,
		_w8699_,
		_w8700_,
		_w24030_
	);
	LUT3 #(
		.INIT('h80)
	) name22130 (
		\m4_data_i[0]_pad ,
		_w8699_,
		_w8700_,
		_w24031_
	);
	LUT4 #(
		.INIT('h9dbf)
	) name22131 (
		_w8694_,
		_w8697_,
		_w24030_,
		_w24031_,
		_w24032_
	);
	LUT3 #(
		.INIT('h80)
	) name22132 (
		\m0_data_i[0]_pad ,
		_w8699_,
		_w8700_,
		_w24033_
	);
	LUT3 #(
		.INIT('h2a)
	) name22133 (
		\m5_data_i[0]_pad ,
		_w8699_,
		_w8700_,
		_w24034_
	);
	LUT4 #(
		.INIT('h5d7f)
	) name22134 (
		_w8694_,
		_w8697_,
		_w24033_,
		_w24034_,
		_w24035_
	);
	LUT3 #(
		.INIT('h2a)
	) name22135 (
		\m7_data_i[0]_pad ,
		_w8699_,
		_w8700_,
		_w24036_
	);
	LUT3 #(
		.INIT('h80)
	) name22136 (
		\m6_data_i[0]_pad ,
		_w8699_,
		_w8700_,
		_w24037_
	);
	LUT3 #(
		.INIT('h57)
	) name22137 (
		_w8712_,
		_w24036_,
		_w24037_,
		_w24038_
	);
	LUT3 #(
		.INIT('h2a)
	) name22138 (
		\m1_data_i[0]_pad ,
		_w8699_,
		_w8700_,
		_w24039_
	);
	LUT3 #(
		.INIT('h80)
	) name22139 (
		\m2_data_i[0]_pad ,
		_w8699_,
		_w8700_,
		_w24040_
	);
	LUT4 #(
		.INIT('h3b7f)
	) name22140 (
		_w8694_,
		_w8697_,
		_w24039_,
		_w24040_,
		_w24041_
	);
	LUT4 #(
		.INIT('h7fff)
	) name22141 (
		_w24032_,
		_w24035_,
		_w24038_,
		_w24041_,
		_w24042_
	);
	LUT3 #(
		.INIT('h2a)
	) name22142 (
		\m3_data_i[10]_pad ,
		_w8699_,
		_w8700_,
		_w24043_
	);
	LUT3 #(
		.INIT('h80)
	) name22143 (
		\m4_data_i[10]_pad ,
		_w8699_,
		_w8700_,
		_w24044_
	);
	LUT4 #(
		.INIT('h9dbf)
	) name22144 (
		_w8694_,
		_w8697_,
		_w24043_,
		_w24044_,
		_w24045_
	);
	LUT3 #(
		.INIT('h80)
	) name22145 (
		\m6_data_i[10]_pad ,
		_w8699_,
		_w8700_,
		_w24046_
	);
	LUT3 #(
		.INIT('h80)
	) name22146 (
		\m2_data_i[10]_pad ,
		_w8699_,
		_w8700_,
		_w24047_
	);
	LUT4 #(
		.INIT('habef)
	) name22147 (
		_w8694_,
		_w8697_,
		_w24046_,
		_w24047_,
		_w24048_
	);
	LUT3 #(
		.INIT('h2a)
	) name22148 (
		\m5_data_i[10]_pad ,
		_w8699_,
		_w8700_,
		_w24049_
	);
	LUT3 #(
		.INIT('h2a)
	) name22149 (
		\m1_data_i[10]_pad ,
		_w8699_,
		_w8700_,
		_w24050_
	);
	LUT4 #(
		.INIT('h57df)
	) name22150 (
		_w8694_,
		_w8697_,
		_w24049_,
		_w24050_,
		_w24051_
	);
	LUT3 #(
		.INIT('h80)
	) name22151 (
		\m0_data_i[10]_pad ,
		_w8699_,
		_w8700_,
		_w24052_
	);
	LUT3 #(
		.INIT('h2a)
	) name22152 (
		\m7_data_i[10]_pad ,
		_w8699_,
		_w8700_,
		_w24053_
	);
	LUT4 #(
		.INIT('h6e7f)
	) name22153 (
		_w8694_,
		_w8697_,
		_w24052_,
		_w24053_,
		_w24054_
	);
	LUT4 #(
		.INIT('h7fff)
	) name22154 (
		_w24045_,
		_w24048_,
		_w24051_,
		_w24054_,
		_w24055_
	);
	LUT3 #(
		.INIT('h2a)
	) name22155 (
		\m3_data_i[11]_pad ,
		_w8699_,
		_w8700_,
		_w24056_
	);
	LUT3 #(
		.INIT('h80)
	) name22156 (
		\m4_data_i[11]_pad ,
		_w8699_,
		_w8700_,
		_w24057_
	);
	LUT4 #(
		.INIT('h9dbf)
	) name22157 (
		_w8694_,
		_w8697_,
		_w24056_,
		_w24057_,
		_w24058_
	);
	LUT3 #(
		.INIT('h80)
	) name22158 (
		\m6_data_i[11]_pad ,
		_w8699_,
		_w8700_,
		_w24059_
	);
	LUT3 #(
		.INIT('h80)
	) name22159 (
		\m2_data_i[11]_pad ,
		_w8699_,
		_w8700_,
		_w24060_
	);
	LUT4 #(
		.INIT('habef)
	) name22160 (
		_w8694_,
		_w8697_,
		_w24059_,
		_w24060_,
		_w24061_
	);
	LUT3 #(
		.INIT('h2a)
	) name22161 (
		\m5_data_i[11]_pad ,
		_w8699_,
		_w8700_,
		_w24062_
	);
	LUT3 #(
		.INIT('h2a)
	) name22162 (
		\m1_data_i[11]_pad ,
		_w8699_,
		_w8700_,
		_w24063_
	);
	LUT4 #(
		.INIT('h57df)
	) name22163 (
		_w8694_,
		_w8697_,
		_w24062_,
		_w24063_,
		_w24064_
	);
	LUT3 #(
		.INIT('h80)
	) name22164 (
		\m0_data_i[11]_pad ,
		_w8699_,
		_w8700_,
		_w24065_
	);
	LUT3 #(
		.INIT('h2a)
	) name22165 (
		\m7_data_i[11]_pad ,
		_w8699_,
		_w8700_,
		_w24066_
	);
	LUT4 #(
		.INIT('h6e7f)
	) name22166 (
		_w8694_,
		_w8697_,
		_w24065_,
		_w24066_,
		_w24067_
	);
	LUT4 #(
		.INIT('h7fff)
	) name22167 (
		_w24058_,
		_w24061_,
		_w24064_,
		_w24067_,
		_w24068_
	);
	LUT3 #(
		.INIT('h2a)
	) name22168 (
		\m3_data_i[12]_pad ,
		_w8699_,
		_w8700_,
		_w24069_
	);
	LUT3 #(
		.INIT('h80)
	) name22169 (
		\m4_data_i[12]_pad ,
		_w8699_,
		_w8700_,
		_w24070_
	);
	LUT4 #(
		.INIT('h9dbf)
	) name22170 (
		_w8694_,
		_w8697_,
		_w24069_,
		_w24070_,
		_w24071_
	);
	LUT3 #(
		.INIT('h80)
	) name22171 (
		\m6_data_i[12]_pad ,
		_w8699_,
		_w8700_,
		_w24072_
	);
	LUT3 #(
		.INIT('h80)
	) name22172 (
		\m2_data_i[12]_pad ,
		_w8699_,
		_w8700_,
		_w24073_
	);
	LUT4 #(
		.INIT('habef)
	) name22173 (
		_w8694_,
		_w8697_,
		_w24072_,
		_w24073_,
		_w24074_
	);
	LUT3 #(
		.INIT('h2a)
	) name22174 (
		\m5_data_i[12]_pad ,
		_w8699_,
		_w8700_,
		_w24075_
	);
	LUT3 #(
		.INIT('h2a)
	) name22175 (
		\m1_data_i[12]_pad ,
		_w8699_,
		_w8700_,
		_w24076_
	);
	LUT4 #(
		.INIT('h57df)
	) name22176 (
		_w8694_,
		_w8697_,
		_w24075_,
		_w24076_,
		_w24077_
	);
	LUT3 #(
		.INIT('h80)
	) name22177 (
		\m0_data_i[12]_pad ,
		_w8699_,
		_w8700_,
		_w24078_
	);
	LUT3 #(
		.INIT('h2a)
	) name22178 (
		\m7_data_i[12]_pad ,
		_w8699_,
		_w8700_,
		_w24079_
	);
	LUT4 #(
		.INIT('h6e7f)
	) name22179 (
		_w8694_,
		_w8697_,
		_w24078_,
		_w24079_,
		_w24080_
	);
	LUT4 #(
		.INIT('h7fff)
	) name22180 (
		_w24071_,
		_w24074_,
		_w24077_,
		_w24080_,
		_w24081_
	);
	LUT3 #(
		.INIT('h2a)
	) name22181 (
		\m3_data_i[13]_pad ,
		_w8699_,
		_w8700_,
		_w24082_
	);
	LUT3 #(
		.INIT('h80)
	) name22182 (
		\m4_data_i[13]_pad ,
		_w8699_,
		_w8700_,
		_w24083_
	);
	LUT4 #(
		.INIT('h9dbf)
	) name22183 (
		_w8694_,
		_w8697_,
		_w24082_,
		_w24083_,
		_w24084_
	);
	LUT3 #(
		.INIT('h80)
	) name22184 (
		\m6_data_i[13]_pad ,
		_w8699_,
		_w8700_,
		_w24085_
	);
	LUT3 #(
		.INIT('h80)
	) name22185 (
		\m2_data_i[13]_pad ,
		_w8699_,
		_w8700_,
		_w24086_
	);
	LUT4 #(
		.INIT('habef)
	) name22186 (
		_w8694_,
		_w8697_,
		_w24085_,
		_w24086_,
		_w24087_
	);
	LUT3 #(
		.INIT('h2a)
	) name22187 (
		\m5_data_i[13]_pad ,
		_w8699_,
		_w8700_,
		_w24088_
	);
	LUT3 #(
		.INIT('h2a)
	) name22188 (
		\m1_data_i[13]_pad ,
		_w8699_,
		_w8700_,
		_w24089_
	);
	LUT4 #(
		.INIT('h57df)
	) name22189 (
		_w8694_,
		_w8697_,
		_w24088_,
		_w24089_,
		_w24090_
	);
	LUT3 #(
		.INIT('h80)
	) name22190 (
		\m0_data_i[13]_pad ,
		_w8699_,
		_w8700_,
		_w24091_
	);
	LUT3 #(
		.INIT('h2a)
	) name22191 (
		\m7_data_i[13]_pad ,
		_w8699_,
		_w8700_,
		_w24092_
	);
	LUT4 #(
		.INIT('h6e7f)
	) name22192 (
		_w8694_,
		_w8697_,
		_w24091_,
		_w24092_,
		_w24093_
	);
	LUT4 #(
		.INIT('h7fff)
	) name22193 (
		_w24084_,
		_w24087_,
		_w24090_,
		_w24093_,
		_w24094_
	);
	LUT3 #(
		.INIT('h2a)
	) name22194 (
		\m3_data_i[14]_pad ,
		_w8699_,
		_w8700_,
		_w24095_
	);
	LUT3 #(
		.INIT('h80)
	) name22195 (
		\m4_data_i[14]_pad ,
		_w8699_,
		_w8700_,
		_w24096_
	);
	LUT4 #(
		.INIT('h9dbf)
	) name22196 (
		_w8694_,
		_w8697_,
		_w24095_,
		_w24096_,
		_w24097_
	);
	LUT3 #(
		.INIT('h80)
	) name22197 (
		\m6_data_i[14]_pad ,
		_w8699_,
		_w8700_,
		_w24098_
	);
	LUT3 #(
		.INIT('h80)
	) name22198 (
		\m2_data_i[14]_pad ,
		_w8699_,
		_w8700_,
		_w24099_
	);
	LUT4 #(
		.INIT('habef)
	) name22199 (
		_w8694_,
		_w8697_,
		_w24098_,
		_w24099_,
		_w24100_
	);
	LUT3 #(
		.INIT('h2a)
	) name22200 (
		\m5_data_i[14]_pad ,
		_w8699_,
		_w8700_,
		_w24101_
	);
	LUT3 #(
		.INIT('h2a)
	) name22201 (
		\m1_data_i[14]_pad ,
		_w8699_,
		_w8700_,
		_w24102_
	);
	LUT4 #(
		.INIT('h57df)
	) name22202 (
		_w8694_,
		_w8697_,
		_w24101_,
		_w24102_,
		_w24103_
	);
	LUT3 #(
		.INIT('h80)
	) name22203 (
		\m0_data_i[14]_pad ,
		_w8699_,
		_w8700_,
		_w24104_
	);
	LUT3 #(
		.INIT('h2a)
	) name22204 (
		\m7_data_i[14]_pad ,
		_w8699_,
		_w8700_,
		_w24105_
	);
	LUT4 #(
		.INIT('h6e7f)
	) name22205 (
		_w8694_,
		_w8697_,
		_w24104_,
		_w24105_,
		_w24106_
	);
	LUT4 #(
		.INIT('h7fff)
	) name22206 (
		_w24097_,
		_w24100_,
		_w24103_,
		_w24106_,
		_w24107_
	);
	LUT3 #(
		.INIT('h2a)
	) name22207 (
		\m3_data_i[15]_pad ,
		_w8699_,
		_w8700_,
		_w24108_
	);
	LUT3 #(
		.INIT('h80)
	) name22208 (
		\m4_data_i[15]_pad ,
		_w8699_,
		_w8700_,
		_w24109_
	);
	LUT4 #(
		.INIT('h9dbf)
	) name22209 (
		_w8694_,
		_w8697_,
		_w24108_,
		_w24109_,
		_w24110_
	);
	LUT3 #(
		.INIT('h80)
	) name22210 (
		\m6_data_i[15]_pad ,
		_w8699_,
		_w8700_,
		_w24111_
	);
	LUT3 #(
		.INIT('h80)
	) name22211 (
		\m2_data_i[15]_pad ,
		_w8699_,
		_w8700_,
		_w24112_
	);
	LUT4 #(
		.INIT('habef)
	) name22212 (
		_w8694_,
		_w8697_,
		_w24111_,
		_w24112_,
		_w24113_
	);
	LUT3 #(
		.INIT('h2a)
	) name22213 (
		\m5_data_i[15]_pad ,
		_w8699_,
		_w8700_,
		_w24114_
	);
	LUT3 #(
		.INIT('h2a)
	) name22214 (
		\m1_data_i[15]_pad ,
		_w8699_,
		_w8700_,
		_w24115_
	);
	LUT4 #(
		.INIT('h57df)
	) name22215 (
		_w8694_,
		_w8697_,
		_w24114_,
		_w24115_,
		_w24116_
	);
	LUT3 #(
		.INIT('h80)
	) name22216 (
		\m0_data_i[15]_pad ,
		_w8699_,
		_w8700_,
		_w24117_
	);
	LUT3 #(
		.INIT('h2a)
	) name22217 (
		\m7_data_i[15]_pad ,
		_w8699_,
		_w8700_,
		_w24118_
	);
	LUT4 #(
		.INIT('h6e7f)
	) name22218 (
		_w8694_,
		_w8697_,
		_w24117_,
		_w24118_,
		_w24119_
	);
	LUT4 #(
		.INIT('h7fff)
	) name22219 (
		_w24110_,
		_w24113_,
		_w24116_,
		_w24119_,
		_w24120_
	);
	LUT3 #(
		.INIT('h2a)
	) name22220 (
		\m3_data_i[16]_pad ,
		_w8699_,
		_w8700_,
		_w24121_
	);
	LUT3 #(
		.INIT('h80)
	) name22221 (
		\m4_data_i[16]_pad ,
		_w8699_,
		_w8700_,
		_w24122_
	);
	LUT4 #(
		.INIT('h9dbf)
	) name22222 (
		_w8694_,
		_w8697_,
		_w24121_,
		_w24122_,
		_w24123_
	);
	LUT3 #(
		.INIT('h80)
	) name22223 (
		\m6_data_i[16]_pad ,
		_w8699_,
		_w8700_,
		_w24124_
	);
	LUT3 #(
		.INIT('h80)
	) name22224 (
		\m2_data_i[16]_pad ,
		_w8699_,
		_w8700_,
		_w24125_
	);
	LUT4 #(
		.INIT('habef)
	) name22225 (
		_w8694_,
		_w8697_,
		_w24124_,
		_w24125_,
		_w24126_
	);
	LUT3 #(
		.INIT('h2a)
	) name22226 (
		\m5_data_i[16]_pad ,
		_w8699_,
		_w8700_,
		_w24127_
	);
	LUT3 #(
		.INIT('h2a)
	) name22227 (
		\m1_data_i[16]_pad ,
		_w8699_,
		_w8700_,
		_w24128_
	);
	LUT4 #(
		.INIT('h57df)
	) name22228 (
		_w8694_,
		_w8697_,
		_w24127_,
		_w24128_,
		_w24129_
	);
	LUT3 #(
		.INIT('h80)
	) name22229 (
		\m0_data_i[16]_pad ,
		_w8699_,
		_w8700_,
		_w24130_
	);
	LUT3 #(
		.INIT('h2a)
	) name22230 (
		\m7_data_i[16]_pad ,
		_w8699_,
		_w8700_,
		_w24131_
	);
	LUT4 #(
		.INIT('h6e7f)
	) name22231 (
		_w8694_,
		_w8697_,
		_w24130_,
		_w24131_,
		_w24132_
	);
	LUT4 #(
		.INIT('h7fff)
	) name22232 (
		_w24123_,
		_w24126_,
		_w24129_,
		_w24132_,
		_w24133_
	);
	LUT3 #(
		.INIT('h2a)
	) name22233 (
		\m3_data_i[17]_pad ,
		_w8699_,
		_w8700_,
		_w24134_
	);
	LUT3 #(
		.INIT('h80)
	) name22234 (
		\m4_data_i[17]_pad ,
		_w8699_,
		_w8700_,
		_w24135_
	);
	LUT4 #(
		.INIT('h9dbf)
	) name22235 (
		_w8694_,
		_w8697_,
		_w24134_,
		_w24135_,
		_w24136_
	);
	LUT3 #(
		.INIT('h80)
	) name22236 (
		\m6_data_i[17]_pad ,
		_w8699_,
		_w8700_,
		_w24137_
	);
	LUT3 #(
		.INIT('h80)
	) name22237 (
		\m2_data_i[17]_pad ,
		_w8699_,
		_w8700_,
		_w24138_
	);
	LUT4 #(
		.INIT('habef)
	) name22238 (
		_w8694_,
		_w8697_,
		_w24137_,
		_w24138_,
		_w24139_
	);
	LUT3 #(
		.INIT('h2a)
	) name22239 (
		\m5_data_i[17]_pad ,
		_w8699_,
		_w8700_,
		_w24140_
	);
	LUT3 #(
		.INIT('h2a)
	) name22240 (
		\m1_data_i[17]_pad ,
		_w8699_,
		_w8700_,
		_w24141_
	);
	LUT4 #(
		.INIT('h57df)
	) name22241 (
		_w8694_,
		_w8697_,
		_w24140_,
		_w24141_,
		_w24142_
	);
	LUT3 #(
		.INIT('h80)
	) name22242 (
		\m0_data_i[17]_pad ,
		_w8699_,
		_w8700_,
		_w24143_
	);
	LUT3 #(
		.INIT('h2a)
	) name22243 (
		\m7_data_i[17]_pad ,
		_w8699_,
		_w8700_,
		_w24144_
	);
	LUT4 #(
		.INIT('h6e7f)
	) name22244 (
		_w8694_,
		_w8697_,
		_w24143_,
		_w24144_,
		_w24145_
	);
	LUT4 #(
		.INIT('h7fff)
	) name22245 (
		_w24136_,
		_w24139_,
		_w24142_,
		_w24145_,
		_w24146_
	);
	LUT3 #(
		.INIT('h2a)
	) name22246 (
		\m3_data_i[18]_pad ,
		_w8699_,
		_w8700_,
		_w24147_
	);
	LUT3 #(
		.INIT('h80)
	) name22247 (
		\m4_data_i[18]_pad ,
		_w8699_,
		_w8700_,
		_w24148_
	);
	LUT4 #(
		.INIT('h9dbf)
	) name22248 (
		_w8694_,
		_w8697_,
		_w24147_,
		_w24148_,
		_w24149_
	);
	LUT3 #(
		.INIT('h80)
	) name22249 (
		\m6_data_i[18]_pad ,
		_w8699_,
		_w8700_,
		_w24150_
	);
	LUT3 #(
		.INIT('h80)
	) name22250 (
		\m2_data_i[18]_pad ,
		_w8699_,
		_w8700_,
		_w24151_
	);
	LUT4 #(
		.INIT('habef)
	) name22251 (
		_w8694_,
		_w8697_,
		_w24150_,
		_w24151_,
		_w24152_
	);
	LUT3 #(
		.INIT('h2a)
	) name22252 (
		\m5_data_i[18]_pad ,
		_w8699_,
		_w8700_,
		_w24153_
	);
	LUT3 #(
		.INIT('h2a)
	) name22253 (
		\m1_data_i[18]_pad ,
		_w8699_,
		_w8700_,
		_w24154_
	);
	LUT4 #(
		.INIT('h57df)
	) name22254 (
		_w8694_,
		_w8697_,
		_w24153_,
		_w24154_,
		_w24155_
	);
	LUT3 #(
		.INIT('h80)
	) name22255 (
		\m0_data_i[18]_pad ,
		_w8699_,
		_w8700_,
		_w24156_
	);
	LUT3 #(
		.INIT('h2a)
	) name22256 (
		\m7_data_i[18]_pad ,
		_w8699_,
		_w8700_,
		_w24157_
	);
	LUT4 #(
		.INIT('h6e7f)
	) name22257 (
		_w8694_,
		_w8697_,
		_w24156_,
		_w24157_,
		_w24158_
	);
	LUT4 #(
		.INIT('h7fff)
	) name22258 (
		_w24149_,
		_w24152_,
		_w24155_,
		_w24158_,
		_w24159_
	);
	LUT3 #(
		.INIT('h2a)
	) name22259 (
		\m3_data_i[19]_pad ,
		_w8699_,
		_w8700_,
		_w24160_
	);
	LUT3 #(
		.INIT('h80)
	) name22260 (
		\m4_data_i[19]_pad ,
		_w8699_,
		_w8700_,
		_w24161_
	);
	LUT4 #(
		.INIT('h9dbf)
	) name22261 (
		_w8694_,
		_w8697_,
		_w24160_,
		_w24161_,
		_w24162_
	);
	LUT3 #(
		.INIT('h80)
	) name22262 (
		\m6_data_i[19]_pad ,
		_w8699_,
		_w8700_,
		_w24163_
	);
	LUT3 #(
		.INIT('h80)
	) name22263 (
		\m2_data_i[19]_pad ,
		_w8699_,
		_w8700_,
		_w24164_
	);
	LUT4 #(
		.INIT('habef)
	) name22264 (
		_w8694_,
		_w8697_,
		_w24163_,
		_w24164_,
		_w24165_
	);
	LUT3 #(
		.INIT('h2a)
	) name22265 (
		\m5_data_i[19]_pad ,
		_w8699_,
		_w8700_,
		_w24166_
	);
	LUT3 #(
		.INIT('h2a)
	) name22266 (
		\m1_data_i[19]_pad ,
		_w8699_,
		_w8700_,
		_w24167_
	);
	LUT4 #(
		.INIT('h57df)
	) name22267 (
		_w8694_,
		_w8697_,
		_w24166_,
		_w24167_,
		_w24168_
	);
	LUT3 #(
		.INIT('h80)
	) name22268 (
		\m0_data_i[19]_pad ,
		_w8699_,
		_w8700_,
		_w24169_
	);
	LUT3 #(
		.INIT('h2a)
	) name22269 (
		\m7_data_i[19]_pad ,
		_w8699_,
		_w8700_,
		_w24170_
	);
	LUT4 #(
		.INIT('h6e7f)
	) name22270 (
		_w8694_,
		_w8697_,
		_w24169_,
		_w24170_,
		_w24171_
	);
	LUT4 #(
		.INIT('h7fff)
	) name22271 (
		_w24162_,
		_w24165_,
		_w24168_,
		_w24171_,
		_w24172_
	);
	LUT3 #(
		.INIT('h2a)
	) name22272 (
		\m1_data_i[1]_pad ,
		_w8699_,
		_w8700_,
		_w24173_
	);
	LUT3 #(
		.INIT('h80)
	) name22273 (
		\m2_data_i[1]_pad ,
		_w8699_,
		_w8700_,
		_w24174_
	);
	LUT4 #(
		.INIT('h3b7f)
	) name22274 (
		_w8694_,
		_w8697_,
		_w24173_,
		_w24174_,
		_w24175_
	);
	LUT3 #(
		.INIT('h80)
	) name22275 (
		\m6_data_i[1]_pad ,
		_w8699_,
		_w8700_,
		_w24176_
	);
	LUT3 #(
		.INIT('h2a)
	) name22276 (
		\m7_data_i[1]_pad ,
		_w8699_,
		_w8700_,
		_w24177_
	);
	LUT3 #(
		.INIT('h57)
	) name22277 (
		_w8712_,
		_w24176_,
		_w24177_,
		_w24178_
	);
	LUT3 #(
		.INIT('h2a)
	) name22278 (
		\m5_data_i[1]_pad ,
		_w8699_,
		_w8700_,
		_w24179_
	);
	LUT3 #(
		.INIT('h80)
	) name22279 (
		\m0_data_i[1]_pad ,
		_w8699_,
		_w8700_,
		_w24180_
	);
	LUT4 #(
		.INIT('h57df)
	) name22280 (
		_w8694_,
		_w8697_,
		_w24179_,
		_w24180_,
		_w24181_
	);
	LUT3 #(
		.INIT('h2a)
	) name22281 (
		\m3_data_i[1]_pad ,
		_w8699_,
		_w8700_,
		_w24182_
	);
	LUT3 #(
		.INIT('h80)
	) name22282 (
		\m4_data_i[1]_pad ,
		_w8699_,
		_w8700_,
		_w24183_
	);
	LUT4 #(
		.INIT('h9dbf)
	) name22283 (
		_w8694_,
		_w8697_,
		_w24182_,
		_w24183_,
		_w24184_
	);
	LUT4 #(
		.INIT('h7fff)
	) name22284 (
		_w24175_,
		_w24178_,
		_w24181_,
		_w24184_,
		_w24185_
	);
	LUT3 #(
		.INIT('h2a)
	) name22285 (
		\m3_data_i[20]_pad ,
		_w8699_,
		_w8700_,
		_w24186_
	);
	LUT3 #(
		.INIT('h80)
	) name22286 (
		\m4_data_i[20]_pad ,
		_w8699_,
		_w8700_,
		_w24187_
	);
	LUT4 #(
		.INIT('h9dbf)
	) name22287 (
		_w8694_,
		_w8697_,
		_w24186_,
		_w24187_,
		_w24188_
	);
	LUT3 #(
		.INIT('h80)
	) name22288 (
		\m6_data_i[20]_pad ,
		_w8699_,
		_w8700_,
		_w24189_
	);
	LUT3 #(
		.INIT('h80)
	) name22289 (
		\m2_data_i[20]_pad ,
		_w8699_,
		_w8700_,
		_w24190_
	);
	LUT4 #(
		.INIT('habef)
	) name22290 (
		_w8694_,
		_w8697_,
		_w24189_,
		_w24190_,
		_w24191_
	);
	LUT3 #(
		.INIT('h2a)
	) name22291 (
		\m5_data_i[20]_pad ,
		_w8699_,
		_w8700_,
		_w24192_
	);
	LUT3 #(
		.INIT('h2a)
	) name22292 (
		\m1_data_i[20]_pad ,
		_w8699_,
		_w8700_,
		_w24193_
	);
	LUT4 #(
		.INIT('h57df)
	) name22293 (
		_w8694_,
		_w8697_,
		_w24192_,
		_w24193_,
		_w24194_
	);
	LUT3 #(
		.INIT('h80)
	) name22294 (
		\m0_data_i[20]_pad ,
		_w8699_,
		_w8700_,
		_w24195_
	);
	LUT3 #(
		.INIT('h2a)
	) name22295 (
		\m7_data_i[20]_pad ,
		_w8699_,
		_w8700_,
		_w24196_
	);
	LUT4 #(
		.INIT('h6e7f)
	) name22296 (
		_w8694_,
		_w8697_,
		_w24195_,
		_w24196_,
		_w24197_
	);
	LUT4 #(
		.INIT('h7fff)
	) name22297 (
		_w24188_,
		_w24191_,
		_w24194_,
		_w24197_,
		_w24198_
	);
	LUT3 #(
		.INIT('h2a)
	) name22298 (
		\m3_data_i[21]_pad ,
		_w8699_,
		_w8700_,
		_w24199_
	);
	LUT3 #(
		.INIT('h80)
	) name22299 (
		\m4_data_i[21]_pad ,
		_w8699_,
		_w8700_,
		_w24200_
	);
	LUT4 #(
		.INIT('h9dbf)
	) name22300 (
		_w8694_,
		_w8697_,
		_w24199_,
		_w24200_,
		_w24201_
	);
	LUT3 #(
		.INIT('h80)
	) name22301 (
		\m6_data_i[21]_pad ,
		_w8699_,
		_w8700_,
		_w24202_
	);
	LUT3 #(
		.INIT('h80)
	) name22302 (
		\m2_data_i[21]_pad ,
		_w8699_,
		_w8700_,
		_w24203_
	);
	LUT4 #(
		.INIT('habef)
	) name22303 (
		_w8694_,
		_w8697_,
		_w24202_,
		_w24203_,
		_w24204_
	);
	LUT3 #(
		.INIT('h2a)
	) name22304 (
		\m5_data_i[21]_pad ,
		_w8699_,
		_w8700_,
		_w24205_
	);
	LUT3 #(
		.INIT('h2a)
	) name22305 (
		\m1_data_i[21]_pad ,
		_w8699_,
		_w8700_,
		_w24206_
	);
	LUT4 #(
		.INIT('h57df)
	) name22306 (
		_w8694_,
		_w8697_,
		_w24205_,
		_w24206_,
		_w24207_
	);
	LUT3 #(
		.INIT('h80)
	) name22307 (
		\m0_data_i[21]_pad ,
		_w8699_,
		_w8700_,
		_w24208_
	);
	LUT3 #(
		.INIT('h2a)
	) name22308 (
		\m7_data_i[21]_pad ,
		_w8699_,
		_w8700_,
		_w24209_
	);
	LUT4 #(
		.INIT('h6e7f)
	) name22309 (
		_w8694_,
		_w8697_,
		_w24208_,
		_w24209_,
		_w24210_
	);
	LUT4 #(
		.INIT('h7fff)
	) name22310 (
		_w24201_,
		_w24204_,
		_w24207_,
		_w24210_,
		_w24211_
	);
	LUT3 #(
		.INIT('h2a)
	) name22311 (
		\m3_data_i[22]_pad ,
		_w8699_,
		_w8700_,
		_w24212_
	);
	LUT3 #(
		.INIT('h80)
	) name22312 (
		\m4_data_i[22]_pad ,
		_w8699_,
		_w8700_,
		_w24213_
	);
	LUT4 #(
		.INIT('h9dbf)
	) name22313 (
		_w8694_,
		_w8697_,
		_w24212_,
		_w24213_,
		_w24214_
	);
	LUT3 #(
		.INIT('h80)
	) name22314 (
		\m6_data_i[22]_pad ,
		_w8699_,
		_w8700_,
		_w24215_
	);
	LUT3 #(
		.INIT('h80)
	) name22315 (
		\m2_data_i[22]_pad ,
		_w8699_,
		_w8700_,
		_w24216_
	);
	LUT4 #(
		.INIT('habef)
	) name22316 (
		_w8694_,
		_w8697_,
		_w24215_,
		_w24216_,
		_w24217_
	);
	LUT3 #(
		.INIT('h2a)
	) name22317 (
		\m5_data_i[22]_pad ,
		_w8699_,
		_w8700_,
		_w24218_
	);
	LUT3 #(
		.INIT('h2a)
	) name22318 (
		\m1_data_i[22]_pad ,
		_w8699_,
		_w8700_,
		_w24219_
	);
	LUT4 #(
		.INIT('h57df)
	) name22319 (
		_w8694_,
		_w8697_,
		_w24218_,
		_w24219_,
		_w24220_
	);
	LUT3 #(
		.INIT('h80)
	) name22320 (
		\m0_data_i[22]_pad ,
		_w8699_,
		_w8700_,
		_w24221_
	);
	LUT3 #(
		.INIT('h2a)
	) name22321 (
		\m7_data_i[22]_pad ,
		_w8699_,
		_w8700_,
		_w24222_
	);
	LUT4 #(
		.INIT('h6e7f)
	) name22322 (
		_w8694_,
		_w8697_,
		_w24221_,
		_w24222_,
		_w24223_
	);
	LUT4 #(
		.INIT('h7fff)
	) name22323 (
		_w24214_,
		_w24217_,
		_w24220_,
		_w24223_,
		_w24224_
	);
	LUT3 #(
		.INIT('h80)
	) name22324 (
		\m6_data_i[23]_pad ,
		_w8699_,
		_w8700_,
		_w24225_
	);
	LUT3 #(
		.INIT('h2a)
	) name22325 (
		\m5_data_i[23]_pad ,
		_w8699_,
		_w8700_,
		_w24226_
	);
	LUT4 #(
		.INIT('hcdef)
	) name22326 (
		_w8694_,
		_w8697_,
		_w24225_,
		_w24226_,
		_w24227_
	);
	LUT3 #(
		.INIT('h80)
	) name22327 (
		\m0_data_i[23]_pad ,
		_w8699_,
		_w8700_,
		_w24228_
	);
	LUT3 #(
		.INIT('h80)
	) name22328 (
		\m4_data_i[23]_pad ,
		_w8699_,
		_w8700_,
		_w24229_
	);
	LUT4 #(
		.INIT('h5d7f)
	) name22329 (
		_w8694_,
		_w8697_,
		_w24228_,
		_w24229_,
		_w24230_
	);
	LUT3 #(
		.INIT('h2a)
	) name22330 (
		\m7_data_i[23]_pad ,
		_w8699_,
		_w8700_,
		_w24231_
	);
	LUT3 #(
		.INIT('h2a)
	) name22331 (
		\m3_data_i[23]_pad ,
		_w8699_,
		_w8700_,
		_w24232_
	);
	LUT4 #(
		.INIT('habef)
	) name22332 (
		_w8694_,
		_w8697_,
		_w24231_,
		_w24232_,
		_w24233_
	);
	LUT3 #(
		.INIT('h2a)
	) name22333 (
		\m1_data_i[23]_pad ,
		_w8699_,
		_w8700_,
		_w24234_
	);
	LUT3 #(
		.INIT('h80)
	) name22334 (
		\m2_data_i[23]_pad ,
		_w8699_,
		_w8700_,
		_w24235_
	);
	LUT4 #(
		.INIT('h3b7f)
	) name22335 (
		_w8694_,
		_w8697_,
		_w24234_,
		_w24235_,
		_w24236_
	);
	LUT4 #(
		.INIT('h7fff)
	) name22336 (
		_w24227_,
		_w24230_,
		_w24233_,
		_w24236_,
		_w24237_
	);
	LUT3 #(
		.INIT('h2a)
	) name22337 (
		\m3_data_i[24]_pad ,
		_w8699_,
		_w8700_,
		_w24238_
	);
	LUT3 #(
		.INIT('h80)
	) name22338 (
		\m4_data_i[24]_pad ,
		_w8699_,
		_w8700_,
		_w24239_
	);
	LUT4 #(
		.INIT('h9dbf)
	) name22339 (
		_w8694_,
		_w8697_,
		_w24238_,
		_w24239_,
		_w24240_
	);
	LUT3 #(
		.INIT('h80)
	) name22340 (
		\m6_data_i[24]_pad ,
		_w8699_,
		_w8700_,
		_w24241_
	);
	LUT3 #(
		.INIT('h80)
	) name22341 (
		\m2_data_i[24]_pad ,
		_w8699_,
		_w8700_,
		_w24242_
	);
	LUT4 #(
		.INIT('habef)
	) name22342 (
		_w8694_,
		_w8697_,
		_w24241_,
		_w24242_,
		_w24243_
	);
	LUT3 #(
		.INIT('h2a)
	) name22343 (
		\m5_data_i[24]_pad ,
		_w8699_,
		_w8700_,
		_w24244_
	);
	LUT3 #(
		.INIT('h2a)
	) name22344 (
		\m1_data_i[24]_pad ,
		_w8699_,
		_w8700_,
		_w24245_
	);
	LUT4 #(
		.INIT('h57df)
	) name22345 (
		_w8694_,
		_w8697_,
		_w24244_,
		_w24245_,
		_w24246_
	);
	LUT3 #(
		.INIT('h80)
	) name22346 (
		\m0_data_i[24]_pad ,
		_w8699_,
		_w8700_,
		_w24247_
	);
	LUT3 #(
		.INIT('h2a)
	) name22347 (
		\m7_data_i[24]_pad ,
		_w8699_,
		_w8700_,
		_w24248_
	);
	LUT4 #(
		.INIT('h6e7f)
	) name22348 (
		_w8694_,
		_w8697_,
		_w24247_,
		_w24248_,
		_w24249_
	);
	LUT4 #(
		.INIT('h7fff)
	) name22349 (
		_w24240_,
		_w24243_,
		_w24246_,
		_w24249_,
		_w24250_
	);
	LUT3 #(
		.INIT('h2a)
	) name22350 (
		\m3_data_i[25]_pad ,
		_w8699_,
		_w8700_,
		_w24251_
	);
	LUT3 #(
		.INIT('h80)
	) name22351 (
		\m4_data_i[25]_pad ,
		_w8699_,
		_w8700_,
		_w24252_
	);
	LUT4 #(
		.INIT('h9dbf)
	) name22352 (
		_w8694_,
		_w8697_,
		_w24251_,
		_w24252_,
		_w24253_
	);
	LUT3 #(
		.INIT('h80)
	) name22353 (
		\m6_data_i[25]_pad ,
		_w8699_,
		_w8700_,
		_w24254_
	);
	LUT3 #(
		.INIT('h80)
	) name22354 (
		\m2_data_i[25]_pad ,
		_w8699_,
		_w8700_,
		_w24255_
	);
	LUT4 #(
		.INIT('habef)
	) name22355 (
		_w8694_,
		_w8697_,
		_w24254_,
		_w24255_,
		_w24256_
	);
	LUT3 #(
		.INIT('h2a)
	) name22356 (
		\m5_data_i[25]_pad ,
		_w8699_,
		_w8700_,
		_w24257_
	);
	LUT3 #(
		.INIT('h2a)
	) name22357 (
		\m1_data_i[25]_pad ,
		_w8699_,
		_w8700_,
		_w24258_
	);
	LUT4 #(
		.INIT('h57df)
	) name22358 (
		_w8694_,
		_w8697_,
		_w24257_,
		_w24258_,
		_w24259_
	);
	LUT3 #(
		.INIT('h80)
	) name22359 (
		\m0_data_i[25]_pad ,
		_w8699_,
		_w8700_,
		_w24260_
	);
	LUT3 #(
		.INIT('h2a)
	) name22360 (
		\m7_data_i[25]_pad ,
		_w8699_,
		_w8700_,
		_w24261_
	);
	LUT4 #(
		.INIT('h6e7f)
	) name22361 (
		_w8694_,
		_w8697_,
		_w24260_,
		_w24261_,
		_w24262_
	);
	LUT4 #(
		.INIT('h7fff)
	) name22362 (
		_w24253_,
		_w24256_,
		_w24259_,
		_w24262_,
		_w24263_
	);
	LUT3 #(
		.INIT('h2a)
	) name22363 (
		\m3_data_i[26]_pad ,
		_w8699_,
		_w8700_,
		_w24264_
	);
	LUT3 #(
		.INIT('h80)
	) name22364 (
		\m4_data_i[26]_pad ,
		_w8699_,
		_w8700_,
		_w24265_
	);
	LUT4 #(
		.INIT('h9dbf)
	) name22365 (
		_w8694_,
		_w8697_,
		_w24264_,
		_w24265_,
		_w24266_
	);
	LUT3 #(
		.INIT('h80)
	) name22366 (
		\m6_data_i[26]_pad ,
		_w8699_,
		_w8700_,
		_w24267_
	);
	LUT3 #(
		.INIT('h80)
	) name22367 (
		\m2_data_i[26]_pad ,
		_w8699_,
		_w8700_,
		_w24268_
	);
	LUT4 #(
		.INIT('habef)
	) name22368 (
		_w8694_,
		_w8697_,
		_w24267_,
		_w24268_,
		_w24269_
	);
	LUT3 #(
		.INIT('h2a)
	) name22369 (
		\m5_data_i[26]_pad ,
		_w8699_,
		_w8700_,
		_w24270_
	);
	LUT3 #(
		.INIT('h2a)
	) name22370 (
		\m1_data_i[26]_pad ,
		_w8699_,
		_w8700_,
		_w24271_
	);
	LUT4 #(
		.INIT('h57df)
	) name22371 (
		_w8694_,
		_w8697_,
		_w24270_,
		_w24271_,
		_w24272_
	);
	LUT3 #(
		.INIT('h80)
	) name22372 (
		\m0_data_i[26]_pad ,
		_w8699_,
		_w8700_,
		_w24273_
	);
	LUT3 #(
		.INIT('h2a)
	) name22373 (
		\m7_data_i[26]_pad ,
		_w8699_,
		_w8700_,
		_w24274_
	);
	LUT4 #(
		.INIT('h6e7f)
	) name22374 (
		_w8694_,
		_w8697_,
		_w24273_,
		_w24274_,
		_w24275_
	);
	LUT4 #(
		.INIT('h7fff)
	) name22375 (
		_w24266_,
		_w24269_,
		_w24272_,
		_w24275_,
		_w24276_
	);
	LUT3 #(
		.INIT('h2a)
	) name22376 (
		\m3_data_i[27]_pad ,
		_w8699_,
		_w8700_,
		_w24277_
	);
	LUT3 #(
		.INIT('h80)
	) name22377 (
		\m4_data_i[27]_pad ,
		_w8699_,
		_w8700_,
		_w24278_
	);
	LUT4 #(
		.INIT('h9dbf)
	) name22378 (
		_w8694_,
		_w8697_,
		_w24277_,
		_w24278_,
		_w24279_
	);
	LUT3 #(
		.INIT('h80)
	) name22379 (
		\m6_data_i[27]_pad ,
		_w8699_,
		_w8700_,
		_w24280_
	);
	LUT3 #(
		.INIT('h80)
	) name22380 (
		\m2_data_i[27]_pad ,
		_w8699_,
		_w8700_,
		_w24281_
	);
	LUT4 #(
		.INIT('habef)
	) name22381 (
		_w8694_,
		_w8697_,
		_w24280_,
		_w24281_,
		_w24282_
	);
	LUT3 #(
		.INIT('h2a)
	) name22382 (
		\m5_data_i[27]_pad ,
		_w8699_,
		_w8700_,
		_w24283_
	);
	LUT3 #(
		.INIT('h2a)
	) name22383 (
		\m1_data_i[27]_pad ,
		_w8699_,
		_w8700_,
		_w24284_
	);
	LUT4 #(
		.INIT('h57df)
	) name22384 (
		_w8694_,
		_w8697_,
		_w24283_,
		_w24284_,
		_w24285_
	);
	LUT3 #(
		.INIT('h80)
	) name22385 (
		\m0_data_i[27]_pad ,
		_w8699_,
		_w8700_,
		_w24286_
	);
	LUT3 #(
		.INIT('h2a)
	) name22386 (
		\m7_data_i[27]_pad ,
		_w8699_,
		_w8700_,
		_w24287_
	);
	LUT4 #(
		.INIT('h6e7f)
	) name22387 (
		_w8694_,
		_w8697_,
		_w24286_,
		_w24287_,
		_w24288_
	);
	LUT4 #(
		.INIT('h7fff)
	) name22388 (
		_w24279_,
		_w24282_,
		_w24285_,
		_w24288_,
		_w24289_
	);
	LUT3 #(
		.INIT('h2a)
	) name22389 (
		\m3_data_i[28]_pad ,
		_w8699_,
		_w8700_,
		_w24290_
	);
	LUT3 #(
		.INIT('h80)
	) name22390 (
		\m4_data_i[28]_pad ,
		_w8699_,
		_w8700_,
		_w24291_
	);
	LUT4 #(
		.INIT('h9dbf)
	) name22391 (
		_w8694_,
		_w8697_,
		_w24290_,
		_w24291_,
		_w24292_
	);
	LUT3 #(
		.INIT('h80)
	) name22392 (
		\m6_data_i[28]_pad ,
		_w8699_,
		_w8700_,
		_w24293_
	);
	LUT3 #(
		.INIT('h80)
	) name22393 (
		\m2_data_i[28]_pad ,
		_w8699_,
		_w8700_,
		_w24294_
	);
	LUT4 #(
		.INIT('habef)
	) name22394 (
		_w8694_,
		_w8697_,
		_w24293_,
		_w24294_,
		_w24295_
	);
	LUT3 #(
		.INIT('h2a)
	) name22395 (
		\m5_data_i[28]_pad ,
		_w8699_,
		_w8700_,
		_w24296_
	);
	LUT3 #(
		.INIT('h2a)
	) name22396 (
		\m1_data_i[28]_pad ,
		_w8699_,
		_w8700_,
		_w24297_
	);
	LUT4 #(
		.INIT('h57df)
	) name22397 (
		_w8694_,
		_w8697_,
		_w24296_,
		_w24297_,
		_w24298_
	);
	LUT3 #(
		.INIT('h80)
	) name22398 (
		\m0_data_i[28]_pad ,
		_w8699_,
		_w8700_,
		_w24299_
	);
	LUT3 #(
		.INIT('h2a)
	) name22399 (
		\m7_data_i[28]_pad ,
		_w8699_,
		_w8700_,
		_w24300_
	);
	LUT4 #(
		.INIT('h6e7f)
	) name22400 (
		_w8694_,
		_w8697_,
		_w24299_,
		_w24300_,
		_w24301_
	);
	LUT4 #(
		.INIT('h7fff)
	) name22401 (
		_w24292_,
		_w24295_,
		_w24298_,
		_w24301_,
		_w24302_
	);
	LUT3 #(
		.INIT('h2a)
	) name22402 (
		\m3_data_i[29]_pad ,
		_w8699_,
		_w8700_,
		_w24303_
	);
	LUT3 #(
		.INIT('h80)
	) name22403 (
		\m4_data_i[29]_pad ,
		_w8699_,
		_w8700_,
		_w24304_
	);
	LUT4 #(
		.INIT('h9dbf)
	) name22404 (
		_w8694_,
		_w8697_,
		_w24303_,
		_w24304_,
		_w24305_
	);
	LUT3 #(
		.INIT('h80)
	) name22405 (
		\m6_data_i[29]_pad ,
		_w8699_,
		_w8700_,
		_w24306_
	);
	LUT3 #(
		.INIT('h80)
	) name22406 (
		\m2_data_i[29]_pad ,
		_w8699_,
		_w8700_,
		_w24307_
	);
	LUT4 #(
		.INIT('habef)
	) name22407 (
		_w8694_,
		_w8697_,
		_w24306_,
		_w24307_,
		_w24308_
	);
	LUT3 #(
		.INIT('h2a)
	) name22408 (
		\m5_data_i[29]_pad ,
		_w8699_,
		_w8700_,
		_w24309_
	);
	LUT3 #(
		.INIT('h2a)
	) name22409 (
		\m1_data_i[29]_pad ,
		_w8699_,
		_w8700_,
		_w24310_
	);
	LUT4 #(
		.INIT('h57df)
	) name22410 (
		_w8694_,
		_w8697_,
		_w24309_,
		_w24310_,
		_w24311_
	);
	LUT3 #(
		.INIT('h80)
	) name22411 (
		\m0_data_i[29]_pad ,
		_w8699_,
		_w8700_,
		_w24312_
	);
	LUT3 #(
		.INIT('h2a)
	) name22412 (
		\m7_data_i[29]_pad ,
		_w8699_,
		_w8700_,
		_w24313_
	);
	LUT4 #(
		.INIT('h6e7f)
	) name22413 (
		_w8694_,
		_w8697_,
		_w24312_,
		_w24313_,
		_w24314_
	);
	LUT4 #(
		.INIT('h7fff)
	) name22414 (
		_w24305_,
		_w24308_,
		_w24311_,
		_w24314_,
		_w24315_
	);
	LUT3 #(
		.INIT('h2a)
	) name22415 (
		\m3_data_i[2]_pad ,
		_w8699_,
		_w8700_,
		_w24316_
	);
	LUT3 #(
		.INIT('h80)
	) name22416 (
		\m4_data_i[2]_pad ,
		_w8699_,
		_w8700_,
		_w24317_
	);
	LUT4 #(
		.INIT('h9dbf)
	) name22417 (
		_w8694_,
		_w8697_,
		_w24316_,
		_w24317_,
		_w24318_
	);
	LUT3 #(
		.INIT('h80)
	) name22418 (
		\m0_data_i[2]_pad ,
		_w8699_,
		_w8700_,
		_w24319_
	);
	LUT3 #(
		.INIT('h2a)
	) name22419 (
		\m5_data_i[2]_pad ,
		_w8699_,
		_w8700_,
		_w24320_
	);
	LUT4 #(
		.INIT('h5d7f)
	) name22420 (
		_w8694_,
		_w8697_,
		_w24319_,
		_w24320_,
		_w24321_
	);
	LUT3 #(
		.INIT('h2a)
	) name22421 (
		\m7_data_i[2]_pad ,
		_w8699_,
		_w8700_,
		_w24322_
	);
	LUT3 #(
		.INIT('h80)
	) name22422 (
		\m6_data_i[2]_pad ,
		_w8699_,
		_w8700_,
		_w24323_
	);
	LUT3 #(
		.INIT('h57)
	) name22423 (
		_w8712_,
		_w24322_,
		_w24323_,
		_w24324_
	);
	LUT3 #(
		.INIT('h2a)
	) name22424 (
		\m1_data_i[2]_pad ,
		_w8699_,
		_w8700_,
		_w24325_
	);
	LUT3 #(
		.INIT('h80)
	) name22425 (
		\m2_data_i[2]_pad ,
		_w8699_,
		_w8700_,
		_w24326_
	);
	LUT4 #(
		.INIT('h3b7f)
	) name22426 (
		_w8694_,
		_w8697_,
		_w24325_,
		_w24326_,
		_w24327_
	);
	LUT4 #(
		.INIT('h7fff)
	) name22427 (
		_w24318_,
		_w24321_,
		_w24324_,
		_w24327_,
		_w24328_
	);
	LUT3 #(
		.INIT('h2a)
	) name22428 (
		\m3_data_i[30]_pad ,
		_w8699_,
		_w8700_,
		_w24329_
	);
	LUT3 #(
		.INIT('h80)
	) name22429 (
		\m4_data_i[30]_pad ,
		_w8699_,
		_w8700_,
		_w24330_
	);
	LUT4 #(
		.INIT('h9dbf)
	) name22430 (
		_w8694_,
		_w8697_,
		_w24329_,
		_w24330_,
		_w24331_
	);
	LUT3 #(
		.INIT('h80)
	) name22431 (
		\m6_data_i[30]_pad ,
		_w8699_,
		_w8700_,
		_w24332_
	);
	LUT3 #(
		.INIT('h80)
	) name22432 (
		\m2_data_i[30]_pad ,
		_w8699_,
		_w8700_,
		_w24333_
	);
	LUT4 #(
		.INIT('habef)
	) name22433 (
		_w8694_,
		_w8697_,
		_w24332_,
		_w24333_,
		_w24334_
	);
	LUT3 #(
		.INIT('h2a)
	) name22434 (
		\m5_data_i[30]_pad ,
		_w8699_,
		_w8700_,
		_w24335_
	);
	LUT3 #(
		.INIT('h2a)
	) name22435 (
		\m1_data_i[30]_pad ,
		_w8699_,
		_w8700_,
		_w24336_
	);
	LUT4 #(
		.INIT('h57df)
	) name22436 (
		_w8694_,
		_w8697_,
		_w24335_,
		_w24336_,
		_w24337_
	);
	LUT3 #(
		.INIT('h80)
	) name22437 (
		\m0_data_i[30]_pad ,
		_w8699_,
		_w8700_,
		_w24338_
	);
	LUT3 #(
		.INIT('h2a)
	) name22438 (
		\m7_data_i[30]_pad ,
		_w8699_,
		_w8700_,
		_w24339_
	);
	LUT4 #(
		.INIT('h6e7f)
	) name22439 (
		_w8694_,
		_w8697_,
		_w24338_,
		_w24339_,
		_w24340_
	);
	LUT4 #(
		.INIT('h7fff)
	) name22440 (
		_w24331_,
		_w24334_,
		_w24337_,
		_w24340_,
		_w24341_
	);
	LUT3 #(
		.INIT('h2a)
	) name22441 (
		\m3_data_i[31]_pad ,
		_w8699_,
		_w8700_,
		_w24342_
	);
	LUT3 #(
		.INIT('h80)
	) name22442 (
		\m4_data_i[31]_pad ,
		_w8699_,
		_w8700_,
		_w24343_
	);
	LUT4 #(
		.INIT('h9dbf)
	) name22443 (
		_w8694_,
		_w8697_,
		_w24342_,
		_w24343_,
		_w24344_
	);
	LUT3 #(
		.INIT('h80)
	) name22444 (
		\m6_data_i[31]_pad ,
		_w8699_,
		_w8700_,
		_w24345_
	);
	LUT3 #(
		.INIT('h80)
	) name22445 (
		\m2_data_i[31]_pad ,
		_w8699_,
		_w8700_,
		_w24346_
	);
	LUT4 #(
		.INIT('habef)
	) name22446 (
		_w8694_,
		_w8697_,
		_w24345_,
		_w24346_,
		_w24347_
	);
	LUT3 #(
		.INIT('h2a)
	) name22447 (
		\m5_data_i[31]_pad ,
		_w8699_,
		_w8700_,
		_w24348_
	);
	LUT3 #(
		.INIT('h2a)
	) name22448 (
		\m1_data_i[31]_pad ,
		_w8699_,
		_w8700_,
		_w24349_
	);
	LUT4 #(
		.INIT('h57df)
	) name22449 (
		_w8694_,
		_w8697_,
		_w24348_,
		_w24349_,
		_w24350_
	);
	LUT3 #(
		.INIT('h80)
	) name22450 (
		\m0_data_i[31]_pad ,
		_w8699_,
		_w8700_,
		_w24351_
	);
	LUT3 #(
		.INIT('h2a)
	) name22451 (
		\m7_data_i[31]_pad ,
		_w8699_,
		_w8700_,
		_w24352_
	);
	LUT4 #(
		.INIT('h6e7f)
	) name22452 (
		_w8694_,
		_w8697_,
		_w24351_,
		_w24352_,
		_w24353_
	);
	LUT4 #(
		.INIT('h7fff)
	) name22453 (
		_w24344_,
		_w24347_,
		_w24350_,
		_w24353_,
		_w24354_
	);
	LUT3 #(
		.INIT('h2a)
	) name22454 (
		\m3_data_i[3]_pad ,
		_w8699_,
		_w8700_,
		_w24355_
	);
	LUT3 #(
		.INIT('h80)
	) name22455 (
		\m4_data_i[3]_pad ,
		_w8699_,
		_w8700_,
		_w24356_
	);
	LUT4 #(
		.INIT('h9dbf)
	) name22456 (
		_w8694_,
		_w8697_,
		_w24355_,
		_w24356_,
		_w24357_
	);
	LUT3 #(
		.INIT('h2a)
	) name22457 (
		\m1_data_i[3]_pad ,
		_w8699_,
		_w8700_,
		_w24358_
	);
	LUT3 #(
		.INIT('h2a)
	) name22458 (
		\m7_data_i[3]_pad ,
		_w8699_,
		_w8700_,
		_w24359_
	);
	LUT4 #(
		.INIT('h6e7f)
	) name22459 (
		_w8694_,
		_w8697_,
		_w24358_,
		_w24359_,
		_w24360_
	);
	LUT3 #(
		.INIT('h80)
	) name22460 (
		\m2_data_i[3]_pad ,
		_w8699_,
		_w8700_,
		_w24361_
	);
	LUT3 #(
		.INIT('h80)
	) name22461 (
		\m0_data_i[3]_pad ,
		_w8699_,
		_w8700_,
		_w24362_
	);
	LUT4 #(
		.INIT('h37bf)
	) name22462 (
		_w8694_,
		_w8697_,
		_w24361_,
		_w24362_,
		_w24363_
	);
	LUT3 #(
		.INIT('h80)
	) name22463 (
		\m6_data_i[3]_pad ,
		_w8699_,
		_w8700_,
		_w24364_
	);
	LUT3 #(
		.INIT('h2a)
	) name22464 (
		\m5_data_i[3]_pad ,
		_w8699_,
		_w8700_,
		_w24365_
	);
	LUT4 #(
		.INIT('hcdef)
	) name22465 (
		_w8694_,
		_w8697_,
		_w24364_,
		_w24365_,
		_w24366_
	);
	LUT4 #(
		.INIT('h7fff)
	) name22466 (
		_w24357_,
		_w24360_,
		_w24363_,
		_w24366_,
		_w24367_
	);
	LUT3 #(
		.INIT('h2a)
	) name22467 (
		\m3_data_i[4]_pad ,
		_w8699_,
		_w8700_,
		_w24368_
	);
	LUT3 #(
		.INIT('h80)
	) name22468 (
		\m4_data_i[4]_pad ,
		_w8699_,
		_w8700_,
		_w24369_
	);
	LUT4 #(
		.INIT('h9dbf)
	) name22469 (
		_w8694_,
		_w8697_,
		_w24368_,
		_w24369_,
		_w24370_
	);
	LUT3 #(
		.INIT('h2a)
	) name22470 (
		\m1_data_i[4]_pad ,
		_w8699_,
		_w8700_,
		_w24371_
	);
	LUT3 #(
		.INIT('h2a)
	) name22471 (
		\m7_data_i[4]_pad ,
		_w8699_,
		_w8700_,
		_w24372_
	);
	LUT4 #(
		.INIT('h6e7f)
	) name22472 (
		_w8694_,
		_w8697_,
		_w24371_,
		_w24372_,
		_w24373_
	);
	LUT3 #(
		.INIT('h80)
	) name22473 (
		\m2_data_i[4]_pad ,
		_w8699_,
		_w8700_,
		_w24374_
	);
	LUT3 #(
		.INIT('h80)
	) name22474 (
		\m0_data_i[4]_pad ,
		_w8699_,
		_w8700_,
		_w24375_
	);
	LUT4 #(
		.INIT('h37bf)
	) name22475 (
		_w8694_,
		_w8697_,
		_w24374_,
		_w24375_,
		_w24376_
	);
	LUT3 #(
		.INIT('h80)
	) name22476 (
		\m6_data_i[4]_pad ,
		_w8699_,
		_w8700_,
		_w24377_
	);
	LUT3 #(
		.INIT('h2a)
	) name22477 (
		\m5_data_i[4]_pad ,
		_w8699_,
		_w8700_,
		_w24378_
	);
	LUT4 #(
		.INIT('hcdef)
	) name22478 (
		_w8694_,
		_w8697_,
		_w24377_,
		_w24378_,
		_w24379_
	);
	LUT4 #(
		.INIT('h7fff)
	) name22479 (
		_w24370_,
		_w24373_,
		_w24376_,
		_w24379_,
		_w24380_
	);
	LUT3 #(
		.INIT('h2a)
	) name22480 (
		\m3_data_i[5]_pad ,
		_w8699_,
		_w8700_,
		_w24381_
	);
	LUT3 #(
		.INIT('h80)
	) name22481 (
		\m4_data_i[5]_pad ,
		_w8699_,
		_w8700_,
		_w24382_
	);
	LUT4 #(
		.INIT('h9dbf)
	) name22482 (
		_w8694_,
		_w8697_,
		_w24381_,
		_w24382_,
		_w24383_
	);
	LUT3 #(
		.INIT('h80)
	) name22483 (
		\m6_data_i[5]_pad ,
		_w8699_,
		_w8700_,
		_w24384_
	);
	LUT3 #(
		.INIT('h80)
	) name22484 (
		\m2_data_i[5]_pad ,
		_w8699_,
		_w8700_,
		_w24385_
	);
	LUT4 #(
		.INIT('habef)
	) name22485 (
		_w8694_,
		_w8697_,
		_w24384_,
		_w24385_,
		_w24386_
	);
	LUT3 #(
		.INIT('h2a)
	) name22486 (
		\m5_data_i[5]_pad ,
		_w8699_,
		_w8700_,
		_w24387_
	);
	LUT3 #(
		.INIT('h2a)
	) name22487 (
		\m1_data_i[5]_pad ,
		_w8699_,
		_w8700_,
		_w24388_
	);
	LUT4 #(
		.INIT('h57df)
	) name22488 (
		_w8694_,
		_w8697_,
		_w24387_,
		_w24388_,
		_w24389_
	);
	LUT3 #(
		.INIT('h80)
	) name22489 (
		\m0_data_i[5]_pad ,
		_w8699_,
		_w8700_,
		_w24390_
	);
	LUT3 #(
		.INIT('h2a)
	) name22490 (
		\m7_data_i[5]_pad ,
		_w8699_,
		_w8700_,
		_w24391_
	);
	LUT4 #(
		.INIT('h6e7f)
	) name22491 (
		_w8694_,
		_w8697_,
		_w24390_,
		_w24391_,
		_w24392_
	);
	LUT4 #(
		.INIT('h7fff)
	) name22492 (
		_w24383_,
		_w24386_,
		_w24389_,
		_w24392_,
		_w24393_
	);
	LUT3 #(
		.INIT('h2a)
	) name22493 (
		\m3_data_i[6]_pad ,
		_w8699_,
		_w8700_,
		_w24394_
	);
	LUT3 #(
		.INIT('h80)
	) name22494 (
		\m4_data_i[6]_pad ,
		_w8699_,
		_w8700_,
		_w24395_
	);
	LUT4 #(
		.INIT('h9dbf)
	) name22495 (
		_w8694_,
		_w8697_,
		_w24394_,
		_w24395_,
		_w24396_
	);
	LUT3 #(
		.INIT('h80)
	) name22496 (
		\m6_data_i[6]_pad ,
		_w8699_,
		_w8700_,
		_w24397_
	);
	LUT3 #(
		.INIT('h80)
	) name22497 (
		\m2_data_i[6]_pad ,
		_w8699_,
		_w8700_,
		_w24398_
	);
	LUT4 #(
		.INIT('habef)
	) name22498 (
		_w8694_,
		_w8697_,
		_w24397_,
		_w24398_,
		_w24399_
	);
	LUT3 #(
		.INIT('h2a)
	) name22499 (
		\m5_data_i[6]_pad ,
		_w8699_,
		_w8700_,
		_w24400_
	);
	LUT3 #(
		.INIT('h2a)
	) name22500 (
		\m1_data_i[6]_pad ,
		_w8699_,
		_w8700_,
		_w24401_
	);
	LUT4 #(
		.INIT('h57df)
	) name22501 (
		_w8694_,
		_w8697_,
		_w24400_,
		_w24401_,
		_w24402_
	);
	LUT3 #(
		.INIT('h80)
	) name22502 (
		\m0_data_i[6]_pad ,
		_w8699_,
		_w8700_,
		_w24403_
	);
	LUT3 #(
		.INIT('h2a)
	) name22503 (
		\m7_data_i[6]_pad ,
		_w8699_,
		_w8700_,
		_w24404_
	);
	LUT4 #(
		.INIT('h6e7f)
	) name22504 (
		_w8694_,
		_w8697_,
		_w24403_,
		_w24404_,
		_w24405_
	);
	LUT4 #(
		.INIT('h7fff)
	) name22505 (
		_w24396_,
		_w24399_,
		_w24402_,
		_w24405_,
		_w24406_
	);
	LUT3 #(
		.INIT('h2a)
	) name22506 (
		\m3_data_i[7]_pad ,
		_w8699_,
		_w8700_,
		_w24407_
	);
	LUT3 #(
		.INIT('h80)
	) name22507 (
		\m4_data_i[7]_pad ,
		_w8699_,
		_w8700_,
		_w24408_
	);
	LUT4 #(
		.INIT('h9dbf)
	) name22508 (
		_w8694_,
		_w8697_,
		_w24407_,
		_w24408_,
		_w24409_
	);
	LUT3 #(
		.INIT('h80)
	) name22509 (
		\m6_data_i[7]_pad ,
		_w8699_,
		_w8700_,
		_w24410_
	);
	LUT3 #(
		.INIT('h80)
	) name22510 (
		\m2_data_i[7]_pad ,
		_w8699_,
		_w8700_,
		_w24411_
	);
	LUT4 #(
		.INIT('habef)
	) name22511 (
		_w8694_,
		_w8697_,
		_w24410_,
		_w24411_,
		_w24412_
	);
	LUT3 #(
		.INIT('h2a)
	) name22512 (
		\m5_data_i[7]_pad ,
		_w8699_,
		_w8700_,
		_w24413_
	);
	LUT3 #(
		.INIT('h2a)
	) name22513 (
		\m1_data_i[7]_pad ,
		_w8699_,
		_w8700_,
		_w24414_
	);
	LUT4 #(
		.INIT('h57df)
	) name22514 (
		_w8694_,
		_w8697_,
		_w24413_,
		_w24414_,
		_w24415_
	);
	LUT3 #(
		.INIT('h80)
	) name22515 (
		\m0_data_i[7]_pad ,
		_w8699_,
		_w8700_,
		_w24416_
	);
	LUT3 #(
		.INIT('h2a)
	) name22516 (
		\m7_data_i[7]_pad ,
		_w8699_,
		_w8700_,
		_w24417_
	);
	LUT4 #(
		.INIT('h6e7f)
	) name22517 (
		_w8694_,
		_w8697_,
		_w24416_,
		_w24417_,
		_w24418_
	);
	LUT4 #(
		.INIT('h7fff)
	) name22518 (
		_w24409_,
		_w24412_,
		_w24415_,
		_w24418_,
		_w24419_
	);
	LUT3 #(
		.INIT('h2a)
	) name22519 (
		\m3_data_i[8]_pad ,
		_w8699_,
		_w8700_,
		_w24420_
	);
	LUT3 #(
		.INIT('h80)
	) name22520 (
		\m4_data_i[8]_pad ,
		_w8699_,
		_w8700_,
		_w24421_
	);
	LUT4 #(
		.INIT('h9dbf)
	) name22521 (
		_w8694_,
		_w8697_,
		_w24420_,
		_w24421_,
		_w24422_
	);
	LUT3 #(
		.INIT('h80)
	) name22522 (
		\m6_data_i[8]_pad ,
		_w8699_,
		_w8700_,
		_w24423_
	);
	LUT3 #(
		.INIT('h80)
	) name22523 (
		\m2_data_i[8]_pad ,
		_w8699_,
		_w8700_,
		_w24424_
	);
	LUT4 #(
		.INIT('habef)
	) name22524 (
		_w8694_,
		_w8697_,
		_w24423_,
		_w24424_,
		_w24425_
	);
	LUT3 #(
		.INIT('h2a)
	) name22525 (
		\m5_data_i[8]_pad ,
		_w8699_,
		_w8700_,
		_w24426_
	);
	LUT3 #(
		.INIT('h2a)
	) name22526 (
		\m1_data_i[8]_pad ,
		_w8699_,
		_w8700_,
		_w24427_
	);
	LUT4 #(
		.INIT('h57df)
	) name22527 (
		_w8694_,
		_w8697_,
		_w24426_,
		_w24427_,
		_w24428_
	);
	LUT3 #(
		.INIT('h80)
	) name22528 (
		\m0_data_i[8]_pad ,
		_w8699_,
		_w8700_,
		_w24429_
	);
	LUT3 #(
		.INIT('h2a)
	) name22529 (
		\m7_data_i[8]_pad ,
		_w8699_,
		_w8700_,
		_w24430_
	);
	LUT4 #(
		.INIT('h6e7f)
	) name22530 (
		_w8694_,
		_w8697_,
		_w24429_,
		_w24430_,
		_w24431_
	);
	LUT4 #(
		.INIT('h7fff)
	) name22531 (
		_w24422_,
		_w24425_,
		_w24428_,
		_w24431_,
		_w24432_
	);
	LUT3 #(
		.INIT('h2a)
	) name22532 (
		\m3_data_i[9]_pad ,
		_w8699_,
		_w8700_,
		_w24433_
	);
	LUT3 #(
		.INIT('h80)
	) name22533 (
		\m4_data_i[9]_pad ,
		_w8699_,
		_w8700_,
		_w24434_
	);
	LUT4 #(
		.INIT('h9dbf)
	) name22534 (
		_w8694_,
		_w8697_,
		_w24433_,
		_w24434_,
		_w24435_
	);
	LUT3 #(
		.INIT('h80)
	) name22535 (
		\m6_data_i[9]_pad ,
		_w8699_,
		_w8700_,
		_w24436_
	);
	LUT3 #(
		.INIT('h80)
	) name22536 (
		\m2_data_i[9]_pad ,
		_w8699_,
		_w8700_,
		_w24437_
	);
	LUT4 #(
		.INIT('habef)
	) name22537 (
		_w8694_,
		_w8697_,
		_w24436_,
		_w24437_,
		_w24438_
	);
	LUT3 #(
		.INIT('h2a)
	) name22538 (
		\m5_data_i[9]_pad ,
		_w8699_,
		_w8700_,
		_w24439_
	);
	LUT3 #(
		.INIT('h2a)
	) name22539 (
		\m1_data_i[9]_pad ,
		_w8699_,
		_w8700_,
		_w24440_
	);
	LUT4 #(
		.INIT('h57df)
	) name22540 (
		_w8694_,
		_w8697_,
		_w24439_,
		_w24440_,
		_w24441_
	);
	LUT3 #(
		.INIT('h80)
	) name22541 (
		\m0_data_i[9]_pad ,
		_w8699_,
		_w8700_,
		_w24442_
	);
	LUT3 #(
		.INIT('h2a)
	) name22542 (
		\m7_data_i[9]_pad ,
		_w8699_,
		_w8700_,
		_w24443_
	);
	LUT4 #(
		.INIT('h6e7f)
	) name22543 (
		_w8694_,
		_w8697_,
		_w24442_,
		_w24443_,
		_w24444_
	);
	LUT4 #(
		.INIT('h7fff)
	) name22544 (
		_w24435_,
		_w24438_,
		_w24441_,
		_w24444_,
		_w24445_
	);
	LUT3 #(
		.INIT('h2a)
	) name22545 (
		\m1_sel_i[0]_pad ,
		_w8699_,
		_w8700_,
		_w24446_
	);
	LUT3 #(
		.INIT('h80)
	) name22546 (
		\m2_sel_i[0]_pad ,
		_w8699_,
		_w8700_,
		_w24447_
	);
	LUT4 #(
		.INIT('h3b7f)
	) name22547 (
		_w8694_,
		_w8697_,
		_w24446_,
		_w24447_,
		_w24448_
	);
	LUT3 #(
		.INIT('h80)
	) name22548 (
		\m0_sel_i[0]_pad ,
		_w8699_,
		_w8700_,
		_w24449_
	);
	LUT3 #(
		.INIT('h80)
	) name22549 (
		\m4_sel_i[0]_pad ,
		_w8699_,
		_w8700_,
		_w24450_
	);
	LUT4 #(
		.INIT('h5d7f)
	) name22550 (
		_w8694_,
		_w8697_,
		_w24449_,
		_w24450_,
		_w24451_
	);
	LUT3 #(
		.INIT('h2a)
	) name22551 (
		\m7_sel_i[0]_pad ,
		_w8699_,
		_w8700_,
		_w24452_
	);
	LUT3 #(
		.INIT('h2a)
	) name22552 (
		\m3_sel_i[0]_pad ,
		_w8699_,
		_w8700_,
		_w24453_
	);
	LUT4 #(
		.INIT('habef)
	) name22553 (
		_w8694_,
		_w8697_,
		_w24452_,
		_w24453_,
		_w24454_
	);
	LUT3 #(
		.INIT('h80)
	) name22554 (
		\m6_sel_i[0]_pad ,
		_w8699_,
		_w8700_,
		_w24455_
	);
	LUT3 #(
		.INIT('h2a)
	) name22555 (
		\m5_sel_i[0]_pad ,
		_w8699_,
		_w8700_,
		_w24456_
	);
	LUT4 #(
		.INIT('hcdef)
	) name22556 (
		_w8694_,
		_w8697_,
		_w24455_,
		_w24456_,
		_w24457_
	);
	LUT4 #(
		.INIT('h7fff)
	) name22557 (
		_w24448_,
		_w24451_,
		_w24454_,
		_w24457_,
		_w24458_
	);
	LUT3 #(
		.INIT('h80)
	) name22558 (
		\m0_sel_i[1]_pad ,
		_w8699_,
		_w8700_,
		_w24459_
	);
	LUT3 #(
		.INIT('h2a)
	) name22559 (
		\m7_sel_i[1]_pad ,
		_w8699_,
		_w8700_,
		_w24460_
	);
	LUT4 #(
		.INIT('h6e7f)
	) name22560 (
		_w8694_,
		_w8697_,
		_w24459_,
		_w24460_,
		_w24461_
	);
	LUT3 #(
		.INIT('h2a)
	) name22561 (
		\m3_sel_i[1]_pad ,
		_w8699_,
		_w8700_,
		_w24462_
	);
	LUT3 #(
		.INIT('h80)
	) name22562 (
		\m2_sel_i[1]_pad ,
		_w8699_,
		_w8700_,
		_w24463_
	);
	LUT3 #(
		.INIT('h57)
	) name22563 (
		_w8698_,
		_w24462_,
		_w24463_,
		_w24464_
	);
	LUT3 #(
		.INIT('h80)
	) name22564 (
		\m4_sel_i[1]_pad ,
		_w8699_,
		_w8700_,
		_w24465_
	);
	LUT3 #(
		.INIT('h2a)
	) name22565 (
		\m1_sel_i[1]_pad ,
		_w8699_,
		_w8700_,
		_w24466_
	);
	LUT4 #(
		.INIT('h57df)
	) name22566 (
		_w8694_,
		_w8697_,
		_w24465_,
		_w24466_,
		_w24467_
	);
	LUT3 #(
		.INIT('h80)
	) name22567 (
		\m6_sel_i[1]_pad ,
		_w8699_,
		_w8700_,
		_w24468_
	);
	LUT3 #(
		.INIT('h2a)
	) name22568 (
		\m5_sel_i[1]_pad ,
		_w8699_,
		_w8700_,
		_w24469_
	);
	LUT4 #(
		.INIT('hcdef)
	) name22569 (
		_w8694_,
		_w8697_,
		_w24468_,
		_w24469_,
		_w24470_
	);
	LUT4 #(
		.INIT('h7fff)
	) name22570 (
		_w24461_,
		_w24464_,
		_w24467_,
		_w24470_,
		_w24471_
	);
	LUT3 #(
		.INIT('h2a)
	) name22571 (
		\m1_sel_i[2]_pad ,
		_w8699_,
		_w8700_,
		_w24472_
	);
	LUT3 #(
		.INIT('h80)
	) name22572 (
		\m2_sel_i[2]_pad ,
		_w8699_,
		_w8700_,
		_w24473_
	);
	LUT4 #(
		.INIT('h3b7f)
	) name22573 (
		_w8694_,
		_w8697_,
		_w24472_,
		_w24473_,
		_w24474_
	);
	LUT3 #(
		.INIT('h80)
	) name22574 (
		\m0_sel_i[2]_pad ,
		_w8699_,
		_w8700_,
		_w24475_
	);
	LUT3 #(
		.INIT('h80)
	) name22575 (
		\m4_sel_i[2]_pad ,
		_w8699_,
		_w8700_,
		_w24476_
	);
	LUT4 #(
		.INIT('h5d7f)
	) name22576 (
		_w8694_,
		_w8697_,
		_w24475_,
		_w24476_,
		_w24477_
	);
	LUT3 #(
		.INIT('h2a)
	) name22577 (
		\m7_sel_i[2]_pad ,
		_w8699_,
		_w8700_,
		_w24478_
	);
	LUT3 #(
		.INIT('h2a)
	) name22578 (
		\m3_sel_i[2]_pad ,
		_w8699_,
		_w8700_,
		_w24479_
	);
	LUT4 #(
		.INIT('habef)
	) name22579 (
		_w8694_,
		_w8697_,
		_w24478_,
		_w24479_,
		_w24480_
	);
	LUT3 #(
		.INIT('h80)
	) name22580 (
		\m6_sel_i[2]_pad ,
		_w8699_,
		_w8700_,
		_w24481_
	);
	LUT3 #(
		.INIT('h2a)
	) name22581 (
		\m5_sel_i[2]_pad ,
		_w8699_,
		_w8700_,
		_w24482_
	);
	LUT4 #(
		.INIT('hcdef)
	) name22582 (
		_w8694_,
		_w8697_,
		_w24481_,
		_w24482_,
		_w24483_
	);
	LUT4 #(
		.INIT('h7fff)
	) name22583 (
		_w24474_,
		_w24477_,
		_w24480_,
		_w24483_,
		_w24484_
	);
	LUT3 #(
		.INIT('h80)
	) name22584 (
		\m0_sel_i[3]_pad ,
		_w8699_,
		_w8700_,
		_w24485_
	);
	LUT3 #(
		.INIT('h2a)
	) name22585 (
		\m7_sel_i[3]_pad ,
		_w8699_,
		_w8700_,
		_w24486_
	);
	LUT4 #(
		.INIT('h6e7f)
	) name22586 (
		_w8694_,
		_w8697_,
		_w24485_,
		_w24486_,
		_w24487_
	);
	LUT3 #(
		.INIT('h80)
	) name22587 (
		\m6_sel_i[3]_pad ,
		_w8699_,
		_w8700_,
		_w24488_
	);
	LUT3 #(
		.INIT('h80)
	) name22588 (
		\m2_sel_i[3]_pad ,
		_w8699_,
		_w8700_,
		_w24489_
	);
	LUT4 #(
		.INIT('habef)
	) name22589 (
		_w8694_,
		_w8697_,
		_w24488_,
		_w24489_,
		_w24490_
	);
	LUT3 #(
		.INIT('h2a)
	) name22590 (
		\m5_sel_i[3]_pad ,
		_w8699_,
		_w8700_,
		_w24491_
	);
	LUT3 #(
		.INIT('h2a)
	) name22591 (
		\m1_sel_i[3]_pad ,
		_w8699_,
		_w8700_,
		_w24492_
	);
	LUT4 #(
		.INIT('h57df)
	) name22592 (
		_w8694_,
		_w8697_,
		_w24491_,
		_w24492_,
		_w24493_
	);
	LUT3 #(
		.INIT('h2a)
	) name22593 (
		\m3_sel_i[3]_pad ,
		_w8699_,
		_w8700_,
		_w24494_
	);
	LUT3 #(
		.INIT('h80)
	) name22594 (
		\m4_sel_i[3]_pad ,
		_w8699_,
		_w8700_,
		_w24495_
	);
	LUT4 #(
		.INIT('h9dbf)
	) name22595 (
		_w8694_,
		_w8697_,
		_w24494_,
		_w24495_,
		_w24496_
	);
	LUT4 #(
		.INIT('h7fff)
	) name22596 (
		_w24487_,
		_w24490_,
		_w24493_,
		_w24496_,
		_w24497_
	);
	LUT4 #(
		.INIT('h2a00)
	) name22597 (
		\m5_stb_i_pad ,
		_w8699_,
		_w8700_,
		_w9547_,
		_w24498_
	);
	LUT4 #(
		.INIT('h8000)
	) name22598 (
		\m4_stb_i_pad ,
		_w8699_,
		_w8700_,
		_w9526_,
		_w24499_
	);
	LUT3 #(
		.INIT('h57)
	) name22599 (
		_w8706_,
		_w24498_,
		_w24499_,
		_w24500_
	);
	LUT4 #(
		.INIT('h8000)
	) name22600 (
		\m2_stb_i_pad ,
		_w8699_,
		_w8700_,
		_w9471_,
		_w24501_
	);
	LUT4 #(
		.INIT('h2a00)
	) name22601 (
		\m1_stb_i_pad ,
		_w8699_,
		_w8700_,
		_w9436_,
		_w24502_
	);
	LUT4 #(
		.INIT('h37bf)
	) name22602 (
		_w8694_,
		_w8697_,
		_w24501_,
		_w24502_,
		_w24503_
	);
	LUT4 #(
		.INIT('h2a00)
	) name22603 (
		\m3_stb_i_pad ,
		_w8699_,
		_w8700_,
		_w9387_,
		_w24504_
	);
	LUT4 #(
		.INIT('h2a00)
	) name22604 (
		\m7_stb_i_pad ,
		_w8699_,
		_w8700_,
		_w9333_,
		_w24505_
	);
	LUT4 #(
		.INIT('haebf)
	) name22605 (
		_w8694_,
		_w8697_,
		_w24504_,
		_w24505_,
		_w24506_
	);
	LUT4 #(
		.INIT('h8000)
	) name22606 (
		\m6_stb_i_pad ,
		_w8699_,
		_w8700_,
		_w9585_,
		_w24507_
	);
	LUT4 #(
		.INIT('h8000)
	) name22607 (
		\m0_stb_i_pad ,
		_w8699_,
		_w8700_,
		_w9401_,
		_w24508_
	);
	LUT4 #(
		.INIT('h67ef)
	) name22608 (
		_w8694_,
		_w8697_,
		_w24507_,
		_w24508_,
		_w24509_
	);
	LUT4 #(
		.INIT('h7fff)
	) name22609 (
		_w24500_,
		_w24503_,
		_w24506_,
		_w24509_,
		_w24510_
	);
	LUT3 #(
		.INIT('h2a)
	) name22610 (
		\m1_we_i_pad ,
		_w8699_,
		_w8700_,
		_w24511_
	);
	LUT3 #(
		.INIT('h80)
	) name22611 (
		\m2_we_i_pad ,
		_w8699_,
		_w8700_,
		_w24512_
	);
	LUT4 #(
		.INIT('h3b7f)
	) name22612 (
		_w8694_,
		_w8697_,
		_w24511_,
		_w24512_,
		_w24513_
	);
	LUT3 #(
		.INIT('h80)
	) name22613 (
		\m0_we_i_pad ,
		_w8699_,
		_w8700_,
		_w24514_
	);
	LUT3 #(
		.INIT('h80)
	) name22614 (
		\m4_we_i_pad ,
		_w8699_,
		_w8700_,
		_w24515_
	);
	LUT4 #(
		.INIT('h5d7f)
	) name22615 (
		_w8694_,
		_w8697_,
		_w24514_,
		_w24515_,
		_w24516_
	);
	LUT3 #(
		.INIT('h2a)
	) name22616 (
		\m7_we_i_pad ,
		_w8699_,
		_w8700_,
		_w24517_
	);
	LUT3 #(
		.INIT('h2a)
	) name22617 (
		\m3_we_i_pad ,
		_w8699_,
		_w8700_,
		_w24518_
	);
	LUT4 #(
		.INIT('habef)
	) name22618 (
		_w8694_,
		_w8697_,
		_w24517_,
		_w24518_,
		_w24519_
	);
	LUT3 #(
		.INIT('h80)
	) name22619 (
		\m6_we_i_pad ,
		_w8699_,
		_w8700_,
		_w24520_
	);
	LUT3 #(
		.INIT('h2a)
	) name22620 (
		\m5_we_i_pad ,
		_w8699_,
		_w8700_,
		_w24521_
	);
	LUT4 #(
		.INIT('hcdef)
	) name22621 (
		_w8694_,
		_w8697_,
		_w24520_,
		_w24521_,
		_w24522_
	);
	LUT4 #(
		.INIT('h7fff)
	) name22622 (
		_w24513_,
		_w24516_,
		_w24519_,
		_w24522_,
		_w24523_
	);
	LUT3 #(
		.INIT('h2a)
	) name22623 (
		\m1_addr_i[0]_pad ,
		_w8743_,
		_w8744_,
		_w24524_
	);
	LUT3 #(
		.INIT('h80)
	) name22624 (
		\m2_addr_i[0]_pad ,
		_w8743_,
		_w8744_,
		_w24525_
	);
	LUT4 #(
		.INIT('h3b7f)
	) name22625 (
		_w8738_,
		_w8741_,
		_w24524_,
		_w24525_,
		_w24526_
	);
	LUT3 #(
		.INIT('h80)
	) name22626 (
		\m6_addr_i[0]_pad ,
		_w8743_,
		_w8744_,
		_w24527_
	);
	LUT3 #(
		.INIT('h2a)
	) name22627 (
		\m7_addr_i[0]_pad ,
		_w8743_,
		_w8744_,
		_w24528_
	);
	LUT3 #(
		.INIT('h57)
	) name22628 (
		_w8756_,
		_w24527_,
		_w24528_,
		_w24529_
	);
	LUT3 #(
		.INIT('h2a)
	) name22629 (
		\m5_addr_i[0]_pad ,
		_w8743_,
		_w8744_,
		_w24530_
	);
	LUT3 #(
		.INIT('h80)
	) name22630 (
		\m0_addr_i[0]_pad ,
		_w8743_,
		_w8744_,
		_w24531_
	);
	LUT4 #(
		.INIT('h57df)
	) name22631 (
		_w8738_,
		_w8741_,
		_w24530_,
		_w24531_,
		_w24532_
	);
	LUT3 #(
		.INIT('h2a)
	) name22632 (
		\m3_addr_i[0]_pad ,
		_w8743_,
		_w8744_,
		_w24533_
	);
	LUT3 #(
		.INIT('h80)
	) name22633 (
		\m4_addr_i[0]_pad ,
		_w8743_,
		_w8744_,
		_w24534_
	);
	LUT4 #(
		.INIT('h9dbf)
	) name22634 (
		_w8738_,
		_w8741_,
		_w24533_,
		_w24534_,
		_w24535_
	);
	LUT4 #(
		.INIT('h7fff)
	) name22635 (
		_w24526_,
		_w24529_,
		_w24532_,
		_w24535_,
		_w24536_
	);
	LUT3 #(
		.INIT('h2a)
	) name22636 (
		\m3_addr_i[10]_pad ,
		_w8743_,
		_w8744_,
		_w24537_
	);
	LUT3 #(
		.INIT('h80)
	) name22637 (
		\m4_addr_i[10]_pad ,
		_w8743_,
		_w8744_,
		_w24538_
	);
	LUT4 #(
		.INIT('h9dbf)
	) name22638 (
		_w8738_,
		_w8741_,
		_w24537_,
		_w24538_,
		_w24539_
	);
	LUT3 #(
		.INIT('h80)
	) name22639 (
		\m6_addr_i[10]_pad ,
		_w8743_,
		_w8744_,
		_w24540_
	);
	LUT3 #(
		.INIT('h80)
	) name22640 (
		\m2_addr_i[10]_pad ,
		_w8743_,
		_w8744_,
		_w24541_
	);
	LUT4 #(
		.INIT('habef)
	) name22641 (
		_w8738_,
		_w8741_,
		_w24540_,
		_w24541_,
		_w24542_
	);
	LUT3 #(
		.INIT('h2a)
	) name22642 (
		\m5_addr_i[10]_pad ,
		_w8743_,
		_w8744_,
		_w24543_
	);
	LUT3 #(
		.INIT('h2a)
	) name22643 (
		\m1_addr_i[10]_pad ,
		_w8743_,
		_w8744_,
		_w24544_
	);
	LUT4 #(
		.INIT('h57df)
	) name22644 (
		_w8738_,
		_w8741_,
		_w24543_,
		_w24544_,
		_w24545_
	);
	LUT3 #(
		.INIT('h80)
	) name22645 (
		\m0_addr_i[10]_pad ,
		_w8743_,
		_w8744_,
		_w24546_
	);
	LUT3 #(
		.INIT('h2a)
	) name22646 (
		\m7_addr_i[10]_pad ,
		_w8743_,
		_w8744_,
		_w24547_
	);
	LUT4 #(
		.INIT('h6e7f)
	) name22647 (
		_w8738_,
		_w8741_,
		_w24546_,
		_w24547_,
		_w24548_
	);
	LUT4 #(
		.INIT('h7fff)
	) name22648 (
		_w24539_,
		_w24542_,
		_w24545_,
		_w24548_,
		_w24549_
	);
	LUT3 #(
		.INIT('h2a)
	) name22649 (
		\m3_addr_i[11]_pad ,
		_w8743_,
		_w8744_,
		_w24550_
	);
	LUT3 #(
		.INIT('h80)
	) name22650 (
		\m4_addr_i[11]_pad ,
		_w8743_,
		_w8744_,
		_w24551_
	);
	LUT4 #(
		.INIT('h9dbf)
	) name22651 (
		_w8738_,
		_w8741_,
		_w24550_,
		_w24551_,
		_w24552_
	);
	LUT3 #(
		.INIT('h80)
	) name22652 (
		\m6_addr_i[11]_pad ,
		_w8743_,
		_w8744_,
		_w24553_
	);
	LUT3 #(
		.INIT('h80)
	) name22653 (
		\m2_addr_i[11]_pad ,
		_w8743_,
		_w8744_,
		_w24554_
	);
	LUT4 #(
		.INIT('habef)
	) name22654 (
		_w8738_,
		_w8741_,
		_w24553_,
		_w24554_,
		_w24555_
	);
	LUT3 #(
		.INIT('h2a)
	) name22655 (
		\m5_addr_i[11]_pad ,
		_w8743_,
		_w8744_,
		_w24556_
	);
	LUT3 #(
		.INIT('h2a)
	) name22656 (
		\m1_addr_i[11]_pad ,
		_w8743_,
		_w8744_,
		_w24557_
	);
	LUT4 #(
		.INIT('h57df)
	) name22657 (
		_w8738_,
		_w8741_,
		_w24556_,
		_w24557_,
		_w24558_
	);
	LUT3 #(
		.INIT('h80)
	) name22658 (
		\m0_addr_i[11]_pad ,
		_w8743_,
		_w8744_,
		_w24559_
	);
	LUT3 #(
		.INIT('h2a)
	) name22659 (
		\m7_addr_i[11]_pad ,
		_w8743_,
		_w8744_,
		_w24560_
	);
	LUT4 #(
		.INIT('h6e7f)
	) name22660 (
		_w8738_,
		_w8741_,
		_w24559_,
		_w24560_,
		_w24561_
	);
	LUT4 #(
		.INIT('h7fff)
	) name22661 (
		_w24552_,
		_w24555_,
		_w24558_,
		_w24561_,
		_w24562_
	);
	LUT3 #(
		.INIT('h2a)
	) name22662 (
		\m3_addr_i[12]_pad ,
		_w8743_,
		_w8744_,
		_w24563_
	);
	LUT3 #(
		.INIT('h80)
	) name22663 (
		\m4_addr_i[12]_pad ,
		_w8743_,
		_w8744_,
		_w24564_
	);
	LUT4 #(
		.INIT('h9dbf)
	) name22664 (
		_w8738_,
		_w8741_,
		_w24563_,
		_w24564_,
		_w24565_
	);
	LUT3 #(
		.INIT('h80)
	) name22665 (
		\m6_addr_i[12]_pad ,
		_w8743_,
		_w8744_,
		_w24566_
	);
	LUT3 #(
		.INIT('h2a)
	) name22666 (
		\m7_addr_i[12]_pad ,
		_w8743_,
		_w8744_,
		_w24567_
	);
	LUT3 #(
		.INIT('h57)
	) name22667 (
		_w8756_,
		_w24566_,
		_w24567_,
		_w24568_
	);
	LUT3 #(
		.INIT('h2a)
	) name22668 (
		\m5_addr_i[12]_pad ,
		_w8743_,
		_w8744_,
		_w24569_
	);
	LUT3 #(
		.INIT('h80)
	) name22669 (
		\m0_addr_i[12]_pad ,
		_w8743_,
		_w8744_,
		_w24570_
	);
	LUT4 #(
		.INIT('h57df)
	) name22670 (
		_w8738_,
		_w8741_,
		_w24569_,
		_w24570_,
		_w24571_
	);
	LUT3 #(
		.INIT('h2a)
	) name22671 (
		\m1_addr_i[12]_pad ,
		_w8743_,
		_w8744_,
		_w24572_
	);
	LUT3 #(
		.INIT('h80)
	) name22672 (
		\m2_addr_i[12]_pad ,
		_w8743_,
		_w8744_,
		_w24573_
	);
	LUT4 #(
		.INIT('h3b7f)
	) name22673 (
		_w8738_,
		_w8741_,
		_w24572_,
		_w24573_,
		_w24574_
	);
	LUT4 #(
		.INIT('h7fff)
	) name22674 (
		_w24565_,
		_w24568_,
		_w24571_,
		_w24574_,
		_w24575_
	);
	LUT3 #(
		.INIT('h2a)
	) name22675 (
		\m3_addr_i[13]_pad ,
		_w8743_,
		_w8744_,
		_w24576_
	);
	LUT3 #(
		.INIT('h80)
	) name22676 (
		\m4_addr_i[13]_pad ,
		_w8743_,
		_w8744_,
		_w24577_
	);
	LUT4 #(
		.INIT('h9dbf)
	) name22677 (
		_w8738_,
		_w8741_,
		_w24576_,
		_w24577_,
		_w24578_
	);
	LUT3 #(
		.INIT('h80)
	) name22678 (
		\m6_addr_i[13]_pad ,
		_w8743_,
		_w8744_,
		_w24579_
	);
	LUT3 #(
		.INIT('h80)
	) name22679 (
		\m2_addr_i[13]_pad ,
		_w8743_,
		_w8744_,
		_w24580_
	);
	LUT4 #(
		.INIT('habef)
	) name22680 (
		_w8738_,
		_w8741_,
		_w24579_,
		_w24580_,
		_w24581_
	);
	LUT3 #(
		.INIT('h2a)
	) name22681 (
		\m5_addr_i[13]_pad ,
		_w8743_,
		_w8744_,
		_w24582_
	);
	LUT3 #(
		.INIT('h2a)
	) name22682 (
		\m1_addr_i[13]_pad ,
		_w8743_,
		_w8744_,
		_w24583_
	);
	LUT4 #(
		.INIT('h57df)
	) name22683 (
		_w8738_,
		_w8741_,
		_w24582_,
		_w24583_,
		_w24584_
	);
	LUT3 #(
		.INIT('h80)
	) name22684 (
		\m0_addr_i[13]_pad ,
		_w8743_,
		_w8744_,
		_w24585_
	);
	LUT3 #(
		.INIT('h2a)
	) name22685 (
		\m7_addr_i[13]_pad ,
		_w8743_,
		_w8744_,
		_w24586_
	);
	LUT4 #(
		.INIT('h6e7f)
	) name22686 (
		_w8738_,
		_w8741_,
		_w24585_,
		_w24586_,
		_w24587_
	);
	LUT4 #(
		.INIT('h7fff)
	) name22687 (
		_w24578_,
		_w24581_,
		_w24584_,
		_w24587_,
		_w24588_
	);
	LUT3 #(
		.INIT('h2a)
	) name22688 (
		\m3_addr_i[14]_pad ,
		_w8743_,
		_w8744_,
		_w24589_
	);
	LUT3 #(
		.INIT('h80)
	) name22689 (
		\m4_addr_i[14]_pad ,
		_w8743_,
		_w8744_,
		_w24590_
	);
	LUT4 #(
		.INIT('h9dbf)
	) name22690 (
		_w8738_,
		_w8741_,
		_w24589_,
		_w24590_,
		_w24591_
	);
	LUT3 #(
		.INIT('h80)
	) name22691 (
		\m6_addr_i[14]_pad ,
		_w8743_,
		_w8744_,
		_w24592_
	);
	LUT3 #(
		.INIT('h80)
	) name22692 (
		\m2_addr_i[14]_pad ,
		_w8743_,
		_w8744_,
		_w24593_
	);
	LUT4 #(
		.INIT('habef)
	) name22693 (
		_w8738_,
		_w8741_,
		_w24592_,
		_w24593_,
		_w24594_
	);
	LUT3 #(
		.INIT('h2a)
	) name22694 (
		\m5_addr_i[14]_pad ,
		_w8743_,
		_w8744_,
		_w24595_
	);
	LUT3 #(
		.INIT('h2a)
	) name22695 (
		\m1_addr_i[14]_pad ,
		_w8743_,
		_w8744_,
		_w24596_
	);
	LUT4 #(
		.INIT('h57df)
	) name22696 (
		_w8738_,
		_w8741_,
		_w24595_,
		_w24596_,
		_w24597_
	);
	LUT3 #(
		.INIT('h80)
	) name22697 (
		\m0_addr_i[14]_pad ,
		_w8743_,
		_w8744_,
		_w24598_
	);
	LUT3 #(
		.INIT('h2a)
	) name22698 (
		\m7_addr_i[14]_pad ,
		_w8743_,
		_w8744_,
		_w24599_
	);
	LUT4 #(
		.INIT('h6e7f)
	) name22699 (
		_w8738_,
		_w8741_,
		_w24598_,
		_w24599_,
		_w24600_
	);
	LUT4 #(
		.INIT('h7fff)
	) name22700 (
		_w24591_,
		_w24594_,
		_w24597_,
		_w24600_,
		_w24601_
	);
	LUT3 #(
		.INIT('h2a)
	) name22701 (
		\m1_addr_i[15]_pad ,
		_w8743_,
		_w8744_,
		_w24602_
	);
	LUT3 #(
		.INIT('h80)
	) name22702 (
		\m2_addr_i[15]_pad ,
		_w8743_,
		_w8744_,
		_w24603_
	);
	LUT4 #(
		.INIT('h3b7f)
	) name22703 (
		_w8738_,
		_w8741_,
		_w24602_,
		_w24603_,
		_w24604_
	);
	LUT3 #(
		.INIT('h2a)
	) name22704 (
		\m3_addr_i[15]_pad ,
		_w8743_,
		_w8744_,
		_w24605_
	);
	LUT3 #(
		.INIT('h2a)
	) name22705 (
		\m7_addr_i[15]_pad ,
		_w8743_,
		_w8744_,
		_w24606_
	);
	LUT4 #(
		.INIT('haebf)
	) name22706 (
		_w8738_,
		_w8741_,
		_w24605_,
		_w24606_,
		_w24607_
	);
	LUT3 #(
		.INIT('h80)
	) name22707 (
		\m4_addr_i[15]_pad ,
		_w8743_,
		_w8744_,
		_w24608_
	);
	LUT3 #(
		.INIT('h80)
	) name22708 (
		\m0_addr_i[15]_pad ,
		_w8743_,
		_w8744_,
		_w24609_
	);
	LUT4 #(
		.INIT('h57df)
	) name22709 (
		_w8738_,
		_w8741_,
		_w24608_,
		_w24609_,
		_w24610_
	);
	LUT3 #(
		.INIT('h80)
	) name22710 (
		\m6_addr_i[15]_pad ,
		_w8743_,
		_w8744_,
		_w24611_
	);
	LUT3 #(
		.INIT('h2a)
	) name22711 (
		\m5_addr_i[15]_pad ,
		_w8743_,
		_w8744_,
		_w24612_
	);
	LUT4 #(
		.INIT('hcdef)
	) name22712 (
		_w8738_,
		_w8741_,
		_w24611_,
		_w24612_,
		_w24613_
	);
	LUT4 #(
		.INIT('h7fff)
	) name22713 (
		_w24604_,
		_w24607_,
		_w24610_,
		_w24613_,
		_w24614_
	);
	LUT3 #(
		.INIT('h2a)
	) name22714 (
		\m3_addr_i[16]_pad ,
		_w8743_,
		_w8744_,
		_w24615_
	);
	LUT3 #(
		.INIT('h80)
	) name22715 (
		\m4_addr_i[16]_pad ,
		_w8743_,
		_w8744_,
		_w24616_
	);
	LUT4 #(
		.INIT('h9dbf)
	) name22716 (
		_w8738_,
		_w8741_,
		_w24615_,
		_w24616_,
		_w24617_
	);
	LUT3 #(
		.INIT('h80)
	) name22717 (
		\m6_addr_i[16]_pad ,
		_w8743_,
		_w8744_,
		_w24618_
	);
	LUT3 #(
		.INIT('h80)
	) name22718 (
		\m2_addr_i[16]_pad ,
		_w8743_,
		_w8744_,
		_w24619_
	);
	LUT4 #(
		.INIT('habef)
	) name22719 (
		_w8738_,
		_w8741_,
		_w24618_,
		_w24619_,
		_w24620_
	);
	LUT3 #(
		.INIT('h2a)
	) name22720 (
		\m5_addr_i[16]_pad ,
		_w8743_,
		_w8744_,
		_w24621_
	);
	LUT3 #(
		.INIT('h2a)
	) name22721 (
		\m1_addr_i[16]_pad ,
		_w8743_,
		_w8744_,
		_w24622_
	);
	LUT4 #(
		.INIT('h57df)
	) name22722 (
		_w8738_,
		_w8741_,
		_w24621_,
		_w24622_,
		_w24623_
	);
	LUT3 #(
		.INIT('h80)
	) name22723 (
		\m0_addr_i[16]_pad ,
		_w8743_,
		_w8744_,
		_w24624_
	);
	LUT3 #(
		.INIT('h2a)
	) name22724 (
		\m7_addr_i[16]_pad ,
		_w8743_,
		_w8744_,
		_w24625_
	);
	LUT4 #(
		.INIT('h6e7f)
	) name22725 (
		_w8738_,
		_w8741_,
		_w24624_,
		_w24625_,
		_w24626_
	);
	LUT4 #(
		.INIT('h7fff)
	) name22726 (
		_w24617_,
		_w24620_,
		_w24623_,
		_w24626_,
		_w24627_
	);
	LUT3 #(
		.INIT('h2a)
	) name22727 (
		\m3_addr_i[17]_pad ,
		_w8743_,
		_w8744_,
		_w24628_
	);
	LUT3 #(
		.INIT('h80)
	) name22728 (
		\m4_addr_i[17]_pad ,
		_w8743_,
		_w8744_,
		_w24629_
	);
	LUT4 #(
		.INIT('h9dbf)
	) name22729 (
		_w8738_,
		_w8741_,
		_w24628_,
		_w24629_,
		_w24630_
	);
	LUT3 #(
		.INIT('h80)
	) name22730 (
		\m6_addr_i[17]_pad ,
		_w8743_,
		_w8744_,
		_w24631_
	);
	LUT3 #(
		.INIT('h80)
	) name22731 (
		\m2_addr_i[17]_pad ,
		_w8743_,
		_w8744_,
		_w24632_
	);
	LUT4 #(
		.INIT('habef)
	) name22732 (
		_w8738_,
		_w8741_,
		_w24631_,
		_w24632_,
		_w24633_
	);
	LUT3 #(
		.INIT('h2a)
	) name22733 (
		\m5_addr_i[17]_pad ,
		_w8743_,
		_w8744_,
		_w24634_
	);
	LUT3 #(
		.INIT('h2a)
	) name22734 (
		\m1_addr_i[17]_pad ,
		_w8743_,
		_w8744_,
		_w24635_
	);
	LUT4 #(
		.INIT('h57df)
	) name22735 (
		_w8738_,
		_w8741_,
		_w24634_,
		_w24635_,
		_w24636_
	);
	LUT3 #(
		.INIT('h80)
	) name22736 (
		\m0_addr_i[17]_pad ,
		_w8743_,
		_w8744_,
		_w24637_
	);
	LUT3 #(
		.INIT('h2a)
	) name22737 (
		\m7_addr_i[17]_pad ,
		_w8743_,
		_w8744_,
		_w24638_
	);
	LUT4 #(
		.INIT('h6e7f)
	) name22738 (
		_w8738_,
		_w8741_,
		_w24637_,
		_w24638_,
		_w24639_
	);
	LUT4 #(
		.INIT('h7fff)
	) name22739 (
		_w24630_,
		_w24633_,
		_w24636_,
		_w24639_,
		_w24640_
	);
	LUT3 #(
		.INIT('h2a)
	) name22740 (
		\m3_addr_i[18]_pad ,
		_w8743_,
		_w8744_,
		_w24641_
	);
	LUT3 #(
		.INIT('h80)
	) name22741 (
		\m4_addr_i[18]_pad ,
		_w8743_,
		_w8744_,
		_w24642_
	);
	LUT4 #(
		.INIT('h9dbf)
	) name22742 (
		_w8738_,
		_w8741_,
		_w24641_,
		_w24642_,
		_w24643_
	);
	LUT3 #(
		.INIT('h80)
	) name22743 (
		\m6_addr_i[18]_pad ,
		_w8743_,
		_w8744_,
		_w24644_
	);
	LUT3 #(
		.INIT('h80)
	) name22744 (
		\m2_addr_i[18]_pad ,
		_w8743_,
		_w8744_,
		_w24645_
	);
	LUT4 #(
		.INIT('habef)
	) name22745 (
		_w8738_,
		_w8741_,
		_w24644_,
		_w24645_,
		_w24646_
	);
	LUT3 #(
		.INIT('h2a)
	) name22746 (
		\m5_addr_i[18]_pad ,
		_w8743_,
		_w8744_,
		_w24647_
	);
	LUT3 #(
		.INIT('h2a)
	) name22747 (
		\m1_addr_i[18]_pad ,
		_w8743_,
		_w8744_,
		_w24648_
	);
	LUT4 #(
		.INIT('h57df)
	) name22748 (
		_w8738_,
		_w8741_,
		_w24647_,
		_w24648_,
		_w24649_
	);
	LUT3 #(
		.INIT('h80)
	) name22749 (
		\m0_addr_i[18]_pad ,
		_w8743_,
		_w8744_,
		_w24650_
	);
	LUT3 #(
		.INIT('h2a)
	) name22750 (
		\m7_addr_i[18]_pad ,
		_w8743_,
		_w8744_,
		_w24651_
	);
	LUT4 #(
		.INIT('h6e7f)
	) name22751 (
		_w8738_,
		_w8741_,
		_w24650_,
		_w24651_,
		_w24652_
	);
	LUT4 #(
		.INIT('h7fff)
	) name22752 (
		_w24643_,
		_w24646_,
		_w24649_,
		_w24652_,
		_w24653_
	);
	LUT3 #(
		.INIT('h2a)
	) name22753 (
		\m3_addr_i[19]_pad ,
		_w8743_,
		_w8744_,
		_w24654_
	);
	LUT3 #(
		.INIT('h80)
	) name22754 (
		\m4_addr_i[19]_pad ,
		_w8743_,
		_w8744_,
		_w24655_
	);
	LUT4 #(
		.INIT('h9dbf)
	) name22755 (
		_w8738_,
		_w8741_,
		_w24654_,
		_w24655_,
		_w24656_
	);
	LUT3 #(
		.INIT('h80)
	) name22756 (
		\m6_addr_i[19]_pad ,
		_w8743_,
		_w8744_,
		_w24657_
	);
	LUT3 #(
		.INIT('h80)
	) name22757 (
		\m2_addr_i[19]_pad ,
		_w8743_,
		_w8744_,
		_w24658_
	);
	LUT4 #(
		.INIT('habef)
	) name22758 (
		_w8738_,
		_w8741_,
		_w24657_,
		_w24658_,
		_w24659_
	);
	LUT3 #(
		.INIT('h2a)
	) name22759 (
		\m5_addr_i[19]_pad ,
		_w8743_,
		_w8744_,
		_w24660_
	);
	LUT3 #(
		.INIT('h2a)
	) name22760 (
		\m1_addr_i[19]_pad ,
		_w8743_,
		_w8744_,
		_w24661_
	);
	LUT4 #(
		.INIT('h57df)
	) name22761 (
		_w8738_,
		_w8741_,
		_w24660_,
		_w24661_,
		_w24662_
	);
	LUT3 #(
		.INIT('h80)
	) name22762 (
		\m0_addr_i[19]_pad ,
		_w8743_,
		_w8744_,
		_w24663_
	);
	LUT3 #(
		.INIT('h2a)
	) name22763 (
		\m7_addr_i[19]_pad ,
		_w8743_,
		_w8744_,
		_w24664_
	);
	LUT4 #(
		.INIT('h6e7f)
	) name22764 (
		_w8738_,
		_w8741_,
		_w24663_,
		_w24664_,
		_w24665_
	);
	LUT4 #(
		.INIT('h7fff)
	) name22765 (
		_w24656_,
		_w24659_,
		_w24662_,
		_w24665_,
		_w24666_
	);
	LUT3 #(
		.INIT('h2a)
	) name22766 (
		\m3_addr_i[1]_pad ,
		_w8743_,
		_w8744_,
		_w24667_
	);
	LUT3 #(
		.INIT('h80)
	) name22767 (
		\m4_addr_i[1]_pad ,
		_w8743_,
		_w8744_,
		_w24668_
	);
	LUT4 #(
		.INIT('h9dbf)
	) name22768 (
		_w8738_,
		_w8741_,
		_w24667_,
		_w24668_,
		_w24669_
	);
	LUT3 #(
		.INIT('h80)
	) name22769 (
		\m6_addr_i[1]_pad ,
		_w8743_,
		_w8744_,
		_w24670_
	);
	LUT3 #(
		.INIT('h2a)
	) name22770 (
		\m7_addr_i[1]_pad ,
		_w8743_,
		_w8744_,
		_w24671_
	);
	LUT3 #(
		.INIT('h57)
	) name22771 (
		_w8756_,
		_w24670_,
		_w24671_,
		_w24672_
	);
	LUT3 #(
		.INIT('h2a)
	) name22772 (
		\m5_addr_i[1]_pad ,
		_w8743_,
		_w8744_,
		_w24673_
	);
	LUT3 #(
		.INIT('h80)
	) name22773 (
		\m0_addr_i[1]_pad ,
		_w8743_,
		_w8744_,
		_w24674_
	);
	LUT4 #(
		.INIT('h57df)
	) name22774 (
		_w8738_,
		_w8741_,
		_w24673_,
		_w24674_,
		_w24675_
	);
	LUT3 #(
		.INIT('h2a)
	) name22775 (
		\m1_addr_i[1]_pad ,
		_w8743_,
		_w8744_,
		_w24676_
	);
	LUT3 #(
		.INIT('h80)
	) name22776 (
		\m2_addr_i[1]_pad ,
		_w8743_,
		_w8744_,
		_w24677_
	);
	LUT4 #(
		.INIT('h3b7f)
	) name22777 (
		_w8738_,
		_w8741_,
		_w24676_,
		_w24677_,
		_w24678_
	);
	LUT4 #(
		.INIT('h7fff)
	) name22778 (
		_w24669_,
		_w24672_,
		_w24675_,
		_w24678_,
		_w24679_
	);
	LUT3 #(
		.INIT('h2a)
	) name22779 (
		\m3_addr_i[20]_pad ,
		_w8743_,
		_w8744_,
		_w24680_
	);
	LUT3 #(
		.INIT('h80)
	) name22780 (
		\m4_addr_i[20]_pad ,
		_w8743_,
		_w8744_,
		_w24681_
	);
	LUT4 #(
		.INIT('h9dbf)
	) name22781 (
		_w8738_,
		_w8741_,
		_w24680_,
		_w24681_,
		_w24682_
	);
	LUT3 #(
		.INIT('h80)
	) name22782 (
		\m6_addr_i[20]_pad ,
		_w8743_,
		_w8744_,
		_w24683_
	);
	LUT3 #(
		.INIT('h80)
	) name22783 (
		\m2_addr_i[20]_pad ,
		_w8743_,
		_w8744_,
		_w24684_
	);
	LUT4 #(
		.INIT('habef)
	) name22784 (
		_w8738_,
		_w8741_,
		_w24683_,
		_w24684_,
		_w24685_
	);
	LUT3 #(
		.INIT('h2a)
	) name22785 (
		\m5_addr_i[20]_pad ,
		_w8743_,
		_w8744_,
		_w24686_
	);
	LUT3 #(
		.INIT('h2a)
	) name22786 (
		\m1_addr_i[20]_pad ,
		_w8743_,
		_w8744_,
		_w24687_
	);
	LUT4 #(
		.INIT('h57df)
	) name22787 (
		_w8738_,
		_w8741_,
		_w24686_,
		_w24687_,
		_w24688_
	);
	LUT3 #(
		.INIT('h80)
	) name22788 (
		\m0_addr_i[20]_pad ,
		_w8743_,
		_w8744_,
		_w24689_
	);
	LUT3 #(
		.INIT('h2a)
	) name22789 (
		\m7_addr_i[20]_pad ,
		_w8743_,
		_w8744_,
		_w24690_
	);
	LUT4 #(
		.INIT('h6e7f)
	) name22790 (
		_w8738_,
		_w8741_,
		_w24689_,
		_w24690_,
		_w24691_
	);
	LUT4 #(
		.INIT('h7fff)
	) name22791 (
		_w24682_,
		_w24685_,
		_w24688_,
		_w24691_,
		_w24692_
	);
	LUT3 #(
		.INIT('h2a)
	) name22792 (
		\m3_addr_i[21]_pad ,
		_w8743_,
		_w8744_,
		_w24693_
	);
	LUT3 #(
		.INIT('h80)
	) name22793 (
		\m4_addr_i[21]_pad ,
		_w8743_,
		_w8744_,
		_w24694_
	);
	LUT4 #(
		.INIT('h9dbf)
	) name22794 (
		_w8738_,
		_w8741_,
		_w24693_,
		_w24694_,
		_w24695_
	);
	LUT3 #(
		.INIT('h80)
	) name22795 (
		\m6_addr_i[21]_pad ,
		_w8743_,
		_w8744_,
		_w24696_
	);
	LUT3 #(
		.INIT('h80)
	) name22796 (
		\m2_addr_i[21]_pad ,
		_w8743_,
		_w8744_,
		_w24697_
	);
	LUT4 #(
		.INIT('habef)
	) name22797 (
		_w8738_,
		_w8741_,
		_w24696_,
		_w24697_,
		_w24698_
	);
	LUT3 #(
		.INIT('h2a)
	) name22798 (
		\m5_addr_i[21]_pad ,
		_w8743_,
		_w8744_,
		_w24699_
	);
	LUT3 #(
		.INIT('h2a)
	) name22799 (
		\m1_addr_i[21]_pad ,
		_w8743_,
		_w8744_,
		_w24700_
	);
	LUT4 #(
		.INIT('h57df)
	) name22800 (
		_w8738_,
		_w8741_,
		_w24699_,
		_w24700_,
		_w24701_
	);
	LUT3 #(
		.INIT('h80)
	) name22801 (
		\m0_addr_i[21]_pad ,
		_w8743_,
		_w8744_,
		_w24702_
	);
	LUT3 #(
		.INIT('h2a)
	) name22802 (
		\m7_addr_i[21]_pad ,
		_w8743_,
		_w8744_,
		_w24703_
	);
	LUT4 #(
		.INIT('h6e7f)
	) name22803 (
		_w8738_,
		_w8741_,
		_w24702_,
		_w24703_,
		_w24704_
	);
	LUT4 #(
		.INIT('h7fff)
	) name22804 (
		_w24695_,
		_w24698_,
		_w24701_,
		_w24704_,
		_w24705_
	);
	LUT3 #(
		.INIT('h2a)
	) name22805 (
		\m1_addr_i[22]_pad ,
		_w8743_,
		_w8744_,
		_w24706_
	);
	LUT3 #(
		.INIT('h80)
	) name22806 (
		\m2_addr_i[22]_pad ,
		_w8743_,
		_w8744_,
		_w24707_
	);
	LUT4 #(
		.INIT('h3b7f)
	) name22807 (
		_w8738_,
		_w8741_,
		_w24706_,
		_w24707_,
		_w24708_
	);
	LUT3 #(
		.INIT('h2a)
	) name22808 (
		\m3_addr_i[22]_pad ,
		_w8743_,
		_w8744_,
		_w24709_
	);
	LUT3 #(
		.INIT('h2a)
	) name22809 (
		\m5_addr_i[22]_pad ,
		_w8743_,
		_w8744_,
		_w24710_
	);
	LUT4 #(
		.INIT('h9dbf)
	) name22810 (
		_w8738_,
		_w8741_,
		_w24709_,
		_w24710_,
		_w24711_
	);
	LUT3 #(
		.INIT('h80)
	) name22811 (
		\m4_addr_i[22]_pad ,
		_w8743_,
		_w8744_,
		_w24712_
	);
	LUT3 #(
		.INIT('h80)
	) name22812 (
		\m6_addr_i[22]_pad ,
		_w8743_,
		_w8744_,
		_w24713_
	);
	LUT4 #(
		.INIT('hcedf)
	) name22813 (
		_w8738_,
		_w8741_,
		_w24712_,
		_w24713_,
		_w24714_
	);
	LUT3 #(
		.INIT('h80)
	) name22814 (
		\m0_addr_i[22]_pad ,
		_w8743_,
		_w8744_,
		_w24715_
	);
	LUT3 #(
		.INIT('h2a)
	) name22815 (
		\m7_addr_i[22]_pad ,
		_w8743_,
		_w8744_,
		_w24716_
	);
	LUT4 #(
		.INIT('h6e7f)
	) name22816 (
		_w8738_,
		_w8741_,
		_w24715_,
		_w24716_,
		_w24717_
	);
	LUT4 #(
		.INIT('h7fff)
	) name22817 (
		_w24708_,
		_w24711_,
		_w24714_,
		_w24717_,
		_w24718_
	);
	LUT3 #(
		.INIT('h2a)
	) name22818 (
		\m3_addr_i[23]_pad ,
		_w8743_,
		_w8744_,
		_w24719_
	);
	LUT3 #(
		.INIT('h80)
	) name22819 (
		\m4_addr_i[23]_pad ,
		_w8743_,
		_w8744_,
		_w24720_
	);
	LUT4 #(
		.INIT('h9dbf)
	) name22820 (
		_w8738_,
		_w8741_,
		_w24719_,
		_w24720_,
		_w24721_
	);
	LUT3 #(
		.INIT('h2a)
	) name22821 (
		\m1_addr_i[23]_pad ,
		_w8743_,
		_w8744_,
		_w24722_
	);
	LUT3 #(
		.INIT('h2a)
	) name22822 (
		\m5_addr_i[23]_pad ,
		_w8743_,
		_w8744_,
		_w24723_
	);
	LUT4 #(
		.INIT('h5d7f)
	) name22823 (
		_w8738_,
		_w8741_,
		_w24722_,
		_w24723_,
		_w24724_
	);
	LUT3 #(
		.INIT('h80)
	) name22824 (
		\m2_addr_i[23]_pad ,
		_w8743_,
		_w8744_,
		_w24725_
	);
	LUT3 #(
		.INIT('h80)
	) name22825 (
		\m6_addr_i[23]_pad ,
		_w8743_,
		_w8744_,
		_w24726_
	);
	LUT4 #(
		.INIT('haebf)
	) name22826 (
		_w8738_,
		_w8741_,
		_w24725_,
		_w24726_,
		_w24727_
	);
	LUT3 #(
		.INIT('h80)
	) name22827 (
		\m0_addr_i[23]_pad ,
		_w8743_,
		_w8744_,
		_w24728_
	);
	LUT3 #(
		.INIT('h2a)
	) name22828 (
		\m7_addr_i[23]_pad ,
		_w8743_,
		_w8744_,
		_w24729_
	);
	LUT4 #(
		.INIT('h6e7f)
	) name22829 (
		_w8738_,
		_w8741_,
		_w24728_,
		_w24729_,
		_w24730_
	);
	LUT4 #(
		.INIT('h7fff)
	) name22830 (
		_w24721_,
		_w24724_,
		_w24727_,
		_w24730_,
		_w24731_
	);
	LUT3 #(
		.INIT('h2a)
	) name22831 (
		\m1_addr_i[24]_pad ,
		_w8743_,
		_w8744_,
		_w24732_
	);
	LUT3 #(
		.INIT('h80)
	) name22832 (
		\m2_addr_i[24]_pad ,
		_w8743_,
		_w8744_,
		_w24733_
	);
	LUT4 #(
		.INIT('h3b7f)
	) name22833 (
		_w8738_,
		_w8741_,
		_w24732_,
		_w24733_,
		_w24734_
	);
	LUT3 #(
		.INIT('h2a)
	) name22834 (
		\m3_addr_i[24]_pad ,
		_w8743_,
		_w8744_,
		_w24735_
	);
	LUT3 #(
		.INIT('h2a)
	) name22835 (
		\m7_addr_i[24]_pad ,
		_w8743_,
		_w8744_,
		_w24736_
	);
	LUT4 #(
		.INIT('haebf)
	) name22836 (
		_w8738_,
		_w8741_,
		_w24735_,
		_w24736_,
		_w24737_
	);
	LUT3 #(
		.INIT('h80)
	) name22837 (
		\m4_addr_i[24]_pad ,
		_w8743_,
		_w8744_,
		_w24738_
	);
	LUT3 #(
		.INIT('h80)
	) name22838 (
		\m0_addr_i[24]_pad ,
		_w8743_,
		_w8744_,
		_w24739_
	);
	LUT4 #(
		.INIT('h57df)
	) name22839 (
		_w8738_,
		_w8741_,
		_w24738_,
		_w24739_,
		_w24740_
	);
	LUT3 #(
		.INIT('h2a)
	) name22840 (
		\m5_addr_i[24]_pad ,
		_w8743_,
		_w8744_,
		_w24741_
	);
	LUT3 #(
		.INIT('h80)
	) name22841 (
		\m6_addr_i[24]_pad ,
		_w8743_,
		_w8744_,
		_w24742_
	);
	LUT4 #(
		.INIT('hcedf)
	) name22842 (
		_w8738_,
		_w8741_,
		_w24741_,
		_w24742_,
		_w24743_
	);
	LUT4 #(
		.INIT('h7fff)
	) name22843 (
		_w24734_,
		_w24737_,
		_w24740_,
		_w24743_,
		_w24744_
	);
	LUT3 #(
		.INIT('h2a)
	) name22844 (
		\m3_addr_i[25]_pad ,
		_w8743_,
		_w8744_,
		_w24745_
	);
	LUT3 #(
		.INIT('h80)
	) name22845 (
		\m4_addr_i[25]_pad ,
		_w8743_,
		_w8744_,
		_w24746_
	);
	LUT4 #(
		.INIT('h9dbf)
	) name22846 (
		_w8738_,
		_w8741_,
		_w24745_,
		_w24746_,
		_w24747_
	);
	LUT3 #(
		.INIT('h80)
	) name22847 (
		\m0_addr_i[25]_pad ,
		_w8743_,
		_w8744_,
		_w24748_
	);
	LUT3 #(
		.INIT('h80)
	) name22848 (
		\m2_addr_i[25]_pad ,
		_w8743_,
		_w8744_,
		_w24749_
	);
	LUT4 #(
		.INIT('h3b7f)
	) name22849 (
		_w8738_,
		_w8741_,
		_w24748_,
		_w24749_,
		_w24750_
	);
	LUT3 #(
		.INIT('h2a)
	) name22850 (
		\m7_addr_i[25]_pad ,
		_w8743_,
		_w8744_,
		_w24751_
	);
	LUT3 #(
		.INIT('h2a)
	) name22851 (
		\m1_addr_i[25]_pad ,
		_w8743_,
		_w8744_,
		_w24752_
	);
	LUT4 #(
		.INIT('h67ef)
	) name22852 (
		_w8738_,
		_w8741_,
		_w24751_,
		_w24752_,
		_w24753_
	);
	LUT3 #(
		.INIT('h2a)
	) name22853 (
		\m5_addr_i[25]_pad ,
		_w8743_,
		_w8744_,
		_w24754_
	);
	LUT3 #(
		.INIT('h80)
	) name22854 (
		\m6_addr_i[25]_pad ,
		_w8743_,
		_w8744_,
		_w24755_
	);
	LUT4 #(
		.INIT('hcedf)
	) name22855 (
		_w8738_,
		_w8741_,
		_w24754_,
		_w24755_,
		_w24756_
	);
	LUT4 #(
		.INIT('h7fff)
	) name22856 (
		_w24747_,
		_w24750_,
		_w24753_,
		_w24756_,
		_w24757_
	);
	LUT3 #(
		.INIT('h2a)
	) name22857 (
		\m1_addr_i[26]_pad ,
		_w8743_,
		_w8744_,
		_w24758_
	);
	LUT3 #(
		.INIT('h80)
	) name22858 (
		\m2_addr_i[26]_pad ,
		_w8743_,
		_w8744_,
		_w24759_
	);
	LUT4 #(
		.INIT('h3b7f)
	) name22859 (
		_w8738_,
		_w8741_,
		_w24758_,
		_w24759_,
		_w24760_
	);
	LUT3 #(
		.INIT('h80)
	) name22860 (
		\m0_addr_i[26]_pad ,
		_w8743_,
		_w8744_,
		_w24761_
	);
	LUT3 #(
		.INIT('h80)
	) name22861 (
		\m4_addr_i[26]_pad ,
		_w8743_,
		_w8744_,
		_w24762_
	);
	LUT4 #(
		.INIT('h5d7f)
	) name22862 (
		_w8738_,
		_w8741_,
		_w24761_,
		_w24762_,
		_w24763_
	);
	LUT3 #(
		.INIT('h2a)
	) name22863 (
		\m7_addr_i[26]_pad ,
		_w8743_,
		_w8744_,
		_w24764_
	);
	LUT3 #(
		.INIT('h2a)
	) name22864 (
		\m3_addr_i[26]_pad ,
		_w8743_,
		_w8744_,
		_w24765_
	);
	LUT4 #(
		.INIT('habef)
	) name22865 (
		_w8738_,
		_w8741_,
		_w24764_,
		_w24765_,
		_w24766_
	);
	LUT3 #(
		.INIT('h2a)
	) name22866 (
		\m5_addr_i[26]_pad ,
		_w8743_,
		_w8744_,
		_w24767_
	);
	LUT3 #(
		.INIT('h80)
	) name22867 (
		\m6_addr_i[26]_pad ,
		_w8743_,
		_w8744_,
		_w24768_
	);
	LUT4 #(
		.INIT('hcedf)
	) name22868 (
		_w8738_,
		_w8741_,
		_w24767_,
		_w24768_,
		_w24769_
	);
	LUT4 #(
		.INIT('h7fff)
	) name22869 (
		_w24760_,
		_w24763_,
		_w24766_,
		_w24769_,
		_w24770_
	);
	LUT3 #(
		.INIT('h2a)
	) name22870 (
		\m3_addr_i[27]_pad ,
		_w8743_,
		_w8744_,
		_w24771_
	);
	LUT3 #(
		.INIT('h80)
	) name22871 (
		\m4_addr_i[27]_pad ,
		_w8743_,
		_w8744_,
		_w24772_
	);
	LUT4 #(
		.INIT('h9dbf)
	) name22872 (
		_w8738_,
		_w8741_,
		_w24771_,
		_w24772_,
		_w24773_
	);
	LUT3 #(
		.INIT('h80)
	) name22873 (
		\m0_addr_i[27]_pad ,
		_w8743_,
		_w8744_,
		_w24774_
	);
	LUT3 #(
		.INIT('h80)
	) name22874 (
		\m6_addr_i[27]_pad ,
		_w8743_,
		_w8744_,
		_w24775_
	);
	LUT4 #(
		.INIT('h6e7f)
	) name22875 (
		_w8738_,
		_w8741_,
		_w24774_,
		_w24775_,
		_w24776_
	);
	LUT3 #(
		.INIT('h2a)
	) name22876 (
		\m7_addr_i[27]_pad ,
		_w8743_,
		_w8744_,
		_w24777_
	);
	LUT3 #(
		.INIT('h2a)
	) name22877 (
		\m5_addr_i[27]_pad ,
		_w8743_,
		_w8744_,
		_w24778_
	);
	LUT4 #(
		.INIT('hcdef)
	) name22878 (
		_w8738_,
		_w8741_,
		_w24777_,
		_w24778_,
		_w24779_
	);
	LUT3 #(
		.INIT('h2a)
	) name22879 (
		\m1_addr_i[27]_pad ,
		_w8743_,
		_w8744_,
		_w24780_
	);
	LUT3 #(
		.INIT('h80)
	) name22880 (
		\m2_addr_i[27]_pad ,
		_w8743_,
		_w8744_,
		_w24781_
	);
	LUT4 #(
		.INIT('h3b7f)
	) name22881 (
		_w8738_,
		_w8741_,
		_w24780_,
		_w24781_,
		_w24782_
	);
	LUT4 #(
		.INIT('h7fff)
	) name22882 (
		_w24773_,
		_w24776_,
		_w24779_,
		_w24782_,
		_w24783_
	);
	LUT3 #(
		.INIT('h2a)
	) name22883 (
		\m1_addr_i[28]_pad ,
		_w8743_,
		_w8744_,
		_w24784_
	);
	LUT3 #(
		.INIT('h80)
	) name22884 (
		\m2_addr_i[28]_pad ,
		_w8743_,
		_w8744_,
		_w24785_
	);
	LUT4 #(
		.INIT('h3b7f)
	) name22885 (
		_w8738_,
		_w8741_,
		_w24784_,
		_w24785_,
		_w24786_
	);
	LUT3 #(
		.INIT('h80)
	) name22886 (
		\m0_addr_i[28]_pad ,
		_w8743_,
		_w8744_,
		_w24787_
	);
	LUT3 #(
		.INIT('h80)
	) name22887 (
		\m6_addr_i[28]_pad ,
		_w8743_,
		_w8744_,
		_w24788_
	);
	LUT4 #(
		.INIT('h6e7f)
	) name22888 (
		_w8738_,
		_w8741_,
		_w24787_,
		_w24788_,
		_w24789_
	);
	LUT3 #(
		.INIT('h2a)
	) name22889 (
		\m7_addr_i[28]_pad ,
		_w8743_,
		_w8744_,
		_w24790_
	);
	LUT3 #(
		.INIT('h2a)
	) name22890 (
		\m5_addr_i[28]_pad ,
		_w8743_,
		_w8744_,
		_w24791_
	);
	LUT4 #(
		.INIT('hcdef)
	) name22891 (
		_w8738_,
		_w8741_,
		_w24790_,
		_w24791_,
		_w24792_
	);
	LUT3 #(
		.INIT('h2a)
	) name22892 (
		\m3_addr_i[28]_pad ,
		_w8743_,
		_w8744_,
		_w24793_
	);
	LUT3 #(
		.INIT('h80)
	) name22893 (
		\m4_addr_i[28]_pad ,
		_w8743_,
		_w8744_,
		_w24794_
	);
	LUT4 #(
		.INIT('h9dbf)
	) name22894 (
		_w8738_,
		_w8741_,
		_w24793_,
		_w24794_,
		_w24795_
	);
	LUT4 #(
		.INIT('h7fff)
	) name22895 (
		_w24786_,
		_w24789_,
		_w24792_,
		_w24795_,
		_w24796_
	);
	LUT3 #(
		.INIT('h80)
	) name22896 (
		\m0_addr_i[29]_pad ,
		_w8743_,
		_w8744_,
		_w24797_
	);
	LUT3 #(
		.INIT('h2a)
	) name22897 (
		\m7_addr_i[29]_pad ,
		_w8743_,
		_w8744_,
		_w24798_
	);
	LUT4 #(
		.INIT('h6e7f)
	) name22898 (
		_w8738_,
		_w8741_,
		_w24797_,
		_w24798_,
		_w24799_
	);
	LUT3 #(
		.INIT('h2a)
	) name22899 (
		\m5_addr_i[29]_pad ,
		_w8743_,
		_w8744_,
		_w24800_
	);
	LUT3 #(
		.INIT('h80)
	) name22900 (
		\m2_addr_i[29]_pad ,
		_w8743_,
		_w8744_,
		_w24801_
	);
	LUT4 #(
		.INIT('h9bdf)
	) name22901 (
		_w8738_,
		_w8741_,
		_w24800_,
		_w24801_,
		_w24802_
	);
	LUT3 #(
		.INIT('h80)
	) name22902 (
		\m6_addr_i[29]_pad ,
		_w8743_,
		_w8744_,
		_w24803_
	);
	LUT3 #(
		.INIT('h2a)
	) name22903 (
		\m1_addr_i[29]_pad ,
		_w8743_,
		_w8744_,
		_w24804_
	);
	LUT4 #(
		.INIT('h67ef)
	) name22904 (
		_w8738_,
		_w8741_,
		_w24803_,
		_w24804_,
		_w24805_
	);
	LUT3 #(
		.INIT('h2a)
	) name22905 (
		\m3_addr_i[29]_pad ,
		_w8743_,
		_w8744_,
		_w24806_
	);
	LUT3 #(
		.INIT('h80)
	) name22906 (
		\m4_addr_i[29]_pad ,
		_w8743_,
		_w8744_,
		_w24807_
	);
	LUT4 #(
		.INIT('h9dbf)
	) name22907 (
		_w8738_,
		_w8741_,
		_w24806_,
		_w24807_,
		_w24808_
	);
	LUT4 #(
		.INIT('h7fff)
	) name22908 (
		_w24799_,
		_w24802_,
		_w24805_,
		_w24808_,
		_w24809_
	);
	LUT3 #(
		.INIT('h2a)
	) name22909 (
		\m3_addr_i[2]_pad ,
		_w8743_,
		_w8744_,
		_w24810_
	);
	LUT3 #(
		.INIT('h80)
	) name22910 (
		\m4_addr_i[2]_pad ,
		_w8743_,
		_w8744_,
		_w24811_
	);
	LUT4 #(
		.INIT('h9dbf)
	) name22911 (
		_w8738_,
		_w8741_,
		_w24810_,
		_w24811_,
		_w24812_
	);
	LUT3 #(
		.INIT('h80)
	) name22912 (
		\m6_addr_i[2]_pad ,
		_w8743_,
		_w8744_,
		_w24813_
	);
	LUT3 #(
		.INIT('h80)
	) name22913 (
		\m2_addr_i[2]_pad ,
		_w8743_,
		_w8744_,
		_w24814_
	);
	LUT4 #(
		.INIT('habef)
	) name22914 (
		_w8738_,
		_w8741_,
		_w24813_,
		_w24814_,
		_w24815_
	);
	LUT3 #(
		.INIT('h2a)
	) name22915 (
		\m5_addr_i[2]_pad ,
		_w8743_,
		_w8744_,
		_w24816_
	);
	LUT3 #(
		.INIT('h2a)
	) name22916 (
		\m1_addr_i[2]_pad ,
		_w8743_,
		_w8744_,
		_w24817_
	);
	LUT4 #(
		.INIT('h57df)
	) name22917 (
		_w8738_,
		_w8741_,
		_w24816_,
		_w24817_,
		_w24818_
	);
	LUT3 #(
		.INIT('h80)
	) name22918 (
		\m0_addr_i[2]_pad ,
		_w8743_,
		_w8744_,
		_w24819_
	);
	LUT3 #(
		.INIT('h2a)
	) name22919 (
		\m7_addr_i[2]_pad ,
		_w8743_,
		_w8744_,
		_w24820_
	);
	LUT4 #(
		.INIT('h6e7f)
	) name22920 (
		_w8738_,
		_w8741_,
		_w24819_,
		_w24820_,
		_w24821_
	);
	LUT4 #(
		.INIT('h7fff)
	) name22921 (
		_w24812_,
		_w24815_,
		_w24818_,
		_w24821_,
		_w24822_
	);
	LUT3 #(
		.INIT('h2a)
	) name22922 (
		\m1_addr_i[30]_pad ,
		_w8743_,
		_w8744_,
		_w24823_
	);
	LUT3 #(
		.INIT('h80)
	) name22923 (
		\m2_addr_i[30]_pad ,
		_w8743_,
		_w8744_,
		_w24824_
	);
	LUT4 #(
		.INIT('h3b7f)
	) name22924 (
		_w8738_,
		_w8741_,
		_w24823_,
		_w24824_,
		_w24825_
	);
	LUT3 #(
		.INIT('h80)
	) name22925 (
		\m0_addr_i[30]_pad ,
		_w8743_,
		_w8744_,
		_w24826_
	);
	LUT3 #(
		.INIT('h80)
	) name22926 (
		\m4_addr_i[30]_pad ,
		_w8743_,
		_w8744_,
		_w24827_
	);
	LUT4 #(
		.INIT('h5d7f)
	) name22927 (
		_w8738_,
		_w8741_,
		_w24826_,
		_w24827_,
		_w24828_
	);
	LUT3 #(
		.INIT('h2a)
	) name22928 (
		\m7_addr_i[30]_pad ,
		_w8743_,
		_w8744_,
		_w24829_
	);
	LUT3 #(
		.INIT('h2a)
	) name22929 (
		\m3_addr_i[30]_pad ,
		_w8743_,
		_w8744_,
		_w24830_
	);
	LUT4 #(
		.INIT('habef)
	) name22930 (
		_w8738_,
		_w8741_,
		_w24829_,
		_w24830_,
		_w24831_
	);
	LUT3 #(
		.INIT('h2a)
	) name22931 (
		\m5_addr_i[30]_pad ,
		_w8743_,
		_w8744_,
		_w24832_
	);
	LUT3 #(
		.INIT('h80)
	) name22932 (
		\m6_addr_i[30]_pad ,
		_w8743_,
		_w8744_,
		_w24833_
	);
	LUT4 #(
		.INIT('hcedf)
	) name22933 (
		_w8738_,
		_w8741_,
		_w24832_,
		_w24833_,
		_w24834_
	);
	LUT4 #(
		.INIT('h7fff)
	) name22934 (
		_w24825_,
		_w24828_,
		_w24831_,
		_w24834_,
		_w24835_
	);
	LUT3 #(
		.INIT('h80)
	) name22935 (
		\m0_addr_i[31]_pad ,
		_w8743_,
		_w8744_,
		_w24836_
	);
	LUT3 #(
		.INIT('h2a)
	) name22936 (
		\m7_addr_i[31]_pad ,
		_w8743_,
		_w8744_,
		_w24837_
	);
	LUT4 #(
		.INIT('h6e7f)
	) name22937 (
		_w8738_,
		_w8741_,
		_w24836_,
		_w24837_,
		_w24838_
	);
	LUT3 #(
		.INIT('h2a)
	) name22938 (
		\m3_addr_i[31]_pad ,
		_w8743_,
		_w8744_,
		_w24839_
	);
	LUT3 #(
		.INIT('h80)
	) name22939 (
		\m2_addr_i[31]_pad ,
		_w8743_,
		_w8744_,
		_w24840_
	);
	LUT3 #(
		.INIT('h57)
	) name22940 (
		_w8750_,
		_w24839_,
		_w24840_,
		_w24841_
	);
	LUT3 #(
		.INIT('h80)
	) name22941 (
		\m4_addr_i[31]_pad ,
		_w8743_,
		_w8744_,
		_w24842_
	);
	LUT3 #(
		.INIT('h2a)
	) name22942 (
		\m1_addr_i[31]_pad ,
		_w8743_,
		_w8744_,
		_w24843_
	);
	LUT4 #(
		.INIT('h57df)
	) name22943 (
		_w8738_,
		_w8741_,
		_w24842_,
		_w24843_,
		_w24844_
	);
	LUT3 #(
		.INIT('h2a)
	) name22944 (
		\m5_addr_i[31]_pad ,
		_w8743_,
		_w8744_,
		_w24845_
	);
	LUT3 #(
		.INIT('h80)
	) name22945 (
		\m6_addr_i[31]_pad ,
		_w8743_,
		_w8744_,
		_w24846_
	);
	LUT4 #(
		.INIT('hcedf)
	) name22946 (
		_w8738_,
		_w8741_,
		_w24845_,
		_w24846_,
		_w24847_
	);
	LUT4 #(
		.INIT('h7fff)
	) name22947 (
		_w24838_,
		_w24841_,
		_w24844_,
		_w24847_,
		_w24848_
	);
	LUT3 #(
		.INIT('h2a)
	) name22948 (
		\m3_addr_i[3]_pad ,
		_w8743_,
		_w8744_,
		_w24849_
	);
	LUT3 #(
		.INIT('h80)
	) name22949 (
		\m4_addr_i[3]_pad ,
		_w8743_,
		_w8744_,
		_w24850_
	);
	LUT4 #(
		.INIT('h9dbf)
	) name22950 (
		_w8738_,
		_w8741_,
		_w24849_,
		_w24850_,
		_w24851_
	);
	LUT3 #(
		.INIT('h80)
	) name22951 (
		\m6_addr_i[3]_pad ,
		_w8743_,
		_w8744_,
		_w24852_
	);
	LUT3 #(
		.INIT('h80)
	) name22952 (
		\m2_addr_i[3]_pad ,
		_w8743_,
		_w8744_,
		_w24853_
	);
	LUT4 #(
		.INIT('habef)
	) name22953 (
		_w8738_,
		_w8741_,
		_w24852_,
		_w24853_,
		_w24854_
	);
	LUT3 #(
		.INIT('h2a)
	) name22954 (
		\m5_addr_i[3]_pad ,
		_w8743_,
		_w8744_,
		_w24855_
	);
	LUT3 #(
		.INIT('h2a)
	) name22955 (
		\m1_addr_i[3]_pad ,
		_w8743_,
		_w8744_,
		_w24856_
	);
	LUT4 #(
		.INIT('h57df)
	) name22956 (
		_w8738_,
		_w8741_,
		_w24855_,
		_w24856_,
		_w24857_
	);
	LUT3 #(
		.INIT('h80)
	) name22957 (
		\m0_addr_i[3]_pad ,
		_w8743_,
		_w8744_,
		_w24858_
	);
	LUT3 #(
		.INIT('h2a)
	) name22958 (
		\m7_addr_i[3]_pad ,
		_w8743_,
		_w8744_,
		_w24859_
	);
	LUT4 #(
		.INIT('h6e7f)
	) name22959 (
		_w8738_,
		_w8741_,
		_w24858_,
		_w24859_,
		_w24860_
	);
	LUT4 #(
		.INIT('h7fff)
	) name22960 (
		_w24851_,
		_w24854_,
		_w24857_,
		_w24860_,
		_w24861_
	);
	LUT3 #(
		.INIT('h2a)
	) name22961 (
		\m3_addr_i[4]_pad ,
		_w8743_,
		_w8744_,
		_w24862_
	);
	LUT3 #(
		.INIT('h80)
	) name22962 (
		\m4_addr_i[4]_pad ,
		_w8743_,
		_w8744_,
		_w24863_
	);
	LUT4 #(
		.INIT('h9dbf)
	) name22963 (
		_w8738_,
		_w8741_,
		_w24862_,
		_w24863_,
		_w24864_
	);
	LUT3 #(
		.INIT('h80)
	) name22964 (
		\m6_addr_i[4]_pad ,
		_w8743_,
		_w8744_,
		_w24865_
	);
	LUT3 #(
		.INIT('h80)
	) name22965 (
		\m2_addr_i[4]_pad ,
		_w8743_,
		_w8744_,
		_w24866_
	);
	LUT4 #(
		.INIT('habef)
	) name22966 (
		_w8738_,
		_w8741_,
		_w24865_,
		_w24866_,
		_w24867_
	);
	LUT3 #(
		.INIT('h2a)
	) name22967 (
		\m5_addr_i[4]_pad ,
		_w8743_,
		_w8744_,
		_w24868_
	);
	LUT3 #(
		.INIT('h2a)
	) name22968 (
		\m1_addr_i[4]_pad ,
		_w8743_,
		_w8744_,
		_w24869_
	);
	LUT4 #(
		.INIT('h57df)
	) name22969 (
		_w8738_,
		_w8741_,
		_w24868_,
		_w24869_,
		_w24870_
	);
	LUT3 #(
		.INIT('h80)
	) name22970 (
		\m0_addr_i[4]_pad ,
		_w8743_,
		_w8744_,
		_w24871_
	);
	LUT3 #(
		.INIT('h2a)
	) name22971 (
		\m7_addr_i[4]_pad ,
		_w8743_,
		_w8744_,
		_w24872_
	);
	LUT4 #(
		.INIT('h6e7f)
	) name22972 (
		_w8738_,
		_w8741_,
		_w24871_,
		_w24872_,
		_w24873_
	);
	LUT4 #(
		.INIT('h7fff)
	) name22973 (
		_w24864_,
		_w24867_,
		_w24870_,
		_w24873_,
		_w24874_
	);
	LUT3 #(
		.INIT('h2a)
	) name22974 (
		\m3_addr_i[5]_pad ,
		_w8743_,
		_w8744_,
		_w24875_
	);
	LUT3 #(
		.INIT('h80)
	) name22975 (
		\m4_addr_i[5]_pad ,
		_w8743_,
		_w8744_,
		_w24876_
	);
	LUT4 #(
		.INIT('h9dbf)
	) name22976 (
		_w8738_,
		_w8741_,
		_w24875_,
		_w24876_,
		_w24877_
	);
	LUT3 #(
		.INIT('h80)
	) name22977 (
		\m6_addr_i[5]_pad ,
		_w8743_,
		_w8744_,
		_w24878_
	);
	LUT3 #(
		.INIT('h80)
	) name22978 (
		\m2_addr_i[5]_pad ,
		_w8743_,
		_w8744_,
		_w24879_
	);
	LUT4 #(
		.INIT('habef)
	) name22979 (
		_w8738_,
		_w8741_,
		_w24878_,
		_w24879_,
		_w24880_
	);
	LUT3 #(
		.INIT('h2a)
	) name22980 (
		\m5_addr_i[5]_pad ,
		_w8743_,
		_w8744_,
		_w24881_
	);
	LUT3 #(
		.INIT('h2a)
	) name22981 (
		\m1_addr_i[5]_pad ,
		_w8743_,
		_w8744_,
		_w24882_
	);
	LUT4 #(
		.INIT('h57df)
	) name22982 (
		_w8738_,
		_w8741_,
		_w24881_,
		_w24882_,
		_w24883_
	);
	LUT3 #(
		.INIT('h80)
	) name22983 (
		\m0_addr_i[5]_pad ,
		_w8743_,
		_w8744_,
		_w24884_
	);
	LUT3 #(
		.INIT('h2a)
	) name22984 (
		\m7_addr_i[5]_pad ,
		_w8743_,
		_w8744_,
		_w24885_
	);
	LUT4 #(
		.INIT('h6e7f)
	) name22985 (
		_w8738_,
		_w8741_,
		_w24884_,
		_w24885_,
		_w24886_
	);
	LUT4 #(
		.INIT('h7fff)
	) name22986 (
		_w24877_,
		_w24880_,
		_w24883_,
		_w24886_,
		_w24887_
	);
	LUT3 #(
		.INIT('h2a)
	) name22987 (
		\m3_addr_i[6]_pad ,
		_w8743_,
		_w8744_,
		_w24888_
	);
	LUT3 #(
		.INIT('h80)
	) name22988 (
		\m4_addr_i[6]_pad ,
		_w8743_,
		_w8744_,
		_w24889_
	);
	LUT4 #(
		.INIT('h9dbf)
	) name22989 (
		_w8738_,
		_w8741_,
		_w24888_,
		_w24889_,
		_w24890_
	);
	LUT3 #(
		.INIT('h80)
	) name22990 (
		\m6_addr_i[6]_pad ,
		_w8743_,
		_w8744_,
		_w24891_
	);
	LUT3 #(
		.INIT('h80)
	) name22991 (
		\m2_addr_i[6]_pad ,
		_w8743_,
		_w8744_,
		_w24892_
	);
	LUT4 #(
		.INIT('habef)
	) name22992 (
		_w8738_,
		_w8741_,
		_w24891_,
		_w24892_,
		_w24893_
	);
	LUT3 #(
		.INIT('h2a)
	) name22993 (
		\m5_addr_i[6]_pad ,
		_w8743_,
		_w8744_,
		_w24894_
	);
	LUT3 #(
		.INIT('h2a)
	) name22994 (
		\m1_addr_i[6]_pad ,
		_w8743_,
		_w8744_,
		_w24895_
	);
	LUT4 #(
		.INIT('h57df)
	) name22995 (
		_w8738_,
		_w8741_,
		_w24894_,
		_w24895_,
		_w24896_
	);
	LUT3 #(
		.INIT('h80)
	) name22996 (
		\m0_addr_i[6]_pad ,
		_w8743_,
		_w8744_,
		_w24897_
	);
	LUT3 #(
		.INIT('h2a)
	) name22997 (
		\m7_addr_i[6]_pad ,
		_w8743_,
		_w8744_,
		_w24898_
	);
	LUT4 #(
		.INIT('h6e7f)
	) name22998 (
		_w8738_,
		_w8741_,
		_w24897_,
		_w24898_,
		_w24899_
	);
	LUT4 #(
		.INIT('h7fff)
	) name22999 (
		_w24890_,
		_w24893_,
		_w24896_,
		_w24899_,
		_w24900_
	);
	LUT3 #(
		.INIT('h2a)
	) name23000 (
		\m3_addr_i[7]_pad ,
		_w8743_,
		_w8744_,
		_w24901_
	);
	LUT3 #(
		.INIT('h80)
	) name23001 (
		\m4_addr_i[7]_pad ,
		_w8743_,
		_w8744_,
		_w24902_
	);
	LUT4 #(
		.INIT('h9dbf)
	) name23002 (
		_w8738_,
		_w8741_,
		_w24901_,
		_w24902_,
		_w24903_
	);
	LUT3 #(
		.INIT('h80)
	) name23003 (
		\m6_addr_i[7]_pad ,
		_w8743_,
		_w8744_,
		_w24904_
	);
	LUT3 #(
		.INIT('h80)
	) name23004 (
		\m2_addr_i[7]_pad ,
		_w8743_,
		_w8744_,
		_w24905_
	);
	LUT4 #(
		.INIT('habef)
	) name23005 (
		_w8738_,
		_w8741_,
		_w24904_,
		_w24905_,
		_w24906_
	);
	LUT3 #(
		.INIT('h2a)
	) name23006 (
		\m5_addr_i[7]_pad ,
		_w8743_,
		_w8744_,
		_w24907_
	);
	LUT3 #(
		.INIT('h2a)
	) name23007 (
		\m1_addr_i[7]_pad ,
		_w8743_,
		_w8744_,
		_w24908_
	);
	LUT4 #(
		.INIT('h57df)
	) name23008 (
		_w8738_,
		_w8741_,
		_w24907_,
		_w24908_,
		_w24909_
	);
	LUT3 #(
		.INIT('h80)
	) name23009 (
		\m0_addr_i[7]_pad ,
		_w8743_,
		_w8744_,
		_w24910_
	);
	LUT3 #(
		.INIT('h2a)
	) name23010 (
		\m7_addr_i[7]_pad ,
		_w8743_,
		_w8744_,
		_w24911_
	);
	LUT4 #(
		.INIT('h6e7f)
	) name23011 (
		_w8738_,
		_w8741_,
		_w24910_,
		_w24911_,
		_w24912_
	);
	LUT4 #(
		.INIT('h7fff)
	) name23012 (
		_w24903_,
		_w24906_,
		_w24909_,
		_w24912_,
		_w24913_
	);
	LUT3 #(
		.INIT('h2a)
	) name23013 (
		\m3_addr_i[8]_pad ,
		_w8743_,
		_w8744_,
		_w24914_
	);
	LUT3 #(
		.INIT('h80)
	) name23014 (
		\m4_addr_i[8]_pad ,
		_w8743_,
		_w8744_,
		_w24915_
	);
	LUT4 #(
		.INIT('h9dbf)
	) name23015 (
		_w8738_,
		_w8741_,
		_w24914_,
		_w24915_,
		_w24916_
	);
	LUT3 #(
		.INIT('h80)
	) name23016 (
		\m6_addr_i[8]_pad ,
		_w8743_,
		_w8744_,
		_w24917_
	);
	LUT3 #(
		.INIT('h80)
	) name23017 (
		\m2_addr_i[8]_pad ,
		_w8743_,
		_w8744_,
		_w24918_
	);
	LUT4 #(
		.INIT('habef)
	) name23018 (
		_w8738_,
		_w8741_,
		_w24917_,
		_w24918_,
		_w24919_
	);
	LUT3 #(
		.INIT('h2a)
	) name23019 (
		\m5_addr_i[8]_pad ,
		_w8743_,
		_w8744_,
		_w24920_
	);
	LUT3 #(
		.INIT('h2a)
	) name23020 (
		\m1_addr_i[8]_pad ,
		_w8743_,
		_w8744_,
		_w24921_
	);
	LUT4 #(
		.INIT('h57df)
	) name23021 (
		_w8738_,
		_w8741_,
		_w24920_,
		_w24921_,
		_w24922_
	);
	LUT3 #(
		.INIT('h80)
	) name23022 (
		\m0_addr_i[8]_pad ,
		_w8743_,
		_w8744_,
		_w24923_
	);
	LUT3 #(
		.INIT('h2a)
	) name23023 (
		\m7_addr_i[8]_pad ,
		_w8743_,
		_w8744_,
		_w24924_
	);
	LUT4 #(
		.INIT('h6e7f)
	) name23024 (
		_w8738_,
		_w8741_,
		_w24923_,
		_w24924_,
		_w24925_
	);
	LUT4 #(
		.INIT('h7fff)
	) name23025 (
		_w24916_,
		_w24919_,
		_w24922_,
		_w24925_,
		_w24926_
	);
	LUT3 #(
		.INIT('h2a)
	) name23026 (
		\m3_addr_i[9]_pad ,
		_w8743_,
		_w8744_,
		_w24927_
	);
	LUT3 #(
		.INIT('h80)
	) name23027 (
		\m4_addr_i[9]_pad ,
		_w8743_,
		_w8744_,
		_w24928_
	);
	LUT4 #(
		.INIT('h9dbf)
	) name23028 (
		_w8738_,
		_w8741_,
		_w24927_,
		_w24928_,
		_w24929_
	);
	LUT3 #(
		.INIT('h80)
	) name23029 (
		\m6_addr_i[9]_pad ,
		_w8743_,
		_w8744_,
		_w24930_
	);
	LUT3 #(
		.INIT('h80)
	) name23030 (
		\m2_addr_i[9]_pad ,
		_w8743_,
		_w8744_,
		_w24931_
	);
	LUT4 #(
		.INIT('habef)
	) name23031 (
		_w8738_,
		_w8741_,
		_w24930_,
		_w24931_,
		_w24932_
	);
	LUT3 #(
		.INIT('h2a)
	) name23032 (
		\m5_addr_i[9]_pad ,
		_w8743_,
		_w8744_,
		_w24933_
	);
	LUT3 #(
		.INIT('h2a)
	) name23033 (
		\m1_addr_i[9]_pad ,
		_w8743_,
		_w8744_,
		_w24934_
	);
	LUT4 #(
		.INIT('h57df)
	) name23034 (
		_w8738_,
		_w8741_,
		_w24933_,
		_w24934_,
		_w24935_
	);
	LUT3 #(
		.INIT('h80)
	) name23035 (
		\m0_addr_i[9]_pad ,
		_w8743_,
		_w8744_,
		_w24936_
	);
	LUT3 #(
		.INIT('h2a)
	) name23036 (
		\m7_addr_i[9]_pad ,
		_w8743_,
		_w8744_,
		_w24937_
	);
	LUT4 #(
		.INIT('h6e7f)
	) name23037 (
		_w8738_,
		_w8741_,
		_w24936_,
		_w24937_,
		_w24938_
	);
	LUT4 #(
		.INIT('h7fff)
	) name23038 (
		_w24929_,
		_w24932_,
		_w24935_,
		_w24938_,
		_w24939_
	);
	LUT3 #(
		.INIT('h80)
	) name23039 (
		\m0_data_i[0]_pad ,
		_w8743_,
		_w8744_,
		_w24940_
	);
	LUT3 #(
		.INIT('h2a)
	) name23040 (
		\m7_data_i[0]_pad ,
		_w8743_,
		_w8744_,
		_w24941_
	);
	LUT4 #(
		.INIT('h6e7f)
	) name23041 (
		_w8738_,
		_w8741_,
		_w24940_,
		_w24941_,
		_w24942_
	);
	LUT3 #(
		.INIT('h80)
	) name23042 (
		\m6_data_i[0]_pad ,
		_w8743_,
		_w8744_,
		_w24943_
	);
	LUT3 #(
		.INIT('h80)
	) name23043 (
		\m2_data_i[0]_pad ,
		_w8743_,
		_w8744_,
		_w24944_
	);
	LUT4 #(
		.INIT('habef)
	) name23044 (
		_w8738_,
		_w8741_,
		_w24943_,
		_w24944_,
		_w24945_
	);
	LUT3 #(
		.INIT('h2a)
	) name23045 (
		\m5_data_i[0]_pad ,
		_w8743_,
		_w8744_,
		_w24946_
	);
	LUT3 #(
		.INIT('h2a)
	) name23046 (
		\m1_data_i[0]_pad ,
		_w8743_,
		_w8744_,
		_w24947_
	);
	LUT4 #(
		.INIT('h57df)
	) name23047 (
		_w8738_,
		_w8741_,
		_w24946_,
		_w24947_,
		_w24948_
	);
	LUT3 #(
		.INIT('h2a)
	) name23048 (
		\m3_data_i[0]_pad ,
		_w8743_,
		_w8744_,
		_w24949_
	);
	LUT3 #(
		.INIT('h80)
	) name23049 (
		\m4_data_i[0]_pad ,
		_w8743_,
		_w8744_,
		_w24950_
	);
	LUT4 #(
		.INIT('h9dbf)
	) name23050 (
		_w8738_,
		_w8741_,
		_w24949_,
		_w24950_,
		_w24951_
	);
	LUT4 #(
		.INIT('h7fff)
	) name23051 (
		_w24942_,
		_w24945_,
		_w24948_,
		_w24951_,
		_w24952_
	);
	LUT3 #(
		.INIT('h80)
	) name23052 (
		\m0_data_i[10]_pad ,
		_w8743_,
		_w8744_,
		_w24953_
	);
	LUT3 #(
		.INIT('h2a)
	) name23053 (
		\m7_data_i[10]_pad ,
		_w8743_,
		_w8744_,
		_w24954_
	);
	LUT4 #(
		.INIT('h6e7f)
	) name23054 (
		_w8738_,
		_w8741_,
		_w24953_,
		_w24954_,
		_w24955_
	);
	LUT3 #(
		.INIT('h80)
	) name23055 (
		\m6_data_i[10]_pad ,
		_w8743_,
		_w8744_,
		_w24956_
	);
	LUT3 #(
		.INIT('h80)
	) name23056 (
		\m2_data_i[10]_pad ,
		_w8743_,
		_w8744_,
		_w24957_
	);
	LUT4 #(
		.INIT('habef)
	) name23057 (
		_w8738_,
		_w8741_,
		_w24956_,
		_w24957_,
		_w24958_
	);
	LUT3 #(
		.INIT('h2a)
	) name23058 (
		\m5_data_i[10]_pad ,
		_w8743_,
		_w8744_,
		_w24959_
	);
	LUT3 #(
		.INIT('h2a)
	) name23059 (
		\m1_data_i[10]_pad ,
		_w8743_,
		_w8744_,
		_w24960_
	);
	LUT4 #(
		.INIT('h57df)
	) name23060 (
		_w8738_,
		_w8741_,
		_w24959_,
		_w24960_,
		_w24961_
	);
	LUT3 #(
		.INIT('h2a)
	) name23061 (
		\m3_data_i[10]_pad ,
		_w8743_,
		_w8744_,
		_w24962_
	);
	LUT3 #(
		.INIT('h80)
	) name23062 (
		\m4_data_i[10]_pad ,
		_w8743_,
		_w8744_,
		_w24963_
	);
	LUT4 #(
		.INIT('h9dbf)
	) name23063 (
		_w8738_,
		_w8741_,
		_w24962_,
		_w24963_,
		_w24964_
	);
	LUT4 #(
		.INIT('h7fff)
	) name23064 (
		_w24955_,
		_w24958_,
		_w24961_,
		_w24964_,
		_w24965_
	);
	LUT3 #(
		.INIT('h2a)
	) name23065 (
		\m3_data_i[11]_pad ,
		_w8743_,
		_w8744_,
		_w24966_
	);
	LUT3 #(
		.INIT('h80)
	) name23066 (
		\m4_data_i[11]_pad ,
		_w8743_,
		_w8744_,
		_w24967_
	);
	LUT4 #(
		.INIT('h9dbf)
	) name23067 (
		_w8738_,
		_w8741_,
		_w24966_,
		_w24967_,
		_w24968_
	);
	LUT3 #(
		.INIT('h80)
	) name23068 (
		\m6_data_i[11]_pad ,
		_w8743_,
		_w8744_,
		_w24969_
	);
	LUT3 #(
		.INIT('h2a)
	) name23069 (
		\m7_data_i[11]_pad ,
		_w8743_,
		_w8744_,
		_w24970_
	);
	LUT3 #(
		.INIT('h57)
	) name23070 (
		_w8756_,
		_w24969_,
		_w24970_,
		_w24971_
	);
	LUT3 #(
		.INIT('h2a)
	) name23071 (
		\m5_data_i[11]_pad ,
		_w8743_,
		_w8744_,
		_w24972_
	);
	LUT3 #(
		.INIT('h80)
	) name23072 (
		\m0_data_i[11]_pad ,
		_w8743_,
		_w8744_,
		_w24973_
	);
	LUT4 #(
		.INIT('h57df)
	) name23073 (
		_w8738_,
		_w8741_,
		_w24972_,
		_w24973_,
		_w24974_
	);
	LUT3 #(
		.INIT('h2a)
	) name23074 (
		\m1_data_i[11]_pad ,
		_w8743_,
		_w8744_,
		_w24975_
	);
	LUT3 #(
		.INIT('h80)
	) name23075 (
		\m2_data_i[11]_pad ,
		_w8743_,
		_w8744_,
		_w24976_
	);
	LUT4 #(
		.INIT('h3b7f)
	) name23076 (
		_w8738_,
		_w8741_,
		_w24975_,
		_w24976_,
		_w24977_
	);
	LUT4 #(
		.INIT('h7fff)
	) name23077 (
		_w24968_,
		_w24971_,
		_w24974_,
		_w24977_,
		_w24978_
	);
	LUT3 #(
		.INIT('h2a)
	) name23078 (
		\m3_data_i[12]_pad ,
		_w8743_,
		_w8744_,
		_w24979_
	);
	LUT3 #(
		.INIT('h80)
	) name23079 (
		\m4_data_i[12]_pad ,
		_w8743_,
		_w8744_,
		_w24980_
	);
	LUT4 #(
		.INIT('h9dbf)
	) name23080 (
		_w8738_,
		_w8741_,
		_w24979_,
		_w24980_,
		_w24981_
	);
	LUT3 #(
		.INIT('h80)
	) name23081 (
		\m6_data_i[12]_pad ,
		_w8743_,
		_w8744_,
		_w24982_
	);
	LUT3 #(
		.INIT('h80)
	) name23082 (
		\m2_data_i[12]_pad ,
		_w8743_,
		_w8744_,
		_w24983_
	);
	LUT4 #(
		.INIT('habef)
	) name23083 (
		_w8738_,
		_w8741_,
		_w24982_,
		_w24983_,
		_w24984_
	);
	LUT3 #(
		.INIT('h2a)
	) name23084 (
		\m5_data_i[12]_pad ,
		_w8743_,
		_w8744_,
		_w24985_
	);
	LUT3 #(
		.INIT('h2a)
	) name23085 (
		\m1_data_i[12]_pad ,
		_w8743_,
		_w8744_,
		_w24986_
	);
	LUT4 #(
		.INIT('h57df)
	) name23086 (
		_w8738_,
		_w8741_,
		_w24985_,
		_w24986_,
		_w24987_
	);
	LUT3 #(
		.INIT('h80)
	) name23087 (
		\m0_data_i[12]_pad ,
		_w8743_,
		_w8744_,
		_w24988_
	);
	LUT3 #(
		.INIT('h2a)
	) name23088 (
		\m7_data_i[12]_pad ,
		_w8743_,
		_w8744_,
		_w24989_
	);
	LUT4 #(
		.INIT('h6e7f)
	) name23089 (
		_w8738_,
		_w8741_,
		_w24988_,
		_w24989_,
		_w24990_
	);
	LUT4 #(
		.INIT('h7fff)
	) name23090 (
		_w24981_,
		_w24984_,
		_w24987_,
		_w24990_,
		_w24991_
	);
	LUT3 #(
		.INIT('h80)
	) name23091 (
		\m0_data_i[13]_pad ,
		_w8743_,
		_w8744_,
		_w24992_
	);
	LUT3 #(
		.INIT('h2a)
	) name23092 (
		\m7_data_i[13]_pad ,
		_w8743_,
		_w8744_,
		_w24993_
	);
	LUT4 #(
		.INIT('h6e7f)
	) name23093 (
		_w8738_,
		_w8741_,
		_w24992_,
		_w24993_,
		_w24994_
	);
	LUT3 #(
		.INIT('h80)
	) name23094 (
		\m6_data_i[13]_pad ,
		_w8743_,
		_w8744_,
		_w24995_
	);
	LUT3 #(
		.INIT('h80)
	) name23095 (
		\m2_data_i[13]_pad ,
		_w8743_,
		_w8744_,
		_w24996_
	);
	LUT4 #(
		.INIT('habef)
	) name23096 (
		_w8738_,
		_w8741_,
		_w24995_,
		_w24996_,
		_w24997_
	);
	LUT3 #(
		.INIT('h2a)
	) name23097 (
		\m5_data_i[13]_pad ,
		_w8743_,
		_w8744_,
		_w24998_
	);
	LUT3 #(
		.INIT('h2a)
	) name23098 (
		\m1_data_i[13]_pad ,
		_w8743_,
		_w8744_,
		_w24999_
	);
	LUT4 #(
		.INIT('h57df)
	) name23099 (
		_w8738_,
		_w8741_,
		_w24998_,
		_w24999_,
		_w25000_
	);
	LUT3 #(
		.INIT('h2a)
	) name23100 (
		\m3_data_i[13]_pad ,
		_w8743_,
		_w8744_,
		_w25001_
	);
	LUT3 #(
		.INIT('h80)
	) name23101 (
		\m4_data_i[13]_pad ,
		_w8743_,
		_w8744_,
		_w25002_
	);
	LUT4 #(
		.INIT('h9dbf)
	) name23102 (
		_w8738_,
		_w8741_,
		_w25001_,
		_w25002_,
		_w25003_
	);
	LUT4 #(
		.INIT('h7fff)
	) name23103 (
		_w24994_,
		_w24997_,
		_w25000_,
		_w25003_,
		_w25004_
	);
	LUT3 #(
		.INIT('h80)
	) name23104 (
		\m0_data_i[14]_pad ,
		_w8743_,
		_w8744_,
		_w25005_
	);
	LUT3 #(
		.INIT('h2a)
	) name23105 (
		\m7_data_i[14]_pad ,
		_w8743_,
		_w8744_,
		_w25006_
	);
	LUT4 #(
		.INIT('h6e7f)
	) name23106 (
		_w8738_,
		_w8741_,
		_w25005_,
		_w25006_,
		_w25007_
	);
	LUT3 #(
		.INIT('h80)
	) name23107 (
		\m6_data_i[14]_pad ,
		_w8743_,
		_w8744_,
		_w25008_
	);
	LUT3 #(
		.INIT('h80)
	) name23108 (
		\m2_data_i[14]_pad ,
		_w8743_,
		_w8744_,
		_w25009_
	);
	LUT4 #(
		.INIT('habef)
	) name23109 (
		_w8738_,
		_w8741_,
		_w25008_,
		_w25009_,
		_w25010_
	);
	LUT3 #(
		.INIT('h2a)
	) name23110 (
		\m5_data_i[14]_pad ,
		_w8743_,
		_w8744_,
		_w25011_
	);
	LUT3 #(
		.INIT('h2a)
	) name23111 (
		\m1_data_i[14]_pad ,
		_w8743_,
		_w8744_,
		_w25012_
	);
	LUT4 #(
		.INIT('h57df)
	) name23112 (
		_w8738_,
		_w8741_,
		_w25011_,
		_w25012_,
		_w25013_
	);
	LUT3 #(
		.INIT('h2a)
	) name23113 (
		\m3_data_i[14]_pad ,
		_w8743_,
		_w8744_,
		_w25014_
	);
	LUT3 #(
		.INIT('h80)
	) name23114 (
		\m4_data_i[14]_pad ,
		_w8743_,
		_w8744_,
		_w25015_
	);
	LUT4 #(
		.INIT('h9dbf)
	) name23115 (
		_w8738_,
		_w8741_,
		_w25014_,
		_w25015_,
		_w25016_
	);
	LUT4 #(
		.INIT('h7fff)
	) name23116 (
		_w25007_,
		_w25010_,
		_w25013_,
		_w25016_,
		_w25017_
	);
	LUT3 #(
		.INIT('h2a)
	) name23117 (
		\m3_data_i[15]_pad ,
		_w8743_,
		_w8744_,
		_w25018_
	);
	LUT3 #(
		.INIT('h80)
	) name23118 (
		\m4_data_i[15]_pad ,
		_w8743_,
		_w8744_,
		_w25019_
	);
	LUT4 #(
		.INIT('h9dbf)
	) name23119 (
		_w8738_,
		_w8741_,
		_w25018_,
		_w25019_,
		_w25020_
	);
	LUT3 #(
		.INIT('h80)
	) name23120 (
		\m6_data_i[15]_pad ,
		_w8743_,
		_w8744_,
		_w25021_
	);
	LUT3 #(
		.INIT('h80)
	) name23121 (
		\m2_data_i[15]_pad ,
		_w8743_,
		_w8744_,
		_w25022_
	);
	LUT4 #(
		.INIT('habef)
	) name23122 (
		_w8738_,
		_w8741_,
		_w25021_,
		_w25022_,
		_w25023_
	);
	LUT3 #(
		.INIT('h2a)
	) name23123 (
		\m5_data_i[15]_pad ,
		_w8743_,
		_w8744_,
		_w25024_
	);
	LUT3 #(
		.INIT('h2a)
	) name23124 (
		\m1_data_i[15]_pad ,
		_w8743_,
		_w8744_,
		_w25025_
	);
	LUT4 #(
		.INIT('h57df)
	) name23125 (
		_w8738_,
		_w8741_,
		_w25024_,
		_w25025_,
		_w25026_
	);
	LUT3 #(
		.INIT('h80)
	) name23126 (
		\m0_data_i[15]_pad ,
		_w8743_,
		_w8744_,
		_w25027_
	);
	LUT3 #(
		.INIT('h2a)
	) name23127 (
		\m7_data_i[15]_pad ,
		_w8743_,
		_w8744_,
		_w25028_
	);
	LUT4 #(
		.INIT('h6e7f)
	) name23128 (
		_w8738_,
		_w8741_,
		_w25027_,
		_w25028_,
		_w25029_
	);
	LUT4 #(
		.INIT('h7fff)
	) name23129 (
		_w25020_,
		_w25023_,
		_w25026_,
		_w25029_,
		_w25030_
	);
	LUT3 #(
		.INIT('h2a)
	) name23130 (
		\m3_data_i[16]_pad ,
		_w8743_,
		_w8744_,
		_w25031_
	);
	LUT3 #(
		.INIT('h80)
	) name23131 (
		\m4_data_i[16]_pad ,
		_w8743_,
		_w8744_,
		_w25032_
	);
	LUT4 #(
		.INIT('h9dbf)
	) name23132 (
		_w8738_,
		_w8741_,
		_w25031_,
		_w25032_,
		_w25033_
	);
	LUT3 #(
		.INIT('h80)
	) name23133 (
		\m6_data_i[16]_pad ,
		_w8743_,
		_w8744_,
		_w25034_
	);
	LUT3 #(
		.INIT('h80)
	) name23134 (
		\m2_data_i[16]_pad ,
		_w8743_,
		_w8744_,
		_w25035_
	);
	LUT4 #(
		.INIT('habef)
	) name23135 (
		_w8738_,
		_w8741_,
		_w25034_,
		_w25035_,
		_w25036_
	);
	LUT3 #(
		.INIT('h2a)
	) name23136 (
		\m5_data_i[16]_pad ,
		_w8743_,
		_w8744_,
		_w25037_
	);
	LUT3 #(
		.INIT('h2a)
	) name23137 (
		\m1_data_i[16]_pad ,
		_w8743_,
		_w8744_,
		_w25038_
	);
	LUT4 #(
		.INIT('h57df)
	) name23138 (
		_w8738_,
		_w8741_,
		_w25037_,
		_w25038_,
		_w25039_
	);
	LUT3 #(
		.INIT('h80)
	) name23139 (
		\m0_data_i[16]_pad ,
		_w8743_,
		_w8744_,
		_w25040_
	);
	LUT3 #(
		.INIT('h2a)
	) name23140 (
		\m7_data_i[16]_pad ,
		_w8743_,
		_w8744_,
		_w25041_
	);
	LUT4 #(
		.INIT('h6e7f)
	) name23141 (
		_w8738_,
		_w8741_,
		_w25040_,
		_w25041_,
		_w25042_
	);
	LUT4 #(
		.INIT('h7fff)
	) name23142 (
		_w25033_,
		_w25036_,
		_w25039_,
		_w25042_,
		_w25043_
	);
	LUT3 #(
		.INIT('h2a)
	) name23143 (
		\m3_data_i[17]_pad ,
		_w8743_,
		_w8744_,
		_w25044_
	);
	LUT3 #(
		.INIT('h80)
	) name23144 (
		\m4_data_i[17]_pad ,
		_w8743_,
		_w8744_,
		_w25045_
	);
	LUT4 #(
		.INIT('h9dbf)
	) name23145 (
		_w8738_,
		_w8741_,
		_w25044_,
		_w25045_,
		_w25046_
	);
	LUT3 #(
		.INIT('h80)
	) name23146 (
		\m6_data_i[17]_pad ,
		_w8743_,
		_w8744_,
		_w25047_
	);
	LUT3 #(
		.INIT('h80)
	) name23147 (
		\m2_data_i[17]_pad ,
		_w8743_,
		_w8744_,
		_w25048_
	);
	LUT4 #(
		.INIT('habef)
	) name23148 (
		_w8738_,
		_w8741_,
		_w25047_,
		_w25048_,
		_w25049_
	);
	LUT3 #(
		.INIT('h2a)
	) name23149 (
		\m5_data_i[17]_pad ,
		_w8743_,
		_w8744_,
		_w25050_
	);
	LUT3 #(
		.INIT('h2a)
	) name23150 (
		\m1_data_i[17]_pad ,
		_w8743_,
		_w8744_,
		_w25051_
	);
	LUT4 #(
		.INIT('h57df)
	) name23151 (
		_w8738_,
		_w8741_,
		_w25050_,
		_w25051_,
		_w25052_
	);
	LUT3 #(
		.INIT('h80)
	) name23152 (
		\m0_data_i[17]_pad ,
		_w8743_,
		_w8744_,
		_w25053_
	);
	LUT3 #(
		.INIT('h2a)
	) name23153 (
		\m7_data_i[17]_pad ,
		_w8743_,
		_w8744_,
		_w25054_
	);
	LUT4 #(
		.INIT('h6e7f)
	) name23154 (
		_w8738_,
		_w8741_,
		_w25053_,
		_w25054_,
		_w25055_
	);
	LUT4 #(
		.INIT('h7fff)
	) name23155 (
		_w25046_,
		_w25049_,
		_w25052_,
		_w25055_,
		_w25056_
	);
	LUT3 #(
		.INIT('h2a)
	) name23156 (
		\m1_data_i[18]_pad ,
		_w8743_,
		_w8744_,
		_w25057_
	);
	LUT3 #(
		.INIT('h80)
	) name23157 (
		\m2_data_i[18]_pad ,
		_w8743_,
		_w8744_,
		_w25058_
	);
	LUT4 #(
		.INIT('h3b7f)
	) name23158 (
		_w8738_,
		_w8741_,
		_w25057_,
		_w25058_,
		_w25059_
	);
	LUT3 #(
		.INIT('h80)
	) name23159 (
		\m6_data_i[18]_pad ,
		_w8743_,
		_w8744_,
		_w25060_
	);
	LUT3 #(
		.INIT('h2a)
	) name23160 (
		\m7_data_i[18]_pad ,
		_w8743_,
		_w8744_,
		_w25061_
	);
	LUT3 #(
		.INIT('h57)
	) name23161 (
		_w8756_,
		_w25060_,
		_w25061_,
		_w25062_
	);
	LUT3 #(
		.INIT('h2a)
	) name23162 (
		\m5_data_i[18]_pad ,
		_w8743_,
		_w8744_,
		_w25063_
	);
	LUT3 #(
		.INIT('h80)
	) name23163 (
		\m0_data_i[18]_pad ,
		_w8743_,
		_w8744_,
		_w25064_
	);
	LUT4 #(
		.INIT('h57df)
	) name23164 (
		_w8738_,
		_w8741_,
		_w25063_,
		_w25064_,
		_w25065_
	);
	LUT3 #(
		.INIT('h2a)
	) name23165 (
		\m3_data_i[18]_pad ,
		_w8743_,
		_w8744_,
		_w25066_
	);
	LUT3 #(
		.INIT('h80)
	) name23166 (
		\m4_data_i[18]_pad ,
		_w8743_,
		_w8744_,
		_w25067_
	);
	LUT4 #(
		.INIT('h9dbf)
	) name23167 (
		_w8738_,
		_w8741_,
		_w25066_,
		_w25067_,
		_w25068_
	);
	LUT4 #(
		.INIT('h7fff)
	) name23168 (
		_w25059_,
		_w25062_,
		_w25065_,
		_w25068_,
		_w25069_
	);
	LUT3 #(
		.INIT('h2a)
	) name23169 (
		\m3_data_i[19]_pad ,
		_w8743_,
		_w8744_,
		_w25070_
	);
	LUT3 #(
		.INIT('h80)
	) name23170 (
		\m4_data_i[19]_pad ,
		_w8743_,
		_w8744_,
		_w25071_
	);
	LUT4 #(
		.INIT('h9dbf)
	) name23171 (
		_w8738_,
		_w8741_,
		_w25070_,
		_w25071_,
		_w25072_
	);
	LUT3 #(
		.INIT('h80)
	) name23172 (
		\m6_data_i[19]_pad ,
		_w8743_,
		_w8744_,
		_w25073_
	);
	LUT3 #(
		.INIT('h80)
	) name23173 (
		\m2_data_i[19]_pad ,
		_w8743_,
		_w8744_,
		_w25074_
	);
	LUT4 #(
		.INIT('habef)
	) name23174 (
		_w8738_,
		_w8741_,
		_w25073_,
		_w25074_,
		_w25075_
	);
	LUT3 #(
		.INIT('h2a)
	) name23175 (
		\m5_data_i[19]_pad ,
		_w8743_,
		_w8744_,
		_w25076_
	);
	LUT3 #(
		.INIT('h2a)
	) name23176 (
		\m1_data_i[19]_pad ,
		_w8743_,
		_w8744_,
		_w25077_
	);
	LUT4 #(
		.INIT('h57df)
	) name23177 (
		_w8738_,
		_w8741_,
		_w25076_,
		_w25077_,
		_w25078_
	);
	LUT3 #(
		.INIT('h80)
	) name23178 (
		\m0_data_i[19]_pad ,
		_w8743_,
		_w8744_,
		_w25079_
	);
	LUT3 #(
		.INIT('h2a)
	) name23179 (
		\m7_data_i[19]_pad ,
		_w8743_,
		_w8744_,
		_w25080_
	);
	LUT4 #(
		.INIT('h6e7f)
	) name23180 (
		_w8738_,
		_w8741_,
		_w25079_,
		_w25080_,
		_w25081_
	);
	LUT4 #(
		.INIT('h7fff)
	) name23181 (
		_w25072_,
		_w25075_,
		_w25078_,
		_w25081_,
		_w25082_
	);
	LUT3 #(
		.INIT('h2a)
	) name23182 (
		\m1_data_i[1]_pad ,
		_w8743_,
		_w8744_,
		_w25083_
	);
	LUT3 #(
		.INIT('h80)
	) name23183 (
		\m2_data_i[1]_pad ,
		_w8743_,
		_w8744_,
		_w25084_
	);
	LUT4 #(
		.INIT('h3b7f)
	) name23184 (
		_w8738_,
		_w8741_,
		_w25083_,
		_w25084_,
		_w25085_
	);
	LUT3 #(
		.INIT('h80)
	) name23185 (
		\m0_data_i[1]_pad ,
		_w8743_,
		_w8744_,
		_w25086_
	);
	LUT3 #(
		.INIT('h80)
	) name23186 (
		\m4_data_i[1]_pad ,
		_w8743_,
		_w8744_,
		_w25087_
	);
	LUT4 #(
		.INIT('h5d7f)
	) name23187 (
		_w8738_,
		_w8741_,
		_w25086_,
		_w25087_,
		_w25088_
	);
	LUT3 #(
		.INIT('h2a)
	) name23188 (
		\m7_data_i[1]_pad ,
		_w8743_,
		_w8744_,
		_w25089_
	);
	LUT3 #(
		.INIT('h2a)
	) name23189 (
		\m3_data_i[1]_pad ,
		_w8743_,
		_w8744_,
		_w25090_
	);
	LUT4 #(
		.INIT('habef)
	) name23190 (
		_w8738_,
		_w8741_,
		_w25089_,
		_w25090_,
		_w25091_
	);
	LUT3 #(
		.INIT('h80)
	) name23191 (
		\m6_data_i[1]_pad ,
		_w8743_,
		_w8744_,
		_w25092_
	);
	LUT3 #(
		.INIT('h2a)
	) name23192 (
		\m5_data_i[1]_pad ,
		_w8743_,
		_w8744_,
		_w25093_
	);
	LUT4 #(
		.INIT('hcdef)
	) name23193 (
		_w8738_,
		_w8741_,
		_w25092_,
		_w25093_,
		_w25094_
	);
	LUT4 #(
		.INIT('h7fff)
	) name23194 (
		_w25085_,
		_w25088_,
		_w25091_,
		_w25094_,
		_w25095_
	);
	LUT3 #(
		.INIT('h2a)
	) name23195 (
		\m3_data_i[20]_pad ,
		_w8743_,
		_w8744_,
		_w25096_
	);
	LUT3 #(
		.INIT('h80)
	) name23196 (
		\m4_data_i[20]_pad ,
		_w8743_,
		_w8744_,
		_w25097_
	);
	LUT4 #(
		.INIT('h9dbf)
	) name23197 (
		_w8738_,
		_w8741_,
		_w25096_,
		_w25097_,
		_w25098_
	);
	LUT3 #(
		.INIT('h80)
	) name23198 (
		\m6_data_i[20]_pad ,
		_w8743_,
		_w8744_,
		_w25099_
	);
	LUT3 #(
		.INIT('h80)
	) name23199 (
		\m2_data_i[20]_pad ,
		_w8743_,
		_w8744_,
		_w25100_
	);
	LUT4 #(
		.INIT('habef)
	) name23200 (
		_w8738_,
		_w8741_,
		_w25099_,
		_w25100_,
		_w25101_
	);
	LUT3 #(
		.INIT('h2a)
	) name23201 (
		\m5_data_i[20]_pad ,
		_w8743_,
		_w8744_,
		_w25102_
	);
	LUT3 #(
		.INIT('h2a)
	) name23202 (
		\m1_data_i[20]_pad ,
		_w8743_,
		_w8744_,
		_w25103_
	);
	LUT4 #(
		.INIT('h57df)
	) name23203 (
		_w8738_,
		_w8741_,
		_w25102_,
		_w25103_,
		_w25104_
	);
	LUT3 #(
		.INIT('h80)
	) name23204 (
		\m0_data_i[20]_pad ,
		_w8743_,
		_w8744_,
		_w25105_
	);
	LUT3 #(
		.INIT('h2a)
	) name23205 (
		\m7_data_i[20]_pad ,
		_w8743_,
		_w8744_,
		_w25106_
	);
	LUT4 #(
		.INIT('h6e7f)
	) name23206 (
		_w8738_,
		_w8741_,
		_w25105_,
		_w25106_,
		_w25107_
	);
	LUT4 #(
		.INIT('h7fff)
	) name23207 (
		_w25098_,
		_w25101_,
		_w25104_,
		_w25107_,
		_w25108_
	);
	LUT3 #(
		.INIT('h2a)
	) name23208 (
		\m3_data_i[21]_pad ,
		_w8743_,
		_w8744_,
		_w25109_
	);
	LUT3 #(
		.INIT('h80)
	) name23209 (
		\m4_data_i[21]_pad ,
		_w8743_,
		_w8744_,
		_w25110_
	);
	LUT4 #(
		.INIT('h9dbf)
	) name23210 (
		_w8738_,
		_w8741_,
		_w25109_,
		_w25110_,
		_w25111_
	);
	LUT3 #(
		.INIT('h80)
	) name23211 (
		\m6_data_i[21]_pad ,
		_w8743_,
		_w8744_,
		_w25112_
	);
	LUT3 #(
		.INIT('h80)
	) name23212 (
		\m2_data_i[21]_pad ,
		_w8743_,
		_w8744_,
		_w25113_
	);
	LUT4 #(
		.INIT('habef)
	) name23213 (
		_w8738_,
		_w8741_,
		_w25112_,
		_w25113_,
		_w25114_
	);
	LUT3 #(
		.INIT('h2a)
	) name23214 (
		\m5_data_i[21]_pad ,
		_w8743_,
		_w8744_,
		_w25115_
	);
	LUT3 #(
		.INIT('h2a)
	) name23215 (
		\m1_data_i[21]_pad ,
		_w8743_,
		_w8744_,
		_w25116_
	);
	LUT4 #(
		.INIT('h57df)
	) name23216 (
		_w8738_,
		_w8741_,
		_w25115_,
		_w25116_,
		_w25117_
	);
	LUT3 #(
		.INIT('h80)
	) name23217 (
		\m0_data_i[21]_pad ,
		_w8743_,
		_w8744_,
		_w25118_
	);
	LUT3 #(
		.INIT('h2a)
	) name23218 (
		\m7_data_i[21]_pad ,
		_w8743_,
		_w8744_,
		_w25119_
	);
	LUT4 #(
		.INIT('h6e7f)
	) name23219 (
		_w8738_,
		_w8741_,
		_w25118_,
		_w25119_,
		_w25120_
	);
	LUT4 #(
		.INIT('h7fff)
	) name23220 (
		_w25111_,
		_w25114_,
		_w25117_,
		_w25120_,
		_w25121_
	);
	LUT3 #(
		.INIT('h2a)
	) name23221 (
		\m3_data_i[22]_pad ,
		_w8743_,
		_w8744_,
		_w25122_
	);
	LUT3 #(
		.INIT('h80)
	) name23222 (
		\m4_data_i[22]_pad ,
		_w8743_,
		_w8744_,
		_w25123_
	);
	LUT4 #(
		.INIT('h9dbf)
	) name23223 (
		_w8738_,
		_w8741_,
		_w25122_,
		_w25123_,
		_w25124_
	);
	LUT3 #(
		.INIT('h80)
	) name23224 (
		\m6_data_i[22]_pad ,
		_w8743_,
		_w8744_,
		_w25125_
	);
	LUT3 #(
		.INIT('h80)
	) name23225 (
		\m2_data_i[22]_pad ,
		_w8743_,
		_w8744_,
		_w25126_
	);
	LUT4 #(
		.INIT('habef)
	) name23226 (
		_w8738_,
		_w8741_,
		_w25125_,
		_w25126_,
		_w25127_
	);
	LUT3 #(
		.INIT('h2a)
	) name23227 (
		\m5_data_i[22]_pad ,
		_w8743_,
		_w8744_,
		_w25128_
	);
	LUT3 #(
		.INIT('h2a)
	) name23228 (
		\m1_data_i[22]_pad ,
		_w8743_,
		_w8744_,
		_w25129_
	);
	LUT4 #(
		.INIT('h57df)
	) name23229 (
		_w8738_,
		_w8741_,
		_w25128_,
		_w25129_,
		_w25130_
	);
	LUT3 #(
		.INIT('h80)
	) name23230 (
		\m0_data_i[22]_pad ,
		_w8743_,
		_w8744_,
		_w25131_
	);
	LUT3 #(
		.INIT('h2a)
	) name23231 (
		\m7_data_i[22]_pad ,
		_w8743_,
		_w8744_,
		_w25132_
	);
	LUT4 #(
		.INIT('h6e7f)
	) name23232 (
		_w8738_,
		_w8741_,
		_w25131_,
		_w25132_,
		_w25133_
	);
	LUT4 #(
		.INIT('h7fff)
	) name23233 (
		_w25124_,
		_w25127_,
		_w25130_,
		_w25133_,
		_w25134_
	);
	LUT3 #(
		.INIT('h80)
	) name23234 (
		\m0_data_i[23]_pad ,
		_w8743_,
		_w8744_,
		_w25135_
	);
	LUT3 #(
		.INIT('h2a)
	) name23235 (
		\m7_data_i[23]_pad ,
		_w8743_,
		_w8744_,
		_w25136_
	);
	LUT4 #(
		.INIT('h6e7f)
	) name23236 (
		_w8738_,
		_w8741_,
		_w25135_,
		_w25136_,
		_w25137_
	);
	LUT3 #(
		.INIT('h2a)
	) name23237 (
		\m3_data_i[23]_pad ,
		_w8743_,
		_w8744_,
		_w25138_
	);
	LUT3 #(
		.INIT('h2a)
	) name23238 (
		\m5_data_i[23]_pad ,
		_w8743_,
		_w8744_,
		_w25139_
	);
	LUT4 #(
		.INIT('h9dbf)
	) name23239 (
		_w8738_,
		_w8741_,
		_w25138_,
		_w25139_,
		_w25140_
	);
	LUT3 #(
		.INIT('h80)
	) name23240 (
		\m4_data_i[23]_pad ,
		_w8743_,
		_w8744_,
		_w25141_
	);
	LUT3 #(
		.INIT('h80)
	) name23241 (
		\m6_data_i[23]_pad ,
		_w8743_,
		_w8744_,
		_w25142_
	);
	LUT4 #(
		.INIT('hcedf)
	) name23242 (
		_w8738_,
		_w8741_,
		_w25141_,
		_w25142_,
		_w25143_
	);
	LUT3 #(
		.INIT('h2a)
	) name23243 (
		\m1_data_i[23]_pad ,
		_w8743_,
		_w8744_,
		_w25144_
	);
	LUT3 #(
		.INIT('h80)
	) name23244 (
		\m2_data_i[23]_pad ,
		_w8743_,
		_w8744_,
		_w25145_
	);
	LUT4 #(
		.INIT('h3b7f)
	) name23245 (
		_w8738_,
		_w8741_,
		_w25144_,
		_w25145_,
		_w25146_
	);
	LUT4 #(
		.INIT('h7fff)
	) name23246 (
		_w25137_,
		_w25140_,
		_w25143_,
		_w25146_,
		_w25147_
	);
	LUT3 #(
		.INIT('h2a)
	) name23247 (
		\m3_data_i[24]_pad ,
		_w8743_,
		_w8744_,
		_w25148_
	);
	LUT3 #(
		.INIT('h80)
	) name23248 (
		\m4_data_i[24]_pad ,
		_w8743_,
		_w8744_,
		_w25149_
	);
	LUT4 #(
		.INIT('h9dbf)
	) name23249 (
		_w8738_,
		_w8741_,
		_w25148_,
		_w25149_,
		_w25150_
	);
	LUT3 #(
		.INIT('h80)
	) name23250 (
		\m6_data_i[24]_pad ,
		_w8743_,
		_w8744_,
		_w25151_
	);
	LUT3 #(
		.INIT('h80)
	) name23251 (
		\m2_data_i[24]_pad ,
		_w8743_,
		_w8744_,
		_w25152_
	);
	LUT4 #(
		.INIT('habef)
	) name23252 (
		_w8738_,
		_w8741_,
		_w25151_,
		_w25152_,
		_w25153_
	);
	LUT3 #(
		.INIT('h2a)
	) name23253 (
		\m5_data_i[24]_pad ,
		_w8743_,
		_w8744_,
		_w25154_
	);
	LUT3 #(
		.INIT('h2a)
	) name23254 (
		\m1_data_i[24]_pad ,
		_w8743_,
		_w8744_,
		_w25155_
	);
	LUT4 #(
		.INIT('h57df)
	) name23255 (
		_w8738_,
		_w8741_,
		_w25154_,
		_w25155_,
		_w25156_
	);
	LUT3 #(
		.INIT('h80)
	) name23256 (
		\m0_data_i[24]_pad ,
		_w8743_,
		_w8744_,
		_w25157_
	);
	LUT3 #(
		.INIT('h2a)
	) name23257 (
		\m7_data_i[24]_pad ,
		_w8743_,
		_w8744_,
		_w25158_
	);
	LUT4 #(
		.INIT('h6e7f)
	) name23258 (
		_w8738_,
		_w8741_,
		_w25157_,
		_w25158_,
		_w25159_
	);
	LUT4 #(
		.INIT('h7fff)
	) name23259 (
		_w25150_,
		_w25153_,
		_w25156_,
		_w25159_,
		_w25160_
	);
	LUT3 #(
		.INIT('h2a)
	) name23260 (
		\m3_data_i[25]_pad ,
		_w8743_,
		_w8744_,
		_w25161_
	);
	LUT3 #(
		.INIT('h80)
	) name23261 (
		\m4_data_i[25]_pad ,
		_w8743_,
		_w8744_,
		_w25162_
	);
	LUT4 #(
		.INIT('h9dbf)
	) name23262 (
		_w8738_,
		_w8741_,
		_w25161_,
		_w25162_,
		_w25163_
	);
	LUT3 #(
		.INIT('h80)
	) name23263 (
		\m6_data_i[25]_pad ,
		_w8743_,
		_w8744_,
		_w25164_
	);
	LUT3 #(
		.INIT('h80)
	) name23264 (
		\m2_data_i[25]_pad ,
		_w8743_,
		_w8744_,
		_w25165_
	);
	LUT4 #(
		.INIT('habef)
	) name23265 (
		_w8738_,
		_w8741_,
		_w25164_,
		_w25165_,
		_w25166_
	);
	LUT3 #(
		.INIT('h2a)
	) name23266 (
		\m5_data_i[25]_pad ,
		_w8743_,
		_w8744_,
		_w25167_
	);
	LUT3 #(
		.INIT('h2a)
	) name23267 (
		\m1_data_i[25]_pad ,
		_w8743_,
		_w8744_,
		_w25168_
	);
	LUT4 #(
		.INIT('h57df)
	) name23268 (
		_w8738_,
		_w8741_,
		_w25167_,
		_w25168_,
		_w25169_
	);
	LUT3 #(
		.INIT('h80)
	) name23269 (
		\m0_data_i[25]_pad ,
		_w8743_,
		_w8744_,
		_w25170_
	);
	LUT3 #(
		.INIT('h2a)
	) name23270 (
		\m7_data_i[25]_pad ,
		_w8743_,
		_w8744_,
		_w25171_
	);
	LUT4 #(
		.INIT('h6e7f)
	) name23271 (
		_w8738_,
		_w8741_,
		_w25170_,
		_w25171_,
		_w25172_
	);
	LUT4 #(
		.INIT('h7fff)
	) name23272 (
		_w25163_,
		_w25166_,
		_w25169_,
		_w25172_,
		_w25173_
	);
	LUT3 #(
		.INIT('h2a)
	) name23273 (
		\m3_data_i[26]_pad ,
		_w8743_,
		_w8744_,
		_w25174_
	);
	LUT3 #(
		.INIT('h80)
	) name23274 (
		\m4_data_i[26]_pad ,
		_w8743_,
		_w8744_,
		_w25175_
	);
	LUT4 #(
		.INIT('h9dbf)
	) name23275 (
		_w8738_,
		_w8741_,
		_w25174_,
		_w25175_,
		_w25176_
	);
	LUT3 #(
		.INIT('h80)
	) name23276 (
		\m6_data_i[26]_pad ,
		_w8743_,
		_w8744_,
		_w25177_
	);
	LUT3 #(
		.INIT('h80)
	) name23277 (
		\m2_data_i[26]_pad ,
		_w8743_,
		_w8744_,
		_w25178_
	);
	LUT4 #(
		.INIT('habef)
	) name23278 (
		_w8738_,
		_w8741_,
		_w25177_,
		_w25178_,
		_w25179_
	);
	LUT3 #(
		.INIT('h2a)
	) name23279 (
		\m5_data_i[26]_pad ,
		_w8743_,
		_w8744_,
		_w25180_
	);
	LUT3 #(
		.INIT('h2a)
	) name23280 (
		\m1_data_i[26]_pad ,
		_w8743_,
		_w8744_,
		_w25181_
	);
	LUT4 #(
		.INIT('h57df)
	) name23281 (
		_w8738_,
		_w8741_,
		_w25180_,
		_w25181_,
		_w25182_
	);
	LUT3 #(
		.INIT('h80)
	) name23282 (
		\m0_data_i[26]_pad ,
		_w8743_,
		_w8744_,
		_w25183_
	);
	LUT3 #(
		.INIT('h2a)
	) name23283 (
		\m7_data_i[26]_pad ,
		_w8743_,
		_w8744_,
		_w25184_
	);
	LUT4 #(
		.INIT('h6e7f)
	) name23284 (
		_w8738_,
		_w8741_,
		_w25183_,
		_w25184_,
		_w25185_
	);
	LUT4 #(
		.INIT('h7fff)
	) name23285 (
		_w25176_,
		_w25179_,
		_w25182_,
		_w25185_,
		_w25186_
	);
	LUT3 #(
		.INIT('h2a)
	) name23286 (
		\m3_data_i[27]_pad ,
		_w8743_,
		_w8744_,
		_w25187_
	);
	LUT3 #(
		.INIT('h80)
	) name23287 (
		\m4_data_i[27]_pad ,
		_w8743_,
		_w8744_,
		_w25188_
	);
	LUT4 #(
		.INIT('h9dbf)
	) name23288 (
		_w8738_,
		_w8741_,
		_w25187_,
		_w25188_,
		_w25189_
	);
	LUT3 #(
		.INIT('h80)
	) name23289 (
		\m6_data_i[27]_pad ,
		_w8743_,
		_w8744_,
		_w25190_
	);
	LUT3 #(
		.INIT('h80)
	) name23290 (
		\m2_data_i[27]_pad ,
		_w8743_,
		_w8744_,
		_w25191_
	);
	LUT4 #(
		.INIT('habef)
	) name23291 (
		_w8738_,
		_w8741_,
		_w25190_,
		_w25191_,
		_w25192_
	);
	LUT3 #(
		.INIT('h2a)
	) name23292 (
		\m5_data_i[27]_pad ,
		_w8743_,
		_w8744_,
		_w25193_
	);
	LUT3 #(
		.INIT('h2a)
	) name23293 (
		\m1_data_i[27]_pad ,
		_w8743_,
		_w8744_,
		_w25194_
	);
	LUT4 #(
		.INIT('h57df)
	) name23294 (
		_w8738_,
		_w8741_,
		_w25193_,
		_w25194_,
		_w25195_
	);
	LUT3 #(
		.INIT('h80)
	) name23295 (
		\m0_data_i[27]_pad ,
		_w8743_,
		_w8744_,
		_w25196_
	);
	LUT3 #(
		.INIT('h2a)
	) name23296 (
		\m7_data_i[27]_pad ,
		_w8743_,
		_w8744_,
		_w25197_
	);
	LUT4 #(
		.INIT('h6e7f)
	) name23297 (
		_w8738_,
		_w8741_,
		_w25196_,
		_w25197_,
		_w25198_
	);
	LUT4 #(
		.INIT('h7fff)
	) name23298 (
		_w25189_,
		_w25192_,
		_w25195_,
		_w25198_,
		_w25199_
	);
	LUT3 #(
		.INIT('h2a)
	) name23299 (
		\m1_data_i[28]_pad ,
		_w8743_,
		_w8744_,
		_w25200_
	);
	LUT3 #(
		.INIT('h80)
	) name23300 (
		\m2_data_i[28]_pad ,
		_w8743_,
		_w8744_,
		_w25201_
	);
	LUT4 #(
		.INIT('h3b7f)
	) name23301 (
		_w8738_,
		_w8741_,
		_w25200_,
		_w25201_,
		_w25202_
	);
	LUT3 #(
		.INIT('h80)
	) name23302 (
		\m0_data_i[28]_pad ,
		_w8743_,
		_w8744_,
		_w25203_
	);
	LUT3 #(
		.INIT('h80)
	) name23303 (
		\m4_data_i[28]_pad ,
		_w8743_,
		_w8744_,
		_w25204_
	);
	LUT4 #(
		.INIT('h5d7f)
	) name23304 (
		_w8738_,
		_w8741_,
		_w25203_,
		_w25204_,
		_w25205_
	);
	LUT3 #(
		.INIT('h2a)
	) name23305 (
		\m7_data_i[28]_pad ,
		_w8743_,
		_w8744_,
		_w25206_
	);
	LUT3 #(
		.INIT('h2a)
	) name23306 (
		\m3_data_i[28]_pad ,
		_w8743_,
		_w8744_,
		_w25207_
	);
	LUT4 #(
		.INIT('habef)
	) name23307 (
		_w8738_,
		_w8741_,
		_w25206_,
		_w25207_,
		_w25208_
	);
	LUT3 #(
		.INIT('h80)
	) name23308 (
		\m6_data_i[28]_pad ,
		_w8743_,
		_w8744_,
		_w25209_
	);
	LUT3 #(
		.INIT('h2a)
	) name23309 (
		\m5_data_i[28]_pad ,
		_w8743_,
		_w8744_,
		_w25210_
	);
	LUT4 #(
		.INIT('hcdef)
	) name23310 (
		_w8738_,
		_w8741_,
		_w25209_,
		_w25210_,
		_w25211_
	);
	LUT4 #(
		.INIT('h7fff)
	) name23311 (
		_w25202_,
		_w25205_,
		_w25208_,
		_w25211_,
		_w25212_
	);
	LUT3 #(
		.INIT('h2a)
	) name23312 (
		\m3_data_i[29]_pad ,
		_w8743_,
		_w8744_,
		_w25213_
	);
	LUT3 #(
		.INIT('h80)
	) name23313 (
		\m4_data_i[29]_pad ,
		_w8743_,
		_w8744_,
		_w25214_
	);
	LUT4 #(
		.INIT('h9dbf)
	) name23314 (
		_w8738_,
		_w8741_,
		_w25213_,
		_w25214_,
		_w25215_
	);
	LUT3 #(
		.INIT('h80)
	) name23315 (
		\m6_data_i[29]_pad ,
		_w8743_,
		_w8744_,
		_w25216_
	);
	LUT3 #(
		.INIT('h2a)
	) name23316 (
		\m7_data_i[29]_pad ,
		_w8743_,
		_w8744_,
		_w25217_
	);
	LUT3 #(
		.INIT('h57)
	) name23317 (
		_w8756_,
		_w25216_,
		_w25217_,
		_w25218_
	);
	LUT3 #(
		.INIT('h2a)
	) name23318 (
		\m5_data_i[29]_pad ,
		_w8743_,
		_w8744_,
		_w25219_
	);
	LUT3 #(
		.INIT('h80)
	) name23319 (
		\m0_data_i[29]_pad ,
		_w8743_,
		_w8744_,
		_w25220_
	);
	LUT4 #(
		.INIT('h57df)
	) name23320 (
		_w8738_,
		_w8741_,
		_w25219_,
		_w25220_,
		_w25221_
	);
	LUT3 #(
		.INIT('h2a)
	) name23321 (
		\m1_data_i[29]_pad ,
		_w8743_,
		_w8744_,
		_w25222_
	);
	LUT3 #(
		.INIT('h80)
	) name23322 (
		\m2_data_i[29]_pad ,
		_w8743_,
		_w8744_,
		_w25223_
	);
	LUT4 #(
		.INIT('h3b7f)
	) name23323 (
		_w8738_,
		_w8741_,
		_w25222_,
		_w25223_,
		_w25224_
	);
	LUT4 #(
		.INIT('h7fff)
	) name23324 (
		_w25215_,
		_w25218_,
		_w25221_,
		_w25224_,
		_w25225_
	);
	LUT3 #(
		.INIT('h2a)
	) name23325 (
		\m1_data_i[2]_pad ,
		_w8743_,
		_w8744_,
		_w25226_
	);
	LUT3 #(
		.INIT('h80)
	) name23326 (
		\m2_data_i[2]_pad ,
		_w8743_,
		_w8744_,
		_w25227_
	);
	LUT4 #(
		.INIT('h3b7f)
	) name23327 (
		_w8738_,
		_w8741_,
		_w25226_,
		_w25227_,
		_w25228_
	);
	LUT3 #(
		.INIT('h80)
	) name23328 (
		\m0_data_i[2]_pad ,
		_w8743_,
		_w8744_,
		_w25229_
	);
	LUT3 #(
		.INIT('h80)
	) name23329 (
		\m4_data_i[2]_pad ,
		_w8743_,
		_w8744_,
		_w25230_
	);
	LUT4 #(
		.INIT('h5d7f)
	) name23330 (
		_w8738_,
		_w8741_,
		_w25229_,
		_w25230_,
		_w25231_
	);
	LUT3 #(
		.INIT('h2a)
	) name23331 (
		\m7_data_i[2]_pad ,
		_w8743_,
		_w8744_,
		_w25232_
	);
	LUT3 #(
		.INIT('h2a)
	) name23332 (
		\m3_data_i[2]_pad ,
		_w8743_,
		_w8744_,
		_w25233_
	);
	LUT4 #(
		.INIT('habef)
	) name23333 (
		_w8738_,
		_w8741_,
		_w25232_,
		_w25233_,
		_w25234_
	);
	LUT3 #(
		.INIT('h80)
	) name23334 (
		\m6_data_i[2]_pad ,
		_w8743_,
		_w8744_,
		_w25235_
	);
	LUT3 #(
		.INIT('h2a)
	) name23335 (
		\m5_data_i[2]_pad ,
		_w8743_,
		_w8744_,
		_w25236_
	);
	LUT4 #(
		.INIT('hcdef)
	) name23336 (
		_w8738_,
		_w8741_,
		_w25235_,
		_w25236_,
		_w25237_
	);
	LUT4 #(
		.INIT('h7fff)
	) name23337 (
		_w25228_,
		_w25231_,
		_w25234_,
		_w25237_,
		_w25238_
	);
	LUT3 #(
		.INIT('h2a)
	) name23338 (
		\m3_data_i[30]_pad ,
		_w8743_,
		_w8744_,
		_w25239_
	);
	LUT3 #(
		.INIT('h80)
	) name23339 (
		\m4_data_i[30]_pad ,
		_w8743_,
		_w8744_,
		_w25240_
	);
	LUT4 #(
		.INIT('h9dbf)
	) name23340 (
		_w8738_,
		_w8741_,
		_w25239_,
		_w25240_,
		_w25241_
	);
	LUT3 #(
		.INIT('h80)
	) name23341 (
		\m6_data_i[30]_pad ,
		_w8743_,
		_w8744_,
		_w25242_
	);
	LUT3 #(
		.INIT('h80)
	) name23342 (
		\m2_data_i[30]_pad ,
		_w8743_,
		_w8744_,
		_w25243_
	);
	LUT4 #(
		.INIT('habef)
	) name23343 (
		_w8738_,
		_w8741_,
		_w25242_,
		_w25243_,
		_w25244_
	);
	LUT3 #(
		.INIT('h2a)
	) name23344 (
		\m5_data_i[30]_pad ,
		_w8743_,
		_w8744_,
		_w25245_
	);
	LUT3 #(
		.INIT('h2a)
	) name23345 (
		\m1_data_i[30]_pad ,
		_w8743_,
		_w8744_,
		_w25246_
	);
	LUT4 #(
		.INIT('h57df)
	) name23346 (
		_w8738_,
		_w8741_,
		_w25245_,
		_w25246_,
		_w25247_
	);
	LUT3 #(
		.INIT('h80)
	) name23347 (
		\m0_data_i[30]_pad ,
		_w8743_,
		_w8744_,
		_w25248_
	);
	LUT3 #(
		.INIT('h2a)
	) name23348 (
		\m7_data_i[30]_pad ,
		_w8743_,
		_w8744_,
		_w25249_
	);
	LUT4 #(
		.INIT('h6e7f)
	) name23349 (
		_w8738_,
		_w8741_,
		_w25248_,
		_w25249_,
		_w25250_
	);
	LUT4 #(
		.INIT('h7fff)
	) name23350 (
		_w25241_,
		_w25244_,
		_w25247_,
		_w25250_,
		_w25251_
	);
	LUT3 #(
		.INIT('h80)
	) name23351 (
		\m0_data_i[31]_pad ,
		_w8743_,
		_w8744_,
		_w25252_
	);
	LUT3 #(
		.INIT('h2a)
	) name23352 (
		\m7_data_i[31]_pad ,
		_w8743_,
		_w8744_,
		_w25253_
	);
	LUT4 #(
		.INIT('h6e7f)
	) name23353 (
		_w8738_,
		_w8741_,
		_w25252_,
		_w25253_,
		_w25254_
	);
	LUT3 #(
		.INIT('h2a)
	) name23354 (
		\m1_data_i[31]_pad ,
		_w8743_,
		_w8744_,
		_w25255_
	);
	LUT3 #(
		.INIT('h80)
	) name23355 (
		\m4_data_i[31]_pad ,
		_w8743_,
		_w8744_,
		_w25256_
	);
	LUT4 #(
		.INIT('h5d7f)
	) name23356 (
		_w8738_,
		_w8741_,
		_w25255_,
		_w25256_,
		_w25257_
	);
	LUT3 #(
		.INIT('h80)
	) name23357 (
		\m2_data_i[31]_pad ,
		_w8743_,
		_w8744_,
		_w25258_
	);
	LUT3 #(
		.INIT('h2a)
	) name23358 (
		\m3_data_i[31]_pad ,
		_w8743_,
		_w8744_,
		_w25259_
	);
	LUT3 #(
		.INIT('h57)
	) name23359 (
		_w8750_,
		_w25258_,
		_w25259_,
		_w25260_
	);
	LUT3 #(
		.INIT('h80)
	) name23360 (
		\m6_data_i[31]_pad ,
		_w8743_,
		_w8744_,
		_w25261_
	);
	LUT3 #(
		.INIT('h2a)
	) name23361 (
		\m5_data_i[31]_pad ,
		_w8743_,
		_w8744_,
		_w25262_
	);
	LUT4 #(
		.INIT('hcdef)
	) name23362 (
		_w8738_,
		_w8741_,
		_w25261_,
		_w25262_,
		_w25263_
	);
	LUT4 #(
		.INIT('h7fff)
	) name23363 (
		_w25254_,
		_w25257_,
		_w25260_,
		_w25263_,
		_w25264_
	);
	LUT3 #(
		.INIT('h2a)
	) name23364 (
		\m1_data_i[3]_pad ,
		_w8743_,
		_w8744_,
		_w25265_
	);
	LUT3 #(
		.INIT('h80)
	) name23365 (
		\m2_data_i[3]_pad ,
		_w8743_,
		_w8744_,
		_w25266_
	);
	LUT4 #(
		.INIT('h3b7f)
	) name23366 (
		_w8738_,
		_w8741_,
		_w25265_,
		_w25266_,
		_w25267_
	);
	LUT3 #(
		.INIT('h80)
	) name23367 (
		\m0_data_i[3]_pad ,
		_w8743_,
		_w8744_,
		_w25268_
	);
	LUT3 #(
		.INIT('h80)
	) name23368 (
		\m4_data_i[3]_pad ,
		_w8743_,
		_w8744_,
		_w25269_
	);
	LUT4 #(
		.INIT('h5d7f)
	) name23369 (
		_w8738_,
		_w8741_,
		_w25268_,
		_w25269_,
		_w25270_
	);
	LUT3 #(
		.INIT('h2a)
	) name23370 (
		\m7_data_i[3]_pad ,
		_w8743_,
		_w8744_,
		_w25271_
	);
	LUT3 #(
		.INIT('h2a)
	) name23371 (
		\m3_data_i[3]_pad ,
		_w8743_,
		_w8744_,
		_w25272_
	);
	LUT4 #(
		.INIT('habef)
	) name23372 (
		_w8738_,
		_w8741_,
		_w25271_,
		_w25272_,
		_w25273_
	);
	LUT3 #(
		.INIT('h80)
	) name23373 (
		\m6_data_i[3]_pad ,
		_w8743_,
		_w8744_,
		_w25274_
	);
	LUT3 #(
		.INIT('h2a)
	) name23374 (
		\m5_data_i[3]_pad ,
		_w8743_,
		_w8744_,
		_w25275_
	);
	LUT4 #(
		.INIT('hcdef)
	) name23375 (
		_w8738_,
		_w8741_,
		_w25274_,
		_w25275_,
		_w25276_
	);
	LUT4 #(
		.INIT('h7fff)
	) name23376 (
		_w25267_,
		_w25270_,
		_w25273_,
		_w25276_,
		_w25277_
	);
	LUT3 #(
		.INIT('h80)
	) name23377 (
		\m0_data_i[4]_pad ,
		_w8743_,
		_w8744_,
		_w25278_
	);
	LUT3 #(
		.INIT('h2a)
	) name23378 (
		\m7_data_i[4]_pad ,
		_w8743_,
		_w8744_,
		_w25279_
	);
	LUT4 #(
		.INIT('h6e7f)
	) name23379 (
		_w8738_,
		_w8741_,
		_w25278_,
		_w25279_,
		_w25280_
	);
	LUT3 #(
		.INIT('h80)
	) name23380 (
		\m6_data_i[4]_pad ,
		_w8743_,
		_w8744_,
		_w25281_
	);
	LUT3 #(
		.INIT('h80)
	) name23381 (
		\m2_data_i[4]_pad ,
		_w8743_,
		_w8744_,
		_w25282_
	);
	LUT4 #(
		.INIT('habef)
	) name23382 (
		_w8738_,
		_w8741_,
		_w25281_,
		_w25282_,
		_w25283_
	);
	LUT3 #(
		.INIT('h2a)
	) name23383 (
		\m5_data_i[4]_pad ,
		_w8743_,
		_w8744_,
		_w25284_
	);
	LUT3 #(
		.INIT('h2a)
	) name23384 (
		\m1_data_i[4]_pad ,
		_w8743_,
		_w8744_,
		_w25285_
	);
	LUT4 #(
		.INIT('h57df)
	) name23385 (
		_w8738_,
		_w8741_,
		_w25284_,
		_w25285_,
		_w25286_
	);
	LUT3 #(
		.INIT('h2a)
	) name23386 (
		\m3_data_i[4]_pad ,
		_w8743_,
		_w8744_,
		_w25287_
	);
	LUT3 #(
		.INIT('h80)
	) name23387 (
		\m4_data_i[4]_pad ,
		_w8743_,
		_w8744_,
		_w25288_
	);
	LUT4 #(
		.INIT('h9dbf)
	) name23388 (
		_w8738_,
		_w8741_,
		_w25287_,
		_w25288_,
		_w25289_
	);
	LUT4 #(
		.INIT('h7fff)
	) name23389 (
		_w25280_,
		_w25283_,
		_w25286_,
		_w25289_,
		_w25290_
	);
	LUT3 #(
		.INIT('h2a)
	) name23390 (
		\m1_data_i[5]_pad ,
		_w8743_,
		_w8744_,
		_w25291_
	);
	LUT3 #(
		.INIT('h80)
	) name23391 (
		\m2_data_i[5]_pad ,
		_w8743_,
		_w8744_,
		_w25292_
	);
	LUT4 #(
		.INIT('h3b7f)
	) name23392 (
		_w8738_,
		_w8741_,
		_w25291_,
		_w25292_,
		_w25293_
	);
	LUT3 #(
		.INIT('h80)
	) name23393 (
		\m0_data_i[5]_pad ,
		_w8743_,
		_w8744_,
		_w25294_
	);
	LUT3 #(
		.INIT('h80)
	) name23394 (
		\m4_data_i[5]_pad ,
		_w8743_,
		_w8744_,
		_w25295_
	);
	LUT4 #(
		.INIT('h5d7f)
	) name23395 (
		_w8738_,
		_w8741_,
		_w25294_,
		_w25295_,
		_w25296_
	);
	LUT3 #(
		.INIT('h2a)
	) name23396 (
		\m7_data_i[5]_pad ,
		_w8743_,
		_w8744_,
		_w25297_
	);
	LUT3 #(
		.INIT('h2a)
	) name23397 (
		\m3_data_i[5]_pad ,
		_w8743_,
		_w8744_,
		_w25298_
	);
	LUT4 #(
		.INIT('habef)
	) name23398 (
		_w8738_,
		_w8741_,
		_w25297_,
		_w25298_,
		_w25299_
	);
	LUT3 #(
		.INIT('h80)
	) name23399 (
		\m6_data_i[5]_pad ,
		_w8743_,
		_w8744_,
		_w25300_
	);
	LUT3 #(
		.INIT('h2a)
	) name23400 (
		\m5_data_i[5]_pad ,
		_w8743_,
		_w8744_,
		_w25301_
	);
	LUT4 #(
		.INIT('hcdef)
	) name23401 (
		_w8738_,
		_w8741_,
		_w25300_,
		_w25301_,
		_w25302_
	);
	LUT4 #(
		.INIT('h7fff)
	) name23402 (
		_w25293_,
		_w25296_,
		_w25299_,
		_w25302_,
		_w25303_
	);
	LUT3 #(
		.INIT('h80)
	) name23403 (
		\m6_data_i[6]_pad ,
		_w8743_,
		_w8744_,
		_w25304_
	);
	LUT3 #(
		.INIT('h2a)
	) name23404 (
		\m5_data_i[6]_pad ,
		_w8743_,
		_w8744_,
		_w25305_
	);
	LUT4 #(
		.INIT('hcdef)
	) name23405 (
		_w8738_,
		_w8741_,
		_w25304_,
		_w25305_,
		_w25306_
	);
	LUT3 #(
		.INIT('h80)
	) name23406 (
		\m0_data_i[6]_pad ,
		_w8743_,
		_w8744_,
		_w25307_
	);
	LUT3 #(
		.INIT('h80)
	) name23407 (
		\m2_data_i[6]_pad ,
		_w8743_,
		_w8744_,
		_w25308_
	);
	LUT4 #(
		.INIT('h3b7f)
	) name23408 (
		_w8738_,
		_w8741_,
		_w25307_,
		_w25308_,
		_w25309_
	);
	LUT3 #(
		.INIT('h2a)
	) name23409 (
		\m7_data_i[6]_pad ,
		_w8743_,
		_w8744_,
		_w25310_
	);
	LUT3 #(
		.INIT('h2a)
	) name23410 (
		\m1_data_i[6]_pad ,
		_w8743_,
		_w8744_,
		_w25311_
	);
	LUT4 #(
		.INIT('h67ef)
	) name23411 (
		_w8738_,
		_w8741_,
		_w25310_,
		_w25311_,
		_w25312_
	);
	LUT3 #(
		.INIT('h2a)
	) name23412 (
		\m3_data_i[6]_pad ,
		_w8743_,
		_w8744_,
		_w25313_
	);
	LUT3 #(
		.INIT('h80)
	) name23413 (
		\m4_data_i[6]_pad ,
		_w8743_,
		_w8744_,
		_w25314_
	);
	LUT4 #(
		.INIT('h9dbf)
	) name23414 (
		_w8738_,
		_w8741_,
		_w25313_,
		_w25314_,
		_w25315_
	);
	LUT4 #(
		.INIT('h7fff)
	) name23415 (
		_w25306_,
		_w25309_,
		_w25312_,
		_w25315_,
		_w25316_
	);
	LUT3 #(
		.INIT('h2a)
	) name23416 (
		\m3_data_i[7]_pad ,
		_w8743_,
		_w8744_,
		_w25317_
	);
	LUT3 #(
		.INIT('h80)
	) name23417 (
		\m4_data_i[7]_pad ,
		_w8743_,
		_w8744_,
		_w25318_
	);
	LUT4 #(
		.INIT('h9dbf)
	) name23418 (
		_w8738_,
		_w8741_,
		_w25317_,
		_w25318_,
		_w25319_
	);
	LUT3 #(
		.INIT('h80)
	) name23419 (
		\m6_data_i[7]_pad ,
		_w8743_,
		_w8744_,
		_w25320_
	);
	LUT3 #(
		.INIT('h2a)
	) name23420 (
		\m7_data_i[7]_pad ,
		_w8743_,
		_w8744_,
		_w25321_
	);
	LUT3 #(
		.INIT('h57)
	) name23421 (
		_w8756_,
		_w25320_,
		_w25321_,
		_w25322_
	);
	LUT3 #(
		.INIT('h2a)
	) name23422 (
		\m5_data_i[7]_pad ,
		_w8743_,
		_w8744_,
		_w25323_
	);
	LUT3 #(
		.INIT('h80)
	) name23423 (
		\m0_data_i[7]_pad ,
		_w8743_,
		_w8744_,
		_w25324_
	);
	LUT4 #(
		.INIT('h57df)
	) name23424 (
		_w8738_,
		_w8741_,
		_w25323_,
		_w25324_,
		_w25325_
	);
	LUT3 #(
		.INIT('h2a)
	) name23425 (
		\m1_data_i[7]_pad ,
		_w8743_,
		_w8744_,
		_w25326_
	);
	LUT3 #(
		.INIT('h80)
	) name23426 (
		\m2_data_i[7]_pad ,
		_w8743_,
		_w8744_,
		_w25327_
	);
	LUT4 #(
		.INIT('h3b7f)
	) name23427 (
		_w8738_,
		_w8741_,
		_w25326_,
		_w25327_,
		_w25328_
	);
	LUT4 #(
		.INIT('h7fff)
	) name23428 (
		_w25319_,
		_w25322_,
		_w25325_,
		_w25328_,
		_w25329_
	);
	LUT3 #(
		.INIT('h2a)
	) name23429 (
		\m1_data_i[8]_pad ,
		_w8743_,
		_w8744_,
		_w25330_
	);
	LUT3 #(
		.INIT('h80)
	) name23430 (
		\m2_data_i[8]_pad ,
		_w8743_,
		_w8744_,
		_w25331_
	);
	LUT4 #(
		.INIT('h3b7f)
	) name23431 (
		_w8738_,
		_w8741_,
		_w25330_,
		_w25331_,
		_w25332_
	);
	LUT3 #(
		.INIT('h80)
	) name23432 (
		\m0_data_i[8]_pad ,
		_w8743_,
		_w8744_,
		_w25333_
	);
	LUT3 #(
		.INIT('h80)
	) name23433 (
		\m4_data_i[8]_pad ,
		_w8743_,
		_w8744_,
		_w25334_
	);
	LUT4 #(
		.INIT('h5d7f)
	) name23434 (
		_w8738_,
		_w8741_,
		_w25333_,
		_w25334_,
		_w25335_
	);
	LUT3 #(
		.INIT('h2a)
	) name23435 (
		\m7_data_i[8]_pad ,
		_w8743_,
		_w8744_,
		_w25336_
	);
	LUT3 #(
		.INIT('h2a)
	) name23436 (
		\m3_data_i[8]_pad ,
		_w8743_,
		_w8744_,
		_w25337_
	);
	LUT4 #(
		.INIT('habef)
	) name23437 (
		_w8738_,
		_w8741_,
		_w25336_,
		_w25337_,
		_w25338_
	);
	LUT3 #(
		.INIT('h80)
	) name23438 (
		\m6_data_i[8]_pad ,
		_w8743_,
		_w8744_,
		_w25339_
	);
	LUT3 #(
		.INIT('h2a)
	) name23439 (
		\m5_data_i[8]_pad ,
		_w8743_,
		_w8744_,
		_w25340_
	);
	LUT4 #(
		.INIT('hcdef)
	) name23440 (
		_w8738_,
		_w8741_,
		_w25339_,
		_w25340_,
		_w25341_
	);
	LUT4 #(
		.INIT('h7fff)
	) name23441 (
		_w25332_,
		_w25335_,
		_w25338_,
		_w25341_,
		_w25342_
	);
	LUT3 #(
		.INIT('h2a)
	) name23442 (
		\m1_data_i[9]_pad ,
		_w8743_,
		_w8744_,
		_w25343_
	);
	LUT3 #(
		.INIT('h80)
	) name23443 (
		\m2_data_i[9]_pad ,
		_w8743_,
		_w8744_,
		_w25344_
	);
	LUT4 #(
		.INIT('h3b7f)
	) name23444 (
		_w8738_,
		_w8741_,
		_w25343_,
		_w25344_,
		_w25345_
	);
	LUT3 #(
		.INIT('h80)
	) name23445 (
		\m0_data_i[9]_pad ,
		_w8743_,
		_w8744_,
		_w25346_
	);
	LUT3 #(
		.INIT('h80)
	) name23446 (
		\m4_data_i[9]_pad ,
		_w8743_,
		_w8744_,
		_w25347_
	);
	LUT4 #(
		.INIT('h5d7f)
	) name23447 (
		_w8738_,
		_w8741_,
		_w25346_,
		_w25347_,
		_w25348_
	);
	LUT3 #(
		.INIT('h2a)
	) name23448 (
		\m7_data_i[9]_pad ,
		_w8743_,
		_w8744_,
		_w25349_
	);
	LUT3 #(
		.INIT('h2a)
	) name23449 (
		\m3_data_i[9]_pad ,
		_w8743_,
		_w8744_,
		_w25350_
	);
	LUT4 #(
		.INIT('habef)
	) name23450 (
		_w8738_,
		_w8741_,
		_w25349_,
		_w25350_,
		_w25351_
	);
	LUT3 #(
		.INIT('h80)
	) name23451 (
		\m6_data_i[9]_pad ,
		_w8743_,
		_w8744_,
		_w25352_
	);
	LUT3 #(
		.INIT('h2a)
	) name23452 (
		\m5_data_i[9]_pad ,
		_w8743_,
		_w8744_,
		_w25353_
	);
	LUT4 #(
		.INIT('hcdef)
	) name23453 (
		_w8738_,
		_w8741_,
		_w25352_,
		_w25353_,
		_w25354_
	);
	LUT4 #(
		.INIT('h7fff)
	) name23454 (
		_w25345_,
		_w25348_,
		_w25351_,
		_w25354_,
		_w25355_
	);
	LUT3 #(
		.INIT('h2a)
	) name23455 (
		\m3_sel_i[0]_pad ,
		_w8743_,
		_w8744_,
		_w25356_
	);
	LUT3 #(
		.INIT('h80)
	) name23456 (
		\m4_sel_i[0]_pad ,
		_w8743_,
		_w8744_,
		_w25357_
	);
	LUT4 #(
		.INIT('h9dbf)
	) name23457 (
		_w8738_,
		_w8741_,
		_w25356_,
		_w25357_,
		_w25358_
	);
	LUT3 #(
		.INIT('h80)
	) name23458 (
		\m6_sel_i[0]_pad ,
		_w8743_,
		_w8744_,
		_w25359_
	);
	LUT3 #(
		.INIT('h80)
	) name23459 (
		\m2_sel_i[0]_pad ,
		_w8743_,
		_w8744_,
		_w25360_
	);
	LUT4 #(
		.INIT('habef)
	) name23460 (
		_w8738_,
		_w8741_,
		_w25359_,
		_w25360_,
		_w25361_
	);
	LUT3 #(
		.INIT('h2a)
	) name23461 (
		\m5_sel_i[0]_pad ,
		_w8743_,
		_w8744_,
		_w25362_
	);
	LUT3 #(
		.INIT('h2a)
	) name23462 (
		\m1_sel_i[0]_pad ,
		_w8743_,
		_w8744_,
		_w25363_
	);
	LUT4 #(
		.INIT('h57df)
	) name23463 (
		_w8738_,
		_w8741_,
		_w25362_,
		_w25363_,
		_w25364_
	);
	LUT3 #(
		.INIT('h80)
	) name23464 (
		\m0_sel_i[0]_pad ,
		_w8743_,
		_w8744_,
		_w25365_
	);
	LUT3 #(
		.INIT('h2a)
	) name23465 (
		\m7_sel_i[0]_pad ,
		_w8743_,
		_w8744_,
		_w25366_
	);
	LUT4 #(
		.INIT('h6e7f)
	) name23466 (
		_w8738_,
		_w8741_,
		_w25365_,
		_w25366_,
		_w25367_
	);
	LUT4 #(
		.INIT('h7fff)
	) name23467 (
		_w25358_,
		_w25361_,
		_w25364_,
		_w25367_,
		_w25368_
	);
	LUT3 #(
		.INIT('h2a)
	) name23468 (
		\m1_sel_i[1]_pad ,
		_w8743_,
		_w8744_,
		_w25369_
	);
	LUT3 #(
		.INIT('h80)
	) name23469 (
		\m2_sel_i[1]_pad ,
		_w8743_,
		_w8744_,
		_w25370_
	);
	LUT4 #(
		.INIT('h3b7f)
	) name23470 (
		_w8738_,
		_w8741_,
		_w25369_,
		_w25370_,
		_w25371_
	);
	LUT3 #(
		.INIT('h80)
	) name23471 (
		\m0_sel_i[1]_pad ,
		_w8743_,
		_w8744_,
		_w25372_
	);
	LUT3 #(
		.INIT('h80)
	) name23472 (
		\m4_sel_i[1]_pad ,
		_w8743_,
		_w8744_,
		_w25373_
	);
	LUT4 #(
		.INIT('h5d7f)
	) name23473 (
		_w8738_,
		_w8741_,
		_w25372_,
		_w25373_,
		_w25374_
	);
	LUT3 #(
		.INIT('h2a)
	) name23474 (
		\m7_sel_i[1]_pad ,
		_w8743_,
		_w8744_,
		_w25375_
	);
	LUT3 #(
		.INIT('h2a)
	) name23475 (
		\m3_sel_i[1]_pad ,
		_w8743_,
		_w8744_,
		_w25376_
	);
	LUT4 #(
		.INIT('habef)
	) name23476 (
		_w8738_,
		_w8741_,
		_w25375_,
		_w25376_,
		_w25377_
	);
	LUT3 #(
		.INIT('h80)
	) name23477 (
		\m6_sel_i[1]_pad ,
		_w8743_,
		_w8744_,
		_w25378_
	);
	LUT3 #(
		.INIT('h2a)
	) name23478 (
		\m5_sel_i[1]_pad ,
		_w8743_,
		_w8744_,
		_w25379_
	);
	LUT4 #(
		.INIT('hcdef)
	) name23479 (
		_w8738_,
		_w8741_,
		_w25378_,
		_w25379_,
		_w25380_
	);
	LUT4 #(
		.INIT('h7fff)
	) name23480 (
		_w25371_,
		_w25374_,
		_w25377_,
		_w25380_,
		_w25381_
	);
	LUT3 #(
		.INIT('h2a)
	) name23481 (
		\m1_sel_i[2]_pad ,
		_w8743_,
		_w8744_,
		_w25382_
	);
	LUT3 #(
		.INIT('h80)
	) name23482 (
		\m2_sel_i[2]_pad ,
		_w8743_,
		_w8744_,
		_w25383_
	);
	LUT4 #(
		.INIT('h3b7f)
	) name23483 (
		_w8738_,
		_w8741_,
		_w25382_,
		_w25383_,
		_w25384_
	);
	LUT3 #(
		.INIT('h80)
	) name23484 (
		\m0_sel_i[2]_pad ,
		_w8743_,
		_w8744_,
		_w25385_
	);
	LUT3 #(
		.INIT('h80)
	) name23485 (
		\m4_sel_i[2]_pad ,
		_w8743_,
		_w8744_,
		_w25386_
	);
	LUT4 #(
		.INIT('h5d7f)
	) name23486 (
		_w8738_,
		_w8741_,
		_w25385_,
		_w25386_,
		_w25387_
	);
	LUT3 #(
		.INIT('h2a)
	) name23487 (
		\m7_sel_i[2]_pad ,
		_w8743_,
		_w8744_,
		_w25388_
	);
	LUT3 #(
		.INIT('h2a)
	) name23488 (
		\m3_sel_i[2]_pad ,
		_w8743_,
		_w8744_,
		_w25389_
	);
	LUT4 #(
		.INIT('habef)
	) name23489 (
		_w8738_,
		_w8741_,
		_w25388_,
		_w25389_,
		_w25390_
	);
	LUT3 #(
		.INIT('h80)
	) name23490 (
		\m6_sel_i[2]_pad ,
		_w8743_,
		_w8744_,
		_w25391_
	);
	LUT3 #(
		.INIT('h2a)
	) name23491 (
		\m5_sel_i[2]_pad ,
		_w8743_,
		_w8744_,
		_w25392_
	);
	LUT4 #(
		.INIT('hcdef)
	) name23492 (
		_w8738_,
		_w8741_,
		_w25391_,
		_w25392_,
		_w25393_
	);
	LUT4 #(
		.INIT('h7fff)
	) name23493 (
		_w25384_,
		_w25387_,
		_w25390_,
		_w25393_,
		_w25394_
	);
	LUT3 #(
		.INIT('h80)
	) name23494 (
		\m0_sel_i[3]_pad ,
		_w8743_,
		_w8744_,
		_w25395_
	);
	LUT3 #(
		.INIT('h2a)
	) name23495 (
		\m7_sel_i[3]_pad ,
		_w8743_,
		_w8744_,
		_w25396_
	);
	LUT4 #(
		.INIT('h6e7f)
	) name23496 (
		_w8738_,
		_w8741_,
		_w25395_,
		_w25396_,
		_w25397_
	);
	LUT3 #(
		.INIT('h2a)
	) name23497 (
		\m3_sel_i[3]_pad ,
		_w8743_,
		_w8744_,
		_w25398_
	);
	LUT3 #(
		.INIT('h80)
	) name23498 (
		\m2_sel_i[3]_pad ,
		_w8743_,
		_w8744_,
		_w25399_
	);
	LUT3 #(
		.INIT('h57)
	) name23499 (
		_w8750_,
		_w25398_,
		_w25399_,
		_w25400_
	);
	LUT3 #(
		.INIT('h80)
	) name23500 (
		\m4_sel_i[3]_pad ,
		_w8743_,
		_w8744_,
		_w25401_
	);
	LUT3 #(
		.INIT('h2a)
	) name23501 (
		\m1_sel_i[3]_pad ,
		_w8743_,
		_w8744_,
		_w25402_
	);
	LUT4 #(
		.INIT('h57df)
	) name23502 (
		_w8738_,
		_w8741_,
		_w25401_,
		_w25402_,
		_w25403_
	);
	LUT3 #(
		.INIT('h80)
	) name23503 (
		\m6_sel_i[3]_pad ,
		_w8743_,
		_w8744_,
		_w25404_
	);
	LUT3 #(
		.INIT('h2a)
	) name23504 (
		\m5_sel_i[3]_pad ,
		_w8743_,
		_w8744_,
		_w25405_
	);
	LUT4 #(
		.INIT('hcdef)
	) name23505 (
		_w8738_,
		_w8741_,
		_w25404_,
		_w25405_,
		_w25406_
	);
	LUT4 #(
		.INIT('h7fff)
	) name23506 (
		_w25397_,
		_w25400_,
		_w25403_,
		_w25406_,
		_w25407_
	);
	LUT4 #(
		.INIT('h2a00)
	) name23507 (
		\m5_stb_i_pad ,
		_w8743_,
		_w8744_,
		_w9550_,
		_w25408_
	);
	LUT4 #(
		.INIT('h8000)
	) name23508 (
		\m4_stb_i_pad ,
		_w8743_,
		_w8744_,
		_w9363_,
		_w25409_
	);
	LUT3 #(
		.INIT('h57)
	) name23509 (
		_w8762_,
		_w25408_,
		_w25409_,
		_w25410_
	);
	LUT4 #(
		.INIT('h8000)
	) name23510 (
		\m2_stb_i_pad ,
		_w8743_,
		_w8744_,
		_w9474_,
		_w25411_
	);
	LUT4 #(
		.INIT('h8000)
	) name23511 (
		\m6_stb_i_pad ,
		_w8743_,
		_w8744_,
		_w9336_,
		_w25412_
	);
	LUT4 #(
		.INIT('haebf)
	) name23512 (
		_w8738_,
		_w8741_,
		_w25411_,
		_w25412_,
		_w25413_
	);
	LUT4 #(
		.INIT('h2a00)
	) name23513 (
		\m3_stb_i_pad ,
		_w8743_,
		_w8744_,
		_w9378_,
		_w25414_
	);
	LUT4 #(
		.INIT('h2a00)
	) name23514 (
		\m7_stb_i_pad ,
		_w8743_,
		_w8744_,
		_w9617_,
		_w25415_
	);
	LUT4 #(
		.INIT('haebf)
	) name23515 (
		_w8738_,
		_w8741_,
		_w25414_,
		_w25415_,
		_w25416_
	);
	LUT4 #(
		.INIT('h2a00)
	) name23516 (
		\m1_stb_i_pad ,
		_w8743_,
		_w8744_,
		_w9439_,
		_w25417_
	);
	LUT4 #(
		.INIT('h8000)
	) name23517 (
		\m0_stb_i_pad ,
		_w8743_,
		_w8744_,
		_w9404_,
		_w25418_
	);
	LUT3 #(
		.INIT('h57)
	) name23518 (
		_w8742_,
		_w25417_,
		_w25418_,
		_w25419_
	);
	LUT4 #(
		.INIT('h7fff)
	) name23519 (
		_w25410_,
		_w25413_,
		_w25416_,
		_w25419_,
		_w25420_
	);
	LUT3 #(
		.INIT('h2a)
	) name23520 (
		\m3_we_i_pad ,
		_w8743_,
		_w8744_,
		_w25421_
	);
	LUT3 #(
		.INIT('h80)
	) name23521 (
		\m4_we_i_pad ,
		_w8743_,
		_w8744_,
		_w25422_
	);
	LUT4 #(
		.INIT('h9dbf)
	) name23522 (
		_w8738_,
		_w8741_,
		_w25421_,
		_w25422_,
		_w25423_
	);
	LUT3 #(
		.INIT('h80)
	) name23523 (
		\m6_we_i_pad ,
		_w8743_,
		_w8744_,
		_w25424_
	);
	LUT3 #(
		.INIT('h2a)
	) name23524 (
		\m7_we_i_pad ,
		_w8743_,
		_w8744_,
		_w25425_
	);
	LUT3 #(
		.INIT('h57)
	) name23525 (
		_w8756_,
		_w25424_,
		_w25425_,
		_w25426_
	);
	LUT3 #(
		.INIT('h2a)
	) name23526 (
		\m5_we_i_pad ,
		_w8743_,
		_w8744_,
		_w25427_
	);
	LUT3 #(
		.INIT('h80)
	) name23527 (
		\m0_we_i_pad ,
		_w8743_,
		_w8744_,
		_w25428_
	);
	LUT4 #(
		.INIT('h57df)
	) name23528 (
		_w8738_,
		_w8741_,
		_w25427_,
		_w25428_,
		_w25429_
	);
	LUT3 #(
		.INIT('h2a)
	) name23529 (
		\m1_we_i_pad ,
		_w8743_,
		_w8744_,
		_w25430_
	);
	LUT3 #(
		.INIT('h80)
	) name23530 (
		\m2_we_i_pad ,
		_w8743_,
		_w8744_,
		_w25431_
	);
	LUT4 #(
		.INIT('h3b7f)
	) name23531 (
		_w8738_,
		_w8741_,
		_w25430_,
		_w25431_,
		_w25432_
	);
	LUT4 #(
		.INIT('h7fff)
	) name23532 (
		_w25423_,
		_w25426_,
		_w25429_,
		_w25432_,
		_w25433_
	);
	LUT3 #(
		.INIT('h80)
	) name23533 (
		\m0_addr_i[0]_pad ,
		_w8782_,
		_w8783_,
		_w25434_
	);
	LUT3 #(
		.INIT('h2a)
	) name23534 (
		\m7_addr_i[0]_pad ,
		_w8782_,
		_w8783_,
		_w25435_
	);
	LUT4 #(
		.INIT('h6e7f)
	) name23535 (
		_w8777_,
		_w8780_,
		_w25434_,
		_w25435_,
		_w25436_
	);
	LUT3 #(
		.INIT('h2a)
	) name23536 (
		\m3_addr_i[0]_pad ,
		_w8782_,
		_w8783_,
		_w25437_
	);
	LUT3 #(
		.INIT('h2a)
	) name23537 (
		\m5_addr_i[0]_pad ,
		_w8782_,
		_w8783_,
		_w25438_
	);
	LUT4 #(
		.INIT('h9dbf)
	) name23538 (
		_w8777_,
		_w8780_,
		_w25437_,
		_w25438_,
		_w25439_
	);
	LUT3 #(
		.INIT('h80)
	) name23539 (
		\m4_addr_i[0]_pad ,
		_w8782_,
		_w8783_,
		_w25440_
	);
	LUT3 #(
		.INIT('h80)
	) name23540 (
		\m6_addr_i[0]_pad ,
		_w8782_,
		_w8783_,
		_w25441_
	);
	LUT4 #(
		.INIT('hcedf)
	) name23541 (
		_w8777_,
		_w8780_,
		_w25440_,
		_w25441_,
		_w25442_
	);
	LUT3 #(
		.INIT('h2a)
	) name23542 (
		\m1_addr_i[0]_pad ,
		_w8782_,
		_w8783_,
		_w25443_
	);
	LUT3 #(
		.INIT('h80)
	) name23543 (
		\m2_addr_i[0]_pad ,
		_w8782_,
		_w8783_,
		_w25444_
	);
	LUT4 #(
		.INIT('h3b7f)
	) name23544 (
		_w8777_,
		_w8780_,
		_w25443_,
		_w25444_,
		_w25445_
	);
	LUT4 #(
		.INIT('h7fff)
	) name23545 (
		_w25436_,
		_w25439_,
		_w25442_,
		_w25445_,
		_w25446_
	);
	LUT3 #(
		.INIT('h2a)
	) name23546 (
		\m3_addr_i[10]_pad ,
		_w8782_,
		_w8783_,
		_w25447_
	);
	LUT3 #(
		.INIT('h80)
	) name23547 (
		\m4_addr_i[10]_pad ,
		_w8782_,
		_w8783_,
		_w25448_
	);
	LUT4 #(
		.INIT('h9dbf)
	) name23548 (
		_w8777_,
		_w8780_,
		_w25447_,
		_w25448_,
		_w25449_
	);
	LUT3 #(
		.INIT('h80)
	) name23549 (
		\m6_addr_i[10]_pad ,
		_w8782_,
		_w8783_,
		_w25450_
	);
	LUT3 #(
		.INIT('h2a)
	) name23550 (
		\m7_addr_i[10]_pad ,
		_w8782_,
		_w8783_,
		_w25451_
	);
	LUT3 #(
		.INIT('h57)
	) name23551 (
		_w8781_,
		_w25450_,
		_w25451_,
		_w25452_
	);
	LUT3 #(
		.INIT('h2a)
	) name23552 (
		\m5_addr_i[10]_pad ,
		_w8782_,
		_w8783_,
		_w25453_
	);
	LUT3 #(
		.INIT('h80)
	) name23553 (
		\m0_addr_i[10]_pad ,
		_w8782_,
		_w8783_,
		_w25454_
	);
	LUT4 #(
		.INIT('h57df)
	) name23554 (
		_w8777_,
		_w8780_,
		_w25453_,
		_w25454_,
		_w25455_
	);
	LUT3 #(
		.INIT('h2a)
	) name23555 (
		\m1_addr_i[10]_pad ,
		_w8782_,
		_w8783_,
		_w25456_
	);
	LUT3 #(
		.INIT('h80)
	) name23556 (
		\m2_addr_i[10]_pad ,
		_w8782_,
		_w8783_,
		_w25457_
	);
	LUT4 #(
		.INIT('h3b7f)
	) name23557 (
		_w8777_,
		_w8780_,
		_w25456_,
		_w25457_,
		_w25458_
	);
	LUT4 #(
		.INIT('h7fff)
	) name23558 (
		_w25449_,
		_w25452_,
		_w25455_,
		_w25458_,
		_w25459_
	);
	LUT3 #(
		.INIT('h2a)
	) name23559 (
		\m1_addr_i[11]_pad ,
		_w8782_,
		_w8783_,
		_w25460_
	);
	LUT3 #(
		.INIT('h80)
	) name23560 (
		\m2_addr_i[11]_pad ,
		_w8782_,
		_w8783_,
		_w25461_
	);
	LUT4 #(
		.INIT('h3b7f)
	) name23561 (
		_w8777_,
		_w8780_,
		_w25460_,
		_w25461_,
		_w25462_
	);
	LUT3 #(
		.INIT('h80)
	) name23562 (
		\m6_addr_i[11]_pad ,
		_w8782_,
		_w8783_,
		_w25463_
	);
	LUT3 #(
		.INIT('h2a)
	) name23563 (
		\m7_addr_i[11]_pad ,
		_w8782_,
		_w8783_,
		_w25464_
	);
	LUT3 #(
		.INIT('h57)
	) name23564 (
		_w8781_,
		_w25463_,
		_w25464_,
		_w25465_
	);
	LUT3 #(
		.INIT('h2a)
	) name23565 (
		\m5_addr_i[11]_pad ,
		_w8782_,
		_w8783_,
		_w25466_
	);
	LUT3 #(
		.INIT('h80)
	) name23566 (
		\m0_addr_i[11]_pad ,
		_w8782_,
		_w8783_,
		_w25467_
	);
	LUT4 #(
		.INIT('h57df)
	) name23567 (
		_w8777_,
		_w8780_,
		_w25466_,
		_w25467_,
		_w25468_
	);
	LUT3 #(
		.INIT('h2a)
	) name23568 (
		\m3_addr_i[11]_pad ,
		_w8782_,
		_w8783_,
		_w25469_
	);
	LUT3 #(
		.INIT('h80)
	) name23569 (
		\m4_addr_i[11]_pad ,
		_w8782_,
		_w8783_,
		_w25470_
	);
	LUT4 #(
		.INIT('h9dbf)
	) name23570 (
		_w8777_,
		_w8780_,
		_w25469_,
		_w25470_,
		_w25471_
	);
	LUT4 #(
		.INIT('h7fff)
	) name23571 (
		_w25462_,
		_w25465_,
		_w25468_,
		_w25471_,
		_w25472_
	);
	LUT3 #(
		.INIT('h2a)
	) name23572 (
		\m1_addr_i[12]_pad ,
		_w8782_,
		_w8783_,
		_w25473_
	);
	LUT3 #(
		.INIT('h80)
	) name23573 (
		\m2_addr_i[12]_pad ,
		_w8782_,
		_w8783_,
		_w25474_
	);
	LUT4 #(
		.INIT('h3b7f)
	) name23574 (
		_w8777_,
		_w8780_,
		_w25473_,
		_w25474_,
		_w25475_
	);
	LUT3 #(
		.INIT('h80)
	) name23575 (
		\m6_addr_i[12]_pad ,
		_w8782_,
		_w8783_,
		_w25476_
	);
	LUT3 #(
		.INIT('h2a)
	) name23576 (
		\m7_addr_i[12]_pad ,
		_w8782_,
		_w8783_,
		_w25477_
	);
	LUT3 #(
		.INIT('h57)
	) name23577 (
		_w8781_,
		_w25476_,
		_w25477_,
		_w25478_
	);
	LUT3 #(
		.INIT('h2a)
	) name23578 (
		\m5_addr_i[12]_pad ,
		_w8782_,
		_w8783_,
		_w25479_
	);
	LUT3 #(
		.INIT('h80)
	) name23579 (
		\m0_addr_i[12]_pad ,
		_w8782_,
		_w8783_,
		_w25480_
	);
	LUT4 #(
		.INIT('h57df)
	) name23580 (
		_w8777_,
		_w8780_,
		_w25479_,
		_w25480_,
		_w25481_
	);
	LUT3 #(
		.INIT('h2a)
	) name23581 (
		\m3_addr_i[12]_pad ,
		_w8782_,
		_w8783_,
		_w25482_
	);
	LUT3 #(
		.INIT('h80)
	) name23582 (
		\m4_addr_i[12]_pad ,
		_w8782_,
		_w8783_,
		_w25483_
	);
	LUT4 #(
		.INIT('h9dbf)
	) name23583 (
		_w8777_,
		_w8780_,
		_w25482_,
		_w25483_,
		_w25484_
	);
	LUT4 #(
		.INIT('h7fff)
	) name23584 (
		_w25475_,
		_w25478_,
		_w25481_,
		_w25484_,
		_w25485_
	);
	LUT3 #(
		.INIT('h2a)
	) name23585 (
		\m3_addr_i[13]_pad ,
		_w8782_,
		_w8783_,
		_w25486_
	);
	LUT3 #(
		.INIT('h80)
	) name23586 (
		\m4_addr_i[13]_pad ,
		_w8782_,
		_w8783_,
		_w25487_
	);
	LUT4 #(
		.INIT('h9dbf)
	) name23587 (
		_w8777_,
		_w8780_,
		_w25486_,
		_w25487_,
		_w25488_
	);
	LUT3 #(
		.INIT('h80)
	) name23588 (
		\m6_addr_i[13]_pad ,
		_w8782_,
		_w8783_,
		_w25489_
	);
	LUT3 #(
		.INIT('h80)
	) name23589 (
		\m2_addr_i[13]_pad ,
		_w8782_,
		_w8783_,
		_w25490_
	);
	LUT4 #(
		.INIT('habef)
	) name23590 (
		_w8777_,
		_w8780_,
		_w25489_,
		_w25490_,
		_w25491_
	);
	LUT3 #(
		.INIT('h2a)
	) name23591 (
		\m5_addr_i[13]_pad ,
		_w8782_,
		_w8783_,
		_w25492_
	);
	LUT3 #(
		.INIT('h2a)
	) name23592 (
		\m1_addr_i[13]_pad ,
		_w8782_,
		_w8783_,
		_w25493_
	);
	LUT4 #(
		.INIT('h57df)
	) name23593 (
		_w8777_,
		_w8780_,
		_w25492_,
		_w25493_,
		_w25494_
	);
	LUT3 #(
		.INIT('h80)
	) name23594 (
		\m0_addr_i[13]_pad ,
		_w8782_,
		_w8783_,
		_w25495_
	);
	LUT3 #(
		.INIT('h2a)
	) name23595 (
		\m7_addr_i[13]_pad ,
		_w8782_,
		_w8783_,
		_w25496_
	);
	LUT4 #(
		.INIT('h6e7f)
	) name23596 (
		_w8777_,
		_w8780_,
		_w25495_,
		_w25496_,
		_w25497_
	);
	LUT4 #(
		.INIT('h7fff)
	) name23597 (
		_w25488_,
		_w25491_,
		_w25494_,
		_w25497_,
		_w25498_
	);
	LUT3 #(
		.INIT('h2a)
	) name23598 (
		\m3_addr_i[14]_pad ,
		_w8782_,
		_w8783_,
		_w25499_
	);
	LUT3 #(
		.INIT('h80)
	) name23599 (
		\m4_addr_i[14]_pad ,
		_w8782_,
		_w8783_,
		_w25500_
	);
	LUT4 #(
		.INIT('h9dbf)
	) name23600 (
		_w8777_,
		_w8780_,
		_w25499_,
		_w25500_,
		_w25501_
	);
	LUT3 #(
		.INIT('h80)
	) name23601 (
		\m6_addr_i[14]_pad ,
		_w8782_,
		_w8783_,
		_w25502_
	);
	LUT3 #(
		.INIT('h80)
	) name23602 (
		\m2_addr_i[14]_pad ,
		_w8782_,
		_w8783_,
		_w25503_
	);
	LUT4 #(
		.INIT('habef)
	) name23603 (
		_w8777_,
		_w8780_,
		_w25502_,
		_w25503_,
		_w25504_
	);
	LUT3 #(
		.INIT('h2a)
	) name23604 (
		\m5_addr_i[14]_pad ,
		_w8782_,
		_w8783_,
		_w25505_
	);
	LUT3 #(
		.INIT('h2a)
	) name23605 (
		\m1_addr_i[14]_pad ,
		_w8782_,
		_w8783_,
		_w25506_
	);
	LUT4 #(
		.INIT('h57df)
	) name23606 (
		_w8777_,
		_w8780_,
		_w25505_,
		_w25506_,
		_w25507_
	);
	LUT3 #(
		.INIT('h80)
	) name23607 (
		\m0_addr_i[14]_pad ,
		_w8782_,
		_w8783_,
		_w25508_
	);
	LUT3 #(
		.INIT('h2a)
	) name23608 (
		\m7_addr_i[14]_pad ,
		_w8782_,
		_w8783_,
		_w25509_
	);
	LUT4 #(
		.INIT('h6e7f)
	) name23609 (
		_w8777_,
		_w8780_,
		_w25508_,
		_w25509_,
		_w25510_
	);
	LUT4 #(
		.INIT('h7fff)
	) name23610 (
		_w25501_,
		_w25504_,
		_w25507_,
		_w25510_,
		_w25511_
	);
	LUT3 #(
		.INIT('h2a)
	) name23611 (
		\m3_addr_i[15]_pad ,
		_w8782_,
		_w8783_,
		_w25512_
	);
	LUT3 #(
		.INIT('h80)
	) name23612 (
		\m4_addr_i[15]_pad ,
		_w8782_,
		_w8783_,
		_w25513_
	);
	LUT4 #(
		.INIT('h9dbf)
	) name23613 (
		_w8777_,
		_w8780_,
		_w25512_,
		_w25513_,
		_w25514_
	);
	LUT3 #(
		.INIT('h80)
	) name23614 (
		\m6_addr_i[15]_pad ,
		_w8782_,
		_w8783_,
		_w25515_
	);
	LUT3 #(
		.INIT('h80)
	) name23615 (
		\m2_addr_i[15]_pad ,
		_w8782_,
		_w8783_,
		_w25516_
	);
	LUT4 #(
		.INIT('habef)
	) name23616 (
		_w8777_,
		_w8780_,
		_w25515_,
		_w25516_,
		_w25517_
	);
	LUT3 #(
		.INIT('h2a)
	) name23617 (
		\m5_addr_i[15]_pad ,
		_w8782_,
		_w8783_,
		_w25518_
	);
	LUT3 #(
		.INIT('h2a)
	) name23618 (
		\m1_addr_i[15]_pad ,
		_w8782_,
		_w8783_,
		_w25519_
	);
	LUT4 #(
		.INIT('h57df)
	) name23619 (
		_w8777_,
		_w8780_,
		_w25518_,
		_w25519_,
		_w25520_
	);
	LUT3 #(
		.INIT('h80)
	) name23620 (
		\m0_addr_i[15]_pad ,
		_w8782_,
		_w8783_,
		_w25521_
	);
	LUT3 #(
		.INIT('h2a)
	) name23621 (
		\m7_addr_i[15]_pad ,
		_w8782_,
		_w8783_,
		_w25522_
	);
	LUT4 #(
		.INIT('h6e7f)
	) name23622 (
		_w8777_,
		_w8780_,
		_w25521_,
		_w25522_,
		_w25523_
	);
	LUT4 #(
		.INIT('h7fff)
	) name23623 (
		_w25514_,
		_w25517_,
		_w25520_,
		_w25523_,
		_w25524_
	);
	LUT3 #(
		.INIT('h2a)
	) name23624 (
		\m3_addr_i[16]_pad ,
		_w8782_,
		_w8783_,
		_w25525_
	);
	LUT3 #(
		.INIT('h80)
	) name23625 (
		\m4_addr_i[16]_pad ,
		_w8782_,
		_w8783_,
		_w25526_
	);
	LUT4 #(
		.INIT('h9dbf)
	) name23626 (
		_w8777_,
		_w8780_,
		_w25525_,
		_w25526_,
		_w25527_
	);
	LUT3 #(
		.INIT('h80)
	) name23627 (
		\m6_addr_i[16]_pad ,
		_w8782_,
		_w8783_,
		_w25528_
	);
	LUT3 #(
		.INIT('h80)
	) name23628 (
		\m2_addr_i[16]_pad ,
		_w8782_,
		_w8783_,
		_w25529_
	);
	LUT4 #(
		.INIT('habef)
	) name23629 (
		_w8777_,
		_w8780_,
		_w25528_,
		_w25529_,
		_w25530_
	);
	LUT3 #(
		.INIT('h2a)
	) name23630 (
		\m5_addr_i[16]_pad ,
		_w8782_,
		_w8783_,
		_w25531_
	);
	LUT3 #(
		.INIT('h2a)
	) name23631 (
		\m1_addr_i[16]_pad ,
		_w8782_,
		_w8783_,
		_w25532_
	);
	LUT4 #(
		.INIT('h57df)
	) name23632 (
		_w8777_,
		_w8780_,
		_w25531_,
		_w25532_,
		_w25533_
	);
	LUT3 #(
		.INIT('h80)
	) name23633 (
		\m0_addr_i[16]_pad ,
		_w8782_,
		_w8783_,
		_w25534_
	);
	LUT3 #(
		.INIT('h2a)
	) name23634 (
		\m7_addr_i[16]_pad ,
		_w8782_,
		_w8783_,
		_w25535_
	);
	LUT4 #(
		.INIT('h6e7f)
	) name23635 (
		_w8777_,
		_w8780_,
		_w25534_,
		_w25535_,
		_w25536_
	);
	LUT4 #(
		.INIT('h7fff)
	) name23636 (
		_w25527_,
		_w25530_,
		_w25533_,
		_w25536_,
		_w25537_
	);
	LUT3 #(
		.INIT('h2a)
	) name23637 (
		\m1_addr_i[17]_pad ,
		_w8782_,
		_w8783_,
		_w25538_
	);
	LUT3 #(
		.INIT('h80)
	) name23638 (
		\m2_addr_i[17]_pad ,
		_w8782_,
		_w8783_,
		_w25539_
	);
	LUT4 #(
		.INIT('h3b7f)
	) name23639 (
		_w8777_,
		_w8780_,
		_w25538_,
		_w25539_,
		_w25540_
	);
	LUT3 #(
		.INIT('h2a)
	) name23640 (
		\m3_addr_i[17]_pad ,
		_w8782_,
		_w8783_,
		_w25541_
	);
	LUT3 #(
		.INIT('h2a)
	) name23641 (
		\m7_addr_i[17]_pad ,
		_w8782_,
		_w8783_,
		_w25542_
	);
	LUT4 #(
		.INIT('haebf)
	) name23642 (
		_w8777_,
		_w8780_,
		_w25541_,
		_w25542_,
		_w25543_
	);
	LUT3 #(
		.INIT('h80)
	) name23643 (
		\m4_addr_i[17]_pad ,
		_w8782_,
		_w8783_,
		_w25544_
	);
	LUT3 #(
		.INIT('h80)
	) name23644 (
		\m0_addr_i[17]_pad ,
		_w8782_,
		_w8783_,
		_w25545_
	);
	LUT4 #(
		.INIT('h57df)
	) name23645 (
		_w8777_,
		_w8780_,
		_w25544_,
		_w25545_,
		_w25546_
	);
	LUT3 #(
		.INIT('h80)
	) name23646 (
		\m6_addr_i[17]_pad ,
		_w8782_,
		_w8783_,
		_w25547_
	);
	LUT3 #(
		.INIT('h2a)
	) name23647 (
		\m5_addr_i[17]_pad ,
		_w8782_,
		_w8783_,
		_w25548_
	);
	LUT4 #(
		.INIT('hcdef)
	) name23648 (
		_w8777_,
		_w8780_,
		_w25547_,
		_w25548_,
		_w25549_
	);
	LUT4 #(
		.INIT('h7fff)
	) name23649 (
		_w25540_,
		_w25543_,
		_w25546_,
		_w25549_,
		_w25550_
	);
	LUT3 #(
		.INIT('h2a)
	) name23650 (
		\m1_addr_i[18]_pad ,
		_w8782_,
		_w8783_,
		_w25551_
	);
	LUT3 #(
		.INIT('h80)
	) name23651 (
		\m2_addr_i[18]_pad ,
		_w8782_,
		_w8783_,
		_w25552_
	);
	LUT4 #(
		.INIT('h3b7f)
	) name23652 (
		_w8777_,
		_w8780_,
		_w25551_,
		_w25552_,
		_w25553_
	);
	LUT3 #(
		.INIT('h2a)
	) name23653 (
		\m3_addr_i[18]_pad ,
		_w8782_,
		_w8783_,
		_w25554_
	);
	LUT3 #(
		.INIT('h2a)
	) name23654 (
		\m7_addr_i[18]_pad ,
		_w8782_,
		_w8783_,
		_w25555_
	);
	LUT4 #(
		.INIT('haebf)
	) name23655 (
		_w8777_,
		_w8780_,
		_w25554_,
		_w25555_,
		_w25556_
	);
	LUT3 #(
		.INIT('h80)
	) name23656 (
		\m4_addr_i[18]_pad ,
		_w8782_,
		_w8783_,
		_w25557_
	);
	LUT3 #(
		.INIT('h80)
	) name23657 (
		\m0_addr_i[18]_pad ,
		_w8782_,
		_w8783_,
		_w25558_
	);
	LUT4 #(
		.INIT('h57df)
	) name23658 (
		_w8777_,
		_w8780_,
		_w25557_,
		_w25558_,
		_w25559_
	);
	LUT3 #(
		.INIT('h80)
	) name23659 (
		\m6_addr_i[18]_pad ,
		_w8782_,
		_w8783_,
		_w25560_
	);
	LUT3 #(
		.INIT('h2a)
	) name23660 (
		\m5_addr_i[18]_pad ,
		_w8782_,
		_w8783_,
		_w25561_
	);
	LUT4 #(
		.INIT('hcdef)
	) name23661 (
		_w8777_,
		_w8780_,
		_w25560_,
		_w25561_,
		_w25562_
	);
	LUT4 #(
		.INIT('h7fff)
	) name23662 (
		_w25553_,
		_w25556_,
		_w25559_,
		_w25562_,
		_w25563_
	);
	LUT3 #(
		.INIT('h2a)
	) name23663 (
		\m3_addr_i[19]_pad ,
		_w8782_,
		_w8783_,
		_w25564_
	);
	LUT3 #(
		.INIT('h80)
	) name23664 (
		\m4_addr_i[19]_pad ,
		_w8782_,
		_w8783_,
		_w25565_
	);
	LUT4 #(
		.INIT('h9dbf)
	) name23665 (
		_w8777_,
		_w8780_,
		_w25564_,
		_w25565_,
		_w25566_
	);
	LUT3 #(
		.INIT('h80)
	) name23666 (
		\m6_addr_i[19]_pad ,
		_w8782_,
		_w8783_,
		_w25567_
	);
	LUT3 #(
		.INIT('h2a)
	) name23667 (
		\m7_addr_i[19]_pad ,
		_w8782_,
		_w8783_,
		_w25568_
	);
	LUT3 #(
		.INIT('h57)
	) name23668 (
		_w8781_,
		_w25567_,
		_w25568_,
		_w25569_
	);
	LUT3 #(
		.INIT('h2a)
	) name23669 (
		\m5_addr_i[19]_pad ,
		_w8782_,
		_w8783_,
		_w25570_
	);
	LUT3 #(
		.INIT('h80)
	) name23670 (
		\m0_addr_i[19]_pad ,
		_w8782_,
		_w8783_,
		_w25571_
	);
	LUT4 #(
		.INIT('h57df)
	) name23671 (
		_w8777_,
		_w8780_,
		_w25570_,
		_w25571_,
		_w25572_
	);
	LUT3 #(
		.INIT('h2a)
	) name23672 (
		\m1_addr_i[19]_pad ,
		_w8782_,
		_w8783_,
		_w25573_
	);
	LUT3 #(
		.INIT('h80)
	) name23673 (
		\m2_addr_i[19]_pad ,
		_w8782_,
		_w8783_,
		_w25574_
	);
	LUT4 #(
		.INIT('h3b7f)
	) name23674 (
		_w8777_,
		_w8780_,
		_w25573_,
		_w25574_,
		_w25575_
	);
	LUT4 #(
		.INIT('h7fff)
	) name23675 (
		_w25566_,
		_w25569_,
		_w25572_,
		_w25575_,
		_w25576_
	);
	LUT3 #(
		.INIT('h2a)
	) name23676 (
		\m3_addr_i[1]_pad ,
		_w8782_,
		_w8783_,
		_w25577_
	);
	LUT3 #(
		.INIT('h80)
	) name23677 (
		\m4_addr_i[1]_pad ,
		_w8782_,
		_w8783_,
		_w25578_
	);
	LUT4 #(
		.INIT('h9dbf)
	) name23678 (
		_w8777_,
		_w8780_,
		_w25577_,
		_w25578_,
		_w25579_
	);
	LUT3 #(
		.INIT('h80)
	) name23679 (
		\m6_addr_i[1]_pad ,
		_w8782_,
		_w8783_,
		_w25580_
	);
	LUT3 #(
		.INIT('h80)
	) name23680 (
		\m2_addr_i[1]_pad ,
		_w8782_,
		_w8783_,
		_w25581_
	);
	LUT4 #(
		.INIT('habef)
	) name23681 (
		_w8777_,
		_w8780_,
		_w25580_,
		_w25581_,
		_w25582_
	);
	LUT3 #(
		.INIT('h2a)
	) name23682 (
		\m5_addr_i[1]_pad ,
		_w8782_,
		_w8783_,
		_w25583_
	);
	LUT3 #(
		.INIT('h2a)
	) name23683 (
		\m1_addr_i[1]_pad ,
		_w8782_,
		_w8783_,
		_w25584_
	);
	LUT4 #(
		.INIT('h57df)
	) name23684 (
		_w8777_,
		_w8780_,
		_w25583_,
		_w25584_,
		_w25585_
	);
	LUT3 #(
		.INIT('h80)
	) name23685 (
		\m0_addr_i[1]_pad ,
		_w8782_,
		_w8783_,
		_w25586_
	);
	LUT3 #(
		.INIT('h2a)
	) name23686 (
		\m7_addr_i[1]_pad ,
		_w8782_,
		_w8783_,
		_w25587_
	);
	LUT4 #(
		.INIT('h6e7f)
	) name23687 (
		_w8777_,
		_w8780_,
		_w25586_,
		_w25587_,
		_w25588_
	);
	LUT4 #(
		.INIT('h7fff)
	) name23688 (
		_w25579_,
		_w25582_,
		_w25585_,
		_w25588_,
		_w25589_
	);
	LUT3 #(
		.INIT('h80)
	) name23689 (
		\m0_addr_i[20]_pad ,
		_w8782_,
		_w8783_,
		_w25590_
	);
	LUT3 #(
		.INIT('h2a)
	) name23690 (
		\m7_addr_i[20]_pad ,
		_w8782_,
		_w8783_,
		_w25591_
	);
	LUT4 #(
		.INIT('h6e7f)
	) name23691 (
		_w8777_,
		_w8780_,
		_w25590_,
		_w25591_,
		_w25592_
	);
	LUT3 #(
		.INIT('h2a)
	) name23692 (
		\m3_addr_i[20]_pad ,
		_w8782_,
		_w8783_,
		_w25593_
	);
	LUT3 #(
		.INIT('h80)
	) name23693 (
		\m2_addr_i[20]_pad ,
		_w8782_,
		_w8783_,
		_w25594_
	);
	LUT3 #(
		.INIT('h57)
	) name23694 (
		_w8795_,
		_w25593_,
		_w25594_,
		_w25595_
	);
	LUT3 #(
		.INIT('h80)
	) name23695 (
		\m4_addr_i[20]_pad ,
		_w8782_,
		_w8783_,
		_w25596_
	);
	LUT3 #(
		.INIT('h2a)
	) name23696 (
		\m1_addr_i[20]_pad ,
		_w8782_,
		_w8783_,
		_w25597_
	);
	LUT4 #(
		.INIT('h57df)
	) name23697 (
		_w8777_,
		_w8780_,
		_w25596_,
		_w25597_,
		_w25598_
	);
	LUT3 #(
		.INIT('h80)
	) name23698 (
		\m6_addr_i[20]_pad ,
		_w8782_,
		_w8783_,
		_w25599_
	);
	LUT3 #(
		.INIT('h2a)
	) name23699 (
		\m5_addr_i[20]_pad ,
		_w8782_,
		_w8783_,
		_w25600_
	);
	LUT4 #(
		.INIT('hcdef)
	) name23700 (
		_w8777_,
		_w8780_,
		_w25599_,
		_w25600_,
		_w25601_
	);
	LUT4 #(
		.INIT('h7fff)
	) name23701 (
		_w25592_,
		_w25595_,
		_w25598_,
		_w25601_,
		_w25602_
	);
	LUT3 #(
		.INIT('h2a)
	) name23702 (
		\m3_addr_i[21]_pad ,
		_w8782_,
		_w8783_,
		_w25603_
	);
	LUT3 #(
		.INIT('h80)
	) name23703 (
		\m4_addr_i[21]_pad ,
		_w8782_,
		_w8783_,
		_w25604_
	);
	LUT4 #(
		.INIT('h9dbf)
	) name23704 (
		_w8777_,
		_w8780_,
		_w25603_,
		_w25604_,
		_w25605_
	);
	LUT3 #(
		.INIT('h80)
	) name23705 (
		\m6_addr_i[21]_pad ,
		_w8782_,
		_w8783_,
		_w25606_
	);
	LUT3 #(
		.INIT('h2a)
	) name23706 (
		\m7_addr_i[21]_pad ,
		_w8782_,
		_w8783_,
		_w25607_
	);
	LUT3 #(
		.INIT('h57)
	) name23707 (
		_w8781_,
		_w25606_,
		_w25607_,
		_w25608_
	);
	LUT3 #(
		.INIT('h2a)
	) name23708 (
		\m5_addr_i[21]_pad ,
		_w8782_,
		_w8783_,
		_w25609_
	);
	LUT3 #(
		.INIT('h80)
	) name23709 (
		\m0_addr_i[21]_pad ,
		_w8782_,
		_w8783_,
		_w25610_
	);
	LUT4 #(
		.INIT('h57df)
	) name23710 (
		_w8777_,
		_w8780_,
		_w25609_,
		_w25610_,
		_w25611_
	);
	LUT3 #(
		.INIT('h2a)
	) name23711 (
		\m1_addr_i[21]_pad ,
		_w8782_,
		_w8783_,
		_w25612_
	);
	LUT3 #(
		.INIT('h80)
	) name23712 (
		\m2_addr_i[21]_pad ,
		_w8782_,
		_w8783_,
		_w25613_
	);
	LUT4 #(
		.INIT('h3b7f)
	) name23713 (
		_w8777_,
		_w8780_,
		_w25612_,
		_w25613_,
		_w25614_
	);
	LUT4 #(
		.INIT('h7fff)
	) name23714 (
		_w25605_,
		_w25608_,
		_w25611_,
		_w25614_,
		_w25615_
	);
	LUT3 #(
		.INIT('h2a)
	) name23715 (
		\m1_addr_i[22]_pad ,
		_w8782_,
		_w8783_,
		_w25616_
	);
	LUT3 #(
		.INIT('h80)
	) name23716 (
		\m2_addr_i[22]_pad ,
		_w8782_,
		_w8783_,
		_w25617_
	);
	LUT4 #(
		.INIT('h3b7f)
	) name23717 (
		_w8777_,
		_w8780_,
		_w25616_,
		_w25617_,
		_w25618_
	);
	LUT3 #(
		.INIT('h2a)
	) name23718 (
		\m3_addr_i[22]_pad ,
		_w8782_,
		_w8783_,
		_w25619_
	);
	LUT3 #(
		.INIT('h2a)
	) name23719 (
		\m7_addr_i[22]_pad ,
		_w8782_,
		_w8783_,
		_w25620_
	);
	LUT4 #(
		.INIT('haebf)
	) name23720 (
		_w8777_,
		_w8780_,
		_w25619_,
		_w25620_,
		_w25621_
	);
	LUT3 #(
		.INIT('h80)
	) name23721 (
		\m4_addr_i[22]_pad ,
		_w8782_,
		_w8783_,
		_w25622_
	);
	LUT3 #(
		.INIT('h80)
	) name23722 (
		\m0_addr_i[22]_pad ,
		_w8782_,
		_w8783_,
		_w25623_
	);
	LUT4 #(
		.INIT('h57df)
	) name23723 (
		_w8777_,
		_w8780_,
		_w25622_,
		_w25623_,
		_w25624_
	);
	LUT3 #(
		.INIT('h80)
	) name23724 (
		\m6_addr_i[22]_pad ,
		_w8782_,
		_w8783_,
		_w25625_
	);
	LUT3 #(
		.INIT('h2a)
	) name23725 (
		\m5_addr_i[22]_pad ,
		_w8782_,
		_w8783_,
		_w25626_
	);
	LUT4 #(
		.INIT('hcdef)
	) name23726 (
		_w8777_,
		_w8780_,
		_w25625_,
		_w25626_,
		_w25627_
	);
	LUT4 #(
		.INIT('h7fff)
	) name23727 (
		_w25618_,
		_w25621_,
		_w25624_,
		_w25627_,
		_w25628_
	);
	LUT3 #(
		.INIT('h2a)
	) name23728 (
		\m1_addr_i[23]_pad ,
		_w8782_,
		_w8783_,
		_w25629_
	);
	LUT3 #(
		.INIT('h80)
	) name23729 (
		\m2_addr_i[23]_pad ,
		_w8782_,
		_w8783_,
		_w25630_
	);
	LUT4 #(
		.INIT('h3b7f)
	) name23730 (
		_w8777_,
		_w8780_,
		_w25629_,
		_w25630_,
		_w25631_
	);
	LUT3 #(
		.INIT('h2a)
	) name23731 (
		\m3_addr_i[23]_pad ,
		_w8782_,
		_w8783_,
		_w25632_
	);
	LUT3 #(
		.INIT('h2a)
	) name23732 (
		\m5_addr_i[23]_pad ,
		_w8782_,
		_w8783_,
		_w25633_
	);
	LUT4 #(
		.INIT('h9dbf)
	) name23733 (
		_w8777_,
		_w8780_,
		_w25632_,
		_w25633_,
		_w25634_
	);
	LUT3 #(
		.INIT('h80)
	) name23734 (
		\m4_addr_i[23]_pad ,
		_w8782_,
		_w8783_,
		_w25635_
	);
	LUT3 #(
		.INIT('h80)
	) name23735 (
		\m6_addr_i[23]_pad ,
		_w8782_,
		_w8783_,
		_w25636_
	);
	LUT4 #(
		.INIT('hcedf)
	) name23736 (
		_w8777_,
		_w8780_,
		_w25635_,
		_w25636_,
		_w25637_
	);
	LUT3 #(
		.INIT('h80)
	) name23737 (
		\m0_addr_i[23]_pad ,
		_w8782_,
		_w8783_,
		_w25638_
	);
	LUT3 #(
		.INIT('h2a)
	) name23738 (
		\m7_addr_i[23]_pad ,
		_w8782_,
		_w8783_,
		_w25639_
	);
	LUT4 #(
		.INIT('h6e7f)
	) name23739 (
		_w8777_,
		_w8780_,
		_w25638_,
		_w25639_,
		_w25640_
	);
	LUT4 #(
		.INIT('h7fff)
	) name23740 (
		_w25631_,
		_w25634_,
		_w25637_,
		_w25640_,
		_w25641_
	);
	LUT3 #(
		.INIT('h2a)
	) name23741 (
		\m1_addr_i[24]_pad ,
		_w8782_,
		_w8783_,
		_w25642_
	);
	LUT3 #(
		.INIT('h80)
	) name23742 (
		\m2_addr_i[24]_pad ,
		_w8782_,
		_w8783_,
		_w25643_
	);
	LUT4 #(
		.INIT('h3b7f)
	) name23743 (
		_w8777_,
		_w8780_,
		_w25642_,
		_w25643_,
		_w25644_
	);
	LUT3 #(
		.INIT('h2a)
	) name23744 (
		\m5_addr_i[24]_pad ,
		_w8782_,
		_w8783_,
		_w25645_
	);
	LUT3 #(
		.INIT('h80)
	) name23745 (
		\m4_addr_i[24]_pad ,
		_w8782_,
		_w8783_,
		_w25646_
	);
	LUT3 #(
		.INIT('h57)
	) name23746 (
		_w8801_,
		_w25645_,
		_w25646_,
		_w25647_
	);
	LUT3 #(
		.INIT('h80)
	) name23747 (
		\m6_addr_i[24]_pad ,
		_w8782_,
		_w8783_,
		_w25648_
	);
	LUT3 #(
		.INIT('h2a)
	) name23748 (
		\m3_addr_i[24]_pad ,
		_w8782_,
		_w8783_,
		_w25649_
	);
	LUT4 #(
		.INIT('habef)
	) name23749 (
		_w8777_,
		_w8780_,
		_w25648_,
		_w25649_,
		_w25650_
	);
	LUT3 #(
		.INIT('h80)
	) name23750 (
		\m0_addr_i[24]_pad ,
		_w8782_,
		_w8783_,
		_w25651_
	);
	LUT3 #(
		.INIT('h2a)
	) name23751 (
		\m7_addr_i[24]_pad ,
		_w8782_,
		_w8783_,
		_w25652_
	);
	LUT4 #(
		.INIT('h6e7f)
	) name23752 (
		_w8777_,
		_w8780_,
		_w25651_,
		_w25652_,
		_w25653_
	);
	LUT4 #(
		.INIT('h7fff)
	) name23753 (
		_w25644_,
		_w25647_,
		_w25650_,
		_w25653_,
		_w25654_
	);
	LUT3 #(
		.INIT('h2a)
	) name23754 (
		\m3_addr_i[25]_pad ,
		_w8782_,
		_w8783_,
		_w25655_
	);
	LUT3 #(
		.INIT('h80)
	) name23755 (
		\m4_addr_i[25]_pad ,
		_w8782_,
		_w8783_,
		_w25656_
	);
	LUT4 #(
		.INIT('h9dbf)
	) name23756 (
		_w8777_,
		_w8780_,
		_w25655_,
		_w25656_,
		_w25657_
	);
	LUT3 #(
		.INIT('h2a)
	) name23757 (
		\m5_addr_i[25]_pad ,
		_w8782_,
		_w8783_,
		_w25658_
	);
	LUT3 #(
		.INIT('h80)
	) name23758 (
		\m2_addr_i[25]_pad ,
		_w8782_,
		_w8783_,
		_w25659_
	);
	LUT4 #(
		.INIT('h9bdf)
	) name23759 (
		_w8777_,
		_w8780_,
		_w25658_,
		_w25659_,
		_w25660_
	);
	LUT3 #(
		.INIT('h80)
	) name23760 (
		\m6_addr_i[25]_pad ,
		_w8782_,
		_w8783_,
		_w25661_
	);
	LUT3 #(
		.INIT('h2a)
	) name23761 (
		\m1_addr_i[25]_pad ,
		_w8782_,
		_w8783_,
		_w25662_
	);
	LUT4 #(
		.INIT('h67ef)
	) name23762 (
		_w8777_,
		_w8780_,
		_w25661_,
		_w25662_,
		_w25663_
	);
	LUT3 #(
		.INIT('h80)
	) name23763 (
		\m0_addr_i[25]_pad ,
		_w8782_,
		_w8783_,
		_w25664_
	);
	LUT3 #(
		.INIT('h2a)
	) name23764 (
		\m7_addr_i[25]_pad ,
		_w8782_,
		_w8783_,
		_w25665_
	);
	LUT4 #(
		.INIT('h6e7f)
	) name23765 (
		_w8777_,
		_w8780_,
		_w25664_,
		_w25665_,
		_w25666_
	);
	LUT4 #(
		.INIT('h7fff)
	) name23766 (
		_w25657_,
		_w25660_,
		_w25663_,
		_w25666_,
		_w25667_
	);
	LUT3 #(
		.INIT('h2a)
	) name23767 (
		\m1_addr_i[26]_pad ,
		_w8782_,
		_w8783_,
		_w25668_
	);
	LUT3 #(
		.INIT('h80)
	) name23768 (
		\m2_addr_i[26]_pad ,
		_w8782_,
		_w8783_,
		_w25669_
	);
	LUT4 #(
		.INIT('h3b7f)
	) name23769 (
		_w8777_,
		_w8780_,
		_w25668_,
		_w25669_,
		_w25670_
	);
	LUT3 #(
		.INIT('h2a)
	) name23770 (
		\m3_addr_i[26]_pad ,
		_w8782_,
		_w8783_,
		_w25671_
	);
	LUT3 #(
		.INIT('h2a)
	) name23771 (
		\m7_addr_i[26]_pad ,
		_w8782_,
		_w8783_,
		_w25672_
	);
	LUT4 #(
		.INIT('haebf)
	) name23772 (
		_w8777_,
		_w8780_,
		_w25671_,
		_w25672_,
		_w25673_
	);
	LUT3 #(
		.INIT('h80)
	) name23773 (
		\m4_addr_i[26]_pad ,
		_w8782_,
		_w8783_,
		_w25674_
	);
	LUT3 #(
		.INIT('h80)
	) name23774 (
		\m0_addr_i[26]_pad ,
		_w8782_,
		_w8783_,
		_w25675_
	);
	LUT4 #(
		.INIT('h57df)
	) name23775 (
		_w8777_,
		_w8780_,
		_w25674_,
		_w25675_,
		_w25676_
	);
	LUT3 #(
		.INIT('h2a)
	) name23776 (
		\m5_addr_i[26]_pad ,
		_w8782_,
		_w8783_,
		_w25677_
	);
	LUT3 #(
		.INIT('h80)
	) name23777 (
		\m6_addr_i[26]_pad ,
		_w8782_,
		_w8783_,
		_w25678_
	);
	LUT4 #(
		.INIT('hcedf)
	) name23778 (
		_w8777_,
		_w8780_,
		_w25677_,
		_w25678_,
		_w25679_
	);
	LUT4 #(
		.INIT('h7fff)
	) name23779 (
		_w25670_,
		_w25673_,
		_w25676_,
		_w25679_,
		_w25680_
	);
	LUT3 #(
		.INIT('h2a)
	) name23780 (
		\m3_addr_i[27]_pad ,
		_w8782_,
		_w8783_,
		_w25681_
	);
	LUT3 #(
		.INIT('h80)
	) name23781 (
		\m4_addr_i[27]_pad ,
		_w8782_,
		_w8783_,
		_w25682_
	);
	LUT4 #(
		.INIT('h9dbf)
	) name23782 (
		_w8777_,
		_w8780_,
		_w25681_,
		_w25682_,
		_w25683_
	);
	LUT3 #(
		.INIT('h2a)
	) name23783 (
		\m5_addr_i[27]_pad ,
		_w8782_,
		_w8783_,
		_w25684_
	);
	LUT3 #(
		.INIT('h2a)
	) name23784 (
		\m7_addr_i[27]_pad ,
		_w8782_,
		_w8783_,
		_w25685_
	);
	LUT4 #(
		.INIT('hcedf)
	) name23785 (
		_w8777_,
		_w8780_,
		_w25684_,
		_w25685_,
		_w25686_
	);
	LUT3 #(
		.INIT('h80)
	) name23786 (
		\m6_addr_i[27]_pad ,
		_w8782_,
		_w8783_,
		_w25687_
	);
	LUT3 #(
		.INIT('h80)
	) name23787 (
		\m0_addr_i[27]_pad ,
		_w8782_,
		_w8783_,
		_w25688_
	);
	LUT4 #(
		.INIT('h67ef)
	) name23788 (
		_w8777_,
		_w8780_,
		_w25687_,
		_w25688_,
		_w25689_
	);
	LUT3 #(
		.INIT('h2a)
	) name23789 (
		\m1_addr_i[27]_pad ,
		_w8782_,
		_w8783_,
		_w25690_
	);
	LUT3 #(
		.INIT('h80)
	) name23790 (
		\m2_addr_i[27]_pad ,
		_w8782_,
		_w8783_,
		_w25691_
	);
	LUT4 #(
		.INIT('h3b7f)
	) name23791 (
		_w8777_,
		_w8780_,
		_w25690_,
		_w25691_,
		_w25692_
	);
	LUT4 #(
		.INIT('h7fff)
	) name23792 (
		_w25683_,
		_w25686_,
		_w25689_,
		_w25692_,
		_w25693_
	);
	LUT3 #(
		.INIT('h2a)
	) name23793 (
		\m1_addr_i[28]_pad ,
		_w8782_,
		_w8783_,
		_w25694_
	);
	LUT3 #(
		.INIT('h80)
	) name23794 (
		\m2_addr_i[28]_pad ,
		_w8782_,
		_w8783_,
		_w25695_
	);
	LUT4 #(
		.INIT('h3b7f)
	) name23795 (
		_w8777_,
		_w8780_,
		_w25694_,
		_w25695_,
		_w25696_
	);
	LUT3 #(
		.INIT('h2a)
	) name23796 (
		\m5_addr_i[28]_pad ,
		_w8782_,
		_w8783_,
		_w25697_
	);
	LUT3 #(
		.INIT('h2a)
	) name23797 (
		\m7_addr_i[28]_pad ,
		_w8782_,
		_w8783_,
		_w25698_
	);
	LUT4 #(
		.INIT('hcedf)
	) name23798 (
		_w8777_,
		_w8780_,
		_w25697_,
		_w25698_,
		_w25699_
	);
	LUT3 #(
		.INIT('h80)
	) name23799 (
		\m6_addr_i[28]_pad ,
		_w8782_,
		_w8783_,
		_w25700_
	);
	LUT3 #(
		.INIT('h80)
	) name23800 (
		\m0_addr_i[28]_pad ,
		_w8782_,
		_w8783_,
		_w25701_
	);
	LUT4 #(
		.INIT('h67ef)
	) name23801 (
		_w8777_,
		_w8780_,
		_w25700_,
		_w25701_,
		_w25702_
	);
	LUT3 #(
		.INIT('h2a)
	) name23802 (
		\m3_addr_i[28]_pad ,
		_w8782_,
		_w8783_,
		_w25703_
	);
	LUT3 #(
		.INIT('h80)
	) name23803 (
		\m4_addr_i[28]_pad ,
		_w8782_,
		_w8783_,
		_w25704_
	);
	LUT4 #(
		.INIT('h9dbf)
	) name23804 (
		_w8777_,
		_w8780_,
		_w25703_,
		_w25704_,
		_w25705_
	);
	LUT4 #(
		.INIT('h7fff)
	) name23805 (
		_w25696_,
		_w25699_,
		_w25702_,
		_w25705_,
		_w25706_
	);
	LUT3 #(
		.INIT('h80)
	) name23806 (
		\m0_addr_i[29]_pad ,
		_w8782_,
		_w8783_,
		_w25707_
	);
	LUT3 #(
		.INIT('h2a)
	) name23807 (
		\m7_addr_i[29]_pad ,
		_w8782_,
		_w8783_,
		_w25708_
	);
	LUT4 #(
		.INIT('h6e7f)
	) name23808 (
		_w8777_,
		_w8780_,
		_w25707_,
		_w25708_,
		_w25709_
	);
	LUT3 #(
		.INIT('h2a)
	) name23809 (
		\m1_addr_i[29]_pad ,
		_w8782_,
		_w8783_,
		_w25710_
	);
	LUT3 #(
		.INIT('h80)
	) name23810 (
		\m4_addr_i[29]_pad ,
		_w8782_,
		_w8783_,
		_w25711_
	);
	LUT4 #(
		.INIT('h5d7f)
	) name23811 (
		_w8777_,
		_w8780_,
		_w25710_,
		_w25711_,
		_w25712_
	);
	LUT3 #(
		.INIT('h80)
	) name23812 (
		\m2_addr_i[29]_pad ,
		_w8782_,
		_w8783_,
		_w25713_
	);
	LUT3 #(
		.INIT('h2a)
	) name23813 (
		\m3_addr_i[29]_pad ,
		_w8782_,
		_w8783_,
		_w25714_
	);
	LUT3 #(
		.INIT('h57)
	) name23814 (
		_w8795_,
		_w25713_,
		_w25714_,
		_w25715_
	);
	LUT3 #(
		.INIT('h2a)
	) name23815 (
		\m5_addr_i[29]_pad ,
		_w8782_,
		_w8783_,
		_w25716_
	);
	LUT3 #(
		.INIT('h80)
	) name23816 (
		\m6_addr_i[29]_pad ,
		_w8782_,
		_w8783_,
		_w25717_
	);
	LUT4 #(
		.INIT('hcedf)
	) name23817 (
		_w8777_,
		_w8780_,
		_w25716_,
		_w25717_,
		_w25718_
	);
	LUT4 #(
		.INIT('h7fff)
	) name23818 (
		_w25709_,
		_w25712_,
		_w25715_,
		_w25718_,
		_w25719_
	);
	LUT3 #(
		.INIT('h2a)
	) name23819 (
		\m3_addr_i[2]_pad ,
		_w8782_,
		_w8783_,
		_w25720_
	);
	LUT3 #(
		.INIT('h80)
	) name23820 (
		\m4_addr_i[2]_pad ,
		_w8782_,
		_w8783_,
		_w25721_
	);
	LUT4 #(
		.INIT('h9dbf)
	) name23821 (
		_w8777_,
		_w8780_,
		_w25720_,
		_w25721_,
		_w25722_
	);
	LUT3 #(
		.INIT('h80)
	) name23822 (
		\m6_addr_i[2]_pad ,
		_w8782_,
		_w8783_,
		_w25723_
	);
	LUT3 #(
		.INIT('h2a)
	) name23823 (
		\m7_addr_i[2]_pad ,
		_w8782_,
		_w8783_,
		_w25724_
	);
	LUT3 #(
		.INIT('h57)
	) name23824 (
		_w8781_,
		_w25723_,
		_w25724_,
		_w25725_
	);
	LUT3 #(
		.INIT('h2a)
	) name23825 (
		\m5_addr_i[2]_pad ,
		_w8782_,
		_w8783_,
		_w25726_
	);
	LUT3 #(
		.INIT('h80)
	) name23826 (
		\m0_addr_i[2]_pad ,
		_w8782_,
		_w8783_,
		_w25727_
	);
	LUT4 #(
		.INIT('h57df)
	) name23827 (
		_w8777_,
		_w8780_,
		_w25726_,
		_w25727_,
		_w25728_
	);
	LUT3 #(
		.INIT('h2a)
	) name23828 (
		\m1_addr_i[2]_pad ,
		_w8782_,
		_w8783_,
		_w25729_
	);
	LUT3 #(
		.INIT('h80)
	) name23829 (
		\m2_addr_i[2]_pad ,
		_w8782_,
		_w8783_,
		_w25730_
	);
	LUT4 #(
		.INIT('h3b7f)
	) name23830 (
		_w8777_,
		_w8780_,
		_w25729_,
		_w25730_,
		_w25731_
	);
	LUT4 #(
		.INIT('h7fff)
	) name23831 (
		_w25722_,
		_w25725_,
		_w25728_,
		_w25731_,
		_w25732_
	);
	LUT3 #(
		.INIT('h2a)
	) name23832 (
		\m1_addr_i[30]_pad ,
		_w8782_,
		_w8783_,
		_w25733_
	);
	LUT3 #(
		.INIT('h80)
	) name23833 (
		\m2_addr_i[30]_pad ,
		_w8782_,
		_w8783_,
		_w25734_
	);
	LUT4 #(
		.INIT('h3b7f)
	) name23834 (
		_w8777_,
		_w8780_,
		_w25733_,
		_w25734_,
		_w25735_
	);
	LUT3 #(
		.INIT('h2a)
	) name23835 (
		\m3_addr_i[30]_pad ,
		_w8782_,
		_w8783_,
		_w25736_
	);
	LUT3 #(
		.INIT('h2a)
	) name23836 (
		\m7_addr_i[30]_pad ,
		_w8782_,
		_w8783_,
		_w25737_
	);
	LUT4 #(
		.INIT('haebf)
	) name23837 (
		_w8777_,
		_w8780_,
		_w25736_,
		_w25737_,
		_w25738_
	);
	LUT3 #(
		.INIT('h80)
	) name23838 (
		\m4_addr_i[30]_pad ,
		_w8782_,
		_w8783_,
		_w25739_
	);
	LUT3 #(
		.INIT('h80)
	) name23839 (
		\m0_addr_i[30]_pad ,
		_w8782_,
		_w8783_,
		_w25740_
	);
	LUT4 #(
		.INIT('h57df)
	) name23840 (
		_w8777_,
		_w8780_,
		_w25739_,
		_w25740_,
		_w25741_
	);
	LUT3 #(
		.INIT('h2a)
	) name23841 (
		\m5_addr_i[30]_pad ,
		_w8782_,
		_w8783_,
		_w25742_
	);
	LUT3 #(
		.INIT('h80)
	) name23842 (
		\m6_addr_i[30]_pad ,
		_w8782_,
		_w8783_,
		_w25743_
	);
	LUT4 #(
		.INIT('hcedf)
	) name23843 (
		_w8777_,
		_w8780_,
		_w25742_,
		_w25743_,
		_w25744_
	);
	LUT4 #(
		.INIT('h7fff)
	) name23844 (
		_w25735_,
		_w25738_,
		_w25741_,
		_w25744_,
		_w25745_
	);
	LUT3 #(
		.INIT('h2a)
	) name23845 (
		\m3_addr_i[31]_pad ,
		_w8782_,
		_w8783_,
		_w25746_
	);
	LUT3 #(
		.INIT('h80)
	) name23846 (
		\m4_addr_i[31]_pad ,
		_w8782_,
		_w8783_,
		_w25747_
	);
	LUT4 #(
		.INIT('h9dbf)
	) name23847 (
		_w8777_,
		_w8780_,
		_w25746_,
		_w25747_,
		_w25748_
	);
	LUT3 #(
		.INIT('h2a)
	) name23848 (
		\m5_addr_i[31]_pad ,
		_w8782_,
		_w8783_,
		_w25749_
	);
	LUT3 #(
		.INIT('h80)
	) name23849 (
		\m2_addr_i[31]_pad ,
		_w8782_,
		_w8783_,
		_w25750_
	);
	LUT4 #(
		.INIT('h9bdf)
	) name23850 (
		_w8777_,
		_w8780_,
		_w25749_,
		_w25750_,
		_w25751_
	);
	LUT3 #(
		.INIT('h80)
	) name23851 (
		\m6_addr_i[31]_pad ,
		_w8782_,
		_w8783_,
		_w25752_
	);
	LUT3 #(
		.INIT('h2a)
	) name23852 (
		\m1_addr_i[31]_pad ,
		_w8782_,
		_w8783_,
		_w25753_
	);
	LUT4 #(
		.INIT('h67ef)
	) name23853 (
		_w8777_,
		_w8780_,
		_w25752_,
		_w25753_,
		_w25754_
	);
	LUT3 #(
		.INIT('h80)
	) name23854 (
		\m0_addr_i[31]_pad ,
		_w8782_,
		_w8783_,
		_w25755_
	);
	LUT3 #(
		.INIT('h2a)
	) name23855 (
		\m7_addr_i[31]_pad ,
		_w8782_,
		_w8783_,
		_w25756_
	);
	LUT4 #(
		.INIT('h6e7f)
	) name23856 (
		_w8777_,
		_w8780_,
		_w25755_,
		_w25756_,
		_w25757_
	);
	LUT4 #(
		.INIT('h7fff)
	) name23857 (
		_w25748_,
		_w25751_,
		_w25754_,
		_w25757_,
		_w25758_
	);
	LUT3 #(
		.INIT('h2a)
	) name23858 (
		\m3_addr_i[3]_pad ,
		_w8782_,
		_w8783_,
		_w25759_
	);
	LUT3 #(
		.INIT('h80)
	) name23859 (
		\m4_addr_i[3]_pad ,
		_w8782_,
		_w8783_,
		_w25760_
	);
	LUT4 #(
		.INIT('h9dbf)
	) name23860 (
		_w8777_,
		_w8780_,
		_w25759_,
		_w25760_,
		_w25761_
	);
	LUT3 #(
		.INIT('h80)
	) name23861 (
		\m6_addr_i[3]_pad ,
		_w8782_,
		_w8783_,
		_w25762_
	);
	LUT3 #(
		.INIT('h80)
	) name23862 (
		\m2_addr_i[3]_pad ,
		_w8782_,
		_w8783_,
		_w25763_
	);
	LUT4 #(
		.INIT('habef)
	) name23863 (
		_w8777_,
		_w8780_,
		_w25762_,
		_w25763_,
		_w25764_
	);
	LUT3 #(
		.INIT('h2a)
	) name23864 (
		\m5_addr_i[3]_pad ,
		_w8782_,
		_w8783_,
		_w25765_
	);
	LUT3 #(
		.INIT('h2a)
	) name23865 (
		\m1_addr_i[3]_pad ,
		_w8782_,
		_w8783_,
		_w25766_
	);
	LUT4 #(
		.INIT('h57df)
	) name23866 (
		_w8777_,
		_w8780_,
		_w25765_,
		_w25766_,
		_w25767_
	);
	LUT3 #(
		.INIT('h80)
	) name23867 (
		\m0_addr_i[3]_pad ,
		_w8782_,
		_w8783_,
		_w25768_
	);
	LUT3 #(
		.INIT('h2a)
	) name23868 (
		\m7_addr_i[3]_pad ,
		_w8782_,
		_w8783_,
		_w25769_
	);
	LUT4 #(
		.INIT('h6e7f)
	) name23869 (
		_w8777_,
		_w8780_,
		_w25768_,
		_w25769_,
		_w25770_
	);
	LUT4 #(
		.INIT('h7fff)
	) name23870 (
		_w25761_,
		_w25764_,
		_w25767_,
		_w25770_,
		_w25771_
	);
	LUT3 #(
		.INIT('h2a)
	) name23871 (
		\m3_addr_i[4]_pad ,
		_w8782_,
		_w8783_,
		_w25772_
	);
	LUT3 #(
		.INIT('h80)
	) name23872 (
		\m4_addr_i[4]_pad ,
		_w8782_,
		_w8783_,
		_w25773_
	);
	LUT4 #(
		.INIT('h9dbf)
	) name23873 (
		_w8777_,
		_w8780_,
		_w25772_,
		_w25773_,
		_w25774_
	);
	LUT3 #(
		.INIT('h80)
	) name23874 (
		\m6_addr_i[4]_pad ,
		_w8782_,
		_w8783_,
		_w25775_
	);
	LUT3 #(
		.INIT('h80)
	) name23875 (
		\m2_addr_i[4]_pad ,
		_w8782_,
		_w8783_,
		_w25776_
	);
	LUT4 #(
		.INIT('habef)
	) name23876 (
		_w8777_,
		_w8780_,
		_w25775_,
		_w25776_,
		_w25777_
	);
	LUT3 #(
		.INIT('h2a)
	) name23877 (
		\m5_addr_i[4]_pad ,
		_w8782_,
		_w8783_,
		_w25778_
	);
	LUT3 #(
		.INIT('h2a)
	) name23878 (
		\m1_addr_i[4]_pad ,
		_w8782_,
		_w8783_,
		_w25779_
	);
	LUT4 #(
		.INIT('h57df)
	) name23879 (
		_w8777_,
		_w8780_,
		_w25778_,
		_w25779_,
		_w25780_
	);
	LUT3 #(
		.INIT('h80)
	) name23880 (
		\m0_addr_i[4]_pad ,
		_w8782_,
		_w8783_,
		_w25781_
	);
	LUT3 #(
		.INIT('h2a)
	) name23881 (
		\m7_addr_i[4]_pad ,
		_w8782_,
		_w8783_,
		_w25782_
	);
	LUT4 #(
		.INIT('h6e7f)
	) name23882 (
		_w8777_,
		_w8780_,
		_w25781_,
		_w25782_,
		_w25783_
	);
	LUT4 #(
		.INIT('h7fff)
	) name23883 (
		_w25774_,
		_w25777_,
		_w25780_,
		_w25783_,
		_w25784_
	);
	LUT3 #(
		.INIT('h2a)
	) name23884 (
		\m3_addr_i[5]_pad ,
		_w8782_,
		_w8783_,
		_w25785_
	);
	LUT3 #(
		.INIT('h80)
	) name23885 (
		\m4_addr_i[5]_pad ,
		_w8782_,
		_w8783_,
		_w25786_
	);
	LUT4 #(
		.INIT('h9dbf)
	) name23886 (
		_w8777_,
		_w8780_,
		_w25785_,
		_w25786_,
		_w25787_
	);
	LUT3 #(
		.INIT('h80)
	) name23887 (
		\m6_addr_i[5]_pad ,
		_w8782_,
		_w8783_,
		_w25788_
	);
	LUT3 #(
		.INIT('h80)
	) name23888 (
		\m2_addr_i[5]_pad ,
		_w8782_,
		_w8783_,
		_w25789_
	);
	LUT4 #(
		.INIT('habef)
	) name23889 (
		_w8777_,
		_w8780_,
		_w25788_,
		_w25789_,
		_w25790_
	);
	LUT3 #(
		.INIT('h2a)
	) name23890 (
		\m5_addr_i[5]_pad ,
		_w8782_,
		_w8783_,
		_w25791_
	);
	LUT3 #(
		.INIT('h2a)
	) name23891 (
		\m1_addr_i[5]_pad ,
		_w8782_,
		_w8783_,
		_w25792_
	);
	LUT4 #(
		.INIT('h57df)
	) name23892 (
		_w8777_,
		_w8780_,
		_w25791_,
		_w25792_,
		_w25793_
	);
	LUT3 #(
		.INIT('h80)
	) name23893 (
		\m0_addr_i[5]_pad ,
		_w8782_,
		_w8783_,
		_w25794_
	);
	LUT3 #(
		.INIT('h2a)
	) name23894 (
		\m7_addr_i[5]_pad ,
		_w8782_,
		_w8783_,
		_w25795_
	);
	LUT4 #(
		.INIT('h6e7f)
	) name23895 (
		_w8777_,
		_w8780_,
		_w25794_,
		_w25795_,
		_w25796_
	);
	LUT4 #(
		.INIT('h7fff)
	) name23896 (
		_w25787_,
		_w25790_,
		_w25793_,
		_w25796_,
		_w25797_
	);
	LUT3 #(
		.INIT('h2a)
	) name23897 (
		\m1_addr_i[6]_pad ,
		_w8782_,
		_w8783_,
		_w25798_
	);
	LUT3 #(
		.INIT('h80)
	) name23898 (
		\m2_addr_i[6]_pad ,
		_w8782_,
		_w8783_,
		_w25799_
	);
	LUT4 #(
		.INIT('h3b7f)
	) name23899 (
		_w8777_,
		_w8780_,
		_w25798_,
		_w25799_,
		_w25800_
	);
	LUT3 #(
		.INIT('h80)
	) name23900 (
		\m6_addr_i[6]_pad ,
		_w8782_,
		_w8783_,
		_w25801_
	);
	LUT3 #(
		.INIT('h2a)
	) name23901 (
		\m7_addr_i[6]_pad ,
		_w8782_,
		_w8783_,
		_w25802_
	);
	LUT3 #(
		.INIT('h57)
	) name23902 (
		_w8781_,
		_w25801_,
		_w25802_,
		_w25803_
	);
	LUT3 #(
		.INIT('h2a)
	) name23903 (
		\m5_addr_i[6]_pad ,
		_w8782_,
		_w8783_,
		_w25804_
	);
	LUT3 #(
		.INIT('h80)
	) name23904 (
		\m0_addr_i[6]_pad ,
		_w8782_,
		_w8783_,
		_w25805_
	);
	LUT4 #(
		.INIT('h57df)
	) name23905 (
		_w8777_,
		_w8780_,
		_w25804_,
		_w25805_,
		_w25806_
	);
	LUT3 #(
		.INIT('h2a)
	) name23906 (
		\m3_addr_i[6]_pad ,
		_w8782_,
		_w8783_,
		_w25807_
	);
	LUT3 #(
		.INIT('h80)
	) name23907 (
		\m4_addr_i[6]_pad ,
		_w8782_,
		_w8783_,
		_w25808_
	);
	LUT4 #(
		.INIT('h9dbf)
	) name23908 (
		_w8777_,
		_w8780_,
		_w25807_,
		_w25808_,
		_w25809_
	);
	LUT4 #(
		.INIT('h7fff)
	) name23909 (
		_w25800_,
		_w25803_,
		_w25806_,
		_w25809_,
		_w25810_
	);
	LUT3 #(
		.INIT('h2a)
	) name23910 (
		\m1_addr_i[7]_pad ,
		_w8782_,
		_w8783_,
		_w25811_
	);
	LUT3 #(
		.INIT('h80)
	) name23911 (
		\m2_addr_i[7]_pad ,
		_w8782_,
		_w8783_,
		_w25812_
	);
	LUT4 #(
		.INIT('h3b7f)
	) name23912 (
		_w8777_,
		_w8780_,
		_w25811_,
		_w25812_,
		_w25813_
	);
	LUT3 #(
		.INIT('h80)
	) name23913 (
		\m6_addr_i[7]_pad ,
		_w8782_,
		_w8783_,
		_w25814_
	);
	LUT3 #(
		.INIT('h80)
	) name23914 (
		\m4_addr_i[7]_pad ,
		_w8782_,
		_w8783_,
		_w25815_
	);
	LUT4 #(
		.INIT('hcdef)
	) name23915 (
		_w8777_,
		_w8780_,
		_w25814_,
		_w25815_,
		_w25816_
	);
	LUT3 #(
		.INIT('h2a)
	) name23916 (
		\m5_addr_i[7]_pad ,
		_w8782_,
		_w8783_,
		_w25817_
	);
	LUT3 #(
		.INIT('h2a)
	) name23917 (
		\m3_addr_i[7]_pad ,
		_w8782_,
		_w8783_,
		_w25818_
	);
	LUT4 #(
		.INIT('h9bdf)
	) name23918 (
		_w8777_,
		_w8780_,
		_w25817_,
		_w25818_,
		_w25819_
	);
	LUT3 #(
		.INIT('h80)
	) name23919 (
		\m0_addr_i[7]_pad ,
		_w8782_,
		_w8783_,
		_w25820_
	);
	LUT3 #(
		.INIT('h2a)
	) name23920 (
		\m7_addr_i[7]_pad ,
		_w8782_,
		_w8783_,
		_w25821_
	);
	LUT4 #(
		.INIT('h6e7f)
	) name23921 (
		_w8777_,
		_w8780_,
		_w25820_,
		_w25821_,
		_w25822_
	);
	LUT4 #(
		.INIT('h7fff)
	) name23922 (
		_w25813_,
		_w25816_,
		_w25819_,
		_w25822_,
		_w25823_
	);
	LUT3 #(
		.INIT('h2a)
	) name23923 (
		\m3_addr_i[8]_pad ,
		_w8782_,
		_w8783_,
		_w25824_
	);
	LUT3 #(
		.INIT('h80)
	) name23924 (
		\m4_addr_i[8]_pad ,
		_w8782_,
		_w8783_,
		_w25825_
	);
	LUT4 #(
		.INIT('h9dbf)
	) name23925 (
		_w8777_,
		_w8780_,
		_w25824_,
		_w25825_,
		_w25826_
	);
	LUT3 #(
		.INIT('h80)
	) name23926 (
		\m6_addr_i[8]_pad ,
		_w8782_,
		_w8783_,
		_w25827_
	);
	LUT3 #(
		.INIT('h80)
	) name23927 (
		\m2_addr_i[8]_pad ,
		_w8782_,
		_w8783_,
		_w25828_
	);
	LUT4 #(
		.INIT('habef)
	) name23928 (
		_w8777_,
		_w8780_,
		_w25827_,
		_w25828_,
		_w25829_
	);
	LUT3 #(
		.INIT('h2a)
	) name23929 (
		\m5_addr_i[8]_pad ,
		_w8782_,
		_w8783_,
		_w25830_
	);
	LUT3 #(
		.INIT('h2a)
	) name23930 (
		\m1_addr_i[8]_pad ,
		_w8782_,
		_w8783_,
		_w25831_
	);
	LUT4 #(
		.INIT('h57df)
	) name23931 (
		_w8777_,
		_w8780_,
		_w25830_,
		_w25831_,
		_w25832_
	);
	LUT3 #(
		.INIT('h80)
	) name23932 (
		\m0_addr_i[8]_pad ,
		_w8782_,
		_w8783_,
		_w25833_
	);
	LUT3 #(
		.INIT('h2a)
	) name23933 (
		\m7_addr_i[8]_pad ,
		_w8782_,
		_w8783_,
		_w25834_
	);
	LUT4 #(
		.INIT('h6e7f)
	) name23934 (
		_w8777_,
		_w8780_,
		_w25833_,
		_w25834_,
		_w25835_
	);
	LUT4 #(
		.INIT('h7fff)
	) name23935 (
		_w25826_,
		_w25829_,
		_w25832_,
		_w25835_,
		_w25836_
	);
	LUT3 #(
		.INIT('h2a)
	) name23936 (
		\m1_addr_i[9]_pad ,
		_w8782_,
		_w8783_,
		_w25837_
	);
	LUT3 #(
		.INIT('h80)
	) name23937 (
		\m2_addr_i[9]_pad ,
		_w8782_,
		_w8783_,
		_w25838_
	);
	LUT4 #(
		.INIT('h3b7f)
	) name23938 (
		_w8777_,
		_w8780_,
		_w25837_,
		_w25838_,
		_w25839_
	);
	LUT3 #(
		.INIT('h80)
	) name23939 (
		\m6_addr_i[9]_pad ,
		_w8782_,
		_w8783_,
		_w25840_
	);
	LUT3 #(
		.INIT('h2a)
	) name23940 (
		\m7_addr_i[9]_pad ,
		_w8782_,
		_w8783_,
		_w25841_
	);
	LUT3 #(
		.INIT('h57)
	) name23941 (
		_w8781_,
		_w25840_,
		_w25841_,
		_w25842_
	);
	LUT3 #(
		.INIT('h2a)
	) name23942 (
		\m5_addr_i[9]_pad ,
		_w8782_,
		_w8783_,
		_w25843_
	);
	LUT3 #(
		.INIT('h80)
	) name23943 (
		\m0_addr_i[9]_pad ,
		_w8782_,
		_w8783_,
		_w25844_
	);
	LUT4 #(
		.INIT('h57df)
	) name23944 (
		_w8777_,
		_w8780_,
		_w25843_,
		_w25844_,
		_w25845_
	);
	LUT3 #(
		.INIT('h2a)
	) name23945 (
		\m3_addr_i[9]_pad ,
		_w8782_,
		_w8783_,
		_w25846_
	);
	LUT3 #(
		.INIT('h80)
	) name23946 (
		\m4_addr_i[9]_pad ,
		_w8782_,
		_w8783_,
		_w25847_
	);
	LUT4 #(
		.INIT('h9dbf)
	) name23947 (
		_w8777_,
		_w8780_,
		_w25846_,
		_w25847_,
		_w25848_
	);
	LUT4 #(
		.INIT('h7fff)
	) name23948 (
		_w25839_,
		_w25842_,
		_w25845_,
		_w25848_,
		_w25849_
	);
	LUT3 #(
		.INIT('h2a)
	) name23949 (
		\m3_data_i[0]_pad ,
		_w8782_,
		_w8783_,
		_w25850_
	);
	LUT3 #(
		.INIT('h80)
	) name23950 (
		\m4_data_i[0]_pad ,
		_w8782_,
		_w8783_,
		_w25851_
	);
	LUT4 #(
		.INIT('h9dbf)
	) name23951 (
		_w8777_,
		_w8780_,
		_w25850_,
		_w25851_,
		_w25852_
	);
	LUT3 #(
		.INIT('h80)
	) name23952 (
		\m6_data_i[0]_pad ,
		_w8782_,
		_w8783_,
		_w25853_
	);
	LUT3 #(
		.INIT('h80)
	) name23953 (
		\m2_data_i[0]_pad ,
		_w8782_,
		_w8783_,
		_w25854_
	);
	LUT4 #(
		.INIT('habef)
	) name23954 (
		_w8777_,
		_w8780_,
		_w25853_,
		_w25854_,
		_w25855_
	);
	LUT3 #(
		.INIT('h2a)
	) name23955 (
		\m5_data_i[0]_pad ,
		_w8782_,
		_w8783_,
		_w25856_
	);
	LUT3 #(
		.INIT('h2a)
	) name23956 (
		\m1_data_i[0]_pad ,
		_w8782_,
		_w8783_,
		_w25857_
	);
	LUT4 #(
		.INIT('h57df)
	) name23957 (
		_w8777_,
		_w8780_,
		_w25856_,
		_w25857_,
		_w25858_
	);
	LUT3 #(
		.INIT('h80)
	) name23958 (
		\m0_data_i[0]_pad ,
		_w8782_,
		_w8783_,
		_w25859_
	);
	LUT3 #(
		.INIT('h2a)
	) name23959 (
		\m7_data_i[0]_pad ,
		_w8782_,
		_w8783_,
		_w25860_
	);
	LUT4 #(
		.INIT('h6e7f)
	) name23960 (
		_w8777_,
		_w8780_,
		_w25859_,
		_w25860_,
		_w25861_
	);
	LUT4 #(
		.INIT('h7fff)
	) name23961 (
		_w25852_,
		_w25855_,
		_w25858_,
		_w25861_,
		_w25862_
	);
	LUT3 #(
		.INIT('h2a)
	) name23962 (
		\m1_data_i[10]_pad ,
		_w8782_,
		_w8783_,
		_w25863_
	);
	LUT3 #(
		.INIT('h80)
	) name23963 (
		\m2_data_i[10]_pad ,
		_w8782_,
		_w8783_,
		_w25864_
	);
	LUT4 #(
		.INIT('h3b7f)
	) name23964 (
		_w8777_,
		_w8780_,
		_w25863_,
		_w25864_,
		_w25865_
	);
	LUT3 #(
		.INIT('h2a)
	) name23965 (
		\m3_data_i[10]_pad ,
		_w8782_,
		_w8783_,
		_w25866_
	);
	LUT3 #(
		.INIT('h2a)
	) name23966 (
		\m5_data_i[10]_pad ,
		_w8782_,
		_w8783_,
		_w25867_
	);
	LUT4 #(
		.INIT('h9dbf)
	) name23967 (
		_w8777_,
		_w8780_,
		_w25866_,
		_w25867_,
		_w25868_
	);
	LUT3 #(
		.INIT('h80)
	) name23968 (
		\m4_data_i[10]_pad ,
		_w8782_,
		_w8783_,
		_w25869_
	);
	LUT3 #(
		.INIT('h80)
	) name23969 (
		\m6_data_i[10]_pad ,
		_w8782_,
		_w8783_,
		_w25870_
	);
	LUT4 #(
		.INIT('hcedf)
	) name23970 (
		_w8777_,
		_w8780_,
		_w25869_,
		_w25870_,
		_w25871_
	);
	LUT3 #(
		.INIT('h80)
	) name23971 (
		\m0_data_i[10]_pad ,
		_w8782_,
		_w8783_,
		_w25872_
	);
	LUT3 #(
		.INIT('h2a)
	) name23972 (
		\m7_data_i[10]_pad ,
		_w8782_,
		_w8783_,
		_w25873_
	);
	LUT4 #(
		.INIT('h6e7f)
	) name23973 (
		_w8777_,
		_w8780_,
		_w25872_,
		_w25873_,
		_w25874_
	);
	LUT4 #(
		.INIT('h7fff)
	) name23974 (
		_w25865_,
		_w25868_,
		_w25871_,
		_w25874_,
		_w25875_
	);
	LUT3 #(
		.INIT('h80)
	) name23975 (
		\m6_data_i[11]_pad ,
		_w8782_,
		_w8783_,
		_w25876_
	);
	LUT3 #(
		.INIT('h2a)
	) name23976 (
		\m5_data_i[11]_pad ,
		_w8782_,
		_w8783_,
		_w25877_
	);
	LUT4 #(
		.INIT('hcdef)
	) name23977 (
		_w8777_,
		_w8780_,
		_w25876_,
		_w25877_,
		_w25878_
	);
	LUT3 #(
		.INIT('h2a)
	) name23978 (
		\m3_data_i[11]_pad ,
		_w8782_,
		_w8783_,
		_w25879_
	);
	LUT3 #(
		.INIT('h80)
	) name23979 (
		\m2_data_i[11]_pad ,
		_w8782_,
		_w8783_,
		_w25880_
	);
	LUT3 #(
		.INIT('h57)
	) name23980 (
		_w8795_,
		_w25879_,
		_w25880_,
		_w25881_
	);
	LUT3 #(
		.INIT('h80)
	) name23981 (
		\m4_data_i[11]_pad ,
		_w8782_,
		_w8783_,
		_w25882_
	);
	LUT3 #(
		.INIT('h2a)
	) name23982 (
		\m1_data_i[11]_pad ,
		_w8782_,
		_w8783_,
		_w25883_
	);
	LUT4 #(
		.INIT('h57df)
	) name23983 (
		_w8777_,
		_w8780_,
		_w25882_,
		_w25883_,
		_w25884_
	);
	LUT3 #(
		.INIT('h80)
	) name23984 (
		\m0_data_i[11]_pad ,
		_w8782_,
		_w8783_,
		_w25885_
	);
	LUT3 #(
		.INIT('h2a)
	) name23985 (
		\m7_data_i[11]_pad ,
		_w8782_,
		_w8783_,
		_w25886_
	);
	LUT4 #(
		.INIT('h6e7f)
	) name23986 (
		_w8777_,
		_w8780_,
		_w25885_,
		_w25886_,
		_w25887_
	);
	LUT4 #(
		.INIT('h7fff)
	) name23987 (
		_w25878_,
		_w25881_,
		_w25884_,
		_w25887_,
		_w25888_
	);
	LUT3 #(
		.INIT('h2a)
	) name23988 (
		\m1_data_i[12]_pad ,
		_w8782_,
		_w8783_,
		_w25889_
	);
	LUT3 #(
		.INIT('h80)
	) name23989 (
		\m2_data_i[12]_pad ,
		_w8782_,
		_w8783_,
		_w25890_
	);
	LUT4 #(
		.INIT('h3b7f)
	) name23990 (
		_w8777_,
		_w8780_,
		_w25889_,
		_w25890_,
		_w25891_
	);
	LUT3 #(
		.INIT('h80)
	) name23991 (
		\m0_data_i[12]_pad ,
		_w8782_,
		_w8783_,
		_w25892_
	);
	LUT3 #(
		.INIT('h80)
	) name23992 (
		\m4_data_i[12]_pad ,
		_w8782_,
		_w8783_,
		_w25893_
	);
	LUT4 #(
		.INIT('h5d7f)
	) name23993 (
		_w8777_,
		_w8780_,
		_w25892_,
		_w25893_,
		_w25894_
	);
	LUT3 #(
		.INIT('h2a)
	) name23994 (
		\m7_data_i[12]_pad ,
		_w8782_,
		_w8783_,
		_w25895_
	);
	LUT3 #(
		.INIT('h2a)
	) name23995 (
		\m3_data_i[12]_pad ,
		_w8782_,
		_w8783_,
		_w25896_
	);
	LUT4 #(
		.INIT('habef)
	) name23996 (
		_w8777_,
		_w8780_,
		_w25895_,
		_w25896_,
		_w25897_
	);
	LUT3 #(
		.INIT('h80)
	) name23997 (
		\m6_data_i[12]_pad ,
		_w8782_,
		_w8783_,
		_w25898_
	);
	LUT3 #(
		.INIT('h2a)
	) name23998 (
		\m5_data_i[12]_pad ,
		_w8782_,
		_w8783_,
		_w25899_
	);
	LUT4 #(
		.INIT('hcdef)
	) name23999 (
		_w8777_,
		_w8780_,
		_w25898_,
		_w25899_,
		_w25900_
	);
	LUT4 #(
		.INIT('h7fff)
	) name24000 (
		_w25891_,
		_w25894_,
		_w25897_,
		_w25900_,
		_w25901_
	);
	LUT3 #(
		.INIT('h2a)
	) name24001 (
		\m1_data_i[13]_pad ,
		_w8782_,
		_w8783_,
		_w25902_
	);
	LUT3 #(
		.INIT('h80)
	) name24002 (
		\m2_data_i[13]_pad ,
		_w8782_,
		_w8783_,
		_w25903_
	);
	LUT4 #(
		.INIT('h3b7f)
	) name24003 (
		_w8777_,
		_w8780_,
		_w25902_,
		_w25903_,
		_w25904_
	);
	LUT3 #(
		.INIT('h80)
	) name24004 (
		\m0_data_i[13]_pad ,
		_w8782_,
		_w8783_,
		_w25905_
	);
	LUT3 #(
		.INIT('h80)
	) name24005 (
		\m4_data_i[13]_pad ,
		_w8782_,
		_w8783_,
		_w25906_
	);
	LUT4 #(
		.INIT('h5d7f)
	) name24006 (
		_w8777_,
		_w8780_,
		_w25905_,
		_w25906_,
		_w25907_
	);
	LUT3 #(
		.INIT('h2a)
	) name24007 (
		\m7_data_i[13]_pad ,
		_w8782_,
		_w8783_,
		_w25908_
	);
	LUT3 #(
		.INIT('h2a)
	) name24008 (
		\m3_data_i[13]_pad ,
		_w8782_,
		_w8783_,
		_w25909_
	);
	LUT4 #(
		.INIT('habef)
	) name24009 (
		_w8777_,
		_w8780_,
		_w25908_,
		_w25909_,
		_w25910_
	);
	LUT3 #(
		.INIT('h80)
	) name24010 (
		\m6_data_i[13]_pad ,
		_w8782_,
		_w8783_,
		_w25911_
	);
	LUT3 #(
		.INIT('h2a)
	) name24011 (
		\m5_data_i[13]_pad ,
		_w8782_,
		_w8783_,
		_w25912_
	);
	LUT4 #(
		.INIT('hcdef)
	) name24012 (
		_w8777_,
		_w8780_,
		_w25911_,
		_w25912_,
		_w25913_
	);
	LUT4 #(
		.INIT('h7fff)
	) name24013 (
		_w25904_,
		_w25907_,
		_w25910_,
		_w25913_,
		_w25914_
	);
	LUT3 #(
		.INIT('h2a)
	) name24014 (
		\m1_data_i[14]_pad ,
		_w8782_,
		_w8783_,
		_w25915_
	);
	LUT3 #(
		.INIT('h80)
	) name24015 (
		\m2_data_i[14]_pad ,
		_w8782_,
		_w8783_,
		_w25916_
	);
	LUT4 #(
		.INIT('h3b7f)
	) name24016 (
		_w8777_,
		_w8780_,
		_w25915_,
		_w25916_,
		_w25917_
	);
	LUT3 #(
		.INIT('h80)
	) name24017 (
		\m0_data_i[14]_pad ,
		_w8782_,
		_w8783_,
		_w25918_
	);
	LUT3 #(
		.INIT('h80)
	) name24018 (
		\m4_data_i[14]_pad ,
		_w8782_,
		_w8783_,
		_w25919_
	);
	LUT4 #(
		.INIT('h5d7f)
	) name24019 (
		_w8777_,
		_w8780_,
		_w25918_,
		_w25919_,
		_w25920_
	);
	LUT3 #(
		.INIT('h2a)
	) name24020 (
		\m7_data_i[14]_pad ,
		_w8782_,
		_w8783_,
		_w25921_
	);
	LUT3 #(
		.INIT('h2a)
	) name24021 (
		\m3_data_i[14]_pad ,
		_w8782_,
		_w8783_,
		_w25922_
	);
	LUT4 #(
		.INIT('habef)
	) name24022 (
		_w8777_,
		_w8780_,
		_w25921_,
		_w25922_,
		_w25923_
	);
	LUT3 #(
		.INIT('h80)
	) name24023 (
		\m6_data_i[14]_pad ,
		_w8782_,
		_w8783_,
		_w25924_
	);
	LUT3 #(
		.INIT('h2a)
	) name24024 (
		\m5_data_i[14]_pad ,
		_w8782_,
		_w8783_,
		_w25925_
	);
	LUT4 #(
		.INIT('hcdef)
	) name24025 (
		_w8777_,
		_w8780_,
		_w25924_,
		_w25925_,
		_w25926_
	);
	LUT4 #(
		.INIT('h7fff)
	) name24026 (
		_w25917_,
		_w25920_,
		_w25923_,
		_w25926_,
		_w25927_
	);
	LUT3 #(
		.INIT('h2a)
	) name24027 (
		\m1_data_i[15]_pad ,
		_w8782_,
		_w8783_,
		_w25928_
	);
	LUT3 #(
		.INIT('h80)
	) name24028 (
		\m2_data_i[15]_pad ,
		_w8782_,
		_w8783_,
		_w25929_
	);
	LUT4 #(
		.INIT('h3b7f)
	) name24029 (
		_w8777_,
		_w8780_,
		_w25928_,
		_w25929_,
		_w25930_
	);
	LUT3 #(
		.INIT('h80)
	) name24030 (
		\m0_data_i[15]_pad ,
		_w8782_,
		_w8783_,
		_w25931_
	);
	LUT3 #(
		.INIT('h80)
	) name24031 (
		\m4_data_i[15]_pad ,
		_w8782_,
		_w8783_,
		_w25932_
	);
	LUT4 #(
		.INIT('h5d7f)
	) name24032 (
		_w8777_,
		_w8780_,
		_w25931_,
		_w25932_,
		_w25933_
	);
	LUT3 #(
		.INIT('h2a)
	) name24033 (
		\m7_data_i[15]_pad ,
		_w8782_,
		_w8783_,
		_w25934_
	);
	LUT3 #(
		.INIT('h2a)
	) name24034 (
		\m3_data_i[15]_pad ,
		_w8782_,
		_w8783_,
		_w25935_
	);
	LUT4 #(
		.INIT('habef)
	) name24035 (
		_w8777_,
		_w8780_,
		_w25934_,
		_w25935_,
		_w25936_
	);
	LUT3 #(
		.INIT('h80)
	) name24036 (
		\m6_data_i[15]_pad ,
		_w8782_,
		_w8783_,
		_w25937_
	);
	LUT3 #(
		.INIT('h2a)
	) name24037 (
		\m5_data_i[15]_pad ,
		_w8782_,
		_w8783_,
		_w25938_
	);
	LUT4 #(
		.INIT('hcdef)
	) name24038 (
		_w8777_,
		_w8780_,
		_w25937_,
		_w25938_,
		_w25939_
	);
	LUT4 #(
		.INIT('h7fff)
	) name24039 (
		_w25930_,
		_w25933_,
		_w25936_,
		_w25939_,
		_w25940_
	);
	LUT3 #(
		.INIT('h2a)
	) name24040 (
		\m3_data_i[16]_pad ,
		_w8782_,
		_w8783_,
		_w25941_
	);
	LUT3 #(
		.INIT('h80)
	) name24041 (
		\m4_data_i[16]_pad ,
		_w8782_,
		_w8783_,
		_w25942_
	);
	LUT4 #(
		.INIT('h9dbf)
	) name24042 (
		_w8777_,
		_w8780_,
		_w25941_,
		_w25942_,
		_w25943_
	);
	LUT3 #(
		.INIT('h80)
	) name24043 (
		\m0_data_i[16]_pad ,
		_w8782_,
		_w8783_,
		_w25944_
	);
	LUT3 #(
		.INIT('h2a)
	) name24044 (
		\m5_data_i[16]_pad ,
		_w8782_,
		_w8783_,
		_w25945_
	);
	LUT4 #(
		.INIT('h5d7f)
	) name24045 (
		_w8777_,
		_w8780_,
		_w25944_,
		_w25945_,
		_w25946_
	);
	LUT3 #(
		.INIT('h2a)
	) name24046 (
		\m7_data_i[16]_pad ,
		_w8782_,
		_w8783_,
		_w25947_
	);
	LUT3 #(
		.INIT('h80)
	) name24047 (
		\m6_data_i[16]_pad ,
		_w8782_,
		_w8783_,
		_w25948_
	);
	LUT3 #(
		.INIT('h57)
	) name24048 (
		_w8781_,
		_w25947_,
		_w25948_,
		_w25949_
	);
	LUT3 #(
		.INIT('h2a)
	) name24049 (
		\m1_data_i[16]_pad ,
		_w8782_,
		_w8783_,
		_w25950_
	);
	LUT3 #(
		.INIT('h80)
	) name24050 (
		\m2_data_i[16]_pad ,
		_w8782_,
		_w8783_,
		_w25951_
	);
	LUT4 #(
		.INIT('h3b7f)
	) name24051 (
		_w8777_,
		_w8780_,
		_w25950_,
		_w25951_,
		_w25952_
	);
	LUT4 #(
		.INIT('h7fff)
	) name24052 (
		_w25943_,
		_w25946_,
		_w25949_,
		_w25952_,
		_w25953_
	);
	LUT3 #(
		.INIT('h2a)
	) name24053 (
		\m1_data_i[17]_pad ,
		_w8782_,
		_w8783_,
		_w25954_
	);
	LUT3 #(
		.INIT('h80)
	) name24054 (
		\m2_data_i[17]_pad ,
		_w8782_,
		_w8783_,
		_w25955_
	);
	LUT4 #(
		.INIT('h3b7f)
	) name24055 (
		_w8777_,
		_w8780_,
		_w25954_,
		_w25955_,
		_w25956_
	);
	LUT3 #(
		.INIT('h80)
	) name24056 (
		\m6_data_i[17]_pad ,
		_w8782_,
		_w8783_,
		_w25957_
	);
	LUT3 #(
		.INIT('h2a)
	) name24057 (
		\m7_data_i[17]_pad ,
		_w8782_,
		_w8783_,
		_w25958_
	);
	LUT3 #(
		.INIT('h57)
	) name24058 (
		_w8781_,
		_w25957_,
		_w25958_,
		_w25959_
	);
	LUT3 #(
		.INIT('h2a)
	) name24059 (
		\m5_data_i[17]_pad ,
		_w8782_,
		_w8783_,
		_w25960_
	);
	LUT3 #(
		.INIT('h80)
	) name24060 (
		\m0_data_i[17]_pad ,
		_w8782_,
		_w8783_,
		_w25961_
	);
	LUT4 #(
		.INIT('h57df)
	) name24061 (
		_w8777_,
		_w8780_,
		_w25960_,
		_w25961_,
		_w25962_
	);
	LUT3 #(
		.INIT('h2a)
	) name24062 (
		\m3_data_i[17]_pad ,
		_w8782_,
		_w8783_,
		_w25963_
	);
	LUT3 #(
		.INIT('h80)
	) name24063 (
		\m4_data_i[17]_pad ,
		_w8782_,
		_w8783_,
		_w25964_
	);
	LUT4 #(
		.INIT('h9dbf)
	) name24064 (
		_w8777_,
		_w8780_,
		_w25963_,
		_w25964_,
		_w25965_
	);
	LUT4 #(
		.INIT('h7fff)
	) name24065 (
		_w25956_,
		_w25959_,
		_w25962_,
		_w25965_,
		_w25966_
	);
	LUT3 #(
		.INIT('h2a)
	) name24066 (
		\m3_data_i[18]_pad ,
		_w8782_,
		_w8783_,
		_w25967_
	);
	LUT3 #(
		.INIT('h80)
	) name24067 (
		\m4_data_i[18]_pad ,
		_w8782_,
		_w8783_,
		_w25968_
	);
	LUT4 #(
		.INIT('h9dbf)
	) name24068 (
		_w8777_,
		_w8780_,
		_w25967_,
		_w25968_,
		_w25969_
	);
	LUT3 #(
		.INIT('h80)
	) name24069 (
		\m6_data_i[18]_pad ,
		_w8782_,
		_w8783_,
		_w25970_
	);
	LUT3 #(
		.INIT('h80)
	) name24070 (
		\m2_data_i[18]_pad ,
		_w8782_,
		_w8783_,
		_w25971_
	);
	LUT4 #(
		.INIT('habef)
	) name24071 (
		_w8777_,
		_w8780_,
		_w25970_,
		_w25971_,
		_w25972_
	);
	LUT3 #(
		.INIT('h2a)
	) name24072 (
		\m5_data_i[18]_pad ,
		_w8782_,
		_w8783_,
		_w25973_
	);
	LUT3 #(
		.INIT('h2a)
	) name24073 (
		\m1_data_i[18]_pad ,
		_w8782_,
		_w8783_,
		_w25974_
	);
	LUT4 #(
		.INIT('h57df)
	) name24074 (
		_w8777_,
		_w8780_,
		_w25973_,
		_w25974_,
		_w25975_
	);
	LUT3 #(
		.INIT('h80)
	) name24075 (
		\m0_data_i[18]_pad ,
		_w8782_,
		_w8783_,
		_w25976_
	);
	LUT3 #(
		.INIT('h2a)
	) name24076 (
		\m7_data_i[18]_pad ,
		_w8782_,
		_w8783_,
		_w25977_
	);
	LUT4 #(
		.INIT('h6e7f)
	) name24077 (
		_w8777_,
		_w8780_,
		_w25976_,
		_w25977_,
		_w25978_
	);
	LUT4 #(
		.INIT('h7fff)
	) name24078 (
		_w25969_,
		_w25972_,
		_w25975_,
		_w25978_,
		_w25979_
	);
	LUT3 #(
		.INIT('h2a)
	) name24079 (
		\m1_data_i[19]_pad ,
		_w8782_,
		_w8783_,
		_w25980_
	);
	LUT3 #(
		.INIT('h80)
	) name24080 (
		\m2_data_i[19]_pad ,
		_w8782_,
		_w8783_,
		_w25981_
	);
	LUT4 #(
		.INIT('h3b7f)
	) name24081 (
		_w8777_,
		_w8780_,
		_w25980_,
		_w25981_,
		_w25982_
	);
	LUT3 #(
		.INIT('h2a)
	) name24082 (
		\m3_data_i[19]_pad ,
		_w8782_,
		_w8783_,
		_w25983_
	);
	LUT3 #(
		.INIT('h2a)
	) name24083 (
		\m7_data_i[19]_pad ,
		_w8782_,
		_w8783_,
		_w25984_
	);
	LUT4 #(
		.INIT('haebf)
	) name24084 (
		_w8777_,
		_w8780_,
		_w25983_,
		_w25984_,
		_w25985_
	);
	LUT3 #(
		.INIT('h80)
	) name24085 (
		\m4_data_i[19]_pad ,
		_w8782_,
		_w8783_,
		_w25986_
	);
	LUT3 #(
		.INIT('h80)
	) name24086 (
		\m0_data_i[19]_pad ,
		_w8782_,
		_w8783_,
		_w25987_
	);
	LUT4 #(
		.INIT('h57df)
	) name24087 (
		_w8777_,
		_w8780_,
		_w25986_,
		_w25987_,
		_w25988_
	);
	LUT3 #(
		.INIT('h80)
	) name24088 (
		\m6_data_i[19]_pad ,
		_w8782_,
		_w8783_,
		_w25989_
	);
	LUT3 #(
		.INIT('h2a)
	) name24089 (
		\m5_data_i[19]_pad ,
		_w8782_,
		_w8783_,
		_w25990_
	);
	LUT4 #(
		.INIT('hcdef)
	) name24090 (
		_w8777_,
		_w8780_,
		_w25989_,
		_w25990_,
		_w25991_
	);
	LUT4 #(
		.INIT('h7fff)
	) name24091 (
		_w25982_,
		_w25985_,
		_w25988_,
		_w25991_,
		_w25992_
	);
	LUT3 #(
		.INIT('h80)
	) name24092 (
		\m0_data_i[1]_pad ,
		_w8782_,
		_w8783_,
		_w25993_
	);
	LUT3 #(
		.INIT('h2a)
	) name24093 (
		\m7_data_i[1]_pad ,
		_w8782_,
		_w8783_,
		_w25994_
	);
	LUT4 #(
		.INIT('h6e7f)
	) name24094 (
		_w8777_,
		_w8780_,
		_w25993_,
		_w25994_,
		_w25995_
	);
	LUT3 #(
		.INIT('h2a)
	) name24095 (
		\m1_data_i[1]_pad ,
		_w8782_,
		_w8783_,
		_w25996_
	);
	LUT3 #(
		.INIT('h80)
	) name24096 (
		\m4_data_i[1]_pad ,
		_w8782_,
		_w8783_,
		_w25997_
	);
	LUT4 #(
		.INIT('h5d7f)
	) name24097 (
		_w8777_,
		_w8780_,
		_w25996_,
		_w25997_,
		_w25998_
	);
	LUT3 #(
		.INIT('h80)
	) name24098 (
		\m2_data_i[1]_pad ,
		_w8782_,
		_w8783_,
		_w25999_
	);
	LUT3 #(
		.INIT('h2a)
	) name24099 (
		\m3_data_i[1]_pad ,
		_w8782_,
		_w8783_,
		_w26000_
	);
	LUT3 #(
		.INIT('h57)
	) name24100 (
		_w8795_,
		_w25999_,
		_w26000_,
		_w26001_
	);
	LUT3 #(
		.INIT('h80)
	) name24101 (
		\m6_data_i[1]_pad ,
		_w8782_,
		_w8783_,
		_w26002_
	);
	LUT3 #(
		.INIT('h2a)
	) name24102 (
		\m5_data_i[1]_pad ,
		_w8782_,
		_w8783_,
		_w26003_
	);
	LUT4 #(
		.INIT('hcdef)
	) name24103 (
		_w8777_,
		_w8780_,
		_w26002_,
		_w26003_,
		_w26004_
	);
	LUT4 #(
		.INIT('h7fff)
	) name24104 (
		_w25995_,
		_w25998_,
		_w26001_,
		_w26004_,
		_w26005_
	);
	LUT3 #(
		.INIT('h2a)
	) name24105 (
		\m1_data_i[20]_pad ,
		_w8782_,
		_w8783_,
		_w26006_
	);
	LUT3 #(
		.INIT('h80)
	) name24106 (
		\m2_data_i[20]_pad ,
		_w8782_,
		_w8783_,
		_w26007_
	);
	LUT4 #(
		.INIT('h3b7f)
	) name24107 (
		_w8777_,
		_w8780_,
		_w26006_,
		_w26007_,
		_w26008_
	);
	LUT3 #(
		.INIT('h80)
	) name24108 (
		\m0_data_i[20]_pad ,
		_w8782_,
		_w8783_,
		_w26009_
	);
	LUT3 #(
		.INIT('h80)
	) name24109 (
		\m4_data_i[20]_pad ,
		_w8782_,
		_w8783_,
		_w26010_
	);
	LUT4 #(
		.INIT('h5d7f)
	) name24110 (
		_w8777_,
		_w8780_,
		_w26009_,
		_w26010_,
		_w26011_
	);
	LUT3 #(
		.INIT('h2a)
	) name24111 (
		\m7_data_i[20]_pad ,
		_w8782_,
		_w8783_,
		_w26012_
	);
	LUT3 #(
		.INIT('h2a)
	) name24112 (
		\m3_data_i[20]_pad ,
		_w8782_,
		_w8783_,
		_w26013_
	);
	LUT4 #(
		.INIT('habef)
	) name24113 (
		_w8777_,
		_w8780_,
		_w26012_,
		_w26013_,
		_w26014_
	);
	LUT3 #(
		.INIT('h80)
	) name24114 (
		\m6_data_i[20]_pad ,
		_w8782_,
		_w8783_,
		_w26015_
	);
	LUT3 #(
		.INIT('h2a)
	) name24115 (
		\m5_data_i[20]_pad ,
		_w8782_,
		_w8783_,
		_w26016_
	);
	LUT4 #(
		.INIT('hcdef)
	) name24116 (
		_w8777_,
		_w8780_,
		_w26015_,
		_w26016_,
		_w26017_
	);
	LUT4 #(
		.INIT('h7fff)
	) name24117 (
		_w26008_,
		_w26011_,
		_w26014_,
		_w26017_,
		_w26018_
	);
	LUT3 #(
		.INIT('h80)
	) name24118 (
		\m6_data_i[21]_pad ,
		_w8782_,
		_w8783_,
		_w26019_
	);
	LUT3 #(
		.INIT('h2a)
	) name24119 (
		\m5_data_i[21]_pad ,
		_w8782_,
		_w8783_,
		_w26020_
	);
	LUT4 #(
		.INIT('hcdef)
	) name24120 (
		_w8777_,
		_w8780_,
		_w26019_,
		_w26020_,
		_w26021_
	);
	LUT3 #(
		.INIT('h2a)
	) name24121 (
		\m1_data_i[21]_pad ,
		_w8782_,
		_w8783_,
		_w26022_
	);
	LUT3 #(
		.INIT('h80)
	) name24122 (
		\m4_data_i[21]_pad ,
		_w8782_,
		_w8783_,
		_w26023_
	);
	LUT4 #(
		.INIT('h5d7f)
	) name24123 (
		_w8777_,
		_w8780_,
		_w26022_,
		_w26023_,
		_w26024_
	);
	LUT3 #(
		.INIT('h80)
	) name24124 (
		\m2_data_i[21]_pad ,
		_w8782_,
		_w8783_,
		_w26025_
	);
	LUT3 #(
		.INIT('h2a)
	) name24125 (
		\m3_data_i[21]_pad ,
		_w8782_,
		_w8783_,
		_w26026_
	);
	LUT3 #(
		.INIT('h57)
	) name24126 (
		_w8795_,
		_w26025_,
		_w26026_,
		_w26027_
	);
	LUT3 #(
		.INIT('h80)
	) name24127 (
		\m0_data_i[21]_pad ,
		_w8782_,
		_w8783_,
		_w26028_
	);
	LUT3 #(
		.INIT('h2a)
	) name24128 (
		\m7_data_i[21]_pad ,
		_w8782_,
		_w8783_,
		_w26029_
	);
	LUT4 #(
		.INIT('h6e7f)
	) name24129 (
		_w8777_,
		_w8780_,
		_w26028_,
		_w26029_,
		_w26030_
	);
	LUT4 #(
		.INIT('h7fff)
	) name24130 (
		_w26021_,
		_w26024_,
		_w26027_,
		_w26030_,
		_w26031_
	);
	LUT3 #(
		.INIT('h2a)
	) name24131 (
		\m3_data_i[22]_pad ,
		_w8782_,
		_w8783_,
		_w26032_
	);
	LUT3 #(
		.INIT('h80)
	) name24132 (
		\m4_data_i[22]_pad ,
		_w8782_,
		_w8783_,
		_w26033_
	);
	LUT4 #(
		.INIT('h9dbf)
	) name24133 (
		_w8777_,
		_w8780_,
		_w26032_,
		_w26033_,
		_w26034_
	);
	LUT3 #(
		.INIT('h80)
	) name24134 (
		\m6_data_i[22]_pad ,
		_w8782_,
		_w8783_,
		_w26035_
	);
	LUT3 #(
		.INIT('h80)
	) name24135 (
		\m2_data_i[22]_pad ,
		_w8782_,
		_w8783_,
		_w26036_
	);
	LUT4 #(
		.INIT('habef)
	) name24136 (
		_w8777_,
		_w8780_,
		_w26035_,
		_w26036_,
		_w26037_
	);
	LUT3 #(
		.INIT('h2a)
	) name24137 (
		\m5_data_i[22]_pad ,
		_w8782_,
		_w8783_,
		_w26038_
	);
	LUT3 #(
		.INIT('h2a)
	) name24138 (
		\m1_data_i[22]_pad ,
		_w8782_,
		_w8783_,
		_w26039_
	);
	LUT4 #(
		.INIT('h57df)
	) name24139 (
		_w8777_,
		_w8780_,
		_w26038_,
		_w26039_,
		_w26040_
	);
	LUT3 #(
		.INIT('h80)
	) name24140 (
		\m0_data_i[22]_pad ,
		_w8782_,
		_w8783_,
		_w26041_
	);
	LUT3 #(
		.INIT('h2a)
	) name24141 (
		\m7_data_i[22]_pad ,
		_w8782_,
		_w8783_,
		_w26042_
	);
	LUT4 #(
		.INIT('h6e7f)
	) name24142 (
		_w8777_,
		_w8780_,
		_w26041_,
		_w26042_,
		_w26043_
	);
	LUT4 #(
		.INIT('h7fff)
	) name24143 (
		_w26034_,
		_w26037_,
		_w26040_,
		_w26043_,
		_w26044_
	);
	LUT3 #(
		.INIT('h80)
	) name24144 (
		\m6_data_i[23]_pad ,
		_w8782_,
		_w8783_,
		_w26045_
	);
	LUT3 #(
		.INIT('h2a)
	) name24145 (
		\m5_data_i[23]_pad ,
		_w8782_,
		_w8783_,
		_w26046_
	);
	LUT4 #(
		.INIT('hcdef)
	) name24146 (
		_w8777_,
		_w8780_,
		_w26045_,
		_w26046_,
		_w26047_
	);
	LUT3 #(
		.INIT('h2a)
	) name24147 (
		\m1_data_i[23]_pad ,
		_w8782_,
		_w8783_,
		_w26048_
	);
	LUT3 #(
		.INIT('h80)
	) name24148 (
		\m4_data_i[23]_pad ,
		_w8782_,
		_w8783_,
		_w26049_
	);
	LUT4 #(
		.INIT('h5d7f)
	) name24149 (
		_w8777_,
		_w8780_,
		_w26048_,
		_w26049_,
		_w26050_
	);
	LUT3 #(
		.INIT('h80)
	) name24150 (
		\m2_data_i[23]_pad ,
		_w8782_,
		_w8783_,
		_w26051_
	);
	LUT3 #(
		.INIT('h2a)
	) name24151 (
		\m3_data_i[23]_pad ,
		_w8782_,
		_w8783_,
		_w26052_
	);
	LUT3 #(
		.INIT('h57)
	) name24152 (
		_w8795_,
		_w26051_,
		_w26052_,
		_w26053_
	);
	LUT3 #(
		.INIT('h80)
	) name24153 (
		\m0_data_i[23]_pad ,
		_w8782_,
		_w8783_,
		_w26054_
	);
	LUT3 #(
		.INIT('h2a)
	) name24154 (
		\m7_data_i[23]_pad ,
		_w8782_,
		_w8783_,
		_w26055_
	);
	LUT4 #(
		.INIT('h6e7f)
	) name24155 (
		_w8777_,
		_w8780_,
		_w26054_,
		_w26055_,
		_w26056_
	);
	LUT4 #(
		.INIT('h7fff)
	) name24156 (
		_w26047_,
		_w26050_,
		_w26053_,
		_w26056_,
		_w26057_
	);
	LUT3 #(
		.INIT('h2a)
	) name24157 (
		\m1_data_i[24]_pad ,
		_w8782_,
		_w8783_,
		_w26058_
	);
	LUT3 #(
		.INIT('h80)
	) name24158 (
		\m2_data_i[24]_pad ,
		_w8782_,
		_w8783_,
		_w26059_
	);
	LUT4 #(
		.INIT('h3b7f)
	) name24159 (
		_w8777_,
		_w8780_,
		_w26058_,
		_w26059_,
		_w26060_
	);
	LUT3 #(
		.INIT('h80)
	) name24160 (
		\m0_data_i[24]_pad ,
		_w8782_,
		_w8783_,
		_w26061_
	);
	LUT3 #(
		.INIT('h80)
	) name24161 (
		\m4_data_i[24]_pad ,
		_w8782_,
		_w8783_,
		_w26062_
	);
	LUT4 #(
		.INIT('h5d7f)
	) name24162 (
		_w8777_,
		_w8780_,
		_w26061_,
		_w26062_,
		_w26063_
	);
	LUT3 #(
		.INIT('h2a)
	) name24163 (
		\m7_data_i[24]_pad ,
		_w8782_,
		_w8783_,
		_w26064_
	);
	LUT3 #(
		.INIT('h2a)
	) name24164 (
		\m3_data_i[24]_pad ,
		_w8782_,
		_w8783_,
		_w26065_
	);
	LUT4 #(
		.INIT('habef)
	) name24165 (
		_w8777_,
		_w8780_,
		_w26064_,
		_w26065_,
		_w26066_
	);
	LUT3 #(
		.INIT('h80)
	) name24166 (
		\m6_data_i[24]_pad ,
		_w8782_,
		_w8783_,
		_w26067_
	);
	LUT3 #(
		.INIT('h2a)
	) name24167 (
		\m5_data_i[24]_pad ,
		_w8782_,
		_w8783_,
		_w26068_
	);
	LUT4 #(
		.INIT('hcdef)
	) name24168 (
		_w8777_,
		_w8780_,
		_w26067_,
		_w26068_,
		_w26069_
	);
	LUT4 #(
		.INIT('h7fff)
	) name24169 (
		_w26060_,
		_w26063_,
		_w26066_,
		_w26069_,
		_w26070_
	);
	LUT3 #(
		.INIT('h2a)
	) name24170 (
		\m1_data_i[25]_pad ,
		_w8782_,
		_w8783_,
		_w26071_
	);
	LUT3 #(
		.INIT('h80)
	) name24171 (
		\m2_data_i[25]_pad ,
		_w8782_,
		_w8783_,
		_w26072_
	);
	LUT4 #(
		.INIT('h3b7f)
	) name24172 (
		_w8777_,
		_w8780_,
		_w26071_,
		_w26072_,
		_w26073_
	);
	LUT3 #(
		.INIT('h80)
	) name24173 (
		\m0_data_i[25]_pad ,
		_w8782_,
		_w8783_,
		_w26074_
	);
	LUT3 #(
		.INIT('h80)
	) name24174 (
		\m4_data_i[25]_pad ,
		_w8782_,
		_w8783_,
		_w26075_
	);
	LUT4 #(
		.INIT('h5d7f)
	) name24175 (
		_w8777_,
		_w8780_,
		_w26074_,
		_w26075_,
		_w26076_
	);
	LUT3 #(
		.INIT('h2a)
	) name24176 (
		\m7_data_i[25]_pad ,
		_w8782_,
		_w8783_,
		_w26077_
	);
	LUT3 #(
		.INIT('h2a)
	) name24177 (
		\m3_data_i[25]_pad ,
		_w8782_,
		_w8783_,
		_w26078_
	);
	LUT4 #(
		.INIT('habef)
	) name24178 (
		_w8777_,
		_w8780_,
		_w26077_,
		_w26078_,
		_w26079_
	);
	LUT3 #(
		.INIT('h80)
	) name24179 (
		\m6_data_i[25]_pad ,
		_w8782_,
		_w8783_,
		_w26080_
	);
	LUT3 #(
		.INIT('h2a)
	) name24180 (
		\m5_data_i[25]_pad ,
		_w8782_,
		_w8783_,
		_w26081_
	);
	LUT4 #(
		.INIT('hcdef)
	) name24181 (
		_w8777_,
		_w8780_,
		_w26080_,
		_w26081_,
		_w26082_
	);
	LUT4 #(
		.INIT('h7fff)
	) name24182 (
		_w26073_,
		_w26076_,
		_w26079_,
		_w26082_,
		_w26083_
	);
	LUT3 #(
		.INIT('h2a)
	) name24183 (
		\m1_data_i[26]_pad ,
		_w8782_,
		_w8783_,
		_w26084_
	);
	LUT3 #(
		.INIT('h80)
	) name24184 (
		\m2_data_i[26]_pad ,
		_w8782_,
		_w8783_,
		_w26085_
	);
	LUT4 #(
		.INIT('h3b7f)
	) name24185 (
		_w8777_,
		_w8780_,
		_w26084_,
		_w26085_,
		_w26086_
	);
	LUT3 #(
		.INIT('h80)
	) name24186 (
		\m6_data_i[26]_pad ,
		_w8782_,
		_w8783_,
		_w26087_
	);
	LUT3 #(
		.INIT('h2a)
	) name24187 (
		\m7_data_i[26]_pad ,
		_w8782_,
		_w8783_,
		_w26088_
	);
	LUT3 #(
		.INIT('h57)
	) name24188 (
		_w8781_,
		_w26087_,
		_w26088_,
		_w26089_
	);
	LUT3 #(
		.INIT('h2a)
	) name24189 (
		\m5_data_i[26]_pad ,
		_w8782_,
		_w8783_,
		_w26090_
	);
	LUT3 #(
		.INIT('h80)
	) name24190 (
		\m0_data_i[26]_pad ,
		_w8782_,
		_w8783_,
		_w26091_
	);
	LUT4 #(
		.INIT('h57df)
	) name24191 (
		_w8777_,
		_w8780_,
		_w26090_,
		_w26091_,
		_w26092_
	);
	LUT3 #(
		.INIT('h2a)
	) name24192 (
		\m3_data_i[26]_pad ,
		_w8782_,
		_w8783_,
		_w26093_
	);
	LUT3 #(
		.INIT('h80)
	) name24193 (
		\m4_data_i[26]_pad ,
		_w8782_,
		_w8783_,
		_w26094_
	);
	LUT4 #(
		.INIT('h9dbf)
	) name24194 (
		_w8777_,
		_w8780_,
		_w26093_,
		_w26094_,
		_w26095_
	);
	LUT4 #(
		.INIT('h7fff)
	) name24195 (
		_w26086_,
		_w26089_,
		_w26092_,
		_w26095_,
		_w26096_
	);
	LUT3 #(
		.INIT('h2a)
	) name24196 (
		\m1_data_i[27]_pad ,
		_w8782_,
		_w8783_,
		_w26097_
	);
	LUT3 #(
		.INIT('h80)
	) name24197 (
		\m2_data_i[27]_pad ,
		_w8782_,
		_w8783_,
		_w26098_
	);
	LUT4 #(
		.INIT('h3b7f)
	) name24198 (
		_w8777_,
		_w8780_,
		_w26097_,
		_w26098_,
		_w26099_
	);
	LUT3 #(
		.INIT('h80)
	) name24199 (
		\m6_data_i[27]_pad ,
		_w8782_,
		_w8783_,
		_w26100_
	);
	LUT3 #(
		.INIT('h2a)
	) name24200 (
		\m7_data_i[27]_pad ,
		_w8782_,
		_w8783_,
		_w26101_
	);
	LUT3 #(
		.INIT('h57)
	) name24201 (
		_w8781_,
		_w26100_,
		_w26101_,
		_w26102_
	);
	LUT3 #(
		.INIT('h2a)
	) name24202 (
		\m5_data_i[27]_pad ,
		_w8782_,
		_w8783_,
		_w26103_
	);
	LUT3 #(
		.INIT('h80)
	) name24203 (
		\m0_data_i[27]_pad ,
		_w8782_,
		_w8783_,
		_w26104_
	);
	LUT4 #(
		.INIT('h57df)
	) name24204 (
		_w8777_,
		_w8780_,
		_w26103_,
		_w26104_,
		_w26105_
	);
	LUT3 #(
		.INIT('h2a)
	) name24205 (
		\m3_data_i[27]_pad ,
		_w8782_,
		_w8783_,
		_w26106_
	);
	LUT3 #(
		.INIT('h80)
	) name24206 (
		\m4_data_i[27]_pad ,
		_w8782_,
		_w8783_,
		_w26107_
	);
	LUT4 #(
		.INIT('h9dbf)
	) name24207 (
		_w8777_,
		_w8780_,
		_w26106_,
		_w26107_,
		_w26108_
	);
	LUT4 #(
		.INIT('h7fff)
	) name24208 (
		_w26099_,
		_w26102_,
		_w26105_,
		_w26108_,
		_w26109_
	);
	LUT3 #(
		.INIT('h2a)
	) name24209 (
		\m3_data_i[28]_pad ,
		_w8782_,
		_w8783_,
		_w26110_
	);
	LUT3 #(
		.INIT('h80)
	) name24210 (
		\m4_data_i[28]_pad ,
		_w8782_,
		_w8783_,
		_w26111_
	);
	LUT4 #(
		.INIT('h9dbf)
	) name24211 (
		_w8777_,
		_w8780_,
		_w26110_,
		_w26111_,
		_w26112_
	);
	LUT3 #(
		.INIT('h80)
	) name24212 (
		\m6_data_i[28]_pad ,
		_w8782_,
		_w8783_,
		_w26113_
	);
	LUT3 #(
		.INIT('h2a)
	) name24213 (
		\m7_data_i[28]_pad ,
		_w8782_,
		_w8783_,
		_w26114_
	);
	LUT3 #(
		.INIT('h57)
	) name24214 (
		_w8781_,
		_w26113_,
		_w26114_,
		_w26115_
	);
	LUT3 #(
		.INIT('h2a)
	) name24215 (
		\m5_data_i[28]_pad ,
		_w8782_,
		_w8783_,
		_w26116_
	);
	LUT3 #(
		.INIT('h80)
	) name24216 (
		\m0_data_i[28]_pad ,
		_w8782_,
		_w8783_,
		_w26117_
	);
	LUT4 #(
		.INIT('h57df)
	) name24217 (
		_w8777_,
		_w8780_,
		_w26116_,
		_w26117_,
		_w26118_
	);
	LUT3 #(
		.INIT('h2a)
	) name24218 (
		\m1_data_i[28]_pad ,
		_w8782_,
		_w8783_,
		_w26119_
	);
	LUT3 #(
		.INIT('h80)
	) name24219 (
		\m2_data_i[28]_pad ,
		_w8782_,
		_w8783_,
		_w26120_
	);
	LUT4 #(
		.INIT('h3b7f)
	) name24220 (
		_w8777_,
		_w8780_,
		_w26119_,
		_w26120_,
		_w26121_
	);
	LUT4 #(
		.INIT('h7fff)
	) name24221 (
		_w26112_,
		_w26115_,
		_w26118_,
		_w26121_,
		_w26122_
	);
	LUT3 #(
		.INIT('h2a)
	) name24222 (
		\m1_data_i[29]_pad ,
		_w8782_,
		_w8783_,
		_w26123_
	);
	LUT3 #(
		.INIT('h80)
	) name24223 (
		\m2_data_i[29]_pad ,
		_w8782_,
		_w8783_,
		_w26124_
	);
	LUT4 #(
		.INIT('h3b7f)
	) name24224 (
		_w8777_,
		_w8780_,
		_w26123_,
		_w26124_,
		_w26125_
	);
	LUT3 #(
		.INIT('h2a)
	) name24225 (
		\m3_data_i[29]_pad ,
		_w8782_,
		_w8783_,
		_w26126_
	);
	LUT3 #(
		.INIT('h2a)
	) name24226 (
		\m7_data_i[29]_pad ,
		_w8782_,
		_w8783_,
		_w26127_
	);
	LUT4 #(
		.INIT('haebf)
	) name24227 (
		_w8777_,
		_w8780_,
		_w26126_,
		_w26127_,
		_w26128_
	);
	LUT3 #(
		.INIT('h80)
	) name24228 (
		\m4_data_i[29]_pad ,
		_w8782_,
		_w8783_,
		_w26129_
	);
	LUT3 #(
		.INIT('h80)
	) name24229 (
		\m0_data_i[29]_pad ,
		_w8782_,
		_w8783_,
		_w26130_
	);
	LUT4 #(
		.INIT('h57df)
	) name24230 (
		_w8777_,
		_w8780_,
		_w26129_,
		_w26130_,
		_w26131_
	);
	LUT3 #(
		.INIT('h80)
	) name24231 (
		\m6_data_i[29]_pad ,
		_w8782_,
		_w8783_,
		_w26132_
	);
	LUT3 #(
		.INIT('h2a)
	) name24232 (
		\m5_data_i[29]_pad ,
		_w8782_,
		_w8783_,
		_w26133_
	);
	LUT4 #(
		.INIT('hcdef)
	) name24233 (
		_w8777_,
		_w8780_,
		_w26132_,
		_w26133_,
		_w26134_
	);
	LUT4 #(
		.INIT('h7fff)
	) name24234 (
		_w26125_,
		_w26128_,
		_w26131_,
		_w26134_,
		_w26135_
	);
	LUT3 #(
		.INIT('h2a)
	) name24235 (
		\m1_data_i[2]_pad ,
		_w8782_,
		_w8783_,
		_w26136_
	);
	LUT3 #(
		.INIT('h80)
	) name24236 (
		\m2_data_i[2]_pad ,
		_w8782_,
		_w8783_,
		_w26137_
	);
	LUT4 #(
		.INIT('h3b7f)
	) name24237 (
		_w8777_,
		_w8780_,
		_w26136_,
		_w26137_,
		_w26138_
	);
	LUT3 #(
		.INIT('h80)
	) name24238 (
		\m0_data_i[2]_pad ,
		_w8782_,
		_w8783_,
		_w26139_
	);
	LUT3 #(
		.INIT('h80)
	) name24239 (
		\m4_data_i[2]_pad ,
		_w8782_,
		_w8783_,
		_w26140_
	);
	LUT4 #(
		.INIT('h5d7f)
	) name24240 (
		_w8777_,
		_w8780_,
		_w26139_,
		_w26140_,
		_w26141_
	);
	LUT3 #(
		.INIT('h2a)
	) name24241 (
		\m7_data_i[2]_pad ,
		_w8782_,
		_w8783_,
		_w26142_
	);
	LUT3 #(
		.INIT('h2a)
	) name24242 (
		\m3_data_i[2]_pad ,
		_w8782_,
		_w8783_,
		_w26143_
	);
	LUT4 #(
		.INIT('habef)
	) name24243 (
		_w8777_,
		_w8780_,
		_w26142_,
		_w26143_,
		_w26144_
	);
	LUT3 #(
		.INIT('h80)
	) name24244 (
		\m6_data_i[2]_pad ,
		_w8782_,
		_w8783_,
		_w26145_
	);
	LUT3 #(
		.INIT('h2a)
	) name24245 (
		\m5_data_i[2]_pad ,
		_w8782_,
		_w8783_,
		_w26146_
	);
	LUT4 #(
		.INIT('hcdef)
	) name24246 (
		_w8777_,
		_w8780_,
		_w26145_,
		_w26146_,
		_w26147_
	);
	LUT4 #(
		.INIT('h7fff)
	) name24247 (
		_w26138_,
		_w26141_,
		_w26144_,
		_w26147_,
		_w26148_
	);
	LUT3 #(
		.INIT('h2a)
	) name24248 (
		\m3_data_i[30]_pad ,
		_w8782_,
		_w8783_,
		_w26149_
	);
	LUT3 #(
		.INIT('h80)
	) name24249 (
		\m4_data_i[30]_pad ,
		_w8782_,
		_w8783_,
		_w26150_
	);
	LUT4 #(
		.INIT('h9dbf)
	) name24250 (
		_w8777_,
		_w8780_,
		_w26149_,
		_w26150_,
		_w26151_
	);
	LUT3 #(
		.INIT('h80)
	) name24251 (
		\m6_data_i[30]_pad ,
		_w8782_,
		_w8783_,
		_w26152_
	);
	LUT3 #(
		.INIT('h2a)
	) name24252 (
		\m7_data_i[30]_pad ,
		_w8782_,
		_w8783_,
		_w26153_
	);
	LUT3 #(
		.INIT('h57)
	) name24253 (
		_w8781_,
		_w26152_,
		_w26153_,
		_w26154_
	);
	LUT3 #(
		.INIT('h2a)
	) name24254 (
		\m5_data_i[30]_pad ,
		_w8782_,
		_w8783_,
		_w26155_
	);
	LUT3 #(
		.INIT('h80)
	) name24255 (
		\m0_data_i[30]_pad ,
		_w8782_,
		_w8783_,
		_w26156_
	);
	LUT4 #(
		.INIT('h57df)
	) name24256 (
		_w8777_,
		_w8780_,
		_w26155_,
		_w26156_,
		_w26157_
	);
	LUT3 #(
		.INIT('h2a)
	) name24257 (
		\m1_data_i[30]_pad ,
		_w8782_,
		_w8783_,
		_w26158_
	);
	LUT3 #(
		.INIT('h80)
	) name24258 (
		\m2_data_i[30]_pad ,
		_w8782_,
		_w8783_,
		_w26159_
	);
	LUT4 #(
		.INIT('h3b7f)
	) name24259 (
		_w8777_,
		_w8780_,
		_w26158_,
		_w26159_,
		_w26160_
	);
	LUT4 #(
		.INIT('h7fff)
	) name24260 (
		_w26151_,
		_w26154_,
		_w26157_,
		_w26160_,
		_w26161_
	);
	LUT3 #(
		.INIT('h2a)
	) name24261 (
		\m3_data_i[31]_pad ,
		_w8782_,
		_w8783_,
		_w26162_
	);
	LUT3 #(
		.INIT('h80)
	) name24262 (
		\m4_data_i[31]_pad ,
		_w8782_,
		_w8783_,
		_w26163_
	);
	LUT4 #(
		.INIT('h9dbf)
	) name24263 (
		_w8777_,
		_w8780_,
		_w26162_,
		_w26163_,
		_w26164_
	);
	LUT3 #(
		.INIT('h80)
	) name24264 (
		\m6_data_i[31]_pad ,
		_w8782_,
		_w8783_,
		_w26165_
	);
	LUT3 #(
		.INIT('h80)
	) name24265 (
		\m2_data_i[31]_pad ,
		_w8782_,
		_w8783_,
		_w26166_
	);
	LUT4 #(
		.INIT('habef)
	) name24266 (
		_w8777_,
		_w8780_,
		_w26165_,
		_w26166_,
		_w26167_
	);
	LUT3 #(
		.INIT('h2a)
	) name24267 (
		\m5_data_i[31]_pad ,
		_w8782_,
		_w8783_,
		_w26168_
	);
	LUT3 #(
		.INIT('h2a)
	) name24268 (
		\m1_data_i[31]_pad ,
		_w8782_,
		_w8783_,
		_w26169_
	);
	LUT4 #(
		.INIT('h57df)
	) name24269 (
		_w8777_,
		_w8780_,
		_w26168_,
		_w26169_,
		_w26170_
	);
	LUT3 #(
		.INIT('h80)
	) name24270 (
		\m0_data_i[31]_pad ,
		_w8782_,
		_w8783_,
		_w26171_
	);
	LUT3 #(
		.INIT('h2a)
	) name24271 (
		\m7_data_i[31]_pad ,
		_w8782_,
		_w8783_,
		_w26172_
	);
	LUT4 #(
		.INIT('h6e7f)
	) name24272 (
		_w8777_,
		_w8780_,
		_w26171_,
		_w26172_,
		_w26173_
	);
	LUT4 #(
		.INIT('h7fff)
	) name24273 (
		_w26164_,
		_w26167_,
		_w26170_,
		_w26173_,
		_w26174_
	);
	LUT3 #(
		.INIT('h2a)
	) name24274 (
		\m3_data_i[3]_pad ,
		_w8782_,
		_w8783_,
		_w26175_
	);
	LUT3 #(
		.INIT('h80)
	) name24275 (
		\m4_data_i[3]_pad ,
		_w8782_,
		_w8783_,
		_w26176_
	);
	LUT4 #(
		.INIT('h9dbf)
	) name24276 (
		_w8777_,
		_w8780_,
		_w26175_,
		_w26176_,
		_w26177_
	);
	LUT3 #(
		.INIT('h80)
	) name24277 (
		\m6_data_i[3]_pad ,
		_w8782_,
		_w8783_,
		_w26178_
	);
	LUT3 #(
		.INIT('h80)
	) name24278 (
		\m2_data_i[3]_pad ,
		_w8782_,
		_w8783_,
		_w26179_
	);
	LUT4 #(
		.INIT('habef)
	) name24279 (
		_w8777_,
		_w8780_,
		_w26178_,
		_w26179_,
		_w26180_
	);
	LUT3 #(
		.INIT('h2a)
	) name24280 (
		\m5_data_i[3]_pad ,
		_w8782_,
		_w8783_,
		_w26181_
	);
	LUT3 #(
		.INIT('h2a)
	) name24281 (
		\m1_data_i[3]_pad ,
		_w8782_,
		_w8783_,
		_w26182_
	);
	LUT4 #(
		.INIT('h57df)
	) name24282 (
		_w8777_,
		_w8780_,
		_w26181_,
		_w26182_,
		_w26183_
	);
	LUT3 #(
		.INIT('h80)
	) name24283 (
		\m0_data_i[3]_pad ,
		_w8782_,
		_w8783_,
		_w26184_
	);
	LUT3 #(
		.INIT('h2a)
	) name24284 (
		\m7_data_i[3]_pad ,
		_w8782_,
		_w8783_,
		_w26185_
	);
	LUT4 #(
		.INIT('h6e7f)
	) name24285 (
		_w8777_,
		_w8780_,
		_w26184_,
		_w26185_,
		_w26186_
	);
	LUT4 #(
		.INIT('h7fff)
	) name24286 (
		_w26177_,
		_w26180_,
		_w26183_,
		_w26186_,
		_w26187_
	);
	LUT3 #(
		.INIT('h2a)
	) name24287 (
		\m1_data_i[4]_pad ,
		_w8782_,
		_w8783_,
		_w26188_
	);
	LUT3 #(
		.INIT('h80)
	) name24288 (
		\m2_data_i[4]_pad ,
		_w8782_,
		_w8783_,
		_w26189_
	);
	LUT4 #(
		.INIT('h3b7f)
	) name24289 (
		_w8777_,
		_w8780_,
		_w26188_,
		_w26189_,
		_w26190_
	);
	LUT3 #(
		.INIT('h80)
	) name24290 (
		\m6_data_i[4]_pad ,
		_w8782_,
		_w8783_,
		_w26191_
	);
	LUT3 #(
		.INIT('h2a)
	) name24291 (
		\m7_data_i[4]_pad ,
		_w8782_,
		_w8783_,
		_w26192_
	);
	LUT3 #(
		.INIT('h57)
	) name24292 (
		_w8781_,
		_w26191_,
		_w26192_,
		_w26193_
	);
	LUT3 #(
		.INIT('h2a)
	) name24293 (
		\m5_data_i[4]_pad ,
		_w8782_,
		_w8783_,
		_w26194_
	);
	LUT3 #(
		.INIT('h80)
	) name24294 (
		\m0_data_i[4]_pad ,
		_w8782_,
		_w8783_,
		_w26195_
	);
	LUT4 #(
		.INIT('h57df)
	) name24295 (
		_w8777_,
		_w8780_,
		_w26194_,
		_w26195_,
		_w26196_
	);
	LUT3 #(
		.INIT('h2a)
	) name24296 (
		\m3_data_i[4]_pad ,
		_w8782_,
		_w8783_,
		_w26197_
	);
	LUT3 #(
		.INIT('h80)
	) name24297 (
		\m4_data_i[4]_pad ,
		_w8782_,
		_w8783_,
		_w26198_
	);
	LUT4 #(
		.INIT('h9dbf)
	) name24298 (
		_w8777_,
		_w8780_,
		_w26197_,
		_w26198_,
		_w26199_
	);
	LUT4 #(
		.INIT('h7fff)
	) name24299 (
		_w26190_,
		_w26193_,
		_w26196_,
		_w26199_,
		_w26200_
	);
	LUT3 #(
		.INIT('h2a)
	) name24300 (
		\m1_data_i[5]_pad ,
		_w8782_,
		_w8783_,
		_w26201_
	);
	LUT3 #(
		.INIT('h80)
	) name24301 (
		\m2_data_i[5]_pad ,
		_w8782_,
		_w8783_,
		_w26202_
	);
	LUT4 #(
		.INIT('h3b7f)
	) name24302 (
		_w8777_,
		_w8780_,
		_w26201_,
		_w26202_,
		_w26203_
	);
	LUT3 #(
		.INIT('h80)
	) name24303 (
		\m0_data_i[5]_pad ,
		_w8782_,
		_w8783_,
		_w26204_
	);
	LUT3 #(
		.INIT('h80)
	) name24304 (
		\m4_data_i[5]_pad ,
		_w8782_,
		_w8783_,
		_w26205_
	);
	LUT4 #(
		.INIT('h5d7f)
	) name24305 (
		_w8777_,
		_w8780_,
		_w26204_,
		_w26205_,
		_w26206_
	);
	LUT3 #(
		.INIT('h2a)
	) name24306 (
		\m7_data_i[5]_pad ,
		_w8782_,
		_w8783_,
		_w26207_
	);
	LUT3 #(
		.INIT('h2a)
	) name24307 (
		\m3_data_i[5]_pad ,
		_w8782_,
		_w8783_,
		_w26208_
	);
	LUT4 #(
		.INIT('habef)
	) name24308 (
		_w8777_,
		_w8780_,
		_w26207_,
		_w26208_,
		_w26209_
	);
	LUT3 #(
		.INIT('h80)
	) name24309 (
		\m6_data_i[5]_pad ,
		_w8782_,
		_w8783_,
		_w26210_
	);
	LUT3 #(
		.INIT('h2a)
	) name24310 (
		\m5_data_i[5]_pad ,
		_w8782_,
		_w8783_,
		_w26211_
	);
	LUT4 #(
		.INIT('hcdef)
	) name24311 (
		_w8777_,
		_w8780_,
		_w26210_,
		_w26211_,
		_w26212_
	);
	LUT4 #(
		.INIT('h7fff)
	) name24312 (
		_w26203_,
		_w26206_,
		_w26209_,
		_w26212_,
		_w26213_
	);
	LUT3 #(
		.INIT('h80)
	) name24313 (
		\m6_data_i[6]_pad ,
		_w8782_,
		_w8783_,
		_w26214_
	);
	LUT3 #(
		.INIT('h2a)
	) name24314 (
		\m5_data_i[6]_pad ,
		_w8782_,
		_w8783_,
		_w26215_
	);
	LUT4 #(
		.INIT('hcdef)
	) name24315 (
		_w8777_,
		_w8780_,
		_w26214_,
		_w26215_,
		_w26216_
	);
	LUT3 #(
		.INIT('h2a)
	) name24316 (
		\m3_data_i[6]_pad ,
		_w8782_,
		_w8783_,
		_w26217_
	);
	LUT3 #(
		.INIT('h2a)
	) name24317 (
		\m7_data_i[6]_pad ,
		_w8782_,
		_w8783_,
		_w26218_
	);
	LUT4 #(
		.INIT('haebf)
	) name24318 (
		_w8777_,
		_w8780_,
		_w26217_,
		_w26218_,
		_w26219_
	);
	LUT3 #(
		.INIT('h80)
	) name24319 (
		\m4_data_i[6]_pad ,
		_w8782_,
		_w8783_,
		_w26220_
	);
	LUT3 #(
		.INIT('h80)
	) name24320 (
		\m0_data_i[6]_pad ,
		_w8782_,
		_w8783_,
		_w26221_
	);
	LUT4 #(
		.INIT('h57df)
	) name24321 (
		_w8777_,
		_w8780_,
		_w26220_,
		_w26221_,
		_w26222_
	);
	LUT3 #(
		.INIT('h2a)
	) name24322 (
		\m1_data_i[6]_pad ,
		_w8782_,
		_w8783_,
		_w26223_
	);
	LUT3 #(
		.INIT('h80)
	) name24323 (
		\m2_data_i[6]_pad ,
		_w8782_,
		_w8783_,
		_w26224_
	);
	LUT4 #(
		.INIT('h3b7f)
	) name24324 (
		_w8777_,
		_w8780_,
		_w26223_,
		_w26224_,
		_w26225_
	);
	LUT4 #(
		.INIT('h7fff)
	) name24325 (
		_w26216_,
		_w26219_,
		_w26222_,
		_w26225_,
		_w26226_
	);
	LUT3 #(
		.INIT('h2a)
	) name24326 (
		\m1_data_i[7]_pad ,
		_w8782_,
		_w8783_,
		_w26227_
	);
	LUT3 #(
		.INIT('h80)
	) name24327 (
		\m2_data_i[7]_pad ,
		_w8782_,
		_w8783_,
		_w26228_
	);
	LUT4 #(
		.INIT('h3b7f)
	) name24328 (
		_w8777_,
		_w8780_,
		_w26227_,
		_w26228_,
		_w26229_
	);
	LUT3 #(
		.INIT('h80)
	) name24329 (
		\m6_data_i[7]_pad ,
		_w8782_,
		_w8783_,
		_w26230_
	);
	LUT3 #(
		.INIT('h2a)
	) name24330 (
		\m7_data_i[7]_pad ,
		_w8782_,
		_w8783_,
		_w26231_
	);
	LUT3 #(
		.INIT('h57)
	) name24331 (
		_w8781_,
		_w26230_,
		_w26231_,
		_w26232_
	);
	LUT3 #(
		.INIT('h2a)
	) name24332 (
		\m5_data_i[7]_pad ,
		_w8782_,
		_w8783_,
		_w26233_
	);
	LUT3 #(
		.INIT('h80)
	) name24333 (
		\m0_data_i[7]_pad ,
		_w8782_,
		_w8783_,
		_w26234_
	);
	LUT4 #(
		.INIT('h57df)
	) name24334 (
		_w8777_,
		_w8780_,
		_w26233_,
		_w26234_,
		_w26235_
	);
	LUT3 #(
		.INIT('h2a)
	) name24335 (
		\m3_data_i[7]_pad ,
		_w8782_,
		_w8783_,
		_w26236_
	);
	LUT3 #(
		.INIT('h80)
	) name24336 (
		\m4_data_i[7]_pad ,
		_w8782_,
		_w8783_,
		_w26237_
	);
	LUT4 #(
		.INIT('h9dbf)
	) name24337 (
		_w8777_,
		_w8780_,
		_w26236_,
		_w26237_,
		_w26238_
	);
	LUT4 #(
		.INIT('h7fff)
	) name24338 (
		_w26229_,
		_w26232_,
		_w26235_,
		_w26238_,
		_w26239_
	);
	LUT3 #(
		.INIT('h2a)
	) name24339 (
		\m1_data_i[8]_pad ,
		_w8782_,
		_w8783_,
		_w26240_
	);
	LUT3 #(
		.INIT('h80)
	) name24340 (
		\m2_data_i[8]_pad ,
		_w8782_,
		_w8783_,
		_w26241_
	);
	LUT4 #(
		.INIT('h3b7f)
	) name24341 (
		_w8777_,
		_w8780_,
		_w26240_,
		_w26241_,
		_w26242_
	);
	LUT3 #(
		.INIT('h2a)
	) name24342 (
		\m3_data_i[8]_pad ,
		_w8782_,
		_w8783_,
		_w26243_
	);
	LUT3 #(
		.INIT('h2a)
	) name24343 (
		\m7_data_i[8]_pad ,
		_w8782_,
		_w8783_,
		_w26244_
	);
	LUT4 #(
		.INIT('haebf)
	) name24344 (
		_w8777_,
		_w8780_,
		_w26243_,
		_w26244_,
		_w26245_
	);
	LUT3 #(
		.INIT('h80)
	) name24345 (
		\m4_data_i[8]_pad ,
		_w8782_,
		_w8783_,
		_w26246_
	);
	LUT3 #(
		.INIT('h80)
	) name24346 (
		\m0_data_i[8]_pad ,
		_w8782_,
		_w8783_,
		_w26247_
	);
	LUT4 #(
		.INIT('h57df)
	) name24347 (
		_w8777_,
		_w8780_,
		_w26246_,
		_w26247_,
		_w26248_
	);
	LUT3 #(
		.INIT('h80)
	) name24348 (
		\m6_data_i[8]_pad ,
		_w8782_,
		_w8783_,
		_w26249_
	);
	LUT3 #(
		.INIT('h2a)
	) name24349 (
		\m5_data_i[8]_pad ,
		_w8782_,
		_w8783_,
		_w26250_
	);
	LUT4 #(
		.INIT('hcdef)
	) name24350 (
		_w8777_,
		_w8780_,
		_w26249_,
		_w26250_,
		_w26251_
	);
	LUT4 #(
		.INIT('h7fff)
	) name24351 (
		_w26242_,
		_w26245_,
		_w26248_,
		_w26251_,
		_w26252_
	);
	LUT3 #(
		.INIT('h80)
	) name24352 (
		\m0_data_i[9]_pad ,
		_w8782_,
		_w8783_,
		_w26253_
	);
	LUT3 #(
		.INIT('h2a)
	) name24353 (
		\m7_data_i[9]_pad ,
		_w8782_,
		_w8783_,
		_w26254_
	);
	LUT4 #(
		.INIT('h6e7f)
	) name24354 (
		_w8777_,
		_w8780_,
		_w26253_,
		_w26254_,
		_w26255_
	);
	LUT3 #(
		.INIT('h2a)
	) name24355 (
		\m3_data_i[9]_pad ,
		_w8782_,
		_w8783_,
		_w26256_
	);
	LUT3 #(
		.INIT('h80)
	) name24356 (
		\m2_data_i[9]_pad ,
		_w8782_,
		_w8783_,
		_w26257_
	);
	LUT3 #(
		.INIT('h57)
	) name24357 (
		_w8795_,
		_w26256_,
		_w26257_,
		_w26258_
	);
	LUT3 #(
		.INIT('h80)
	) name24358 (
		\m4_data_i[9]_pad ,
		_w8782_,
		_w8783_,
		_w26259_
	);
	LUT3 #(
		.INIT('h2a)
	) name24359 (
		\m1_data_i[9]_pad ,
		_w8782_,
		_w8783_,
		_w26260_
	);
	LUT4 #(
		.INIT('h57df)
	) name24360 (
		_w8777_,
		_w8780_,
		_w26259_,
		_w26260_,
		_w26261_
	);
	LUT3 #(
		.INIT('h80)
	) name24361 (
		\m6_data_i[9]_pad ,
		_w8782_,
		_w8783_,
		_w26262_
	);
	LUT3 #(
		.INIT('h2a)
	) name24362 (
		\m5_data_i[9]_pad ,
		_w8782_,
		_w8783_,
		_w26263_
	);
	LUT4 #(
		.INIT('hcdef)
	) name24363 (
		_w8777_,
		_w8780_,
		_w26262_,
		_w26263_,
		_w26264_
	);
	LUT4 #(
		.INIT('h7fff)
	) name24364 (
		_w26255_,
		_w26258_,
		_w26261_,
		_w26264_,
		_w26265_
	);
	LUT3 #(
		.INIT('h2a)
	) name24365 (
		\m3_sel_i[0]_pad ,
		_w8782_,
		_w8783_,
		_w26266_
	);
	LUT3 #(
		.INIT('h80)
	) name24366 (
		\m4_sel_i[0]_pad ,
		_w8782_,
		_w8783_,
		_w26267_
	);
	LUT4 #(
		.INIT('h9dbf)
	) name24367 (
		_w8777_,
		_w8780_,
		_w26266_,
		_w26267_,
		_w26268_
	);
	LUT3 #(
		.INIT('h80)
	) name24368 (
		\m6_sel_i[0]_pad ,
		_w8782_,
		_w8783_,
		_w26269_
	);
	LUT3 #(
		.INIT('h80)
	) name24369 (
		\m2_sel_i[0]_pad ,
		_w8782_,
		_w8783_,
		_w26270_
	);
	LUT4 #(
		.INIT('habef)
	) name24370 (
		_w8777_,
		_w8780_,
		_w26269_,
		_w26270_,
		_w26271_
	);
	LUT3 #(
		.INIT('h2a)
	) name24371 (
		\m5_sel_i[0]_pad ,
		_w8782_,
		_w8783_,
		_w26272_
	);
	LUT3 #(
		.INIT('h2a)
	) name24372 (
		\m1_sel_i[0]_pad ,
		_w8782_,
		_w8783_,
		_w26273_
	);
	LUT4 #(
		.INIT('h57df)
	) name24373 (
		_w8777_,
		_w8780_,
		_w26272_,
		_w26273_,
		_w26274_
	);
	LUT3 #(
		.INIT('h80)
	) name24374 (
		\m0_sel_i[0]_pad ,
		_w8782_,
		_w8783_,
		_w26275_
	);
	LUT3 #(
		.INIT('h2a)
	) name24375 (
		\m7_sel_i[0]_pad ,
		_w8782_,
		_w8783_,
		_w26276_
	);
	LUT4 #(
		.INIT('h6e7f)
	) name24376 (
		_w8777_,
		_w8780_,
		_w26275_,
		_w26276_,
		_w26277_
	);
	LUT4 #(
		.INIT('h7fff)
	) name24377 (
		_w26268_,
		_w26271_,
		_w26274_,
		_w26277_,
		_w26278_
	);
	LUT3 #(
		.INIT('h2a)
	) name24378 (
		\m1_sel_i[1]_pad ,
		_w8782_,
		_w8783_,
		_w26279_
	);
	LUT3 #(
		.INIT('h80)
	) name24379 (
		\m2_sel_i[1]_pad ,
		_w8782_,
		_w8783_,
		_w26280_
	);
	LUT4 #(
		.INIT('h3b7f)
	) name24380 (
		_w8777_,
		_w8780_,
		_w26279_,
		_w26280_,
		_w26281_
	);
	LUT3 #(
		.INIT('h80)
	) name24381 (
		\m6_sel_i[1]_pad ,
		_w8782_,
		_w8783_,
		_w26282_
	);
	LUT3 #(
		.INIT('h2a)
	) name24382 (
		\m7_sel_i[1]_pad ,
		_w8782_,
		_w8783_,
		_w26283_
	);
	LUT3 #(
		.INIT('h57)
	) name24383 (
		_w8781_,
		_w26282_,
		_w26283_,
		_w26284_
	);
	LUT3 #(
		.INIT('h2a)
	) name24384 (
		\m5_sel_i[1]_pad ,
		_w8782_,
		_w8783_,
		_w26285_
	);
	LUT3 #(
		.INIT('h80)
	) name24385 (
		\m0_sel_i[1]_pad ,
		_w8782_,
		_w8783_,
		_w26286_
	);
	LUT4 #(
		.INIT('h57df)
	) name24386 (
		_w8777_,
		_w8780_,
		_w26285_,
		_w26286_,
		_w26287_
	);
	LUT3 #(
		.INIT('h2a)
	) name24387 (
		\m3_sel_i[1]_pad ,
		_w8782_,
		_w8783_,
		_w26288_
	);
	LUT3 #(
		.INIT('h80)
	) name24388 (
		\m4_sel_i[1]_pad ,
		_w8782_,
		_w8783_,
		_w26289_
	);
	LUT4 #(
		.INIT('h9dbf)
	) name24389 (
		_w8777_,
		_w8780_,
		_w26288_,
		_w26289_,
		_w26290_
	);
	LUT4 #(
		.INIT('h7fff)
	) name24390 (
		_w26281_,
		_w26284_,
		_w26287_,
		_w26290_,
		_w26291_
	);
	LUT3 #(
		.INIT('h2a)
	) name24391 (
		\m3_sel_i[2]_pad ,
		_w8782_,
		_w8783_,
		_w26292_
	);
	LUT3 #(
		.INIT('h80)
	) name24392 (
		\m4_sel_i[2]_pad ,
		_w8782_,
		_w8783_,
		_w26293_
	);
	LUT4 #(
		.INIT('h9dbf)
	) name24393 (
		_w8777_,
		_w8780_,
		_w26292_,
		_w26293_,
		_w26294_
	);
	LUT3 #(
		.INIT('h80)
	) name24394 (
		\m6_sel_i[2]_pad ,
		_w8782_,
		_w8783_,
		_w26295_
	);
	LUT3 #(
		.INIT('h80)
	) name24395 (
		\m2_sel_i[2]_pad ,
		_w8782_,
		_w8783_,
		_w26296_
	);
	LUT4 #(
		.INIT('habef)
	) name24396 (
		_w8777_,
		_w8780_,
		_w26295_,
		_w26296_,
		_w26297_
	);
	LUT3 #(
		.INIT('h2a)
	) name24397 (
		\m5_sel_i[2]_pad ,
		_w8782_,
		_w8783_,
		_w26298_
	);
	LUT3 #(
		.INIT('h2a)
	) name24398 (
		\m1_sel_i[2]_pad ,
		_w8782_,
		_w8783_,
		_w26299_
	);
	LUT4 #(
		.INIT('h57df)
	) name24399 (
		_w8777_,
		_w8780_,
		_w26298_,
		_w26299_,
		_w26300_
	);
	LUT3 #(
		.INIT('h80)
	) name24400 (
		\m0_sel_i[2]_pad ,
		_w8782_,
		_w8783_,
		_w26301_
	);
	LUT3 #(
		.INIT('h2a)
	) name24401 (
		\m7_sel_i[2]_pad ,
		_w8782_,
		_w8783_,
		_w26302_
	);
	LUT4 #(
		.INIT('h6e7f)
	) name24402 (
		_w8777_,
		_w8780_,
		_w26301_,
		_w26302_,
		_w26303_
	);
	LUT4 #(
		.INIT('h7fff)
	) name24403 (
		_w26294_,
		_w26297_,
		_w26300_,
		_w26303_,
		_w26304_
	);
	LUT3 #(
		.INIT('h2a)
	) name24404 (
		\m3_sel_i[3]_pad ,
		_w8782_,
		_w8783_,
		_w26305_
	);
	LUT3 #(
		.INIT('h80)
	) name24405 (
		\m4_sel_i[3]_pad ,
		_w8782_,
		_w8783_,
		_w26306_
	);
	LUT4 #(
		.INIT('h9dbf)
	) name24406 (
		_w8777_,
		_w8780_,
		_w26305_,
		_w26306_,
		_w26307_
	);
	LUT3 #(
		.INIT('h80)
	) name24407 (
		\m6_sel_i[3]_pad ,
		_w8782_,
		_w8783_,
		_w26308_
	);
	LUT3 #(
		.INIT('h80)
	) name24408 (
		\m2_sel_i[3]_pad ,
		_w8782_,
		_w8783_,
		_w26309_
	);
	LUT4 #(
		.INIT('habef)
	) name24409 (
		_w8777_,
		_w8780_,
		_w26308_,
		_w26309_,
		_w26310_
	);
	LUT3 #(
		.INIT('h2a)
	) name24410 (
		\m5_sel_i[3]_pad ,
		_w8782_,
		_w8783_,
		_w26311_
	);
	LUT3 #(
		.INIT('h2a)
	) name24411 (
		\m1_sel_i[3]_pad ,
		_w8782_,
		_w8783_,
		_w26312_
	);
	LUT4 #(
		.INIT('h57df)
	) name24412 (
		_w8777_,
		_w8780_,
		_w26311_,
		_w26312_,
		_w26313_
	);
	LUT3 #(
		.INIT('h80)
	) name24413 (
		\m0_sel_i[3]_pad ,
		_w8782_,
		_w8783_,
		_w26314_
	);
	LUT3 #(
		.INIT('h2a)
	) name24414 (
		\m7_sel_i[3]_pad ,
		_w8782_,
		_w8783_,
		_w26315_
	);
	LUT4 #(
		.INIT('h6e7f)
	) name24415 (
		_w8777_,
		_w8780_,
		_w26314_,
		_w26315_,
		_w26316_
	);
	LUT4 #(
		.INIT('h7fff)
	) name24416 (
		_w26307_,
		_w26310_,
		_w26313_,
		_w26316_,
		_w26317_
	);
	LUT4 #(
		.INIT('h2a00)
	) name24417 (
		\m5_stb_i_pad ,
		_w8782_,
		_w8783_,
		_w9345_,
		_w26318_
	);
	LUT4 #(
		.INIT('h8000)
	) name24418 (
		\m4_stb_i_pad ,
		_w8782_,
		_w8783_,
		_w9529_,
		_w26319_
	);
	LUT3 #(
		.INIT('h57)
	) name24419 (
		_w8801_,
		_w26318_,
		_w26319_,
		_w26320_
	);
	LUT4 #(
		.INIT('h8000)
	) name24420 (
		\m6_stb_i_pad ,
		_w8782_,
		_w8783_,
		_w9588_,
		_w26321_
	);
	LUT4 #(
		.INIT('h2a00)
	) name24421 (
		\m1_stb_i_pad ,
		_w8782_,
		_w8783_,
		_w9442_,
		_w26322_
	);
	LUT4 #(
		.INIT('h67ef)
	) name24422 (
		_w8777_,
		_w8780_,
		_w26321_,
		_w26322_,
		_w26323_
	);
	LUT4 #(
		.INIT('h2a00)
	) name24423 (
		\m7_stb_i_pad ,
		_w8782_,
		_w8783_,
		_w9330_,
		_w26324_
	);
	LUT4 #(
		.INIT('h2a00)
	) name24424 (
		\m3_stb_i_pad ,
		_w8782_,
		_w8783_,
		_w9375_,
		_w26325_
	);
	LUT4 #(
		.INIT('habef)
	) name24425 (
		_w8777_,
		_w8780_,
		_w26324_,
		_w26325_,
		_w26326_
	);
	LUT4 #(
		.INIT('h8000)
	) name24426 (
		\m2_stb_i_pad ,
		_w8782_,
		_w8783_,
		_w9626_,
		_w26327_
	);
	LUT4 #(
		.INIT('h8000)
	) name24427 (
		\m0_stb_i_pad ,
		_w8782_,
		_w8783_,
		_w9407_,
		_w26328_
	);
	LUT4 #(
		.INIT('h37bf)
	) name24428 (
		_w8777_,
		_w8780_,
		_w26327_,
		_w26328_,
		_w26329_
	);
	LUT4 #(
		.INIT('h7fff)
	) name24429 (
		_w26320_,
		_w26323_,
		_w26326_,
		_w26329_,
		_w26330_
	);
	LUT3 #(
		.INIT('h2a)
	) name24430 (
		\m1_we_i_pad ,
		_w8782_,
		_w8783_,
		_w26331_
	);
	LUT3 #(
		.INIT('h80)
	) name24431 (
		\m2_we_i_pad ,
		_w8782_,
		_w8783_,
		_w26332_
	);
	LUT4 #(
		.INIT('h3b7f)
	) name24432 (
		_w8777_,
		_w8780_,
		_w26331_,
		_w26332_,
		_w26333_
	);
	LUT3 #(
		.INIT('h80)
	) name24433 (
		\m6_we_i_pad ,
		_w8782_,
		_w8783_,
		_w26334_
	);
	LUT3 #(
		.INIT('h2a)
	) name24434 (
		\m7_we_i_pad ,
		_w8782_,
		_w8783_,
		_w26335_
	);
	LUT3 #(
		.INIT('h57)
	) name24435 (
		_w8781_,
		_w26334_,
		_w26335_,
		_w26336_
	);
	LUT3 #(
		.INIT('h2a)
	) name24436 (
		\m5_we_i_pad ,
		_w8782_,
		_w8783_,
		_w26337_
	);
	LUT3 #(
		.INIT('h80)
	) name24437 (
		\m0_we_i_pad ,
		_w8782_,
		_w8783_,
		_w26338_
	);
	LUT4 #(
		.INIT('h57df)
	) name24438 (
		_w8777_,
		_w8780_,
		_w26337_,
		_w26338_,
		_w26339_
	);
	LUT3 #(
		.INIT('h2a)
	) name24439 (
		\m3_we_i_pad ,
		_w8782_,
		_w8783_,
		_w26340_
	);
	LUT3 #(
		.INIT('h80)
	) name24440 (
		\m4_we_i_pad ,
		_w8782_,
		_w8783_,
		_w26341_
	);
	LUT4 #(
		.INIT('h9dbf)
	) name24441 (
		_w8777_,
		_w8780_,
		_w26340_,
		_w26341_,
		_w26342_
	);
	LUT4 #(
		.INIT('h7fff)
	) name24442 (
		_w26333_,
		_w26336_,
		_w26339_,
		_w26342_,
		_w26343_
	);
	LUT3 #(
		.INIT('h2a)
	) name24443 (
		\m1_addr_i[0]_pad ,
		_w8821_,
		_w8822_,
		_w26344_
	);
	LUT3 #(
		.INIT('h80)
	) name24444 (
		\m2_addr_i[0]_pad ,
		_w8821_,
		_w8822_,
		_w26345_
	);
	LUT4 #(
		.INIT('h3b7f)
	) name24445 (
		_w8816_,
		_w8819_,
		_w26344_,
		_w26345_,
		_w26346_
	);
	LUT3 #(
		.INIT('h80)
	) name24446 (
		\m6_addr_i[0]_pad ,
		_w8821_,
		_w8822_,
		_w26347_
	);
	LUT3 #(
		.INIT('h2a)
	) name24447 (
		\m7_addr_i[0]_pad ,
		_w8821_,
		_w8822_,
		_w26348_
	);
	LUT3 #(
		.INIT('h57)
	) name24448 (
		_w8834_,
		_w26347_,
		_w26348_,
		_w26349_
	);
	LUT3 #(
		.INIT('h2a)
	) name24449 (
		\m5_addr_i[0]_pad ,
		_w8821_,
		_w8822_,
		_w26350_
	);
	LUT3 #(
		.INIT('h80)
	) name24450 (
		\m0_addr_i[0]_pad ,
		_w8821_,
		_w8822_,
		_w26351_
	);
	LUT4 #(
		.INIT('h57df)
	) name24451 (
		_w8816_,
		_w8819_,
		_w26350_,
		_w26351_,
		_w26352_
	);
	LUT3 #(
		.INIT('h2a)
	) name24452 (
		\m3_addr_i[0]_pad ,
		_w8821_,
		_w8822_,
		_w26353_
	);
	LUT3 #(
		.INIT('h80)
	) name24453 (
		\m4_addr_i[0]_pad ,
		_w8821_,
		_w8822_,
		_w26354_
	);
	LUT4 #(
		.INIT('h9dbf)
	) name24454 (
		_w8816_,
		_w8819_,
		_w26353_,
		_w26354_,
		_w26355_
	);
	LUT4 #(
		.INIT('h7fff)
	) name24455 (
		_w26346_,
		_w26349_,
		_w26352_,
		_w26355_,
		_w26356_
	);
	LUT3 #(
		.INIT('h2a)
	) name24456 (
		\m3_addr_i[10]_pad ,
		_w8821_,
		_w8822_,
		_w26357_
	);
	LUT3 #(
		.INIT('h80)
	) name24457 (
		\m4_addr_i[10]_pad ,
		_w8821_,
		_w8822_,
		_w26358_
	);
	LUT4 #(
		.INIT('h9dbf)
	) name24458 (
		_w8816_,
		_w8819_,
		_w26357_,
		_w26358_,
		_w26359_
	);
	LUT3 #(
		.INIT('h80)
	) name24459 (
		\m6_addr_i[10]_pad ,
		_w8821_,
		_w8822_,
		_w26360_
	);
	LUT3 #(
		.INIT('h2a)
	) name24460 (
		\m7_addr_i[10]_pad ,
		_w8821_,
		_w8822_,
		_w26361_
	);
	LUT3 #(
		.INIT('h57)
	) name24461 (
		_w8834_,
		_w26360_,
		_w26361_,
		_w26362_
	);
	LUT3 #(
		.INIT('h2a)
	) name24462 (
		\m5_addr_i[10]_pad ,
		_w8821_,
		_w8822_,
		_w26363_
	);
	LUT3 #(
		.INIT('h80)
	) name24463 (
		\m0_addr_i[10]_pad ,
		_w8821_,
		_w8822_,
		_w26364_
	);
	LUT4 #(
		.INIT('h57df)
	) name24464 (
		_w8816_,
		_w8819_,
		_w26363_,
		_w26364_,
		_w26365_
	);
	LUT3 #(
		.INIT('h2a)
	) name24465 (
		\m1_addr_i[10]_pad ,
		_w8821_,
		_w8822_,
		_w26366_
	);
	LUT3 #(
		.INIT('h80)
	) name24466 (
		\m2_addr_i[10]_pad ,
		_w8821_,
		_w8822_,
		_w26367_
	);
	LUT4 #(
		.INIT('h3b7f)
	) name24467 (
		_w8816_,
		_w8819_,
		_w26366_,
		_w26367_,
		_w26368_
	);
	LUT4 #(
		.INIT('h7fff)
	) name24468 (
		_w26359_,
		_w26362_,
		_w26365_,
		_w26368_,
		_w26369_
	);
	LUT3 #(
		.INIT('h2a)
	) name24469 (
		\m3_addr_i[11]_pad ,
		_w8821_,
		_w8822_,
		_w26370_
	);
	LUT3 #(
		.INIT('h80)
	) name24470 (
		\m4_addr_i[11]_pad ,
		_w8821_,
		_w8822_,
		_w26371_
	);
	LUT4 #(
		.INIT('h9dbf)
	) name24471 (
		_w8816_,
		_w8819_,
		_w26370_,
		_w26371_,
		_w26372_
	);
	LUT3 #(
		.INIT('h80)
	) name24472 (
		\m6_addr_i[11]_pad ,
		_w8821_,
		_w8822_,
		_w26373_
	);
	LUT3 #(
		.INIT('h80)
	) name24473 (
		\m2_addr_i[11]_pad ,
		_w8821_,
		_w8822_,
		_w26374_
	);
	LUT4 #(
		.INIT('habef)
	) name24474 (
		_w8816_,
		_w8819_,
		_w26373_,
		_w26374_,
		_w26375_
	);
	LUT3 #(
		.INIT('h2a)
	) name24475 (
		\m5_addr_i[11]_pad ,
		_w8821_,
		_w8822_,
		_w26376_
	);
	LUT3 #(
		.INIT('h2a)
	) name24476 (
		\m1_addr_i[11]_pad ,
		_w8821_,
		_w8822_,
		_w26377_
	);
	LUT4 #(
		.INIT('h57df)
	) name24477 (
		_w8816_,
		_w8819_,
		_w26376_,
		_w26377_,
		_w26378_
	);
	LUT3 #(
		.INIT('h80)
	) name24478 (
		\m0_addr_i[11]_pad ,
		_w8821_,
		_w8822_,
		_w26379_
	);
	LUT3 #(
		.INIT('h2a)
	) name24479 (
		\m7_addr_i[11]_pad ,
		_w8821_,
		_w8822_,
		_w26380_
	);
	LUT4 #(
		.INIT('h6e7f)
	) name24480 (
		_w8816_,
		_w8819_,
		_w26379_,
		_w26380_,
		_w26381_
	);
	LUT4 #(
		.INIT('h7fff)
	) name24481 (
		_w26372_,
		_w26375_,
		_w26378_,
		_w26381_,
		_w26382_
	);
	LUT3 #(
		.INIT('h2a)
	) name24482 (
		\m1_addr_i[12]_pad ,
		_w8821_,
		_w8822_,
		_w26383_
	);
	LUT3 #(
		.INIT('h80)
	) name24483 (
		\m2_addr_i[12]_pad ,
		_w8821_,
		_w8822_,
		_w26384_
	);
	LUT4 #(
		.INIT('h3b7f)
	) name24484 (
		_w8816_,
		_w8819_,
		_w26383_,
		_w26384_,
		_w26385_
	);
	LUT3 #(
		.INIT('h2a)
	) name24485 (
		\m3_addr_i[12]_pad ,
		_w8821_,
		_w8822_,
		_w26386_
	);
	LUT3 #(
		.INIT('h2a)
	) name24486 (
		\m7_addr_i[12]_pad ,
		_w8821_,
		_w8822_,
		_w26387_
	);
	LUT4 #(
		.INIT('haebf)
	) name24487 (
		_w8816_,
		_w8819_,
		_w26386_,
		_w26387_,
		_w26388_
	);
	LUT3 #(
		.INIT('h80)
	) name24488 (
		\m4_addr_i[12]_pad ,
		_w8821_,
		_w8822_,
		_w26389_
	);
	LUT3 #(
		.INIT('h80)
	) name24489 (
		\m0_addr_i[12]_pad ,
		_w8821_,
		_w8822_,
		_w26390_
	);
	LUT4 #(
		.INIT('h57df)
	) name24490 (
		_w8816_,
		_w8819_,
		_w26389_,
		_w26390_,
		_w26391_
	);
	LUT3 #(
		.INIT('h80)
	) name24491 (
		\m6_addr_i[12]_pad ,
		_w8821_,
		_w8822_,
		_w26392_
	);
	LUT3 #(
		.INIT('h2a)
	) name24492 (
		\m5_addr_i[12]_pad ,
		_w8821_,
		_w8822_,
		_w26393_
	);
	LUT4 #(
		.INIT('hcdef)
	) name24493 (
		_w8816_,
		_w8819_,
		_w26392_,
		_w26393_,
		_w26394_
	);
	LUT4 #(
		.INIT('h7fff)
	) name24494 (
		_w26385_,
		_w26388_,
		_w26391_,
		_w26394_,
		_w26395_
	);
	LUT3 #(
		.INIT('h2a)
	) name24495 (
		\m3_addr_i[13]_pad ,
		_w8821_,
		_w8822_,
		_w26396_
	);
	LUT3 #(
		.INIT('h80)
	) name24496 (
		\m4_addr_i[13]_pad ,
		_w8821_,
		_w8822_,
		_w26397_
	);
	LUT4 #(
		.INIT('h9dbf)
	) name24497 (
		_w8816_,
		_w8819_,
		_w26396_,
		_w26397_,
		_w26398_
	);
	LUT3 #(
		.INIT('h80)
	) name24498 (
		\m6_addr_i[13]_pad ,
		_w8821_,
		_w8822_,
		_w26399_
	);
	LUT3 #(
		.INIT('h80)
	) name24499 (
		\m2_addr_i[13]_pad ,
		_w8821_,
		_w8822_,
		_w26400_
	);
	LUT4 #(
		.INIT('habef)
	) name24500 (
		_w8816_,
		_w8819_,
		_w26399_,
		_w26400_,
		_w26401_
	);
	LUT3 #(
		.INIT('h2a)
	) name24501 (
		\m5_addr_i[13]_pad ,
		_w8821_,
		_w8822_,
		_w26402_
	);
	LUT3 #(
		.INIT('h2a)
	) name24502 (
		\m1_addr_i[13]_pad ,
		_w8821_,
		_w8822_,
		_w26403_
	);
	LUT4 #(
		.INIT('h57df)
	) name24503 (
		_w8816_,
		_w8819_,
		_w26402_,
		_w26403_,
		_w26404_
	);
	LUT3 #(
		.INIT('h80)
	) name24504 (
		\m0_addr_i[13]_pad ,
		_w8821_,
		_w8822_,
		_w26405_
	);
	LUT3 #(
		.INIT('h2a)
	) name24505 (
		\m7_addr_i[13]_pad ,
		_w8821_,
		_w8822_,
		_w26406_
	);
	LUT4 #(
		.INIT('h6e7f)
	) name24506 (
		_w8816_,
		_w8819_,
		_w26405_,
		_w26406_,
		_w26407_
	);
	LUT4 #(
		.INIT('h7fff)
	) name24507 (
		_w26398_,
		_w26401_,
		_w26404_,
		_w26407_,
		_w26408_
	);
	LUT3 #(
		.INIT('h2a)
	) name24508 (
		\m3_addr_i[14]_pad ,
		_w8821_,
		_w8822_,
		_w26409_
	);
	LUT3 #(
		.INIT('h80)
	) name24509 (
		\m4_addr_i[14]_pad ,
		_w8821_,
		_w8822_,
		_w26410_
	);
	LUT4 #(
		.INIT('h9dbf)
	) name24510 (
		_w8816_,
		_w8819_,
		_w26409_,
		_w26410_,
		_w26411_
	);
	LUT3 #(
		.INIT('h80)
	) name24511 (
		\m6_addr_i[14]_pad ,
		_w8821_,
		_w8822_,
		_w26412_
	);
	LUT3 #(
		.INIT('h80)
	) name24512 (
		\m2_addr_i[14]_pad ,
		_w8821_,
		_w8822_,
		_w26413_
	);
	LUT4 #(
		.INIT('habef)
	) name24513 (
		_w8816_,
		_w8819_,
		_w26412_,
		_w26413_,
		_w26414_
	);
	LUT3 #(
		.INIT('h2a)
	) name24514 (
		\m5_addr_i[14]_pad ,
		_w8821_,
		_w8822_,
		_w26415_
	);
	LUT3 #(
		.INIT('h2a)
	) name24515 (
		\m1_addr_i[14]_pad ,
		_w8821_,
		_w8822_,
		_w26416_
	);
	LUT4 #(
		.INIT('h57df)
	) name24516 (
		_w8816_,
		_w8819_,
		_w26415_,
		_w26416_,
		_w26417_
	);
	LUT3 #(
		.INIT('h80)
	) name24517 (
		\m0_addr_i[14]_pad ,
		_w8821_,
		_w8822_,
		_w26418_
	);
	LUT3 #(
		.INIT('h2a)
	) name24518 (
		\m7_addr_i[14]_pad ,
		_w8821_,
		_w8822_,
		_w26419_
	);
	LUT4 #(
		.INIT('h6e7f)
	) name24519 (
		_w8816_,
		_w8819_,
		_w26418_,
		_w26419_,
		_w26420_
	);
	LUT4 #(
		.INIT('h7fff)
	) name24520 (
		_w26411_,
		_w26414_,
		_w26417_,
		_w26420_,
		_w26421_
	);
	LUT3 #(
		.INIT('h2a)
	) name24521 (
		\m1_addr_i[15]_pad ,
		_w8821_,
		_w8822_,
		_w26422_
	);
	LUT3 #(
		.INIT('h80)
	) name24522 (
		\m2_addr_i[15]_pad ,
		_w8821_,
		_w8822_,
		_w26423_
	);
	LUT4 #(
		.INIT('h3b7f)
	) name24523 (
		_w8816_,
		_w8819_,
		_w26422_,
		_w26423_,
		_w26424_
	);
	LUT3 #(
		.INIT('h80)
	) name24524 (
		\m6_addr_i[15]_pad ,
		_w8821_,
		_w8822_,
		_w26425_
	);
	LUT3 #(
		.INIT('h2a)
	) name24525 (
		\m7_addr_i[15]_pad ,
		_w8821_,
		_w8822_,
		_w26426_
	);
	LUT3 #(
		.INIT('h57)
	) name24526 (
		_w8834_,
		_w26425_,
		_w26426_,
		_w26427_
	);
	LUT3 #(
		.INIT('h2a)
	) name24527 (
		\m5_addr_i[15]_pad ,
		_w8821_,
		_w8822_,
		_w26428_
	);
	LUT3 #(
		.INIT('h80)
	) name24528 (
		\m0_addr_i[15]_pad ,
		_w8821_,
		_w8822_,
		_w26429_
	);
	LUT4 #(
		.INIT('h57df)
	) name24529 (
		_w8816_,
		_w8819_,
		_w26428_,
		_w26429_,
		_w26430_
	);
	LUT3 #(
		.INIT('h2a)
	) name24530 (
		\m3_addr_i[15]_pad ,
		_w8821_,
		_w8822_,
		_w26431_
	);
	LUT3 #(
		.INIT('h80)
	) name24531 (
		\m4_addr_i[15]_pad ,
		_w8821_,
		_w8822_,
		_w26432_
	);
	LUT4 #(
		.INIT('h9dbf)
	) name24532 (
		_w8816_,
		_w8819_,
		_w26431_,
		_w26432_,
		_w26433_
	);
	LUT4 #(
		.INIT('h7fff)
	) name24533 (
		_w26424_,
		_w26427_,
		_w26430_,
		_w26433_,
		_w26434_
	);
	LUT3 #(
		.INIT('h2a)
	) name24534 (
		\m3_addr_i[16]_pad ,
		_w8821_,
		_w8822_,
		_w26435_
	);
	LUT3 #(
		.INIT('h80)
	) name24535 (
		\m4_addr_i[16]_pad ,
		_w8821_,
		_w8822_,
		_w26436_
	);
	LUT4 #(
		.INIT('h9dbf)
	) name24536 (
		_w8816_,
		_w8819_,
		_w26435_,
		_w26436_,
		_w26437_
	);
	LUT3 #(
		.INIT('h80)
	) name24537 (
		\m6_addr_i[16]_pad ,
		_w8821_,
		_w8822_,
		_w26438_
	);
	LUT3 #(
		.INIT('h2a)
	) name24538 (
		\m7_addr_i[16]_pad ,
		_w8821_,
		_w8822_,
		_w26439_
	);
	LUT3 #(
		.INIT('h57)
	) name24539 (
		_w8834_,
		_w26438_,
		_w26439_,
		_w26440_
	);
	LUT3 #(
		.INIT('h2a)
	) name24540 (
		\m5_addr_i[16]_pad ,
		_w8821_,
		_w8822_,
		_w26441_
	);
	LUT3 #(
		.INIT('h80)
	) name24541 (
		\m0_addr_i[16]_pad ,
		_w8821_,
		_w8822_,
		_w26442_
	);
	LUT4 #(
		.INIT('h57df)
	) name24542 (
		_w8816_,
		_w8819_,
		_w26441_,
		_w26442_,
		_w26443_
	);
	LUT3 #(
		.INIT('h2a)
	) name24543 (
		\m1_addr_i[16]_pad ,
		_w8821_,
		_w8822_,
		_w26444_
	);
	LUT3 #(
		.INIT('h80)
	) name24544 (
		\m2_addr_i[16]_pad ,
		_w8821_,
		_w8822_,
		_w26445_
	);
	LUT4 #(
		.INIT('h3b7f)
	) name24545 (
		_w8816_,
		_w8819_,
		_w26444_,
		_w26445_,
		_w26446_
	);
	LUT4 #(
		.INIT('h7fff)
	) name24546 (
		_w26437_,
		_w26440_,
		_w26443_,
		_w26446_,
		_w26447_
	);
	LUT3 #(
		.INIT('h80)
	) name24547 (
		\m0_addr_i[17]_pad ,
		_w8821_,
		_w8822_,
		_w26448_
	);
	LUT3 #(
		.INIT('h2a)
	) name24548 (
		\m7_addr_i[17]_pad ,
		_w8821_,
		_w8822_,
		_w26449_
	);
	LUT4 #(
		.INIT('h6e7f)
	) name24549 (
		_w8816_,
		_w8819_,
		_w26448_,
		_w26449_,
		_w26450_
	);
	LUT3 #(
		.INIT('h80)
	) name24550 (
		\m6_addr_i[17]_pad ,
		_w8821_,
		_w8822_,
		_w26451_
	);
	LUT3 #(
		.INIT('h80)
	) name24551 (
		\m2_addr_i[17]_pad ,
		_w8821_,
		_w8822_,
		_w26452_
	);
	LUT4 #(
		.INIT('habef)
	) name24552 (
		_w8816_,
		_w8819_,
		_w26451_,
		_w26452_,
		_w26453_
	);
	LUT3 #(
		.INIT('h2a)
	) name24553 (
		\m5_addr_i[17]_pad ,
		_w8821_,
		_w8822_,
		_w26454_
	);
	LUT3 #(
		.INIT('h2a)
	) name24554 (
		\m1_addr_i[17]_pad ,
		_w8821_,
		_w8822_,
		_w26455_
	);
	LUT4 #(
		.INIT('h57df)
	) name24555 (
		_w8816_,
		_w8819_,
		_w26454_,
		_w26455_,
		_w26456_
	);
	LUT3 #(
		.INIT('h2a)
	) name24556 (
		\m3_addr_i[17]_pad ,
		_w8821_,
		_w8822_,
		_w26457_
	);
	LUT3 #(
		.INIT('h80)
	) name24557 (
		\m4_addr_i[17]_pad ,
		_w8821_,
		_w8822_,
		_w26458_
	);
	LUT4 #(
		.INIT('h9dbf)
	) name24558 (
		_w8816_,
		_w8819_,
		_w26457_,
		_w26458_,
		_w26459_
	);
	LUT4 #(
		.INIT('h7fff)
	) name24559 (
		_w26450_,
		_w26453_,
		_w26456_,
		_w26459_,
		_w26460_
	);
	LUT3 #(
		.INIT('h2a)
	) name24560 (
		\m3_addr_i[18]_pad ,
		_w8821_,
		_w8822_,
		_w26461_
	);
	LUT3 #(
		.INIT('h80)
	) name24561 (
		\m4_addr_i[18]_pad ,
		_w8821_,
		_w8822_,
		_w26462_
	);
	LUT4 #(
		.INIT('h9dbf)
	) name24562 (
		_w8816_,
		_w8819_,
		_w26461_,
		_w26462_,
		_w26463_
	);
	LUT3 #(
		.INIT('h80)
	) name24563 (
		\m6_addr_i[18]_pad ,
		_w8821_,
		_w8822_,
		_w26464_
	);
	LUT3 #(
		.INIT('h2a)
	) name24564 (
		\m7_addr_i[18]_pad ,
		_w8821_,
		_w8822_,
		_w26465_
	);
	LUT3 #(
		.INIT('h57)
	) name24565 (
		_w8834_,
		_w26464_,
		_w26465_,
		_w26466_
	);
	LUT3 #(
		.INIT('h2a)
	) name24566 (
		\m5_addr_i[18]_pad ,
		_w8821_,
		_w8822_,
		_w26467_
	);
	LUT3 #(
		.INIT('h80)
	) name24567 (
		\m0_addr_i[18]_pad ,
		_w8821_,
		_w8822_,
		_w26468_
	);
	LUT4 #(
		.INIT('h57df)
	) name24568 (
		_w8816_,
		_w8819_,
		_w26467_,
		_w26468_,
		_w26469_
	);
	LUT3 #(
		.INIT('h2a)
	) name24569 (
		\m1_addr_i[18]_pad ,
		_w8821_,
		_w8822_,
		_w26470_
	);
	LUT3 #(
		.INIT('h80)
	) name24570 (
		\m2_addr_i[18]_pad ,
		_w8821_,
		_w8822_,
		_w26471_
	);
	LUT4 #(
		.INIT('h3b7f)
	) name24571 (
		_w8816_,
		_w8819_,
		_w26470_,
		_w26471_,
		_w26472_
	);
	LUT4 #(
		.INIT('h7fff)
	) name24572 (
		_w26463_,
		_w26466_,
		_w26469_,
		_w26472_,
		_w26473_
	);
	LUT3 #(
		.INIT('h2a)
	) name24573 (
		\m1_addr_i[19]_pad ,
		_w8821_,
		_w8822_,
		_w26474_
	);
	LUT3 #(
		.INIT('h80)
	) name24574 (
		\m2_addr_i[19]_pad ,
		_w8821_,
		_w8822_,
		_w26475_
	);
	LUT4 #(
		.INIT('h3b7f)
	) name24575 (
		_w8816_,
		_w8819_,
		_w26474_,
		_w26475_,
		_w26476_
	);
	LUT3 #(
		.INIT('h2a)
	) name24576 (
		\m3_addr_i[19]_pad ,
		_w8821_,
		_w8822_,
		_w26477_
	);
	LUT3 #(
		.INIT('h2a)
	) name24577 (
		\m7_addr_i[19]_pad ,
		_w8821_,
		_w8822_,
		_w26478_
	);
	LUT4 #(
		.INIT('haebf)
	) name24578 (
		_w8816_,
		_w8819_,
		_w26477_,
		_w26478_,
		_w26479_
	);
	LUT3 #(
		.INIT('h80)
	) name24579 (
		\m4_addr_i[19]_pad ,
		_w8821_,
		_w8822_,
		_w26480_
	);
	LUT3 #(
		.INIT('h80)
	) name24580 (
		\m0_addr_i[19]_pad ,
		_w8821_,
		_w8822_,
		_w26481_
	);
	LUT4 #(
		.INIT('h57df)
	) name24581 (
		_w8816_,
		_w8819_,
		_w26480_,
		_w26481_,
		_w26482_
	);
	LUT3 #(
		.INIT('h80)
	) name24582 (
		\m6_addr_i[19]_pad ,
		_w8821_,
		_w8822_,
		_w26483_
	);
	LUT3 #(
		.INIT('h2a)
	) name24583 (
		\m5_addr_i[19]_pad ,
		_w8821_,
		_w8822_,
		_w26484_
	);
	LUT4 #(
		.INIT('hcdef)
	) name24584 (
		_w8816_,
		_w8819_,
		_w26483_,
		_w26484_,
		_w26485_
	);
	LUT4 #(
		.INIT('h7fff)
	) name24585 (
		_w26476_,
		_w26479_,
		_w26482_,
		_w26485_,
		_w26486_
	);
	LUT3 #(
		.INIT('h2a)
	) name24586 (
		\m3_addr_i[1]_pad ,
		_w8821_,
		_w8822_,
		_w26487_
	);
	LUT3 #(
		.INIT('h80)
	) name24587 (
		\m4_addr_i[1]_pad ,
		_w8821_,
		_w8822_,
		_w26488_
	);
	LUT4 #(
		.INIT('h9dbf)
	) name24588 (
		_w8816_,
		_w8819_,
		_w26487_,
		_w26488_,
		_w26489_
	);
	LUT3 #(
		.INIT('h80)
	) name24589 (
		\m6_addr_i[1]_pad ,
		_w8821_,
		_w8822_,
		_w26490_
	);
	LUT3 #(
		.INIT('h2a)
	) name24590 (
		\m7_addr_i[1]_pad ,
		_w8821_,
		_w8822_,
		_w26491_
	);
	LUT3 #(
		.INIT('h57)
	) name24591 (
		_w8834_,
		_w26490_,
		_w26491_,
		_w26492_
	);
	LUT3 #(
		.INIT('h2a)
	) name24592 (
		\m5_addr_i[1]_pad ,
		_w8821_,
		_w8822_,
		_w26493_
	);
	LUT3 #(
		.INIT('h80)
	) name24593 (
		\m0_addr_i[1]_pad ,
		_w8821_,
		_w8822_,
		_w26494_
	);
	LUT4 #(
		.INIT('h57df)
	) name24594 (
		_w8816_,
		_w8819_,
		_w26493_,
		_w26494_,
		_w26495_
	);
	LUT3 #(
		.INIT('h2a)
	) name24595 (
		\m1_addr_i[1]_pad ,
		_w8821_,
		_w8822_,
		_w26496_
	);
	LUT3 #(
		.INIT('h80)
	) name24596 (
		\m2_addr_i[1]_pad ,
		_w8821_,
		_w8822_,
		_w26497_
	);
	LUT4 #(
		.INIT('h3b7f)
	) name24597 (
		_w8816_,
		_w8819_,
		_w26496_,
		_w26497_,
		_w26498_
	);
	LUT4 #(
		.INIT('h7fff)
	) name24598 (
		_w26489_,
		_w26492_,
		_w26495_,
		_w26498_,
		_w26499_
	);
	LUT3 #(
		.INIT('h80)
	) name24599 (
		\m0_addr_i[20]_pad ,
		_w8821_,
		_w8822_,
		_w26500_
	);
	LUT3 #(
		.INIT('h2a)
	) name24600 (
		\m7_addr_i[20]_pad ,
		_w8821_,
		_w8822_,
		_w26501_
	);
	LUT4 #(
		.INIT('h6e7f)
	) name24601 (
		_w8816_,
		_w8819_,
		_w26500_,
		_w26501_,
		_w26502_
	);
	LUT3 #(
		.INIT('h2a)
	) name24602 (
		\m1_addr_i[20]_pad ,
		_w8821_,
		_w8822_,
		_w26503_
	);
	LUT3 #(
		.INIT('h80)
	) name24603 (
		\m4_addr_i[20]_pad ,
		_w8821_,
		_w8822_,
		_w26504_
	);
	LUT4 #(
		.INIT('h5d7f)
	) name24604 (
		_w8816_,
		_w8819_,
		_w26503_,
		_w26504_,
		_w26505_
	);
	LUT3 #(
		.INIT('h80)
	) name24605 (
		\m2_addr_i[20]_pad ,
		_w8821_,
		_w8822_,
		_w26506_
	);
	LUT3 #(
		.INIT('h2a)
	) name24606 (
		\m3_addr_i[20]_pad ,
		_w8821_,
		_w8822_,
		_w26507_
	);
	LUT3 #(
		.INIT('h57)
	) name24607 (
		_w8828_,
		_w26506_,
		_w26507_,
		_w26508_
	);
	LUT3 #(
		.INIT('h80)
	) name24608 (
		\m6_addr_i[20]_pad ,
		_w8821_,
		_w8822_,
		_w26509_
	);
	LUT3 #(
		.INIT('h2a)
	) name24609 (
		\m5_addr_i[20]_pad ,
		_w8821_,
		_w8822_,
		_w26510_
	);
	LUT4 #(
		.INIT('hcdef)
	) name24610 (
		_w8816_,
		_w8819_,
		_w26509_,
		_w26510_,
		_w26511_
	);
	LUT4 #(
		.INIT('h7fff)
	) name24611 (
		_w26502_,
		_w26505_,
		_w26508_,
		_w26511_,
		_w26512_
	);
	LUT3 #(
		.INIT('h2a)
	) name24612 (
		\m3_addr_i[21]_pad ,
		_w8821_,
		_w8822_,
		_w26513_
	);
	LUT3 #(
		.INIT('h80)
	) name24613 (
		\m4_addr_i[21]_pad ,
		_w8821_,
		_w8822_,
		_w26514_
	);
	LUT4 #(
		.INIT('h9dbf)
	) name24614 (
		_w8816_,
		_w8819_,
		_w26513_,
		_w26514_,
		_w26515_
	);
	LUT3 #(
		.INIT('h80)
	) name24615 (
		\m6_addr_i[21]_pad ,
		_w8821_,
		_w8822_,
		_w26516_
	);
	LUT3 #(
		.INIT('h80)
	) name24616 (
		\m2_addr_i[21]_pad ,
		_w8821_,
		_w8822_,
		_w26517_
	);
	LUT4 #(
		.INIT('habef)
	) name24617 (
		_w8816_,
		_w8819_,
		_w26516_,
		_w26517_,
		_w26518_
	);
	LUT3 #(
		.INIT('h2a)
	) name24618 (
		\m5_addr_i[21]_pad ,
		_w8821_,
		_w8822_,
		_w26519_
	);
	LUT3 #(
		.INIT('h2a)
	) name24619 (
		\m1_addr_i[21]_pad ,
		_w8821_,
		_w8822_,
		_w26520_
	);
	LUT4 #(
		.INIT('h57df)
	) name24620 (
		_w8816_,
		_w8819_,
		_w26519_,
		_w26520_,
		_w26521_
	);
	LUT3 #(
		.INIT('h80)
	) name24621 (
		\m0_addr_i[21]_pad ,
		_w8821_,
		_w8822_,
		_w26522_
	);
	LUT3 #(
		.INIT('h2a)
	) name24622 (
		\m7_addr_i[21]_pad ,
		_w8821_,
		_w8822_,
		_w26523_
	);
	LUT4 #(
		.INIT('h6e7f)
	) name24623 (
		_w8816_,
		_w8819_,
		_w26522_,
		_w26523_,
		_w26524_
	);
	LUT4 #(
		.INIT('h7fff)
	) name24624 (
		_w26515_,
		_w26518_,
		_w26521_,
		_w26524_,
		_w26525_
	);
	LUT3 #(
		.INIT('h2a)
	) name24625 (
		\m1_addr_i[22]_pad ,
		_w8821_,
		_w8822_,
		_w26526_
	);
	LUT3 #(
		.INIT('h80)
	) name24626 (
		\m2_addr_i[22]_pad ,
		_w8821_,
		_w8822_,
		_w26527_
	);
	LUT4 #(
		.INIT('h3b7f)
	) name24627 (
		_w8816_,
		_w8819_,
		_w26526_,
		_w26527_,
		_w26528_
	);
	LUT3 #(
		.INIT('h2a)
	) name24628 (
		\m3_addr_i[22]_pad ,
		_w8821_,
		_w8822_,
		_w26529_
	);
	LUT3 #(
		.INIT('h2a)
	) name24629 (
		\m7_addr_i[22]_pad ,
		_w8821_,
		_w8822_,
		_w26530_
	);
	LUT4 #(
		.INIT('haebf)
	) name24630 (
		_w8816_,
		_w8819_,
		_w26529_,
		_w26530_,
		_w26531_
	);
	LUT3 #(
		.INIT('h80)
	) name24631 (
		\m4_addr_i[22]_pad ,
		_w8821_,
		_w8822_,
		_w26532_
	);
	LUT3 #(
		.INIT('h80)
	) name24632 (
		\m0_addr_i[22]_pad ,
		_w8821_,
		_w8822_,
		_w26533_
	);
	LUT4 #(
		.INIT('h57df)
	) name24633 (
		_w8816_,
		_w8819_,
		_w26532_,
		_w26533_,
		_w26534_
	);
	LUT3 #(
		.INIT('h80)
	) name24634 (
		\m6_addr_i[22]_pad ,
		_w8821_,
		_w8822_,
		_w26535_
	);
	LUT3 #(
		.INIT('h2a)
	) name24635 (
		\m5_addr_i[22]_pad ,
		_w8821_,
		_w8822_,
		_w26536_
	);
	LUT4 #(
		.INIT('hcdef)
	) name24636 (
		_w8816_,
		_w8819_,
		_w26535_,
		_w26536_,
		_w26537_
	);
	LUT4 #(
		.INIT('h7fff)
	) name24637 (
		_w26528_,
		_w26531_,
		_w26534_,
		_w26537_,
		_w26538_
	);
	LUT3 #(
		.INIT('h2a)
	) name24638 (
		\m1_addr_i[23]_pad ,
		_w8821_,
		_w8822_,
		_w26539_
	);
	LUT3 #(
		.INIT('h80)
	) name24639 (
		\m2_addr_i[23]_pad ,
		_w8821_,
		_w8822_,
		_w26540_
	);
	LUT4 #(
		.INIT('h3b7f)
	) name24640 (
		_w8816_,
		_w8819_,
		_w26539_,
		_w26540_,
		_w26541_
	);
	LUT3 #(
		.INIT('h80)
	) name24641 (
		\m6_addr_i[23]_pad ,
		_w8821_,
		_w8822_,
		_w26542_
	);
	LUT3 #(
		.INIT('h2a)
	) name24642 (
		\m7_addr_i[23]_pad ,
		_w8821_,
		_w8822_,
		_w26543_
	);
	LUT3 #(
		.INIT('h57)
	) name24643 (
		_w8834_,
		_w26542_,
		_w26543_,
		_w26544_
	);
	LUT3 #(
		.INIT('h2a)
	) name24644 (
		\m5_addr_i[23]_pad ,
		_w8821_,
		_w8822_,
		_w26545_
	);
	LUT3 #(
		.INIT('h80)
	) name24645 (
		\m0_addr_i[23]_pad ,
		_w8821_,
		_w8822_,
		_w26546_
	);
	LUT4 #(
		.INIT('h57df)
	) name24646 (
		_w8816_,
		_w8819_,
		_w26545_,
		_w26546_,
		_w26547_
	);
	LUT3 #(
		.INIT('h2a)
	) name24647 (
		\m3_addr_i[23]_pad ,
		_w8821_,
		_w8822_,
		_w26548_
	);
	LUT3 #(
		.INIT('h80)
	) name24648 (
		\m4_addr_i[23]_pad ,
		_w8821_,
		_w8822_,
		_w26549_
	);
	LUT4 #(
		.INIT('h9dbf)
	) name24649 (
		_w8816_,
		_w8819_,
		_w26548_,
		_w26549_,
		_w26550_
	);
	LUT4 #(
		.INIT('h7fff)
	) name24650 (
		_w26541_,
		_w26544_,
		_w26547_,
		_w26550_,
		_w26551_
	);
	LUT3 #(
		.INIT('h2a)
	) name24651 (
		\m1_addr_i[24]_pad ,
		_w8821_,
		_w8822_,
		_w26552_
	);
	LUT3 #(
		.INIT('h80)
	) name24652 (
		\m2_addr_i[24]_pad ,
		_w8821_,
		_w8822_,
		_w26553_
	);
	LUT4 #(
		.INIT('h3b7f)
	) name24653 (
		_w8816_,
		_w8819_,
		_w26552_,
		_w26553_,
		_w26554_
	);
	LUT3 #(
		.INIT('h2a)
	) name24654 (
		\m3_addr_i[24]_pad ,
		_w8821_,
		_w8822_,
		_w26555_
	);
	LUT3 #(
		.INIT('h2a)
	) name24655 (
		\m7_addr_i[24]_pad ,
		_w8821_,
		_w8822_,
		_w26556_
	);
	LUT4 #(
		.INIT('haebf)
	) name24656 (
		_w8816_,
		_w8819_,
		_w26555_,
		_w26556_,
		_w26557_
	);
	LUT3 #(
		.INIT('h80)
	) name24657 (
		\m4_addr_i[24]_pad ,
		_w8821_,
		_w8822_,
		_w26558_
	);
	LUT3 #(
		.INIT('h80)
	) name24658 (
		\m0_addr_i[24]_pad ,
		_w8821_,
		_w8822_,
		_w26559_
	);
	LUT4 #(
		.INIT('h57df)
	) name24659 (
		_w8816_,
		_w8819_,
		_w26558_,
		_w26559_,
		_w26560_
	);
	LUT3 #(
		.INIT('h2a)
	) name24660 (
		\m5_addr_i[24]_pad ,
		_w8821_,
		_w8822_,
		_w26561_
	);
	LUT3 #(
		.INIT('h80)
	) name24661 (
		\m6_addr_i[24]_pad ,
		_w8821_,
		_w8822_,
		_w26562_
	);
	LUT4 #(
		.INIT('hcedf)
	) name24662 (
		_w8816_,
		_w8819_,
		_w26561_,
		_w26562_,
		_w26563_
	);
	LUT4 #(
		.INIT('h7fff)
	) name24663 (
		_w26554_,
		_w26557_,
		_w26560_,
		_w26563_,
		_w26564_
	);
	LUT3 #(
		.INIT('h2a)
	) name24664 (
		\m3_addr_i[25]_pad ,
		_w8821_,
		_w8822_,
		_w26565_
	);
	LUT3 #(
		.INIT('h80)
	) name24665 (
		\m4_addr_i[25]_pad ,
		_w8821_,
		_w8822_,
		_w26566_
	);
	LUT4 #(
		.INIT('h9dbf)
	) name24666 (
		_w8816_,
		_w8819_,
		_w26565_,
		_w26566_,
		_w26567_
	);
	LUT3 #(
		.INIT('h2a)
	) name24667 (
		\m5_addr_i[25]_pad ,
		_w8821_,
		_w8822_,
		_w26568_
	);
	LUT3 #(
		.INIT('h80)
	) name24668 (
		\m2_addr_i[25]_pad ,
		_w8821_,
		_w8822_,
		_w26569_
	);
	LUT4 #(
		.INIT('h9bdf)
	) name24669 (
		_w8816_,
		_w8819_,
		_w26568_,
		_w26569_,
		_w26570_
	);
	LUT3 #(
		.INIT('h80)
	) name24670 (
		\m6_addr_i[25]_pad ,
		_w8821_,
		_w8822_,
		_w26571_
	);
	LUT3 #(
		.INIT('h2a)
	) name24671 (
		\m1_addr_i[25]_pad ,
		_w8821_,
		_w8822_,
		_w26572_
	);
	LUT4 #(
		.INIT('h67ef)
	) name24672 (
		_w8816_,
		_w8819_,
		_w26571_,
		_w26572_,
		_w26573_
	);
	LUT3 #(
		.INIT('h80)
	) name24673 (
		\m0_addr_i[25]_pad ,
		_w8821_,
		_w8822_,
		_w26574_
	);
	LUT3 #(
		.INIT('h2a)
	) name24674 (
		\m7_addr_i[25]_pad ,
		_w8821_,
		_w8822_,
		_w26575_
	);
	LUT4 #(
		.INIT('h6e7f)
	) name24675 (
		_w8816_,
		_w8819_,
		_w26574_,
		_w26575_,
		_w26576_
	);
	LUT4 #(
		.INIT('h7fff)
	) name24676 (
		_w26567_,
		_w26570_,
		_w26573_,
		_w26576_,
		_w26577_
	);
	LUT3 #(
		.INIT('h80)
	) name24677 (
		\m0_addr_i[26]_pad ,
		_w8821_,
		_w8822_,
		_w26578_
	);
	LUT3 #(
		.INIT('h2a)
	) name24678 (
		\m7_addr_i[26]_pad ,
		_w8821_,
		_w8822_,
		_w26579_
	);
	LUT4 #(
		.INIT('h6e7f)
	) name24679 (
		_w8816_,
		_w8819_,
		_w26578_,
		_w26579_,
		_w26580_
	);
	LUT3 #(
		.INIT('h2a)
	) name24680 (
		\m5_addr_i[26]_pad ,
		_w8821_,
		_w8822_,
		_w26581_
	);
	LUT3 #(
		.INIT('h80)
	) name24681 (
		\m2_addr_i[26]_pad ,
		_w8821_,
		_w8822_,
		_w26582_
	);
	LUT4 #(
		.INIT('h9bdf)
	) name24682 (
		_w8816_,
		_w8819_,
		_w26581_,
		_w26582_,
		_w26583_
	);
	LUT3 #(
		.INIT('h80)
	) name24683 (
		\m6_addr_i[26]_pad ,
		_w8821_,
		_w8822_,
		_w26584_
	);
	LUT3 #(
		.INIT('h2a)
	) name24684 (
		\m1_addr_i[26]_pad ,
		_w8821_,
		_w8822_,
		_w26585_
	);
	LUT4 #(
		.INIT('h67ef)
	) name24685 (
		_w8816_,
		_w8819_,
		_w26584_,
		_w26585_,
		_w26586_
	);
	LUT3 #(
		.INIT('h2a)
	) name24686 (
		\m3_addr_i[26]_pad ,
		_w8821_,
		_w8822_,
		_w26587_
	);
	LUT3 #(
		.INIT('h80)
	) name24687 (
		\m4_addr_i[26]_pad ,
		_w8821_,
		_w8822_,
		_w26588_
	);
	LUT4 #(
		.INIT('h9dbf)
	) name24688 (
		_w8816_,
		_w8819_,
		_w26587_,
		_w26588_,
		_w26589_
	);
	LUT4 #(
		.INIT('h7fff)
	) name24689 (
		_w26580_,
		_w26583_,
		_w26586_,
		_w26589_,
		_w26590_
	);
	LUT3 #(
		.INIT('h2a)
	) name24690 (
		\m3_addr_i[27]_pad ,
		_w8821_,
		_w8822_,
		_w26591_
	);
	LUT3 #(
		.INIT('h80)
	) name24691 (
		\m4_addr_i[27]_pad ,
		_w8821_,
		_w8822_,
		_w26592_
	);
	LUT4 #(
		.INIT('h9dbf)
	) name24692 (
		_w8816_,
		_w8819_,
		_w26591_,
		_w26592_,
		_w26593_
	);
	LUT3 #(
		.INIT('h2a)
	) name24693 (
		\m5_addr_i[27]_pad ,
		_w8821_,
		_w8822_,
		_w26594_
	);
	LUT3 #(
		.INIT('h80)
	) name24694 (
		\m2_addr_i[27]_pad ,
		_w8821_,
		_w8822_,
		_w26595_
	);
	LUT4 #(
		.INIT('h9bdf)
	) name24695 (
		_w8816_,
		_w8819_,
		_w26594_,
		_w26595_,
		_w26596_
	);
	LUT3 #(
		.INIT('h80)
	) name24696 (
		\m6_addr_i[27]_pad ,
		_w8821_,
		_w8822_,
		_w26597_
	);
	LUT3 #(
		.INIT('h2a)
	) name24697 (
		\m1_addr_i[27]_pad ,
		_w8821_,
		_w8822_,
		_w26598_
	);
	LUT4 #(
		.INIT('h67ef)
	) name24698 (
		_w8816_,
		_w8819_,
		_w26597_,
		_w26598_,
		_w26599_
	);
	LUT3 #(
		.INIT('h80)
	) name24699 (
		\m0_addr_i[27]_pad ,
		_w8821_,
		_w8822_,
		_w26600_
	);
	LUT3 #(
		.INIT('h2a)
	) name24700 (
		\m7_addr_i[27]_pad ,
		_w8821_,
		_w8822_,
		_w26601_
	);
	LUT4 #(
		.INIT('h6e7f)
	) name24701 (
		_w8816_,
		_w8819_,
		_w26600_,
		_w26601_,
		_w26602_
	);
	LUT4 #(
		.INIT('h7fff)
	) name24702 (
		_w26593_,
		_w26596_,
		_w26599_,
		_w26602_,
		_w26603_
	);
	LUT3 #(
		.INIT('h2a)
	) name24703 (
		\m3_addr_i[28]_pad ,
		_w8821_,
		_w8822_,
		_w26604_
	);
	LUT3 #(
		.INIT('h80)
	) name24704 (
		\m4_addr_i[28]_pad ,
		_w8821_,
		_w8822_,
		_w26605_
	);
	LUT4 #(
		.INIT('h9dbf)
	) name24705 (
		_w8816_,
		_w8819_,
		_w26604_,
		_w26605_,
		_w26606_
	);
	LUT3 #(
		.INIT('h2a)
	) name24706 (
		\m5_addr_i[28]_pad ,
		_w8821_,
		_w8822_,
		_w26607_
	);
	LUT3 #(
		.INIT('h2a)
	) name24707 (
		\m7_addr_i[28]_pad ,
		_w8821_,
		_w8822_,
		_w26608_
	);
	LUT4 #(
		.INIT('hcedf)
	) name24708 (
		_w8816_,
		_w8819_,
		_w26607_,
		_w26608_,
		_w26609_
	);
	LUT3 #(
		.INIT('h80)
	) name24709 (
		\m6_addr_i[28]_pad ,
		_w8821_,
		_w8822_,
		_w26610_
	);
	LUT3 #(
		.INIT('h80)
	) name24710 (
		\m0_addr_i[28]_pad ,
		_w8821_,
		_w8822_,
		_w26611_
	);
	LUT4 #(
		.INIT('h67ef)
	) name24711 (
		_w8816_,
		_w8819_,
		_w26610_,
		_w26611_,
		_w26612_
	);
	LUT3 #(
		.INIT('h2a)
	) name24712 (
		\m1_addr_i[28]_pad ,
		_w8821_,
		_w8822_,
		_w26613_
	);
	LUT3 #(
		.INIT('h80)
	) name24713 (
		\m2_addr_i[28]_pad ,
		_w8821_,
		_w8822_,
		_w26614_
	);
	LUT4 #(
		.INIT('h3b7f)
	) name24714 (
		_w8816_,
		_w8819_,
		_w26613_,
		_w26614_,
		_w26615_
	);
	LUT4 #(
		.INIT('h7fff)
	) name24715 (
		_w26606_,
		_w26609_,
		_w26612_,
		_w26615_,
		_w26616_
	);
	LUT3 #(
		.INIT('h2a)
	) name24716 (
		\m1_addr_i[29]_pad ,
		_w8821_,
		_w8822_,
		_w26617_
	);
	LUT3 #(
		.INIT('h80)
	) name24717 (
		\m2_addr_i[29]_pad ,
		_w8821_,
		_w8822_,
		_w26618_
	);
	LUT4 #(
		.INIT('h3b7f)
	) name24718 (
		_w8816_,
		_w8819_,
		_w26617_,
		_w26618_,
		_w26619_
	);
	LUT3 #(
		.INIT('h2a)
	) name24719 (
		\m3_addr_i[29]_pad ,
		_w8821_,
		_w8822_,
		_w26620_
	);
	LUT3 #(
		.INIT('h80)
	) name24720 (
		\m6_addr_i[29]_pad ,
		_w8821_,
		_w8822_,
		_w26621_
	);
	LUT4 #(
		.INIT('haebf)
	) name24721 (
		_w8816_,
		_w8819_,
		_w26620_,
		_w26621_,
		_w26622_
	);
	LUT3 #(
		.INIT('h80)
	) name24722 (
		\m4_addr_i[29]_pad ,
		_w8821_,
		_w8822_,
		_w26623_
	);
	LUT3 #(
		.INIT('h2a)
	) name24723 (
		\m5_addr_i[29]_pad ,
		_w8821_,
		_w8822_,
		_w26624_
	);
	LUT3 #(
		.INIT('h57)
	) name24724 (
		_w8840_,
		_w26623_,
		_w26624_,
		_w26625_
	);
	LUT3 #(
		.INIT('h80)
	) name24725 (
		\m0_addr_i[29]_pad ,
		_w8821_,
		_w8822_,
		_w26626_
	);
	LUT3 #(
		.INIT('h2a)
	) name24726 (
		\m7_addr_i[29]_pad ,
		_w8821_,
		_w8822_,
		_w26627_
	);
	LUT4 #(
		.INIT('h6e7f)
	) name24727 (
		_w8816_,
		_w8819_,
		_w26626_,
		_w26627_,
		_w26628_
	);
	LUT4 #(
		.INIT('h7fff)
	) name24728 (
		_w26619_,
		_w26622_,
		_w26625_,
		_w26628_,
		_w26629_
	);
	LUT3 #(
		.INIT('h80)
	) name24729 (
		\m6_addr_i[2]_pad ,
		_w8821_,
		_w8822_,
		_w26630_
	);
	LUT3 #(
		.INIT('h2a)
	) name24730 (
		\m5_addr_i[2]_pad ,
		_w8821_,
		_w8822_,
		_w26631_
	);
	LUT4 #(
		.INIT('hcdef)
	) name24731 (
		_w8816_,
		_w8819_,
		_w26630_,
		_w26631_,
		_w26632_
	);
	LUT3 #(
		.INIT('h2a)
	) name24732 (
		\m1_addr_i[2]_pad ,
		_w8821_,
		_w8822_,
		_w26633_
	);
	LUT3 #(
		.INIT('h80)
	) name24733 (
		\m4_addr_i[2]_pad ,
		_w8821_,
		_w8822_,
		_w26634_
	);
	LUT4 #(
		.INIT('h5d7f)
	) name24734 (
		_w8816_,
		_w8819_,
		_w26633_,
		_w26634_,
		_w26635_
	);
	LUT3 #(
		.INIT('h80)
	) name24735 (
		\m2_addr_i[2]_pad ,
		_w8821_,
		_w8822_,
		_w26636_
	);
	LUT3 #(
		.INIT('h2a)
	) name24736 (
		\m3_addr_i[2]_pad ,
		_w8821_,
		_w8822_,
		_w26637_
	);
	LUT3 #(
		.INIT('h57)
	) name24737 (
		_w8828_,
		_w26636_,
		_w26637_,
		_w26638_
	);
	LUT3 #(
		.INIT('h80)
	) name24738 (
		\m0_addr_i[2]_pad ,
		_w8821_,
		_w8822_,
		_w26639_
	);
	LUT3 #(
		.INIT('h2a)
	) name24739 (
		\m7_addr_i[2]_pad ,
		_w8821_,
		_w8822_,
		_w26640_
	);
	LUT4 #(
		.INIT('h6e7f)
	) name24740 (
		_w8816_,
		_w8819_,
		_w26639_,
		_w26640_,
		_w26641_
	);
	LUT4 #(
		.INIT('h7fff)
	) name24741 (
		_w26632_,
		_w26635_,
		_w26638_,
		_w26641_,
		_w26642_
	);
	LUT3 #(
		.INIT('h2a)
	) name24742 (
		\m3_addr_i[30]_pad ,
		_w8821_,
		_w8822_,
		_w26643_
	);
	LUT3 #(
		.INIT('h80)
	) name24743 (
		\m4_addr_i[30]_pad ,
		_w8821_,
		_w8822_,
		_w26644_
	);
	LUT4 #(
		.INIT('h9dbf)
	) name24744 (
		_w8816_,
		_w8819_,
		_w26643_,
		_w26644_,
		_w26645_
	);
	LUT3 #(
		.INIT('h2a)
	) name24745 (
		\m5_addr_i[30]_pad ,
		_w8821_,
		_w8822_,
		_w26646_
	);
	LUT3 #(
		.INIT('h2a)
	) name24746 (
		\m7_addr_i[30]_pad ,
		_w8821_,
		_w8822_,
		_w26647_
	);
	LUT4 #(
		.INIT('hcedf)
	) name24747 (
		_w8816_,
		_w8819_,
		_w26646_,
		_w26647_,
		_w26648_
	);
	LUT3 #(
		.INIT('h80)
	) name24748 (
		\m6_addr_i[30]_pad ,
		_w8821_,
		_w8822_,
		_w26649_
	);
	LUT3 #(
		.INIT('h80)
	) name24749 (
		\m0_addr_i[30]_pad ,
		_w8821_,
		_w8822_,
		_w26650_
	);
	LUT4 #(
		.INIT('h67ef)
	) name24750 (
		_w8816_,
		_w8819_,
		_w26649_,
		_w26650_,
		_w26651_
	);
	LUT3 #(
		.INIT('h2a)
	) name24751 (
		\m1_addr_i[30]_pad ,
		_w8821_,
		_w8822_,
		_w26652_
	);
	LUT3 #(
		.INIT('h80)
	) name24752 (
		\m2_addr_i[30]_pad ,
		_w8821_,
		_w8822_,
		_w26653_
	);
	LUT4 #(
		.INIT('h3b7f)
	) name24753 (
		_w8816_,
		_w8819_,
		_w26652_,
		_w26653_,
		_w26654_
	);
	LUT4 #(
		.INIT('h7fff)
	) name24754 (
		_w26645_,
		_w26648_,
		_w26651_,
		_w26654_,
		_w26655_
	);
	LUT3 #(
		.INIT('h2a)
	) name24755 (
		\m1_addr_i[31]_pad ,
		_w8821_,
		_w8822_,
		_w26656_
	);
	LUT3 #(
		.INIT('h80)
	) name24756 (
		\m2_addr_i[31]_pad ,
		_w8821_,
		_w8822_,
		_w26657_
	);
	LUT4 #(
		.INIT('h3b7f)
	) name24757 (
		_w8816_,
		_w8819_,
		_w26656_,
		_w26657_,
		_w26658_
	);
	LUT3 #(
		.INIT('h2a)
	) name24758 (
		\m5_addr_i[31]_pad ,
		_w8821_,
		_w8822_,
		_w26659_
	);
	LUT3 #(
		.INIT('h2a)
	) name24759 (
		\m7_addr_i[31]_pad ,
		_w8821_,
		_w8822_,
		_w26660_
	);
	LUT4 #(
		.INIT('hcedf)
	) name24760 (
		_w8816_,
		_w8819_,
		_w26659_,
		_w26660_,
		_w26661_
	);
	LUT3 #(
		.INIT('h80)
	) name24761 (
		\m6_addr_i[31]_pad ,
		_w8821_,
		_w8822_,
		_w26662_
	);
	LUT3 #(
		.INIT('h80)
	) name24762 (
		\m0_addr_i[31]_pad ,
		_w8821_,
		_w8822_,
		_w26663_
	);
	LUT4 #(
		.INIT('h67ef)
	) name24763 (
		_w8816_,
		_w8819_,
		_w26662_,
		_w26663_,
		_w26664_
	);
	LUT3 #(
		.INIT('h2a)
	) name24764 (
		\m3_addr_i[31]_pad ,
		_w8821_,
		_w8822_,
		_w26665_
	);
	LUT3 #(
		.INIT('h80)
	) name24765 (
		\m4_addr_i[31]_pad ,
		_w8821_,
		_w8822_,
		_w26666_
	);
	LUT4 #(
		.INIT('h9dbf)
	) name24766 (
		_w8816_,
		_w8819_,
		_w26665_,
		_w26666_,
		_w26667_
	);
	LUT4 #(
		.INIT('h7fff)
	) name24767 (
		_w26658_,
		_w26661_,
		_w26664_,
		_w26667_,
		_w26668_
	);
	LUT3 #(
		.INIT('h2a)
	) name24768 (
		\m3_addr_i[3]_pad ,
		_w8821_,
		_w8822_,
		_w26669_
	);
	LUT3 #(
		.INIT('h80)
	) name24769 (
		\m4_addr_i[3]_pad ,
		_w8821_,
		_w8822_,
		_w26670_
	);
	LUT4 #(
		.INIT('h9dbf)
	) name24770 (
		_w8816_,
		_w8819_,
		_w26669_,
		_w26670_,
		_w26671_
	);
	LUT3 #(
		.INIT('h80)
	) name24771 (
		\m6_addr_i[3]_pad ,
		_w8821_,
		_w8822_,
		_w26672_
	);
	LUT3 #(
		.INIT('h80)
	) name24772 (
		\m2_addr_i[3]_pad ,
		_w8821_,
		_w8822_,
		_w26673_
	);
	LUT4 #(
		.INIT('habef)
	) name24773 (
		_w8816_,
		_w8819_,
		_w26672_,
		_w26673_,
		_w26674_
	);
	LUT3 #(
		.INIT('h2a)
	) name24774 (
		\m5_addr_i[3]_pad ,
		_w8821_,
		_w8822_,
		_w26675_
	);
	LUT3 #(
		.INIT('h2a)
	) name24775 (
		\m1_addr_i[3]_pad ,
		_w8821_,
		_w8822_,
		_w26676_
	);
	LUT4 #(
		.INIT('h57df)
	) name24776 (
		_w8816_,
		_w8819_,
		_w26675_,
		_w26676_,
		_w26677_
	);
	LUT3 #(
		.INIT('h80)
	) name24777 (
		\m0_addr_i[3]_pad ,
		_w8821_,
		_w8822_,
		_w26678_
	);
	LUT3 #(
		.INIT('h2a)
	) name24778 (
		\m7_addr_i[3]_pad ,
		_w8821_,
		_w8822_,
		_w26679_
	);
	LUT4 #(
		.INIT('h6e7f)
	) name24779 (
		_w8816_,
		_w8819_,
		_w26678_,
		_w26679_,
		_w26680_
	);
	LUT4 #(
		.INIT('h7fff)
	) name24780 (
		_w26671_,
		_w26674_,
		_w26677_,
		_w26680_,
		_w26681_
	);
	LUT3 #(
		.INIT('h2a)
	) name24781 (
		\m1_addr_i[4]_pad ,
		_w8821_,
		_w8822_,
		_w26682_
	);
	LUT3 #(
		.INIT('h80)
	) name24782 (
		\m2_addr_i[4]_pad ,
		_w8821_,
		_w8822_,
		_w26683_
	);
	LUT4 #(
		.INIT('h3b7f)
	) name24783 (
		_w8816_,
		_w8819_,
		_w26682_,
		_w26683_,
		_w26684_
	);
	LUT3 #(
		.INIT('h80)
	) name24784 (
		\m6_addr_i[4]_pad ,
		_w8821_,
		_w8822_,
		_w26685_
	);
	LUT3 #(
		.INIT('h2a)
	) name24785 (
		\m7_addr_i[4]_pad ,
		_w8821_,
		_w8822_,
		_w26686_
	);
	LUT3 #(
		.INIT('h57)
	) name24786 (
		_w8834_,
		_w26685_,
		_w26686_,
		_w26687_
	);
	LUT3 #(
		.INIT('h2a)
	) name24787 (
		\m5_addr_i[4]_pad ,
		_w8821_,
		_w8822_,
		_w26688_
	);
	LUT3 #(
		.INIT('h80)
	) name24788 (
		\m0_addr_i[4]_pad ,
		_w8821_,
		_w8822_,
		_w26689_
	);
	LUT4 #(
		.INIT('h57df)
	) name24789 (
		_w8816_,
		_w8819_,
		_w26688_,
		_w26689_,
		_w26690_
	);
	LUT3 #(
		.INIT('h2a)
	) name24790 (
		\m3_addr_i[4]_pad ,
		_w8821_,
		_w8822_,
		_w26691_
	);
	LUT3 #(
		.INIT('h80)
	) name24791 (
		\m4_addr_i[4]_pad ,
		_w8821_,
		_w8822_,
		_w26692_
	);
	LUT4 #(
		.INIT('h9dbf)
	) name24792 (
		_w8816_,
		_w8819_,
		_w26691_,
		_w26692_,
		_w26693_
	);
	LUT4 #(
		.INIT('h7fff)
	) name24793 (
		_w26684_,
		_w26687_,
		_w26690_,
		_w26693_,
		_w26694_
	);
	LUT3 #(
		.INIT('h2a)
	) name24794 (
		\m3_addr_i[5]_pad ,
		_w8821_,
		_w8822_,
		_w26695_
	);
	LUT3 #(
		.INIT('h80)
	) name24795 (
		\m4_addr_i[5]_pad ,
		_w8821_,
		_w8822_,
		_w26696_
	);
	LUT4 #(
		.INIT('h9dbf)
	) name24796 (
		_w8816_,
		_w8819_,
		_w26695_,
		_w26696_,
		_w26697_
	);
	LUT3 #(
		.INIT('h80)
	) name24797 (
		\m6_addr_i[5]_pad ,
		_w8821_,
		_w8822_,
		_w26698_
	);
	LUT3 #(
		.INIT('h80)
	) name24798 (
		\m2_addr_i[5]_pad ,
		_w8821_,
		_w8822_,
		_w26699_
	);
	LUT4 #(
		.INIT('habef)
	) name24799 (
		_w8816_,
		_w8819_,
		_w26698_,
		_w26699_,
		_w26700_
	);
	LUT3 #(
		.INIT('h2a)
	) name24800 (
		\m5_addr_i[5]_pad ,
		_w8821_,
		_w8822_,
		_w26701_
	);
	LUT3 #(
		.INIT('h2a)
	) name24801 (
		\m1_addr_i[5]_pad ,
		_w8821_,
		_w8822_,
		_w26702_
	);
	LUT4 #(
		.INIT('h57df)
	) name24802 (
		_w8816_,
		_w8819_,
		_w26701_,
		_w26702_,
		_w26703_
	);
	LUT3 #(
		.INIT('h80)
	) name24803 (
		\m0_addr_i[5]_pad ,
		_w8821_,
		_w8822_,
		_w26704_
	);
	LUT3 #(
		.INIT('h2a)
	) name24804 (
		\m7_addr_i[5]_pad ,
		_w8821_,
		_w8822_,
		_w26705_
	);
	LUT4 #(
		.INIT('h6e7f)
	) name24805 (
		_w8816_,
		_w8819_,
		_w26704_,
		_w26705_,
		_w26706_
	);
	LUT4 #(
		.INIT('h7fff)
	) name24806 (
		_w26697_,
		_w26700_,
		_w26703_,
		_w26706_,
		_w26707_
	);
	LUT3 #(
		.INIT('h2a)
	) name24807 (
		\m3_addr_i[6]_pad ,
		_w8821_,
		_w8822_,
		_w26708_
	);
	LUT3 #(
		.INIT('h80)
	) name24808 (
		\m4_addr_i[6]_pad ,
		_w8821_,
		_w8822_,
		_w26709_
	);
	LUT4 #(
		.INIT('h9dbf)
	) name24809 (
		_w8816_,
		_w8819_,
		_w26708_,
		_w26709_,
		_w26710_
	);
	LUT3 #(
		.INIT('h80)
	) name24810 (
		\m6_addr_i[6]_pad ,
		_w8821_,
		_w8822_,
		_w26711_
	);
	LUT3 #(
		.INIT('h80)
	) name24811 (
		\m2_addr_i[6]_pad ,
		_w8821_,
		_w8822_,
		_w26712_
	);
	LUT4 #(
		.INIT('habef)
	) name24812 (
		_w8816_,
		_w8819_,
		_w26711_,
		_w26712_,
		_w26713_
	);
	LUT3 #(
		.INIT('h2a)
	) name24813 (
		\m5_addr_i[6]_pad ,
		_w8821_,
		_w8822_,
		_w26714_
	);
	LUT3 #(
		.INIT('h2a)
	) name24814 (
		\m1_addr_i[6]_pad ,
		_w8821_,
		_w8822_,
		_w26715_
	);
	LUT4 #(
		.INIT('h57df)
	) name24815 (
		_w8816_,
		_w8819_,
		_w26714_,
		_w26715_,
		_w26716_
	);
	LUT3 #(
		.INIT('h80)
	) name24816 (
		\m0_addr_i[6]_pad ,
		_w8821_,
		_w8822_,
		_w26717_
	);
	LUT3 #(
		.INIT('h2a)
	) name24817 (
		\m7_addr_i[6]_pad ,
		_w8821_,
		_w8822_,
		_w26718_
	);
	LUT4 #(
		.INIT('h6e7f)
	) name24818 (
		_w8816_,
		_w8819_,
		_w26717_,
		_w26718_,
		_w26719_
	);
	LUT4 #(
		.INIT('h7fff)
	) name24819 (
		_w26710_,
		_w26713_,
		_w26716_,
		_w26719_,
		_w26720_
	);
	LUT3 #(
		.INIT('h2a)
	) name24820 (
		\m3_addr_i[7]_pad ,
		_w8821_,
		_w8822_,
		_w26721_
	);
	LUT3 #(
		.INIT('h80)
	) name24821 (
		\m4_addr_i[7]_pad ,
		_w8821_,
		_w8822_,
		_w26722_
	);
	LUT4 #(
		.INIT('h9dbf)
	) name24822 (
		_w8816_,
		_w8819_,
		_w26721_,
		_w26722_,
		_w26723_
	);
	LUT3 #(
		.INIT('h80)
	) name24823 (
		\m6_addr_i[7]_pad ,
		_w8821_,
		_w8822_,
		_w26724_
	);
	LUT3 #(
		.INIT('h80)
	) name24824 (
		\m2_addr_i[7]_pad ,
		_w8821_,
		_w8822_,
		_w26725_
	);
	LUT4 #(
		.INIT('habef)
	) name24825 (
		_w8816_,
		_w8819_,
		_w26724_,
		_w26725_,
		_w26726_
	);
	LUT3 #(
		.INIT('h2a)
	) name24826 (
		\m5_addr_i[7]_pad ,
		_w8821_,
		_w8822_,
		_w26727_
	);
	LUT3 #(
		.INIT('h2a)
	) name24827 (
		\m1_addr_i[7]_pad ,
		_w8821_,
		_w8822_,
		_w26728_
	);
	LUT4 #(
		.INIT('h57df)
	) name24828 (
		_w8816_,
		_w8819_,
		_w26727_,
		_w26728_,
		_w26729_
	);
	LUT3 #(
		.INIT('h80)
	) name24829 (
		\m0_addr_i[7]_pad ,
		_w8821_,
		_w8822_,
		_w26730_
	);
	LUT3 #(
		.INIT('h2a)
	) name24830 (
		\m7_addr_i[7]_pad ,
		_w8821_,
		_w8822_,
		_w26731_
	);
	LUT4 #(
		.INIT('h6e7f)
	) name24831 (
		_w8816_,
		_w8819_,
		_w26730_,
		_w26731_,
		_w26732_
	);
	LUT4 #(
		.INIT('h7fff)
	) name24832 (
		_w26723_,
		_w26726_,
		_w26729_,
		_w26732_,
		_w26733_
	);
	LUT3 #(
		.INIT('h80)
	) name24833 (
		\m6_addr_i[8]_pad ,
		_w8821_,
		_w8822_,
		_w26734_
	);
	LUT3 #(
		.INIT('h2a)
	) name24834 (
		\m5_addr_i[8]_pad ,
		_w8821_,
		_w8822_,
		_w26735_
	);
	LUT4 #(
		.INIT('hcdef)
	) name24835 (
		_w8816_,
		_w8819_,
		_w26734_,
		_w26735_,
		_w26736_
	);
	LUT3 #(
		.INIT('h80)
	) name24836 (
		\m0_addr_i[8]_pad ,
		_w8821_,
		_w8822_,
		_w26737_
	);
	LUT3 #(
		.INIT('h80)
	) name24837 (
		\m4_addr_i[8]_pad ,
		_w8821_,
		_w8822_,
		_w26738_
	);
	LUT4 #(
		.INIT('h5d7f)
	) name24838 (
		_w8816_,
		_w8819_,
		_w26737_,
		_w26738_,
		_w26739_
	);
	LUT3 #(
		.INIT('h2a)
	) name24839 (
		\m7_addr_i[8]_pad ,
		_w8821_,
		_w8822_,
		_w26740_
	);
	LUT3 #(
		.INIT('h2a)
	) name24840 (
		\m3_addr_i[8]_pad ,
		_w8821_,
		_w8822_,
		_w26741_
	);
	LUT4 #(
		.INIT('habef)
	) name24841 (
		_w8816_,
		_w8819_,
		_w26740_,
		_w26741_,
		_w26742_
	);
	LUT3 #(
		.INIT('h2a)
	) name24842 (
		\m1_addr_i[8]_pad ,
		_w8821_,
		_w8822_,
		_w26743_
	);
	LUT3 #(
		.INIT('h80)
	) name24843 (
		\m2_addr_i[8]_pad ,
		_w8821_,
		_w8822_,
		_w26744_
	);
	LUT4 #(
		.INIT('h3b7f)
	) name24844 (
		_w8816_,
		_w8819_,
		_w26743_,
		_w26744_,
		_w26745_
	);
	LUT4 #(
		.INIT('h7fff)
	) name24845 (
		_w26736_,
		_w26739_,
		_w26742_,
		_w26745_,
		_w26746_
	);
	LUT3 #(
		.INIT('h2a)
	) name24846 (
		\m3_addr_i[9]_pad ,
		_w8821_,
		_w8822_,
		_w26747_
	);
	LUT3 #(
		.INIT('h80)
	) name24847 (
		\m4_addr_i[9]_pad ,
		_w8821_,
		_w8822_,
		_w26748_
	);
	LUT4 #(
		.INIT('h9dbf)
	) name24848 (
		_w8816_,
		_w8819_,
		_w26747_,
		_w26748_,
		_w26749_
	);
	LUT3 #(
		.INIT('h80)
	) name24849 (
		\m6_addr_i[9]_pad ,
		_w8821_,
		_w8822_,
		_w26750_
	);
	LUT3 #(
		.INIT('h80)
	) name24850 (
		\m2_addr_i[9]_pad ,
		_w8821_,
		_w8822_,
		_w26751_
	);
	LUT4 #(
		.INIT('habef)
	) name24851 (
		_w8816_,
		_w8819_,
		_w26750_,
		_w26751_,
		_w26752_
	);
	LUT3 #(
		.INIT('h2a)
	) name24852 (
		\m5_addr_i[9]_pad ,
		_w8821_,
		_w8822_,
		_w26753_
	);
	LUT3 #(
		.INIT('h2a)
	) name24853 (
		\m1_addr_i[9]_pad ,
		_w8821_,
		_w8822_,
		_w26754_
	);
	LUT4 #(
		.INIT('h57df)
	) name24854 (
		_w8816_,
		_w8819_,
		_w26753_,
		_w26754_,
		_w26755_
	);
	LUT3 #(
		.INIT('h80)
	) name24855 (
		\m0_addr_i[9]_pad ,
		_w8821_,
		_w8822_,
		_w26756_
	);
	LUT3 #(
		.INIT('h2a)
	) name24856 (
		\m7_addr_i[9]_pad ,
		_w8821_,
		_w8822_,
		_w26757_
	);
	LUT4 #(
		.INIT('h6e7f)
	) name24857 (
		_w8816_,
		_w8819_,
		_w26756_,
		_w26757_,
		_w26758_
	);
	LUT4 #(
		.INIT('h7fff)
	) name24858 (
		_w26749_,
		_w26752_,
		_w26755_,
		_w26758_,
		_w26759_
	);
	LUT3 #(
		.INIT('h2a)
	) name24859 (
		\m1_data_i[0]_pad ,
		_w8821_,
		_w8822_,
		_w26760_
	);
	LUT3 #(
		.INIT('h80)
	) name24860 (
		\m2_data_i[0]_pad ,
		_w8821_,
		_w8822_,
		_w26761_
	);
	LUT4 #(
		.INIT('h3b7f)
	) name24861 (
		_w8816_,
		_w8819_,
		_w26760_,
		_w26761_,
		_w26762_
	);
	LUT3 #(
		.INIT('h2a)
	) name24862 (
		\m3_data_i[0]_pad ,
		_w8821_,
		_w8822_,
		_w26763_
	);
	LUT3 #(
		.INIT('h2a)
	) name24863 (
		\m7_data_i[0]_pad ,
		_w8821_,
		_w8822_,
		_w26764_
	);
	LUT4 #(
		.INIT('haebf)
	) name24864 (
		_w8816_,
		_w8819_,
		_w26763_,
		_w26764_,
		_w26765_
	);
	LUT3 #(
		.INIT('h80)
	) name24865 (
		\m4_data_i[0]_pad ,
		_w8821_,
		_w8822_,
		_w26766_
	);
	LUT3 #(
		.INIT('h80)
	) name24866 (
		\m0_data_i[0]_pad ,
		_w8821_,
		_w8822_,
		_w26767_
	);
	LUT4 #(
		.INIT('h57df)
	) name24867 (
		_w8816_,
		_w8819_,
		_w26766_,
		_w26767_,
		_w26768_
	);
	LUT3 #(
		.INIT('h80)
	) name24868 (
		\m6_data_i[0]_pad ,
		_w8821_,
		_w8822_,
		_w26769_
	);
	LUT3 #(
		.INIT('h2a)
	) name24869 (
		\m5_data_i[0]_pad ,
		_w8821_,
		_w8822_,
		_w26770_
	);
	LUT4 #(
		.INIT('hcdef)
	) name24870 (
		_w8816_,
		_w8819_,
		_w26769_,
		_w26770_,
		_w26771_
	);
	LUT4 #(
		.INIT('h7fff)
	) name24871 (
		_w26762_,
		_w26765_,
		_w26768_,
		_w26771_,
		_w26772_
	);
	LUT3 #(
		.INIT('h2a)
	) name24872 (
		\m3_data_i[10]_pad ,
		_w8821_,
		_w8822_,
		_w26773_
	);
	LUT3 #(
		.INIT('h80)
	) name24873 (
		\m4_data_i[10]_pad ,
		_w8821_,
		_w8822_,
		_w26774_
	);
	LUT4 #(
		.INIT('h9dbf)
	) name24874 (
		_w8816_,
		_w8819_,
		_w26773_,
		_w26774_,
		_w26775_
	);
	LUT3 #(
		.INIT('h80)
	) name24875 (
		\m6_data_i[10]_pad ,
		_w8821_,
		_w8822_,
		_w26776_
	);
	LUT3 #(
		.INIT('h2a)
	) name24876 (
		\m7_data_i[10]_pad ,
		_w8821_,
		_w8822_,
		_w26777_
	);
	LUT3 #(
		.INIT('h57)
	) name24877 (
		_w8834_,
		_w26776_,
		_w26777_,
		_w26778_
	);
	LUT3 #(
		.INIT('h2a)
	) name24878 (
		\m5_data_i[10]_pad ,
		_w8821_,
		_w8822_,
		_w26779_
	);
	LUT3 #(
		.INIT('h80)
	) name24879 (
		\m0_data_i[10]_pad ,
		_w8821_,
		_w8822_,
		_w26780_
	);
	LUT4 #(
		.INIT('h57df)
	) name24880 (
		_w8816_,
		_w8819_,
		_w26779_,
		_w26780_,
		_w26781_
	);
	LUT3 #(
		.INIT('h2a)
	) name24881 (
		\m1_data_i[10]_pad ,
		_w8821_,
		_w8822_,
		_w26782_
	);
	LUT3 #(
		.INIT('h80)
	) name24882 (
		\m2_data_i[10]_pad ,
		_w8821_,
		_w8822_,
		_w26783_
	);
	LUT4 #(
		.INIT('h3b7f)
	) name24883 (
		_w8816_,
		_w8819_,
		_w26782_,
		_w26783_,
		_w26784_
	);
	LUT4 #(
		.INIT('h7fff)
	) name24884 (
		_w26775_,
		_w26778_,
		_w26781_,
		_w26784_,
		_w26785_
	);
	LUT3 #(
		.INIT('h2a)
	) name24885 (
		\m3_data_i[11]_pad ,
		_w8821_,
		_w8822_,
		_w26786_
	);
	LUT3 #(
		.INIT('h80)
	) name24886 (
		\m4_data_i[11]_pad ,
		_w8821_,
		_w8822_,
		_w26787_
	);
	LUT4 #(
		.INIT('h9dbf)
	) name24887 (
		_w8816_,
		_w8819_,
		_w26786_,
		_w26787_,
		_w26788_
	);
	LUT3 #(
		.INIT('h80)
	) name24888 (
		\m6_data_i[11]_pad ,
		_w8821_,
		_w8822_,
		_w26789_
	);
	LUT3 #(
		.INIT('h2a)
	) name24889 (
		\m7_data_i[11]_pad ,
		_w8821_,
		_w8822_,
		_w26790_
	);
	LUT3 #(
		.INIT('h57)
	) name24890 (
		_w8834_,
		_w26789_,
		_w26790_,
		_w26791_
	);
	LUT3 #(
		.INIT('h2a)
	) name24891 (
		\m5_data_i[11]_pad ,
		_w8821_,
		_w8822_,
		_w26792_
	);
	LUT3 #(
		.INIT('h80)
	) name24892 (
		\m0_data_i[11]_pad ,
		_w8821_,
		_w8822_,
		_w26793_
	);
	LUT4 #(
		.INIT('h57df)
	) name24893 (
		_w8816_,
		_w8819_,
		_w26792_,
		_w26793_,
		_w26794_
	);
	LUT3 #(
		.INIT('h2a)
	) name24894 (
		\m1_data_i[11]_pad ,
		_w8821_,
		_w8822_,
		_w26795_
	);
	LUT3 #(
		.INIT('h80)
	) name24895 (
		\m2_data_i[11]_pad ,
		_w8821_,
		_w8822_,
		_w26796_
	);
	LUT4 #(
		.INIT('h3b7f)
	) name24896 (
		_w8816_,
		_w8819_,
		_w26795_,
		_w26796_,
		_w26797_
	);
	LUT4 #(
		.INIT('h7fff)
	) name24897 (
		_w26788_,
		_w26791_,
		_w26794_,
		_w26797_,
		_w26798_
	);
	LUT3 #(
		.INIT('h2a)
	) name24898 (
		\m3_data_i[12]_pad ,
		_w8821_,
		_w8822_,
		_w26799_
	);
	LUT3 #(
		.INIT('h80)
	) name24899 (
		\m4_data_i[12]_pad ,
		_w8821_,
		_w8822_,
		_w26800_
	);
	LUT4 #(
		.INIT('h9dbf)
	) name24900 (
		_w8816_,
		_w8819_,
		_w26799_,
		_w26800_,
		_w26801_
	);
	LUT3 #(
		.INIT('h80)
	) name24901 (
		\m6_data_i[12]_pad ,
		_w8821_,
		_w8822_,
		_w26802_
	);
	LUT3 #(
		.INIT('h2a)
	) name24902 (
		\m7_data_i[12]_pad ,
		_w8821_,
		_w8822_,
		_w26803_
	);
	LUT3 #(
		.INIT('h57)
	) name24903 (
		_w8834_,
		_w26802_,
		_w26803_,
		_w26804_
	);
	LUT3 #(
		.INIT('h2a)
	) name24904 (
		\m5_data_i[12]_pad ,
		_w8821_,
		_w8822_,
		_w26805_
	);
	LUT3 #(
		.INIT('h80)
	) name24905 (
		\m0_data_i[12]_pad ,
		_w8821_,
		_w8822_,
		_w26806_
	);
	LUT4 #(
		.INIT('h57df)
	) name24906 (
		_w8816_,
		_w8819_,
		_w26805_,
		_w26806_,
		_w26807_
	);
	LUT3 #(
		.INIT('h2a)
	) name24907 (
		\m1_data_i[12]_pad ,
		_w8821_,
		_w8822_,
		_w26808_
	);
	LUT3 #(
		.INIT('h80)
	) name24908 (
		\m2_data_i[12]_pad ,
		_w8821_,
		_w8822_,
		_w26809_
	);
	LUT4 #(
		.INIT('h3b7f)
	) name24909 (
		_w8816_,
		_w8819_,
		_w26808_,
		_w26809_,
		_w26810_
	);
	LUT4 #(
		.INIT('h7fff)
	) name24910 (
		_w26801_,
		_w26804_,
		_w26807_,
		_w26810_,
		_w26811_
	);
	LUT3 #(
		.INIT('h2a)
	) name24911 (
		\m3_data_i[13]_pad ,
		_w8821_,
		_w8822_,
		_w26812_
	);
	LUT3 #(
		.INIT('h80)
	) name24912 (
		\m4_data_i[13]_pad ,
		_w8821_,
		_w8822_,
		_w26813_
	);
	LUT4 #(
		.INIT('h9dbf)
	) name24913 (
		_w8816_,
		_w8819_,
		_w26812_,
		_w26813_,
		_w26814_
	);
	LUT3 #(
		.INIT('h80)
	) name24914 (
		\m6_data_i[13]_pad ,
		_w8821_,
		_w8822_,
		_w26815_
	);
	LUT3 #(
		.INIT('h80)
	) name24915 (
		\m2_data_i[13]_pad ,
		_w8821_,
		_w8822_,
		_w26816_
	);
	LUT4 #(
		.INIT('habef)
	) name24916 (
		_w8816_,
		_w8819_,
		_w26815_,
		_w26816_,
		_w26817_
	);
	LUT3 #(
		.INIT('h2a)
	) name24917 (
		\m5_data_i[13]_pad ,
		_w8821_,
		_w8822_,
		_w26818_
	);
	LUT3 #(
		.INIT('h2a)
	) name24918 (
		\m1_data_i[13]_pad ,
		_w8821_,
		_w8822_,
		_w26819_
	);
	LUT4 #(
		.INIT('h57df)
	) name24919 (
		_w8816_,
		_w8819_,
		_w26818_,
		_w26819_,
		_w26820_
	);
	LUT3 #(
		.INIT('h80)
	) name24920 (
		\m0_data_i[13]_pad ,
		_w8821_,
		_w8822_,
		_w26821_
	);
	LUT3 #(
		.INIT('h2a)
	) name24921 (
		\m7_data_i[13]_pad ,
		_w8821_,
		_w8822_,
		_w26822_
	);
	LUT4 #(
		.INIT('h6e7f)
	) name24922 (
		_w8816_,
		_w8819_,
		_w26821_,
		_w26822_,
		_w26823_
	);
	LUT4 #(
		.INIT('h7fff)
	) name24923 (
		_w26814_,
		_w26817_,
		_w26820_,
		_w26823_,
		_w26824_
	);
	LUT3 #(
		.INIT('h2a)
	) name24924 (
		\m1_data_i[14]_pad ,
		_w8821_,
		_w8822_,
		_w26825_
	);
	LUT3 #(
		.INIT('h80)
	) name24925 (
		\m2_data_i[14]_pad ,
		_w8821_,
		_w8822_,
		_w26826_
	);
	LUT4 #(
		.INIT('h3b7f)
	) name24926 (
		_w8816_,
		_w8819_,
		_w26825_,
		_w26826_,
		_w26827_
	);
	LUT3 #(
		.INIT('h80)
	) name24927 (
		\m6_data_i[14]_pad ,
		_w8821_,
		_w8822_,
		_w26828_
	);
	LUT3 #(
		.INIT('h2a)
	) name24928 (
		\m7_data_i[14]_pad ,
		_w8821_,
		_w8822_,
		_w26829_
	);
	LUT3 #(
		.INIT('h57)
	) name24929 (
		_w8834_,
		_w26828_,
		_w26829_,
		_w26830_
	);
	LUT3 #(
		.INIT('h2a)
	) name24930 (
		\m5_data_i[14]_pad ,
		_w8821_,
		_w8822_,
		_w26831_
	);
	LUT3 #(
		.INIT('h80)
	) name24931 (
		\m0_data_i[14]_pad ,
		_w8821_,
		_w8822_,
		_w26832_
	);
	LUT4 #(
		.INIT('h57df)
	) name24932 (
		_w8816_,
		_w8819_,
		_w26831_,
		_w26832_,
		_w26833_
	);
	LUT3 #(
		.INIT('h2a)
	) name24933 (
		\m3_data_i[14]_pad ,
		_w8821_,
		_w8822_,
		_w26834_
	);
	LUT3 #(
		.INIT('h80)
	) name24934 (
		\m4_data_i[14]_pad ,
		_w8821_,
		_w8822_,
		_w26835_
	);
	LUT4 #(
		.INIT('h9dbf)
	) name24935 (
		_w8816_,
		_w8819_,
		_w26834_,
		_w26835_,
		_w26836_
	);
	LUT4 #(
		.INIT('h7fff)
	) name24936 (
		_w26827_,
		_w26830_,
		_w26833_,
		_w26836_,
		_w26837_
	);
	LUT3 #(
		.INIT('h2a)
	) name24937 (
		\m3_data_i[15]_pad ,
		_w8821_,
		_w8822_,
		_w26838_
	);
	LUT3 #(
		.INIT('h80)
	) name24938 (
		\m4_data_i[15]_pad ,
		_w8821_,
		_w8822_,
		_w26839_
	);
	LUT4 #(
		.INIT('h9dbf)
	) name24939 (
		_w8816_,
		_w8819_,
		_w26838_,
		_w26839_,
		_w26840_
	);
	LUT3 #(
		.INIT('h80)
	) name24940 (
		\m6_data_i[15]_pad ,
		_w8821_,
		_w8822_,
		_w26841_
	);
	LUT3 #(
		.INIT('h80)
	) name24941 (
		\m2_data_i[15]_pad ,
		_w8821_,
		_w8822_,
		_w26842_
	);
	LUT4 #(
		.INIT('habef)
	) name24942 (
		_w8816_,
		_w8819_,
		_w26841_,
		_w26842_,
		_w26843_
	);
	LUT3 #(
		.INIT('h2a)
	) name24943 (
		\m5_data_i[15]_pad ,
		_w8821_,
		_w8822_,
		_w26844_
	);
	LUT3 #(
		.INIT('h2a)
	) name24944 (
		\m1_data_i[15]_pad ,
		_w8821_,
		_w8822_,
		_w26845_
	);
	LUT4 #(
		.INIT('h57df)
	) name24945 (
		_w8816_,
		_w8819_,
		_w26844_,
		_w26845_,
		_w26846_
	);
	LUT3 #(
		.INIT('h80)
	) name24946 (
		\m0_data_i[15]_pad ,
		_w8821_,
		_w8822_,
		_w26847_
	);
	LUT3 #(
		.INIT('h2a)
	) name24947 (
		\m7_data_i[15]_pad ,
		_w8821_,
		_w8822_,
		_w26848_
	);
	LUT4 #(
		.INIT('h6e7f)
	) name24948 (
		_w8816_,
		_w8819_,
		_w26847_,
		_w26848_,
		_w26849_
	);
	LUT4 #(
		.INIT('h7fff)
	) name24949 (
		_w26840_,
		_w26843_,
		_w26846_,
		_w26849_,
		_w26850_
	);
	LUT3 #(
		.INIT('h2a)
	) name24950 (
		\m3_data_i[16]_pad ,
		_w8821_,
		_w8822_,
		_w26851_
	);
	LUT3 #(
		.INIT('h80)
	) name24951 (
		\m4_data_i[16]_pad ,
		_w8821_,
		_w8822_,
		_w26852_
	);
	LUT4 #(
		.INIT('h9dbf)
	) name24952 (
		_w8816_,
		_w8819_,
		_w26851_,
		_w26852_,
		_w26853_
	);
	LUT3 #(
		.INIT('h80)
	) name24953 (
		\m6_data_i[16]_pad ,
		_w8821_,
		_w8822_,
		_w26854_
	);
	LUT3 #(
		.INIT('h80)
	) name24954 (
		\m2_data_i[16]_pad ,
		_w8821_,
		_w8822_,
		_w26855_
	);
	LUT4 #(
		.INIT('habef)
	) name24955 (
		_w8816_,
		_w8819_,
		_w26854_,
		_w26855_,
		_w26856_
	);
	LUT3 #(
		.INIT('h2a)
	) name24956 (
		\m5_data_i[16]_pad ,
		_w8821_,
		_w8822_,
		_w26857_
	);
	LUT3 #(
		.INIT('h2a)
	) name24957 (
		\m1_data_i[16]_pad ,
		_w8821_,
		_w8822_,
		_w26858_
	);
	LUT4 #(
		.INIT('h57df)
	) name24958 (
		_w8816_,
		_w8819_,
		_w26857_,
		_w26858_,
		_w26859_
	);
	LUT3 #(
		.INIT('h80)
	) name24959 (
		\m0_data_i[16]_pad ,
		_w8821_,
		_w8822_,
		_w26860_
	);
	LUT3 #(
		.INIT('h2a)
	) name24960 (
		\m7_data_i[16]_pad ,
		_w8821_,
		_w8822_,
		_w26861_
	);
	LUT4 #(
		.INIT('h6e7f)
	) name24961 (
		_w8816_,
		_w8819_,
		_w26860_,
		_w26861_,
		_w26862_
	);
	LUT4 #(
		.INIT('h7fff)
	) name24962 (
		_w26853_,
		_w26856_,
		_w26859_,
		_w26862_,
		_w26863_
	);
	LUT3 #(
		.INIT('h2a)
	) name24963 (
		\m3_data_i[17]_pad ,
		_w8821_,
		_w8822_,
		_w26864_
	);
	LUT3 #(
		.INIT('h80)
	) name24964 (
		\m4_data_i[17]_pad ,
		_w8821_,
		_w8822_,
		_w26865_
	);
	LUT4 #(
		.INIT('h9dbf)
	) name24965 (
		_w8816_,
		_w8819_,
		_w26864_,
		_w26865_,
		_w26866_
	);
	LUT3 #(
		.INIT('h80)
	) name24966 (
		\m6_data_i[17]_pad ,
		_w8821_,
		_w8822_,
		_w26867_
	);
	LUT3 #(
		.INIT('h2a)
	) name24967 (
		\m7_data_i[17]_pad ,
		_w8821_,
		_w8822_,
		_w26868_
	);
	LUT3 #(
		.INIT('h57)
	) name24968 (
		_w8834_,
		_w26867_,
		_w26868_,
		_w26869_
	);
	LUT3 #(
		.INIT('h2a)
	) name24969 (
		\m5_data_i[17]_pad ,
		_w8821_,
		_w8822_,
		_w26870_
	);
	LUT3 #(
		.INIT('h80)
	) name24970 (
		\m0_data_i[17]_pad ,
		_w8821_,
		_w8822_,
		_w26871_
	);
	LUT4 #(
		.INIT('h57df)
	) name24971 (
		_w8816_,
		_w8819_,
		_w26870_,
		_w26871_,
		_w26872_
	);
	LUT3 #(
		.INIT('h2a)
	) name24972 (
		\m1_data_i[17]_pad ,
		_w8821_,
		_w8822_,
		_w26873_
	);
	LUT3 #(
		.INIT('h80)
	) name24973 (
		\m2_data_i[17]_pad ,
		_w8821_,
		_w8822_,
		_w26874_
	);
	LUT4 #(
		.INIT('h3b7f)
	) name24974 (
		_w8816_,
		_w8819_,
		_w26873_,
		_w26874_,
		_w26875_
	);
	LUT4 #(
		.INIT('h7fff)
	) name24975 (
		_w26866_,
		_w26869_,
		_w26872_,
		_w26875_,
		_w26876_
	);
	LUT3 #(
		.INIT('h2a)
	) name24976 (
		\m1_data_i[18]_pad ,
		_w8821_,
		_w8822_,
		_w26877_
	);
	LUT3 #(
		.INIT('h80)
	) name24977 (
		\m2_data_i[18]_pad ,
		_w8821_,
		_w8822_,
		_w26878_
	);
	LUT4 #(
		.INIT('h3b7f)
	) name24978 (
		_w8816_,
		_w8819_,
		_w26877_,
		_w26878_,
		_w26879_
	);
	LUT3 #(
		.INIT('h2a)
	) name24979 (
		\m3_data_i[18]_pad ,
		_w8821_,
		_w8822_,
		_w26880_
	);
	LUT3 #(
		.INIT('h2a)
	) name24980 (
		\m7_data_i[18]_pad ,
		_w8821_,
		_w8822_,
		_w26881_
	);
	LUT4 #(
		.INIT('haebf)
	) name24981 (
		_w8816_,
		_w8819_,
		_w26880_,
		_w26881_,
		_w26882_
	);
	LUT3 #(
		.INIT('h80)
	) name24982 (
		\m4_data_i[18]_pad ,
		_w8821_,
		_w8822_,
		_w26883_
	);
	LUT3 #(
		.INIT('h80)
	) name24983 (
		\m0_data_i[18]_pad ,
		_w8821_,
		_w8822_,
		_w26884_
	);
	LUT4 #(
		.INIT('h57df)
	) name24984 (
		_w8816_,
		_w8819_,
		_w26883_,
		_w26884_,
		_w26885_
	);
	LUT3 #(
		.INIT('h80)
	) name24985 (
		\m6_data_i[18]_pad ,
		_w8821_,
		_w8822_,
		_w26886_
	);
	LUT3 #(
		.INIT('h2a)
	) name24986 (
		\m5_data_i[18]_pad ,
		_w8821_,
		_w8822_,
		_w26887_
	);
	LUT4 #(
		.INIT('hcdef)
	) name24987 (
		_w8816_,
		_w8819_,
		_w26886_,
		_w26887_,
		_w26888_
	);
	LUT4 #(
		.INIT('h7fff)
	) name24988 (
		_w26879_,
		_w26882_,
		_w26885_,
		_w26888_,
		_w26889_
	);
	LUT3 #(
		.INIT('h2a)
	) name24989 (
		\m1_data_i[19]_pad ,
		_w8821_,
		_w8822_,
		_w26890_
	);
	LUT3 #(
		.INIT('h80)
	) name24990 (
		\m2_data_i[19]_pad ,
		_w8821_,
		_w8822_,
		_w26891_
	);
	LUT4 #(
		.INIT('h3b7f)
	) name24991 (
		_w8816_,
		_w8819_,
		_w26890_,
		_w26891_,
		_w26892_
	);
	LUT3 #(
		.INIT('h80)
	) name24992 (
		\m6_data_i[19]_pad ,
		_w8821_,
		_w8822_,
		_w26893_
	);
	LUT3 #(
		.INIT('h2a)
	) name24993 (
		\m7_data_i[19]_pad ,
		_w8821_,
		_w8822_,
		_w26894_
	);
	LUT3 #(
		.INIT('h57)
	) name24994 (
		_w8834_,
		_w26893_,
		_w26894_,
		_w26895_
	);
	LUT3 #(
		.INIT('h2a)
	) name24995 (
		\m5_data_i[19]_pad ,
		_w8821_,
		_w8822_,
		_w26896_
	);
	LUT3 #(
		.INIT('h80)
	) name24996 (
		\m0_data_i[19]_pad ,
		_w8821_,
		_w8822_,
		_w26897_
	);
	LUT4 #(
		.INIT('h57df)
	) name24997 (
		_w8816_,
		_w8819_,
		_w26896_,
		_w26897_,
		_w26898_
	);
	LUT3 #(
		.INIT('h2a)
	) name24998 (
		\m3_data_i[19]_pad ,
		_w8821_,
		_w8822_,
		_w26899_
	);
	LUT3 #(
		.INIT('h80)
	) name24999 (
		\m4_data_i[19]_pad ,
		_w8821_,
		_w8822_,
		_w26900_
	);
	LUT4 #(
		.INIT('h9dbf)
	) name25000 (
		_w8816_,
		_w8819_,
		_w26899_,
		_w26900_,
		_w26901_
	);
	LUT4 #(
		.INIT('h7fff)
	) name25001 (
		_w26892_,
		_w26895_,
		_w26898_,
		_w26901_,
		_w26902_
	);
	LUT3 #(
		.INIT('h80)
	) name25002 (
		\m0_data_i[1]_pad ,
		_w8821_,
		_w8822_,
		_w26903_
	);
	LUT3 #(
		.INIT('h2a)
	) name25003 (
		\m7_data_i[1]_pad ,
		_w8821_,
		_w8822_,
		_w26904_
	);
	LUT4 #(
		.INIT('h6e7f)
	) name25004 (
		_w8816_,
		_w8819_,
		_w26903_,
		_w26904_,
		_w26905_
	);
	LUT3 #(
		.INIT('h2a)
	) name25005 (
		\m3_data_i[1]_pad ,
		_w8821_,
		_w8822_,
		_w26906_
	);
	LUT3 #(
		.INIT('h80)
	) name25006 (
		\m2_data_i[1]_pad ,
		_w8821_,
		_w8822_,
		_w26907_
	);
	LUT3 #(
		.INIT('h57)
	) name25007 (
		_w8828_,
		_w26906_,
		_w26907_,
		_w26908_
	);
	LUT3 #(
		.INIT('h80)
	) name25008 (
		\m4_data_i[1]_pad ,
		_w8821_,
		_w8822_,
		_w26909_
	);
	LUT3 #(
		.INIT('h2a)
	) name25009 (
		\m1_data_i[1]_pad ,
		_w8821_,
		_w8822_,
		_w26910_
	);
	LUT4 #(
		.INIT('h57df)
	) name25010 (
		_w8816_,
		_w8819_,
		_w26909_,
		_w26910_,
		_w26911_
	);
	LUT3 #(
		.INIT('h80)
	) name25011 (
		\m6_data_i[1]_pad ,
		_w8821_,
		_w8822_,
		_w26912_
	);
	LUT3 #(
		.INIT('h2a)
	) name25012 (
		\m5_data_i[1]_pad ,
		_w8821_,
		_w8822_,
		_w26913_
	);
	LUT4 #(
		.INIT('hcdef)
	) name25013 (
		_w8816_,
		_w8819_,
		_w26912_,
		_w26913_,
		_w26914_
	);
	LUT4 #(
		.INIT('h7fff)
	) name25014 (
		_w26905_,
		_w26908_,
		_w26911_,
		_w26914_,
		_w26915_
	);
	LUT3 #(
		.INIT('h80)
	) name25015 (
		\m0_data_i[20]_pad ,
		_w8821_,
		_w8822_,
		_w26916_
	);
	LUT3 #(
		.INIT('h2a)
	) name25016 (
		\m7_data_i[20]_pad ,
		_w8821_,
		_w8822_,
		_w26917_
	);
	LUT4 #(
		.INIT('h6e7f)
	) name25017 (
		_w8816_,
		_w8819_,
		_w26916_,
		_w26917_,
		_w26918_
	);
	LUT3 #(
		.INIT('h2a)
	) name25018 (
		\m3_data_i[20]_pad ,
		_w8821_,
		_w8822_,
		_w26919_
	);
	LUT3 #(
		.INIT('h80)
	) name25019 (
		\m2_data_i[20]_pad ,
		_w8821_,
		_w8822_,
		_w26920_
	);
	LUT3 #(
		.INIT('h57)
	) name25020 (
		_w8828_,
		_w26919_,
		_w26920_,
		_w26921_
	);
	LUT3 #(
		.INIT('h80)
	) name25021 (
		\m4_data_i[20]_pad ,
		_w8821_,
		_w8822_,
		_w26922_
	);
	LUT3 #(
		.INIT('h2a)
	) name25022 (
		\m1_data_i[20]_pad ,
		_w8821_,
		_w8822_,
		_w26923_
	);
	LUT4 #(
		.INIT('h57df)
	) name25023 (
		_w8816_,
		_w8819_,
		_w26922_,
		_w26923_,
		_w26924_
	);
	LUT3 #(
		.INIT('h80)
	) name25024 (
		\m6_data_i[20]_pad ,
		_w8821_,
		_w8822_,
		_w26925_
	);
	LUT3 #(
		.INIT('h2a)
	) name25025 (
		\m5_data_i[20]_pad ,
		_w8821_,
		_w8822_,
		_w26926_
	);
	LUT4 #(
		.INIT('hcdef)
	) name25026 (
		_w8816_,
		_w8819_,
		_w26925_,
		_w26926_,
		_w26927_
	);
	LUT4 #(
		.INIT('h7fff)
	) name25027 (
		_w26918_,
		_w26921_,
		_w26924_,
		_w26927_,
		_w26928_
	);
	LUT3 #(
		.INIT('h2a)
	) name25028 (
		\m1_data_i[21]_pad ,
		_w8821_,
		_w8822_,
		_w26929_
	);
	LUT3 #(
		.INIT('h80)
	) name25029 (
		\m2_data_i[21]_pad ,
		_w8821_,
		_w8822_,
		_w26930_
	);
	LUT4 #(
		.INIT('h3b7f)
	) name25030 (
		_w8816_,
		_w8819_,
		_w26929_,
		_w26930_,
		_w26931_
	);
	LUT3 #(
		.INIT('h2a)
	) name25031 (
		\m3_data_i[21]_pad ,
		_w8821_,
		_w8822_,
		_w26932_
	);
	LUT3 #(
		.INIT('h2a)
	) name25032 (
		\m7_data_i[21]_pad ,
		_w8821_,
		_w8822_,
		_w26933_
	);
	LUT4 #(
		.INIT('haebf)
	) name25033 (
		_w8816_,
		_w8819_,
		_w26932_,
		_w26933_,
		_w26934_
	);
	LUT3 #(
		.INIT('h80)
	) name25034 (
		\m4_data_i[21]_pad ,
		_w8821_,
		_w8822_,
		_w26935_
	);
	LUT3 #(
		.INIT('h80)
	) name25035 (
		\m0_data_i[21]_pad ,
		_w8821_,
		_w8822_,
		_w26936_
	);
	LUT4 #(
		.INIT('h57df)
	) name25036 (
		_w8816_,
		_w8819_,
		_w26935_,
		_w26936_,
		_w26937_
	);
	LUT3 #(
		.INIT('h80)
	) name25037 (
		\m6_data_i[21]_pad ,
		_w8821_,
		_w8822_,
		_w26938_
	);
	LUT3 #(
		.INIT('h2a)
	) name25038 (
		\m5_data_i[21]_pad ,
		_w8821_,
		_w8822_,
		_w26939_
	);
	LUT4 #(
		.INIT('hcdef)
	) name25039 (
		_w8816_,
		_w8819_,
		_w26938_,
		_w26939_,
		_w26940_
	);
	LUT4 #(
		.INIT('h7fff)
	) name25040 (
		_w26931_,
		_w26934_,
		_w26937_,
		_w26940_,
		_w26941_
	);
	LUT3 #(
		.INIT('h2a)
	) name25041 (
		\m1_data_i[22]_pad ,
		_w8821_,
		_w8822_,
		_w26942_
	);
	LUT3 #(
		.INIT('h80)
	) name25042 (
		\m2_data_i[22]_pad ,
		_w8821_,
		_w8822_,
		_w26943_
	);
	LUT4 #(
		.INIT('h3b7f)
	) name25043 (
		_w8816_,
		_w8819_,
		_w26942_,
		_w26943_,
		_w26944_
	);
	LUT3 #(
		.INIT('h80)
	) name25044 (
		\m6_data_i[22]_pad ,
		_w8821_,
		_w8822_,
		_w26945_
	);
	LUT3 #(
		.INIT('h2a)
	) name25045 (
		\m7_data_i[22]_pad ,
		_w8821_,
		_w8822_,
		_w26946_
	);
	LUT3 #(
		.INIT('h57)
	) name25046 (
		_w8834_,
		_w26945_,
		_w26946_,
		_w26947_
	);
	LUT3 #(
		.INIT('h2a)
	) name25047 (
		\m5_data_i[22]_pad ,
		_w8821_,
		_w8822_,
		_w26948_
	);
	LUT3 #(
		.INIT('h80)
	) name25048 (
		\m0_data_i[22]_pad ,
		_w8821_,
		_w8822_,
		_w26949_
	);
	LUT4 #(
		.INIT('h57df)
	) name25049 (
		_w8816_,
		_w8819_,
		_w26948_,
		_w26949_,
		_w26950_
	);
	LUT3 #(
		.INIT('h2a)
	) name25050 (
		\m3_data_i[22]_pad ,
		_w8821_,
		_w8822_,
		_w26951_
	);
	LUT3 #(
		.INIT('h80)
	) name25051 (
		\m4_data_i[22]_pad ,
		_w8821_,
		_w8822_,
		_w26952_
	);
	LUT4 #(
		.INIT('h9dbf)
	) name25052 (
		_w8816_,
		_w8819_,
		_w26951_,
		_w26952_,
		_w26953_
	);
	LUT4 #(
		.INIT('h7fff)
	) name25053 (
		_w26944_,
		_w26947_,
		_w26950_,
		_w26953_,
		_w26954_
	);
	LUT3 #(
		.INIT('h2a)
	) name25054 (
		\m3_data_i[23]_pad ,
		_w8821_,
		_w8822_,
		_w26955_
	);
	LUT3 #(
		.INIT('h80)
	) name25055 (
		\m4_data_i[23]_pad ,
		_w8821_,
		_w8822_,
		_w26956_
	);
	LUT4 #(
		.INIT('h9dbf)
	) name25056 (
		_w8816_,
		_w8819_,
		_w26955_,
		_w26956_,
		_w26957_
	);
	LUT3 #(
		.INIT('h80)
	) name25057 (
		\m6_data_i[23]_pad ,
		_w8821_,
		_w8822_,
		_w26958_
	);
	LUT3 #(
		.INIT('h80)
	) name25058 (
		\m2_data_i[23]_pad ,
		_w8821_,
		_w8822_,
		_w26959_
	);
	LUT4 #(
		.INIT('habef)
	) name25059 (
		_w8816_,
		_w8819_,
		_w26958_,
		_w26959_,
		_w26960_
	);
	LUT3 #(
		.INIT('h2a)
	) name25060 (
		\m5_data_i[23]_pad ,
		_w8821_,
		_w8822_,
		_w26961_
	);
	LUT3 #(
		.INIT('h2a)
	) name25061 (
		\m1_data_i[23]_pad ,
		_w8821_,
		_w8822_,
		_w26962_
	);
	LUT4 #(
		.INIT('h57df)
	) name25062 (
		_w8816_,
		_w8819_,
		_w26961_,
		_w26962_,
		_w26963_
	);
	LUT3 #(
		.INIT('h80)
	) name25063 (
		\m0_data_i[23]_pad ,
		_w8821_,
		_w8822_,
		_w26964_
	);
	LUT3 #(
		.INIT('h2a)
	) name25064 (
		\m7_data_i[23]_pad ,
		_w8821_,
		_w8822_,
		_w26965_
	);
	LUT4 #(
		.INIT('h6e7f)
	) name25065 (
		_w8816_,
		_w8819_,
		_w26964_,
		_w26965_,
		_w26966_
	);
	LUT4 #(
		.INIT('h7fff)
	) name25066 (
		_w26957_,
		_w26960_,
		_w26963_,
		_w26966_,
		_w26967_
	);
	LUT3 #(
		.INIT('h2a)
	) name25067 (
		\m1_data_i[24]_pad ,
		_w8821_,
		_w8822_,
		_w26968_
	);
	LUT3 #(
		.INIT('h80)
	) name25068 (
		\m2_data_i[24]_pad ,
		_w8821_,
		_w8822_,
		_w26969_
	);
	LUT4 #(
		.INIT('h3b7f)
	) name25069 (
		_w8816_,
		_w8819_,
		_w26968_,
		_w26969_,
		_w26970_
	);
	LUT3 #(
		.INIT('h2a)
	) name25070 (
		\m3_data_i[24]_pad ,
		_w8821_,
		_w8822_,
		_w26971_
	);
	LUT3 #(
		.INIT('h2a)
	) name25071 (
		\m7_data_i[24]_pad ,
		_w8821_,
		_w8822_,
		_w26972_
	);
	LUT4 #(
		.INIT('haebf)
	) name25072 (
		_w8816_,
		_w8819_,
		_w26971_,
		_w26972_,
		_w26973_
	);
	LUT3 #(
		.INIT('h80)
	) name25073 (
		\m4_data_i[24]_pad ,
		_w8821_,
		_w8822_,
		_w26974_
	);
	LUT3 #(
		.INIT('h80)
	) name25074 (
		\m0_data_i[24]_pad ,
		_w8821_,
		_w8822_,
		_w26975_
	);
	LUT4 #(
		.INIT('h57df)
	) name25075 (
		_w8816_,
		_w8819_,
		_w26974_,
		_w26975_,
		_w26976_
	);
	LUT3 #(
		.INIT('h80)
	) name25076 (
		\m6_data_i[24]_pad ,
		_w8821_,
		_w8822_,
		_w26977_
	);
	LUT3 #(
		.INIT('h2a)
	) name25077 (
		\m5_data_i[24]_pad ,
		_w8821_,
		_w8822_,
		_w26978_
	);
	LUT4 #(
		.INIT('hcdef)
	) name25078 (
		_w8816_,
		_w8819_,
		_w26977_,
		_w26978_,
		_w26979_
	);
	LUT4 #(
		.INIT('h7fff)
	) name25079 (
		_w26970_,
		_w26973_,
		_w26976_,
		_w26979_,
		_w26980_
	);
	LUT3 #(
		.INIT('h2a)
	) name25080 (
		\m3_data_i[25]_pad ,
		_w8821_,
		_w8822_,
		_w26981_
	);
	LUT3 #(
		.INIT('h80)
	) name25081 (
		\m4_data_i[25]_pad ,
		_w8821_,
		_w8822_,
		_w26982_
	);
	LUT4 #(
		.INIT('h9dbf)
	) name25082 (
		_w8816_,
		_w8819_,
		_w26981_,
		_w26982_,
		_w26983_
	);
	LUT3 #(
		.INIT('h80)
	) name25083 (
		\m6_data_i[25]_pad ,
		_w8821_,
		_w8822_,
		_w26984_
	);
	LUT3 #(
		.INIT('h2a)
	) name25084 (
		\m7_data_i[25]_pad ,
		_w8821_,
		_w8822_,
		_w26985_
	);
	LUT3 #(
		.INIT('h57)
	) name25085 (
		_w8834_,
		_w26984_,
		_w26985_,
		_w26986_
	);
	LUT3 #(
		.INIT('h2a)
	) name25086 (
		\m5_data_i[25]_pad ,
		_w8821_,
		_w8822_,
		_w26987_
	);
	LUT3 #(
		.INIT('h80)
	) name25087 (
		\m0_data_i[25]_pad ,
		_w8821_,
		_w8822_,
		_w26988_
	);
	LUT4 #(
		.INIT('h57df)
	) name25088 (
		_w8816_,
		_w8819_,
		_w26987_,
		_w26988_,
		_w26989_
	);
	LUT3 #(
		.INIT('h2a)
	) name25089 (
		\m1_data_i[25]_pad ,
		_w8821_,
		_w8822_,
		_w26990_
	);
	LUT3 #(
		.INIT('h80)
	) name25090 (
		\m2_data_i[25]_pad ,
		_w8821_,
		_w8822_,
		_w26991_
	);
	LUT4 #(
		.INIT('h3b7f)
	) name25091 (
		_w8816_,
		_w8819_,
		_w26990_,
		_w26991_,
		_w26992_
	);
	LUT4 #(
		.INIT('h7fff)
	) name25092 (
		_w26983_,
		_w26986_,
		_w26989_,
		_w26992_,
		_w26993_
	);
	LUT3 #(
		.INIT('h80)
	) name25093 (
		\m0_data_i[26]_pad ,
		_w8821_,
		_w8822_,
		_w26994_
	);
	LUT3 #(
		.INIT('h2a)
	) name25094 (
		\m7_data_i[26]_pad ,
		_w8821_,
		_w8822_,
		_w26995_
	);
	LUT4 #(
		.INIT('h6e7f)
	) name25095 (
		_w8816_,
		_w8819_,
		_w26994_,
		_w26995_,
		_w26996_
	);
	LUT3 #(
		.INIT('h2a)
	) name25096 (
		\m3_data_i[26]_pad ,
		_w8821_,
		_w8822_,
		_w26997_
	);
	LUT3 #(
		.INIT('h80)
	) name25097 (
		\m2_data_i[26]_pad ,
		_w8821_,
		_w8822_,
		_w26998_
	);
	LUT3 #(
		.INIT('h57)
	) name25098 (
		_w8828_,
		_w26997_,
		_w26998_,
		_w26999_
	);
	LUT3 #(
		.INIT('h80)
	) name25099 (
		\m4_data_i[26]_pad ,
		_w8821_,
		_w8822_,
		_w27000_
	);
	LUT3 #(
		.INIT('h2a)
	) name25100 (
		\m1_data_i[26]_pad ,
		_w8821_,
		_w8822_,
		_w27001_
	);
	LUT4 #(
		.INIT('h57df)
	) name25101 (
		_w8816_,
		_w8819_,
		_w27000_,
		_w27001_,
		_w27002_
	);
	LUT3 #(
		.INIT('h80)
	) name25102 (
		\m6_data_i[26]_pad ,
		_w8821_,
		_w8822_,
		_w27003_
	);
	LUT3 #(
		.INIT('h2a)
	) name25103 (
		\m5_data_i[26]_pad ,
		_w8821_,
		_w8822_,
		_w27004_
	);
	LUT4 #(
		.INIT('hcdef)
	) name25104 (
		_w8816_,
		_w8819_,
		_w27003_,
		_w27004_,
		_w27005_
	);
	LUT4 #(
		.INIT('h7fff)
	) name25105 (
		_w26996_,
		_w26999_,
		_w27002_,
		_w27005_,
		_w27006_
	);
	LUT3 #(
		.INIT('h2a)
	) name25106 (
		\m3_data_i[27]_pad ,
		_w8821_,
		_w8822_,
		_w27007_
	);
	LUT3 #(
		.INIT('h80)
	) name25107 (
		\m4_data_i[27]_pad ,
		_w8821_,
		_w8822_,
		_w27008_
	);
	LUT4 #(
		.INIT('h9dbf)
	) name25108 (
		_w8816_,
		_w8819_,
		_w27007_,
		_w27008_,
		_w27009_
	);
	LUT3 #(
		.INIT('h80)
	) name25109 (
		\m6_data_i[27]_pad ,
		_w8821_,
		_w8822_,
		_w27010_
	);
	LUT3 #(
		.INIT('h80)
	) name25110 (
		\m2_data_i[27]_pad ,
		_w8821_,
		_w8822_,
		_w27011_
	);
	LUT4 #(
		.INIT('habef)
	) name25111 (
		_w8816_,
		_w8819_,
		_w27010_,
		_w27011_,
		_w27012_
	);
	LUT3 #(
		.INIT('h2a)
	) name25112 (
		\m5_data_i[27]_pad ,
		_w8821_,
		_w8822_,
		_w27013_
	);
	LUT3 #(
		.INIT('h2a)
	) name25113 (
		\m1_data_i[27]_pad ,
		_w8821_,
		_w8822_,
		_w27014_
	);
	LUT4 #(
		.INIT('h57df)
	) name25114 (
		_w8816_,
		_w8819_,
		_w27013_,
		_w27014_,
		_w27015_
	);
	LUT3 #(
		.INIT('h80)
	) name25115 (
		\m0_data_i[27]_pad ,
		_w8821_,
		_w8822_,
		_w27016_
	);
	LUT3 #(
		.INIT('h2a)
	) name25116 (
		\m7_data_i[27]_pad ,
		_w8821_,
		_w8822_,
		_w27017_
	);
	LUT4 #(
		.INIT('h6e7f)
	) name25117 (
		_w8816_,
		_w8819_,
		_w27016_,
		_w27017_,
		_w27018_
	);
	LUT4 #(
		.INIT('h7fff)
	) name25118 (
		_w27009_,
		_w27012_,
		_w27015_,
		_w27018_,
		_w27019_
	);
	LUT3 #(
		.INIT('h2a)
	) name25119 (
		\m1_data_i[28]_pad ,
		_w8821_,
		_w8822_,
		_w27020_
	);
	LUT3 #(
		.INIT('h80)
	) name25120 (
		\m2_data_i[28]_pad ,
		_w8821_,
		_w8822_,
		_w27021_
	);
	LUT4 #(
		.INIT('h3b7f)
	) name25121 (
		_w8816_,
		_w8819_,
		_w27020_,
		_w27021_,
		_w27022_
	);
	LUT3 #(
		.INIT('h80)
	) name25122 (
		\m6_data_i[28]_pad ,
		_w8821_,
		_w8822_,
		_w27023_
	);
	LUT3 #(
		.INIT('h2a)
	) name25123 (
		\m7_data_i[28]_pad ,
		_w8821_,
		_w8822_,
		_w27024_
	);
	LUT3 #(
		.INIT('h57)
	) name25124 (
		_w8834_,
		_w27023_,
		_w27024_,
		_w27025_
	);
	LUT3 #(
		.INIT('h2a)
	) name25125 (
		\m5_data_i[28]_pad ,
		_w8821_,
		_w8822_,
		_w27026_
	);
	LUT3 #(
		.INIT('h80)
	) name25126 (
		\m0_data_i[28]_pad ,
		_w8821_,
		_w8822_,
		_w27027_
	);
	LUT4 #(
		.INIT('h57df)
	) name25127 (
		_w8816_,
		_w8819_,
		_w27026_,
		_w27027_,
		_w27028_
	);
	LUT3 #(
		.INIT('h2a)
	) name25128 (
		\m3_data_i[28]_pad ,
		_w8821_,
		_w8822_,
		_w27029_
	);
	LUT3 #(
		.INIT('h80)
	) name25129 (
		\m4_data_i[28]_pad ,
		_w8821_,
		_w8822_,
		_w27030_
	);
	LUT4 #(
		.INIT('h9dbf)
	) name25130 (
		_w8816_,
		_w8819_,
		_w27029_,
		_w27030_,
		_w27031_
	);
	LUT4 #(
		.INIT('h7fff)
	) name25131 (
		_w27022_,
		_w27025_,
		_w27028_,
		_w27031_,
		_w27032_
	);
	LUT3 #(
		.INIT('h2a)
	) name25132 (
		\m3_data_i[29]_pad ,
		_w8821_,
		_w8822_,
		_w27033_
	);
	LUT3 #(
		.INIT('h80)
	) name25133 (
		\m4_data_i[29]_pad ,
		_w8821_,
		_w8822_,
		_w27034_
	);
	LUT4 #(
		.INIT('h9dbf)
	) name25134 (
		_w8816_,
		_w8819_,
		_w27033_,
		_w27034_,
		_w27035_
	);
	LUT3 #(
		.INIT('h80)
	) name25135 (
		\m6_data_i[29]_pad ,
		_w8821_,
		_w8822_,
		_w27036_
	);
	LUT3 #(
		.INIT('h80)
	) name25136 (
		\m2_data_i[29]_pad ,
		_w8821_,
		_w8822_,
		_w27037_
	);
	LUT4 #(
		.INIT('habef)
	) name25137 (
		_w8816_,
		_w8819_,
		_w27036_,
		_w27037_,
		_w27038_
	);
	LUT3 #(
		.INIT('h2a)
	) name25138 (
		\m5_data_i[29]_pad ,
		_w8821_,
		_w8822_,
		_w27039_
	);
	LUT3 #(
		.INIT('h2a)
	) name25139 (
		\m1_data_i[29]_pad ,
		_w8821_,
		_w8822_,
		_w27040_
	);
	LUT4 #(
		.INIT('h57df)
	) name25140 (
		_w8816_,
		_w8819_,
		_w27039_,
		_w27040_,
		_w27041_
	);
	LUT3 #(
		.INIT('h80)
	) name25141 (
		\m0_data_i[29]_pad ,
		_w8821_,
		_w8822_,
		_w27042_
	);
	LUT3 #(
		.INIT('h2a)
	) name25142 (
		\m7_data_i[29]_pad ,
		_w8821_,
		_w8822_,
		_w27043_
	);
	LUT4 #(
		.INIT('h6e7f)
	) name25143 (
		_w8816_,
		_w8819_,
		_w27042_,
		_w27043_,
		_w27044_
	);
	LUT4 #(
		.INIT('h7fff)
	) name25144 (
		_w27035_,
		_w27038_,
		_w27041_,
		_w27044_,
		_w27045_
	);
	LUT3 #(
		.INIT('h2a)
	) name25145 (
		\m3_data_i[2]_pad ,
		_w8821_,
		_w8822_,
		_w27046_
	);
	LUT3 #(
		.INIT('h80)
	) name25146 (
		\m4_data_i[2]_pad ,
		_w8821_,
		_w8822_,
		_w27047_
	);
	LUT4 #(
		.INIT('h9dbf)
	) name25147 (
		_w8816_,
		_w8819_,
		_w27046_,
		_w27047_,
		_w27048_
	);
	LUT3 #(
		.INIT('h80)
	) name25148 (
		\m6_data_i[2]_pad ,
		_w8821_,
		_w8822_,
		_w27049_
	);
	LUT3 #(
		.INIT('h80)
	) name25149 (
		\m2_data_i[2]_pad ,
		_w8821_,
		_w8822_,
		_w27050_
	);
	LUT4 #(
		.INIT('habef)
	) name25150 (
		_w8816_,
		_w8819_,
		_w27049_,
		_w27050_,
		_w27051_
	);
	LUT3 #(
		.INIT('h2a)
	) name25151 (
		\m5_data_i[2]_pad ,
		_w8821_,
		_w8822_,
		_w27052_
	);
	LUT3 #(
		.INIT('h2a)
	) name25152 (
		\m1_data_i[2]_pad ,
		_w8821_,
		_w8822_,
		_w27053_
	);
	LUT4 #(
		.INIT('h57df)
	) name25153 (
		_w8816_,
		_w8819_,
		_w27052_,
		_w27053_,
		_w27054_
	);
	LUT3 #(
		.INIT('h80)
	) name25154 (
		\m0_data_i[2]_pad ,
		_w8821_,
		_w8822_,
		_w27055_
	);
	LUT3 #(
		.INIT('h2a)
	) name25155 (
		\m7_data_i[2]_pad ,
		_w8821_,
		_w8822_,
		_w27056_
	);
	LUT4 #(
		.INIT('h6e7f)
	) name25156 (
		_w8816_,
		_w8819_,
		_w27055_,
		_w27056_,
		_w27057_
	);
	LUT4 #(
		.INIT('h7fff)
	) name25157 (
		_w27048_,
		_w27051_,
		_w27054_,
		_w27057_,
		_w27058_
	);
	LUT3 #(
		.INIT('h80)
	) name25158 (
		\m0_data_i[30]_pad ,
		_w8821_,
		_w8822_,
		_w27059_
	);
	LUT3 #(
		.INIT('h2a)
	) name25159 (
		\m7_data_i[30]_pad ,
		_w8821_,
		_w8822_,
		_w27060_
	);
	LUT4 #(
		.INIT('h6e7f)
	) name25160 (
		_w8816_,
		_w8819_,
		_w27059_,
		_w27060_,
		_w27061_
	);
	LUT3 #(
		.INIT('h2a)
	) name25161 (
		\m3_data_i[30]_pad ,
		_w8821_,
		_w8822_,
		_w27062_
	);
	LUT3 #(
		.INIT('h2a)
	) name25162 (
		\m5_data_i[30]_pad ,
		_w8821_,
		_w8822_,
		_w27063_
	);
	LUT4 #(
		.INIT('h9dbf)
	) name25163 (
		_w8816_,
		_w8819_,
		_w27062_,
		_w27063_,
		_w27064_
	);
	LUT3 #(
		.INIT('h80)
	) name25164 (
		\m4_data_i[30]_pad ,
		_w8821_,
		_w8822_,
		_w27065_
	);
	LUT3 #(
		.INIT('h80)
	) name25165 (
		\m6_data_i[30]_pad ,
		_w8821_,
		_w8822_,
		_w27066_
	);
	LUT4 #(
		.INIT('hcedf)
	) name25166 (
		_w8816_,
		_w8819_,
		_w27065_,
		_w27066_,
		_w27067_
	);
	LUT3 #(
		.INIT('h2a)
	) name25167 (
		\m1_data_i[30]_pad ,
		_w8821_,
		_w8822_,
		_w27068_
	);
	LUT3 #(
		.INIT('h80)
	) name25168 (
		\m2_data_i[30]_pad ,
		_w8821_,
		_w8822_,
		_w27069_
	);
	LUT4 #(
		.INIT('h3b7f)
	) name25169 (
		_w8816_,
		_w8819_,
		_w27068_,
		_w27069_,
		_w27070_
	);
	LUT4 #(
		.INIT('h7fff)
	) name25170 (
		_w27061_,
		_w27064_,
		_w27067_,
		_w27070_,
		_w27071_
	);
	LUT3 #(
		.INIT('h2a)
	) name25171 (
		\m1_data_i[31]_pad ,
		_w8821_,
		_w8822_,
		_w27072_
	);
	LUT3 #(
		.INIT('h80)
	) name25172 (
		\m2_data_i[31]_pad ,
		_w8821_,
		_w8822_,
		_w27073_
	);
	LUT4 #(
		.INIT('h3b7f)
	) name25173 (
		_w8816_,
		_w8819_,
		_w27072_,
		_w27073_,
		_w27074_
	);
	LUT3 #(
		.INIT('h2a)
	) name25174 (
		\m3_data_i[31]_pad ,
		_w8821_,
		_w8822_,
		_w27075_
	);
	LUT3 #(
		.INIT('h2a)
	) name25175 (
		\m7_data_i[31]_pad ,
		_w8821_,
		_w8822_,
		_w27076_
	);
	LUT4 #(
		.INIT('haebf)
	) name25176 (
		_w8816_,
		_w8819_,
		_w27075_,
		_w27076_,
		_w27077_
	);
	LUT3 #(
		.INIT('h80)
	) name25177 (
		\m4_data_i[31]_pad ,
		_w8821_,
		_w8822_,
		_w27078_
	);
	LUT3 #(
		.INIT('h80)
	) name25178 (
		\m0_data_i[31]_pad ,
		_w8821_,
		_w8822_,
		_w27079_
	);
	LUT4 #(
		.INIT('h57df)
	) name25179 (
		_w8816_,
		_w8819_,
		_w27078_,
		_w27079_,
		_w27080_
	);
	LUT3 #(
		.INIT('h80)
	) name25180 (
		\m6_data_i[31]_pad ,
		_w8821_,
		_w8822_,
		_w27081_
	);
	LUT3 #(
		.INIT('h2a)
	) name25181 (
		\m5_data_i[31]_pad ,
		_w8821_,
		_w8822_,
		_w27082_
	);
	LUT4 #(
		.INIT('hcdef)
	) name25182 (
		_w8816_,
		_w8819_,
		_w27081_,
		_w27082_,
		_w27083_
	);
	LUT4 #(
		.INIT('h7fff)
	) name25183 (
		_w27074_,
		_w27077_,
		_w27080_,
		_w27083_,
		_w27084_
	);
	LUT3 #(
		.INIT('h2a)
	) name25184 (
		\m1_data_i[3]_pad ,
		_w8821_,
		_w8822_,
		_w27085_
	);
	LUT3 #(
		.INIT('h80)
	) name25185 (
		\m2_data_i[3]_pad ,
		_w8821_,
		_w8822_,
		_w27086_
	);
	LUT4 #(
		.INIT('h3b7f)
	) name25186 (
		_w8816_,
		_w8819_,
		_w27085_,
		_w27086_,
		_w27087_
	);
	LUT3 #(
		.INIT('h80)
	) name25187 (
		\m6_data_i[3]_pad ,
		_w8821_,
		_w8822_,
		_w27088_
	);
	LUT3 #(
		.INIT('h2a)
	) name25188 (
		\m7_data_i[3]_pad ,
		_w8821_,
		_w8822_,
		_w27089_
	);
	LUT3 #(
		.INIT('h57)
	) name25189 (
		_w8834_,
		_w27088_,
		_w27089_,
		_w27090_
	);
	LUT3 #(
		.INIT('h2a)
	) name25190 (
		\m5_data_i[3]_pad ,
		_w8821_,
		_w8822_,
		_w27091_
	);
	LUT3 #(
		.INIT('h80)
	) name25191 (
		\m0_data_i[3]_pad ,
		_w8821_,
		_w8822_,
		_w27092_
	);
	LUT4 #(
		.INIT('h57df)
	) name25192 (
		_w8816_,
		_w8819_,
		_w27091_,
		_w27092_,
		_w27093_
	);
	LUT3 #(
		.INIT('h2a)
	) name25193 (
		\m3_data_i[3]_pad ,
		_w8821_,
		_w8822_,
		_w27094_
	);
	LUT3 #(
		.INIT('h80)
	) name25194 (
		\m4_data_i[3]_pad ,
		_w8821_,
		_w8822_,
		_w27095_
	);
	LUT4 #(
		.INIT('h9dbf)
	) name25195 (
		_w8816_,
		_w8819_,
		_w27094_,
		_w27095_,
		_w27096_
	);
	LUT4 #(
		.INIT('h7fff)
	) name25196 (
		_w27087_,
		_w27090_,
		_w27093_,
		_w27096_,
		_w27097_
	);
	LUT3 #(
		.INIT('h80)
	) name25197 (
		\m0_data_i[4]_pad ,
		_w8821_,
		_w8822_,
		_w27098_
	);
	LUT3 #(
		.INIT('h2a)
	) name25198 (
		\m7_data_i[4]_pad ,
		_w8821_,
		_w8822_,
		_w27099_
	);
	LUT4 #(
		.INIT('h6e7f)
	) name25199 (
		_w8816_,
		_w8819_,
		_w27098_,
		_w27099_,
		_w27100_
	);
	LUT3 #(
		.INIT('h2a)
	) name25200 (
		\m3_data_i[4]_pad ,
		_w8821_,
		_w8822_,
		_w27101_
	);
	LUT3 #(
		.INIT('h80)
	) name25201 (
		\m2_data_i[4]_pad ,
		_w8821_,
		_w8822_,
		_w27102_
	);
	LUT3 #(
		.INIT('h57)
	) name25202 (
		_w8828_,
		_w27101_,
		_w27102_,
		_w27103_
	);
	LUT3 #(
		.INIT('h80)
	) name25203 (
		\m4_data_i[4]_pad ,
		_w8821_,
		_w8822_,
		_w27104_
	);
	LUT3 #(
		.INIT('h2a)
	) name25204 (
		\m1_data_i[4]_pad ,
		_w8821_,
		_w8822_,
		_w27105_
	);
	LUT4 #(
		.INIT('h57df)
	) name25205 (
		_w8816_,
		_w8819_,
		_w27104_,
		_w27105_,
		_w27106_
	);
	LUT3 #(
		.INIT('h80)
	) name25206 (
		\m6_data_i[4]_pad ,
		_w8821_,
		_w8822_,
		_w27107_
	);
	LUT3 #(
		.INIT('h2a)
	) name25207 (
		\m5_data_i[4]_pad ,
		_w8821_,
		_w8822_,
		_w27108_
	);
	LUT4 #(
		.INIT('hcdef)
	) name25208 (
		_w8816_,
		_w8819_,
		_w27107_,
		_w27108_,
		_w27109_
	);
	LUT4 #(
		.INIT('h7fff)
	) name25209 (
		_w27100_,
		_w27103_,
		_w27106_,
		_w27109_,
		_w27110_
	);
	LUT3 #(
		.INIT('h2a)
	) name25210 (
		\m3_data_i[5]_pad ,
		_w8821_,
		_w8822_,
		_w27111_
	);
	LUT3 #(
		.INIT('h80)
	) name25211 (
		\m4_data_i[5]_pad ,
		_w8821_,
		_w8822_,
		_w27112_
	);
	LUT4 #(
		.INIT('h9dbf)
	) name25212 (
		_w8816_,
		_w8819_,
		_w27111_,
		_w27112_,
		_w27113_
	);
	LUT3 #(
		.INIT('h80)
	) name25213 (
		\m6_data_i[5]_pad ,
		_w8821_,
		_w8822_,
		_w27114_
	);
	LUT3 #(
		.INIT('h80)
	) name25214 (
		\m2_data_i[5]_pad ,
		_w8821_,
		_w8822_,
		_w27115_
	);
	LUT4 #(
		.INIT('habef)
	) name25215 (
		_w8816_,
		_w8819_,
		_w27114_,
		_w27115_,
		_w27116_
	);
	LUT3 #(
		.INIT('h2a)
	) name25216 (
		\m5_data_i[5]_pad ,
		_w8821_,
		_w8822_,
		_w27117_
	);
	LUT3 #(
		.INIT('h2a)
	) name25217 (
		\m1_data_i[5]_pad ,
		_w8821_,
		_w8822_,
		_w27118_
	);
	LUT4 #(
		.INIT('h57df)
	) name25218 (
		_w8816_,
		_w8819_,
		_w27117_,
		_w27118_,
		_w27119_
	);
	LUT3 #(
		.INIT('h80)
	) name25219 (
		\m0_data_i[5]_pad ,
		_w8821_,
		_w8822_,
		_w27120_
	);
	LUT3 #(
		.INIT('h2a)
	) name25220 (
		\m7_data_i[5]_pad ,
		_w8821_,
		_w8822_,
		_w27121_
	);
	LUT4 #(
		.INIT('h6e7f)
	) name25221 (
		_w8816_,
		_w8819_,
		_w27120_,
		_w27121_,
		_w27122_
	);
	LUT4 #(
		.INIT('h7fff)
	) name25222 (
		_w27113_,
		_w27116_,
		_w27119_,
		_w27122_,
		_w27123_
	);
	LUT3 #(
		.INIT('h2a)
	) name25223 (
		\m3_data_i[6]_pad ,
		_w8821_,
		_w8822_,
		_w27124_
	);
	LUT3 #(
		.INIT('h80)
	) name25224 (
		\m4_data_i[6]_pad ,
		_w8821_,
		_w8822_,
		_w27125_
	);
	LUT4 #(
		.INIT('h9dbf)
	) name25225 (
		_w8816_,
		_w8819_,
		_w27124_,
		_w27125_,
		_w27126_
	);
	LUT3 #(
		.INIT('h80)
	) name25226 (
		\m6_data_i[6]_pad ,
		_w8821_,
		_w8822_,
		_w27127_
	);
	LUT3 #(
		.INIT('h2a)
	) name25227 (
		\m7_data_i[6]_pad ,
		_w8821_,
		_w8822_,
		_w27128_
	);
	LUT3 #(
		.INIT('h57)
	) name25228 (
		_w8834_,
		_w27127_,
		_w27128_,
		_w27129_
	);
	LUT3 #(
		.INIT('h2a)
	) name25229 (
		\m5_data_i[6]_pad ,
		_w8821_,
		_w8822_,
		_w27130_
	);
	LUT3 #(
		.INIT('h80)
	) name25230 (
		\m0_data_i[6]_pad ,
		_w8821_,
		_w8822_,
		_w27131_
	);
	LUT4 #(
		.INIT('h57df)
	) name25231 (
		_w8816_,
		_w8819_,
		_w27130_,
		_w27131_,
		_w27132_
	);
	LUT3 #(
		.INIT('h2a)
	) name25232 (
		\m1_data_i[6]_pad ,
		_w8821_,
		_w8822_,
		_w27133_
	);
	LUT3 #(
		.INIT('h80)
	) name25233 (
		\m2_data_i[6]_pad ,
		_w8821_,
		_w8822_,
		_w27134_
	);
	LUT4 #(
		.INIT('h3b7f)
	) name25234 (
		_w8816_,
		_w8819_,
		_w27133_,
		_w27134_,
		_w27135_
	);
	LUT4 #(
		.INIT('h7fff)
	) name25235 (
		_w27126_,
		_w27129_,
		_w27132_,
		_w27135_,
		_w27136_
	);
	LUT3 #(
		.INIT('h2a)
	) name25236 (
		\m3_data_i[7]_pad ,
		_w8821_,
		_w8822_,
		_w27137_
	);
	LUT3 #(
		.INIT('h80)
	) name25237 (
		\m4_data_i[7]_pad ,
		_w8821_,
		_w8822_,
		_w27138_
	);
	LUT4 #(
		.INIT('h9dbf)
	) name25238 (
		_w8816_,
		_w8819_,
		_w27137_,
		_w27138_,
		_w27139_
	);
	LUT3 #(
		.INIT('h80)
	) name25239 (
		\m6_data_i[7]_pad ,
		_w8821_,
		_w8822_,
		_w27140_
	);
	LUT3 #(
		.INIT('h80)
	) name25240 (
		\m2_data_i[7]_pad ,
		_w8821_,
		_w8822_,
		_w27141_
	);
	LUT4 #(
		.INIT('habef)
	) name25241 (
		_w8816_,
		_w8819_,
		_w27140_,
		_w27141_,
		_w27142_
	);
	LUT3 #(
		.INIT('h2a)
	) name25242 (
		\m5_data_i[7]_pad ,
		_w8821_,
		_w8822_,
		_w27143_
	);
	LUT3 #(
		.INIT('h2a)
	) name25243 (
		\m1_data_i[7]_pad ,
		_w8821_,
		_w8822_,
		_w27144_
	);
	LUT4 #(
		.INIT('h57df)
	) name25244 (
		_w8816_,
		_w8819_,
		_w27143_,
		_w27144_,
		_w27145_
	);
	LUT3 #(
		.INIT('h80)
	) name25245 (
		\m0_data_i[7]_pad ,
		_w8821_,
		_w8822_,
		_w27146_
	);
	LUT3 #(
		.INIT('h2a)
	) name25246 (
		\m7_data_i[7]_pad ,
		_w8821_,
		_w8822_,
		_w27147_
	);
	LUT4 #(
		.INIT('h6e7f)
	) name25247 (
		_w8816_,
		_w8819_,
		_w27146_,
		_w27147_,
		_w27148_
	);
	LUT4 #(
		.INIT('h7fff)
	) name25248 (
		_w27139_,
		_w27142_,
		_w27145_,
		_w27148_,
		_w27149_
	);
	LUT3 #(
		.INIT('h2a)
	) name25249 (
		\m1_data_i[8]_pad ,
		_w8821_,
		_w8822_,
		_w27150_
	);
	LUT3 #(
		.INIT('h80)
	) name25250 (
		\m2_data_i[8]_pad ,
		_w8821_,
		_w8822_,
		_w27151_
	);
	LUT4 #(
		.INIT('h3b7f)
	) name25251 (
		_w8816_,
		_w8819_,
		_w27150_,
		_w27151_,
		_w27152_
	);
	LUT3 #(
		.INIT('h2a)
	) name25252 (
		\m3_data_i[8]_pad ,
		_w8821_,
		_w8822_,
		_w27153_
	);
	LUT3 #(
		.INIT('h2a)
	) name25253 (
		\m7_data_i[8]_pad ,
		_w8821_,
		_w8822_,
		_w27154_
	);
	LUT4 #(
		.INIT('haebf)
	) name25254 (
		_w8816_,
		_w8819_,
		_w27153_,
		_w27154_,
		_w27155_
	);
	LUT3 #(
		.INIT('h80)
	) name25255 (
		\m4_data_i[8]_pad ,
		_w8821_,
		_w8822_,
		_w27156_
	);
	LUT3 #(
		.INIT('h80)
	) name25256 (
		\m0_data_i[8]_pad ,
		_w8821_,
		_w8822_,
		_w27157_
	);
	LUT4 #(
		.INIT('h57df)
	) name25257 (
		_w8816_,
		_w8819_,
		_w27156_,
		_w27157_,
		_w27158_
	);
	LUT3 #(
		.INIT('h80)
	) name25258 (
		\m6_data_i[8]_pad ,
		_w8821_,
		_w8822_,
		_w27159_
	);
	LUT3 #(
		.INIT('h2a)
	) name25259 (
		\m5_data_i[8]_pad ,
		_w8821_,
		_w8822_,
		_w27160_
	);
	LUT4 #(
		.INIT('hcdef)
	) name25260 (
		_w8816_,
		_w8819_,
		_w27159_,
		_w27160_,
		_w27161_
	);
	LUT4 #(
		.INIT('h7fff)
	) name25261 (
		_w27152_,
		_w27155_,
		_w27158_,
		_w27161_,
		_w27162_
	);
	LUT3 #(
		.INIT('h2a)
	) name25262 (
		\m3_data_i[9]_pad ,
		_w8821_,
		_w8822_,
		_w27163_
	);
	LUT3 #(
		.INIT('h80)
	) name25263 (
		\m4_data_i[9]_pad ,
		_w8821_,
		_w8822_,
		_w27164_
	);
	LUT4 #(
		.INIT('h9dbf)
	) name25264 (
		_w8816_,
		_w8819_,
		_w27163_,
		_w27164_,
		_w27165_
	);
	LUT3 #(
		.INIT('h80)
	) name25265 (
		\m6_data_i[9]_pad ,
		_w8821_,
		_w8822_,
		_w27166_
	);
	LUT3 #(
		.INIT('h2a)
	) name25266 (
		\m7_data_i[9]_pad ,
		_w8821_,
		_w8822_,
		_w27167_
	);
	LUT3 #(
		.INIT('h57)
	) name25267 (
		_w8834_,
		_w27166_,
		_w27167_,
		_w27168_
	);
	LUT3 #(
		.INIT('h2a)
	) name25268 (
		\m5_data_i[9]_pad ,
		_w8821_,
		_w8822_,
		_w27169_
	);
	LUT3 #(
		.INIT('h80)
	) name25269 (
		\m0_data_i[9]_pad ,
		_w8821_,
		_w8822_,
		_w27170_
	);
	LUT4 #(
		.INIT('h57df)
	) name25270 (
		_w8816_,
		_w8819_,
		_w27169_,
		_w27170_,
		_w27171_
	);
	LUT3 #(
		.INIT('h2a)
	) name25271 (
		\m1_data_i[9]_pad ,
		_w8821_,
		_w8822_,
		_w27172_
	);
	LUT3 #(
		.INIT('h80)
	) name25272 (
		\m2_data_i[9]_pad ,
		_w8821_,
		_w8822_,
		_w27173_
	);
	LUT4 #(
		.INIT('h3b7f)
	) name25273 (
		_w8816_,
		_w8819_,
		_w27172_,
		_w27173_,
		_w27174_
	);
	LUT4 #(
		.INIT('h7fff)
	) name25274 (
		_w27165_,
		_w27168_,
		_w27171_,
		_w27174_,
		_w27175_
	);
	LUT3 #(
		.INIT('h2a)
	) name25275 (
		\m1_sel_i[0]_pad ,
		_w8821_,
		_w8822_,
		_w27176_
	);
	LUT3 #(
		.INIT('h80)
	) name25276 (
		\m2_sel_i[0]_pad ,
		_w8821_,
		_w8822_,
		_w27177_
	);
	LUT4 #(
		.INIT('h3b7f)
	) name25277 (
		_w8816_,
		_w8819_,
		_w27176_,
		_w27177_,
		_w27178_
	);
	LUT3 #(
		.INIT('h80)
	) name25278 (
		\m6_sel_i[0]_pad ,
		_w8821_,
		_w8822_,
		_w27179_
	);
	LUT3 #(
		.INIT('h2a)
	) name25279 (
		\m7_sel_i[0]_pad ,
		_w8821_,
		_w8822_,
		_w27180_
	);
	LUT3 #(
		.INIT('h57)
	) name25280 (
		_w8834_,
		_w27179_,
		_w27180_,
		_w27181_
	);
	LUT3 #(
		.INIT('h2a)
	) name25281 (
		\m5_sel_i[0]_pad ,
		_w8821_,
		_w8822_,
		_w27182_
	);
	LUT3 #(
		.INIT('h80)
	) name25282 (
		\m0_sel_i[0]_pad ,
		_w8821_,
		_w8822_,
		_w27183_
	);
	LUT4 #(
		.INIT('h57df)
	) name25283 (
		_w8816_,
		_w8819_,
		_w27182_,
		_w27183_,
		_w27184_
	);
	LUT3 #(
		.INIT('h2a)
	) name25284 (
		\m3_sel_i[0]_pad ,
		_w8821_,
		_w8822_,
		_w27185_
	);
	LUT3 #(
		.INIT('h80)
	) name25285 (
		\m4_sel_i[0]_pad ,
		_w8821_,
		_w8822_,
		_w27186_
	);
	LUT4 #(
		.INIT('h9dbf)
	) name25286 (
		_w8816_,
		_w8819_,
		_w27185_,
		_w27186_,
		_w27187_
	);
	LUT4 #(
		.INIT('h7fff)
	) name25287 (
		_w27178_,
		_w27181_,
		_w27184_,
		_w27187_,
		_w27188_
	);
	LUT3 #(
		.INIT('h2a)
	) name25288 (
		\m3_sel_i[1]_pad ,
		_w8821_,
		_w8822_,
		_w27189_
	);
	LUT3 #(
		.INIT('h80)
	) name25289 (
		\m4_sel_i[1]_pad ,
		_w8821_,
		_w8822_,
		_w27190_
	);
	LUT4 #(
		.INIT('h9dbf)
	) name25290 (
		_w8816_,
		_w8819_,
		_w27189_,
		_w27190_,
		_w27191_
	);
	LUT3 #(
		.INIT('h80)
	) name25291 (
		\m6_sel_i[1]_pad ,
		_w8821_,
		_w8822_,
		_w27192_
	);
	LUT3 #(
		.INIT('h2a)
	) name25292 (
		\m7_sel_i[1]_pad ,
		_w8821_,
		_w8822_,
		_w27193_
	);
	LUT3 #(
		.INIT('h57)
	) name25293 (
		_w8834_,
		_w27192_,
		_w27193_,
		_w27194_
	);
	LUT3 #(
		.INIT('h2a)
	) name25294 (
		\m5_sel_i[1]_pad ,
		_w8821_,
		_w8822_,
		_w27195_
	);
	LUT3 #(
		.INIT('h80)
	) name25295 (
		\m0_sel_i[1]_pad ,
		_w8821_,
		_w8822_,
		_w27196_
	);
	LUT4 #(
		.INIT('h57df)
	) name25296 (
		_w8816_,
		_w8819_,
		_w27195_,
		_w27196_,
		_w27197_
	);
	LUT3 #(
		.INIT('h2a)
	) name25297 (
		\m1_sel_i[1]_pad ,
		_w8821_,
		_w8822_,
		_w27198_
	);
	LUT3 #(
		.INIT('h80)
	) name25298 (
		\m2_sel_i[1]_pad ,
		_w8821_,
		_w8822_,
		_w27199_
	);
	LUT4 #(
		.INIT('h3b7f)
	) name25299 (
		_w8816_,
		_w8819_,
		_w27198_,
		_w27199_,
		_w27200_
	);
	LUT4 #(
		.INIT('h7fff)
	) name25300 (
		_w27191_,
		_w27194_,
		_w27197_,
		_w27200_,
		_w27201_
	);
	LUT3 #(
		.INIT('h80)
	) name25301 (
		\m0_sel_i[2]_pad ,
		_w8821_,
		_w8822_,
		_w27202_
	);
	LUT3 #(
		.INIT('h2a)
	) name25302 (
		\m7_sel_i[2]_pad ,
		_w8821_,
		_w8822_,
		_w27203_
	);
	LUT4 #(
		.INIT('h6e7f)
	) name25303 (
		_w8816_,
		_w8819_,
		_w27202_,
		_w27203_,
		_w27204_
	);
	LUT3 #(
		.INIT('h2a)
	) name25304 (
		\m3_sel_i[2]_pad ,
		_w8821_,
		_w8822_,
		_w27205_
	);
	LUT3 #(
		.INIT('h80)
	) name25305 (
		\m2_sel_i[2]_pad ,
		_w8821_,
		_w8822_,
		_w27206_
	);
	LUT3 #(
		.INIT('h57)
	) name25306 (
		_w8828_,
		_w27205_,
		_w27206_,
		_w27207_
	);
	LUT3 #(
		.INIT('h80)
	) name25307 (
		\m4_sel_i[2]_pad ,
		_w8821_,
		_w8822_,
		_w27208_
	);
	LUT3 #(
		.INIT('h2a)
	) name25308 (
		\m1_sel_i[2]_pad ,
		_w8821_,
		_w8822_,
		_w27209_
	);
	LUT4 #(
		.INIT('h57df)
	) name25309 (
		_w8816_,
		_w8819_,
		_w27208_,
		_w27209_,
		_w27210_
	);
	LUT3 #(
		.INIT('h80)
	) name25310 (
		\m6_sel_i[2]_pad ,
		_w8821_,
		_w8822_,
		_w27211_
	);
	LUT3 #(
		.INIT('h2a)
	) name25311 (
		\m5_sel_i[2]_pad ,
		_w8821_,
		_w8822_,
		_w27212_
	);
	LUT4 #(
		.INIT('hcdef)
	) name25312 (
		_w8816_,
		_w8819_,
		_w27211_,
		_w27212_,
		_w27213_
	);
	LUT4 #(
		.INIT('h7fff)
	) name25313 (
		_w27204_,
		_w27207_,
		_w27210_,
		_w27213_,
		_w27214_
	);
	LUT3 #(
		.INIT('h2a)
	) name25314 (
		\m1_sel_i[3]_pad ,
		_w8821_,
		_w8822_,
		_w27215_
	);
	LUT3 #(
		.INIT('h80)
	) name25315 (
		\m2_sel_i[3]_pad ,
		_w8821_,
		_w8822_,
		_w27216_
	);
	LUT4 #(
		.INIT('h3b7f)
	) name25316 (
		_w8816_,
		_w8819_,
		_w27215_,
		_w27216_,
		_w27217_
	);
	LUT3 #(
		.INIT('h2a)
	) name25317 (
		\m3_sel_i[3]_pad ,
		_w8821_,
		_w8822_,
		_w27218_
	);
	LUT3 #(
		.INIT('h2a)
	) name25318 (
		\m7_sel_i[3]_pad ,
		_w8821_,
		_w8822_,
		_w27219_
	);
	LUT4 #(
		.INIT('haebf)
	) name25319 (
		_w8816_,
		_w8819_,
		_w27218_,
		_w27219_,
		_w27220_
	);
	LUT3 #(
		.INIT('h80)
	) name25320 (
		\m4_sel_i[3]_pad ,
		_w8821_,
		_w8822_,
		_w27221_
	);
	LUT3 #(
		.INIT('h80)
	) name25321 (
		\m0_sel_i[3]_pad ,
		_w8821_,
		_w8822_,
		_w27222_
	);
	LUT4 #(
		.INIT('h57df)
	) name25322 (
		_w8816_,
		_w8819_,
		_w27221_,
		_w27222_,
		_w27223_
	);
	LUT3 #(
		.INIT('h80)
	) name25323 (
		\m6_sel_i[3]_pad ,
		_w8821_,
		_w8822_,
		_w27224_
	);
	LUT3 #(
		.INIT('h2a)
	) name25324 (
		\m5_sel_i[3]_pad ,
		_w8821_,
		_w8822_,
		_w27225_
	);
	LUT4 #(
		.INIT('hcdef)
	) name25325 (
		_w8816_,
		_w8819_,
		_w27224_,
		_w27225_,
		_w27226_
	);
	LUT4 #(
		.INIT('h7fff)
	) name25326 (
		_w27217_,
		_w27220_,
		_w27223_,
		_w27226_,
		_w27227_
	);
	LUT4 #(
		.INIT('h2a00)
	) name25327 (
		\m5_stb_i_pad ,
		_w8821_,
		_w8822_,
		_w9553_,
		_w27228_
	);
	LUT4 #(
		.INIT('h8000)
	) name25328 (
		\m4_stb_i_pad ,
		_w8821_,
		_w8822_,
		_w9360_,
		_w27229_
	);
	LUT3 #(
		.INIT('h57)
	) name25329 (
		_w8840_,
		_w27228_,
		_w27229_,
		_w27230_
	);
	LUT4 #(
		.INIT('h8000)
	) name25330 (
		\m6_stb_i_pad ,
		_w8821_,
		_w8822_,
		_w9342_,
		_w27231_
	);
	LUT4 #(
		.INIT('h2a00)
	) name25331 (
		\m1_stb_i_pad ,
		_w8821_,
		_w8822_,
		_w9445_,
		_w27232_
	);
	LUT4 #(
		.INIT('h67ef)
	) name25332 (
		_w8816_,
		_w8819_,
		_w27231_,
		_w27232_,
		_w27233_
	);
	LUT4 #(
		.INIT('h2a00)
	) name25333 (
		\m7_stb_i_pad ,
		_w8821_,
		_w8822_,
		_w9623_,
		_w27234_
	);
	LUT4 #(
		.INIT('h2a00)
	) name25334 (
		\m3_stb_i_pad ,
		_w8821_,
		_w8822_,
		_w9503_,
		_w27235_
	);
	LUT4 #(
		.INIT('habef)
	) name25335 (
		_w8816_,
		_w8819_,
		_w27234_,
		_w27235_,
		_w27236_
	);
	LUT4 #(
		.INIT('h8000)
	) name25336 (
		\m2_stb_i_pad ,
		_w8821_,
		_w8822_,
		_w9620_,
		_w27237_
	);
	LUT4 #(
		.INIT('h8000)
	) name25337 (
		\m0_stb_i_pad ,
		_w8821_,
		_w8822_,
		_w9410_,
		_w27238_
	);
	LUT4 #(
		.INIT('h37bf)
	) name25338 (
		_w8816_,
		_w8819_,
		_w27237_,
		_w27238_,
		_w27239_
	);
	LUT4 #(
		.INIT('h7fff)
	) name25339 (
		_w27230_,
		_w27233_,
		_w27236_,
		_w27239_,
		_w27240_
	);
	LUT3 #(
		.INIT('h80)
	) name25340 (
		\m6_we_i_pad ,
		_w8821_,
		_w8822_,
		_w27241_
	);
	LUT3 #(
		.INIT('h2a)
	) name25341 (
		\m5_we_i_pad ,
		_w8821_,
		_w8822_,
		_w27242_
	);
	LUT4 #(
		.INIT('hcdef)
	) name25342 (
		_w8816_,
		_w8819_,
		_w27241_,
		_w27242_,
		_w27243_
	);
	LUT3 #(
		.INIT('h2a)
	) name25343 (
		\m3_we_i_pad ,
		_w8821_,
		_w8822_,
		_w27244_
	);
	LUT3 #(
		.INIT('h80)
	) name25344 (
		\m2_we_i_pad ,
		_w8821_,
		_w8822_,
		_w27245_
	);
	LUT3 #(
		.INIT('h57)
	) name25345 (
		_w8828_,
		_w27244_,
		_w27245_,
		_w27246_
	);
	LUT3 #(
		.INIT('h80)
	) name25346 (
		\m4_we_i_pad ,
		_w8821_,
		_w8822_,
		_w27247_
	);
	LUT3 #(
		.INIT('h2a)
	) name25347 (
		\m1_we_i_pad ,
		_w8821_,
		_w8822_,
		_w27248_
	);
	LUT4 #(
		.INIT('h57df)
	) name25348 (
		_w8816_,
		_w8819_,
		_w27247_,
		_w27248_,
		_w27249_
	);
	LUT3 #(
		.INIT('h80)
	) name25349 (
		\m0_we_i_pad ,
		_w8821_,
		_w8822_,
		_w27250_
	);
	LUT3 #(
		.INIT('h2a)
	) name25350 (
		\m7_we_i_pad ,
		_w8821_,
		_w8822_,
		_w27251_
	);
	LUT4 #(
		.INIT('h6e7f)
	) name25351 (
		_w8816_,
		_w8819_,
		_w27250_,
		_w27251_,
		_w27252_
	);
	LUT4 #(
		.INIT('h7fff)
	) name25352 (
		_w27243_,
		_w27246_,
		_w27249_,
		_w27252_,
		_w27253_
	);
	LUT3 #(
		.INIT('h2a)
	) name25353 (
		\m3_addr_i[0]_pad ,
		_w8865_,
		_w8866_,
		_w27254_
	);
	LUT3 #(
		.INIT('h80)
	) name25354 (
		\m4_addr_i[0]_pad ,
		_w8865_,
		_w8866_,
		_w27255_
	);
	LUT4 #(
		.INIT('h9dbf)
	) name25355 (
		_w8860_,
		_w8863_,
		_w27254_,
		_w27255_,
		_w27256_
	);
	LUT3 #(
		.INIT('h80)
	) name25356 (
		\m6_addr_i[0]_pad ,
		_w8865_,
		_w8866_,
		_w27257_
	);
	LUT3 #(
		.INIT('h80)
	) name25357 (
		\m2_addr_i[0]_pad ,
		_w8865_,
		_w8866_,
		_w27258_
	);
	LUT4 #(
		.INIT('habef)
	) name25358 (
		_w8860_,
		_w8863_,
		_w27257_,
		_w27258_,
		_w27259_
	);
	LUT3 #(
		.INIT('h2a)
	) name25359 (
		\m5_addr_i[0]_pad ,
		_w8865_,
		_w8866_,
		_w27260_
	);
	LUT3 #(
		.INIT('h2a)
	) name25360 (
		\m1_addr_i[0]_pad ,
		_w8865_,
		_w8866_,
		_w27261_
	);
	LUT4 #(
		.INIT('h57df)
	) name25361 (
		_w8860_,
		_w8863_,
		_w27260_,
		_w27261_,
		_w27262_
	);
	LUT3 #(
		.INIT('h80)
	) name25362 (
		\m0_addr_i[0]_pad ,
		_w8865_,
		_w8866_,
		_w27263_
	);
	LUT3 #(
		.INIT('h2a)
	) name25363 (
		\m7_addr_i[0]_pad ,
		_w8865_,
		_w8866_,
		_w27264_
	);
	LUT4 #(
		.INIT('h6e7f)
	) name25364 (
		_w8860_,
		_w8863_,
		_w27263_,
		_w27264_,
		_w27265_
	);
	LUT4 #(
		.INIT('h7fff)
	) name25365 (
		_w27256_,
		_w27259_,
		_w27262_,
		_w27265_,
		_w27266_
	);
	LUT3 #(
		.INIT('h2a)
	) name25366 (
		\m3_addr_i[10]_pad ,
		_w8865_,
		_w8866_,
		_w27267_
	);
	LUT3 #(
		.INIT('h80)
	) name25367 (
		\m4_addr_i[10]_pad ,
		_w8865_,
		_w8866_,
		_w27268_
	);
	LUT4 #(
		.INIT('h9dbf)
	) name25368 (
		_w8860_,
		_w8863_,
		_w27267_,
		_w27268_,
		_w27269_
	);
	LUT3 #(
		.INIT('h2a)
	) name25369 (
		\m1_addr_i[10]_pad ,
		_w8865_,
		_w8866_,
		_w27270_
	);
	LUT3 #(
		.INIT('h2a)
	) name25370 (
		\m5_addr_i[10]_pad ,
		_w8865_,
		_w8866_,
		_w27271_
	);
	LUT4 #(
		.INIT('h5d7f)
	) name25371 (
		_w8860_,
		_w8863_,
		_w27270_,
		_w27271_,
		_w27272_
	);
	LUT3 #(
		.INIT('h80)
	) name25372 (
		\m2_addr_i[10]_pad ,
		_w8865_,
		_w8866_,
		_w27273_
	);
	LUT3 #(
		.INIT('h80)
	) name25373 (
		\m6_addr_i[10]_pad ,
		_w8865_,
		_w8866_,
		_w27274_
	);
	LUT4 #(
		.INIT('haebf)
	) name25374 (
		_w8860_,
		_w8863_,
		_w27273_,
		_w27274_,
		_w27275_
	);
	LUT3 #(
		.INIT('h80)
	) name25375 (
		\m0_addr_i[10]_pad ,
		_w8865_,
		_w8866_,
		_w27276_
	);
	LUT3 #(
		.INIT('h2a)
	) name25376 (
		\m7_addr_i[10]_pad ,
		_w8865_,
		_w8866_,
		_w27277_
	);
	LUT4 #(
		.INIT('h6e7f)
	) name25377 (
		_w8860_,
		_w8863_,
		_w27276_,
		_w27277_,
		_w27278_
	);
	LUT4 #(
		.INIT('h7fff)
	) name25378 (
		_w27269_,
		_w27272_,
		_w27275_,
		_w27278_,
		_w27279_
	);
	LUT3 #(
		.INIT('h2a)
	) name25379 (
		\m3_addr_i[11]_pad ,
		_w8865_,
		_w8866_,
		_w27280_
	);
	LUT3 #(
		.INIT('h80)
	) name25380 (
		\m4_addr_i[11]_pad ,
		_w8865_,
		_w8866_,
		_w27281_
	);
	LUT4 #(
		.INIT('h9dbf)
	) name25381 (
		_w8860_,
		_w8863_,
		_w27280_,
		_w27281_,
		_w27282_
	);
	LUT3 #(
		.INIT('h2a)
	) name25382 (
		\m1_addr_i[11]_pad ,
		_w8865_,
		_w8866_,
		_w27283_
	);
	LUT3 #(
		.INIT('h2a)
	) name25383 (
		\m5_addr_i[11]_pad ,
		_w8865_,
		_w8866_,
		_w27284_
	);
	LUT4 #(
		.INIT('h5d7f)
	) name25384 (
		_w8860_,
		_w8863_,
		_w27283_,
		_w27284_,
		_w27285_
	);
	LUT3 #(
		.INIT('h80)
	) name25385 (
		\m2_addr_i[11]_pad ,
		_w8865_,
		_w8866_,
		_w27286_
	);
	LUT3 #(
		.INIT('h80)
	) name25386 (
		\m6_addr_i[11]_pad ,
		_w8865_,
		_w8866_,
		_w27287_
	);
	LUT4 #(
		.INIT('haebf)
	) name25387 (
		_w8860_,
		_w8863_,
		_w27286_,
		_w27287_,
		_w27288_
	);
	LUT3 #(
		.INIT('h80)
	) name25388 (
		\m0_addr_i[11]_pad ,
		_w8865_,
		_w8866_,
		_w27289_
	);
	LUT3 #(
		.INIT('h2a)
	) name25389 (
		\m7_addr_i[11]_pad ,
		_w8865_,
		_w8866_,
		_w27290_
	);
	LUT4 #(
		.INIT('h6e7f)
	) name25390 (
		_w8860_,
		_w8863_,
		_w27289_,
		_w27290_,
		_w27291_
	);
	LUT4 #(
		.INIT('h7fff)
	) name25391 (
		_w27282_,
		_w27285_,
		_w27288_,
		_w27291_,
		_w27292_
	);
	LUT3 #(
		.INIT('h2a)
	) name25392 (
		\m1_addr_i[12]_pad ,
		_w8865_,
		_w8866_,
		_w27293_
	);
	LUT3 #(
		.INIT('h80)
	) name25393 (
		\m2_addr_i[12]_pad ,
		_w8865_,
		_w8866_,
		_w27294_
	);
	LUT4 #(
		.INIT('h3b7f)
	) name25394 (
		_w8860_,
		_w8863_,
		_w27293_,
		_w27294_,
		_w27295_
	);
	LUT3 #(
		.INIT('h80)
	) name25395 (
		\m0_addr_i[12]_pad ,
		_w8865_,
		_w8866_,
		_w27296_
	);
	LUT3 #(
		.INIT('h80)
	) name25396 (
		\m4_addr_i[12]_pad ,
		_w8865_,
		_w8866_,
		_w27297_
	);
	LUT4 #(
		.INIT('h5d7f)
	) name25397 (
		_w8860_,
		_w8863_,
		_w27296_,
		_w27297_,
		_w27298_
	);
	LUT3 #(
		.INIT('h2a)
	) name25398 (
		\m7_addr_i[12]_pad ,
		_w8865_,
		_w8866_,
		_w27299_
	);
	LUT3 #(
		.INIT('h2a)
	) name25399 (
		\m3_addr_i[12]_pad ,
		_w8865_,
		_w8866_,
		_w27300_
	);
	LUT4 #(
		.INIT('habef)
	) name25400 (
		_w8860_,
		_w8863_,
		_w27299_,
		_w27300_,
		_w27301_
	);
	LUT3 #(
		.INIT('h80)
	) name25401 (
		\m6_addr_i[12]_pad ,
		_w8865_,
		_w8866_,
		_w27302_
	);
	LUT3 #(
		.INIT('h2a)
	) name25402 (
		\m5_addr_i[12]_pad ,
		_w8865_,
		_w8866_,
		_w27303_
	);
	LUT4 #(
		.INIT('hcdef)
	) name25403 (
		_w8860_,
		_w8863_,
		_w27302_,
		_w27303_,
		_w27304_
	);
	LUT4 #(
		.INIT('h7fff)
	) name25404 (
		_w27295_,
		_w27298_,
		_w27301_,
		_w27304_,
		_w27305_
	);
	LUT3 #(
		.INIT('h80)
	) name25405 (
		\m0_addr_i[13]_pad ,
		_w8865_,
		_w8866_,
		_w27306_
	);
	LUT3 #(
		.INIT('h2a)
	) name25406 (
		\m7_addr_i[13]_pad ,
		_w8865_,
		_w8866_,
		_w27307_
	);
	LUT4 #(
		.INIT('h6e7f)
	) name25407 (
		_w8860_,
		_w8863_,
		_w27306_,
		_w27307_,
		_w27308_
	);
	LUT3 #(
		.INIT('h2a)
	) name25408 (
		\m1_addr_i[13]_pad ,
		_w8865_,
		_w8866_,
		_w27309_
	);
	LUT3 #(
		.INIT('h2a)
	) name25409 (
		\m5_addr_i[13]_pad ,
		_w8865_,
		_w8866_,
		_w27310_
	);
	LUT4 #(
		.INIT('h5d7f)
	) name25410 (
		_w8860_,
		_w8863_,
		_w27309_,
		_w27310_,
		_w27311_
	);
	LUT3 #(
		.INIT('h80)
	) name25411 (
		\m2_addr_i[13]_pad ,
		_w8865_,
		_w8866_,
		_w27312_
	);
	LUT3 #(
		.INIT('h80)
	) name25412 (
		\m6_addr_i[13]_pad ,
		_w8865_,
		_w8866_,
		_w27313_
	);
	LUT4 #(
		.INIT('haebf)
	) name25413 (
		_w8860_,
		_w8863_,
		_w27312_,
		_w27313_,
		_w27314_
	);
	LUT3 #(
		.INIT('h2a)
	) name25414 (
		\m3_addr_i[13]_pad ,
		_w8865_,
		_w8866_,
		_w27315_
	);
	LUT3 #(
		.INIT('h80)
	) name25415 (
		\m4_addr_i[13]_pad ,
		_w8865_,
		_w8866_,
		_w27316_
	);
	LUT4 #(
		.INIT('h9dbf)
	) name25416 (
		_w8860_,
		_w8863_,
		_w27315_,
		_w27316_,
		_w27317_
	);
	LUT4 #(
		.INIT('h7fff)
	) name25417 (
		_w27308_,
		_w27311_,
		_w27314_,
		_w27317_,
		_w27318_
	);
	LUT3 #(
		.INIT('h80)
	) name25418 (
		\m6_addr_i[14]_pad ,
		_w8865_,
		_w8866_,
		_w27319_
	);
	LUT3 #(
		.INIT('h2a)
	) name25419 (
		\m5_addr_i[14]_pad ,
		_w8865_,
		_w8866_,
		_w27320_
	);
	LUT4 #(
		.INIT('hcdef)
	) name25420 (
		_w8860_,
		_w8863_,
		_w27319_,
		_w27320_,
		_w27321_
	);
	LUT3 #(
		.INIT('h2a)
	) name25421 (
		\m3_addr_i[14]_pad ,
		_w8865_,
		_w8866_,
		_w27322_
	);
	LUT3 #(
		.INIT('h2a)
	) name25422 (
		\m7_addr_i[14]_pad ,
		_w8865_,
		_w8866_,
		_w27323_
	);
	LUT4 #(
		.INIT('haebf)
	) name25423 (
		_w8860_,
		_w8863_,
		_w27322_,
		_w27323_,
		_w27324_
	);
	LUT3 #(
		.INIT('h80)
	) name25424 (
		\m4_addr_i[14]_pad ,
		_w8865_,
		_w8866_,
		_w27325_
	);
	LUT3 #(
		.INIT('h80)
	) name25425 (
		\m0_addr_i[14]_pad ,
		_w8865_,
		_w8866_,
		_w27326_
	);
	LUT4 #(
		.INIT('h57df)
	) name25426 (
		_w8860_,
		_w8863_,
		_w27325_,
		_w27326_,
		_w27327_
	);
	LUT3 #(
		.INIT('h2a)
	) name25427 (
		\m1_addr_i[14]_pad ,
		_w8865_,
		_w8866_,
		_w27328_
	);
	LUT3 #(
		.INIT('h80)
	) name25428 (
		\m2_addr_i[14]_pad ,
		_w8865_,
		_w8866_,
		_w27329_
	);
	LUT4 #(
		.INIT('h3b7f)
	) name25429 (
		_w8860_,
		_w8863_,
		_w27328_,
		_w27329_,
		_w27330_
	);
	LUT4 #(
		.INIT('h7fff)
	) name25430 (
		_w27321_,
		_w27324_,
		_w27327_,
		_w27330_,
		_w27331_
	);
	LUT3 #(
		.INIT('h2a)
	) name25431 (
		\m1_addr_i[15]_pad ,
		_w8865_,
		_w8866_,
		_w27332_
	);
	LUT3 #(
		.INIT('h80)
	) name25432 (
		\m2_addr_i[15]_pad ,
		_w8865_,
		_w8866_,
		_w27333_
	);
	LUT4 #(
		.INIT('h3b7f)
	) name25433 (
		_w8860_,
		_w8863_,
		_w27332_,
		_w27333_,
		_w27334_
	);
	LUT3 #(
		.INIT('h80)
	) name25434 (
		\m0_addr_i[15]_pad ,
		_w8865_,
		_w8866_,
		_w27335_
	);
	LUT3 #(
		.INIT('h80)
	) name25435 (
		\m4_addr_i[15]_pad ,
		_w8865_,
		_w8866_,
		_w27336_
	);
	LUT4 #(
		.INIT('h5d7f)
	) name25436 (
		_w8860_,
		_w8863_,
		_w27335_,
		_w27336_,
		_w27337_
	);
	LUT3 #(
		.INIT('h2a)
	) name25437 (
		\m7_addr_i[15]_pad ,
		_w8865_,
		_w8866_,
		_w27338_
	);
	LUT3 #(
		.INIT('h2a)
	) name25438 (
		\m3_addr_i[15]_pad ,
		_w8865_,
		_w8866_,
		_w27339_
	);
	LUT4 #(
		.INIT('habef)
	) name25439 (
		_w8860_,
		_w8863_,
		_w27338_,
		_w27339_,
		_w27340_
	);
	LUT3 #(
		.INIT('h80)
	) name25440 (
		\m6_addr_i[15]_pad ,
		_w8865_,
		_w8866_,
		_w27341_
	);
	LUT3 #(
		.INIT('h2a)
	) name25441 (
		\m5_addr_i[15]_pad ,
		_w8865_,
		_w8866_,
		_w27342_
	);
	LUT4 #(
		.INIT('hcdef)
	) name25442 (
		_w8860_,
		_w8863_,
		_w27341_,
		_w27342_,
		_w27343_
	);
	LUT4 #(
		.INIT('h7fff)
	) name25443 (
		_w27334_,
		_w27337_,
		_w27340_,
		_w27343_,
		_w27344_
	);
	LUT3 #(
		.INIT('h2a)
	) name25444 (
		\m1_addr_i[16]_pad ,
		_w8865_,
		_w8866_,
		_w27345_
	);
	LUT3 #(
		.INIT('h80)
	) name25445 (
		\m2_addr_i[16]_pad ,
		_w8865_,
		_w8866_,
		_w27346_
	);
	LUT4 #(
		.INIT('h3b7f)
	) name25446 (
		_w8860_,
		_w8863_,
		_w27345_,
		_w27346_,
		_w27347_
	);
	LUT3 #(
		.INIT('h80)
	) name25447 (
		\m0_addr_i[16]_pad ,
		_w8865_,
		_w8866_,
		_w27348_
	);
	LUT3 #(
		.INIT('h2a)
	) name25448 (
		\m5_addr_i[16]_pad ,
		_w8865_,
		_w8866_,
		_w27349_
	);
	LUT4 #(
		.INIT('h5d7f)
	) name25449 (
		_w8860_,
		_w8863_,
		_w27348_,
		_w27349_,
		_w27350_
	);
	LUT3 #(
		.INIT('h2a)
	) name25450 (
		\m7_addr_i[16]_pad ,
		_w8865_,
		_w8866_,
		_w27351_
	);
	LUT3 #(
		.INIT('h80)
	) name25451 (
		\m6_addr_i[16]_pad ,
		_w8865_,
		_w8866_,
		_w27352_
	);
	LUT3 #(
		.INIT('h57)
	) name25452 (
		_w8878_,
		_w27351_,
		_w27352_,
		_w27353_
	);
	LUT3 #(
		.INIT('h2a)
	) name25453 (
		\m3_addr_i[16]_pad ,
		_w8865_,
		_w8866_,
		_w27354_
	);
	LUT3 #(
		.INIT('h80)
	) name25454 (
		\m4_addr_i[16]_pad ,
		_w8865_,
		_w8866_,
		_w27355_
	);
	LUT4 #(
		.INIT('h9dbf)
	) name25455 (
		_w8860_,
		_w8863_,
		_w27354_,
		_w27355_,
		_w27356_
	);
	LUT4 #(
		.INIT('h7fff)
	) name25456 (
		_w27347_,
		_w27350_,
		_w27353_,
		_w27356_,
		_w27357_
	);
	LUT3 #(
		.INIT('h2a)
	) name25457 (
		\m1_addr_i[17]_pad ,
		_w8865_,
		_w8866_,
		_w27358_
	);
	LUT3 #(
		.INIT('h80)
	) name25458 (
		\m2_addr_i[17]_pad ,
		_w8865_,
		_w8866_,
		_w27359_
	);
	LUT4 #(
		.INIT('h3b7f)
	) name25459 (
		_w8860_,
		_w8863_,
		_w27358_,
		_w27359_,
		_w27360_
	);
	LUT3 #(
		.INIT('h80)
	) name25460 (
		\m0_addr_i[17]_pad ,
		_w8865_,
		_w8866_,
		_w27361_
	);
	LUT3 #(
		.INIT('h2a)
	) name25461 (
		\m5_addr_i[17]_pad ,
		_w8865_,
		_w8866_,
		_w27362_
	);
	LUT4 #(
		.INIT('h5d7f)
	) name25462 (
		_w8860_,
		_w8863_,
		_w27361_,
		_w27362_,
		_w27363_
	);
	LUT3 #(
		.INIT('h2a)
	) name25463 (
		\m7_addr_i[17]_pad ,
		_w8865_,
		_w8866_,
		_w27364_
	);
	LUT3 #(
		.INIT('h80)
	) name25464 (
		\m6_addr_i[17]_pad ,
		_w8865_,
		_w8866_,
		_w27365_
	);
	LUT3 #(
		.INIT('h57)
	) name25465 (
		_w8878_,
		_w27364_,
		_w27365_,
		_w27366_
	);
	LUT3 #(
		.INIT('h2a)
	) name25466 (
		\m3_addr_i[17]_pad ,
		_w8865_,
		_w8866_,
		_w27367_
	);
	LUT3 #(
		.INIT('h80)
	) name25467 (
		\m4_addr_i[17]_pad ,
		_w8865_,
		_w8866_,
		_w27368_
	);
	LUT4 #(
		.INIT('h9dbf)
	) name25468 (
		_w8860_,
		_w8863_,
		_w27367_,
		_w27368_,
		_w27369_
	);
	LUT4 #(
		.INIT('h7fff)
	) name25469 (
		_w27360_,
		_w27363_,
		_w27366_,
		_w27369_,
		_w27370_
	);
	LUT3 #(
		.INIT('h80)
	) name25470 (
		\m6_addr_i[18]_pad ,
		_w8865_,
		_w8866_,
		_w27371_
	);
	LUT3 #(
		.INIT('h2a)
	) name25471 (
		\m5_addr_i[18]_pad ,
		_w8865_,
		_w8866_,
		_w27372_
	);
	LUT4 #(
		.INIT('hcdef)
	) name25472 (
		_w8860_,
		_w8863_,
		_w27371_,
		_w27372_,
		_w27373_
	);
	LUT3 #(
		.INIT('h2a)
	) name25473 (
		\m1_addr_i[18]_pad ,
		_w8865_,
		_w8866_,
		_w27374_
	);
	LUT3 #(
		.INIT('h80)
	) name25474 (
		\m4_addr_i[18]_pad ,
		_w8865_,
		_w8866_,
		_w27375_
	);
	LUT4 #(
		.INIT('h5d7f)
	) name25475 (
		_w8860_,
		_w8863_,
		_w27374_,
		_w27375_,
		_w27376_
	);
	LUT3 #(
		.INIT('h80)
	) name25476 (
		\m2_addr_i[18]_pad ,
		_w8865_,
		_w8866_,
		_w27377_
	);
	LUT3 #(
		.INIT('h2a)
	) name25477 (
		\m3_addr_i[18]_pad ,
		_w8865_,
		_w8866_,
		_w27378_
	);
	LUT3 #(
		.INIT('h57)
	) name25478 (
		_w8864_,
		_w27377_,
		_w27378_,
		_w27379_
	);
	LUT3 #(
		.INIT('h80)
	) name25479 (
		\m0_addr_i[18]_pad ,
		_w8865_,
		_w8866_,
		_w27380_
	);
	LUT3 #(
		.INIT('h2a)
	) name25480 (
		\m7_addr_i[18]_pad ,
		_w8865_,
		_w8866_,
		_w27381_
	);
	LUT4 #(
		.INIT('h6e7f)
	) name25481 (
		_w8860_,
		_w8863_,
		_w27380_,
		_w27381_,
		_w27382_
	);
	LUT4 #(
		.INIT('h7fff)
	) name25482 (
		_w27373_,
		_w27376_,
		_w27379_,
		_w27382_,
		_w27383_
	);
	LUT3 #(
		.INIT('h2a)
	) name25483 (
		\m3_addr_i[19]_pad ,
		_w8865_,
		_w8866_,
		_w27384_
	);
	LUT3 #(
		.INIT('h80)
	) name25484 (
		\m4_addr_i[19]_pad ,
		_w8865_,
		_w8866_,
		_w27385_
	);
	LUT4 #(
		.INIT('h9dbf)
	) name25485 (
		_w8860_,
		_w8863_,
		_w27384_,
		_w27385_,
		_w27386_
	);
	LUT3 #(
		.INIT('h80)
	) name25486 (
		\m0_addr_i[19]_pad ,
		_w8865_,
		_w8866_,
		_w27387_
	);
	LUT3 #(
		.INIT('h2a)
	) name25487 (
		\m5_addr_i[19]_pad ,
		_w8865_,
		_w8866_,
		_w27388_
	);
	LUT4 #(
		.INIT('h5d7f)
	) name25488 (
		_w8860_,
		_w8863_,
		_w27387_,
		_w27388_,
		_w27389_
	);
	LUT3 #(
		.INIT('h2a)
	) name25489 (
		\m7_addr_i[19]_pad ,
		_w8865_,
		_w8866_,
		_w27390_
	);
	LUT3 #(
		.INIT('h80)
	) name25490 (
		\m6_addr_i[19]_pad ,
		_w8865_,
		_w8866_,
		_w27391_
	);
	LUT3 #(
		.INIT('h57)
	) name25491 (
		_w8878_,
		_w27390_,
		_w27391_,
		_w27392_
	);
	LUT3 #(
		.INIT('h2a)
	) name25492 (
		\m1_addr_i[19]_pad ,
		_w8865_,
		_w8866_,
		_w27393_
	);
	LUT3 #(
		.INIT('h80)
	) name25493 (
		\m2_addr_i[19]_pad ,
		_w8865_,
		_w8866_,
		_w27394_
	);
	LUT4 #(
		.INIT('h3b7f)
	) name25494 (
		_w8860_,
		_w8863_,
		_w27393_,
		_w27394_,
		_w27395_
	);
	LUT4 #(
		.INIT('h7fff)
	) name25495 (
		_w27386_,
		_w27389_,
		_w27392_,
		_w27395_,
		_w27396_
	);
	LUT3 #(
		.INIT('h2a)
	) name25496 (
		\m3_addr_i[1]_pad ,
		_w8865_,
		_w8866_,
		_w27397_
	);
	LUT3 #(
		.INIT('h80)
	) name25497 (
		\m4_addr_i[1]_pad ,
		_w8865_,
		_w8866_,
		_w27398_
	);
	LUT4 #(
		.INIT('h9dbf)
	) name25498 (
		_w8860_,
		_w8863_,
		_w27397_,
		_w27398_,
		_w27399_
	);
	LUT3 #(
		.INIT('h80)
	) name25499 (
		\m6_addr_i[1]_pad ,
		_w8865_,
		_w8866_,
		_w27400_
	);
	LUT3 #(
		.INIT('h80)
	) name25500 (
		\m2_addr_i[1]_pad ,
		_w8865_,
		_w8866_,
		_w27401_
	);
	LUT4 #(
		.INIT('habef)
	) name25501 (
		_w8860_,
		_w8863_,
		_w27400_,
		_w27401_,
		_w27402_
	);
	LUT3 #(
		.INIT('h2a)
	) name25502 (
		\m5_addr_i[1]_pad ,
		_w8865_,
		_w8866_,
		_w27403_
	);
	LUT3 #(
		.INIT('h2a)
	) name25503 (
		\m1_addr_i[1]_pad ,
		_w8865_,
		_w8866_,
		_w27404_
	);
	LUT4 #(
		.INIT('h57df)
	) name25504 (
		_w8860_,
		_w8863_,
		_w27403_,
		_w27404_,
		_w27405_
	);
	LUT3 #(
		.INIT('h80)
	) name25505 (
		\m0_addr_i[1]_pad ,
		_w8865_,
		_w8866_,
		_w27406_
	);
	LUT3 #(
		.INIT('h2a)
	) name25506 (
		\m7_addr_i[1]_pad ,
		_w8865_,
		_w8866_,
		_w27407_
	);
	LUT4 #(
		.INIT('h6e7f)
	) name25507 (
		_w8860_,
		_w8863_,
		_w27406_,
		_w27407_,
		_w27408_
	);
	LUT4 #(
		.INIT('h7fff)
	) name25508 (
		_w27399_,
		_w27402_,
		_w27405_,
		_w27408_,
		_w27409_
	);
	LUT3 #(
		.INIT('h80)
	) name25509 (
		\m0_addr_i[20]_pad ,
		_w8865_,
		_w8866_,
		_w27410_
	);
	LUT3 #(
		.INIT('h2a)
	) name25510 (
		\m7_addr_i[20]_pad ,
		_w8865_,
		_w8866_,
		_w27411_
	);
	LUT4 #(
		.INIT('h6e7f)
	) name25511 (
		_w8860_,
		_w8863_,
		_w27410_,
		_w27411_,
		_w27412_
	);
	LUT3 #(
		.INIT('h2a)
	) name25512 (
		\m1_addr_i[20]_pad ,
		_w8865_,
		_w8866_,
		_w27413_
	);
	LUT3 #(
		.INIT('h2a)
	) name25513 (
		\m5_addr_i[20]_pad ,
		_w8865_,
		_w8866_,
		_w27414_
	);
	LUT4 #(
		.INIT('h5d7f)
	) name25514 (
		_w8860_,
		_w8863_,
		_w27413_,
		_w27414_,
		_w27415_
	);
	LUT3 #(
		.INIT('h80)
	) name25515 (
		\m2_addr_i[20]_pad ,
		_w8865_,
		_w8866_,
		_w27416_
	);
	LUT3 #(
		.INIT('h80)
	) name25516 (
		\m6_addr_i[20]_pad ,
		_w8865_,
		_w8866_,
		_w27417_
	);
	LUT4 #(
		.INIT('haebf)
	) name25517 (
		_w8860_,
		_w8863_,
		_w27416_,
		_w27417_,
		_w27418_
	);
	LUT3 #(
		.INIT('h2a)
	) name25518 (
		\m3_addr_i[20]_pad ,
		_w8865_,
		_w8866_,
		_w27419_
	);
	LUT3 #(
		.INIT('h80)
	) name25519 (
		\m4_addr_i[20]_pad ,
		_w8865_,
		_w8866_,
		_w27420_
	);
	LUT4 #(
		.INIT('h9dbf)
	) name25520 (
		_w8860_,
		_w8863_,
		_w27419_,
		_w27420_,
		_w27421_
	);
	LUT4 #(
		.INIT('h7fff)
	) name25521 (
		_w27412_,
		_w27415_,
		_w27418_,
		_w27421_,
		_w27422_
	);
	LUT3 #(
		.INIT('h80)
	) name25522 (
		\m6_addr_i[21]_pad ,
		_w8865_,
		_w8866_,
		_w27423_
	);
	LUT3 #(
		.INIT('h2a)
	) name25523 (
		\m5_addr_i[21]_pad ,
		_w8865_,
		_w8866_,
		_w27424_
	);
	LUT4 #(
		.INIT('hcdef)
	) name25524 (
		_w8860_,
		_w8863_,
		_w27423_,
		_w27424_,
		_w27425_
	);
	LUT3 #(
		.INIT('h2a)
	) name25525 (
		\m3_addr_i[21]_pad ,
		_w8865_,
		_w8866_,
		_w27426_
	);
	LUT3 #(
		.INIT('h80)
	) name25526 (
		\m2_addr_i[21]_pad ,
		_w8865_,
		_w8866_,
		_w27427_
	);
	LUT3 #(
		.INIT('h57)
	) name25527 (
		_w8864_,
		_w27426_,
		_w27427_,
		_w27428_
	);
	LUT3 #(
		.INIT('h80)
	) name25528 (
		\m4_addr_i[21]_pad ,
		_w8865_,
		_w8866_,
		_w27429_
	);
	LUT3 #(
		.INIT('h2a)
	) name25529 (
		\m1_addr_i[21]_pad ,
		_w8865_,
		_w8866_,
		_w27430_
	);
	LUT4 #(
		.INIT('h57df)
	) name25530 (
		_w8860_,
		_w8863_,
		_w27429_,
		_w27430_,
		_w27431_
	);
	LUT3 #(
		.INIT('h80)
	) name25531 (
		\m0_addr_i[21]_pad ,
		_w8865_,
		_w8866_,
		_w27432_
	);
	LUT3 #(
		.INIT('h2a)
	) name25532 (
		\m7_addr_i[21]_pad ,
		_w8865_,
		_w8866_,
		_w27433_
	);
	LUT4 #(
		.INIT('h6e7f)
	) name25533 (
		_w8860_,
		_w8863_,
		_w27432_,
		_w27433_,
		_w27434_
	);
	LUT4 #(
		.INIT('h7fff)
	) name25534 (
		_w27425_,
		_w27428_,
		_w27431_,
		_w27434_,
		_w27435_
	);
	LUT3 #(
		.INIT('h2a)
	) name25535 (
		\m1_addr_i[22]_pad ,
		_w8865_,
		_w8866_,
		_w27436_
	);
	LUT3 #(
		.INIT('h80)
	) name25536 (
		\m2_addr_i[22]_pad ,
		_w8865_,
		_w8866_,
		_w27437_
	);
	LUT4 #(
		.INIT('h3b7f)
	) name25537 (
		_w8860_,
		_w8863_,
		_w27436_,
		_w27437_,
		_w27438_
	);
	LUT3 #(
		.INIT('h80)
	) name25538 (
		\m0_addr_i[22]_pad ,
		_w8865_,
		_w8866_,
		_w27439_
	);
	LUT3 #(
		.INIT('h2a)
	) name25539 (
		\m5_addr_i[22]_pad ,
		_w8865_,
		_w8866_,
		_w27440_
	);
	LUT4 #(
		.INIT('h5d7f)
	) name25540 (
		_w8860_,
		_w8863_,
		_w27439_,
		_w27440_,
		_w27441_
	);
	LUT3 #(
		.INIT('h2a)
	) name25541 (
		\m7_addr_i[22]_pad ,
		_w8865_,
		_w8866_,
		_w27442_
	);
	LUT3 #(
		.INIT('h80)
	) name25542 (
		\m6_addr_i[22]_pad ,
		_w8865_,
		_w8866_,
		_w27443_
	);
	LUT3 #(
		.INIT('h57)
	) name25543 (
		_w8878_,
		_w27442_,
		_w27443_,
		_w27444_
	);
	LUT3 #(
		.INIT('h2a)
	) name25544 (
		\m3_addr_i[22]_pad ,
		_w8865_,
		_w8866_,
		_w27445_
	);
	LUT3 #(
		.INIT('h80)
	) name25545 (
		\m4_addr_i[22]_pad ,
		_w8865_,
		_w8866_,
		_w27446_
	);
	LUT4 #(
		.INIT('h9dbf)
	) name25546 (
		_w8860_,
		_w8863_,
		_w27445_,
		_w27446_,
		_w27447_
	);
	LUT4 #(
		.INIT('h7fff)
	) name25547 (
		_w27438_,
		_w27441_,
		_w27444_,
		_w27447_,
		_w27448_
	);
	LUT3 #(
		.INIT('h80)
	) name25548 (
		\m6_addr_i[23]_pad ,
		_w8865_,
		_w8866_,
		_w27449_
	);
	LUT3 #(
		.INIT('h2a)
	) name25549 (
		\m5_addr_i[23]_pad ,
		_w8865_,
		_w8866_,
		_w27450_
	);
	LUT4 #(
		.INIT('hcdef)
	) name25550 (
		_w8860_,
		_w8863_,
		_w27449_,
		_w27450_,
		_w27451_
	);
	LUT3 #(
		.INIT('h2a)
	) name25551 (
		\m3_addr_i[23]_pad ,
		_w8865_,
		_w8866_,
		_w27452_
	);
	LUT3 #(
		.INIT('h2a)
	) name25552 (
		\m7_addr_i[23]_pad ,
		_w8865_,
		_w8866_,
		_w27453_
	);
	LUT4 #(
		.INIT('haebf)
	) name25553 (
		_w8860_,
		_w8863_,
		_w27452_,
		_w27453_,
		_w27454_
	);
	LUT3 #(
		.INIT('h80)
	) name25554 (
		\m4_addr_i[23]_pad ,
		_w8865_,
		_w8866_,
		_w27455_
	);
	LUT3 #(
		.INIT('h80)
	) name25555 (
		\m0_addr_i[23]_pad ,
		_w8865_,
		_w8866_,
		_w27456_
	);
	LUT4 #(
		.INIT('h57df)
	) name25556 (
		_w8860_,
		_w8863_,
		_w27455_,
		_w27456_,
		_w27457_
	);
	LUT3 #(
		.INIT('h2a)
	) name25557 (
		\m1_addr_i[23]_pad ,
		_w8865_,
		_w8866_,
		_w27458_
	);
	LUT3 #(
		.INIT('h80)
	) name25558 (
		\m2_addr_i[23]_pad ,
		_w8865_,
		_w8866_,
		_w27459_
	);
	LUT4 #(
		.INIT('h3b7f)
	) name25559 (
		_w8860_,
		_w8863_,
		_w27458_,
		_w27459_,
		_w27460_
	);
	LUT4 #(
		.INIT('h7fff)
	) name25560 (
		_w27451_,
		_w27454_,
		_w27457_,
		_w27460_,
		_w27461_
	);
	LUT3 #(
		.INIT('h80)
	) name25561 (
		\m0_addr_i[24]_pad ,
		_w8865_,
		_w8866_,
		_w27462_
	);
	LUT3 #(
		.INIT('h2a)
	) name25562 (
		\m7_addr_i[24]_pad ,
		_w8865_,
		_w8866_,
		_w27463_
	);
	LUT4 #(
		.INIT('h6e7f)
	) name25563 (
		_w8860_,
		_w8863_,
		_w27462_,
		_w27463_,
		_w27464_
	);
	LUT3 #(
		.INIT('h2a)
	) name25564 (
		\m1_addr_i[24]_pad ,
		_w8865_,
		_w8866_,
		_w27465_
	);
	LUT3 #(
		.INIT('h80)
	) name25565 (
		\m6_addr_i[24]_pad ,
		_w8865_,
		_w8866_,
		_w27466_
	);
	LUT4 #(
		.INIT('h6e7f)
	) name25566 (
		_w8860_,
		_w8863_,
		_w27465_,
		_w27466_,
		_w27467_
	);
	LUT3 #(
		.INIT('h80)
	) name25567 (
		\m2_addr_i[24]_pad ,
		_w8865_,
		_w8866_,
		_w27468_
	);
	LUT3 #(
		.INIT('h2a)
	) name25568 (
		\m5_addr_i[24]_pad ,
		_w8865_,
		_w8866_,
		_w27469_
	);
	LUT4 #(
		.INIT('h9dbf)
	) name25569 (
		_w8860_,
		_w8863_,
		_w27468_,
		_w27469_,
		_w27470_
	);
	LUT3 #(
		.INIT('h2a)
	) name25570 (
		\m3_addr_i[24]_pad ,
		_w8865_,
		_w8866_,
		_w27471_
	);
	LUT3 #(
		.INIT('h80)
	) name25571 (
		\m4_addr_i[24]_pad ,
		_w8865_,
		_w8866_,
		_w27472_
	);
	LUT4 #(
		.INIT('h9dbf)
	) name25572 (
		_w8860_,
		_w8863_,
		_w27471_,
		_w27472_,
		_w27473_
	);
	LUT4 #(
		.INIT('h7fff)
	) name25573 (
		_w27464_,
		_w27467_,
		_w27470_,
		_w27473_,
		_w27474_
	);
	LUT3 #(
		.INIT('h80)
	) name25574 (
		\m0_addr_i[25]_pad ,
		_w8865_,
		_w8866_,
		_w27475_
	);
	LUT3 #(
		.INIT('h2a)
	) name25575 (
		\m7_addr_i[25]_pad ,
		_w8865_,
		_w8866_,
		_w27476_
	);
	LUT4 #(
		.INIT('h6e7f)
	) name25576 (
		_w8860_,
		_w8863_,
		_w27475_,
		_w27476_,
		_w27477_
	);
	LUT3 #(
		.INIT('h2a)
	) name25577 (
		\m5_addr_i[25]_pad ,
		_w8865_,
		_w8866_,
		_w27478_
	);
	LUT3 #(
		.INIT('h80)
	) name25578 (
		\m2_addr_i[25]_pad ,
		_w8865_,
		_w8866_,
		_w27479_
	);
	LUT4 #(
		.INIT('h9bdf)
	) name25579 (
		_w8860_,
		_w8863_,
		_w27478_,
		_w27479_,
		_w27480_
	);
	LUT3 #(
		.INIT('h80)
	) name25580 (
		\m6_addr_i[25]_pad ,
		_w8865_,
		_w8866_,
		_w27481_
	);
	LUT3 #(
		.INIT('h2a)
	) name25581 (
		\m1_addr_i[25]_pad ,
		_w8865_,
		_w8866_,
		_w27482_
	);
	LUT4 #(
		.INIT('h67ef)
	) name25582 (
		_w8860_,
		_w8863_,
		_w27481_,
		_w27482_,
		_w27483_
	);
	LUT3 #(
		.INIT('h2a)
	) name25583 (
		\m3_addr_i[25]_pad ,
		_w8865_,
		_w8866_,
		_w27484_
	);
	LUT3 #(
		.INIT('h80)
	) name25584 (
		\m4_addr_i[25]_pad ,
		_w8865_,
		_w8866_,
		_w27485_
	);
	LUT4 #(
		.INIT('h9dbf)
	) name25585 (
		_w8860_,
		_w8863_,
		_w27484_,
		_w27485_,
		_w27486_
	);
	LUT4 #(
		.INIT('h7fff)
	) name25586 (
		_w27477_,
		_w27480_,
		_w27483_,
		_w27486_,
		_w27487_
	);
	LUT3 #(
		.INIT('h2a)
	) name25587 (
		\m1_addr_i[26]_pad ,
		_w8865_,
		_w8866_,
		_w27488_
	);
	LUT3 #(
		.INIT('h80)
	) name25588 (
		\m2_addr_i[26]_pad ,
		_w8865_,
		_w8866_,
		_w27489_
	);
	LUT4 #(
		.INIT('h3b7f)
	) name25589 (
		_w8860_,
		_w8863_,
		_w27488_,
		_w27489_,
		_w27490_
	);
	LUT3 #(
		.INIT('h2a)
	) name25590 (
		\m5_addr_i[26]_pad ,
		_w8865_,
		_w8866_,
		_w27491_
	);
	LUT3 #(
		.INIT('h2a)
	) name25591 (
		\m7_addr_i[26]_pad ,
		_w8865_,
		_w8866_,
		_w27492_
	);
	LUT4 #(
		.INIT('hcedf)
	) name25592 (
		_w8860_,
		_w8863_,
		_w27491_,
		_w27492_,
		_w27493_
	);
	LUT3 #(
		.INIT('h80)
	) name25593 (
		\m6_addr_i[26]_pad ,
		_w8865_,
		_w8866_,
		_w27494_
	);
	LUT3 #(
		.INIT('h80)
	) name25594 (
		\m0_addr_i[26]_pad ,
		_w8865_,
		_w8866_,
		_w27495_
	);
	LUT4 #(
		.INIT('h67ef)
	) name25595 (
		_w8860_,
		_w8863_,
		_w27494_,
		_w27495_,
		_w27496_
	);
	LUT3 #(
		.INIT('h2a)
	) name25596 (
		\m3_addr_i[26]_pad ,
		_w8865_,
		_w8866_,
		_w27497_
	);
	LUT3 #(
		.INIT('h80)
	) name25597 (
		\m4_addr_i[26]_pad ,
		_w8865_,
		_w8866_,
		_w27498_
	);
	LUT4 #(
		.INIT('h9dbf)
	) name25598 (
		_w8860_,
		_w8863_,
		_w27497_,
		_w27498_,
		_w27499_
	);
	LUT4 #(
		.INIT('h7fff)
	) name25599 (
		_w27490_,
		_w27493_,
		_w27496_,
		_w27499_,
		_w27500_
	);
	LUT3 #(
		.INIT('h2a)
	) name25600 (
		\m1_addr_i[27]_pad ,
		_w8865_,
		_w8866_,
		_w27501_
	);
	LUT3 #(
		.INIT('h80)
	) name25601 (
		\m2_addr_i[27]_pad ,
		_w8865_,
		_w8866_,
		_w27502_
	);
	LUT4 #(
		.INIT('h3b7f)
	) name25602 (
		_w8860_,
		_w8863_,
		_w27501_,
		_w27502_,
		_w27503_
	);
	LUT3 #(
		.INIT('h2a)
	) name25603 (
		\m3_addr_i[27]_pad ,
		_w8865_,
		_w8866_,
		_w27504_
	);
	LUT3 #(
		.INIT('h2a)
	) name25604 (
		\m7_addr_i[27]_pad ,
		_w8865_,
		_w8866_,
		_w27505_
	);
	LUT4 #(
		.INIT('haebf)
	) name25605 (
		_w8860_,
		_w8863_,
		_w27504_,
		_w27505_,
		_w27506_
	);
	LUT3 #(
		.INIT('h80)
	) name25606 (
		\m4_addr_i[27]_pad ,
		_w8865_,
		_w8866_,
		_w27507_
	);
	LUT3 #(
		.INIT('h80)
	) name25607 (
		\m0_addr_i[27]_pad ,
		_w8865_,
		_w8866_,
		_w27508_
	);
	LUT4 #(
		.INIT('h57df)
	) name25608 (
		_w8860_,
		_w8863_,
		_w27507_,
		_w27508_,
		_w27509_
	);
	LUT3 #(
		.INIT('h2a)
	) name25609 (
		\m5_addr_i[27]_pad ,
		_w8865_,
		_w8866_,
		_w27510_
	);
	LUT3 #(
		.INIT('h80)
	) name25610 (
		\m6_addr_i[27]_pad ,
		_w8865_,
		_w8866_,
		_w27511_
	);
	LUT4 #(
		.INIT('hcedf)
	) name25611 (
		_w8860_,
		_w8863_,
		_w27510_,
		_w27511_,
		_w27512_
	);
	LUT4 #(
		.INIT('h7fff)
	) name25612 (
		_w27503_,
		_w27506_,
		_w27509_,
		_w27512_,
		_w27513_
	);
	LUT3 #(
		.INIT('h2a)
	) name25613 (
		\m5_addr_i[28]_pad ,
		_w8865_,
		_w8866_,
		_w27514_
	);
	LUT3 #(
		.INIT('h80)
	) name25614 (
		\m6_addr_i[28]_pad ,
		_w8865_,
		_w8866_,
		_w27515_
	);
	LUT4 #(
		.INIT('hcedf)
	) name25615 (
		_w8860_,
		_w8863_,
		_w27514_,
		_w27515_,
		_w27516_
	);
	LUT3 #(
		.INIT('h2a)
	) name25616 (
		\m3_addr_i[28]_pad ,
		_w8865_,
		_w8866_,
		_w27517_
	);
	LUT3 #(
		.INIT('h80)
	) name25617 (
		\m2_addr_i[28]_pad ,
		_w8865_,
		_w8866_,
		_w27518_
	);
	LUT3 #(
		.INIT('h57)
	) name25618 (
		_w8864_,
		_w27517_,
		_w27518_,
		_w27519_
	);
	LUT3 #(
		.INIT('h80)
	) name25619 (
		\m4_addr_i[28]_pad ,
		_w8865_,
		_w8866_,
		_w27520_
	);
	LUT3 #(
		.INIT('h2a)
	) name25620 (
		\m1_addr_i[28]_pad ,
		_w8865_,
		_w8866_,
		_w27521_
	);
	LUT4 #(
		.INIT('h57df)
	) name25621 (
		_w8860_,
		_w8863_,
		_w27520_,
		_w27521_,
		_w27522_
	);
	LUT3 #(
		.INIT('h80)
	) name25622 (
		\m0_addr_i[28]_pad ,
		_w8865_,
		_w8866_,
		_w27523_
	);
	LUT3 #(
		.INIT('h2a)
	) name25623 (
		\m7_addr_i[28]_pad ,
		_w8865_,
		_w8866_,
		_w27524_
	);
	LUT4 #(
		.INIT('h6e7f)
	) name25624 (
		_w8860_,
		_w8863_,
		_w27523_,
		_w27524_,
		_w27525_
	);
	LUT4 #(
		.INIT('h7fff)
	) name25625 (
		_w27516_,
		_w27519_,
		_w27522_,
		_w27525_,
		_w27526_
	);
	LUT3 #(
		.INIT('h2a)
	) name25626 (
		\m1_addr_i[29]_pad ,
		_w8865_,
		_w8866_,
		_w27527_
	);
	LUT3 #(
		.INIT('h80)
	) name25627 (
		\m2_addr_i[29]_pad ,
		_w8865_,
		_w8866_,
		_w27528_
	);
	LUT4 #(
		.INIT('h3b7f)
	) name25628 (
		_w8860_,
		_w8863_,
		_w27527_,
		_w27528_,
		_w27529_
	);
	LUT3 #(
		.INIT('h2a)
	) name25629 (
		\m5_addr_i[29]_pad ,
		_w8865_,
		_w8866_,
		_w27530_
	);
	LUT3 #(
		.INIT('h2a)
	) name25630 (
		\m7_addr_i[29]_pad ,
		_w8865_,
		_w8866_,
		_w27531_
	);
	LUT4 #(
		.INIT('hcedf)
	) name25631 (
		_w8860_,
		_w8863_,
		_w27530_,
		_w27531_,
		_w27532_
	);
	LUT3 #(
		.INIT('h80)
	) name25632 (
		\m6_addr_i[29]_pad ,
		_w8865_,
		_w8866_,
		_w27533_
	);
	LUT3 #(
		.INIT('h80)
	) name25633 (
		\m0_addr_i[29]_pad ,
		_w8865_,
		_w8866_,
		_w27534_
	);
	LUT4 #(
		.INIT('h67ef)
	) name25634 (
		_w8860_,
		_w8863_,
		_w27533_,
		_w27534_,
		_w27535_
	);
	LUT3 #(
		.INIT('h2a)
	) name25635 (
		\m3_addr_i[29]_pad ,
		_w8865_,
		_w8866_,
		_w27536_
	);
	LUT3 #(
		.INIT('h80)
	) name25636 (
		\m4_addr_i[29]_pad ,
		_w8865_,
		_w8866_,
		_w27537_
	);
	LUT4 #(
		.INIT('h9dbf)
	) name25637 (
		_w8860_,
		_w8863_,
		_w27536_,
		_w27537_,
		_w27538_
	);
	LUT4 #(
		.INIT('h7fff)
	) name25638 (
		_w27529_,
		_w27532_,
		_w27535_,
		_w27538_,
		_w27539_
	);
	LUT3 #(
		.INIT('h2a)
	) name25639 (
		\m3_addr_i[2]_pad ,
		_w8865_,
		_w8866_,
		_w27540_
	);
	LUT3 #(
		.INIT('h80)
	) name25640 (
		\m4_addr_i[2]_pad ,
		_w8865_,
		_w8866_,
		_w27541_
	);
	LUT4 #(
		.INIT('h9dbf)
	) name25641 (
		_w8860_,
		_w8863_,
		_w27540_,
		_w27541_,
		_w27542_
	);
	LUT3 #(
		.INIT('h80)
	) name25642 (
		\m6_addr_i[2]_pad ,
		_w8865_,
		_w8866_,
		_w27543_
	);
	LUT3 #(
		.INIT('h2a)
	) name25643 (
		\m7_addr_i[2]_pad ,
		_w8865_,
		_w8866_,
		_w27544_
	);
	LUT3 #(
		.INIT('h57)
	) name25644 (
		_w8878_,
		_w27543_,
		_w27544_,
		_w27545_
	);
	LUT3 #(
		.INIT('h2a)
	) name25645 (
		\m5_addr_i[2]_pad ,
		_w8865_,
		_w8866_,
		_w27546_
	);
	LUT3 #(
		.INIT('h80)
	) name25646 (
		\m0_addr_i[2]_pad ,
		_w8865_,
		_w8866_,
		_w27547_
	);
	LUT4 #(
		.INIT('h57df)
	) name25647 (
		_w8860_,
		_w8863_,
		_w27546_,
		_w27547_,
		_w27548_
	);
	LUT3 #(
		.INIT('h2a)
	) name25648 (
		\m1_addr_i[2]_pad ,
		_w8865_,
		_w8866_,
		_w27549_
	);
	LUT3 #(
		.INIT('h80)
	) name25649 (
		\m2_addr_i[2]_pad ,
		_w8865_,
		_w8866_,
		_w27550_
	);
	LUT4 #(
		.INIT('h3b7f)
	) name25650 (
		_w8860_,
		_w8863_,
		_w27549_,
		_w27550_,
		_w27551_
	);
	LUT4 #(
		.INIT('h7fff)
	) name25651 (
		_w27542_,
		_w27545_,
		_w27548_,
		_w27551_,
		_w27552_
	);
	LUT3 #(
		.INIT('h80)
	) name25652 (
		\m0_addr_i[30]_pad ,
		_w8865_,
		_w8866_,
		_w27553_
	);
	LUT3 #(
		.INIT('h2a)
	) name25653 (
		\m7_addr_i[30]_pad ,
		_w8865_,
		_w8866_,
		_w27554_
	);
	LUT4 #(
		.INIT('h6e7f)
	) name25654 (
		_w8860_,
		_w8863_,
		_w27553_,
		_w27554_,
		_w27555_
	);
	LUT3 #(
		.INIT('h2a)
	) name25655 (
		\m3_addr_i[30]_pad ,
		_w8865_,
		_w8866_,
		_w27556_
	);
	LUT3 #(
		.INIT('h80)
	) name25656 (
		\m6_addr_i[30]_pad ,
		_w8865_,
		_w8866_,
		_w27557_
	);
	LUT4 #(
		.INIT('haebf)
	) name25657 (
		_w8860_,
		_w8863_,
		_w27556_,
		_w27557_,
		_w27558_
	);
	LUT3 #(
		.INIT('h80)
	) name25658 (
		\m4_addr_i[30]_pad ,
		_w8865_,
		_w8866_,
		_w27559_
	);
	LUT3 #(
		.INIT('h2a)
	) name25659 (
		\m5_addr_i[30]_pad ,
		_w8865_,
		_w8866_,
		_w27560_
	);
	LUT3 #(
		.INIT('h57)
	) name25660 (
		_w8884_,
		_w27559_,
		_w27560_,
		_w27561_
	);
	LUT3 #(
		.INIT('h2a)
	) name25661 (
		\m1_addr_i[30]_pad ,
		_w8865_,
		_w8866_,
		_w27562_
	);
	LUT3 #(
		.INIT('h80)
	) name25662 (
		\m2_addr_i[30]_pad ,
		_w8865_,
		_w8866_,
		_w27563_
	);
	LUT4 #(
		.INIT('h3b7f)
	) name25663 (
		_w8860_,
		_w8863_,
		_w27562_,
		_w27563_,
		_w27564_
	);
	LUT4 #(
		.INIT('h7fff)
	) name25664 (
		_w27555_,
		_w27558_,
		_w27561_,
		_w27564_,
		_w27565_
	);
	LUT3 #(
		.INIT('h2a)
	) name25665 (
		\m1_addr_i[31]_pad ,
		_w8865_,
		_w8866_,
		_w27566_
	);
	LUT3 #(
		.INIT('h80)
	) name25666 (
		\m2_addr_i[31]_pad ,
		_w8865_,
		_w8866_,
		_w27567_
	);
	LUT4 #(
		.INIT('h3b7f)
	) name25667 (
		_w8860_,
		_w8863_,
		_w27566_,
		_w27567_,
		_w27568_
	);
	LUT3 #(
		.INIT('h80)
	) name25668 (
		\m0_addr_i[31]_pad ,
		_w8865_,
		_w8866_,
		_w27569_
	);
	LUT3 #(
		.INIT('h80)
	) name25669 (
		\m4_addr_i[31]_pad ,
		_w8865_,
		_w8866_,
		_w27570_
	);
	LUT4 #(
		.INIT('h5d7f)
	) name25670 (
		_w8860_,
		_w8863_,
		_w27569_,
		_w27570_,
		_w27571_
	);
	LUT3 #(
		.INIT('h2a)
	) name25671 (
		\m7_addr_i[31]_pad ,
		_w8865_,
		_w8866_,
		_w27572_
	);
	LUT3 #(
		.INIT('h2a)
	) name25672 (
		\m3_addr_i[31]_pad ,
		_w8865_,
		_w8866_,
		_w27573_
	);
	LUT4 #(
		.INIT('habef)
	) name25673 (
		_w8860_,
		_w8863_,
		_w27572_,
		_w27573_,
		_w27574_
	);
	LUT3 #(
		.INIT('h2a)
	) name25674 (
		\m5_addr_i[31]_pad ,
		_w8865_,
		_w8866_,
		_w27575_
	);
	LUT3 #(
		.INIT('h80)
	) name25675 (
		\m6_addr_i[31]_pad ,
		_w8865_,
		_w8866_,
		_w27576_
	);
	LUT4 #(
		.INIT('hcedf)
	) name25676 (
		_w8860_,
		_w8863_,
		_w27575_,
		_w27576_,
		_w27577_
	);
	LUT4 #(
		.INIT('h7fff)
	) name25677 (
		_w27568_,
		_w27571_,
		_w27574_,
		_w27577_,
		_w27578_
	);
	LUT3 #(
		.INIT('h2a)
	) name25678 (
		\m3_addr_i[3]_pad ,
		_w8865_,
		_w8866_,
		_w27579_
	);
	LUT3 #(
		.INIT('h80)
	) name25679 (
		\m4_addr_i[3]_pad ,
		_w8865_,
		_w8866_,
		_w27580_
	);
	LUT4 #(
		.INIT('h9dbf)
	) name25680 (
		_w8860_,
		_w8863_,
		_w27579_,
		_w27580_,
		_w27581_
	);
	LUT3 #(
		.INIT('h80)
	) name25681 (
		\m6_addr_i[3]_pad ,
		_w8865_,
		_w8866_,
		_w27582_
	);
	LUT3 #(
		.INIT('h80)
	) name25682 (
		\m2_addr_i[3]_pad ,
		_w8865_,
		_w8866_,
		_w27583_
	);
	LUT4 #(
		.INIT('habef)
	) name25683 (
		_w8860_,
		_w8863_,
		_w27582_,
		_w27583_,
		_w27584_
	);
	LUT3 #(
		.INIT('h2a)
	) name25684 (
		\m5_addr_i[3]_pad ,
		_w8865_,
		_w8866_,
		_w27585_
	);
	LUT3 #(
		.INIT('h2a)
	) name25685 (
		\m1_addr_i[3]_pad ,
		_w8865_,
		_w8866_,
		_w27586_
	);
	LUT4 #(
		.INIT('h57df)
	) name25686 (
		_w8860_,
		_w8863_,
		_w27585_,
		_w27586_,
		_w27587_
	);
	LUT3 #(
		.INIT('h80)
	) name25687 (
		\m0_addr_i[3]_pad ,
		_w8865_,
		_w8866_,
		_w27588_
	);
	LUT3 #(
		.INIT('h2a)
	) name25688 (
		\m7_addr_i[3]_pad ,
		_w8865_,
		_w8866_,
		_w27589_
	);
	LUT4 #(
		.INIT('h6e7f)
	) name25689 (
		_w8860_,
		_w8863_,
		_w27588_,
		_w27589_,
		_w27590_
	);
	LUT4 #(
		.INIT('h7fff)
	) name25690 (
		_w27581_,
		_w27584_,
		_w27587_,
		_w27590_,
		_w27591_
	);
	LUT3 #(
		.INIT('h2a)
	) name25691 (
		\m3_addr_i[4]_pad ,
		_w8865_,
		_w8866_,
		_w27592_
	);
	LUT3 #(
		.INIT('h80)
	) name25692 (
		\m4_addr_i[4]_pad ,
		_w8865_,
		_w8866_,
		_w27593_
	);
	LUT4 #(
		.INIT('h9dbf)
	) name25693 (
		_w8860_,
		_w8863_,
		_w27592_,
		_w27593_,
		_w27594_
	);
	LUT3 #(
		.INIT('h80)
	) name25694 (
		\m6_addr_i[4]_pad ,
		_w8865_,
		_w8866_,
		_w27595_
	);
	LUT3 #(
		.INIT('h80)
	) name25695 (
		\m2_addr_i[4]_pad ,
		_w8865_,
		_w8866_,
		_w27596_
	);
	LUT4 #(
		.INIT('habef)
	) name25696 (
		_w8860_,
		_w8863_,
		_w27595_,
		_w27596_,
		_w27597_
	);
	LUT3 #(
		.INIT('h2a)
	) name25697 (
		\m5_addr_i[4]_pad ,
		_w8865_,
		_w8866_,
		_w27598_
	);
	LUT3 #(
		.INIT('h2a)
	) name25698 (
		\m1_addr_i[4]_pad ,
		_w8865_,
		_w8866_,
		_w27599_
	);
	LUT4 #(
		.INIT('h57df)
	) name25699 (
		_w8860_,
		_w8863_,
		_w27598_,
		_w27599_,
		_w27600_
	);
	LUT3 #(
		.INIT('h80)
	) name25700 (
		\m0_addr_i[4]_pad ,
		_w8865_,
		_w8866_,
		_w27601_
	);
	LUT3 #(
		.INIT('h2a)
	) name25701 (
		\m7_addr_i[4]_pad ,
		_w8865_,
		_w8866_,
		_w27602_
	);
	LUT4 #(
		.INIT('h6e7f)
	) name25702 (
		_w8860_,
		_w8863_,
		_w27601_,
		_w27602_,
		_w27603_
	);
	LUT4 #(
		.INIT('h7fff)
	) name25703 (
		_w27594_,
		_w27597_,
		_w27600_,
		_w27603_,
		_w27604_
	);
	LUT3 #(
		.INIT('h2a)
	) name25704 (
		\m1_addr_i[5]_pad ,
		_w8865_,
		_w8866_,
		_w27605_
	);
	LUT3 #(
		.INIT('h80)
	) name25705 (
		\m2_addr_i[5]_pad ,
		_w8865_,
		_w8866_,
		_w27606_
	);
	LUT4 #(
		.INIT('h3b7f)
	) name25706 (
		_w8860_,
		_w8863_,
		_w27605_,
		_w27606_,
		_w27607_
	);
	LUT3 #(
		.INIT('h2a)
	) name25707 (
		\m3_addr_i[5]_pad ,
		_w8865_,
		_w8866_,
		_w27608_
	);
	LUT3 #(
		.INIT('h2a)
	) name25708 (
		\m7_addr_i[5]_pad ,
		_w8865_,
		_w8866_,
		_w27609_
	);
	LUT4 #(
		.INIT('haebf)
	) name25709 (
		_w8860_,
		_w8863_,
		_w27608_,
		_w27609_,
		_w27610_
	);
	LUT3 #(
		.INIT('h80)
	) name25710 (
		\m4_addr_i[5]_pad ,
		_w8865_,
		_w8866_,
		_w27611_
	);
	LUT3 #(
		.INIT('h80)
	) name25711 (
		\m0_addr_i[5]_pad ,
		_w8865_,
		_w8866_,
		_w27612_
	);
	LUT4 #(
		.INIT('h57df)
	) name25712 (
		_w8860_,
		_w8863_,
		_w27611_,
		_w27612_,
		_w27613_
	);
	LUT3 #(
		.INIT('h80)
	) name25713 (
		\m6_addr_i[5]_pad ,
		_w8865_,
		_w8866_,
		_w27614_
	);
	LUT3 #(
		.INIT('h2a)
	) name25714 (
		\m5_addr_i[5]_pad ,
		_w8865_,
		_w8866_,
		_w27615_
	);
	LUT4 #(
		.INIT('hcdef)
	) name25715 (
		_w8860_,
		_w8863_,
		_w27614_,
		_w27615_,
		_w27616_
	);
	LUT4 #(
		.INIT('h7fff)
	) name25716 (
		_w27607_,
		_w27610_,
		_w27613_,
		_w27616_,
		_w27617_
	);
	LUT3 #(
		.INIT('h2a)
	) name25717 (
		\m1_addr_i[6]_pad ,
		_w8865_,
		_w8866_,
		_w27618_
	);
	LUT3 #(
		.INIT('h80)
	) name25718 (
		\m2_addr_i[6]_pad ,
		_w8865_,
		_w8866_,
		_w27619_
	);
	LUT4 #(
		.INIT('h3b7f)
	) name25719 (
		_w8860_,
		_w8863_,
		_w27618_,
		_w27619_,
		_w27620_
	);
	LUT3 #(
		.INIT('h80)
	) name25720 (
		\m0_addr_i[6]_pad ,
		_w8865_,
		_w8866_,
		_w27621_
	);
	LUT3 #(
		.INIT('h80)
	) name25721 (
		\m4_addr_i[6]_pad ,
		_w8865_,
		_w8866_,
		_w27622_
	);
	LUT4 #(
		.INIT('h5d7f)
	) name25722 (
		_w8860_,
		_w8863_,
		_w27621_,
		_w27622_,
		_w27623_
	);
	LUT3 #(
		.INIT('h2a)
	) name25723 (
		\m7_addr_i[6]_pad ,
		_w8865_,
		_w8866_,
		_w27624_
	);
	LUT3 #(
		.INIT('h2a)
	) name25724 (
		\m3_addr_i[6]_pad ,
		_w8865_,
		_w8866_,
		_w27625_
	);
	LUT4 #(
		.INIT('habef)
	) name25725 (
		_w8860_,
		_w8863_,
		_w27624_,
		_w27625_,
		_w27626_
	);
	LUT3 #(
		.INIT('h80)
	) name25726 (
		\m6_addr_i[6]_pad ,
		_w8865_,
		_w8866_,
		_w27627_
	);
	LUT3 #(
		.INIT('h2a)
	) name25727 (
		\m5_addr_i[6]_pad ,
		_w8865_,
		_w8866_,
		_w27628_
	);
	LUT4 #(
		.INIT('hcdef)
	) name25728 (
		_w8860_,
		_w8863_,
		_w27627_,
		_w27628_,
		_w27629_
	);
	LUT4 #(
		.INIT('h7fff)
	) name25729 (
		_w27620_,
		_w27623_,
		_w27626_,
		_w27629_,
		_w27630_
	);
	LUT3 #(
		.INIT('h80)
	) name25730 (
		\m6_addr_i[7]_pad ,
		_w8865_,
		_w8866_,
		_w27631_
	);
	LUT3 #(
		.INIT('h2a)
	) name25731 (
		\m5_addr_i[7]_pad ,
		_w8865_,
		_w8866_,
		_w27632_
	);
	LUT4 #(
		.INIT('hcdef)
	) name25732 (
		_w8860_,
		_w8863_,
		_w27631_,
		_w27632_,
		_w27633_
	);
	LUT3 #(
		.INIT('h2a)
	) name25733 (
		\m1_addr_i[7]_pad ,
		_w8865_,
		_w8866_,
		_w27634_
	);
	LUT3 #(
		.INIT('h80)
	) name25734 (
		\m4_addr_i[7]_pad ,
		_w8865_,
		_w8866_,
		_w27635_
	);
	LUT4 #(
		.INIT('h5d7f)
	) name25735 (
		_w8860_,
		_w8863_,
		_w27634_,
		_w27635_,
		_w27636_
	);
	LUT3 #(
		.INIT('h80)
	) name25736 (
		\m2_addr_i[7]_pad ,
		_w8865_,
		_w8866_,
		_w27637_
	);
	LUT3 #(
		.INIT('h2a)
	) name25737 (
		\m3_addr_i[7]_pad ,
		_w8865_,
		_w8866_,
		_w27638_
	);
	LUT3 #(
		.INIT('h57)
	) name25738 (
		_w8864_,
		_w27637_,
		_w27638_,
		_w27639_
	);
	LUT3 #(
		.INIT('h80)
	) name25739 (
		\m0_addr_i[7]_pad ,
		_w8865_,
		_w8866_,
		_w27640_
	);
	LUT3 #(
		.INIT('h2a)
	) name25740 (
		\m7_addr_i[7]_pad ,
		_w8865_,
		_w8866_,
		_w27641_
	);
	LUT4 #(
		.INIT('h6e7f)
	) name25741 (
		_w8860_,
		_w8863_,
		_w27640_,
		_w27641_,
		_w27642_
	);
	LUT4 #(
		.INIT('h7fff)
	) name25742 (
		_w27633_,
		_w27636_,
		_w27639_,
		_w27642_,
		_w27643_
	);
	LUT3 #(
		.INIT('h2a)
	) name25743 (
		\m1_addr_i[8]_pad ,
		_w8865_,
		_w8866_,
		_w27644_
	);
	LUT3 #(
		.INIT('h80)
	) name25744 (
		\m2_addr_i[8]_pad ,
		_w8865_,
		_w8866_,
		_w27645_
	);
	LUT4 #(
		.INIT('h3b7f)
	) name25745 (
		_w8860_,
		_w8863_,
		_w27644_,
		_w27645_,
		_w27646_
	);
	LUT3 #(
		.INIT('h2a)
	) name25746 (
		\m3_addr_i[8]_pad ,
		_w8865_,
		_w8866_,
		_w27647_
	);
	LUT3 #(
		.INIT('h2a)
	) name25747 (
		\m7_addr_i[8]_pad ,
		_w8865_,
		_w8866_,
		_w27648_
	);
	LUT4 #(
		.INIT('haebf)
	) name25748 (
		_w8860_,
		_w8863_,
		_w27647_,
		_w27648_,
		_w27649_
	);
	LUT3 #(
		.INIT('h80)
	) name25749 (
		\m4_addr_i[8]_pad ,
		_w8865_,
		_w8866_,
		_w27650_
	);
	LUT3 #(
		.INIT('h80)
	) name25750 (
		\m0_addr_i[8]_pad ,
		_w8865_,
		_w8866_,
		_w27651_
	);
	LUT4 #(
		.INIT('h57df)
	) name25751 (
		_w8860_,
		_w8863_,
		_w27650_,
		_w27651_,
		_w27652_
	);
	LUT3 #(
		.INIT('h80)
	) name25752 (
		\m6_addr_i[8]_pad ,
		_w8865_,
		_w8866_,
		_w27653_
	);
	LUT3 #(
		.INIT('h2a)
	) name25753 (
		\m5_addr_i[8]_pad ,
		_w8865_,
		_w8866_,
		_w27654_
	);
	LUT4 #(
		.INIT('hcdef)
	) name25754 (
		_w8860_,
		_w8863_,
		_w27653_,
		_w27654_,
		_w27655_
	);
	LUT4 #(
		.INIT('h7fff)
	) name25755 (
		_w27646_,
		_w27649_,
		_w27652_,
		_w27655_,
		_w27656_
	);
	LUT3 #(
		.INIT('h80)
	) name25756 (
		\m0_addr_i[9]_pad ,
		_w8865_,
		_w8866_,
		_w27657_
	);
	LUT3 #(
		.INIT('h2a)
	) name25757 (
		\m7_addr_i[9]_pad ,
		_w8865_,
		_w8866_,
		_w27658_
	);
	LUT4 #(
		.INIT('h6e7f)
	) name25758 (
		_w8860_,
		_w8863_,
		_w27657_,
		_w27658_,
		_w27659_
	);
	LUT3 #(
		.INIT('h2a)
	) name25759 (
		\m1_addr_i[9]_pad ,
		_w8865_,
		_w8866_,
		_w27660_
	);
	LUT3 #(
		.INIT('h80)
	) name25760 (
		\m4_addr_i[9]_pad ,
		_w8865_,
		_w8866_,
		_w27661_
	);
	LUT4 #(
		.INIT('h5d7f)
	) name25761 (
		_w8860_,
		_w8863_,
		_w27660_,
		_w27661_,
		_w27662_
	);
	LUT3 #(
		.INIT('h80)
	) name25762 (
		\m2_addr_i[9]_pad ,
		_w8865_,
		_w8866_,
		_w27663_
	);
	LUT3 #(
		.INIT('h2a)
	) name25763 (
		\m3_addr_i[9]_pad ,
		_w8865_,
		_w8866_,
		_w27664_
	);
	LUT3 #(
		.INIT('h57)
	) name25764 (
		_w8864_,
		_w27663_,
		_w27664_,
		_w27665_
	);
	LUT3 #(
		.INIT('h80)
	) name25765 (
		\m6_addr_i[9]_pad ,
		_w8865_,
		_w8866_,
		_w27666_
	);
	LUT3 #(
		.INIT('h2a)
	) name25766 (
		\m5_addr_i[9]_pad ,
		_w8865_,
		_w8866_,
		_w27667_
	);
	LUT4 #(
		.INIT('hcdef)
	) name25767 (
		_w8860_,
		_w8863_,
		_w27666_,
		_w27667_,
		_w27668_
	);
	LUT4 #(
		.INIT('h7fff)
	) name25768 (
		_w27659_,
		_w27662_,
		_w27665_,
		_w27668_,
		_w27669_
	);
	LUT3 #(
		.INIT('h80)
	) name25769 (
		\m0_data_i[0]_pad ,
		_w8865_,
		_w8866_,
		_w27670_
	);
	LUT3 #(
		.INIT('h2a)
	) name25770 (
		\m7_data_i[0]_pad ,
		_w8865_,
		_w8866_,
		_w27671_
	);
	LUT4 #(
		.INIT('h6e7f)
	) name25771 (
		_w8860_,
		_w8863_,
		_w27670_,
		_w27671_,
		_w27672_
	);
	LUT3 #(
		.INIT('h80)
	) name25772 (
		\m6_data_i[0]_pad ,
		_w8865_,
		_w8866_,
		_w27673_
	);
	LUT3 #(
		.INIT('h80)
	) name25773 (
		\m2_data_i[0]_pad ,
		_w8865_,
		_w8866_,
		_w27674_
	);
	LUT4 #(
		.INIT('habef)
	) name25774 (
		_w8860_,
		_w8863_,
		_w27673_,
		_w27674_,
		_w27675_
	);
	LUT3 #(
		.INIT('h2a)
	) name25775 (
		\m5_data_i[0]_pad ,
		_w8865_,
		_w8866_,
		_w27676_
	);
	LUT3 #(
		.INIT('h2a)
	) name25776 (
		\m1_data_i[0]_pad ,
		_w8865_,
		_w8866_,
		_w27677_
	);
	LUT4 #(
		.INIT('h57df)
	) name25777 (
		_w8860_,
		_w8863_,
		_w27676_,
		_w27677_,
		_w27678_
	);
	LUT3 #(
		.INIT('h2a)
	) name25778 (
		\m3_data_i[0]_pad ,
		_w8865_,
		_w8866_,
		_w27679_
	);
	LUT3 #(
		.INIT('h80)
	) name25779 (
		\m4_data_i[0]_pad ,
		_w8865_,
		_w8866_,
		_w27680_
	);
	LUT4 #(
		.INIT('h9dbf)
	) name25780 (
		_w8860_,
		_w8863_,
		_w27679_,
		_w27680_,
		_w27681_
	);
	LUT4 #(
		.INIT('h7fff)
	) name25781 (
		_w27672_,
		_w27675_,
		_w27678_,
		_w27681_,
		_w27682_
	);
	LUT3 #(
		.INIT('h80)
	) name25782 (
		\m6_data_i[10]_pad ,
		_w8865_,
		_w8866_,
		_w27683_
	);
	LUT3 #(
		.INIT('h2a)
	) name25783 (
		\m5_data_i[10]_pad ,
		_w8865_,
		_w8866_,
		_w27684_
	);
	LUT4 #(
		.INIT('hcdef)
	) name25784 (
		_w8860_,
		_w8863_,
		_w27683_,
		_w27684_,
		_w27685_
	);
	LUT3 #(
		.INIT('h2a)
	) name25785 (
		\m1_data_i[10]_pad ,
		_w8865_,
		_w8866_,
		_w27686_
	);
	LUT3 #(
		.INIT('h2a)
	) name25786 (
		\m7_data_i[10]_pad ,
		_w8865_,
		_w8866_,
		_w27687_
	);
	LUT4 #(
		.INIT('h6e7f)
	) name25787 (
		_w8860_,
		_w8863_,
		_w27686_,
		_w27687_,
		_w27688_
	);
	LUT3 #(
		.INIT('h80)
	) name25788 (
		\m2_data_i[10]_pad ,
		_w8865_,
		_w8866_,
		_w27689_
	);
	LUT3 #(
		.INIT('h80)
	) name25789 (
		\m0_data_i[10]_pad ,
		_w8865_,
		_w8866_,
		_w27690_
	);
	LUT4 #(
		.INIT('h37bf)
	) name25790 (
		_w8860_,
		_w8863_,
		_w27689_,
		_w27690_,
		_w27691_
	);
	LUT3 #(
		.INIT('h2a)
	) name25791 (
		\m3_data_i[10]_pad ,
		_w8865_,
		_w8866_,
		_w27692_
	);
	LUT3 #(
		.INIT('h80)
	) name25792 (
		\m4_data_i[10]_pad ,
		_w8865_,
		_w8866_,
		_w27693_
	);
	LUT4 #(
		.INIT('h9dbf)
	) name25793 (
		_w8860_,
		_w8863_,
		_w27692_,
		_w27693_,
		_w27694_
	);
	LUT4 #(
		.INIT('h7fff)
	) name25794 (
		_w27685_,
		_w27688_,
		_w27691_,
		_w27694_,
		_w27695_
	);
	LUT3 #(
		.INIT('h2a)
	) name25795 (
		\m1_data_i[11]_pad ,
		_w8865_,
		_w8866_,
		_w27696_
	);
	LUT3 #(
		.INIT('h80)
	) name25796 (
		\m2_data_i[11]_pad ,
		_w8865_,
		_w8866_,
		_w27697_
	);
	LUT4 #(
		.INIT('h3b7f)
	) name25797 (
		_w8860_,
		_w8863_,
		_w27696_,
		_w27697_,
		_w27698_
	);
	LUT3 #(
		.INIT('h80)
	) name25798 (
		\m6_data_i[11]_pad ,
		_w8865_,
		_w8866_,
		_w27699_
	);
	LUT3 #(
		.INIT('h80)
	) name25799 (
		\m4_data_i[11]_pad ,
		_w8865_,
		_w8866_,
		_w27700_
	);
	LUT4 #(
		.INIT('hcdef)
	) name25800 (
		_w8860_,
		_w8863_,
		_w27699_,
		_w27700_,
		_w27701_
	);
	LUT3 #(
		.INIT('h2a)
	) name25801 (
		\m5_data_i[11]_pad ,
		_w8865_,
		_w8866_,
		_w27702_
	);
	LUT3 #(
		.INIT('h2a)
	) name25802 (
		\m3_data_i[11]_pad ,
		_w8865_,
		_w8866_,
		_w27703_
	);
	LUT4 #(
		.INIT('h9bdf)
	) name25803 (
		_w8860_,
		_w8863_,
		_w27702_,
		_w27703_,
		_w27704_
	);
	LUT3 #(
		.INIT('h80)
	) name25804 (
		\m0_data_i[11]_pad ,
		_w8865_,
		_w8866_,
		_w27705_
	);
	LUT3 #(
		.INIT('h2a)
	) name25805 (
		\m7_data_i[11]_pad ,
		_w8865_,
		_w8866_,
		_w27706_
	);
	LUT4 #(
		.INIT('h6e7f)
	) name25806 (
		_w8860_,
		_w8863_,
		_w27705_,
		_w27706_,
		_w27707_
	);
	LUT4 #(
		.INIT('h7fff)
	) name25807 (
		_w27698_,
		_w27701_,
		_w27704_,
		_w27707_,
		_w27708_
	);
	LUT3 #(
		.INIT('h2a)
	) name25808 (
		\m1_data_i[12]_pad ,
		_w8865_,
		_w8866_,
		_w27709_
	);
	LUT3 #(
		.INIT('h80)
	) name25809 (
		\m2_data_i[12]_pad ,
		_w8865_,
		_w8866_,
		_w27710_
	);
	LUT4 #(
		.INIT('h3b7f)
	) name25810 (
		_w8860_,
		_w8863_,
		_w27709_,
		_w27710_,
		_w27711_
	);
	LUT3 #(
		.INIT('h80)
	) name25811 (
		\m6_data_i[12]_pad ,
		_w8865_,
		_w8866_,
		_w27712_
	);
	LUT3 #(
		.INIT('h2a)
	) name25812 (
		\m7_data_i[12]_pad ,
		_w8865_,
		_w8866_,
		_w27713_
	);
	LUT3 #(
		.INIT('h57)
	) name25813 (
		_w8878_,
		_w27712_,
		_w27713_,
		_w27714_
	);
	LUT3 #(
		.INIT('h2a)
	) name25814 (
		\m5_data_i[12]_pad ,
		_w8865_,
		_w8866_,
		_w27715_
	);
	LUT3 #(
		.INIT('h80)
	) name25815 (
		\m0_data_i[12]_pad ,
		_w8865_,
		_w8866_,
		_w27716_
	);
	LUT4 #(
		.INIT('h57df)
	) name25816 (
		_w8860_,
		_w8863_,
		_w27715_,
		_w27716_,
		_w27717_
	);
	LUT3 #(
		.INIT('h2a)
	) name25817 (
		\m3_data_i[12]_pad ,
		_w8865_,
		_w8866_,
		_w27718_
	);
	LUT3 #(
		.INIT('h80)
	) name25818 (
		\m4_data_i[12]_pad ,
		_w8865_,
		_w8866_,
		_w27719_
	);
	LUT4 #(
		.INIT('h9dbf)
	) name25819 (
		_w8860_,
		_w8863_,
		_w27718_,
		_w27719_,
		_w27720_
	);
	LUT4 #(
		.INIT('h7fff)
	) name25820 (
		_w27711_,
		_w27714_,
		_w27717_,
		_w27720_,
		_w27721_
	);
	LUT3 #(
		.INIT('h2a)
	) name25821 (
		\m1_data_i[13]_pad ,
		_w8865_,
		_w8866_,
		_w27722_
	);
	LUT3 #(
		.INIT('h80)
	) name25822 (
		\m2_data_i[13]_pad ,
		_w8865_,
		_w8866_,
		_w27723_
	);
	LUT4 #(
		.INIT('h3b7f)
	) name25823 (
		_w8860_,
		_w8863_,
		_w27722_,
		_w27723_,
		_w27724_
	);
	LUT3 #(
		.INIT('h80)
	) name25824 (
		\m6_data_i[13]_pad ,
		_w8865_,
		_w8866_,
		_w27725_
	);
	LUT3 #(
		.INIT('h2a)
	) name25825 (
		\m7_data_i[13]_pad ,
		_w8865_,
		_w8866_,
		_w27726_
	);
	LUT3 #(
		.INIT('h57)
	) name25826 (
		_w8878_,
		_w27725_,
		_w27726_,
		_w27727_
	);
	LUT3 #(
		.INIT('h2a)
	) name25827 (
		\m5_data_i[13]_pad ,
		_w8865_,
		_w8866_,
		_w27728_
	);
	LUT3 #(
		.INIT('h80)
	) name25828 (
		\m0_data_i[13]_pad ,
		_w8865_,
		_w8866_,
		_w27729_
	);
	LUT4 #(
		.INIT('h57df)
	) name25829 (
		_w8860_,
		_w8863_,
		_w27728_,
		_w27729_,
		_w27730_
	);
	LUT3 #(
		.INIT('h2a)
	) name25830 (
		\m3_data_i[13]_pad ,
		_w8865_,
		_w8866_,
		_w27731_
	);
	LUT3 #(
		.INIT('h80)
	) name25831 (
		\m4_data_i[13]_pad ,
		_w8865_,
		_w8866_,
		_w27732_
	);
	LUT4 #(
		.INIT('h9dbf)
	) name25832 (
		_w8860_,
		_w8863_,
		_w27731_,
		_w27732_,
		_w27733_
	);
	LUT4 #(
		.INIT('h7fff)
	) name25833 (
		_w27724_,
		_w27727_,
		_w27730_,
		_w27733_,
		_w27734_
	);
	LUT3 #(
		.INIT('h2a)
	) name25834 (
		\m3_data_i[14]_pad ,
		_w8865_,
		_w8866_,
		_w27735_
	);
	LUT3 #(
		.INIT('h80)
	) name25835 (
		\m4_data_i[14]_pad ,
		_w8865_,
		_w8866_,
		_w27736_
	);
	LUT4 #(
		.INIT('h9dbf)
	) name25836 (
		_w8860_,
		_w8863_,
		_w27735_,
		_w27736_,
		_w27737_
	);
	LUT3 #(
		.INIT('h80)
	) name25837 (
		\m6_data_i[14]_pad ,
		_w8865_,
		_w8866_,
		_w27738_
	);
	LUT3 #(
		.INIT('h2a)
	) name25838 (
		\m7_data_i[14]_pad ,
		_w8865_,
		_w8866_,
		_w27739_
	);
	LUT3 #(
		.INIT('h57)
	) name25839 (
		_w8878_,
		_w27738_,
		_w27739_,
		_w27740_
	);
	LUT3 #(
		.INIT('h2a)
	) name25840 (
		\m5_data_i[14]_pad ,
		_w8865_,
		_w8866_,
		_w27741_
	);
	LUT3 #(
		.INIT('h80)
	) name25841 (
		\m0_data_i[14]_pad ,
		_w8865_,
		_w8866_,
		_w27742_
	);
	LUT4 #(
		.INIT('h57df)
	) name25842 (
		_w8860_,
		_w8863_,
		_w27741_,
		_w27742_,
		_w27743_
	);
	LUT3 #(
		.INIT('h2a)
	) name25843 (
		\m1_data_i[14]_pad ,
		_w8865_,
		_w8866_,
		_w27744_
	);
	LUT3 #(
		.INIT('h80)
	) name25844 (
		\m2_data_i[14]_pad ,
		_w8865_,
		_w8866_,
		_w27745_
	);
	LUT4 #(
		.INIT('h3b7f)
	) name25845 (
		_w8860_,
		_w8863_,
		_w27744_,
		_w27745_,
		_w27746_
	);
	LUT4 #(
		.INIT('h7fff)
	) name25846 (
		_w27737_,
		_w27740_,
		_w27743_,
		_w27746_,
		_w27747_
	);
	LUT3 #(
		.INIT('h80)
	) name25847 (
		\m6_data_i[15]_pad ,
		_w8865_,
		_w8866_,
		_w27748_
	);
	LUT3 #(
		.INIT('h2a)
	) name25848 (
		\m5_data_i[15]_pad ,
		_w8865_,
		_w8866_,
		_w27749_
	);
	LUT4 #(
		.INIT('hcdef)
	) name25849 (
		_w8860_,
		_w8863_,
		_w27748_,
		_w27749_,
		_w27750_
	);
	LUT3 #(
		.INIT('h2a)
	) name25850 (
		\m3_data_i[15]_pad ,
		_w8865_,
		_w8866_,
		_w27751_
	);
	LUT3 #(
		.INIT('h80)
	) name25851 (
		\m2_data_i[15]_pad ,
		_w8865_,
		_w8866_,
		_w27752_
	);
	LUT3 #(
		.INIT('h57)
	) name25852 (
		_w8864_,
		_w27751_,
		_w27752_,
		_w27753_
	);
	LUT3 #(
		.INIT('h80)
	) name25853 (
		\m4_data_i[15]_pad ,
		_w8865_,
		_w8866_,
		_w27754_
	);
	LUT3 #(
		.INIT('h2a)
	) name25854 (
		\m1_data_i[15]_pad ,
		_w8865_,
		_w8866_,
		_w27755_
	);
	LUT4 #(
		.INIT('h57df)
	) name25855 (
		_w8860_,
		_w8863_,
		_w27754_,
		_w27755_,
		_w27756_
	);
	LUT3 #(
		.INIT('h80)
	) name25856 (
		\m0_data_i[15]_pad ,
		_w8865_,
		_w8866_,
		_w27757_
	);
	LUT3 #(
		.INIT('h2a)
	) name25857 (
		\m7_data_i[15]_pad ,
		_w8865_,
		_w8866_,
		_w27758_
	);
	LUT4 #(
		.INIT('h6e7f)
	) name25858 (
		_w8860_,
		_w8863_,
		_w27757_,
		_w27758_,
		_w27759_
	);
	LUT4 #(
		.INIT('h7fff)
	) name25859 (
		_w27750_,
		_w27753_,
		_w27756_,
		_w27759_,
		_w27760_
	);
	LUT3 #(
		.INIT('h2a)
	) name25860 (
		\m1_data_i[16]_pad ,
		_w8865_,
		_w8866_,
		_w27761_
	);
	LUT3 #(
		.INIT('h80)
	) name25861 (
		\m2_data_i[16]_pad ,
		_w8865_,
		_w8866_,
		_w27762_
	);
	LUT4 #(
		.INIT('h3b7f)
	) name25862 (
		_w8860_,
		_w8863_,
		_w27761_,
		_w27762_,
		_w27763_
	);
	LUT3 #(
		.INIT('h80)
	) name25863 (
		\m0_data_i[16]_pad ,
		_w8865_,
		_w8866_,
		_w27764_
	);
	LUT3 #(
		.INIT('h80)
	) name25864 (
		\m4_data_i[16]_pad ,
		_w8865_,
		_w8866_,
		_w27765_
	);
	LUT4 #(
		.INIT('h5d7f)
	) name25865 (
		_w8860_,
		_w8863_,
		_w27764_,
		_w27765_,
		_w27766_
	);
	LUT3 #(
		.INIT('h2a)
	) name25866 (
		\m7_data_i[16]_pad ,
		_w8865_,
		_w8866_,
		_w27767_
	);
	LUT3 #(
		.INIT('h2a)
	) name25867 (
		\m3_data_i[16]_pad ,
		_w8865_,
		_w8866_,
		_w27768_
	);
	LUT4 #(
		.INIT('habef)
	) name25868 (
		_w8860_,
		_w8863_,
		_w27767_,
		_w27768_,
		_w27769_
	);
	LUT3 #(
		.INIT('h80)
	) name25869 (
		\m6_data_i[16]_pad ,
		_w8865_,
		_w8866_,
		_w27770_
	);
	LUT3 #(
		.INIT('h2a)
	) name25870 (
		\m5_data_i[16]_pad ,
		_w8865_,
		_w8866_,
		_w27771_
	);
	LUT4 #(
		.INIT('hcdef)
	) name25871 (
		_w8860_,
		_w8863_,
		_w27770_,
		_w27771_,
		_w27772_
	);
	LUT4 #(
		.INIT('h7fff)
	) name25872 (
		_w27763_,
		_w27766_,
		_w27769_,
		_w27772_,
		_w27773_
	);
	LUT3 #(
		.INIT('h2a)
	) name25873 (
		\m3_data_i[17]_pad ,
		_w8865_,
		_w8866_,
		_w27774_
	);
	LUT3 #(
		.INIT('h80)
	) name25874 (
		\m4_data_i[17]_pad ,
		_w8865_,
		_w8866_,
		_w27775_
	);
	LUT4 #(
		.INIT('h9dbf)
	) name25875 (
		_w8860_,
		_w8863_,
		_w27774_,
		_w27775_,
		_w27776_
	);
	LUT3 #(
		.INIT('h80)
	) name25876 (
		\m0_data_i[17]_pad ,
		_w8865_,
		_w8866_,
		_w27777_
	);
	LUT3 #(
		.INIT('h2a)
	) name25877 (
		\m5_data_i[17]_pad ,
		_w8865_,
		_w8866_,
		_w27778_
	);
	LUT4 #(
		.INIT('h5d7f)
	) name25878 (
		_w8860_,
		_w8863_,
		_w27777_,
		_w27778_,
		_w27779_
	);
	LUT3 #(
		.INIT('h2a)
	) name25879 (
		\m7_data_i[17]_pad ,
		_w8865_,
		_w8866_,
		_w27780_
	);
	LUT3 #(
		.INIT('h80)
	) name25880 (
		\m6_data_i[17]_pad ,
		_w8865_,
		_w8866_,
		_w27781_
	);
	LUT3 #(
		.INIT('h57)
	) name25881 (
		_w8878_,
		_w27780_,
		_w27781_,
		_w27782_
	);
	LUT3 #(
		.INIT('h2a)
	) name25882 (
		\m1_data_i[17]_pad ,
		_w8865_,
		_w8866_,
		_w27783_
	);
	LUT3 #(
		.INIT('h80)
	) name25883 (
		\m2_data_i[17]_pad ,
		_w8865_,
		_w8866_,
		_w27784_
	);
	LUT4 #(
		.INIT('h3b7f)
	) name25884 (
		_w8860_,
		_w8863_,
		_w27783_,
		_w27784_,
		_w27785_
	);
	LUT4 #(
		.INIT('h7fff)
	) name25885 (
		_w27776_,
		_w27779_,
		_w27782_,
		_w27785_,
		_w27786_
	);
	LUT3 #(
		.INIT('h2a)
	) name25886 (
		\m3_data_i[18]_pad ,
		_w8865_,
		_w8866_,
		_w27787_
	);
	LUT3 #(
		.INIT('h80)
	) name25887 (
		\m4_data_i[18]_pad ,
		_w8865_,
		_w8866_,
		_w27788_
	);
	LUT4 #(
		.INIT('h9dbf)
	) name25888 (
		_w8860_,
		_w8863_,
		_w27787_,
		_w27788_,
		_w27789_
	);
	LUT3 #(
		.INIT('h80)
	) name25889 (
		\m6_data_i[18]_pad ,
		_w8865_,
		_w8866_,
		_w27790_
	);
	LUT3 #(
		.INIT('h80)
	) name25890 (
		\m2_data_i[18]_pad ,
		_w8865_,
		_w8866_,
		_w27791_
	);
	LUT4 #(
		.INIT('habef)
	) name25891 (
		_w8860_,
		_w8863_,
		_w27790_,
		_w27791_,
		_w27792_
	);
	LUT3 #(
		.INIT('h2a)
	) name25892 (
		\m5_data_i[18]_pad ,
		_w8865_,
		_w8866_,
		_w27793_
	);
	LUT3 #(
		.INIT('h2a)
	) name25893 (
		\m1_data_i[18]_pad ,
		_w8865_,
		_w8866_,
		_w27794_
	);
	LUT4 #(
		.INIT('h57df)
	) name25894 (
		_w8860_,
		_w8863_,
		_w27793_,
		_w27794_,
		_w27795_
	);
	LUT3 #(
		.INIT('h80)
	) name25895 (
		\m0_data_i[18]_pad ,
		_w8865_,
		_w8866_,
		_w27796_
	);
	LUT3 #(
		.INIT('h2a)
	) name25896 (
		\m7_data_i[18]_pad ,
		_w8865_,
		_w8866_,
		_w27797_
	);
	LUT4 #(
		.INIT('h6e7f)
	) name25897 (
		_w8860_,
		_w8863_,
		_w27796_,
		_w27797_,
		_w27798_
	);
	LUT4 #(
		.INIT('h7fff)
	) name25898 (
		_w27789_,
		_w27792_,
		_w27795_,
		_w27798_,
		_w27799_
	);
	LUT3 #(
		.INIT('h80)
	) name25899 (
		\m0_data_i[19]_pad ,
		_w8865_,
		_w8866_,
		_w27800_
	);
	LUT3 #(
		.INIT('h2a)
	) name25900 (
		\m7_data_i[19]_pad ,
		_w8865_,
		_w8866_,
		_w27801_
	);
	LUT4 #(
		.INIT('h6e7f)
	) name25901 (
		_w8860_,
		_w8863_,
		_w27800_,
		_w27801_,
		_w27802_
	);
	LUT3 #(
		.INIT('h2a)
	) name25902 (
		\m1_data_i[19]_pad ,
		_w8865_,
		_w8866_,
		_w27803_
	);
	LUT3 #(
		.INIT('h80)
	) name25903 (
		\m4_data_i[19]_pad ,
		_w8865_,
		_w8866_,
		_w27804_
	);
	LUT4 #(
		.INIT('h5d7f)
	) name25904 (
		_w8860_,
		_w8863_,
		_w27803_,
		_w27804_,
		_w27805_
	);
	LUT3 #(
		.INIT('h80)
	) name25905 (
		\m2_data_i[19]_pad ,
		_w8865_,
		_w8866_,
		_w27806_
	);
	LUT3 #(
		.INIT('h2a)
	) name25906 (
		\m3_data_i[19]_pad ,
		_w8865_,
		_w8866_,
		_w27807_
	);
	LUT3 #(
		.INIT('h57)
	) name25907 (
		_w8864_,
		_w27806_,
		_w27807_,
		_w27808_
	);
	LUT3 #(
		.INIT('h80)
	) name25908 (
		\m6_data_i[19]_pad ,
		_w8865_,
		_w8866_,
		_w27809_
	);
	LUT3 #(
		.INIT('h2a)
	) name25909 (
		\m5_data_i[19]_pad ,
		_w8865_,
		_w8866_,
		_w27810_
	);
	LUT4 #(
		.INIT('hcdef)
	) name25910 (
		_w8860_,
		_w8863_,
		_w27809_,
		_w27810_,
		_w27811_
	);
	LUT4 #(
		.INIT('h7fff)
	) name25911 (
		_w27802_,
		_w27805_,
		_w27808_,
		_w27811_,
		_w27812_
	);
	LUT3 #(
		.INIT('h2a)
	) name25912 (
		\m3_data_i[1]_pad ,
		_w8865_,
		_w8866_,
		_w27813_
	);
	LUT3 #(
		.INIT('h80)
	) name25913 (
		\m4_data_i[1]_pad ,
		_w8865_,
		_w8866_,
		_w27814_
	);
	LUT4 #(
		.INIT('h9dbf)
	) name25914 (
		_w8860_,
		_w8863_,
		_w27813_,
		_w27814_,
		_w27815_
	);
	LUT3 #(
		.INIT('h80)
	) name25915 (
		\m6_data_i[1]_pad ,
		_w8865_,
		_w8866_,
		_w27816_
	);
	LUT3 #(
		.INIT('h80)
	) name25916 (
		\m2_data_i[1]_pad ,
		_w8865_,
		_w8866_,
		_w27817_
	);
	LUT4 #(
		.INIT('habef)
	) name25917 (
		_w8860_,
		_w8863_,
		_w27816_,
		_w27817_,
		_w27818_
	);
	LUT3 #(
		.INIT('h2a)
	) name25918 (
		\m5_data_i[1]_pad ,
		_w8865_,
		_w8866_,
		_w27819_
	);
	LUT3 #(
		.INIT('h2a)
	) name25919 (
		\m1_data_i[1]_pad ,
		_w8865_,
		_w8866_,
		_w27820_
	);
	LUT4 #(
		.INIT('h57df)
	) name25920 (
		_w8860_,
		_w8863_,
		_w27819_,
		_w27820_,
		_w27821_
	);
	LUT3 #(
		.INIT('h80)
	) name25921 (
		\m0_data_i[1]_pad ,
		_w8865_,
		_w8866_,
		_w27822_
	);
	LUT3 #(
		.INIT('h2a)
	) name25922 (
		\m7_data_i[1]_pad ,
		_w8865_,
		_w8866_,
		_w27823_
	);
	LUT4 #(
		.INIT('h6e7f)
	) name25923 (
		_w8860_,
		_w8863_,
		_w27822_,
		_w27823_,
		_w27824_
	);
	LUT4 #(
		.INIT('h7fff)
	) name25924 (
		_w27815_,
		_w27818_,
		_w27821_,
		_w27824_,
		_w27825_
	);
	LUT3 #(
		.INIT('h2a)
	) name25925 (
		\m3_data_i[20]_pad ,
		_w8865_,
		_w8866_,
		_w27826_
	);
	LUT3 #(
		.INIT('h80)
	) name25926 (
		\m4_data_i[20]_pad ,
		_w8865_,
		_w8866_,
		_w27827_
	);
	LUT4 #(
		.INIT('h9dbf)
	) name25927 (
		_w8860_,
		_w8863_,
		_w27826_,
		_w27827_,
		_w27828_
	);
	LUT3 #(
		.INIT('h80)
	) name25928 (
		\m6_data_i[20]_pad ,
		_w8865_,
		_w8866_,
		_w27829_
	);
	LUT3 #(
		.INIT('h80)
	) name25929 (
		\m2_data_i[20]_pad ,
		_w8865_,
		_w8866_,
		_w27830_
	);
	LUT4 #(
		.INIT('habef)
	) name25930 (
		_w8860_,
		_w8863_,
		_w27829_,
		_w27830_,
		_w27831_
	);
	LUT3 #(
		.INIT('h2a)
	) name25931 (
		\m5_data_i[20]_pad ,
		_w8865_,
		_w8866_,
		_w27832_
	);
	LUT3 #(
		.INIT('h2a)
	) name25932 (
		\m1_data_i[20]_pad ,
		_w8865_,
		_w8866_,
		_w27833_
	);
	LUT4 #(
		.INIT('h57df)
	) name25933 (
		_w8860_,
		_w8863_,
		_w27832_,
		_w27833_,
		_w27834_
	);
	LUT3 #(
		.INIT('h80)
	) name25934 (
		\m0_data_i[20]_pad ,
		_w8865_,
		_w8866_,
		_w27835_
	);
	LUT3 #(
		.INIT('h2a)
	) name25935 (
		\m7_data_i[20]_pad ,
		_w8865_,
		_w8866_,
		_w27836_
	);
	LUT4 #(
		.INIT('h6e7f)
	) name25936 (
		_w8860_,
		_w8863_,
		_w27835_,
		_w27836_,
		_w27837_
	);
	LUT4 #(
		.INIT('h7fff)
	) name25937 (
		_w27828_,
		_w27831_,
		_w27834_,
		_w27837_,
		_w27838_
	);
	LUT3 #(
		.INIT('h2a)
	) name25938 (
		\m1_data_i[21]_pad ,
		_w8865_,
		_w8866_,
		_w27839_
	);
	LUT3 #(
		.INIT('h80)
	) name25939 (
		\m2_data_i[21]_pad ,
		_w8865_,
		_w8866_,
		_w27840_
	);
	LUT4 #(
		.INIT('h3b7f)
	) name25940 (
		_w8860_,
		_w8863_,
		_w27839_,
		_w27840_,
		_w27841_
	);
	LUT3 #(
		.INIT('h80)
	) name25941 (
		\m6_data_i[21]_pad ,
		_w8865_,
		_w8866_,
		_w27842_
	);
	LUT3 #(
		.INIT('h2a)
	) name25942 (
		\m7_data_i[21]_pad ,
		_w8865_,
		_w8866_,
		_w27843_
	);
	LUT3 #(
		.INIT('h57)
	) name25943 (
		_w8878_,
		_w27842_,
		_w27843_,
		_w27844_
	);
	LUT3 #(
		.INIT('h2a)
	) name25944 (
		\m5_data_i[21]_pad ,
		_w8865_,
		_w8866_,
		_w27845_
	);
	LUT3 #(
		.INIT('h80)
	) name25945 (
		\m0_data_i[21]_pad ,
		_w8865_,
		_w8866_,
		_w27846_
	);
	LUT4 #(
		.INIT('h57df)
	) name25946 (
		_w8860_,
		_w8863_,
		_w27845_,
		_w27846_,
		_w27847_
	);
	LUT3 #(
		.INIT('h2a)
	) name25947 (
		\m3_data_i[21]_pad ,
		_w8865_,
		_w8866_,
		_w27848_
	);
	LUT3 #(
		.INIT('h80)
	) name25948 (
		\m4_data_i[21]_pad ,
		_w8865_,
		_w8866_,
		_w27849_
	);
	LUT4 #(
		.INIT('h9dbf)
	) name25949 (
		_w8860_,
		_w8863_,
		_w27848_,
		_w27849_,
		_w27850_
	);
	LUT4 #(
		.INIT('h7fff)
	) name25950 (
		_w27841_,
		_w27844_,
		_w27847_,
		_w27850_,
		_w27851_
	);
	LUT3 #(
		.INIT('h2a)
	) name25951 (
		\m3_data_i[22]_pad ,
		_w8865_,
		_w8866_,
		_w27852_
	);
	LUT3 #(
		.INIT('h80)
	) name25952 (
		\m4_data_i[22]_pad ,
		_w8865_,
		_w8866_,
		_w27853_
	);
	LUT4 #(
		.INIT('h9dbf)
	) name25953 (
		_w8860_,
		_w8863_,
		_w27852_,
		_w27853_,
		_w27854_
	);
	LUT3 #(
		.INIT('h80)
	) name25954 (
		\m6_data_i[22]_pad ,
		_w8865_,
		_w8866_,
		_w27855_
	);
	LUT3 #(
		.INIT('h80)
	) name25955 (
		\m2_data_i[22]_pad ,
		_w8865_,
		_w8866_,
		_w27856_
	);
	LUT4 #(
		.INIT('habef)
	) name25956 (
		_w8860_,
		_w8863_,
		_w27855_,
		_w27856_,
		_w27857_
	);
	LUT3 #(
		.INIT('h2a)
	) name25957 (
		\m5_data_i[22]_pad ,
		_w8865_,
		_w8866_,
		_w27858_
	);
	LUT3 #(
		.INIT('h2a)
	) name25958 (
		\m1_data_i[22]_pad ,
		_w8865_,
		_w8866_,
		_w27859_
	);
	LUT4 #(
		.INIT('h57df)
	) name25959 (
		_w8860_,
		_w8863_,
		_w27858_,
		_w27859_,
		_w27860_
	);
	LUT3 #(
		.INIT('h80)
	) name25960 (
		\m0_data_i[22]_pad ,
		_w8865_,
		_w8866_,
		_w27861_
	);
	LUT3 #(
		.INIT('h2a)
	) name25961 (
		\m7_data_i[22]_pad ,
		_w8865_,
		_w8866_,
		_w27862_
	);
	LUT4 #(
		.INIT('h6e7f)
	) name25962 (
		_w8860_,
		_w8863_,
		_w27861_,
		_w27862_,
		_w27863_
	);
	LUT4 #(
		.INIT('h7fff)
	) name25963 (
		_w27854_,
		_w27857_,
		_w27860_,
		_w27863_,
		_w27864_
	);
	LUT3 #(
		.INIT('h2a)
	) name25964 (
		\m3_data_i[23]_pad ,
		_w8865_,
		_w8866_,
		_w27865_
	);
	LUT3 #(
		.INIT('h80)
	) name25965 (
		\m4_data_i[23]_pad ,
		_w8865_,
		_w8866_,
		_w27866_
	);
	LUT4 #(
		.INIT('h9dbf)
	) name25966 (
		_w8860_,
		_w8863_,
		_w27865_,
		_w27866_,
		_w27867_
	);
	LUT3 #(
		.INIT('h80)
	) name25967 (
		\m6_data_i[23]_pad ,
		_w8865_,
		_w8866_,
		_w27868_
	);
	LUT3 #(
		.INIT('h80)
	) name25968 (
		\m2_data_i[23]_pad ,
		_w8865_,
		_w8866_,
		_w27869_
	);
	LUT4 #(
		.INIT('habef)
	) name25969 (
		_w8860_,
		_w8863_,
		_w27868_,
		_w27869_,
		_w27870_
	);
	LUT3 #(
		.INIT('h2a)
	) name25970 (
		\m5_data_i[23]_pad ,
		_w8865_,
		_w8866_,
		_w27871_
	);
	LUT3 #(
		.INIT('h2a)
	) name25971 (
		\m1_data_i[23]_pad ,
		_w8865_,
		_w8866_,
		_w27872_
	);
	LUT4 #(
		.INIT('h57df)
	) name25972 (
		_w8860_,
		_w8863_,
		_w27871_,
		_w27872_,
		_w27873_
	);
	LUT3 #(
		.INIT('h80)
	) name25973 (
		\m0_data_i[23]_pad ,
		_w8865_,
		_w8866_,
		_w27874_
	);
	LUT3 #(
		.INIT('h2a)
	) name25974 (
		\m7_data_i[23]_pad ,
		_w8865_,
		_w8866_,
		_w27875_
	);
	LUT4 #(
		.INIT('h6e7f)
	) name25975 (
		_w8860_,
		_w8863_,
		_w27874_,
		_w27875_,
		_w27876_
	);
	LUT4 #(
		.INIT('h7fff)
	) name25976 (
		_w27867_,
		_w27870_,
		_w27873_,
		_w27876_,
		_w27877_
	);
	LUT3 #(
		.INIT('h2a)
	) name25977 (
		\m3_data_i[24]_pad ,
		_w8865_,
		_w8866_,
		_w27878_
	);
	LUT3 #(
		.INIT('h80)
	) name25978 (
		\m4_data_i[24]_pad ,
		_w8865_,
		_w8866_,
		_w27879_
	);
	LUT4 #(
		.INIT('h9dbf)
	) name25979 (
		_w8860_,
		_w8863_,
		_w27878_,
		_w27879_,
		_w27880_
	);
	LUT3 #(
		.INIT('h80)
	) name25980 (
		\m6_data_i[24]_pad ,
		_w8865_,
		_w8866_,
		_w27881_
	);
	LUT3 #(
		.INIT('h80)
	) name25981 (
		\m2_data_i[24]_pad ,
		_w8865_,
		_w8866_,
		_w27882_
	);
	LUT4 #(
		.INIT('habef)
	) name25982 (
		_w8860_,
		_w8863_,
		_w27881_,
		_w27882_,
		_w27883_
	);
	LUT3 #(
		.INIT('h2a)
	) name25983 (
		\m5_data_i[24]_pad ,
		_w8865_,
		_w8866_,
		_w27884_
	);
	LUT3 #(
		.INIT('h2a)
	) name25984 (
		\m1_data_i[24]_pad ,
		_w8865_,
		_w8866_,
		_w27885_
	);
	LUT4 #(
		.INIT('h57df)
	) name25985 (
		_w8860_,
		_w8863_,
		_w27884_,
		_w27885_,
		_w27886_
	);
	LUT3 #(
		.INIT('h80)
	) name25986 (
		\m0_data_i[24]_pad ,
		_w8865_,
		_w8866_,
		_w27887_
	);
	LUT3 #(
		.INIT('h2a)
	) name25987 (
		\m7_data_i[24]_pad ,
		_w8865_,
		_w8866_,
		_w27888_
	);
	LUT4 #(
		.INIT('h6e7f)
	) name25988 (
		_w8860_,
		_w8863_,
		_w27887_,
		_w27888_,
		_w27889_
	);
	LUT4 #(
		.INIT('h7fff)
	) name25989 (
		_w27880_,
		_w27883_,
		_w27886_,
		_w27889_,
		_w27890_
	);
	LUT3 #(
		.INIT('h2a)
	) name25990 (
		\m3_data_i[25]_pad ,
		_w8865_,
		_w8866_,
		_w27891_
	);
	LUT3 #(
		.INIT('h80)
	) name25991 (
		\m4_data_i[25]_pad ,
		_w8865_,
		_w8866_,
		_w27892_
	);
	LUT4 #(
		.INIT('h9dbf)
	) name25992 (
		_w8860_,
		_w8863_,
		_w27891_,
		_w27892_,
		_w27893_
	);
	LUT3 #(
		.INIT('h80)
	) name25993 (
		\m6_data_i[25]_pad ,
		_w8865_,
		_w8866_,
		_w27894_
	);
	LUT3 #(
		.INIT('h2a)
	) name25994 (
		\m7_data_i[25]_pad ,
		_w8865_,
		_w8866_,
		_w27895_
	);
	LUT3 #(
		.INIT('h57)
	) name25995 (
		_w8878_,
		_w27894_,
		_w27895_,
		_w27896_
	);
	LUT3 #(
		.INIT('h2a)
	) name25996 (
		\m5_data_i[25]_pad ,
		_w8865_,
		_w8866_,
		_w27897_
	);
	LUT3 #(
		.INIT('h80)
	) name25997 (
		\m0_data_i[25]_pad ,
		_w8865_,
		_w8866_,
		_w27898_
	);
	LUT4 #(
		.INIT('h57df)
	) name25998 (
		_w8860_,
		_w8863_,
		_w27897_,
		_w27898_,
		_w27899_
	);
	LUT3 #(
		.INIT('h2a)
	) name25999 (
		\m1_data_i[25]_pad ,
		_w8865_,
		_w8866_,
		_w27900_
	);
	LUT3 #(
		.INIT('h80)
	) name26000 (
		\m2_data_i[25]_pad ,
		_w8865_,
		_w8866_,
		_w27901_
	);
	LUT4 #(
		.INIT('h3b7f)
	) name26001 (
		_w8860_,
		_w8863_,
		_w27900_,
		_w27901_,
		_w27902_
	);
	LUT4 #(
		.INIT('h7fff)
	) name26002 (
		_w27893_,
		_w27896_,
		_w27899_,
		_w27902_,
		_w27903_
	);
	LUT3 #(
		.INIT('h2a)
	) name26003 (
		\m1_data_i[26]_pad ,
		_w8865_,
		_w8866_,
		_w27904_
	);
	LUT3 #(
		.INIT('h80)
	) name26004 (
		\m2_data_i[26]_pad ,
		_w8865_,
		_w8866_,
		_w27905_
	);
	LUT4 #(
		.INIT('h3b7f)
	) name26005 (
		_w8860_,
		_w8863_,
		_w27904_,
		_w27905_,
		_w27906_
	);
	LUT3 #(
		.INIT('h80)
	) name26006 (
		\m0_data_i[26]_pad ,
		_w8865_,
		_w8866_,
		_w27907_
	);
	LUT3 #(
		.INIT('h80)
	) name26007 (
		\m4_data_i[26]_pad ,
		_w8865_,
		_w8866_,
		_w27908_
	);
	LUT4 #(
		.INIT('h5d7f)
	) name26008 (
		_w8860_,
		_w8863_,
		_w27907_,
		_w27908_,
		_w27909_
	);
	LUT3 #(
		.INIT('h2a)
	) name26009 (
		\m7_data_i[26]_pad ,
		_w8865_,
		_w8866_,
		_w27910_
	);
	LUT3 #(
		.INIT('h2a)
	) name26010 (
		\m3_data_i[26]_pad ,
		_w8865_,
		_w8866_,
		_w27911_
	);
	LUT4 #(
		.INIT('habef)
	) name26011 (
		_w8860_,
		_w8863_,
		_w27910_,
		_w27911_,
		_w27912_
	);
	LUT3 #(
		.INIT('h80)
	) name26012 (
		\m6_data_i[26]_pad ,
		_w8865_,
		_w8866_,
		_w27913_
	);
	LUT3 #(
		.INIT('h2a)
	) name26013 (
		\m5_data_i[26]_pad ,
		_w8865_,
		_w8866_,
		_w27914_
	);
	LUT4 #(
		.INIT('hcdef)
	) name26014 (
		_w8860_,
		_w8863_,
		_w27913_,
		_w27914_,
		_w27915_
	);
	LUT4 #(
		.INIT('h7fff)
	) name26015 (
		_w27906_,
		_w27909_,
		_w27912_,
		_w27915_,
		_w27916_
	);
	LUT3 #(
		.INIT('h2a)
	) name26016 (
		\m3_data_i[27]_pad ,
		_w8865_,
		_w8866_,
		_w27917_
	);
	LUT3 #(
		.INIT('h80)
	) name26017 (
		\m4_data_i[27]_pad ,
		_w8865_,
		_w8866_,
		_w27918_
	);
	LUT4 #(
		.INIT('h9dbf)
	) name26018 (
		_w8860_,
		_w8863_,
		_w27917_,
		_w27918_,
		_w27919_
	);
	LUT3 #(
		.INIT('h80)
	) name26019 (
		\m0_data_i[27]_pad ,
		_w8865_,
		_w8866_,
		_w27920_
	);
	LUT3 #(
		.INIT('h80)
	) name26020 (
		\m2_data_i[27]_pad ,
		_w8865_,
		_w8866_,
		_w27921_
	);
	LUT4 #(
		.INIT('h3b7f)
	) name26021 (
		_w8860_,
		_w8863_,
		_w27920_,
		_w27921_,
		_w27922_
	);
	LUT3 #(
		.INIT('h2a)
	) name26022 (
		\m7_data_i[27]_pad ,
		_w8865_,
		_w8866_,
		_w27923_
	);
	LUT3 #(
		.INIT('h2a)
	) name26023 (
		\m1_data_i[27]_pad ,
		_w8865_,
		_w8866_,
		_w27924_
	);
	LUT4 #(
		.INIT('h67ef)
	) name26024 (
		_w8860_,
		_w8863_,
		_w27923_,
		_w27924_,
		_w27925_
	);
	LUT3 #(
		.INIT('h80)
	) name26025 (
		\m6_data_i[27]_pad ,
		_w8865_,
		_w8866_,
		_w27926_
	);
	LUT3 #(
		.INIT('h2a)
	) name26026 (
		\m5_data_i[27]_pad ,
		_w8865_,
		_w8866_,
		_w27927_
	);
	LUT4 #(
		.INIT('hcdef)
	) name26027 (
		_w8860_,
		_w8863_,
		_w27926_,
		_w27927_,
		_w27928_
	);
	LUT4 #(
		.INIT('h7fff)
	) name26028 (
		_w27919_,
		_w27922_,
		_w27925_,
		_w27928_,
		_w27929_
	);
	LUT3 #(
		.INIT('h2a)
	) name26029 (
		\m3_data_i[28]_pad ,
		_w8865_,
		_w8866_,
		_w27930_
	);
	LUT3 #(
		.INIT('h80)
	) name26030 (
		\m4_data_i[28]_pad ,
		_w8865_,
		_w8866_,
		_w27931_
	);
	LUT4 #(
		.INIT('h9dbf)
	) name26031 (
		_w8860_,
		_w8863_,
		_w27930_,
		_w27931_,
		_w27932_
	);
	LUT3 #(
		.INIT('h80)
	) name26032 (
		\m0_data_i[28]_pad ,
		_w8865_,
		_w8866_,
		_w27933_
	);
	LUT3 #(
		.INIT('h2a)
	) name26033 (
		\m5_data_i[28]_pad ,
		_w8865_,
		_w8866_,
		_w27934_
	);
	LUT4 #(
		.INIT('h5d7f)
	) name26034 (
		_w8860_,
		_w8863_,
		_w27933_,
		_w27934_,
		_w27935_
	);
	LUT3 #(
		.INIT('h2a)
	) name26035 (
		\m7_data_i[28]_pad ,
		_w8865_,
		_w8866_,
		_w27936_
	);
	LUT3 #(
		.INIT('h80)
	) name26036 (
		\m6_data_i[28]_pad ,
		_w8865_,
		_w8866_,
		_w27937_
	);
	LUT3 #(
		.INIT('h57)
	) name26037 (
		_w8878_,
		_w27936_,
		_w27937_,
		_w27938_
	);
	LUT3 #(
		.INIT('h2a)
	) name26038 (
		\m1_data_i[28]_pad ,
		_w8865_,
		_w8866_,
		_w27939_
	);
	LUT3 #(
		.INIT('h80)
	) name26039 (
		\m2_data_i[28]_pad ,
		_w8865_,
		_w8866_,
		_w27940_
	);
	LUT4 #(
		.INIT('h3b7f)
	) name26040 (
		_w8860_,
		_w8863_,
		_w27939_,
		_w27940_,
		_w27941_
	);
	LUT4 #(
		.INIT('h7fff)
	) name26041 (
		_w27932_,
		_w27935_,
		_w27938_,
		_w27941_,
		_w27942_
	);
	LUT3 #(
		.INIT('h2a)
	) name26042 (
		\m1_data_i[29]_pad ,
		_w8865_,
		_w8866_,
		_w27943_
	);
	LUT3 #(
		.INIT('h80)
	) name26043 (
		\m2_data_i[29]_pad ,
		_w8865_,
		_w8866_,
		_w27944_
	);
	LUT4 #(
		.INIT('h3b7f)
	) name26044 (
		_w8860_,
		_w8863_,
		_w27943_,
		_w27944_,
		_w27945_
	);
	LUT3 #(
		.INIT('h2a)
	) name26045 (
		\m3_data_i[29]_pad ,
		_w8865_,
		_w8866_,
		_w27946_
	);
	LUT3 #(
		.INIT('h2a)
	) name26046 (
		\m5_data_i[29]_pad ,
		_w8865_,
		_w8866_,
		_w27947_
	);
	LUT4 #(
		.INIT('h9dbf)
	) name26047 (
		_w8860_,
		_w8863_,
		_w27946_,
		_w27947_,
		_w27948_
	);
	LUT3 #(
		.INIT('h80)
	) name26048 (
		\m4_data_i[29]_pad ,
		_w8865_,
		_w8866_,
		_w27949_
	);
	LUT3 #(
		.INIT('h80)
	) name26049 (
		\m6_data_i[29]_pad ,
		_w8865_,
		_w8866_,
		_w27950_
	);
	LUT4 #(
		.INIT('hcedf)
	) name26050 (
		_w8860_,
		_w8863_,
		_w27949_,
		_w27950_,
		_w27951_
	);
	LUT3 #(
		.INIT('h80)
	) name26051 (
		\m0_data_i[29]_pad ,
		_w8865_,
		_w8866_,
		_w27952_
	);
	LUT3 #(
		.INIT('h2a)
	) name26052 (
		\m7_data_i[29]_pad ,
		_w8865_,
		_w8866_,
		_w27953_
	);
	LUT4 #(
		.INIT('h6e7f)
	) name26053 (
		_w8860_,
		_w8863_,
		_w27952_,
		_w27953_,
		_w27954_
	);
	LUT4 #(
		.INIT('h7fff)
	) name26054 (
		_w27945_,
		_w27948_,
		_w27951_,
		_w27954_,
		_w27955_
	);
	LUT3 #(
		.INIT('h2a)
	) name26055 (
		\m1_data_i[2]_pad ,
		_w8865_,
		_w8866_,
		_w27956_
	);
	LUT3 #(
		.INIT('h80)
	) name26056 (
		\m2_data_i[2]_pad ,
		_w8865_,
		_w8866_,
		_w27957_
	);
	LUT4 #(
		.INIT('h3b7f)
	) name26057 (
		_w8860_,
		_w8863_,
		_w27956_,
		_w27957_,
		_w27958_
	);
	LUT3 #(
		.INIT('h80)
	) name26058 (
		\m6_data_i[2]_pad ,
		_w8865_,
		_w8866_,
		_w27959_
	);
	LUT3 #(
		.INIT('h2a)
	) name26059 (
		\m7_data_i[2]_pad ,
		_w8865_,
		_w8866_,
		_w27960_
	);
	LUT3 #(
		.INIT('h57)
	) name26060 (
		_w8878_,
		_w27959_,
		_w27960_,
		_w27961_
	);
	LUT3 #(
		.INIT('h2a)
	) name26061 (
		\m5_data_i[2]_pad ,
		_w8865_,
		_w8866_,
		_w27962_
	);
	LUT3 #(
		.INIT('h80)
	) name26062 (
		\m0_data_i[2]_pad ,
		_w8865_,
		_w8866_,
		_w27963_
	);
	LUT4 #(
		.INIT('h57df)
	) name26063 (
		_w8860_,
		_w8863_,
		_w27962_,
		_w27963_,
		_w27964_
	);
	LUT3 #(
		.INIT('h2a)
	) name26064 (
		\m3_data_i[2]_pad ,
		_w8865_,
		_w8866_,
		_w27965_
	);
	LUT3 #(
		.INIT('h80)
	) name26065 (
		\m4_data_i[2]_pad ,
		_w8865_,
		_w8866_,
		_w27966_
	);
	LUT4 #(
		.INIT('h9dbf)
	) name26066 (
		_w8860_,
		_w8863_,
		_w27965_,
		_w27966_,
		_w27967_
	);
	LUT4 #(
		.INIT('h7fff)
	) name26067 (
		_w27958_,
		_w27961_,
		_w27964_,
		_w27967_,
		_w27968_
	);
	LUT3 #(
		.INIT('h80)
	) name26068 (
		\m0_data_i[30]_pad ,
		_w8865_,
		_w8866_,
		_w27969_
	);
	LUT3 #(
		.INIT('h2a)
	) name26069 (
		\m7_data_i[30]_pad ,
		_w8865_,
		_w8866_,
		_w27970_
	);
	LUT4 #(
		.INIT('h6e7f)
	) name26070 (
		_w8860_,
		_w8863_,
		_w27969_,
		_w27970_,
		_w27971_
	);
	LUT3 #(
		.INIT('h2a)
	) name26071 (
		\m3_data_i[30]_pad ,
		_w8865_,
		_w8866_,
		_w27972_
	);
	LUT3 #(
		.INIT('h80)
	) name26072 (
		\m2_data_i[30]_pad ,
		_w8865_,
		_w8866_,
		_w27973_
	);
	LUT3 #(
		.INIT('h57)
	) name26073 (
		_w8864_,
		_w27972_,
		_w27973_,
		_w27974_
	);
	LUT3 #(
		.INIT('h80)
	) name26074 (
		\m4_data_i[30]_pad ,
		_w8865_,
		_w8866_,
		_w27975_
	);
	LUT3 #(
		.INIT('h2a)
	) name26075 (
		\m1_data_i[30]_pad ,
		_w8865_,
		_w8866_,
		_w27976_
	);
	LUT4 #(
		.INIT('h57df)
	) name26076 (
		_w8860_,
		_w8863_,
		_w27975_,
		_w27976_,
		_w27977_
	);
	LUT3 #(
		.INIT('h80)
	) name26077 (
		\m6_data_i[30]_pad ,
		_w8865_,
		_w8866_,
		_w27978_
	);
	LUT3 #(
		.INIT('h2a)
	) name26078 (
		\m5_data_i[30]_pad ,
		_w8865_,
		_w8866_,
		_w27979_
	);
	LUT4 #(
		.INIT('hcdef)
	) name26079 (
		_w8860_,
		_w8863_,
		_w27978_,
		_w27979_,
		_w27980_
	);
	LUT4 #(
		.INIT('h7fff)
	) name26080 (
		_w27971_,
		_w27974_,
		_w27977_,
		_w27980_,
		_w27981_
	);
	LUT3 #(
		.INIT('h80)
	) name26081 (
		\m0_data_i[31]_pad ,
		_w8865_,
		_w8866_,
		_w27982_
	);
	LUT3 #(
		.INIT('h2a)
	) name26082 (
		\m7_data_i[31]_pad ,
		_w8865_,
		_w8866_,
		_w27983_
	);
	LUT4 #(
		.INIT('h6e7f)
	) name26083 (
		_w8860_,
		_w8863_,
		_w27982_,
		_w27983_,
		_w27984_
	);
	LUT3 #(
		.INIT('h2a)
	) name26084 (
		\m1_data_i[31]_pad ,
		_w8865_,
		_w8866_,
		_w27985_
	);
	LUT3 #(
		.INIT('h2a)
	) name26085 (
		\m5_data_i[31]_pad ,
		_w8865_,
		_w8866_,
		_w27986_
	);
	LUT4 #(
		.INIT('h5d7f)
	) name26086 (
		_w8860_,
		_w8863_,
		_w27985_,
		_w27986_,
		_w27987_
	);
	LUT3 #(
		.INIT('h80)
	) name26087 (
		\m2_data_i[31]_pad ,
		_w8865_,
		_w8866_,
		_w27988_
	);
	LUT3 #(
		.INIT('h80)
	) name26088 (
		\m6_data_i[31]_pad ,
		_w8865_,
		_w8866_,
		_w27989_
	);
	LUT4 #(
		.INIT('haebf)
	) name26089 (
		_w8860_,
		_w8863_,
		_w27988_,
		_w27989_,
		_w27990_
	);
	LUT3 #(
		.INIT('h2a)
	) name26090 (
		\m3_data_i[31]_pad ,
		_w8865_,
		_w8866_,
		_w27991_
	);
	LUT3 #(
		.INIT('h80)
	) name26091 (
		\m4_data_i[31]_pad ,
		_w8865_,
		_w8866_,
		_w27992_
	);
	LUT4 #(
		.INIT('h9dbf)
	) name26092 (
		_w8860_,
		_w8863_,
		_w27991_,
		_w27992_,
		_w27993_
	);
	LUT4 #(
		.INIT('h7fff)
	) name26093 (
		_w27984_,
		_w27987_,
		_w27990_,
		_w27993_,
		_w27994_
	);
	LUT3 #(
		.INIT('h80)
	) name26094 (
		\m0_data_i[3]_pad ,
		_w8865_,
		_w8866_,
		_w27995_
	);
	LUT3 #(
		.INIT('h2a)
	) name26095 (
		\m7_data_i[3]_pad ,
		_w8865_,
		_w8866_,
		_w27996_
	);
	LUT4 #(
		.INIT('h6e7f)
	) name26096 (
		_w8860_,
		_w8863_,
		_w27995_,
		_w27996_,
		_w27997_
	);
	LUT3 #(
		.INIT('h2a)
	) name26097 (
		\m3_data_i[3]_pad ,
		_w8865_,
		_w8866_,
		_w27998_
	);
	LUT3 #(
		.INIT('h2a)
	) name26098 (
		\m5_data_i[3]_pad ,
		_w8865_,
		_w8866_,
		_w27999_
	);
	LUT4 #(
		.INIT('h9dbf)
	) name26099 (
		_w8860_,
		_w8863_,
		_w27998_,
		_w27999_,
		_w28000_
	);
	LUT3 #(
		.INIT('h80)
	) name26100 (
		\m4_data_i[3]_pad ,
		_w8865_,
		_w8866_,
		_w28001_
	);
	LUT3 #(
		.INIT('h80)
	) name26101 (
		\m6_data_i[3]_pad ,
		_w8865_,
		_w8866_,
		_w28002_
	);
	LUT4 #(
		.INIT('hcedf)
	) name26102 (
		_w8860_,
		_w8863_,
		_w28001_,
		_w28002_,
		_w28003_
	);
	LUT3 #(
		.INIT('h2a)
	) name26103 (
		\m1_data_i[3]_pad ,
		_w8865_,
		_w8866_,
		_w28004_
	);
	LUT3 #(
		.INIT('h80)
	) name26104 (
		\m2_data_i[3]_pad ,
		_w8865_,
		_w8866_,
		_w28005_
	);
	LUT4 #(
		.INIT('h3b7f)
	) name26105 (
		_w8860_,
		_w8863_,
		_w28004_,
		_w28005_,
		_w28006_
	);
	LUT4 #(
		.INIT('h7fff)
	) name26106 (
		_w27997_,
		_w28000_,
		_w28003_,
		_w28006_,
		_w28007_
	);
	LUT3 #(
		.INIT('h2a)
	) name26107 (
		\m1_data_i[4]_pad ,
		_w8865_,
		_w8866_,
		_w28008_
	);
	LUT3 #(
		.INIT('h80)
	) name26108 (
		\m2_data_i[4]_pad ,
		_w8865_,
		_w8866_,
		_w28009_
	);
	LUT4 #(
		.INIT('h3b7f)
	) name26109 (
		_w8860_,
		_w8863_,
		_w28008_,
		_w28009_,
		_w28010_
	);
	LUT3 #(
		.INIT('h80)
	) name26110 (
		\m6_data_i[4]_pad ,
		_w8865_,
		_w8866_,
		_w28011_
	);
	LUT3 #(
		.INIT('h80)
	) name26111 (
		\m4_data_i[4]_pad ,
		_w8865_,
		_w8866_,
		_w28012_
	);
	LUT4 #(
		.INIT('hcdef)
	) name26112 (
		_w8860_,
		_w8863_,
		_w28011_,
		_w28012_,
		_w28013_
	);
	LUT3 #(
		.INIT('h2a)
	) name26113 (
		\m5_data_i[4]_pad ,
		_w8865_,
		_w8866_,
		_w28014_
	);
	LUT3 #(
		.INIT('h2a)
	) name26114 (
		\m3_data_i[4]_pad ,
		_w8865_,
		_w8866_,
		_w28015_
	);
	LUT4 #(
		.INIT('h9bdf)
	) name26115 (
		_w8860_,
		_w8863_,
		_w28014_,
		_w28015_,
		_w28016_
	);
	LUT3 #(
		.INIT('h80)
	) name26116 (
		\m0_data_i[4]_pad ,
		_w8865_,
		_w8866_,
		_w28017_
	);
	LUT3 #(
		.INIT('h2a)
	) name26117 (
		\m7_data_i[4]_pad ,
		_w8865_,
		_w8866_,
		_w28018_
	);
	LUT4 #(
		.INIT('h6e7f)
	) name26118 (
		_w8860_,
		_w8863_,
		_w28017_,
		_w28018_,
		_w28019_
	);
	LUT4 #(
		.INIT('h7fff)
	) name26119 (
		_w28010_,
		_w28013_,
		_w28016_,
		_w28019_,
		_w28020_
	);
	LUT3 #(
		.INIT('h2a)
	) name26120 (
		\m1_data_i[5]_pad ,
		_w8865_,
		_w8866_,
		_w28021_
	);
	LUT3 #(
		.INIT('h80)
	) name26121 (
		\m2_data_i[5]_pad ,
		_w8865_,
		_w8866_,
		_w28022_
	);
	LUT4 #(
		.INIT('h3b7f)
	) name26122 (
		_w8860_,
		_w8863_,
		_w28021_,
		_w28022_,
		_w28023_
	);
	LUT3 #(
		.INIT('h80)
	) name26123 (
		\m0_data_i[5]_pad ,
		_w8865_,
		_w8866_,
		_w28024_
	);
	LUT3 #(
		.INIT('h2a)
	) name26124 (
		\m5_data_i[5]_pad ,
		_w8865_,
		_w8866_,
		_w28025_
	);
	LUT4 #(
		.INIT('h5d7f)
	) name26125 (
		_w8860_,
		_w8863_,
		_w28024_,
		_w28025_,
		_w28026_
	);
	LUT3 #(
		.INIT('h2a)
	) name26126 (
		\m7_data_i[5]_pad ,
		_w8865_,
		_w8866_,
		_w28027_
	);
	LUT3 #(
		.INIT('h80)
	) name26127 (
		\m6_data_i[5]_pad ,
		_w8865_,
		_w8866_,
		_w28028_
	);
	LUT3 #(
		.INIT('h57)
	) name26128 (
		_w8878_,
		_w28027_,
		_w28028_,
		_w28029_
	);
	LUT3 #(
		.INIT('h2a)
	) name26129 (
		\m3_data_i[5]_pad ,
		_w8865_,
		_w8866_,
		_w28030_
	);
	LUT3 #(
		.INIT('h80)
	) name26130 (
		\m4_data_i[5]_pad ,
		_w8865_,
		_w8866_,
		_w28031_
	);
	LUT4 #(
		.INIT('h9dbf)
	) name26131 (
		_w8860_,
		_w8863_,
		_w28030_,
		_w28031_,
		_w28032_
	);
	LUT4 #(
		.INIT('h7fff)
	) name26132 (
		_w28023_,
		_w28026_,
		_w28029_,
		_w28032_,
		_w28033_
	);
	LUT3 #(
		.INIT('h80)
	) name26133 (
		\m6_data_i[6]_pad ,
		_w8865_,
		_w8866_,
		_w28034_
	);
	LUT3 #(
		.INIT('h2a)
	) name26134 (
		\m5_data_i[6]_pad ,
		_w8865_,
		_w8866_,
		_w28035_
	);
	LUT4 #(
		.INIT('hcdef)
	) name26135 (
		_w8860_,
		_w8863_,
		_w28034_,
		_w28035_,
		_w28036_
	);
	LUT3 #(
		.INIT('h80)
	) name26136 (
		\m0_data_i[6]_pad ,
		_w8865_,
		_w8866_,
		_w28037_
	);
	LUT3 #(
		.INIT('h80)
	) name26137 (
		\m2_data_i[6]_pad ,
		_w8865_,
		_w8866_,
		_w28038_
	);
	LUT4 #(
		.INIT('h3b7f)
	) name26138 (
		_w8860_,
		_w8863_,
		_w28037_,
		_w28038_,
		_w28039_
	);
	LUT3 #(
		.INIT('h2a)
	) name26139 (
		\m7_data_i[6]_pad ,
		_w8865_,
		_w8866_,
		_w28040_
	);
	LUT3 #(
		.INIT('h2a)
	) name26140 (
		\m1_data_i[6]_pad ,
		_w8865_,
		_w8866_,
		_w28041_
	);
	LUT4 #(
		.INIT('h67ef)
	) name26141 (
		_w8860_,
		_w8863_,
		_w28040_,
		_w28041_,
		_w28042_
	);
	LUT3 #(
		.INIT('h2a)
	) name26142 (
		\m3_data_i[6]_pad ,
		_w8865_,
		_w8866_,
		_w28043_
	);
	LUT3 #(
		.INIT('h80)
	) name26143 (
		\m4_data_i[6]_pad ,
		_w8865_,
		_w8866_,
		_w28044_
	);
	LUT4 #(
		.INIT('h9dbf)
	) name26144 (
		_w8860_,
		_w8863_,
		_w28043_,
		_w28044_,
		_w28045_
	);
	LUT4 #(
		.INIT('h7fff)
	) name26145 (
		_w28036_,
		_w28039_,
		_w28042_,
		_w28045_,
		_w28046_
	);
	LUT3 #(
		.INIT('h80)
	) name26146 (
		\m6_data_i[7]_pad ,
		_w8865_,
		_w8866_,
		_w28047_
	);
	LUT3 #(
		.INIT('h2a)
	) name26147 (
		\m5_data_i[7]_pad ,
		_w8865_,
		_w8866_,
		_w28048_
	);
	LUT4 #(
		.INIT('hcdef)
	) name26148 (
		_w8860_,
		_w8863_,
		_w28047_,
		_w28048_,
		_w28049_
	);
	LUT3 #(
		.INIT('h2a)
	) name26149 (
		\m1_data_i[7]_pad ,
		_w8865_,
		_w8866_,
		_w28050_
	);
	LUT3 #(
		.INIT('h2a)
	) name26150 (
		\m7_data_i[7]_pad ,
		_w8865_,
		_w8866_,
		_w28051_
	);
	LUT4 #(
		.INIT('h6e7f)
	) name26151 (
		_w8860_,
		_w8863_,
		_w28050_,
		_w28051_,
		_w28052_
	);
	LUT3 #(
		.INIT('h80)
	) name26152 (
		\m2_data_i[7]_pad ,
		_w8865_,
		_w8866_,
		_w28053_
	);
	LUT3 #(
		.INIT('h80)
	) name26153 (
		\m0_data_i[7]_pad ,
		_w8865_,
		_w8866_,
		_w28054_
	);
	LUT4 #(
		.INIT('h37bf)
	) name26154 (
		_w8860_,
		_w8863_,
		_w28053_,
		_w28054_,
		_w28055_
	);
	LUT3 #(
		.INIT('h2a)
	) name26155 (
		\m3_data_i[7]_pad ,
		_w8865_,
		_w8866_,
		_w28056_
	);
	LUT3 #(
		.INIT('h80)
	) name26156 (
		\m4_data_i[7]_pad ,
		_w8865_,
		_w8866_,
		_w28057_
	);
	LUT4 #(
		.INIT('h9dbf)
	) name26157 (
		_w8860_,
		_w8863_,
		_w28056_,
		_w28057_,
		_w28058_
	);
	LUT4 #(
		.INIT('h7fff)
	) name26158 (
		_w28049_,
		_w28052_,
		_w28055_,
		_w28058_,
		_w28059_
	);
	LUT3 #(
		.INIT('h2a)
	) name26159 (
		\m3_data_i[8]_pad ,
		_w8865_,
		_w8866_,
		_w28060_
	);
	LUT3 #(
		.INIT('h80)
	) name26160 (
		\m4_data_i[8]_pad ,
		_w8865_,
		_w8866_,
		_w28061_
	);
	LUT4 #(
		.INIT('h9dbf)
	) name26161 (
		_w8860_,
		_w8863_,
		_w28060_,
		_w28061_,
		_w28062_
	);
	LUT3 #(
		.INIT('h80)
	) name26162 (
		\m6_data_i[8]_pad ,
		_w8865_,
		_w8866_,
		_w28063_
	);
	LUT3 #(
		.INIT('h2a)
	) name26163 (
		\m7_data_i[8]_pad ,
		_w8865_,
		_w8866_,
		_w28064_
	);
	LUT3 #(
		.INIT('h57)
	) name26164 (
		_w8878_,
		_w28063_,
		_w28064_,
		_w28065_
	);
	LUT3 #(
		.INIT('h2a)
	) name26165 (
		\m5_data_i[8]_pad ,
		_w8865_,
		_w8866_,
		_w28066_
	);
	LUT3 #(
		.INIT('h80)
	) name26166 (
		\m0_data_i[8]_pad ,
		_w8865_,
		_w8866_,
		_w28067_
	);
	LUT4 #(
		.INIT('h57df)
	) name26167 (
		_w8860_,
		_w8863_,
		_w28066_,
		_w28067_,
		_w28068_
	);
	LUT3 #(
		.INIT('h2a)
	) name26168 (
		\m1_data_i[8]_pad ,
		_w8865_,
		_w8866_,
		_w28069_
	);
	LUT3 #(
		.INIT('h80)
	) name26169 (
		\m2_data_i[8]_pad ,
		_w8865_,
		_w8866_,
		_w28070_
	);
	LUT4 #(
		.INIT('h3b7f)
	) name26170 (
		_w8860_,
		_w8863_,
		_w28069_,
		_w28070_,
		_w28071_
	);
	LUT4 #(
		.INIT('h7fff)
	) name26171 (
		_w28062_,
		_w28065_,
		_w28068_,
		_w28071_,
		_w28072_
	);
	LUT3 #(
		.INIT('h2a)
	) name26172 (
		\m3_data_i[9]_pad ,
		_w8865_,
		_w8866_,
		_w28073_
	);
	LUT3 #(
		.INIT('h80)
	) name26173 (
		\m4_data_i[9]_pad ,
		_w8865_,
		_w8866_,
		_w28074_
	);
	LUT4 #(
		.INIT('h9dbf)
	) name26174 (
		_w8860_,
		_w8863_,
		_w28073_,
		_w28074_,
		_w28075_
	);
	LUT3 #(
		.INIT('h80)
	) name26175 (
		\m6_data_i[9]_pad ,
		_w8865_,
		_w8866_,
		_w28076_
	);
	LUT3 #(
		.INIT('h80)
	) name26176 (
		\m2_data_i[9]_pad ,
		_w8865_,
		_w8866_,
		_w28077_
	);
	LUT4 #(
		.INIT('habef)
	) name26177 (
		_w8860_,
		_w8863_,
		_w28076_,
		_w28077_,
		_w28078_
	);
	LUT3 #(
		.INIT('h2a)
	) name26178 (
		\m5_data_i[9]_pad ,
		_w8865_,
		_w8866_,
		_w28079_
	);
	LUT3 #(
		.INIT('h2a)
	) name26179 (
		\m1_data_i[9]_pad ,
		_w8865_,
		_w8866_,
		_w28080_
	);
	LUT4 #(
		.INIT('h57df)
	) name26180 (
		_w8860_,
		_w8863_,
		_w28079_,
		_w28080_,
		_w28081_
	);
	LUT3 #(
		.INIT('h80)
	) name26181 (
		\m0_data_i[9]_pad ,
		_w8865_,
		_w8866_,
		_w28082_
	);
	LUT3 #(
		.INIT('h2a)
	) name26182 (
		\m7_data_i[9]_pad ,
		_w8865_,
		_w8866_,
		_w28083_
	);
	LUT4 #(
		.INIT('h6e7f)
	) name26183 (
		_w8860_,
		_w8863_,
		_w28082_,
		_w28083_,
		_w28084_
	);
	LUT4 #(
		.INIT('h7fff)
	) name26184 (
		_w28075_,
		_w28078_,
		_w28081_,
		_w28084_,
		_w28085_
	);
	LUT3 #(
		.INIT('h2a)
	) name26185 (
		\m1_sel_i[0]_pad ,
		_w8865_,
		_w8866_,
		_w28086_
	);
	LUT3 #(
		.INIT('h80)
	) name26186 (
		\m2_sel_i[0]_pad ,
		_w8865_,
		_w8866_,
		_w28087_
	);
	LUT4 #(
		.INIT('h3b7f)
	) name26187 (
		_w8860_,
		_w8863_,
		_w28086_,
		_w28087_,
		_w28088_
	);
	LUT3 #(
		.INIT('h80)
	) name26188 (
		\m6_sel_i[0]_pad ,
		_w8865_,
		_w8866_,
		_w28089_
	);
	LUT3 #(
		.INIT('h80)
	) name26189 (
		\m4_sel_i[0]_pad ,
		_w8865_,
		_w8866_,
		_w28090_
	);
	LUT4 #(
		.INIT('hcdef)
	) name26190 (
		_w8860_,
		_w8863_,
		_w28089_,
		_w28090_,
		_w28091_
	);
	LUT3 #(
		.INIT('h2a)
	) name26191 (
		\m5_sel_i[0]_pad ,
		_w8865_,
		_w8866_,
		_w28092_
	);
	LUT3 #(
		.INIT('h2a)
	) name26192 (
		\m3_sel_i[0]_pad ,
		_w8865_,
		_w8866_,
		_w28093_
	);
	LUT4 #(
		.INIT('h9bdf)
	) name26193 (
		_w8860_,
		_w8863_,
		_w28092_,
		_w28093_,
		_w28094_
	);
	LUT3 #(
		.INIT('h80)
	) name26194 (
		\m0_sel_i[0]_pad ,
		_w8865_,
		_w8866_,
		_w28095_
	);
	LUT3 #(
		.INIT('h2a)
	) name26195 (
		\m7_sel_i[0]_pad ,
		_w8865_,
		_w8866_,
		_w28096_
	);
	LUT4 #(
		.INIT('h6e7f)
	) name26196 (
		_w8860_,
		_w8863_,
		_w28095_,
		_w28096_,
		_w28097_
	);
	LUT4 #(
		.INIT('h7fff)
	) name26197 (
		_w28088_,
		_w28091_,
		_w28094_,
		_w28097_,
		_w28098_
	);
	LUT3 #(
		.INIT('h2a)
	) name26198 (
		\m1_sel_i[1]_pad ,
		_w8865_,
		_w8866_,
		_w28099_
	);
	LUT3 #(
		.INIT('h80)
	) name26199 (
		\m2_sel_i[1]_pad ,
		_w8865_,
		_w8866_,
		_w28100_
	);
	LUT4 #(
		.INIT('h3b7f)
	) name26200 (
		_w8860_,
		_w8863_,
		_w28099_,
		_w28100_,
		_w28101_
	);
	LUT3 #(
		.INIT('h80)
	) name26201 (
		\m6_sel_i[1]_pad ,
		_w8865_,
		_w8866_,
		_w28102_
	);
	LUT3 #(
		.INIT('h2a)
	) name26202 (
		\m7_sel_i[1]_pad ,
		_w8865_,
		_w8866_,
		_w28103_
	);
	LUT3 #(
		.INIT('h57)
	) name26203 (
		_w8878_,
		_w28102_,
		_w28103_,
		_w28104_
	);
	LUT3 #(
		.INIT('h2a)
	) name26204 (
		\m5_sel_i[1]_pad ,
		_w8865_,
		_w8866_,
		_w28105_
	);
	LUT3 #(
		.INIT('h80)
	) name26205 (
		\m0_sel_i[1]_pad ,
		_w8865_,
		_w8866_,
		_w28106_
	);
	LUT4 #(
		.INIT('h57df)
	) name26206 (
		_w8860_,
		_w8863_,
		_w28105_,
		_w28106_,
		_w28107_
	);
	LUT3 #(
		.INIT('h2a)
	) name26207 (
		\m3_sel_i[1]_pad ,
		_w8865_,
		_w8866_,
		_w28108_
	);
	LUT3 #(
		.INIT('h80)
	) name26208 (
		\m4_sel_i[1]_pad ,
		_w8865_,
		_w8866_,
		_w28109_
	);
	LUT4 #(
		.INIT('h9dbf)
	) name26209 (
		_w8860_,
		_w8863_,
		_w28108_,
		_w28109_,
		_w28110_
	);
	LUT4 #(
		.INIT('h7fff)
	) name26210 (
		_w28101_,
		_w28104_,
		_w28107_,
		_w28110_,
		_w28111_
	);
	LUT3 #(
		.INIT('h80)
	) name26211 (
		\m0_sel_i[2]_pad ,
		_w8865_,
		_w8866_,
		_w28112_
	);
	LUT3 #(
		.INIT('h2a)
	) name26212 (
		\m7_sel_i[2]_pad ,
		_w8865_,
		_w8866_,
		_w28113_
	);
	LUT4 #(
		.INIT('h6e7f)
	) name26213 (
		_w8860_,
		_w8863_,
		_w28112_,
		_w28113_,
		_w28114_
	);
	LUT3 #(
		.INIT('h80)
	) name26214 (
		\m6_sel_i[2]_pad ,
		_w8865_,
		_w8866_,
		_w28115_
	);
	LUT3 #(
		.INIT('h80)
	) name26215 (
		\m4_sel_i[2]_pad ,
		_w8865_,
		_w8866_,
		_w28116_
	);
	LUT4 #(
		.INIT('hcdef)
	) name26216 (
		_w8860_,
		_w8863_,
		_w28115_,
		_w28116_,
		_w28117_
	);
	LUT3 #(
		.INIT('h2a)
	) name26217 (
		\m5_sel_i[2]_pad ,
		_w8865_,
		_w8866_,
		_w28118_
	);
	LUT3 #(
		.INIT('h2a)
	) name26218 (
		\m3_sel_i[2]_pad ,
		_w8865_,
		_w8866_,
		_w28119_
	);
	LUT4 #(
		.INIT('h9bdf)
	) name26219 (
		_w8860_,
		_w8863_,
		_w28118_,
		_w28119_,
		_w28120_
	);
	LUT3 #(
		.INIT('h2a)
	) name26220 (
		\m1_sel_i[2]_pad ,
		_w8865_,
		_w8866_,
		_w28121_
	);
	LUT3 #(
		.INIT('h80)
	) name26221 (
		\m2_sel_i[2]_pad ,
		_w8865_,
		_w8866_,
		_w28122_
	);
	LUT4 #(
		.INIT('h3b7f)
	) name26222 (
		_w8860_,
		_w8863_,
		_w28121_,
		_w28122_,
		_w28123_
	);
	LUT4 #(
		.INIT('h7fff)
	) name26223 (
		_w28114_,
		_w28117_,
		_w28120_,
		_w28123_,
		_w28124_
	);
	LUT3 #(
		.INIT('h2a)
	) name26224 (
		\m1_sel_i[3]_pad ,
		_w8865_,
		_w8866_,
		_w28125_
	);
	LUT3 #(
		.INIT('h80)
	) name26225 (
		\m2_sel_i[3]_pad ,
		_w8865_,
		_w8866_,
		_w28126_
	);
	LUT4 #(
		.INIT('h3b7f)
	) name26226 (
		_w8860_,
		_w8863_,
		_w28125_,
		_w28126_,
		_w28127_
	);
	LUT3 #(
		.INIT('h80)
	) name26227 (
		\m0_sel_i[3]_pad ,
		_w8865_,
		_w8866_,
		_w28128_
	);
	LUT3 #(
		.INIT('h80)
	) name26228 (
		\m4_sel_i[3]_pad ,
		_w8865_,
		_w8866_,
		_w28129_
	);
	LUT4 #(
		.INIT('h5d7f)
	) name26229 (
		_w8860_,
		_w8863_,
		_w28128_,
		_w28129_,
		_w28130_
	);
	LUT3 #(
		.INIT('h2a)
	) name26230 (
		\m7_sel_i[3]_pad ,
		_w8865_,
		_w8866_,
		_w28131_
	);
	LUT3 #(
		.INIT('h2a)
	) name26231 (
		\m3_sel_i[3]_pad ,
		_w8865_,
		_w8866_,
		_w28132_
	);
	LUT4 #(
		.INIT('habef)
	) name26232 (
		_w8860_,
		_w8863_,
		_w28131_,
		_w28132_,
		_w28133_
	);
	LUT3 #(
		.INIT('h80)
	) name26233 (
		\m6_sel_i[3]_pad ,
		_w8865_,
		_w8866_,
		_w28134_
	);
	LUT3 #(
		.INIT('h2a)
	) name26234 (
		\m5_sel_i[3]_pad ,
		_w8865_,
		_w8866_,
		_w28135_
	);
	LUT4 #(
		.INIT('hcdef)
	) name26235 (
		_w8860_,
		_w8863_,
		_w28134_,
		_w28135_,
		_w28136_
	);
	LUT4 #(
		.INIT('h7fff)
	) name26236 (
		_w28127_,
		_w28130_,
		_w28133_,
		_w28136_,
		_w28137_
	);
	LUT4 #(
		.INIT('h2a00)
	) name26237 (
		\m3_stb_i_pad ,
		_w8865_,
		_w8866_,
		_w9506_,
		_w28138_
	);
	LUT4 #(
		.INIT('h8000)
	) name26238 (
		\m2_stb_i_pad ,
		_w8865_,
		_w8866_,
		_w9477_,
		_w28139_
	);
	LUT3 #(
		.INIT('h57)
	) name26239 (
		_w8864_,
		_w28138_,
		_w28139_,
		_w28140_
	);
	LUT4 #(
		.INIT('h8000)
	) name26240 (
		\m6_stb_i_pad ,
		_w8865_,
		_w8866_,
		_w9591_,
		_w28141_
	);
	LUT4 #(
		.INIT('h2a00)
	) name26241 (
		\m1_stb_i_pad ,
		_w8865_,
		_w8866_,
		_w9448_,
		_w28142_
	);
	LUT4 #(
		.INIT('h67ef)
	) name26242 (
		_w8860_,
		_w8863_,
		_w28141_,
		_w28142_,
		_w28143_
	);
	LUT4 #(
		.INIT('h2a00)
	) name26243 (
		\m7_stb_i_pad ,
		_w8865_,
		_w8866_,
		_w9327_,
		_w28144_
	);
	LUT4 #(
		.INIT('h2a00)
	) name26244 (
		\m5_stb_i_pad ,
		_w8865_,
		_w8866_,
		_w9556_,
		_w28145_
	);
	LUT4 #(
		.INIT('hcdef)
	) name26245 (
		_w8860_,
		_w8863_,
		_w28144_,
		_w28145_,
		_w28146_
	);
	LUT4 #(
		.INIT('h8000)
	) name26246 (
		\m4_stb_i_pad ,
		_w8865_,
		_w8866_,
		_w9357_,
		_w28147_
	);
	LUT4 #(
		.INIT('h8000)
	) name26247 (
		\m0_stb_i_pad ,
		_w8865_,
		_w8866_,
		_w9641_,
		_w28148_
	);
	LUT4 #(
		.INIT('h57df)
	) name26248 (
		_w8860_,
		_w8863_,
		_w28147_,
		_w28148_,
		_w28149_
	);
	LUT4 #(
		.INIT('h7fff)
	) name26249 (
		_w28140_,
		_w28143_,
		_w28146_,
		_w28149_,
		_w28150_
	);
	LUT3 #(
		.INIT('h2a)
	) name26250 (
		\m3_we_i_pad ,
		_w8865_,
		_w8866_,
		_w28151_
	);
	LUT3 #(
		.INIT('h80)
	) name26251 (
		\m4_we_i_pad ,
		_w8865_,
		_w8866_,
		_w28152_
	);
	LUT4 #(
		.INIT('h9dbf)
	) name26252 (
		_w8860_,
		_w8863_,
		_w28151_,
		_w28152_,
		_w28153_
	);
	LUT3 #(
		.INIT('h80)
	) name26253 (
		\m6_we_i_pad ,
		_w8865_,
		_w8866_,
		_w28154_
	);
	LUT3 #(
		.INIT('h80)
	) name26254 (
		\m2_we_i_pad ,
		_w8865_,
		_w8866_,
		_w28155_
	);
	LUT4 #(
		.INIT('habef)
	) name26255 (
		_w8860_,
		_w8863_,
		_w28154_,
		_w28155_,
		_w28156_
	);
	LUT3 #(
		.INIT('h2a)
	) name26256 (
		\m5_we_i_pad ,
		_w8865_,
		_w8866_,
		_w28157_
	);
	LUT3 #(
		.INIT('h2a)
	) name26257 (
		\m1_we_i_pad ,
		_w8865_,
		_w8866_,
		_w28158_
	);
	LUT4 #(
		.INIT('h57df)
	) name26258 (
		_w8860_,
		_w8863_,
		_w28157_,
		_w28158_,
		_w28159_
	);
	LUT3 #(
		.INIT('h80)
	) name26259 (
		\m0_we_i_pad ,
		_w8865_,
		_w8866_,
		_w28160_
	);
	LUT3 #(
		.INIT('h2a)
	) name26260 (
		\m7_we_i_pad ,
		_w8865_,
		_w8866_,
		_w28161_
	);
	LUT4 #(
		.INIT('h6e7f)
	) name26261 (
		_w8860_,
		_w8863_,
		_w28160_,
		_w28161_,
		_w28162_
	);
	LUT4 #(
		.INIT('h7fff)
	) name26262 (
		_w28153_,
		_w28156_,
		_w28159_,
		_w28162_,
		_w28163_
	);
	assign \_al_n0  = 1'b0;
	assign \_al_n1  = 1'b1;
	assign \g106655/_1_  = _w2099_ ;
	assign \g106703/_1_  = _w1955_ ;
	assign \g69412/_0_  = _w2110_ ;
	assign \g69413/_0_  = _w2121_ ;
	assign \g69417/_1_  = _w2132_ ;
	assign \g69418/_0_  = _w2143_ ;
	assign \g69420/_1_  = _w2154_ ;
	assign \g69421/_0_  = _w2165_ ;
	assign \g69423/_1_  = _w2176_ ;
	assign \g69424/_0_  = _w2187_ ;
	assign \g69426/_1_  = _w2198_ ;
	assign \g69428/_1_  = _w2209_ ;
	assign \g69430/_1_  = _w2220_ ;
	assign \g69432/_1_  = _w2231_ ;
	assign \g69434/_1_  = _w2242_ ;
	assign \g69436/_1_  = _w2253_ ;
	assign \g69438/_1_  = _w2264_ ;
	assign \g69757/_2_  = _w2301_ ;
	assign \g69758/_2_  = _w2338_ ;
	assign \g69759/_2_  = _w2375_ ;
	assign \g69760/_2_  = _w2412_ ;
	assign \g69761/_0_  = _w2458_ ;
	assign \g69762/_2_  = _w2495_ ;
	assign \g69763/_2_  = _w2532_ ;
	assign \g69764/_2_  = _w2569_ ;
	assign \g69765/_2_  = _w2606_ ;
	assign \g69766/_2_  = _w2643_ ;
	assign \g69767/_0_  = _w2682_ ;
	assign \g69768/_0_  = _w2721_ ;
	assign \g69769/_0_  = _w2760_ ;
	assign \g69770/_0_  = _w2799_ ;
	assign \g69771/_0_  = _w2838_ ;
	assign \g69772/_0_  = _w2877_ ;
	assign \g70206/_0_  = _w2919_ ;
	assign \g70392/_0_  = _w2930_ ;
	assign \g70393/_0_  = _w2942_ ;
	assign \g70394/_0_  = _w2972_ ;
	assign \g70395/_0_  = _w3002_ ;
	assign \g70396/_0_  = _w3032_ ;
	assign \g70397/_0_  = _w3054_ ;
	assign \g70398/_0_  = _w3086_ ;
	assign \g70399/_0_  = _w3108_ ;
	assign \g70400/_0_  = _w3130_ ;
	assign \g70401/_0_  = _w3152_ ;
	assign \g70402/_0_  = _w3182_ ;
	assign \g70403/_0_  = _w3204_ ;
	assign \g70404/_0_  = _w3236_ ;
	assign \g70405/_0_  = _w3266_ ;
	assign \g70406/_0_  = _w3298_ ;
	assign \g70407/_0_  = _w3320_ ;
	assign \g70408/_0_  = _w3352_ ;
	assign \g70409/_0_  = _w3384_ ;
	assign \g70410/_0_  = _w3406_ ;
	assign \g70411/_0_  = _w3436_ ;
	assign \g70412/_0_  = _w3466_ ;
	assign \g70413/_0_  = _w3496_ ;
	assign \g70414/_0_  = _w3528_ ;
	assign \g70415/_0_  = _w3558_ ;
	assign \g70416/_0_  = _w3583_ ;
	assign \g70417/_0_  = _w3618_ ;
	assign \g70418/_0_  = _w3644_ ;
	assign \g70419/_0_  = _w3669_ ;
	assign \g70420/_0_  = _w3695_ ;
	assign \g70421/_0_  = _w3721_ ;
	assign \g70422/_0_  = _w3746_ ;
	assign \g70423/_0_  = _w3775_ ;
	assign \g70424/_0_  = _w3801_ ;
	assign \g70425/_0_  = _w3832_ ;
	assign \g70426/_0_  = _w3863_ ;
	assign \g70427/_0_  = _w3889_ ;
	assign \g70428/_0_  = _w3920_ ;
	assign \g70429/_0_  = _w3951_ ;
	assign \g70430/_0_  = _w3982_ ;
	assign \g70431/_0_  = _w4025_ ;
	assign \g70432/_0_  = _w4080_ ;
	assign \g70433/_0_  = _w4121_ ;
	assign \g70434/_0_  = _w4169_ ;
	assign \g70435/_0_  = _w4201_ ;
	assign \g70436/_0_  = _w4244_ ;
	assign \g70437/_0_  = _w4286_ ;
	assign \g70438/_0_  = _w4334_ ;
	assign \g70439/_0_  = _w4363_ ;
	assign \g70440/_0_  = _w4418_ ;
	assign \g70441/_0_  = _w4459_ ;
	assign \g70442/_0_  = _w4507_ ;
	assign \g70443/_0_  = _w4550_ ;
	assign \g70444/_0_  = _w4599_ ;
	assign \g70445/_0_  = _w4640_ ;
	assign \g70446/_0_  = _w4688_ ;
	assign \g70447/_0_  = _w4726_ ;
	assign \g70448/_0_  = _w4767_ ;
	assign \g70449/_0_  = _w4809_ ;
	assign \g70450/_0_  = _w4837_ ;
	assign \g70451/_0_  = _w4884_ ;
	assign \g70452/_0_  = _w4895_ ;
	assign \g70453/_0_  = _w4939_ ;
	assign \g70454/_0_  = _w4978_ ;
	assign \g70455/_0_  = _w5016_ ;
	assign \g70456/_0_  = _w5059_ ;
	assign \g70457/_0_  = _w5101_ ;
	assign \g70458/_0_  = _w5140_ ;
	assign \g70459/_0_  = _w5183_ ;
	assign \g70460/_0_  = _w5232_ ;
	assign \g70461/_0_  = _w5273_ ;
	assign \g70462/_0_  = _w5321_ ;
	assign \g70463/_0_  = _w5363_ ;
	assign \g70464/_0_  = _w5406_ ;
	assign \g70465/_0_  = _w5448_ ;
	assign \g70466/_0_  = _w5496_ ;
	assign \g70467/_0_  = _w5534_ ;
	assign \g70468/_0_  = _w5583_ ;
	assign \g70469/_0_  = _w5625_ ;
	assign \g70470/_0_  = _w5673_ ;
	assign \g70471/_0_  = _w5703_ ;
	assign \g70472/_0_  = _w5746_ ;
	assign \g70473/_0_  = _w5787_ ;
	assign \g70474/_0_  = _w5835_ ;
	assign \g70475/_0_  = _w5865_ ;
	assign \g70476/_0_  = _w5908_ ;
	assign \g70477/_0_  = _w5949_ ;
	assign \g70478/_0_  = _w5988_ ;
	assign \g70479/_0_  = _w6037_ ;
	assign \g70480/_0_  = _w6092_ ;
	assign \g70481/_0_  = _w6133_ ;
	assign \g70482/_0_  = _w6181_ ;
	assign \g70483/_0_  = _w6211_ ;
	assign \g70484/_0_  = _w6254_ ;
	assign \g70485/_0_  = _w6296_ ;
	assign \g70486/_0_  = _w6335_ ;
	assign \g70487/_0_  = _w6365_ ;
	assign \g70488/_0_  = _w6420_ ;
	assign \g70489/_0_  = _w6469_ ;
	assign \g70490/_0_  = _w6508_ ;
	assign \g70491/_0_  = _w6538_ ;
	assign \g70492/_0_  = _w6581_ ;
	assign \g70493/_0_  = _w6622_ ;
	assign \g70494/_0_  = _w6661_ ;
	assign \g70495/_0_  = _w6679_ ;
	assign \g70496/_0_  = _w6697_ ;
	assign \g70497/_0_  = _w6712_ ;
	assign \g70498/_0_  = _w6727_ ;
	assign \g70499/_0_  = _w6742_ ;
	assign \g70500/_0_  = _w6760_ ;
	assign \g70501/_0_  = _w6778_ ;
	assign \g70502/_0_  = _w6793_ ;
	assign \g70503/_0_  = _w6803_ ;
	assign \g70504/_0_  = _w6823_ ;
	assign \g70505/_0_  = _w6843_ ;
	assign \g70506/_0_  = _w6863_ ;
	assign \g70507/_0_  = _w6883_ ;
	assign \g70508/_0_  = _w6933_ ;
	assign \g70509/_0_  = _w6950_ ;
	assign \g70510/_0_  = _w6964_ ;
	assign \g70511/_0_  = _w6982_ ;
	assign \g70513/_0_  = _w6992_ ;
	assign \g70515/_0_  = _w7002_ ;
	assign \g70516/_0_  = _w7022_ ;
	assign \g70517/_0_  = _w7042_ ;
	assign \g70518/_0_  = _w7062_ ;
	assign \g70519/_0_  = _w7082_ ;
	assign \g70521/_0_  = _w7092_ ;
	assign \g70522/_0_  = _w7112_ ;
	assign \g70524/_0_  = _w7122_ ;
	assign \g70557/_0_  = _w7132_ ;
	assign \g70559/_0_  = _w7158_ ;
	assign \g70560/_0_  = _w7179_ ;
	assign \g70561/_0_  = _w7206_ ;
	assign \g70562/_0_  = _w7229_ ;
	assign \g70563/_0_  = _w7255_ ;
	assign \g70564/_0_  = _w7276_ ;
	assign \g70565/_0_  = _w7297_ ;
	assign \g70566/_0_  = _w7318_ ;
	assign \g70567/_0_  = _w7339_ ;
	assign \g70568/_0_  = _w7362_ ;
	assign \g70569/_0_  = _w7389_ ;
	assign \g70570/_0_  = _w7412_ ;
	assign \g70571/_0_  = _w7433_ ;
	assign \g70572/_0_  = _w7454_ ;
	assign \g70573/_0_  = _w7481_ ;
	assign \g70574/_0_  = _w7504_ ;
	assign \g70575/_0_  = _w7525_ ;
	assign \g70576/_0_  = _w7548_ ;
	assign \g70577/_0_  = _w7575_ ;
	assign \g70578/_0_  = _w7596_ ;
	assign \g70579/_0_  = _w7623_ ;
	assign \g70580/_0_  = _w7644_ ;
	assign \g70581/_0_  = _w7670_ ;
	assign \g70582/_0_  = _w7691_ ;
	assign \g70583/_0_  = _w7718_ ;
	assign \g70584/_0_  = _w7741_ ;
	assign \g70585/_0_  = _w7767_ ;
	assign \g70586/_0_  = _w7788_ ;
	assign \g70587/_0_  = _w7815_ ;
	assign \g70588/_0_  = _w7836_ ;
	assign \g70589/_0_  = _w7861_ ;
	assign \g70590/_0_  = _w7881_ ;
	assign \g70591/_0_  = _w7902_ ;
	assign \g70592/_0_  = _w7927_ ;
	assign \g70593/_0_  = _w7945_ ;
	assign \g70594/_0_  = _w7971_ ;
	assign \g70595/_0_  = _w7989_ ;
	assign \g70596/_0_  = _w8014_ ;
	assign \g70597/_0_  = _w8040_ ;
	assign \g70598/_0_  = _w8058_ ;
	assign \g70599/_0_  = _w8072_ ;
	assign \g70600/_0_  = _w8086_ ;
	assign \g70601/_0_  = _w8105_ ;
	assign \g70602/_0_  = _w8119_ ;
	assign \g70603/_0_  = _w8133_ ;
	assign \g70604/_0_  = _w8147_ ;
	assign \g70605/_0_  = _w8149_ ;
	assign \g70606/_0_  = _w8164_ ;
	assign \g70607/_0_  = _w8179_ ;
	assign \g70608/_0_  = _w8194_ ;
	assign \g70609/_0_  = _w8209_ ;
	assign \g70610/_0_  = _w8224_ ;
	assign \g70611/_0_  = _w8239_ ;
	assign \g70612/_0_  = _w8254_ ;
	assign \g70613/_0_  = _w8269_ ;
	assign \g70614/_0_  = _w8284_ ;
	assign \g70615/_0_  = _w8299_ ;
	assign \g70616/_0_  = _w8314_ ;
	assign \g70617/_0_  = _w8329_ ;
	assign \g70618/_0_  = _w8344_ ;
	assign \g70619/_0_  = _w8359_ ;
	assign \g70620/_0_  = _w8374_ ;
	assign \g70621/_0_  = _w8389_ ;
	assign \g70622/_0_  = _w8390_ ;
	assign \g70623/_0_  = _w8391_ ;
	assign \g70624/_0_  = _w8392_ ;
	assign \g70625/_0_  = _w8393_ ;
	assign \g70626/_0_  = _w8394_ ;
	assign \g70627/_0_  = _w8395_ ;
	assign \g70628/_0_  = _w8396_ ;
	assign \g70629/_0_  = _w8397_ ;
	assign \g70630/_0_  = _w8398_ ;
	assign \g70631/_0_  = _w8399_ ;
	assign \g70632/_0_  = _w8400_ ;
	assign \g70633/_0_  = _w8401_ ;
	assign \g70634/_0_  = _w8402_ ;
	assign \g70635/_0_  = _w8403_ ;
	assign \g70636/_0_  = _w8404_ ;
	assign \g70637/_0_  = _w8405_ ;
	assign \g70638/_0_  = _w8406_ ;
	assign \g70639/_0_  = _w8407_ ;
	assign \g70640/_0_  = _w8408_ ;
	assign \g70641/_0_  = _w8409_ ;
	assign \g70642/_0_  = _w8410_ ;
	assign \g70643/_0_  = _w8411_ ;
	assign \g70644/_0_  = _w8412_ ;
	assign \g70645/_0_  = _w8413_ ;
	assign \g70646/_0_  = _w8414_ ;
	assign \g70647/_0_  = _w8415_ ;
	assign \g70648/_0_  = _w8416_ ;
	assign \g70649/_0_  = _w8417_ ;
	assign \g70650/_0_  = _w8418_ ;
	assign \g70651/_0_  = _w8419_ ;
	assign \g70652/_0_  = _w8420_ ;
	assign \g70653/_0_  = _w8421_ ;
	assign \g70654/_0_  = _w8422_ ;
	assign \g70655/_0_  = _w8423_ ;
	assign \g70656/_0_  = _w8424_ ;
	assign \g70657/_0_  = _w8425_ ;
	assign \g70658/_0_  = _w8426_ ;
	assign \g70659/_0_  = _w8427_ ;
	assign \g70660/_0_  = _w8428_ ;
	assign \g70661/_0_  = _w8429_ ;
	assign \g70662/_0_  = _w8430_ ;
	assign \g70663/_0_  = _w8431_ ;
	assign \g70664/_0_  = _w8432_ ;
	assign \g70665/_0_  = _w8433_ ;
	assign \g70666/_0_  = _w8434_ ;
	assign \g70667/_0_  = _w8435_ ;
	assign \g70668/_0_  = _w8436_ ;
	assign \g70669/_0_  = _w8437_ ;
	assign \g70670/_0_  = _w8438_ ;
	assign \g70671/_0_  = _w8439_ ;
	assign \g70672/_0_  = _w8440_ ;
	assign \g70673/_0_  = _w8441_ ;
	assign \g70674/_0_  = _w8442_ ;
	assign \g70675/_0_  = _w8443_ ;
	assign \g70676/_0_  = _w8444_ ;
	assign \g70677/_0_  = _w8445_ ;
	assign \g70678/_0_  = _w8446_ ;
	assign \g70679/_0_  = _w8447_ ;
	assign \g70680/_0_  = _w8448_ ;
	assign \g70681/_0_  = _w8449_ ;
	assign \g70682/_0_  = _w8450_ ;
	assign \g70683/_0_  = _w8451_ ;
	assign \g70684/_0_  = _w8452_ ;
	assign \g70685/_0_  = _w8453_ ;
	assign \g70686/_0_  = _w8454_ ;
	assign \g70687/_0_  = _w8455_ ;
	assign \g70688/_0_  = _w8456_ ;
	assign \g70689/_0_  = _w8457_ ;
	assign \g70690/_0_  = _w8458_ ;
	assign \g70691/_0_  = _w8459_ ;
	assign \g70692/_0_  = _w8460_ ;
	assign \g70693/_0_  = _w8461_ ;
	assign \g70694/_0_  = _w8462_ ;
	assign \g70695/_0_  = _w8463_ ;
	assign \g70696/_0_  = _w8464_ ;
	assign \g70697/_0_  = _w8465_ ;
	assign \g70698/_0_  = _w8466_ ;
	assign \g70699/_0_  = _w8467_ ;
	assign \g70700/_0_  = _w8468_ ;
	assign \g70701/_0_  = _w8469_ ;
	assign \g70702/_0_  = _w8470_ ;
	assign \g70703/_0_  = _w8471_ ;
	assign \g70704/_0_  = _w8472_ ;
	assign \g70705/_0_  = _w8473_ ;
	assign \g70706/_0_  = _w8474_ ;
	assign \g70707/_0_  = _w8475_ ;
	assign \g70708/_0_  = _w8476_ ;
	assign \g70709/_0_  = _w8477_ ;
	assign \g70710/_0_  = _w8478_ ;
	assign \g70711/_0_  = _w8479_ ;
	assign \g70712/_0_  = _w8480_ ;
	assign \g70713/_0_  = _w8481_ ;
	assign \g70714/_0_  = _w8482_ ;
	assign \g70715/_0_  = _w8483_ ;
	assign \g70716/_0_  = _w8484_ ;
	assign \g70717/_0_  = _w8485_ ;
	assign \g70718/_0_  = _w8486_ ;
	assign \g70719/_0_  = _w8487_ ;
	assign \g70720/_0_  = _w8488_ ;
	assign \g70721/_0_  = _w8489_ ;
	assign \g70722/_0_  = _w8490_ ;
	assign \g70723/_0_  = _w8491_ ;
	assign \g70724/_0_  = _w8492_ ;
	assign \g70725/_0_  = _w8493_ ;
	assign \g70726/_0_  = _w8494_ ;
	assign \g70727/_0_  = _w8495_ ;
	assign \g70728/_0_  = _w8496_ ;
	assign \g70729/_0_  = _w8497_ ;
	assign \g70730/_0_  = _w8498_ ;
	assign \g70731/_0_  = _w8499_ ;
	assign \g70732/_0_  = _w8500_ ;
	assign \g70733/_0_  = _w8501_ ;
	assign \g70734/_0_  = _w8502_ ;
	assign \g70735/_0_  = _w8503_ ;
	assign \g70736/_0_  = _w8504_ ;
	assign \g70737/_0_  = _w8505_ ;
	assign \g70738/_0_  = _w8506_ ;
	assign \g70739/_0_  = _w8507_ ;
	assign \g70740/_0_  = _w8508_ ;
	assign \g70741/_0_  = _w8509_ ;
	assign \g70742/_0_  = _w8510_ ;
	assign \g70743/_0_  = _w8511_ ;
	assign \g70744/_0_  = _w8512_ ;
	assign \g70745/_0_  = _w8513_ ;
	assign \g70746/_0_  = _w8514_ ;
	assign \g70747/_0_  = _w8515_ ;
	assign \g70748/_0_  = _w8516_ ;
	assign \g70749/_0_  = _w8517_ ;
	assign \g70750/_0_  = _w8518_ ;
	assign \g70751/_0_  = _w8519_ ;
	assign \g70752/_0_  = _w8520_ ;
	assign \g70753/_0_  = _w8521_ ;
	assign \g70754/_0_  = _w8522_ ;
	assign \g70755/_0_  = _w8523_ ;
	assign \g70756/_0_  = _w8524_ ;
	assign \g70757/_0_  = _w8525_ ;
	assign \g70758/_0_  = _w8526_ ;
	assign \g70759/_0_  = _w8527_ ;
	assign \g70760/_0_  = _w8528_ ;
	assign \g70761/_0_  = _w8529_ ;
	assign \g70762/_0_  = _w8530_ ;
	assign \g70763/_0_  = _w8531_ ;
	assign \g70764/_0_  = _w8532_ ;
	assign \g70765/_0_  = _w8533_ ;
	assign \g70766/_0_  = _w8534_ ;
	assign \g70767/_0_  = _w8535_ ;
	assign \g70768/_0_  = _w8536_ ;
	assign \g70769/_0_  = _w8537_ ;
	assign \g70770/_0_  = _w8538_ ;
	assign \g70771/_0_  = _w8539_ ;
	assign \g70772/_0_  = _w8540_ ;
	assign \g70773/_0_  = _w8541_ ;
	assign \g70774/_0_  = _w8542_ ;
	assign \g70775/_0_  = _w8543_ ;
	assign \g70776/_0_  = _w8544_ ;
	assign \g70777/_0_  = _w8545_ ;
	assign \g70778/_0_  = _w8546_ ;
	assign \g70779/_0_  = _w8547_ ;
	assign \g70780/_0_  = _w8548_ ;
	assign \g70781/_0_  = _w8549_ ;
	assign \g70782/_0_  = _w8550_ ;
	assign \g70783/_0_  = _w8551_ ;
	assign \g70784/_0_  = _w8552_ ;
	assign \g70785/_0_  = _w8553_ ;
	assign \g70786/_0_  = _w8554_ ;
	assign \g70787/_0_  = _w8555_ ;
	assign \g70788/_0_  = _w8556_ ;
	assign \g70789/_0_  = _w8557_ ;
	assign \g70790/_0_  = _w8558_ ;
	assign \g70791/_0_  = _w8559_ ;
	assign \g70792/_0_  = _w8560_ ;
	assign \g70793/_0_  = _w8561_ ;
	assign \g70794/_0_  = _w8562_ ;
	assign \g70795/_0_  = _w8563_ ;
	assign \g70796/_0_  = _w8564_ ;
	assign \g70797/_0_  = _w8565_ ;
	assign \g70798/_0_  = _w8566_ ;
	assign \g70799/_0_  = _w8567_ ;
	assign \g70800/_0_  = _w8568_ ;
	assign \g70801/_0_  = _w8569_ ;
	assign \g70802/_0_  = _w8570_ ;
	assign \g70803/_0_  = _w8571_ ;
	assign \g70804/_0_  = _w8572_ ;
	assign \g70805/_0_  = _w8573_ ;
	assign \g70806/_0_  = _w8574_ ;
	assign \g70807/_0_  = _w8575_ ;
	assign \g70808/_0_  = _w8576_ ;
	assign \g70809/_0_  = _w8577_ ;
	assign \g70810/_0_  = _w8578_ ;
	assign \g70811/_0_  = _w8579_ ;
	assign \g70812/_0_  = _w8580_ ;
	assign \g70813/_0_  = _w8581_ ;
	assign \g70814/_0_  = _w8582_ ;
	assign \g70815/_0_  = _w8583_ ;
	assign \g70816/_0_  = _w8584_ ;
	assign \g70817/_0_  = _w8585_ ;
	assign \g70818/_0_  = _w8586_ ;
	assign \g70819/_0_  = _w8587_ ;
	assign \g70820/_0_  = _w8588_ ;
	assign \g70821/_0_  = _w8589_ ;
	assign \g70822/_0_  = _w8590_ ;
	assign \g70823/_0_  = _w8591_ ;
	assign \g70824/_0_  = _w8592_ ;
	assign \g70825/_0_  = _w8593_ ;
	assign \g70826/_0_  = _w8594_ ;
	assign \g70827/_0_  = _w8595_ ;
	assign \g70828/_0_  = _w8596_ ;
	assign \g70829/_0_  = _w8597_ ;
	assign \g70830/_0_  = _w8598_ ;
	assign \g70831/_0_  = _w8599_ ;
	assign \g70832/_0_  = _w8600_ ;
	assign \g70833/_0_  = _w8601_ ;
	assign \g70834/_0_  = _w8602_ ;
	assign \g70835/_0_  = _w8603_ ;
	assign \g70836/_0_  = _w8604_ ;
	assign \g70837/_0_  = _w8605_ ;
	assign \g70838/_0_  = _w8606_ ;
	assign \g70839/_0_  = _w8607_ ;
	assign \g70840/_0_  = _w8608_ ;
	assign \g70841/_0_  = _w8609_ ;
	assign \g70842/_0_  = _w8610_ ;
	assign \g70843/_0_  = _w8611_ ;
	assign \g70844/_0_  = _w8612_ ;
	assign \g70845/_0_  = _w8613_ ;
	assign \g70846/_0_  = _w8614_ ;
	assign \g70847/_0_  = _w8615_ ;
	assign \g70848/_0_  = _w8616_ ;
	assign \g70849/_0_  = _w8617_ ;
	assign \g70850/_0_  = _w8618_ ;
	assign \g70851/_0_  = _w8619_ ;
	assign \g70852/_0_  = _w8620_ ;
	assign \g70853/_0_  = _w8621_ ;
	assign \g70854/_0_  = _w8622_ ;
	assign \g70855/_0_  = _w8623_ ;
	assign \g70856/_0_  = _w8624_ ;
	assign \g70857/_0_  = _w8625_ ;
	assign \g70858/_0_  = _w8626_ ;
	assign \g70859/_0_  = _w8627_ ;
	assign \g70860/_0_  = _w8628_ ;
	assign \g70861/_0_  = _w8629_ ;
	assign \g71404/_0_  = _w8631_ ;
	assign \g71407/_0_  = _w8647_ ;
	assign \g72631/_0_  = _w8680_ ;
	assign \g72631/_1_  = _w8681_ ;
	assign \g72633/_0_  = _w8686_ ;
	assign \g72642/_0_  = _w8691_ ;
	assign \g72649/_0_  = _w8724_ ;
	assign \g72649/_1_  = _w8725_ ;
	assign \g72652/_0_  = _w8730_ ;
	assign \g72660/_0_  = _w8735_ ;
	assign \g72666/_0_  = _w8768_ ;
	assign \g72666/_1_  = _w8769_ ;
	assign \g72671/_0_  = _w8774_ ;
	assign \g72681/_0_  = _w8807_ ;
	assign \g72681/_1_  = _w8808_ ;
	assign \g72689/_0_  = _w8813_ ;
	assign \g72696/_0_  = _w8846_ ;
	assign \g72696/_1_  = _w8847_ ;
	assign \g72698/_0_  = _w8852_ ;
	assign \g72707/_0_  = _w8857_ ;
	assign \g72715/_0_  = _w8890_ ;
	assign \g72715/_1_  = _w8891_ ;
	assign \g72718/_0_  = _w8896_ ;
	assign \g72726/_0_  = _w8902_ ;
	assign \g72732/_0_  = _w8935_ ;
	assign \g72732/_1_  = _w8936_ ;
	assign \g72736/_0_  = _w8942_ ;
	assign \g72743/_0_  = _w8947_ ;
	assign \g72745/_0_  = _w8980_ ;
	assign \g72745/_1_  = _w8981_ ;
	assign \g72752/_0_  = _w9014_ ;
	assign \g72752/_1_  = _w9015_ ;
	assign \g72756/_0_  = _w9021_ ;
	assign \g72763/_0_  = _w9054_ ;
	assign \g72763/_1_  = _w9055_ ;
	assign \g72765/_0_  = _w9061_ ;
	assign \g72767/_0_  = _w9094_ ;
	assign \g72767/_1_  = _w9095_ ;
	assign \g72769/_0_  = _w9128_ ;
	assign \g72769/_1_  = _w9129_ ;
	assign \g72772/_0_  = _w9162_ ;
	assign \g72772/_1_  = _w9163_ ;
	assign \g72774/_0_  = _w9196_ ;
	assign \g72774/_1_  = _w9197_ ;
	assign \g72790/_0_  = _w9230_ ;
	assign \g72790/_1_  = _w9231_ ;
	assign \g72797/_0_  = _w9237_ ;
	assign \g73807/_0_  = _w9239_ ;
	assign \g73820/_0_  = _w9241_ ;
	assign \g73832/_0_  = _w9243_ ;
	assign \g73844/_0_  = _w9245_ ;
	assign \g73856/_0_  = _w9247_ ;
	assign \g73871/_0_  = _w9249_ ;
	assign \g73883/_0_  = _w9251_ ;
	assign \g73895/_0_  = _w9253_ ;
	assign \g73905/_3_  = _w2016_ ;
	assign \g73910/_0_  = _w9255_ ;
	assign \g73922/_0_  = _w9257_ ;
	assign \g73934/_0_  = _w9259_ ;
	assign \g73946/_0_  = _w9261_ ;
	assign \g73958/_0_  = _w9263_ ;
	assign \g73970/_0_  = _w9265_ ;
	assign \g73982/_0_  = _w9267_ ;
	assign \g87036/_0_  = _w9271_ ;
	assign \g87042/_0_  = _w9275_ ;
	assign \g87043/_0_  = _w9278_ ;
	assign \g87044/_0_  = _w9282_ ;
	assign \g87045/_0_  = _w9286_ ;
	assign \g87046/_0_  = _w9289_ ;
	assign \g87047/_0_  = _w9293_ ;
	assign \g87048/_0_  = _w9296_ ;
	assign \g87049/_0_  = _w9300_ ;
	assign \g87050/_0_  = _w9303_ ;
	assign \g87051/_0_  = _w9306_ ;
	assign \g87052/_0_  = _w9310_ ;
	assign \g87053/_0_  = _w9313_ ;
	assign \g87054/_0_  = _w9317_ ;
	assign \g87055/_0_  = _w9320_ ;
	assign \g87062/_0_  = _w9323_ ;
	assign \g88572/_0_  = _w9325_ ;
	assign \g88681/_0_  = _w9328_ ;
	assign \g88682/_0_  = _w9331_ ;
	assign \g88683/_0_  = _w9334_ ;
	assign \g88684/_0_  = _w9337_ ;
	assign \g88685/_0_  = _w9340_ ;
	assign \g88686/_0_  = _w9343_ ;
	assign \g88687/_0_  = _w9346_ ;
	assign \g88688/_0_  = _w9349_ ;
	assign \g88689/_0_  = _w9352_ ;
	assign \g88690/_0_  = _w9355_ ;
	assign \g88691/_0_  = _w9358_ ;
	assign \g88692/_0_  = _w9361_ ;
	assign \g88693/_0_  = _w9364_ ;
	assign \g88695/_0_  = _w9367_ ;
	assign \g88697/_0_  = _w9370_ ;
	assign \g88698/_0_  = _w9373_ ;
	assign \g88700/_0_  = _w9376_ ;
	assign \g88701/_0_  = _w9379_ ;
	assign \g88703/_0_  = _w9382_ ;
	assign \g88704/_0_  = _w9385_ ;
	assign \g88705/_0_  = _w9388_ ;
	assign \g88706/_0_  = _w9391_ ;
	assign \g88707/_0_  = _w9393_ ;
	assign \g88709/_0_  = _w9396_ ;
	assign \g88710/_0_  = _w9399_ ;
	assign \g88711/_0_  = _w9402_ ;
	assign \g88712/_0_  = _w9405_ ;
	assign \g88713/_0_  = _w9408_ ;
	assign \g88714/_0_  = _w9411_ ;
	assign \g88716/_0_  = _w9414_ ;
	assign \g88717/_0_  = _w9417_ ;
	assign \g88718/_0_  = _w9420_ ;
	assign \g88719/_0_  = _w9423_ ;
	assign \g88720/_0_  = _w9425_ ;
	assign \g88722/_0_  = _w9428_ ;
	assign \g88723/_0_  = _w9431_ ;
	assign \g88724/_0_  = _w9434_ ;
	assign \g88725/_0_  = _w9437_ ;
	assign \g88726/_0_  = _w9440_ ;
	assign \g88727/_0_  = _w9443_ ;
	assign \g88728/_0_  = _w9446_ ;
	assign \g88729/_0_  = _w9449_ ;
	assign \g88731/_0_  = _w9452_ ;
	assign \g88732/_0_  = _w9455_ ;
	assign \g88733/_0_  = _w9458_ ;
	assign \g88734/_0_  = _w9460_ ;
	assign \g88736/_0_  = _w9463_ ;
	assign \g88737/_0_  = _w9466_ ;
	assign \g88738/_0_  = _w9469_ ;
	assign \g88739/_0_  = _w9472_ ;
	assign \g88740/_0_  = _w9475_ ;
	assign \g88741/_0_  = _w9478_ ;
	assign \g88742/_0_  = _w9481_ ;
	assign \g88743/_0_  = _w9484_ ;
	assign \g88744/_0_  = _w9487_ ;
	assign \g88745/_0_  = _w9490_ ;
	assign \g88746/_0_  = _w9492_ ;
	assign \g88748/_0_  = _w9495_ ;
	assign \g88749/_0_  = _w9498_ ;
	assign \g88750/_0_  = _w9501_ ;
	assign \g88752/_0_  = _w9504_ ;
	assign \g88753/_0_  = _w9507_ ;
	assign \g88754/_0_  = _w9510_ ;
	assign \g88755/_0_  = _w9513_ ;
	assign \g88756/_0_  = _w9516_ ;
	assign \g88757/_0_  = _w9518_ ;
	assign \g88759/_0_  = _w9521_ ;
	assign \g88760/_0_  = _w9524_ ;
	assign \g88761/_0_  = _w9527_ ;
	assign \g88762/_0_  = _w9530_ ;
	assign \g88764/_0_  = _w9533_ ;
	assign \g88765/_0_  = _w9536_ ;
	assign \g88766/_0_  = _w9539_ ;
	assign \g88768/_0_  = _w9542_ ;
	assign \g88769/_0_  = _w9545_ ;
	assign \g88770/_0_  = _w9548_ ;
	assign \g88771/_0_  = _w9551_ ;
	assign \g88772/_0_  = _w9554_ ;
	assign \g88773/_0_  = _w9557_ ;
	assign \g88775/_0_  = _w9560_ ;
	assign \g88776/_0_  = _w9563_ ;
	assign \g88777/_0_  = _w9566_ ;
	assign \g88778/_0_  = _w9569_ ;
	assign \g88779/_0_  = _w9572_ ;
	assign \g88780/_0_  = _w9574_ ;
	assign \g88782/_0_  = _w9577_ ;
	assign \g88783/_0_  = _w9580_ ;
	assign \g88784/_0_  = _w9583_ ;
	assign \g88785/_0_  = _w9586_ ;
	assign \g88786/_0_  = _w9589_ ;
	assign \g88787/_0_  = _w9592_ ;
	assign \g88789/_0_  = _w9595_ ;
	assign \g88790/_0_  = _w9598_ ;
	assign \g88791/_0_  = _w9601_ ;
	assign \g88792/_0_  = _w9604_ ;
	assign \g88793/_0_  = _w9606_ ;
	assign \g88795/_0_  = _w9609_ ;
	assign \g88796/_0_  = _w9612_ ;
	assign \g88797/_0_  = _w9615_ ;
	assign \g88799/_0_  = _w9618_ ;
	assign \g88800/_0_  = _w9621_ ;
	assign \g88801/_0_  = _w9624_ ;
	assign \g88802/_0_  = _w9627_ ;
	assign \g88806/_0_  = _w9630_ ;
	assign \g88807/_0_  = _w9633_ ;
	assign \g88808/_0_  = _w9636_ ;
	assign \g88809/_0_  = _w9639_ ;
	assign \g88810/_0_  = _w9642_ ;
	assign \g88813/_0_  = _w9645_ ;
	assign \g88814/_0_  = _w9648_ ;
	assign \g88815/_0_  = _w9651_ ;
	assign \m0_ack_o_pad  = _w9682_ ;
	assign \m0_data_o[0]_pad  = _w9698_ ;
	assign \m0_data_o[10]_pad  = _w9714_ ;
	assign \m0_data_o[11]_pad  = _w9730_ ;
	assign \m0_data_o[12]_pad  = _w9746_ ;
	assign \m0_data_o[13]_pad  = _w9762_ ;
	assign \m0_data_o[14]_pad  = _w9778_ ;
	assign \m0_data_o[15]_pad  = _w9794_ ;
	assign \m0_data_o[16]_pad  = _w9807_ ;
	assign \m0_data_o[17]_pad  = _w9820_ ;
	assign \m0_data_o[18]_pad  = _w9833_ ;
	assign \m0_data_o[19]_pad  = _w9846_ ;
	assign \m0_data_o[1]_pad  = _w9862_ ;
	assign \m0_data_o[20]_pad  = _w9875_ ;
	assign \m0_data_o[21]_pad  = _w9888_ ;
	assign \m0_data_o[22]_pad  = _w9901_ ;
	assign \m0_data_o[23]_pad  = _w9914_ ;
	assign \m0_data_o[24]_pad  = _w9927_ ;
	assign \m0_data_o[25]_pad  = _w9940_ ;
	assign \m0_data_o[26]_pad  = _w9953_ ;
	assign \m0_data_o[27]_pad  = _w9966_ ;
	assign \m0_data_o[28]_pad  = _w9979_ ;
	assign \m0_data_o[29]_pad  = _w9992_ ;
	assign \m0_data_o[2]_pad  = _w10008_ ;
	assign \m0_data_o[30]_pad  = _w10021_ ;
	assign \m0_data_o[31]_pad  = _w10034_ ;
	assign \m0_data_o[3]_pad  = _w10050_ ;
	assign \m0_data_o[4]_pad  = _w10066_ ;
	assign \m0_data_o[5]_pad  = _w10082_ ;
	assign \m0_data_o[6]_pad  = _w10098_ ;
	assign \m0_data_o[7]_pad  = _w10114_ ;
	assign \m0_data_o[8]_pad  = _w10130_ ;
	assign \m0_data_o[9]_pad  = _w10146_ ;
	assign \m0_err_o_pad  = _w10174_ ;
	assign \m0_rty_o_pad  = _w10202_ ;
	assign \m1_ack_o_pad  = _w10232_ ;
	assign \m1_data_o[0]_pad  = _w10247_ ;
	assign \m1_data_o[10]_pad  = _w10262_ ;
	assign \m1_data_o[11]_pad  = _w10277_ ;
	assign \m1_data_o[12]_pad  = _w10292_ ;
	assign \m1_data_o[13]_pad  = _w10307_ ;
	assign \m1_data_o[14]_pad  = _w10322_ ;
	assign \m1_data_o[15]_pad  = _w10337_ ;
	assign \m1_data_o[16]_pad  = _w10350_ ;
	assign \m1_data_o[17]_pad  = _w10363_ ;
	assign \m1_data_o[18]_pad  = _w10376_ ;
	assign \m1_data_o[19]_pad  = _w10389_ ;
	assign \m1_data_o[1]_pad  = _w10404_ ;
	assign \m1_data_o[20]_pad  = _w10417_ ;
	assign \m1_data_o[21]_pad  = _w10430_ ;
	assign \m1_data_o[22]_pad  = _w10443_ ;
	assign \m1_data_o[23]_pad  = _w10456_ ;
	assign \m1_data_o[24]_pad  = _w10469_ ;
	assign \m1_data_o[25]_pad  = _w10482_ ;
	assign \m1_data_o[26]_pad  = _w10495_ ;
	assign \m1_data_o[27]_pad  = _w10508_ ;
	assign \m1_data_o[28]_pad  = _w10521_ ;
	assign \m1_data_o[29]_pad  = _w10534_ ;
	assign \m1_data_o[2]_pad  = _w10549_ ;
	assign \m1_data_o[30]_pad  = _w10562_ ;
	assign \m1_data_o[31]_pad  = _w10575_ ;
	assign \m1_data_o[3]_pad  = _w10590_ ;
	assign \m1_data_o[4]_pad  = _w10605_ ;
	assign \m1_data_o[5]_pad  = _w10620_ ;
	assign \m1_data_o[6]_pad  = _w10635_ ;
	assign \m1_data_o[7]_pad  = _w10650_ ;
	assign \m1_data_o[8]_pad  = _w10665_ ;
	assign \m1_data_o[9]_pad  = _w10680_ ;
	assign \m1_err_o_pad  = _w10708_ ;
	assign \m1_rty_o_pad  = _w10736_ ;
	assign \m2_ack_o_pad  = _w10766_ ;
	assign \m2_data_o[0]_pad  = _w10781_ ;
	assign \m2_data_o[10]_pad  = _w10796_ ;
	assign \m2_data_o[11]_pad  = _w10811_ ;
	assign \m2_data_o[12]_pad  = _w10826_ ;
	assign \m2_data_o[13]_pad  = _w10841_ ;
	assign \m2_data_o[14]_pad  = _w10856_ ;
	assign \m2_data_o[15]_pad  = _w10871_ ;
	assign \m2_data_o[16]_pad  = _w10884_ ;
	assign \m2_data_o[17]_pad  = _w10897_ ;
	assign \m2_data_o[18]_pad  = _w10910_ ;
	assign \m2_data_o[19]_pad  = _w10923_ ;
	assign \m2_data_o[1]_pad  = _w10938_ ;
	assign \m2_data_o[20]_pad  = _w10951_ ;
	assign \m2_data_o[21]_pad  = _w10964_ ;
	assign \m2_data_o[22]_pad  = _w10977_ ;
	assign \m2_data_o[23]_pad  = _w10990_ ;
	assign \m2_data_o[24]_pad  = _w11003_ ;
	assign \m2_data_o[25]_pad  = _w11016_ ;
	assign \m2_data_o[26]_pad  = _w11029_ ;
	assign \m2_data_o[27]_pad  = _w11042_ ;
	assign \m2_data_o[28]_pad  = _w11055_ ;
	assign \m2_data_o[29]_pad  = _w11068_ ;
	assign \m2_data_o[2]_pad  = _w11083_ ;
	assign \m2_data_o[30]_pad  = _w11096_ ;
	assign \m2_data_o[31]_pad  = _w11109_ ;
	assign \m2_data_o[3]_pad  = _w11124_ ;
	assign \m2_data_o[4]_pad  = _w11139_ ;
	assign \m2_data_o[5]_pad  = _w11154_ ;
	assign \m2_data_o[6]_pad  = _w11169_ ;
	assign \m2_data_o[7]_pad  = _w11184_ ;
	assign \m2_data_o[8]_pad  = _w11199_ ;
	assign \m2_data_o[9]_pad  = _w11214_ ;
	assign \m2_err_o_pad  = _w11242_ ;
	assign \m2_rty_o_pad  = _w11270_ ;
	assign \m3_ack_o_pad  = _w11300_ ;
	assign \m3_data_o[0]_pad  = _w11315_ ;
	assign \m3_data_o[10]_pad  = _w11330_ ;
	assign \m3_data_o[11]_pad  = _w11345_ ;
	assign \m3_data_o[12]_pad  = _w11360_ ;
	assign \m3_data_o[13]_pad  = _w11375_ ;
	assign \m3_data_o[14]_pad  = _w11390_ ;
	assign \m3_data_o[15]_pad  = _w11405_ ;
	assign \m3_data_o[16]_pad  = _w11418_ ;
	assign \m3_data_o[17]_pad  = _w11431_ ;
	assign \m3_data_o[18]_pad  = _w11444_ ;
	assign \m3_data_o[19]_pad  = _w11457_ ;
	assign \m3_data_o[1]_pad  = _w11472_ ;
	assign \m3_data_o[20]_pad  = _w11485_ ;
	assign \m3_data_o[21]_pad  = _w11498_ ;
	assign \m3_data_o[22]_pad  = _w11511_ ;
	assign \m3_data_o[23]_pad  = _w11524_ ;
	assign \m3_data_o[24]_pad  = _w11537_ ;
	assign \m3_data_o[25]_pad  = _w11550_ ;
	assign \m3_data_o[26]_pad  = _w11563_ ;
	assign \m3_data_o[27]_pad  = _w11576_ ;
	assign \m3_data_o[28]_pad  = _w11589_ ;
	assign \m3_data_o[29]_pad  = _w11602_ ;
	assign \m3_data_o[2]_pad  = _w11617_ ;
	assign \m3_data_o[30]_pad  = _w11630_ ;
	assign \m3_data_o[31]_pad  = _w11643_ ;
	assign \m3_data_o[3]_pad  = _w11658_ ;
	assign \m3_data_o[4]_pad  = _w11673_ ;
	assign \m3_data_o[5]_pad  = _w11688_ ;
	assign \m3_data_o[6]_pad  = _w11703_ ;
	assign \m3_data_o[7]_pad  = _w11718_ ;
	assign \m3_data_o[8]_pad  = _w11733_ ;
	assign \m3_data_o[9]_pad  = _w11748_ ;
	assign \m3_err_o_pad  = _w11776_ ;
	assign \m3_rty_o_pad  = _w11804_ ;
	assign \m4_ack_o_pad  = _w11834_ ;
	assign \m4_data_o[0]_pad  = _w11849_ ;
	assign \m4_data_o[10]_pad  = _w11864_ ;
	assign \m4_data_o[11]_pad  = _w11879_ ;
	assign \m4_data_o[12]_pad  = _w11894_ ;
	assign \m4_data_o[13]_pad  = _w11909_ ;
	assign \m4_data_o[14]_pad  = _w11924_ ;
	assign \m4_data_o[15]_pad  = _w11939_ ;
	assign \m4_data_o[16]_pad  = _w11952_ ;
	assign \m4_data_o[17]_pad  = _w11965_ ;
	assign \m4_data_o[18]_pad  = _w11978_ ;
	assign \m4_data_o[19]_pad  = _w11991_ ;
	assign \m4_data_o[1]_pad  = _w12006_ ;
	assign \m4_data_o[20]_pad  = _w12019_ ;
	assign \m4_data_o[21]_pad  = _w12032_ ;
	assign \m4_data_o[22]_pad  = _w12045_ ;
	assign \m4_data_o[23]_pad  = _w12058_ ;
	assign \m4_data_o[24]_pad  = _w12071_ ;
	assign \m4_data_o[25]_pad  = _w12084_ ;
	assign \m4_data_o[26]_pad  = _w12097_ ;
	assign \m4_data_o[27]_pad  = _w12110_ ;
	assign \m4_data_o[28]_pad  = _w12123_ ;
	assign \m4_data_o[29]_pad  = _w12136_ ;
	assign \m4_data_o[2]_pad  = _w12151_ ;
	assign \m4_data_o[30]_pad  = _w12164_ ;
	assign \m4_data_o[31]_pad  = _w12177_ ;
	assign \m4_data_o[3]_pad  = _w12192_ ;
	assign \m4_data_o[4]_pad  = _w12207_ ;
	assign \m4_data_o[5]_pad  = _w12222_ ;
	assign \m4_data_o[6]_pad  = _w12237_ ;
	assign \m4_data_o[7]_pad  = _w12252_ ;
	assign \m4_data_o[8]_pad  = _w12267_ ;
	assign \m4_data_o[9]_pad  = _w12282_ ;
	assign \m4_err_o_pad  = _w12310_ ;
	assign \m4_rty_o_pad  = _w12338_ ;
	assign \m5_ack_o_pad  = _w12368_ ;
	assign \m5_data_o[0]_pad  = _w12383_ ;
	assign \m5_data_o[10]_pad  = _w12398_ ;
	assign \m5_data_o[11]_pad  = _w12413_ ;
	assign \m5_data_o[12]_pad  = _w12428_ ;
	assign \m5_data_o[13]_pad  = _w12443_ ;
	assign \m5_data_o[14]_pad  = _w12458_ ;
	assign \m5_data_o[15]_pad  = _w12473_ ;
	assign \m5_data_o[16]_pad  = _w12486_ ;
	assign \m5_data_o[17]_pad  = _w12499_ ;
	assign \m5_data_o[18]_pad  = _w12512_ ;
	assign \m5_data_o[19]_pad  = _w12525_ ;
	assign \m5_data_o[1]_pad  = _w12540_ ;
	assign \m5_data_o[20]_pad  = _w12553_ ;
	assign \m5_data_o[21]_pad  = _w12566_ ;
	assign \m5_data_o[22]_pad  = _w12579_ ;
	assign \m5_data_o[23]_pad  = _w12592_ ;
	assign \m5_data_o[24]_pad  = _w12605_ ;
	assign \m5_data_o[25]_pad  = _w12618_ ;
	assign \m5_data_o[26]_pad  = _w12631_ ;
	assign \m5_data_o[27]_pad  = _w12644_ ;
	assign \m5_data_o[28]_pad  = _w12657_ ;
	assign \m5_data_o[29]_pad  = _w12670_ ;
	assign \m5_data_o[2]_pad  = _w12685_ ;
	assign \m5_data_o[30]_pad  = _w12698_ ;
	assign \m5_data_o[31]_pad  = _w12711_ ;
	assign \m5_data_o[3]_pad  = _w12726_ ;
	assign \m5_data_o[4]_pad  = _w12741_ ;
	assign \m5_data_o[5]_pad  = _w12756_ ;
	assign \m5_data_o[6]_pad  = _w12771_ ;
	assign \m5_data_o[7]_pad  = _w12786_ ;
	assign \m5_data_o[8]_pad  = _w12801_ ;
	assign \m5_data_o[9]_pad  = _w12816_ ;
	assign \m5_err_o_pad  = _w12844_ ;
	assign \m5_rty_o_pad  = _w12872_ ;
	assign \m6_ack_o_pad  = _w12902_ ;
	assign \m6_data_o[0]_pad  = _w12917_ ;
	assign \m6_data_o[10]_pad  = _w12932_ ;
	assign \m6_data_o[11]_pad  = _w12947_ ;
	assign \m6_data_o[12]_pad  = _w12962_ ;
	assign \m6_data_o[13]_pad  = _w12977_ ;
	assign \m6_data_o[14]_pad  = _w12992_ ;
	assign \m6_data_o[15]_pad  = _w13007_ ;
	assign \m6_data_o[16]_pad  = _w13020_ ;
	assign \m6_data_o[17]_pad  = _w13033_ ;
	assign \m6_data_o[18]_pad  = _w13046_ ;
	assign \m6_data_o[19]_pad  = _w13059_ ;
	assign \m6_data_o[1]_pad  = _w13074_ ;
	assign \m6_data_o[20]_pad  = _w13087_ ;
	assign \m6_data_o[21]_pad  = _w13100_ ;
	assign \m6_data_o[22]_pad  = _w13113_ ;
	assign \m6_data_o[23]_pad  = _w13126_ ;
	assign \m6_data_o[24]_pad  = _w13139_ ;
	assign \m6_data_o[25]_pad  = _w13152_ ;
	assign \m6_data_o[26]_pad  = _w13165_ ;
	assign \m6_data_o[27]_pad  = _w13178_ ;
	assign \m6_data_o[28]_pad  = _w13191_ ;
	assign \m6_data_o[29]_pad  = _w13204_ ;
	assign \m6_data_o[2]_pad  = _w13219_ ;
	assign \m6_data_o[30]_pad  = _w13232_ ;
	assign \m6_data_o[31]_pad  = _w13245_ ;
	assign \m6_data_o[3]_pad  = _w13260_ ;
	assign \m6_data_o[4]_pad  = _w13275_ ;
	assign \m6_data_o[5]_pad  = _w13290_ ;
	assign \m6_data_o[6]_pad  = _w13305_ ;
	assign \m6_data_o[7]_pad  = _w13320_ ;
	assign \m6_data_o[8]_pad  = _w13335_ ;
	assign \m6_data_o[9]_pad  = _w13350_ ;
	assign \m6_err_o_pad  = _w13378_ ;
	assign \m6_rty_o_pad  = _w13406_ ;
	assign \m7_ack_o_pad  = _w13436_ ;
	assign \m7_data_o[0]_pad  = _w13451_ ;
	assign \m7_data_o[10]_pad  = _w13466_ ;
	assign \m7_data_o[11]_pad  = _w13481_ ;
	assign \m7_data_o[12]_pad  = _w13496_ ;
	assign \m7_data_o[13]_pad  = _w13511_ ;
	assign \m7_data_o[14]_pad  = _w13526_ ;
	assign \m7_data_o[15]_pad  = _w13541_ ;
	assign \m7_data_o[16]_pad  = _w13554_ ;
	assign \m7_data_o[17]_pad  = _w13567_ ;
	assign \m7_data_o[18]_pad  = _w13580_ ;
	assign \m7_data_o[19]_pad  = _w13593_ ;
	assign \m7_data_o[1]_pad  = _w13608_ ;
	assign \m7_data_o[20]_pad  = _w13621_ ;
	assign \m7_data_o[21]_pad  = _w13634_ ;
	assign \m7_data_o[22]_pad  = _w13647_ ;
	assign \m7_data_o[23]_pad  = _w13660_ ;
	assign \m7_data_o[24]_pad  = _w13673_ ;
	assign \m7_data_o[25]_pad  = _w13686_ ;
	assign \m7_data_o[26]_pad  = _w13699_ ;
	assign \m7_data_o[27]_pad  = _w13712_ ;
	assign \m7_data_o[28]_pad  = _w13725_ ;
	assign \m7_data_o[29]_pad  = _w13738_ ;
	assign \m7_data_o[2]_pad  = _w13753_ ;
	assign \m7_data_o[30]_pad  = _w13766_ ;
	assign \m7_data_o[31]_pad  = _w13779_ ;
	assign \m7_data_o[3]_pad  = _w13794_ ;
	assign \m7_data_o[4]_pad  = _w13809_ ;
	assign \m7_data_o[5]_pad  = _w13824_ ;
	assign \m7_data_o[6]_pad  = _w13839_ ;
	assign \m7_data_o[7]_pad  = _w13854_ ;
	assign \m7_data_o[8]_pad  = _w13869_ ;
	assign \m7_data_o[9]_pad  = _w13884_ ;
	assign \m7_err_o_pad  = _w13912_ ;
	assign \m7_rty_o_pad  = _w13940_ ;
	assign \s0_addr_o[0]_pad  = _w13953_ ;
	assign \s0_addr_o[10]_pad  = _w13966_ ;
	assign \s0_addr_o[11]_pad  = _w13979_ ;
	assign \s0_addr_o[12]_pad  = _w13992_ ;
	assign \s0_addr_o[13]_pad  = _w14005_ ;
	assign \s0_addr_o[14]_pad  = _w14018_ ;
	assign \s0_addr_o[15]_pad  = _w14031_ ;
	assign \s0_addr_o[16]_pad  = _w14044_ ;
	assign \s0_addr_o[17]_pad  = _w14057_ ;
	assign \s0_addr_o[18]_pad  = _w14070_ ;
	assign \s0_addr_o[19]_pad  = _w14083_ ;
	assign \s0_addr_o[1]_pad  = _w14096_ ;
	assign \s0_addr_o[20]_pad  = _w14109_ ;
	assign \s0_addr_o[21]_pad  = _w14122_ ;
	assign \s0_addr_o[22]_pad  = _w14135_ ;
	assign \s0_addr_o[23]_pad  = _w14148_ ;
	assign \s0_addr_o[24]_pad  = _w14161_ ;
	assign \s0_addr_o[25]_pad  = _w14174_ ;
	assign \s0_addr_o[26]_pad  = _w14187_ ;
	assign \s0_addr_o[27]_pad  = _w14200_ ;
	assign \s0_addr_o[28]_pad  = _w14213_ ;
	assign \s0_addr_o[29]_pad  = _w14226_ ;
	assign \s0_addr_o[2]_pad  = _w14239_ ;
	assign \s0_addr_o[30]_pad  = _w14252_ ;
	assign \s0_addr_o[31]_pad  = _w14265_ ;
	assign \s0_addr_o[3]_pad  = _w14278_ ;
	assign \s0_addr_o[4]_pad  = _w14291_ ;
	assign \s0_addr_o[5]_pad  = _w14304_ ;
	assign \s0_addr_o[6]_pad  = _w14317_ ;
	assign \s0_addr_o[7]_pad  = _w14330_ ;
	assign \s0_addr_o[8]_pad  = _w14343_ ;
	assign \s0_addr_o[9]_pad  = _w14356_ ;
	assign \s0_data_o[0]_pad  = _w14369_ ;
	assign \s0_data_o[10]_pad  = _w14382_ ;
	assign \s0_data_o[11]_pad  = _w14395_ ;
	assign \s0_data_o[12]_pad  = _w14408_ ;
	assign \s0_data_o[13]_pad  = _w14421_ ;
	assign \s0_data_o[14]_pad  = _w14434_ ;
	assign \s0_data_o[15]_pad  = _w14447_ ;
	assign \s0_data_o[16]_pad  = _w14460_ ;
	assign \s0_data_o[17]_pad  = _w14473_ ;
	assign \s0_data_o[18]_pad  = _w14486_ ;
	assign \s0_data_o[19]_pad  = _w14499_ ;
	assign \s0_data_o[1]_pad  = _w14512_ ;
	assign \s0_data_o[20]_pad  = _w14525_ ;
	assign \s0_data_o[21]_pad  = _w14538_ ;
	assign \s0_data_o[22]_pad  = _w14551_ ;
	assign \s0_data_o[23]_pad  = _w14564_ ;
	assign \s0_data_o[24]_pad  = _w14577_ ;
	assign \s0_data_o[25]_pad  = _w14590_ ;
	assign \s0_data_o[26]_pad  = _w14603_ ;
	assign \s0_data_o[27]_pad  = _w14616_ ;
	assign \s0_data_o[28]_pad  = _w14629_ ;
	assign \s0_data_o[29]_pad  = _w14642_ ;
	assign \s0_data_o[2]_pad  = _w14655_ ;
	assign \s0_data_o[30]_pad  = _w14668_ ;
	assign \s0_data_o[31]_pad  = _w14681_ ;
	assign \s0_data_o[3]_pad  = _w14694_ ;
	assign \s0_data_o[4]_pad  = _w14707_ ;
	assign \s0_data_o[5]_pad  = _w14720_ ;
	assign \s0_data_o[6]_pad  = _w14733_ ;
	assign \s0_data_o[7]_pad  = _w14746_ ;
	assign \s0_data_o[8]_pad  = _w14759_ ;
	assign \s0_data_o[9]_pad  = _w14772_ ;
	assign \s0_sel_o[0]_pad  = _w14785_ ;
	assign \s0_sel_o[1]_pad  = _w14798_ ;
	assign \s0_sel_o[2]_pad  = _w14811_ ;
	assign \s0_sel_o[3]_pad  = _w14824_ ;
	assign \s0_stb_o_pad  = _w14837_ ;
	assign \s0_we_o_pad  = _w14850_ ;
	assign \s10_addr_o[0]_pad  = _w14863_ ;
	assign \s10_addr_o[10]_pad  = _w14876_ ;
	assign \s10_addr_o[11]_pad  = _w14889_ ;
	assign \s10_addr_o[12]_pad  = _w14902_ ;
	assign \s10_addr_o[13]_pad  = _w14915_ ;
	assign \s10_addr_o[14]_pad  = _w14928_ ;
	assign \s10_addr_o[15]_pad  = _w14941_ ;
	assign \s10_addr_o[16]_pad  = _w14954_ ;
	assign \s10_addr_o[17]_pad  = _w14967_ ;
	assign \s10_addr_o[18]_pad  = _w14980_ ;
	assign \s10_addr_o[19]_pad  = _w14993_ ;
	assign \s10_addr_o[1]_pad  = _w15006_ ;
	assign \s10_addr_o[20]_pad  = _w15019_ ;
	assign \s10_addr_o[21]_pad  = _w15032_ ;
	assign \s10_addr_o[22]_pad  = _w15045_ ;
	assign \s10_addr_o[23]_pad  = _w15058_ ;
	assign \s10_addr_o[24]_pad  = _w15071_ ;
	assign \s10_addr_o[25]_pad  = _w15084_ ;
	assign \s10_addr_o[26]_pad  = _w15097_ ;
	assign \s10_addr_o[27]_pad  = _w15110_ ;
	assign \s10_addr_o[28]_pad  = _w15123_ ;
	assign \s10_addr_o[29]_pad  = _w15136_ ;
	assign \s10_addr_o[2]_pad  = _w15149_ ;
	assign \s10_addr_o[30]_pad  = _w15162_ ;
	assign \s10_addr_o[31]_pad  = _w15175_ ;
	assign \s10_addr_o[3]_pad  = _w15188_ ;
	assign \s10_addr_o[4]_pad  = _w15201_ ;
	assign \s10_addr_o[5]_pad  = _w15214_ ;
	assign \s10_addr_o[6]_pad  = _w15227_ ;
	assign \s10_addr_o[7]_pad  = _w15240_ ;
	assign \s10_addr_o[8]_pad  = _w15253_ ;
	assign \s10_addr_o[9]_pad  = _w15266_ ;
	assign \s10_data_o[0]_pad  = _w15279_ ;
	assign \s10_data_o[10]_pad  = _w15292_ ;
	assign \s10_data_o[11]_pad  = _w15305_ ;
	assign \s10_data_o[12]_pad  = _w15318_ ;
	assign \s10_data_o[13]_pad  = _w15331_ ;
	assign \s10_data_o[14]_pad  = _w15344_ ;
	assign \s10_data_o[15]_pad  = _w15357_ ;
	assign \s10_data_o[16]_pad  = _w15370_ ;
	assign \s10_data_o[17]_pad  = _w15383_ ;
	assign \s10_data_o[18]_pad  = _w15396_ ;
	assign \s10_data_o[19]_pad  = _w15409_ ;
	assign \s10_data_o[1]_pad  = _w15422_ ;
	assign \s10_data_o[20]_pad  = _w15435_ ;
	assign \s10_data_o[21]_pad  = _w15448_ ;
	assign \s10_data_o[22]_pad  = _w15461_ ;
	assign \s10_data_o[23]_pad  = _w15474_ ;
	assign \s10_data_o[24]_pad  = _w15487_ ;
	assign \s10_data_o[25]_pad  = _w15500_ ;
	assign \s10_data_o[26]_pad  = _w15513_ ;
	assign \s10_data_o[27]_pad  = _w15526_ ;
	assign \s10_data_o[28]_pad  = _w15539_ ;
	assign \s10_data_o[29]_pad  = _w15552_ ;
	assign \s10_data_o[2]_pad  = _w15565_ ;
	assign \s10_data_o[30]_pad  = _w15578_ ;
	assign \s10_data_o[31]_pad  = _w15591_ ;
	assign \s10_data_o[3]_pad  = _w15604_ ;
	assign \s10_data_o[4]_pad  = _w15617_ ;
	assign \s10_data_o[5]_pad  = _w15630_ ;
	assign \s10_data_o[6]_pad  = _w15643_ ;
	assign \s10_data_o[7]_pad  = _w15656_ ;
	assign \s10_data_o[8]_pad  = _w15669_ ;
	assign \s10_data_o[9]_pad  = _w15682_ ;
	assign \s10_sel_o[0]_pad  = _w15695_ ;
	assign \s10_sel_o[1]_pad  = _w15708_ ;
	assign \s10_sel_o[2]_pad  = _w15721_ ;
	assign \s10_sel_o[3]_pad  = _w15734_ ;
	assign \s10_stb_o_pad  = _w15747_ ;
	assign \s10_we_o_pad  = _w15760_ ;
	assign \s11_addr_o[0]_pad  = _w15773_ ;
	assign \s11_addr_o[10]_pad  = _w15786_ ;
	assign \s11_addr_o[11]_pad  = _w15799_ ;
	assign \s11_addr_o[12]_pad  = _w15812_ ;
	assign \s11_addr_o[13]_pad  = _w15825_ ;
	assign \s11_addr_o[14]_pad  = _w15838_ ;
	assign \s11_addr_o[15]_pad  = _w15851_ ;
	assign \s11_addr_o[16]_pad  = _w15864_ ;
	assign \s11_addr_o[17]_pad  = _w15877_ ;
	assign \s11_addr_o[18]_pad  = _w15890_ ;
	assign \s11_addr_o[19]_pad  = _w15903_ ;
	assign \s11_addr_o[1]_pad  = _w15916_ ;
	assign \s11_addr_o[20]_pad  = _w15929_ ;
	assign \s11_addr_o[21]_pad  = _w15942_ ;
	assign \s11_addr_o[22]_pad  = _w15955_ ;
	assign \s11_addr_o[23]_pad  = _w15968_ ;
	assign \s11_addr_o[24]_pad  = _w15981_ ;
	assign \s11_addr_o[25]_pad  = _w15994_ ;
	assign \s11_addr_o[26]_pad  = _w16007_ ;
	assign \s11_addr_o[27]_pad  = _w16020_ ;
	assign \s11_addr_o[28]_pad  = _w16033_ ;
	assign \s11_addr_o[29]_pad  = _w16046_ ;
	assign \s11_addr_o[2]_pad  = _w16059_ ;
	assign \s11_addr_o[30]_pad  = _w16072_ ;
	assign \s11_addr_o[31]_pad  = _w16085_ ;
	assign \s11_addr_o[3]_pad  = _w16098_ ;
	assign \s11_addr_o[4]_pad  = _w16111_ ;
	assign \s11_addr_o[5]_pad  = _w16124_ ;
	assign \s11_addr_o[6]_pad  = _w16137_ ;
	assign \s11_addr_o[7]_pad  = _w16150_ ;
	assign \s11_addr_o[8]_pad  = _w16163_ ;
	assign \s11_addr_o[9]_pad  = _w16176_ ;
	assign \s11_data_o[0]_pad  = _w16189_ ;
	assign \s11_data_o[10]_pad  = _w16202_ ;
	assign \s11_data_o[11]_pad  = _w16215_ ;
	assign \s11_data_o[12]_pad  = _w16228_ ;
	assign \s11_data_o[13]_pad  = _w16241_ ;
	assign \s11_data_o[14]_pad  = _w16254_ ;
	assign \s11_data_o[15]_pad  = _w16267_ ;
	assign \s11_data_o[16]_pad  = _w16280_ ;
	assign \s11_data_o[17]_pad  = _w16293_ ;
	assign \s11_data_o[18]_pad  = _w16306_ ;
	assign \s11_data_o[19]_pad  = _w16319_ ;
	assign \s11_data_o[1]_pad  = _w16332_ ;
	assign \s11_data_o[20]_pad  = _w16345_ ;
	assign \s11_data_o[21]_pad  = _w16358_ ;
	assign \s11_data_o[22]_pad  = _w16371_ ;
	assign \s11_data_o[23]_pad  = _w16384_ ;
	assign \s11_data_o[24]_pad  = _w16397_ ;
	assign \s11_data_o[25]_pad  = _w16410_ ;
	assign \s11_data_o[26]_pad  = _w16423_ ;
	assign \s11_data_o[27]_pad  = _w16436_ ;
	assign \s11_data_o[28]_pad  = _w16449_ ;
	assign \s11_data_o[29]_pad  = _w16462_ ;
	assign \s11_data_o[2]_pad  = _w16475_ ;
	assign \s11_data_o[30]_pad  = _w16488_ ;
	assign \s11_data_o[31]_pad  = _w16501_ ;
	assign \s11_data_o[3]_pad  = _w16514_ ;
	assign \s11_data_o[4]_pad  = _w16527_ ;
	assign \s11_data_o[5]_pad  = _w16540_ ;
	assign \s11_data_o[6]_pad  = _w16553_ ;
	assign \s11_data_o[7]_pad  = _w16566_ ;
	assign \s11_data_o[8]_pad  = _w16579_ ;
	assign \s11_data_o[9]_pad  = _w16592_ ;
	assign \s11_sel_o[0]_pad  = _w16605_ ;
	assign \s11_sel_o[1]_pad  = _w16618_ ;
	assign \s11_sel_o[2]_pad  = _w16631_ ;
	assign \s11_sel_o[3]_pad  = _w16644_ ;
	assign \s11_stb_o_pad  = _w16657_ ;
	assign \s11_we_o_pad  = _w16670_ ;
	assign \s12_addr_o[0]_pad  = _w16683_ ;
	assign \s12_addr_o[10]_pad  = _w16696_ ;
	assign \s12_addr_o[11]_pad  = _w16709_ ;
	assign \s12_addr_o[12]_pad  = _w16722_ ;
	assign \s12_addr_o[13]_pad  = _w16735_ ;
	assign \s12_addr_o[14]_pad  = _w16748_ ;
	assign \s12_addr_o[15]_pad  = _w16761_ ;
	assign \s12_addr_o[16]_pad  = _w16774_ ;
	assign \s12_addr_o[17]_pad  = _w16787_ ;
	assign \s12_addr_o[18]_pad  = _w16800_ ;
	assign \s12_addr_o[19]_pad  = _w16813_ ;
	assign \s12_addr_o[1]_pad  = _w16826_ ;
	assign \s12_addr_o[20]_pad  = _w16839_ ;
	assign \s12_addr_o[21]_pad  = _w16852_ ;
	assign \s12_addr_o[22]_pad  = _w16865_ ;
	assign \s12_addr_o[23]_pad  = _w16878_ ;
	assign \s12_addr_o[24]_pad  = _w16891_ ;
	assign \s12_addr_o[25]_pad  = _w16904_ ;
	assign \s12_addr_o[26]_pad  = _w16917_ ;
	assign \s12_addr_o[27]_pad  = _w16930_ ;
	assign \s12_addr_o[28]_pad  = _w16943_ ;
	assign \s12_addr_o[29]_pad  = _w16956_ ;
	assign \s12_addr_o[2]_pad  = _w16969_ ;
	assign \s12_addr_o[30]_pad  = _w16982_ ;
	assign \s12_addr_o[31]_pad  = _w16995_ ;
	assign \s12_addr_o[3]_pad  = _w17008_ ;
	assign \s12_addr_o[4]_pad  = _w17021_ ;
	assign \s12_addr_o[5]_pad  = _w17034_ ;
	assign \s12_addr_o[6]_pad  = _w17047_ ;
	assign \s12_addr_o[7]_pad  = _w17060_ ;
	assign \s12_addr_o[8]_pad  = _w17073_ ;
	assign \s12_addr_o[9]_pad  = _w17086_ ;
	assign \s12_data_o[0]_pad  = _w17099_ ;
	assign \s12_data_o[10]_pad  = _w17112_ ;
	assign \s12_data_o[11]_pad  = _w17125_ ;
	assign \s12_data_o[12]_pad  = _w17138_ ;
	assign \s12_data_o[13]_pad  = _w17151_ ;
	assign \s12_data_o[14]_pad  = _w17164_ ;
	assign \s12_data_o[15]_pad  = _w17177_ ;
	assign \s12_data_o[16]_pad  = _w17190_ ;
	assign \s12_data_o[17]_pad  = _w17203_ ;
	assign \s12_data_o[18]_pad  = _w17216_ ;
	assign \s12_data_o[19]_pad  = _w17229_ ;
	assign \s12_data_o[1]_pad  = _w17242_ ;
	assign \s12_data_o[20]_pad  = _w17255_ ;
	assign \s12_data_o[21]_pad  = _w17268_ ;
	assign \s12_data_o[22]_pad  = _w17281_ ;
	assign \s12_data_o[23]_pad  = _w17294_ ;
	assign \s12_data_o[24]_pad  = _w17307_ ;
	assign \s12_data_o[25]_pad  = _w17320_ ;
	assign \s12_data_o[26]_pad  = _w17333_ ;
	assign \s12_data_o[27]_pad  = _w17346_ ;
	assign \s12_data_o[28]_pad  = _w17359_ ;
	assign \s12_data_o[29]_pad  = _w17372_ ;
	assign \s12_data_o[2]_pad  = _w17385_ ;
	assign \s12_data_o[30]_pad  = _w17398_ ;
	assign \s12_data_o[31]_pad  = _w17411_ ;
	assign \s12_data_o[3]_pad  = _w17424_ ;
	assign \s12_data_o[4]_pad  = _w17437_ ;
	assign \s12_data_o[5]_pad  = _w17450_ ;
	assign \s12_data_o[6]_pad  = _w17463_ ;
	assign \s12_data_o[7]_pad  = _w17476_ ;
	assign \s12_data_o[8]_pad  = _w17489_ ;
	assign \s12_data_o[9]_pad  = _w17502_ ;
	assign \s12_sel_o[0]_pad  = _w17515_ ;
	assign \s12_sel_o[1]_pad  = _w17528_ ;
	assign \s12_sel_o[2]_pad  = _w17541_ ;
	assign \s12_sel_o[3]_pad  = _w17554_ ;
	assign \s12_stb_o_pad  = _w17567_ ;
	assign \s12_we_o_pad  = _w17580_ ;
	assign \s13_addr_o[0]_pad  = _w17593_ ;
	assign \s13_addr_o[10]_pad  = _w17606_ ;
	assign \s13_addr_o[11]_pad  = _w17619_ ;
	assign \s13_addr_o[12]_pad  = _w17632_ ;
	assign \s13_addr_o[13]_pad  = _w17645_ ;
	assign \s13_addr_o[14]_pad  = _w17658_ ;
	assign \s13_addr_o[15]_pad  = _w17671_ ;
	assign \s13_addr_o[16]_pad  = _w17684_ ;
	assign \s13_addr_o[17]_pad  = _w17697_ ;
	assign \s13_addr_o[18]_pad  = _w17710_ ;
	assign \s13_addr_o[19]_pad  = _w17723_ ;
	assign \s13_addr_o[1]_pad  = _w17736_ ;
	assign \s13_addr_o[20]_pad  = _w17749_ ;
	assign \s13_addr_o[21]_pad  = _w17762_ ;
	assign \s13_addr_o[22]_pad  = _w17775_ ;
	assign \s13_addr_o[23]_pad  = _w17788_ ;
	assign \s13_addr_o[24]_pad  = _w17801_ ;
	assign \s13_addr_o[25]_pad  = _w17814_ ;
	assign \s13_addr_o[26]_pad  = _w17827_ ;
	assign \s13_addr_o[27]_pad  = _w17840_ ;
	assign \s13_addr_o[28]_pad  = _w17853_ ;
	assign \s13_addr_o[29]_pad  = _w17866_ ;
	assign \s13_addr_o[2]_pad  = _w17879_ ;
	assign \s13_addr_o[30]_pad  = _w17892_ ;
	assign \s13_addr_o[31]_pad  = _w17905_ ;
	assign \s13_addr_o[3]_pad  = _w17918_ ;
	assign \s13_addr_o[4]_pad  = _w17931_ ;
	assign \s13_addr_o[5]_pad  = _w17944_ ;
	assign \s13_addr_o[6]_pad  = _w17957_ ;
	assign \s13_addr_o[7]_pad  = _w17970_ ;
	assign \s13_addr_o[8]_pad  = _w17983_ ;
	assign \s13_addr_o[9]_pad  = _w17996_ ;
	assign \s13_data_o[0]_pad  = _w18009_ ;
	assign \s13_data_o[10]_pad  = _w18022_ ;
	assign \s13_data_o[11]_pad  = _w18035_ ;
	assign \s13_data_o[12]_pad  = _w18048_ ;
	assign \s13_data_o[13]_pad  = _w18061_ ;
	assign \s13_data_o[14]_pad  = _w18074_ ;
	assign \s13_data_o[15]_pad  = _w18087_ ;
	assign \s13_data_o[16]_pad  = _w18100_ ;
	assign \s13_data_o[17]_pad  = _w18113_ ;
	assign \s13_data_o[18]_pad  = _w18126_ ;
	assign \s13_data_o[19]_pad  = _w18139_ ;
	assign \s13_data_o[1]_pad  = _w18152_ ;
	assign \s13_data_o[20]_pad  = _w18165_ ;
	assign \s13_data_o[21]_pad  = _w18178_ ;
	assign \s13_data_o[22]_pad  = _w18191_ ;
	assign \s13_data_o[23]_pad  = _w18204_ ;
	assign \s13_data_o[24]_pad  = _w18217_ ;
	assign \s13_data_o[25]_pad  = _w18230_ ;
	assign \s13_data_o[26]_pad  = _w18243_ ;
	assign \s13_data_o[27]_pad  = _w18256_ ;
	assign \s13_data_o[28]_pad  = _w18269_ ;
	assign \s13_data_o[29]_pad  = _w18282_ ;
	assign \s13_data_o[2]_pad  = _w18295_ ;
	assign \s13_data_o[30]_pad  = _w18308_ ;
	assign \s13_data_o[31]_pad  = _w18321_ ;
	assign \s13_data_o[3]_pad  = _w18334_ ;
	assign \s13_data_o[4]_pad  = _w18347_ ;
	assign \s13_data_o[5]_pad  = _w18360_ ;
	assign \s13_data_o[6]_pad  = _w18373_ ;
	assign \s13_data_o[7]_pad  = _w18386_ ;
	assign \s13_data_o[8]_pad  = _w18399_ ;
	assign \s13_data_o[9]_pad  = _w18412_ ;
	assign \s13_sel_o[0]_pad  = _w18425_ ;
	assign \s13_sel_o[1]_pad  = _w18438_ ;
	assign \s13_sel_o[2]_pad  = _w18451_ ;
	assign \s13_sel_o[3]_pad  = _w18464_ ;
	assign \s13_stb_o_pad  = _w18477_ ;
	assign \s13_we_o_pad  = _w18490_ ;
	assign \s14_addr_o[0]_pad  = _w18503_ ;
	assign \s14_addr_o[10]_pad  = _w18516_ ;
	assign \s14_addr_o[11]_pad  = _w18529_ ;
	assign \s14_addr_o[12]_pad  = _w18542_ ;
	assign \s14_addr_o[13]_pad  = _w18555_ ;
	assign \s14_addr_o[14]_pad  = _w18568_ ;
	assign \s14_addr_o[15]_pad  = _w18581_ ;
	assign \s14_addr_o[16]_pad  = _w18594_ ;
	assign \s14_addr_o[17]_pad  = _w18607_ ;
	assign \s14_addr_o[18]_pad  = _w18620_ ;
	assign \s14_addr_o[19]_pad  = _w18633_ ;
	assign \s14_addr_o[1]_pad  = _w18646_ ;
	assign \s14_addr_o[20]_pad  = _w18659_ ;
	assign \s14_addr_o[21]_pad  = _w18672_ ;
	assign \s14_addr_o[22]_pad  = _w18685_ ;
	assign \s14_addr_o[23]_pad  = _w18698_ ;
	assign \s14_addr_o[24]_pad  = _w18711_ ;
	assign \s14_addr_o[25]_pad  = _w18724_ ;
	assign \s14_addr_o[26]_pad  = _w18737_ ;
	assign \s14_addr_o[27]_pad  = _w18750_ ;
	assign \s14_addr_o[28]_pad  = _w18763_ ;
	assign \s14_addr_o[29]_pad  = _w18776_ ;
	assign \s14_addr_o[2]_pad  = _w18789_ ;
	assign \s14_addr_o[30]_pad  = _w18802_ ;
	assign \s14_addr_o[31]_pad  = _w18815_ ;
	assign \s14_addr_o[3]_pad  = _w18828_ ;
	assign \s14_addr_o[4]_pad  = _w18841_ ;
	assign \s14_addr_o[5]_pad  = _w18854_ ;
	assign \s14_addr_o[6]_pad  = _w18867_ ;
	assign \s14_addr_o[7]_pad  = _w18880_ ;
	assign \s14_addr_o[8]_pad  = _w18893_ ;
	assign \s14_addr_o[9]_pad  = _w18906_ ;
	assign \s14_data_o[0]_pad  = _w18919_ ;
	assign \s14_data_o[10]_pad  = _w18932_ ;
	assign \s14_data_o[11]_pad  = _w18945_ ;
	assign \s14_data_o[12]_pad  = _w18958_ ;
	assign \s14_data_o[13]_pad  = _w18971_ ;
	assign \s14_data_o[14]_pad  = _w18984_ ;
	assign \s14_data_o[15]_pad  = _w18997_ ;
	assign \s14_data_o[16]_pad  = _w19010_ ;
	assign \s14_data_o[17]_pad  = _w19023_ ;
	assign \s14_data_o[18]_pad  = _w19036_ ;
	assign \s14_data_o[19]_pad  = _w19049_ ;
	assign \s14_data_o[1]_pad  = _w19062_ ;
	assign \s14_data_o[20]_pad  = _w19075_ ;
	assign \s14_data_o[21]_pad  = _w19088_ ;
	assign \s14_data_o[22]_pad  = _w19101_ ;
	assign \s14_data_o[23]_pad  = _w19114_ ;
	assign \s14_data_o[24]_pad  = _w19127_ ;
	assign \s14_data_o[25]_pad  = _w19140_ ;
	assign \s14_data_o[26]_pad  = _w19153_ ;
	assign \s14_data_o[27]_pad  = _w19166_ ;
	assign \s14_data_o[28]_pad  = _w19179_ ;
	assign \s14_data_o[29]_pad  = _w19192_ ;
	assign \s14_data_o[2]_pad  = _w19205_ ;
	assign \s14_data_o[30]_pad  = _w19218_ ;
	assign \s14_data_o[31]_pad  = _w19231_ ;
	assign \s14_data_o[3]_pad  = _w19244_ ;
	assign \s14_data_o[4]_pad  = _w19257_ ;
	assign \s14_data_o[5]_pad  = _w19270_ ;
	assign \s14_data_o[6]_pad  = _w19283_ ;
	assign \s14_data_o[7]_pad  = _w19296_ ;
	assign \s14_data_o[8]_pad  = _w19309_ ;
	assign \s14_data_o[9]_pad  = _w19322_ ;
	assign \s14_sel_o[0]_pad  = _w19335_ ;
	assign \s14_sel_o[1]_pad  = _w19348_ ;
	assign \s14_sel_o[2]_pad  = _w19361_ ;
	assign \s14_sel_o[3]_pad  = _w19374_ ;
	assign \s14_stb_o_pad  = _w19387_ ;
	assign \s14_we_o_pad  = _w19400_ ;
	assign \s15_addr_o[0]_pad  = _w19413_ ;
	assign \s15_addr_o[10]_pad  = _w19426_ ;
	assign \s15_addr_o[11]_pad  = _w19439_ ;
	assign \s15_addr_o[12]_pad  = _w19452_ ;
	assign \s15_addr_o[13]_pad  = _w19465_ ;
	assign \s15_addr_o[14]_pad  = _w19478_ ;
	assign \s15_addr_o[15]_pad  = _w19491_ ;
	assign \s15_addr_o[16]_pad  = _w19504_ ;
	assign \s15_addr_o[17]_pad  = _w19517_ ;
	assign \s15_addr_o[18]_pad  = _w19530_ ;
	assign \s15_addr_o[19]_pad  = _w19543_ ;
	assign \s15_addr_o[1]_pad  = _w19556_ ;
	assign \s15_addr_o[20]_pad  = _w19569_ ;
	assign \s15_addr_o[21]_pad  = _w19582_ ;
	assign \s15_addr_o[22]_pad  = _w19595_ ;
	assign \s15_addr_o[23]_pad  = _w19608_ ;
	assign \s15_addr_o[24]_pad  = _w2044_ ;
	assign \s15_addr_o[25]_pad  = _w2082_ ;
	assign \s15_addr_o[26]_pad  = _w2096_ ;
	assign \s15_addr_o[27]_pad  = _w2030_ ;
	assign \s15_addr_o[28]_pad  = _w19621_ ;
	assign \s15_addr_o[29]_pad  = _w19634_ ;
	assign \s15_addr_o[2]_pad  = _w1927_ ;
	assign \s15_addr_o[30]_pad  = _w19647_ ;
	assign \s15_addr_o[31]_pad  = _w19660_ ;
	assign \s15_addr_o[3]_pad  = _w1941_ ;
	assign \s15_addr_o[4]_pad  = _w1969_ ;
	assign \s15_addr_o[6]_pad  = _w19673_ ;
	assign \s15_addr_o[7]_pad  = _w19686_ ;
	assign \s15_addr_o[8]_pad  = _w19699_ ;
	assign \s15_addr_o[9]_pad  = _w19712_ ;
	assign \s15_cyc_o_pad  = _w19713_ ;
	assign \s15_data_o[0]_pad  = _w8163_ ;
	assign \s15_data_o[10]_pad  = _w8178_ ;
	assign \s15_data_o[11]_pad  = _w8193_ ;
	assign \s15_data_o[12]_pad  = _w8208_ ;
	assign \s15_data_o[13]_pad  = _w8223_ ;
	assign \s15_data_o[14]_pad  = _w8238_ ;
	assign \s15_data_o[15]_pad  = _w8253_ ;
	assign \s15_data_o[16]_pad  = _w19726_ ;
	assign \s15_data_o[17]_pad  = _w19739_ ;
	assign \s15_data_o[18]_pad  = _w19752_ ;
	assign \s15_data_o[19]_pad  = _w19765_ ;
	assign \s15_data_o[1]_pad  = _w8268_ ;
	assign \s15_data_o[20]_pad  = _w19778_ ;
	assign \s15_data_o[21]_pad  = _w19791_ ;
	assign \s15_data_o[22]_pad  = _w19804_ ;
	assign \s15_data_o[23]_pad  = _w19817_ ;
	assign \s15_data_o[24]_pad  = _w19830_ ;
	assign \s15_data_o[25]_pad  = _w19843_ ;
	assign \s15_data_o[26]_pad  = _w19856_ ;
	assign \s15_data_o[27]_pad  = _w19869_ ;
	assign \s15_data_o[28]_pad  = _w19882_ ;
	assign \s15_data_o[29]_pad  = _w19895_ ;
	assign \s15_data_o[2]_pad  = _w8283_ ;
	assign \s15_data_o[30]_pad  = _w19908_ ;
	assign \s15_data_o[31]_pad  = _w19921_ ;
	assign \s15_data_o[3]_pad  = _w8298_ ;
	assign \s15_data_o[4]_pad  = _w8313_ ;
	assign \s15_data_o[5]_pad  = _w8328_ ;
	assign \s15_data_o[6]_pad  = _w8343_ ;
	assign \s15_data_o[7]_pad  = _w8358_ ;
	assign \s15_data_o[8]_pad  = _w8373_ ;
	assign \s15_data_o[9]_pad  = _w8388_ ;
	assign \s15_sel_o[0]_pad  = _w19934_ ;
	assign \s15_sel_o[1]_pad  = _w19947_ ;
	assign \s15_sel_o[2]_pad  = _w19960_ ;
	assign \s15_sel_o[3]_pad  = _w19973_ ;
	assign \s15_stb_o_pad  = _w2068_ ;
	assign \s15_we_o_pad  = _w8645_ ;
	assign \s1_addr_o[0]_pad  = _w19986_ ;
	assign \s1_addr_o[10]_pad  = _w19999_ ;
	assign \s1_addr_o[11]_pad  = _w20012_ ;
	assign \s1_addr_o[12]_pad  = _w20025_ ;
	assign \s1_addr_o[13]_pad  = _w20038_ ;
	assign \s1_addr_o[14]_pad  = _w20051_ ;
	assign \s1_addr_o[15]_pad  = _w20064_ ;
	assign \s1_addr_o[16]_pad  = _w20077_ ;
	assign \s1_addr_o[17]_pad  = _w20090_ ;
	assign \s1_addr_o[18]_pad  = _w20103_ ;
	assign \s1_addr_o[19]_pad  = _w20116_ ;
	assign \s1_addr_o[1]_pad  = _w20129_ ;
	assign \s1_addr_o[20]_pad  = _w20142_ ;
	assign \s1_addr_o[21]_pad  = _w20155_ ;
	assign \s1_addr_o[22]_pad  = _w20168_ ;
	assign \s1_addr_o[23]_pad  = _w20181_ ;
	assign \s1_addr_o[24]_pad  = _w20194_ ;
	assign \s1_addr_o[25]_pad  = _w20207_ ;
	assign \s1_addr_o[26]_pad  = _w20220_ ;
	assign \s1_addr_o[27]_pad  = _w20233_ ;
	assign \s1_addr_o[28]_pad  = _w20246_ ;
	assign \s1_addr_o[29]_pad  = _w20259_ ;
	assign \s1_addr_o[2]_pad  = _w20272_ ;
	assign \s1_addr_o[30]_pad  = _w20285_ ;
	assign \s1_addr_o[31]_pad  = _w20298_ ;
	assign \s1_addr_o[3]_pad  = _w20311_ ;
	assign \s1_addr_o[4]_pad  = _w20324_ ;
	assign \s1_addr_o[5]_pad  = _w20337_ ;
	assign \s1_addr_o[6]_pad  = _w20350_ ;
	assign \s1_addr_o[7]_pad  = _w20363_ ;
	assign \s1_addr_o[8]_pad  = _w20376_ ;
	assign \s1_addr_o[9]_pad  = _w20389_ ;
	assign \s1_data_o[0]_pad  = _w20402_ ;
	assign \s1_data_o[10]_pad  = _w20415_ ;
	assign \s1_data_o[11]_pad  = _w20428_ ;
	assign \s1_data_o[12]_pad  = _w20441_ ;
	assign \s1_data_o[13]_pad  = _w20454_ ;
	assign \s1_data_o[14]_pad  = _w20467_ ;
	assign \s1_data_o[15]_pad  = _w20480_ ;
	assign \s1_data_o[16]_pad  = _w20493_ ;
	assign \s1_data_o[17]_pad  = _w20506_ ;
	assign \s1_data_o[18]_pad  = _w20519_ ;
	assign \s1_data_o[19]_pad  = _w20532_ ;
	assign \s1_data_o[1]_pad  = _w20545_ ;
	assign \s1_data_o[20]_pad  = _w20558_ ;
	assign \s1_data_o[21]_pad  = _w20571_ ;
	assign \s1_data_o[22]_pad  = _w20584_ ;
	assign \s1_data_o[23]_pad  = _w20597_ ;
	assign \s1_data_o[24]_pad  = _w20610_ ;
	assign \s1_data_o[25]_pad  = _w20623_ ;
	assign \s1_data_o[26]_pad  = _w20636_ ;
	assign \s1_data_o[27]_pad  = _w20649_ ;
	assign \s1_data_o[28]_pad  = _w20662_ ;
	assign \s1_data_o[29]_pad  = _w20675_ ;
	assign \s1_data_o[2]_pad  = _w20688_ ;
	assign \s1_data_o[30]_pad  = _w20701_ ;
	assign \s1_data_o[31]_pad  = _w20714_ ;
	assign \s1_data_o[3]_pad  = _w20727_ ;
	assign \s1_data_o[4]_pad  = _w20740_ ;
	assign \s1_data_o[5]_pad  = _w20753_ ;
	assign \s1_data_o[6]_pad  = _w20766_ ;
	assign \s1_data_o[7]_pad  = _w20779_ ;
	assign \s1_data_o[8]_pad  = _w20792_ ;
	assign \s1_data_o[9]_pad  = _w20805_ ;
	assign \s1_sel_o[0]_pad  = _w20818_ ;
	assign \s1_sel_o[1]_pad  = _w20831_ ;
	assign \s1_sel_o[2]_pad  = _w20844_ ;
	assign \s1_sel_o[3]_pad  = _w20857_ ;
	assign \s1_stb_o_pad  = _w20870_ ;
	assign \s1_we_o_pad  = _w20883_ ;
	assign \s2_addr_o[0]_pad  = _w20896_ ;
	assign \s2_addr_o[10]_pad  = _w20909_ ;
	assign \s2_addr_o[11]_pad  = _w20922_ ;
	assign \s2_addr_o[12]_pad  = _w20935_ ;
	assign \s2_addr_o[13]_pad  = _w20948_ ;
	assign \s2_addr_o[14]_pad  = _w20961_ ;
	assign \s2_addr_o[15]_pad  = _w20974_ ;
	assign \s2_addr_o[16]_pad  = _w20987_ ;
	assign \s2_addr_o[17]_pad  = _w21000_ ;
	assign \s2_addr_o[18]_pad  = _w21013_ ;
	assign \s2_addr_o[19]_pad  = _w21026_ ;
	assign \s2_addr_o[1]_pad  = _w21039_ ;
	assign \s2_addr_o[20]_pad  = _w21052_ ;
	assign \s2_addr_o[21]_pad  = _w21065_ ;
	assign \s2_addr_o[22]_pad  = _w21078_ ;
	assign \s2_addr_o[23]_pad  = _w21091_ ;
	assign \s2_addr_o[24]_pad  = _w21104_ ;
	assign \s2_addr_o[25]_pad  = _w21117_ ;
	assign \s2_addr_o[26]_pad  = _w21130_ ;
	assign \s2_addr_o[27]_pad  = _w21143_ ;
	assign \s2_addr_o[28]_pad  = _w21156_ ;
	assign \s2_addr_o[29]_pad  = _w21169_ ;
	assign \s2_addr_o[2]_pad  = _w21182_ ;
	assign \s2_addr_o[30]_pad  = _w21195_ ;
	assign \s2_addr_o[31]_pad  = _w21208_ ;
	assign \s2_addr_o[3]_pad  = _w21221_ ;
	assign \s2_addr_o[4]_pad  = _w21234_ ;
	assign \s2_addr_o[5]_pad  = _w21247_ ;
	assign \s2_addr_o[6]_pad  = _w21260_ ;
	assign \s2_addr_o[7]_pad  = _w21273_ ;
	assign \s2_addr_o[8]_pad  = _w21286_ ;
	assign \s2_addr_o[9]_pad  = _w21299_ ;
	assign \s2_data_o[0]_pad  = _w21312_ ;
	assign \s2_data_o[10]_pad  = _w21325_ ;
	assign \s2_data_o[11]_pad  = _w21338_ ;
	assign \s2_data_o[12]_pad  = _w21351_ ;
	assign \s2_data_o[13]_pad  = _w21364_ ;
	assign \s2_data_o[14]_pad  = _w21377_ ;
	assign \s2_data_o[15]_pad  = _w21390_ ;
	assign \s2_data_o[16]_pad  = _w21403_ ;
	assign \s2_data_o[17]_pad  = _w21416_ ;
	assign \s2_data_o[18]_pad  = _w21429_ ;
	assign \s2_data_o[19]_pad  = _w21442_ ;
	assign \s2_data_o[1]_pad  = _w21455_ ;
	assign \s2_data_o[20]_pad  = _w21468_ ;
	assign \s2_data_o[21]_pad  = _w21481_ ;
	assign \s2_data_o[22]_pad  = _w21494_ ;
	assign \s2_data_o[23]_pad  = _w21507_ ;
	assign \s2_data_o[24]_pad  = _w21520_ ;
	assign \s2_data_o[25]_pad  = _w21533_ ;
	assign \s2_data_o[26]_pad  = _w21546_ ;
	assign \s2_data_o[27]_pad  = _w21559_ ;
	assign \s2_data_o[28]_pad  = _w21572_ ;
	assign \s2_data_o[29]_pad  = _w21585_ ;
	assign \s2_data_o[2]_pad  = _w21598_ ;
	assign \s2_data_o[30]_pad  = _w21611_ ;
	assign \s2_data_o[31]_pad  = _w21624_ ;
	assign \s2_data_o[3]_pad  = _w21637_ ;
	assign \s2_data_o[4]_pad  = _w21650_ ;
	assign \s2_data_o[5]_pad  = _w21663_ ;
	assign \s2_data_o[6]_pad  = _w21676_ ;
	assign \s2_data_o[7]_pad  = _w21689_ ;
	assign \s2_data_o[8]_pad  = _w21702_ ;
	assign \s2_data_o[9]_pad  = _w21715_ ;
	assign \s2_sel_o[0]_pad  = _w21728_ ;
	assign \s2_sel_o[1]_pad  = _w21741_ ;
	assign \s2_sel_o[2]_pad  = _w21754_ ;
	assign \s2_sel_o[3]_pad  = _w21767_ ;
	assign \s2_stb_o_pad  = _w21780_ ;
	assign \s2_we_o_pad  = _w21793_ ;
	assign \s3_addr_o[0]_pad  = _w21806_ ;
	assign \s3_addr_o[10]_pad  = _w21819_ ;
	assign \s3_addr_o[11]_pad  = _w21832_ ;
	assign \s3_addr_o[12]_pad  = _w21845_ ;
	assign \s3_addr_o[13]_pad  = _w21858_ ;
	assign \s3_addr_o[14]_pad  = _w21871_ ;
	assign \s3_addr_o[15]_pad  = _w21884_ ;
	assign \s3_addr_o[16]_pad  = _w21897_ ;
	assign \s3_addr_o[17]_pad  = _w21910_ ;
	assign \s3_addr_o[18]_pad  = _w21923_ ;
	assign \s3_addr_o[19]_pad  = _w21936_ ;
	assign \s3_addr_o[1]_pad  = _w21949_ ;
	assign \s3_addr_o[20]_pad  = _w21962_ ;
	assign \s3_addr_o[21]_pad  = _w21975_ ;
	assign \s3_addr_o[22]_pad  = _w21988_ ;
	assign \s3_addr_o[23]_pad  = _w22001_ ;
	assign \s3_addr_o[24]_pad  = _w22014_ ;
	assign \s3_addr_o[25]_pad  = _w22027_ ;
	assign \s3_addr_o[26]_pad  = _w22040_ ;
	assign \s3_addr_o[27]_pad  = _w22053_ ;
	assign \s3_addr_o[28]_pad  = _w22066_ ;
	assign \s3_addr_o[29]_pad  = _w22079_ ;
	assign \s3_addr_o[2]_pad  = _w22092_ ;
	assign \s3_addr_o[30]_pad  = _w22105_ ;
	assign \s3_addr_o[31]_pad  = _w22118_ ;
	assign \s3_addr_o[3]_pad  = _w22131_ ;
	assign \s3_addr_o[4]_pad  = _w22144_ ;
	assign \s3_addr_o[5]_pad  = _w22157_ ;
	assign \s3_addr_o[6]_pad  = _w22170_ ;
	assign \s3_addr_o[7]_pad  = _w22183_ ;
	assign \s3_addr_o[8]_pad  = _w22196_ ;
	assign \s3_addr_o[9]_pad  = _w22209_ ;
	assign \s3_data_o[0]_pad  = _w22222_ ;
	assign \s3_data_o[10]_pad  = _w22235_ ;
	assign \s3_data_o[11]_pad  = _w22248_ ;
	assign \s3_data_o[12]_pad  = _w22261_ ;
	assign \s3_data_o[13]_pad  = _w22274_ ;
	assign \s3_data_o[14]_pad  = _w22287_ ;
	assign \s3_data_o[15]_pad  = _w22300_ ;
	assign \s3_data_o[16]_pad  = _w22313_ ;
	assign \s3_data_o[17]_pad  = _w22326_ ;
	assign \s3_data_o[18]_pad  = _w22339_ ;
	assign \s3_data_o[19]_pad  = _w22352_ ;
	assign \s3_data_o[1]_pad  = _w22365_ ;
	assign \s3_data_o[20]_pad  = _w22378_ ;
	assign \s3_data_o[21]_pad  = _w22391_ ;
	assign \s3_data_o[22]_pad  = _w22404_ ;
	assign \s3_data_o[23]_pad  = _w22417_ ;
	assign \s3_data_o[24]_pad  = _w22430_ ;
	assign \s3_data_o[25]_pad  = _w22443_ ;
	assign \s3_data_o[26]_pad  = _w22456_ ;
	assign \s3_data_o[27]_pad  = _w22469_ ;
	assign \s3_data_o[28]_pad  = _w22482_ ;
	assign \s3_data_o[29]_pad  = _w22495_ ;
	assign \s3_data_o[2]_pad  = _w22508_ ;
	assign \s3_data_o[30]_pad  = _w22521_ ;
	assign \s3_data_o[31]_pad  = _w22534_ ;
	assign \s3_data_o[3]_pad  = _w22547_ ;
	assign \s3_data_o[4]_pad  = _w22560_ ;
	assign \s3_data_o[5]_pad  = _w22573_ ;
	assign \s3_data_o[6]_pad  = _w22586_ ;
	assign \s3_data_o[7]_pad  = _w22599_ ;
	assign \s3_data_o[8]_pad  = _w22612_ ;
	assign \s3_data_o[9]_pad  = _w22625_ ;
	assign \s3_sel_o[0]_pad  = _w22638_ ;
	assign \s3_sel_o[1]_pad  = _w22651_ ;
	assign \s3_sel_o[2]_pad  = _w22664_ ;
	assign \s3_sel_o[3]_pad  = _w22677_ ;
	assign \s3_stb_o_pad  = _w22690_ ;
	assign \s3_we_o_pad  = _w22703_ ;
	assign \s4_addr_o[0]_pad  = _w22716_ ;
	assign \s4_addr_o[10]_pad  = _w22729_ ;
	assign \s4_addr_o[11]_pad  = _w22742_ ;
	assign \s4_addr_o[12]_pad  = _w22755_ ;
	assign \s4_addr_o[13]_pad  = _w22768_ ;
	assign \s4_addr_o[14]_pad  = _w22781_ ;
	assign \s4_addr_o[15]_pad  = _w22794_ ;
	assign \s4_addr_o[16]_pad  = _w22807_ ;
	assign \s4_addr_o[17]_pad  = _w22820_ ;
	assign \s4_addr_o[18]_pad  = _w22833_ ;
	assign \s4_addr_o[19]_pad  = _w22846_ ;
	assign \s4_addr_o[1]_pad  = _w22859_ ;
	assign \s4_addr_o[20]_pad  = _w22872_ ;
	assign \s4_addr_o[21]_pad  = _w22885_ ;
	assign \s4_addr_o[22]_pad  = _w22898_ ;
	assign \s4_addr_o[23]_pad  = _w22911_ ;
	assign \s4_addr_o[24]_pad  = _w22924_ ;
	assign \s4_addr_o[25]_pad  = _w22937_ ;
	assign \s4_addr_o[26]_pad  = _w22950_ ;
	assign \s4_addr_o[27]_pad  = _w22963_ ;
	assign \s4_addr_o[28]_pad  = _w22976_ ;
	assign \s4_addr_o[29]_pad  = _w22989_ ;
	assign \s4_addr_o[2]_pad  = _w23002_ ;
	assign \s4_addr_o[30]_pad  = _w23015_ ;
	assign \s4_addr_o[31]_pad  = _w23028_ ;
	assign \s4_addr_o[3]_pad  = _w23041_ ;
	assign \s4_addr_o[4]_pad  = _w23054_ ;
	assign \s4_addr_o[5]_pad  = _w23067_ ;
	assign \s4_addr_o[6]_pad  = _w23080_ ;
	assign \s4_addr_o[7]_pad  = _w23093_ ;
	assign \s4_addr_o[8]_pad  = _w23106_ ;
	assign \s4_addr_o[9]_pad  = _w23119_ ;
	assign \s4_data_o[0]_pad  = _w23132_ ;
	assign \s4_data_o[10]_pad  = _w23145_ ;
	assign \s4_data_o[11]_pad  = _w23158_ ;
	assign \s4_data_o[12]_pad  = _w23171_ ;
	assign \s4_data_o[13]_pad  = _w23184_ ;
	assign \s4_data_o[14]_pad  = _w23197_ ;
	assign \s4_data_o[15]_pad  = _w23210_ ;
	assign \s4_data_o[16]_pad  = _w23223_ ;
	assign \s4_data_o[17]_pad  = _w23236_ ;
	assign \s4_data_o[18]_pad  = _w23249_ ;
	assign \s4_data_o[19]_pad  = _w23262_ ;
	assign \s4_data_o[1]_pad  = _w23275_ ;
	assign \s4_data_o[20]_pad  = _w23288_ ;
	assign \s4_data_o[21]_pad  = _w23301_ ;
	assign \s4_data_o[22]_pad  = _w23314_ ;
	assign \s4_data_o[23]_pad  = _w23327_ ;
	assign \s4_data_o[24]_pad  = _w23340_ ;
	assign \s4_data_o[25]_pad  = _w23353_ ;
	assign \s4_data_o[26]_pad  = _w23366_ ;
	assign \s4_data_o[27]_pad  = _w23379_ ;
	assign \s4_data_o[28]_pad  = _w23392_ ;
	assign \s4_data_o[29]_pad  = _w23405_ ;
	assign \s4_data_o[2]_pad  = _w23418_ ;
	assign \s4_data_o[30]_pad  = _w23431_ ;
	assign \s4_data_o[31]_pad  = _w23444_ ;
	assign \s4_data_o[3]_pad  = _w23457_ ;
	assign \s4_data_o[4]_pad  = _w23470_ ;
	assign \s4_data_o[5]_pad  = _w23483_ ;
	assign \s4_data_o[6]_pad  = _w23496_ ;
	assign \s4_data_o[7]_pad  = _w23509_ ;
	assign \s4_data_o[8]_pad  = _w23522_ ;
	assign \s4_data_o[9]_pad  = _w23535_ ;
	assign \s4_sel_o[0]_pad  = _w23548_ ;
	assign \s4_sel_o[1]_pad  = _w23561_ ;
	assign \s4_sel_o[2]_pad  = _w23574_ ;
	assign \s4_sel_o[3]_pad  = _w23587_ ;
	assign \s4_stb_o_pad  = _w23600_ ;
	assign \s4_we_o_pad  = _w23613_ ;
	assign \s5_addr_o[0]_pad  = _w23626_ ;
	assign \s5_addr_o[10]_pad  = _w23639_ ;
	assign \s5_addr_o[11]_pad  = _w23652_ ;
	assign \s5_addr_o[12]_pad  = _w23665_ ;
	assign \s5_addr_o[13]_pad  = _w23678_ ;
	assign \s5_addr_o[14]_pad  = _w23691_ ;
	assign \s5_addr_o[15]_pad  = _w23704_ ;
	assign \s5_addr_o[16]_pad  = _w23717_ ;
	assign \s5_addr_o[17]_pad  = _w23730_ ;
	assign \s5_addr_o[18]_pad  = _w23743_ ;
	assign \s5_addr_o[19]_pad  = _w23756_ ;
	assign \s5_addr_o[1]_pad  = _w23769_ ;
	assign \s5_addr_o[20]_pad  = _w23782_ ;
	assign \s5_addr_o[21]_pad  = _w23795_ ;
	assign \s5_addr_o[22]_pad  = _w23808_ ;
	assign \s5_addr_o[23]_pad  = _w23821_ ;
	assign \s5_addr_o[24]_pad  = _w23834_ ;
	assign \s5_addr_o[25]_pad  = _w23847_ ;
	assign \s5_addr_o[26]_pad  = _w23860_ ;
	assign \s5_addr_o[27]_pad  = _w23873_ ;
	assign \s5_addr_o[28]_pad  = _w23886_ ;
	assign \s5_addr_o[29]_pad  = _w23899_ ;
	assign \s5_addr_o[2]_pad  = _w23912_ ;
	assign \s5_addr_o[30]_pad  = _w23925_ ;
	assign \s5_addr_o[31]_pad  = _w23938_ ;
	assign \s5_addr_o[3]_pad  = _w23951_ ;
	assign \s5_addr_o[4]_pad  = _w23964_ ;
	assign \s5_addr_o[5]_pad  = _w23977_ ;
	assign \s5_addr_o[6]_pad  = _w23990_ ;
	assign \s5_addr_o[7]_pad  = _w24003_ ;
	assign \s5_addr_o[8]_pad  = _w24016_ ;
	assign \s5_addr_o[9]_pad  = _w24029_ ;
	assign \s5_data_o[0]_pad  = _w24042_ ;
	assign \s5_data_o[10]_pad  = _w24055_ ;
	assign \s5_data_o[11]_pad  = _w24068_ ;
	assign \s5_data_o[12]_pad  = _w24081_ ;
	assign \s5_data_o[13]_pad  = _w24094_ ;
	assign \s5_data_o[14]_pad  = _w24107_ ;
	assign \s5_data_o[15]_pad  = _w24120_ ;
	assign \s5_data_o[16]_pad  = _w24133_ ;
	assign \s5_data_o[17]_pad  = _w24146_ ;
	assign \s5_data_o[18]_pad  = _w24159_ ;
	assign \s5_data_o[19]_pad  = _w24172_ ;
	assign \s5_data_o[1]_pad  = _w24185_ ;
	assign \s5_data_o[20]_pad  = _w24198_ ;
	assign \s5_data_o[21]_pad  = _w24211_ ;
	assign \s5_data_o[22]_pad  = _w24224_ ;
	assign \s5_data_o[23]_pad  = _w24237_ ;
	assign \s5_data_o[24]_pad  = _w24250_ ;
	assign \s5_data_o[25]_pad  = _w24263_ ;
	assign \s5_data_o[26]_pad  = _w24276_ ;
	assign \s5_data_o[27]_pad  = _w24289_ ;
	assign \s5_data_o[28]_pad  = _w24302_ ;
	assign \s5_data_o[29]_pad  = _w24315_ ;
	assign \s5_data_o[2]_pad  = _w24328_ ;
	assign \s5_data_o[30]_pad  = _w24341_ ;
	assign \s5_data_o[31]_pad  = _w24354_ ;
	assign \s5_data_o[3]_pad  = _w24367_ ;
	assign \s5_data_o[4]_pad  = _w24380_ ;
	assign \s5_data_o[5]_pad  = _w24393_ ;
	assign \s5_data_o[6]_pad  = _w24406_ ;
	assign \s5_data_o[7]_pad  = _w24419_ ;
	assign \s5_data_o[8]_pad  = _w24432_ ;
	assign \s5_data_o[9]_pad  = _w24445_ ;
	assign \s5_sel_o[0]_pad  = _w24458_ ;
	assign \s5_sel_o[1]_pad  = _w24471_ ;
	assign \s5_sel_o[2]_pad  = _w24484_ ;
	assign \s5_sel_o[3]_pad  = _w24497_ ;
	assign \s5_stb_o_pad  = _w24510_ ;
	assign \s5_we_o_pad  = _w24523_ ;
	assign \s6_addr_o[0]_pad  = _w24536_ ;
	assign \s6_addr_o[10]_pad  = _w24549_ ;
	assign \s6_addr_o[11]_pad  = _w24562_ ;
	assign \s6_addr_o[12]_pad  = _w24575_ ;
	assign \s6_addr_o[13]_pad  = _w24588_ ;
	assign \s6_addr_o[14]_pad  = _w24601_ ;
	assign \s6_addr_o[15]_pad  = _w24614_ ;
	assign \s6_addr_o[16]_pad  = _w24627_ ;
	assign \s6_addr_o[17]_pad  = _w24640_ ;
	assign \s6_addr_o[18]_pad  = _w24653_ ;
	assign \s6_addr_o[19]_pad  = _w24666_ ;
	assign \s6_addr_o[1]_pad  = _w24679_ ;
	assign \s6_addr_o[20]_pad  = _w24692_ ;
	assign \s6_addr_o[21]_pad  = _w24705_ ;
	assign \s6_addr_o[22]_pad  = _w24718_ ;
	assign \s6_addr_o[23]_pad  = _w24731_ ;
	assign \s6_addr_o[24]_pad  = _w24744_ ;
	assign \s6_addr_o[25]_pad  = _w24757_ ;
	assign \s6_addr_o[26]_pad  = _w24770_ ;
	assign \s6_addr_o[27]_pad  = _w24783_ ;
	assign \s6_addr_o[28]_pad  = _w24796_ ;
	assign \s6_addr_o[29]_pad  = _w24809_ ;
	assign \s6_addr_o[2]_pad  = _w24822_ ;
	assign \s6_addr_o[30]_pad  = _w24835_ ;
	assign \s6_addr_o[31]_pad  = _w24848_ ;
	assign \s6_addr_o[3]_pad  = _w24861_ ;
	assign \s6_addr_o[4]_pad  = _w24874_ ;
	assign \s6_addr_o[5]_pad  = _w24887_ ;
	assign \s6_addr_o[6]_pad  = _w24900_ ;
	assign \s6_addr_o[7]_pad  = _w24913_ ;
	assign \s6_addr_o[8]_pad  = _w24926_ ;
	assign \s6_addr_o[9]_pad  = _w24939_ ;
	assign \s6_data_o[0]_pad  = _w24952_ ;
	assign \s6_data_o[10]_pad  = _w24965_ ;
	assign \s6_data_o[11]_pad  = _w24978_ ;
	assign \s6_data_o[12]_pad  = _w24991_ ;
	assign \s6_data_o[13]_pad  = _w25004_ ;
	assign \s6_data_o[14]_pad  = _w25017_ ;
	assign \s6_data_o[15]_pad  = _w25030_ ;
	assign \s6_data_o[16]_pad  = _w25043_ ;
	assign \s6_data_o[17]_pad  = _w25056_ ;
	assign \s6_data_o[18]_pad  = _w25069_ ;
	assign \s6_data_o[19]_pad  = _w25082_ ;
	assign \s6_data_o[1]_pad  = _w25095_ ;
	assign \s6_data_o[20]_pad  = _w25108_ ;
	assign \s6_data_o[21]_pad  = _w25121_ ;
	assign \s6_data_o[22]_pad  = _w25134_ ;
	assign \s6_data_o[23]_pad  = _w25147_ ;
	assign \s6_data_o[24]_pad  = _w25160_ ;
	assign \s6_data_o[25]_pad  = _w25173_ ;
	assign \s6_data_o[26]_pad  = _w25186_ ;
	assign \s6_data_o[27]_pad  = _w25199_ ;
	assign \s6_data_o[28]_pad  = _w25212_ ;
	assign \s6_data_o[29]_pad  = _w25225_ ;
	assign \s6_data_o[2]_pad  = _w25238_ ;
	assign \s6_data_o[30]_pad  = _w25251_ ;
	assign \s6_data_o[31]_pad  = _w25264_ ;
	assign \s6_data_o[3]_pad  = _w25277_ ;
	assign \s6_data_o[4]_pad  = _w25290_ ;
	assign \s6_data_o[5]_pad  = _w25303_ ;
	assign \s6_data_o[6]_pad  = _w25316_ ;
	assign \s6_data_o[7]_pad  = _w25329_ ;
	assign \s6_data_o[8]_pad  = _w25342_ ;
	assign \s6_data_o[9]_pad  = _w25355_ ;
	assign \s6_sel_o[0]_pad  = _w25368_ ;
	assign \s6_sel_o[1]_pad  = _w25381_ ;
	assign \s6_sel_o[2]_pad  = _w25394_ ;
	assign \s6_sel_o[3]_pad  = _w25407_ ;
	assign \s6_stb_o_pad  = _w25420_ ;
	assign \s6_we_o_pad  = _w25433_ ;
	assign \s7_addr_o[0]_pad  = _w25446_ ;
	assign \s7_addr_o[10]_pad  = _w25459_ ;
	assign \s7_addr_o[11]_pad  = _w25472_ ;
	assign \s7_addr_o[12]_pad  = _w25485_ ;
	assign \s7_addr_o[13]_pad  = _w25498_ ;
	assign \s7_addr_o[14]_pad  = _w25511_ ;
	assign \s7_addr_o[15]_pad  = _w25524_ ;
	assign \s7_addr_o[16]_pad  = _w25537_ ;
	assign \s7_addr_o[17]_pad  = _w25550_ ;
	assign \s7_addr_o[18]_pad  = _w25563_ ;
	assign \s7_addr_o[19]_pad  = _w25576_ ;
	assign \s7_addr_o[1]_pad  = _w25589_ ;
	assign \s7_addr_o[20]_pad  = _w25602_ ;
	assign \s7_addr_o[21]_pad  = _w25615_ ;
	assign \s7_addr_o[22]_pad  = _w25628_ ;
	assign \s7_addr_o[23]_pad  = _w25641_ ;
	assign \s7_addr_o[24]_pad  = _w25654_ ;
	assign \s7_addr_o[25]_pad  = _w25667_ ;
	assign \s7_addr_o[26]_pad  = _w25680_ ;
	assign \s7_addr_o[27]_pad  = _w25693_ ;
	assign \s7_addr_o[28]_pad  = _w25706_ ;
	assign \s7_addr_o[29]_pad  = _w25719_ ;
	assign \s7_addr_o[2]_pad  = _w25732_ ;
	assign \s7_addr_o[30]_pad  = _w25745_ ;
	assign \s7_addr_o[31]_pad  = _w25758_ ;
	assign \s7_addr_o[3]_pad  = _w25771_ ;
	assign \s7_addr_o[4]_pad  = _w25784_ ;
	assign \s7_addr_o[5]_pad  = _w25797_ ;
	assign \s7_addr_o[6]_pad  = _w25810_ ;
	assign \s7_addr_o[7]_pad  = _w25823_ ;
	assign \s7_addr_o[8]_pad  = _w25836_ ;
	assign \s7_addr_o[9]_pad  = _w25849_ ;
	assign \s7_data_o[0]_pad  = _w25862_ ;
	assign \s7_data_o[10]_pad  = _w25875_ ;
	assign \s7_data_o[11]_pad  = _w25888_ ;
	assign \s7_data_o[12]_pad  = _w25901_ ;
	assign \s7_data_o[13]_pad  = _w25914_ ;
	assign \s7_data_o[14]_pad  = _w25927_ ;
	assign \s7_data_o[15]_pad  = _w25940_ ;
	assign \s7_data_o[16]_pad  = _w25953_ ;
	assign \s7_data_o[17]_pad  = _w25966_ ;
	assign \s7_data_o[18]_pad  = _w25979_ ;
	assign \s7_data_o[19]_pad  = _w25992_ ;
	assign \s7_data_o[1]_pad  = _w26005_ ;
	assign \s7_data_o[20]_pad  = _w26018_ ;
	assign \s7_data_o[21]_pad  = _w26031_ ;
	assign \s7_data_o[22]_pad  = _w26044_ ;
	assign \s7_data_o[23]_pad  = _w26057_ ;
	assign \s7_data_o[24]_pad  = _w26070_ ;
	assign \s7_data_o[25]_pad  = _w26083_ ;
	assign \s7_data_o[26]_pad  = _w26096_ ;
	assign \s7_data_o[27]_pad  = _w26109_ ;
	assign \s7_data_o[28]_pad  = _w26122_ ;
	assign \s7_data_o[29]_pad  = _w26135_ ;
	assign \s7_data_o[2]_pad  = _w26148_ ;
	assign \s7_data_o[30]_pad  = _w26161_ ;
	assign \s7_data_o[31]_pad  = _w26174_ ;
	assign \s7_data_o[3]_pad  = _w26187_ ;
	assign \s7_data_o[4]_pad  = _w26200_ ;
	assign \s7_data_o[5]_pad  = _w26213_ ;
	assign \s7_data_o[6]_pad  = _w26226_ ;
	assign \s7_data_o[7]_pad  = _w26239_ ;
	assign \s7_data_o[8]_pad  = _w26252_ ;
	assign \s7_data_o[9]_pad  = _w26265_ ;
	assign \s7_sel_o[0]_pad  = _w26278_ ;
	assign \s7_sel_o[1]_pad  = _w26291_ ;
	assign \s7_sel_o[2]_pad  = _w26304_ ;
	assign \s7_sel_o[3]_pad  = _w26317_ ;
	assign \s7_stb_o_pad  = _w26330_ ;
	assign \s7_we_o_pad  = _w26343_ ;
	assign \s8_addr_o[0]_pad  = _w26356_ ;
	assign \s8_addr_o[10]_pad  = _w26369_ ;
	assign \s8_addr_o[11]_pad  = _w26382_ ;
	assign \s8_addr_o[12]_pad  = _w26395_ ;
	assign \s8_addr_o[13]_pad  = _w26408_ ;
	assign \s8_addr_o[14]_pad  = _w26421_ ;
	assign \s8_addr_o[15]_pad  = _w26434_ ;
	assign \s8_addr_o[16]_pad  = _w26447_ ;
	assign \s8_addr_o[17]_pad  = _w26460_ ;
	assign \s8_addr_o[18]_pad  = _w26473_ ;
	assign \s8_addr_o[19]_pad  = _w26486_ ;
	assign \s8_addr_o[1]_pad  = _w26499_ ;
	assign \s8_addr_o[20]_pad  = _w26512_ ;
	assign \s8_addr_o[21]_pad  = _w26525_ ;
	assign \s8_addr_o[22]_pad  = _w26538_ ;
	assign \s8_addr_o[23]_pad  = _w26551_ ;
	assign \s8_addr_o[24]_pad  = _w26564_ ;
	assign \s8_addr_o[25]_pad  = _w26577_ ;
	assign \s8_addr_o[26]_pad  = _w26590_ ;
	assign \s8_addr_o[27]_pad  = _w26603_ ;
	assign \s8_addr_o[28]_pad  = _w26616_ ;
	assign \s8_addr_o[29]_pad  = _w26629_ ;
	assign \s8_addr_o[2]_pad  = _w26642_ ;
	assign \s8_addr_o[30]_pad  = _w26655_ ;
	assign \s8_addr_o[31]_pad  = _w26668_ ;
	assign \s8_addr_o[3]_pad  = _w26681_ ;
	assign \s8_addr_o[4]_pad  = _w26694_ ;
	assign \s8_addr_o[5]_pad  = _w26707_ ;
	assign \s8_addr_o[6]_pad  = _w26720_ ;
	assign \s8_addr_o[7]_pad  = _w26733_ ;
	assign \s8_addr_o[8]_pad  = _w26746_ ;
	assign \s8_addr_o[9]_pad  = _w26759_ ;
	assign \s8_data_o[0]_pad  = _w26772_ ;
	assign \s8_data_o[10]_pad  = _w26785_ ;
	assign \s8_data_o[11]_pad  = _w26798_ ;
	assign \s8_data_o[12]_pad  = _w26811_ ;
	assign \s8_data_o[13]_pad  = _w26824_ ;
	assign \s8_data_o[14]_pad  = _w26837_ ;
	assign \s8_data_o[15]_pad  = _w26850_ ;
	assign \s8_data_o[16]_pad  = _w26863_ ;
	assign \s8_data_o[17]_pad  = _w26876_ ;
	assign \s8_data_o[18]_pad  = _w26889_ ;
	assign \s8_data_o[19]_pad  = _w26902_ ;
	assign \s8_data_o[1]_pad  = _w26915_ ;
	assign \s8_data_o[20]_pad  = _w26928_ ;
	assign \s8_data_o[21]_pad  = _w26941_ ;
	assign \s8_data_o[22]_pad  = _w26954_ ;
	assign \s8_data_o[23]_pad  = _w26967_ ;
	assign \s8_data_o[24]_pad  = _w26980_ ;
	assign \s8_data_o[25]_pad  = _w26993_ ;
	assign \s8_data_o[26]_pad  = _w27006_ ;
	assign \s8_data_o[27]_pad  = _w27019_ ;
	assign \s8_data_o[28]_pad  = _w27032_ ;
	assign \s8_data_o[29]_pad  = _w27045_ ;
	assign \s8_data_o[2]_pad  = _w27058_ ;
	assign \s8_data_o[30]_pad  = _w27071_ ;
	assign \s8_data_o[31]_pad  = _w27084_ ;
	assign \s8_data_o[3]_pad  = _w27097_ ;
	assign \s8_data_o[4]_pad  = _w27110_ ;
	assign \s8_data_o[5]_pad  = _w27123_ ;
	assign \s8_data_o[6]_pad  = _w27136_ ;
	assign \s8_data_o[7]_pad  = _w27149_ ;
	assign \s8_data_o[8]_pad  = _w27162_ ;
	assign \s8_data_o[9]_pad  = _w27175_ ;
	assign \s8_sel_o[0]_pad  = _w27188_ ;
	assign \s8_sel_o[1]_pad  = _w27201_ ;
	assign \s8_sel_o[2]_pad  = _w27214_ ;
	assign \s8_sel_o[3]_pad  = _w27227_ ;
	assign \s8_stb_o_pad  = _w27240_ ;
	assign \s8_we_o_pad  = _w27253_ ;
	assign \s9_addr_o[0]_pad  = _w27266_ ;
	assign \s9_addr_o[10]_pad  = _w27279_ ;
	assign \s9_addr_o[11]_pad  = _w27292_ ;
	assign \s9_addr_o[12]_pad  = _w27305_ ;
	assign \s9_addr_o[13]_pad  = _w27318_ ;
	assign \s9_addr_o[14]_pad  = _w27331_ ;
	assign \s9_addr_o[15]_pad  = _w27344_ ;
	assign \s9_addr_o[16]_pad  = _w27357_ ;
	assign \s9_addr_o[17]_pad  = _w27370_ ;
	assign \s9_addr_o[18]_pad  = _w27383_ ;
	assign \s9_addr_o[19]_pad  = _w27396_ ;
	assign \s9_addr_o[1]_pad  = _w27409_ ;
	assign \s9_addr_o[20]_pad  = _w27422_ ;
	assign \s9_addr_o[21]_pad  = _w27435_ ;
	assign \s9_addr_o[22]_pad  = _w27448_ ;
	assign \s9_addr_o[23]_pad  = _w27461_ ;
	assign \s9_addr_o[24]_pad  = _w27474_ ;
	assign \s9_addr_o[25]_pad  = _w27487_ ;
	assign \s9_addr_o[26]_pad  = _w27500_ ;
	assign \s9_addr_o[27]_pad  = _w27513_ ;
	assign \s9_addr_o[28]_pad  = _w27526_ ;
	assign \s9_addr_o[29]_pad  = _w27539_ ;
	assign \s9_addr_o[2]_pad  = _w27552_ ;
	assign \s9_addr_o[30]_pad  = _w27565_ ;
	assign \s9_addr_o[31]_pad  = _w27578_ ;
	assign \s9_addr_o[3]_pad  = _w27591_ ;
	assign \s9_addr_o[4]_pad  = _w27604_ ;
	assign \s9_addr_o[5]_pad  = _w27617_ ;
	assign \s9_addr_o[6]_pad  = _w27630_ ;
	assign \s9_addr_o[7]_pad  = _w27643_ ;
	assign \s9_addr_o[8]_pad  = _w27656_ ;
	assign \s9_addr_o[9]_pad  = _w27669_ ;
	assign \s9_data_o[0]_pad  = _w27682_ ;
	assign \s9_data_o[10]_pad  = _w27695_ ;
	assign \s9_data_o[11]_pad  = _w27708_ ;
	assign \s9_data_o[12]_pad  = _w27721_ ;
	assign \s9_data_o[13]_pad  = _w27734_ ;
	assign \s9_data_o[14]_pad  = _w27747_ ;
	assign \s9_data_o[15]_pad  = _w27760_ ;
	assign \s9_data_o[16]_pad  = _w27773_ ;
	assign \s9_data_o[17]_pad  = _w27786_ ;
	assign \s9_data_o[18]_pad  = _w27799_ ;
	assign \s9_data_o[19]_pad  = _w27812_ ;
	assign \s9_data_o[1]_pad  = _w27825_ ;
	assign \s9_data_o[20]_pad  = _w27838_ ;
	assign \s9_data_o[21]_pad  = _w27851_ ;
	assign \s9_data_o[22]_pad  = _w27864_ ;
	assign \s9_data_o[23]_pad  = _w27877_ ;
	assign \s9_data_o[24]_pad  = _w27890_ ;
	assign \s9_data_o[25]_pad  = _w27903_ ;
	assign \s9_data_o[26]_pad  = _w27916_ ;
	assign \s9_data_o[27]_pad  = _w27929_ ;
	assign \s9_data_o[28]_pad  = _w27942_ ;
	assign \s9_data_o[29]_pad  = _w27955_ ;
	assign \s9_data_o[2]_pad  = _w27968_ ;
	assign \s9_data_o[30]_pad  = _w27981_ ;
	assign \s9_data_o[31]_pad  = _w27994_ ;
	assign \s9_data_o[3]_pad  = _w28007_ ;
	assign \s9_data_o[4]_pad  = _w28020_ ;
	assign \s9_data_o[5]_pad  = _w28033_ ;
	assign \s9_data_o[6]_pad  = _w28046_ ;
	assign \s9_data_o[7]_pad  = _w28059_ ;
	assign \s9_data_o[8]_pad  = _w28072_ ;
	assign \s9_data_o[9]_pad  = _w28085_ ;
	assign \s9_sel_o[0]_pad  = _w28098_ ;
	assign \s9_sel_o[1]_pad  = _w28111_ ;
	assign \s9_sel_o[2]_pad  = _w28124_ ;
	assign \s9_sel_o[3]_pad  = _w28137_ ;
	assign \s9_stb_o_pad  = _w28150_ ;
	assign \s9_we_o_pad  = _w28163_ ;
endmodule;