module top (\C_0_pad , \C_10_pad , \C_11_pad , \C_12_pad , \C_13_pad , \C_14_pad , \C_15_pad , \C_16_pad , \C_1_pad , \C_2_pad , \C_3_pad , \C_4_pad , \C_5_pad , \C_6_pad , \C_7_pad , \C_8_pad , \C_9_pad , \P_0_pad , \X_10_reg/NET0131 , \X_11_reg/NET0131 , \X_12_reg/NET0131 , \X_13_reg/NET0131 , \X_14_reg/NET0131 , \X_15_reg/NET0131 , \X_16_reg/P0002 , \X_1_reg/NET0131 , \X_2_reg/NET0131 , \X_3_reg/NET0131 , \X_4_reg/NET0131 , \X_5_reg/NET0131 , \X_6_reg/NET0131 , \X_7_reg/NET0131 , \X_8_reg/NET0131 , \X_9_reg/NET0131 , \X_12_reg/P0001 , \X_13_reg/P0001 , \X_14_reg/P0001 , \X_15_reg/P0001 , \X_16_reg/P0000 , \X_9_reg/P0001 , Z_pad, \_al_n0 , \_al_n1 , \g1160/_3_ , \g1169/_0_ , \g1185/_0_ , \g1212/_2_ , \g1218/_0_ , \g1234/_0_ , \g16/_1_ , \g17/_0_ , \g27/_2_ , \g29/_3_ , \g669/_1__syn_2 , \g714/_0_ , \g721/_0_ , \g734/_0_ , \g743/_0_ , \g763/_0_ );
	input \C_0_pad  ;
	input \C_10_pad  ;
	input \C_11_pad  ;
	input \C_12_pad  ;
	input \C_13_pad  ;
	input \C_14_pad  ;
	input \C_15_pad  ;
	input \C_16_pad  ;
	input \C_1_pad  ;
	input \C_2_pad  ;
	input \C_3_pad  ;
	input \C_4_pad  ;
	input \C_5_pad  ;
	input \C_6_pad  ;
	input \C_7_pad  ;
	input \C_8_pad  ;
	input \C_9_pad  ;
	input \P_0_pad  ;
	input \X_10_reg/NET0131  ;
	input \X_11_reg/NET0131  ;
	input \X_12_reg/NET0131  ;
	input \X_13_reg/NET0131  ;
	input \X_14_reg/NET0131  ;
	input \X_15_reg/NET0131  ;
	input \X_16_reg/P0002  ;
	input \X_1_reg/NET0131  ;
	input \X_2_reg/NET0131  ;
	input \X_3_reg/NET0131  ;
	input \X_4_reg/NET0131  ;
	input \X_5_reg/NET0131  ;
	input \X_6_reg/NET0131  ;
	input \X_7_reg/NET0131  ;
	input \X_8_reg/NET0131  ;
	input \X_9_reg/NET0131  ;
	output \X_12_reg/P0001  ;
	output \X_13_reg/P0001  ;
	output \X_14_reg/P0001  ;
	output \X_15_reg/P0001  ;
	output \X_16_reg/P0000  ;
	output \X_9_reg/P0001  ;
	output Z_pad ;
	output \_al_n0  ;
	output \_al_n1  ;
	output \g1160/_3_  ;
	output \g1169/_0_  ;
	output \g1185/_0_  ;
	output \g1212/_2_  ;
	output \g1218/_0_  ;
	output \g1234/_0_  ;
	output \g16/_1_  ;
	output \g17/_0_  ;
	output \g27/_2_  ;
	output \g29/_3_  ;
	output \g669/_1__syn_2  ;
	output \g714/_0_  ;
	output \g721/_0_  ;
	output \g734/_0_  ;
	output \g743/_0_  ;
	output \g763/_0_  ;
	wire _w145_ ;
	wire _w144_ ;
	wire _w143_ ;
	wire _w142_ ;
	wire _w141_ ;
	wire _w140_ ;
	wire _w139_ ;
	wire _w138_ ;
	wire _w137_ ;
	wire _w136_ ;
	wire _w135_ ;
	wire _w134_ ;
	wire _w133_ ;
	wire _w132_ ;
	wire _w131_ ;
	wire _w130_ ;
	wire _w129_ ;
	wire _w128_ ;
	wire _w127_ ;
	wire _w126_ ;
	wire _w125_ ;
	wire _w124_ ;
	wire _w123_ ;
	wire _w122_ ;
	wire _w121_ ;
	wire _w120_ ;
	wire _w119_ ;
	wire _w118_ ;
	wire _w117_ ;
	wire _w116_ ;
	wire _w115_ ;
	wire _w114_ ;
	wire _w113_ ;
	wire _w112_ ;
	wire _w111_ ;
	wire _w110_ ;
	wire _w109_ ;
	wire _w108_ ;
	wire _w107_ ;
	wire _w106_ ;
	wire _w105_ ;
	wire _w104_ ;
	wire _w103_ ;
	wire _w102_ ;
	wire _w101_ ;
	wire _w100_ ;
	wire _w99_ ;
	wire _w98_ ;
	wire _w97_ ;
	wire _w96_ ;
	wire _w95_ ;
	wire _w94_ ;
	wire _w63_ ;
	wire _w62_ ;
	wire _w61_ ;
	wire _w60_ ;
	wire _w59_ ;
	wire _w58_ ;
	wire _w57_ ;
	wire _w56_ ;
	wire _w55_ ;
	wire _w54_ ;
	wire _w53_ ;
	wire _w52_ ;
	wire _w51_ ;
	wire _w50_ ;
	wire _w49_ ;
	wire _w48_ ;
	wire _w35_ ;
	wire _w36_ ;
	wire _w37_ ;
	wire _w38_ ;
	wire _w39_ ;
	wire _w40_ ;
	wire _w41_ ;
	wire _w42_ ;
	wire _w43_ ;
	wire _w44_ ;
	wire _w45_ ;
	wire _w46_ ;
	wire _w47_ ;
	wire _w64_ ;
	wire _w65_ ;
	wire _w66_ ;
	wire _w67_ ;
	wire _w68_ ;
	wire _w69_ ;
	wire _w70_ ;
	wire _w71_ ;
	wire _w72_ ;
	wire _w73_ ;
	wire _w74_ ;
	wire _w75_ ;
	wire _w76_ ;
	wire _w77_ ;
	wire _w78_ ;
	wire _w79_ ;
	wire _w80_ ;
	wire _w81_ ;
	wire _w82_ ;
	wire _w83_ ;
	wire _w84_ ;
	wire _w85_ ;
	wire _w86_ ;
	wire _w87_ ;
	wire _w88_ ;
	wire _w89_ ;
	wire _w90_ ;
	wire _w91_ ;
	wire _w92_ ;
	wire _w93_ ;
	LUT2 #(
		.INIT('h8)
	) name0 (
		\C_13_pad ,
		\X_13_reg/NET0131 ,
		_w35_
	);
	LUT2 #(
		.INIT('h2)
	) name1 (
		\C_14_pad ,
		\X_13_reg/NET0131 ,
		_w36_
	);
	LUT2 #(
		.INIT('h8)
	) name2 (
		\X_14_reg/NET0131 ,
		_w36_,
		_w37_
	);
	LUT2 #(
		.INIT('h1)
	) name3 (
		_w35_,
		_w37_,
		_w38_
	);
	LUT2 #(
		.INIT('h2)
	) name4 (
		\P_0_pad ,
		_w38_,
		_w39_
	);
	LUT2 #(
		.INIT('h8)
	) name5 (
		\C_15_pad ,
		\X_15_reg/NET0131 ,
		_w40_
	);
	LUT2 #(
		.INIT('h2)
	) name6 (
		\C_16_pad ,
		\X_15_reg/NET0131 ,
		_w41_
	);
	LUT2 #(
		.INIT('h8)
	) name7 (
		\X_16_reg/P0002 ,
		_w41_,
		_w42_
	);
	LUT2 #(
		.INIT('h1)
	) name8 (
		_w40_,
		_w42_,
		_w43_
	);
	LUT2 #(
		.INIT('h2)
	) name9 (
		\P_0_pad ,
		\X_13_reg/NET0131 ,
		_w44_
	);
	LUT2 #(
		.INIT('h4)
	) name10 (
		\X_14_reg/NET0131 ,
		_w44_,
		_w45_
	);
	LUT2 #(
		.INIT('h4)
	) name11 (
		_w43_,
		_w45_,
		_w46_
	);
	LUT2 #(
		.INIT('h1)
	) name12 (
		_w39_,
		_w46_,
		_w47_
	);
	LUT2 #(
		.INIT('h1)
	) name13 (
		\X_10_reg/NET0131 ,
		\X_11_reg/NET0131 ,
		_w48_
	);
	LUT2 #(
		.INIT('h1)
	) name14 (
		\X_12_reg/NET0131 ,
		\X_9_reg/NET0131 ,
		_w49_
	);
	LUT2 #(
		.INIT('h8)
	) name15 (
		_w48_,
		_w49_,
		_w50_
	);
	LUT2 #(
		.INIT('h4)
	) name16 (
		_w47_,
		_w50_,
		_w51_
	);
	LUT2 #(
		.INIT('h2)
	) name17 (
		\P_0_pad ,
		\X_9_reg/NET0131 ,
		_w52_
	);
	LUT2 #(
		.INIT('h4)
	) name18 (
		\X_10_reg/NET0131 ,
		_w52_,
		_w53_
	);
	LUT2 #(
		.INIT('h8)
	) name19 (
		\C_11_pad ,
		\X_11_reg/NET0131 ,
		_w54_
	);
	LUT2 #(
		.INIT('h8)
	) name20 (
		_w53_,
		_w54_,
		_w55_
	);
	LUT2 #(
		.INIT('h8)
	) name21 (
		\C_10_pad ,
		\X_10_reg/NET0131 ,
		_w56_
	);
	LUT2 #(
		.INIT('h8)
	) name22 (
		_w52_,
		_w56_,
		_w57_
	);
	LUT2 #(
		.INIT('h1)
	) name23 (
		_w55_,
		_w57_,
		_w58_
	);
	LUT2 #(
		.INIT('h4)
	) name24 (
		_w51_,
		_w58_,
		_w59_
	);
	LUT2 #(
		.INIT('h1)
	) name25 (
		\X_1_reg/NET0131 ,
		\X_2_reg/NET0131 ,
		_w60_
	);
	LUT2 #(
		.INIT('h1)
	) name26 (
		\X_3_reg/NET0131 ,
		\X_4_reg/NET0131 ,
		_w61_
	);
	LUT2 #(
		.INIT('h8)
	) name27 (
		_w60_,
		_w61_,
		_w62_
	);
	LUT2 #(
		.INIT('h4)
	) name28 (
		\X_6_reg/NET0131 ,
		_w62_,
		_w63_
	);
	LUT2 #(
		.INIT('h1)
	) name29 (
		\X_7_reg/NET0131 ,
		\X_8_reg/NET0131 ,
		_w64_
	);
	LUT2 #(
		.INIT('h4)
	) name30 (
		\X_5_reg/NET0131 ,
		_w64_,
		_w65_
	);
	LUT2 #(
		.INIT('h8)
	) name31 (
		_w63_,
		_w65_,
		_w66_
	);
	LUT2 #(
		.INIT('h4)
	) name32 (
		_w59_,
		_w66_,
		_w67_
	);
	LUT2 #(
		.INIT('h8)
	) name33 (
		\C_5_pad ,
		\X_5_reg/NET0131 ,
		_w68_
	);
	LUT2 #(
		.INIT('h2)
	) name34 (
		\C_6_pad ,
		\X_5_reg/NET0131 ,
		_w69_
	);
	LUT2 #(
		.INIT('h8)
	) name35 (
		\X_6_reg/NET0131 ,
		_w69_,
		_w70_
	);
	LUT2 #(
		.INIT('h1)
	) name36 (
		_w68_,
		_w70_,
		_w71_
	);
	LUT2 #(
		.INIT('h2)
	) name37 (
		_w62_,
		_w71_,
		_w72_
	);
	LUT2 #(
		.INIT('h8)
	) name38 (
		\C_3_pad ,
		\X_3_reg/NET0131 ,
		_w73_
	);
	LUT2 #(
		.INIT('h2)
	) name39 (
		\C_4_pad ,
		\X_3_reg/NET0131 ,
		_w74_
	);
	LUT2 #(
		.INIT('h8)
	) name40 (
		\X_4_reg/NET0131 ,
		_w74_,
		_w75_
	);
	LUT2 #(
		.INIT('h1)
	) name41 (
		_w73_,
		_w75_,
		_w76_
	);
	LUT2 #(
		.INIT('h2)
	) name42 (
		_w60_,
		_w76_,
		_w77_
	);
	LUT2 #(
		.INIT('h8)
	) name43 (
		\C_1_pad ,
		\X_1_reg/NET0131 ,
		_w78_
	);
	LUT2 #(
		.INIT('h2)
	) name44 (
		\C_2_pad ,
		\X_1_reg/NET0131 ,
		_w79_
	);
	LUT2 #(
		.INIT('h8)
	) name45 (
		\X_2_reg/NET0131 ,
		_w79_,
		_w80_
	);
	LUT2 #(
		.INIT('h1)
	) name46 (
		\C_0_pad ,
		_w78_,
		_w81_
	);
	LUT2 #(
		.INIT('h4)
	) name47 (
		_w80_,
		_w81_,
		_w82_
	);
	LUT2 #(
		.INIT('h4)
	) name48 (
		_w72_,
		_w82_,
		_w83_
	);
	LUT2 #(
		.INIT('h4)
	) name49 (
		_w77_,
		_w83_,
		_w84_
	);
	LUT2 #(
		.INIT('h2)
	) name50 (
		\P_0_pad ,
		_w84_,
		_w85_
	);
	LUT2 #(
		.INIT('h8)
	) name51 (
		\C_9_pad ,
		\P_0_pad ,
		_w86_
	);
	LUT2 #(
		.INIT('h8)
	) name52 (
		\X_9_reg/NET0131 ,
		_w86_,
		_w87_
	);
	LUT2 #(
		.INIT('h2)
	) name53 (
		\C_12_pad ,
		\X_11_reg/NET0131 ,
		_w88_
	);
	LUT2 #(
		.INIT('h8)
	) name54 (
		\X_12_reg/NET0131 ,
		_w88_,
		_w89_
	);
	LUT2 #(
		.INIT('h8)
	) name55 (
		_w53_,
		_w89_,
		_w90_
	);
	LUT2 #(
		.INIT('h1)
	) name56 (
		_w87_,
		_w90_,
		_w91_
	);
	LUT2 #(
		.INIT('h2)
	) name57 (
		_w66_,
		_w91_,
		_w92_
	);
	LUT2 #(
		.INIT('h8)
	) name58 (
		\C_7_pad ,
		\X_7_reg/NET0131 ,
		_w93_
	);
	LUT2 #(
		.INIT('h2)
	) name59 (
		\C_8_pad ,
		\X_7_reg/NET0131 ,
		_w94_
	);
	LUT2 #(
		.INIT('h8)
	) name60 (
		\X_8_reg/NET0131 ,
		_w94_,
		_w95_
	);
	LUT2 #(
		.INIT('h1)
	) name61 (
		_w93_,
		_w95_,
		_w96_
	);
	LUT2 #(
		.INIT('h2)
	) name62 (
		\P_0_pad ,
		\X_5_reg/NET0131 ,
		_w97_
	);
	LUT2 #(
		.INIT('h8)
	) name63 (
		_w63_,
		_w97_,
		_w98_
	);
	LUT2 #(
		.INIT('h4)
	) name64 (
		_w96_,
		_w98_,
		_w99_
	);
	LUT2 #(
		.INIT('h1)
	) name65 (
		_w92_,
		_w99_,
		_w100_
	);
	LUT2 #(
		.INIT('h4)
	) name66 (
		_w85_,
		_w100_,
		_w101_
	);
	LUT2 #(
		.INIT('h4)
	) name67 (
		_w67_,
		_w101_,
		_w102_
	);
	LUT2 #(
		.INIT('h8)
	) name68 (
		\X_7_reg/NET0131 ,
		\X_8_reg/NET0131 ,
		_w103_
	);
	LUT2 #(
		.INIT('h8)
	) name69 (
		\P_0_pad ,
		\X_1_reg/NET0131 ,
		_w104_
	);
	LUT2 #(
		.INIT('h8)
	) name70 (
		\X_2_reg/NET0131 ,
		_w104_,
		_w105_
	);
	LUT2 #(
		.INIT('h8)
	) name71 (
		\X_3_reg/NET0131 ,
		_w105_,
		_w106_
	);
	LUT2 #(
		.INIT('h8)
	) name72 (
		\X_4_reg/NET0131 ,
		_w106_,
		_w107_
	);
	LUT2 #(
		.INIT('h8)
	) name73 (
		\X_5_reg/NET0131 ,
		\X_6_reg/NET0131 ,
		_w108_
	);
	LUT2 #(
		.INIT('h8)
	) name74 (
		_w107_,
		_w108_,
		_w109_
	);
	LUT2 #(
		.INIT('h8)
	) name75 (
		_w103_,
		_w109_,
		_w110_
	);
	LUT2 #(
		.INIT('h8)
	) name76 (
		\X_10_reg/NET0131 ,
		\X_4_reg/NET0131 ,
		_w111_
	);
	LUT2 #(
		.INIT('h8)
	) name77 (
		\X_9_reg/NET0131 ,
		_w111_,
		_w112_
	);
	LUT2 #(
		.INIT('h8)
	) name78 (
		_w103_,
		_w108_,
		_w113_
	);
	LUT2 #(
		.INIT('h8)
	) name79 (
		_w112_,
		_w113_,
		_w114_
	);
	LUT2 #(
		.INIT('h8)
	) name80 (
		_w106_,
		_w114_,
		_w115_
	);
	LUT2 #(
		.INIT('h8)
	) name81 (
		\X_11_reg/NET0131 ,
		_w115_,
		_w116_
	);
	LUT2 #(
		.INIT('h1)
	) name82 (
		\X_11_reg/NET0131 ,
		_w115_,
		_w117_
	);
	LUT2 #(
		.INIT('h1)
	) name83 (
		_w116_,
		_w117_,
		_w118_
	);
	LUT2 #(
		.INIT('h2)
	) name84 (
		\X_7_reg/NET0131 ,
		_w109_,
		_w119_
	);
	LUT2 #(
		.INIT('h1)
	) name85 (
		_w64_,
		_w103_,
		_w120_
	);
	LUT2 #(
		.INIT('h1)
	) name86 (
		_w119_,
		_w120_,
		_w121_
	);
	LUT2 #(
		.INIT('h8)
	) name87 (
		_w119_,
		_w120_,
		_w122_
	);
	LUT2 #(
		.INIT('h1)
	) name88 (
		_w121_,
		_w122_,
		_w123_
	);
	LUT2 #(
		.INIT('h8)
	) name89 (
		\X_12_reg/NET0131 ,
		_w116_,
		_w124_
	);
	LUT2 #(
		.INIT('h8)
	) name90 (
		\X_13_reg/NET0131 ,
		_w124_,
		_w125_
	);
	LUT2 #(
		.INIT('h1)
	) name91 (
		\X_2_reg/NET0131 ,
		_w104_,
		_w126_
	);
	LUT2 #(
		.INIT('h1)
	) name92 (
		_w105_,
		_w126_,
		_w127_
	);
	LUT2 #(
		.INIT('h8)
	) name93 (
		\X_9_reg/NET0131 ,
		_w110_,
		_w128_
	);
	LUT2 #(
		.INIT('h1)
	) name94 (
		\X_10_reg/NET0131 ,
		_w128_,
		_w129_
	);
	LUT2 #(
		.INIT('h1)
	) name95 (
		_w115_,
		_w129_,
		_w130_
	);
	LUT2 #(
		.INIT('h8)
	) name96 (
		\X_14_reg/NET0131 ,
		_w125_,
		_w131_
	);
	LUT2 #(
		.INIT('h8)
	) name97 (
		\X_5_reg/NET0131 ,
		_w107_,
		_w132_
	);
	LUT2 #(
		.INIT('h1)
	) name98 (
		\X_6_reg/NET0131 ,
		_w132_,
		_w133_
	);
	LUT2 #(
		.INIT('h1)
	) name99 (
		_w109_,
		_w133_,
		_w134_
	);
	LUT2 #(
		.INIT('h8)
	) name100 (
		\X_15_reg/NET0131 ,
		_w131_,
		_w135_
	);
	LUT2 #(
		.INIT('h1)
	) name101 (
		\X_4_reg/NET0131 ,
		_w106_,
		_w136_
	);
	LUT2 #(
		.INIT('h1)
	) name102 (
		_w107_,
		_w136_,
		_w137_
	);
	LUT2 #(
		.INIT('h4)
	) name103 (
		\X_7_reg/NET0131 ,
		_w109_,
		_w138_
	);
	LUT2 #(
		.INIT('h1)
	) name104 (
		_w119_,
		_w138_,
		_w139_
	);
	LUT2 #(
		.INIT('h1)
	) name105 (
		\X_5_reg/NET0131 ,
		_w107_,
		_w140_
	);
	LUT2 #(
		.INIT('h1)
	) name106 (
		_w132_,
		_w140_,
		_w141_
	);
	LUT2 #(
		.INIT('h1)
	) name107 (
		\X_3_reg/NET0131 ,
		_w105_,
		_w142_
	);
	LUT2 #(
		.INIT('h1)
	) name108 (
		_w106_,
		_w142_,
		_w143_
	);
	LUT2 #(
		.INIT('h1)
	) name109 (
		\P_0_pad ,
		\X_1_reg/NET0131 ,
		_w144_
	);
	LUT2 #(
		.INIT('h1)
	) name110 (
		_w104_,
		_w144_,
		_w145_
	);
	assign \X_12_reg/P0001  = \X_12_reg/NET0131 ;
	assign \X_13_reg/P0001  = \X_13_reg/NET0131 ;
	assign \X_14_reg/P0001  = \X_14_reg/NET0131 ;
	assign \X_15_reg/P0001  = \X_15_reg/NET0131 ;
	assign \X_16_reg/P0000  = \X_16_reg/P0002 ;
	assign \X_9_reg/P0001  = \X_9_reg/NET0131 ;
	assign Z_pad = _w102_ ;
	assign \_al_n0  = 1'b0;
	assign \_al_n1  = 1'b0;
	assign \g1160/_3_  = _w110_ ;
	assign \g1169/_0_  = _w118_ ;
	assign \g1185/_0_  = _w123_ ;
	assign \g1212/_2_  = _w125_ ;
	assign \g1218/_0_  = _w127_ ;
	assign \g1234/_0_  = _w130_ ;
	assign \g16/_1_  = _w131_ ;
	assign \g17/_0_  = _w134_ ;
	assign \g27/_2_  = _w124_ ;
	assign \g29/_3_  = _w116_ ;
	assign \g669/_1__syn_2  = _w135_ ;
	assign \g714/_0_  = _w137_ ;
	assign \g721/_0_  = _w139_ ;
	assign \g734/_0_  = _w141_ ;
	assign \g743/_0_  = _w143_ ;
	assign \g763/_0_  = _w145_ ;
endmodule;