module top( \B[0]  , \B[1]  , \B[2]  , \B[3]  , \B[4]  , \B[5]  , \B[6]  , \B[7]  , \B[8]  , \B[9]  , \B[10]  , \M[0]  , \M[1]  , \M[2]  , \M[3]  , \E[0]  , \E[1]  , \E[2]  );
  input \B[0]  ;
  input \B[1]  ;
  input \B[2]  ;
  input \B[3]  ;
  input \B[4]  ;
  input \B[5]  ;
  input \B[6]  ;
  input \B[7]  ;
  input \B[8]  ;
  input \B[9]  ;
  input \B[10]  ;
  output \M[0]  ;
  output \M[1]  ;
  output \M[2]  ;
  output \M[3]  ;
  output \E[0]  ;
  output \E[1]  ;
  output \E[2]  ;
  wire n12 , n13 , n14 , n15 , n16 , n17 , n18 , n19 , n20 , n21 , n22 , n23 , n24 , n25 , n26 , n27 , n28 , n29 , n30 , n31 , n32 , n33 , n34 , n35 , n36 , n37 , n38 , n39 , n40 , n41 , n42 , n43 , n44 , n45 , n46 , n47 , n48 , n49 , n50 , n51 , n52 , n53 , n54 , n55 , n56 , n57 , n58 , n59 , n60 , n61 , n62 , n63 , n64 , n65 , n66 , n67 , n68 , n69 , n70 , n71 , n72 , n73 , n74 , n75 , n76 , n77 , n78 , n79 , n80 , n81 , n82 , n83 , n84 , n85 , n86 , n87 , n88 , n89 , n90 , n91 , n92 , n93 , n94 , n95 , n96 , n97 , n98 , n99 , n100 , n101 , n102 , n103 , n104 , n105 , n106 , n107 , n108 , n109 , n110 , n111 , n112 , n113 , n114 , n115 , n116 , n117 , n118 , n119 , n120 , n121 , n122 , n123 , n124 , n125 , n126 , n127 , n128 , n129 , n130 , n131 , n132 , n133 , n134 , n135 , n136 , n137 , n138 , n139 , n140 , n141 , n142 , n143 , n144 , n145 , n146 , n147 , n148 , n149 , n150 , n151 , n152 , n153 , n154 , n155 , n156 , n157 , n158 , n159 , n160 , n161 , n162 , n163 , n164 , n165 , n166 , n167 , n168 , n169 , n170 , n171 , n172 , n173 , n174 , n175 , n176 , n177 , n178 , n179 , n180 , n181 , n182 , n183 , n184 , n185 , n186 , n187 , n188 , n189 , n190 , n191 , n192 , n193 , n194 , n195 , n196 , n197 , n198 , n199 , n200 , n201 , n202 , n203 , n204 , n205 , n206 , n207 , n208 , n209 , n210 , n211 , n212 , n213 , n214 , n215 , n216 , n217 , n218 , n219 , n220 , n221 , n222 , n223 , n224 , n225 , n226 , n227 , n228 , n229 , n230 , n231 , n232 , n233 , n234 , n235 , n236 , n237 , n238 , n239 , n240 , n241 , n242 , n243 , n244 , n245 ;
  assign n12 = ~\B[6]  & ~\B[10]  ;
  assign n13 = ~\B[6]  & ~\B[7]  ;
  assign n14 = ~n12 & ~n13 ;
  assign n15 = \B[10]  & ~n14 ;
  assign n16 = ~\B[7]  & \B[10]  ;
  assign n17 = ~\B[2]  & ~\B[3]  ;
  assign n18 = \B[2]  & \B[3]  ;
  assign n19 = ~n17 & ~n18 ;
  assign n20 = ~\B[8]  & ~\B[9]  ;
  assign n21 = ~\B[7]  & n20 ;
  assign n22 = n19 & n21 ;
  assign n23 = ~n16 & ~n22 ;
  assign n24 = ~\B[6]  & \B[7]  ;
  assign n25 = \B[10]  & n24 ;
  assign n26 = \B[8]  & \B[10]  ;
  assign n27 = \B[9]  & n26 ;
  assign n28 = ~n25 & ~n27 ;
  assign n29 = \B[10]  & n28 ;
  assign n30 = n23 & n29 ;
  assign n31 = ~n15 & ~n30 ;
  assign n32 = ~\B[3]  & \B[4]  ;
  assign n33 = \B[7]  & ~\B[8]  ;
  assign n34 = n32 & n33 ;
  assign n35 = ~\B[9]  & n34 ;
  assign n36 = ~\B[4]  & \B[7]  ;
  assign n37 = ~\B[2]  & ~\B[7]  ;
  assign n38 = \B[1]  & \B[5]  ;
  assign n39 = n37 & n38 ;
  assign n40 = ~n36 & ~n39 ;
  assign n41 = \B[3]  & ~\B[8]  ;
  assign n42 = ~\B[9]  & n41 ;
  assign n43 = ~n40 & n42 ;
  assign n44 = ~n35 & ~n43 ;
  assign n45 = ~\B[4]  & \B[8]  ;
  assign n46 = \B[1]  & \B[4]  ;
  assign n47 = ~n45 & ~n46 ;
  assign n48 = \B[0]  & ~n47 ;
  assign n49 = ~\B[0]  & ~n46 ;
  assign n50 = n13 & ~n49 ;
  assign n51 = ~n48 & n50 ;
  assign n52 = \B[4]  & \B[8]  ;
  assign n53 = ~\B[5]  & ~n52 ;
  assign n54 = ~n51 & n53 ;
  assign n55 = \B[5]  & ~n45 ;
  assign n56 = ~\B[9]  & ~n55 ;
  assign n57 = ~n54 & n56 ;
  assign n58 = n44 & ~n57 ;
  assign n59 = n23 & n28 ;
  assign n60 = n14 & ~n59 ;
  assign n61 = ~\B[5]  & \B[6]  ;
  assign n62 = \B[9]  & n61 ;
  assign n63 = \B[5]  & ~\B[6]  ;
  assign n64 = \B[1]  & ~\B[2]  ;
  assign n65 = ~n36 & n64 ;
  assign n66 = \B[3]  & \B[4]  ;
  assign n67 = ~n52 & ~n66 ;
  assign n68 = n65 & n67 ;
  assign n69 = ~\B[7]  & ~\B[8]  ;
  assign n70 = ~\B[1]  & \B[2]  ;
  assign n71 = n69 & n70 ;
  assign n72 = ~\B[9]  & ~n71 ;
  assign n73 = ~n68 & n72 ;
  assign n74 = n63 & ~n73 ;
  assign n75 = ~n62 & ~n74 ;
  assign n76 = ~n60 & n75 ;
  assign n77 = n58 & n76 ;
  assign n78 = n31 & ~n77 ;
  assign n79 = \B[7]  & ~\B[10]  ;
  assign n80 = \B[6]  & ~\B[9]  ;
  assign n81 = \B[2]  & n66 ;
  assign n82 = n80 & n81 ;
  assign n83 = ~\B[4]  & n80 ;
  assign n84 = ~\B[3]  & \B[5]  ;
  assign n85 = ~\B[6]  & n84 ;
  assign n86 = ~n83 & ~n85 ;
  assign n87 = ~\B[2]  & ~n86 ;
  assign n88 = ~n82 & ~n87 ;
  assign n89 = ~\B[1]  & n63 ;
  assign n90 = ~n83 & ~n89 ;
  assign n91 = ~\B[3]  & ~n90 ;
  assign n92 = ~\B[10]  & ~n91 ;
  assign n93 = n88 & n92 ;
  assign n94 = ~n79 & ~n93 ;
  assign n95 = \B[6]  & \B[7]  ;
  assign n96 = ~\B[8]  & ~n95 ;
  assign n97 = n94 & n96 ;
  assign n98 = ~\B[9]  & n95 ;
  assign n99 = n26 & n98 ;
  assign n100 = \B[10]  & ~n99 ;
  assign n101 = ~\B[7]  & \B[9]  ;
  assign n102 = ~\B[5]  & n101 ;
  assign n103 = \B[7]  & ~n66 ;
  assign n104 = ~\B[5]  & n20 ;
  assign n105 = n103 & n104 ;
  assign n106 = ~n102 & ~n105 ;
  assign n107 = \B[1]  & \B[2]  ;
  assign n108 = \B[0]  & ~n107 ;
  assign n109 = \B[4]  & ~\B[7]  ;
  assign n110 = ~\B[0]  & \B[2]  ;
  assign n111 = n109 & ~n110 ;
  assign n112 = ~n108 & n111 ;
  assign n113 = \B[8]  & ~\B[9]  ;
  assign n114 = ~\B[4]  & ~\B[9]  ;
  assign n115 = ~n37 & ~n114 ;
  assign n116 = ~\B[1]  & ~n115 ;
  assign n117 = ~n113 & ~n116 ;
  assign n118 = ~n112 & n117 ;
  assign n119 = ~\B[5]  & ~\B[6]  ;
  assign n120 = ~n118 & n119 ;
  assign n121 = n106 & ~n120 ;
  assign n122 = ~\B[4]  & ~\B[6]  ;
  assign n123 = n113 & n122 ;
  assign n124 = \B[9]  & n13 ;
  assign n125 = ~n123 & ~n124 ;
  assign n126 = ~\B[5]  & n125 ;
  assign n127 = ~\B[4]  & ~n13 ;
  assign n128 = \B[3]  & ~n127 ;
  assign n129 = \B[4]  & ~n20 ;
  assign n130 = ~\B[7]  & ~n107 ;
  assign n131 = ~n129 & ~n130 ;
  assign n132 = n128 & n131 ;
  assign n133 = \B[6]  & ~n20 ;
  assign n134 = ~n101 & ~n114 ;
  assign n135 = n133 & n134 ;
  assign n136 = n125 & ~n135 ;
  assign n137 = ~n132 & n136 ;
  assign n138 = ~n126 & ~n137 ;
  assign n139 = ~n99 & ~n138 ;
  assign n140 = n121 & n139 ;
  assign n141 = ~n100 & ~n140 ;
  assign n142 = ~n97 & ~n141 ;
  assign n143 = \B[4]  & \B[5]  ;
  assign n144 = ~n95 & ~n143 ;
  assign n145 = \B[8]  & n144 ;
  assign n146 = \B[3]  & ~\B[6]  ;
  assign n147 = ~n37 & ~n146 ;
  assign n148 = ~n13 & ~n147 ;
  assign n149 = \B[8]  & n143 ;
  assign n150 = ~n148 & n149 ;
  assign n151 = ~n145 & ~n150 ;
  assign n152 = ~\B[9]  & ~\B[10]  ;
  assign n153 = n151 & n152 ;
  assign n154 = \B[5]  & \B[6]  ;
  assign n155 = n109 & n154 ;
  assign n156 = ~n24 & ~n155 ;
  assign n157 = \B[8]  & ~\B[10]  ;
  assign n158 = ~n156 & n157 ;
  assign n159 = ~n153 & ~n158 ;
  assign n160 = \B[4]  & n84 ;
  assign n161 = ~\B[2]  & ~\B[6]  ;
  assign n162 = n66 & n161 ;
  assign n163 = ~n160 & ~n162 ;
  assign n164 = ~\B[7]  & ~n163 ;
  assign n165 = \B[0]  & ~\B[6]  ;
  assign n166 = n32 & n165 ;
  assign n167 = \B[3]  & ~\B[4]  ;
  assign n168 = \B[5]  & n167 ;
  assign n169 = ~n166 & ~n168 ;
  assign n170 = \B[1]  & ~n169 ;
  assign n171 = \B[0]  & \B[1]  ;
  assign n172 = n66 & ~n171 ;
  assign n173 = ~n122 & ~n172 ;
  assign n174 = ~\B[5]  & ~n173 ;
  assign n175 = ~n170 & ~n174 ;
  assign n176 = \B[2]  & ~\B[7]  ;
  assign n177 = ~n175 & n176 ;
  assign n178 = ~n164 & ~n177 ;
  assign n179 = n143 & ~n148 ;
  assign n180 = ~n144 & ~n179 ;
  assign n181 = ~n66 & n154 ;
  assign n182 = \B[2]  & n61 ;
  assign n183 = ~n89 & ~n182 ;
  assign n184 = n66 & ~n183 ;
  assign n185 = ~n181 & ~n184 ;
  assign n186 = ~n180 & n185 ;
  assign n187 = ~n158 & n186 ;
  assign n188 = n178 & n187 ;
  assign n189 = ~n159 & ~n188 ;
  assign n190 = \B[9]  & \B[10]  ;
  assign n191 = \B[5]  & \B[7]  ;
  assign n192 = \B[8]  & \B[9]  ;
  assign n193 = ~n191 & n192 ;
  assign n194 = ~n190 & ~n193 ;
  assign n195 = \B[5]  & ~\B[8]  ;
  assign n196 = \B[9]  & n195 ;
  assign n197 = ~n26 & ~n196 ;
  assign n198 = n95 & ~n197 ;
  assign n199 = n194 & ~n198 ;
  assign n200 = ~n189 & n199 ;
  assign n201 = ~\B[5]  & n69 ;
  assign n202 = n122 & n201 ;
  assign n203 = ~\B[2]  & \B[7]  ;
  assign n204 = n154 & n203 ;
  assign n205 = n52 & n204 ;
  assign n206 = ~n202 & ~n205 ;
  assign n207 = ~\B[3]  & n152 ;
  assign n208 = ~n206 & n207 ;
  assign n209 = \B[5]  & \B[8]  ;
  assign n210 = n95 & n209 ;
  assign n211 = \B[9]  & ~n210 ;
  assign n212 = ~\B[10]  & n211 ;
  assign n213 = ~n17 & n143 ;
  assign n214 = ~n41 & n213 ;
  assign n215 = ~\B[10]  & n98 ;
  assign n216 = n214 & n215 ;
  assign n217 = ~n212 & ~n216 ;
  assign n218 = ~\B[8]  & ~\B[10]  ;
  assign n219 = \B[4]  & ~n84 ;
  assign n220 = ~\B[6]  & ~n219 ;
  assign n221 = n119 & n171 ;
  assign n222 = ~n155 & ~n221 ;
  assign n223 = n18 & ~n222 ;
  assign n224 = \B[5]  & ~n107 ;
  assign n225 = ~\B[7]  & ~n224 ;
  assign n226 = ~n103 & n154 ;
  assign n227 = ~n225 & ~n226 ;
  assign n228 = ~n223 & ~n227 ;
  assign n229 = ~n220 & n228 ;
  assign n230 = n218 & ~n229 ;
  assign n231 = n217 & ~n230 ;
  assign n232 = ~n17 & n210 ;
  assign n233 = n18 & n171 ;
  assign n234 = n201 & n233 ;
  assign n235 = ~n232 & ~n234 ;
  assign n236 = \B[4]  & ~n235 ;
  assign n237 = n69 & ~n119 ;
  assign n238 = n152 & ~n237 ;
  assign n239 = n152 & n154 ;
  assign n240 = n81 & n239 ;
  assign n241 = ~n238 & ~n240 ;
  assign n242 = ~n236 & ~n241 ;
  assign n243 = n81 & n154 ;
  assign n244 = n69 & n152 ;
  assign n245 = ~n243 & n244 ;
  assign \M[0]  = n78 ;
  assign \M[1]  = n142 ;
  assign \M[2]  = ~n200 ;
  assign \M[3]  = ~n208 ;
  assign \E[0]  = n231 ;
  assign \E[1]  = ~n242 ;
  assign \E[2]  = ~n245 ;
endmodule
