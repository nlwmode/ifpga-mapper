module top (\103GAT(6)_pad , \120GAT(7)_pad , \137GAT(8)_pad , \154GAT(9)_pad , \171GAT(10)_pad , \188GAT(11)_pad , \18GAT(1)_pad , \1GAT(0)_pad , \205GAT(12)_pad , \222GAT(13)_pad , \239GAT(14)_pad , \256GAT(15)_pad , \273GAT(16)_pad , \290GAT(17)_pad , \307GAT(18)_pad , \324GAT(19)_pad , \341GAT(20)_pad , \358GAT(21)_pad , \35GAT(2)_pad , \375GAT(22)_pad , \392GAT(23)_pad , \409GAT(24)_pad , \426GAT(25)_pad , \443GAT(26)_pad , \460GAT(27)_pad , \477GAT(28)_pad , \494GAT(29)_pad , \511GAT(30)_pad , \528GAT(31)_pad , \52GAT(3)_pad , \69GAT(4)_pad , \86GAT(5)_pad , \1581GAT(423)_pad , \1901GAT(561)_pad , \2223GAT(700)_pad , \2548GAT(840)_pad , \2877GAT(983)_pad , \3211GAT(1128)_pad , \3552GAT(1275)_pad , \3895GAT(1423)_pad , \4241GAT(1572)_pad , \4591GAT(1722)_pad , \4946GAT(1876)_pad , \5308GAT(2031)_pad , \545GAT(287)_pad , \5672GAT(2187)_pad , \5971GAT(2309)_pad , \6123GAT(2368)_pad , \6150GAT(2378)_pad , \6160GAT(2383)_pad , \6170GAT(2388)_pad , \6180GAT(2393)_pad , \6190GAT(2398)_pad , \6200GAT(2403)_pad , \6210GAT(2408)_pad , \6220GAT(2413)_pad , \6230GAT(2418)_pad , \6240GAT(2423)_pad , \6250GAT(2428)_pad , \6260GAT(2433)_pad , \6270GAT(2438)_pad , \6280GAT(2443)_pad , \6287GAT(2444)_pad , \6288GAT(2447)_pad );
	input \103GAT(6)_pad  ;
	input \120GAT(7)_pad  ;
	input \137GAT(8)_pad  ;
	input \154GAT(9)_pad  ;
	input \171GAT(10)_pad  ;
	input \188GAT(11)_pad  ;
	input \18GAT(1)_pad  ;
	input \1GAT(0)_pad  ;
	input \205GAT(12)_pad  ;
	input \222GAT(13)_pad  ;
	input \239GAT(14)_pad  ;
	input \256GAT(15)_pad  ;
	input \273GAT(16)_pad  ;
	input \290GAT(17)_pad  ;
	input \307GAT(18)_pad  ;
	input \324GAT(19)_pad  ;
	input \341GAT(20)_pad  ;
	input \358GAT(21)_pad  ;
	input \35GAT(2)_pad  ;
	input \375GAT(22)_pad  ;
	input \392GAT(23)_pad  ;
	input \409GAT(24)_pad  ;
	input \426GAT(25)_pad  ;
	input \443GAT(26)_pad  ;
	input \460GAT(27)_pad  ;
	input \477GAT(28)_pad  ;
	input \494GAT(29)_pad  ;
	input \511GAT(30)_pad  ;
	input \528GAT(31)_pad  ;
	input \52GAT(3)_pad  ;
	input \69GAT(4)_pad  ;
	input \86GAT(5)_pad  ;
	output \1581GAT(423)_pad  ;
	output \1901GAT(561)_pad  ;
	output \2223GAT(700)_pad  ;
	output \2548GAT(840)_pad  ;
	output \2877GAT(983)_pad  ;
	output \3211GAT(1128)_pad  ;
	output \3552GAT(1275)_pad  ;
	output \3895GAT(1423)_pad  ;
	output \4241GAT(1572)_pad  ;
	output \4591GAT(1722)_pad  ;
	output \4946GAT(1876)_pad  ;
	output \5308GAT(2031)_pad  ;
	output \545GAT(287)_pad  ;
	output \5672GAT(2187)_pad  ;
	output \5971GAT(2309)_pad  ;
	output \6123GAT(2368)_pad  ;
	output \6150GAT(2378)_pad  ;
	output \6160GAT(2383)_pad  ;
	output \6170GAT(2388)_pad  ;
	output \6180GAT(2393)_pad  ;
	output \6190GAT(2398)_pad  ;
	output \6200GAT(2403)_pad  ;
	output \6210GAT(2408)_pad  ;
	output \6220GAT(2413)_pad  ;
	output \6230GAT(2418)_pad  ;
	output \6240GAT(2423)_pad  ;
	output \6250GAT(2428)_pad  ;
	output \6260GAT(2433)_pad  ;
	output \6270GAT(2438)_pad  ;
	output \6280GAT(2443)_pad  ;
	output \6287GAT(2444)_pad  ;
	output \6288GAT(2447)_pad  ;
	wire _w1902_ ;
	wire _w1901_ ;
	wire _w1900_ ;
	wire _w1899_ ;
	wire _w1898_ ;
	wire _w1897_ ;
	wire _w1896_ ;
	wire _w1895_ ;
	wire _w1894_ ;
	wire _w1893_ ;
	wire _w1892_ ;
	wire _w1891_ ;
	wire _w1890_ ;
	wire _w1889_ ;
	wire _w1888_ ;
	wire _w1887_ ;
	wire _w1886_ ;
	wire _w1885_ ;
	wire _w1884_ ;
	wire _w1883_ ;
	wire _w1882_ ;
	wire _w1881_ ;
	wire _w1880_ ;
	wire _w1879_ ;
	wire _w1878_ ;
	wire _w1877_ ;
	wire _w1876_ ;
	wire _w1875_ ;
	wire _w1874_ ;
	wire _w1873_ ;
	wire _w1872_ ;
	wire _w1871_ ;
	wire _w1870_ ;
	wire _w1869_ ;
	wire _w1868_ ;
	wire _w1867_ ;
	wire _w1866_ ;
	wire _w1865_ ;
	wire _w1864_ ;
	wire _w1863_ ;
	wire _w1862_ ;
	wire _w1861_ ;
	wire _w1860_ ;
	wire _w1859_ ;
	wire _w1858_ ;
	wire _w1857_ ;
	wire _w1856_ ;
	wire _w1855_ ;
	wire _w1854_ ;
	wire _w1853_ ;
	wire _w1852_ ;
	wire _w1851_ ;
	wire _w1850_ ;
	wire _w1849_ ;
	wire _w1848_ ;
	wire _w1847_ ;
	wire _w1846_ ;
	wire _w1845_ ;
	wire _w1844_ ;
	wire _w1843_ ;
	wire _w1842_ ;
	wire _w1841_ ;
	wire _w1840_ ;
	wire _w1839_ ;
	wire _w1838_ ;
	wire _w1837_ ;
	wire _w1836_ ;
	wire _w1835_ ;
	wire _w1834_ ;
	wire _w1833_ ;
	wire _w1832_ ;
	wire _w1831_ ;
	wire _w1830_ ;
	wire _w1829_ ;
	wire _w1828_ ;
	wire _w1827_ ;
	wire _w1826_ ;
	wire _w1825_ ;
	wire _w1824_ ;
	wire _w1823_ ;
	wire _w1822_ ;
	wire _w1821_ ;
	wire _w1820_ ;
	wire _w1819_ ;
	wire _w1818_ ;
	wire _w1817_ ;
	wire _w1816_ ;
	wire _w1815_ ;
	wire _w1814_ ;
	wire _w1813_ ;
	wire _w1812_ ;
	wire _w1811_ ;
	wire _w1810_ ;
	wire _w1809_ ;
	wire _w1808_ ;
	wire _w1807_ ;
	wire _w1806_ ;
	wire _w1805_ ;
	wire _w1804_ ;
	wire _w1803_ ;
	wire _w1802_ ;
	wire _w1801_ ;
	wire _w1800_ ;
	wire _w1799_ ;
	wire _w1798_ ;
	wire _w1797_ ;
	wire _w1796_ ;
	wire _w1795_ ;
	wire _w1794_ ;
	wire _w1793_ ;
	wire _w1792_ ;
	wire _w1791_ ;
	wire _w1790_ ;
	wire _w1789_ ;
	wire _w1788_ ;
	wire _w1787_ ;
	wire _w1786_ ;
	wire _w1785_ ;
	wire _w1784_ ;
	wire _w1783_ ;
	wire _w1782_ ;
	wire _w1781_ ;
	wire _w1780_ ;
	wire _w1779_ ;
	wire _w1778_ ;
	wire _w1777_ ;
	wire _w1776_ ;
	wire _w1775_ ;
	wire _w1774_ ;
	wire _w1773_ ;
	wire _w1772_ ;
	wire _w1771_ ;
	wire _w1770_ ;
	wire _w1769_ ;
	wire _w1768_ ;
	wire _w1767_ ;
	wire _w1766_ ;
	wire _w1765_ ;
	wire _w1764_ ;
	wire _w1763_ ;
	wire _w1762_ ;
	wire _w1761_ ;
	wire _w1760_ ;
	wire _w1759_ ;
	wire _w1758_ ;
	wire _w1757_ ;
	wire _w1756_ ;
	wire _w1755_ ;
	wire _w1754_ ;
	wire _w1753_ ;
	wire _w1752_ ;
	wire _w1751_ ;
	wire _w1750_ ;
	wire _w1749_ ;
	wire _w1748_ ;
	wire _w1747_ ;
	wire _w1746_ ;
	wire _w1745_ ;
	wire _w1744_ ;
	wire _w1743_ ;
	wire _w1742_ ;
	wire _w1741_ ;
	wire _w1740_ ;
	wire _w1739_ ;
	wire _w1738_ ;
	wire _w1737_ ;
	wire _w1736_ ;
	wire _w1735_ ;
	wire _w1734_ ;
	wire _w1733_ ;
	wire _w1732_ ;
	wire _w1731_ ;
	wire _w1730_ ;
	wire _w1729_ ;
	wire _w1728_ ;
	wire _w1727_ ;
	wire _w1726_ ;
	wire _w1725_ ;
	wire _w1724_ ;
	wire _w1723_ ;
	wire _w1722_ ;
	wire _w1721_ ;
	wire _w1720_ ;
	wire _w1719_ ;
	wire _w1718_ ;
	wire _w1717_ ;
	wire _w1716_ ;
	wire _w1715_ ;
	wire _w1714_ ;
	wire _w1713_ ;
	wire _w1712_ ;
	wire _w1711_ ;
	wire _w1710_ ;
	wire _w1709_ ;
	wire _w1708_ ;
	wire _w1707_ ;
	wire _w1706_ ;
	wire _w1705_ ;
	wire _w1704_ ;
	wire _w1703_ ;
	wire _w1702_ ;
	wire _w1701_ ;
	wire _w1700_ ;
	wire _w1699_ ;
	wire _w1698_ ;
	wire _w1697_ ;
	wire _w1696_ ;
	wire _w1695_ ;
	wire _w1694_ ;
	wire _w1693_ ;
	wire _w1692_ ;
	wire _w1691_ ;
	wire _w1690_ ;
	wire _w1689_ ;
	wire _w1688_ ;
	wire _w1687_ ;
	wire _w1686_ ;
	wire _w1685_ ;
	wire _w1684_ ;
	wire _w1683_ ;
	wire _w1682_ ;
	wire _w1681_ ;
	wire _w1680_ ;
	wire _w1679_ ;
	wire _w1678_ ;
	wire _w1677_ ;
	wire _w1676_ ;
	wire _w1675_ ;
	wire _w1674_ ;
	wire _w1673_ ;
	wire _w1672_ ;
	wire _w1671_ ;
	wire _w1670_ ;
	wire _w1669_ ;
	wire _w1668_ ;
	wire _w1667_ ;
	wire _w1666_ ;
	wire _w1665_ ;
	wire _w1664_ ;
	wire _w1663_ ;
	wire _w1662_ ;
	wire _w1661_ ;
	wire _w1660_ ;
	wire _w1659_ ;
	wire _w1658_ ;
	wire _w1657_ ;
	wire _w1656_ ;
	wire _w1655_ ;
	wire _w1654_ ;
	wire _w1653_ ;
	wire _w1652_ ;
	wire _w1651_ ;
	wire _w1650_ ;
	wire _w1649_ ;
	wire _w1648_ ;
	wire _w1647_ ;
	wire _w1646_ ;
	wire _w1645_ ;
	wire _w1644_ ;
	wire _w1643_ ;
	wire _w1642_ ;
	wire _w1641_ ;
	wire _w1640_ ;
	wire _w1639_ ;
	wire _w1638_ ;
	wire _w1637_ ;
	wire _w1636_ ;
	wire _w1635_ ;
	wire _w1634_ ;
	wire _w1633_ ;
	wire _w1632_ ;
	wire _w1631_ ;
	wire _w1630_ ;
	wire _w1629_ ;
	wire _w1628_ ;
	wire _w1627_ ;
	wire _w1626_ ;
	wire _w1625_ ;
	wire _w1624_ ;
	wire _w1623_ ;
	wire _w1622_ ;
	wire _w1621_ ;
	wire _w1620_ ;
	wire _w1619_ ;
	wire _w1618_ ;
	wire _w1617_ ;
	wire _w1616_ ;
	wire _w1615_ ;
	wire _w1614_ ;
	wire _w1613_ ;
	wire _w1612_ ;
	wire _w1611_ ;
	wire _w1610_ ;
	wire _w1609_ ;
	wire _w1608_ ;
	wire _w1607_ ;
	wire _w1606_ ;
	wire _w1605_ ;
	wire _w1604_ ;
	wire _w1603_ ;
	wire _w1602_ ;
	wire _w1601_ ;
	wire _w1600_ ;
	wire _w1599_ ;
	wire _w1598_ ;
	wire _w1597_ ;
	wire _w1596_ ;
	wire _w1595_ ;
	wire _w1594_ ;
	wire _w1593_ ;
	wire _w1592_ ;
	wire _w1591_ ;
	wire _w1590_ ;
	wire _w1589_ ;
	wire _w1588_ ;
	wire _w1587_ ;
	wire _w1586_ ;
	wire _w1585_ ;
	wire _w1584_ ;
	wire _w1583_ ;
	wire _w1582_ ;
	wire _w1581_ ;
	wire _w1580_ ;
	wire _w1579_ ;
	wire _w1578_ ;
	wire _w1577_ ;
	wire _w1576_ ;
	wire _w1575_ ;
	wire _w1574_ ;
	wire _w1573_ ;
	wire _w1572_ ;
	wire _w1571_ ;
	wire _w1570_ ;
	wire _w1569_ ;
	wire _w1568_ ;
	wire _w1567_ ;
	wire _w1566_ ;
	wire _w1565_ ;
	wire _w1564_ ;
	wire _w1563_ ;
	wire _w1562_ ;
	wire _w1561_ ;
	wire _w1560_ ;
	wire _w1559_ ;
	wire _w1558_ ;
	wire _w1557_ ;
	wire _w1556_ ;
	wire _w1555_ ;
	wire _w1554_ ;
	wire _w1553_ ;
	wire _w1552_ ;
	wire _w1551_ ;
	wire _w1550_ ;
	wire _w1549_ ;
	wire _w1548_ ;
	wire _w1547_ ;
	wire _w1546_ ;
	wire _w1545_ ;
	wire _w1544_ ;
	wire _w1543_ ;
	wire _w1542_ ;
	wire _w1541_ ;
	wire _w1540_ ;
	wire _w1539_ ;
	wire _w1538_ ;
	wire _w1537_ ;
	wire _w1536_ ;
	wire _w1535_ ;
	wire _w1534_ ;
	wire _w1533_ ;
	wire _w1532_ ;
	wire _w1531_ ;
	wire _w1530_ ;
	wire _w1529_ ;
	wire _w1528_ ;
	wire _w1527_ ;
	wire _w1526_ ;
	wire _w1525_ ;
	wire _w1524_ ;
	wire _w1523_ ;
	wire _w1522_ ;
	wire _w1521_ ;
	wire _w1520_ ;
	wire _w1519_ ;
	wire _w1518_ ;
	wire _w1517_ ;
	wire _w1516_ ;
	wire _w1515_ ;
	wire _w1514_ ;
	wire _w1513_ ;
	wire _w1512_ ;
	wire _w1511_ ;
	wire _w1510_ ;
	wire _w1509_ ;
	wire _w1508_ ;
	wire _w1507_ ;
	wire _w1506_ ;
	wire _w1505_ ;
	wire _w1504_ ;
	wire _w1503_ ;
	wire _w1502_ ;
	wire _w1501_ ;
	wire _w1500_ ;
	wire _w1499_ ;
	wire _w1498_ ;
	wire _w1497_ ;
	wire _w1496_ ;
	wire _w1495_ ;
	wire _w1494_ ;
	wire _w1493_ ;
	wire _w1492_ ;
	wire _w1491_ ;
	wire _w1490_ ;
	wire _w1489_ ;
	wire _w1488_ ;
	wire _w1487_ ;
	wire _w1486_ ;
	wire _w1485_ ;
	wire _w1484_ ;
	wire _w1483_ ;
	wire _w1482_ ;
	wire _w1481_ ;
	wire _w1480_ ;
	wire _w1479_ ;
	wire _w1478_ ;
	wire _w1477_ ;
	wire _w1476_ ;
	wire _w1475_ ;
	wire _w1474_ ;
	wire _w1473_ ;
	wire _w1472_ ;
	wire _w1471_ ;
	wire _w1470_ ;
	wire _w1469_ ;
	wire _w1468_ ;
	wire _w1467_ ;
	wire _w1466_ ;
	wire _w1465_ ;
	wire _w1464_ ;
	wire _w1463_ ;
	wire _w1462_ ;
	wire _w1461_ ;
	wire _w1460_ ;
	wire _w1459_ ;
	wire _w1458_ ;
	wire _w1457_ ;
	wire _w1456_ ;
	wire _w1455_ ;
	wire _w1454_ ;
	wire _w1453_ ;
	wire _w1452_ ;
	wire _w1451_ ;
	wire _w1450_ ;
	wire _w1449_ ;
	wire _w1448_ ;
	wire _w1447_ ;
	wire _w1446_ ;
	wire _w1445_ ;
	wire _w1444_ ;
	wire _w1443_ ;
	wire _w1442_ ;
	wire _w1441_ ;
	wire _w1440_ ;
	wire _w1439_ ;
	wire _w1438_ ;
	wire _w1437_ ;
	wire _w1436_ ;
	wire _w1435_ ;
	wire _w1434_ ;
	wire _w1433_ ;
	wire _w1432_ ;
	wire _w1431_ ;
	wire _w1430_ ;
	wire _w1429_ ;
	wire _w1428_ ;
	wire _w1427_ ;
	wire _w1426_ ;
	wire _w1425_ ;
	wire _w1424_ ;
	wire _w1423_ ;
	wire _w1422_ ;
	wire _w1421_ ;
	wire _w1420_ ;
	wire _w1419_ ;
	wire _w1418_ ;
	wire _w1417_ ;
	wire _w1416_ ;
	wire _w1415_ ;
	wire _w1414_ ;
	wire _w1413_ ;
	wire _w1412_ ;
	wire _w1411_ ;
	wire _w1410_ ;
	wire _w1409_ ;
	wire _w1408_ ;
	wire _w1407_ ;
	wire _w1406_ ;
	wire _w1405_ ;
	wire _w1404_ ;
	wire _w1403_ ;
	wire _w1402_ ;
	wire _w1401_ ;
	wire _w1400_ ;
	wire _w1399_ ;
	wire _w1398_ ;
	wire _w1397_ ;
	wire _w1396_ ;
	wire _w1395_ ;
	wire _w1394_ ;
	wire _w1393_ ;
	wire _w1392_ ;
	wire _w1391_ ;
	wire _w1390_ ;
	wire _w1389_ ;
	wire _w1388_ ;
	wire _w1387_ ;
	wire _w1386_ ;
	wire _w1385_ ;
	wire _w1384_ ;
	wire _w1383_ ;
	wire _w1382_ ;
	wire _w1381_ ;
	wire _w1380_ ;
	wire _w1379_ ;
	wire _w1378_ ;
	wire _w1377_ ;
	wire _w1376_ ;
	wire _w1375_ ;
	wire _w1374_ ;
	wire _w1373_ ;
	wire _w1372_ ;
	wire _w1371_ ;
	wire _w1370_ ;
	wire _w1369_ ;
	wire _w1368_ ;
	wire _w1367_ ;
	wire _w1366_ ;
	wire _w1365_ ;
	wire _w1364_ ;
	wire _w1363_ ;
	wire _w1362_ ;
	wire _w1361_ ;
	wire _w1360_ ;
	wire _w1359_ ;
	wire _w1358_ ;
	wire _w1357_ ;
	wire _w1356_ ;
	wire _w1355_ ;
	wire _w1354_ ;
	wire _w1353_ ;
	wire _w1352_ ;
	wire _w1351_ ;
	wire _w1350_ ;
	wire _w1349_ ;
	wire _w1348_ ;
	wire _w1347_ ;
	wire _w1346_ ;
	wire _w1345_ ;
	wire _w1344_ ;
	wire _w1343_ ;
	wire _w1342_ ;
	wire _w1341_ ;
	wire _w1340_ ;
	wire _w1339_ ;
	wire _w1338_ ;
	wire _w1337_ ;
	wire _w1336_ ;
	wire _w1335_ ;
	wire _w1334_ ;
	wire _w1333_ ;
	wire _w1332_ ;
	wire _w1331_ ;
	wire _w1330_ ;
	wire _w1329_ ;
	wire _w1328_ ;
	wire _w1327_ ;
	wire _w1326_ ;
	wire _w1325_ ;
	wire _w1324_ ;
	wire _w1323_ ;
	wire _w1322_ ;
	wire _w1321_ ;
	wire _w1320_ ;
	wire _w1319_ ;
	wire _w1318_ ;
	wire _w1317_ ;
	wire _w1316_ ;
	wire _w1315_ ;
	wire _w1314_ ;
	wire _w1313_ ;
	wire _w1312_ ;
	wire _w1311_ ;
	wire _w1310_ ;
	wire _w1309_ ;
	wire _w1308_ ;
	wire _w1307_ ;
	wire _w1306_ ;
	wire _w1305_ ;
	wire _w1304_ ;
	wire _w1303_ ;
	wire _w1302_ ;
	wire _w1301_ ;
	wire _w1300_ ;
	wire _w1299_ ;
	wire _w1298_ ;
	wire _w1297_ ;
	wire _w1296_ ;
	wire _w1295_ ;
	wire _w1294_ ;
	wire _w1293_ ;
	wire _w1292_ ;
	wire _w1291_ ;
	wire _w1290_ ;
	wire _w1289_ ;
	wire _w1288_ ;
	wire _w1287_ ;
	wire _w1286_ ;
	wire _w1285_ ;
	wire _w1284_ ;
	wire _w1283_ ;
	wire _w1282_ ;
	wire _w1281_ ;
	wire _w1280_ ;
	wire _w1279_ ;
	wire _w1278_ ;
	wire _w1277_ ;
	wire _w1276_ ;
	wire _w1275_ ;
	wire _w1274_ ;
	wire _w1273_ ;
	wire _w1272_ ;
	wire _w1271_ ;
	wire _w1270_ ;
	wire _w1269_ ;
	wire _w1268_ ;
	wire _w1267_ ;
	wire _w1266_ ;
	wire _w1265_ ;
	wire _w1264_ ;
	wire _w1263_ ;
	wire _w1262_ ;
	wire _w1261_ ;
	wire _w1260_ ;
	wire _w1259_ ;
	wire _w1258_ ;
	wire _w1257_ ;
	wire _w1256_ ;
	wire _w1255_ ;
	wire _w1254_ ;
	wire _w1253_ ;
	wire _w1252_ ;
	wire _w1251_ ;
	wire _w1250_ ;
	wire _w1249_ ;
	wire _w1248_ ;
	wire _w1247_ ;
	wire _w1246_ ;
	wire _w1245_ ;
	wire _w1244_ ;
	wire _w1243_ ;
	wire _w1242_ ;
	wire _w1241_ ;
	wire _w1240_ ;
	wire _w1239_ ;
	wire _w1238_ ;
	wire _w1237_ ;
	wire _w1236_ ;
	wire _w1235_ ;
	wire _w1234_ ;
	wire _w1233_ ;
	wire _w1232_ ;
	wire _w1231_ ;
	wire _w1230_ ;
	wire _w1229_ ;
	wire _w1228_ ;
	wire _w1227_ ;
	wire _w1226_ ;
	wire _w1225_ ;
	wire _w1224_ ;
	wire _w1223_ ;
	wire _w1222_ ;
	wire _w1221_ ;
	wire _w1220_ ;
	wire _w1219_ ;
	wire _w1218_ ;
	wire _w1217_ ;
	wire _w1216_ ;
	wire _w1215_ ;
	wire _w1214_ ;
	wire _w1213_ ;
	wire _w1212_ ;
	wire _w1211_ ;
	wire _w1210_ ;
	wire _w1209_ ;
	wire _w1208_ ;
	wire _w1207_ ;
	wire _w1206_ ;
	wire _w1205_ ;
	wire _w1204_ ;
	wire _w1203_ ;
	wire _w1202_ ;
	wire _w1201_ ;
	wire _w1200_ ;
	wire _w1199_ ;
	wire _w1198_ ;
	wire _w1197_ ;
	wire _w1196_ ;
	wire _w1195_ ;
	wire _w1194_ ;
	wire _w1193_ ;
	wire _w1192_ ;
	wire _w1191_ ;
	wire _w1190_ ;
	wire _w1189_ ;
	wire _w1188_ ;
	wire _w1187_ ;
	wire _w1186_ ;
	wire _w1185_ ;
	wire _w1184_ ;
	wire _w1183_ ;
	wire _w1182_ ;
	wire _w1181_ ;
	wire _w1180_ ;
	wire _w1179_ ;
	wire _w1178_ ;
	wire _w1177_ ;
	wire _w1176_ ;
	wire _w1175_ ;
	wire _w1174_ ;
	wire _w1173_ ;
	wire _w1172_ ;
	wire _w1171_ ;
	wire _w1170_ ;
	wire _w1169_ ;
	wire _w1168_ ;
	wire _w1167_ ;
	wire _w1166_ ;
	wire _w1165_ ;
	wire _w1164_ ;
	wire _w1163_ ;
	wire _w1162_ ;
	wire _w1161_ ;
	wire _w1160_ ;
	wire _w1159_ ;
	wire _w1158_ ;
	wire _w1157_ ;
	wire _w1156_ ;
	wire _w1155_ ;
	wire _w1154_ ;
	wire _w1153_ ;
	wire _w1152_ ;
	wire _w1151_ ;
	wire _w1150_ ;
	wire _w1149_ ;
	wire _w1148_ ;
	wire _w1147_ ;
	wire _w1146_ ;
	wire _w1145_ ;
	wire _w1144_ ;
	wire _w1143_ ;
	wire _w1142_ ;
	wire _w573_ ;
	wire _w572_ ;
	wire _w571_ ;
	wire _w570_ ;
	wire _w569_ ;
	wire _w568_ ;
	wire _w567_ ;
	wire _w566_ ;
	wire _w565_ ;
	wire _w564_ ;
	wire _w563_ ;
	wire _w562_ ;
	wire _w561_ ;
	wire _w560_ ;
	wire _w559_ ;
	wire _w558_ ;
	wire _w557_ ;
	wire _w556_ ;
	wire _w555_ ;
	wire _w554_ ;
	wire _w553_ ;
	wire _w552_ ;
	wire _w551_ ;
	wire _w550_ ;
	wire _w549_ ;
	wire _w548_ ;
	wire _w547_ ;
	wire _w546_ ;
	wire _w545_ ;
	wire _w544_ ;
	wire _w543_ ;
	wire _w542_ ;
	wire _w541_ ;
	wire _w540_ ;
	wire _w539_ ;
	wire _w538_ ;
	wire _w537_ ;
	wire _w536_ ;
	wire _w535_ ;
	wire _w534_ ;
	wire _w533_ ;
	wire _w532_ ;
	wire _w531_ ;
	wire _w530_ ;
	wire _w529_ ;
	wire _w528_ ;
	wire _w527_ ;
	wire _w526_ ;
	wire _w525_ ;
	wire _w524_ ;
	wire _w523_ ;
	wire _w522_ ;
	wire _w521_ ;
	wire _w520_ ;
	wire _w519_ ;
	wire _w518_ ;
	wire _w517_ ;
	wire _w516_ ;
	wire _w515_ ;
	wire _w514_ ;
	wire _w513_ ;
	wire _w512_ ;
	wire _w511_ ;
	wire _w510_ ;
	wire _w509_ ;
	wire _w508_ ;
	wire _w507_ ;
	wire _w506_ ;
	wire _w505_ ;
	wire _w504_ ;
	wire _w503_ ;
	wire _w502_ ;
	wire _w501_ ;
	wire _w500_ ;
	wire _w499_ ;
	wire _w498_ ;
	wire _w497_ ;
	wire _w496_ ;
	wire _w495_ ;
	wire _w494_ ;
	wire _w493_ ;
	wire _w492_ ;
	wire _w491_ ;
	wire _w490_ ;
	wire _w489_ ;
	wire _w488_ ;
	wire _w487_ ;
	wire _w486_ ;
	wire _w485_ ;
	wire _w484_ ;
	wire _w483_ ;
	wire _w482_ ;
	wire _w481_ ;
	wire _w480_ ;
	wire _w479_ ;
	wire _w478_ ;
	wire _w477_ ;
	wire _w476_ ;
	wire _w475_ ;
	wire _w474_ ;
	wire _w473_ ;
	wire _w472_ ;
	wire _w471_ ;
	wire _w470_ ;
	wire _w469_ ;
	wire _w468_ ;
	wire _w467_ ;
	wire _w466_ ;
	wire _w465_ ;
	wire _w464_ ;
	wire _w463_ ;
	wire _w462_ ;
	wire _w461_ ;
	wire _w460_ ;
	wire _w459_ ;
	wire _w458_ ;
	wire _w457_ ;
	wire _w456_ ;
	wire _w455_ ;
	wire _w454_ ;
	wire _w453_ ;
	wire _w452_ ;
	wire _w451_ ;
	wire _w450_ ;
	wire _w449_ ;
	wire _w448_ ;
	wire _w447_ ;
	wire _w446_ ;
	wire _w445_ ;
	wire _w444_ ;
	wire _w443_ ;
	wire _w442_ ;
	wire _w441_ ;
	wire _w440_ ;
	wire _w439_ ;
	wire _w438_ ;
	wire _w437_ ;
	wire _w436_ ;
	wire _w435_ ;
	wire _w434_ ;
	wire _w433_ ;
	wire _w432_ ;
	wire _w431_ ;
	wire _w430_ ;
	wire _w429_ ;
	wire _w428_ ;
	wire _w427_ ;
	wire _w426_ ;
	wire _w425_ ;
	wire _w424_ ;
	wire _w423_ ;
	wire _w422_ ;
	wire _w421_ ;
	wire _w420_ ;
	wire _w419_ ;
	wire _w418_ ;
	wire _w417_ ;
	wire _w416_ ;
	wire _w415_ ;
	wire _w414_ ;
	wire _w413_ ;
	wire _w412_ ;
	wire _w411_ ;
	wire _w410_ ;
	wire _w409_ ;
	wire _w408_ ;
	wire _w407_ ;
	wire _w406_ ;
	wire _w405_ ;
	wire _w404_ ;
	wire _w403_ ;
	wire _w402_ ;
	wire _w401_ ;
	wire _w400_ ;
	wire _w399_ ;
	wire _w398_ ;
	wire _w397_ ;
	wire _w396_ ;
	wire _w395_ ;
	wire _w394_ ;
	wire _w393_ ;
	wire _w392_ ;
	wire _w391_ ;
	wire _w390_ ;
	wire _w389_ ;
	wire _w388_ ;
	wire _w387_ ;
	wire _w386_ ;
	wire _w385_ ;
	wire _w384_ ;
	wire _w383_ ;
	wire _w382_ ;
	wire _w381_ ;
	wire _w380_ ;
	wire _w379_ ;
	wire _w378_ ;
	wire _w377_ ;
	wire _w376_ ;
	wire _w375_ ;
	wire _w374_ ;
	wire _w373_ ;
	wire _w372_ ;
	wire _w371_ ;
	wire _w370_ ;
	wire _w369_ ;
	wire _w368_ ;
	wire _w367_ ;
	wire _w366_ ;
	wire _w365_ ;
	wire _w364_ ;
	wire _w363_ ;
	wire _w362_ ;
	wire _w361_ ;
	wire _w360_ ;
	wire _w359_ ;
	wire _w358_ ;
	wire _w357_ ;
	wire _w356_ ;
	wire _w355_ ;
	wire _w354_ ;
	wire _w353_ ;
	wire _w352_ ;
	wire _w351_ ;
	wire _w350_ ;
	wire _w349_ ;
	wire _w348_ ;
	wire _w347_ ;
	wire _w346_ ;
	wire _w345_ ;
	wire _w344_ ;
	wire _w343_ ;
	wire _w342_ ;
	wire _w341_ ;
	wire _w340_ ;
	wire _w339_ ;
	wire _w338_ ;
	wire _w337_ ;
	wire _w336_ ;
	wire _w335_ ;
	wire _w334_ ;
	wire _w333_ ;
	wire _w332_ ;
	wire _w331_ ;
	wire _w330_ ;
	wire _w329_ ;
	wire _w328_ ;
	wire _w327_ ;
	wire _w326_ ;
	wire _w325_ ;
	wire _w324_ ;
	wire _w323_ ;
	wire _w322_ ;
	wire _w321_ ;
	wire _w320_ ;
	wire _w319_ ;
	wire _w318_ ;
	wire _w317_ ;
	wire _w316_ ;
	wire _w315_ ;
	wire _w314_ ;
	wire _w313_ ;
	wire _w312_ ;
	wire _w311_ ;
	wire _w310_ ;
	wire _w309_ ;
	wire _w308_ ;
	wire _w307_ ;
	wire _w306_ ;
	wire _w305_ ;
	wire _w304_ ;
	wire _w303_ ;
	wire _w302_ ;
	wire _w301_ ;
	wire _w300_ ;
	wire _w299_ ;
	wire _w298_ ;
	wire _w297_ ;
	wire _w296_ ;
	wire _w295_ ;
	wire _w294_ ;
	wire _w293_ ;
	wire _w292_ ;
	wire _w291_ ;
	wire _w290_ ;
	wire _w159_ ;
	wire _w158_ ;
	wire _w157_ ;
	wire _w156_ ;
	wire _w155_ ;
	wire _w154_ ;
	wire _w153_ ;
	wire _w152_ ;
	wire _w151_ ;
	wire _w150_ ;
	wire _w149_ ;
	wire _w148_ ;
	wire _w147_ ;
	wire _w146_ ;
	wire _w145_ ;
	wire _w144_ ;
	wire _w143_ ;
	wire _w142_ ;
	wire _w141_ ;
	wire _w140_ ;
	wire _w139_ ;
	wire _w138_ ;
	wire _w137_ ;
	wire _w136_ ;
	wire _w135_ ;
	wire _w134_ ;
	wire _w133_ ;
	wire _w132_ ;
	wire _w131_ ;
	wire _w130_ ;
	wire _w129_ ;
	wire _w128_ ;
	wire _w127_ ;
	wire _w126_ ;
	wire _w125_ ;
	wire _w124_ ;
	wire _w123_ ;
	wire _w122_ ;
	wire _w121_ ;
	wire _w120_ ;
	wire _w119_ ;
	wire _w118_ ;
	wire _w117_ ;
	wire _w116_ ;
	wire _w115_ ;
	wire _w114_ ;
	wire _w113_ ;
	wire _w112_ ;
	wire _w111_ ;
	wire _w110_ ;
	wire _w109_ ;
	wire _w108_ ;
	wire _w107_ ;
	wire _w106_ ;
	wire _w105_ ;
	wire _w104_ ;
	wire _w103_ ;
	wire _w102_ ;
	wire _w101_ ;
	wire _w100_ ;
	wire _w99_ ;
	wire _w98_ ;
	wire _w97_ ;
	wire _w96_ ;
	wire _w95_ ;
	wire _w94_ ;
	wire _w93_ ;
	wire _w92_ ;
	wire _w61_ ;
	wire _w60_ ;
	wire _w59_ ;
	wire _w58_ ;
	wire _w57_ ;
	wire _w56_ ;
	wire _w55_ ;
	wire _w54_ ;
	wire _w53_ ;
	wire _w52_ ;
	wire _w51_ ;
	wire _w50_ ;
	wire _w49_ ;
	wire _w48_ ;
	wire _w47_ ;
	wire _w46_ ;
	wire _w33_ ;
	wire _w34_ ;
	wire _w35_ ;
	wire _w36_ ;
	wire _w37_ ;
	wire _w38_ ;
	wire _w39_ ;
	wire _w40_ ;
	wire _w41_ ;
	wire _w42_ ;
	wire _w43_ ;
	wire _w44_ ;
	wire _w45_ ;
	wire _w62_ ;
	wire _w63_ ;
	wire _w64_ ;
	wire _w65_ ;
	wire _w66_ ;
	wire _w67_ ;
	wire _w68_ ;
	wire _w69_ ;
	wire _w70_ ;
	wire _w71_ ;
	wire _w72_ ;
	wire _w73_ ;
	wire _w74_ ;
	wire _w75_ ;
	wire _w76_ ;
	wire _w77_ ;
	wire _w78_ ;
	wire _w79_ ;
	wire _w80_ ;
	wire _w81_ ;
	wire _w82_ ;
	wire _w83_ ;
	wire _w84_ ;
	wire _w85_ ;
	wire _w86_ ;
	wire _w87_ ;
	wire _w88_ ;
	wire _w89_ ;
	wire _w90_ ;
	wire _w91_ ;
	wire _w160_ ;
	wire _w161_ ;
	wire _w162_ ;
	wire _w163_ ;
	wire _w164_ ;
	wire _w165_ ;
	wire _w166_ ;
	wire _w167_ ;
	wire _w168_ ;
	wire _w169_ ;
	wire _w170_ ;
	wire _w171_ ;
	wire _w172_ ;
	wire _w173_ ;
	wire _w174_ ;
	wire _w175_ ;
	wire _w176_ ;
	wire _w177_ ;
	wire _w178_ ;
	wire _w179_ ;
	wire _w180_ ;
	wire _w181_ ;
	wire _w182_ ;
	wire _w183_ ;
	wire _w184_ ;
	wire _w185_ ;
	wire _w186_ ;
	wire _w187_ ;
	wire _w188_ ;
	wire _w189_ ;
	wire _w190_ ;
	wire _w191_ ;
	wire _w192_ ;
	wire _w193_ ;
	wire _w194_ ;
	wire _w195_ ;
	wire _w196_ ;
	wire _w197_ ;
	wire _w198_ ;
	wire _w199_ ;
	wire _w200_ ;
	wire _w201_ ;
	wire _w202_ ;
	wire _w203_ ;
	wire _w204_ ;
	wire _w205_ ;
	wire _w206_ ;
	wire _w207_ ;
	wire _w208_ ;
	wire _w209_ ;
	wire _w210_ ;
	wire _w211_ ;
	wire _w212_ ;
	wire _w213_ ;
	wire _w214_ ;
	wire _w215_ ;
	wire _w216_ ;
	wire _w217_ ;
	wire _w218_ ;
	wire _w219_ ;
	wire _w220_ ;
	wire _w221_ ;
	wire _w222_ ;
	wire _w223_ ;
	wire _w224_ ;
	wire _w225_ ;
	wire _w226_ ;
	wire _w227_ ;
	wire _w228_ ;
	wire _w229_ ;
	wire _w230_ ;
	wire _w231_ ;
	wire _w232_ ;
	wire _w233_ ;
	wire _w234_ ;
	wire _w235_ ;
	wire _w236_ ;
	wire _w237_ ;
	wire _w238_ ;
	wire _w239_ ;
	wire _w240_ ;
	wire _w241_ ;
	wire _w242_ ;
	wire _w243_ ;
	wire _w244_ ;
	wire _w245_ ;
	wire _w246_ ;
	wire _w247_ ;
	wire _w248_ ;
	wire _w249_ ;
	wire _w250_ ;
	wire _w251_ ;
	wire _w252_ ;
	wire _w253_ ;
	wire _w254_ ;
	wire _w255_ ;
	wire _w256_ ;
	wire _w257_ ;
	wire _w258_ ;
	wire _w259_ ;
	wire _w260_ ;
	wire _w261_ ;
	wire _w262_ ;
	wire _w263_ ;
	wire _w264_ ;
	wire _w265_ ;
	wire _w266_ ;
	wire _w267_ ;
	wire _w268_ ;
	wire _w269_ ;
	wire _w270_ ;
	wire _w271_ ;
	wire _w272_ ;
	wire _w273_ ;
	wire _w274_ ;
	wire _w275_ ;
	wire _w276_ ;
	wire _w277_ ;
	wire _w278_ ;
	wire _w279_ ;
	wire _w280_ ;
	wire _w281_ ;
	wire _w282_ ;
	wire _w283_ ;
	wire _w284_ ;
	wire _w285_ ;
	wire _w286_ ;
	wire _w287_ ;
	wire _w288_ ;
	wire _w289_ ;
	wire _w574_ ;
	wire _w575_ ;
	wire _w576_ ;
	wire _w577_ ;
	wire _w578_ ;
	wire _w579_ ;
	wire _w580_ ;
	wire _w581_ ;
	wire _w582_ ;
	wire _w583_ ;
	wire _w584_ ;
	wire _w585_ ;
	wire _w586_ ;
	wire _w587_ ;
	wire _w588_ ;
	wire _w589_ ;
	wire _w590_ ;
	wire _w591_ ;
	wire _w592_ ;
	wire _w593_ ;
	wire _w594_ ;
	wire _w595_ ;
	wire _w596_ ;
	wire _w597_ ;
	wire _w598_ ;
	wire _w599_ ;
	wire _w600_ ;
	wire _w601_ ;
	wire _w602_ ;
	wire _w603_ ;
	wire _w604_ ;
	wire _w605_ ;
	wire _w606_ ;
	wire _w607_ ;
	wire _w608_ ;
	wire _w609_ ;
	wire _w610_ ;
	wire _w611_ ;
	wire _w612_ ;
	wire _w613_ ;
	wire _w614_ ;
	wire _w615_ ;
	wire _w616_ ;
	wire _w617_ ;
	wire _w618_ ;
	wire _w619_ ;
	wire _w620_ ;
	wire _w621_ ;
	wire _w622_ ;
	wire _w623_ ;
	wire _w624_ ;
	wire _w625_ ;
	wire _w626_ ;
	wire _w627_ ;
	wire _w628_ ;
	wire _w629_ ;
	wire _w630_ ;
	wire _w631_ ;
	wire _w632_ ;
	wire _w633_ ;
	wire _w634_ ;
	wire _w635_ ;
	wire _w636_ ;
	wire _w637_ ;
	wire _w638_ ;
	wire _w639_ ;
	wire _w640_ ;
	wire _w641_ ;
	wire _w642_ ;
	wire _w643_ ;
	wire _w644_ ;
	wire _w645_ ;
	wire _w646_ ;
	wire _w647_ ;
	wire _w648_ ;
	wire _w649_ ;
	wire _w650_ ;
	wire _w651_ ;
	wire _w652_ ;
	wire _w653_ ;
	wire _w654_ ;
	wire _w655_ ;
	wire _w656_ ;
	wire _w657_ ;
	wire _w658_ ;
	wire _w659_ ;
	wire _w660_ ;
	wire _w661_ ;
	wire _w662_ ;
	wire _w663_ ;
	wire _w664_ ;
	wire _w665_ ;
	wire _w666_ ;
	wire _w667_ ;
	wire _w668_ ;
	wire _w669_ ;
	wire _w670_ ;
	wire _w671_ ;
	wire _w672_ ;
	wire _w673_ ;
	wire _w674_ ;
	wire _w675_ ;
	wire _w676_ ;
	wire _w677_ ;
	wire _w678_ ;
	wire _w679_ ;
	wire _w680_ ;
	wire _w681_ ;
	wire _w682_ ;
	wire _w683_ ;
	wire _w684_ ;
	wire _w685_ ;
	wire _w686_ ;
	wire _w687_ ;
	wire _w688_ ;
	wire _w689_ ;
	wire _w690_ ;
	wire _w691_ ;
	wire _w692_ ;
	wire _w693_ ;
	wire _w694_ ;
	wire _w695_ ;
	wire _w696_ ;
	wire _w697_ ;
	wire _w698_ ;
	wire _w699_ ;
	wire _w700_ ;
	wire _w701_ ;
	wire _w702_ ;
	wire _w703_ ;
	wire _w704_ ;
	wire _w705_ ;
	wire _w706_ ;
	wire _w707_ ;
	wire _w708_ ;
	wire _w709_ ;
	wire _w710_ ;
	wire _w711_ ;
	wire _w712_ ;
	wire _w713_ ;
	wire _w714_ ;
	wire _w715_ ;
	wire _w716_ ;
	wire _w717_ ;
	wire _w718_ ;
	wire _w719_ ;
	wire _w720_ ;
	wire _w721_ ;
	wire _w722_ ;
	wire _w723_ ;
	wire _w724_ ;
	wire _w725_ ;
	wire _w726_ ;
	wire _w727_ ;
	wire _w728_ ;
	wire _w729_ ;
	wire _w730_ ;
	wire _w731_ ;
	wire _w732_ ;
	wire _w733_ ;
	wire _w734_ ;
	wire _w735_ ;
	wire _w736_ ;
	wire _w737_ ;
	wire _w738_ ;
	wire _w739_ ;
	wire _w740_ ;
	wire _w741_ ;
	wire _w742_ ;
	wire _w743_ ;
	wire _w744_ ;
	wire _w745_ ;
	wire _w746_ ;
	wire _w747_ ;
	wire _w748_ ;
	wire _w749_ ;
	wire _w750_ ;
	wire _w751_ ;
	wire _w752_ ;
	wire _w753_ ;
	wire _w754_ ;
	wire _w755_ ;
	wire _w756_ ;
	wire _w757_ ;
	wire _w758_ ;
	wire _w759_ ;
	wire _w760_ ;
	wire _w761_ ;
	wire _w762_ ;
	wire _w763_ ;
	wire _w764_ ;
	wire _w765_ ;
	wire _w766_ ;
	wire _w767_ ;
	wire _w768_ ;
	wire _w769_ ;
	wire _w770_ ;
	wire _w771_ ;
	wire _w772_ ;
	wire _w773_ ;
	wire _w774_ ;
	wire _w775_ ;
	wire _w776_ ;
	wire _w777_ ;
	wire _w778_ ;
	wire _w779_ ;
	wire _w780_ ;
	wire _w781_ ;
	wire _w782_ ;
	wire _w783_ ;
	wire _w784_ ;
	wire _w785_ ;
	wire _w786_ ;
	wire _w787_ ;
	wire _w788_ ;
	wire _w789_ ;
	wire _w790_ ;
	wire _w791_ ;
	wire _w792_ ;
	wire _w793_ ;
	wire _w794_ ;
	wire _w795_ ;
	wire _w796_ ;
	wire _w797_ ;
	wire _w798_ ;
	wire _w799_ ;
	wire _w800_ ;
	wire _w801_ ;
	wire _w802_ ;
	wire _w803_ ;
	wire _w804_ ;
	wire _w805_ ;
	wire _w806_ ;
	wire _w807_ ;
	wire _w808_ ;
	wire _w809_ ;
	wire _w810_ ;
	wire _w811_ ;
	wire _w812_ ;
	wire _w813_ ;
	wire _w814_ ;
	wire _w815_ ;
	wire _w816_ ;
	wire _w817_ ;
	wire _w818_ ;
	wire _w819_ ;
	wire _w820_ ;
	wire _w821_ ;
	wire _w822_ ;
	wire _w823_ ;
	wire _w824_ ;
	wire _w825_ ;
	wire _w826_ ;
	wire _w827_ ;
	wire _w828_ ;
	wire _w829_ ;
	wire _w830_ ;
	wire _w831_ ;
	wire _w832_ ;
	wire _w833_ ;
	wire _w834_ ;
	wire _w835_ ;
	wire _w836_ ;
	wire _w837_ ;
	wire _w838_ ;
	wire _w839_ ;
	wire _w840_ ;
	wire _w841_ ;
	wire _w842_ ;
	wire _w843_ ;
	wire _w844_ ;
	wire _w845_ ;
	wire _w846_ ;
	wire _w847_ ;
	wire _w848_ ;
	wire _w849_ ;
	wire _w850_ ;
	wire _w851_ ;
	wire _w852_ ;
	wire _w853_ ;
	wire _w854_ ;
	wire _w855_ ;
	wire _w856_ ;
	wire _w857_ ;
	wire _w858_ ;
	wire _w859_ ;
	wire _w860_ ;
	wire _w861_ ;
	wire _w862_ ;
	wire _w863_ ;
	wire _w864_ ;
	wire _w865_ ;
	wire _w866_ ;
	wire _w867_ ;
	wire _w868_ ;
	wire _w869_ ;
	wire _w870_ ;
	wire _w871_ ;
	wire _w872_ ;
	wire _w873_ ;
	wire _w874_ ;
	wire _w875_ ;
	wire _w876_ ;
	wire _w877_ ;
	wire _w878_ ;
	wire _w879_ ;
	wire _w880_ ;
	wire _w881_ ;
	wire _w882_ ;
	wire _w883_ ;
	wire _w884_ ;
	wire _w885_ ;
	wire _w886_ ;
	wire _w887_ ;
	wire _w888_ ;
	wire _w889_ ;
	wire _w890_ ;
	wire _w891_ ;
	wire _w892_ ;
	wire _w893_ ;
	wire _w894_ ;
	wire _w895_ ;
	wire _w896_ ;
	wire _w897_ ;
	wire _w898_ ;
	wire _w899_ ;
	wire _w900_ ;
	wire _w901_ ;
	wire _w902_ ;
	wire _w903_ ;
	wire _w904_ ;
	wire _w905_ ;
	wire _w906_ ;
	wire _w907_ ;
	wire _w908_ ;
	wire _w909_ ;
	wire _w910_ ;
	wire _w911_ ;
	wire _w912_ ;
	wire _w913_ ;
	wire _w914_ ;
	wire _w915_ ;
	wire _w916_ ;
	wire _w917_ ;
	wire _w918_ ;
	wire _w919_ ;
	wire _w920_ ;
	wire _w921_ ;
	wire _w922_ ;
	wire _w923_ ;
	wire _w924_ ;
	wire _w925_ ;
	wire _w926_ ;
	wire _w927_ ;
	wire _w928_ ;
	wire _w929_ ;
	wire _w930_ ;
	wire _w931_ ;
	wire _w932_ ;
	wire _w933_ ;
	wire _w934_ ;
	wire _w935_ ;
	wire _w936_ ;
	wire _w937_ ;
	wire _w938_ ;
	wire _w939_ ;
	wire _w940_ ;
	wire _w941_ ;
	wire _w942_ ;
	wire _w943_ ;
	wire _w944_ ;
	wire _w945_ ;
	wire _w946_ ;
	wire _w947_ ;
	wire _w948_ ;
	wire _w949_ ;
	wire _w950_ ;
	wire _w951_ ;
	wire _w952_ ;
	wire _w953_ ;
	wire _w954_ ;
	wire _w955_ ;
	wire _w956_ ;
	wire _w957_ ;
	wire _w958_ ;
	wire _w959_ ;
	wire _w960_ ;
	wire _w961_ ;
	wire _w962_ ;
	wire _w963_ ;
	wire _w964_ ;
	wire _w965_ ;
	wire _w966_ ;
	wire _w967_ ;
	wire _w968_ ;
	wire _w969_ ;
	wire _w970_ ;
	wire _w971_ ;
	wire _w972_ ;
	wire _w973_ ;
	wire _w974_ ;
	wire _w975_ ;
	wire _w976_ ;
	wire _w977_ ;
	wire _w978_ ;
	wire _w979_ ;
	wire _w980_ ;
	wire _w981_ ;
	wire _w982_ ;
	wire _w983_ ;
	wire _w984_ ;
	wire _w985_ ;
	wire _w986_ ;
	wire _w987_ ;
	wire _w988_ ;
	wire _w989_ ;
	wire _w990_ ;
	wire _w991_ ;
	wire _w992_ ;
	wire _w993_ ;
	wire _w994_ ;
	wire _w995_ ;
	wire _w996_ ;
	wire _w997_ ;
	wire _w998_ ;
	wire _w999_ ;
	wire _w1000_ ;
	wire _w1001_ ;
	wire _w1002_ ;
	wire _w1003_ ;
	wire _w1004_ ;
	wire _w1005_ ;
	wire _w1006_ ;
	wire _w1007_ ;
	wire _w1008_ ;
	wire _w1009_ ;
	wire _w1010_ ;
	wire _w1011_ ;
	wire _w1012_ ;
	wire _w1013_ ;
	wire _w1014_ ;
	wire _w1015_ ;
	wire _w1016_ ;
	wire _w1017_ ;
	wire _w1018_ ;
	wire _w1019_ ;
	wire _w1020_ ;
	wire _w1021_ ;
	wire _w1022_ ;
	wire _w1023_ ;
	wire _w1024_ ;
	wire _w1025_ ;
	wire _w1026_ ;
	wire _w1027_ ;
	wire _w1028_ ;
	wire _w1029_ ;
	wire _w1030_ ;
	wire _w1031_ ;
	wire _w1032_ ;
	wire _w1033_ ;
	wire _w1034_ ;
	wire _w1035_ ;
	wire _w1036_ ;
	wire _w1037_ ;
	wire _w1038_ ;
	wire _w1039_ ;
	wire _w1040_ ;
	wire _w1041_ ;
	wire _w1042_ ;
	wire _w1043_ ;
	wire _w1044_ ;
	wire _w1045_ ;
	wire _w1046_ ;
	wire _w1047_ ;
	wire _w1048_ ;
	wire _w1049_ ;
	wire _w1050_ ;
	wire _w1051_ ;
	wire _w1052_ ;
	wire _w1053_ ;
	wire _w1054_ ;
	wire _w1055_ ;
	wire _w1056_ ;
	wire _w1057_ ;
	wire _w1058_ ;
	wire _w1059_ ;
	wire _w1060_ ;
	wire _w1061_ ;
	wire _w1062_ ;
	wire _w1063_ ;
	wire _w1064_ ;
	wire _w1065_ ;
	wire _w1066_ ;
	wire _w1067_ ;
	wire _w1068_ ;
	wire _w1069_ ;
	wire _w1070_ ;
	wire _w1071_ ;
	wire _w1072_ ;
	wire _w1073_ ;
	wire _w1074_ ;
	wire _w1075_ ;
	wire _w1076_ ;
	wire _w1077_ ;
	wire _w1078_ ;
	wire _w1079_ ;
	wire _w1080_ ;
	wire _w1081_ ;
	wire _w1082_ ;
	wire _w1083_ ;
	wire _w1084_ ;
	wire _w1085_ ;
	wire _w1086_ ;
	wire _w1087_ ;
	wire _w1088_ ;
	wire _w1089_ ;
	wire _w1090_ ;
	wire _w1091_ ;
	wire _w1092_ ;
	wire _w1093_ ;
	wire _w1094_ ;
	wire _w1095_ ;
	wire _w1096_ ;
	wire _w1097_ ;
	wire _w1098_ ;
	wire _w1099_ ;
	wire _w1100_ ;
	wire _w1101_ ;
	wire _w1102_ ;
	wire _w1103_ ;
	wire _w1104_ ;
	wire _w1105_ ;
	wire _w1106_ ;
	wire _w1107_ ;
	wire _w1108_ ;
	wire _w1109_ ;
	wire _w1110_ ;
	wire _w1111_ ;
	wire _w1112_ ;
	wire _w1113_ ;
	wire _w1114_ ;
	wire _w1115_ ;
	wire _w1116_ ;
	wire _w1117_ ;
	wire _w1118_ ;
	wire _w1119_ ;
	wire _w1120_ ;
	wire _w1121_ ;
	wire _w1122_ ;
	wire _w1123_ ;
	wire _w1124_ ;
	wire _w1125_ ;
	wire _w1126_ ;
	wire _w1127_ ;
	wire _w1128_ ;
	wire _w1129_ ;
	wire _w1130_ ;
	wire _w1131_ ;
	wire _w1132_ ;
	wire _w1133_ ;
	wire _w1134_ ;
	wire _w1135_ ;
	wire _w1136_ ;
	wire _w1137_ ;
	wire _w1138_ ;
	wire _w1139_ ;
	wire _w1140_ ;
	wire _w1141_ ;
	LUT2 #(
		.INIT('h8)
	) name0 (
		\1GAT(0)_pad ,
		\290GAT(17)_pad ,
		_w33_
	);
	LUT2 #(
		.INIT('h8)
	) name1 (
		\18GAT(1)_pad ,
		\273GAT(16)_pad ,
		_w34_
	);
	LUT2 #(
		.INIT('h1)
	) name2 (
		_w33_,
		_w34_,
		_w35_
	);
	LUT2 #(
		.INIT('h8)
	) name3 (
		_w33_,
		_w34_,
		_w36_
	);
	LUT2 #(
		.INIT('h1)
	) name4 (
		_w35_,
		_w36_,
		_w37_
	);
	LUT2 #(
		.INIT('h8)
	) name5 (
		\1GAT(0)_pad ,
		\307GAT(18)_pad ,
		_w38_
	);
	LUT2 #(
		.INIT('h4)
	) name6 (
		\35GAT(2)_pad ,
		_w36_,
		_w39_
	);
	LUT2 #(
		.INIT('h8)
	) name7 (
		\18GAT(1)_pad ,
		\290GAT(17)_pad ,
		_w40_
	);
	LUT2 #(
		.INIT('h8)
	) name8 (
		\273GAT(16)_pad ,
		\35GAT(2)_pad ,
		_w41_
	);
	LUT2 #(
		.INIT('h4)
	) name9 (
		_w40_,
		_w41_,
		_w42_
	);
	LUT2 #(
		.INIT('h4)
	) name10 (
		\1GAT(0)_pad ,
		_w41_,
		_w43_
	);
	LUT2 #(
		.INIT('h2)
	) name11 (
		_w40_,
		_w43_,
		_w44_
	);
	LUT2 #(
		.INIT('h1)
	) name12 (
		_w42_,
		_w44_,
		_w45_
	);
	LUT2 #(
		.INIT('h1)
	) name13 (
		_w39_,
		_w45_,
		_w46_
	);
	LUT2 #(
		.INIT('h4)
	) name14 (
		_w38_,
		_w46_,
		_w47_
	);
	LUT2 #(
		.INIT('h2)
	) name15 (
		_w38_,
		_w46_,
		_w48_
	);
	LUT2 #(
		.INIT('h1)
	) name16 (
		_w47_,
		_w48_,
		_w49_
	);
	LUT2 #(
		.INIT('h8)
	) name17 (
		\1GAT(0)_pad ,
		\324GAT(19)_pad ,
		_w50_
	);
	LUT2 #(
		.INIT('h1)
	) name18 (
		_w45_,
		_w47_,
		_w51_
	);
	LUT2 #(
		.INIT('h8)
	) name19 (
		\18GAT(1)_pad ,
		\307GAT(18)_pad ,
		_w52_
	);
	LUT2 #(
		.INIT('h4)
	) name20 (
		\52GAT(3)_pad ,
		_w34_,
		_w53_
	);
	LUT2 #(
		.INIT('h8)
	) name21 (
		\273GAT(16)_pad ,
		\52GAT(3)_pad ,
		_w54_
	);
	LUT2 #(
		.INIT('h8)
	) name22 (
		\290GAT(17)_pad ,
		\35GAT(2)_pad ,
		_w55_
	);
	LUT2 #(
		.INIT('h1)
	) name23 (
		_w54_,
		_w55_,
		_w56_
	);
	LUT2 #(
		.INIT('h4)
	) name24 (
		\18GAT(1)_pad ,
		_w54_,
		_w57_
	);
	LUT2 #(
		.INIT('h8)
	) name25 (
		_w55_,
		_w57_,
		_w58_
	);
	LUT2 #(
		.INIT('h1)
	) name26 (
		_w56_,
		_w58_,
		_w59_
	);
	LUT2 #(
		.INIT('h4)
	) name27 (
		_w53_,
		_w59_,
		_w60_
	);
	LUT2 #(
		.INIT('h4)
	) name28 (
		_w52_,
		_w60_,
		_w61_
	);
	LUT2 #(
		.INIT('h2)
	) name29 (
		_w52_,
		_w60_,
		_w62_
	);
	LUT2 #(
		.INIT('h1)
	) name30 (
		_w61_,
		_w62_,
		_w63_
	);
	LUT2 #(
		.INIT('h4)
	) name31 (
		_w51_,
		_w63_,
		_w64_
	);
	LUT2 #(
		.INIT('h2)
	) name32 (
		_w51_,
		_w63_,
		_w65_
	);
	LUT2 #(
		.INIT('h1)
	) name33 (
		_w64_,
		_w65_,
		_w66_
	);
	LUT2 #(
		.INIT('h4)
	) name34 (
		_w50_,
		_w66_,
		_w67_
	);
	LUT2 #(
		.INIT('h2)
	) name35 (
		_w50_,
		_w66_,
		_w68_
	);
	LUT2 #(
		.INIT('h1)
	) name36 (
		_w67_,
		_w68_,
		_w69_
	);
	LUT2 #(
		.INIT('h8)
	) name37 (
		\1GAT(0)_pad ,
		\341GAT(20)_pad ,
		_w70_
	);
	LUT2 #(
		.INIT('h1)
	) name38 (
		_w64_,
		_w67_,
		_w71_
	);
	LUT2 #(
		.INIT('h8)
	) name39 (
		\18GAT(1)_pad ,
		\324GAT(19)_pad ,
		_w72_
	);
	LUT2 #(
		.INIT('h2)
	) name40 (
		_w59_,
		_w61_,
		_w73_
	);
	LUT2 #(
		.INIT('h8)
	) name41 (
		\307GAT(18)_pad ,
		\35GAT(2)_pad ,
		_w74_
	);
	LUT2 #(
		.INIT('h4)
	) name42 (
		\69GAT(4)_pad ,
		_w41_,
		_w75_
	);
	LUT2 #(
		.INIT('h8)
	) name43 (
		\273GAT(16)_pad ,
		\69GAT(4)_pad ,
		_w76_
	);
	LUT2 #(
		.INIT('h8)
	) name44 (
		\290GAT(17)_pad ,
		\52GAT(3)_pad ,
		_w77_
	);
	LUT2 #(
		.INIT('h1)
	) name45 (
		_w76_,
		_w77_,
		_w78_
	);
	LUT2 #(
		.INIT('h4)
	) name46 (
		\35GAT(2)_pad ,
		_w76_,
		_w79_
	);
	LUT2 #(
		.INIT('h8)
	) name47 (
		_w77_,
		_w79_,
		_w80_
	);
	LUT2 #(
		.INIT('h1)
	) name48 (
		_w78_,
		_w80_,
		_w81_
	);
	LUT2 #(
		.INIT('h4)
	) name49 (
		_w75_,
		_w81_,
		_w82_
	);
	LUT2 #(
		.INIT('h4)
	) name50 (
		_w74_,
		_w82_,
		_w83_
	);
	LUT2 #(
		.INIT('h2)
	) name51 (
		_w74_,
		_w82_,
		_w84_
	);
	LUT2 #(
		.INIT('h1)
	) name52 (
		_w83_,
		_w84_,
		_w85_
	);
	LUT2 #(
		.INIT('h4)
	) name53 (
		_w73_,
		_w85_,
		_w86_
	);
	LUT2 #(
		.INIT('h2)
	) name54 (
		_w73_,
		_w85_,
		_w87_
	);
	LUT2 #(
		.INIT('h1)
	) name55 (
		_w86_,
		_w87_,
		_w88_
	);
	LUT2 #(
		.INIT('h4)
	) name56 (
		_w72_,
		_w88_,
		_w89_
	);
	LUT2 #(
		.INIT('h2)
	) name57 (
		_w72_,
		_w88_,
		_w90_
	);
	LUT2 #(
		.INIT('h1)
	) name58 (
		_w89_,
		_w90_,
		_w91_
	);
	LUT2 #(
		.INIT('h4)
	) name59 (
		_w71_,
		_w91_,
		_w92_
	);
	LUT2 #(
		.INIT('h2)
	) name60 (
		_w71_,
		_w91_,
		_w93_
	);
	LUT2 #(
		.INIT('h1)
	) name61 (
		_w92_,
		_w93_,
		_w94_
	);
	LUT2 #(
		.INIT('h4)
	) name62 (
		_w70_,
		_w94_,
		_w95_
	);
	LUT2 #(
		.INIT('h2)
	) name63 (
		_w70_,
		_w94_,
		_w96_
	);
	LUT2 #(
		.INIT('h1)
	) name64 (
		_w95_,
		_w96_,
		_w97_
	);
	LUT2 #(
		.INIT('h8)
	) name65 (
		\1GAT(0)_pad ,
		\358GAT(21)_pad ,
		_w98_
	);
	LUT2 #(
		.INIT('h1)
	) name66 (
		_w92_,
		_w95_,
		_w99_
	);
	LUT2 #(
		.INIT('h8)
	) name67 (
		\18GAT(1)_pad ,
		\341GAT(20)_pad ,
		_w100_
	);
	LUT2 #(
		.INIT('h1)
	) name68 (
		_w86_,
		_w89_,
		_w101_
	);
	LUT2 #(
		.INIT('h8)
	) name69 (
		\324GAT(19)_pad ,
		\35GAT(2)_pad ,
		_w102_
	);
	LUT2 #(
		.INIT('h2)
	) name70 (
		_w81_,
		_w83_,
		_w103_
	);
	LUT2 #(
		.INIT('h8)
	) name71 (
		\307GAT(18)_pad ,
		\52GAT(3)_pad ,
		_w104_
	);
	LUT2 #(
		.INIT('h4)
	) name72 (
		\86GAT(5)_pad ,
		_w54_,
		_w105_
	);
	LUT2 #(
		.INIT('h8)
	) name73 (
		\273GAT(16)_pad ,
		\86GAT(5)_pad ,
		_w106_
	);
	LUT2 #(
		.INIT('h8)
	) name74 (
		\290GAT(17)_pad ,
		\69GAT(4)_pad ,
		_w107_
	);
	LUT2 #(
		.INIT('h1)
	) name75 (
		_w106_,
		_w107_,
		_w108_
	);
	LUT2 #(
		.INIT('h8)
	) name76 (
		\290GAT(17)_pad ,
		\86GAT(5)_pad ,
		_w109_
	);
	LUT2 #(
		.INIT('h8)
	) name77 (
		_w76_,
		_w109_,
		_w110_
	);
	LUT2 #(
		.INIT('h4)
	) name78 (
		\52GAT(3)_pad ,
		_w110_,
		_w111_
	);
	LUT2 #(
		.INIT('h1)
	) name79 (
		_w108_,
		_w111_,
		_w112_
	);
	LUT2 #(
		.INIT('h4)
	) name80 (
		_w105_,
		_w112_,
		_w113_
	);
	LUT2 #(
		.INIT('h4)
	) name81 (
		_w104_,
		_w113_,
		_w114_
	);
	LUT2 #(
		.INIT('h2)
	) name82 (
		_w104_,
		_w113_,
		_w115_
	);
	LUT2 #(
		.INIT('h1)
	) name83 (
		_w114_,
		_w115_,
		_w116_
	);
	LUT2 #(
		.INIT('h4)
	) name84 (
		_w103_,
		_w116_,
		_w117_
	);
	LUT2 #(
		.INIT('h2)
	) name85 (
		_w103_,
		_w116_,
		_w118_
	);
	LUT2 #(
		.INIT('h1)
	) name86 (
		_w117_,
		_w118_,
		_w119_
	);
	LUT2 #(
		.INIT('h4)
	) name87 (
		_w102_,
		_w119_,
		_w120_
	);
	LUT2 #(
		.INIT('h2)
	) name88 (
		_w102_,
		_w119_,
		_w121_
	);
	LUT2 #(
		.INIT('h1)
	) name89 (
		_w120_,
		_w121_,
		_w122_
	);
	LUT2 #(
		.INIT('h4)
	) name90 (
		_w101_,
		_w122_,
		_w123_
	);
	LUT2 #(
		.INIT('h2)
	) name91 (
		_w101_,
		_w122_,
		_w124_
	);
	LUT2 #(
		.INIT('h1)
	) name92 (
		_w123_,
		_w124_,
		_w125_
	);
	LUT2 #(
		.INIT('h4)
	) name93 (
		_w100_,
		_w125_,
		_w126_
	);
	LUT2 #(
		.INIT('h2)
	) name94 (
		_w100_,
		_w125_,
		_w127_
	);
	LUT2 #(
		.INIT('h1)
	) name95 (
		_w126_,
		_w127_,
		_w128_
	);
	LUT2 #(
		.INIT('h4)
	) name96 (
		_w99_,
		_w128_,
		_w129_
	);
	LUT2 #(
		.INIT('h2)
	) name97 (
		_w99_,
		_w128_,
		_w130_
	);
	LUT2 #(
		.INIT('h1)
	) name98 (
		_w129_,
		_w130_,
		_w131_
	);
	LUT2 #(
		.INIT('h4)
	) name99 (
		_w98_,
		_w131_,
		_w132_
	);
	LUT2 #(
		.INIT('h2)
	) name100 (
		_w98_,
		_w131_,
		_w133_
	);
	LUT2 #(
		.INIT('h1)
	) name101 (
		_w132_,
		_w133_,
		_w134_
	);
	LUT2 #(
		.INIT('h8)
	) name102 (
		\1GAT(0)_pad ,
		\375GAT(22)_pad ,
		_w135_
	);
	LUT2 #(
		.INIT('h1)
	) name103 (
		_w129_,
		_w132_,
		_w136_
	);
	LUT2 #(
		.INIT('h8)
	) name104 (
		\18GAT(1)_pad ,
		\358GAT(21)_pad ,
		_w137_
	);
	LUT2 #(
		.INIT('h1)
	) name105 (
		_w123_,
		_w126_,
		_w138_
	);
	LUT2 #(
		.INIT('h8)
	) name106 (
		\341GAT(20)_pad ,
		\35GAT(2)_pad ,
		_w139_
	);
	LUT2 #(
		.INIT('h1)
	) name107 (
		_w117_,
		_w120_,
		_w140_
	);
	LUT2 #(
		.INIT('h8)
	) name108 (
		\324GAT(19)_pad ,
		\52GAT(3)_pad ,
		_w141_
	);
	LUT2 #(
		.INIT('h2)
	) name109 (
		_w112_,
		_w114_,
		_w142_
	);
	LUT2 #(
		.INIT('h8)
	) name110 (
		\307GAT(18)_pad ,
		\69GAT(4)_pad ,
		_w143_
	);
	LUT2 #(
		.INIT('h8)
	) name111 (
		\103GAT(6)_pad ,
		\273GAT(16)_pad ,
		_w144_
	);
	LUT2 #(
		.INIT('h1)
	) name112 (
		_w109_,
		_w144_,
		_w145_
	);
	LUT2 #(
		.INIT('h8)
	) name113 (
		_w109_,
		_w144_,
		_w146_
	);
	LUT2 #(
		.INIT('h1)
	) name114 (
		_w145_,
		_w146_,
		_w147_
	);
	LUT2 #(
		.INIT('h1)
	) name115 (
		_w110_,
		_w147_,
		_w148_
	);
	LUT2 #(
		.INIT('h8)
	) name116 (
		_w110_,
		_w147_,
		_w149_
	);
	LUT2 #(
		.INIT('h1)
	) name117 (
		_w148_,
		_w149_,
		_w150_
	);
	LUT2 #(
		.INIT('h4)
	) name118 (
		_w143_,
		_w150_,
		_w151_
	);
	LUT2 #(
		.INIT('h2)
	) name119 (
		_w143_,
		_w150_,
		_w152_
	);
	LUT2 #(
		.INIT('h1)
	) name120 (
		_w151_,
		_w152_,
		_w153_
	);
	LUT2 #(
		.INIT('h4)
	) name121 (
		_w142_,
		_w153_,
		_w154_
	);
	LUT2 #(
		.INIT('h2)
	) name122 (
		_w142_,
		_w153_,
		_w155_
	);
	LUT2 #(
		.INIT('h1)
	) name123 (
		_w154_,
		_w155_,
		_w156_
	);
	LUT2 #(
		.INIT('h4)
	) name124 (
		_w141_,
		_w156_,
		_w157_
	);
	LUT2 #(
		.INIT('h2)
	) name125 (
		_w141_,
		_w156_,
		_w158_
	);
	LUT2 #(
		.INIT('h1)
	) name126 (
		_w157_,
		_w158_,
		_w159_
	);
	LUT2 #(
		.INIT('h4)
	) name127 (
		_w140_,
		_w159_,
		_w160_
	);
	LUT2 #(
		.INIT('h2)
	) name128 (
		_w140_,
		_w159_,
		_w161_
	);
	LUT2 #(
		.INIT('h1)
	) name129 (
		_w160_,
		_w161_,
		_w162_
	);
	LUT2 #(
		.INIT('h4)
	) name130 (
		_w139_,
		_w162_,
		_w163_
	);
	LUT2 #(
		.INIT('h2)
	) name131 (
		_w139_,
		_w162_,
		_w164_
	);
	LUT2 #(
		.INIT('h1)
	) name132 (
		_w163_,
		_w164_,
		_w165_
	);
	LUT2 #(
		.INIT('h4)
	) name133 (
		_w138_,
		_w165_,
		_w166_
	);
	LUT2 #(
		.INIT('h2)
	) name134 (
		_w138_,
		_w165_,
		_w167_
	);
	LUT2 #(
		.INIT('h1)
	) name135 (
		_w166_,
		_w167_,
		_w168_
	);
	LUT2 #(
		.INIT('h4)
	) name136 (
		_w137_,
		_w168_,
		_w169_
	);
	LUT2 #(
		.INIT('h2)
	) name137 (
		_w137_,
		_w168_,
		_w170_
	);
	LUT2 #(
		.INIT('h1)
	) name138 (
		_w169_,
		_w170_,
		_w171_
	);
	LUT2 #(
		.INIT('h4)
	) name139 (
		_w136_,
		_w171_,
		_w172_
	);
	LUT2 #(
		.INIT('h2)
	) name140 (
		_w136_,
		_w171_,
		_w173_
	);
	LUT2 #(
		.INIT('h1)
	) name141 (
		_w172_,
		_w173_,
		_w174_
	);
	LUT2 #(
		.INIT('h4)
	) name142 (
		_w135_,
		_w174_,
		_w175_
	);
	LUT2 #(
		.INIT('h2)
	) name143 (
		_w135_,
		_w174_,
		_w176_
	);
	LUT2 #(
		.INIT('h1)
	) name144 (
		_w175_,
		_w176_,
		_w177_
	);
	LUT2 #(
		.INIT('h8)
	) name145 (
		\1GAT(0)_pad ,
		\392GAT(23)_pad ,
		_w178_
	);
	LUT2 #(
		.INIT('h1)
	) name146 (
		_w172_,
		_w175_,
		_w179_
	);
	LUT2 #(
		.INIT('h8)
	) name147 (
		\18GAT(1)_pad ,
		\375GAT(22)_pad ,
		_w180_
	);
	LUT2 #(
		.INIT('h1)
	) name148 (
		_w166_,
		_w169_,
		_w181_
	);
	LUT2 #(
		.INIT('h8)
	) name149 (
		\358GAT(21)_pad ,
		\35GAT(2)_pad ,
		_w182_
	);
	LUT2 #(
		.INIT('h1)
	) name150 (
		_w160_,
		_w163_,
		_w183_
	);
	LUT2 #(
		.INIT('h8)
	) name151 (
		\341GAT(20)_pad ,
		\52GAT(3)_pad ,
		_w184_
	);
	LUT2 #(
		.INIT('h1)
	) name152 (
		_w154_,
		_w157_,
		_w185_
	);
	LUT2 #(
		.INIT('h8)
	) name153 (
		\324GAT(19)_pad ,
		\69GAT(4)_pad ,
		_w186_
	);
	LUT2 #(
		.INIT('h1)
	) name154 (
		_w148_,
		_w151_,
		_w187_
	);
	LUT2 #(
		.INIT('h8)
	) name155 (
		\307GAT(18)_pad ,
		\86GAT(5)_pad ,
		_w188_
	);
	LUT2 #(
		.INIT('h4)
	) name156 (
		\120GAT(7)_pad ,
		_w146_,
		_w189_
	);
	LUT2 #(
		.INIT('h8)
	) name157 (
		\103GAT(6)_pad ,
		\290GAT(17)_pad ,
		_w190_
	);
	LUT2 #(
		.INIT('h8)
	) name158 (
		\120GAT(7)_pad ,
		\273GAT(16)_pad ,
		_w191_
	);
	LUT2 #(
		.INIT('h4)
	) name159 (
		_w190_,
		_w191_,
		_w192_
	);
	LUT2 #(
		.INIT('h4)
	) name160 (
		\86GAT(5)_pad ,
		_w191_,
		_w193_
	);
	LUT2 #(
		.INIT('h2)
	) name161 (
		_w190_,
		_w193_,
		_w194_
	);
	LUT2 #(
		.INIT('h1)
	) name162 (
		_w192_,
		_w194_,
		_w195_
	);
	LUT2 #(
		.INIT('h1)
	) name163 (
		_w189_,
		_w195_,
		_w196_
	);
	LUT2 #(
		.INIT('h4)
	) name164 (
		_w188_,
		_w196_,
		_w197_
	);
	LUT2 #(
		.INIT('h2)
	) name165 (
		_w188_,
		_w196_,
		_w198_
	);
	LUT2 #(
		.INIT('h1)
	) name166 (
		_w197_,
		_w198_,
		_w199_
	);
	LUT2 #(
		.INIT('h4)
	) name167 (
		_w187_,
		_w199_,
		_w200_
	);
	LUT2 #(
		.INIT('h2)
	) name168 (
		_w187_,
		_w199_,
		_w201_
	);
	LUT2 #(
		.INIT('h1)
	) name169 (
		_w200_,
		_w201_,
		_w202_
	);
	LUT2 #(
		.INIT('h4)
	) name170 (
		_w186_,
		_w202_,
		_w203_
	);
	LUT2 #(
		.INIT('h2)
	) name171 (
		_w186_,
		_w202_,
		_w204_
	);
	LUT2 #(
		.INIT('h1)
	) name172 (
		_w203_,
		_w204_,
		_w205_
	);
	LUT2 #(
		.INIT('h4)
	) name173 (
		_w185_,
		_w205_,
		_w206_
	);
	LUT2 #(
		.INIT('h2)
	) name174 (
		_w185_,
		_w205_,
		_w207_
	);
	LUT2 #(
		.INIT('h1)
	) name175 (
		_w206_,
		_w207_,
		_w208_
	);
	LUT2 #(
		.INIT('h4)
	) name176 (
		_w184_,
		_w208_,
		_w209_
	);
	LUT2 #(
		.INIT('h2)
	) name177 (
		_w184_,
		_w208_,
		_w210_
	);
	LUT2 #(
		.INIT('h1)
	) name178 (
		_w209_,
		_w210_,
		_w211_
	);
	LUT2 #(
		.INIT('h4)
	) name179 (
		_w183_,
		_w211_,
		_w212_
	);
	LUT2 #(
		.INIT('h2)
	) name180 (
		_w183_,
		_w211_,
		_w213_
	);
	LUT2 #(
		.INIT('h1)
	) name181 (
		_w212_,
		_w213_,
		_w214_
	);
	LUT2 #(
		.INIT('h4)
	) name182 (
		_w182_,
		_w214_,
		_w215_
	);
	LUT2 #(
		.INIT('h2)
	) name183 (
		_w182_,
		_w214_,
		_w216_
	);
	LUT2 #(
		.INIT('h1)
	) name184 (
		_w215_,
		_w216_,
		_w217_
	);
	LUT2 #(
		.INIT('h4)
	) name185 (
		_w181_,
		_w217_,
		_w218_
	);
	LUT2 #(
		.INIT('h2)
	) name186 (
		_w181_,
		_w217_,
		_w219_
	);
	LUT2 #(
		.INIT('h1)
	) name187 (
		_w218_,
		_w219_,
		_w220_
	);
	LUT2 #(
		.INIT('h4)
	) name188 (
		_w180_,
		_w220_,
		_w221_
	);
	LUT2 #(
		.INIT('h2)
	) name189 (
		_w180_,
		_w220_,
		_w222_
	);
	LUT2 #(
		.INIT('h1)
	) name190 (
		_w221_,
		_w222_,
		_w223_
	);
	LUT2 #(
		.INIT('h4)
	) name191 (
		_w179_,
		_w223_,
		_w224_
	);
	LUT2 #(
		.INIT('h2)
	) name192 (
		_w179_,
		_w223_,
		_w225_
	);
	LUT2 #(
		.INIT('h1)
	) name193 (
		_w224_,
		_w225_,
		_w226_
	);
	LUT2 #(
		.INIT('h4)
	) name194 (
		_w178_,
		_w226_,
		_w227_
	);
	LUT2 #(
		.INIT('h2)
	) name195 (
		_w178_,
		_w226_,
		_w228_
	);
	LUT2 #(
		.INIT('h1)
	) name196 (
		_w227_,
		_w228_,
		_w229_
	);
	LUT2 #(
		.INIT('h8)
	) name197 (
		\1GAT(0)_pad ,
		\409GAT(24)_pad ,
		_w230_
	);
	LUT2 #(
		.INIT('h1)
	) name198 (
		_w224_,
		_w227_,
		_w231_
	);
	LUT2 #(
		.INIT('h8)
	) name199 (
		\18GAT(1)_pad ,
		\392GAT(23)_pad ,
		_w232_
	);
	LUT2 #(
		.INIT('h1)
	) name200 (
		_w218_,
		_w221_,
		_w233_
	);
	LUT2 #(
		.INIT('h8)
	) name201 (
		\35GAT(2)_pad ,
		\375GAT(22)_pad ,
		_w234_
	);
	LUT2 #(
		.INIT('h1)
	) name202 (
		_w212_,
		_w215_,
		_w235_
	);
	LUT2 #(
		.INIT('h8)
	) name203 (
		\358GAT(21)_pad ,
		\52GAT(3)_pad ,
		_w236_
	);
	LUT2 #(
		.INIT('h1)
	) name204 (
		_w206_,
		_w209_,
		_w237_
	);
	LUT2 #(
		.INIT('h8)
	) name205 (
		\341GAT(20)_pad ,
		\69GAT(4)_pad ,
		_w238_
	);
	LUT2 #(
		.INIT('h1)
	) name206 (
		_w200_,
		_w203_,
		_w239_
	);
	LUT2 #(
		.INIT('h8)
	) name207 (
		\324GAT(19)_pad ,
		\86GAT(5)_pad ,
		_w240_
	);
	LUT2 #(
		.INIT('h1)
	) name208 (
		_w195_,
		_w197_,
		_w241_
	);
	LUT2 #(
		.INIT('h8)
	) name209 (
		\103GAT(6)_pad ,
		\307GAT(18)_pad ,
		_w242_
	);
	LUT2 #(
		.INIT('h4)
	) name210 (
		\137GAT(8)_pad ,
		_w144_,
		_w243_
	);
	LUT2 #(
		.INIT('h8)
	) name211 (
		\137GAT(8)_pad ,
		\273GAT(16)_pad ,
		_w244_
	);
	LUT2 #(
		.INIT('h8)
	) name212 (
		\120GAT(7)_pad ,
		\290GAT(17)_pad ,
		_w245_
	);
	LUT2 #(
		.INIT('h1)
	) name213 (
		_w244_,
		_w245_,
		_w246_
	);
	LUT2 #(
		.INIT('h4)
	) name214 (
		\103GAT(6)_pad ,
		_w244_,
		_w247_
	);
	LUT2 #(
		.INIT('h8)
	) name215 (
		_w245_,
		_w247_,
		_w248_
	);
	LUT2 #(
		.INIT('h1)
	) name216 (
		_w246_,
		_w248_,
		_w249_
	);
	LUT2 #(
		.INIT('h4)
	) name217 (
		_w243_,
		_w249_,
		_w250_
	);
	LUT2 #(
		.INIT('h4)
	) name218 (
		_w242_,
		_w250_,
		_w251_
	);
	LUT2 #(
		.INIT('h2)
	) name219 (
		_w242_,
		_w250_,
		_w252_
	);
	LUT2 #(
		.INIT('h1)
	) name220 (
		_w251_,
		_w252_,
		_w253_
	);
	LUT2 #(
		.INIT('h4)
	) name221 (
		_w241_,
		_w253_,
		_w254_
	);
	LUT2 #(
		.INIT('h2)
	) name222 (
		_w241_,
		_w253_,
		_w255_
	);
	LUT2 #(
		.INIT('h1)
	) name223 (
		_w254_,
		_w255_,
		_w256_
	);
	LUT2 #(
		.INIT('h4)
	) name224 (
		_w240_,
		_w256_,
		_w257_
	);
	LUT2 #(
		.INIT('h2)
	) name225 (
		_w240_,
		_w256_,
		_w258_
	);
	LUT2 #(
		.INIT('h1)
	) name226 (
		_w257_,
		_w258_,
		_w259_
	);
	LUT2 #(
		.INIT('h4)
	) name227 (
		_w239_,
		_w259_,
		_w260_
	);
	LUT2 #(
		.INIT('h2)
	) name228 (
		_w239_,
		_w259_,
		_w261_
	);
	LUT2 #(
		.INIT('h1)
	) name229 (
		_w260_,
		_w261_,
		_w262_
	);
	LUT2 #(
		.INIT('h4)
	) name230 (
		_w238_,
		_w262_,
		_w263_
	);
	LUT2 #(
		.INIT('h2)
	) name231 (
		_w238_,
		_w262_,
		_w264_
	);
	LUT2 #(
		.INIT('h1)
	) name232 (
		_w263_,
		_w264_,
		_w265_
	);
	LUT2 #(
		.INIT('h4)
	) name233 (
		_w237_,
		_w265_,
		_w266_
	);
	LUT2 #(
		.INIT('h2)
	) name234 (
		_w237_,
		_w265_,
		_w267_
	);
	LUT2 #(
		.INIT('h1)
	) name235 (
		_w266_,
		_w267_,
		_w268_
	);
	LUT2 #(
		.INIT('h4)
	) name236 (
		_w236_,
		_w268_,
		_w269_
	);
	LUT2 #(
		.INIT('h2)
	) name237 (
		_w236_,
		_w268_,
		_w270_
	);
	LUT2 #(
		.INIT('h1)
	) name238 (
		_w269_,
		_w270_,
		_w271_
	);
	LUT2 #(
		.INIT('h4)
	) name239 (
		_w235_,
		_w271_,
		_w272_
	);
	LUT2 #(
		.INIT('h2)
	) name240 (
		_w235_,
		_w271_,
		_w273_
	);
	LUT2 #(
		.INIT('h1)
	) name241 (
		_w272_,
		_w273_,
		_w274_
	);
	LUT2 #(
		.INIT('h4)
	) name242 (
		_w234_,
		_w274_,
		_w275_
	);
	LUT2 #(
		.INIT('h2)
	) name243 (
		_w234_,
		_w274_,
		_w276_
	);
	LUT2 #(
		.INIT('h1)
	) name244 (
		_w275_,
		_w276_,
		_w277_
	);
	LUT2 #(
		.INIT('h4)
	) name245 (
		_w233_,
		_w277_,
		_w278_
	);
	LUT2 #(
		.INIT('h2)
	) name246 (
		_w233_,
		_w277_,
		_w279_
	);
	LUT2 #(
		.INIT('h1)
	) name247 (
		_w278_,
		_w279_,
		_w280_
	);
	LUT2 #(
		.INIT('h4)
	) name248 (
		_w232_,
		_w280_,
		_w281_
	);
	LUT2 #(
		.INIT('h2)
	) name249 (
		_w232_,
		_w280_,
		_w282_
	);
	LUT2 #(
		.INIT('h1)
	) name250 (
		_w281_,
		_w282_,
		_w283_
	);
	LUT2 #(
		.INIT('h4)
	) name251 (
		_w231_,
		_w283_,
		_w284_
	);
	LUT2 #(
		.INIT('h2)
	) name252 (
		_w231_,
		_w283_,
		_w285_
	);
	LUT2 #(
		.INIT('h1)
	) name253 (
		_w284_,
		_w285_,
		_w286_
	);
	LUT2 #(
		.INIT('h4)
	) name254 (
		_w230_,
		_w286_,
		_w287_
	);
	LUT2 #(
		.INIT('h2)
	) name255 (
		_w230_,
		_w286_,
		_w288_
	);
	LUT2 #(
		.INIT('h1)
	) name256 (
		_w287_,
		_w288_,
		_w289_
	);
	LUT2 #(
		.INIT('h8)
	) name257 (
		\1GAT(0)_pad ,
		\426GAT(25)_pad ,
		_w290_
	);
	LUT2 #(
		.INIT('h1)
	) name258 (
		_w284_,
		_w287_,
		_w291_
	);
	LUT2 #(
		.INIT('h8)
	) name259 (
		\18GAT(1)_pad ,
		\409GAT(24)_pad ,
		_w292_
	);
	LUT2 #(
		.INIT('h1)
	) name260 (
		_w278_,
		_w281_,
		_w293_
	);
	LUT2 #(
		.INIT('h8)
	) name261 (
		\35GAT(2)_pad ,
		\392GAT(23)_pad ,
		_w294_
	);
	LUT2 #(
		.INIT('h1)
	) name262 (
		_w272_,
		_w275_,
		_w295_
	);
	LUT2 #(
		.INIT('h8)
	) name263 (
		\375GAT(22)_pad ,
		\52GAT(3)_pad ,
		_w296_
	);
	LUT2 #(
		.INIT('h1)
	) name264 (
		_w266_,
		_w269_,
		_w297_
	);
	LUT2 #(
		.INIT('h8)
	) name265 (
		\358GAT(21)_pad ,
		\69GAT(4)_pad ,
		_w298_
	);
	LUT2 #(
		.INIT('h1)
	) name266 (
		_w260_,
		_w263_,
		_w299_
	);
	LUT2 #(
		.INIT('h8)
	) name267 (
		\341GAT(20)_pad ,
		\86GAT(5)_pad ,
		_w300_
	);
	LUT2 #(
		.INIT('h1)
	) name268 (
		_w254_,
		_w257_,
		_w301_
	);
	LUT2 #(
		.INIT('h8)
	) name269 (
		\103GAT(6)_pad ,
		\324GAT(19)_pad ,
		_w302_
	);
	LUT2 #(
		.INIT('h2)
	) name270 (
		_w249_,
		_w251_,
		_w303_
	);
	LUT2 #(
		.INIT('h8)
	) name271 (
		\120GAT(7)_pad ,
		\307GAT(18)_pad ,
		_w304_
	);
	LUT2 #(
		.INIT('h4)
	) name272 (
		\154GAT(9)_pad ,
		_w191_,
		_w305_
	);
	LUT2 #(
		.INIT('h8)
	) name273 (
		\154GAT(9)_pad ,
		\273GAT(16)_pad ,
		_w306_
	);
	LUT2 #(
		.INIT('h8)
	) name274 (
		\137GAT(8)_pad ,
		\290GAT(17)_pad ,
		_w307_
	);
	LUT2 #(
		.INIT('h1)
	) name275 (
		_w306_,
		_w307_,
		_w308_
	);
	LUT2 #(
		.INIT('h4)
	) name276 (
		\120GAT(7)_pad ,
		_w306_,
		_w309_
	);
	LUT2 #(
		.INIT('h8)
	) name277 (
		_w307_,
		_w309_,
		_w310_
	);
	LUT2 #(
		.INIT('h1)
	) name278 (
		_w308_,
		_w310_,
		_w311_
	);
	LUT2 #(
		.INIT('h4)
	) name279 (
		_w305_,
		_w311_,
		_w312_
	);
	LUT2 #(
		.INIT('h4)
	) name280 (
		_w304_,
		_w312_,
		_w313_
	);
	LUT2 #(
		.INIT('h2)
	) name281 (
		_w304_,
		_w312_,
		_w314_
	);
	LUT2 #(
		.INIT('h1)
	) name282 (
		_w313_,
		_w314_,
		_w315_
	);
	LUT2 #(
		.INIT('h4)
	) name283 (
		_w303_,
		_w315_,
		_w316_
	);
	LUT2 #(
		.INIT('h2)
	) name284 (
		_w303_,
		_w315_,
		_w317_
	);
	LUT2 #(
		.INIT('h1)
	) name285 (
		_w316_,
		_w317_,
		_w318_
	);
	LUT2 #(
		.INIT('h4)
	) name286 (
		_w302_,
		_w318_,
		_w319_
	);
	LUT2 #(
		.INIT('h2)
	) name287 (
		_w302_,
		_w318_,
		_w320_
	);
	LUT2 #(
		.INIT('h1)
	) name288 (
		_w319_,
		_w320_,
		_w321_
	);
	LUT2 #(
		.INIT('h4)
	) name289 (
		_w301_,
		_w321_,
		_w322_
	);
	LUT2 #(
		.INIT('h2)
	) name290 (
		_w301_,
		_w321_,
		_w323_
	);
	LUT2 #(
		.INIT('h1)
	) name291 (
		_w322_,
		_w323_,
		_w324_
	);
	LUT2 #(
		.INIT('h4)
	) name292 (
		_w300_,
		_w324_,
		_w325_
	);
	LUT2 #(
		.INIT('h2)
	) name293 (
		_w300_,
		_w324_,
		_w326_
	);
	LUT2 #(
		.INIT('h1)
	) name294 (
		_w325_,
		_w326_,
		_w327_
	);
	LUT2 #(
		.INIT('h4)
	) name295 (
		_w299_,
		_w327_,
		_w328_
	);
	LUT2 #(
		.INIT('h2)
	) name296 (
		_w299_,
		_w327_,
		_w329_
	);
	LUT2 #(
		.INIT('h1)
	) name297 (
		_w328_,
		_w329_,
		_w330_
	);
	LUT2 #(
		.INIT('h4)
	) name298 (
		_w298_,
		_w330_,
		_w331_
	);
	LUT2 #(
		.INIT('h2)
	) name299 (
		_w298_,
		_w330_,
		_w332_
	);
	LUT2 #(
		.INIT('h1)
	) name300 (
		_w331_,
		_w332_,
		_w333_
	);
	LUT2 #(
		.INIT('h4)
	) name301 (
		_w297_,
		_w333_,
		_w334_
	);
	LUT2 #(
		.INIT('h2)
	) name302 (
		_w297_,
		_w333_,
		_w335_
	);
	LUT2 #(
		.INIT('h1)
	) name303 (
		_w334_,
		_w335_,
		_w336_
	);
	LUT2 #(
		.INIT('h4)
	) name304 (
		_w296_,
		_w336_,
		_w337_
	);
	LUT2 #(
		.INIT('h2)
	) name305 (
		_w296_,
		_w336_,
		_w338_
	);
	LUT2 #(
		.INIT('h1)
	) name306 (
		_w337_,
		_w338_,
		_w339_
	);
	LUT2 #(
		.INIT('h4)
	) name307 (
		_w295_,
		_w339_,
		_w340_
	);
	LUT2 #(
		.INIT('h2)
	) name308 (
		_w295_,
		_w339_,
		_w341_
	);
	LUT2 #(
		.INIT('h1)
	) name309 (
		_w340_,
		_w341_,
		_w342_
	);
	LUT2 #(
		.INIT('h4)
	) name310 (
		_w294_,
		_w342_,
		_w343_
	);
	LUT2 #(
		.INIT('h2)
	) name311 (
		_w294_,
		_w342_,
		_w344_
	);
	LUT2 #(
		.INIT('h1)
	) name312 (
		_w343_,
		_w344_,
		_w345_
	);
	LUT2 #(
		.INIT('h4)
	) name313 (
		_w293_,
		_w345_,
		_w346_
	);
	LUT2 #(
		.INIT('h2)
	) name314 (
		_w293_,
		_w345_,
		_w347_
	);
	LUT2 #(
		.INIT('h1)
	) name315 (
		_w346_,
		_w347_,
		_w348_
	);
	LUT2 #(
		.INIT('h4)
	) name316 (
		_w292_,
		_w348_,
		_w349_
	);
	LUT2 #(
		.INIT('h2)
	) name317 (
		_w292_,
		_w348_,
		_w350_
	);
	LUT2 #(
		.INIT('h1)
	) name318 (
		_w349_,
		_w350_,
		_w351_
	);
	LUT2 #(
		.INIT('h4)
	) name319 (
		_w291_,
		_w351_,
		_w352_
	);
	LUT2 #(
		.INIT('h2)
	) name320 (
		_w291_,
		_w351_,
		_w353_
	);
	LUT2 #(
		.INIT('h1)
	) name321 (
		_w352_,
		_w353_,
		_w354_
	);
	LUT2 #(
		.INIT('h4)
	) name322 (
		_w290_,
		_w354_,
		_w355_
	);
	LUT2 #(
		.INIT('h2)
	) name323 (
		_w290_,
		_w354_,
		_w356_
	);
	LUT2 #(
		.INIT('h1)
	) name324 (
		_w355_,
		_w356_,
		_w357_
	);
	LUT2 #(
		.INIT('h8)
	) name325 (
		\1GAT(0)_pad ,
		\443GAT(26)_pad ,
		_w358_
	);
	LUT2 #(
		.INIT('h1)
	) name326 (
		_w352_,
		_w355_,
		_w359_
	);
	LUT2 #(
		.INIT('h8)
	) name327 (
		\18GAT(1)_pad ,
		\426GAT(25)_pad ,
		_w360_
	);
	LUT2 #(
		.INIT('h1)
	) name328 (
		_w346_,
		_w349_,
		_w361_
	);
	LUT2 #(
		.INIT('h8)
	) name329 (
		\35GAT(2)_pad ,
		\409GAT(24)_pad ,
		_w362_
	);
	LUT2 #(
		.INIT('h1)
	) name330 (
		_w340_,
		_w343_,
		_w363_
	);
	LUT2 #(
		.INIT('h8)
	) name331 (
		\392GAT(23)_pad ,
		\52GAT(3)_pad ,
		_w364_
	);
	LUT2 #(
		.INIT('h1)
	) name332 (
		_w334_,
		_w337_,
		_w365_
	);
	LUT2 #(
		.INIT('h8)
	) name333 (
		\375GAT(22)_pad ,
		\69GAT(4)_pad ,
		_w366_
	);
	LUT2 #(
		.INIT('h1)
	) name334 (
		_w328_,
		_w331_,
		_w367_
	);
	LUT2 #(
		.INIT('h8)
	) name335 (
		\358GAT(21)_pad ,
		\86GAT(5)_pad ,
		_w368_
	);
	LUT2 #(
		.INIT('h1)
	) name336 (
		_w322_,
		_w325_,
		_w369_
	);
	LUT2 #(
		.INIT('h8)
	) name337 (
		\103GAT(6)_pad ,
		\341GAT(20)_pad ,
		_w370_
	);
	LUT2 #(
		.INIT('h1)
	) name338 (
		_w316_,
		_w319_,
		_w371_
	);
	LUT2 #(
		.INIT('h8)
	) name339 (
		\120GAT(7)_pad ,
		\324GAT(19)_pad ,
		_w372_
	);
	LUT2 #(
		.INIT('h2)
	) name340 (
		_w311_,
		_w313_,
		_w373_
	);
	LUT2 #(
		.INIT('h8)
	) name341 (
		\137GAT(8)_pad ,
		\307GAT(18)_pad ,
		_w374_
	);
	LUT2 #(
		.INIT('h4)
	) name342 (
		\171GAT(10)_pad ,
		_w244_,
		_w375_
	);
	LUT2 #(
		.INIT('h8)
	) name343 (
		\171GAT(10)_pad ,
		\273GAT(16)_pad ,
		_w376_
	);
	LUT2 #(
		.INIT('h8)
	) name344 (
		\154GAT(9)_pad ,
		\290GAT(17)_pad ,
		_w377_
	);
	LUT2 #(
		.INIT('h1)
	) name345 (
		_w376_,
		_w377_,
		_w378_
	);
	LUT2 #(
		.INIT('h4)
	) name346 (
		\137GAT(8)_pad ,
		_w376_,
		_w379_
	);
	LUT2 #(
		.INIT('h8)
	) name347 (
		_w377_,
		_w379_,
		_w380_
	);
	LUT2 #(
		.INIT('h1)
	) name348 (
		_w378_,
		_w380_,
		_w381_
	);
	LUT2 #(
		.INIT('h4)
	) name349 (
		_w375_,
		_w381_,
		_w382_
	);
	LUT2 #(
		.INIT('h4)
	) name350 (
		_w374_,
		_w382_,
		_w383_
	);
	LUT2 #(
		.INIT('h2)
	) name351 (
		_w374_,
		_w382_,
		_w384_
	);
	LUT2 #(
		.INIT('h1)
	) name352 (
		_w383_,
		_w384_,
		_w385_
	);
	LUT2 #(
		.INIT('h4)
	) name353 (
		_w373_,
		_w385_,
		_w386_
	);
	LUT2 #(
		.INIT('h2)
	) name354 (
		_w373_,
		_w385_,
		_w387_
	);
	LUT2 #(
		.INIT('h1)
	) name355 (
		_w386_,
		_w387_,
		_w388_
	);
	LUT2 #(
		.INIT('h4)
	) name356 (
		_w372_,
		_w388_,
		_w389_
	);
	LUT2 #(
		.INIT('h2)
	) name357 (
		_w372_,
		_w388_,
		_w390_
	);
	LUT2 #(
		.INIT('h1)
	) name358 (
		_w389_,
		_w390_,
		_w391_
	);
	LUT2 #(
		.INIT('h4)
	) name359 (
		_w371_,
		_w391_,
		_w392_
	);
	LUT2 #(
		.INIT('h2)
	) name360 (
		_w371_,
		_w391_,
		_w393_
	);
	LUT2 #(
		.INIT('h1)
	) name361 (
		_w392_,
		_w393_,
		_w394_
	);
	LUT2 #(
		.INIT('h4)
	) name362 (
		_w370_,
		_w394_,
		_w395_
	);
	LUT2 #(
		.INIT('h2)
	) name363 (
		_w370_,
		_w394_,
		_w396_
	);
	LUT2 #(
		.INIT('h1)
	) name364 (
		_w395_,
		_w396_,
		_w397_
	);
	LUT2 #(
		.INIT('h4)
	) name365 (
		_w369_,
		_w397_,
		_w398_
	);
	LUT2 #(
		.INIT('h2)
	) name366 (
		_w369_,
		_w397_,
		_w399_
	);
	LUT2 #(
		.INIT('h1)
	) name367 (
		_w398_,
		_w399_,
		_w400_
	);
	LUT2 #(
		.INIT('h4)
	) name368 (
		_w368_,
		_w400_,
		_w401_
	);
	LUT2 #(
		.INIT('h2)
	) name369 (
		_w368_,
		_w400_,
		_w402_
	);
	LUT2 #(
		.INIT('h1)
	) name370 (
		_w401_,
		_w402_,
		_w403_
	);
	LUT2 #(
		.INIT('h4)
	) name371 (
		_w367_,
		_w403_,
		_w404_
	);
	LUT2 #(
		.INIT('h2)
	) name372 (
		_w367_,
		_w403_,
		_w405_
	);
	LUT2 #(
		.INIT('h1)
	) name373 (
		_w404_,
		_w405_,
		_w406_
	);
	LUT2 #(
		.INIT('h4)
	) name374 (
		_w366_,
		_w406_,
		_w407_
	);
	LUT2 #(
		.INIT('h2)
	) name375 (
		_w366_,
		_w406_,
		_w408_
	);
	LUT2 #(
		.INIT('h1)
	) name376 (
		_w407_,
		_w408_,
		_w409_
	);
	LUT2 #(
		.INIT('h4)
	) name377 (
		_w365_,
		_w409_,
		_w410_
	);
	LUT2 #(
		.INIT('h2)
	) name378 (
		_w365_,
		_w409_,
		_w411_
	);
	LUT2 #(
		.INIT('h1)
	) name379 (
		_w410_,
		_w411_,
		_w412_
	);
	LUT2 #(
		.INIT('h4)
	) name380 (
		_w364_,
		_w412_,
		_w413_
	);
	LUT2 #(
		.INIT('h2)
	) name381 (
		_w364_,
		_w412_,
		_w414_
	);
	LUT2 #(
		.INIT('h1)
	) name382 (
		_w413_,
		_w414_,
		_w415_
	);
	LUT2 #(
		.INIT('h4)
	) name383 (
		_w363_,
		_w415_,
		_w416_
	);
	LUT2 #(
		.INIT('h2)
	) name384 (
		_w363_,
		_w415_,
		_w417_
	);
	LUT2 #(
		.INIT('h1)
	) name385 (
		_w416_,
		_w417_,
		_w418_
	);
	LUT2 #(
		.INIT('h4)
	) name386 (
		_w362_,
		_w418_,
		_w419_
	);
	LUT2 #(
		.INIT('h2)
	) name387 (
		_w362_,
		_w418_,
		_w420_
	);
	LUT2 #(
		.INIT('h1)
	) name388 (
		_w419_,
		_w420_,
		_w421_
	);
	LUT2 #(
		.INIT('h4)
	) name389 (
		_w361_,
		_w421_,
		_w422_
	);
	LUT2 #(
		.INIT('h2)
	) name390 (
		_w361_,
		_w421_,
		_w423_
	);
	LUT2 #(
		.INIT('h1)
	) name391 (
		_w422_,
		_w423_,
		_w424_
	);
	LUT2 #(
		.INIT('h4)
	) name392 (
		_w360_,
		_w424_,
		_w425_
	);
	LUT2 #(
		.INIT('h2)
	) name393 (
		_w360_,
		_w424_,
		_w426_
	);
	LUT2 #(
		.INIT('h1)
	) name394 (
		_w425_,
		_w426_,
		_w427_
	);
	LUT2 #(
		.INIT('h4)
	) name395 (
		_w359_,
		_w427_,
		_w428_
	);
	LUT2 #(
		.INIT('h2)
	) name396 (
		_w359_,
		_w427_,
		_w429_
	);
	LUT2 #(
		.INIT('h1)
	) name397 (
		_w428_,
		_w429_,
		_w430_
	);
	LUT2 #(
		.INIT('h4)
	) name398 (
		_w358_,
		_w430_,
		_w431_
	);
	LUT2 #(
		.INIT('h2)
	) name399 (
		_w358_,
		_w430_,
		_w432_
	);
	LUT2 #(
		.INIT('h1)
	) name400 (
		_w431_,
		_w432_,
		_w433_
	);
	LUT2 #(
		.INIT('h8)
	) name401 (
		\1GAT(0)_pad ,
		\460GAT(27)_pad ,
		_w434_
	);
	LUT2 #(
		.INIT('h1)
	) name402 (
		_w428_,
		_w431_,
		_w435_
	);
	LUT2 #(
		.INIT('h8)
	) name403 (
		\18GAT(1)_pad ,
		\443GAT(26)_pad ,
		_w436_
	);
	LUT2 #(
		.INIT('h1)
	) name404 (
		_w422_,
		_w425_,
		_w437_
	);
	LUT2 #(
		.INIT('h8)
	) name405 (
		\35GAT(2)_pad ,
		\426GAT(25)_pad ,
		_w438_
	);
	LUT2 #(
		.INIT('h1)
	) name406 (
		_w416_,
		_w419_,
		_w439_
	);
	LUT2 #(
		.INIT('h8)
	) name407 (
		\409GAT(24)_pad ,
		\52GAT(3)_pad ,
		_w440_
	);
	LUT2 #(
		.INIT('h1)
	) name408 (
		_w410_,
		_w413_,
		_w441_
	);
	LUT2 #(
		.INIT('h8)
	) name409 (
		\392GAT(23)_pad ,
		\69GAT(4)_pad ,
		_w442_
	);
	LUT2 #(
		.INIT('h1)
	) name410 (
		_w404_,
		_w407_,
		_w443_
	);
	LUT2 #(
		.INIT('h8)
	) name411 (
		\375GAT(22)_pad ,
		\86GAT(5)_pad ,
		_w444_
	);
	LUT2 #(
		.INIT('h1)
	) name412 (
		_w398_,
		_w401_,
		_w445_
	);
	LUT2 #(
		.INIT('h8)
	) name413 (
		\103GAT(6)_pad ,
		\358GAT(21)_pad ,
		_w446_
	);
	LUT2 #(
		.INIT('h1)
	) name414 (
		_w392_,
		_w395_,
		_w447_
	);
	LUT2 #(
		.INIT('h8)
	) name415 (
		\120GAT(7)_pad ,
		\341GAT(20)_pad ,
		_w448_
	);
	LUT2 #(
		.INIT('h1)
	) name416 (
		_w386_,
		_w389_,
		_w449_
	);
	LUT2 #(
		.INIT('h8)
	) name417 (
		\137GAT(8)_pad ,
		\324GAT(19)_pad ,
		_w450_
	);
	LUT2 #(
		.INIT('h2)
	) name418 (
		_w381_,
		_w383_,
		_w451_
	);
	LUT2 #(
		.INIT('h8)
	) name419 (
		\154GAT(9)_pad ,
		\307GAT(18)_pad ,
		_w452_
	);
	LUT2 #(
		.INIT('h4)
	) name420 (
		\188GAT(11)_pad ,
		_w306_,
		_w453_
	);
	LUT2 #(
		.INIT('h8)
	) name421 (
		\188GAT(11)_pad ,
		\273GAT(16)_pad ,
		_w454_
	);
	LUT2 #(
		.INIT('h8)
	) name422 (
		\171GAT(10)_pad ,
		\290GAT(17)_pad ,
		_w455_
	);
	LUT2 #(
		.INIT('h1)
	) name423 (
		_w454_,
		_w455_,
		_w456_
	);
	LUT2 #(
		.INIT('h4)
	) name424 (
		\154GAT(9)_pad ,
		_w454_,
		_w457_
	);
	LUT2 #(
		.INIT('h8)
	) name425 (
		_w455_,
		_w457_,
		_w458_
	);
	LUT2 #(
		.INIT('h1)
	) name426 (
		_w456_,
		_w458_,
		_w459_
	);
	LUT2 #(
		.INIT('h4)
	) name427 (
		_w453_,
		_w459_,
		_w460_
	);
	LUT2 #(
		.INIT('h4)
	) name428 (
		_w452_,
		_w460_,
		_w461_
	);
	LUT2 #(
		.INIT('h2)
	) name429 (
		_w452_,
		_w460_,
		_w462_
	);
	LUT2 #(
		.INIT('h1)
	) name430 (
		_w461_,
		_w462_,
		_w463_
	);
	LUT2 #(
		.INIT('h4)
	) name431 (
		_w451_,
		_w463_,
		_w464_
	);
	LUT2 #(
		.INIT('h2)
	) name432 (
		_w451_,
		_w463_,
		_w465_
	);
	LUT2 #(
		.INIT('h1)
	) name433 (
		_w464_,
		_w465_,
		_w466_
	);
	LUT2 #(
		.INIT('h4)
	) name434 (
		_w450_,
		_w466_,
		_w467_
	);
	LUT2 #(
		.INIT('h2)
	) name435 (
		_w450_,
		_w466_,
		_w468_
	);
	LUT2 #(
		.INIT('h1)
	) name436 (
		_w467_,
		_w468_,
		_w469_
	);
	LUT2 #(
		.INIT('h4)
	) name437 (
		_w449_,
		_w469_,
		_w470_
	);
	LUT2 #(
		.INIT('h2)
	) name438 (
		_w449_,
		_w469_,
		_w471_
	);
	LUT2 #(
		.INIT('h1)
	) name439 (
		_w470_,
		_w471_,
		_w472_
	);
	LUT2 #(
		.INIT('h4)
	) name440 (
		_w448_,
		_w472_,
		_w473_
	);
	LUT2 #(
		.INIT('h2)
	) name441 (
		_w448_,
		_w472_,
		_w474_
	);
	LUT2 #(
		.INIT('h1)
	) name442 (
		_w473_,
		_w474_,
		_w475_
	);
	LUT2 #(
		.INIT('h4)
	) name443 (
		_w447_,
		_w475_,
		_w476_
	);
	LUT2 #(
		.INIT('h2)
	) name444 (
		_w447_,
		_w475_,
		_w477_
	);
	LUT2 #(
		.INIT('h1)
	) name445 (
		_w476_,
		_w477_,
		_w478_
	);
	LUT2 #(
		.INIT('h4)
	) name446 (
		_w446_,
		_w478_,
		_w479_
	);
	LUT2 #(
		.INIT('h2)
	) name447 (
		_w446_,
		_w478_,
		_w480_
	);
	LUT2 #(
		.INIT('h1)
	) name448 (
		_w479_,
		_w480_,
		_w481_
	);
	LUT2 #(
		.INIT('h4)
	) name449 (
		_w445_,
		_w481_,
		_w482_
	);
	LUT2 #(
		.INIT('h2)
	) name450 (
		_w445_,
		_w481_,
		_w483_
	);
	LUT2 #(
		.INIT('h1)
	) name451 (
		_w482_,
		_w483_,
		_w484_
	);
	LUT2 #(
		.INIT('h4)
	) name452 (
		_w444_,
		_w484_,
		_w485_
	);
	LUT2 #(
		.INIT('h2)
	) name453 (
		_w444_,
		_w484_,
		_w486_
	);
	LUT2 #(
		.INIT('h1)
	) name454 (
		_w485_,
		_w486_,
		_w487_
	);
	LUT2 #(
		.INIT('h4)
	) name455 (
		_w443_,
		_w487_,
		_w488_
	);
	LUT2 #(
		.INIT('h2)
	) name456 (
		_w443_,
		_w487_,
		_w489_
	);
	LUT2 #(
		.INIT('h1)
	) name457 (
		_w488_,
		_w489_,
		_w490_
	);
	LUT2 #(
		.INIT('h4)
	) name458 (
		_w442_,
		_w490_,
		_w491_
	);
	LUT2 #(
		.INIT('h2)
	) name459 (
		_w442_,
		_w490_,
		_w492_
	);
	LUT2 #(
		.INIT('h1)
	) name460 (
		_w491_,
		_w492_,
		_w493_
	);
	LUT2 #(
		.INIT('h4)
	) name461 (
		_w441_,
		_w493_,
		_w494_
	);
	LUT2 #(
		.INIT('h2)
	) name462 (
		_w441_,
		_w493_,
		_w495_
	);
	LUT2 #(
		.INIT('h1)
	) name463 (
		_w494_,
		_w495_,
		_w496_
	);
	LUT2 #(
		.INIT('h4)
	) name464 (
		_w440_,
		_w496_,
		_w497_
	);
	LUT2 #(
		.INIT('h2)
	) name465 (
		_w440_,
		_w496_,
		_w498_
	);
	LUT2 #(
		.INIT('h1)
	) name466 (
		_w497_,
		_w498_,
		_w499_
	);
	LUT2 #(
		.INIT('h4)
	) name467 (
		_w439_,
		_w499_,
		_w500_
	);
	LUT2 #(
		.INIT('h2)
	) name468 (
		_w439_,
		_w499_,
		_w501_
	);
	LUT2 #(
		.INIT('h1)
	) name469 (
		_w500_,
		_w501_,
		_w502_
	);
	LUT2 #(
		.INIT('h4)
	) name470 (
		_w438_,
		_w502_,
		_w503_
	);
	LUT2 #(
		.INIT('h2)
	) name471 (
		_w438_,
		_w502_,
		_w504_
	);
	LUT2 #(
		.INIT('h1)
	) name472 (
		_w503_,
		_w504_,
		_w505_
	);
	LUT2 #(
		.INIT('h4)
	) name473 (
		_w437_,
		_w505_,
		_w506_
	);
	LUT2 #(
		.INIT('h2)
	) name474 (
		_w437_,
		_w505_,
		_w507_
	);
	LUT2 #(
		.INIT('h1)
	) name475 (
		_w506_,
		_w507_,
		_w508_
	);
	LUT2 #(
		.INIT('h4)
	) name476 (
		_w436_,
		_w508_,
		_w509_
	);
	LUT2 #(
		.INIT('h2)
	) name477 (
		_w436_,
		_w508_,
		_w510_
	);
	LUT2 #(
		.INIT('h1)
	) name478 (
		_w509_,
		_w510_,
		_w511_
	);
	LUT2 #(
		.INIT('h4)
	) name479 (
		_w435_,
		_w511_,
		_w512_
	);
	LUT2 #(
		.INIT('h2)
	) name480 (
		_w435_,
		_w511_,
		_w513_
	);
	LUT2 #(
		.INIT('h1)
	) name481 (
		_w512_,
		_w513_,
		_w514_
	);
	LUT2 #(
		.INIT('h4)
	) name482 (
		_w434_,
		_w514_,
		_w515_
	);
	LUT2 #(
		.INIT('h2)
	) name483 (
		_w434_,
		_w514_,
		_w516_
	);
	LUT2 #(
		.INIT('h1)
	) name484 (
		_w515_,
		_w516_,
		_w517_
	);
	LUT2 #(
		.INIT('h8)
	) name485 (
		\1GAT(0)_pad ,
		\477GAT(28)_pad ,
		_w518_
	);
	LUT2 #(
		.INIT('h1)
	) name486 (
		_w512_,
		_w515_,
		_w519_
	);
	LUT2 #(
		.INIT('h8)
	) name487 (
		\18GAT(1)_pad ,
		\460GAT(27)_pad ,
		_w520_
	);
	LUT2 #(
		.INIT('h1)
	) name488 (
		_w506_,
		_w509_,
		_w521_
	);
	LUT2 #(
		.INIT('h8)
	) name489 (
		\35GAT(2)_pad ,
		\443GAT(26)_pad ,
		_w522_
	);
	LUT2 #(
		.INIT('h1)
	) name490 (
		_w500_,
		_w503_,
		_w523_
	);
	LUT2 #(
		.INIT('h8)
	) name491 (
		\426GAT(25)_pad ,
		\52GAT(3)_pad ,
		_w524_
	);
	LUT2 #(
		.INIT('h1)
	) name492 (
		_w494_,
		_w497_,
		_w525_
	);
	LUT2 #(
		.INIT('h8)
	) name493 (
		\409GAT(24)_pad ,
		\69GAT(4)_pad ,
		_w526_
	);
	LUT2 #(
		.INIT('h1)
	) name494 (
		_w488_,
		_w491_,
		_w527_
	);
	LUT2 #(
		.INIT('h8)
	) name495 (
		\392GAT(23)_pad ,
		\86GAT(5)_pad ,
		_w528_
	);
	LUT2 #(
		.INIT('h1)
	) name496 (
		_w482_,
		_w485_,
		_w529_
	);
	LUT2 #(
		.INIT('h8)
	) name497 (
		\103GAT(6)_pad ,
		\375GAT(22)_pad ,
		_w530_
	);
	LUT2 #(
		.INIT('h1)
	) name498 (
		_w476_,
		_w479_,
		_w531_
	);
	LUT2 #(
		.INIT('h8)
	) name499 (
		\120GAT(7)_pad ,
		\358GAT(21)_pad ,
		_w532_
	);
	LUT2 #(
		.INIT('h1)
	) name500 (
		_w470_,
		_w473_,
		_w533_
	);
	LUT2 #(
		.INIT('h8)
	) name501 (
		\137GAT(8)_pad ,
		\341GAT(20)_pad ,
		_w534_
	);
	LUT2 #(
		.INIT('h1)
	) name502 (
		_w464_,
		_w467_,
		_w535_
	);
	LUT2 #(
		.INIT('h8)
	) name503 (
		\154GAT(9)_pad ,
		\324GAT(19)_pad ,
		_w536_
	);
	LUT2 #(
		.INIT('h2)
	) name504 (
		_w459_,
		_w461_,
		_w537_
	);
	LUT2 #(
		.INIT('h8)
	) name505 (
		\171GAT(10)_pad ,
		\307GAT(18)_pad ,
		_w538_
	);
	LUT2 #(
		.INIT('h4)
	) name506 (
		\205GAT(12)_pad ,
		_w376_,
		_w539_
	);
	LUT2 #(
		.INIT('h8)
	) name507 (
		\205GAT(12)_pad ,
		\273GAT(16)_pad ,
		_w540_
	);
	LUT2 #(
		.INIT('h8)
	) name508 (
		\188GAT(11)_pad ,
		\290GAT(17)_pad ,
		_w541_
	);
	LUT2 #(
		.INIT('h1)
	) name509 (
		_w540_,
		_w541_,
		_w542_
	);
	LUT2 #(
		.INIT('h4)
	) name510 (
		\171GAT(10)_pad ,
		_w540_,
		_w543_
	);
	LUT2 #(
		.INIT('h8)
	) name511 (
		_w541_,
		_w543_,
		_w544_
	);
	LUT2 #(
		.INIT('h1)
	) name512 (
		_w542_,
		_w544_,
		_w545_
	);
	LUT2 #(
		.INIT('h4)
	) name513 (
		_w539_,
		_w545_,
		_w546_
	);
	LUT2 #(
		.INIT('h4)
	) name514 (
		_w538_,
		_w546_,
		_w547_
	);
	LUT2 #(
		.INIT('h2)
	) name515 (
		_w538_,
		_w546_,
		_w548_
	);
	LUT2 #(
		.INIT('h1)
	) name516 (
		_w547_,
		_w548_,
		_w549_
	);
	LUT2 #(
		.INIT('h4)
	) name517 (
		_w537_,
		_w549_,
		_w550_
	);
	LUT2 #(
		.INIT('h2)
	) name518 (
		_w537_,
		_w549_,
		_w551_
	);
	LUT2 #(
		.INIT('h1)
	) name519 (
		_w550_,
		_w551_,
		_w552_
	);
	LUT2 #(
		.INIT('h4)
	) name520 (
		_w536_,
		_w552_,
		_w553_
	);
	LUT2 #(
		.INIT('h2)
	) name521 (
		_w536_,
		_w552_,
		_w554_
	);
	LUT2 #(
		.INIT('h1)
	) name522 (
		_w553_,
		_w554_,
		_w555_
	);
	LUT2 #(
		.INIT('h4)
	) name523 (
		_w535_,
		_w555_,
		_w556_
	);
	LUT2 #(
		.INIT('h2)
	) name524 (
		_w535_,
		_w555_,
		_w557_
	);
	LUT2 #(
		.INIT('h1)
	) name525 (
		_w556_,
		_w557_,
		_w558_
	);
	LUT2 #(
		.INIT('h4)
	) name526 (
		_w534_,
		_w558_,
		_w559_
	);
	LUT2 #(
		.INIT('h2)
	) name527 (
		_w534_,
		_w558_,
		_w560_
	);
	LUT2 #(
		.INIT('h1)
	) name528 (
		_w559_,
		_w560_,
		_w561_
	);
	LUT2 #(
		.INIT('h4)
	) name529 (
		_w533_,
		_w561_,
		_w562_
	);
	LUT2 #(
		.INIT('h2)
	) name530 (
		_w533_,
		_w561_,
		_w563_
	);
	LUT2 #(
		.INIT('h1)
	) name531 (
		_w562_,
		_w563_,
		_w564_
	);
	LUT2 #(
		.INIT('h4)
	) name532 (
		_w532_,
		_w564_,
		_w565_
	);
	LUT2 #(
		.INIT('h2)
	) name533 (
		_w532_,
		_w564_,
		_w566_
	);
	LUT2 #(
		.INIT('h1)
	) name534 (
		_w565_,
		_w566_,
		_w567_
	);
	LUT2 #(
		.INIT('h4)
	) name535 (
		_w531_,
		_w567_,
		_w568_
	);
	LUT2 #(
		.INIT('h2)
	) name536 (
		_w531_,
		_w567_,
		_w569_
	);
	LUT2 #(
		.INIT('h1)
	) name537 (
		_w568_,
		_w569_,
		_w570_
	);
	LUT2 #(
		.INIT('h4)
	) name538 (
		_w530_,
		_w570_,
		_w571_
	);
	LUT2 #(
		.INIT('h2)
	) name539 (
		_w530_,
		_w570_,
		_w572_
	);
	LUT2 #(
		.INIT('h1)
	) name540 (
		_w571_,
		_w572_,
		_w573_
	);
	LUT2 #(
		.INIT('h4)
	) name541 (
		_w529_,
		_w573_,
		_w574_
	);
	LUT2 #(
		.INIT('h2)
	) name542 (
		_w529_,
		_w573_,
		_w575_
	);
	LUT2 #(
		.INIT('h1)
	) name543 (
		_w574_,
		_w575_,
		_w576_
	);
	LUT2 #(
		.INIT('h4)
	) name544 (
		_w528_,
		_w576_,
		_w577_
	);
	LUT2 #(
		.INIT('h2)
	) name545 (
		_w528_,
		_w576_,
		_w578_
	);
	LUT2 #(
		.INIT('h1)
	) name546 (
		_w577_,
		_w578_,
		_w579_
	);
	LUT2 #(
		.INIT('h4)
	) name547 (
		_w527_,
		_w579_,
		_w580_
	);
	LUT2 #(
		.INIT('h2)
	) name548 (
		_w527_,
		_w579_,
		_w581_
	);
	LUT2 #(
		.INIT('h1)
	) name549 (
		_w580_,
		_w581_,
		_w582_
	);
	LUT2 #(
		.INIT('h4)
	) name550 (
		_w526_,
		_w582_,
		_w583_
	);
	LUT2 #(
		.INIT('h2)
	) name551 (
		_w526_,
		_w582_,
		_w584_
	);
	LUT2 #(
		.INIT('h1)
	) name552 (
		_w583_,
		_w584_,
		_w585_
	);
	LUT2 #(
		.INIT('h4)
	) name553 (
		_w525_,
		_w585_,
		_w586_
	);
	LUT2 #(
		.INIT('h2)
	) name554 (
		_w525_,
		_w585_,
		_w587_
	);
	LUT2 #(
		.INIT('h1)
	) name555 (
		_w586_,
		_w587_,
		_w588_
	);
	LUT2 #(
		.INIT('h4)
	) name556 (
		_w524_,
		_w588_,
		_w589_
	);
	LUT2 #(
		.INIT('h2)
	) name557 (
		_w524_,
		_w588_,
		_w590_
	);
	LUT2 #(
		.INIT('h1)
	) name558 (
		_w589_,
		_w590_,
		_w591_
	);
	LUT2 #(
		.INIT('h4)
	) name559 (
		_w523_,
		_w591_,
		_w592_
	);
	LUT2 #(
		.INIT('h2)
	) name560 (
		_w523_,
		_w591_,
		_w593_
	);
	LUT2 #(
		.INIT('h1)
	) name561 (
		_w592_,
		_w593_,
		_w594_
	);
	LUT2 #(
		.INIT('h4)
	) name562 (
		_w522_,
		_w594_,
		_w595_
	);
	LUT2 #(
		.INIT('h2)
	) name563 (
		_w522_,
		_w594_,
		_w596_
	);
	LUT2 #(
		.INIT('h1)
	) name564 (
		_w595_,
		_w596_,
		_w597_
	);
	LUT2 #(
		.INIT('h4)
	) name565 (
		_w521_,
		_w597_,
		_w598_
	);
	LUT2 #(
		.INIT('h2)
	) name566 (
		_w521_,
		_w597_,
		_w599_
	);
	LUT2 #(
		.INIT('h1)
	) name567 (
		_w598_,
		_w599_,
		_w600_
	);
	LUT2 #(
		.INIT('h4)
	) name568 (
		_w520_,
		_w600_,
		_w601_
	);
	LUT2 #(
		.INIT('h2)
	) name569 (
		_w520_,
		_w600_,
		_w602_
	);
	LUT2 #(
		.INIT('h1)
	) name570 (
		_w601_,
		_w602_,
		_w603_
	);
	LUT2 #(
		.INIT('h4)
	) name571 (
		_w519_,
		_w603_,
		_w604_
	);
	LUT2 #(
		.INIT('h2)
	) name572 (
		_w519_,
		_w603_,
		_w605_
	);
	LUT2 #(
		.INIT('h1)
	) name573 (
		_w604_,
		_w605_,
		_w606_
	);
	LUT2 #(
		.INIT('h4)
	) name574 (
		_w518_,
		_w606_,
		_w607_
	);
	LUT2 #(
		.INIT('h2)
	) name575 (
		_w518_,
		_w606_,
		_w608_
	);
	LUT2 #(
		.INIT('h1)
	) name576 (
		_w607_,
		_w608_,
		_w609_
	);
	LUT2 #(
		.INIT('h8)
	) name577 (
		\1GAT(0)_pad ,
		\273GAT(16)_pad ,
		_w610_
	);
	LUT2 #(
		.INIT('h8)
	) name578 (
		\1GAT(0)_pad ,
		\494GAT(29)_pad ,
		_w611_
	);
	LUT2 #(
		.INIT('h1)
	) name579 (
		_w604_,
		_w607_,
		_w612_
	);
	LUT2 #(
		.INIT('h8)
	) name580 (
		\18GAT(1)_pad ,
		\477GAT(28)_pad ,
		_w613_
	);
	LUT2 #(
		.INIT('h1)
	) name581 (
		_w598_,
		_w601_,
		_w614_
	);
	LUT2 #(
		.INIT('h8)
	) name582 (
		\35GAT(2)_pad ,
		\460GAT(27)_pad ,
		_w615_
	);
	LUT2 #(
		.INIT('h1)
	) name583 (
		_w592_,
		_w595_,
		_w616_
	);
	LUT2 #(
		.INIT('h8)
	) name584 (
		\443GAT(26)_pad ,
		\52GAT(3)_pad ,
		_w617_
	);
	LUT2 #(
		.INIT('h1)
	) name585 (
		_w586_,
		_w589_,
		_w618_
	);
	LUT2 #(
		.INIT('h8)
	) name586 (
		\426GAT(25)_pad ,
		\69GAT(4)_pad ,
		_w619_
	);
	LUT2 #(
		.INIT('h1)
	) name587 (
		_w580_,
		_w583_,
		_w620_
	);
	LUT2 #(
		.INIT('h8)
	) name588 (
		\409GAT(24)_pad ,
		\86GAT(5)_pad ,
		_w621_
	);
	LUT2 #(
		.INIT('h1)
	) name589 (
		_w574_,
		_w577_,
		_w622_
	);
	LUT2 #(
		.INIT('h8)
	) name590 (
		\103GAT(6)_pad ,
		\392GAT(23)_pad ,
		_w623_
	);
	LUT2 #(
		.INIT('h1)
	) name591 (
		_w568_,
		_w571_,
		_w624_
	);
	LUT2 #(
		.INIT('h8)
	) name592 (
		\120GAT(7)_pad ,
		\375GAT(22)_pad ,
		_w625_
	);
	LUT2 #(
		.INIT('h1)
	) name593 (
		_w562_,
		_w565_,
		_w626_
	);
	LUT2 #(
		.INIT('h8)
	) name594 (
		\137GAT(8)_pad ,
		\358GAT(21)_pad ,
		_w627_
	);
	LUT2 #(
		.INIT('h1)
	) name595 (
		_w556_,
		_w559_,
		_w628_
	);
	LUT2 #(
		.INIT('h8)
	) name596 (
		\154GAT(9)_pad ,
		\341GAT(20)_pad ,
		_w629_
	);
	LUT2 #(
		.INIT('h1)
	) name597 (
		_w550_,
		_w553_,
		_w630_
	);
	LUT2 #(
		.INIT('h8)
	) name598 (
		\171GAT(10)_pad ,
		\324GAT(19)_pad ,
		_w631_
	);
	LUT2 #(
		.INIT('h2)
	) name599 (
		_w545_,
		_w547_,
		_w632_
	);
	LUT2 #(
		.INIT('h8)
	) name600 (
		\188GAT(11)_pad ,
		\307GAT(18)_pad ,
		_w633_
	);
	LUT2 #(
		.INIT('h4)
	) name601 (
		\222GAT(13)_pad ,
		_w454_,
		_w634_
	);
	LUT2 #(
		.INIT('h8)
	) name602 (
		\222GAT(13)_pad ,
		\273GAT(16)_pad ,
		_w635_
	);
	LUT2 #(
		.INIT('h8)
	) name603 (
		\205GAT(12)_pad ,
		\290GAT(17)_pad ,
		_w636_
	);
	LUT2 #(
		.INIT('h1)
	) name604 (
		_w635_,
		_w636_,
		_w637_
	);
	LUT2 #(
		.INIT('h4)
	) name605 (
		\188GAT(11)_pad ,
		_w635_,
		_w638_
	);
	LUT2 #(
		.INIT('h8)
	) name606 (
		_w636_,
		_w638_,
		_w639_
	);
	LUT2 #(
		.INIT('h1)
	) name607 (
		_w637_,
		_w639_,
		_w640_
	);
	LUT2 #(
		.INIT('h4)
	) name608 (
		_w634_,
		_w640_,
		_w641_
	);
	LUT2 #(
		.INIT('h4)
	) name609 (
		_w633_,
		_w641_,
		_w642_
	);
	LUT2 #(
		.INIT('h2)
	) name610 (
		_w633_,
		_w641_,
		_w643_
	);
	LUT2 #(
		.INIT('h1)
	) name611 (
		_w642_,
		_w643_,
		_w644_
	);
	LUT2 #(
		.INIT('h4)
	) name612 (
		_w632_,
		_w644_,
		_w645_
	);
	LUT2 #(
		.INIT('h2)
	) name613 (
		_w632_,
		_w644_,
		_w646_
	);
	LUT2 #(
		.INIT('h1)
	) name614 (
		_w645_,
		_w646_,
		_w647_
	);
	LUT2 #(
		.INIT('h4)
	) name615 (
		_w631_,
		_w647_,
		_w648_
	);
	LUT2 #(
		.INIT('h2)
	) name616 (
		_w631_,
		_w647_,
		_w649_
	);
	LUT2 #(
		.INIT('h1)
	) name617 (
		_w648_,
		_w649_,
		_w650_
	);
	LUT2 #(
		.INIT('h4)
	) name618 (
		_w630_,
		_w650_,
		_w651_
	);
	LUT2 #(
		.INIT('h2)
	) name619 (
		_w630_,
		_w650_,
		_w652_
	);
	LUT2 #(
		.INIT('h1)
	) name620 (
		_w651_,
		_w652_,
		_w653_
	);
	LUT2 #(
		.INIT('h4)
	) name621 (
		_w629_,
		_w653_,
		_w654_
	);
	LUT2 #(
		.INIT('h2)
	) name622 (
		_w629_,
		_w653_,
		_w655_
	);
	LUT2 #(
		.INIT('h1)
	) name623 (
		_w654_,
		_w655_,
		_w656_
	);
	LUT2 #(
		.INIT('h4)
	) name624 (
		_w628_,
		_w656_,
		_w657_
	);
	LUT2 #(
		.INIT('h2)
	) name625 (
		_w628_,
		_w656_,
		_w658_
	);
	LUT2 #(
		.INIT('h1)
	) name626 (
		_w657_,
		_w658_,
		_w659_
	);
	LUT2 #(
		.INIT('h4)
	) name627 (
		_w627_,
		_w659_,
		_w660_
	);
	LUT2 #(
		.INIT('h2)
	) name628 (
		_w627_,
		_w659_,
		_w661_
	);
	LUT2 #(
		.INIT('h1)
	) name629 (
		_w660_,
		_w661_,
		_w662_
	);
	LUT2 #(
		.INIT('h4)
	) name630 (
		_w626_,
		_w662_,
		_w663_
	);
	LUT2 #(
		.INIT('h2)
	) name631 (
		_w626_,
		_w662_,
		_w664_
	);
	LUT2 #(
		.INIT('h1)
	) name632 (
		_w663_,
		_w664_,
		_w665_
	);
	LUT2 #(
		.INIT('h4)
	) name633 (
		_w625_,
		_w665_,
		_w666_
	);
	LUT2 #(
		.INIT('h2)
	) name634 (
		_w625_,
		_w665_,
		_w667_
	);
	LUT2 #(
		.INIT('h1)
	) name635 (
		_w666_,
		_w667_,
		_w668_
	);
	LUT2 #(
		.INIT('h4)
	) name636 (
		_w624_,
		_w668_,
		_w669_
	);
	LUT2 #(
		.INIT('h2)
	) name637 (
		_w624_,
		_w668_,
		_w670_
	);
	LUT2 #(
		.INIT('h1)
	) name638 (
		_w669_,
		_w670_,
		_w671_
	);
	LUT2 #(
		.INIT('h4)
	) name639 (
		_w623_,
		_w671_,
		_w672_
	);
	LUT2 #(
		.INIT('h2)
	) name640 (
		_w623_,
		_w671_,
		_w673_
	);
	LUT2 #(
		.INIT('h1)
	) name641 (
		_w672_,
		_w673_,
		_w674_
	);
	LUT2 #(
		.INIT('h4)
	) name642 (
		_w622_,
		_w674_,
		_w675_
	);
	LUT2 #(
		.INIT('h2)
	) name643 (
		_w622_,
		_w674_,
		_w676_
	);
	LUT2 #(
		.INIT('h1)
	) name644 (
		_w675_,
		_w676_,
		_w677_
	);
	LUT2 #(
		.INIT('h4)
	) name645 (
		_w621_,
		_w677_,
		_w678_
	);
	LUT2 #(
		.INIT('h2)
	) name646 (
		_w621_,
		_w677_,
		_w679_
	);
	LUT2 #(
		.INIT('h1)
	) name647 (
		_w678_,
		_w679_,
		_w680_
	);
	LUT2 #(
		.INIT('h4)
	) name648 (
		_w620_,
		_w680_,
		_w681_
	);
	LUT2 #(
		.INIT('h2)
	) name649 (
		_w620_,
		_w680_,
		_w682_
	);
	LUT2 #(
		.INIT('h1)
	) name650 (
		_w681_,
		_w682_,
		_w683_
	);
	LUT2 #(
		.INIT('h4)
	) name651 (
		_w619_,
		_w683_,
		_w684_
	);
	LUT2 #(
		.INIT('h2)
	) name652 (
		_w619_,
		_w683_,
		_w685_
	);
	LUT2 #(
		.INIT('h1)
	) name653 (
		_w684_,
		_w685_,
		_w686_
	);
	LUT2 #(
		.INIT('h4)
	) name654 (
		_w618_,
		_w686_,
		_w687_
	);
	LUT2 #(
		.INIT('h2)
	) name655 (
		_w618_,
		_w686_,
		_w688_
	);
	LUT2 #(
		.INIT('h1)
	) name656 (
		_w687_,
		_w688_,
		_w689_
	);
	LUT2 #(
		.INIT('h4)
	) name657 (
		_w617_,
		_w689_,
		_w690_
	);
	LUT2 #(
		.INIT('h2)
	) name658 (
		_w617_,
		_w689_,
		_w691_
	);
	LUT2 #(
		.INIT('h1)
	) name659 (
		_w690_,
		_w691_,
		_w692_
	);
	LUT2 #(
		.INIT('h4)
	) name660 (
		_w616_,
		_w692_,
		_w693_
	);
	LUT2 #(
		.INIT('h2)
	) name661 (
		_w616_,
		_w692_,
		_w694_
	);
	LUT2 #(
		.INIT('h1)
	) name662 (
		_w693_,
		_w694_,
		_w695_
	);
	LUT2 #(
		.INIT('h4)
	) name663 (
		_w615_,
		_w695_,
		_w696_
	);
	LUT2 #(
		.INIT('h2)
	) name664 (
		_w615_,
		_w695_,
		_w697_
	);
	LUT2 #(
		.INIT('h1)
	) name665 (
		_w696_,
		_w697_,
		_w698_
	);
	LUT2 #(
		.INIT('h4)
	) name666 (
		_w614_,
		_w698_,
		_w699_
	);
	LUT2 #(
		.INIT('h2)
	) name667 (
		_w614_,
		_w698_,
		_w700_
	);
	LUT2 #(
		.INIT('h1)
	) name668 (
		_w699_,
		_w700_,
		_w701_
	);
	LUT2 #(
		.INIT('h4)
	) name669 (
		_w613_,
		_w701_,
		_w702_
	);
	LUT2 #(
		.INIT('h2)
	) name670 (
		_w613_,
		_w701_,
		_w703_
	);
	LUT2 #(
		.INIT('h1)
	) name671 (
		_w702_,
		_w703_,
		_w704_
	);
	LUT2 #(
		.INIT('h4)
	) name672 (
		_w612_,
		_w704_,
		_w705_
	);
	LUT2 #(
		.INIT('h2)
	) name673 (
		_w612_,
		_w704_,
		_w706_
	);
	LUT2 #(
		.INIT('h1)
	) name674 (
		_w705_,
		_w706_,
		_w707_
	);
	LUT2 #(
		.INIT('h4)
	) name675 (
		_w611_,
		_w707_,
		_w708_
	);
	LUT2 #(
		.INIT('h2)
	) name676 (
		_w611_,
		_w707_,
		_w709_
	);
	LUT2 #(
		.INIT('h1)
	) name677 (
		_w708_,
		_w709_,
		_w710_
	);
	LUT2 #(
		.INIT('h8)
	) name678 (
		\1GAT(0)_pad ,
		\511GAT(30)_pad ,
		_w711_
	);
	LUT2 #(
		.INIT('h1)
	) name679 (
		_w705_,
		_w708_,
		_w712_
	);
	LUT2 #(
		.INIT('h8)
	) name680 (
		\18GAT(1)_pad ,
		\494GAT(29)_pad ,
		_w713_
	);
	LUT2 #(
		.INIT('h1)
	) name681 (
		_w699_,
		_w702_,
		_w714_
	);
	LUT2 #(
		.INIT('h8)
	) name682 (
		\35GAT(2)_pad ,
		\477GAT(28)_pad ,
		_w715_
	);
	LUT2 #(
		.INIT('h1)
	) name683 (
		_w693_,
		_w696_,
		_w716_
	);
	LUT2 #(
		.INIT('h8)
	) name684 (
		\460GAT(27)_pad ,
		\52GAT(3)_pad ,
		_w717_
	);
	LUT2 #(
		.INIT('h1)
	) name685 (
		_w687_,
		_w690_,
		_w718_
	);
	LUT2 #(
		.INIT('h8)
	) name686 (
		\443GAT(26)_pad ,
		\69GAT(4)_pad ,
		_w719_
	);
	LUT2 #(
		.INIT('h1)
	) name687 (
		_w681_,
		_w684_,
		_w720_
	);
	LUT2 #(
		.INIT('h8)
	) name688 (
		\426GAT(25)_pad ,
		\86GAT(5)_pad ,
		_w721_
	);
	LUT2 #(
		.INIT('h1)
	) name689 (
		_w675_,
		_w678_,
		_w722_
	);
	LUT2 #(
		.INIT('h8)
	) name690 (
		\103GAT(6)_pad ,
		\409GAT(24)_pad ,
		_w723_
	);
	LUT2 #(
		.INIT('h1)
	) name691 (
		_w669_,
		_w672_,
		_w724_
	);
	LUT2 #(
		.INIT('h8)
	) name692 (
		\120GAT(7)_pad ,
		\392GAT(23)_pad ,
		_w725_
	);
	LUT2 #(
		.INIT('h1)
	) name693 (
		_w663_,
		_w666_,
		_w726_
	);
	LUT2 #(
		.INIT('h8)
	) name694 (
		\137GAT(8)_pad ,
		\375GAT(22)_pad ,
		_w727_
	);
	LUT2 #(
		.INIT('h1)
	) name695 (
		_w657_,
		_w660_,
		_w728_
	);
	LUT2 #(
		.INIT('h8)
	) name696 (
		\154GAT(9)_pad ,
		\358GAT(21)_pad ,
		_w729_
	);
	LUT2 #(
		.INIT('h1)
	) name697 (
		_w651_,
		_w654_,
		_w730_
	);
	LUT2 #(
		.INIT('h8)
	) name698 (
		\171GAT(10)_pad ,
		\341GAT(20)_pad ,
		_w731_
	);
	LUT2 #(
		.INIT('h1)
	) name699 (
		_w645_,
		_w648_,
		_w732_
	);
	LUT2 #(
		.INIT('h8)
	) name700 (
		\188GAT(11)_pad ,
		\324GAT(19)_pad ,
		_w733_
	);
	LUT2 #(
		.INIT('h2)
	) name701 (
		_w640_,
		_w642_,
		_w734_
	);
	LUT2 #(
		.INIT('h8)
	) name702 (
		\205GAT(12)_pad ,
		\307GAT(18)_pad ,
		_w735_
	);
	LUT2 #(
		.INIT('h4)
	) name703 (
		\239GAT(14)_pad ,
		_w540_,
		_w736_
	);
	LUT2 #(
		.INIT('h8)
	) name704 (
		\239GAT(14)_pad ,
		\273GAT(16)_pad ,
		_w737_
	);
	LUT2 #(
		.INIT('h8)
	) name705 (
		\222GAT(13)_pad ,
		\290GAT(17)_pad ,
		_w738_
	);
	LUT2 #(
		.INIT('h1)
	) name706 (
		_w737_,
		_w738_,
		_w739_
	);
	LUT2 #(
		.INIT('h4)
	) name707 (
		\205GAT(12)_pad ,
		_w737_,
		_w740_
	);
	LUT2 #(
		.INIT('h8)
	) name708 (
		_w738_,
		_w740_,
		_w741_
	);
	LUT2 #(
		.INIT('h1)
	) name709 (
		_w739_,
		_w741_,
		_w742_
	);
	LUT2 #(
		.INIT('h4)
	) name710 (
		_w736_,
		_w742_,
		_w743_
	);
	LUT2 #(
		.INIT('h4)
	) name711 (
		_w735_,
		_w743_,
		_w744_
	);
	LUT2 #(
		.INIT('h2)
	) name712 (
		_w735_,
		_w743_,
		_w745_
	);
	LUT2 #(
		.INIT('h1)
	) name713 (
		_w744_,
		_w745_,
		_w746_
	);
	LUT2 #(
		.INIT('h4)
	) name714 (
		_w734_,
		_w746_,
		_w747_
	);
	LUT2 #(
		.INIT('h2)
	) name715 (
		_w734_,
		_w746_,
		_w748_
	);
	LUT2 #(
		.INIT('h1)
	) name716 (
		_w747_,
		_w748_,
		_w749_
	);
	LUT2 #(
		.INIT('h4)
	) name717 (
		_w733_,
		_w749_,
		_w750_
	);
	LUT2 #(
		.INIT('h2)
	) name718 (
		_w733_,
		_w749_,
		_w751_
	);
	LUT2 #(
		.INIT('h1)
	) name719 (
		_w750_,
		_w751_,
		_w752_
	);
	LUT2 #(
		.INIT('h4)
	) name720 (
		_w732_,
		_w752_,
		_w753_
	);
	LUT2 #(
		.INIT('h2)
	) name721 (
		_w732_,
		_w752_,
		_w754_
	);
	LUT2 #(
		.INIT('h1)
	) name722 (
		_w753_,
		_w754_,
		_w755_
	);
	LUT2 #(
		.INIT('h4)
	) name723 (
		_w731_,
		_w755_,
		_w756_
	);
	LUT2 #(
		.INIT('h2)
	) name724 (
		_w731_,
		_w755_,
		_w757_
	);
	LUT2 #(
		.INIT('h1)
	) name725 (
		_w756_,
		_w757_,
		_w758_
	);
	LUT2 #(
		.INIT('h4)
	) name726 (
		_w730_,
		_w758_,
		_w759_
	);
	LUT2 #(
		.INIT('h2)
	) name727 (
		_w730_,
		_w758_,
		_w760_
	);
	LUT2 #(
		.INIT('h1)
	) name728 (
		_w759_,
		_w760_,
		_w761_
	);
	LUT2 #(
		.INIT('h4)
	) name729 (
		_w729_,
		_w761_,
		_w762_
	);
	LUT2 #(
		.INIT('h2)
	) name730 (
		_w729_,
		_w761_,
		_w763_
	);
	LUT2 #(
		.INIT('h1)
	) name731 (
		_w762_,
		_w763_,
		_w764_
	);
	LUT2 #(
		.INIT('h4)
	) name732 (
		_w728_,
		_w764_,
		_w765_
	);
	LUT2 #(
		.INIT('h2)
	) name733 (
		_w728_,
		_w764_,
		_w766_
	);
	LUT2 #(
		.INIT('h1)
	) name734 (
		_w765_,
		_w766_,
		_w767_
	);
	LUT2 #(
		.INIT('h4)
	) name735 (
		_w727_,
		_w767_,
		_w768_
	);
	LUT2 #(
		.INIT('h2)
	) name736 (
		_w727_,
		_w767_,
		_w769_
	);
	LUT2 #(
		.INIT('h1)
	) name737 (
		_w768_,
		_w769_,
		_w770_
	);
	LUT2 #(
		.INIT('h4)
	) name738 (
		_w726_,
		_w770_,
		_w771_
	);
	LUT2 #(
		.INIT('h2)
	) name739 (
		_w726_,
		_w770_,
		_w772_
	);
	LUT2 #(
		.INIT('h1)
	) name740 (
		_w771_,
		_w772_,
		_w773_
	);
	LUT2 #(
		.INIT('h4)
	) name741 (
		_w725_,
		_w773_,
		_w774_
	);
	LUT2 #(
		.INIT('h2)
	) name742 (
		_w725_,
		_w773_,
		_w775_
	);
	LUT2 #(
		.INIT('h1)
	) name743 (
		_w774_,
		_w775_,
		_w776_
	);
	LUT2 #(
		.INIT('h4)
	) name744 (
		_w724_,
		_w776_,
		_w777_
	);
	LUT2 #(
		.INIT('h2)
	) name745 (
		_w724_,
		_w776_,
		_w778_
	);
	LUT2 #(
		.INIT('h1)
	) name746 (
		_w777_,
		_w778_,
		_w779_
	);
	LUT2 #(
		.INIT('h4)
	) name747 (
		_w723_,
		_w779_,
		_w780_
	);
	LUT2 #(
		.INIT('h2)
	) name748 (
		_w723_,
		_w779_,
		_w781_
	);
	LUT2 #(
		.INIT('h1)
	) name749 (
		_w780_,
		_w781_,
		_w782_
	);
	LUT2 #(
		.INIT('h4)
	) name750 (
		_w722_,
		_w782_,
		_w783_
	);
	LUT2 #(
		.INIT('h2)
	) name751 (
		_w722_,
		_w782_,
		_w784_
	);
	LUT2 #(
		.INIT('h1)
	) name752 (
		_w783_,
		_w784_,
		_w785_
	);
	LUT2 #(
		.INIT('h4)
	) name753 (
		_w721_,
		_w785_,
		_w786_
	);
	LUT2 #(
		.INIT('h2)
	) name754 (
		_w721_,
		_w785_,
		_w787_
	);
	LUT2 #(
		.INIT('h1)
	) name755 (
		_w786_,
		_w787_,
		_w788_
	);
	LUT2 #(
		.INIT('h4)
	) name756 (
		_w720_,
		_w788_,
		_w789_
	);
	LUT2 #(
		.INIT('h2)
	) name757 (
		_w720_,
		_w788_,
		_w790_
	);
	LUT2 #(
		.INIT('h1)
	) name758 (
		_w789_,
		_w790_,
		_w791_
	);
	LUT2 #(
		.INIT('h4)
	) name759 (
		_w719_,
		_w791_,
		_w792_
	);
	LUT2 #(
		.INIT('h2)
	) name760 (
		_w719_,
		_w791_,
		_w793_
	);
	LUT2 #(
		.INIT('h1)
	) name761 (
		_w792_,
		_w793_,
		_w794_
	);
	LUT2 #(
		.INIT('h4)
	) name762 (
		_w718_,
		_w794_,
		_w795_
	);
	LUT2 #(
		.INIT('h2)
	) name763 (
		_w718_,
		_w794_,
		_w796_
	);
	LUT2 #(
		.INIT('h1)
	) name764 (
		_w795_,
		_w796_,
		_w797_
	);
	LUT2 #(
		.INIT('h4)
	) name765 (
		_w717_,
		_w797_,
		_w798_
	);
	LUT2 #(
		.INIT('h2)
	) name766 (
		_w717_,
		_w797_,
		_w799_
	);
	LUT2 #(
		.INIT('h1)
	) name767 (
		_w798_,
		_w799_,
		_w800_
	);
	LUT2 #(
		.INIT('h4)
	) name768 (
		_w716_,
		_w800_,
		_w801_
	);
	LUT2 #(
		.INIT('h2)
	) name769 (
		_w716_,
		_w800_,
		_w802_
	);
	LUT2 #(
		.INIT('h1)
	) name770 (
		_w801_,
		_w802_,
		_w803_
	);
	LUT2 #(
		.INIT('h4)
	) name771 (
		_w715_,
		_w803_,
		_w804_
	);
	LUT2 #(
		.INIT('h2)
	) name772 (
		_w715_,
		_w803_,
		_w805_
	);
	LUT2 #(
		.INIT('h1)
	) name773 (
		_w804_,
		_w805_,
		_w806_
	);
	LUT2 #(
		.INIT('h4)
	) name774 (
		_w714_,
		_w806_,
		_w807_
	);
	LUT2 #(
		.INIT('h2)
	) name775 (
		_w714_,
		_w806_,
		_w808_
	);
	LUT2 #(
		.INIT('h1)
	) name776 (
		_w807_,
		_w808_,
		_w809_
	);
	LUT2 #(
		.INIT('h4)
	) name777 (
		_w713_,
		_w809_,
		_w810_
	);
	LUT2 #(
		.INIT('h2)
	) name778 (
		_w713_,
		_w809_,
		_w811_
	);
	LUT2 #(
		.INIT('h1)
	) name779 (
		_w810_,
		_w811_,
		_w812_
	);
	LUT2 #(
		.INIT('h4)
	) name780 (
		_w712_,
		_w812_,
		_w813_
	);
	LUT2 #(
		.INIT('h2)
	) name781 (
		_w712_,
		_w812_,
		_w814_
	);
	LUT2 #(
		.INIT('h1)
	) name782 (
		_w813_,
		_w814_,
		_w815_
	);
	LUT2 #(
		.INIT('h4)
	) name783 (
		_w711_,
		_w815_,
		_w816_
	);
	LUT2 #(
		.INIT('h2)
	) name784 (
		_w711_,
		_w815_,
		_w817_
	);
	LUT2 #(
		.INIT('h1)
	) name785 (
		_w816_,
		_w817_,
		_w818_
	);
	LUT2 #(
		.INIT('h8)
	) name786 (
		\1GAT(0)_pad ,
		\528GAT(31)_pad ,
		_w819_
	);
	LUT2 #(
		.INIT('h1)
	) name787 (
		_w813_,
		_w816_,
		_w820_
	);
	LUT2 #(
		.INIT('h8)
	) name788 (
		\18GAT(1)_pad ,
		\511GAT(30)_pad ,
		_w821_
	);
	LUT2 #(
		.INIT('h1)
	) name789 (
		_w807_,
		_w810_,
		_w822_
	);
	LUT2 #(
		.INIT('h8)
	) name790 (
		\35GAT(2)_pad ,
		\494GAT(29)_pad ,
		_w823_
	);
	LUT2 #(
		.INIT('h1)
	) name791 (
		_w801_,
		_w804_,
		_w824_
	);
	LUT2 #(
		.INIT('h8)
	) name792 (
		\477GAT(28)_pad ,
		\52GAT(3)_pad ,
		_w825_
	);
	LUT2 #(
		.INIT('h1)
	) name793 (
		_w795_,
		_w798_,
		_w826_
	);
	LUT2 #(
		.INIT('h8)
	) name794 (
		\460GAT(27)_pad ,
		\69GAT(4)_pad ,
		_w827_
	);
	LUT2 #(
		.INIT('h1)
	) name795 (
		_w789_,
		_w792_,
		_w828_
	);
	LUT2 #(
		.INIT('h8)
	) name796 (
		\443GAT(26)_pad ,
		\86GAT(5)_pad ,
		_w829_
	);
	LUT2 #(
		.INIT('h1)
	) name797 (
		_w783_,
		_w786_,
		_w830_
	);
	LUT2 #(
		.INIT('h8)
	) name798 (
		\103GAT(6)_pad ,
		\426GAT(25)_pad ,
		_w831_
	);
	LUT2 #(
		.INIT('h1)
	) name799 (
		_w777_,
		_w780_,
		_w832_
	);
	LUT2 #(
		.INIT('h8)
	) name800 (
		\120GAT(7)_pad ,
		\409GAT(24)_pad ,
		_w833_
	);
	LUT2 #(
		.INIT('h1)
	) name801 (
		_w771_,
		_w774_,
		_w834_
	);
	LUT2 #(
		.INIT('h8)
	) name802 (
		\137GAT(8)_pad ,
		\392GAT(23)_pad ,
		_w835_
	);
	LUT2 #(
		.INIT('h1)
	) name803 (
		_w765_,
		_w768_,
		_w836_
	);
	LUT2 #(
		.INIT('h8)
	) name804 (
		\154GAT(9)_pad ,
		\375GAT(22)_pad ,
		_w837_
	);
	LUT2 #(
		.INIT('h1)
	) name805 (
		_w759_,
		_w762_,
		_w838_
	);
	LUT2 #(
		.INIT('h8)
	) name806 (
		\171GAT(10)_pad ,
		\358GAT(21)_pad ,
		_w839_
	);
	LUT2 #(
		.INIT('h1)
	) name807 (
		_w753_,
		_w756_,
		_w840_
	);
	LUT2 #(
		.INIT('h8)
	) name808 (
		\188GAT(11)_pad ,
		\341GAT(20)_pad ,
		_w841_
	);
	LUT2 #(
		.INIT('h1)
	) name809 (
		_w747_,
		_w750_,
		_w842_
	);
	LUT2 #(
		.INIT('h8)
	) name810 (
		\205GAT(12)_pad ,
		\324GAT(19)_pad ,
		_w843_
	);
	LUT2 #(
		.INIT('h2)
	) name811 (
		_w742_,
		_w744_,
		_w844_
	);
	LUT2 #(
		.INIT('h8)
	) name812 (
		\222GAT(13)_pad ,
		\307GAT(18)_pad ,
		_w845_
	);
	LUT2 #(
		.INIT('h4)
	) name813 (
		\256GAT(15)_pad ,
		_w635_,
		_w846_
	);
	LUT2 #(
		.INIT('h8)
	) name814 (
		\256GAT(15)_pad ,
		\273GAT(16)_pad ,
		_w847_
	);
	LUT2 #(
		.INIT('h8)
	) name815 (
		\239GAT(14)_pad ,
		\290GAT(17)_pad ,
		_w848_
	);
	LUT2 #(
		.INIT('h1)
	) name816 (
		_w847_,
		_w848_,
		_w849_
	);
	LUT2 #(
		.INIT('h4)
	) name817 (
		\222GAT(13)_pad ,
		_w847_,
		_w850_
	);
	LUT2 #(
		.INIT('h8)
	) name818 (
		_w848_,
		_w850_,
		_w851_
	);
	LUT2 #(
		.INIT('h1)
	) name819 (
		_w849_,
		_w851_,
		_w852_
	);
	LUT2 #(
		.INIT('h4)
	) name820 (
		_w846_,
		_w852_,
		_w853_
	);
	LUT2 #(
		.INIT('h4)
	) name821 (
		_w845_,
		_w853_,
		_w854_
	);
	LUT2 #(
		.INIT('h2)
	) name822 (
		_w845_,
		_w853_,
		_w855_
	);
	LUT2 #(
		.INIT('h1)
	) name823 (
		_w854_,
		_w855_,
		_w856_
	);
	LUT2 #(
		.INIT('h4)
	) name824 (
		_w844_,
		_w856_,
		_w857_
	);
	LUT2 #(
		.INIT('h2)
	) name825 (
		_w844_,
		_w856_,
		_w858_
	);
	LUT2 #(
		.INIT('h1)
	) name826 (
		_w857_,
		_w858_,
		_w859_
	);
	LUT2 #(
		.INIT('h4)
	) name827 (
		_w843_,
		_w859_,
		_w860_
	);
	LUT2 #(
		.INIT('h2)
	) name828 (
		_w843_,
		_w859_,
		_w861_
	);
	LUT2 #(
		.INIT('h1)
	) name829 (
		_w860_,
		_w861_,
		_w862_
	);
	LUT2 #(
		.INIT('h4)
	) name830 (
		_w842_,
		_w862_,
		_w863_
	);
	LUT2 #(
		.INIT('h2)
	) name831 (
		_w842_,
		_w862_,
		_w864_
	);
	LUT2 #(
		.INIT('h1)
	) name832 (
		_w863_,
		_w864_,
		_w865_
	);
	LUT2 #(
		.INIT('h4)
	) name833 (
		_w841_,
		_w865_,
		_w866_
	);
	LUT2 #(
		.INIT('h2)
	) name834 (
		_w841_,
		_w865_,
		_w867_
	);
	LUT2 #(
		.INIT('h1)
	) name835 (
		_w866_,
		_w867_,
		_w868_
	);
	LUT2 #(
		.INIT('h4)
	) name836 (
		_w840_,
		_w868_,
		_w869_
	);
	LUT2 #(
		.INIT('h2)
	) name837 (
		_w840_,
		_w868_,
		_w870_
	);
	LUT2 #(
		.INIT('h1)
	) name838 (
		_w869_,
		_w870_,
		_w871_
	);
	LUT2 #(
		.INIT('h4)
	) name839 (
		_w839_,
		_w871_,
		_w872_
	);
	LUT2 #(
		.INIT('h2)
	) name840 (
		_w839_,
		_w871_,
		_w873_
	);
	LUT2 #(
		.INIT('h1)
	) name841 (
		_w872_,
		_w873_,
		_w874_
	);
	LUT2 #(
		.INIT('h4)
	) name842 (
		_w838_,
		_w874_,
		_w875_
	);
	LUT2 #(
		.INIT('h2)
	) name843 (
		_w838_,
		_w874_,
		_w876_
	);
	LUT2 #(
		.INIT('h1)
	) name844 (
		_w875_,
		_w876_,
		_w877_
	);
	LUT2 #(
		.INIT('h4)
	) name845 (
		_w837_,
		_w877_,
		_w878_
	);
	LUT2 #(
		.INIT('h2)
	) name846 (
		_w837_,
		_w877_,
		_w879_
	);
	LUT2 #(
		.INIT('h1)
	) name847 (
		_w878_,
		_w879_,
		_w880_
	);
	LUT2 #(
		.INIT('h4)
	) name848 (
		_w836_,
		_w880_,
		_w881_
	);
	LUT2 #(
		.INIT('h2)
	) name849 (
		_w836_,
		_w880_,
		_w882_
	);
	LUT2 #(
		.INIT('h1)
	) name850 (
		_w881_,
		_w882_,
		_w883_
	);
	LUT2 #(
		.INIT('h4)
	) name851 (
		_w835_,
		_w883_,
		_w884_
	);
	LUT2 #(
		.INIT('h2)
	) name852 (
		_w835_,
		_w883_,
		_w885_
	);
	LUT2 #(
		.INIT('h1)
	) name853 (
		_w884_,
		_w885_,
		_w886_
	);
	LUT2 #(
		.INIT('h4)
	) name854 (
		_w834_,
		_w886_,
		_w887_
	);
	LUT2 #(
		.INIT('h2)
	) name855 (
		_w834_,
		_w886_,
		_w888_
	);
	LUT2 #(
		.INIT('h1)
	) name856 (
		_w887_,
		_w888_,
		_w889_
	);
	LUT2 #(
		.INIT('h4)
	) name857 (
		_w833_,
		_w889_,
		_w890_
	);
	LUT2 #(
		.INIT('h2)
	) name858 (
		_w833_,
		_w889_,
		_w891_
	);
	LUT2 #(
		.INIT('h1)
	) name859 (
		_w890_,
		_w891_,
		_w892_
	);
	LUT2 #(
		.INIT('h4)
	) name860 (
		_w832_,
		_w892_,
		_w893_
	);
	LUT2 #(
		.INIT('h2)
	) name861 (
		_w832_,
		_w892_,
		_w894_
	);
	LUT2 #(
		.INIT('h1)
	) name862 (
		_w893_,
		_w894_,
		_w895_
	);
	LUT2 #(
		.INIT('h4)
	) name863 (
		_w831_,
		_w895_,
		_w896_
	);
	LUT2 #(
		.INIT('h2)
	) name864 (
		_w831_,
		_w895_,
		_w897_
	);
	LUT2 #(
		.INIT('h1)
	) name865 (
		_w896_,
		_w897_,
		_w898_
	);
	LUT2 #(
		.INIT('h4)
	) name866 (
		_w830_,
		_w898_,
		_w899_
	);
	LUT2 #(
		.INIT('h2)
	) name867 (
		_w830_,
		_w898_,
		_w900_
	);
	LUT2 #(
		.INIT('h1)
	) name868 (
		_w899_,
		_w900_,
		_w901_
	);
	LUT2 #(
		.INIT('h4)
	) name869 (
		_w829_,
		_w901_,
		_w902_
	);
	LUT2 #(
		.INIT('h2)
	) name870 (
		_w829_,
		_w901_,
		_w903_
	);
	LUT2 #(
		.INIT('h1)
	) name871 (
		_w902_,
		_w903_,
		_w904_
	);
	LUT2 #(
		.INIT('h4)
	) name872 (
		_w828_,
		_w904_,
		_w905_
	);
	LUT2 #(
		.INIT('h2)
	) name873 (
		_w828_,
		_w904_,
		_w906_
	);
	LUT2 #(
		.INIT('h1)
	) name874 (
		_w905_,
		_w906_,
		_w907_
	);
	LUT2 #(
		.INIT('h4)
	) name875 (
		_w827_,
		_w907_,
		_w908_
	);
	LUT2 #(
		.INIT('h2)
	) name876 (
		_w827_,
		_w907_,
		_w909_
	);
	LUT2 #(
		.INIT('h1)
	) name877 (
		_w908_,
		_w909_,
		_w910_
	);
	LUT2 #(
		.INIT('h4)
	) name878 (
		_w826_,
		_w910_,
		_w911_
	);
	LUT2 #(
		.INIT('h2)
	) name879 (
		_w826_,
		_w910_,
		_w912_
	);
	LUT2 #(
		.INIT('h1)
	) name880 (
		_w911_,
		_w912_,
		_w913_
	);
	LUT2 #(
		.INIT('h4)
	) name881 (
		_w825_,
		_w913_,
		_w914_
	);
	LUT2 #(
		.INIT('h2)
	) name882 (
		_w825_,
		_w913_,
		_w915_
	);
	LUT2 #(
		.INIT('h1)
	) name883 (
		_w914_,
		_w915_,
		_w916_
	);
	LUT2 #(
		.INIT('h4)
	) name884 (
		_w824_,
		_w916_,
		_w917_
	);
	LUT2 #(
		.INIT('h2)
	) name885 (
		_w824_,
		_w916_,
		_w918_
	);
	LUT2 #(
		.INIT('h1)
	) name886 (
		_w917_,
		_w918_,
		_w919_
	);
	LUT2 #(
		.INIT('h4)
	) name887 (
		_w823_,
		_w919_,
		_w920_
	);
	LUT2 #(
		.INIT('h2)
	) name888 (
		_w823_,
		_w919_,
		_w921_
	);
	LUT2 #(
		.INIT('h1)
	) name889 (
		_w920_,
		_w921_,
		_w922_
	);
	LUT2 #(
		.INIT('h4)
	) name890 (
		_w822_,
		_w922_,
		_w923_
	);
	LUT2 #(
		.INIT('h2)
	) name891 (
		_w822_,
		_w922_,
		_w924_
	);
	LUT2 #(
		.INIT('h1)
	) name892 (
		_w923_,
		_w924_,
		_w925_
	);
	LUT2 #(
		.INIT('h4)
	) name893 (
		_w821_,
		_w925_,
		_w926_
	);
	LUT2 #(
		.INIT('h2)
	) name894 (
		_w821_,
		_w925_,
		_w927_
	);
	LUT2 #(
		.INIT('h1)
	) name895 (
		_w926_,
		_w927_,
		_w928_
	);
	LUT2 #(
		.INIT('h4)
	) name896 (
		_w820_,
		_w928_,
		_w929_
	);
	LUT2 #(
		.INIT('h2)
	) name897 (
		_w820_,
		_w928_,
		_w930_
	);
	LUT2 #(
		.INIT('h1)
	) name898 (
		_w929_,
		_w930_,
		_w931_
	);
	LUT2 #(
		.INIT('h4)
	) name899 (
		_w819_,
		_w931_,
		_w932_
	);
	LUT2 #(
		.INIT('h2)
	) name900 (
		_w819_,
		_w931_,
		_w933_
	);
	LUT2 #(
		.INIT('h1)
	) name901 (
		_w932_,
		_w933_,
		_w934_
	);
	LUT2 #(
		.INIT('h1)
	) name902 (
		_w929_,
		_w932_,
		_w935_
	);
	LUT2 #(
		.INIT('h8)
	) name903 (
		\18GAT(1)_pad ,
		\528GAT(31)_pad ,
		_w936_
	);
	LUT2 #(
		.INIT('h1)
	) name904 (
		_w923_,
		_w926_,
		_w937_
	);
	LUT2 #(
		.INIT('h8)
	) name905 (
		\35GAT(2)_pad ,
		\511GAT(30)_pad ,
		_w938_
	);
	LUT2 #(
		.INIT('h1)
	) name906 (
		_w917_,
		_w920_,
		_w939_
	);
	LUT2 #(
		.INIT('h8)
	) name907 (
		\494GAT(29)_pad ,
		\52GAT(3)_pad ,
		_w940_
	);
	LUT2 #(
		.INIT('h1)
	) name908 (
		_w911_,
		_w914_,
		_w941_
	);
	LUT2 #(
		.INIT('h8)
	) name909 (
		\477GAT(28)_pad ,
		\69GAT(4)_pad ,
		_w942_
	);
	LUT2 #(
		.INIT('h1)
	) name910 (
		_w905_,
		_w908_,
		_w943_
	);
	LUT2 #(
		.INIT('h8)
	) name911 (
		\460GAT(27)_pad ,
		\86GAT(5)_pad ,
		_w944_
	);
	LUT2 #(
		.INIT('h1)
	) name912 (
		_w899_,
		_w902_,
		_w945_
	);
	LUT2 #(
		.INIT('h8)
	) name913 (
		\103GAT(6)_pad ,
		\443GAT(26)_pad ,
		_w946_
	);
	LUT2 #(
		.INIT('h1)
	) name914 (
		_w893_,
		_w896_,
		_w947_
	);
	LUT2 #(
		.INIT('h8)
	) name915 (
		\120GAT(7)_pad ,
		\426GAT(25)_pad ,
		_w948_
	);
	LUT2 #(
		.INIT('h1)
	) name916 (
		_w887_,
		_w890_,
		_w949_
	);
	LUT2 #(
		.INIT('h8)
	) name917 (
		\137GAT(8)_pad ,
		\409GAT(24)_pad ,
		_w950_
	);
	LUT2 #(
		.INIT('h1)
	) name918 (
		_w881_,
		_w884_,
		_w951_
	);
	LUT2 #(
		.INIT('h8)
	) name919 (
		\154GAT(9)_pad ,
		\392GAT(23)_pad ,
		_w952_
	);
	LUT2 #(
		.INIT('h1)
	) name920 (
		_w875_,
		_w878_,
		_w953_
	);
	LUT2 #(
		.INIT('h8)
	) name921 (
		\171GAT(10)_pad ,
		\375GAT(22)_pad ,
		_w954_
	);
	LUT2 #(
		.INIT('h1)
	) name922 (
		_w869_,
		_w872_,
		_w955_
	);
	LUT2 #(
		.INIT('h8)
	) name923 (
		\188GAT(11)_pad ,
		\358GAT(21)_pad ,
		_w956_
	);
	LUT2 #(
		.INIT('h1)
	) name924 (
		_w863_,
		_w866_,
		_w957_
	);
	LUT2 #(
		.INIT('h8)
	) name925 (
		\205GAT(12)_pad ,
		\341GAT(20)_pad ,
		_w958_
	);
	LUT2 #(
		.INIT('h1)
	) name926 (
		_w857_,
		_w860_,
		_w959_
	);
	LUT2 #(
		.INIT('h8)
	) name927 (
		\222GAT(13)_pad ,
		\324GAT(19)_pad ,
		_w960_
	);
	LUT2 #(
		.INIT('h2)
	) name928 (
		_w852_,
		_w854_,
		_w961_
	);
	LUT2 #(
		.INIT('h8)
	) name929 (
		\239GAT(14)_pad ,
		\307GAT(18)_pad ,
		_w962_
	);
	LUT2 #(
		.INIT('h8)
	) name930 (
		\256GAT(15)_pad ,
		\290GAT(17)_pad ,
		_w963_
	);
	LUT2 #(
		.INIT('h4)
	) name931 (
		_w737_,
		_w963_,
		_w964_
	);
	LUT2 #(
		.INIT('h4)
	) name932 (
		_w962_,
		_w964_,
		_w965_
	);
	LUT2 #(
		.INIT('h2)
	) name933 (
		_w962_,
		_w964_,
		_w966_
	);
	LUT2 #(
		.INIT('h1)
	) name934 (
		_w965_,
		_w966_,
		_w967_
	);
	LUT2 #(
		.INIT('h4)
	) name935 (
		_w961_,
		_w967_,
		_w968_
	);
	LUT2 #(
		.INIT('h2)
	) name936 (
		_w961_,
		_w967_,
		_w969_
	);
	LUT2 #(
		.INIT('h1)
	) name937 (
		_w968_,
		_w969_,
		_w970_
	);
	LUT2 #(
		.INIT('h4)
	) name938 (
		_w960_,
		_w970_,
		_w971_
	);
	LUT2 #(
		.INIT('h2)
	) name939 (
		_w960_,
		_w970_,
		_w972_
	);
	LUT2 #(
		.INIT('h1)
	) name940 (
		_w971_,
		_w972_,
		_w973_
	);
	LUT2 #(
		.INIT('h4)
	) name941 (
		_w959_,
		_w973_,
		_w974_
	);
	LUT2 #(
		.INIT('h2)
	) name942 (
		_w959_,
		_w973_,
		_w975_
	);
	LUT2 #(
		.INIT('h1)
	) name943 (
		_w974_,
		_w975_,
		_w976_
	);
	LUT2 #(
		.INIT('h4)
	) name944 (
		_w958_,
		_w976_,
		_w977_
	);
	LUT2 #(
		.INIT('h2)
	) name945 (
		_w958_,
		_w976_,
		_w978_
	);
	LUT2 #(
		.INIT('h1)
	) name946 (
		_w977_,
		_w978_,
		_w979_
	);
	LUT2 #(
		.INIT('h4)
	) name947 (
		_w957_,
		_w979_,
		_w980_
	);
	LUT2 #(
		.INIT('h2)
	) name948 (
		_w957_,
		_w979_,
		_w981_
	);
	LUT2 #(
		.INIT('h1)
	) name949 (
		_w980_,
		_w981_,
		_w982_
	);
	LUT2 #(
		.INIT('h4)
	) name950 (
		_w956_,
		_w982_,
		_w983_
	);
	LUT2 #(
		.INIT('h2)
	) name951 (
		_w956_,
		_w982_,
		_w984_
	);
	LUT2 #(
		.INIT('h1)
	) name952 (
		_w983_,
		_w984_,
		_w985_
	);
	LUT2 #(
		.INIT('h4)
	) name953 (
		_w955_,
		_w985_,
		_w986_
	);
	LUT2 #(
		.INIT('h2)
	) name954 (
		_w955_,
		_w985_,
		_w987_
	);
	LUT2 #(
		.INIT('h1)
	) name955 (
		_w986_,
		_w987_,
		_w988_
	);
	LUT2 #(
		.INIT('h4)
	) name956 (
		_w954_,
		_w988_,
		_w989_
	);
	LUT2 #(
		.INIT('h2)
	) name957 (
		_w954_,
		_w988_,
		_w990_
	);
	LUT2 #(
		.INIT('h1)
	) name958 (
		_w989_,
		_w990_,
		_w991_
	);
	LUT2 #(
		.INIT('h4)
	) name959 (
		_w953_,
		_w991_,
		_w992_
	);
	LUT2 #(
		.INIT('h2)
	) name960 (
		_w953_,
		_w991_,
		_w993_
	);
	LUT2 #(
		.INIT('h1)
	) name961 (
		_w992_,
		_w993_,
		_w994_
	);
	LUT2 #(
		.INIT('h4)
	) name962 (
		_w952_,
		_w994_,
		_w995_
	);
	LUT2 #(
		.INIT('h2)
	) name963 (
		_w952_,
		_w994_,
		_w996_
	);
	LUT2 #(
		.INIT('h1)
	) name964 (
		_w995_,
		_w996_,
		_w997_
	);
	LUT2 #(
		.INIT('h4)
	) name965 (
		_w951_,
		_w997_,
		_w998_
	);
	LUT2 #(
		.INIT('h2)
	) name966 (
		_w951_,
		_w997_,
		_w999_
	);
	LUT2 #(
		.INIT('h1)
	) name967 (
		_w998_,
		_w999_,
		_w1000_
	);
	LUT2 #(
		.INIT('h4)
	) name968 (
		_w950_,
		_w1000_,
		_w1001_
	);
	LUT2 #(
		.INIT('h2)
	) name969 (
		_w950_,
		_w1000_,
		_w1002_
	);
	LUT2 #(
		.INIT('h1)
	) name970 (
		_w1001_,
		_w1002_,
		_w1003_
	);
	LUT2 #(
		.INIT('h4)
	) name971 (
		_w949_,
		_w1003_,
		_w1004_
	);
	LUT2 #(
		.INIT('h2)
	) name972 (
		_w949_,
		_w1003_,
		_w1005_
	);
	LUT2 #(
		.INIT('h1)
	) name973 (
		_w1004_,
		_w1005_,
		_w1006_
	);
	LUT2 #(
		.INIT('h4)
	) name974 (
		_w948_,
		_w1006_,
		_w1007_
	);
	LUT2 #(
		.INIT('h2)
	) name975 (
		_w948_,
		_w1006_,
		_w1008_
	);
	LUT2 #(
		.INIT('h1)
	) name976 (
		_w1007_,
		_w1008_,
		_w1009_
	);
	LUT2 #(
		.INIT('h4)
	) name977 (
		_w947_,
		_w1009_,
		_w1010_
	);
	LUT2 #(
		.INIT('h2)
	) name978 (
		_w947_,
		_w1009_,
		_w1011_
	);
	LUT2 #(
		.INIT('h1)
	) name979 (
		_w1010_,
		_w1011_,
		_w1012_
	);
	LUT2 #(
		.INIT('h4)
	) name980 (
		_w946_,
		_w1012_,
		_w1013_
	);
	LUT2 #(
		.INIT('h2)
	) name981 (
		_w946_,
		_w1012_,
		_w1014_
	);
	LUT2 #(
		.INIT('h1)
	) name982 (
		_w1013_,
		_w1014_,
		_w1015_
	);
	LUT2 #(
		.INIT('h4)
	) name983 (
		_w945_,
		_w1015_,
		_w1016_
	);
	LUT2 #(
		.INIT('h2)
	) name984 (
		_w945_,
		_w1015_,
		_w1017_
	);
	LUT2 #(
		.INIT('h1)
	) name985 (
		_w1016_,
		_w1017_,
		_w1018_
	);
	LUT2 #(
		.INIT('h4)
	) name986 (
		_w944_,
		_w1018_,
		_w1019_
	);
	LUT2 #(
		.INIT('h2)
	) name987 (
		_w944_,
		_w1018_,
		_w1020_
	);
	LUT2 #(
		.INIT('h1)
	) name988 (
		_w1019_,
		_w1020_,
		_w1021_
	);
	LUT2 #(
		.INIT('h4)
	) name989 (
		_w943_,
		_w1021_,
		_w1022_
	);
	LUT2 #(
		.INIT('h2)
	) name990 (
		_w943_,
		_w1021_,
		_w1023_
	);
	LUT2 #(
		.INIT('h1)
	) name991 (
		_w1022_,
		_w1023_,
		_w1024_
	);
	LUT2 #(
		.INIT('h4)
	) name992 (
		_w942_,
		_w1024_,
		_w1025_
	);
	LUT2 #(
		.INIT('h2)
	) name993 (
		_w942_,
		_w1024_,
		_w1026_
	);
	LUT2 #(
		.INIT('h1)
	) name994 (
		_w1025_,
		_w1026_,
		_w1027_
	);
	LUT2 #(
		.INIT('h4)
	) name995 (
		_w941_,
		_w1027_,
		_w1028_
	);
	LUT2 #(
		.INIT('h2)
	) name996 (
		_w941_,
		_w1027_,
		_w1029_
	);
	LUT2 #(
		.INIT('h1)
	) name997 (
		_w1028_,
		_w1029_,
		_w1030_
	);
	LUT2 #(
		.INIT('h4)
	) name998 (
		_w940_,
		_w1030_,
		_w1031_
	);
	LUT2 #(
		.INIT('h2)
	) name999 (
		_w940_,
		_w1030_,
		_w1032_
	);
	LUT2 #(
		.INIT('h1)
	) name1000 (
		_w1031_,
		_w1032_,
		_w1033_
	);
	LUT2 #(
		.INIT('h4)
	) name1001 (
		_w939_,
		_w1033_,
		_w1034_
	);
	LUT2 #(
		.INIT('h2)
	) name1002 (
		_w939_,
		_w1033_,
		_w1035_
	);
	LUT2 #(
		.INIT('h1)
	) name1003 (
		_w1034_,
		_w1035_,
		_w1036_
	);
	LUT2 #(
		.INIT('h4)
	) name1004 (
		_w938_,
		_w1036_,
		_w1037_
	);
	LUT2 #(
		.INIT('h2)
	) name1005 (
		_w938_,
		_w1036_,
		_w1038_
	);
	LUT2 #(
		.INIT('h1)
	) name1006 (
		_w1037_,
		_w1038_,
		_w1039_
	);
	LUT2 #(
		.INIT('h4)
	) name1007 (
		_w937_,
		_w1039_,
		_w1040_
	);
	LUT2 #(
		.INIT('h2)
	) name1008 (
		_w937_,
		_w1039_,
		_w1041_
	);
	LUT2 #(
		.INIT('h1)
	) name1009 (
		_w1040_,
		_w1041_,
		_w1042_
	);
	LUT2 #(
		.INIT('h4)
	) name1010 (
		_w936_,
		_w1042_,
		_w1043_
	);
	LUT2 #(
		.INIT('h2)
	) name1011 (
		_w936_,
		_w1042_,
		_w1044_
	);
	LUT2 #(
		.INIT('h1)
	) name1012 (
		_w1043_,
		_w1044_,
		_w1045_
	);
	LUT2 #(
		.INIT('h4)
	) name1013 (
		_w935_,
		_w1045_,
		_w1046_
	);
	LUT2 #(
		.INIT('h2)
	) name1014 (
		_w935_,
		_w1045_,
		_w1047_
	);
	LUT2 #(
		.INIT('h1)
	) name1015 (
		_w1046_,
		_w1047_,
		_w1048_
	);
	LUT2 #(
		.INIT('h1)
	) name1016 (
		_w1040_,
		_w1043_,
		_w1049_
	);
	LUT2 #(
		.INIT('h8)
	) name1017 (
		\35GAT(2)_pad ,
		\528GAT(31)_pad ,
		_w1050_
	);
	LUT2 #(
		.INIT('h1)
	) name1018 (
		_w1034_,
		_w1037_,
		_w1051_
	);
	LUT2 #(
		.INIT('h8)
	) name1019 (
		\511GAT(30)_pad ,
		\52GAT(3)_pad ,
		_w1052_
	);
	LUT2 #(
		.INIT('h1)
	) name1020 (
		_w1028_,
		_w1031_,
		_w1053_
	);
	LUT2 #(
		.INIT('h8)
	) name1021 (
		\494GAT(29)_pad ,
		\69GAT(4)_pad ,
		_w1054_
	);
	LUT2 #(
		.INIT('h1)
	) name1022 (
		_w1022_,
		_w1025_,
		_w1055_
	);
	LUT2 #(
		.INIT('h8)
	) name1023 (
		\477GAT(28)_pad ,
		\86GAT(5)_pad ,
		_w1056_
	);
	LUT2 #(
		.INIT('h1)
	) name1024 (
		_w1016_,
		_w1019_,
		_w1057_
	);
	LUT2 #(
		.INIT('h8)
	) name1025 (
		\103GAT(6)_pad ,
		\460GAT(27)_pad ,
		_w1058_
	);
	LUT2 #(
		.INIT('h1)
	) name1026 (
		_w1010_,
		_w1013_,
		_w1059_
	);
	LUT2 #(
		.INIT('h8)
	) name1027 (
		\120GAT(7)_pad ,
		\443GAT(26)_pad ,
		_w1060_
	);
	LUT2 #(
		.INIT('h1)
	) name1028 (
		_w1004_,
		_w1007_,
		_w1061_
	);
	LUT2 #(
		.INIT('h8)
	) name1029 (
		\137GAT(8)_pad ,
		\426GAT(25)_pad ,
		_w1062_
	);
	LUT2 #(
		.INIT('h1)
	) name1030 (
		_w998_,
		_w1001_,
		_w1063_
	);
	LUT2 #(
		.INIT('h8)
	) name1031 (
		\154GAT(9)_pad ,
		\409GAT(24)_pad ,
		_w1064_
	);
	LUT2 #(
		.INIT('h1)
	) name1032 (
		_w992_,
		_w995_,
		_w1065_
	);
	LUT2 #(
		.INIT('h8)
	) name1033 (
		\171GAT(10)_pad ,
		\392GAT(23)_pad ,
		_w1066_
	);
	LUT2 #(
		.INIT('h1)
	) name1034 (
		_w986_,
		_w989_,
		_w1067_
	);
	LUT2 #(
		.INIT('h8)
	) name1035 (
		\188GAT(11)_pad ,
		\375GAT(22)_pad ,
		_w1068_
	);
	LUT2 #(
		.INIT('h1)
	) name1036 (
		_w980_,
		_w983_,
		_w1069_
	);
	LUT2 #(
		.INIT('h8)
	) name1037 (
		\205GAT(12)_pad ,
		\358GAT(21)_pad ,
		_w1070_
	);
	LUT2 #(
		.INIT('h1)
	) name1038 (
		_w974_,
		_w977_,
		_w1071_
	);
	LUT2 #(
		.INIT('h8)
	) name1039 (
		\222GAT(13)_pad ,
		\341GAT(20)_pad ,
		_w1072_
	);
	LUT2 #(
		.INIT('h1)
	) name1040 (
		_w968_,
		_w971_,
		_w1073_
	);
	LUT2 #(
		.INIT('h8)
	) name1041 (
		\239GAT(14)_pad ,
		\324GAT(19)_pad ,
		_w1074_
	);
	LUT2 #(
		.INIT('h8)
	) name1042 (
		\273GAT(16)_pad ,
		_w848_,
		_w1075_
	);
	LUT2 #(
		.INIT('h1)
	) name1043 (
		\307GAT(18)_pad ,
		_w1075_,
		_w1076_
	);
	LUT2 #(
		.INIT('h2)
	) name1044 (
		\256GAT(15)_pad ,
		_w1076_,
		_w1077_
	);
	LUT2 #(
		.INIT('h8)
	) name1045 (
		\290GAT(17)_pad ,
		_w962_,
		_w1078_
	);
	LUT2 #(
		.INIT('h2)
	) name1046 (
		_w1077_,
		_w1078_,
		_w1079_
	);
	LUT2 #(
		.INIT('h4)
	) name1047 (
		_w1074_,
		_w1079_,
		_w1080_
	);
	LUT2 #(
		.INIT('h2)
	) name1048 (
		_w1074_,
		_w1079_,
		_w1081_
	);
	LUT2 #(
		.INIT('h1)
	) name1049 (
		_w1080_,
		_w1081_,
		_w1082_
	);
	LUT2 #(
		.INIT('h4)
	) name1050 (
		_w1073_,
		_w1082_,
		_w1083_
	);
	LUT2 #(
		.INIT('h2)
	) name1051 (
		_w1073_,
		_w1082_,
		_w1084_
	);
	LUT2 #(
		.INIT('h1)
	) name1052 (
		_w1083_,
		_w1084_,
		_w1085_
	);
	LUT2 #(
		.INIT('h4)
	) name1053 (
		_w1072_,
		_w1085_,
		_w1086_
	);
	LUT2 #(
		.INIT('h2)
	) name1054 (
		_w1072_,
		_w1085_,
		_w1087_
	);
	LUT2 #(
		.INIT('h1)
	) name1055 (
		_w1086_,
		_w1087_,
		_w1088_
	);
	LUT2 #(
		.INIT('h4)
	) name1056 (
		_w1071_,
		_w1088_,
		_w1089_
	);
	LUT2 #(
		.INIT('h2)
	) name1057 (
		_w1071_,
		_w1088_,
		_w1090_
	);
	LUT2 #(
		.INIT('h1)
	) name1058 (
		_w1089_,
		_w1090_,
		_w1091_
	);
	LUT2 #(
		.INIT('h4)
	) name1059 (
		_w1070_,
		_w1091_,
		_w1092_
	);
	LUT2 #(
		.INIT('h2)
	) name1060 (
		_w1070_,
		_w1091_,
		_w1093_
	);
	LUT2 #(
		.INIT('h1)
	) name1061 (
		_w1092_,
		_w1093_,
		_w1094_
	);
	LUT2 #(
		.INIT('h4)
	) name1062 (
		_w1069_,
		_w1094_,
		_w1095_
	);
	LUT2 #(
		.INIT('h2)
	) name1063 (
		_w1069_,
		_w1094_,
		_w1096_
	);
	LUT2 #(
		.INIT('h1)
	) name1064 (
		_w1095_,
		_w1096_,
		_w1097_
	);
	LUT2 #(
		.INIT('h4)
	) name1065 (
		_w1068_,
		_w1097_,
		_w1098_
	);
	LUT2 #(
		.INIT('h2)
	) name1066 (
		_w1068_,
		_w1097_,
		_w1099_
	);
	LUT2 #(
		.INIT('h1)
	) name1067 (
		_w1098_,
		_w1099_,
		_w1100_
	);
	LUT2 #(
		.INIT('h4)
	) name1068 (
		_w1067_,
		_w1100_,
		_w1101_
	);
	LUT2 #(
		.INIT('h2)
	) name1069 (
		_w1067_,
		_w1100_,
		_w1102_
	);
	LUT2 #(
		.INIT('h1)
	) name1070 (
		_w1101_,
		_w1102_,
		_w1103_
	);
	LUT2 #(
		.INIT('h4)
	) name1071 (
		_w1066_,
		_w1103_,
		_w1104_
	);
	LUT2 #(
		.INIT('h2)
	) name1072 (
		_w1066_,
		_w1103_,
		_w1105_
	);
	LUT2 #(
		.INIT('h1)
	) name1073 (
		_w1104_,
		_w1105_,
		_w1106_
	);
	LUT2 #(
		.INIT('h4)
	) name1074 (
		_w1065_,
		_w1106_,
		_w1107_
	);
	LUT2 #(
		.INIT('h2)
	) name1075 (
		_w1065_,
		_w1106_,
		_w1108_
	);
	LUT2 #(
		.INIT('h1)
	) name1076 (
		_w1107_,
		_w1108_,
		_w1109_
	);
	LUT2 #(
		.INIT('h4)
	) name1077 (
		_w1064_,
		_w1109_,
		_w1110_
	);
	LUT2 #(
		.INIT('h2)
	) name1078 (
		_w1064_,
		_w1109_,
		_w1111_
	);
	LUT2 #(
		.INIT('h1)
	) name1079 (
		_w1110_,
		_w1111_,
		_w1112_
	);
	LUT2 #(
		.INIT('h4)
	) name1080 (
		_w1063_,
		_w1112_,
		_w1113_
	);
	LUT2 #(
		.INIT('h2)
	) name1081 (
		_w1063_,
		_w1112_,
		_w1114_
	);
	LUT2 #(
		.INIT('h1)
	) name1082 (
		_w1113_,
		_w1114_,
		_w1115_
	);
	LUT2 #(
		.INIT('h4)
	) name1083 (
		_w1062_,
		_w1115_,
		_w1116_
	);
	LUT2 #(
		.INIT('h2)
	) name1084 (
		_w1062_,
		_w1115_,
		_w1117_
	);
	LUT2 #(
		.INIT('h1)
	) name1085 (
		_w1116_,
		_w1117_,
		_w1118_
	);
	LUT2 #(
		.INIT('h4)
	) name1086 (
		_w1061_,
		_w1118_,
		_w1119_
	);
	LUT2 #(
		.INIT('h2)
	) name1087 (
		_w1061_,
		_w1118_,
		_w1120_
	);
	LUT2 #(
		.INIT('h1)
	) name1088 (
		_w1119_,
		_w1120_,
		_w1121_
	);
	LUT2 #(
		.INIT('h4)
	) name1089 (
		_w1060_,
		_w1121_,
		_w1122_
	);
	LUT2 #(
		.INIT('h2)
	) name1090 (
		_w1060_,
		_w1121_,
		_w1123_
	);
	LUT2 #(
		.INIT('h1)
	) name1091 (
		_w1122_,
		_w1123_,
		_w1124_
	);
	LUT2 #(
		.INIT('h4)
	) name1092 (
		_w1059_,
		_w1124_,
		_w1125_
	);
	LUT2 #(
		.INIT('h2)
	) name1093 (
		_w1059_,
		_w1124_,
		_w1126_
	);
	LUT2 #(
		.INIT('h1)
	) name1094 (
		_w1125_,
		_w1126_,
		_w1127_
	);
	LUT2 #(
		.INIT('h4)
	) name1095 (
		_w1058_,
		_w1127_,
		_w1128_
	);
	LUT2 #(
		.INIT('h2)
	) name1096 (
		_w1058_,
		_w1127_,
		_w1129_
	);
	LUT2 #(
		.INIT('h1)
	) name1097 (
		_w1128_,
		_w1129_,
		_w1130_
	);
	LUT2 #(
		.INIT('h4)
	) name1098 (
		_w1057_,
		_w1130_,
		_w1131_
	);
	LUT2 #(
		.INIT('h2)
	) name1099 (
		_w1057_,
		_w1130_,
		_w1132_
	);
	LUT2 #(
		.INIT('h1)
	) name1100 (
		_w1131_,
		_w1132_,
		_w1133_
	);
	LUT2 #(
		.INIT('h4)
	) name1101 (
		_w1056_,
		_w1133_,
		_w1134_
	);
	LUT2 #(
		.INIT('h2)
	) name1102 (
		_w1056_,
		_w1133_,
		_w1135_
	);
	LUT2 #(
		.INIT('h1)
	) name1103 (
		_w1134_,
		_w1135_,
		_w1136_
	);
	LUT2 #(
		.INIT('h4)
	) name1104 (
		_w1055_,
		_w1136_,
		_w1137_
	);
	LUT2 #(
		.INIT('h2)
	) name1105 (
		_w1055_,
		_w1136_,
		_w1138_
	);
	LUT2 #(
		.INIT('h1)
	) name1106 (
		_w1137_,
		_w1138_,
		_w1139_
	);
	LUT2 #(
		.INIT('h4)
	) name1107 (
		_w1054_,
		_w1139_,
		_w1140_
	);
	LUT2 #(
		.INIT('h2)
	) name1108 (
		_w1054_,
		_w1139_,
		_w1141_
	);
	LUT2 #(
		.INIT('h1)
	) name1109 (
		_w1140_,
		_w1141_,
		_w1142_
	);
	LUT2 #(
		.INIT('h4)
	) name1110 (
		_w1053_,
		_w1142_,
		_w1143_
	);
	LUT2 #(
		.INIT('h2)
	) name1111 (
		_w1053_,
		_w1142_,
		_w1144_
	);
	LUT2 #(
		.INIT('h1)
	) name1112 (
		_w1143_,
		_w1144_,
		_w1145_
	);
	LUT2 #(
		.INIT('h4)
	) name1113 (
		_w1052_,
		_w1145_,
		_w1146_
	);
	LUT2 #(
		.INIT('h2)
	) name1114 (
		_w1052_,
		_w1145_,
		_w1147_
	);
	LUT2 #(
		.INIT('h1)
	) name1115 (
		_w1146_,
		_w1147_,
		_w1148_
	);
	LUT2 #(
		.INIT('h4)
	) name1116 (
		_w1051_,
		_w1148_,
		_w1149_
	);
	LUT2 #(
		.INIT('h2)
	) name1117 (
		_w1051_,
		_w1148_,
		_w1150_
	);
	LUT2 #(
		.INIT('h1)
	) name1118 (
		_w1149_,
		_w1150_,
		_w1151_
	);
	LUT2 #(
		.INIT('h4)
	) name1119 (
		_w1050_,
		_w1151_,
		_w1152_
	);
	LUT2 #(
		.INIT('h2)
	) name1120 (
		_w1050_,
		_w1151_,
		_w1153_
	);
	LUT2 #(
		.INIT('h1)
	) name1121 (
		_w1152_,
		_w1153_,
		_w1154_
	);
	LUT2 #(
		.INIT('h4)
	) name1122 (
		_w1049_,
		_w1154_,
		_w1155_
	);
	LUT2 #(
		.INIT('h2)
	) name1123 (
		_w1049_,
		_w1154_,
		_w1156_
	);
	LUT2 #(
		.INIT('h1)
	) name1124 (
		_w1155_,
		_w1156_,
		_w1157_
	);
	LUT2 #(
		.INIT('h4)
	) name1125 (
		_w1047_,
		_w1157_,
		_w1158_
	);
	LUT2 #(
		.INIT('h2)
	) name1126 (
		_w1047_,
		_w1157_,
		_w1159_
	);
	LUT2 #(
		.INIT('h1)
	) name1127 (
		_w1158_,
		_w1159_,
		_w1160_
	);
	LUT2 #(
		.INIT('h1)
	) name1128 (
		_w1155_,
		_w1158_,
		_w1161_
	);
	LUT2 #(
		.INIT('h1)
	) name1129 (
		_w1149_,
		_w1152_,
		_w1162_
	);
	LUT2 #(
		.INIT('h8)
	) name1130 (
		\528GAT(31)_pad ,
		\52GAT(3)_pad ,
		_w1163_
	);
	LUT2 #(
		.INIT('h1)
	) name1131 (
		_w1143_,
		_w1146_,
		_w1164_
	);
	LUT2 #(
		.INIT('h8)
	) name1132 (
		\511GAT(30)_pad ,
		\69GAT(4)_pad ,
		_w1165_
	);
	LUT2 #(
		.INIT('h1)
	) name1133 (
		_w1137_,
		_w1140_,
		_w1166_
	);
	LUT2 #(
		.INIT('h8)
	) name1134 (
		\494GAT(29)_pad ,
		\86GAT(5)_pad ,
		_w1167_
	);
	LUT2 #(
		.INIT('h1)
	) name1135 (
		_w1131_,
		_w1134_,
		_w1168_
	);
	LUT2 #(
		.INIT('h8)
	) name1136 (
		\103GAT(6)_pad ,
		\477GAT(28)_pad ,
		_w1169_
	);
	LUT2 #(
		.INIT('h1)
	) name1137 (
		_w1125_,
		_w1128_,
		_w1170_
	);
	LUT2 #(
		.INIT('h8)
	) name1138 (
		\120GAT(7)_pad ,
		\460GAT(27)_pad ,
		_w1171_
	);
	LUT2 #(
		.INIT('h1)
	) name1139 (
		_w1119_,
		_w1122_,
		_w1172_
	);
	LUT2 #(
		.INIT('h8)
	) name1140 (
		\137GAT(8)_pad ,
		\443GAT(26)_pad ,
		_w1173_
	);
	LUT2 #(
		.INIT('h1)
	) name1141 (
		_w1113_,
		_w1116_,
		_w1174_
	);
	LUT2 #(
		.INIT('h8)
	) name1142 (
		\154GAT(9)_pad ,
		\426GAT(25)_pad ,
		_w1175_
	);
	LUT2 #(
		.INIT('h1)
	) name1143 (
		_w1107_,
		_w1110_,
		_w1176_
	);
	LUT2 #(
		.INIT('h8)
	) name1144 (
		\171GAT(10)_pad ,
		\409GAT(24)_pad ,
		_w1177_
	);
	LUT2 #(
		.INIT('h1)
	) name1145 (
		_w1101_,
		_w1104_,
		_w1178_
	);
	LUT2 #(
		.INIT('h8)
	) name1146 (
		\188GAT(11)_pad ,
		\392GAT(23)_pad ,
		_w1179_
	);
	LUT2 #(
		.INIT('h1)
	) name1147 (
		_w1095_,
		_w1098_,
		_w1180_
	);
	LUT2 #(
		.INIT('h8)
	) name1148 (
		\205GAT(12)_pad ,
		\375GAT(22)_pad ,
		_w1181_
	);
	LUT2 #(
		.INIT('h1)
	) name1149 (
		_w1089_,
		_w1092_,
		_w1182_
	);
	LUT2 #(
		.INIT('h8)
	) name1150 (
		\222GAT(13)_pad ,
		\358GAT(21)_pad ,
		_w1183_
	);
	LUT2 #(
		.INIT('h1)
	) name1151 (
		_w1083_,
		_w1086_,
		_w1184_
	);
	LUT2 #(
		.INIT('h8)
	) name1152 (
		\239GAT(14)_pad ,
		\341GAT(20)_pad ,
		_w1185_
	);
	LUT2 #(
		.INIT('h2)
	) name1153 (
		_w1077_,
		_w1080_,
		_w1186_
	);
	LUT2 #(
		.INIT('h8)
	) name1154 (
		\256GAT(15)_pad ,
		\324GAT(19)_pad ,
		_w1187_
	);
	LUT2 #(
		.INIT('h1)
	) name1155 (
		_w1186_,
		_w1187_,
		_w1188_
	);
	LUT2 #(
		.INIT('h8)
	) name1156 (
		\324GAT(19)_pad ,
		_w1186_,
		_w1189_
	);
	LUT2 #(
		.INIT('h1)
	) name1157 (
		_w1188_,
		_w1189_,
		_w1190_
	);
	LUT2 #(
		.INIT('h4)
	) name1158 (
		_w1185_,
		_w1190_,
		_w1191_
	);
	LUT2 #(
		.INIT('h2)
	) name1159 (
		_w1185_,
		_w1190_,
		_w1192_
	);
	LUT2 #(
		.INIT('h1)
	) name1160 (
		_w1191_,
		_w1192_,
		_w1193_
	);
	LUT2 #(
		.INIT('h4)
	) name1161 (
		_w1184_,
		_w1193_,
		_w1194_
	);
	LUT2 #(
		.INIT('h2)
	) name1162 (
		_w1184_,
		_w1193_,
		_w1195_
	);
	LUT2 #(
		.INIT('h1)
	) name1163 (
		_w1194_,
		_w1195_,
		_w1196_
	);
	LUT2 #(
		.INIT('h4)
	) name1164 (
		_w1183_,
		_w1196_,
		_w1197_
	);
	LUT2 #(
		.INIT('h2)
	) name1165 (
		_w1183_,
		_w1196_,
		_w1198_
	);
	LUT2 #(
		.INIT('h1)
	) name1166 (
		_w1197_,
		_w1198_,
		_w1199_
	);
	LUT2 #(
		.INIT('h4)
	) name1167 (
		_w1182_,
		_w1199_,
		_w1200_
	);
	LUT2 #(
		.INIT('h2)
	) name1168 (
		_w1182_,
		_w1199_,
		_w1201_
	);
	LUT2 #(
		.INIT('h1)
	) name1169 (
		_w1200_,
		_w1201_,
		_w1202_
	);
	LUT2 #(
		.INIT('h4)
	) name1170 (
		_w1181_,
		_w1202_,
		_w1203_
	);
	LUT2 #(
		.INIT('h2)
	) name1171 (
		_w1181_,
		_w1202_,
		_w1204_
	);
	LUT2 #(
		.INIT('h1)
	) name1172 (
		_w1203_,
		_w1204_,
		_w1205_
	);
	LUT2 #(
		.INIT('h4)
	) name1173 (
		_w1180_,
		_w1205_,
		_w1206_
	);
	LUT2 #(
		.INIT('h2)
	) name1174 (
		_w1180_,
		_w1205_,
		_w1207_
	);
	LUT2 #(
		.INIT('h1)
	) name1175 (
		_w1206_,
		_w1207_,
		_w1208_
	);
	LUT2 #(
		.INIT('h4)
	) name1176 (
		_w1179_,
		_w1208_,
		_w1209_
	);
	LUT2 #(
		.INIT('h2)
	) name1177 (
		_w1179_,
		_w1208_,
		_w1210_
	);
	LUT2 #(
		.INIT('h1)
	) name1178 (
		_w1209_,
		_w1210_,
		_w1211_
	);
	LUT2 #(
		.INIT('h4)
	) name1179 (
		_w1178_,
		_w1211_,
		_w1212_
	);
	LUT2 #(
		.INIT('h2)
	) name1180 (
		_w1178_,
		_w1211_,
		_w1213_
	);
	LUT2 #(
		.INIT('h1)
	) name1181 (
		_w1212_,
		_w1213_,
		_w1214_
	);
	LUT2 #(
		.INIT('h4)
	) name1182 (
		_w1177_,
		_w1214_,
		_w1215_
	);
	LUT2 #(
		.INIT('h2)
	) name1183 (
		_w1177_,
		_w1214_,
		_w1216_
	);
	LUT2 #(
		.INIT('h1)
	) name1184 (
		_w1215_,
		_w1216_,
		_w1217_
	);
	LUT2 #(
		.INIT('h4)
	) name1185 (
		_w1176_,
		_w1217_,
		_w1218_
	);
	LUT2 #(
		.INIT('h2)
	) name1186 (
		_w1176_,
		_w1217_,
		_w1219_
	);
	LUT2 #(
		.INIT('h1)
	) name1187 (
		_w1218_,
		_w1219_,
		_w1220_
	);
	LUT2 #(
		.INIT('h4)
	) name1188 (
		_w1175_,
		_w1220_,
		_w1221_
	);
	LUT2 #(
		.INIT('h2)
	) name1189 (
		_w1175_,
		_w1220_,
		_w1222_
	);
	LUT2 #(
		.INIT('h1)
	) name1190 (
		_w1221_,
		_w1222_,
		_w1223_
	);
	LUT2 #(
		.INIT('h4)
	) name1191 (
		_w1174_,
		_w1223_,
		_w1224_
	);
	LUT2 #(
		.INIT('h2)
	) name1192 (
		_w1174_,
		_w1223_,
		_w1225_
	);
	LUT2 #(
		.INIT('h1)
	) name1193 (
		_w1224_,
		_w1225_,
		_w1226_
	);
	LUT2 #(
		.INIT('h4)
	) name1194 (
		_w1173_,
		_w1226_,
		_w1227_
	);
	LUT2 #(
		.INIT('h2)
	) name1195 (
		_w1173_,
		_w1226_,
		_w1228_
	);
	LUT2 #(
		.INIT('h1)
	) name1196 (
		_w1227_,
		_w1228_,
		_w1229_
	);
	LUT2 #(
		.INIT('h4)
	) name1197 (
		_w1172_,
		_w1229_,
		_w1230_
	);
	LUT2 #(
		.INIT('h2)
	) name1198 (
		_w1172_,
		_w1229_,
		_w1231_
	);
	LUT2 #(
		.INIT('h1)
	) name1199 (
		_w1230_,
		_w1231_,
		_w1232_
	);
	LUT2 #(
		.INIT('h4)
	) name1200 (
		_w1171_,
		_w1232_,
		_w1233_
	);
	LUT2 #(
		.INIT('h2)
	) name1201 (
		_w1171_,
		_w1232_,
		_w1234_
	);
	LUT2 #(
		.INIT('h1)
	) name1202 (
		_w1233_,
		_w1234_,
		_w1235_
	);
	LUT2 #(
		.INIT('h4)
	) name1203 (
		_w1170_,
		_w1235_,
		_w1236_
	);
	LUT2 #(
		.INIT('h2)
	) name1204 (
		_w1170_,
		_w1235_,
		_w1237_
	);
	LUT2 #(
		.INIT('h1)
	) name1205 (
		_w1236_,
		_w1237_,
		_w1238_
	);
	LUT2 #(
		.INIT('h4)
	) name1206 (
		_w1169_,
		_w1238_,
		_w1239_
	);
	LUT2 #(
		.INIT('h2)
	) name1207 (
		_w1169_,
		_w1238_,
		_w1240_
	);
	LUT2 #(
		.INIT('h1)
	) name1208 (
		_w1239_,
		_w1240_,
		_w1241_
	);
	LUT2 #(
		.INIT('h4)
	) name1209 (
		_w1168_,
		_w1241_,
		_w1242_
	);
	LUT2 #(
		.INIT('h2)
	) name1210 (
		_w1168_,
		_w1241_,
		_w1243_
	);
	LUT2 #(
		.INIT('h1)
	) name1211 (
		_w1242_,
		_w1243_,
		_w1244_
	);
	LUT2 #(
		.INIT('h4)
	) name1212 (
		_w1167_,
		_w1244_,
		_w1245_
	);
	LUT2 #(
		.INIT('h2)
	) name1213 (
		_w1167_,
		_w1244_,
		_w1246_
	);
	LUT2 #(
		.INIT('h1)
	) name1214 (
		_w1245_,
		_w1246_,
		_w1247_
	);
	LUT2 #(
		.INIT('h4)
	) name1215 (
		_w1166_,
		_w1247_,
		_w1248_
	);
	LUT2 #(
		.INIT('h2)
	) name1216 (
		_w1166_,
		_w1247_,
		_w1249_
	);
	LUT2 #(
		.INIT('h1)
	) name1217 (
		_w1248_,
		_w1249_,
		_w1250_
	);
	LUT2 #(
		.INIT('h4)
	) name1218 (
		_w1165_,
		_w1250_,
		_w1251_
	);
	LUT2 #(
		.INIT('h2)
	) name1219 (
		_w1165_,
		_w1250_,
		_w1252_
	);
	LUT2 #(
		.INIT('h1)
	) name1220 (
		_w1251_,
		_w1252_,
		_w1253_
	);
	LUT2 #(
		.INIT('h4)
	) name1221 (
		_w1164_,
		_w1253_,
		_w1254_
	);
	LUT2 #(
		.INIT('h2)
	) name1222 (
		_w1164_,
		_w1253_,
		_w1255_
	);
	LUT2 #(
		.INIT('h1)
	) name1223 (
		_w1254_,
		_w1255_,
		_w1256_
	);
	LUT2 #(
		.INIT('h4)
	) name1224 (
		_w1163_,
		_w1256_,
		_w1257_
	);
	LUT2 #(
		.INIT('h2)
	) name1225 (
		_w1163_,
		_w1256_,
		_w1258_
	);
	LUT2 #(
		.INIT('h1)
	) name1226 (
		_w1257_,
		_w1258_,
		_w1259_
	);
	LUT2 #(
		.INIT('h4)
	) name1227 (
		_w1162_,
		_w1259_,
		_w1260_
	);
	LUT2 #(
		.INIT('h2)
	) name1228 (
		_w1162_,
		_w1259_,
		_w1261_
	);
	LUT2 #(
		.INIT('h1)
	) name1229 (
		_w1260_,
		_w1261_,
		_w1262_
	);
	LUT2 #(
		.INIT('h4)
	) name1230 (
		_w1161_,
		_w1262_,
		_w1263_
	);
	LUT2 #(
		.INIT('h2)
	) name1231 (
		_w1161_,
		_w1262_,
		_w1264_
	);
	LUT2 #(
		.INIT('h1)
	) name1232 (
		_w1263_,
		_w1264_,
		_w1265_
	);
	LUT2 #(
		.INIT('h1)
	) name1233 (
		_w1260_,
		_w1263_,
		_w1266_
	);
	LUT2 #(
		.INIT('h1)
	) name1234 (
		_w1254_,
		_w1257_,
		_w1267_
	);
	LUT2 #(
		.INIT('h8)
	) name1235 (
		\528GAT(31)_pad ,
		\69GAT(4)_pad ,
		_w1268_
	);
	LUT2 #(
		.INIT('h1)
	) name1236 (
		_w1248_,
		_w1251_,
		_w1269_
	);
	LUT2 #(
		.INIT('h8)
	) name1237 (
		\511GAT(30)_pad ,
		\86GAT(5)_pad ,
		_w1270_
	);
	LUT2 #(
		.INIT('h1)
	) name1238 (
		_w1242_,
		_w1245_,
		_w1271_
	);
	LUT2 #(
		.INIT('h8)
	) name1239 (
		\103GAT(6)_pad ,
		\494GAT(29)_pad ,
		_w1272_
	);
	LUT2 #(
		.INIT('h1)
	) name1240 (
		_w1236_,
		_w1239_,
		_w1273_
	);
	LUT2 #(
		.INIT('h8)
	) name1241 (
		\120GAT(7)_pad ,
		\477GAT(28)_pad ,
		_w1274_
	);
	LUT2 #(
		.INIT('h1)
	) name1242 (
		_w1230_,
		_w1233_,
		_w1275_
	);
	LUT2 #(
		.INIT('h8)
	) name1243 (
		\137GAT(8)_pad ,
		\460GAT(27)_pad ,
		_w1276_
	);
	LUT2 #(
		.INIT('h1)
	) name1244 (
		_w1224_,
		_w1227_,
		_w1277_
	);
	LUT2 #(
		.INIT('h8)
	) name1245 (
		\154GAT(9)_pad ,
		\443GAT(26)_pad ,
		_w1278_
	);
	LUT2 #(
		.INIT('h1)
	) name1246 (
		_w1218_,
		_w1221_,
		_w1279_
	);
	LUT2 #(
		.INIT('h8)
	) name1247 (
		\171GAT(10)_pad ,
		\426GAT(25)_pad ,
		_w1280_
	);
	LUT2 #(
		.INIT('h1)
	) name1248 (
		_w1212_,
		_w1215_,
		_w1281_
	);
	LUT2 #(
		.INIT('h8)
	) name1249 (
		\188GAT(11)_pad ,
		\409GAT(24)_pad ,
		_w1282_
	);
	LUT2 #(
		.INIT('h1)
	) name1250 (
		_w1206_,
		_w1209_,
		_w1283_
	);
	LUT2 #(
		.INIT('h8)
	) name1251 (
		\205GAT(12)_pad ,
		\392GAT(23)_pad ,
		_w1284_
	);
	LUT2 #(
		.INIT('h1)
	) name1252 (
		_w1200_,
		_w1203_,
		_w1285_
	);
	LUT2 #(
		.INIT('h8)
	) name1253 (
		\222GAT(13)_pad ,
		\375GAT(22)_pad ,
		_w1286_
	);
	LUT2 #(
		.INIT('h1)
	) name1254 (
		_w1194_,
		_w1197_,
		_w1287_
	);
	LUT2 #(
		.INIT('h8)
	) name1255 (
		\239GAT(14)_pad ,
		\358GAT(21)_pad ,
		_w1288_
	);
	LUT2 #(
		.INIT('h1)
	) name1256 (
		_w1188_,
		_w1191_,
		_w1289_
	);
	LUT2 #(
		.INIT('h8)
	) name1257 (
		\256GAT(15)_pad ,
		\341GAT(20)_pad ,
		_w1290_
	);
	LUT2 #(
		.INIT('h1)
	) name1258 (
		_w1289_,
		_w1290_,
		_w1291_
	);
	LUT2 #(
		.INIT('h8)
	) name1259 (
		_w1289_,
		_w1290_,
		_w1292_
	);
	LUT2 #(
		.INIT('h1)
	) name1260 (
		_w1291_,
		_w1292_,
		_w1293_
	);
	LUT2 #(
		.INIT('h4)
	) name1261 (
		_w1288_,
		_w1293_,
		_w1294_
	);
	LUT2 #(
		.INIT('h2)
	) name1262 (
		_w1288_,
		_w1293_,
		_w1295_
	);
	LUT2 #(
		.INIT('h1)
	) name1263 (
		_w1294_,
		_w1295_,
		_w1296_
	);
	LUT2 #(
		.INIT('h4)
	) name1264 (
		_w1287_,
		_w1296_,
		_w1297_
	);
	LUT2 #(
		.INIT('h2)
	) name1265 (
		_w1287_,
		_w1296_,
		_w1298_
	);
	LUT2 #(
		.INIT('h1)
	) name1266 (
		_w1297_,
		_w1298_,
		_w1299_
	);
	LUT2 #(
		.INIT('h4)
	) name1267 (
		_w1286_,
		_w1299_,
		_w1300_
	);
	LUT2 #(
		.INIT('h2)
	) name1268 (
		_w1286_,
		_w1299_,
		_w1301_
	);
	LUT2 #(
		.INIT('h1)
	) name1269 (
		_w1300_,
		_w1301_,
		_w1302_
	);
	LUT2 #(
		.INIT('h4)
	) name1270 (
		_w1285_,
		_w1302_,
		_w1303_
	);
	LUT2 #(
		.INIT('h2)
	) name1271 (
		_w1285_,
		_w1302_,
		_w1304_
	);
	LUT2 #(
		.INIT('h1)
	) name1272 (
		_w1303_,
		_w1304_,
		_w1305_
	);
	LUT2 #(
		.INIT('h4)
	) name1273 (
		_w1284_,
		_w1305_,
		_w1306_
	);
	LUT2 #(
		.INIT('h2)
	) name1274 (
		_w1284_,
		_w1305_,
		_w1307_
	);
	LUT2 #(
		.INIT('h1)
	) name1275 (
		_w1306_,
		_w1307_,
		_w1308_
	);
	LUT2 #(
		.INIT('h4)
	) name1276 (
		_w1283_,
		_w1308_,
		_w1309_
	);
	LUT2 #(
		.INIT('h2)
	) name1277 (
		_w1283_,
		_w1308_,
		_w1310_
	);
	LUT2 #(
		.INIT('h1)
	) name1278 (
		_w1309_,
		_w1310_,
		_w1311_
	);
	LUT2 #(
		.INIT('h4)
	) name1279 (
		_w1282_,
		_w1311_,
		_w1312_
	);
	LUT2 #(
		.INIT('h2)
	) name1280 (
		_w1282_,
		_w1311_,
		_w1313_
	);
	LUT2 #(
		.INIT('h1)
	) name1281 (
		_w1312_,
		_w1313_,
		_w1314_
	);
	LUT2 #(
		.INIT('h4)
	) name1282 (
		_w1281_,
		_w1314_,
		_w1315_
	);
	LUT2 #(
		.INIT('h2)
	) name1283 (
		_w1281_,
		_w1314_,
		_w1316_
	);
	LUT2 #(
		.INIT('h1)
	) name1284 (
		_w1315_,
		_w1316_,
		_w1317_
	);
	LUT2 #(
		.INIT('h4)
	) name1285 (
		_w1280_,
		_w1317_,
		_w1318_
	);
	LUT2 #(
		.INIT('h2)
	) name1286 (
		_w1280_,
		_w1317_,
		_w1319_
	);
	LUT2 #(
		.INIT('h1)
	) name1287 (
		_w1318_,
		_w1319_,
		_w1320_
	);
	LUT2 #(
		.INIT('h4)
	) name1288 (
		_w1279_,
		_w1320_,
		_w1321_
	);
	LUT2 #(
		.INIT('h2)
	) name1289 (
		_w1279_,
		_w1320_,
		_w1322_
	);
	LUT2 #(
		.INIT('h1)
	) name1290 (
		_w1321_,
		_w1322_,
		_w1323_
	);
	LUT2 #(
		.INIT('h4)
	) name1291 (
		_w1278_,
		_w1323_,
		_w1324_
	);
	LUT2 #(
		.INIT('h2)
	) name1292 (
		_w1278_,
		_w1323_,
		_w1325_
	);
	LUT2 #(
		.INIT('h1)
	) name1293 (
		_w1324_,
		_w1325_,
		_w1326_
	);
	LUT2 #(
		.INIT('h4)
	) name1294 (
		_w1277_,
		_w1326_,
		_w1327_
	);
	LUT2 #(
		.INIT('h2)
	) name1295 (
		_w1277_,
		_w1326_,
		_w1328_
	);
	LUT2 #(
		.INIT('h1)
	) name1296 (
		_w1327_,
		_w1328_,
		_w1329_
	);
	LUT2 #(
		.INIT('h4)
	) name1297 (
		_w1276_,
		_w1329_,
		_w1330_
	);
	LUT2 #(
		.INIT('h2)
	) name1298 (
		_w1276_,
		_w1329_,
		_w1331_
	);
	LUT2 #(
		.INIT('h1)
	) name1299 (
		_w1330_,
		_w1331_,
		_w1332_
	);
	LUT2 #(
		.INIT('h4)
	) name1300 (
		_w1275_,
		_w1332_,
		_w1333_
	);
	LUT2 #(
		.INIT('h2)
	) name1301 (
		_w1275_,
		_w1332_,
		_w1334_
	);
	LUT2 #(
		.INIT('h1)
	) name1302 (
		_w1333_,
		_w1334_,
		_w1335_
	);
	LUT2 #(
		.INIT('h4)
	) name1303 (
		_w1274_,
		_w1335_,
		_w1336_
	);
	LUT2 #(
		.INIT('h2)
	) name1304 (
		_w1274_,
		_w1335_,
		_w1337_
	);
	LUT2 #(
		.INIT('h1)
	) name1305 (
		_w1336_,
		_w1337_,
		_w1338_
	);
	LUT2 #(
		.INIT('h4)
	) name1306 (
		_w1273_,
		_w1338_,
		_w1339_
	);
	LUT2 #(
		.INIT('h2)
	) name1307 (
		_w1273_,
		_w1338_,
		_w1340_
	);
	LUT2 #(
		.INIT('h1)
	) name1308 (
		_w1339_,
		_w1340_,
		_w1341_
	);
	LUT2 #(
		.INIT('h4)
	) name1309 (
		_w1272_,
		_w1341_,
		_w1342_
	);
	LUT2 #(
		.INIT('h2)
	) name1310 (
		_w1272_,
		_w1341_,
		_w1343_
	);
	LUT2 #(
		.INIT('h1)
	) name1311 (
		_w1342_,
		_w1343_,
		_w1344_
	);
	LUT2 #(
		.INIT('h4)
	) name1312 (
		_w1271_,
		_w1344_,
		_w1345_
	);
	LUT2 #(
		.INIT('h2)
	) name1313 (
		_w1271_,
		_w1344_,
		_w1346_
	);
	LUT2 #(
		.INIT('h1)
	) name1314 (
		_w1345_,
		_w1346_,
		_w1347_
	);
	LUT2 #(
		.INIT('h4)
	) name1315 (
		_w1270_,
		_w1347_,
		_w1348_
	);
	LUT2 #(
		.INIT('h2)
	) name1316 (
		_w1270_,
		_w1347_,
		_w1349_
	);
	LUT2 #(
		.INIT('h1)
	) name1317 (
		_w1348_,
		_w1349_,
		_w1350_
	);
	LUT2 #(
		.INIT('h4)
	) name1318 (
		_w1269_,
		_w1350_,
		_w1351_
	);
	LUT2 #(
		.INIT('h2)
	) name1319 (
		_w1269_,
		_w1350_,
		_w1352_
	);
	LUT2 #(
		.INIT('h1)
	) name1320 (
		_w1351_,
		_w1352_,
		_w1353_
	);
	LUT2 #(
		.INIT('h4)
	) name1321 (
		_w1268_,
		_w1353_,
		_w1354_
	);
	LUT2 #(
		.INIT('h2)
	) name1322 (
		_w1268_,
		_w1353_,
		_w1355_
	);
	LUT2 #(
		.INIT('h1)
	) name1323 (
		_w1354_,
		_w1355_,
		_w1356_
	);
	LUT2 #(
		.INIT('h4)
	) name1324 (
		_w1267_,
		_w1356_,
		_w1357_
	);
	LUT2 #(
		.INIT('h2)
	) name1325 (
		_w1267_,
		_w1356_,
		_w1358_
	);
	LUT2 #(
		.INIT('h1)
	) name1326 (
		_w1357_,
		_w1358_,
		_w1359_
	);
	LUT2 #(
		.INIT('h4)
	) name1327 (
		_w1266_,
		_w1359_,
		_w1360_
	);
	LUT2 #(
		.INIT('h2)
	) name1328 (
		_w1266_,
		_w1359_,
		_w1361_
	);
	LUT2 #(
		.INIT('h1)
	) name1329 (
		_w1360_,
		_w1361_,
		_w1362_
	);
	LUT2 #(
		.INIT('h1)
	) name1330 (
		_w1357_,
		_w1360_,
		_w1363_
	);
	LUT2 #(
		.INIT('h1)
	) name1331 (
		_w1351_,
		_w1354_,
		_w1364_
	);
	LUT2 #(
		.INIT('h8)
	) name1332 (
		\528GAT(31)_pad ,
		\86GAT(5)_pad ,
		_w1365_
	);
	LUT2 #(
		.INIT('h1)
	) name1333 (
		_w1345_,
		_w1348_,
		_w1366_
	);
	LUT2 #(
		.INIT('h8)
	) name1334 (
		\103GAT(6)_pad ,
		\511GAT(30)_pad ,
		_w1367_
	);
	LUT2 #(
		.INIT('h1)
	) name1335 (
		_w1339_,
		_w1342_,
		_w1368_
	);
	LUT2 #(
		.INIT('h8)
	) name1336 (
		\120GAT(7)_pad ,
		\494GAT(29)_pad ,
		_w1369_
	);
	LUT2 #(
		.INIT('h1)
	) name1337 (
		_w1333_,
		_w1336_,
		_w1370_
	);
	LUT2 #(
		.INIT('h8)
	) name1338 (
		\137GAT(8)_pad ,
		\477GAT(28)_pad ,
		_w1371_
	);
	LUT2 #(
		.INIT('h1)
	) name1339 (
		_w1327_,
		_w1330_,
		_w1372_
	);
	LUT2 #(
		.INIT('h8)
	) name1340 (
		\154GAT(9)_pad ,
		\460GAT(27)_pad ,
		_w1373_
	);
	LUT2 #(
		.INIT('h1)
	) name1341 (
		_w1321_,
		_w1324_,
		_w1374_
	);
	LUT2 #(
		.INIT('h8)
	) name1342 (
		\171GAT(10)_pad ,
		\443GAT(26)_pad ,
		_w1375_
	);
	LUT2 #(
		.INIT('h1)
	) name1343 (
		_w1315_,
		_w1318_,
		_w1376_
	);
	LUT2 #(
		.INIT('h8)
	) name1344 (
		\188GAT(11)_pad ,
		\426GAT(25)_pad ,
		_w1377_
	);
	LUT2 #(
		.INIT('h1)
	) name1345 (
		_w1309_,
		_w1312_,
		_w1378_
	);
	LUT2 #(
		.INIT('h8)
	) name1346 (
		\205GAT(12)_pad ,
		\409GAT(24)_pad ,
		_w1379_
	);
	LUT2 #(
		.INIT('h1)
	) name1347 (
		_w1303_,
		_w1306_,
		_w1380_
	);
	LUT2 #(
		.INIT('h8)
	) name1348 (
		\222GAT(13)_pad ,
		\392GAT(23)_pad ,
		_w1381_
	);
	LUT2 #(
		.INIT('h1)
	) name1349 (
		_w1297_,
		_w1300_,
		_w1382_
	);
	LUT2 #(
		.INIT('h8)
	) name1350 (
		\239GAT(14)_pad ,
		\375GAT(22)_pad ,
		_w1383_
	);
	LUT2 #(
		.INIT('h1)
	) name1351 (
		_w1291_,
		_w1294_,
		_w1384_
	);
	LUT2 #(
		.INIT('h8)
	) name1352 (
		\256GAT(15)_pad ,
		\358GAT(21)_pad ,
		_w1385_
	);
	LUT2 #(
		.INIT('h1)
	) name1353 (
		_w1384_,
		_w1385_,
		_w1386_
	);
	LUT2 #(
		.INIT('h8)
	) name1354 (
		_w1384_,
		_w1385_,
		_w1387_
	);
	LUT2 #(
		.INIT('h1)
	) name1355 (
		_w1386_,
		_w1387_,
		_w1388_
	);
	LUT2 #(
		.INIT('h4)
	) name1356 (
		_w1383_,
		_w1388_,
		_w1389_
	);
	LUT2 #(
		.INIT('h2)
	) name1357 (
		_w1383_,
		_w1388_,
		_w1390_
	);
	LUT2 #(
		.INIT('h1)
	) name1358 (
		_w1389_,
		_w1390_,
		_w1391_
	);
	LUT2 #(
		.INIT('h4)
	) name1359 (
		_w1382_,
		_w1391_,
		_w1392_
	);
	LUT2 #(
		.INIT('h2)
	) name1360 (
		_w1382_,
		_w1391_,
		_w1393_
	);
	LUT2 #(
		.INIT('h1)
	) name1361 (
		_w1392_,
		_w1393_,
		_w1394_
	);
	LUT2 #(
		.INIT('h4)
	) name1362 (
		_w1381_,
		_w1394_,
		_w1395_
	);
	LUT2 #(
		.INIT('h2)
	) name1363 (
		_w1381_,
		_w1394_,
		_w1396_
	);
	LUT2 #(
		.INIT('h1)
	) name1364 (
		_w1395_,
		_w1396_,
		_w1397_
	);
	LUT2 #(
		.INIT('h4)
	) name1365 (
		_w1380_,
		_w1397_,
		_w1398_
	);
	LUT2 #(
		.INIT('h2)
	) name1366 (
		_w1380_,
		_w1397_,
		_w1399_
	);
	LUT2 #(
		.INIT('h1)
	) name1367 (
		_w1398_,
		_w1399_,
		_w1400_
	);
	LUT2 #(
		.INIT('h4)
	) name1368 (
		_w1379_,
		_w1400_,
		_w1401_
	);
	LUT2 #(
		.INIT('h2)
	) name1369 (
		_w1379_,
		_w1400_,
		_w1402_
	);
	LUT2 #(
		.INIT('h1)
	) name1370 (
		_w1401_,
		_w1402_,
		_w1403_
	);
	LUT2 #(
		.INIT('h4)
	) name1371 (
		_w1378_,
		_w1403_,
		_w1404_
	);
	LUT2 #(
		.INIT('h2)
	) name1372 (
		_w1378_,
		_w1403_,
		_w1405_
	);
	LUT2 #(
		.INIT('h1)
	) name1373 (
		_w1404_,
		_w1405_,
		_w1406_
	);
	LUT2 #(
		.INIT('h4)
	) name1374 (
		_w1377_,
		_w1406_,
		_w1407_
	);
	LUT2 #(
		.INIT('h2)
	) name1375 (
		_w1377_,
		_w1406_,
		_w1408_
	);
	LUT2 #(
		.INIT('h1)
	) name1376 (
		_w1407_,
		_w1408_,
		_w1409_
	);
	LUT2 #(
		.INIT('h4)
	) name1377 (
		_w1376_,
		_w1409_,
		_w1410_
	);
	LUT2 #(
		.INIT('h2)
	) name1378 (
		_w1376_,
		_w1409_,
		_w1411_
	);
	LUT2 #(
		.INIT('h1)
	) name1379 (
		_w1410_,
		_w1411_,
		_w1412_
	);
	LUT2 #(
		.INIT('h4)
	) name1380 (
		_w1375_,
		_w1412_,
		_w1413_
	);
	LUT2 #(
		.INIT('h2)
	) name1381 (
		_w1375_,
		_w1412_,
		_w1414_
	);
	LUT2 #(
		.INIT('h1)
	) name1382 (
		_w1413_,
		_w1414_,
		_w1415_
	);
	LUT2 #(
		.INIT('h4)
	) name1383 (
		_w1374_,
		_w1415_,
		_w1416_
	);
	LUT2 #(
		.INIT('h2)
	) name1384 (
		_w1374_,
		_w1415_,
		_w1417_
	);
	LUT2 #(
		.INIT('h1)
	) name1385 (
		_w1416_,
		_w1417_,
		_w1418_
	);
	LUT2 #(
		.INIT('h4)
	) name1386 (
		_w1373_,
		_w1418_,
		_w1419_
	);
	LUT2 #(
		.INIT('h2)
	) name1387 (
		_w1373_,
		_w1418_,
		_w1420_
	);
	LUT2 #(
		.INIT('h1)
	) name1388 (
		_w1419_,
		_w1420_,
		_w1421_
	);
	LUT2 #(
		.INIT('h4)
	) name1389 (
		_w1372_,
		_w1421_,
		_w1422_
	);
	LUT2 #(
		.INIT('h2)
	) name1390 (
		_w1372_,
		_w1421_,
		_w1423_
	);
	LUT2 #(
		.INIT('h1)
	) name1391 (
		_w1422_,
		_w1423_,
		_w1424_
	);
	LUT2 #(
		.INIT('h4)
	) name1392 (
		_w1371_,
		_w1424_,
		_w1425_
	);
	LUT2 #(
		.INIT('h2)
	) name1393 (
		_w1371_,
		_w1424_,
		_w1426_
	);
	LUT2 #(
		.INIT('h1)
	) name1394 (
		_w1425_,
		_w1426_,
		_w1427_
	);
	LUT2 #(
		.INIT('h4)
	) name1395 (
		_w1370_,
		_w1427_,
		_w1428_
	);
	LUT2 #(
		.INIT('h2)
	) name1396 (
		_w1370_,
		_w1427_,
		_w1429_
	);
	LUT2 #(
		.INIT('h1)
	) name1397 (
		_w1428_,
		_w1429_,
		_w1430_
	);
	LUT2 #(
		.INIT('h4)
	) name1398 (
		_w1369_,
		_w1430_,
		_w1431_
	);
	LUT2 #(
		.INIT('h2)
	) name1399 (
		_w1369_,
		_w1430_,
		_w1432_
	);
	LUT2 #(
		.INIT('h1)
	) name1400 (
		_w1431_,
		_w1432_,
		_w1433_
	);
	LUT2 #(
		.INIT('h4)
	) name1401 (
		_w1368_,
		_w1433_,
		_w1434_
	);
	LUT2 #(
		.INIT('h2)
	) name1402 (
		_w1368_,
		_w1433_,
		_w1435_
	);
	LUT2 #(
		.INIT('h1)
	) name1403 (
		_w1434_,
		_w1435_,
		_w1436_
	);
	LUT2 #(
		.INIT('h4)
	) name1404 (
		_w1367_,
		_w1436_,
		_w1437_
	);
	LUT2 #(
		.INIT('h2)
	) name1405 (
		_w1367_,
		_w1436_,
		_w1438_
	);
	LUT2 #(
		.INIT('h1)
	) name1406 (
		_w1437_,
		_w1438_,
		_w1439_
	);
	LUT2 #(
		.INIT('h4)
	) name1407 (
		_w1366_,
		_w1439_,
		_w1440_
	);
	LUT2 #(
		.INIT('h2)
	) name1408 (
		_w1366_,
		_w1439_,
		_w1441_
	);
	LUT2 #(
		.INIT('h1)
	) name1409 (
		_w1440_,
		_w1441_,
		_w1442_
	);
	LUT2 #(
		.INIT('h4)
	) name1410 (
		_w1365_,
		_w1442_,
		_w1443_
	);
	LUT2 #(
		.INIT('h2)
	) name1411 (
		_w1365_,
		_w1442_,
		_w1444_
	);
	LUT2 #(
		.INIT('h1)
	) name1412 (
		_w1443_,
		_w1444_,
		_w1445_
	);
	LUT2 #(
		.INIT('h4)
	) name1413 (
		_w1364_,
		_w1445_,
		_w1446_
	);
	LUT2 #(
		.INIT('h2)
	) name1414 (
		_w1364_,
		_w1445_,
		_w1447_
	);
	LUT2 #(
		.INIT('h1)
	) name1415 (
		_w1446_,
		_w1447_,
		_w1448_
	);
	LUT2 #(
		.INIT('h4)
	) name1416 (
		_w1363_,
		_w1448_,
		_w1449_
	);
	LUT2 #(
		.INIT('h2)
	) name1417 (
		_w1363_,
		_w1448_,
		_w1450_
	);
	LUT2 #(
		.INIT('h1)
	) name1418 (
		_w1449_,
		_w1450_,
		_w1451_
	);
	LUT2 #(
		.INIT('h1)
	) name1419 (
		_w1446_,
		_w1449_,
		_w1452_
	);
	LUT2 #(
		.INIT('h1)
	) name1420 (
		_w1440_,
		_w1443_,
		_w1453_
	);
	LUT2 #(
		.INIT('h8)
	) name1421 (
		\103GAT(6)_pad ,
		\528GAT(31)_pad ,
		_w1454_
	);
	LUT2 #(
		.INIT('h1)
	) name1422 (
		_w1434_,
		_w1437_,
		_w1455_
	);
	LUT2 #(
		.INIT('h8)
	) name1423 (
		\120GAT(7)_pad ,
		\511GAT(30)_pad ,
		_w1456_
	);
	LUT2 #(
		.INIT('h1)
	) name1424 (
		_w1428_,
		_w1431_,
		_w1457_
	);
	LUT2 #(
		.INIT('h8)
	) name1425 (
		\137GAT(8)_pad ,
		\494GAT(29)_pad ,
		_w1458_
	);
	LUT2 #(
		.INIT('h1)
	) name1426 (
		_w1422_,
		_w1425_,
		_w1459_
	);
	LUT2 #(
		.INIT('h8)
	) name1427 (
		\154GAT(9)_pad ,
		\477GAT(28)_pad ,
		_w1460_
	);
	LUT2 #(
		.INIT('h1)
	) name1428 (
		_w1416_,
		_w1419_,
		_w1461_
	);
	LUT2 #(
		.INIT('h8)
	) name1429 (
		\171GAT(10)_pad ,
		\460GAT(27)_pad ,
		_w1462_
	);
	LUT2 #(
		.INIT('h1)
	) name1430 (
		_w1410_,
		_w1413_,
		_w1463_
	);
	LUT2 #(
		.INIT('h8)
	) name1431 (
		\188GAT(11)_pad ,
		\443GAT(26)_pad ,
		_w1464_
	);
	LUT2 #(
		.INIT('h1)
	) name1432 (
		_w1404_,
		_w1407_,
		_w1465_
	);
	LUT2 #(
		.INIT('h8)
	) name1433 (
		\205GAT(12)_pad ,
		\426GAT(25)_pad ,
		_w1466_
	);
	LUT2 #(
		.INIT('h1)
	) name1434 (
		_w1398_,
		_w1401_,
		_w1467_
	);
	LUT2 #(
		.INIT('h8)
	) name1435 (
		\222GAT(13)_pad ,
		\409GAT(24)_pad ,
		_w1468_
	);
	LUT2 #(
		.INIT('h1)
	) name1436 (
		_w1392_,
		_w1395_,
		_w1469_
	);
	LUT2 #(
		.INIT('h8)
	) name1437 (
		\239GAT(14)_pad ,
		\392GAT(23)_pad ,
		_w1470_
	);
	LUT2 #(
		.INIT('h1)
	) name1438 (
		_w1386_,
		_w1389_,
		_w1471_
	);
	LUT2 #(
		.INIT('h8)
	) name1439 (
		\256GAT(15)_pad ,
		\375GAT(22)_pad ,
		_w1472_
	);
	LUT2 #(
		.INIT('h1)
	) name1440 (
		_w1471_,
		_w1472_,
		_w1473_
	);
	LUT2 #(
		.INIT('h8)
	) name1441 (
		_w1471_,
		_w1472_,
		_w1474_
	);
	LUT2 #(
		.INIT('h1)
	) name1442 (
		_w1473_,
		_w1474_,
		_w1475_
	);
	LUT2 #(
		.INIT('h4)
	) name1443 (
		_w1470_,
		_w1475_,
		_w1476_
	);
	LUT2 #(
		.INIT('h2)
	) name1444 (
		_w1470_,
		_w1475_,
		_w1477_
	);
	LUT2 #(
		.INIT('h1)
	) name1445 (
		_w1476_,
		_w1477_,
		_w1478_
	);
	LUT2 #(
		.INIT('h4)
	) name1446 (
		_w1469_,
		_w1478_,
		_w1479_
	);
	LUT2 #(
		.INIT('h2)
	) name1447 (
		_w1469_,
		_w1478_,
		_w1480_
	);
	LUT2 #(
		.INIT('h1)
	) name1448 (
		_w1479_,
		_w1480_,
		_w1481_
	);
	LUT2 #(
		.INIT('h4)
	) name1449 (
		_w1468_,
		_w1481_,
		_w1482_
	);
	LUT2 #(
		.INIT('h2)
	) name1450 (
		_w1468_,
		_w1481_,
		_w1483_
	);
	LUT2 #(
		.INIT('h1)
	) name1451 (
		_w1482_,
		_w1483_,
		_w1484_
	);
	LUT2 #(
		.INIT('h4)
	) name1452 (
		_w1467_,
		_w1484_,
		_w1485_
	);
	LUT2 #(
		.INIT('h2)
	) name1453 (
		_w1467_,
		_w1484_,
		_w1486_
	);
	LUT2 #(
		.INIT('h1)
	) name1454 (
		_w1485_,
		_w1486_,
		_w1487_
	);
	LUT2 #(
		.INIT('h4)
	) name1455 (
		_w1466_,
		_w1487_,
		_w1488_
	);
	LUT2 #(
		.INIT('h2)
	) name1456 (
		_w1466_,
		_w1487_,
		_w1489_
	);
	LUT2 #(
		.INIT('h1)
	) name1457 (
		_w1488_,
		_w1489_,
		_w1490_
	);
	LUT2 #(
		.INIT('h4)
	) name1458 (
		_w1465_,
		_w1490_,
		_w1491_
	);
	LUT2 #(
		.INIT('h2)
	) name1459 (
		_w1465_,
		_w1490_,
		_w1492_
	);
	LUT2 #(
		.INIT('h1)
	) name1460 (
		_w1491_,
		_w1492_,
		_w1493_
	);
	LUT2 #(
		.INIT('h4)
	) name1461 (
		_w1464_,
		_w1493_,
		_w1494_
	);
	LUT2 #(
		.INIT('h2)
	) name1462 (
		_w1464_,
		_w1493_,
		_w1495_
	);
	LUT2 #(
		.INIT('h1)
	) name1463 (
		_w1494_,
		_w1495_,
		_w1496_
	);
	LUT2 #(
		.INIT('h4)
	) name1464 (
		_w1463_,
		_w1496_,
		_w1497_
	);
	LUT2 #(
		.INIT('h2)
	) name1465 (
		_w1463_,
		_w1496_,
		_w1498_
	);
	LUT2 #(
		.INIT('h1)
	) name1466 (
		_w1497_,
		_w1498_,
		_w1499_
	);
	LUT2 #(
		.INIT('h4)
	) name1467 (
		_w1462_,
		_w1499_,
		_w1500_
	);
	LUT2 #(
		.INIT('h2)
	) name1468 (
		_w1462_,
		_w1499_,
		_w1501_
	);
	LUT2 #(
		.INIT('h1)
	) name1469 (
		_w1500_,
		_w1501_,
		_w1502_
	);
	LUT2 #(
		.INIT('h4)
	) name1470 (
		_w1461_,
		_w1502_,
		_w1503_
	);
	LUT2 #(
		.INIT('h2)
	) name1471 (
		_w1461_,
		_w1502_,
		_w1504_
	);
	LUT2 #(
		.INIT('h1)
	) name1472 (
		_w1503_,
		_w1504_,
		_w1505_
	);
	LUT2 #(
		.INIT('h4)
	) name1473 (
		_w1460_,
		_w1505_,
		_w1506_
	);
	LUT2 #(
		.INIT('h2)
	) name1474 (
		_w1460_,
		_w1505_,
		_w1507_
	);
	LUT2 #(
		.INIT('h1)
	) name1475 (
		_w1506_,
		_w1507_,
		_w1508_
	);
	LUT2 #(
		.INIT('h4)
	) name1476 (
		_w1459_,
		_w1508_,
		_w1509_
	);
	LUT2 #(
		.INIT('h2)
	) name1477 (
		_w1459_,
		_w1508_,
		_w1510_
	);
	LUT2 #(
		.INIT('h1)
	) name1478 (
		_w1509_,
		_w1510_,
		_w1511_
	);
	LUT2 #(
		.INIT('h4)
	) name1479 (
		_w1458_,
		_w1511_,
		_w1512_
	);
	LUT2 #(
		.INIT('h2)
	) name1480 (
		_w1458_,
		_w1511_,
		_w1513_
	);
	LUT2 #(
		.INIT('h1)
	) name1481 (
		_w1512_,
		_w1513_,
		_w1514_
	);
	LUT2 #(
		.INIT('h4)
	) name1482 (
		_w1457_,
		_w1514_,
		_w1515_
	);
	LUT2 #(
		.INIT('h2)
	) name1483 (
		_w1457_,
		_w1514_,
		_w1516_
	);
	LUT2 #(
		.INIT('h1)
	) name1484 (
		_w1515_,
		_w1516_,
		_w1517_
	);
	LUT2 #(
		.INIT('h4)
	) name1485 (
		_w1456_,
		_w1517_,
		_w1518_
	);
	LUT2 #(
		.INIT('h2)
	) name1486 (
		_w1456_,
		_w1517_,
		_w1519_
	);
	LUT2 #(
		.INIT('h1)
	) name1487 (
		_w1518_,
		_w1519_,
		_w1520_
	);
	LUT2 #(
		.INIT('h4)
	) name1488 (
		_w1455_,
		_w1520_,
		_w1521_
	);
	LUT2 #(
		.INIT('h2)
	) name1489 (
		_w1455_,
		_w1520_,
		_w1522_
	);
	LUT2 #(
		.INIT('h1)
	) name1490 (
		_w1521_,
		_w1522_,
		_w1523_
	);
	LUT2 #(
		.INIT('h4)
	) name1491 (
		_w1454_,
		_w1523_,
		_w1524_
	);
	LUT2 #(
		.INIT('h2)
	) name1492 (
		_w1454_,
		_w1523_,
		_w1525_
	);
	LUT2 #(
		.INIT('h1)
	) name1493 (
		_w1524_,
		_w1525_,
		_w1526_
	);
	LUT2 #(
		.INIT('h4)
	) name1494 (
		_w1453_,
		_w1526_,
		_w1527_
	);
	LUT2 #(
		.INIT('h2)
	) name1495 (
		_w1453_,
		_w1526_,
		_w1528_
	);
	LUT2 #(
		.INIT('h1)
	) name1496 (
		_w1527_,
		_w1528_,
		_w1529_
	);
	LUT2 #(
		.INIT('h4)
	) name1497 (
		_w1452_,
		_w1529_,
		_w1530_
	);
	LUT2 #(
		.INIT('h2)
	) name1498 (
		_w1452_,
		_w1529_,
		_w1531_
	);
	LUT2 #(
		.INIT('h1)
	) name1499 (
		_w1530_,
		_w1531_,
		_w1532_
	);
	LUT2 #(
		.INIT('h1)
	) name1500 (
		_w1527_,
		_w1530_,
		_w1533_
	);
	LUT2 #(
		.INIT('h1)
	) name1501 (
		_w1521_,
		_w1524_,
		_w1534_
	);
	LUT2 #(
		.INIT('h8)
	) name1502 (
		\120GAT(7)_pad ,
		\528GAT(31)_pad ,
		_w1535_
	);
	LUT2 #(
		.INIT('h1)
	) name1503 (
		_w1515_,
		_w1518_,
		_w1536_
	);
	LUT2 #(
		.INIT('h8)
	) name1504 (
		\137GAT(8)_pad ,
		\511GAT(30)_pad ,
		_w1537_
	);
	LUT2 #(
		.INIT('h1)
	) name1505 (
		_w1509_,
		_w1512_,
		_w1538_
	);
	LUT2 #(
		.INIT('h8)
	) name1506 (
		\154GAT(9)_pad ,
		\494GAT(29)_pad ,
		_w1539_
	);
	LUT2 #(
		.INIT('h1)
	) name1507 (
		_w1503_,
		_w1506_,
		_w1540_
	);
	LUT2 #(
		.INIT('h8)
	) name1508 (
		\171GAT(10)_pad ,
		\477GAT(28)_pad ,
		_w1541_
	);
	LUT2 #(
		.INIT('h1)
	) name1509 (
		_w1497_,
		_w1500_,
		_w1542_
	);
	LUT2 #(
		.INIT('h8)
	) name1510 (
		\188GAT(11)_pad ,
		\460GAT(27)_pad ,
		_w1543_
	);
	LUT2 #(
		.INIT('h1)
	) name1511 (
		_w1491_,
		_w1494_,
		_w1544_
	);
	LUT2 #(
		.INIT('h8)
	) name1512 (
		\205GAT(12)_pad ,
		\443GAT(26)_pad ,
		_w1545_
	);
	LUT2 #(
		.INIT('h1)
	) name1513 (
		_w1485_,
		_w1488_,
		_w1546_
	);
	LUT2 #(
		.INIT('h8)
	) name1514 (
		\222GAT(13)_pad ,
		\426GAT(25)_pad ,
		_w1547_
	);
	LUT2 #(
		.INIT('h1)
	) name1515 (
		_w1479_,
		_w1482_,
		_w1548_
	);
	LUT2 #(
		.INIT('h8)
	) name1516 (
		\239GAT(14)_pad ,
		\409GAT(24)_pad ,
		_w1549_
	);
	LUT2 #(
		.INIT('h1)
	) name1517 (
		_w1473_,
		_w1476_,
		_w1550_
	);
	LUT2 #(
		.INIT('h8)
	) name1518 (
		\256GAT(15)_pad ,
		\392GAT(23)_pad ,
		_w1551_
	);
	LUT2 #(
		.INIT('h1)
	) name1519 (
		_w1550_,
		_w1551_,
		_w1552_
	);
	LUT2 #(
		.INIT('h8)
	) name1520 (
		_w1550_,
		_w1551_,
		_w1553_
	);
	LUT2 #(
		.INIT('h1)
	) name1521 (
		_w1552_,
		_w1553_,
		_w1554_
	);
	LUT2 #(
		.INIT('h4)
	) name1522 (
		_w1549_,
		_w1554_,
		_w1555_
	);
	LUT2 #(
		.INIT('h2)
	) name1523 (
		_w1549_,
		_w1554_,
		_w1556_
	);
	LUT2 #(
		.INIT('h1)
	) name1524 (
		_w1555_,
		_w1556_,
		_w1557_
	);
	LUT2 #(
		.INIT('h4)
	) name1525 (
		_w1548_,
		_w1557_,
		_w1558_
	);
	LUT2 #(
		.INIT('h2)
	) name1526 (
		_w1548_,
		_w1557_,
		_w1559_
	);
	LUT2 #(
		.INIT('h1)
	) name1527 (
		_w1558_,
		_w1559_,
		_w1560_
	);
	LUT2 #(
		.INIT('h4)
	) name1528 (
		_w1547_,
		_w1560_,
		_w1561_
	);
	LUT2 #(
		.INIT('h2)
	) name1529 (
		_w1547_,
		_w1560_,
		_w1562_
	);
	LUT2 #(
		.INIT('h1)
	) name1530 (
		_w1561_,
		_w1562_,
		_w1563_
	);
	LUT2 #(
		.INIT('h4)
	) name1531 (
		_w1546_,
		_w1563_,
		_w1564_
	);
	LUT2 #(
		.INIT('h2)
	) name1532 (
		_w1546_,
		_w1563_,
		_w1565_
	);
	LUT2 #(
		.INIT('h1)
	) name1533 (
		_w1564_,
		_w1565_,
		_w1566_
	);
	LUT2 #(
		.INIT('h4)
	) name1534 (
		_w1545_,
		_w1566_,
		_w1567_
	);
	LUT2 #(
		.INIT('h2)
	) name1535 (
		_w1545_,
		_w1566_,
		_w1568_
	);
	LUT2 #(
		.INIT('h1)
	) name1536 (
		_w1567_,
		_w1568_,
		_w1569_
	);
	LUT2 #(
		.INIT('h4)
	) name1537 (
		_w1544_,
		_w1569_,
		_w1570_
	);
	LUT2 #(
		.INIT('h2)
	) name1538 (
		_w1544_,
		_w1569_,
		_w1571_
	);
	LUT2 #(
		.INIT('h1)
	) name1539 (
		_w1570_,
		_w1571_,
		_w1572_
	);
	LUT2 #(
		.INIT('h4)
	) name1540 (
		_w1543_,
		_w1572_,
		_w1573_
	);
	LUT2 #(
		.INIT('h2)
	) name1541 (
		_w1543_,
		_w1572_,
		_w1574_
	);
	LUT2 #(
		.INIT('h1)
	) name1542 (
		_w1573_,
		_w1574_,
		_w1575_
	);
	LUT2 #(
		.INIT('h4)
	) name1543 (
		_w1542_,
		_w1575_,
		_w1576_
	);
	LUT2 #(
		.INIT('h2)
	) name1544 (
		_w1542_,
		_w1575_,
		_w1577_
	);
	LUT2 #(
		.INIT('h1)
	) name1545 (
		_w1576_,
		_w1577_,
		_w1578_
	);
	LUT2 #(
		.INIT('h4)
	) name1546 (
		_w1541_,
		_w1578_,
		_w1579_
	);
	LUT2 #(
		.INIT('h2)
	) name1547 (
		_w1541_,
		_w1578_,
		_w1580_
	);
	LUT2 #(
		.INIT('h1)
	) name1548 (
		_w1579_,
		_w1580_,
		_w1581_
	);
	LUT2 #(
		.INIT('h4)
	) name1549 (
		_w1540_,
		_w1581_,
		_w1582_
	);
	LUT2 #(
		.INIT('h2)
	) name1550 (
		_w1540_,
		_w1581_,
		_w1583_
	);
	LUT2 #(
		.INIT('h1)
	) name1551 (
		_w1582_,
		_w1583_,
		_w1584_
	);
	LUT2 #(
		.INIT('h4)
	) name1552 (
		_w1539_,
		_w1584_,
		_w1585_
	);
	LUT2 #(
		.INIT('h2)
	) name1553 (
		_w1539_,
		_w1584_,
		_w1586_
	);
	LUT2 #(
		.INIT('h1)
	) name1554 (
		_w1585_,
		_w1586_,
		_w1587_
	);
	LUT2 #(
		.INIT('h4)
	) name1555 (
		_w1538_,
		_w1587_,
		_w1588_
	);
	LUT2 #(
		.INIT('h2)
	) name1556 (
		_w1538_,
		_w1587_,
		_w1589_
	);
	LUT2 #(
		.INIT('h1)
	) name1557 (
		_w1588_,
		_w1589_,
		_w1590_
	);
	LUT2 #(
		.INIT('h4)
	) name1558 (
		_w1537_,
		_w1590_,
		_w1591_
	);
	LUT2 #(
		.INIT('h2)
	) name1559 (
		_w1537_,
		_w1590_,
		_w1592_
	);
	LUT2 #(
		.INIT('h1)
	) name1560 (
		_w1591_,
		_w1592_,
		_w1593_
	);
	LUT2 #(
		.INIT('h4)
	) name1561 (
		_w1536_,
		_w1593_,
		_w1594_
	);
	LUT2 #(
		.INIT('h2)
	) name1562 (
		_w1536_,
		_w1593_,
		_w1595_
	);
	LUT2 #(
		.INIT('h1)
	) name1563 (
		_w1594_,
		_w1595_,
		_w1596_
	);
	LUT2 #(
		.INIT('h4)
	) name1564 (
		_w1535_,
		_w1596_,
		_w1597_
	);
	LUT2 #(
		.INIT('h2)
	) name1565 (
		_w1535_,
		_w1596_,
		_w1598_
	);
	LUT2 #(
		.INIT('h1)
	) name1566 (
		_w1597_,
		_w1598_,
		_w1599_
	);
	LUT2 #(
		.INIT('h4)
	) name1567 (
		_w1534_,
		_w1599_,
		_w1600_
	);
	LUT2 #(
		.INIT('h2)
	) name1568 (
		_w1534_,
		_w1599_,
		_w1601_
	);
	LUT2 #(
		.INIT('h1)
	) name1569 (
		_w1600_,
		_w1601_,
		_w1602_
	);
	LUT2 #(
		.INIT('h4)
	) name1570 (
		_w1533_,
		_w1602_,
		_w1603_
	);
	LUT2 #(
		.INIT('h2)
	) name1571 (
		_w1533_,
		_w1602_,
		_w1604_
	);
	LUT2 #(
		.INIT('h1)
	) name1572 (
		_w1603_,
		_w1604_,
		_w1605_
	);
	LUT2 #(
		.INIT('h1)
	) name1573 (
		_w1600_,
		_w1603_,
		_w1606_
	);
	LUT2 #(
		.INIT('h1)
	) name1574 (
		_w1594_,
		_w1597_,
		_w1607_
	);
	LUT2 #(
		.INIT('h8)
	) name1575 (
		\137GAT(8)_pad ,
		\528GAT(31)_pad ,
		_w1608_
	);
	LUT2 #(
		.INIT('h1)
	) name1576 (
		_w1588_,
		_w1591_,
		_w1609_
	);
	LUT2 #(
		.INIT('h8)
	) name1577 (
		\154GAT(9)_pad ,
		\511GAT(30)_pad ,
		_w1610_
	);
	LUT2 #(
		.INIT('h1)
	) name1578 (
		_w1582_,
		_w1585_,
		_w1611_
	);
	LUT2 #(
		.INIT('h8)
	) name1579 (
		\171GAT(10)_pad ,
		\494GAT(29)_pad ,
		_w1612_
	);
	LUT2 #(
		.INIT('h1)
	) name1580 (
		_w1576_,
		_w1579_,
		_w1613_
	);
	LUT2 #(
		.INIT('h8)
	) name1581 (
		\188GAT(11)_pad ,
		\477GAT(28)_pad ,
		_w1614_
	);
	LUT2 #(
		.INIT('h1)
	) name1582 (
		_w1570_,
		_w1573_,
		_w1615_
	);
	LUT2 #(
		.INIT('h8)
	) name1583 (
		\205GAT(12)_pad ,
		\460GAT(27)_pad ,
		_w1616_
	);
	LUT2 #(
		.INIT('h1)
	) name1584 (
		_w1564_,
		_w1567_,
		_w1617_
	);
	LUT2 #(
		.INIT('h8)
	) name1585 (
		\222GAT(13)_pad ,
		\443GAT(26)_pad ,
		_w1618_
	);
	LUT2 #(
		.INIT('h1)
	) name1586 (
		_w1558_,
		_w1561_,
		_w1619_
	);
	LUT2 #(
		.INIT('h8)
	) name1587 (
		\239GAT(14)_pad ,
		\426GAT(25)_pad ,
		_w1620_
	);
	LUT2 #(
		.INIT('h1)
	) name1588 (
		_w1552_,
		_w1555_,
		_w1621_
	);
	LUT2 #(
		.INIT('h8)
	) name1589 (
		\256GAT(15)_pad ,
		\409GAT(24)_pad ,
		_w1622_
	);
	LUT2 #(
		.INIT('h1)
	) name1590 (
		_w1621_,
		_w1622_,
		_w1623_
	);
	LUT2 #(
		.INIT('h8)
	) name1591 (
		_w1621_,
		_w1622_,
		_w1624_
	);
	LUT2 #(
		.INIT('h1)
	) name1592 (
		_w1623_,
		_w1624_,
		_w1625_
	);
	LUT2 #(
		.INIT('h4)
	) name1593 (
		_w1620_,
		_w1625_,
		_w1626_
	);
	LUT2 #(
		.INIT('h2)
	) name1594 (
		_w1620_,
		_w1625_,
		_w1627_
	);
	LUT2 #(
		.INIT('h1)
	) name1595 (
		_w1626_,
		_w1627_,
		_w1628_
	);
	LUT2 #(
		.INIT('h4)
	) name1596 (
		_w1619_,
		_w1628_,
		_w1629_
	);
	LUT2 #(
		.INIT('h2)
	) name1597 (
		_w1619_,
		_w1628_,
		_w1630_
	);
	LUT2 #(
		.INIT('h1)
	) name1598 (
		_w1629_,
		_w1630_,
		_w1631_
	);
	LUT2 #(
		.INIT('h4)
	) name1599 (
		_w1618_,
		_w1631_,
		_w1632_
	);
	LUT2 #(
		.INIT('h2)
	) name1600 (
		_w1618_,
		_w1631_,
		_w1633_
	);
	LUT2 #(
		.INIT('h1)
	) name1601 (
		_w1632_,
		_w1633_,
		_w1634_
	);
	LUT2 #(
		.INIT('h4)
	) name1602 (
		_w1617_,
		_w1634_,
		_w1635_
	);
	LUT2 #(
		.INIT('h2)
	) name1603 (
		_w1617_,
		_w1634_,
		_w1636_
	);
	LUT2 #(
		.INIT('h1)
	) name1604 (
		_w1635_,
		_w1636_,
		_w1637_
	);
	LUT2 #(
		.INIT('h4)
	) name1605 (
		_w1616_,
		_w1637_,
		_w1638_
	);
	LUT2 #(
		.INIT('h2)
	) name1606 (
		_w1616_,
		_w1637_,
		_w1639_
	);
	LUT2 #(
		.INIT('h1)
	) name1607 (
		_w1638_,
		_w1639_,
		_w1640_
	);
	LUT2 #(
		.INIT('h4)
	) name1608 (
		_w1615_,
		_w1640_,
		_w1641_
	);
	LUT2 #(
		.INIT('h2)
	) name1609 (
		_w1615_,
		_w1640_,
		_w1642_
	);
	LUT2 #(
		.INIT('h1)
	) name1610 (
		_w1641_,
		_w1642_,
		_w1643_
	);
	LUT2 #(
		.INIT('h4)
	) name1611 (
		_w1614_,
		_w1643_,
		_w1644_
	);
	LUT2 #(
		.INIT('h2)
	) name1612 (
		_w1614_,
		_w1643_,
		_w1645_
	);
	LUT2 #(
		.INIT('h1)
	) name1613 (
		_w1644_,
		_w1645_,
		_w1646_
	);
	LUT2 #(
		.INIT('h4)
	) name1614 (
		_w1613_,
		_w1646_,
		_w1647_
	);
	LUT2 #(
		.INIT('h2)
	) name1615 (
		_w1613_,
		_w1646_,
		_w1648_
	);
	LUT2 #(
		.INIT('h1)
	) name1616 (
		_w1647_,
		_w1648_,
		_w1649_
	);
	LUT2 #(
		.INIT('h4)
	) name1617 (
		_w1612_,
		_w1649_,
		_w1650_
	);
	LUT2 #(
		.INIT('h2)
	) name1618 (
		_w1612_,
		_w1649_,
		_w1651_
	);
	LUT2 #(
		.INIT('h1)
	) name1619 (
		_w1650_,
		_w1651_,
		_w1652_
	);
	LUT2 #(
		.INIT('h4)
	) name1620 (
		_w1611_,
		_w1652_,
		_w1653_
	);
	LUT2 #(
		.INIT('h2)
	) name1621 (
		_w1611_,
		_w1652_,
		_w1654_
	);
	LUT2 #(
		.INIT('h1)
	) name1622 (
		_w1653_,
		_w1654_,
		_w1655_
	);
	LUT2 #(
		.INIT('h4)
	) name1623 (
		_w1610_,
		_w1655_,
		_w1656_
	);
	LUT2 #(
		.INIT('h2)
	) name1624 (
		_w1610_,
		_w1655_,
		_w1657_
	);
	LUT2 #(
		.INIT('h1)
	) name1625 (
		_w1656_,
		_w1657_,
		_w1658_
	);
	LUT2 #(
		.INIT('h4)
	) name1626 (
		_w1609_,
		_w1658_,
		_w1659_
	);
	LUT2 #(
		.INIT('h2)
	) name1627 (
		_w1609_,
		_w1658_,
		_w1660_
	);
	LUT2 #(
		.INIT('h1)
	) name1628 (
		_w1659_,
		_w1660_,
		_w1661_
	);
	LUT2 #(
		.INIT('h4)
	) name1629 (
		_w1608_,
		_w1661_,
		_w1662_
	);
	LUT2 #(
		.INIT('h2)
	) name1630 (
		_w1608_,
		_w1661_,
		_w1663_
	);
	LUT2 #(
		.INIT('h1)
	) name1631 (
		_w1662_,
		_w1663_,
		_w1664_
	);
	LUT2 #(
		.INIT('h4)
	) name1632 (
		_w1607_,
		_w1664_,
		_w1665_
	);
	LUT2 #(
		.INIT('h2)
	) name1633 (
		_w1607_,
		_w1664_,
		_w1666_
	);
	LUT2 #(
		.INIT('h1)
	) name1634 (
		_w1665_,
		_w1666_,
		_w1667_
	);
	LUT2 #(
		.INIT('h4)
	) name1635 (
		_w1606_,
		_w1667_,
		_w1668_
	);
	LUT2 #(
		.INIT('h2)
	) name1636 (
		_w1606_,
		_w1667_,
		_w1669_
	);
	LUT2 #(
		.INIT('h1)
	) name1637 (
		_w1668_,
		_w1669_,
		_w1670_
	);
	LUT2 #(
		.INIT('h1)
	) name1638 (
		_w1665_,
		_w1668_,
		_w1671_
	);
	LUT2 #(
		.INIT('h1)
	) name1639 (
		_w1659_,
		_w1662_,
		_w1672_
	);
	LUT2 #(
		.INIT('h8)
	) name1640 (
		\154GAT(9)_pad ,
		\528GAT(31)_pad ,
		_w1673_
	);
	LUT2 #(
		.INIT('h1)
	) name1641 (
		_w1653_,
		_w1656_,
		_w1674_
	);
	LUT2 #(
		.INIT('h8)
	) name1642 (
		\171GAT(10)_pad ,
		\511GAT(30)_pad ,
		_w1675_
	);
	LUT2 #(
		.INIT('h1)
	) name1643 (
		_w1647_,
		_w1650_,
		_w1676_
	);
	LUT2 #(
		.INIT('h8)
	) name1644 (
		\188GAT(11)_pad ,
		\494GAT(29)_pad ,
		_w1677_
	);
	LUT2 #(
		.INIT('h1)
	) name1645 (
		_w1641_,
		_w1644_,
		_w1678_
	);
	LUT2 #(
		.INIT('h8)
	) name1646 (
		\205GAT(12)_pad ,
		\477GAT(28)_pad ,
		_w1679_
	);
	LUT2 #(
		.INIT('h1)
	) name1647 (
		_w1635_,
		_w1638_,
		_w1680_
	);
	LUT2 #(
		.INIT('h8)
	) name1648 (
		\222GAT(13)_pad ,
		\460GAT(27)_pad ,
		_w1681_
	);
	LUT2 #(
		.INIT('h1)
	) name1649 (
		_w1629_,
		_w1632_,
		_w1682_
	);
	LUT2 #(
		.INIT('h8)
	) name1650 (
		\239GAT(14)_pad ,
		\443GAT(26)_pad ,
		_w1683_
	);
	LUT2 #(
		.INIT('h1)
	) name1651 (
		_w1623_,
		_w1626_,
		_w1684_
	);
	LUT2 #(
		.INIT('h8)
	) name1652 (
		\256GAT(15)_pad ,
		\426GAT(25)_pad ,
		_w1685_
	);
	LUT2 #(
		.INIT('h1)
	) name1653 (
		_w1684_,
		_w1685_,
		_w1686_
	);
	LUT2 #(
		.INIT('h8)
	) name1654 (
		_w1684_,
		_w1685_,
		_w1687_
	);
	LUT2 #(
		.INIT('h1)
	) name1655 (
		_w1686_,
		_w1687_,
		_w1688_
	);
	LUT2 #(
		.INIT('h4)
	) name1656 (
		_w1683_,
		_w1688_,
		_w1689_
	);
	LUT2 #(
		.INIT('h2)
	) name1657 (
		_w1683_,
		_w1688_,
		_w1690_
	);
	LUT2 #(
		.INIT('h1)
	) name1658 (
		_w1689_,
		_w1690_,
		_w1691_
	);
	LUT2 #(
		.INIT('h4)
	) name1659 (
		_w1682_,
		_w1691_,
		_w1692_
	);
	LUT2 #(
		.INIT('h2)
	) name1660 (
		_w1682_,
		_w1691_,
		_w1693_
	);
	LUT2 #(
		.INIT('h1)
	) name1661 (
		_w1692_,
		_w1693_,
		_w1694_
	);
	LUT2 #(
		.INIT('h4)
	) name1662 (
		_w1681_,
		_w1694_,
		_w1695_
	);
	LUT2 #(
		.INIT('h2)
	) name1663 (
		_w1681_,
		_w1694_,
		_w1696_
	);
	LUT2 #(
		.INIT('h1)
	) name1664 (
		_w1695_,
		_w1696_,
		_w1697_
	);
	LUT2 #(
		.INIT('h4)
	) name1665 (
		_w1680_,
		_w1697_,
		_w1698_
	);
	LUT2 #(
		.INIT('h2)
	) name1666 (
		_w1680_,
		_w1697_,
		_w1699_
	);
	LUT2 #(
		.INIT('h1)
	) name1667 (
		_w1698_,
		_w1699_,
		_w1700_
	);
	LUT2 #(
		.INIT('h4)
	) name1668 (
		_w1679_,
		_w1700_,
		_w1701_
	);
	LUT2 #(
		.INIT('h2)
	) name1669 (
		_w1679_,
		_w1700_,
		_w1702_
	);
	LUT2 #(
		.INIT('h1)
	) name1670 (
		_w1701_,
		_w1702_,
		_w1703_
	);
	LUT2 #(
		.INIT('h4)
	) name1671 (
		_w1678_,
		_w1703_,
		_w1704_
	);
	LUT2 #(
		.INIT('h2)
	) name1672 (
		_w1678_,
		_w1703_,
		_w1705_
	);
	LUT2 #(
		.INIT('h1)
	) name1673 (
		_w1704_,
		_w1705_,
		_w1706_
	);
	LUT2 #(
		.INIT('h4)
	) name1674 (
		_w1677_,
		_w1706_,
		_w1707_
	);
	LUT2 #(
		.INIT('h2)
	) name1675 (
		_w1677_,
		_w1706_,
		_w1708_
	);
	LUT2 #(
		.INIT('h1)
	) name1676 (
		_w1707_,
		_w1708_,
		_w1709_
	);
	LUT2 #(
		.INIT('h4)
	) name1677 (
		_w1676_,
		_w1709_,
		_w1710_
	);
	LUT2 #(
		.INIT('h2)
	) name1678 (
		_w1676_,
		_w1709_,
		_w1711_
	);
	LUT2 #(
		.INIT('h1)
	) name1679 (
		_w1710_,
		_w1711_,
		_w1712_
	);
	LUT2 #(
		.INIT('h4)
	) name1680 (
		_w1675_,
		_w1712_,
		_w1713_
	);
	LUT2 #(
		.INIT('h2)
	) name1681 (
		_w1675_,
		_w1712_,
		_w1714_
	);
	LUT2 #(
		.INIT('h1)
	) name1682 (
		_w1713_,
		_w1714_,
		_w1715_
	);
	LUT2 #(
		.INIT('h4)
	) name1683 (
		_w1674_,
		_w1715_,
		_w1716_
	);
	LUT2 #(
		.INIT('h2)
	) name1684 (
		_w1674_,
		_w1715_,
		_w1717_
	);
	LUT2 #(
		.INIT('h1)
	) name1685 (
		_w1716_,
		_w1717_,
		_w1718_
	);
	LUT2 #(
		.INIT('h4)
	) name1686 (
		_w1673_,
		_w1718_,
		_w1719_
	);
	LUT2 #(
		.INIT('h2)
	) name1687 (
		_w1673_,
		_w1718_,
		_w1720_
	);
	LUT2 #(
		.INIT('h1)
	) name1688 (
		_w1719_,
		_w1720_,
		_w1721_
	);
	LUT2 #(
		.INIT('h4)
	) name1689 (
		_w1672_,
		_w1721_,
		_w1722_
	);
	LUT2 #(
		.INIT('h2)
	) name1690 (
		_w1672_,
		_w1721_,
		_w1723_
	);
	LUT2 #(
		.INIT('h1)
	) name1691 (
		_w1722_,
		_w1723_,
		_w1724_
	);
	LUT2 #(
		.INIT('h4)
	) name1692 (
		_w1671_,
		_w1724_,
		_w1725_
	);
	LUT2 #(
		.INIT('h2)
	) name1693 (
		_w1671_,
		_w1724_,
		_w1726_
	);
	LUT2 #(
		.INIT('h1)
	) name1694 (
		_w1725_,
		_w1726_,
		_w1727_
	);
	LUT2 #(
		.INIT('h1)
	) name1695 (
		_w1722_,
		_w1725_,
		_w1728_
	);
	LUT2 #(
		.INIT('h1)
	) name1696 (
		_w1716_,
		_w1719_,
		_w1729_
	);
	LUT2 #(
		.INIT('h8)
	) name1697 (
		\171GAT(10)_pad ,
		\528GAT(31)_pad ,
		_w1730_
	);
	LUT2 #(
		.INIT('h1)
	) name1698 (
		_w1710_,
		_w1713_,
		_w1731_
	);
	LUT2 #(
		.INIT('h8)
	) name1699 (
		\188GAT(11)_pad ,
		\511GAT(30)_pad ,
		_w1732_
	);
	LUT2 #(
		.INIT('h1)
	) name1700 (
		_w1704_,
		_w1707_,
		_w1733_
	);
	LUT2 #(
		.INIT('h8)
	) name1701 (
		\205GAT(12)_pad ,
		\494GAT(29)_pad ,
		_w1734_
	);
	LUT2 #(
		.INIT('h1)
	) name1702 (
		_w1698_,
		_w1701_,
		_w1735_
	);
	LUT2 #(
		.INIT('h8)
	) name1703 (
		\222GAT(13)_pad ,
		\477GAT(28)_pad ,
		_w1736_
	);
	LUT2 #(
		.INIT('h1)
	) name1704 (
		_w1692_,
		_w1695_,
		_w1737_
	);
	LUT2 #(
		.INIT('h8)
	) name1705 (
		\239GAT(14)_pad ,
		\460GAT(27)_pad ,
		_w1738_
	);
	LUT2 #(
		.INIT('h1)
	) name1706 (
		_w1686_,
		_w1689_,
		_w1739_
	);
	LUT2 #(
		.INIT('h8)
	) name1707 (
		\256GAT(15)_pad ,
		\443GAT(26)_pad ,
		_w1740_
	);
	LUT2 #(
		.INIT('h1)
	) name1708 (
		_w1739_,
		_w1740_,
		_w1741_
	);
	LUT2 #(
		.INIT('h8)
	) name1709 (
		_w1739_,
		_w1740_,
		_w1742_
	);
	LUT2 #(
		.INIT('h1)
	) name1710 (
		_w1741_,
		_w1742_,
		_w1743_
	);
	LUT2 #(
		.INIT('h4)
	) name1711 (
		_w1738_,
		_w1743_,
		_w1744_
	);
	LUT2 #(
		.INIT('h2)
	) name1712 (
		_w1738_,
		_w1743_,
		_w1745_
	);
	LUT2 #(
		.INIT('h1)
	) name1713 (
		_w1744_,
		_w1745_,
		_w1746_
	);
	LUT2 #(
		.INIT('h4)
	) name1714 (
		_w1737_,
		_w1746_,
		_w1747_
	);
	LUT2 #(
		.INIT('h2)
	) name1715 (
		_w1737_,
		_w1746_,
		_w1748_
	);
	LUT2 #(
		.INIT('h1)
	) name1716 (
		_w1747_,
		_w1748_,
		_w1749_
	);
	LUT2 #(
		.INIT('h4)
	) name1717 (
		_w1736_,
		_w1749_,
		_w1750_
	);
	LUT2 #(
		.INIT('h2)
	) name1718 (
		_w1736_,
		_w1749_,
		_w1751_
	);
	LUT2 #(
		.INIT('h1)
	) name1719 (
		_w1750_,
		_w1751_,
		_w1752_
	);
	LUT2 #(
		.INIT('h4)
	) name1720 (
		_w1735_,
		_w1752_,
		_w1753_
	);
	LUT2 #(
		.INIT('h2)
	) name1721 (
		_w1735_,
		_w1752_,
		_w1754_
	);
	LUT2 #(
		.INIT('h1)
	) name1722 (
		_w1753_,
		_w1754_,
		_w1755_
	);
	LUT2 #(
		.INIT('h4)
	) name1723 (
		_w1734_,
		_w1755_,
		_w1756_
	);
	LUT2 #(
		.INIT('h2)
	) name1724 (
		_w1734_,
		_w1755_,
		_w1757_
	);
	LUT2 #(
		.INIT('h1)
	) name1725 (
		_w1756_,
		_w1757_,
		_w1758_
	);
	LUT2 #(
		.INIT('h4)
	) name1726 (
		_w1733_,
		_w1758_,
		_w1759_
	);
	LUT2 #(
		.INIT('h2)
	) name1727 (
		_w1733_,
		_w1758_,
		_w1760_
	);
	LUT2 #(
		.INIT('h1)
	) name1728 (
		_w1759_,
		_w1760_,
		_w1761_
	);
	LUT2 #(
		.INIT('h4)
	) name1729 (
		_w1732_,
		_w1761_,
		_w1762_
	);
	LUT2 #(
		.INIT('h2)
	) name1730 (
		_w1732_,
		_w1761_,
		_w1763_
	);
	LUT2 #(
		.INIT('h1)
	) name1731 (
		_w1762_,
		_w1763_,
		_w1764_
	);
	LUT2 #(
		.INIT('h4)
	) name1732 (
		_w1731_,
		_w1764_,
		_w1765_
	);
	LUT2 #(
		.INIT('h2)
	) name1733 (
		_w1731_,
		_w1764_,
		_w1766_
	);
	LUT2 #(
		.INIT('h1)
	) name1734 (
		_w1765_,
		_w1766_,
		_w1767_
	);
	LUT2 #(
		.INIT('h4)
	) name1735 (
		_w1730_,
		_w1767_,
		_w1768_
	);
	LUT2 #(
		.INIT('h2)
	) name1736 (
		_w1730_,
		_w1767_,
		_w1769_
	);
	LUT2 #(
		.INIT('h1)
	) name1737 (
		_w1768_,
		_w1769_,
		_w1770_
	);
	LUT2 #(
		.INIT('h4)
	) name1738 (
		_w1729_,
		_w1770_,
		_w1771_
	);
	LUT2 #(
		.INIT('h2)
	) name1739 (
		_w1729_,
		_w1770_,
		_w1772_
	);
	LUT2 #(
		.INIT('h1)
	) name1740 (
		_w1771_,
		_w1772_,
		_w1773_
	);
	LUT2 #(
		.INIT('h4)
	) name1741 (
		_w1728_,
		_w1773_,
		_w1774_
	);
	LUT2 #(
		.INIT('h2)
	) name1742 (
		_w1728_,
		_w1773_,
		_w1775_
	);
	LUT2 #(
		.INIT('h1)
	) name1743 (
		_w1774_,
		_w1775_,
		_w1776_
	);
	LUT2 #(
		.INIT('h1)
	) name1744 (
		_w1771_,
		_w1774_,
		_w1777_
	);
	LUT2 #(
		.INIT('h1)
	) name1745 (
		_w1765_,
		_w1768_,
		_w1778_
	);
	LUT2 #(
		.INIT('h8)
	) name1746 (
		\188GAT(11)_pad ,
		\528GAT(31)_pad ,
		_w1779_
	);
	LUT2 #(
		.INIT('h1)
	) name1747 (
		_w1759_,
		_w1762_,
		_w1780_
	);
	LUT2 #(
		.INIT('h8)
	) name1748 (
		\205GAT(12)_pad ,
		\511GAT(30)_pad ,
		_w1781_
	);
	LUT2 #(
		.INIT('h1)
	) name1749 (
		_w1753_,
		_w1756_,
		_w1782_
	);
	LUT2 #(
		.INIT('h8)
	) name1750 (
		\222GAT(13)_pad ,
		\494GAT(29)_pad ,
		_w1783_
	);
	LUT2 #(
		.INIT('h1)
	) name1751 (
		_w1747_,
		_w1750_,
		_w1784_
	);
	LUT2 #(
		.INIT('h8)
	) name1752 (
		\239GAT(14)_pad ,
		\477GAT(28)_pad ,
		_w1785_
	);
	LUT2 #(
		.INIT('h1)
	) name1753 (
		_w1741_,
		_w1744_,
		_w1786_
	);
	LUT2 #(
		.INIT('h8)
	) name1754 (
		\256GAT(15)_pad ,
		\460GAT(27)_pad ,
		_w1787_
	);
	LUT2 #(
		.INIT('h1)
	) name1755 (
		_w1786_,
		_w1787_,
		_w1788_
	);
	LUT2 #(
		.INIT('h8)
	) name1756 (
		_w1786_,
		_w1787_,
		_w1789_
	);
	LUT2 #(
		.INIT('h1)
	) name1757 (
		_w1788_,
		_w1789_,
		_w1790_
	);
	LUT2 #(
		.INIT('h4)
	) name1758 (
		_w1785_,
		_w1790_,
		_w1791_
	);
	LUT2 #(
		.INIT('h2)
	) name1759 (
		_w1785_,
		_w1790_,
		_w1792_
	);
	LUT2 #(
		.INIT('h1)
	) name1760 (
		_w1791_,
		_w1792_,
		_w1793_
	);
	LUT2 #(
		.INIT('h4)
	) name1761 (
		_w1784_,
		_w1793_,
		_w1794_
	);
	LUT2 #(
		.INIT('h2)
	) name1762 (
		_w1784_,
		_w1793_,
		_w1795_
	);
	LUT2 #(
		.INIT('h1)
	) name1763 (
		_w1794_,
		_w1795_,
		_w1796_
	);
	LUT2 #(
		.INIT('h4)
	) name1764 (
		_w1783_,
		_w1796_,
		_w1797_
	);
	LUT2 #(
		.INIT('h2)
	) name1765 (
		_w1783_,
		_w1796_,
		_w1798_
	);
	LUT2 #(
		.INIT('h1)
	) name1766 (
		_w1797_,
		_w1798_,
		_w1799_
	);
	LUT2 #(
		.INIT('h4)
	) name1767 (
		_w1782_,
		_w1799_,
		_w1800_
	);
	LUT2 #(
		.INIT('h2)
	) name1768 (
		_w1782_,
		_w1799_,
		_w1801_
	);
	LUT2 #(
		.INIT('h1)
	) name1769 (
		_w1800_,
		_w1801_,
		_w1802_
	);
	LUT2 #(
		.INIT('h4)
	) name1770 (
		_w1781_,
		_w1802_,
		_w1803_
	);
	LUT2 #(
		.INIT('h2)
	) name1771 (
		_w1781_,
		_w1802_,
		_w1804_
	);
	LUT2 #(
		.INIT('h1)
	) name1772 (
		_w1803_,
		_w1804_,
		_w1805_
	);
	LUT2 #(
		.INIT('h4)
	) name1773 (
		_w1780_,
		_w1805_,
		_w1806_
	);
	LUT2 #(
		.INIT('h2)
	) name1774 (
		_w1780_,
		_w1805_,
		_w1807_
	);
	LUT2 #(
		.INIT('h1)
	) name1775 (
		_w1806_,
		_w1807_,
		_w1808_
	);
	LUT2 #(
		.INIT('h4)
	) name1776 (
		_w1779_,
		_w1808_,
		_w1809_
	);
	LUT2 #(
		.INIT('h2)
	) name1777 (
		_w1779_,
		_w1808_,
		_w1810_
	);
	LUT2 #(
		.INIT('h1)
	) name1778 (
		_w1809_,
		_w1810_,
		_w1811_
	);
	LUT2 #(
		.INIT('h4)
	) name1779 (
		_w1778_,
		_w1811_,
		_w1812_
	);
	LUT2 #(
		.INIT('h2)
	) name1780 (
		_w1778_,
		_w1811_,
		_w1813_
	);
	LUT2 #(
		.INIT('h1)
	) name1781 (
		_w1812_,
		_w1813_,
		_w1814_
	);
	LUT2 #(
		.INIT('h4)
	) name1782 (
		_w1777_,
		_w1814_,
		_w1815_
	);
	LUT2 #(
		.INIT('h2)
	) name1783 (
		_w1777_,
		_w1814_,
		_w1816_
	);
	LUT2 #(
		.INIT('h1)
	) name1784 (
		_w1815_,
		_w1816_,
		_w1817_
	);
	LUT2 #(
		.INIT('h1)
	) name1785 (
		_w1812_,
		_w1815_,
		_w1818_
	);
	LUT2 #(
		.INIT('h1)
	) name1786 (
		_w1806_,
		_w1809_,
		_w1819_
	);
	LUT2 #(
		.INIT('h8)
	) name1787 (
		\205GAT(12)_pad ,
		\528GAT(31)_pad ,
		_w1820_
	);
	LUT2 #(
		.INIT('h1)
	) name1788 (
		_w1800_,
		_w1803_,
		_w1821_
	);
	LUT2 #(
		.INIT('h8)
	) name1789 (
		\222GAT(13)_pad ,
		\511GAT(30)_pad ,
		_w1822_
	);
	LUT2 #(
		.INIT('h1)
	) name1790 (
		_w1794_,
		_w1797_,
		_w1823_
	);
	LUT2 #(
		.INIT('h8)
	) name1791 (
		\239GAT(14)_pad ,
		\494GAT(29)_pad ,
		_w1824_
	);
	LUT2 #(
		.INIT('h1)
	) name1792 (
		_w1788_,
		_w1791_,
		_w1825_
	);
	LUT2 #(
		.INIT('h8)
	) name1793 (
		\256GAT(15)_pad ,
		\477GAT(28)_pad ,
		_w1826_
	);
	LUT2 #(
		.INIT('h1)
	) name1794 (
		_w1825_,
		_w1826_,
		_w1827_
	);
	LUT2 #(
		.INIT('h8)
	) name1795 (
		_w1825_,
		_w1826_,
		_w1828_
	);
	LUT2 #(
		.INIT('h1)
	) name1796 (
		_w1827_,
		_w1828_,
		_w1829_
	);
	LUT2 #(
		.INIT('h4)
	) name1797 (
		_w1824_,
		_w1829_,
		_w1830_
	);
	LUT2 #(
		.INIT('h2)
	) name1798 (
		_w1824_,
		_w1829_,
		_w1831_
	);
	LUT2 #(
		.INIT('h1)
	) name1799 (
		_w1830_,
		_w1831_,
		_w1832_
	);
	LUT2 #(
		.INIT('h4)
	) name1800 (
		_w1823_,
		_w1832_,
		_w1833_
	);
	LUT2 #(
		.INIT('h2)
	) name1801 (
		_w1823_,
		_w1832_,
		_w1834_
	);
	LUT2 #(
		.INIT('h1)
	) name1802 (
		_w1833_,
		_w1834_,
		_w1835_
	);
	LUT2 #(
		.INIT('h4)
	) name1803 (
		_w1822_,
		_w1835_,
		_w1836_
	);
	LUT2 #(
		.INIT('h2)
	) name1804 (
		_w1822_,
		_w1835_,
		_w1837_
	);
	LUT2 #(
		.INIT('h1)
	) name1805 (
		_w1836_,
		_w1837_,
		_w1838_
	);
	LUT2 #(
		.INIT('h4)
	) name1806 (
		_w1821_,
		_w1838_,
		_w1839_
	);
	LUT2 #(
		.INIT('h2)
	) name1807 (
		_w1821_,
		_w1838_,
		_w1840_
	);
	LUT2 #(
		.INIT('h1)
	) name1808 (
		_w1839_,
		_w1840_,
		_w1841_
	);
	LUT2 #(
		.INIT('h4)
	) name1809 (
		_w1820_,
		_w1841_,
		_w1842_
	);
	LUT2 #(
		.INIT('h2)
	) name1810 (
		_w1820_,
		_w1841_,
		_w1843_
	);
	LUT2 #(
		.INIT('h1)
	) name1811 (
		_w1842_,
		_w1843_,
		_w1844_
	);
	LUT2 #(
		.INIT('h4)
	) name1812 (
		_w1819_,
		_w1844_,
		_w1845_
	);
	LUT2 #(
		.INIT('h2)
	) name1813 (
		_w1819_,
		_w1844_,
		_w1846_
	);
	LUT2 #(
		.INIT('h1)
	) name1814 (
		_w1845_,
		_w1846_,
		_w1847_
	);
	LUT2 #(
		.INIT('h4)
	) name1815 (
		_w1818_,
		_w1847_,
		_w1848_
	);
	LUT2 #(
		.INIT('h2)
	) name1816 (
		_w1818_,
		_w1847_,
		_w1849_
	);
	LUT2 #(
		.INIT('h1)
	) name1817 (
		_w1848_,
		_w1849_,
		_w1850_
	);
	LUT2 #(
		.INIT('h1)
	) name1818 (
		_w1845_,
		_w1848_,
		_w1851_
	);
	LUT2 #(
		.INIT('h1)
	) name1819 (
		_w1839_,
		_w1842_,
		_w1852_
	);
	LUT2 #(
		.INIT('h8)
	) name1820 (
		\222GAT(13)_pad ,
		\528GAT(31)_pad ,
		_w1853_
	);
	LUT2 #(
		.INIT('h1)
	) name1821 (
		_w1833_,
		_w1836_,
		_w1854_
	);
	LUT2 #(
		.INIT('h8)
	) name1822 (
		\239GAT(14)_pad ,
		\511GAT(30)_pad ,
		_w1855_
	);
	LUT2 #(
		.INIT('h1)
	) name1823 (
		_w1827_,
		_w1830_,
		_w1856_
	);
	LUT2 #(
		.INIT('h8)
	) name1824 (
		\256GAT(15)_pad ,
		\494GAT(29)_pad ,
		_w1857_
	);
	LUT2 #(
		.INIT('h1)
	) name1825 (
		_w1856_,
		_w1857_,
		_w1858_
	);
	LUT2 #(
		.INIT('h8)
	) name1826 (
		_w1856_,
		_w1857_,
		_w1859_
	);
	LUT2 #(
		.INIT('h1)
	) name1827 (
		_w1858_,
		_w1859_,
		_w1860_
	);
	LUT2 #(
		.INIT('h4)
	) name1828 (
		_w1855_,
		_w1860_,
		_w1861_
	);
	LUT2 #(
		.INIT('h2)
	) name1829 (
		_w1855_,
		_w1860_,
		_w1862_
	);
	LUT2 #(
		.INIT('h1)
	) name1830 (
		_w1861_,
		_w1862_,
		_w1863_
	);
	LUT2 #(
		.INIT('h4)
	) name1831 (
		_w1854_,
		_w1863_,
		_w1864_
	);
	LUT2 #(
		.INIT('h2)
	) name1832 (
		_w1854_,
		_w1863_,
		_w1865_
	);
	LUT2 #(
		.INIT('h1)
	) name1833 (
		_w1864_,
		_w1865_,
		_w1866_
	);
	LUT2 #(
		.INIT('h4)
	) name1834 (
		_w1853_,
		_w1866_,
		_w1867_
	);
	LUT2 #(
		.INIT('h2)
	) name1835 (
		_w1853_,
		_w1866_,
		_w1868_
	);
	LUT2 #(
		.INIT('h1)
	) name1836 (
		_w1867_,
		_w1868_,
		_w1869_
	);
	LUT2 #(
		.INIT('h4)
	) name1837 (
		_w1852_,
		_w1869_,
		_w1870_
	);
	LUT2 #(
		.INIT('h2)
	) name1838 (
		_w1852_,
		_w1869_,
		_w1871_
	);
	LUT2 #(
		.INIT('h1)
	) name1839 (
		_w1870_,
		_w1871_,
		_w1872_
	);
	LUT2 #(
		.INIT('h4)
	) name1840 (
		_w1851_,
		_w1872_,
		_w1873_
	);
	LUT2 #(
		.INIT('h2)
	) name1841 (
		_w1851_,
		_w1872_,
		_w1874_
	);
	LUT2 #(
		.INIT('h1)
	) name1842 (
		_w1873_,
		_w1874_,
		_w1875_
	);
	LUT2 #(
		.INIT('h1)
	) name1843 (
		_w1870_,
		_w1873_,
		_w1876_
	);
	LUT2 #(
		.INIT('h1)
	) name1844 (
		_w1864_,
		_w1867_,
		_w1877_
	);
	LUT2 #(
		.INIT('h8)
	) name1845 (
		\239GAT(14)_pad ,
		\528GAT(31)_pad ,
		_w1878_
	);
	LUT2 #(
		.INIT('h1)
	) name1846 (
		_w1858_,
		_w1861_,
		_w1879_
	);
	LUT2 #(
		.INIT('h8)
	) name1847 (
		\256GAT(15)_pad ,
		\511GAT(30)_pad ,
		_w1880_
	);
	LUT2 #(
		.INIT('h1)
	) name1848 (
		_w1879_,
		_w1880_,
		_w1881_
	);
	LUT2 #(
		.INIT('h8)
	) name1849 (
		_w1879_,
		_w1880_,
		_w1882_
	);
	LUT2 #(
		.INIT('h1)
	) name1850 (
		_w1881_,
		_w1882_,
		_w1883_
	);
	LUT2 #(
		.INIT('h4)
	) name1851 (
		_w1878_,
		_w1883_,
		_w1884_
	);
	LUT2 #(
		.INIT('h2)
	) name1852 (
		_w1878_,
		_w1883_,
		_w1885_
	);
	LUT2 #(
		.INIT('h1)
	) name1853 (
		_w1884_,
		_w1885_,
		_w1886_
	);
	LUT2 #(
		.INIT('h4)
	) name1854 (
		_w1877_,
		_w1886_,
		_w1887_
	);
	LUT2 #(
		.INIT('h2)
	) name1855 (
		_w1877_,
		_w1886_,
		_w1888_
	);
	LUT2 #(
		.INIT('h1)
	) name1856 (
		_w1887_,
		_w1888_,
		_w1889_
	);
	LUT2 #(
		.INIT('h4)
	) name1857 (
		_w1876_,
		_w1889_,
		_w1890_
	);
	LUT2 #(
		.INIT('h2)
	) name1858 (
		_w1876_,
		_w1889_,
		_w1891_
	);
	LUT2 #(
		.INIT('h1)
	) name1859 (
		_w1890_,
		_w1891_,
		_w1892_
	);
	LUT2 #(
		.INIT('h1)
	) name1860 (
		_w1881_,
		_w1884_,
		_w1893_
	);
	LUT2 #(
		.INIT('h8)
	) name1861 (
		\256GAT(15)_pad ,
		\528GAT(31)_pad ,
		_w1894_
	);
	LUT2 #(
		.INIT('h1)
	) name1862 (
		_w1893_,
		_w1894_,
		_w1895_
	);
	LUT2 #(
		.INIT('h1)
	) name1863 (
		_w1887_,
		_w1890_,
		_w1896_
	);
	LUT2 #(
		.INIT('h8)
	) name1864 (
		_w1893_,
		_w1894_,
		_w1897_
	);
	LUT2 #(
		.INIT('h1)
	) name1865 (
		_w1895_,
		_w1897_,
		_w1898_
	);
	LUT2 #(
		.INIT('h4)
	) name1866 (
		_w1896_,
		_w1898_,
		_w1899_
	);
	LUT2 #(
		.INIT('h1)
	) name1867 (
		_w1895_,
		_w1899_,
		_w1900_
	);
	LUT2 #(
		.INIT('h2)
	) name1868 (
		_w1896_,
		_w1898_,
		_w1901_
	);
	LUT2 #(
		.INIT('h1)
	) name1869 (
		_w1899_,
		_w1901_,
		_w1902_
	);
	assign \1581GAT(423)_pad  = _w37_ ;
	assign \1901GAT(561)_pad  = _w49_ ;
	assign \2223GAT(700)_pad  = _w69_ ;
	assign \2548GAT(840)_pad  = _w97_ ;
	assign \2877GAT(983)_pad  = _w134_ ;
	assign \3211GAT(1128)_pad  = _w177_ ;
	assign \3552GAT(1275)_pad  = _w229_ ;
	assign \3895GAT(1423)_pad  = _w289_ ;
	assign \4241GAT(1572)_pad  = _w357_ ;
	assign \4591GAT(1722)_pad  = _w433_ ;
	assign \4946GAT(1876)_pad  = _w517_ ;
	assign \5308GAT(2031)_pad  = _w609_ ;
	assign \545GAT(287)_pad  = _w610_ ;
	assign \5672GAT(2187)_pad  = _w710_ ;
	assign \5971GAT(2309)_pad  = _w818_ ;
	assign \6123GAT(2368)_pad  = _w934_ ;
	assign \6150GAT(2378)_pad  = _w1048_ ;
	assign \6160GAT(2383)_pad  = _w1160_ ;
	assign \6170GAT(2388)_pad  = _w1265_ ;
	assign \6180GAT(2393)_pad  = _w1362_ ;
	assign \6190GAT(2398)_pad  = _w1451_ ;
	assign \6200GAT(2403)_pad  = _w1532_ ;
	assign \6210GAT(2408)_pad  = _w1605_ ;
	assign \6220GAT(2413)_pad  = _w1670_ ;
	assign \6230GAT(2418)_pad  = _w1727_ ;
	assign \6240GAT(2423)_pad  = _w1776_ ;
	assign \6250GAT(2428)_pad  = _w1817_ ;
	assign \6260GAT(2433)_pad  = _w1850_ ;
	assign \6270GAT(2438)_pad  = _w1875_ ;
	assign \6280GAT(2443)_pad  = _w1892_ ;
	assign \6287GAT(2444)_pad  = _w1900_ ;
	assign \6288GAT(2447)_pad  = _w1902_ ;
endmodule;