module top( \a[0]  , \a[1]  , \a[2]  , \a[3]  , \a[4]  , \a[5]  , \a[6]  , \a[7]  , \a[8]  , \a[9]  , \a[10]  , \a[11]  , \a[12]  , \a[13]  , \a[14]  , \a[15]  , \a[16]  , \a[17]  , \a[18]  , \a[19]  , \a[20]  , \a[21]  , \a[22]  , \a[23]  , \a[24]  , \a[25]  , \a[26]  , \a[27]  , \a[28]  , \a[29]  , \a[30]  , \a[31]  , \a[32]  , \a[33]  , \a[34]  , \a[35]  , \a[36]  , \a[37]  , \a[38]  , \a[39]  , \a[40]  , \a[41]  , \a[42]  , \a[43]  , \a[44]  , \a[45]  , \a[46]  , \a[47]  , \a[48]  , \a[49]  , \a[50]  , \a[51]  , \a[52]  , \a[53]  , \a[54]  , \a[55]  , \a[56]  , \a[57]  , \a[58]  , \a[59]  , \a[60]  , \a[61]  , \a[62]  , \a[63]  , \a[64]  , \a[65]  , \a[66]  , \a[67]  , \a[68]  , \a[69]  , \a[70]  , \a[71]  , \a[72]  , \a[73]  , \a[74]  , \a[75]  , \a[76]  , \a[77]  , \a[78]  , \a[79]  , \a[80]  , \a[81]  , \a[82]  , \a[83]  , \a[84]  , \a[85]  , \a[86]  , \a[87]  , \a[88]  , \a[89]  , \a[90]  , \a[91]  , \a[92]  , \a[93]  , \a[94]  , \a[95]  , \a[96]  , \a[97]  , \a[98]  , \a[99]  , \a[100]  , \a[101]  , \a[102]  , \a[103]  , \a[104]  , \a[105]  , \a[106]  , \a[107]  , \a[108]  , \a[109]  , \a[110]  , \a[111]  , \a[112]  , \a[113]  , \a[114]  , \a[115]  , \a[116]  , \a[117]  , \a[118]  , \a[119]  , \a[120]  , \a[121]  , \a[122]  , \a[123]  , \a[124]  , \a[125]  , \a[126]  , \a[127]  , \b[0]  , \b[1]  , \b[2]  , \b[3]  , \b[4]  , \b[5]  , \b[6]  , \b[7]  , \b[8]  , \b[9]  , \b[10]  , \b[11]  , \b[12]  , \b[13]  , \b[14]  , \b[15]  , \b[16]  , \b[17]  , \b[18]  , \b[19]  , \b[20]  , \b[21]  , \b[22]  , \b[23]  , \b[24]  , \b[25]  , \b[26]  , \b[27]  , \b[28]  , \b[29]  , \b[30]  , \b[31]  , \b[32]  , \b[33]  , \b[34]  , \b[35]  , \b[36]  , \b[37]  , \b[38]  , \b[39]  , \b[40]  , \b[41]  , \b[42]  , \b[43]  , \b[44]  , \b[45]  , \b[46]  , \b[47]  , \b[48]  , \b[49]  , \b[50]  , \b[51]  , \b[52]  , \b[53]  , \b[54]  , \b[55]  , \b[56]  , \b[57]  , \b[58]  , \b[59]  , \b[60]  , \b[61]  , \b[62]  , \b[63]  , \b[64]  , \b[65]  , \b[66]  , \b[67]  , \b[68]  , \b[69]  , \b[70]  , \b[71]  , \b[72]  , \b[73]  , \b[74]  , \b[75]  , \b[76]  , \b[77]  , \b[78]  , \b[79]  , \b[80]  , \b[81]  , \b[82]  , \b[83]  , \b[84]  , \b[85]  , \b[86]  , \b[87]  , \b[88]  , \b[89]  , \b[90]  , \b[91]  , \b[92]  , \b[93]  , \b[94]  , \b[95]  , \b[96]  , \b[97]  , \b[98]  , \b[99]  , \b[100]  , \b[101]  , \b[102]  , \b[103]  , \b[104]  , \b[105]  , \b[106]  , \b[107]  , \b[108]  , \b[109]  , \b[110]  , \b[111]  , \b[112]  , \b[113]  , \b[114]  , \b[115]  , \b[116]  , \b[117]  , \b[118]  , \b[119]  , \b[120]  , \b[121]  , \b[122]  , \b[123]  , \b[124]  , \b[125]  , \b[126]  , \b[127]  , \f[0]  , \f[1]  , \f[2]  , \f[3]  , \f[4]  , \f[5]  , \f[6]  , \f[7]  , \f[8]  , \f[9]  , \f[10]  , \f[11]  , \f[12]  , \f[13]  , \f[14]  , \f[15]  , \f[16]  , \f[17]  , \f[18]  , \f[19]  , \f[20]  , \f[21]  , \f[22]  , \f[23]  , \f[24]  , \f[25]  , \f[26]  , \f[27]  , \f[28]  , \f[29]  , \f[30]  , \f[31]  , \f[32]  , \f[33]  , \f[34]  , \f[35]  , \f[36]  , \f[37]  , \f[38]  , \f[39]  , \f[40]  , \f[41]  , \f[42]  , \f[43]  , \f[44]  , \f[45]  , \f[46]  , \f[47]  , \f[48]  , \f[49]  , \f[50]  , \f[51]  , \f[52]  , \f[53]  , \f[54]  , \f[55]  , \f[56]  , \f[57]  , \f[58]  , \f[59]  , \f[60]  , \f[61]  , \f[62]  , \f[63]  , \f[64]  , \f[65]  , \f[66]  , \f[67]  , \f[68]  , \f[69]  , \f[70]  , \f[71]  , \f[72]  , \f[73]  , \f[74]  , \f[75]  , \f[76]  , \f[77]  , \f[78]  , \f[79]  , \f[80]  , \f[81]  , \f[82]  , \f[83]  , \f[84]  , \f[85]  , \f[86]  , \f[87]  , \f[88]  , \f[89]  , \f[90]  , \f[91]  , \f[92]  , \f[93]  , \f[94]  , \f[95]  , \f[96]  , \f[97]  , \f[98]  , \f[99]  , \f[100]  , \f[101]  , \f[102]  , \f[103]  , \f[104]  , \f[105]  , \f[106]  , \f[107]  , \f[108]  , \f[109]  , \f[110]  , \f[111]  , \f[112]  , \f[113]  , \f[114]  , \f[115]  , \f[116]  , \f[117]  , \f[118]  , \f[119]  , \f[120]  , \f[121]  , \f[122]  , \f[123]  , \f[124]  , \f[125]  , \f[126]  , \f[127]  , cOut );
  input \a[0]  ;
  input \a[1]  ;
  input \a[2]  ;
  input \a[3]  ;
  input \a[4]  ;
  input \a[5]  ;
  input \a[6]  ;
  input \a[7]  ;
  input \a[8]  ;
  input \a[9]  ;
  input \a[10]  ;
  input \a[11]  ;
  input \a[12]  ;
  input \a[13]  ;
  input \a[14]  ;
  input \a[15]  ;
  input \a[16]  ;
  input \a[17]  ;
  input \a[18]  ;
  input \a[19]  ;
  input \a[20]  ;
  input \a[21]  ;
  input \a[22]  ;
  input \a[23]  ;
  input \a[24]  ;
  input \a[25]  ;
  input \a[26]  ;
  input \a[27]  ;
  input \a[28]  ;
  input \a[29]  ;
  input \a[30]  ;
  input \a[31]  ;
  input \a[32]  ;
  input \a[33]  ;
  input \a[34]  ;
  input \a[35]  ;
  input \a[36]  ;
  input \a[37]  ;
  input \a[38]  ;
  input \a[39]  ;
  input \a[40]  ;
  input \a[41]  ;
  input \a[42]  ;
  input \a[43]  ;
  input \a[44]  ;
  input \a[45]  ;
  input \a[46]  ;
  input \a[47]  ;
  input \a[48]  ;
  input \a[49]  ;
  input \a[50]  ;
  input \a[51]  ;
  input \a[52]  ;
  input \a[53]  ;
  input \a[54]  ;
  input \a[55]  ;
  input \a[56]  ;
  input \a[57]  ;
  input \a[58]  ;
  input \a[59]  ;
  input \a[60]  ;
  input \a[61]  ;
  input \a[62]  ;
  input \a[63]  ;
  input \a[64]  ;
  input \a[65]  ;
  input \a[66]  ;
  input \a[67]  ;
  input \a[68]  ;
  input \a[69]  ;
  input \a[70]  ;
  input \a[71]  ;
  input \a[72]  ;
  input \a[73]  ;
  input \a[74]  ;
  input \a[75]  ;
  input \a[76]  ;
  input \a[77]  ;
  input \a[78]  ;
  input \a[79]  ;
  input \a[80]  ;
  input \a[81]  ;
  input \a[82]  ;
  input \a[83]  ;
  input \a[84]  ;
  input \a[85]  ;
  input \a[86]  ;
  input \a[87]  ;
  input \a[88]  ;
  input \a[89]  ;
  input \a[90]  ;
  input \a[91]  ;
  input \a[92]  ;
  input \a[93]  ;
  input \a[94]  ;
  input \a[95]  ;
  input \a[96]  ;
  input \a[97]  ;
  input \a[98]  ;
  input \a[99]  ;
  input \a[100]  ;
  input \a[101]  ;
  input \a[102]  ;
  input \a[103]  ;
  input \a[104]  ;
  input \a[105]  ;
  input \a[106]  ;
  input \a[107]  ;
  input \a[108]  ;
  input \a[109]  ;
  input \a[110]  ;
  input \a[111]  ;
  input \a[112]  ;
  input \a[113]  ;
  input \a[114]  ;
  input \a[115]  ;
  input \a[116]  ;
  input \a[117]  ;
  input \a[118]  ;
  input \a[119]  ;
  input \a[120]  ;
  input \a[121]  ;
  input \a[122]  ;
  input \a[123]  ;
  input \a[124]  ;
  input \a[125]  ;
  input \a[126]  ;
  input \a[127]  ;
  input \b[0]  ;
  input \b[1]  ;
  input \b[2]  ;
  input \b[3]  ;
  input \b[4]  ;
  input \b[5]  ;
  input \b[6]  ;
  input \b[7]  ;
  input \b[8]  ;
  input \b[9]  ;
  input \b[10]  ;
  input \b[11]  ;
  input \b[12]  ;
  input \b[13]  ;
  input \b[14]  ;
  input \b[15]  ;
  input \b[16]  ;
  input \b[17]  ;
  input \b[18]  ;
  input \b[19]  ;
  input \b[20]  ;
  input \b[21]  ;
  input \b[22]  ;
  input \b[23]  ;
  input \b[24]  ;
  input \b[25]  ;
  input \b[26]  ;
  input \b[27]  ;
  input \b[28]  ;
  input \b[29]  ;
  input \b[30]  ;
  input \b[31]  ;
  input \b[32]  ;
  input \b[33]  ;
  input \b[34]  ;
  input \b[35]  ;
  input \b[36]  ;
  input \b[37]  ;
  input \b[38]  ;
  input \b[39]  ;
  input \b[40]  ;
  input \b[41]  ;
  input \b[42]  ;
  input \b[43]  ;
  input \b[44]  ;
  input \b[45]  ;
  input \b[46]  ;
  input \b[47]  ;
  input \b[48]  ;
  input \b[49]  ;
  input \b[50]  ;
  input \b[51]  ;
  input \b[52]  ;
  input \b[53]  ;
  input \b[54]  ;
  input \b[55]  ;
  input \b[56]  ;
  input \b[57]  ;
  input \b[58]  ;
  input \b[59]  ;
  input \b[60]  ;
  input \b[61]  ;
  input \b[62]  ;
  input \b[63]  ;
  input \b[64]  ;
  input \b[65]  ;
  input \b[66]  ;
  input \b[67]  ;
  input \b[68]  ;
  input \b[69]  ;
  input \b[70]  ;
  input \b[71]  ;
  input \b[72]  ;
  input \b[73]  ;
  input \b[74]  ;
  input \b[75]  ;
  input \b[76]  ;
  input \b[77]  ;
  input \b[78]  ;
  input \b[79]  ;
  input \b[80]  ;
  input \b[81]  ;
  input \b[82]  ;
  input \b[83]  ;
  input \b[84]  ;
  input \b[85]  ;
  input \b[86]  ;
  input \b[87]  ;
  input \b[88]  ;
  input \b[89]  ;
  input \b[90]  ;
  input \b[91]  ;
  input \b[92]  ;
  input \b[93]  ;
  input \b[94]  ;
  input \b[95]  ;
  input \b[96]  ;
  input \b[97]  ;
  input \b[98]  ;
  input \b[99]  ;
  input \b[100]  ;
  input \b[101]  ;
  input \b[102]  ;
  input \b[103]  ;
  input \b[104]  ;
  input \b[105]  ;
  input \b[106]  ;
  input \b[107]  ;
  input \b[108]  ;
  input \b[109]  ;
  input \b[110]  ;
  input \b[111]  ;
  input \b[112]  ;
  input \b[113]  ;
  input \b[114]  ;
  input \b[115]  ;
  input \b[116]  ;
  input \b[117]  ;
  input \b[118]  ;
  input \b[119]  ;
  input \b[120]  ;
  input \b[121]  ;
  input \b[122]  ;
  input \b[123]  ;
  input \b[124]  ;
  input \b[125]  ;
  input \b[126]  ;
  input \b[127]  ;
  output \f[0]  ;
  output \f[1]  ;
  output \f[2]  ;
  output \f[3]  ;
  output \f[4]  ;
  output \f[5]  ;
  output \f[6]  ;
  output \f[7]  ;
  output \f[8]  ;
  output \f[9]  ;
  output \f[10]  ;
  output \f[11]  ;
  output \f[12]  ;
  output \f[13]  ;
  output \f[14]  ;
  output \f[15]  ;
  output \f[16]  ;
  output \f[17]  ;
  output \f[18]  ;
  output \f[19]  ;
  output \f[20]  ;
  output \f[21]  ;
  output \f[22]  ;
  output \f[23]  ;
  output \f[24]  ;
  output \f[25]  ;
  output \f[26]  ;
  output \f[27]  ;
  output \f[28]  ;
  output \f[29]  ;
  output \f[30]  ;
  output \f[31]  ;
  output \f[32]  ;
  output \f[33]  ;
  output \f[34]  ;
  output \f[35]  ;
  output \f[36]  ;
  output \f[37]  ;
  output \f[38]  ;
  output \f[39]  ;
  output \f[40]  ;
  output \f[41]  ;
  output \f[42]  ;
  output \f[43]  ;
  output \f[44]  ;
  output \f[45]  ;
  output \f[46]  ;
  output \f[47]  ;
  output \f[48]  ;
  output \f[49]  ;
  output \f[50]  ;
  output \f[51]  ;
  output \f[52]  ;
  output \f[53]  ;
  output \f[54]  ;
  output \f[55]  ;
  output \f[56]  ;
  output \f[57]  ;
  output \f[58]  ;
  output \f[59]  ;
  output \f[60]  ;
  output \f[61]  ;
  output \f[62]  ;
  output \f[63]  ;
  output \f[64]  ;
  output \f[65]  ;
  output \f[66]  ;
  output \f[67]  ;
  output \f[68]  ;
  output \f[69]  ;
  output \f[70]  ;
  output \f[71]  ;
  output \f[72]  ;
  output \f[73]  ;
  output \f[74]  ;
  output \f[75]  ;
  output \f[76]  ;
  output \f[77]  ;
  output \f[78]  ;
  output \f[79]  ;
  output \f[80]  ;
  output \f[81]  ;
  output \f[82]  ;
  output \f[83]  ;
  output \f[84]  ;
  output \f[85]  ;
  output \f[86]  ;
  output \f[87]  ;
  output \f[88]  ;
  output \f[89]  ;
  output \f[90]  ;
  output \f[91]  ;
  output \f[92]  ;
  output \f[93]  ;
  output \f[94]  ;
  output \f[95]  ;
  output \f[96]  ;
  output \f[97]  ;
  output \f[98]  ;
  output \f[99]  ;
  output \f[100]  ;
  output \f[101]  ;
  output \f[102]  ;
  output \f[103]  ;
  output \f[104]  ;
  output \f[105]  ;
  output \f[106]  ;
  output \f[107]  ;
  output \f[108]  ;
  output \f[109]  ;
  output \f[110]  ;
  output \f[111]  ;
  output \f[112]  ;
  output \f[113]  ;
  output \f[114]  ;
  output \f[115]  ;
  output \f[116]  ;
  output \f[117]  ;
  output \f[118]  ;
  output \f[119]  ;
  output \f[120]  ;
  output \f[121]  ;
  output \f[122]  ;
  output \f[123]  ;
  output \f[124]  ;
  output \f[125]  ;
  output \f[126]  ;
  output \f[127]  ;
  output cOut ;
  wire n257 , n258 , n259 , n260 , n261 , n262 , n263 , n264 , n265 , n266 , n267 , n268 , n269 , n270 , n271 , n272 , n273 , n274 , n275 , n276 , n277 , n278 , n279 , n280 , n281 , n282 , n283 , n284 , n285 , n286 , n287 , n288 , n289 , n290 , n291 , n292 , n293 , n294 , n295 , n296 , n297 , n298 , n299 , n300 , n301 , n302 , n303 , n304 , n305 , n306 , n307 , n308 , n309 , n310 , n311 , n312 , n313 , n314 , n315 , n316 , n317 , n318 , n319 , n320 , n321 , n322 , n323 , n324 , n325 , n326 , n327 , n328 , n329 , n330 , n331 , n332 , n333 , n334 , n335 , n336 , n337 , n338 , n339 , n340 , n341 , n342 , n343 , n344 , n345 , n346 , n347 , n348 , n349 , n350 , n351 , n352 , n353 , n354 , n355 , n356 , n357 , n358 , n359 , n360 , n361 , n362 , n363 , n364 , n365 , n366 , n367 , n368 , n369 , n370 , n371 , n372 , n373 , n374 , n375 , n376 , n377 , n378 , n379 , n380 , n381 , n382 , n383 , n384 , n385 , n386 , n387 , n388 , n389 , n390 , n391 , n392 , n393 , n394 , n395 , n396 , n397 , n398 , n399 , n400 , n401 , n402 , n403 , n404 , n405 , n406 , n407 , n408 , n409 , n410 , n411 , n412 , n413 , n414 , n415 , n416 , n417 , n418 , n419 , n420 , n421 , n422 , n423 , n424 , n425 , n426 , n427 , n428 , n429 , n430 , n431 , n432 , n433 , n434 , n435 , n436 , n437 , n438 , n439 , n440 , n441 , n442 , n443 , n444 , n445 , n446 , n447 , n448 , n449 , n450 , n451 , n452 , n453 , n454 , n455 , n456 , n457 , n458 , n459 , n460 , n461 , n462 , n463 , n464 , n465 , n466 , n467 , n468 , n469 , n470 , n471 , n472 , n473 , n474 , n475 , n476 , n477 , n478 , n479 , n480 , n481 , n482 , n483 , n484 , n485 , n486 , n487 , n488 , n489 , n490 , n491 , n492 , n493 , n494 , n495 , n496 , n497 , n498 , n499 , n500 , n501 , n502 , n503 , n504 , n505 , n506 , n507 , n508 , n509 , n510 , n511 , n512 , n513 , n514 , n515 , n516 , n517 , n518 , n519 , n520 , n521 , n522 , n523 , n524 , n525 , n526 , n527 , n528 , n529 , n530 , n531 , n532 , n533 , n534 , n535 , n536 , n537 , n538 , n539 , n540 , n541 , n542 , n543 , n544 , n545 , n546 , n547 , n548 , n549 , n550 , n551 , n552 , n553 , n554 , n555 , n556 , n557 , n558 , n559 , n560 , n561 , n562 , n563 , n564 , n565 , n566 , n567 , n568 , n569 , n570 , n571 , n572 , n573 , n574 , n575 , n576 , n577 , n578 , n579 , n580 , n581 , n582 , n583 , n584 , n585 , n586 , n587 , n588 , n589 , n590 , n591 , n592 , n593 , n594 , n595 , n596 , n597 , n598 , n599 , n600 , n601 , n602 , n603 , n604 , n605 , n606 , n607 , n608 , n609 , n610 , n611 , n612 , n613 , n614 , n615 , n616 , n617 , n618 , n619 , n620 , n621 , n622 , n623 , n624 , n625 , n626 , n627 , n628 , n629 , n630 , n631 , n632 , n633 , n634 , n635 , n636 , n637 , n638 , n639 , n640 , n641 , n642 , n643 , n644 , n645 , n646 , n647 , n648 , n649 , n650 , n651 , n652 , n653 , n654 , n655 , n656 , n657 , n658 , n659 , n660 , n661 , n662 , n663 , n664 , n665 , n666 , n667 , n668 , n669 , n670 , n671 , n672 , n673 , n674 , n675 , n676 , n677 , n678 , n679 , n680 , n681 , n682 , n683 , n684 , n685 , n686 , n687 , n688 , n689 , n690 , n691 , n692 , n693 , n694 , n695 , n696 , n697 , n698 , n699 , n700 , n701 , n702 , n703 , n704 , n705 , n706 , n707 , n708 , n709 , n710 , n711 , n712 , n713 , n714 , n715 , n716 , n717 , n718 , n719 , n720 , n721 , n722 , n723 , n724 , n725 , n726 , n727 , n728 , n729 , n730 , n731 , n732 , n733 , n734 , n735 , n736 , n737 , n738 , n739 , n740 , n741 , n742 , n743 , n744 , n745 , n746 , n747 , n748 , n749 , n750 , n751 , n752 , n753 , n754 , n755 , n756 , n757 , n758 , n759 , n760 , n761 , n762 , n763 , n764 , n765 , n766 , n767 , n768 , n769 , n770 , n771 , n772 , n773 , n774 , n775 , n776 , n777 , n778 , n779 , n780 , n781 , n782 , n783 , n784 , n785 , n786 , n787 , n788 , n789 , n790 , n791 , n792 , n793 , n794 , n795 , n796 , n797 , n798 , n799 , n800 , n801 , n802 , n803 , n804 , n805 , n806 , n807 , n808 , n809 , n810 , n811 , n812 , n813 , n814 , n815 , n816 , n817 , n818 , n819 , n820 , n821 , n822 , n823 , n824 , n825 , n826 , n827 , n828 , n829 , n830 , n831 , n832 , n833 , n834 , n835 , n836 , n837 , n838 , n839 , n840 , n841 , n842 , n843 , n844 , n845 , n846 , n847 , n848 , n849 , n850 , n851 , n852 , n853 , n854 , n855 , n856 , n857 , n858 , n859 , n860 , n861 , n862 , n863 , n864 , n865 , n866 , n867 , n868 , n869 , n870 , n871 , n872 , n873 , n874 , n875 , n876 , n877 , n878 , n879 , n880 , n881 , n882 , n883 , n884 , n885 , n886 , n887 , n888 , n889 , n890 , n891 , n892 , n893 , n894 , n895 , n896 , n897 , n898 , n899 , n900 , n901 , n902 , n903 , n904 , n905 , n906 , n907 , n908 , n909 , n910 , n911 , n912 , n913 , n914 , n915 , n916 , n917 , n918 , n919 , n920 , n921 , n922 , n923 , n924 , n925 , n926 , n927 , n928 , n929 , n930 , n931 , n932 , n933 , n934 , n935 , n936 , n937 , n938 , n939 , n940 , n941 , n942 , n943 , n944 , n945 , n946 , n947 , n948 , n949 , n950 , n951 , n952 , n953 , n954 , n955 , n956 , n957 , n958 , n959 , n960 , n961 , n962 , n963 , n964 , n965 , n966 , n967 , n968 , n969 , n970 , n971 , n972 , n973 , n974 , n975 , n976 , n977 , n978 , n979 , n980 , n981 , n982 , n983 , n984 , n985 , n986 , n987 , n988 , n989 , n990 , n991 , n992 , n993 , n994 , n995 , n996 , n997 , n998 , n999 , n1000 , n1001 , n1002 , n1003 , n1004 , n1005 , n1006 , n1007 , n1008 , n1009 , n1010 , n1011 , n1012 , n1013 , n1014 , n1015 , n1016 , n1017 , n1018 , n1019 , n1020 , n1021 , n1022 , n1023 , n1024 , n1025 , n1026 , n1027 , n1028 , n1029 , n1030 , n1031 , n1032 , n1033 , n1034 , n1035 , n1036 , n1037 , n1038 , n1039 , n1040 , n1041 , n1042 , n1043 , n1044 , n1045 , n1046 , n1047 , n1048 , n1049 , n1050 , n1051 , n1052 , n1053 , n1054 , n1055 , n1056 , n1057 , n1058 , n1059 , n1060 , n1061 , n1062 , n1063 , n1064 , n1065 , n1066 , n1067 , n1068 , n1069 , n1070 , n1071 , n1072 , n1073 , n1074 , n1075 , n1076 , n1077 , n1078 , n1079 , n1080 , n1081 , n1082 , n1083 , n1084 , n1085 , n1086 , n1087 , n1088 , n1089 , n1090 , n1091 , n1092 , n1093 , n1094 , n1095 , n1096 , n1097 , n1098 , n1099 , n1100 , n1101 , n1102 , n1103 , n1104 , n1105 , n1106 , n1107 , n1108 , n1109 , n1110 , n1111 , n1112 , n1113 , n1114 , n1115 , n1116 , n1117 , n1118 , n1119 , n1120 , n1121 , n1122 , n1123 , n1124 , n1125 , n1126 , n1127 , n1128 , n1129 , n1130 , n1131 , n1132 , n1133 , n1134 , n1135 , n1136 , n1137 , n1138 , n1139 , n1140 , n1141 , n1142 , n1143 , n1144 , n1145 , n1146 , n1147 , n1148 , n1149 , n1150 , n1151 , n1152 , n1153 , n1154 , n1155 , n1156 , n1157 , n1158 , n1159 , n1160 , n1161 , n1162 , n1163 , n1164 , n1165 , n1166 , n1167 , n1168 , n1169 , n1170 , n1171 , n1172 , n1173 , n1174 , n1175 , n1176 , n1177 , n1178 , n1179 , n1180 , n1181 , n1182 , n1183 , n1184 , n1185 , n1186 , n1187 , n1188 , n1189 , n1190 , n1191 , n1192 , n1193 , n1194 , n1195 , n1196 , n1197 , n1198 , n1199 , n1200 , n1201 , n1202 , n1203 , n1204 , n1205 , n1206 , n1207 , n1208 , n1209 , n1210 , n1211 , n1212 , n1213 , n1214 , n1215 , n1216 , n1217 , n1218 , n1219 , n1220 , n1221 , n1222 , n1223 , n1224 , n1225 , n1226 , n1227 , n1228 , n1229 , n1230 , n1231 , n1232 , n1233 , n1234 , n1235 , n1236 , n1237 , n1238 , n1239 , n1240 , n1241 , n1242 , n1243 , n1244 , n1245 , n1246 , n1247 , n1248 , n1249 , n1250 , n1251 , n1252 , n1253 , n1254 , n1255 , n1256 , n1257 , n1258 , n1259 , n1260 , n1261 , n1262 , n1263 , n1264 , n1265 , n1266 , n1267 , n1268 , n1269 , n1270 , n1271 , n1272 , n1273 , n1274 , n1275 , n1276 , n1277 , n1278 , n1279 , n1280 , n1281 , n1282 , n1283 , n1284 , n1285 , n1286 , n1287 , n1288 , n1289 , n1290 , n1291 , n1292 , n1293 , n1294 , n1295 , n1296 , n1297 , n1298 , n1299 , n1300 , n1301 , n1302 , n1303 , n1304 , n1305 , n1306 , n1307 , n1308 , n1309 , n1310 , n1311 , n1312 , n1313 , n1314 , n1315 , n1316 , n1317 , n1318 , n1319 , n1320 , n1321 , n1322 , n1323 , n1324 , n1325 , n1326 , n1327 , n1328 , n1329 , n1330 , n1331 , n1332 , n1333 , n1334 , n1335 , n1336 , n1337 , n1338 , n1339 , n1340 , n1341 , n1342 , n1343 , n1344 , n1345 , n1346 , n1347 , n1348 , n1349 , n1350 , n1351 , n1352 , n1353 , n1354 , n1355 , n1356 , n1357 , n1358 , n1359 , n1360 , n1361 , n1362 , n1363 , n1364 , n1365 , n1366 , n1367 , n1368 , n1369 , n1370 , n1371 , n1372 , n1373 , n1374 , n1375 , n1376 , n1377 , n1378 , n1379 , n1380 , n1381 , n1382 , n1383 , n1384 , n1385 , n1386 , n1387 , n1388 , n1389 , n1390 , n1391 , n1392 , n1393 , n1394 , n1395 , n1396 , n1397 , n1398 , n1399 , n1400 , n1401 , n1402 , n1403 , n1404 , n1405 , n1406 , n1407 , n1408 , n1409 , n1410 , n1411 , n1412 , n1413 , n1414 , n1415 , n1416 , n1417 , n1418 , n1419 , n1420 , n1421 , n1422 , n1423 , n1424 , n1425 , n1426 , n1427 , n1428 , n1429 , n1430 , n1431 , n1432 , n1433 , n1434 , n1435 , n1436 , n1437 , n1438 , n1439 , n1440 , n1441 , n1442 , n1443 , n1444 , n1445 , n1446 , n1447 , n1448 , n1449 , n1450 , n1451 , n1452 , n1453 , n1454 , n1455 , n1456 , n1457 , n1458 , n1459 , n1460 , n1461 , n1462 , n1463 , n1464 , n1465 , n1466 , n1467 , n1468 , n1469 , n1470 , n1471 , n1472 , n1473 , n1474 , n1475 , n1476 , n1477 , n1478 , n1479 , n1480 , n1481 , n1482 , n1483 , n1484 , n1485 , n1486 , n1487 , n1488 , n1489 , n1490 , n1491 , n1492 , n1493 , n1494 , n1495 , n1496 , n1497 , n1498 , n1499 , n1500 , n1501 , n1502 , n1503 , n1504 , n1505 , n1506 , n1507 , n1508 , n1509 , n1510 , n1511 , n1512 , n1513 , n1514 , n1515 , n1516 , n1517 , n1518 , n1519 , n1520 , n1521 , n1522 , n1523 , n1524 , n1525 , n1526 , n1527 , n1528 , n1529 , n1530 , n1531 , n1532 , n1533 , n1534 , n1535 , n1536 , n1537 , n1538 , n1539 , n1540 , n1541 , n1542 , n1543 , n1544 , n1545 , n1546 , n1547 , n1548 , n1549 , n1550 , n1551 , n1552 , n1553 , n1554 , n1555 , n1556 , n1557 , n1558 , n1559 , n1560 , n1561 , n1562 , n1563 , n1564 , n1565 , n1566 , n1567 , n1568 , n1569 , n1570 , n1571 , n1572 , n1573 , n1574 , n1575 , n1576 , n1577 , n1578 , n1579 , n1580 , n1581 , n1582 , n1583 , n1584 , n1585 , n1586 , n1587 , n1588 , n1589 , n1590 , n1591 , n1592 , n1593 , n1594 , n1595 , n1596 , n1597 , n1598 , n1599 , n1600 , n1601 , n1602 , n1603 , n1604 , n1605 , n1606 , n1607 , n1608 , n1609 , n1610 , n1611 , n1612 , n1613 , n1614 , n1615 , n1616 , n1617 , n1618 , n1619 , n1620 , n1621 , n1622 , n1623 , n1624 , n1625 , n1626 , n1627 , n1628 , n1629 , n1630 , n1631 , n1632 , n1633 , n1634 , n1635 , n1636 , n1637 , n1638 , n1639 , n1640 , n1641 , n1642 , n1643 , n1644 , n1645 , n1646 , n1647 , n1648 , n1649 , n1650 , n1651 , n1652 , n1653 , n1654 , n1655 , n1656 , n1657 , n1658 , n1659 , n1660 , n1661 , n1662 , n1663 , n1664 , n1665 , n1666 , n1667 , n1668 , n1669 , n1670 , n1671 , n1672 , n1673 , n1674 , n1675 , n1676 , n1677 , n1678 , n1679 , n1680 , n1681 , n1682 , n1683 , n1684 , n1685 , n1686 , n1687 , n1688 , n1689 , n1690 , n1691 , n1692 , n1693 , n1694 , n1695 , n1696 , n1697 , n1698 , n1699 , n1700 , n1701 , n1702 , n1703 , n1704 , n1705 , n1706 , n1707 , n1708 , n1709 , n1710 , n1711 , n1712 , n1713 , n1714 , n1715 , n1716 , n1717 , n1718 , n1719 , n1720 , n1721 , n1722 , n1723 , n1724 , n1725 , n1726 , n1727 , n1728 , n1729 , n1730 , n1731 , n1732 , n1733 , n1734 , n1735 , n1736 , n1737 , n1738 , n1739 , n1740 , n1741 , n1742 , n1743 , n1744 , n1745 , n1746 , n1747 , n1748 , n1749 , n1750 , n1751 , n1752 , n1753 , n1754 , n1755 , n1756 , n1757 , n1758 , n1759 , n1760 , n1761 , n1762 , n1763 , n1764 , n1765 , n1766 , n1767 , n1768 , n1769 , n1770 , n1771 , n1772 , n1773 , n1774 ;
  assign n257 = \a[0]  & \b[0]  ;
  assign n258 = ~\a[0]  & ~\b[0]  ;
  assign n259 = ~n257 & ~n258 ;
  assign n260 = ~\a[1]  & ~\b[1]  ;
  assign n261 = \a[1]  & \b[1]  ;
  assign n262 = ~n260 & ~n261 ;
  assign n263 = ~n257 & ~n262 ;
  assign n264 = n257 & n262 ;
  assign n265 = ~n263 & ~n264 ;
  assign n266 = ~\a[2]  & ~\b[2]  ;
  assign n267 = \a[2]  & \b[2]  ;
  assign n268 = ~n266 & ~n267 ;
  assign n269 = ~n257 & ~n261 ;
  assign n270 = ~n260 & ~n269 ;
  assign n271 = ~n268 & ~n270 ;
  assign n272 = n268 & n270 ;
  assign n273 = ~n271 & ~n272 ;
  assign n274 = ~\a[3]  & ~\b[3]  ;
  assign n275 = \a[3]  & \b[3]  ;
  assign n276 = ~n274 & ~n275 ;
  assign n277 = ~n260 & ~n266 ;
  assign n278 = ~n269 & n277 ;
  assign n279 = ~n267 & ~n278 ;
  assign n280 = ~n276 & ~n279 ;
  assign n281 = ~n267 & n276 ;
  assign n282 = ~n278 & n281 ;
  assign n283 = ~n280 & ~n282 ;
  assign n284 = ~n267 & ~n275 ;
  assign n285 = ~n278 & n284 ;
  assign n286 = ~\a[4]  & ~\b[4]  ;
  assign n287 = \a[4]  & \b[4]  ;
  assign n288 = ~n286 & ~n287 ;
  assign n289 = ~n274 & ~n288 ;
  assign n290 = ~n285 & n289 ;
  assign n291 = n274 & n288 ;
  assign n292 = n284 & n288 ;
  assign n293 = ~n278 & n292 ;
  assign n294 = ~n291 & ~n293 ;
  assign n295 = ~n290 & n294 ;
  assign n296 = n284 & ~n287 ;
  assign n297 = ~n278 & n296 ;
  assign n298 = n274 & ~n287 ;
  assign n299 = ~\a[5]  & ~\b[5]  ;
  assign n300 = \a[5]  & \b[5]  ;
  assign n301 = ~n299 & ~n300 ;
  assign n302 = ~n286 & ~n301 ;
  assign n303 = ~n298 & n302 ;
  assign n304 = ~n297 & n303 ;
  assign n305 = ~n286 & ~n298 ;
  assign n306 = ~n297 & n305 ;
  assign n307 = n301 & ~n306 ;
  assign n308 = ~n304 & ~n307 ;
  assign n309 = ~\a[6]  & ~\b[6]  ;
  assign n310 = \a[6]  & \b[6]  ;
  assign n311 = ~n309 & ~n310 ;
  assign n312 = ~n286 & ~n299 ;
  assign n313 = ~n298 & n312 ;
  assign n314 = ~n297 & n313 ;
  assign n315 = ~n300 & ~n314 ;
  assign n316 = ~n311 & ~n315 ;
  assign n317 = ~n300 & n311 ;
  assign n318 = ~n314 & n317 ;
  assign n319 = ~n316 & ~n318 ;
  assign n320 = ~n300 & ~n310 ;
  assign n321 = ~n314 & n320 ;
  assign n322 = ~\a[7]  & ~\b[7]  ;
  assign n323 = \a[7]  & \b[7]  ;
  assign n324 = ~n322 & ~n323 ;
  assign n325 = ~n309 & ~n324 ;
  assign n326 = ~n321 & n325 ;
  assign n327 = n309 & n324 ;
  assign n328 = n320 & n324 ;
  assign n329 = ~n314 & n328 ;
  assign n330 = ~n327 & ~n329 ;
  assign n331 = ~n326 & n330 ;
  assign n332 = n320 & ~n323 ;
  assign n333 = ~n314 & n332 ;
  assign n334 = n309 & ~n323 ;
  assign n335 = ~\a[8]  & ~\b[8]  ;
  assign n336 = \a[8]  & \b[8]  ;
  assign n337 = ~n335 & ~n336 ;
  assign n338 = ~n322 & ~n337 ;
  assign n339 = ~n334 & n338 ;
  assign n340 = ~n333 & n339 ;
  assign n341 = ~n322 & ~n334 ;
  assign n342 = ~n333 & n341 ;
  assign n343 = n337 & ~n342 ;
  assign n344 = ~n340 & ~n343 ;
  assign n345 = ~\a[9]  & ~\b[9]  ;
  assign n346 = \a[9]  & \b[9]  ;
  assign n347 = ~n345 & ~n346 ;
  assign n348 = ~n322 & ~n335 ;
  assign n349 = ~n334 & n348 ;
  assign n350 = ~n333 & n349 ;
  assign n351 = ~n336 & ~n350 ;
  assign n352 = ~n347 & ~n351 ;
  assign n353 = ~n336 & n347 ;
  assign n354 = ~n350 & n353 ;
  assign n355 = ~n352 & ~n354 ;
  assign n356 = ~n336 & ~n346 ;
  assign n357 = ~n350 & n356 ;
  assign n358 = ~\a[10]  & ~\b[10]  ;
  assign n359 = \a[10]  & \b[10]  ;
  assign n360 = ~n358 & ~n359 ;
  assign n361 = ~n345 & ~n360 ;
  assign n362 = ~n357 & n361 ;
  assign n363 = n345 & n360 ;
  assign n364 = n356 & n360 ;
  assign n365 = ~n350 & n364 ;
  assign n366 = ~n363 & ~n365 ;
  assign n367 = ~n362 & n366 ;
  assign n368 = n356 & ~n359 ;
  assign n369 = ~n350 & n368 ;
  assign n370 = n345 & ~n359 ;
  assign n371 = ~\a[11]  & ~\b[11]  ;
  assign n372 = \a[11]  & \b[11]  ;
  assign n373 = ~n371 & ~n372 ;
  assign n374 = ~n358 & ~n373 ;
  assign n375 = ~n370 & n374 ;
  assign n376 = ~n369 & n375 ;
  assign n377 = ~n358 & ~n370 ;
  assign n378 = ~n369 & n377 ;
  assign n379 = n373 & ~n378 ;
  assign n380 = ~n376 & ~n379 ;
  assign n381 = ~\a[12]  & ~\b[12]  ;
  assign n382 = \a[12]  & \b[12]  ;
  assign n383 = ~n381 & ~n382 ;
  assign n384 = ~n358 & ~n371 ;
  assign n385 = ~n370 & n384 ;
  assign n386 = ~n369 & n385 ;
  assign n387 = ~n372 & ~n386 ;
  assign n388 = ~n383 & ~n387 ;
  assign n389 = ~n372 & n383 ;
  assign n390 = ~n386 & n389 ;
  assign n391 = ~n388 & ~n390 ;
  assign n392 = ~n372 & ~n382 ;
  assign n393 = ~n386 & n392 ;
  assign n394 = ~\a[13]  & ~\b[13]  ;
  assign n395 = \a[13]  & \b[13]  ;
  assign n396 = ~n394 & ~n395 ;
  assign n397 = ~n381 & ~n396 ;
  assign n398 = ~n393 & n397 ;
  assign n399 = n381 & n396 ;
  assign n400 = n392 & n396 ;
  assign n401 = ~n386 & n400 ;
  assign n402 = ~n399 & ~n401 ;
  assign n403 = ~n398 & n402 ;
  assign n404 = n392 & ~n395 ;
  assign n405 = ~n386 & n404 ;
  assign n406 = n381 & ~n395 ;
  assign n407 = ~\a[14]  & ~\b[14]  ;
  assign n408 = \a[14]  & \b[14]  ;
  assign n409 = ~n407 & ~n408 ;
  assign n410 = ~n394 & ~n409 ;
  assign n411 = ~n406 & n410 ;
  assign n412 = ~n405 & n411 ;
  assign n413 = ~n394 & ~n406 ;
  assign n414 = ~n405 & n413 ;
  assign n415 = n409 & ~n414 ;
  assign n416 = ~n412 & ~n415 ;
  assign n417 = ~\a[15]  & ~\b[15]  ;
  assign n418 = \a[15]  & \b[15]  ;
  assign n419 = ~n417 & ~n418 ;
  assign n420 = ~n394 & ~n407 ;
  assign n421 = ~n406 & n420 ;
  assign n422 = ~n405 & n421 ;
  assign n423 = ~n408 & ~n422 ;
  assign n424 = ~n419 & ~n423 ;
  assign n425 = ~n408 & n419 ;
  assign n426 = ~n422 & n425 ;
  assign n427 = ~n424 & ~n426 ;
  assign n428 = ~n408 & ~n418 ;
  assign n429 = ~n422 & n428 ;
  assign n430 = ~\a[16]  & ~\b[16]  ;
  assign n431 = \a[16]  & \b[16]  ;
  assign n432 = ~n430 & ~n431 ;
  assign n433 = ~n417 & ~n432 ;
  assign n434 = ~n429 & n433 ;
  assign n435 = n417 & n432 ;
  assign n436 = n428 & n432 ;
  assign n437 = ~n422 & n436 ;
  assign n438 = ~n435 & ~n437 ;
  assign n439 = ~n434 & n438 ;
  assign n440 = n428 & ~n431 ;
  assign n441 = ~n422 & n440 ;
  assign n442 = n417 & ~n431 ;
  assign n443 = ~\a[17]  & ~\b[17]  ;
  assign n444 = \a[17]  & \b[17]  ;
  assign n445 = ~n443 & ~n444 ;
  assign n446 = ~n430 & ~n445 ;
  assign n447 = ~n442 & n446 ;
  assign n448 = ~n441 & n447 ;
  assign n449 = ~n430 & ~n442 ;
  assign n450 = ~n441 & n449 ;
  assign n451 = n445 & ~n450 ;
  assign n452 = ~n448 & ~n451 ;
  assign n453 = ~\a[18]  & ~\b[18]  ;
  assign n454 = \a[18]  & \b[18]  ;
  assign n455 = ~n453 & ~n454 ;
  assign n456 = ~n430 & ~n443 ;
  assign n457 = ~n442 & n456 ;
  assign n458 = ~n441 & n457 ;
  assign n459 = ~n444 & ~n458 ;
  assign n460 = ~n455 & ~n459 ;
  assign n461 = ~n444 & n455 ;
  assign n462 = ~n458 & n461 ;
  assign n463 = ~n460 & ~n462 ;
  assign n464 = ~n444 & ~n454 ;
  assign n465 = ~n458 & n464 ;
  assign n466 = ~\a[19]  & ~\b[19]  ;
  assign n467 = \a[19]  & \b[19]  ;
  assign n468 = ~n466 & ~n467 ;
  assign n469 = ~n453 & ~n468 ;
  assign n470 = ~n465 & n469 ;
  assign n471 = n453 & n468 ;
  assign n472 = n464 & n468 ;
  assign n473 = ~n458 & n472 ;
  assign n474 = ~n471 & ~n473 ;
  assign n475 = ~n470 & n474 ;
  assign n476 = n464 & ~n467 ;
  assign n477 = ~n458 & n476 ;
  assign n478 = n453 & ~n467 ;
  assign n479 = ~\a[20]  & ~\b[20]  ;
  assign n480 = \a[20]  & \b[20]  ;
  assign n481 = ~n479 & ~n480 ;
  assign n482 = ~n466 & ~n481 ;
  assign n483 = ~n478 & n482 ;
  assign n484 = ~n477 & n483 ;
  assign n485 = ~n466 & ~n478 ;
  assign n486 = ~n477 & n485 ;
  assign n487 = n481 & ~n486 ;
  assign n488 = ~n484 & ~n487 ;
  assign n489 = ~\a[21]  & ~\b[21]  ;
  assign n490 = \a[21]  & \b[21]  ;
  assign n491 = ~n489 & ~n490 ;
  assign n492 = ~n466 & ~n479 ;
  assign n493 = ~n478 & n492 ;
  assign n494 = ~n477 & n493 ;
  assign n495 = ~n480 & ~n494 ;
  assign n496 = ~n491 & ~n495 ;
  assign n497 = ~n480 & n491 ;
  assign n498 = ~n494 & n497 ;
  assign n499 = ~n496 & ~n498 ;
  assign n500 = ~n480 & ~n490 ;
  assign n501 = ~n494 & n500 ;
  assign n502 = ~\a[22]  & ~\b[22]  ;
  assign n503 = \a[22]  & \b[22]  ;
  assign n504 = ~n502 & ~n503 ;
  assign n505 = ~n489 & ~n504 ;
  assign n506 = ~n501 & n505 ;
  assign n507 = n489 & n504 ;
  assign n508 = n500 & n504 ;
  assign n509 = ~n494 & n508 ;
  assign n510 = ~n507 & ~n509 ;
  assign n511 = ~n506 & n510 ;
  assign n512 = n500 & ~n503 ;
  assign n513 = ~n494 & n512 ;
  assign n514 = n489 & ~n503 ;
  assign n515 = ~\a[23]  & ~\b[23]  ;
  assign n516 = \a[23]  & \b[23]  ;
  assign n517 = ~n515 & ~n516 ;
  assign n518 = ~n502 & ~n517 ;
  assign n519 = ~n514 & n518 ;
  assign n520 = ~n513 & n519 ;
  assign n521 = ~n502 & ~n514 ;
  assign n522 = ~n513 & n521 ;
  assign n523 = n517 & ~n522 ;
  assign n524 = ~n520 & ~n523 ;
  assign n525 = ~\a[24]  & ~\b[24]  ;
  assign n526 = \a[24]  & \b[24]  ;
  assign n527 = ~n525 & ~n526 ;
  assign n528 = ~n502 & ~n515 ;
  assign n529 = ~n514 & n528 ;
  assign n530 = ~n513 & n529 ;
  assign n531 = ~n516 & ~n530 ;
  assign n532 = ~n527 & ~n531 ;
  assign n533 = ~n516 & n527 ;
  assign n534 = ~n530 & n533 ;
  assign n535 = ~n532 & ~n534 ;
  assign n536 = ~n516 & ~n526 ;
  assign n537 = ~n530 & n536 ;
  assign n538 = ~\a[25]  & ~\b[25]  ;
  assign n539 = \a[25]  & \b[25]  ;
  assign n540 = ~n538 & ~n539 ;
  assign n541 = ~n525 & ~n540 ;
  assign n542 = ~n537 & n541 ;
  assign n543 = n525 & n540 ;
  assign n544 = n536 & n540 ;
  assign n545 = ~n530 & n544 ;
  assign n546 = ~n543 & ~n545 ;
  assign n547 = ~n542 & n546 ;
  assign n548 = n536 & ~n539 ;
  assign n549 = ~n530 & n548 ;
  assign n550 = n525 & ~n539 ;
  assign n551 = ~\a[26]  & ~\b[26]  ;
  assign n552 = \a[26]  & \b[26]  ;
  assign n553 = ~n551 & ~n552 ;
  assign n554 = ~n538 & ~n553 ;
  assign n555 = ~n550 & n554 ;
  assign n556 = ~n549 & n555 ;
  assign n557 = ~n538 & ~n550 ;
  assign n558 = ~n549 & n557 ;
  assign n559 = n553 & ~n558 ;
  assign n560 = ~n556 & ~n559 ;
  assign n561 = ~\a[27]  & ~\b[27]  ;
  assign n562 = \a[27]  & \b[27]  ;
  assign n563 = ~n561 & ~n562 ;
  assign n564 = ~n538 & ~n551 ;
  assign n565 = ~n550 & n564 ;
  assign n566 = ~n549 & n565 ;
  assign n567 = ~n552 & ~n566 ;
  assign n568 = ~n563 & ~n567 ;
  assign n569 = ~n552 & n563 ;
  assign n570 = ~n566 & n569 ;
  assign n571 = ~n568 & ~n570 ;
  assign n572 = ~n552 & ~n562 ;
  assign n573 = ~n566 & n572 ;
  assign n574 = ~\a[28]  & ~\b[28]  ;
  assign n575 = \a[28]  & \b[28]  ;
  assign n576 = ~n574 & ~n575 ;
  assign n577 = ~n561 & ~n576 ;
  assign n578 = ~n573 & n577 ;
  assign n579 = n561 & n576 ;
  assign n580 = n572 & n576 ;
  assign n581 = ~n566 & n580 ;
  assign n582 = ~n579 & ~n581 ;
  assign n583 = ~n578 & n582 ;
  assign n584 = n572 & ~n575 ;
  assign n585 = ~n566 & n584 ;
  assign n586 = n561 & ~n575 ;
  assign n587 = ~\a[29]  & ~\b[29]  ;
  assign n588 = \a[29]  & \b[29]  ;
  assign n589 = ~n587 & ~n588 ;
  assign n590 = ~n574 & ~n589 ;
  assign n591 = ~n586 & n590 ;
  assign n592 = ~n585 & n591 ;
  assign n593 = ~n574 & ~n586 ;
  assign n594 = ~n585 & n593 ;
  assign n595 = n589 & ~n594 ;
  assign n596 = ~n592 & ~n595 ;
  assign n597 = ~\a[30]  & ~\b[30]  ;
  assign n598 = \a[30]  & \b[30]  ;
  assign n599 = ~n597 & ~n598 ;
  assign n600 = ~n574 & ~n587 ;
  assign n601 = ~n586 & n600 ;
  assign n602 = ~n585 & n601 ;
  assign n603 = ~n588 & ~n602 ;
  assign n604 = ~n599 & ~n603 ;
  assign n605 = ~n588 & n599 ;
  assign n606 = ~n602 & n605 ;
  assign n607 = ~n604 & ~n606 ;
  assign n608 = ~n588 & ~n598 ;
  assign n609 = ~n602 & n608 ;
  assign n610 = ~\a[31]  & ~\b[31]  ;
  assign n611 = \a[31]  & \b[31]  ;
  assign n612 = ~n610 & ~n611 ;
  assign n613 = ~n597 & ~n612 ;
  assign n614 = ~n609 & n613 ;
  assign n615 = n597 & n612 ;
  assign n616 = n608 & n612 ;
  assign n617 = ~n602 & n616 ;
  assign n618 = ~n615 & ~n617 ;
  assign n619 = ~n614 & n618 ;
  assign n620 = n608 & ~n611 ;
  assign n621 = ~n602 & n620 ;
  assign n622 = n597 & ~n611 ;
  assign n623 = ~\a[32]  & ~\b[32]  ;
  assign n624 = \a[32]  & \b[32]  ;
  assign n625 = ~n623 & ~n624 ;
  assign n626 = ~n610 & ~n625 ;
  assign n627 = ~n622 & n626 ;
  assign n628 = ~n621 & n627 ;
  assign n629 = ~n610 & ~n622 ;
  assign n630 = ~n621 & n629 ;
  assign n631 = n625 & ~n630 ;
  assign n632 = ~n628 & ~n631 ;
  assign n633 = ~\a[33]  & ~\b[33]  ;
  assign n634 = \a[33]  & \b[33]  ;
  assign n635 = ~n633 & ~n634 ;
  assign n636 = ~n610 & ~n623 ;
  assign n637 = ~n622 & n636 ;
  assign n638 = ~n621 & n637 ;
  assign n639 = ~n624 & ~n638 ;
  assign n640 = ~n635 & ~n639 ;
  assign n641 = ~n624 & n635 ;
  assign n642 = ~n638 & n641 ;
  assign n643 = ~n640 & ~n642 ;
  assign n644 = ~n624 & ~n634 ;
  assign n645 = ~n638 & n644 ;
  assign n646 = ~\a[34]  & ~\b[34]  ;
  assign n647 = \a[34]  & \b[34]  ;
  assign n648 = ~n646 & ~n647 ;
  assign n649 = ~n633 & ~n648 ;
  assign n650 = ~n645 & n649 ;
  assign n651 = n633 & n648 ;
  assign n652 = n644 & n648 ;
  assign n653 = ~n638 & n652 ;
  assign n654 = ~n651 & ~n653 ;
  assign n655 = ~n650 & n654 ;
  assign n656 = n644 & ~n647 ;
  assign n657 = ~n638 & n656 ;
  assign n658 = n633 & ~n647 ;
  assign n659 = ~\a[35]  & ~\b[35]  ;
  assign n660 = \a[35]  & \b[35]  ;
  assign n661 = ~n659 & ~n660 ;
  assign n662 = ~n646 & ~n661 ;
  assign n663 = ~n658 & n662 ;
  assign n664 = ~n657 & n663 ;
  assign n665 = ~n646 & ~n658 ;
  assign n666 = ~n657 & n665 ;
  assign n667 = n661 & ~n666 ;
  assign n668 = ~n664 & ~n667 ;
  assign n669 = ~\a[36]  & ~\b[36]  ;
  assign n670 = \a[36]  & \b[36]  ;
  assign n671 = ~n669 & ~n670 ;
  assign n672 = ~n646 & ~n659 ;
  assign n673 = ~n658 & n672 ;
  assign n674 = ~n657 & n673 ;
  assign n675 = ~n660 & ~n674 ;
  assign n676 = ~n671 & ~n675 ;
  assign n677 = ~n660 & n671 ;
  assign n678 = ~n674 & n677 ;
  assign n679 = ~n676 & ~n678 ;
  assign n680 = ~n660 & ~n670 ;
  assign n681 = ~n674 & n680 ;
  assign n682 = ~\a[37]  & ~\b[37]  ;
  assign n683 = \a[37]  & \b[37]  ;
  assign n684 = ~n682 & ~n683 ;
  assign n685 = ~n669 & ~n684 ;
  assign n686 = ~n681 & n685 ;
  assign n687 = n669 & n684 ;
  assign n688 = n680 & n684 ;
  assign n689 = ~n674 & n688 ;
  assign n690 = ~n687 & ~n689 ;
  assign n691 = ~n686 & n690 ;
  assign n692 = n680 & ~n683 ;
  assign n693 = ~n674 & n692 ;
  assign n694 = n669 & ~n683 ;
  assign n695 = ~\a[38]  & ~\b[38]  ;
  assign n696 = \a[38]  & \b[38]  ;
  assign n697 = ~n695 & ~n696 ;
  assign n698 = ~n682 & ~n697 ;
  assign n699 = ~n694 & n698 ;
  assign n700 = ~n693 & n699 ;
  assign n701 = ~n682 & ~n694 ;
  assign n702 = ~n693 & n701 ;
  assign n703 = n697 & ~n702 ;
  assign n704 = ~n700 & ~n703 ;
  assign n705 = ~\a[39]  & ~\b[39]  ;
  assign n706 = \a[39]  & \b[39]  ;
  assign n707 = ~n705 & ~n706 ;
  assign n708 = ~n682 & ~n695 ;
  assign n709 = ~n694 & n708 ;
  assign n710 = ~n693 & n709 ;
  assign n711 = ~n696 & ~n710 ;
  assign n712 = ~n707 & ~n711 ;
  assign n713 = ~n696 & n707 ;
  assign n714 = ~n710 & n713 ;
  assign n715 = ~n712 & ~n714 ;
  assign n716 = ~n696 & ~n706 ;
  assign n717 = ~n710 & n716 ;
  assign n718 = ~\a[40]  & ~\b[40]  ;
  assign n719 = \a[40]  & \b[40]  ;
  assign n720 = ~n718 & ~n719 ;
  assign n721 = ~n705 & ~n720 ;
  assign n722 = ~n717 & n721 ;
  assign n723 = n705 & n720 ;
  assign n724 = n716 & n720 ;
  assign n725 = ~n710 & n724 ;
  assign n726 = ~n723 & ~n725 ;
  assign n727 = ~n722 & n726 ;
  assign n728 = n716 & ~n719 ;
  assign n729 = ~n710 & n728 ;
  assign n730 = n705 & ~n719 ;
  assign n731 = ~\a[41]  & ~\b[41]  ;
  assign n732 = \a[41]  & \b[41]  ;
  assign n733 = ~n731 & ~n732 ;
  assign n734 = ~n718 & ~n733 ;
  assign n735 = ~n730 & n734 ;
  assign n736 = ~n729 & n735 ;
  assign n737 = ~n718 & ~n730 ;
  assign n738 = ~n729 & n737 ;
  assign n739 = n733 & ~n738 ;
  assign n740 = ~n736 & ~n739 ;
  assign n741 = ~\a[42]  & ~\b[42]  ;
  assign n742 = \a[42]  & \b[42]  ;
  assign n743 = ~n741 & ~n742 ;
  assign n744 = ~n718 & ~n731 ;
  assign n745 = ~n730 & n744 ;
  assign n746 = ~n729 & n745 ;
  assign n747 = ~n732 & ~n746 ;
  assign n748 = ~n743 & ~n747 ;
  assign n749 = ~n732 & n743 ;
  assign n750 = ~n746 & n749 ;
  assign n751 = ~n748 & ~n750 ;
  assign n752 = ~n732 & ~n742 ;
  assign n753 = ~n746 & n752 ;
  assign n754 = ~\a[43]  & ~\b[43]  ;
  assign n755 = \a[43]  & \b[43]  ;
  assign n756 = ~n754 & ~n755 ;
  assign n757 = ~n741 & ~n756 ;
  assign n758 = ~n753 & n757 ;
  assign n759 = n741 & n756 ;
  assign n760 = n752 & n756 ;
  assign n761 = ~n746 & n760 ;
  assign n762 = ~n759 & ~n761 ;
  assign n763 = ~n758 & n762 ;
  assign n764 = n752 & ~n755 ;
  assign n765 = ~n746 & n764 ;
  assign n766 = n741 & ~n755 ;
  assign n767 = ~\a[44]  & ~\b[44]  ;
  assign n768 = \a[44]  & \b[44]  ;
  assign n769 = ~n767 & ~n768 ;
  assign n770 = ~n754 & ~n769 ;
  assign n771 = ~n766 & n770 ;
  assign n772 = ~n765 & n771 ;
  assign n773 = ~n754 & ~n766 ;
  assign n774 = ~n765 & n773 ;
  assign n775 = n769 & ~n774 ;
  assign n776 = ~n772 & ~n775 ;
  assign n777 = ~\a[45]  & ~\b[45]  ;
  assign n778 = \a[45]  & \b[45]  ;
  assign n779 = ~n777 & ~n778 ;
  assign n780 = ~n754 & ~n767 ;
  assign n781 = ~n766 & n780 ;
  assign n782 = ~n765 & n781 ;
  assign n783 = ~n768 & ~n782 ;
  assign n784 = ~n779 & ~n783 ;
  assign n785 = ~n768 & n779 ;
  assign n786 = ~n782 & n785 ;
  assign n787 = ~n784 & ~n786 ;
  assign n788 = ~n768 & ~n778 ;
  assign n789 = ~n782 & n788 ;
  assign n790 = ~\a[46]  & ~\b[46]  ;
  assign n791 = \a[46]  & \b[46]  ;
  assign n792 = ~n790 & ~n791 ;
  assign n793 = ~n777 & ~n792 ;
  assign n794 = ~n789 & n793 ;
  assign n795 = n777 & n792 ;
  assign n796 = n788 & n792 ;
  assign n797 = ~n782 & n796 ;
  assign n798 = ~n795 & ~n797 ;
  assign n799 = ~n794 & n798 ;
  assign n800 = n788 & ~n791 ;
  assign n801 = ~n782 & n800 ;
  assign n802 = n777 & ~n791 ;
  assign n803 = ~\a[47]  & ~\b[47]  ;
  assign n804 = \a[47]  & \b[47]  ;
  assign n805 = ~n803 & ~n804 ;
  assign n806 = ~n790 & ~n805 ;
  assign n807 = ~n802 & n806 ;
  assign n808 = ~n801 & n807 ;
  assign n809 = ~n790 & ~n802 ;
  assign n810 = ~n801 & n809 ;
  assign n811 = n805 & ~n810 ;
  assign n812 = ~n808 & ~n811 ;
  assign n813 = ~\a[48]  & ~\b[48]  ;
  assign n814 = \a[48]  & \b[48]  ;
  assign n815 = ~n813 & ~n814 ;
  assign n816 = ~n790 & ~n803 ;
  assign n817 = ~n802 & n816 ;
  assign n818 = ~n801 & n817 ;
  assign n819 = ~n804 & ~n818 ;
  assign n820 = ~n815 & ~n819 ;
  assign n821 = ~n804 & n815 ;
  assign n822 = ~n818 & n821 ;
  assign n823 = ~n820 & ~n822 ;
  assign n824 = ~n804 & ~n814 ;
  assign n825 = ~n818 & n824 ;
  assign n826 = ~\a[49]  & ~\b[49]  ;
  assign n827 = \a[49]  & \b[49]  ;
  assign n828 = ~n826 & ~n827 ;
  assign n829 = ~n813 & ~n828 ;
  assign n830 = ~n825 & n829 ;
  assign n831 = n813 & n828 ;
  assign n832 = n824 & n828 ;
  assign n833 = ~n818 & n832 ;
  assign n834 = ~n831 & ~n833 ;
  assign n835 = ~n830 & n834 ;
  assign n836 = n824 & ~n827 ;
  assign n837 = ~n818 & n836 ;
  assign n838 = n813 & ~n827 ;
  assign n839 = ~\a[50]  & ~\b[50]  ;
  assign n840 = \a[50]  & \b[50]  ;
  assign n841 = ~n839 & ~n840 ;
  assign n842 = ~n826 & ~n841 ;
  assign n843 = ~n838 & n842 ;
  assign n844 = ~n837 & n843 ;
  assign n845 = ~n826 & ~n838 ;
  assign n846 = ~n837 & n845 ;
  assign n847 = n841 & ~n846 ;
  assign n848 = ~n844 & ~n847 ;
  assign n849 = ~\a[51]  & ~\b[51]  ;
  assign n850 = \a[51]  & \b[51]  ;
  assign n851 = ~n849 & ~n850 ;
  assign n852 = ~n826 & ~n839 ;
  assign n853 = ~n838 & n852 ;
  assign n854 = ~n837 & n853 ;
  assign n855 = ~n840 & ~n854 ;
  assign n856 = ~n851 & ~n855 ;
  assign n857 = ~n840 & n851 ;
  assign n858 = ~n854 & n857 ;
  assign n859 = ~n856 & ~n858 ;
  assign n860 = ~n840 & ~n850 ;
  assign n861 = ~n854 & n860 ;
  assign n862 = ~\a[52]  & ~\b[52]  ;
  assign n863 = \a[52]  & \b[52]  ;
  assign n864 = ~n862 & ~n863 ;
  assign n865 = ~n849 & ~n864 ;
  assign n866 = ~n861 & n865 ;
  assign n867 = n849 & n864 ;
  assign n868 = n860 & n864 ;
  assign n869 = ~n854 & n868 ;
  assign n870 = ~n867 & ~n869 ;
  assign n871 = ~n866 & n870 ;
  assign n872 = n860 & ~n863 ;
  assign n873 = ~n854 & n872 ;
  assign n874 = n849 & ~n863 ;
  assign n875 = ~\a[53]  & ~\b[53]  ;
  assign n876 = \a[53]  & \b[53]  ;
  assign n877 = ~n875 & ~n876 ;
  assign n878 = ~n862 & ~n877 ;
  assign n879 = ~n874 & n878 ;
  assign n880 = ~n873 & n879 ;
  assign n881 = ~n862 & ~n874 ;
  assign n882 = ~n873 & n881 ;
  assign n883 = n877 & ~n882 ;
  assign n884 = ~n880 & ~n883 ;
  assign n885 = ~\a[54]  & ~\b[54]  ;
  assign n886 = \a[54]  & \b[54]  ;
  assign n887 = ~n885 & ~n886 ;
  assign n888 = ~n862 & ~n875 ;
  assign n889 = ~n874 & n888 ;
  assign n890 = ~n873 & n889 ;
  assign n891 = ~n876 & ~n890 ;
  assign n892 = ~n887 & ~n891 ;
  assign n893 = ~n876 & n887 ;
  assign n894 = ~n890 & n893 ;
  assign n895 = ~n892 & ~n894 ;
  assign n896 = ~n876 & ~n886 ;
  assign n897 = ~n890 & n896 ;
  assign n898 = ~\a[55]  & ~\b[55]  ;
  assign n899 = \a[55]  & \b[55]  ;
  assign n900 = ~n898 & ~n899 ;
  assign n901 = ~n885 & ~n900 ;
  assign n902 = ~n897 & n901 ;
  assign n903 = n885 & n900 ;
  assign n904 = n896 & n900 ;
  assign n905 = ~n890 & n904 ;
  assign n906 = ~n903 & ~n905 ;
  assign n907 = ~n902 & n906 ;
  assign n908 = n896 & ~n899 ;
  assign n909 = ~n890 & n908 ;
  assign n910 = n885 & ~n899 ;
  assign n911 = ~\a[56]  & ~\b[56]  ;
  assign n912 = \a[56]  & \b[56]  ;
  assign n913 = ~n911 & ~n912 ;
  assign n914 = ~n898 & ~n913 ;
  assign n915 = ~n910 & n914 ;
  assign n916 = ~n909 & n915 ;
  assign n917 = ~n898 & ~n910 ;
  assign n918 = ~n909 & n917 ;
  assign n919 = n913 & ~n918 ;
  assign n920 = ~n916 & ~n919 ;
  assign n921 = ~\a[57]  & ~\b[57]  ;
  assign n922 = \a[57]  & \b[57]  ;
  assign n923 = ~n921 & ~n922 ;
  assign n924 = ~n898 & ~n911 ;
  assign n925 = ~n910 & n924 ;
  assign n926 = ~n909 & n925 ;
  assign n927 = ~n912 & ~n926 ;
  assign n928 = ~n923 & ~n927 ;
  assign n929 = ~n912 & n923 ;
  assign n930 = ~n926 & n929 ;
  assign n931 = ~n928 & ~n930 ;
  assign n932 = ~n912 & ~n922 ;
  assign n933 = ~n926 & n932 ;
  assign n934 = ~\a[58]  & ~\b[58]  ;
  assign n935 = \a[58]  & \b[58]  ;
  assign n936 = ~n934 & ~n935 ;
  assign n937 = ~n921 & ~n936 ;
  assign n938 = ~n933 & n937 ;
  assign n939 = n921 & n936 ;
  assign n940 = n932 & n936 ;
  assign n941 = ~n926 & n940 ;
  assign n942 = ~n939 & ~n941 ;
  assign n943 = ~n938 & n942 ;
  assign n944 = n932 & ~n935 ;
  assign n945 = ~n926 & n944 ;
  assign n946 = n921 & ~n935 ;
  assign n947 = ~\a[59]  & ~\b[59]  ;
  assign n948 = \a[59]  & \b[59]  ;
  assign n949 = ~n947 & ~n948 ;
  assign n950 = ~n934 & ~n949 ;
  assign n951 = ~n946 & n950 ;
  assign n952 = ~n945 & n951 ;
  assign n953 = ~n934 & ~n946 ;
  assign n954 = ~n945 & n953 ;
  assign n955 = n949 & ~n954 ;
  assign n956 = ~n952 & ~n955 ;
  assign n957 = ~\a[60]  & ~\b[60]  ;
  assign n958 = \a[60]  & \b[60]  ;
  assign n959 = ~n957 & ~n958 ;
  assign n960 = ~n934 & ~n947 ;
  assign n961 = ~n946 & n960 ;
  assign n962 = ~n945 & n961 ;
  assign n963 = ~n948 & ~n962 ;
  assign n964 = ~n959 & ~n963 ;
  assign n965 = ~n948 & n959 ;
  assign n966 = ~n962 & n965 ;
  assign n967 = ~n964 & ~n966 ;
  assign n968 = ~n948 & ~n958 ;
  assign n969 = ~n962 & n968 ;
  assign n970 = ~\a[61]  & ~\b[61]  ;
  assign n971 = \a[61]  & \b[61]  ;
  assign n972 = ~n970 & ~n971 ;
  assign n973 = ~n957 & ~n972 ;
  assign n974 = ~n969 & n973 ;
  assign n975 = n957 & n972 ;
  assign n976 = n968 & n972 ;
  assign n977 = ~n962 & n976 ;
  assign n978 = ~n975 & ~n977 ;
  assign n979 = ~n974 & n978 ;
  assign n980 = n968 & ~n971 ;
  assign n981 = ~n962 & n980 ;
  assign n982 = n957 & ~n971 ;
  assign n983 = ~\a[62]  & ~\b[62]  ;
  assign n984 = \a[62]  & \b[62]  ;
  assign n985 = ~n983 & ~n984 ;
  assign n986 = ~n970 & ~n985 ;
  assign n987 = ~n982 & n986 ;
  assign n988 = ~n981 & n987 ;
  assign n989 = ~n970 & ~n982 ;
  assign n990 = ~n981 & n989 ;
  assign n991 = n985 & ~n990 ;
  assign n992 = ~n988 & ~n991 ;
  assign n993 = ~\a[63]  & ~\b[63]  ;
  assign n994 = \a[63]  & \b[63]  ;
  assign n995 = ~n993 & ~n994 ;
  assign n996 = ~n970 & ~n983 ;
  assign n997 = ~n982 & n996 ;
  assign n998 = ~n981 & n997 ;
  assign n999 = ~n984 & ~n998 ;
  assign n1000 = ~n995 & ~n999 ;
  assign n1001 = ~n984 & n995 ;
  assign n1002 = ~n998 & n1001 ;
  assign n1003 = ~n1000 & ~n1002 ;
  assign n1004 = ~n984 & ~n994 ;
  assign n1005 = ~n998 & n1004 ;
  assign n1006 = ~\a[64]  & ~\b[64]  ;
  assign n1007 = \a[64]  & \b[64]  ;
  assign n1008 = ~n1006 & ~n1007 ;
  assign n1009 = ~n993 & ~n1008 ;
  assign n1010 = ~n1005 & n1009 ;
  assign n1011 = n993 & n1008 ;
  assign n1012 = n1004 & n1008 ;
  assign n1013 = ~n998 & n1012 ;
  assign n1014 = ~n1011 & ~n1013 ;
  assign n1015 = ~n1010 & n1014 ;
  assign n1016 = n1004 & ~n1007 ;
  assign n1017 = ~n998 & n1016 ;
  assign n1018 = n993 & ~n1007 ;
  assign n1019 = ~\a[65]  & ~\b[65]  ;
  assign n1020 = \a[65]  & \b[65]  ;
  assign n1021 = ~n1019 & ~n1020 ;
  assign n1022 = ~n1006 & ~n1021 ;
  assign n1023 = ~n1018 & n1022 ;
  assign n1024 = ~n1017 & n1023 ;
  assign n1025 = ~n1006 & ~n1018 ;
  assign n1026 = ~n1017 & n1025 ;
  assign n1027 = n1021 & ~n1026 ;
  assign n1028 = ~n1024 & ~n1027 ;
  assign n1029 = ~\a[66]  & ~\b[66]  ;
  assign n1030 = \a[66]  & \b[66]  ;
  assign n1031 = ~n1029 & ~n1030 ;
  assign n1032 = ~n1006 & ~n1019 ;
  assign n1033 = ~n1018 & n1032 ;
  assign n1034 = ~n1017 & n1033 ;
  assign n1035 = ~n1020 & ~n1034 ;
  assign n1036 = ~n1031 & ~n1035 ;
  assign n1037 = ~n1020 & n1031 ;
  assign n1038 = ~n1034 & n1037 ;
  assign n1039 = ~n1036 & ~n1038 ;
  assign n1040 = ~n1020 & ~n1030 ;
  assign n1041 = ~n1034 & n1040 ;
  assign n1042 = ~\a[67]  & ~\b[67]  ;
  assign n1043 = \a[67]  & \b[67]  ;
  assign n1044 = ~n1042 & ~n1043 ;
  assign n1045 = ~n1029 & ~n1044 ;
  assign n1046 = ~n1041 & n1045 ;
  assign n1047 = n1029 & n1044 ;
  assign n1048 = n1040 & n1044 ;
  assign n1049 = ~n1034 & n1048 ;
  assign n1050 = ~n1047 & ~n1049 ;
  assign n1051 = ~n1046 & n1050 ;
  assign n1052 = n1040 & ~n1043 ;
  assign n1053 = ~n1034 & n1052 ;
  assign n1054 = n1029 & ~n1043 ;
  assign n1055 = ~\a[68]  & ~\b[68]  ;
  assign n1056 = \a[68]  & \b[68]  ;
  assign n1057 = ~n1055 & ~n1056 ;
  assign n1058 = ~n1042 & ~n1057 ;
  assign n1059 = ~n1054 & n1058 ;
  assign n1060 = ~n1053 & n1059 ;
  assign n1061 = ~n1042 & ~n1054 ;
  assign n1062 = ~n1053 & n1061 ;
  assign n1063 = n1057 & ~n1062 ;
  assign n1064 = ~n1060 & ~n1063 ;
  assign n1065 = ~\a[69]  & ~\b[69]  ;
  assign n1066 = \a[69]  & \b[69]  ;
  assign n1067 = ~n1065 & ~n1066 ;
  assign n1068 = ~n1042 & ~n1055 ;
  assign n1069 = ~n1054 & n1068 ;
  assign n1070 = ~n1053 & n1069 ;
  assign n1071 = ~n1056 & ~n1070 ;
  assign n1072 = ~n1067 & ~n1071 ;
  assign n1073 = ~n1056 & n1067 ;
  assign n1074 = ~n1070 & n1073 ;
  assign n1075 = ~n1072 & ~n1074 ;
  assign n1076 = ~n1056 & ~n1066 ;
  assign n1077 = ~n1070 & n1076 ;
  assign n1078 = ~\a[70]  & ~\b[70]  ;
  assign n1079 = \a[70]  & \b[70]  ;
  assign n1080 = ~n1078 & ~n1079 ;
  assign n1081 = ~n1065 & ~n1080 ;
  assign n1082 = ~n1077 & n1081 ;
  assign n1083 = n1065 & n1080 ;
  assign n1084 = n1076 & n1080 ;
  assign n1085 = ~n1070 & n1084 ;
  assign n1086 = ~n1083 & ~n1085 ;
  assign n1087 = ~n1082 & n1086 ;
  assign n1088 = n1076 & ~n1079 ;
  assign n1089 = ~n1070 & n1088 ;
  assign n1090 = n1065 & ~n1079 ;
  assign n1091 = ~\a[71]  & ~\b[71]  ;
  assign n1092 = \a[71]  & \b[71]  ;
  assign n1093 = ~n1091 & ~n1092 ;
  assign n1094 = ~n1078 & ~n1093 ;
  assign n1095 = ~n1090 & n1094 ;
  assign n1096 = ~n1089 & n1095 ;
  assign n1097 = ~n1078 & ~n1090 ;
  assign n1098 = ~n1089 & n1097 ;
  assign n1099 = n1093 & ~n1098 ;
  assign n1100 = ~n1096 & ~n1099 ;
  assign n1101 = ~\a[72]  & ~\b[72]  ;
  assign n1102 = \a[72]  & \b[72]  ;
  assign n1103 = ~n1101 & ~n1102 ;
  assign n1104 = ~n1078 & ~n1091 ;
  assign n1105 = ~n1090 & n1104 ;
  assign n1106 = ~n1089 & n1105 ;
  assign n1107 = ~n1092 & ~n1106 ;
  assign n1108 = ~n1103 & ~n1107 ;
  assign n1109 = ~n1092 & n1103 ;
  assign n1110 = ~n1106 & n1109 ;
  assign n1111 = ~n1108 & ~n1110 ;
  assign n1112 = ~n1092 & ~n1102 ;
  assign n1113 = ~n1106 & n1112 ;
  assign n1114 = ~\a[73]  & ~\b[73]  ;
  assign n1115 = \a[73]  & \b[73]  ;
  assign n1116 = ~n1114 & ~n1115 ;
  assign n1117 = ~n1101 & ~n1116 ;
  assign n1118 = ~n1113 & n1117 ;
  assign n1119 = n1101 & n1116 ;
  assign n1120 = n1112 & n1116 ;
  assign n1121 = ~n1106 & n1120 ;
  assign n1122 = ~n1119 & ~n1121 ;
  assign n1123 = ~n1118 & n1122 ;
  assign n1124 = n1112 & ~n1115 ;
  assign n1125 = ~n1106 & n1124 ;
  assign n1126 = n1101 & ~n1115 ;
  assign n1127 = ~\a[74]  & ~\b[74]  ;
  assign n1128 = \a[74]  & \b[74]  ;
  assign n1129 = ~n1127 & ~n1128 ;
  assign n1130 = ~n1114 & ~n1129 ;
  assign n1131 = ~n1126 & n1130 ;
  assign n1132 = ~n1125 & n1131 ;
  assign n1133 = ~n1114 & ~n1126 ;
  assign n1134 = ~n1125 & n1133 ;
  assign n1135 = n1129 & ~n1134 ;
  assign n1136 = ~n1132 & ~n1135 ;
  assign n1137 = ~\a[75]  & ~\b[75]  ;
  assign n1138 = \a[75]  & \b[75]  ;
  assign n1139 = ~n1137 & ~n1138 ;
  assign n1140 = ~n1114 & ~n1127 ;
  assign n1141 = ~n1126 & n1140 ;
  assign n1142 = ~n1125 & n1141 ;
  assign n1143 = ~n1128 & ~n1142 ;
  assign n1144 = ~n1139 & ~n1143 ;
  assign n1145 = ~n1128 & n1139 ;
  assign n1146 = ~n1142 & n1145 ;
  assign n1147 = ~n1144 & ~n1146 ;
  assign n1148 = ~n1128 & ~n1138 ;
  assign n1149 = ~n1142 & n1148 ;
  assign n1150 = ~\a[76]  & ~\b[76]  ;
  assign n1151 = \a[76]  & \b[76]  ;
  assign n1152 = ~n1150 & ~n1151 ;
  assign n1153 = ~n1137 & ~n1152 ;
  assign n1154 = ~n1149 & n1153 ;
  assign n1155 = n1137 & n1152 ;
  assign n1156 = n1148 & n1152 ;
  assign n1157 = ~n1142 & n1156 ;
  assign n1158 = ~n1155 & ~n1157 ;
  assign n1159 = ~n1154 & n1158 ;
  assign n1160 = n1148 & ~n1151 ;
  assign n1161 = ~n1142 & n1160 ;
  assign n1162 = n1137 & ~n1151 ;
  assign n1163 = ~\a[77]  & ~\b[77]  ;
  assign n1164 = \a[77]  & \b[77]  ;
  assign n1165 = ~n1163 & ~n1164 ;
  assign n1166 = ~n1150 & ~n1165 ;
  assign n1167 = ~n1162 & n1166 ;
  assign n1168 = ~n1161 & n1167 ;
  assign n1169 = ~n1150 & ~n1162 ;
  assign n1170 = ~n1161 & n1169 ;
  assign n1171 = n1165 & ~n1170 ;
  assign n1172 = ~n1168 & ~n1171 ;
  assign n1173 = ~\a[78]  & ~\b[78]  ;
  assign n1174 = \a[78]  & \b[78]  ;
  assign n1175 = ~n1173 & ~n1174 ;
  assign n1176 = ~n1150 & ~n1163 ;
  assign n1177 = ~n1162 & n1176 ;
  assign n1178 = ~n1161 & n1177 ;
  assign n1179 = ~n1164 & ~n1178 ;
  assign n1180 = ~n1175 & ~n1179 ;
  assign n1181 = ~n1164 & n1175 ;
  assign n1182 = ~n1178 & n1181 ;
  assign n1183 = ~n1180 & ~n1182 ;
  assign n1184 = ~n1164 & ~n1174 ;
  assign n1185 = ~n1178 & n1184 ;
  assign n1186 = ~\a[79]  & ~\b[79]  ;
  assign n1187 = \a[79]  & \b[79]  ;
  assign n1188 = ~n1186 & ~n1187 ;
  assign n1189 = ~n1173 & ~n1188 ;
  assign n1190 = ~n1185 & n1189 ;
  assign n1191 = n1173 & n1188 ;
  assign n1192 = n1184 & n1188 ;
  assign n1193 = ~n1178 & n1192 ;
  assign n1194 = ~n1191 & ~n1193 ;
  assign n1195 = ~n1190 & n1194 ;
  assign n1196 = n1184 & ~n1187 ;
  assign n1197 = ~n1178 & n1196 ;
  assign n1198 = n1173 & ~n1187 ;
  assign n1199 = ~\a[80]  & ~\b[80]  ;
  assign n1200 = \a[80]  & \b[80]  ;
  assign n1201 = ~n1199 & ~n1200 ;
  assign n1202 = ~n1186 & ~n1201 ;
  assign n1203 = ~n1198 & n1202 ;
  assign n1204 = ~n1197 & n1203 ;
  assign n1205 = ~n1186 & ~n1198 ;
  assign n1206 = ~n1197 & n1205 ;
  assign n1207 = n1201 & ~n1206 ;
  assign n1208 = ~n1204 & ~n1207 ;
  assign n1209 = ~\a[81]  & ~\b[81]  ;
  assign n1210 = \a[81]  & \b[81]  ;
  assign n1211 = ~n1209 & ~n1210 ;
  assign n1212 = ~n1186 & ~n1199 ;
  assign n1213 = ~n1198 & n1212 ;
  assign n1214 = ~n1197 & n1213 ;
  assign n1215 = ~n1200 & ~n1214 ;
  assign n1216 = ~n1211 & ~n1215 ;
  assign n1217 = ~n1200 & n1211 ;
  assign n1218 = ~n1214 & n1217 ;
  assign n1219 = ~n1216 & ~n1218 ;
  assign n1220 = ~n1200 & ~n1210 ;
  assign n1221 = ~n1214 & n1220 ;
  assign n1222 = ~\a[82]  & ~\b[82]  ;
  assign n1223 = \a[82]  & \b[82]  ;
  assign n1224 = ~n1222 & ~n1223 ;
  assign n1225 = ~n1209 & ~n1224 ;
  assign n1226 = ~n1221 & n1225 ;
  assign n1227 = n1209 & n1224 ;
  assign n1228 = n1220 & n1224 ;
  assign n1229 = ~n1214 & n1228 ;
  assign n1230 = ~n1227 & ~n1229 ;
  assign n1231 = ~n1226 & n1230 ;
  assign n1232 = n1220 & ~n1223 ;
  assign n1233 = ~n1214 & n1232 ;
  assign n1234 = n1209 & ~n1223 ;
  assign n1235 = ~\a[83]  & ~\b[83]  ;
  assign n1236 = \a[83]  & \b[83]  ;
  assign n1237 = ~n1235 & ~n1236 ;
  assign n1238 = ~n1222 & ~n1237 ;
  assign n1239 = ~n1234 & n1238 ;
  assign n1240 = ~n1233 & n1239 ;
  assign n1241 = ~n1222 & ~n1234 ;
  assign n1242 = ~n1233 & n1241 ;
  assign n1243 = n1237 & ~n1242 ;
  assign n1244 = ~n1240 & ~n1243 ;
  assign n1245 = ~\a[84]  & ~\b[84]  ;
  assign n1246 = \a[84]  & \b[84]  ;
  assign n1247 = ~n1245 & ~n1246 ;
  assign n1248 = ~n1222 & ~n1235 ;
  assign n1249 = ~n1234 & n1248 ;
  assign n1250 = ~n1233 & n1249 ;
  assign n1251 = ~n1236 & ~n1250 ;
  assign n1252 = ~n1247 & ~n1251 ;
  assign n1253 = ~n1236 & n1247 ;
  assign n1254 = ~n1250 & n1253 ;
  assign n1255 = ~n1252 & ~n1254 ;
  assign n1256 = ~n1236 & ~n1246 ;
  assign n1257 = ~n1250 & n1256 ;
  assign n1258 = ~\a[85]  & ~\b[85]  ;
  assign n1259 = \a[85]  & \b[85]  ;
  assign n1260 = ~n1258 & ~n1259 ;
  assign n1261 = ~n1245 & ~n1260 ;
  assign n1262 = ~n1257 & n1261 ;
  assign n1263 = n1245 & n1260 ;
  assign n1264 = n1256 & n1260 ;
  assign n1265 = ~n1250 & n1264 ;
  assign n1266 = ~n1263 & ~n1265 ;
  assign n1267 = ~n1262 & n1266 ;
  assign n1268 = n1256 & ~n1259 ;
  assign n1269 = ~n1250 & n1268 ;
  assign n1270 = n1245 & ~n1259 ;
  assign n1271 = ~\a[86]  & ~\b[86]  ;
  assign n1272 = \a[86]  & \b[86]  ;
  assign n1273 = ~n1271 & ~n1272 ;
  assign n1274 = ~n1258 & ~n1273 ;
  assign n1275 = ~n1270 & n1274 ;
  assign n1276 = ~n1269 & n1275 ;
  assign n1277 = ~n1258 & ~n1270 ;
  assign n1278 = ~n1269 & n1277 ;
  assign n1279 = n1273 & ~n1278 ;
  assign n1280 = ~n1276 & ~n1279 ;
  assign n1281 = ~\a[87]  & ~\b[87]  ;
  assign n1282 = \a[87]  & \b[87]  ;
  assign n1283 = ~n1281 & ~n1282 ;
  assign n1284 = ~n1258 & ~n1271 ;
  assign n1285 = ~n1270 & n1284 ;
  assign n1286 = ~n1269 & n1285 ;
  assign n1287 = ~n1272 & ~n1286 ;
  assign n1288 = ~n1283 & ~n1287 ;
  assign n1289 = ~n1272 & n1283 ;
  assign n1290 = ~n1286 & n1289 ;
  assign n1291 = ~n1288 & ~n1290 ;
  assign n1292 = ~n1272 & ~n1282 ;
  assign n1293 = ~n1286 & n1292 ;
  assign n1294 = ~\a[88]  & ~\b[88]  ;
  assign n1295 = \a[88]  & \b[88]  ;
  assign n1296 = ~n1294 & ~n1295 ;
  assign n1297 = ~n1281 & ~n1296 ;
  assign n1298 = ~n1293 & n1297 ;
  assign n1299 = n1281 & n1296 ;
  assign n1300 = n1292 & n1296 ;
  assign n1301 = ~n1286 & n1300 ;
  assign n1302 = ~n1299 & ~n1301 ;
  assign n1303 = ~n1298 & n1302 ;
  assign n1304 = n1292 & ~n1295 ;
  assign n1305 = ~n1286 & n1304 ;
  assign n1306 = n1281 & ~n1295 ;
  assign n1307 = ~\a[89]  & ~\b[89]  ;
  assign n1308 = \a[89]  & \b[89]  ;
  assign n1309 = ~n1307 & ~n1308 ;
  assign n1310 = ~n1294 & ~n1309 ;
  assign n1311 = ~n1306 & n1310 ;
  assign n1312 = ~n1305 & n1311 ;
  assign n1313 = ~n1294 & ~n1306 ;
  assign n1314 = ~n1305 & n1313 ;
  assign n1315 = n1309 & ~n1314 ;
  assign n1316 = ~n1312 & ~n1315 ;
  assign n1317 = ~\a[90]  & ~\b[90]  ;
  assign n1318 = \a[90]  & \b[90]  ;
  assign n1319 = ~n1317 & ~n1318 ;
  assign n1320 = ~n1294 & ~n1307 ;
  assign n1321 = ~n1306 & n1320 ;
  assign n1322 = ~n1305 & n1321 ;
  assign n1323 = ~n1308 & ~n1322 ;
  assign n1324 = ~n1319 & ~n1323 ;
  assign n1325 = ~n1308 & n1319 ;
  assign n1326 = ~n1322 & n1325 ;
  assign n1327 = ~n1324 & ~n1326 ;
  assign n1328 = ~n1308 & ~n1318 ;
  assign n1329 = ~n1322 & n1328 ;
  assign n1330 = ~\a[91]  & ~\b[91]  ;
  assign n1331 = \a[91]  & \b[91]  ;
  assign n1332 = ~n1330 & ~n1331 ;
  assign n1333 = ~n1317 & ~n1332 ;
  assign n1334 = ~n1329 & n1333 ;
  assign n1335 = n1317 & n1332 ;
  assign n1336 = n1328 & n1332 ;
  assign n1337 = ~n1322 & n1336 ;
  assign n1338 = ~n1335 & ~n1337 ;
  assign n1339 = ~n1334 & n1338 ;
  assign n1340 = n1328 & ~n1331 ;
  assign n1341 = ~n1322 & n1340 ;
  assign n1342 = n1317 & ~n1331 ;
  assign n1343 = ~\a[92]  & ~\b[92]  ;
  assign n1344 = \a[92]  & \b[92]  ;
  assign n1345 = ~n1343 & ~n1344 ;
  assign n1346 = ~n1330 & ~n1345 ;
  assign n1347 = ~n1342 & n1346 ;
  assign n1348 = ~n1341 & n1347 ;
  assign n1349 = ~n1330 & ~n1342 ;
  assign n1350 = ~n1341 & n1349 ;
  assign n1351 = n1345 & ~n1350 ;
  assign n1352 = ~n1348 & ~n1351 ;
  assign n1353 = ~\a[93]  & ~\b[93]  ;
  assign n1354 = \a[93]  & \b[93]  ;
  assign n1355 = ~n1353 & ~n1354 ;
  assign n1356 = ~n1330 & ~n1343 ;
  assign n1357 = ~n1342 & n1356 ;
  assign n1358 = ~n1341 & n1357 ;
  assign n1359 = ~n1344 & ~n1358 ;
  assign n1360 = ~n1355 & ~n1359 ;
  assign n1361 = ~n1344 & n1355 ;
  assign n1362 = ~n1358 & n1361 ;
  assign n1363 = ~n1360 & ~n1362 ;
  assign n1364 = ~n1344 & ~n1354 ;
  assign n1365 = ~n1358 & n1364 ;
  assign n1366 = ~\a[94]  & ~\b[94]  ;
  assign n1367 = \a[94]  & \b[94]  ;
  assign n1368 = ~n1366 & ~n1367 ;
  assign n1369 = ~n1353 & ~n1368 ;
  assign n1370 = ~n1365 & n1369 ;
  assign n1371 = n1353 & n1368 ;
  assign n1372 = n1364 & n1368 ;
  assign n1373 = ~n1358 & n1372 ;
  assign n1374 = ~n1371 & ~n1373 ;
  assign n1375 = ~n1370 & n1374 ;
  assign n1376 = n1364 & ~n1367 ;
  assign n1377 = ~n1358 & n1376 ;
  assign n1378 = n1353 & ~n1367 ;
  assign n1379 = ~\a[95]  & ~\b[95]  ;
  assign n1380 = \a[95]  & \b[95]  ;
  assign n1381 = ~n1379 & ~n1380 ;
  assign n1382 = ~n1366 & ~n1381 ;
  assign n1383 = ~n1378 & n1382 ;
  assign n1384 = ~n1377 & n1383 ;
  assign n1385 = ~n1366 & ~n1378 ;
  assign n1386 = ~n1377 & n1385 ;
  assign n1387 = n1381 & ~n1386 ;
  assign n1388 = ~n1384 & ~n1387 ;
  assign n1389 = ~\a[96]  & ~\b[96]  ;
  assign n1390 = \a[96]  & \b[96]  ;
  assign n1391 = ~n1389 & ~n1390 ;
  assign n1392 = ~n1366 & ~n1379 ;
  assign n1393 = ~n1378 & n1392 ;
  assign n1394 = ~n1377 & n1393 ;
  assign n1395 = ~n1380 & ~n1394 ;
  assign n1396 = ~n1391 & ~n1395 ;
  assign n1397 = ~n1380 & n1391 ;
  assign n1398 = ~n1394 & n1397 ;
  assign n1399 = ~n1396 & ~n1398 ;
  assign n1400 = ~n1380 & ~n1390 ;
  assign n1401 = ~n1394 & n1400 ;
  assign n1402 = ~\a[97]  & ~\b[97]  ;
  assign n1403 = \a[97]  & \b[97]  ;
  assign n1404 = ~n1402 & ~n1403 ;
  assign n1405 = ~n1389 & ~n1404 ;
  assign n1406 = ~n1401 & n1405 ;
  assign n1407 = n1389 & n1404 ;
  assign n1408 = n1400 & n1404 ;
  assign n1409 = ~n1394 & n1408 ;
  assign n1410 = ~n1407 & ~n1409 ;
  assign n1411 = ~n1406 & n1410 ;
  assign n1412 = n1400 & ~n1403 ;
  assign n1413 = ~n1394 & n1412 ;
  assign n1414 = n1389 & ~n1403 ;
  assign n1415 = ~\a[98]  & ~\b[98]  ;
  assign n1416 = \a[98]  & \b[98]  ;
  assign n1417 = ~n1415 & ~n1416 ;
  assign n1418 = ~n1402 & ~n1417 ;
  assign n1419 = ~n1414 & n1418 ;
  assign n1420 = ~n1413 & n1419 ;
  assign n1421 = ~n1402 & ~n1414 ;
  assign n1422 = ~n1413 & n1421 ;
  assign n1423 = n1417 & ~n1422 ;
  assign n1424 = ~n1420 & ~n1423 ;
  assign n1425 = ~\a[99]  & ~\b[99]  ;
  assign n1426 = \a[99]  & \b[99]  ;
  assign n1427 = ~n1425 & ~n1426 ;
  assign n1428 = ~n1402 & ~n1415 ;
  assign n1429 = ~n1414 & n1428 ;
  assign n1430 = ~n1413 & n1429 ;
  assign n1431 = ~n1416 & ~n1430 ;
  assign n1432 = ~n1427 & ~n1431 ;
  assign n1433 = ~n1416 & n1427 ;
  assign n1434 = ~n1430 & n1433 ;
  assign n1435 = ~n1432 & ~n1434 ;
  assign n1436 = ~n1416 & ~n1426 ;
  assign n1437 = ~n1430 & n1436 ;
  assign n1438 = ~\a[100]  & ~\b[100]  ;
  assign n1439 = \a[100]  & \b[100]  ;
  assign n1440 = ~n1438 & ~n1439 ;
  assign n1441 = ~n1425 & ~n1440 ;
  assign n1442 = ~n1437 & n1441 ;
  assign n1443 = n1425 & n1440 ;
  assign n1444 = n1436 & n1440 ;
  assign n1445 = ~n1430 & n1444 ;
  assign n1446 = ~n1443 & ~n1445 ;
  assign n1447 = ~n1442 & n1446 ;
  assign n1448 = n1436 & ~n1439 ;
  assign n1449 = ~n1430 & n1448 ;
  assign n1450 = n1425 & ~n1439 ;
  assign n1451 = ~\a[101]  & ~\b[101]  ;
  assign n1452 = \a[101]  & \b[101]  ;
  assign n1453 = ~n1451 & ~n1452 ;
  assign n1454 = ~n1438 & ~n1453 ;
  assign n1455 = ~n1450 & n1454 ;
  assign n1456 = ~n1449 & n1455 ;
  assign n1457 = ~n1438 & ~n1450 ;
  assign n1458 = ~n1449 & n1457 ;
  assign n1459 = n1453 & ~n1458 ;
  assign n1460 = ~n1456 & ~n1459 ;
  assign n1461 = ~\a[102]  & ~\b[102]  ;
  assign n1462 = \a[102]  & \b[102]  ;
  assign n1463 = ~n1461 & ~n1462 ;
  assign n1464 = ~n1438 & ~n1451 ;
  assign n1465 = ~n1450 & n1464 ;
  assign n1466 = ~n1449 & n1465 ;
  assign n1467 = ~n1452 & ~n1466 ;
  assign n1468 = ~n1463 & ~n1467 ;
  assign n1469 = ~n1452 & n1463 ;
  assign n1470 = ~n1466 & n1469 ;
  assign n1471 = ~n1468 & ~n1470 ;
  assign n1472 = ~n1452 & ~n1462 ;
  assign n1473 = ~n1466 & n1472 ;
  assign n1474 = ~\a[103]  & ~\b[103]  ;
  assign n1475 = \a[103]  & \b[103]  ;
  assign n1476 = ~n1474 & ~n1475 ;
  assign n1477 = ~n1461 & ~n1476 ;
  assign n1478 = ~n1473 & n1477 ;
  assign n1479 = n1461 & n1476 ;
  assign n1480 = n1472 & n1476 ;
  assign n1481 = ~n1466 & n1480 ;
  assign n1482 = ~n1479 & ~n1481 ;
  assign n1483 = ~n1478 & n1482 ;
  assign n1484 = n1472 & ~n1475 ;
  assign n1485 = ~n1466 & n1484 ;
  assign n1486 = n1461 & ~n1475 ;
  assign n1487 = ~\a[104]  & ~\b[104]  ;
  assign n1488 = \a[104]  & \b[104]  ;
  assign n1489 = ~n1487 & ~n1488 ;
  assign n1490 = ~n1474 & ~n1489 ;
  assign n1491 = ~n1486 & n1490 ;
  assign n1492 = ~n1485 & n1491 ;
  assign n1493 = ~n1474 & ~n1486 ;
  assign n1494 = ~n1485 & n1493 ;
  assign n1495 = n1489 & ~n1494 ;
  assign n1496 = ~n1492 & ~n1495 ;
  assign n1497 = ~\a[105]  & ~\b[105]  ;
  assign n1498 = \a[105]  & \b[105]  ;
  assign n1499 = ~n1497 & ~n1498 ;
  assign n1500 = ~n1474 & ~n1487 ;
  assign n1501 = ~n1486 & n1500 ;
  assign n1502 = ~n1485 & n1501 ;
  assign n1503 = ~n1488 & ~n1502 ;
  assign n1504 = ~n1499 & ~n1503 ;
  assign n1505 = ~n1488 & n1499 ;
  assign n1506 = ~n1502 & n1505 ;
  assign n1507 = ~n1504 & ~n1506 ;
  assign n1508 = ~n1488 & ~n1498 ;
  assign n1509 = ~n1502 & n1508 ;
  assign n1510 = ~\a[106]  & ~\b[106]  ;
  assign n1511 = \a[106]  & \b[106]  ;
  assign n1512 = ~n1510 & ~n1511 ;
  assign n1513 = ~n1497 & ~n1512 ;
  assign n1514 = ~n1509 & n1513 ;
  assign n1515 = n1497 & n1512 ;
  assign n1516 = n1508 & n1512 ;
  assign n1517 = ~n1502 & n1516 ;
  assign n1518 = ~n1515 & ~n1517 ;
  assign n1519 = ~n1514 & n1518 ;
  assign n1520 = n1508 & ~n1511 ;
  assign n1521 = ~n1502 & n1520 ;
  assign n1522 = n1497 & ~n1511 ;
  assign n1523 = ~\a[107]  & ~\b[107]  ;
  assign n1524 = \a[107]  & \b[107]  ;
  assign n1525 = ~n1523 & ~n1524 ;
  assign n1526 = ~n1510 & ~n1525 ;
  assign n1527 = ~n1522 & n1526 ;
  assign n1528 = ~n1521 & n1527 ;
  assign n1529 = ~n1510 & ~n1522 ;
  assign n1530 = ~n1521 & n1529 ;
  assign n1531 = n1525 & ~n1530 ;
  assign n1532 = ~n1528 & ~n1531 ;
  assign n1533 = ~\a[108]  & ~\b[108]  ;
  assign n1534 = \a[108]  & \b[108]  ;
  assign n1535 = ~n1533 & ~n1534 ;
  assign n1536 = ~n1510 & ~n1523 ;
  assign n1537 = ~n1522 & n1536 ;
  assign n1538 = ~n1521 & n1537 ;
  assign n1539 = ~n1524 & ~n1538 ;
  assign n1540 = ~n1535 & ~n1539 ;
  assign n1541 = ~n1524 & n1535 ;
  assign n1542 = ~n1538 & n1541 ;
  assign n1543 = ~n1540 & ~n1542 ;
  assign n1544 = ~n1524 & ~n1534 ;
  assign n1545 = ~n1538 & n1544 ;
  assign n1546 = ~\a[109]  & ~\b[109]  ;
  assign n1547 = \a[109]  & \b[109]  ;
  assign n1548 = ~n1546 & ~n1547 ;
  assign n1549 = ~n1533 & ~n1548 ;
  assign n1550 = ~n1545 & n1549 ;
  assign n1551 = n1533 & n1548 ;
  assign n1552 = n1544 & n1548 ;
  assign n1553 = ~n1538 & n1552 ;
  assign n1554 = ~n1551 & ~n1553 ;
  assign n1555 = ~n1550 & n1554 ;
  assign n1556 = n1544 & ~n1547 ;
  assign n1557 = ~n1538 & n1556 ;
  assign n1558 = n1533 & ~n1547 ;
  assign n1559 = ~\a[110]  & ~\b[110]  ;
  assign n1560 = \a[110]  & \b[110]  ;
  assign n1561 = ~n1559 & ~n1560 ;
  assign n1562 = ~n1546 & ~n1561 ;
  assign n1563 = ~n1558 & n1562 ;
  assign n1564 = ~n1557 & n1563 ;
  assign n1565 = ~n1546 & ~n1558 ;
  assign n1566 = ~n1557 & n1565 ;
  assign n1567 = n1561 & ~n1566 ;
  assign n1568 = ~n1564 & ~n1567 ;
  assign n1569 = ~\a[111]  & ~\b[111]  ;
  assign n1570 = \a[111]  & \b[111]  ;
  assign n1571 = ~n1569 & ~n1570 ;
  assign n1572 = ~n1546 & ~n1559 ;
  assign n1573 = ~n1558 & n1572 ;
  assign n1574 = ~n1557 & n1573 ;
  assign n1575 = ~n1560 & ~n1574 ;
  assign n1576 = ~n1571 & ~n1575 ;
  assign n1577 = ~n1560 & n1571 ;
  assign n1578 = ~n1574 & n1577 ;
  assign n1579 = ~n1576 & ~n1578 ;
  assign n1580 = ~n1560 & ~n1570 ;
  assign n1581 = ~n1574 & n1580 ;
  assign n1582 = ~\a[112]  & ~\b[112]  ;
  assign n1583 = \a[112]  & \b[112]  ;
  assign n1584 = ~n1582 & ~n1583 ;
  assign n1585 = ~n1569 & ~n1584 ;
  assign n1586 = ~n1581 & n1585 ;
  assign n1587 = n1569 & n1584 ;
  assign n1588 = n1580 & n1584 ;
  assign n1589 = ~n1574 & n1588 ;
  assign n1590 = ~n1587 & ~n1589 ;
  assign n1591 = ~n1586 & n1590 ;
  assign n1592 = n1580 & ~n1583 ;
  assign n1593 = ~n1574 & n1592 ;
  assign n1594 = n1569 & ~n1583 ;
  assign n1595 = ~\a[113]  & ~\b[113]  ;
  assign n1596 = \a[113]  & \b[113]  ;
  assign n1597 = ~n1595 & ~n1596 ;
  assign n1598 = ~n1582 & ~n1597 ;
  assign n1599 = ~n1594 & n1598 ;
  assign n1600 = ~n1593 & n1599 ;
  assign n1601 = ~n1582 & ~n1594 ;
  assign n1602 = ~n1593 & n1601 ;
  assign n1603 = n1597 & ~n1602 ;
  assign n1604 = ~n1600 & ~n1603 ;
  assign n1605 = ~\a[114]  & ~\b[114]  ;
  assign n1606 = \a[114]  & \b[114]  ;
  assign n1607 = ~n1605 & ~n1606 ;
  assign n1608 = ~n1582 & ~n1595 ;
  assign n1609 = ~n1594 & n1608 ;
  assign n1610 = ~n1593 & n1609 ;
  assign n1611 = ~n1596 & ~n1610 ;
  assign n1612 = ~n1607 & ~n1611 ;
  assign n1613 = ~n1596 & n1607 ;
  assign n1614 = ~n1610 & n1613 ;
  assign n1615 = ~n1612 & ~n1614 ;
  assign n1616 = ~n1596 & ~n1606 ;
  assign n1617 = ~n1610 & n1616 ;
  assign n1618 = ~\a[115]  & ~\b[115]  ;
  assign n1619 = \a[115]  & \b[115]  ;
  assign n1620 = ~n1618 & ~n1619 ;
  assign n1621 = ~n1605 & ~n1620 ;
  assign n1622 = ~n1617 & n1621 ;
  assign n1623 = n1605 & n1620 ;
  assign n1624 = n1616 & n1620 ;
  assign n1625 = ~n1610 & n1624 ;
  assign n1626 = ~n1623 & ~n1625 ;
  assign n1627 = ~n1622 & n1626 ;
  assign n1628 = n1616 & ~n1619 ;
  assign n1629 = ~n1610 & n1628 ;
  assign n1630 = n1605 & ~n1619 ;
  assign n1631 = ~\a[116]  & ~\b[116]  ;
  assign n1632 = \a[116]  & \b[116]  ;
  assign n1633 = ~n1631 & ~n1632 ;
  assign n1634 = ~n1618 & ~n1633 ;
  assign n1635 = ~n1630 & n1634 ;
  assign n1636 = ~n1629 & n1635 ;
  assign n1637 = ~n1618 & ~n1630 ;
  assign n1638 = ~n1629 & n1637 ;
  assign n1639 = n1633 & ~n1638 ;
  assign n1640 = ~n1636 & ~n1639 ;
  assign n1641 = ~\a[117]  & ~\b[117]  ;
  assign n1642 = \a[117]  & \b[117]  ;
  assign n1643 = ~n1641 & ~n1642 ;
  assign n1644 = ~n1618 & ~n1631 ;
  assign n1645 = ~n1630 & n1644 ;
  assign n1646 = ~n1629 & n1645 ;
  assign n1647 = ~n1632 & ~n1646 ;
  assign n1648 = ~n1643 & ~n1647 ;
  assign n1649 = ~n1632 & n1643 ;
  assign n1650 = ~n1646 & n1649 ;
  assign n1651 = ~n1648 & ~n1650 ;
  assign n1652 = ~n1632 & ~n1642 ;
  assign n1653 = ~n1646 & n1652 ;
  assign n1654 = ~\a[118]  & ~\b[118]  ;
  assign n1655 = \a[118]  & \b[118]  ;
  assign n1656 = ~n1654 & ~n1655 ;
  assign n1657 = ~n1641 & ~n1656 ;
  assign n1658 = ~n1653 & n1657 ;
  assign n1659 = n1641 & n1656 ;
  assign n1660 = n1652 & n1656 ;
  assign n1661 = ~n1646 & n1660 ;
  assign n1662 = ~n1659 & ~n1661 ;
  assign n1663 = ~n1658 & n1662 ;
  assign n1664 = n1652 & ~n1655 ;
  assign n1665 = ~n1646 & n1664 ;
  assign n1666 = n1641 & ~n1655 ;
  assign n1667 = ~\a[119]  & ~\b[119]  ;
  assign n1668 = \a[119]  & \b[119]  ;
  assign n1669 = ~n1667 & ~n1668 ;
  assign n1670 = ~n1654 & ~n1669 ;
  assign n1671 = ~n1666 & n1670 ;
  assign n1672 = ~n1665 & n1671 ;
  assign n1673 = ~n1654 & ~n1666 ;
  assign n1674 = ~n1665 & n1673 ;
  assign n1675 = n1669 & ~n1674 ;
  assign n1676 = ~n1672 & ~n1675 ;
  assign n1677 = ~\a[120]  & ~\b[120]  ;
  assign n1678 = \a[120]  & \b[120]  ;
  assign n1679 = ~n1677 & ~n1678 ;
  assign n1680 = ~n1654 & ~n1667 ;
  assign n1681 = ~n1666 & n1680 ;
  assign n1682 = ~n1665 & n1681 ;
  assign n1683 = ~n1668 & ~n1682 ;
  assign n1684 = ~n1679 & ~n1683 ;
  assign n1685 = ~n1668 & n1679 ;
  assign n1686 = ~n1682 & n1685 ;
  assign n1687 = ~n1684 & ~n1686 ;
  assign n1688 = ~n1668 & ~n1678 ;
  assign n1689 = ~n1682 & n1688 ;
  assign n1690 = ~\a[121]  & ~\b[121]  ;
  assign n1691 = \a[121]  & \b[121]  ;
  assign n1692 = ~n1690 & ~n1691 ;
  assign n1693 = ~n1677 & ~n1692 ;
  assign n1694 = ~n1689 & n1693 ;
  assign n1695 = n1677 & n1692 ;
  assign n1696 = n1688 & n1692 ;
  assign n1697 = ~n1682 & n1696 ;
  assign n1698 = ~n1695 & ~n1697 ;
  assign n1699 = ~n1694 & n1698 ;
  assign n1700 = n1688 & ~n1691 ;
  assign n1701 = ~n1682 & n1700 ;
  assign n1702 = n1677 & ~n1691 ;
  assign n1703 = ~\a[122]  & ~\b[122]  ;
  assign n1704 = \a[122]  & \b[122]  ;
  assign n1705 = ~n1703 & ~n1704 ;
  assign n1706 = ~n1690 & ~n1705 ;
  assign n1707 = ~n1702 & n1706 ;
  assign n1708 = ~n1701 & n1707 ;
  assign n1709 = ~n1690 & ~n1702 ;
  assign n1710 = ~n1701 & n1709 ;
  assign n1711 = n1705 & ~n1710 ;
  assign n1712 = ~n1708 & ~n1711 ;
  assign n1713 = ~\a[123]  & ~\b[123]  ;
  assign n1714 = \a[123]  & \b[123]  ;
  assign n1715 = ~n1713 & ~n1714 ;
  assign n1716 = ~n1690 & ~n1703 ;
  assign n1717 = ~n1702 & n1716 ;
  assign n1718 = ~n1701 & n1717 ;
  assign n1719 = ~n1704 & ~n1718 ;
  assign n1720 = ~n1715 & ~n1719 ;
  assign n1721 = ~n1704 & n1715 ;
  assign n1722 = ~n1718 & n1721 ;
  assign n1723 = ~n1720 & ~n1722 ;
  assign n1724 = ~n1704 & ~n1714 ;
  assign n1725 = ~n1718 & n1724 ;
  assign n1726 = ~\a[124]  & ~\b[124]  ;
  assign n1727 = \a[124]  & \b[124]  ;
  assign n1728 = ~n1726 & ~n1727 ;
  assign n1729 = ~n1713 & ~n1728 ;
  assign n1730 = ~n1725 & n1729 ;
  assign n1731 = n1713 & n1728 ;
  assign n1732 = n1724 & n1728 ;
  assign n1733 = ~n1718 & n1732 ;
  assign n1734 = ~n1731 & ~n1733 ;
  assign n1735 = ~n1730 & n1734 ;
  assign n1736 = n1724 & ~n1727 ;
  assign n1737 = ~n1718 & n1736 ;
  assign n1738 = n1713 & ~n1727 ;
  assign n1739 = ~\a[125]  & ~\b[125]  ;
  assign n1740 = \a[125]  & \b[125]  ;
  assign n1741 = ~n1739 & ~n1740 ;
  assign n1742 = ~n1726 & ~n1741 ;
  assign n1743 = ~n1738 & n1742 ;
  assign n1744 = ~n1737 & n1743 ;
  assign n1745 = ~n1726 & ~n1738 ;
  assign n1746 = ~n1737 & n1745 ;
  assign n1747 = n1741 & ~n1746 ;
  assign n1748 = ~n1744 & ~n1747 ;
  assign n1749 = ~\a[126]  & ~\b[126]  ;
  assign n1750 = \a[126]  & \b[126]  ;
  assign n1751 = ~n1749 & ~n1750 ;
  assign n1752 = ~n1726 & ~n1739 ;
  assign n1753 = ~n1738 & n1752 ;
  assign n1754 = ~n1737 & n1753 ;
  assign n1755 = ~n1740 & ~n1754 ;
  assign n1756 = ~n1751 & ~n1755 ;
  assign n1757 = ~n1740 & n1751 ;
  assign n1758 = ~n1754 & n1757 ;
  assign n1759 = ~n1756 & ~n1758 ;
  assign n1760 = ~n1740 & ~n1750 ;
  assign n1761 = ~n1754 & n1760 ;
  assign n1762 = ~\a[127]  & ~\b[127]  ;
  assign n1763 = \a[127]  & \b[127]  ;
  assign n1764 = ~n1762 & ~n1763 ;
  assign n1765 = ~n1749 & n1764 ;
  assign n1766 = ~n1761 & n1765 ;
  assign n1767 = ~n1749 & ~n1761 ;
  assign n1768 = ~n1764 & ~n1767 ;
  assign n1769 = ~n1766 & ~n1768 ;
  assign n1770 = n1760 & ~n1763 ;
  assign n1771 = ~n1754 & n1770 ;
  assign n1772 = n1749 & ~n1763 ;
  assign n1773 = ~n1762 & ~n1772 ;
  assign n1774 = ~n1771 & n1773 ;
  assign \f[0]  = n259 ;
  assign \f[1]  = n265 ;
  assign \f[2]  = n273 ;
  assign \f[3]  = ~n283 ;
  assign \f[4]  = ~n295 ;
  assign \f[5]  = ~n308 ;
  assign \f[6]  = ~n319 ;
  assign \f[7]  = ~n331 ;
  assign \f[8]  = ~n344 ;
  assign \f[9]  = ~n355 ;
  assign \f[10]  = ~n367 ;
  assign \f[11]  = ~n380 ;
  assign \f[12]  = ~n391 ;
  assign \f[13]  = ~n403 ;
  assign \f[14]  = ~n416 ;
  assign \f[15]  = ~n427 ;
  assign \f[16]  = ~n439 ;
  assign \f[17]  = ~n452 ;
  assign \f[18]  = ~n463 ;
  assign \f[19]  = ~n475 ;
  assign \f[20]  = ~n488 ;
  assign \f[21]  = ~n499 ;
  assign \f[22]  = ~n511 ;
  assign \f[23]  = ~n524 ;
  assign \f[24]  = ~n535 ;
  assign \f[25]  = ~n547 ;
  assign \f[26]  = ~n560 ;
  assign \f[27]  = ~n571 ;
  assign \f[28]  = ~n583 ;
  assign \f[29]  = ~n596 ;
  assign \f[30]  = ~n607 ;
  assign \f[31]  = ~n619 ;
  assign \f[32]  = ~n632 ;
  assign \f[33]  = ~n643 ;
  assign \f[34]  = ~n655 ;
  assign \f[35]  = ~n668 ;
  assign \f[36]  = ~n679 ;
  assign \f[37]  = ~n691 ;
  assign \f[38]  = ~n704 ;
  assign \f[39]  = ~n715 ;
  assign \f[40]  = ~n727 ;
  assign \f[41]  = ~n740 ;
  assign \f[42]  = ~n751 ;
  assign \f[43]  = ~n763 ;
  assign \f[44]  = ~n776 ;
  assign \f[45]  = ~n787 ;
  assign \f[46]  = ~n799 ;
  assign \f[47]  = ~n812 ;
  assign \f[48]  = ~n823 ;
  assign \f[49]  = ~n835 ;
  assign \f[50]  = ~n848 ;
  assign \f[51]  = ~n859 ;
  assign \f[52]  = ~n871 ;
  assign \f[53]  = ~n884 ;
  assign \f[54]  = ~n895 ;
  assign \f[55]  = ~n907 ;
  assign \f[56]  = ~n920 ;
  assign \f[57]  = ~n931 ;
  assign \f[58]  = ~n943 ;
  assign \f[59]  = ~n956 ;
  assign \f[60]  = ~n967 ;
  assign \f[61]  = ~n979 ;
  assign \f[62]  = ~n992 ;
  assign \f[63]  = ~n1003 ;
  assign \f[64]  = ~n1015 ;
  assign \f[65]  = ~n1028 ;
  assign \f[66]  = ~n1039 ;
  assign \f[67]  = ~n1051 ;
  assign \f[68]  = ~n1064 ;
  assign \f[69]  = ~n1075 ;
  assign \f[70]  = ~n1087 ;
  assign \f[71]  = ~n1100 ;
  assign \f[72]  = ~n1111 ;
  assign \f[73]  = ~n1123 ;
  assign \f[74]  = ~n1136 ;
  assign \f[75]  = ~n1147 ;
  assign \f[76]  = ~n1159 ;
  assign \f[77]  = ~n1172 ;
  assign \f[78]  = ~n1183 ;
  assign \f[79]  = ~n1195 ;
  assign \f[80]  = ~n1208 ;
  assign \f[81]  = ~n1219 ;
  assign \f[82]  = ~n1231 ;
  assign \f[83]  = ~n1244 ;
  assign \f[84]  = ~n1255 ;
  assign \f[85]  = ~n1267 ;
  assign \f[86]  = ~n1280 ;
  assign \f[87]  = ~n1291 ;
  assign \f[88]  = ~n1303 ;
  assign \f[89]  = ~n1316 ;
  assign \f[90]  = ~n1327 ;
  assign \f[91]  = ~n1339 ;
  assign \f[92]  = ~n1352 ;
  assign \f[93]  = ~n1363 ;
  assign \f[94]  = ~n1375 ;
  assign \f[95]  = ~n1388 ;
  assign \f[96]  = ~n1399 ;
  assign \f[97]  = ~n1411 ;
  assign \f[98]  = ~n1424 ;
  assign \f[99]  = ~n1435 ;
  assign \f[100]  = ~n1447 ;
  assign \f[101]  = ~n1460 ;
  assign \f[102]  = ~n1471 ;
  assign \f[103]  = ~n1483 ;
  assign \f[104]  = ~n1496 ;
  assign \f[105]  = ~n1507 ;
  assign \f[106]  = ~n1519 ;
  assign \f[107]  = ~n1532 ;
  assign \f[108]  = ~n1543 ;
  assign \f[109]  = ~n1555 ;
  assign \f[110]  = ~n1568 ;
  assign \f[111]  = ~n1579 ;
  assign \f[112]  = ~n1591 ;
  assign \f[113]  = ~n1604 ;
  assign \f[114]  = ~n1615 ;
  assign \f[115]  = ~n1627 ;
  assign \f[116]  = ~n1640 ;
  assign \f[117]  = ~n1651 ;
  assign \f[118]  = ~n1663 ;
  assign \f[119]  = ~n1676 ;
  assign \f[120]  = ~n1687 ;
  assign \f[121]  = ~n1699 ;
  assign \f[122]  = ~n1712 ;
  assign \f[123]  = ~n1723 ;
  assign \f[124]  = ~n1735 ;
  assign \f[125]  = ~n1748 ;
  assign \f[126]  = ~n1759 ;
  assign \f[127]  = n1769 ;
  assign cOut = n1774 ;
endmodule
