module top( \A[0]  , \A[1]  , \A[2]  , \A[3]  , \A[4]  , \A[5]  , \A[6]  , \A[7]  , \A[8]  , \A[9]  , \A[10]  , \A[11]  , \A[12]  , \A[13]  , \A[14]  , \A[15]  , \A[16]  , \A[17]  , \A[18]  , \A[19]  , \A[20]  , \A[21]  , \A[22]  , \A[23]  , \A[24]  , \A[25]  , \A[26]  , \A[27]  , \A[28]  , \A[29]  , \A[30]  , \A[31]  , \A[32]  , \A[33]  , \A[34]  , \A[35]  , \A[36]  , \A[37]  , \A[38]  , \A[39]  , \A[40]  , \A[41]  , \A[42]  , \A[43]  , \A[44]  , \A[45]  , \A[46]  , \A[47]  , \A[48]  , \A[49]  , \A[50]  , \A[51]  , \A[52]  , \A[53]  , \A[54]  , \A[55]  , \A[56]  , \A[57]  , \A[58]  , \A[59]  , \A[60]  , \A[61]  , \A[62]  , \A[63]  , \A[64]  , \A[65]  , \A[66]  , \A[67]  , \A[68]  , \A[69]  , \A[70]  , \A[71]  , \A[72]  , \A[73]  , \A[74]  , \A[75]  , \A[76]  , \A[77]  , \A[78]  , \A[79]  , \A[80]  , \A[81]  , \A[82]  , \A[83]  , \A[84]  , \A[85]  , \A[86]  , \A[87]  , \A[88]  , \A[89]  , \A[90]  , \A[91]  , \A[92]  , \A[93]  , \A[94]  , \A[95]  , \A[96]  , \A[97]  , \A[98]  , \A[99]  , \A[100]  , \A[101]  , \A[102]  , \A[103]  , \A[104]  , \A[105]  , \A[106]  , \A[107]  , \A[108]  , \A[109]  , \A[110]  , \A[111]  , \A[112]  , \A[113]  , \A[114]  , \A[115]  , \A[116]  , \A[117]  , \A[118]  , \A[119]  , \A[120]  , \A[121]  , \A[122]  , \A[123]  , \A[124]  , \A[125]  , \A[126]  , \A[127]  , \P[0]  , \P[1]  , \P[2]  , \P[3]  , \P[4]  , \P[5]  , \P[6]  , F );
  input \A[0]  ;
  input \A[1]  ;
  input \A[2]  ;
  input \A[3]  ;
  input \A[4]  ;
  input \A[5]  ;
  input \A[6]  ;
  input \A[7]  ;
  input \A[8]  ;
  input \A[9]  ;
  input \A[10]  ;
  input \A[11]  ;
  input \A[12]  ;
  input \A[13]  ;
  input \A[14]  ;
  input \A[15]  ;
  input \A[16]  ;
  input \A[17]  ;
  input \A[18]  ;
  input \A[19]  ;
  input \A[20]  ;
  input \A[21]  ;
  input \A[22]  ;
  input \A[23]  ;
  input \A[24]  ;
  input \A[25]  ;
  input \A[26]  ;
  input \A[27]  ;
  input \A[28]  ;
  input \A[29]  ;
  input \A[30]  ;
  input \A[31]  ;
  input \A[32]  ;
  input \A[33]  ;
  input \A[34]  ;
  input \A[35]  ;
  input \A[36]  ;
  input \A[37]  ;
  input \A[38]  ;
  input \A[39]  ;
  input \A[40]  ;
  input \A[41]  ;
  input \A[42]  ;
  input \A[43]  ;
  input \A[44]  ;
  input \A[45]  ;
  input \A[46]  ;
  input \A[47]  ;
  input \A[48]  ;
  input \A[49]  ;
  input \A[50]  ;
  input \A[51]  ;
  input \A[52]  ;
  input \A[53]  ;
  input \A[54]  ;
  input \A[55]  ;
  input \A[56]  ;
  input \A[57]  ;
  input \A[58]  ;
  input \A[59]  ;
  input \A[60]  ;
  input \A[61]  ;
  input \A[62]  ;
  input \A[63]  ;
  input \A[64]  ;
  input \A[65]  ;
  input \A[66]  ;
  input \A[67]  ;
  input \A[68]  ;
  input \A[69]  ;
  input \A[70]  ;
  input \A[71]  ;
  input \A[72]  ;
  input \A[73]  ;
  input \A[74]  ;
  input \A[75]  ;
  input \A[76]  ;
  input \A[77]  ;
  input \A[78]  ;
  input \A[79]  ;
  input \A[80]  ;
  input \A[81]  ;
  input \A[82]  ;
  input \A[83]  ;
  input \A[84]  ;
  input \A[85]  ;
  input \A[86]  ;
  input \A[87]  ;
  input \A[88]  ;
  input \A[89]  ;
  input \A[90]  ;
  input \A[91]  ;
  input \A[92]  ;
  input \A[93]  ;
  input \A[94]  ;
  input \A[95]  ;
  input \A[96]  ;
  input \A[97]  ;
  input \A[98]  ;
  input \A[99]  ;
  input \A[100]  ;
  input \A[101]  ;
  input \A[102]  ;
  input \A[103]  ;
  input \A[104]  ;
  input \A[105]  ;
  input \A[106]  ;
  input \A[107]  ;
  input \A[108]  ;
  input \A[109]  ;
  input \A[110]  ;
  input \A[111]  ;
  input \A[112]  ;
  input \A[113]  ;
  input \A[114]  ;
  input \A[115]  ;
  input \A[116]  ;
  input \A[117]  ;
  input \A[118]  ;
  input \A[119]  ;
  input \A[120]  ;
  input \A[121]  ;
  input \A[122]  ;
  input \A[123]  ;
  input \A[124]  ;
  input \A[125]  ;
  input \A[126]  ;
  input \A[127]  ;
  output \P[0]  ;
  output \P[1]  ;
  output \P[2]  ;
  output \P[3]  ;
  output \P[4]  ;
  output \P[5]  ;
  output \P[6]  ;
  output F ;
  wire n129 , n130 , n131 , n132 , n133 , n134 , n135 , n136 , n137 , n138 , n139 , n140 , n141 , n142 , n143 , n144 , n145 , n146 , n147 , n148 , n149 , n150 , n151 , n152 , n153 , n154 , n155 , n156 , n157 , n158 , n159 , n160 , n161 , n162 , n163 , n164 , n165 , n166 , n167 , n168 , n169 , n170 , n171 , n172 , n173 , n174 , n175 , n176 , n177 , n178 , n179 , n180 , n181 , n182 , n183 , n184 , n185 , n186 , n187 , n188 , n189 , n190 , n191 , n192 , n193 , n194 , n195 , n196 , n197 , n198 , n199 , n200 , n201 , n202 , n203 , n204 , n205 , n206 , n207 , n208 , n209 , n210 , n211 , n212 , n213 , n214 , n215 , n216 , n217 , n218 , n219 , n220 , n221 , n222 , n223 , n224 , n225 , n226 , n227 , n228 , n229 , n230 , n231 , n232 , n233 , n234 , n235 , n236 , n237 , n238 , n239 , n240 , n241 , n242 , n243 , n244 , n245 , n246 , n247 , n248 , n249 , n250 , n251 , n252 , n253 , n254 , n255 , n256 , n257 , n258 , n259 , n260 , n261 , n262 , n263 , n264 , n265 , n266 , n267 , n268 , n269 , n270 , n271 , n272 , n273 , n274 , n275 , n276 , n277 , n278 , n279 , n280 , n281 , n282 , n283 , n284 , n285 , n286 , n287 , n288 , n289 , n290 , n291 , n292 , n293 , n294 , n295 , n296 , n297 , n298 , n299 , n300 , n301 , n302 , n303 , n304 , n305 , n306 , n307 , n308 , n309 , n310 , n311 , n312 , n313 , n314 , n315 , n316 , n317 , n318 , n319 , n320 , n321 , n322 , n323 , n324 , n325 , n326 , n327 , n328 , n329 , n330 , n331 , n332 , n333 , n334 , n335 , n336 , n337 , n338 , n339 , n340 , n341 , n342 , n343 , n344 , n345 , n346 , n347 , n348 , n349 , n350 , n351 , n352 , n353 , n354 , n355 , n356 , n357 , n358 , n359 , n360 , n361 , n362 , n363 , n364 , n365 , n366 , n367 , n368 , n369 , n370 , n371 , n372 , n373 , n374 , n375 , n376 , n377 , n378 , n379 , n380 , n381 , n382 , n383 , n384 , n385 , n386 , n387 , n388 , n389 , n390 , n391 , n392 , n393 , n394 , n395 , n396 , n397 , n398 , n399 , n400 , n401 , n402 , n403 , n404 , n405 , n406 , n407 , n408 , n409 , n410 , n411 , n412 , n413 , n414 , n415 , n416 , n417 , n418 , n419 , n420 , n421 , n422 , n423 , n424 , n425 , n426 , n427 , n428 , n429 , n430 , n431 , n432 , n433 , n434 , n435 , n436 , n437 , n438 , n439 , n440 , n441 , n442 , n443 , n444 , n445 , n446 , n447 , n448 , n449 , n450 , n451 , n452 , n453 , n454 , n455 , n456 , n457 , n458 , n459 , n460 , n461 , n462 , n463 , n464 , n465 , n466 , n467 , n468 , n469 , n470 , n471 , n472 , n473 , n474 , n475 , n476 , n477 , n478 , n479 , n480 , n481 , n482 , n483 , n484 , n485 , n486 , n487 , n488 , n489 , n490 , n491 , n492 , n493 , n494 , n495 , n496 , n497 , n498 , n499 , n500 , n501 , n502 , n503 , n504 , n505 , n506 , n507 , n508 , n509 , n510 , n511 , n512 , n513 , n514 , n515 , n516 , n517 , n518 , n519 , n520 , n521 , n522 , n523 , n524 , n525 , n526 , n527 , n528 , n529 , n530 , n531 , n532 , n533 , n534 , n535 , n536 , n537 , n538 , n539 , n540 , n541 , n542 , n543 , n544 , n545 , n546 , n547 , n548 , n549 , n550 , n551 , n552 , n553 , n554 , n555 , n556 , n557 , n558 , n559 , n560 , n561 , n562 , n563 , n564 , n565 , n566 , n567 , n568 , n569 , n570 , n571 , n572 , n573 , n574 , n575 , n576 , n577 , n578 , n579 , n580 , n581 , n582 , n583 , n584 , n585 , n586 , n587 , n588 , n589 , n590 , n591 , n592 , n593 , n594 , n595 , n596 , n597 , n598 , n599 , n600 , n601 , n602 , n603 , n604 , n605 , n606 , n607 , n608 , n609 , n610 , n611 , n612 , n613 , n614 , n615 , n616 , n617 , n618 , n619 , n620 , n621 , n622 , n623 , n624 , n625 , n626 , n627 , n628 , n629 , n630 , n631 , n632 , n633 , n634 , n635 , n636 , n637 , n638 , n639 , n640 , n641 , n642 , n643 , n644 , n645 , n646 , n647 , n648 , n649 , n650 , n651 , n652 , n653 , n654 , n655 , n656 , n657 , n658 , n659 , n660 , n661 , n662 , n663 , n664 , n665 , n666 , n667 , n668 , n669 , n670 ;
  assign n129 = \A[76]  & ~\A[77]  ;
  assign n130 = \A[73]  & ~\A[74]  ;
  assign n131 = ~\A[75]  & ~\A[77]  ;
  assign n132 = ~n130 & n131 ;
  assign n133 = ~n129 & ~n132 ;
  assign n134 = \A[64]  & ~\A[65]  ;
  assign n135 = ~\A[66]  & ~\A[68]  ;
  assign n136 = ~n134 & n135 ;
  assign n137 = \A[67]  & ~\A[68]  ;
  assign n138 = ~\A[69]  & ~\A[71]  ;
  assign n139 = ~n137 & n138 ;
  assign n140 = ~n136 & n139 ;
  assign n141 = \A[55]  & ~\A[56]  ;
  assign n142 = ~\A[57]  & ~\A[59]  ;
  assign n143 = ~n141 & n142 ;
  assign n144 = \A[58]  & ~\A[59]  ;
  assign n145 = ~\A[60]  & ~\A[62]  ;
  assign n146 = ~n144 & n145 ;
  assign n147 = ~n143 & n146 ;
  assign n148 = \A[46]  & ~\A[47]  ;
  assign n149 = ~\A[48]  & ~\A[50]  ;
  assign n150 = ~n148 & n149 ;
  assign n151 = \A[49]  & ~\A[50]  ;
  assign n152 = ~\A[51]  & ~\A[53]  ;
  assign n153 = ~n151 & n152 ;
  assign n154 = ~n150 & n153 ;
  assign n155 = \A[37]  & ~\A[38]  ;
  assign n156 = ~\A[39]  & ~\A[41]  ;
  assign n157 = ~n155 & n156 ;
  assign n158 = \A[40]  & ~\A[41]  ;
  assign n159 = ~\A[42]  & ~\A[44]  ;
  assign n160 = ~n158 & n159 ;
  assign n161 = ~n157 & n160 ;
  assign n162 = \A[28]  & ~\A[29]  ;
  assign n163 = ~\A[30]  & ~\A[32]  ;
  assign n164 = ~n162 & n163 ;
  assign n165 = \A[31]  & ~\A[32]  ;
  assign n166 = ~\A[33]  & ~\A[35]  ;
  assign n167 = ~n165 & n166 ;
  assign n168 = ~n164 & n167 ;
  assign n169 = \A[19]  & ~\A[20]  ;
  assign n170 = ~\A[21]  & ~\A[23]  ;
  assign n171 = ~n169 & n170 ;
  assign n172 = \A[22]  & ~\A[23]  ;
  assign n173 = ~\A[24]  & ~\A[26]  ;
  assign n174 = ~n172 & n173 ;
  assign n175 = ~n171 & n174 ;
  assign n176 = \A[10]  & ~\A[11]  ;
  assign n177 = ~\A[12]  & ~\A[14]  ;
  assign n178 = ~n176 & n177 ;
  assign n179 = \A[13]  & ~\A[14]  ;
  assign n180 = ~\A[15]  & ~\A[17]  ;
  assign n181 = ~n179 & n180 ;
  assign n182 = ~n178 & n181 ;
  assign n183 = \A[1]  & ~\A[2]  ;
  assign n184 = ~\A[3]  & ~\A[5]  ;
  assign n185 = ~n183 & n184 ;
  assign n186 = \A[4]  & ~\A[5]  ;
  assign n187 = ~\A[6]  & ~\A[8]  ;
  assign n188 = ~n186 & n187 ;
  assign n189 = ~n185 & n188 ;
  assign n190 = \A[7]  & ~\A[8]  ;
  assign n191 = ~\A[9]  & ~\A[11]  ;
  assign n192 = ~n190 & n191 ;
  assign n193 = n181 & n192 ;
  assign n194 = ~n189 & n193 ;
  assign n195 = ~n182 & ~n194 ;
  assign n196 = \A[16]  & ~\A[17]  ;
  assign n197 = ~\A[18]  & ~\A[20]  ;
  assign n198 = ~n196 & n197 ;
  assign n199 = n174 & n198 ;
  assign n200 = n195 & n199 ;
  assign n201 = ~n175 & ~n200 ;
  assign n202 = \A[25]  & ~\A[26]  ;
  assign n203 = ~\A[27]  & ~\A[29]  ;
  assign n204 = ~n202 & n203 ;
  assign n205 = n167 & n204 ;
  assign n206 = n201 & n205 ;
  assign n207 = ~n168 & ~n206 ;
  assign n208 = \A[34]  & ~\A[35]  ;
  assign n209 = ~\A[36]  & ~\A[38]  ;
  assign n210 = ~n208 & n209 ;
  assign n211 = n160 & n210 ;
  assign n212 = n207 & n211 ;
  assign n213 = ~n161 & ~n212 ;
  assign n214 = \A[43]  & ~\A[44]  ;
  assign n215 = ~\A[45]  & ~\A[47]  ;
  assign n216 = ~n214 & n215 ;
  assign n217 = n153 & n216 ;
  assign n218 = n213 & n217 ;
  assign n219 = ~n154 & ~n218 ;
  assign n220 = \A[52]  & ~\A[53]  ;
  assign n221 = ~\A[54]  & ~\A[56]  ;
  assign n222 = ~n220 & n221 ;
  assign n223 = n146 & n222 ;
  assign n224 = n219 & n223 ;
  assign n225 = ~n147 & ~n224 ;
  assign n226 = \A[61]  & ~\A[62]  ;
  assign n227 = ~\A[63]  & ~\A[65]  ;
  assign n228 = ~n226 & n227 ;
  assign n229 = n139 & n228 ;
  assign n230 = n225 & n229 ;
  assign n231 = ~n140 & ~n230 ;
  assign n232 = \A[70]  & ~\A[71]  ;
  assign n233 = ~\A[72]  & ~\A[74]  ;
  assign n234 = ~n232 & n233 ;
  assign n235 = ~n129 & n234 ;
  assign n236 = n231 & n235 ;
  assign n237 = ~n133 & ~n236 ;
  assign n238 = ~\A[78]  & ~\A[80]  ;
  assign n239 = ~n237 & n238 ;
  assign n240 = \A[79]  & ~\A[80]  ;
  assign n241 = ~\A[81]  & ~\A[83]  ;
  assign n242 = ~n240 & n241 ;
  assign n243 = ~n239 & n242 ;
  assign n244 = \A[82]  & ~\A[83]  ;
  assign n245 = ~\A[84]  & ~n244 ;
  assign n246 = ~n243 & n245 ;
  assign n247 = \A[126]  & ~\A[127]  ;
  assign n248 = \A[120]  & ~\A[121]  ;
  assign n249 = ~\A[122]  & ~\A[124]  ;
  assign n250 = ~n248 & n249 ;
  assign n251 = \A[123]  & ~\A[124]  ;
  assign n252 = ~\A[125]  & ~\A[127]  ;
  assign n253 = ~n251 & n252 ;
  assign n254 = ~n250 & n253 ;
  assign n255 = \A[111]  & ~\A[112]  ;
  assign n256 = ~\A[113]  & ~\A[115]  ;
  assign n257 = ~n255 & n256 ;
  assign n258 = \A[114]  & ~\A[115]  ;
  assign n259 = ~\A[116]  & ~\A[118]  ;
  assign n260 = ~n258 & n259 ;
  assign n261 = ~n257 & n260 ;
  assign n262 = \A[102]  & ~\A[103]  ;
  assign n263 = ~\A[104]  & ~\A[106]  ;
  assign n264 = ~n262 & n263 ;
  assign n265 = \A[105]  & ~\A[106]  ;
  assign n266 = ~\A[107]  & ~\A[109]  ;
  assign n267 = ~n265 & n266 ;
  assign n268 = ~n264 & n267 ;
  assign n269 = \A[93]  & ~\A[94]  ;
  assign n270 = ~\A[95]  & ~\A[97]  ;
  assign n271 = ~n269 & n270 ;
  assign n272 = \A[96]  & ~\A[97]  ;
  assign n273 = ~\A[98]  & ~\A[100]  ;
  assign n274 = ~n272 & n273 ;
  assign n275 = ~n271 & n274 ;
  assign n276 = ~\A[85]  & \A[87]  ;
  assign n277 = ~\A[88]  & n276 ;
  assign n278 = ~\A[89]  & ~n277 ;
  assign n279 = \A[86]  & ~\A[87]  ;
  assign n280 = \A[85]  & ~\A[88]  ;
  assign n281 = ~n279 & n280 ;
  assign n282 = ~\A[91]  & ~n281 ;
  assign n283 = n278 & n282 ;
  assign n284 = \A[90]  & ~\A[91]  ;
  assign n285 = ~\A[92]  & ~\A[94]  ;
  assign n286 = ~n284 & n285 ;
  assign n287 = n274 & n286 ;
  assign n288 = ~n283 & n287 ;
  assign n289 = ~n275 & ~n288 ;
  assign n290 = \A[99]  & ~\A[100]  ;
  assign n291 = ~\A[101]  & ~\A[103]  ;
  assign n292 = ~n290 & n291 ;
  assign n293 = n267 & n292 ;
  assign n294 = n289 & n293 ;
  assign n295 = ~n268 & ~n294 ;
  assign n296 = \A[108]  & ~\A[109]  ;
  assign n297 = ~\A[110]  & ~\A[112]  ;
  assign n298 = ~n296 & n297 ;
  assign n299 = n260 & n298 ;
  assign n300 = n295 & n299 ;
  assign n301 = ~n261 & ~n300 ;
  assign n302 = \A[117]  & ~\A[118]  ;
  assign n303 = ~\A[119]  & ~\A[121]  ;
  assign n304 = ~n302 & n303 ;
  assign n305 = n253 & n304 ;
  assign n306 = n301 & n305 ;
  assign n307 = ~n254 & ~n306 ;
  assign n308 = ~n247 & n307 ;
  assign n309 = ~n246 & n308 ;
  assign n310 = \A[116]  & ~\A[117]  ;
  assign n311 = ~\A[118]  & ~\A[120]  ;
  assign n312 = ~n310 & n311 ;
  assign n313 = \A[119]  & ~\A[120]  ;
  assign n314 = ~\A[121]  & ~\A[123]  ;
  assign n315 = ~n313 & n314 ;
  assign n316 = ~n312 & n315 ;
  assign n317 = \A[107]  & ~\A[108]  ;
  assign n318 = ~\A[109]  & ~\A[111]  ;
  assign n319 = ~n317 & n318 ;
  assign n320 = \A[110]  & ~\A[111]  ;
  assign n321 = ~\A[112]  & ~\A[114]  ;
  assign n322 = ~n320 & n321 ;
  assign n323 = ~n319 & n322 ;
  assign n324 = \A[98]  & ~\A[99]  ;
  assign n325 = \A[95]  & ~\A[96]  ;
  assign n326 = ~\A[97]  & ~\A[99]  ;
  assign n327 = ~n325 & n326 ;
  assign n328 = ~\A[100]  & ~\A[102]  ;
  assign n329 = ~n327 & n328 ;
  assign n330 = ~\A[88]  & ~\A[90]  ;
  assign n331 = ~n279 & n330 ;
  assign n332 = \A[89]  & ~\A[90]  ;
  assign n333 = ~\A[91]  & ~\A[93]  ;
  assign n334 = ~n332 & n333 ;
  assign n335 = ~n331 & n334 ;
  assign n336 = \A[92]  & ~\A[93]  ;
  assign n337 = ~\A[94]  & ~\A[96]  ;
  assign n338 = ~n336 & n337 ;
  assign n339 = n328 & n338 ;
  assign n340 = ~n335 & n339 ;
  assign n341 = ~n329 & ~n340 ;
  assign n342 = ~n324 & ~n341 ;
  assign n343 = \A[101]  & ~\A[102]  ;
  assign n344 = ~\A[103]  & ~\A[105]  ;
  assign n345 = ~n343 & n344 ;
  assign n346 = ~n342 & n345 ;
  assign n347 = \A[104]  & ~\A[105]  ;
  assign n348 = ~\A[106]  & ~\A[108]  ;
  assign n349 = ~n347 & n348 ;
  assign n350 = n322 & n349 ;
  assign n351 = ~n346 & n350 ;
  assign n352 = ~n323 & ~n351 ;
  assign n353 = \A[113]  & ~\A[114]  ;
  assign n354 = ~\A[115]  & ~\A[117]  ;
  assign n355 = ~n353 & n354 ;
  assign n356 = n315 & n355 ;
  assign n357 = n352 & n356 ;
  assign n358 = ~n316 & ~n357 ;
  assign n359 = \A[122]  & ~\A[123]  ;
  assign n360 = ~\A[124]  & ~\A[126]  ;
  assign n361 = ~n359 & n360 ;
  assign n362 = n358 & n361 ;
  assign n363 = \A[125]  & ~\A[126]  ;
  assign n364 = ~\A[127]  & ~n363 ;
  assign n365 = ~n362 & n364 ;
  assign n366 = n245 & ~n365 ;
  assign n367 = ~n243 & n366 ;
  assign n368 = ~n309 & ~n367 ;
  assign n369 = ~\A[124]  & ~\A[125]  ;
  assign n370 = ~\A[118]  & ~\A[119]  ;
  assign n371 = ~\A[120]  & ~\A[121]  ;
  assign n372 = ~n370 & n371 ;
  assign n373 = ~\A[112]  & ~\A[113]  ;
  assign n374 = ~\A[114]  & ~\A[115]  ;
  assign n375 = ~n373 & n374 ;
  assign n376 = ~\A[106]  & ~\A[107]  ;
  assign n377 = ~\A[108]  & ~\A[109]  ;
  assign n378 = ~n376 & n377 ;
  assign n379 = ~\A[100]  & ~\A[101]  ;
  assign n380 = ~\A[94]  & ~\A[95]  ;
  assign n381 = ~\A[96]  & ~\A[97]  ;
  assign n382 = ~n380 & n381 ;
  assign n383 = ~\A[84]  & ~\A[85]  ;
  assign n384 = ~\A[88]  & ~\A[89]  ;
  assign n385 = ~\A[82]  & ~\A[83]  ;
  assign n386 = n384 & ~n385 ;
  assign n387 = ~\A[76]  & ~\A[77]  ;
  assign n388 = ~\A[78]  & ~\A[79]  ;
  assign n389 = ~n387 & n388 ;
  assign n390 = ~\A[70]  & ~\A[71]  ;
  assign n391 = ~\A[72]  & ~\A[73]  ;
  assign n392 = ~n390 & n391 ;
  assign n393 = ~\A[64]  & ~\A[65]  ;
  assign n394 = ~\A[66]  & ~\A[67]  ;
  assign n395 = ~n393 & n394 ;
  assign n396 = ~\A[58]  & ~\A[59]  ;
  assign n397 = ~\A[60]  & ~\A[61]  ;
  assign n398 = ~n396 & n397 ;
  assign n399 = ~\A[52]  & ~\A[53]  ;
  assign n400 = ~\A[54]  & ~\A[55]  ;
  assign n401 = ~n399 & n400 ;
  assign n402 = ~\A[28]  & ~\A[29]  ;
  assign n403 = ~\A[26]  & ~\A[27]  ;
  assign n404 = n402 & ~n403 ;
  assign n405 = ~\A[22]  & ~\A[23]  ;
  assign n406 = ~\A[20]  & ~\A[21]  ;
  assign n407 = n405 & ~n406 ;
  assign n408 = ~\A[16]  & ~\A[17]  ;
  assign n409 = ~\A[14]  & ~\A[15]  ;
  assign n410 = n408 & ~n409 ;
  assign n411 = ~\A[10]  & ~\A[11]  ;
  assign n412 = ~\A[8]  & ~\A[9]  ;
  assign n413 = n411 & ~n412 ;
  assign n414 = ~\A[4]  & ~\A[5]  ;
  assign n415 = ~\A[2]  & ~\A[3]  ;
  assign n416 = n414 & ~n415 ;
  assign n417 = ~\A[6]  & ~\A[7]  ;
  assign n418 = n411 & n417 ;
  assign n419 = ~n416 & n418 ;
  assign n420 = ~n413 & ~n419 ;
  assign n421 = ~\A[12]  & ~\A[13]  ;
  assign n422 = n408 & n421 ;
  assign n423 = n420 & n422 ;
  assign n424 = ~n410 & ~n423 ;
  assign n425 = ~\A[18]  & ~\A[19]  ;
  assign n426 = n405 & n425 ;
  assign n427 = n424 & n426 ;
  assign n428 = ~n407 & ~n427 ;
  assign n429 = ~\A[24]  & ~\A[25]  ;
  assign n430 = n402 & n429 ;
  assign n431 = n428 & n430 ;
  assign n432 = ~n404 & ~n431 ;
  assign n433 = ~\A[36]  & ~\A[37]  ;
  assign n434 = ~\A[34]  & ~\A[35]  ;
  assign n435 = n433 & ~n434 ;
  assign n436 = ~\A[42]  & ~\A[43]  ;
  assign n437 = ~\A[38]  & ~\A[39]  ;
  assign n438 = n436 & n437 ;
  assign n439 = ~n435 & n438 ;
  assign n440 = ~\A[44]  & ~\A[45]  ;
  assign n441 = ~\A[40]  & ~\A[41]  ;
  assign n442 = n436 & ~n441 ;
  assign n443 = n440 & ~n442 ;
  assign n444 = ~n439 & n443 ;
  assign n445 = ~\A[46]  & ~\A[47]  ;
  assign n446 = ~\A[30]  & ~\A[31]  ;
  assign n447 = n445 & n446 ;
  assign n448 = ~n444 & n447 ;
  assign n449 = n432 & n448 ;
  assign n450 = ~\A[48]  & ~\A[49]  ;
  assign n451 = ~\A[32]  & ~\A[33]  ;
  assign n452 = n445 & ~n451 ;
  assign n453 = ~n444 & n452 ;
  assign n454 = n450 & ~n453 ;
  assign n455 = ~n449 & n454 ;
  assign n456 = n432 & n446 ;
  assign n457 = ~n433 & n437 ;
  assign n458 = n440 & n441 ;
  assign n459 = ~n457 & n458 ;
  assign n460 = ~n436 & n440 ;
  assign n461 = n445 & n451 ;
  assign n462 = ~n460 & n461 ;
  assign n463 = ~n459 & n462 ;
  assign n464 = ~n456 & n463 ;
  assign n465 = n455 & ~n464 ;
  assign n466 = ~\A[50]  & ~\A[51]  ;
  assign n467 = n400 & n466 ;
  assign n468 = ~n465 & n467 ;
  assign n469 = ~n401 & ~n468 ;
  assign n470 = ~\A[56]  & ~\A[57]  ;
  assign n471 = n397 & n470 ;
  assign n472 = n469 & n471 ;
  assign n473 = ~n398 & ~n472 ;
  assign n474 = ~\A[62]  & ~\A[63]  ;
  assign n475 = n394 & n474 ;
  assign n476 = n473 & n475 ;
  assign n477 = ~n395 & ~n476 ;
  assign n478 = ~\A[68]  & ~\A[69]  ;
  assign n479 = n391 & n478 ;
  assign n480 = n477 & n479 ;
  assign n481 = ~n392 & ~n480 ;
  assign n482 = ~\A[74]  & ~\A[75]  ;
  assign n483 = n388 & n482 ;
  assign n484 = n481 & n483 ;
  assign n485 = ~n389 & ~n484 ;
  assign n486 = ~\A[80]  & ~\A[81]  ;
  assign n487 = n384 & n486 ;
  assign n488 = n485 & n487 ;
  assign n489 = ~n386 & ~n488 ;
  assign n490 = n383 & ~n489 ;
  assign n491 = ~\A[86]  & ~\A[87]  ;
  assign n492 = n384 & ~n491 ;
  assign n493 = ~\A[90]  & ~\A[91]  ;
  assign n494 = ~n492 & n493 ;
  assign n495 = ~n490 & n494 ;
  assign n496 = ~\A[92]  & ~\A[93]  ;
  assign n497 = n381 & n496 ;
  assign n498 = ~n495 & n497 ;
  assign n499 = ~n382 & ~n498 ;
  assign n500 = n379 & ~n499 ;
  assign n501 = ~\A[98]  & ~\A[99]  ;
  assign n502 = n379 & ~n501 ;
  assign n503 = ~\A[102]  & ~\A[103]  ;
  assign n504 = ~n502 & n503 ;
  assign n505 = ~n500 & n504 ;
  assign n506 = ~\A[104]  & ~\A[105]  ;
  assign n507 = n377 & n506 ;
  assign n508 = ~n505 & n507 ;
  assign n509 = ~n378 & ~n508 ;
  assign n510 = ~\A[110]  & ~\A[111]  ;
  assign n511 = n374 & n510 ;
  assign n512 = n509 & n511 ;
  assign n513 = ~n375 & ~n512 ;
  assign n514 = ~\A[116]  & ~\A[117]  ;
  assign n515 = n371 & n514 ;
  assign n516 = n513 & n515 ;
  assign n517 = ~n372 & ~n516 ;
  assign n518 = n369 & ~n517 ;
  assign n519 = ~\A[126]  & ~\A[127]  ;
  assign n520 = ~\A[122]  & ~\A[123]  ;
  assign n521 = n369 & ~n520 ;
  assign n522 = n519 & ~n521 ;
  assign n523 = ~n518 & n522 ;
  assign n524 = n390 & n478 ;
  assign n525 = n393 & n394 ;
  assign n526 = n524 & ~n525 ;
  assign n527 = n396 & n470 ;
  assign n528 = n399 & n400 ;
  assign n529 = n527 & ~n528 ;
  assign n530 = n440 & n445 ;
  assign n531 = n436 & n441 ;
  assign n532 = n530 & ~n531 ;
  assign n533 = n434 & n451 ;
  assign n534 = n402 & n446 ;
  assign n535 = n533 & ~n534 ;
  assign n536 = n405 & n406 ;
  assign n537 = n408 & n425 ;
  assign n538 = n536 & ~n537 ;
  assign n539 = n411 & n412 ;
  assign n540 = n414 & n417 ;
  assign n541 = n539 & ~n540 ;
  assign n542 = n409 & n421 ;
  assign n543 = n536 & n542 ;
  assign n544 = ~n541 & n543 ;
  assign n545 = ~n538 & ~n544 ;
  assign n546 = n403 & n429 ;
  assign n547 = n533 & n546 ;
  assign n548 = n545 & n547 ;
  assign n549 = ~n535 & ~n548 ;
  assign n550 = n433 & n437 ;
  assign n551 = n530 & n550 ;
  assign n552 = n549 & n551 ;
  assign n553 = ~n532 & ~n552 ;
  assign n554 = n450 & n466 ;
  assign n555 = n527 & n554 ;
  assign n556 = n553 & n555 ;
  assign n557 = ~n529 & ~n556 ;
  assign n558 = n397 & n474 ;
  assign n559 = n524 & n558 ;
  assign n560 = n557 & n559 ;
  assign n561 = ~n526 & ~n560 ;
  assign n562 = n391 & n482 ;
  assign n563 = n561 & n562 ;
  assign n564 = n383 & n491 ;
  assign n565 = n384 & n493 ;
  assign n566 = ~n564 & n565 ;
  assign n567 = n380 & n496 ;
  assign n568 = n379 & n503 ;
  assign n569 = n567 & n568 ;
  assign n570 = ~n566 & n569 ;
  assign n571 = n376 & n506 ;
  assign n572 = n373 & n374 ;
  assign n573 = n571 & n572 ;
  assign n574 = n381 & n501 ;
  assign n575 = n568 & ~n574 ;
  assign n576 = n573 & ~n575 ;
  assign n577 = ~n570 & n576 ;
  assign n578 = n387 & n388 ;
  assign n579 = n370 & n514 ;
  assign n580 = n377 & n510 ;
  assign n581 = n572 & ~n580 ;
  assign n582 = n579 & ~n581 ;
  assign n583 = n578 & n582 ;
  assign n584 = ~n577 & n583 ;
  assign n585 = ~n563 & n584 ;
  assign n586 = ~n571 & n580 ;
  assign n587 = ~n567 & n574 ;
  assign n588 = n385 & n486 ;
  assign n589 = n564 & ~n588 ;
  assign n590 = n565 & n574 ;
  assign n591 = ~n589 & n590 ;
  assign n592 = ~n587 & ~n591 ;
  assign n593 = n568 & n580 ;
  assign n594 = n592 & n593 ;
  assign n595 = ~n586 & ~n594 ;
  assign n596 = n572 & n595 ;
  assign n597 = n562 & n579 ;
  assign n598 = ~n596 & n597 ;
  assign n599 = n561 & n598 ;
  assign n600 = n371 & n520 ;
  assign n601 = ~n578 & n579 ;
  assign n602 = ~n596 & n601 ;
  assign n603 = n600 & ~n602 ;
  assign n604 = ~n599 & n603 ;
  assign n605 = ~n585 & n604 ;
  assign n606 = n369 & n519 ;
  assign n607 = ~n605 & n606 ;
  assign n608 = n565 & n567 ;
  assign n609 = n564 & n588 ;
  assign n610 = n608 & ~n609 ;
  assign n611 = n524 & n525 ;
  assign n612 = n527 & n558 ;
  assign n613 = n611 & ~n612 ;
  assign n614 = n530 & n531 ;
  assign n615 = n533 & n550 ;
  assign n616 = n614 & ~n615 ;
  assign n617 = n536 & n537 ;
  assign n618 = n539 & n542 ;
  assign n619 = n617 & ~n618 ;
  assign n620 = n534 & n546 ;
  assign n621 = n614 & n620 ;
  assign n622 = ~n619 & n621 ;
  assign n623 = ~n616 & ~n622 ;
  assign n624 = n528 & n554 ;
  assign n625 = n611 & n624 ;
  assign n626 = n623 & n625 ;
  assign n627 = ~n613 & ~n626 ;
  assign n628 = n562 & n578 ;
  assign n629 = n608 & n628 ;
  assign n630 = n627 & n629 ;
  assign n631 = ~n610 & ~n630 ;
  assign n632 = n600 & n606 ;
  assign n633 = n572 & n579 ;
  assign n634 = n571 & n580 ;
  assign n635 = n568 & n574 ;
  assign n636 = n634 & ~n635 ;
  assign n637 = n633 & ~n636 ;
  assign n638 = n632 & ~n637 ;
  assign n639 = n631 & n638 ;
  assign n640 = n633 & ~n634 ;
  assign n641 = n632 & ~n640 ;
  assign n642 = ~n631 & n641 ;
  assign n643 = ~n639 & ~n642 ;
  assign n644 = n632 & n633 ;
  assign n645 = n608 & n609 ;
  assign n646 = n611 & n628 ;
  assign n647 = n645 & ~n646 ;
  assign n648 = n614 & n615 ;
  assign n649 = n617 & n620 ;
  assign n650 = n648 & ~n649 ;
  assign n651 = n612 & n624 ;
  assign n652 = n645 & n651 ;
  assign n653 = ~n650 & n652 ;
  assign n654 = ~n647 & ~n653 ;
  assign n655 = n634 & n635 ;
  assign n656 = n654 & n655 ;
  assign n657 = n644 & ~n656 ;
  assign n658 = n644 & n655 ;
  assign n659 = n648 & n651 ;
  assign n660 = n645 & n646 ;
  assign n661 = ~n659 & n660 ;
  assign n662 = n658 & ~n661 ;
  assign n663 = n658 & n660 ;
  assign n664 = ~\A[0]  & ~\A[1]  ;
  assign n665 = n415 & n664 ;
  assign n666 = n540 & n665 ;
  assign n667 = n618 & n666 ;
  assign n668 = n649 & n667 ;
  assign n669 = n659 & n668 ;
  assign n670 = n663 & n669 ;
  assign \P[0]  = ~n368 ;
  assign \P[1]  = ~n523 ;
  assign \P[2]  = ~n607 ;
  assign \P[3]  = n643 ;
  assign \P[4]  = ~n657 ;
  assign \P[5]  = ~n662 ;
  assign \P[6]  = ~n663 ;
  assign F = ~n670 ;
endmodule
