module top( \P1_B_reg/NET0131  , \P1_IR_reg[0]/NET0131  , \P1_IR_reg[10]/NET0131  , \P1_IR_reg[11]/NET0131  , \P1_IR_reg[12]/NET0131  , \P1_IR_reg[13]/NET0131  , \P1_IR_reg[14]/NET0131  , \P1_IR_reg[15]/NET0131  , \P1_IR_reg[16]/NET0131  , \P1_IR_reg[17]/NET0131  , \P1_IR_reg[18]/NET0131  , \P1_IR_reg[19]/NET0131  , \P1_IR_reg[1]/NET0131  , \P1_IR_reg[20]/NET0131  , \P1_IR_reg[21]/NET0131  , \P1_IR_reg[22]/NET0131  , \P1_IR_reg[23]/NET0131  , \P1_IR_reg[24]/NET0131  , \P1_IR_reg[25]/NET0131  , \P1_IR_reg[26]/NET0131  , \P1_IR_reg[27]/NET0131  , \P1_IR_reg[28]/NET0131  , \P1_IR_reg[29]/NET0131  , \P1_IR_reg[2]/NET0131  , \P1_IR_reg[30]/NET0131  , \P1_IR_reg[31]/NET0131  , \P1_IR_reg[3]/NET0131  , \P1_IR_reg[4]/NET0131  , \P1_IR_reg[5]/NET0131  , \P1_IR_reg[6]/NET0131  , \P1_IR_reg[7]/NET0131  , \P1_IR_reg[8]/NET0131  , \P1_IR_reg[9]/NET0131  , \P1_addr_reg[0]/NET0131  , \P1_addr_reg[10]/NET0131  , \P1_addr_reg[11]/NET0131  , \P1_addr_reg[12]/NET0131  , \P1_addr_reg[13]/NET0131  , \P1_addr_reg[14]/NET0131  , \P1_addr_reg[15]/NET0131  , \P1_addr_reg[16]/NET0131  , \P1_addr_reg[17]/NET0131  , \P1_addr_reg[18]/NET0131  , \P1_addr_reg[19]/NET0131  , \P1_addr_reg[1]/NET0131  , \P1_addr_reg[2]/NET0131  , \P1_addr_reg[3]/NET0131  , \P1_addr_reg[4]/NET0131  , \P1_addr_reg[5]/NET0131  , \P1_addr_reg[6]/NET0131  , \P1_addr_reg[7]/NET0131  , \P1_addr_reg[8]/NET0131  , \P1_addr_reg[9]/NET0131  , \P1_d_reg[0]/NET0131  , \P1_d_reg[1]/NET0131  , \P1_datao_reg[0]/NET0131  , \P1_datao_reg[10]/NET0131  , \P1_datao_reg[11]/NET0131  , \P1_datao_reg[12]/NET0131  , \P1_datao_reg[13]/NET0131  , \P1_datao_reg[14]/NET0131  , \P1_datao_reg[15]/NET0131  , \P1_datao_reg[16]/NET0131  , \P1_datao_reg[17]/NET0131  , \P1_datao_reg[18]/NET0131  , \P1_datao_reg[19]/NET0131  , \P1_datao_reg[1]/NET0131  , \P1_datao_reg[20]/NET0131  , \P1_datao_reg[21]/NET0131  , \P1_datao_reg[22]/NET0131  , \P1_datao_reg[23]/NET0131  , \P1_datao_reg[24]/NET0131  , \P1_datao_reg[25]/NET0131  , \P1_datao_reg[26]/NET0131  , \P1_datao_reg[27]/NET0131  , \P1_datao_reg[28]/NET0131  , \P1_datao_reg[29]/NET0131  , \P1_datao_reg[2]/NET0131  , \P1_datao_reg[30]/NET0131  , \P1_datao_reg[31]/NET0131  , \P1_datao_reg[3]/NET0131  , \P1_datao_reg[4]/NET0131  , \P1_datao_reg[5]/NET0131  , \P1_datao_reg[6]/NET0131  , \P1_datao_reg[7]/NET0131  , \P1_datao_reg[8]/NET0131  , \P1_datao_reg[9]/NET0131  , \P1_rd_reg/NET0131  , \P1_reg0_reg[0]/NET0131  , \P1_reg0_reg[10]/NET0131  , \P1_reg0_reg[11]/NET0131  , \P1_reg0_reg[12]/NET0131  , \P1_reg0_reg[13]/NET0131  , \P1_reg0_reg[14]/NET0131  , \P1_reg0_reg[15]/NET0131  , \P1_reg0_reg[16]/NET0131  , \P1_reg0_reg[17]/NET0131  , \P1_reg0_reg[18]/NET0131  , \P1_reg0_reg[19]/NET0131  , \P1_reg0_reg[1]/NET0131  , \P1_reg0_reg[20]/NET0131  , \P1_reg0_reg[21]/NET0131  , \P1_reg0_reg[22]/NET0131  , \P1_reg0_reg[23]/NET0131  , \P1_reg0_reg[24]/NET0131  , \P1_reg0_reg[25]/NET0131  , \P1_reg0_reg[26]/NET0131  , \P1_reg0_reg[27]/NET0131  , \P1_reg0_reg[28]/NET0131  , \P1_reg0_reg[29]/NET0131  , \P1_reg0_reg[2]/NET0131  , \P1_reg0_reg[30]/NET0131  , \P1_reg0_reg[31]/NET0131  , \P1_reg0_reg[3]/NET0131  , \P1_reg0_reg[4]/NET0131  , \P1_reg0_reg[5]/NET0131  , \P1_reg0_reg[6]/NET0131  , \P1_reg0_reg[7]/NET0131  , \P1_reg0_reg[8]/NET0131  , \P1_reg0_reg[9]/NET0131  , \P1_reg1_reg[0]/NET0131  , \P1_reg1_reg[10]/NET0131  , \P1_reg1_reg[11]/NET0131  , \P1_reg1_reg[12]/NET0131  , \P1_reg1_reg[13]/NET0131  , \P1_reg1_reg[14]/NET0131  , \P1_reg1_reg[15]/NET0131  , \P1_reg1_reg[16]/NET0131  , \P1_reg1_reg[17]/NET0131  , \P1_reg1_reg[18]/NET0131  , \P1_reg1_reg[19]/NET0131  , \P1_reg1_reg[1]/NET0131  , \P1_reg1_reg[20]/NET0131  , \P1_reg1_reg[21]/NET0131  , \P1_reg1_reg[22]/NET0131  , \P1_reg1_reg[23]/NET0131  , \P1_reg1_reg[24]/NET0131  , \P1_reg1_reg[25]/NET0131  , \P1_reg1_reg[26]/NET0131  , \P1_reg1_reg[27]/NET0131  , \P1_reg1_reg[28]/NET0131  , \P1_reg1_reg[29]/NET0131  , \P1_reg1_reg[2]/NET0131  , \P1_reg1_reg[30]/NET0131  , \P1_reg1_reg[31]/NET0131  , \P1_reg1_reg[3]/NET0131  , \P1_reg1_reg[4]/NET0131  , \P1_reg1_reg[5]/NET0131  , \P1_reg1_reg[6]/NET0131  , \P1_reg1_reg[7]/NET0131  , \P1_reg1_reg[8]/NET0131  , \P1_reg1_reg[9]/NET0131  , \P1_reg2_reg[0]/NET0131  , \P1_reg2_reg[10]/NET0131  , \P1_reg2_reg[11]/NET0131  , \P1_reg2_reg[12]/NET0131  , \P1_reg2_reg[13]/NET0131  , \P1_reg2_reg[14]/NET0131  , \P1_reg2_reg[15]/NET0131  , \P1_reg2_reg[16]/NET0131  , \P1_reg2_reg[17]/NET0131  , \P1_reg2_reg[18]/NET0131  , \P1_reg2_reg[19]/NET0131  , \P1_reg2_reg[1]/NET0131  , \P1_reg2_reg[20]/NET0131  , \P1_reg2_reg[21]/NET0131  , \P1_reg2_reg[22]/NET0131  , \P1_reg2_reg[23]/NET0131  , \P1_reg2_reg[24]/NET0131  , \P1_reg2_reg[25]/NET0131  , \P1_reg2_reg[26]/NET0131  , \P1_reg2_reg[27]/NET0131  , \P1_reg2_reg[28]/NET0131  , \P1_reg2_reg[29]/NET0131  , \P1_reg2_reg[2]/NET0131  , \P1_reg2_reg[30]/NET0131  , \P1_reg2_reg[31]/NET0131  , \P1_reg2_reg[3]/NET0131  , \P1_reg2_reg[4]/NET0131  , \P1_reg2_reg[5]/NET0131  , \P1_reg2_reg[6]/NET0131  , \P1_reg2_reg[7]/NET0131  , \P1_reg2_reg[8]/NET0131  , \P1_reg2_reg[9]/NET0131  , \P1_reg3_reg[0]/NET0131  , \P1_reg3_reg[10]/NET0131  , \P1_reg3_reg[11]/NET0131  , \P1_reg3_reg[12]/NET0131  , \P1_reg3_reg[13]/NET0131  , \P1_reg3_reg[14]/NET0131  , \P1_reg3_reg[15]/NET0131  , \P1_reg3_reg[16]/NET0131  , \P1_reg3_reg[17]/NET0131  , \P1_reg3_reg[18]/NET0131  , \P1_reg3_reg[19]/NET0131  , \P1_reg3_reg[1]/NET0131  , \P1_reg3_reg[20]/NET0131  , \P1_reg3_reg[21]/NET0131  , \P1_reg3_reg[22]/NET0131  , \P1_reg3_reg[23]/NET0131  , \P1_reg3_reg[24]/NET0131  , \P1_reg3_reg[25]/NET0131  , \P1_reg3_reg[26]/NET0131  , \P1_reg3_reg[27]/NET0131  , \P1_reg3_reg[28]/NET0131  , \P1_reg3_reg[2]/NET0131  , \P1_reg3_reg[3]/NET0131  , \P1_reg3_reg[4]/NET0131  , \P1_reg3_reg[5]/NET0131  , \P1_reg3_reg[6]/NET0131  , \P1_reg3_reg[7]/NET0131  , \P1_reg3_reg[8]/NET0131  , \P1_reg3_reg[9]/NET0131  , \P1_state_reg[0]/NET0131  , \P1_wr_reg/NET0131  , \P2_B_reg/NET0131  , \P2_IR_reg[0]/NET0131  , \P2_IR_reg[10]/NET0131  , \P2_IR_reg[11]/NET0131  , \P2_IR_reg[12]/NET0131  , \P2_IR_reg[13]/NET0131  , \P2_IR_reg[14]/NET0131  , \P2_IR_reg[15]/NET0131  , \P2_IR_reg[16]/NET0131  , \P2_IR_reg[17]/NET0131  , \P2_IR_reg[18]/NET0131  , \P2_IR_reg[19]/NET0131  , \P2_IR_reg[1]/NET0131  , \P2_IR_reg[20]/NET0131  , \P2_IR_reg[21]/NET0131  , \P2_IR_reg[22]/NET0131  , \P2_IR_reg[23]/NET0131  , \P2_IR_reg[24]/NET0131  , \P2_IR_reg[25]/NET0131  , \P2_IR_reg[26]/NET0131  , \P2_IR_reg[27]/NET0131  , \P2_IR_reg[28]/NET0131  , \P2_IR_reg[29]/NET0131  , \P2_IR_reg[2]/NET0131  , \P2_IR_reg[30]/NET0131  , \P2_IR_reg[31]/NET0131  , \P2_IR_reg[3]/NET0131  , \P2_IR_reg[4]/NET0131  , \P2_IR_reg[5]/NET0131  , \P2_IR_reg[6]/NET0131  , \P2_IR_reg[7]/NET0131  , \P2_IR_reg[8]/NET0131  , \P2_IR_reg[9]/NET0131  , \P2_addr_reg[0]/NET0131  , \P2_addr_reg[10]/NET0131  , \P2_addr_reg[11]/NET0131  , \P2_addr_reg[12]/NET0131  , \P2_addr_reg[13]/NET0131  , \P2_addr_reg[14]/NET0131  , \P2_addr_reg[15]/NET0131  , \P2_addr_reg[16]/NET0131  , \P2_addr_reg[17]/NET0131  , \P2_addr_reg[18]/NET0131  , \P2_addr_reg[19]/NET0131  , \P2_addr_reg[1]/NET0131  , \P2_addr_reg[2]/NET0131  , \P2_addr_reg[3]/NET0131  , \P2_addr_reg[4]/NET0131  , \P2_addr_reg[5]/NET0131  , \P2_addr_reg[6]/NET0131  , \P2_addr_reg[7]/NET0131  , \P2_addr_reg[8]/NET0131  , \P2_addr_reg[9]/NET0131  , \P2_d_reg[0]/NET0131  , \P2_d_reg[1]/NET0131  , \P2_datao_reg[0]/NET0131  , \P2_datao_reg[10]/NET0131  , \P2_datao_reg[11]/NET0131  , \P2_datao_reg[12]/NET0131  , \P2_datao_reg[13]/NET0131  , \P2_datao_reg[14]/NET0131  , \P2_datao_reg[15]/NET0131  , \P2_datao_reg[16]/NET0131  , \P2_datao_reg[17]/NET0131  , \P2_datao_reg[18]/NET0131  , \P2_datao_reg[19]/NET0131  , \P2_datao_reg[1]/NET0131  , \P2_datao_reg[20]/NET0131  , \P2_datao_reg[21]/NET0131  , \P2_datao_reg[22]/NET0131  , \P2_datao_reg[23]/NET0131  , \P2_datao_reg[24]/NET0131  , \P2_datao_reg[25]/NET0131  , \P2_datao_reg[26]/NET0131  , \P2_datao_reg[27]/NET0131  , \P2_datao_reg[28]/NET0131  , \P2_datao_reg[29]/NET0131  , \P2_datao_reg[2]/NET0131  , \P2_datao_reg[30]/NET0131  , \P2_datao_reg[31]/NET0131  , \P2_datao_reg[3]/NET0131  , \P2_datao_reg[4]/NET0131  , \P2_datao_reg[5]/NET0131  , \P2_datao_reg[6]/NET0131  , \P2_datao_reg[7]/NET0131  , \P2_datao_reg[8]/NET0131  , \P2_datao_reg[9]/NET0131  , \P2_rd_reg/NET0131  , \P2_reg0_reg[0]/NET0131  , \P2_reg0_reg[10]/NET0131  , \P2_reg0_reg[11]/NET0131  , \P2_reg0_reg[12]/NET0131  , \P2_reg0_reg[13]/NET0131  , \P2_reg0_reg[14]/NET0131  , \P2_reg0_reg[15]/NET0131  , \P2_reg0_reg[16]/NET0131  , \P2_reg0_reg[17]/NET0131  , \P2_reg0_reg[18]/NET0131  , \P2_reg0_reg[19]/NET0131  , \P2_reg0_reg[1]/NET0131  , \P2_reg0_reg[20]/NET0131  , \P2_reg0_reg[21]/NET0131  , \P2_reg0_reg[22]/NET0131  , \P2_reg0_reg[23]/NET0131  , \P2_reg0_reg[24]/NET0131  , \P2_reg0_reg[25]/NET0131  , \P2_reg0_reg[26]/NET0131  , \P2_reg0_reg[27]/NET0131  , \P2_reg0_reg[28]/NET0131  , \P2_reg0_reg[29]/NET0131  , \P2_reg0_reg[2]/NET0131  , \P2_reg0_reg[30]/NET0131  , \P2_reg0_reg[31]/NET0131  , \P2_reg0_reg[3]/NET0131  , \P2_reg0_reg[4]/NET0131  , \P2_reg0_reg[5]/NET0131  , \P2_reg0_reg[6]/NET0131  , \P2_reg0_reg[7]/NET0131  , \P2_reg0_reg[8]/NET0131  , \P2_reg0_reg[9]/NET0131  , \P2_reg1_reg[0]/NET0131  , \P2_reg1_reg[10]/NET0131  , \P2_reg1_reg[11]/NET0131  , \P2_reg1_reg[12]/NET0131  , \P2_reg1_reg[13]/NET0131  , \P2_reg1_reg[14]/NET0131  , \P2_reg1_reg[15]/NET0131  , \P2_reg1_reg[16]/NET0131  , \P2_reg1_reg[17]/NET0131  , \P2_reg1_reg[18]/NET0131  , \P2_reg1_reg[19]/NET0131  , \P2_reg1_reg[1]/NET0131  , \P2_reg1_reg[20]/NET0131  , \P2_reg1_reg[21]/NET0131  , \P2_reg1_reg[22]/NET0131  , \P2_reg1_reg[23]/NET0131  , \P2_reg1_reg[24]/NET0131  , \P2_reg1_reg[25]/NET0131  , \P2_reg1_reg[26]/NET0131  , \P2_reg1_reg[27]/NET0131  , \P2_reg1_reg[28]/NET0131  , \P2_reg1_reg[29]/NET0131  , \P2_reg1_reg[2]/NET0131  , \P2_reg1_reg[30]/NET0131  , \P2_reg1_reg[31]/NET0131  , \P2_reg1_reg[3]/NET0131  , \P2_reg1_reg[4]/NET0131  , \P2_reg1_reg[5]/NET0131  , \P2_reg1_reg[6]/NET0131  , \P2_reg1_reg[7]/NET0131  , \P2_reg1_reg[8]/NET0131  , \P2_reg1_reg[9]/NET0131  , \P2_reg2_reg[0]/NET0131  , \P2_reg2_reg[10]/NET0131  , \P2_reg2_reg[11]/NET0131  , \P2_reg2_reg[12]/NET0131  , \P2_reg2_reg[13]/NET0131  , \P2_reg2_reg[14]/NET0131  , \P2_reg2_reg[15]/NET0131  , \P2_reg2_reg[16]/NET0131  , \P2_reg2_reg[17]/NET0131  , \P2_reg2_reg[18]/NET0131  , \P2_reg2_reg[19]/NET0131  , \P2_reg2_reg[1]/NET0131  , \P2_reg2_reg[20]/NET0131  , \P2_reg2_reg[21]/NET0131  , \P2_reg2_reg[22]/NET0131  , \P2_reg2_reg[23]/NET0131  , \P2_reg2_reg[24]/NET0131  , \P2_reg2_reg[25]/NET0131  , \P2_reg2_reg[26]/NET0131  , \P2_reg2_reg[27]/NET0131  , \P2_reg2_reg[28]/NET0131  , \P2_reg2_reg[29]/NET0131  , \P2_reg2_reg[2]/NET0131  , \P2_reg2_reg[30]/NET0131  , \P2_reg2_reg[31]/NET0131  , \P2_reg2_reg[3]/NET0131  , \P2_reg2_reg[4]/NET0131  , \P2_reg2_reg[5]/NET0131  , \P2_reg2_reg[6]/NET0131  , \P2_reg2_reg[7]/NET0131  , \P2_reg2_reg[8]/NET0131  , \P2_reg2_reg[9]/NET0131  , \P2_reg3_reg[0]/NET0131  , \P2_reg3_reg[10]/NET0131  , \P2_reg3_reg[11]/NET0131  , \P2_reg3_reg[12]/NET0131  , \P2_reg3_reg[13]/NET0131  , \P2_reg3_reg[14]/NET0131  , \P2_reg3_reg[15]/NET0131  , \P2_reg3_reg[16]/NET0131  , \P2_reg3_reg[17]/NET0131  , \P2_reg3_reg[18]/NET0131  , \P2_reg3_reg[19]/NET0131  , \P2_reg3_reg[1]/NET0131  , \P2_reg3_reg[20]/NET0131  , \P2_reg3_reg[21]/NET0131  , \P2_reg3_reg[22]/NET0131  , \P2_reg3_reg[23]/NET0131  , \P2_reg3_reg[24]/NET0131  , \P2_reg3_reg[25]/NET0131  , \P2_reg3_reg[26]/NET0131  , \P2_reg3_reg[27]/NET0131  , \P2_reg3_reg[28]/NET0131  , \P2_reg3_reg[2]/NET0131  , \P2_reg3_reg[3]/NET0131  , \P2_reg3_reg[4]/NET0131  , \P2_reg3_reg[5]/NET0131  , \P2_reg3_reg[6]/NET0131  , \P2_reg3_reg[7]/NET0131  , \P2_reg3_reg[8]/NET0131  , \P2_reg3_reg[9]/NET0131  , \P2_wr_reg/NET0131  , \si[0]_pad  , \si[10]_pad  , \si[11]_pad  , \si[12]_pad  , \si[13]_pad  , \si[14]_pad  , \si[15]_pad  , \si[16]_pad  , \si[17]_pad  , \si[18]_pad  , \si[19]_pad  , \si[1]_pad  , \si[20]_pad  , \si[21]_pad  , \si[22]_pad  , \si[23]_pad  , \si[24]_pad  , \si[25]_pad  , \si[26]_pad  , \si[27]_pad  , \si[28]_pad  , \si[29]_pad  , \si[2]_pad  , \si[30]_pad  , \si[31]_pad  , \si[3]_pad  , \si[4]_pad  , \si[5]_pad  , \si[6]_pad  , \si[7]_pad  , \si[8]_pad  , \si[9]_pad  , \P1_state_reg[0]/NET0131_syn_2  , \_al_n0  , \_al_n1  , \g73521/_0_  , \g73537/_0_  , \g73538/_0_  , \g73539/_0_  , \g73540/_0_  , \g73570/_0_  , \g73571/_0_  , \g73572/_0_  , \g73573/_0_  , \g73574/_0_  , \g73575/_0_  , \g73576/_0_  , \g73577/_0_  , \g73578/_0_  , \g73579/_0_  , \g73609/_0_  , \g73610/_0_  , \g73611/_0_  , \g73613/_0_  , \g73614/_0_  , \g73615/_0_  , \g73617/_0_  , \g73618/_0_  , \g73619/_0_  , \g73620/_0_  , \g73621/_0_  , \g73622/_0_  , \g73623/_0_  , \g73624/_0_  , \g73625/_0_  , \g73626/_0_  , \g73627/_0_  , \g73628/_0_  , \g73629/_0_  , \g73630/_0_  , \g73631/_0_  , \g73632/_0_  , \g73633/_0_  , \g73692/_0_  , \g73693/_0_  , \g73694/_0_  , \g73696/_0_  , \g73697/_0_  , \g73703/_0_  , \g73704/_0_  , \g73709/_0_  , \g73710/_0_  , \g73711/_0_  , \g73712/_0_  , \g73713/_0_  , \g73714/_0_  , \g73715/_0_  , \g73716/_0_  , \g73717/_0_  , \g73718/_0_  , \g73719/_0_  , \g73720/_0_  , \g73774/_0_  , \g73775/_0_  , \g73776/_0_  , \g73777/_0_  , \g73806/_0_  , \g73807/_0_  , \g73808/_0_  , \g73809/_0_  , \g73810/_0_  , \g73811/_0_  , \g73812/_0_  , \g73813/_0_  , \g73814/_0_  , \g73815/_0_  , \g73816/_0_  , \g73817/_0_  , \g73818/_0_  , \g73819/_0_  , \g73820/_0_  , \g73821/_0_  , \g73822/_0_  , \g73823/_0_  , \g73824/_0_  , \g73825/_0_  , \g73826/_0_  , \g73827/_0_  , \g73828/_0_  , \g73829/_0_  , \g73830/_0_  , \g73831/_0_  , \g73832/_0_  , \g73833/_0_  , \g73834/_0_  , \g73835/_0_  , \g73836/_0_  , \g73908/_0_  , \g73909/_0_  , \g73911/_0_  , \g73912/_0_  , \g73915/_0_  , \g73916/_0_  , \g73946/_0_  , \g73950/_0_  , \g73957/_0_  , \g73958/_0_  , \g73959/_0_  , \g73960/_0_  , \g73961/_0_  , \g73962/_0_  , \g73963/_0_  , \g73964/_0_  , \g73965/_0_  , \g73966/_0_  , \g73968/_0_  , \g73969/_0_  , \g73970/_0_  , \g73971/_0_  , \g73972/_0_  , \g73973/_0_  , \g73974/_0_  , \g73975/_0_  , \g73976/_0_  , \g73977/_0_  , \g73978/_0_  , \g73979/_0_  , \g73980/_0_  , \g73981/_0_  , \g73982/_0_  , \g73983/_0_  , \g73984/_0_  , \g73985/_0_  , \g74044/_0_  , \g74045/_0_  , \g74046/_0_  , \g74047/_0_  , \g74048/_0_  , \g74049/_0_  , \g74051/_0_  , \g74052/_0_  , \g74099/_0_  , \g74100/_0_  , \g74101/_0_  , \g74102/_0_  , \g74103/_0_  , \g74104/_0_  , \g74105/_0_  , \g74106/_0_  , \g74107/_0_  , \g74108/_0_  , \g74109/_0_  , \g74110/_0_  , \g74111/_0_  , \g74112/_0_  , \g74113/_0_  , \g74114/_0_  , \g74115/_0_  , \g74116/_0_  , \g74117/_0_  , \g74118/_0_  , \g74119/_0_  , \g74120/_0_  , \g74121/_0_  , \g74122/_0_  , \g74199/_0_  , \g74200/_0_  , \g74201/_0_  , \g74202/_0_  , \g74279/_0_  , \g74280/_0_  , \g74284/_0_  , \g74285/_0_  , \g74287/_0_  , \g74288/_0_  , \g74289/_0_  , \g74290/_0_  , \g74291/_0_  , \g74292/_0_  , \g74293/_0_  , \g74294/_0_  , \g74295/_0_  , \g74296/_0_  , \g74298/_0_  , \g74299/_0_  , \g74300/_0_  , \g74301/_0_  , \g74302/_0_  , \g74382/_0_  , \g74383/_0_  , \g74384/_0_  , \g74385/_0_  , \g74386/_0_  , \g74387/_0_  , \g74456/_0_  , \g74457/_0_  , \g74458/_0_  , \g74459/_0_  , \g74460/_0_  , \g74461/_0_  , \g74462/_0_  , \g74463/_0_  , \g74464/_0_  , \g74465/_0_  , \g74466/_0_  , \g74467/_0_  , \g74468/_0_  , \g74469/_0_  , \g74470/_0_  , \g74471/_0_  , \g74661/_0_  , \g74662/_0_  , \g74663/_0_  , \g74664/_0_  , \g74665/_0_  , \g74666/_0_  , \g74667/_0_  , \g74668/_0_  , \g74669/_0_  , \g74670/_0_  , \g74671/_0_  , \g74672/_0_  , \g74673/_0_  , \g74674/_0_  , \g74899/_0_  , \g74900/_0_  , \g74901/_0_  , \g74902/_0_  , \g75002/_0_  , \g75005/_0_  , \g75191/_0_  , \g75192/_0_  , \g75193/_0_  , \g75194/_0_  , \g75195/_0_  , \g75392/_0_  , \g75399/_0_  , \g75606/_0_  , \g75607/_0_  , \g75608/_0_  , \g75609/_0_  , \g75610/_0_  , \g76007/_0_  , \g76008/_0_  , \g76685/_0_  , \g76696/_0_  , \g77574/_0_  , \g77575/_0_  , \g77576/_0_  , \g77577/_0_  , \g77578/_0_  , \g77579/_0_  , \g82699/_3_  , \g82700/_3_  , \g82701/_3_  , \g82702/_3_  , \g82703/_3_  , \g82704/_3_  , \g83319/_0_  , \g83320/_0_  , \g83321/_0_  , \g83322/_0_  , \g83323/_3_  , \g83324/_0_  , \g83325/_0_  , \g83326/_0_  , \g83327/_0_  , \g83328/_0_  , \g83329/_0_  , \g83330/_0_  , \g83331/_0_  , \g83332/_0_  , \g83333/_0_  , \g83334/_0_  , \g83335/_0_  , \g83336/_3_  , \g83337/_0_  , \g83338/_0_  , \g83339/_0_  , \g83340/_0_  , \g83341/_0_  , \g83342/_0_  , \g83343/_0_  , \g83344/_0_  , \g83345/_0_  , \g83347/_3_  , \g83348/_3_  , \g83349/_3_  , \g83350/_3_  , \g83351/_3_  , \g83352/_3_  , \g83353/_3_  , \g83354/_3_  , \g83355/_3_  , \g83356/_3_  , \g83357/_0_  , \g83358/_3_  , \g83359/_3_  , \g83360/_3_  , \g83361/_3_  , \g83362/_3_  , \g83363/_3_  , \g83364/_3_  , \g83365/_0_  , \g83366/_3_  , \g83367/_0_  , \g83368/_3_  , \g83369/_3_  , \g83370/_0_  , \g83371/_3_  , \g83372/_3_  , \g83373/_3_  , \g83374/_3_  , \g83376/_0_  , \g83778/_0_  , \g83784/_0_  , \g84388/_0_  , \g84389/_0_  , \g84391/_0_  , \g84395/_0_  , \g84397/_0_  , \g84398/_0_  , \g84399/_0_  , \g84400/_0_  , \g84401/_0_  , \g84402/_0_  , \g84403/_0_  , \g84405/_0_  , \g84406/_0_  , \g84407/_0_  , \g84408/_0_  , \g84409/_0_  , \g84410/_0_  , \g84411/_0_  , \g84412/_0_  , \g84413/_0_  , \g84414/_0_  , \g84415/_0_  , \g84416/_0_  , \g84417/_0_  , \g84418/_0_  , \g84419/_0_  , \g84420/_0_  , \g84421/_0_  , \g84422/_0_  , \g84423/_0_  , \g84424/_0_  , \g84425/_0_  , \g84426/_0_  , \g84427/_0_  , \g84429/_0_  , \g84430/_0_  , \g84442/_0_  , \g84443/_0_  , \g84444/_0_  , \g84445/_0_  , \g84908/_0_  , \g84961/_0_  , \g84984/u3_syn_4  , \g84985/u3_syn_4  , \g85802/_0_  , \g86055/_1_  , \g86073/_0_  , \g86298/u3_syn_4  , \g86300/u3_syn_4  , \g87397/_0_  , \g87409/_0_  , \g87480/_0_  , \g87494/_0_  , \g87544/_0_  , \g87555/_0_  , \g87567/_0_  , \g87576/_0_  , \g87894/_0_  , \g87905/_0_  , \g87914/_0_  , \g87955/_1_  , \g88030/_0_  , \g88039/_0_  , \g88054/_0_  , \g88079/_0_  , \g88094/_0_  , \g88111/_0_  , \g88122/_0_  , \g88129/_0_  , \g88162/_0_  , \g88185/_0_  , \g88196/_0_  , \g88204/_0_  , \g88220/_0_  , \g88226/_0_  , \g88243/_0_  , \g88252/_0_  , \g88261/_0_  , \g88269/_0_  , \g88288/_0_  , \g88299/_0_  , \g88310/_0_  , \g88321/_0_  , \g88328/_0_  , \g88335/_0_  , \g88356/_0_  , \g88366/_0_  , \g88372/_0_  , \g88380/_0_  , \g88395_dup/_0_  , \g88403/_0_  , \g88414/_0_  , \g88425/_0_  , \g88443/_0_  , \g88453/_0_  , \g88471/_0_  , \g88524/_0_  , \g88546/_0_  , \g88556/_0_  , \g88563/_0_  , \g89966/_1_  , \g89999/_1_  , \g95209/_0_  , \g95269/_0_  , \g95319/_0_  , \g95354/_0_  , \g95786/_0_  , \g95909/_0_  , \g95914/_0_  , \g95918/_0_  , \g95984/_0_  , \g96009/_0_  , \g96124/_0_  , \g96218/_0_  , \g96286/_0_  , \g96335/_0_  , \g96465/_0_  , \g96694/_0_  , \g96713/_0_  , \g96830/_0_  , \g96875/_0_  , rd_pad , \so[0]_pad  , \so[10]_pad  , \so[11]_pad  , \so[12]_pad  , \so[13]_pad  , \so[14]_pad  , \so[15]_pad  , \so[16]_pad  , \so[17]_pad  , \so[18]_pad  , \so[19]_pad  , \so[1]_pad  , \so[2]_pad  , \so[3]_pad  , \so[4]_pad  , \so[5]_pad  , \so[6]_pad  , \so[7]_pad  , \so[8]_pad  , \so[9]_pad  , wr_pad );
  input \P1_B_reg/NET0131  ;
  input \P1_IR_reg[0]/NET0131  ;
  input \P1_IR_reg[10]/NET0131  ;
  input \P1_IR_reg[11]/NET0131  ;
  input \P1_IR_reg[12]/NET0131  ;
  input \P1_IR_reg[13]/NET0131  ;
  input \P1_IR_reg[14]/NET0131  ;
  input \P1_IR_reg[15]/NET0131  ;
  input \P1_IR_reg[16]/NET0131  ;
  input \P1_IR_reg[17]/NET0131  ;
  input \P1_IR_reg[18]/NET0131  ;
  input \P1_IR_reg[19]/NET0131  ;
  input \P1_IR_reg[1]/NET0131  ;
  input \P1_IR_reg[20]/NET0131  ;
  input \P1_IR_reg[21]/NET0131  ;
  input \P1_IR_reg[22]/NET0131  ;
  input \P1_IR_reg[23]/NET0131  ;
  input \P1_IR_reg[24]/NET0131  ;
  input \P1_IR_reg[25]/NET0131  ;
  input \P1_IR_reg[26]/NET0131  ;
  input \P1_IR_reg[27]/NET0131  ;
  input \P1_IR_reg[28]/NET0131  ;
  input \P1_IR_reg[29]/NET0131  ;
  input \P1_IR_reg[2]/NET0131  ;
  input \P1_IR_reg[30]/NET0131  ;
  input \P1_IR_reg[31]/NET0131  ;
  input \P1_IR_reg[3]/NET0131  ;
  input \P1_IR_reg[4]/NET0131  ;
  input \P1_IR_reg[5]/NET0131  ;
  input \P1_IR_reg[6]/NET0131  ;
  input \P1_IR_reg[7]/NET0131  ;
  input \P1_IR_reg[8]/NET0131  ;
  input \P1_IR_reg[9]/NET0131  ;
  input \P1_addr_reg[0]/NET0131  ;
  input \P1_addr_reg[10]/NET0131  ;
  input \P1_addr_reg[11]/NET0131  ;
  input \P1_addr_reg[12]/NET0131  ;
  input \P1_addr_reg[13]/NET0131  ;
  input \P1_addr_reg[14]/NET0131  ;
  input \P1_addr_reg[15]/NET0131  ;
  input \P1_addr_reg[16]/NET0131  ;
  input \P1_addr_reg[17]/NET0131  ;
  input \P1_addr_reg[18]/NET0131  ;
  input \P1_addr_reg[19]/NET0131  ;
  input \P1_addr_reg[1]/NET0131  ;
  input \P1_addr_reg[2]/NET0131  ;
  input \P1_addr_reg[3]/NET0131  ;
  input \P1_addr_reg[4]/NET0131  ;
  input \P1_addr_reg[5]/NET0131  ;
  input \P1_addr_reg[6]/NET0131  ;
  input \P1_addr_reg[7]/NET0131  ;
  input \P1_addr_reg[8]/NET0131  ;
  input \P1_addr_reg[9]/NET0131  ;
  input \P1_d_reg[0]/NET0131  ;
  input \P1_d_reg[1]/NET0131  ;
  input \P1_datao_reg[0]/NET0131  ;
  input \P1_datao_reg[10]/NET0131  ;
  input \P1_datao_reg[11]/NET0131  ;
  input \P1_datao_reg[12]/NET0131  ;
  input \P1_datao_reg[13]/NET0131  ;
  input \P1_datao_reg[14]/NET0131  ;
  input \P1_datao_reg[15]/NET0131  ;
  input \P1_datao_reg[16]/NET0131  ;
  input \P1_datao_reg[17]/NET0131  ;
  input \P1_datao_reg[18]/NET0131  ;
  input \P1_datao_reg[19]/NET0131  ;
  input \P1_datao_reg[1]/NET0131  ;
  input \P1_datao_reg[20]/NET0131  ;
  input \P1_datao_reg[21]/NET0131  ;
  input \P1_datao_reg[22]/NET0131  ;
  input \P1_datao_reg[23]/NET0131  ;
  input \P1_datao_reg[24]/NET0131  ;
  input \P1_datao_reg[25]/NET0131  ;
  input \P1_datao_reg[26]/NET0131  ;
  input \P1_datao_reg[27]/NET0131  ;
  input \P1_datao_reg[28]/NET0131  ;
  input \P1_datao_reg[29]/NET0131  ;
  input \P1_datao_reg[2]/NET0131  ;
  input \P1_datao_reg[30]/NET0131  ;
  input \P1_datao_reg[31]/NET0131  ;
  input \P1_datao_reg[3]/NET0131  ;
  input \P1_datao_reg[4]/NET0131  ;
  input \P1_datao_reg[5]/NET0131  ;
  input \P1_datao_reg[6]/NET0131  ;
  input \P1_datao_reg[7]/NET0131  ;
  input \P1_datao_reg[8]/NET0131  ;
  input \P1_datao_reg[9]/NET0131  ;
  input \P1_rd_reg/NET0131  ;
  input \P1_reg0_reg[0]/NET0131  ;
  input \P1_reg0_reg[10]/NET0131  ;
  input \P1_reg0_reg[11]/NET0131  ;
  input \P1_reg0_reg[12]/NET0131  ;
  input \P1_reg0_reg[13]/NET0131  ;
  input \P1_reg0_reg[14]/NET0131  ;
  input \P1_reg0_reg[15]/NET0131  ;
  input \P1_reg0_reg[16]/NET0131  ;
  input \P1_reg0_reg[17]/NET0131  ;
  input \P1_reg0_reg[18]/NET0131  ;
  input \P1_reg0_reg[19]/NET0131  ;
  input \P1_reg0_reg[1]/NET0131  ;
  input \P1_reg0_reg[20]/NET0131  ;
  input \P1_reg0_reg[21]/NET0131  ;
  input \P1_reg0_reg[22]/NET0131  ;
  input \P1_reg0_reg[23]/NET0131  ;
  input \P1_reg0_reg[24]/NET0131  ;
  input \P1_reg0_reg[25]/NET0131  ;
  input \P1_reg0_reg[26]/NET0131  ;
  input \P1_reg0_reg[27]/NET0131  ;
  input \P1_reg0_reg[28]/NET0131  ;
  input \P1_reg0_reg[29]/NET0131  ;
  input \P1_reg0_reg[2]/NET0131  ;
  input \P1_reg0_reg[30]/NET0131  ;
  input \P1_reg0_reg[31]/NET0131  ;
  input \P1_reg0_reg[3]/NET0131  ;
  input \P1_reg0_reg[4]/NET0131  ;
  input \P1_reg0_reg[5]/NET0131  ;
  input \P1_reg0_reg[6]/NET0131  ;
  input \P1_reg0_reg[7]/NET0131  ;
  input \P1_reg0_reg[8]/NET0131  ;
  input \P1_reg0_reg[9]/NET0131  ;
  input \P1_reg1_reg[0]/NET0131  ;
  input \P1_reg1_reg[10]/NET0131  ;
  input \P1_reg1_reg[11]/NET0131  ;
  input \P1_reg1_reg[12]/NET0131  ;
  input \P1_reg1_reg[13]/NET0131  ;
  input \P1_reg1_reg[14]/NET0131  ;
  input \P1_reg1_reg[15]/NET0131  ;
  input \P1_reg1_reg[16]/NET0131  ;
  input \P1_reg1_reg[17]/NET0131  ;
  input \P1_reg1_reg[18]/NET0131  ;
  input \P1_reg1_reg[19]/NET0131  ;
  input \P1_reg1_reg[1]/NET0131  ;
  input \P1_reg1_reg[20]/NET0131  ;
  input \P1_reg1_reg[21]/NET0131  ;
  input \P1_reg1_reg[22]/NET0131  ;
  input \P1_reg1_reg[23]/NET0131  ;
  input \P1_reg1_reg[24]/NET0131  ;
  input \P1_reg1_reg[25]/NET0131  ;
  input \P1_reg1_reg[26]/NET0131  ;
  input \P1_reg1_reg[27]/NET0131  ;
  input \P1_reg1_reg[28]/NET0131  ;
  input \P1_reg1_reg[29]/NET0131  ;
  input \P1_reg1_reg[2]/NET0131  ;
  input \P1_reg1_reg[30]/NET0131  ;
  input \P1_reg1_reg[31]/NET0131  ;
  input \P1_reg1_reg[3]/NET0131  ;
  input \P1_reg1_reg[4]/NET0131  ;
  input \P1_reg1_reg[5]/NET0131  ;
  input \P1_reg1_reg[6]/NET0131  ;
  input \P1_reg1_reg[7]/NET0131  ;
  input \P1_reg1_reg[8]/NET0131  ;
  input \P1_reg1_reg[9]/NET0131  ;
  input \P1_reg2_reg[0]/NET0131  ;
  input \P1_reg2_reg[10]/NET0131  ;
  input \P1_reg2_reg[11]/NET0131  ;
  input \P1_reg2_reg[12]/NET0131  ;
  input \P1_reg2_reg[13]/NET0131  ;
  input \P1_reg2_reg[14]/NET0131  ;
  input \P1_reg2_reg[15]/NET0131  ;
  input \P1_reg2_reg[16]/NET0131  ;
  input \P1_reg2_reg[17]/NET0131  ;
  input \P1_reg2_reg[18]/NET0131  ;
  input \P1_reg2_reg[19]/NET0131  ;
  input \P1_reg2_reg[1]/NET0131  ;
  input \P1_reg2_reg[20]/NET0131  ;
  input \P1_reg2_reg[21]/NET0131  ;
  input \P1_reg2_reg[22]/NET0131  ;
  input \P1_reg2_reg[23]/NET0131  ;
  input \P1_reg2_reg[24]/NET0131  ;
  input \P1_reg2_reg[25]/NET0131  ;
  input \P1_reg2_reg[26]/NET0131  ;
  input \P1_reg2_reg[27]/NET0131  ;
  input \P1_reg2_reg[28]/NET0131  ;
  input \P1_reg2_reg[29]/NET0131  ;
  input \P1_reg2_reg[2]/NET0131  ;
  input \P1_reg2_reg[30]/NET0131  ;
  input \P1_reg2_reg[31]/NET0131  ;
  input \P1_reg2_reg[3]/NET0131  ;
  input \P1_reg2_reg[4]/NET0131  ;
  input \P1_reg2_reg[5]/NET0131  ;
  input \P1_reg2_reg[6]/NET0131  ;
  input \P1_reg2_reg[7]/NET0131  ;
  input \P1_reg2_reg[8]/NET0131  ;
  input \P1_reg2_reg[9]/NET0131  ;
  input \P1_reg3_reg[0]/NET0131  ;
  input \P1_reg3_reg[10]/NET0131  ;
  input \P1_reg3_reg[11]/NET0131  ;
  input \P1_reg3_reg[12]/NET0131  ;
  input \P1_reg3_reg[13]/NET0131  ;
  input \P1_reg3_reg[14]/NET0131  ;
  input \P1_reg3_reg[15]/NET0131  ;
  input \P1_reg3_reg[16]/NET0131  ;
  input \P1_reg3_reg[17]/NET0131  ;
  input \P1_reg3_reg[18]/NET0131  ;
  input \P1_reg3_reg[19]/NET0131  ;
  input \P1_reg3_reg[1]/NET0131  ;
  input \P1_reg3_reg[20]/NET0131  ;
  input \P1_reg3_reg[21]/NET0131  ;
  input \P1_reg3_reg[22]/NET0131  ;
  input \P1_reg3_reg[23]/NET0131  ;
  input \P1_reg3_reg[24]/NET0131  ;
  input \P1_reg3_reg[25]/NET0131  ;
  input \P1_reg3_reg[26]/NET0131  ;
  input \P1_reg3_reg[27]/NET0131  ;
  input \P1_reg3_reg[28]/NET0131  ;
  input \P1_reg3_reg[2]/NET0131  ;
  input \P1_reg3_reg[3]/NET0131  ;
  input \P1_reg3_reg[4]/NET0131  ;
  input \P1_reg3_reg[5]/NET0131  ;
  input \P1_reg3_reg[6]/NET0131  ;
  input \P1_reg3_reg[7]/NET0131  ;
  input \P1_reg3_reg[8]/NET0131  ;
  input \P1_reg3_reg[9]/NET0131  ;
  input \P1_state_reg[0]/NET0131  ;
  input \P1_wr_reg/NET0131  ;
  input \P2_B_reg/NET0131  ;
  input \P2_IR_reg[0]/NET0131  ;
  input \P2_IR_reg[10]/NET0131  ;
  input \P2_IR_reg[11]/NET0131  ;
  input \P2_IR_reg[12]/NET0131  ;
  input \P2_IR_reg[13]/NET0131  ;
  input \P2_IR_reg[14]/NET0131  ;
  input \P2_IR_reg[15]/NET0131  ;
  input \P2_IR_reg[16]/NET0131  ;
  input \P2_IR_reg[17]/NET0131  ;
  input \P2_IR_reg[18]/NET0131  ;
  input \P2_IR_reg[19]/NET0131  ;
  input \P2_IR_reg[1]/NET0131  ;
  input \P2_IR_reg[20]/NET0131  ;
  input \P2_IR_reg[21]/NET0131  ;
  input \P2_IR_reg[22]/NET0131  ;
  input \P2_IR_reg[23]/NET0131  ;
  input \P2_IR_reg[24]/NET0131  ;
  input \P2_IR_reg[25]/NET0131  ;
  input \P2_IR_reg[26]/NET0131  ;
  input \P2_IR_reg[27]/NET0131  ;
  input \P2_IR_reg[28]/NET0131  ;
  input \P2_IR_reg[29]/NET0131  ;
  input \P2_IR_reg[2]/NET0131  ;
  input \P2_IR_reg[30]/NET0131  ;
  input \P2_IR_reg[31]/NET0131  ;
  input \P2_IR_reg[3]/NET0131  ;
  input \P2_IR_reg[4]/NET0131  ;
  input \P2_IR_reg[5]/NET0131  ;
  input \P2_IR_reg[6]/NET0131  ;
  input \P2_IR_reg[7]/NET0131  ;
  input \P2_IR_reg[8]/NET0131  ;
  input \P2_IR_reg[9]/NET0131  ;
  input \P2_addr_reg[0]/NET0131  ;
  input \P2_addr_reg[10]/NET0131  ;
  input \P2_addr_reg[11]/NET0131  ;
  input \P2_addr_reg[12]/NET0131  ;
  input \P2_addr_reg[13]/NET0131  ;
  input \P2_addr_reg[14]/NET0131  ;
  input \P2_addr_reg[15]/NET0131  ;
  input \P2_addr_reg[16]/NET0131  ;
  input \P2_addr_reg[17]/NET0131  ;
  input \P2_addr_reg[18]/NET0131  ;
  input \P2_addr_reg[19]/NET0131  ;
  input \P2_addr_reg[1]/NET0131  ;
  input \P2_addr_reg[2]/NET0131  ;
  input \P2_addr_reg[3]/NET0131  ;
  input \P2_addr_reg[4]/NET0131  ;
  input \P2_addr_reg[5]/NET0131  ;
  input \P2_addr_reg[6]/NET0131  ;
  input \P2_addr_reg[7]/NET0131  ;
  input \P2_addr_reg[8]/NET0131  ;
  input \P2_addr_reg[9]/NET0131  ;
  input \P2_d_reg[0]/NET0131  ;
  input \P2_d_reg[1]/NET0131  ;
  input \P2_datao_reg[0]/NET0131  ;
  input \P2_datao_reg[10]/NET0131  ;
  input \P2_datao_reg[11]/NET0131  ;
  input \P2_datao_reg[12]/NET0131  ;
  input \P2_datao_reg[13]/NET0131  ;
  input \P2_datao_reg[14]/NET0131  ;
  input \P2_datao_reg[15]/NET0131  ;
  input \P2_datao_reg[16]/NET0131  ;
  input \P2_datao_reg[17]/NET0131  ;
  input \P2_datao_reg[18]/NET0131  ;
  input \P2_datao_reg[19]/NET0131  ;
  input \P2_datao_reg[1]/NET0131  ;
  input \P2_datao_reg[20]/NET0131  ;
  input \P2_datao_reg[21]/NET0131  ;
  input \P2_datao_reg[22]/NET0131  ;
  input \P2_datao_reg[23]/NET0131  ;
  input \P2_datao_reg[24]/NET0131  ;
  input \P2_datao_reg[25]/NET0131  ;
  input \P2_datao_reg[26]/NET0131  ;
  input \P2_datao_reg[27]/NET0131  ;
  input \P2_datao_reg[28]/NET0131  ;
  input \P2_datao_reg[29]/NET0131  ;
  input \P2_datao_reg[2]/NET0131  ;
  input \P2_datao_reg[30]/NET0131  ;
  input \P2_datao_reg[31]/NET0131  ;
  input \P2_datao_reg[3]/NET0131  ;
  input \P2_datao_reg[4]/NET0131  ;
  input \P2_datao_reg[5]/NET0131  ;
  input \P2_datao_reg[6]/NET0131  ;
  input \P2_datao_reg[7]/NET0131  ;
  input \P2_datao_reg[8]/NET0131  ;
  input \P2_datao_reg[9]/NET0131  ;
  input \P2_rd_reg/NET0131  ;
  input \P2_reg0_reg[0]/NET0131  ;
  input \P2_reg0_reg[10]/NET0131  ;
  input \P2_reg0_reg[11]/NET0131  ;
  input \P2_reg0_reg[12]/NET0131  ;
  input \P2_reg0_reg[13]/NET0131  ;
  input \P2_reg0_reg[14]/NET0131  ;
  input \P2_reg0_reg[15]/NET0131  ;
  input \P2_reg0_reg[16]/NET0131  ;
  input \P2_reg0_reg[17]/NET0131  ;
  input \P2_reg0_reg[18]/NET0131  ;
  input \P2_reg0_reg[19]/NET0131  ;
  input \P2_reg0_reg[1]/NET0131  ;
  input \P2_reg0_reg[20]/NET0131  ;
  input \P2_reg0_reg[21]/NET0131  ;
  input \P2_reg0_reg[22]/NET0131  ;
  input \P2_reg0_reg[23]/NET0131  ;
  input \P2_reg0_reg[24]/NET0131  ;
  input \P2_reg0_reg[25]/NET0131  ;
  input \P2_reg0_reg[26]/NET0131  ;
  input \P2_reg0_reg[27]/NET0131  ;
  input \P2_reg0_reg[28]/NET0131  ;
  input \P2_reg0_reg[29]/NET0131  ;
  input \P2_reg0_reg[2]/NET0131  ;
  input \P2_reg0_reg[30]/NET0131  ;
  input \P2_reg0_reg[31]/NET0131  ;
  input \P2_reg0_reg[3]/NET0131  ;
  input \P2_reg0_reg[4]/NET0131  ;
  input \P2_reg0_reg[5]/NET0131  ;
  input \P2_reg0_reg[6]/NET0131  ;
  input \P2_reg0_reg[7]/NET0131  ;
  input \P2_reg0_reg[8]/NET0131  ;
  input \P2_reg0_reg[9]/NET0131  ;
  input \P2_reg1_reg[0]/NET0131  ;
  input \P2_reg1_reg[10]/NET0131  ;
  input \P2_reg1_reg[11]/NET0131  ;
  input \P2_reg1_reg[12]/NET0131  ;
  input \P2_reg1_reg[13]/NET0131  ;
  input \P2_reg1_reg[14]/NET0131  ;
  input \P2_reg1_reg[15]/NET0131  ;
  input \P2_reg1_reg[16]/NET0131  ;
  input \P2_reg1_reg[17]/NET0131  ;
  input \P2_reg1_reg[18]/NET0131  ;
  input \P2_reg1_reg[19]/NET0131  ;
  input \P2_reg1_reg[1]/NET0131  ;
  input \P2_reg1_reg[20]/NET0131  ;
  input \P2_reg1_reg[21]/NET0131  ;
  input \P2_reg1_reg[22]/NET0131  ;
  input \P2_reg1_reg[23]/NET0131  ;
  input \P2_reg1_reg[24]/NET0131  ;
  input \P2_reg1_reg[25]/NET0131  ;
  input \P2_reg1_reg[26]/NET0131  ;
  input \P2_reg1_reg[27]/NET0131  ;
  input \P2_reg1_reg[28]/NET0131  ;
  input \P2_reg1_reg[29]/NET0131  ;
  input \P2_reg1_reg[2]/NET0131  ;
  input \P2_reg1_reg[30]/NET0131  ;
  input \P2_reg1_reg[31]/NET0131  ;
  input \P2_reg1_reg[3]/NET0131  ;
  input \P2_reg1_reg[4]/NET0131  ;
  input \P2_reg1_reg[5]/NET0131  ;
  input \P2_reg1_reg[6]/NET0131  ;
  input \P2_reg1_reg[7]/NET0131  ;
  input \P2_reg1_reg[8]/NET0131  ;
  input \P2_reg1_reg[9]/NET0131  ;
  input \P2_reg2_reg[0]/NET0131  ;
  input \P2_reg2_reg[10]/NET0131  ;
  input \P2_reg2_reg[11]/NET0131  ;
  input \P2_reg2_reg[12]/NET0131  ;
  input \P2_reg2_reg[13]/NET0131  ;
  input \P2_reg2_reg[14]/NET0131  ;
  input \P2_reg2_reg[15]/NET0131  ;
  input \P2_reg2_reg[16]/NET0131  ;
  input \P2_reg2_reg[17]/NET0131  ;
  input \P2_reg2_reg[18]/NET0131  ;
  input \P2_reg2_reg[19]/NET0131  ;
  input \P2_reg2_reg[1]/NET0131  ;
  input \P2_reg2_reg[20]/NET0131  ;
  input \P2_reg2_reg[21]/NET0131  ;
  input \P2_reg2_reg[22]/NET0131  ;
  input \P2_reg2_reg[23]/NET0131  ;
  input \P2_reg2_reg[24]/NET0131  ;
  input \P2_reg2_reg[25]/NET0131  ;
  input \P2_reg2_reg[26]/NET0131  ;
  input \P2_reg2_reg[27]/NET0131  ;
  input \P2_reg2_reg[28]/NET0131  ;
  input \P2_reg2_reg[29]/NET0131  ;
  input \P2_reg2_reg[2]/NET0131  ;
  input \P2_reg2_reg[30]/NET0131  ;
  input \P2_reg2_reg[31]/NET0131  ;
  input \P2_reg2_reg[3]/NET0131  ;
  input \P2_reg2_reg[4]/NET0131  ;
  input \P2_reg2_reg[5]/NET0131  ;
  input \P2_reg2_reg[6]/NET0131  ;
  input \P2_reg2_reg[7]/NET0131  ;
  input \P2_reg2_reg[8]/NET0131  ;
  input \P2_reg2_reg[9]/NET0131  ;
  input \P2_reg3_reg[0]/NET0131  ;
  input \P2_reg3_reg[10]/NET0131  ;
  input \P2_reg3_reg[11]/NET0131  ;
  input \P2_reg3_reg[12]/NET0131  ;
  input \P2_reg3_reg[13]/NET0131  ;
  input \P2_reg3_reg[14]/NET0131  ;
  input \P2_reg3_reg[15]/NET0131  ;
  input \P2_reg3_reg[16]/NET0131  ;
  input \P2_reg3_reg[17]/NET0131  ;
  input \P2_reg3_reg[18]/NET0131  ;
  input \P2_reg3_reg[19]/NET0131  ;
  input \P2_reg3_reg[1]/NET0131  ;
  input \P2_reg3_reg[20]/NET0131  ;
  input \P2_reg3_reg[21]/NET0131  ;
  input \P2_reg3_reg[22]/NET0131  ;
  input \P2_reg3_reg[23]/NET0131  ;
  input \P2_reg3_reg[24]/NET0131  ;
  input \P2_reg3_reg[25]/NET0131  ;
  input \P2_reg3_reg[26]/NET0131  ;
  input \P2_reg3_reg[27]/NET0131  ;
  input \P2_reg3_reg[28]/NET0131  ;
  input \P2_reg3_reg[2]/NET0131  ;
  input \P2_reg3_reg[3]/NET0131  ;
  input \P2_reg3_reg[4]/NET0131  ;
  input \P2_reg3_reg[5]/NET0131  ;
  input \P2_reg3_reg[6]/NET0131  ;
  input \P2_reg3_reg[7]/NET0131  ;
  input \P2_reg3_reg[8]/NET0131  ;
  input \P2_reg3_reg[9]/NET0131  ;
  input \P2_wr_reg/NET0131  ;
  input \si[0]_pad  ;
  input \si[10]_pad  ;
  input \si[11]_pad  ;
  input \si[12]_pad  ;
  input \si[13]_pad  ;
  input \si[14]_pad  ;
  input \si[15]_pad  ;
  input \si[16]_pad  ;
  input \si[17]_pad  ;
  input \si[18]_pad  ;
  input \si[19]_pad  ;
  input \si[1]_pad  ;
  input \si[20]_pad  ;
  input \si[21]_pad  ;
  input \si[22]_pad  ;
  input \si[23]_pad  ;
  input \si[24]_pad  ;
  input \si[25]_pad  ;
  input \si[26]_pad  ;
  input \si[27]_pad  ;
  input \si[28]_pad  ;
  input \si[29]_pad  ;
  input \si[2]_pad  ;
  input \si[30]_pad  ;
  input \si[31]_pad  ;
  input \si[3]_pad  ;
  input \si[4]_pad  ;
  input \si[5]_pad  ;
  input \si[6]_pad  ;
  input \si[7]_pad  ;
  input \si[8]_pad  ;
  input \si[9]_pad  ;
  output \P1_state_reg[0]/NET0131_syn_2  ;
  output \_al_n0  ;
  output \_al_n1  ;
  output \g73521/_0_  ;
  output \g73537/_0_  ;
  output \g73538/_0_  ;
  output \g73539/_0_  ;
  output \g73540/_0_  ;
  output \g73570/_0_  ;
  output \g73571/_0_  ;
  output \g73572/_0_  ;
  output \g73573/_0_  ;
  output \g73574/_0_  ;
  output \g73575/_0_  ;
  output \g73576/_0_  ;
  output \g73577/_0_  ;
  output \g73578/_0_  ;
  output \g73579/_0_  ;
  output \g73609/_0_  ;
  output \g73610/_0_  ;
  output \g73611/_0_  ;
  output \g73613/_0_  ;
  output \g73614/_0_  ;
  output \g73615/_0_  ;
  output \g73617/_0_  ;
  output \g73618/_0_  ;
  output \g73619/_0_  ;
  output \g73620/_0_  ;
  output \g73621/_0_  ;
  output \g73622/_0_  ;
  output \g73623/_0_  ;
  output \g73624/_0_  ;
  output \g73625/_0_  ;
  output \g73626/_0_  ;
  output \g73627/_0_  ;
  output \g73628/_0_  ;
  output \g73629/_0_  ;
  output \g73630/_0_  ;
  output \g73631/_0_  ;
  output \g73632/_0_  ;
  output \g73633/_0_  ;
  output \g73692/_0_  ;
  output \g73693/_0_  ;
  output \g73694/_0_  ;
  output \g73696/_0_  ;
  output \g73697/_0_  ;
  output \g73703/_0_  ;
  output \g73704/_0_  ;
  output \g73709/_0_  ;
  output \g73710/_0_  ;
  output \g73711/_0_  ;
  output \g73712/_0_  ;
  output \g73713/_0_  ;
  output \g73714/_0_  ;
  output \g73715/_0_  ;
  output \g73716/_0_  ;
  output \g73717/_0_  ;
  output \g73718/_0_  ;
  output \g73719/_0_  ;
  output \g73720/_0_  ;
  output \g73774/_0_  ;
  output \g73775/_0_  ;
  output \g73776/_0_  ;
  output \g73777/_0_  ;
  output \g73806/_0_  ;
  output \g73807/_0_  ;
  output \g73808/_0_  ;
  output \g73809/_0_  ;
  output \g73810/_0_  ;
  output \g73811/_0_  ;
  output \g73812/_0_  ;
  output \g73813/_0_  ;
  output \g73814/_0_  ;
  output \g73815/_0_  ;
  output \g73816/_0_  ;
  output \g73817/_0_  ;
  output \g73818/_0_  ;
  output \g73819/_0_  ;
  output \g73820/_0_  ;
  output \g73821/_0_  ;
  output \g73822/_0_  ;
  output \g73823/_0_  ;
  output \g73824/_0_  ;
  output \g73825/_0_  ;
  output \g73826/_0_  ;
  output \g73827/_0_  ;
  output \g73828/_0_  ;
  output \g73829/_0_  ;
  output \g73830/_0_  ;
  output \g73831/_0_  ;
  output \g73832/_0_  ;
  output \g73833/_0_  ;
  output \g73834/_0_  ;
  output \g73835/_0_  ;
  output \g73836/_0_  ;
  output \g73908/_0_  ;
  output \g73909/_0_  ;
  output \g73911/_0_  ;
  output \g73912/_0_  ;
  output \g73915/_0_  ;
  output \g73916/_0_  ;
  output \g73946/_0_  ;
  output \g73950/_0_  ;
  output \g73957/_0_  ;
  output \g73958/_0_  ;
  output \g73959/_0_  ;
  output \g73960/_0_  ;
  output \g73961/_0_  ;
  output \g73962/_0_  ;
  output \g73963/_0_  ;
  output \g73964/_0_  ;
  output \g73965/_0_  ;
  output \g73966/_0_  ;
  output \g73968/_0_  ;
  output \g73969/_0_  ;
  output \g73970/_0_  ;
  output \g73971/_0_  ;
  output \g73972/_0_  ;
  output \g73973/_0_  ;
  output \g73974/_0_  ;
  output \g73975/_0_  ;
  output \g73976/_0_  ;
  output \g73977/_0_  ;
  output \g73978/_0_  ;
  output \g73979/_0_  ;
  output \g73980/_0_  ;
  output \g73981/_0_  ;
  output \g73982/_0_  ;
  output \g73983/_0_  ;
  output \g73984/_0_  ;
  output \g73985/_0_  ;
  output \g74044/_0_  ;
  output \g74045/_0_  ;
  output \g74046/_0_  ;
  output \g74047/_0_  ;
  output \g74048/_0_  ;
  output \g74049/_0_  ;
  output \g74051/_0_  ;
  output \g74052/_0_  ;
  output \g74099/_0_  ;
  output \g74100/_0_  ;
  output \g74101/_0_  ;
  output \g74102/_0_  ;
  output \g74103/_0_  ;
  output \g74104/_0_  ;
  output \g74105/_0_  ;
  output \g74106/_0_  ;
  output \g74107/_0_  ;
  output \g74108/_0_  ;
  output \g74109/_0_  ;
  output \g74110/_0_  ;
  output \g74111/_0_  ;
  output \g74112/_0_  ;
  output \g74113/_0_  ;
  output \g74114/_0_  ;
  output \g74115/_0_  ;
  output \g74116/_0_  ;
  output \g74117/_0_  ;
  output \g74118/_0_  ;
  output \g74119/_0_  ;
  output \g74120/_0_  ;
  output \g74121/_0_  ;
  output \g74122/_0_  ;
  output \g74199/_0_  ;
  output \g74200/_0_  ;
  output \g74201/_0_  ;
  output \g74202/_0_  ;
  output \g74279/_0_  ;
  output \g74280/_0_  ;
  output \g74284/_0_  ;
  output \g74285/_0_  ;
  output \g74287/_0_  ;
  output \g74288/_0_  ;
  output \g74289/_0_  ;
  output \g74290/_0_  ;
  output \g74291/_0_  ;
  output \g74292/_0_  ;
  output \g74293/_0_  ;
  output \g74294/_0_  ;
  output \g74295/_0_  ;
  output \g74296/_0_  ;
  output \g74298/_0_  ;
  output \g74299/_0_  ;
  output \g74300/_0_  ;
  output \g74301/_0_  ;
  output \g74302/_0_  ;
  output \g74382/_0_  ;
  output \g74383/_0_  ;
  output \g74384/_0_  ;
  output \g74385/_0_  ;
  output \g74386/_0_  ;
  output \g74387/_0_  ;
  output \g74456/_0_  ;
  output \g74457/_0_  ;
  output \g74458/_0_  ;
  output \g74459/_0_  ;
  output \g74460/_0_  ;
  output \g74461/_0_  ;
  output \g74462/_0_  ;
  output \g74463/_0_  ;
  output \g74464/_0_  ;
  output \g74465/_0_  ;
  output \g74466/_0_  ;
  output \g74467/_0_  ;
  output \g74468/_0_  ;
  output \g74469/_0_  ;
  output \g74470/_0_  ;
  output \g74471/_0_  ;
  output \g74661/_0_  ;
  output \g74662/_0_  ;
  output \g74663/_0_  ;
  output \g74664/_0_  ;
  output \g74665/_0_  ;
  output \g74666/_0_  ;
  output \g74667/_0_  ;
  output \g74668/_0_  ;
  output \g74669/_0_  ;
  output \g74670/_0_  ;
  output \g74671/_0_  ;
  output \g74672/_0_  ;
  output \g74673/_0_  ;
  output \g74674/_0_  ;
  output \g74899/_0_  ;
  output \g74900/_0_  ;
  output \g74901/_0_  ;
  output \g74902/_0_  ;
  output \g75002/_0_  ;
  output \g75005/_0_  ;
  output \g75191/_0_  ;
  output \g75192/_0_  ;
  output \g75193/_0_  ;
  output \g75194/_0_  ;
  output \g75195/_0_  ;
  output \g75392/_0_  ;
  output \g75399/_0_  ;
  output \g75606/_0_  ;
  output \g75607/_0_  ;
  output \g75608/_0_  ;
  output \g75609/_0_  ;
  output \g75610/_0_  ;
  output \g76007/_0_  ;
  output \g76008/_0_  ;
  output \g76685/_0_  ;
  output \g76696/_0_  ;
  output \g77574/_0_  ;
  output \g77575/_0_  ;
  output \g77576/_0_  ;
  output \g77577/_0_  ;
  output \g77578/_0_  ;
  output \g77579/_0_  ;
  output \g82699/_3_  ;
  output \g82700/_3_  ;
  output \g82701/_3_  ;
  output \g82702/_3_  ;
  output \g82703/_3_  ;
  output \g82704/_3_  ;
  output \g83319/_0_  ;
  output \g83320/_0_  ;
  output \g83321/_0_  ;
  output \g83322/_0_  ;
  output \g83323/_3_  ;
  output \g83324/_0_  ;
  output \g83325/_0_  ;
  output \g83326/_0_  ;
  output \g83327/_0_  ;
  output \g83328/_0_  ;
  output \g83329/_0_  ;
  output \g83330/_0_  ;
  output \g83331/_0_  ;
  output \g83332/_0_  ;
  output \g83333/_0_  ;
  output \g83334/_0_  ;
  output \g83335/_0_  ;
  output \g83336/_3_  ;
  output \g83337/_0_  ;
  output \g83338/_0_  ;
  output \g83339/_0_  ;
  output \g83340/_0_  ;
  output \g83341/_0_  ;
  output \g83342/_0_  ;
  output \g83343/_0_  ;
  output \g83344/_0_  ;
  output \g83345/_0_  ;
  output \g83347/_3_  ;
  output \g83348/_3_  ;
  output \g83349/_3_  ;
  output \g83350/_3_  ;
  output \g83351/_3_  ;
  output \g83352/_3_  ;
  output \g83353/_3_  ;
  output \g83354/_3_  ;
  output \g83355/_3_  ;
  output \g83356/_3_  ;
  output \g83357/_0_  ;
  output \g83358/_3_  ;
  output \g83359/_3_  ;
  output \g83360/_3_  ;
  output \g83361/_3_  ;
  output \g83362/_3_  ;
  output \g83363/_3_  ;
  output \g83364/_3_  ;
  output \g83365/_0_  ;
  output \g83366/_3_  ;
  output \g83367/_0_  ;
  output \g83368/_3_  ;
  output \g83369/_3_  ;
  output \g83370/_0_  ;
  output \g83371/_3_  ;
  output \g83372/_3_  ;
  output \g83373/_3_  ;
  output \g83374/_3_  ;
  output \g83376/_0_  ;
  output \g83778/_0_  ;
  output \g83784/_0_  ;
  output \g84388/_0_  ;
  output \g84389/_0_  ;
  output \g84391/_0_  ;
  output \g84395/_0_  ;
  output \g84397/_0_  ;
  output \g84398/_0_  ;
  output \g84399/_0_  ;
  output \g84400/_0_  ;
  output \g84401/_0_  ;
  output \g84402/_0_  ;
  output \g84403/_0_  ;
  output \g84405/_0_  ;
  output \g84406/_0_  ;
  output \g84407/_0_  ;
  output \g84408/_0_  ;
  output \g84409/_0_  ;
  output \g84410/_0_  ;
  output \g84411/_0_  ;
  output \g84412/_0_  ;
  output \g84413/_0_  ;
  output \g84414/_0_  ;
  output \g84415/_0_  ;
  output \g84416/_0_  ;
  output \g84417/_0_  ;
  output \g84418/_0_  ;
  output \g84419/_0_  ;
  output \g84420/_0_  ;
  output \g84421/_0_  ;
  output \g84422/_0_  ;
  output \g84423/_0_  ;
  output \g84424/_0_  ;
  output \g84425/_0_  ;
  output \g84426/_0_  ;
  output \g84427/_0_  ;
  output \g84429/_0_  ;
  output \g84430/_0_  ;
  output \g84442/_0_  ;
  output \g84443/_0_  ;
  output \g84444/_0_  ;
  output \g84445/_0_  ;
  output \g84908/_0_  ;
  output \g84961/_0_  ;
  output \g84984/u3_syn_4  ;
  output \g84985/u3_syn_4  ;
  output \g85802/_0_  ;
  output \g86055/_1_  ;
  output \g86073/_0_  ;
  output \g86298/u3_syn_4  ;
  output \g86300/u3_syn_4  ;
  output \g87397/_0_  ;
  output \g87409/_0_  ;
  output \g87480/_0_  ;
  output \g87494/_0_  ;
  output \g87544/_0_  ;
  output \g87555/_0_  ;
  output \g87567/_0_  ;
  output \g87576/_0_  ;
  output \g87894/_0_  ;
  output \g87905/_0_  ;
  output \g87914/_0_  ;
  output \g87955/_1_  ;
  output \g88030/_0_  ;
  output \g88039/_0_  ;
  output \g88054/_0_  ;
  output \g88079/_0_  ;
  output \g88094/_0_  ;
  output \g88111/_0_  ;
  output \g88122/_0_  ;
  output \g88129/_0_  ;
  output \g88162/_0_  ;
  output \g88185/_0_  ;
  output \g88196/_0_  ;
  output \g88204/_0_  ;
  output \g88220/_0_  ;
  output \g88226/_0_  ;
  output \g88243/_0_  ;
  output \g88252/_0_  ;
  output \g88261/_0_  ;
  output \g88269/_0_  ;
  output \g88288/_0_  ;
  output \g88299/_0_  ;
  output \g88310/_0_  ;
  output \g88321/_0_  ;
  output \g88328/_0_  ;
  output \g88335/_0_  ;
  output \g88356/_0_  ;
  output \g88366/_0_  ;
  output \g88372/_0_  ;
  output \g88380/_0_  ;
  output \g88395_dup/_0_  ;
  output \g88403/_0_  ;
  output \g88414/_0_  ;
  output \g88425/_0_  ;
  output \g88443/_0_  ;
  output \g88453/_0_  ;
  output \g88471/_0_  ;
  output \g88524/_0_  ;
  output \g88546/_0_  ;
  output \g88556/_0_  ;
  output \g88563/_0_  ;
  output \g89966/_1_  ;
  output \g89999/_1_  ;
  output \g95209/_0_  ;
  output \g95269/_0_  ;
  output \g95319/_0_  ;
  output \g95354/_0_  ;
  output \g95786/_0_  ;
  output \g95909/_0_  ;
  output \g95914/_0_  ;
  output \g95918/_0_  ;
  output \g95984/_0_  ;
  output \g96009/_0_  ;
  output \g96124/_0_  ;
  output \g96218/_0_  ;
  output \g96286/_0_  ;
  output \g96335/_0_  ;
  output \g96465/_0_  ;
  output \g96694/_0_  ;
  output \g96713/_0_  ;
  output \g96830/_0_  ;
  output \g96875/_0_  ;
  output rd_pad ;
  output \so[0]_pad  ;
  output \so[10]_pad  ;
  output \so[11]_pad  ;
  output \so[12]_pad  ;
  output \so[13]_pad  ;
  output \so[14]_pad  ;
  output \so[15]_pad  ;
  output \so[16]_pad  ;
  output \so[17]_pad  ;
  output \so[18]_pad  ;
  output \so[19]_pad  ;
  output \so[1]_pad  ;
  output \so[2]_pad  ;
  output \so[3]_pad  ;
  output \so[4]_pad  ;
  output \so[5]_pad  ;
  output \so[6]_pad  ;
  output \so[7]_pad  ;
  output \so[8]_pad  ;
  output \so[9]_pad  ;
  output wr_pad ;
  wire n462 , n463 , n464 , n465 , n466 , n467 , n468 , n469 , n470 , n471 , n472 , n473 , n474 , n475 , n476 , n477 , n478 , n479 , n480 , n481 , n482 , n483 , n484 , n485 , n486 , n487 , n488 , n489 , n490 , n491 , n492 , n493 , n494 , n495 , n496 , n497 , n498 , n499 , n500 , n501 , n502 , n503 , n504 , n505 , n506 , n507 , n508 , n509 , n510 , n511 , n512 , n513 , n514 , n515 , n516 , n517 , n518 , n519 , n520 , n521 , n522 , n523 , n524 , n525 , n526 , n527 , n528 , n529 , n530 , n531 , n532 , n533 , n534 , n535 , n536 , n537 , n538 , n539 , n540 , n541 , n542 , n543 , n544 , n545 , n546 , n547 , n548 , n549 , n550 , n551 , n552 , n553 , n554 , n555 , n556 , n557 , n558 , n559 , n560 , n561 , n562 , n563 , n564 , n565 , n566 , n567 , n568 , n569 , n570 , n571 , n572 , n573 , n574 , n575 , n576 , n577 , n578 , n579 , n580 , n581 , n582 , n583 , n584 , n585 , n586 , n587 , n588 , n589 , n590 , n591 , n592 , n593 , n594 , n595 , n596 , n597 , n598 , n599 , n600 , n601 , n602 , n603 , n604 , n605 , n606 , n607 , n608 , n609 , n610 , n611 , n612 , n613 , n614 , n615 , n616 , n617 , n618 , n619 , n620 , n621 , n622 , n623 , n624 , n625 , n626 , n627 , n628 , n629 , n630 , n631 , n632 , n633 , n634 , n635 , n636 , n637 , n638 , n639 , n640 , n641 , n642 , n643 , n644 , n645 , n646 , n647 , n648 , n649 , n650 , n651 , n652 , n653 , n654 , n655 , n656 , n657 , n658 , n659 , n660 , n661 , n662 , n663 , n664 , n665 , n666 , n667 , n668 , n669 , n670 , n671 , n672 , n673 , n674 , n675 , n676 , n677 , n678 , n679 , n680 , n681 , n682 , n683 , n684 , n685 , n686 , n687 , n688 , n689 , n690 , n691 , n692 , n693 , n694 , n695 , n696 , n697 , n698 , n699 , n700 , n701 , n702 , n703 , n704 , n705 , n706 , n707 , n708 , n709 , n710 , n711 , n712 , n713 , n714 , n715 , n716 , n717 , n718 , n719 , n720 , n721 , n722 , n723 , n724 , n725 , n726 , n727 , n728 , n729 , n730 , n731 , n732 , n733 , n734 , n735 , n736 , n737 , n738 , n739 , n740 , n741 , n742 , n743 , n744 , n745 , n746 , n747 , n748 , n749 , n750 , n751 , n752 , n753 , n754 , n755 , n756 , n757 , n758 , n759 , n760 , n761 , n762 , n763 , n764 , n765 , n766 , n767 , n768 , n769 , n770 , n771 , n772 , n773 , n774 , n775 , n776 , n777 , n778 , n779 , n780 , n781 , n782 , n783 , n784 , n785 , n786 , n787 , n788 , n789 , n790 , n791 , n792 , n793 , n794 , n795 , n796 , n797 , n798 , n799 , n800 , n801 , n802 , n803 , n804 , n805 , n806 , n807 , n808 , n809 , n810 , n811 , n812 , n813 , n814 , n815 , n816 , n817 , n818 , n819 , n820 , n821 , n822 , n823 , n824 , n825 , n826 , n827 , n828 , n829 , n830 , n831 , n832 , n833 , n834 , n835 , n836 , n837 , n838 , n839 , n840 , n841 , n842 , n843 , n844 , n845 , n846 , n847 , n848 , n849 , n850 , n851 , n852 , n853 , n854 , n855 , n856 , n857 , n858 , n859 , n860 , n861 , n862 , n863 , n864 , n865 , n866 , n867 , n868 , n869 , n870 , n871 , n872 , n873 , n874 , n875 , n876 , n877 , n878 , n879 , n880 , n881 , n882 , n883 , n884 , n885 , n886 , n887 , n888 , n889 , n890 , n891 , n892 , n893 , n894 , n895 , n896 , n897 , n898 , n899 , n900 , n901 , n902 , n903 , n904 , n905 , n906 , n907 , n908 , n909 , n910 , n911 , n912 , n913 , n914 , n915 , n916 , n917 , n918 , n919 , n920 , n921 , n922 , n923 , n924 , n925 , n926 , n927 , n928 , n929 , n930 , n931 , n932 , n933 , n934 , n935 , n936 , n937 , n938 , n939 , n940 , n941 , n942 , n943 , n944 , n945 , n946 , n947 , n948 , n949 , n950 , n951 , n952 , n953 , n954 , n955 , n956 , n957 , n958 , n959 , n960 , n961 , n962 , n963 , n964 , n965 , n966 , n967 , n968 , n969 , n970 , n971 , n972 , n973 , n974 , n975 , n976 , n977 , n978 , n979 , n980 , n981 , n982 , n983 , n984 , n985 , n986 , n987 , n988 , n989 , n990 , n991 , n992 , n993 , n994 , n995 , n996 , n997 , n998 , n999 , n1000 , n1001 , n1002 , n1003 , n1004 , n1005 , n1006 , n1007 , n1008 , n1009 , n1010 , n1011 , n1012 , n1013 , n1014 , n1015 , n1016 , n1017 , n1018 , n1019 , n1020 , n1021 , n1022 , n1023 , n1024 , n1025 , n1026 , n1027 , n1028 , n1029 , n1030 , n1031 , n1032 , n1033 , n1034 , n1035 , n1036 , n1037 , n1038 , n1039 , n1040 , n1041 , n1042 , n1043 , n1044 , n1045 , n1046 , n1047 , n1048 , n1049 , n1050 , n1051 , n1052 , n1053 , n1054 , n1055 , n1056 , n1057 , n1058 , n1059 , n1060 , n1061 , n1062 , n1063 , n1064 , n1065 , n1066 , n1067 , n1068 , n1069 , n1070 , n1071 , n1072 , n1073 , n1074 , n1075 , n1076 , n1077 , n1078 , n1079 , n1080 , n1081 , n1082 , n1083 , n1084 , n1085 , n1086 , n1087 , n1088 , n1089 , n1090 , n1091 , n1092 , n1093 , n1094 , n1095 , n1096 , n1097 , n1098 , n1099 , n1100 , n1101 , n1102 , n1103 , n1104 , n1105 , n1106 , n1107 , n1108 , n1109 , n1110 , n1111 , n1112 , n1113 , n1114 , n1115 , n1116 , n1117 , n1118 , n1119 , n1120 , n1121 , n1122 , n1123 , n1124 , n1125 , n1126 , n1127 , n1128 , n1129 , n1130 , n1131 , n1132 , n1133 , n1134 , n1135 , n1136 , n1137 , n1138 , n1139 , n1140 , n1141 , n1142 , n1143 , n1144 , n1145 , n1146 , n1147 , n1148 , n1149 , n1150 , n1151 , n1152 , n1153 , n1154 , n1155 , n1156 , n1157 , n1158 , n1159 , n1160 , n1161 , n1162 , n1163 , n1164 , n1165 , n1166 , n1167 , n1168 , n1169 , n1170 , n1171 , n1172 , n1173 , n1174 , n1175 , n1176 , n1177 , n1178 , n1179 , n1180 , n1181 , n1182 , n1183 , n1184 , n1185 , n1186 , n1187 , n1188 , n1189 , n1190 , n1191 , n1192 , n1193 , n1194 , n1195 , n1196 , n1197 , n1198 , n1199 , n1200 , n1201 , n1202 , n1203 , n1204 , n1205 , n1206 , n1207 , n1208 , n1209 , n1210 , n1211 , n1212 , n1213 , n1214 , n1215 , n1216 , n1217 , n1218 , n1219 , n1220 , n1221 , n1222 , n1223 , n1224 , n1225 , n1226 , n1227 , n1228 , n1229 , n1230 , n1231 , n1232 , n1233 , n1234 , n1235 , n1236 , n1237 , n1238 , n1239 , n1240 , n1241 , n1242 , n1243 , n1244 , n1245 , n1246 , n1247 , n1248 , n1249 , n1250 , n1251 , n1252 , n1253 , n1254 , n1255 , n1256 , n1257 , n1258 , n1259 , n1260 , n1261 , n1262 , n1263 , n1264 , n1265 , n1266 , n1267 , n1268 , n1269 , n1270 , n1271 , n1272 , n1273 , n1274 , n1275 , n1276 , n1277 , n1278 , n1279 , n1280 , n1281 , n1282 , n1283 , n1284 , n1285 , n1286 , n1287 , n1288 , n1289 , n1290 , n1291 , n1292 , n1293 , n1294 , n1295 , n1296 , n1297 , n1298 , n1299 , n1300 , n1301 , n1302 , n1303 , n1304 , n1305 , n1306 , n1307 , n1308 , n1309 , n1310 , n1311 , n1312 , n1313 , n1314 , n1315 , n1316 , n1317 , n1318 , n1319 , n1320 , n1321 , n1322 , n1323 , n1324 , n1325 , n1326 , n1327 , n1328 , n1329 , n1330 , n1331 , n1332 , n1333 , n1334 , n1335 , n1336 , n1337 , n1338 , n1339 , n1340 , n1341 , n1342 , n1343 , n1344 , n1345 , n1346 , n1347 , n1348 , n1349 , n1350 , n1351 , n1352 , n1353 , n1354 , n1355 , n1356 , n1357 , n1358 , n1359 , n1360 , n1361 , n1362 , n1363 , n1364 , n1365 , n1366 , n1367 , n1368 , n1369 , n1370 , n1371 , n1372 , n1373 , n1374 , n1375 , n1376 , n1377 , n1378 , n1379 , n1380 , n1381 , n1382 , n1383 , n1384 , n1385 , n1386 , n1387 , n1388 , n1389 , n1390 , n1391 , n1392 , n1393 , n1394 , n1395 , n1396 , n1397 , n1398 , n1399 , n1400 , n1401 , n1402 , n1403 , n1404 , n1405 , n1406 , n1407 , n1408 , n1409 , n1410 , n1411 , n1412 , n1413 , n1414 , n1415 , n1416 , n1417 , n1418 , n1419 , n1420 , n1421 , n1422 , n1423 , n1424 , n1425 , n1426 , n1427 , n1428 , n1429 , n1430 , n1431 , n1432 , n1433 , n1434 , n1435 , n1436 , n1437 , n1438 , n1439 , n1440 , n1441 , n1442 , n1443 , n1444 , n1445 , n1446 , n1447 , n1448 , n1449 , n1450 , n1451 , n1452 , n1453 , n1454 , n1455 , n1456 , n1457 , n1458 , n1459 , n1460 , n1461 , n1462 , n1463 , n1464 , n1465 , n1466 , n1467 , n1468 , n1469 , n1470 , n1471 , n1472 , n1473 , n1474 , n1475 , n1476 , n1477 , n1478 , n1479 , n1480 , n1481 , n1482 , n1483 , n1484 , n1485 , n1486 , n1487 , n1488 , n1489 , n1490 , n1491 , n1492 , n1493 , n1494 , n1495 , n1496 , n1497 , n1498 , n1499 , n1500 , n1501 , n1502 , n1503 , n1504 , n1505 , n1506 , n1507 , n1508 , n1509 , n1510 , n1511 , n1512 , n1513 , n1514 , n1515 , n1516 , n1517 , n1518 , n1519 , n1520 , n1521 , n1522 , n1523 , n1524 , n1525 , n1526 , n1527 , n1528 , n1529 , n1530 , n1531 , n1532 , n1533 , n1534 , n1535 , n1536 , n1537 , n1538 , n1539 , n1540 , n1541 , n1542 , n1543 , n1544 , n1545 , n1546 , n1547 , n1548 , n1549 , n1550 , n1551 , n1552 , n1553 , n1554 , n1555 , n1556 , n1557 , n1558 , n1559 , n1560 , n1561 , n1562 , n1563 , n1564 , n1565 , n1566 , n1567 , n1568 , n1569 , n1570 , n1571 , n1572 , n1573 , n1574 , n1575 , n1576 , n1577 , n1578 , n1579 , n1580 , n1581 , n1582 , n1583 , n1584 , n1585 , n1586 , n1587 , n1588 , n1589 , n1590 , n1591 , n1592 , n1593 , n1594 , n1595 , n1596 , n1597 , n1598 , n1599 , n1600 , n1601 , n1602 , n1603 , n1604 , n1605 , n1606 , n1607 , n1608 , n1609 , n1610 , n1611 , n1612 , n1613 , n1614 , n1615 , n1616 , n1617 , n1618 , n1619 , n1620 , n1621 , n1622 , n1623 , n1624 , n1625 , n1626 , n1627 , n1628 , n1629 , n1630 , n1631 , n1632 , n1633 , n1634 , n1635 , n1636 , n1637 , n1638 , n1639 , n1640 , n1641 , n1642 , n1643 , n1644 , n1645 , n1646 , n1647 , n1648 , n1649 , n1650 , n1651 , n1652 , n1653 , n1654 , n1655 , n1656 , n1657 , n1658 , n1659 , n1660 , n1661 , n1662 , n1663 , n1664 , n1665 , n1666 , n1667 , n1668 , n1669 , n1670 , n1671 , n1672 , n1673 , n1674 , n1675 , n1676 , n1677 , n1678 , n1679 , n1680 , n1681 , n1682 , n1683 , n1684 , n1685 , n1686 , n1687 , n1688 , n1689 , n1690 , n1691 , n1692 , n1693 , n1694 , n1695 , n1696 , n1697 , n1698 , n1699 , n1700 , n1701 , n1702 , n1703 , n1704 , n1705 , n1706 , n1707 , n1708 , n1709 , n1710 , n1711 , n1712 , n1713 , n1714 , n1715 , n1716 , n1717 , n1718 , n1719 , n1720 , n1721 , n1722 , n1723 , n1724 , n1725 , n1726 , n1727 , n1728 , n1729 , n1730 , n1731 , n1732 , n1733 , n1734 , n1735 , n1736 , n1737 , n1738 , n1739 , n1740 , n1741 , n1742 , n1743 , n1744 , n1745 , n1746 , n1747 , n1748 , n1749 , n1750 , n1751 , n1752 , n1753 , n1754 , n1755 , n1756 , n1757 , n1758 , n1759 , n1760 , n1761 , n1762 , n1763 , n1764 , n1765 , n1766 , n1767 , n1768 , n1769 , n1770 , n1771 , n1772 , n1773 , n1774 , n1775 , n1776 , n1777 , n1778 , n1779 , n1780 , n1781 , n1782 , n1783 , n1784 , n1785 , n1786 , n1787 , n1788 , n1789 , n1790 , n1791 , n1792 , n1793 , n1794 , n1795 , n1796 , n1797 , n1798 , n1799 , n1800 , n1801 , n1802 , n1803 , n1804 , n1805 , n1806 , n1807 , n1808 , n1809 , n1810 , n1811 , n1812 , n1813 , n1814 , n1815 , n1816 , n1817 , n1818 , n1819 , n1820 , n1821 , n1822 , n1823 , n1824 , n1825 , n1826 , n1827 , n1828 , n1829 , n1830 , n1831 , n1832 , n1833 , n1834 , n1835 , n1836 , n1837 , n1838 , n1839 , n1840 , n1841 , n1842 , n1843 , n1844 , n1845 , n1846 , n1847 , n1848 , n1849 , n1850 , n1851 , n1852 , n1853 , n1854 , n1855 , n1856 , n1857 , n1858 , n1859 , n1860 , n1861 , n1862 , n1863 , n1864 , n1865 , n1866 , n1867 , n1868 , n1869 , n1870 , n1871 , n1872 , n1873 , n1874 , n1875 , n1876 , n1877 , n1878 , n1879 , n1880 , n1881 , n1882 , n1883 , n1884 , n1885 , n1886 , n1887 , n1888 , n1889 , n1890 , n1891 , n1892 , n1893 , n1894 , n1895 , n1896 , n1897 , n1898 , n1899 , n1900 , n1901 , n1902 , n1903 , n1904 , n1905 , n1906 , n1907 , n1908 , n1909 , n1910 , n1911 , n1912 , n1913 , n1914 , n1915 , n1916 , n1917 , n1918 , n1919 , n1920 , n1921 , n1922 , n1923 , n1924 , n1925 , n1926 , n1927 , n1928 , n1929 , n1930 , n1931 , n1932 , n1933 , n1934 , n1935 , n1936 , n1937 , n1938 , n1939 , n1940 , n1941 , n1942 , n1943 , n1944 , n1945 , n1946 , n1947 , n1948 , n1949 , n1950 , n1951 , n1952 , n1953 , n1954 , n1955 , n1956 , n1957 , n1958 , n1959 , n1960 , n1961 , n1962 , n1963 , n1964 , n1965 , n1966 , n1967 , n1968 , n1969 , n1970 , n1971 , n1972 , n1973 , n1974 , n1975 , n1976 , n1977 , n1978 , n1979 , n1980 , n1981 , n1982 , n1983 , n1984 , n1985 , n1986 , n1987 , n1988 , n1989 , n1990 , n1991 , n1992 , n1993 , n1994 , n1995 , n1996 , n1997 , n1998 , n1999 , n2000 , n2001 , n2002 , n2003 , n2004 , n2005 , n2006 , n2007 , n2008 , n2009 , n2010 , n2011 , n2012 , n2013 , n2014 , n2015 , n2016 , n2017 , n2018 , n2019 , n2020 , n2021 , n2022 , n2023 , n2024 , n2025 , n2026 , n2027 , n2028 , n2029 , n2030 , n2031 , n2032 , n2033 , n2034 , n2035 , n2036 , n2037 , n2038 , n2039 , n2040 , n2041 , n2042 , n2043 , n2044 , n2045 , n2046 , n2047 , n2048 , n2049 , n2050 , n2051 , n2052 , n2053 , n2054 , n2055 , n2056 , n2057 , n2058 , n2059 , n2060 , n2061 , n2062 , n2063 , n2064 , n2065 , n2066 , n2067 , n2068 , n2069 , n2070 , n2071 , n2072 , n2073 , n2074 , n2075 , n2076 , n2077 , n2078 , n2079 , n2080 , n2081 , n2082 , n2083 , n2084 , n2085 , n2086 , n2087 , n2088 , n2089 , n2090 , n2091 , n2092 , n2093 , n2094 , n2095 , n2096 , n2097 , n2098 , n2099 , n2100 , n2101 , n2102 , n2103 , n2104 , n2105 , n2106 , n2107 , n2108 , n2109 , n2110 , n2111 , n2112 , n2113 , n2114 , n2115 , n2116 , n2117 , n2118 , n2119 , n2120 , n2121 , n2122 , n2123 , n2124 , n2125 , n2126 , n2127 , n2128 , n2129 , n2130 , n2131 , n2132 , n2133 , n2134 , n2135 , n2136 , n2137 , n2138 , n2139 , n2140 , n2141 , n2142 , n2143 , n2144 , n2145 , n2146 , n2147 , n2148 , n2149 , n2150 , n2151 , n2152 , n2153 , n2154 , n2155 , n2156 , n2157 , n2158 , n2159 , n2160 , n2161 , n2162 , n2163 , n2164 , n2165 , n2166 , n2167 , n2168 , n2169 , n2170 , n2171 , n2172 , n2173 , n2174 , n2175 , n2176 , n2177 , n2178 , n2179 , n2180 , n2181 , n2182 , n2183 , n2184 , n2185 , n2186 , n2187 , n2188 , n2189 , n2190 , n2191 , n2192 , n2193 , n2194 , n2195 , n2196 , n2197 , n2198 , n2199 , n2200 , n2201 , n2202 , n2203 , n2204 , n2205 , n2206 , n2207 , n2208 , n2209 , n2210 , n2211 , n2212 , n2213 , n2214 , n2215 , n2216 , n2217 , n2218 , n2219 , n2220 , n2221 , n2222 , n2223 , n2224 , n2225 , n2226 , n2227 , n2228 , n2229 , n2230 , n2231 , n2232 , n2233 , n2234 , n2235 , n2236 , n2237 , n2238 , n2239 , n2240 , n2241 , n2242 , n2243 , n2244 , n2245 , n2246 , n2247 , n2248 , n2249 , n2250 , n2251 , n2252 , n2253 , n2254 , n2255 , n2256 , n2257 , n2258 , n2259 , n2260 , n2261 , n2262 , n2263 , n2264 , n2265 , n2266 , n2267 , n2268 , n2269 , n2270 , n2271 , n2272 , n2273 , n2274 , n2275 , n2276 , n2277 , n2278 , n2279 , n2280 , n2281 , n2282 , n2283 , n2284 , n2285 , n2286 , n2287 , n2288 , n2289 , n2290 , n2291 , n2292 , n2293 , n2294 , n2295 , n2296 , n2297 , n2298 , n2299 , n2300 , n2301 , n2302 , n2303 , n2304 , n2305 , n2306 , n2307 , n2308 , n2309 , n2310 , n2311 , n2312 , n2313 , n2314 , n2315 , n2316 , n2317 , n2318 , n2319 , n2320 , n2321 , n2322 , n2323 , n2324 , n2325 , n2326 , n2327 , n2328 , n2329 , n2330 , n2331 , n2332 , n2333 , n2334 , n2335 , n2336 , n2337 , n2338 , n2339 , n2340 , n2341 , n2342 , n2343 , n2344 , n2345 , n2346 , n2347 , n2348 , n2349 , n2350 , n2351 , n2352 , n2353 , n2354 , n2355 , n2356 , n2357 , n2358 , n2359 , n2360 , n2361 , n2362 , n2363 , n2364 , n2365 , n2366 , n2367 , n2368 , n2369 , n2370 , n2371 , n2372 , n2373 , n2374 , n2375 , n2376 , n2377 , n2378 , n2379 , n2380 , n2381 , n2382 , n2383 , n2384 , n2385 , n2386 , n2387 , n2388 , n2389 , n2390 , n2391 , n2392 , n2393 , n2394 , n2395 , n2396 , n2397 , n2398 , n2399 , n2400 , n2401 , n2402 , n2403 , n2404 , n2405 , n2406 , n2407 , n2408 , n2409 , n2410 , n2411 , n2412 , n2413 , n2414 , n2415 , n2416 , n2417 , n2418 , n2419 , n2420 , n2421 , n2422 , n2423 , n2424 , n2425 , n2426 , n2427 , n2428 , n2429 , n2430 , n2431 , n2432 , n2433 , n2434 , n2435 , n2436 , n2437 , n2438 , n2439 , n2440 , n2441 , n2442 , n2443 , n2444 , n2445 , n2446 , n2447 , n2448 , n2449 , n2450 , n2451 , n2452 , n2453 , n2454 , n2455 , n2456 , n2457 , n2458 , n2459 , n2460 , n2461 , n2462 , n2463 , n2464 , n2465 , n2466 , n2467 , n2468 , n2469 , n2470 , n2471 , n2472 , n2473 , n2474 , n2475 , n2476 , n2477 , n2478 , n2479 , n2480 , n2481 , n2482 , n2483 , n2484 , n2485 , n2486 , n2487 , n2488 , n2489 , n2490 , n2491 , n2492 , n2493 , n2494 , n2495 , n2496 , n2497 , n2498 , n2499 , n2500 , n2501 , n2502 , n2503 , n2504 , n2505 , n2506 , n2507 , n2508 , n2509 , n2510 , n2511 , n2512 , n2513 , n2514 , n2515 , n2516 , n2517 , n2518 , n2519 , n2520 , n2521 , n2522 , n2523 , n2524 , n2525 , n2526 , n2527 , n2528 , n2529 , n2530 , n2531 , n2532 , n2533 , n2534 , n2535 , n2536 , n2537 , n2538 , n2539 , n2540 , n2541 , n2542 , n2543 , n2544 , n2545 , n2546 , n2547 , n2548 , n2549 , n2550 , n2551 , n2552 , n2553 , n2554 , n2555 , n2556 , n2557 , n2558 , n2559 , n2560 , n2561 , n2562 , n2563 , n2564 , n2565 , n2566 , n2567 , n2568 , n2569 , n2570 , n2571 , n2572 , n2573 , n2574 , n2575 , n2576 , n2577 , n2578 , n2579 , n2580 , n2581 , n2582 , n2583 , n2584 , n2585 , n2586 , n2587 , n2588 , n2589 , n2590 , n2591 , n2592 , n2593 , n2594 , n2595 , n2596 , n2597 , n2598 , n2599 , n2600 , n2601 , n2602 , n2603 , n2604 , n2605 , n2606 , n2607 , n2608 , n2609 , n2610 , n2611 , n2612 , n2613 , n2614 , n2615 , n2616 , n2617 , n2618 , n2619 , n2620 , n2621 , n2622 , n2623 , n2624 , n2625 , n2626 , n2627 , n2628 , n2629 , n2630 , n2631 , n2632 , n2633 , n2634 , n2635 , n2636 , n2637 , n2638 , n2639 , n2640 , n2641 , n2642 , n2643 , n2644 , n2645 , n2646 , n2647 , n2648 , n2649 , n2650 , n2651 , n2652 , n2653 , n2654 , n2655 , n2656 , n2657 , n2658 , n2659 , n2660 , n2661 , n2662 , n2663 , n2664 , n2665 , n2666 , n2667 , n2668 , n2669 , n2670 , n2671 , n2672 , n2673 , n2674 , n2675 , n2676 , n2677 , n2678 , n2679 , n2680 , n2681 , n2682 , n2683 , n2684 , n2685 , n2686 , n2687 , n2688 , n2689 , n2690 , n2691 , n2692 , n2693 , n2694 , n2695 , n2696 , n2697 , n2698 , n2699 , n2700 , n2701 , n2702 , n2703 , n2704 , n2705 , n2706 , n2707 , n2708 , n2709 , n2710 , n2711 , n2712 , n2713 , n2714 , n2715 , n2716 , n2717 , n2718 , n2719 , n2720 , n2721 , n2722 , n2723 , n2724 , n2725 , n2726 , n2727 , n2728 , n2729 , n2730 , n2731 , n2732 , n2733 , n2734 , n2735 , n2736 , n2737 , n2738 , n2739 , n2740 , n2741 , n2742 , n2743 , n2744 , n2745 , n2746 , n2747 , n2748 , n2749 , n2750 , n2751 , n2752 , n2753 , n2754 , n2755 , n2756 , n2757 , n2758 , n2759 , n2760 , n2761 , n2762 , n2763 , n2764 , n2765 , n2766 , n2767 , n2768 , n2769 , n2770 , n2771 , n2772 , n2773 , n2774 , n2775 , n2776 , n2777 , n2778 , n2779 , n2780 , n2781 , n2782 , n2783 , n2784 , n2785 , n2786 , n2787 , n2788 , n2789 , n2790 , n2791 , n2792 , n2793 , n2794 , n2795 , n2796 , n2797 , n2798 , n2799 , n2800 , n2801 , n2802 , n2803 , n2804 , n2805 , n2806 , n2807 , n2808 , n2809 , n2810 , n2811 , n2812 , n2813 , n2814 , n2815 , n2816 , n2817 , n2818 , n2819 , n2820 , n2821 , n2822 , n2823 , n2824 , n2825 , n2826 , n2827 , n2828 , n2829 , n2830 , n2831 , n2832 , n2833 , n2834 , n2835 , n2836 , n2837 , n2838 , n2839 , n2840 , n2841 , n2842 , n2843 , n2844 , n2845 , n2846 , n2847 , n2848 , n2849 , n2850 , n2851 , n2852 , n2853 , n2854 , n2855 , n2856 , n2857 , n2858 , n2859 , n2860 , n2861 , n2862 , n2863 , n2864 , n2865 , n2866 , n2867 , n2868 , n2869 , n2870 , n2871 , n2872 , n2873 , n2874 , n2875 , n2876 , n2877 , n2878 , n2879 , n2880 , n2881 , n2882 , n2883 , n2884 , n2885 , n2886 , n2887 , n2888 , n2889 , n2890 , n2891 , n2892 , n2893 , n2894 , n2895 , n2896 , n2897 , n2898 , n2899 , n2900 , n2901 , n2902 , n2903 , n2904 , n2905 , n2906 , n2907 , n2908 , n2909 , n2910 , n2911 , n2912 , n2913 , n2914 , n2915 , n2916 , n2917 , n2918 , n2919 , n2920 , n2921 , n2922 , n2923 , n2924 , n2925 , n2926 , n2927 , n2928 , n2929 , n2930 , n2931 , n2932 , n2933 , n2934 , n2935 , n2936 , n2937 , n2938 , n2939 , n2940 , n2941 , n2942 , n2943 , n2944 , n2945 , n2946 , n2947 , n2948 , n2949 , n2950 , n2951 , n2952 , n2953 , n2954 , n2955 , n2956 , n2957 , n2958 , n2959 , n2960 , n2961 , n2962 , n2963 , n2964 , n2965 , n2966 , n2967 , n2968 , n2969 , n2970 , n2971 , n2972 , n2973 , n2974 , n2975 , n2976 , n2977 , n2978 , n2979 , n2980 , n2981 , n2982 , n2983 , n2984 , n2985 , n2986 , n2987 , n2988 , n2989 , n2990 , n2991 , n2992 , n2993 , n2994 , n2995 , n2996 , n2997 , n2998 , n2999 , n3000 , n3001 , n3002 , n3003 , n3004 , n3005 , n3006 , n3007 , n3008 , n3009 , n3010 , n3011 , n3012 , n3013 , n3014 , n3015 , n3016 , n3017 , n3018 , n3019 , n3020 , n3021 , n3022 , n3023 , n3024 , n3025 , n3026 , n3027 , n3028 , n3029 , n3030 , n3031 , n3032 , n3033 , n3034 , n3035 , n3036 , n3037 , n3038 , n3039 , n3040 , n3041 , n3042 , n3043 , n3044 , n3045 , n3046 , n3047 , n3048 , n3049 , n3050 , n3051 , n3052 , n3053 , n3054 , n3055 , n3056 , n3057 , n3058 , n3059 , n3060 , n3061 , n3062 , n3063 , n3064 , n3065 , n3066 , n3067 , n3068 , n3069 , n3070 , n3071 , n3072 , n3073 , n3074 , n3075 , n3076 , n3077 , n3078 , n3079 , n3080 , n3081 , n3082 , n3083 , n3084 , n3085 , n3086 , n3087 , n3088 , n3089 , n3090 , n3091 , n3092 , n3093 , n3094 , n3095 , n3096 , n3097 , n3098 , n3099 , n3100 , n3101 , n3102 , n3103 , n3104 , n3105 , n3106 , n3107 , n3108 , n3109 , n3110 , n3111 , n3112 , n3113 , n3114 , n3115 , n3116 , n3117 , n3118 , n3119 , n3120 , n3121 , n3122 , n3123 , n3124 , n3125 , n3126 , n3127 , n3128 , n3129 , n3130 , n3131 , n3132 , n3133 , n3134 , n3135 , n3136 , n3137 , n3138 , n3139 , n3140 , n3141 , n3142 , n3143 , n3144 , n3145 , n3146 , n3147 , n3148 , n3149 , n3150 , n3151 , n3152 , n3153 , n3154 , n3155 , n3156 , n3157 , n3158 , n3159 , n3160 , n3161 , n3162 , n3163 , n3164 , n3165 , n3166 , n3167 , n3168 , n3169 , n3170 , n3171 , n3172 , n3173 , n3174 , n3175 , n3176 , n3177 , n3178 , n3179 , n3180 , n3181 , n3182 , n3183 , n3184 , n3185 , n3186 , n3187 , n3188 , n3189 , n3190 , n3191 , n3192 , n3193 , n3194 , n3195 , n3196 , n3197 , n3198 , n3199 , n3200 , n3201 , n3202 , n3203 , n3204 , n3205 , n3206 , n3207 , n3208 , n3209 , n3210 , n3211 , n3212 , n3213 , n3214 , n3215 , n3216 , n3217 , n3218 , n3219 , n3220 , n3221 , n3222 , n3223 , n3224 , n3225 , n3226 , n3227 , n3228 , n3229 , n3230 , n3231 , n3232 , n3233 , n3234 , n3235 , n3236 , n3237 , n3238 , n3239 , n3240 , n3241 , n3242 , n3243 , n3244 , n3245 , n3246 , n3247 , n3248 , n3249 , n3250 , n3251 , n3252 , n3253 , n3254 , n3255 , n3256 , n3257 , n3258 , n3259 , n3260 , n3261 , n3262 , n3263 , n3264 , n3265 , n3266 , n3267 , n3268 , n3269 , n3270 , n3271 , n3272 , n3273 , n3274 , n3275 , n3276 , n3277 , n3278 , n3279 , n3280 , n3281 , n3282 , n3283 , n3284 , n3285 , n3286 , n3287 , n3288 , n3289 , n3290 , n3291 , n3292 , n3293 , n3294 , n3295 , n3296 , n3297 , n3298 , n3299 , n3300 , n3301 , n3302 , n3303 , n3304 , n3305 , n3306 , n3307 , n3308 , n3309 , n3310 , n3311 , n3312 , n3313 , n3314 , n3315 , n3316 , n3317 , n3318 , n3319 , n3320 , n3321 , n3322 , n3323 , n3324 , n3325 , n3326 , n3327 , n3328 , n3329 , n3330 , n3331 , n3332 , n3333 , n3334 , n3335 , n3336 , n3337 , n3338 , n3339 , n3340 , n3341 , n3342 , n3343 , n3344 , n3345 , n3346 , n3347 , n3348 , n3349 , n3350 , n3351 , n3352 , n3353 , n3354 , n3355 , n3356 , n3357 , n3358 , n3359 , n3360 , n3361 , n3362 , n3363 , n3364 , n3365 , n3366 , n3367 , n3368 , n3369 , n3370 , n3371 , n3372 , n3373 , n3374 , n3375 , n3376 , n3377 , n3378 , n3379 , n3380 , n3381 , n3382 , n3383 , n3384 , n3385 , n3386 , n3387 , n3388 , n3389 , n3390 , n3391 , n3392 , n3393 , n3394 , n3395 , n3396 , n3397 , n3398 , n3399 , n3400 , n3401 , n3402 , n3403 , n3404 , n3405 , n3406 , n3407 , n3408 , n3409 , n3410 , n3411 , n3412 , n3413 , n3414 , n3415 , n3416 , n3417 , n3418 , n3419 , n3420 , n3421 , n3422 , n3423 , n3424 , n3425 , n3426 , n3427 , n3428 , n3429 , n3430 , n3431 , n3432 , n3433 , n3434 , n3435 , n3436 , n3437 , n3438 , n3439 , n3440 , n3441 , n3442 , n3443 , n3444 , n3445 , n3446 , n3447 , n3448 , n3449 , n3450 , n3451 , n3452 , n3453 , n3454 , n3455 , n3456 , n3457 , n3458 , n3459 , n3460 , n3461 , n3462 , n3463 , n3464 , n3465 , n3466 , n3467 , n3468 , n3469 , n3470 , n3471 , n3472 , n3473 , n3474 , n3475 , n3476 , n3477 , n3478 , n3479 , n3480 , n3481 , n3482 , n3483 , n3484 , n3485 , n3486 , n3487 , n3488 , n3489 , n3490 , n3491 , n3492 , n3493 , n3494 , n3495 , n3496 , n3497 , n3498 , n3499 , n3500 , n3501 , n3502 , n3503 , n3504 , n3505 , n3506 , n3507 , n3508 , n3509 , n3510 , n3511 , n3512 , n3513 , n3514 , n3515 , n3516 , n3517 , n3518 , n3519 , n3520 , n3521 , n3522 , n3523 , n3524 , n3525 , n3526 , n3527 , n3528 , n3529 , n3530 , n3531 , n3532 , n3533 , n3534 , n3535 , n3536 , n3537 , n3538 , n3539 , n3540 , n3541 , n3542 , n3543 , n3544 , n3545 , n3546 , n3547 , n3548 , n3549 , n3550 , n3551 , n3552 , n3553 , n3554 , n3555 , n3556 , n3557 , n3558 , n3559 , n3560 , n3561 , n3562 , n3563 , n3564 , n3565 , n3566 , n3567 , n3568 , n3569 , n3570 , n3571 , n3572 , n3573 , n3574 , n3575 , n3576 , n3577 , n3578 , n3579 , n3580 , n3581 , n3582 , n3583 , n3584 , n3585 , n3586 , n3587 , n3588 , n3589 , n3590 , n3591 , n3592 , n3593 , n3594 , n3595 , n3596 , n3597 , n3598 , n3599 , n3600 , n3601 , n3602 , n3603 , n3604 , n3605 , n3606 , n3607 , n3608 , n3609 , n3610 , n3611 , n3612 , n3613 , n3614 , n3615 , n3616 , n3617 , n3618 , n3619 , n3620 , n3621 , n3622 , n3623 , n3624 , n3625 , n3626 , n3627 , n3628 , n3629 , n3630 , n3631 , n3632 , n3633 , n3634 , n3635 , n3636 , n3637 , n3638 , n3639 , n3640 , n3641 , n3642 , n3643 , n3644 , n3645 , n3646 , n3647 , n3648 , n3649 , n3650 , n3651 , n3652 , n3653 , n3654 , n3655 , n3656 , n3657 , n3658 , n3659 , n3660 , n3661 , n3662 , n3663 , n3664 , n3665 , n3666 , n3667 , n3668 , n3669 , n3670 , n3671 , n3672 , n3673 , n3674 , n3675 , n3676 , n3677 , n3678 , n3679 , n3680 , n3681 , n3682 , n3683 , n3684 , n3685 , n3686 , n3687 , n3688 , n3689 , n3690 , n3691 , n3692 , n3693 , n3694 , n3695 , n3696 , n3697 , n3698 , n3699 , n3700 , n3701 , n3702 , n3703 , n3704 , n3705 , n3706 , n3707 , n3708 , n3709 , n3710 , n3711 , n3712 , n3713 , n3714 , n3715 , n3716 , n3717 , n3718 , n3719 , n3720 , n3721 , n3722 , n3723 , n3724 , n3725 , n3726 , n3727 , n3728 , n3729 , n3730 , n3731 , n3732 , n3733 , n3734 , n3735 , n3736 , n3737 , n3738 , n3739 , n3740 , n3741 , n3742 , n3743 , n3744 , n3745 , n3746 , n3747 , n3748 , n3749 , n3750 , n3751 , n3752 , n3753 , n3754 , n3755 , n3756 , n3757 , n3758 , n3759 , n3760 , n3761 , n3762 , n3763 , n3764 , n3765 , n3766 , n3767 , n3768 , n3769 , n3770 , n3771 , n3772 , n3773 , n3774 , n3775 , n3776 , n3777 , n3778 , n3779 , n3780 , n3781 , n3782 , n3783 , n3784 , n3785 , n3786 , n3787 , n3788 , n3789 , n3790 , n3791 , n3792 , n3793 , n3794 , n3795 , n3796 , n3797 , n3798 , n3799 , n3800 , n3801 , n3802 , n3803 , n3804 , n3805 , n3806 , n3807 , n3808 , n3809 , n3810 , n3811 , n3812 , n3813 , n3814 , n3815 , n3816 , n3817 , n3818 , n3819 , n3820 , n3821 , n3822 , n3823 , n3824 , n3825 , n3826 , n3827 , n3828 , n3829 , n3830 , n3831 , n3832 , n3833 , n3834 , n3835 , n3836 , n3837 , n3838 , n3839 , n3840 , n3841 , n3842 , n3843 , n3844 , n3845 , n3846 , n3847 , n3848 , n3849 , n3850 , n3851 , n3852 , n3853 , n3854 , n3855 , n3856 , n3857 , n3858 , n3859 , n3860 , n3861 , n3862 , n3863 , n3864 , n3865 , n3866 , n3867 , n3868 , n3869 , n3870 , n3871 , n3872 , n3873 , n3874 , n3875 , n3876 , n3877 , n3878 , n3879 , n3880 , n3881 , n3882 , n3883 , n3884 , n3885 , n3886 , n3887 , n3888 , n3889 , n3890 , n3891 , n3892 , n3893 , n3894 , n3895 , n3896 , n3897 , n3898 , n3899 , n3900 , n3901 , n3902 , n3903 , n3904 , n3905 , n3906 , n3907 , n3908 , n3909 , n3910 , n3911 , n3912 , n3913 , n3914 , n3915 , n3916 , n3917 , n3918 , n3919 , n3920 , n3921 , n3922 , n3923 , n3924 , n3925 , n3926 , n3927 , n3928 , n3929 , n3930 , n3931 , n3932 , n3933 , n3934 , n3935 , n3936 , n3937 , n3938 , n3939 , n3940 , n3941 , n3942 , n3943 , n3944 , n3945 , n3946 , n3947 , n3948 , n3949 , n3950 , n3951 , n3952 , n3953 , n3954 , n3955 , n3956 , n3957 , n3958 , n3959 , n3960 , n3961 , n3962 , n3963 , n3964 , n3965 , n3966 , n3967 , n3968 , n3969 , n3970 , n3971 , n3972 , n3973 , n3974 , n3975 , n3976 , n3977 , n3978 , n3979 , n3980 , n3981 , n3982 , n3983 , n3984 , n3985 , n3986 , n3987 , n3988 , n3989 , n3990 , n3991 , n3992 , n3993 , n3994 , n3995 , n3996 , n3997 , n3998 , n3999 , n4000 , n4001 , n4002 , n4003 , n4004 , n4005 , n4006 , n4007 , n4008 , n4009 , n4010 , n4011 , n4012 , n4013 , n4014 , n4015 , n4016 , n4017 , n4018 , n4019 , n4020 , n4021 , n4022 , n4023 , n4024 , n4025 , n4026 , n4027 , n4028 , n4029 , n4030 , n4031 , n4032 , n4033 , n4034 , n4035 , n4036 , n4037 , n4038 , n4039 , n4040 , n4041 , n4042 , n4043 , n4044 , n4045 , n4046 , n4047 , n4048 , n4049 , n4050 , n4051 , n4052 , n4053 , n4054 , n4055 , n4056 , n4057 , n4058 , n4059 , n4060 , n4061 , n4062 , n4063 , n4064 , n4065 , n4066 , n4067 , n4068 , n4069 , n4070 , n4071 , n4072 , n4073 , n4074 , n4075 , n4076 , n4077 , n4078 , n4079 , n4080 , n4081 , n4082 , n4083 , n4084 , n4085 , n4086 , n4087 , n4088 , n4089 , n4090 , n4091 , n4092 , n4093 , n4094 , n4095 , n4096 , n4097 , n4098 , n4099 , n4100 , n4101 , n4102 , n4103 , n4104 , n4105 , n4106 , n4107 , n4108 , n4109 , n4110 , n4111 , n4112 , n4113 , n4114 , n4115 , n4116 , n4117 , n4118 , n4119 , n4120 , n4121 , n4122 , n4123 , n4124 , n4125 , n4126 , n4127 , n4128 , n4129 , n4130 , n4131 , n4132 , n4133 , n4134 , n4135 , n4136 , n4137 , n4138 , n4139 , n4140 , n4141 , n4142 , n4143 , n4144 , n4145 , n4146 , n4147 , n4148 , n4149 , n4150 , n4151 , n4152 , n4153 , n4154 , n4155 , n4156 , n4157 , n4158 , n4159 , n4160 , n4161 , n4162 , n4163 , n4164 , n4165 , n4166 , n4167 , n4168 , n4169 , n4170 , n4171 , n4172 , n4173 , n4174 , n4175 , n4176 , n4177 , n4178 , n4179 , n4180 , n4181 , n4182 , n4183 , n4184 , n4185 , n4186 , n4187 , n4188 , n4189 , n4190 , n4191 , n4192 , n4193 , n4194 , n4195 , n4196 , n4197 , n4198 , n4199 , n4200 , n4201 , n4202 , n4203 , n4204 , n4205 , n4206 , n4207 , n4208 , n4209 , n4210 , n4211 , n4212 , n4213 , n4214 , n4215 , n4216 , n4217 , n4218 , n4219 , n4220 , n4221 , n4222 , n4223 , n4224 , n4225 , n4226 , n4227 , n4228 , n4229 , n4230 , n4231 , n4232 , n4233 , n4234 , n4235 , n4236 , n4237 , n4238 , n4239 , n4240 , n4241 , n4242 , n4243 , n4244 , n4245 , n4246 , n4247 , n4248 , n4249 , n4250 , n4251 , n4252 , n4253 , n4254 , n4255 , n4256 , n4257 , n4258 , n4259 , n4260 , n4261 , n4262 , n4263 , n4264 , n4265 , n4266 , n4267 , n4268 , n4269 , n4270 , n4271 , n4272 , n4273 , n4274 , n4275 , n4276 , n4277 , n4278 , n4279 , n4280 , n4281 , n4282 , n4283 , n4284 , n4285 , n4286 , n4287 , n4288 , n4289 , n4290 , n4291 , n4292 , n4293 , n4294 , n4295 , n4296 , n4297 , n4298 , n4299 , n4300 , n4301 , n4302 , n4303 , n4304 , n4305 , n4306 , n4307 , n4308 , n4309 , n4310 , n4311 , n4312 , n4313 , n4314 , n4315 , n4316 , n4317 , n4318 , n4319 , n4320 , n4321 , n4322 , n4323 , n4324 , n4325 , n4326 , n4327 , n4328 , n4329 , n4330 , n4331 , n4332 , n4333 , n4334 , n4335 , n4336 , n4337 , n4338 , n4339 , n4340 , n4341 , n4342 , n4343 , n4344 , n4345 , n4346 , n4347 , n4348 , n4349 , n4350 , n4351 , n4352 , n4353 , n4354 , n4355 , n4356 , n4357 , n4358 , n4359 , n4360 , n4361 , n4362 , n4363 , n4364 , n4365 , n4366 , n4367 , n4368 , n4369 , n4370 , n4371 , n4372 , n4373 , n4374 , n4375 , n4376 , n4377 , n4378 , n4379 , n4380 , n4381 , n4382 , n4383 , n4384 , n4385 , n4386 , n4387 , n4388 , n4389 , n4390 , n4391 , n4392 , n4393 , n4394 , n4395 , n4396 , n4397 , n4398 , n4399 , n4400 , n4401 , n4402 , n4403 , n4404 , n4405 , n4406 , n4407 , n4408 , n4409 , n4410 , n4411 , n4412 , n4413 , n4414 , n4415 , n4416 , n4417 , n4418 , n4419 , n4420 , n4421 , n4422 , n4423 , n4424 , n4425 , n4426 , n4427 , n4428 , n4429 , n4430 , n4431 , n4432 , n4433 , n4434 , n4435 , n4436 , n4437 , n4438 , n4439 , n4440 , n4441 , n4442 , n4443 , n4444 , n4445 , n4446 , n4447 , n4448 , n4449 , n4450 , n4451 , n4452 , n4453 , n4454 , n4455 , n4456 , n4457 , n4458 , n4459 , n4460 , n4461 , n4462 , n4463 , n4464 , n4465 , n4466 , n4467 , n4468 , n4469 , n4470 , n4471 , n4472 , n4473 , n4474 , n4475 , n4476 , n4477 , n4478 , n4479 , n4480 , n4481 , n4482 , n4483 , n4484 , n4485 , n4486 , n4487 , n4488 , n4489 , n4490 , n4491 , n4492 , n4493 , n4494 , n4495 , n4496 , n4497 , n4498 , n4499 , n4500 , n4501 , n4502 , n4503 , n4504 , n4505 , n4506 , n4507 , n4508 , n4509 , n4510 , n4511 , n4512 , n4513 , n4514 , n4515 , n4516 , n4517 , n4518 , n4519 , n4520 , n4521 , n4522 , n4523 , n4524 , n4525 , n4526 , n4527 , n4528 , n4529 , n4530 , n4531 , n4532 , n4533 , n4534 , n4535 , n4536 , n4537 , n4538 , n4539 , n4540 , n4541 , n4542 , n4543 , n4544 , n4545 , n4546 , n4547 , n4548 , n4549 , n4550 , n4551 , n4552 , n4553 , n4554 , n4555 , n4556 , n4557 , n4558 , n4559 , n4560 , n4561 , n4562 , n4563 , n4564 , n4565 , n4566 , n4567 , n4568 , n4569 , n4570 , n4571 , n4572 , n4573 , n4574 , n4575 , n4576 , n4577 , n4578 , n4579 , n4580 , n4581 , n4582 , n4583 , n4584 , n4585 , n4586 , n4587 , n4588 , n4589 , n4590 , n4591 , n4592 , n4593 , n4594 , n4595 , n4596 , n4597 , n4598 , n4599 , n4600 , n4601 , n4602 , n4603 , n4604 , n4605 , n4606 , n4607 , n4608 , n4609 , n4610 , n4611 , n4612 , n4613 , n4614 , n4615 , n4616 , n4617 , n4618 , n4619 , n4620 , n4621 , n4622 , n4623 , n4624 , n4625 , n4626 , n4627 , n4628 , n4629 , n4630 , n4631 , n4632 , n4633 , n4634 , n4635 , n4636 , n4637 , n4638 , n4639 , n4640 , n4641 , n4642 , n4643 , n4644 , n4645 , n4646 , n4647 , n4648 , n4649 , n4650 , n4651 , n4652 , n4653 , n4654 , n4655 , n4656 , n4657 , n4658 , n4659 , n4660 , n4661 , n4662 , n4663 , n4664 , n4665 , n4666 , n4667 , n4668 , n4669 , n4670 , n4671 , n4672 , n4673 , n4674 , n4675 , n4676 , n4677 , n4678 , n4679 , n4680 , n4681 , n4682 , n4683 , n4684 , n4685 , n4686 , n4687 , n4688 , n4689 , n4690 , n4691 , n4692 , n4693 , n4694 , n4695 , n4696 , n4697 , n4698 , n4699 , n4700 , n4701 , n4702 , n4703 , n4704 , n4705 , n4706 , n4707 , n4708 , n4709 , n4710 , n4711 , n4712 , n4713 , n4714 , n4715 , n4716 , n4717 , n4718 , n4719 , n4720 , n4721 , n4722 , n4723 , n4724 , n4725 , n4726 , n4727 , n4728 , n4729 , n4730 , n4731 , n4732 , n4733 , n4734 , n4735 , n4736 , n4737 , n4738 , n4739 , n4740 , n4741 , n4742 , n4743 , n4744 , n4745 , n4746 , n4747 , n4748 , n4749 , n4750 , n4751 , n4752 , n4753 , n4754 , n4755 , n4756 , n4757 , n4758 , n4759 , n4760 , n4761 , n4762 , n4763 , n4764 , n4765 , n4766 , n4767 , n4768 , n4769 , n4770 , n4771 , n4772 , n4773 , n4774 , n4775 , n4776 , n4777 , n4778 , n4779 , n4780 , n4781 , n4782 , n4783 , n4784 , n4785 , n4786 , n4787 , n4788 , n4789 , n4790 , n4791 , n4792 , n4793 , n4794 , n4795 , n4796 , n4797 , n4798 , n4799 , n4800 , n4801 , n4802 , n4803 , n4804 , n4805 , n4806 , n4807 , n4808 , n4809 , n4810 , n4811 , n4812 , n4813 , n4814 , n4815 , n4816 , n4817 , n4818 , n4819 , n4820 , n4821 , n4822 , n4823 , n4824 , n4825 , n4826 , n4827 , n4828 , n4829 , n4830 , n4831 , n4832 , n4833 , n4834 , n4835 , n4836 , n4837 , n4838 , n4839 , n4840 , n4841 , n4842 , n4843 , n4844 , n4845 , n4846 , n4847 , n4848 , n4849 , n4850 , n4851 , n4852 , n4853 , n4854 , n4855 , n4856 , n4857 , n4858 , n4859 , n4860 , n4861 , n4862 , n4863 , n4864 , n4865 , n4866 , n4867 , n4868 , n4869 , n4870 , n4871 , n4872 , n4873 , n4874 , n4875 , n4876 , n4877 , n4878 , n4879 , n4880 , n4881 , n4882 , n4883 , n4884 , n4885 , n4886 , n4887 , n4888 , n4889 , n4890 , n4891 , n4892 , n4893 , n4894 , n4895 , n4896 , n4897 , n4898 , n4899 , n4900 , n4901 , n4902 , n4903 , n4904 , n4905 , n4906 , n4907 , n4908 , n4909 , n4910 , n4911 , n4912 , n4913 , n4914 , n4915 , n4916 , n4917 , n4918 , n4919 , n4920 , n4921 , n4922 , n4923 , n4924 , n4925 , n4926 , n4927 , n4928 , n4929 , n4930 , n4931 , n4932 , n4933 , n4934 , n4935 , n4936 , n4937 , n4938 , n4939 , n4940 , n4941 , n4942 , n4943 , n4944 , n4945 , n4946 , n4947 , n4948 , n4949 , n4950 , n4951 , n4952 , n4953 , n4954 , n4955 , n4956 , n4957 , n4958 , n4959 , n4960 , n4961 , n4962 , n4963 , n4964 , n4965 , n4966 , n4967 , n4968 , n4969 , n4970 , n4971 , n4972 , n4973 , n4974 , n4975 , n4976 , n4977 , n4978 , n4979 , n4980 , n4981 , n4982 , n4983 , n4984 , n4985 , n4986 , n4987 , n4988 , n4989 , n4990 , n4991 , n4992 , n4993 , n4994 , n4995 , n4996 , n4997 , n4998 , n4999 , n5000 , n5001 , n5002 , n5003 , n5004 , n5005 , n5006 , n5007 , n5008 , n5009 , n5010 , n5011 , n5012 , n5013 , n5014 , n5015 , n5016 , n5017 , n5018 , n5019 , n5020 , n5021 , n5022 , n5023 , n5024 , n5025 , n5026 , n5027 , n5028 , n5029 , n5030 , n5031 , n5032 , n5033 , n5034 , n5035 , n5036 , n5037 , n5038 , n5039 , n5040 , n5041 , n5042 , n5043 , n5044 , n5045 , n5046 , n5047 , n5048 , n5049 , n5050 , n5051 , n5052 , n5053 , n5054 , n5055 , n5056 , n5057 , n5058 , n5059 , n5060 , n5061 , n5062 , n5063 , n5064 , n5065 , n5066 , n5067 , n5068 , n5069 , n5070 , n5071 , n5072 , n5073 , n5074 , n5075 , n5076 , n5077 , n5078 , n5079 , n5080 , n5081 , n5082 , n5083 , n5084 , n5085 , n5086 , n5087 , n5088 , n5089 , n5090 , n5091 , n5092 , n5093 , n5094 , n5095 , n5096 , n5097 , n5098 , n5099 , n5100 , n5101 , n5102 , n5103 , n5104 , n5105 , n5106 , n5107 , n5108 , n5109 , n5110 , n5111 , n5112 , n5113 , n5114 , n5115 , n5116 , n5117 , n5118 , n5119 , n5120 , n5121 , n5122 , n5123 , n5124 , n5125 , n5126 , n5127 , n5128 , n5129 , n5130 , n5131 , n5132 , n5133 , n5134 , n5135 , n5136 , n5137 , n5138 , n5139 , n5140 , n5141 , n5142 , n5143 , n5144 , n5145 , n5146 , n5147 , n5148 , n5149 , n5150 , n5151 , n5152 , n5153 , n5154 , n5155 , n5156 , n5157 , n5158 , n5159 , n5160 , n5161 , n5162 , n5163 , n5164 , n5165 , n5166 , n5167 , n5168 , n5169 , n5170 , n5171 , n5172 , n5173 , n5174 , n5175 , n5176 , n5177 , n5178 , n5179 , n5180 , n5181 , n5182 , n5183 , n5184 , n5185 , n5186 , n5187 , n5188 , n5189 , n5190 , n5191 , n5192 , n5193 , n5194 , n5195 , n5196 , n5197 , n5198 , n5199 , n5200 , n5201 , n5202 , n5203 , n5204 , n5205 , n5206 , n5207 , n5208 , n5209 , n5210 , n5211 , n5212 , n5213 , n5214 , n5215 , n5216 , n5217 , n5218 , n5219 , n5220 , n5221 , n5222 , n5223 , n5224 , n5225 , n5226 , n5227 , n5228 , n5229 , n5230 , n5231 , n5232 , n5233 , n5234 , n5235 , n5236 , n5237 , n5238 , n5239 , n5240 , n5241 , n5242 , n5243 , n5244 , n5245 , n5246 , n5247 , n5248 , n5249 , n5250 , n5251 , n5252 , n5253 , n5254 , n5255 , n5256 , n5257 , n5258 , n5259 , n5260 , n5261 , n5262 , n5263 , n5264 , n5265 , n5266 , n5267 , n5268 , n5269 , n5270 , n5271 , n5272 , n5273 , n5274 , n5275 , n5276 , n5277 , n5278 , n5279 , n5280 , n5281 , n5282 , n5283 , n5284 , n5285 , n5286 , n5287 , n5288 , n5289 , n5290 , n5291 , n5292 , n5293 , n5294 , n5295 , n5296 , n5297 , n5298 , n5299 , n5300 , n5301 , n5302 , n5303 , n5304 , n5305 , n5306 , n5307 , n5308 , n5309 , n5310 , n5311 , n5312 , n5313 , n5314 , n5315 , n5316 , n5317 , n5318 , n5319 , n5320 , n5321 , n5322 , n5323 , n5324 , n5325 , n5326 , n5327 , n5328 , n5329 , n5330 , n5331 , n5332 , n5333 , n5334 , n5335 , n5336 , n5337 , n5338 , n5339 , n5340 , n5341 , n5342 , n5343 , n5344 , n5345 , n5346 , n5347 , n5348 , n5349 , n5350 , n5351 , n5352 , n5353 , n5354 , n5355 , n5356 , n5357 , n5358 , n5359 , n5360 , n5361 , n5362 , n5363 , n5364 , n5365 , n5366 , n5367 , n5368 , n5369 , n5370 , n5371 , n5372 , n5373 , n5374 , n5375 , n5376 , n5377 , n5378 , n5379 , n5380 , n5381 , n5382 , n5383 , n5384 , n5385 , n5386 , n5387 , n5388 , n5389 , n5390 , n5391 , n5392 , n5393 , n5394 , n5395 , n5396 , n5397 , n5398 , n5399 , n5400 , n5401 , n5402 , n5403 , n5404 , n5405 , n5406 , n5407 , n5408 , n5409 , n5410 , n5411 , n5412 , n5413 , n5414 , n5415 , n5416 , n5417 , n5418 , n5419 , n5420 , n5421 , n5422 , n5423 , n5424 , n5425 , n5426 , n5427 , n5428 , n5429 , n5430 , n5431 , n5432 , n5433 , n5434 , n5435 , n5436 , n5437 , n5438 , n5439 , n5440 , n5441 , n5442 , n5443 , n5444 , n5445 , n5446 , n5447 , n5448 , n5449 , n5450 , n5451 , n5452 , n5453 , n5454 , n5455 , n5456 , n5457 , n5458 , n5459 , n5460 , n5461 , n5462 , n5463 , n5464 , n5465 , n5466 , n5467 , n5468 , n5469 , n5470 , n5471 , n5472 , n5473 , n5474 , n5475 , n5476 , n5477 , n5478 , n5479 , n5480 , n5481 , n5482 , n5483 , n5484 , n5485 , n5486 , n5487 , n5488 , n5489 , n5490 , n5491 , n5492 , n5493 , n5494 , n5495 , n5496 , n5497 , n5498 , n5499 , n5500 , n5501 , n5502 , n5503 , n5504 , n5505 , n5506 , n5507 , n5508 , n5509 , n5510 , n5511 , n5512 , n5513 , n5514 , n5515 , n5516 , n5517 , n5518 , n5519 , n5520 , n5521 , n5522 , n5523 , n5524 , n5525 , n5526 , n5527 , n5528 , n5529 , n5530 , n5531 , n5532 , n5533 , n5534 , n5535 , n5536 , n5537 , n5538 , n5539 , n5540 , n5541 , n5542 , n5543 , n5544 , n5545 , n5546 , n5547 , n5548 , n5549 , n5550 , n5551 , n5552 , n5553 , n5554 , n5555 , n5556 , n5557 , n5558 , n5559 , n5560 , n5561 , n5562 , n5563 , n5564 , n5565 , n5566 , n5567 , n5568 , n5569 , n5570 , n5571 , n5572 , n5573 , n5574 , n5575 , n5576 , n5577 , n5578 , n5579 , n5580 , n5581 , n5582 , n5583 , n5584 , n5585 , n5586 , n5587 , n5588 , n5589 , n5590 , n5591 , n5592 , n5593 , n5594 , n5595 , n5596 , n5597 , n5598 , n5599 , n5600 , n5601 , n5602 , n5603 , n5604 , n5605 , n5606 , n5607 , n5608 , n5609 , n5610 , n5611 , n5612 , n5613 , n5614 , n5615 , n5616 , n5617 , n5618 , n5619 , n5620 , n5621 , n5622 , n5623 , n5624 , n5625 , n5626 , n5627 , n5628 , n5629 , n5630 , n5631 , n5632 , n5633 , n5634 , n5635 , n5636 , n5637 , n5638 , n5639 , n5640 , n5641 , n5642 , n5643 , n5644 , n5645 , n5646 , n5647 , n5648 , n5649 , n5650 , n5651 , n5652 , n5653 , n5654 , n5655 , n5656 , n5657 , n5658 , n5659 , n5660 , n5661 , n5662 , n5663 , n5664 , n5665 , n5666 , n5667 , n5668 , n5669 , n5670 , n5671 , n5672 , n5673 , n5674 , n5675 , n5676 , n5677 , n5678 , n5679 , n5680 , n5681 , n5682 , n5683 , n5684 , n5685 , n5686 , n5687 , n5688 , n5689 , n5690 , n5691 , n5692 , n5693 , n5694 , n5695 , n5696 , n5697 , n5698 , n5699 , n5700 , n5701 , n5702 , n5703 , n5704 , n5705 , n5706 , n5707 , n5708 , n5709 , n5710 , n5711 , n5712 , n5713 , n5714 , n5715 , n5716 , n5717 , n5718 , n5719 , n5720 , n5721 , n5722 , n5723 , n5724 , n5725 , n5726 , n5727 , n5728 , n5729 , n5730 , n5731 , n5732 , n5733 , n5734 , n5735 , n5736 , n5737 , n5738 , n5739 , n5740 , n5741 , n5742 , n5743 , n5744 , n5745 , n5746 , n5747 , n5748 , n5749 , n5750 , n5751 , n5752 , n5753 , n5754 , n5755 , n5756 , n5757 , n5758 , n5759 , n5760 , n5761 , n5762 , n5763 , n5764 , n5765 , n5766 , n5767 , n5768 , n5769 , n5770 , n5771 , n5772 , n5773 , n5774 , n5775 , n5776 , n5777 , n5778 , n5779 , n5780 , n5781 , n5782 , n5783 , n5784 , n5785 , n5786 , n5787 , n5788 , n5789 , n5790 , n5791 , n5792 , n5793 , n5794 , n5795 , n5796 , n5797 , n5798 , n5799 , n5800 , n5801 , n5802 , n5803 , n5804 , n5805 , n5806 , n5807 , n5808 , n5809 , n5810 , n5811 , n5812 , n5813 , n5814 , n5815 , n5816 , n5817 , n5818 , n5819 , n5820 , n5821 , n5822 , n5823 , n5824 , n5825 , n5826 , n5827 , n5828 , n5829 , n5830 , n5831 , n5832 , n5833 , n5834 , n5835 , n5836 , n5837 , n5838 , n5839 , n5840 , n5841 , n5842 , n5843 , n5844 , n5845 , n5846 , n5847 , n5848 , n5849 , n5850 , n5851 , n5852 , n5853 , n5854 , n5855 , n5856 , n5857 , n5858 , n5859 , n5860 , n5861 , n5862 , n5863 , n5864 , n5865 , n5866 , n5867 , n5868 , n5869 , n5870 , n5871 , n5872 , n5873 , n5874 , n5875 , n5876 , n5877 , n5878 , n5879 , n5880 , n5881 , n5882 , n5883 , n5884 , n5885 , n5886 , n5887 , n5888 , n5889 , n5890 , n5891 , n5892 , n5893 , n5894 , n5895 , n5896 , n5897 , n5898 , n5899 , n5900 , n5901 , n5902 , n5903 , n5904 , n5905 , n5906 , n5907 , n5908 , n5909 , n5910 , n5911 , n5912 , n5913 , n5914 , n5915 , n5916 , n5917 , n5918 , n5919 , n5920 , n5921 , n5922 , n5923 , n5924 , n5925 , n5926 , n5927 , n5928 , n5929 , n5930 , n5931 , n5932 , n5933 , n5934 , n5935 , n5936 , n5937 , n5938 , n5939 , n5940 , n5941 , n5942 , n5943 , n5944 , n5945 , n5946 , n5947 , n5948 , n5949 , n5950 , n5951 , n5952 , n5953 , n5954 , n5955 , n5956 , n5957 , n5958 , n5959 , n5960 , n5961 , n5962 , n5963 , n5964 , n5965 , n5966 , n5967 , n5968 , n5969 , n5970 , n5971 , n5972 , n5973 , n5974 , n5975 , n5976 , n5977 , n5978 , n5979 , n5980 , n5981 , n5982 , n5983 , n5984 , n5985 , n5986 , n5987 , n5988 , n5989 , n5990 , n5991 , n5992 , n5993 , n5994 , n5995 , n5996 , n5997 , n5998 , n5999 , n6000 , n6001 , n6002 , n6003 , n6004 , n6005 , n6006 , n6007 , n6008 , n6009 , n6010 , n6011 , n6012 , n6013 , n6014 , n6015 , n6016 , n6017 , n6018 , n6019 , n6020 , n6021 , n6022 , n6023 , n6024 , n6025 , n6026 , n6027 , n6028 , n6029 , n6030 , n6031 , n6032 , n6033 , n6034 , n6035 , n6036 , n6037 , n6038 , n6039 , n6040 , n6041 , n6042 , n6043 , n6044 , n6045 , n6046 , n6047 , n6048 , n6049 , n6050 , n6051 , n6052 , n6053 , n6054 , n6055 , n6056 , n6057 , n6058 , n6059 , n6060 , n6061 , n6062 , n6063 , n6064 , n6065 , n6066 , n6067 , n6068 , n6069 , n6070 , n6071 , n6072 , n6073 , n6074 , n6075 , n6076 , n6077 , n6078 , n6079 , n6080 , n6081 , n6082 , n6083 , n6084 , n6085 , n6086 , n6087 , n6088 , n6089 , n6090 , n6091 , n6092 , n6093 , n6094 , n6095 , n6096 , n6097 , n6098 , n6099 , n6100 , n6101 , n6102 , n6103 , n6104 , n6105 , n6106 , n6107 , n6108 , n6109 , n6110 , n6111 , n6112 , n6113 , n6114 , n6115 , n6116 , n6117 , n6118 , n6119 , n6120 , n6121 , n6122 , n6123 , n6124 , n6125 , n6126 , n6127 , n6128 , n6129 , n6130 , n6131 , n6132 , n6133 , n6134 , n6135 , n6136 , n6137 , n6138 , n6139 , n6140 , n6141 , n6142 , n6143 , n6144 , n6145 , n6146 , n6147 , n6148 , n6149 , n6150 , n6151 , n6152 , n6153 , n6154 , n6155 , n6156 , n6157 , n6158 , n6159 , n6160 , n6161 , n6162 , n6163 , n6164 , n6165 , n6166 , n6167 , n6168 , n6169 , n6170 , n6171 , n6172 , n6173 , n6174 , n6175 , n6176 , n6177 , n6178 , n6179 , n6180 , n6181 , n6182 , n6183 , n6184 , n6185 , n6186 , n6187 , n6188 , n6189 , n6190 , n6191 , n6192 , n6193 , n6194 , n6195 , n6196 , n6197 , n6198 , n6199 , n6200 , n6201 , n6202 , n6203 , n6204 , n6205 , n6206 , n6207 , n6208 , n6209 , n6210 , n6211 , n6212 , n6213 , n6214 , n6215 , n6216 , n6217 , n6218 , n6219 , n6220 , n6221 , n6222 , n6223 , n6224 , n6225 , n6226 , n6227 , n6228 , n6229 , n6230 , n6231 , n6232 , n6233 , n6234 , n6235 , n6236 , n6237 , n6238 , n6239 , n6240 , n6241 , n6242 , n6243 , n6244 , n6245 , n6246 , n6247 , n6248 , n6249 , n6250 , n6251 , n6252 , n6253 , n6254 , n6255 , n6256 , n6257 , n6258 , n6259 , n6260 , n6261 , n6262 , n6263 , n6264 , n6265 , n6266 , n6267 , n6268 , n6269 , n6270 , n6271 , n6272 , n6273 , n6274 , n6275 , n6276 , n6277 , n6278 , n6279 , n6280 , n6281 , n6282 , n6283 , n6284 , n6285 , n6286 , n6287 , n6288 , n6289 , n6290 , n6291 , n6292 , n6293 , n6294 , n6295 , n6296 , n6297 , n6298 , n6299 , n6300 , n6301 , n6302 , n6303 , n6304 , n6305 , n6306 , n6307 , n6308 , n6309 , n6310 , n6311 , n6312 , n6313 , n6314 , n6315 , n6316 , n6317 , n6318 , n6319 , n6320 , n6321 , n6322 , n6323 , n6324 , n6325 , n6326 , n6327 , n6328 , n6329 , n6330 , n6331 , n6332 , n6333 , n6334 , n6335 , n6336 , n6337 , n6338 , n6339 , n6340 , n6341 , n6342 , n6343 , n6344 , n6345 , n6346 , n6347 , n6348 , n6349 , n6350 , n6351 , n6352 , n6353 , n6354 , n6355 , n6356 , n6357 , n6358 , n6359 , n6360 , n6361 , n6362 , n6363 , n6364 , n6365 , n6366 , n6367 , n6368 , n6369 , n6370 , n6371 , n6372 , n6373 , n6374 , n6375 , n6376 , n6377 , n6378 , n6379 , n6380 , n6381 , n6382 , n6383 , n6384 , n6385 , n6386 , n6387 , n6388 , n6389 , n6390 , n6391 , n6392 , n6393 , n6394 , n6395 , n6396 , n6397 , n6398 , n6399 , n6400 , n6401 , n6402 , n6403 , n6404 , n6405 , n6406 , n6407 , n6408 , n6409 , n6410 , n6411 , n6412 , n6413 , n6414 , n6415 , n6416 , n6417 , n6418 , n6419 , n6420 , n6421 , n6422 , n6423 , n6424 , n6425 , n6426 , n6427 , n6428 , n6429 , n6430 , n6431 , n6432 , n6433 , n6434 , n6435 , n6436 , n6437 , n6438 , n6439 , n6440 , n6441 , n6442 , n6443 , n6444 , n6445 , n6446 , n6447 , n6448 , n6449 , n6450 , n6451 , n6452 , n6453 , n6454 , n6455 , n6456 , n6457 , n6458 , n6459 , n6460 , n6461 , n6462 , n6463 , n6464 , n6465 , n6466 , n6467 , n6468 , n6469 , n6470 , n6471 , n6472 , n6473 , n6474 , n6475 , n6476 , n6477 , n6478 , n6479 , n6480 , n6481 , n6482 , n6483 , n6484 , n6485 , n6486 , n6487 , n6488 , n6489 , n6490 , n6491 , n6492 , n6493 , n6494 , n6495 , n6496 , n6497 , n6498 , n6499 , n6500 , n6501 , n6502 , n6503 , n6504 , n6505 , n6506 , n6507 , n6508 , n6509 , n6510 , n6511 , n6512 , n6513 , n6514 , n6515 , n6516 , n6517 , n6518 , n6519 , n6520 , n6521 , n6522 , n6523 , n6524 , n6525 , n6526 , n6527 , n6528 , n6529 , n6530 , n6531 , n6532 , n6533 , n6534 , n6535 , n6536 , n6537 , n6538 , n6539 , n6540 , n6541 , n6542 , n6543 , n6544 , n6545 , n6546 , n6547 , n6548 , n6549 , n6550 , n6551 , n6552 , n6553 , n6554 , n6555 , n6556 , n6557 , n6558 , n6559 , n6560 , n6561 , n6562 , n6563 , n6564 , n6565 , n6566 , n6567 , n6568 , n6569 , n6570 , n6571 , n6572 , n6573 , n6574 , n6575 , n6576 , n6577 , n6578 , n6579 , n6580 , n6581 , n6582 , n6583 , n6584 , n6585 , n6586 , n6587 , n6588 , n6589 , n6590 , n6591 , n6592 , n6593 , n6594 , n6595 , n6596 , n6597 , n6598 , n6599 , n6600 , n6601 , n6602 , n6603 , n6604 , n6605 , n6606 , n6607 , n6608 , n6609 , n6610 , n6611 , n6612 , n6613 , n6614 , n6615 , n6616 , n6617 , n6618 , n6619 , n6620 , n6621 , n6622 , n6623 , n6624 , n6625 , n6626 , n6627 , n6628 , n6629 , n6630 , n6631 , n6632 , n6633 , n6634 , n6635 , n6636 , n6637 , n6638 , n6639 , n6640 , n6641 , n6642 , n6643 , n6644 , n6645 , n6646 , n6647 , n6648 , n6649 , n6650 , n6651 , n6652 , n6653 , n6654 , n6655 , n6656 , n6657 , n6658 , n6659 , n6660 , n6661 , n6662 , n6663 , n6664 , n6665 , n6666 , n6667 , n6668 , n6669 , n6670 , n6671 , n6672 , n6673 , n6674 , n6675 , n6676 , n6677 , n6678 , n6679 , n6680 , n6681 , n6682 , n6683 , n6684 , n6685 , n6686 , n6687 , n6688 , n6689 , n6690 , n6691 , n6692 , n6693 , n6694 , n6695 , n6696 , n6697 , n6698 , n6699 , n6700 , n6701 , n6702 , n6703 , n6704 , n6705 , n6706 , n6707 , n6708 , n6709 , n6710 , n6711 , n6712 , n6713 , n6714 , n6715 , n6716 , n6717 , n6718 , n6719 , n6720 , n6721 , n6722 , n6723 , n6724 , n6725 , n6726 , n6727 , n6728 , n6729 , n6730 , n6731 , n6732 , n6733 , n6734 , n6735 , n6736 , n6737 , n6738 , n6739 , n6740 , n6741 , n6742 , n6743 , n6744 , n6745 , n6746 , n6747 , n6748 , n6749 , n6750 , n6751 , n6752 , n6753 , n6754 , n6755 , n6756 , n6757 , n6758 , n6759 , n6760 , n6761 , n6762 , n6763 , n6764 , n6765 , n6766 , n6767 , n6768 , n6769 , n6770 , n6771 , n6772 , n6773 , n6774 , n6775 , n6776 , n6777 , n6778 , n6779 , n6780 , n6781 , n6782 , n6783 , n6784 , n6785 , n6786 , n6787 , n6788 , n6789 , n6790 , n6791 , n6792 , n6793 , n6794 , n6795 , n6796 , n6797 , n6798 , n6799 , n6800 , n6801 , n6802 , n6803 , n6804 , n6805 , n6806 , n6807 , n6808 , n6809 , n6810 , n6811 , n6812 , n6813 , n6814 , n6815 , n6816 , n6817 , n6818 , n6819 , n6820 , n6821 , n6822 , n6823 , n6824 , n6825 , n6826 , n6827 , n6828 , n6829 , n6830 , n6831 , n6832 , n6833 , n6834 , n6835 , n6836 , n6837 , n6838 , n6839 , n6840 , n6841 , n6842 , n6843 , n6844 , n6845 , n6846 , n6847 , n6848 , n6849 , n6850 , n6851 , n6852 , n6853 , n6854 , n6855 , n6856 , n6857 , n6858 , n6859 , n6860 , n6861 , n6862 , n6863 , n6864 , n6865 , n6866 , n6867 , n6868 , n6869 , n6870 , n6871 , n6872 , n6873 , n6874 , n6875 , n6876 , n6877 , n6878 , n6879 , n6880 , n6881 , n6882 , n6883 , n6884 , n6885 , n6886 , n6887 , n6888 , n6889 , n6890 , n6891 , n6892 , n6893 , n6894 , n6895 , n6896 , n6897 , n6898 , n6899 , n6900 , n6901 , n6902 , n6903 , n6904 , n6905 , n6906 , n6907 , n6908 , n6909 , n6910 , n6911 , n6912 , n6913 , n6914 , n6915 , n6916 , n6917 , n6918 , n6919 , n6920 , n6921 , n6922 , n6923 , n6924 , n6925 , n6926 , n6927 , n6928 , n6929 , n6930 , n6931 , n6932 , n6933 , n6934 , n6935 , n6936 , n6937 , n6938 , n6939 , n6940 , n6941 , n6942 , n6943 , n6944 , n6945 , n6946 , n6947 , n6948 , n6949 , n6950 , n6951 , n6952 , n6953 , n6954 , n6955 , n6956 , n6957 , n6958 , n6959 , n6960 , n6961 , n6962 , n6963 , n6964 , n6965 , n6966 , n6967 , n6968 , n6969 , n6970 , n6971 , n6972 , n6973 , n6974 , n6975 , n6976 , n6977 , n6978 , n6979 , n6980 , n6981 , n6982 , n6983 , n6984 , n6985 , n6986 , n6987 , n6988 , n6989 , n6990 , n6991 , n6992 , n6993 , n6994 , n6995 , n6996 , n6997 , n6998 , n6999 , n7000 , n7001 , n7002 , n7003 , n7004 , n7005 , n7006 , n7007 , n7008 , n7009 , n7010 , n7011 , n7012 , n7013 , n7014 , n7015 , n7016 , n7017 , n7018 , n7019 , n7020 , n7021 , n7022 , n7023 , n7024 , n7025 , n7026 , n7027 , n7028 , n7029 , n7030 , n7031 , n7032 , n7033 , n7034 , n7035 , n7036 , n7037 , n7038 , n7039 , n7040 , n7041 , n7042 , n7043 , n7044 , n7045 , n7046 , n7047 , n7048 , n7049 , n7050 , n7051 , n7052 , n7053 , n7054 , n7055 , n7056 , n7057 , n7058 , n7059 , n7060 , n7061 , n7062 , n7063 , n7064 , n7065 , n7066 , n7067 , n7068 , n7069 , n7070 , n7071 , n7072 , n7073 , n7074 , n7075 , n7076 , n7077 , n7078 , n7079 , n7080 , n7081 , n7082 , n7083 , n7084 , n7085 , n7086 , n7087 , n7088 , n7089 , n7090 , n7091 , n7092 , n7093 , n7094 , n7095 , n7096 , n7097 , n7098 , n7099 , n7100 , n7101 , n7102 , n7103 , n7104 , n7105 , n7106 , n7107 , n7108 , n7109 , n7110 , n7111 , n7112 , n7113 , n7114 , n7115 , n7116 , n7117 , n7118 , n7119 , n7120 , n7121 , n7122 , n7123 , n7124 , n7125 , n7126 , n7127 , n7128 , n7129 , n7130 , n7131 , n7132 , n7133 , n7134 , n7135 , n7136 , n7137 , n7138 , n7139 , n7140 , n7141 , n7142 , n7143 , n7144 , n7145 , n7146 , n7147 , n7148 , n7149 , n7150 , n7151 , n7152 , n7153 , n7154 , n7155 , n7156 , n7157 , n7158 , n7159 , n7160 , n7161 , n7162 , n7163 , n7164 , n7165 , n7166 , n7167 , n7168 , n7169 , n7170 , n7171 , n7172 , n7173 , n7174 , n7175 , n7176 , n7177 , n7178 , n7179 , n7180 , n7181 , n7182 , n7183 , n7184 , n7185 , n7186 , n7187 , n7188 , n7189 , n7190 , n7191 , n7192 , n7193 , n7194 , n7195 , n7196 , n7197 , n7198 , n7199 , n7200 , n7201 , n7202 , n7203 , n7204 , n7205 , n7206 , n7207 , n7208 , n7209 , n7210 , n7211 , n7212 , n7213 , n7214 , n7215 , n7216 , n7217 , n7218 , n7219 , n7220 , n7221 , n7222 , n7223 , n7224 , n7225 , n7226 , n7227 , n7228 , n7229 , n7230 , n7231 , n7232 , n7233 , n7234 , n7235 , n7236 , n7237 , n7238 , n7239 , n7240 , n7241 , n7242 , n7243 , n7244 , n7245 , n7246 , n7247 , n7248 , n7249 , n7250 , n7251 , n7252 , n7253 , n7254 , n7255 , n7256 , n7257 , n7258 , n7259 , n7260 , n7261 , n7262 , n7263 , n7264 , n7265 , n7266 , n7267 , n7268 , n7269 , n7270 , n7271 , n7272 , n7273 , n7274 , n7275 , n7276 , n7277 , n7278 , n7279 , n7280 , n7281 , n7282 , n7283 , n7284 , n7285 , n7286 , n7287 , n7288 , n7289 , n7290 , n7291 , n7292 , n7293 , n7294 , n7295 , n7296 , n7297 , n7298 , n7299 , n7300 , n7301 , n7302 , n7303 , n7304 , n7305 , n7306 , n7307 , n7308 , n7309 , n7310 , n7311 , n7312 , n7313 , n7314 , n7315 , n7316 , n7317 , n7318 , n7319 , n7320 , n7321 , n7322 , n7323 , n7324 , n7325 , n7326 , n7327 , n7328 , n7329 , n7330 , n7331 , n7332 , n7333 , n7334 , n7335 , n7336 , n7337 , n7338 , n7339 , n7340 , n7341 , n7342 , n7343 , n7344 , n7345 , n7346 , n7347 , n7348 , n7349 , n7350 , n7351 , n7352 , n7353 , n7354 , n7355 , n7356 , n7357 , n7358 , n7359 , n7360 , n7361 , n7362 , n7363 , n7364 , n7365 , n7366 , n7367 , n7368 , n7369 , n7370 , n7371 , n7372 , n7373 , n7374 , n7375 , n7376 , n7377 , n7378 , n7379 , n7380 , n7381 , n7382 , n7383 , n7384 , n7385 , n7386 , n7387 , n7388 , n7389 , n7390 , n7391 , n7392 , n7393 , n7394 , n7395 , n7396 , n7397 , n7398 , n7399 , n7400 , n7401 , n7402 , n7403 , n7404 , n7405 , n7406 , n7407 , n7408 , n7409 , n7410 , n7411 , n7412 , n7413 , n7414 , n7415 , n7416 , n7417 , n7418 , n7419 , n7420 , n7421 , n7422 , n7423 , n7424 , n7425 , n7426 , n7427 , n7428 , n7429 , n7430 , n7431 , n7432 , n7433 , n7434 , n7435 , n7436 , n7437 , n7438 , n7439 , n7440 , n7441 , n7442 , n7443 , n7444 , n7445 , n7446 , n7447 , n7448 , n7449 , n7450 , n7451 , n7452 , n7453 , n7454 , n7455 , n7456 , n7457 , n7458 , n7459 , n7460 , n7461 , n7462 , n7463 , n7464 , n7465 , n7466 , n7467 , n7468 , n7469 , n7470 , n7471 , n7472 , n7473 , n7474 , n7475 , n7476 , n7477 , n7478 , n7479 , n7480 , n7481 , n7482 , n7483 , n7484 , n7485 , n7486 , n7487 , n7488 , n7489 , n7490 , n7491 , n7492 , n7493 , n7494 , n7495 , n7496 , n7497 , n7498 , n7499 , n7500 , n7501 , n7502 , n7503 , n7504 , n7505 , n7506 , n7507 , n7508 , n7509 , n7510 , n7511 , n7512 , n7513 , n7514 , n7515 , n7516 , n7517 , n7518 , n7519 , n7520 , n7521 , n7522 , n7523 , n7524 , n7525 , n7526 , n7527 , n7528 , n7529 , n7530 , n7531 , n7532 , n7533 , n7534 , n7535 , n7536 , n7537 , n7538 , n7539 , n7540 , n7541 , n7542 , n7543 , n7544 , n7545 , n7546 , n7547 , n7548 , n7549 , n7550 , n7551 , n7552 , n7553 , n7554 , n7555 , n7556 , n7557 , n7558 , n7559 , n7560 , n7561 , n7562 , n7563 , n7564 , n7565 , n7566 , n7567 , n7568 , n7569 , n7570 , n7571 , n7572 , n7573 , n7574 , n7575 , n7576 , n7577 , n7578 , n7579 , n7580 , n7581 , n7582 , n7583 , n7584 , n7585 , n7586 , n7587 , n7588 , n7589 , n7590 , n7591 , n7592 , n7593 , n7594 , n7595 , n7596 , n7597 , n7598 , n7599 , n7600 , n7601 , n7602 , n7603 , n7604 , n7605 , n7606 , n7607 , n7608 , n7609 , n7610 , n7611 , n7612 , n7613 , n7614 , n7615 , n7616 , n7617 , n7618 , n7619 , n7620 , n7621 , n7622 , n7623 , n7624 , n7625 , n7626 , n7627 , n7628 , n7629 , n7630 , n7631 , n7632 , n7633 , n7634 , n7635 , n7636 , n7637 , n7638 , n7639 , n7640 , n7641 , n7642 , n7643 , n7644 , n7645 , n7646 , n7647 , n7648 , n7649 , n7650 , n7651 , n7652 , n7653 , n7654 , n7655 , n7656 , n7657 , n7658 , n7659 , n7660 , n7661 , n7662 , n7663 , n7664 , n7665 , n7666 , n7667 , n7668 , n7669 , n7670 , n7671 , n7672 , n7673 , n7674 , n7675 , n7676 , n7677 , n7678 , n7679 , n7680 , n7681 , n7682 , n7683 , n7684 , n7685 , n7686 , n7687 , n7688 , n7689 , n7690 , n7691 , n7692 , n7693 , n7694 , n7695 , n7696 , n7697 , n7698 , n7699 , n7700 , n7701 , n7702 , n7703 , n7704 , n7705 , n7706 , n7707 , n7708 , n7709 , n7710 , n7711 , n7712 , n7713 , n7714 , n7715 , n7716 , n7717 , n7718 , n7719 , n7720 , n7721 , n7722 , n7723 , n7724 , n7725 , n7726 , n7727 , n7728 , n7729 , n7730 , n7731 , n7732 , n7733 , n7734 , n7735 , n7736 , n7737 , n7738 , n7739 , n7740 , n7741 , n7742 , n7743 , n7744 , n7745 , n7746 , n7747 , n7748 , n7749 , n7750 , n7751 , n7752 , n7753 , n7754 , n7755 , n7756 , n7757 , n7758 , n7759 , n7760 , n7761 , n7762 , n7763 , n7764 , n7765 , n7766 , n7767 , n7768 , n7769 , n7770 , n7771 , n7772 , n7773 , n7774 , n7775 , n7776 , n7777 , n7778 , n7779 , n7780 , n7781 , n7782 , n7783 , n7784 , n7785 , n7786 , n7787 , n7788 , n7789 , n7790 , n7791 , n7792 , n7793 , n7794 , n7795 , n7796 , n7797 , n7798 , n7799 , n7800 , n7801 , n7802 , n7803 , n7804 , n7805 , n7806 , n7807 , n7808 , n7809 , n7810 , n7811 , n7812 , n7813 , n7814 , n7815 , n7816 , n7817 , n7818 , n7819 , n7820 , n7821 , n7822 , n7823 , n7824 , n7825 , n7826 , n7827 , n7828 , n7829 , n7830 , n7831 , n7832 , n7833 , n7834 , n7835 , n7836 , n7837 , n7838 , n7839 , n7840 , n7841 , n7842 , n7843 , n7844 , n7845 , n7846 , n7847 , n7848 , n7849 , n7850 , n7851 , n7852 , n7853 , n7854 , n7855 , n7856 , n7857 , n7858 , n7859 , n7860 , n7861 , n7862 , n7863 , n7864 , n7865 , n7866 , n7867 , n7868 , n7869 , n7870 , n7871 , n7872 , n7873 , n7874 , n7875 , n7876 , n7877 , n7878 , n7879 , n7880 , n7881 , n7882 , n7883 , n7884 , n7885 , n7886 , n7887 , n7888 , n7889 , n7890 , n7891 , n7892 , n7893 , n7894 , n7895 , n7896 , n7897 , n7898 , n7899 , n7900 , n7901 , n7902 , n7903 , n7904 , n7905 , n7906 , n7907 , n7908 , n7909 , n7910 , n7911 , n7912 , n7913 , n7914 , n7915 , n7916 , n7917 , n7918 , n7919 , n7920 , n7921 , n7922 , n7923 , n7924 , n7925 , n7926 , n7927 , n7928 , n7929 , n7930 , n7931 , n7932 , n7933 , n7934 , n7935 , n7936 , n7937 , n7938 , n7939 , n7940 , n7941 , n7942 , n7943 , n7944 , n7945 , n7946 , n7947 , n7948 , n7949 , n7950 , n7951 , n7952 , n7953 , n7954 , n7955 , n7956 , n7957 , n7958 , n7959 , n7960 , n7961 , n7962 , n7963 , n7964 , n7965 , n7966 , n7967 , n7968 , n7969 , n7970 , n7971 , n7972 , n7973 , n7974 , n7975 , n7976 , n7977 , n7978 , n7979 , n7980 , n7981 , n7982 , n7983 , n7984 , n7985 , n7986 , n7987 , n7988 , n7989 , n7990 , n7991 , n7992 , n7993 , n7994 , n7995 , n7996 , n7997 , n7998 , n7999 , n8000 , n8001 , n8002 , n8003 , n8004 , n8005 , n8006 , n8007 , n8008 , n8009 , n8010 , n8011 , n8012 , n8013 , n8014 , n8015 , n8016 , n8017 , n8018 , n8019 , n8020 , n8021 , n8022 , n8023 , n8024 , n8025 , n8026 , n8027 , n8028 , n8029 , n8030 , n8031 , n8032 , n8033 , n8034 , n8035 , n8036 , n8037 , n8038 , n8039 , n8040 , n8041 , n8042 , n8043 , n8044 , n8045 , n8046 , n8047 , n8048 , n8049 , n8050 , n8051 , n8052 , n8053 , n8054 , n8055 , n8056 , n8057 , n8058 , n8059 , n8060 , n8061 , n8062 , n8063 , n8064 , n8065 , n8066 , n8067 , n8068 , n8069 , n8070 , n8071 , n8072 , n8073 , n8074 , n8075 , n8076 , n8077 , n8078 , n8079 , n8080 , n8081 , n8082 , n8083 , n8084 , n8085 , n8086 , n8087 , n8088 , n8089 , n8090 , n8091 , n8092 , n8093 , n8094 , n8095 , n8096 , n8097 , n8098 , n8099 , n8100 , n8101 , n8102 , n8103 , n8104 , n8105 , n8106 , n8107 , n8108 , n8109 , n8110 , n8111 , n8112 , n8113 , n8114 , n8115 , n8116 , n8117 , n8118 , n8119 , n8120 , n8121 , n8122 , n8123 , n8124 , n8125 , n8126 , n8127 , n8128 , n8129 , n8130 , n8131 , n8132 , n8133 , n8134 , n8135 , n8136 , n8137 , n8138 , n8139 , n8140 , n8141 , n8142 , n8143 , n8144 , n8145 , n8146 , n8147 , n8148 , n8149 , n8150 , n8151 , n8152 , n8153 , n8154 , n8155 , n8156 , n8157 , n8158 , n8159 , n8160 , n8161 , n8162 , n8163 , n8164 , n8165 , n8166 , n8167 , n8168 , n8169 , n8170 , n8171 , n8172 , n8173 , n8174 , n8175 , n8176 , n8177 , n8178 , n8179 , n8180 , n8181 , n8182 , n8183 , n8184 , n8185 , n8186 , n8187 , n8188 , n8189 , n8190 , n8191 , n8192 , n8193 , n8194 , n8195 , n8196 , n8197 , n8198 , n8199 , n8200 , n8201 , n8202 , n8203 , n8204 , n8205 , n8206 , n8207 , n8208 , n8209 , n8210 , n8211 , n8212 , n8213 , n8214 , n8215 , n8216 , n8217 , n8218 , n8219 , n8220 , n8221 , n8222 , n8223 , n8224 , n8225 , n8226 , n8227 , n8228 , n8229 , n8230 , n8231 , n8232 , n8233 , n8234 , n8235 , n8236 , n8237 , n8238 , n8239 , n8240 , n8241 , n8242 , n8243 , n8244 , n8245 , n8246 , n8247 , n8248 , n8249 , n8250 , n8251 , n8252 , n8253 , n8254 , n8255 , n8256 , n8257 , n8258 , n8259 , n8260 , n8261 , n8262 , n8263 , n8264 , n8265 , n8266 , n8267 , n8268 , n8269 , n8270 , n8271 , n8272 , n8273 , n8274 , n8275 , n8276 , n8277 , n8278 , n8279 , n8280 , n8281 , n8282 , n8283 , n8284 , n8285 , n8286 , n8287 , n8288 , n8289 , n8290 , n8291 , n8292 , n8293 , n8294 , n8295 , n8296 , n8297 , n8298 , n8299 , n8300 , n8301 , n8302 , n8303 , n8304 , n8305 , n8306 , n8307 , n8308 , n8309 , n8310 , n8311 , n8312 , n8313 , n8314 , n8315 , n8316 , n8317 , n8318 , n8319 , n8320 , n8321 , n8322 , n8323 , n8324 , n8325 , n8326 , n8327 , n8328 , n8329 , n8330 , n8331 , n8332 , n8333 , n8334 , n8335 , n8336 , n8337 , n8338 , n8339 , n8340 , n8341 , n8342 , n8343 , n8344 , n8345 , n8346 , n8347 , n8348 , n8349 , n8350 , n8351 , n8352 , n8353 , n8354 , n8355 , n8356 , n8357 , n8358 , n8359 , n8360 , n8361 , n8362 , n8363 , n8364 , n8365 , n8366 , n8367 , n8368 , n8369 , n8370 , n8371 , n8372 , n8373 , n8374 , n8375 , n8376 , n8377 , n8378 , n8379 , n8380 , n8381 , n8382 , n8383 , n8384 , n8385 , n8386 , n8387 , n8388 , n8389 , n8390 , n8391 , n8392 , n8393 , n8394 , n8395 , n8396 , n8397 , n8398 , n8399 , n8400 , n8401 , n8402 , n8403 , n8404 , n8405 , n8406 , n8407 , n8408 , n8409 , n8410 , n8411 , n8412 , n8413 , n8414 , n8415 , n8416 , n8417 , n8418 , n8419 , n8420 , n8421 , n8422 , n8423 , n8424 , n8425 , n8426 , n8427 , n8428 , n8429 , n8430 , n8431 , n8432 , n8433 , n8434 , n8435 , n8436 , n8437 , n8438 , n8439 , n8440 , n8441 , n8442 , n8443 , n8444 , n8445 , n8446 , n8447 , n8448 , n8449 , n8450 , n8451 , n8452 , n8453 , n8454 , n8455 , n8456 , n8457 , n8458 , n8459 , n8460 , n8461 , n8462 , n8463 , n8464 , n8465 , n8466 , n8467 , n8468 , n8469 , n8470 , n8471 , n8472 , n8473 , n8474 , n8475 , n8476 , n8477 , n8478 , n8479 , n8480 , n8481 , n8482 , n8483 , n8484 , n8485 , n8486 , n8487 , n8488 , n8489 , n8490 , n8491 , n8492 , n8493 , n8494 , n8495 , n8496 , n8497 , n8498 , n8499 , n8500 , n8501 , n8502 , n8503 , n8504 , n8505 , n8506 , n8507 , n8508 , n8509 , n8510 , n8511 , n8512 , n8513 , n8514 , n8515 , n8516 , n8517 , n8518 , n8519 , n8520 , n8521 , n8522 , n8523 , n8524 , n8525 , n8526 , n8527 , n8528 , n8529 , n8530 , n8531 , n8532 , n8533 , n8534 , n8535 , n8536 , n8537 , n8538 , n8539 , n8540 , n8541 , n8542 , n8543 , n8544 , n8545 , n8546 , n8547 , n8548 , n8549 , n8550 , n8551 , n8552 , n8553 , n8554 , n8555 , n8556 , n8557 , n8558 , n8559 , n8560 , n8561 , n8562 , n8563 , n8564 , n8565 , n8566 , n8567 , n8568 , n8569 , n8570 , n8571 , n8572 , n8573 , n8574 , n8575 , n8576 , n8577 , n8578 , n8579 , n8580 , n8581 , n8582 , n8583 , n8584 , n8585 , n8586 , n8587 , n8588 , n8589 , n8590 , n8591 , n8592 , n8593 , n8594 , n8595 , n8596 , n8597 , n8598 , n8599 , n8600 , n8601 , n8602 , n8603 , n8604 , n8605 , n8606 , n8607 , n8608 , n8609 , n8610 , n8611 , n8612 , n8613 , n8614 , n8615 , n8616 , n8617 , n8618 , n8619 , n8620 , n8621 , n8622 , n8623 , n8624 , n8625 , n8626 , n8627 , n8628 , n8629 , n8630 , n8631 , n8632 , n8633 , n8634 , n8635 , n8636 , n8637 , n8638 , n8639 , n8640 , n8641 , n8642 , n8643 , n8644 , n8645 , n8646 , n8647 , n8648 , n8649 , n8650 , n8651 , n8652 , n8653 , n8654 , n8655 , n8656 , n8657 , n8658 , n8659 , n8660 , n8661 , n8662 , n8663 , n8664 , n8665 , n8666 , n8667 , n8668 , n8669 , n8670 , n8671 , n8672 , n8673 , n8674 , n8675 , n8676 , n8677 , n8678 , n8679 , n8680 , n8681 , n8682 , n8683 , n8684 , n8685 , n8686 , n8687 , n8688 , n8689 , n8690 , n8691 , n8692 , n8693 , n8694 , n8695 , n8696 , n8697 , n8698 , n8699 , n8700 , n8701 , n8702 , n8703 , n8704 , n8705 , n8706 , n8707 , n8708 , n8709 , n8710 , n8711 , n8712 , n8713 , n8714 , n8715 , n8716 , n8717 , n8718 , n8719 , n8720 , n8721 , n8722 , n8723 , n8724 , n8725 , n8726 , n8727 , n8728 , n8729 , n8730 , n8731 , n8732 , n8733 , n8734 , n8735 , n8736 , n8737 , n8738 , n8739 , n8740 , n8741 , n8742 , n8743 , n8744 , n8745 , n8746 , n8747 , n8748 , n8749 , n8750 , n8751 , n8752 , n8753 , n8754 , n8755 , n8756 , n8757 , n8758 , n8759 , n8760 , n8761 , n8762 , n8763 , n8764 , n8765 , n8766 , n8767 , n8768 , n8769 , n8770 , n8771 , n8772 , n8773 , n8774 , n8775 , n8776 , n8777 , n8778 , n8779 , n8780 , n8781 , n8782 , n8783 , n8784 , n8785 , n8786 , n8787 , n8788 , n8789 , n8790 , n8791 , n8792 , n8793 , n8794 , n8795 , n8796 , n8797 , n8798 , n8799 , n8800 , n8801 , n8802 , n8803 , n8804 , n8805 , n8806 , n8807 , n8808 , n8809 , n8810 , n8811 , n8812 , n8813 , n8814 , n8815 , n8816 , n8817 , n8818 , n8819 , n8820 , n8821 , n8822 , n8823 , n8824 , n8825 , n8826 , n8827 , n8828 , n8829 , n8830 , n8831 , n8832 , n8833 , n8834 , n8835 , n8836 , n8837 , n8838 , n8839 , n8840 , n8841 , n8842 , n8843 , n8844 , n8845 , n8846 , n8847 , n8848 , n8849 , n8850 , n8851 , n8852 , n8853 , n8854 , n8855 , n8856 , n8857 , n8858 , n8859 , n8860 , n8861 , n8862 , n8863 , n8864 , n8865 , n8866 , n8867 , n8868 , n8869 , n8870 , n8871 , n8872 , n8873 , n8874 , n8875 , n8876 , n8877 , n8878 , n8879 , n8880 , n8881 , n8882 , n8883 , n8884 , n8885 , n8886 , n8887 , n8888 , n8889 , n8890 , n8891 , n8892 , n8893 , n8894 , n8895 , n8896 , n8897 , n8898 , n8899 , n8900 , n8901 , n8902 , n8903 , n8904 , n8905 , n8906 , n8907 , n8908 , n8909 , n8910 , n8911 , n8912 , n8913 , n8914 , n8915 , n8916 , n8917 , n8918 , n8919 , n8920 , n8921 , n8922 , n8923 , n8924 , n8925 , n8926 , n8927 , n8928 , n8929 , n8930 , n8931 , n8932 , n8933 , n8934 , n8935 , n8936 , n8937 , n8938 , n8939 , n8940 , n8941 , n8942 , n8943 , n8944 , n8945 , n8946 , n8947 , n8948 , n8949 , n8950 , n8951 , n8952 , n8953 , n8954 , n8955 , n8956 , n8957 , n8958 , n8959 , n8960 , n8961 , n8962 , n8963 , n8964 , n8965 , n8966 , n8967 , n8968 , n8969 , n8970 , n8971 , n8972 , n8973 , n8974 , n8975 , n8976 , n8977 , n8978 , n8979 , n8980 , n8981 , n8982 , n8983 , n8984 , n8985 , n8986 , n8987 , n8988 , n8989 , n8990 , n8991 , n8992 , n8993 , n8994 , n8995 , n8996 , n8997 , n8998 , n8999 , n9000 , n9001 , n9002 , n9003 , n9004 , n9005 , n9006 , n9007 , n9008 , n9009 , n9010 , n9011 , n9012 , n9013 , n9014 , n9015 , n9016 , n9017 , n9018 , n9019 , n9020 , n9021 , n9022 , n9023 , n9024 , n9025 , n9026 , n9027 , n9028 , n9029 , n9030 , n9031 , n9032 , n9033 , n9034 , n9035 , n9036 , n9037 , n9038 , n9039 , n9040 , n9041 , n9042 , n9043 , n9044 , n9045 , n9046 , n9047 , n9048 , n9049 , n9050 , n9051 , n9052 , n9053 , n9054 , n9055 , n9056 , n9057 , n9058 , n9059 , n9060 , n9061 , n9062 , n9063 , n9064 , n9065 , n9066 , n9067 , n9068 , n9069 , n9070 , n9071 , n9072 , n9073 , n9074 , n9075 , n9076 , n9077 , n9078 , n9079 , n9080 , n9081 , n9082 , n9083 , n9084 , n9085 , n9086 , n9087 , n9088 , n9089 , n9090 , n9091 , n9092 , n9093 , n9094 , n9095 , n9096 , n9097 , n9098 , n9099 , n9100 , n9101 , n9102 , n9103 , n9104 , n9105 , n9106 , n9107 , n9108 , n9109 , n9110 , n9111 , n9112 , n9113 , n9114 , n9115 , n9116 , n9117 , n9118 , n9119 , n9120 , n9121 , n9122 , n9123 , n9124 , n9125 , n9126 , n9127 , n9128 , n9129 , n9130 , n9131 , n9132 , n9133 , n9134 , n9135 , n9136 , n9137 , n9138 , n9139 , n9140 , n9141 , n9142 , n9143 , n9144 , n9145 , n9146 , n9147 , n9148 , n9149 , n9150 , n9151 , n9152 , n9153 , n9154 , n9155 , n9156 , n9157 , n9158 , n9159 , n9160 , n9161 , n9162 , n9163 , n9164 , n9165 , n9166 , n9167 , n9168 , n9169 , n9170 , n9171 , n9172 , n9173 , n9174 , n9175 , n9176 , n9177 , n9178 , n9179 , n9180 , n9181 , n9182 , n9183 , n9184 , n9185 , n9186 , n9187 , n9188 , n9189 , n9190 , n9191 , n9192 , n9193 , n9194 , n9195 , n9196 , n9197 , n9198 , n9199 , n9200 , n9201 , n9202 , n9203 , n9204 , n9205 , n9206 , n9207 , n9208 , n9209 , n9210 , n9211 , n9212 , n9213 , n9214 , n9215 , n9216 , n9217 , n9218 , n9219 , n9220 , n9221 , n9222 , n9223 , n9224 , n9225 , n9226 , n9227 , n9228 , n9229 , n9230 , n9231 , n9232 , n9233 , n9234 , n9235 , n9236 , n9237 , n9238 , n9239 , n9240 , n9241 , n9242 , n9243 , n9244 , n9245 , n9246 , n9247 , n9248 , n9249 , n9250 , n9251 , n9252 , n9253 , n9254 , n9255 , n9256 , n9257 , n9258 , n9259 , n9260 , n9261 , n9262 , n9263 , n9264 , n9265 , n9266 , n9267 , n9268 , n9269 , n9270 , n9271 , n9272 , n9273 , n9274 , n9275 , n9276 , n9277 , n9278 , n9279 , n9280 , n9281 , n9282 , n9283 , n9284 , n9285 , n9286 , n9287 , n9288 , n9289 , n9290 , n9291 , n9292 , n9293 , n9294 , n9295 , n9296 , n9297 , n9298 , n9299 , n9300 , n9301 , n9302 , n9303 , n9304 , n9305 , n9306 , n9307 , n9308 , n9309 , n9310 , n9311 , n9312 , n9313 , n9314 , n9315 , n9316 , n9317 , n9318 , n9319 , n9320 , n9321 , n9322 , n9323 , n9324 , n9325 , n9326 , n9327 , n9328 , n9329 , n9330 , n9331 , n9332 , n9333 , n9334 , n9335 , n9336 , n9337 , n9338 , n9339 , n9340 , n9341 , n9342 , n9343 , n9344 , n9345 , n9346 , n9347 , n9348 , n9349 , n9350 , n9351 , n9352 , n9353 , n9354 , n9355 , n9356 , n9357 , n9358 , n9359 , n9360 , n9361 , n9362 , n9363 , n9364 , n9365 , n9366 , n9367 , n9368 , n9369 , n9370 , n9371 , n9372 , n9373 , n9374 , n9375 , n9376 , n9377 , n9378 , n9379 , n9380 , n9381 , n9382 , n9383 , n9384 , n9385 , n9386 , n9387 , n9388 , n9389 , n9390 , n9391 , n9392 , n9393 , n9394 , n9395 , n9396 , n9397 , n9398 , n9399 , n9400 , n9401 , n9402 , n9403 , n9404 , n9405 , n9406 , n9407 , n9408 , n9409 , n9410 , n9411 , n9412 , n9413 , n9414 , n9415 , n9416 , n9417 , n9418 , n9419 , n9420 , n9421 , n9422 , n9423 , n9424 , n9425 , n9426 , n9427 , n9428 , n9429 , n9430 , n9431 , n9432 , n9433 , n9434 , n9435 , n9436 , n9437 , n9438 , n9439 , n9440 , n9441 , n9442 , n9443 , n9444 , n9445 , n9446 , n9447 , n9448 , n9449 , n9450 , n9451 , n9452 , n9453 , n9454 , n9455 , n9456 , n9457 , n9458 , n9459 , n9460 , n9461 , n9462 , n9463 , n9464 , n9465 , n9466 , n9467 , n9468 , n9469 , n9470 , n9471 , n9472 , n9473 , n9474 , n9475 , n9476 , n9477 , n9478 , n9479 , n9480 , n9481 , n9482 , n9483 , n9484 , n9485 , n9486 , n9487 , n9488 , n9489 , n9490 , n9491 , n9492 , n9493 , n9494 , n9495 , n9496 , n9497 , n9498 , n9499 , n9500 , n9501 , n9502 , n9503 , n9504 , n9505 , n9506 , n9507 , n9508 , n9509 , n9510 , n9511 , n9512 , n9513 , n9514 , n9515 , n9516 , n9517 , n9518 , n9519 , n9520 , n9521 , n9522 , n9523 , n9524 , n9525 , n9526 , n9527 , n9528 , n9529 , n9530 , n9531 , n9532 , n9533 , n9534 , n9535 , n9536 , n9537 , n9538 , n9539 , n9540 , n9541 , n9542 , n9543 , n9544 , n9545 , n9546 , n9547 , n9548 , n9549 , n9550 , n9551 , n9552 , n9553 , n9554 , n9555 , n9556 , n9557 , n9558 , n9559 , n9560 , n9561 , n9562 , n9563 , n9564 , n9565 , n9566 , n9567 , n9568 , n9569 , n9570 , n9571 , n9572 , n9573 , n9574 , n9575 , n9576 , n9577 , n9578 , n9579 , n9580 , n9581 , n9582 , n9583 , n9584 , n9585 , n9586 , n9587 , n9588 , n9589 , n9590 , n9591 , n9592 , n9593 , n9594 , n9595 , n9596 , n9597 , n9598 , n9599 , n9600 , n9601 , n9602 , n9603 , n9604 , n9605 , n9606 , n9607 , n9608 , n9609 , n9610 , n9611 , n9612 , n9613 , n9614 , n9615 , n9616 , n9617 , n9618 , n9619 , n9620 , n9621 , n9622 , n9623 , n9624 , n9625 , n9626 , n9627 , n9628 , n9629 , n9630 , n9631 , n9632 , n9633 , n9634 , n9635 , n9636 , n9637 , n9638 , n9639 , n9640 , n9641 , n9642 , n9643 , n9644 , n9645 , n9646 , n9647 , n9648 , n9649 , n9650 , n9651 , n9652 , n9653 , n9654 , n9655 , n9656 , n9657 , n9658 , n9659 , n9660 , n9661 , n9662 , n9663 , n9664 , n9665 , n9666 , n9667 , n9668 , n9669 , n9670 , n9671 , n9672 , n9673 , n9674 , n9675 , n9676 , n9677 , n9678 , n9679 , n9680 , n9681 , n9682 , n9683 , n9684 , n9685 , n9686 , n9687 , n9688 , n9689 , n9690 , n9691 , n9692 , n9693 , n9694 , n9695 , n9696 , n9697 , n9698 , n9699 , n9700 , n9701 , n9702 , n9703 , n9704 , n9705 , n9706 , n9707 , n9708 , n9709 , n9710 , n9711 , n9712 , n9713 , n9714 , n9715 , n9716 , n9717 , n9718 , n9719 , n9720 , n9721 , n9722 , n9723 , n9724 , n9725 , n9726 , n9727 , n9728 , n9729 , n9730 , n9731 , n9732 , n9733 , n9734 , n9735 , n9736 , n9737 , n9738 , n9739 , n9740 , n9741 , n9742 , n9743 , n9744 , n9745 , n9746 , n9747 , n9748 , n9749 , n9750 , n9751 , n9752 , n9753 , n9754 , n9755 , n9756 , n9757 , n9758 , n9759 , n9760 , n9761 , n9762 , n9763 , n9764 , n9765 , n9766 , n9767 , n9768 , n9769 , n9770 , n9771 , n9772 , n9773 , n9774 , n9775 , n9776 , n9777 , n9778 , n9779 , n9780 , n9781 , n9782 , n9783 , n9784 , n9785 , n9786 , n9787 , n9788 , n9789 , n9790 , n9791 , n9792 , n9793 , n9794 , n9795 , n9796 , n9797 , n9798 , n9799 , n9800 , n9801 , n9802 , n9803 , n9804 , n9805 , n9806 , n9807 , n9808 , n9809 , n9810 , n9811 , n9812 , n9813 , n9814 , n9815 , n9816 , n9817 , n9818 , n9819 , n9820 , n9821 , n9822 , n9823 , n9824 , n9825 , n9826 , n9827 , n9828 , n9829 , n9830 , n9831 , n9832 , n9833 , n9834 , n9835 , n9836 , n9837 , n9838 , n9839 , n9840 , n9841 , n9842 , n9843 , n9844 , n9845 , n9846 , n9847 , n9848 , n9849 , n9850 , n9851 , n9852 , n9853 , n9854 , n9855 , n9856 , n9857 , n9858 , n9859 , n9860 , n9861 , n9862 , n9863 , n9864 , n9865 , n9866 , n9867 , n9868 , n9869 , n9870 , n9871 , n9872 , n9873 , n9874 , n9875 , n9876 , n9877 , n9878 , n9879 , n9880 , n9881 , n9882 , n9883 , n9884 , n9885 , n9886 , n9887 , n9888 , n9889 , n9890 , n9891 , n9892 , n9893 , n9894 , n9895 , n9896 , n9897 , n9898 , n9899 , n9900 , n9901 , n9902 , n9903 , n9904 , n9905 , n9906 , n9907 , n9908 , n9909 , n9910 , n9911 , n9912 , n9913 , n9914 , n9915 , n9916 , n9917 , n9918 , n9919 , n9920 , n9921 , n9922 , n9923 , n9924 , n9925 , n9926 , n9927 , n9928 , n9929 , n9930 , n9931 , n9932 , n9933 , n9934 , n9935 , n9936 , n9937 , n9938 , n9939 , n9940 , n9941 , n9942 , n9943 , n9944 , n9945 , n9946 , n9947 , n9948 , n9949 , n9950 , n9951 , n9952 , n9953 , n9954 , n9955 , n9956 , n9957 , n9958 , n9959 , n9960 , n9961 , n9962 , n9963 , n9964 , n9965 , n9966 , n9967 , n9968 , n9969 , n9970 , n9971 , n9972 , n9973 , n9974 , n9975 , n9976 , n9977 , n9978 , n9979 , n9980 , n9981 , n9982 , n9983 , n9984 , n9985 , n9986 , n9987 , n9988 , n9989 , n9990 , n9991 , n9992 , n9993 , n9994 , n9995 , n9996 , n9997 , n9998 , n9999 , n10000 , n10001 , n10002 , n10003 , n10004 , n10005 , n10006 , n10007 , n10008 , n10009 , n10010 , n10011 , n10012 , n10013 , n10014 , n10015 , n10016 , n10017 , n10018 , n10019 , n10020 , n10021 , n10022 , n10023 , n10024 , n10025 , n10026 , n10027 , n10028 , n10029 , n10030 , n10031 , n10032 , n10033 , n10034 , n10035 , n10036 , n10037 , n10038 , n10039 , n10040 , n10041 , n10042 , n10043 , n10044 , n10045 , n10046 , n10047 , n10048 , n10049 , n10050 , n10051 , n10052 , n10053 , n10054 , n10055 , n10056 , n10057 , n10058 , n10059 , n10060 , n10061 , n10062 , n10063 , n10064 , n10065 , n10066 , n10067 , n10068 , n10069 , n10070 , n10071 , n10072 , n10073 , n10074 , n10075 , n10076 , n10077 , n10078 , n10079 , n10080 , n10081 , n10082 , n10083 , n10084 , n10085 , n10086 , n10087 , n10088 , n10089 , n10090 , n10091 , n10092 , n10093 , n10094 , n10095 , n10096 , n10097 , n10098 , n10099 , n10100 , n10101 , n10102 , n10103 , n10104 , n10105 , n10106 , n10107 , n10108 , n10109 , n10110 , n10111 , n10112 , n10113 , n10114 , n10115 , n10116 , n10117 , n10118 , n10119 , n10120 , n10121 , n10122 , n10123 , n10124 , n10125 , n10126 , n10127 , n10128 , n10129 , n10130 , n10131 , n10132 , n10133 , n10134 , n10135 , n10136 , n10137 , n10138 , n10139 , n10140 , n10141 , n10142 , n10143 , n10144 , n10145 , n10146 , n10147 , n10148 , n10149 , n10150 , n10151 , n10152 , n10153 , n10154 , n10155 , n10156 , n10157 , n10158 , n10159 , n10160 , n10161 , n10162 , n10163 , n10164 , n10165 , n10166 , n10167 , n10168 , n10169 , n10170 , n10171 , n10172 , n10173 , n10174 , n10175 , n10176 , n10177 , n10178 , n10179 , n10180 , n10181 , n10182 , n10183 , n10184 , n10185 , n10186 , n10187 , n10188 , n10189 , n10190 , n10191 , n10192 , n10193 , n10194 , n10195 , n10196 , n10197 , n10198 , n10199 , n10200 , n10201 , n10202 , n10203 , n10204 , n10205 , n10206 , n10207 , n10208 , n10209 , n10210 , n10211 , n10212 , n10213 , n10214 , n10215 , n10216 , n10217 , n10218 , n10219 , n10220 , n10221 , n10222 , n10223 , n10224 , n10225 , n10226 , n10227 , n10228 , n10229 , n10230 , n10231 , n10232 , n10233 , n10234 , n10235 , n10236 , n10237 , n10238 , n10239 , n10240 , n10241 , n10242 , n10243 , n10244 , n10245 , n10246 , n10247 , n10248 , n10249 , n10250 , n10251 , n10252 , n10253 , n10254 , n10255 , n10256 , n10257 , n10258 , n10259 , n10260 , n10261 , n10262 , n10263 , n10264 , n10265 , n10266 , n10267 , n10268 , n10269 , n10270 , n10271 , n10272 , n10273 , n10274 , n10275 , n10276 , n10277 , n10278 , n10279 , n10280 , n10281 , n10282 , n10283 , n10284 , n10285 , n10286 , n10287 , n10288 , n10289 , n10290 , n10291 , n10292 , n10293 , n10294 , n10295 , n10296 , n10297 , n10298 , n10299 , n10300 , n10301 , n10302 , n10303 , n10304 , n10305 , n10306 , n10307 , n10308 , n10309 , n10310 , n10311 , n10312 , n10313 , n10314 , n10315 , n10316 , n10317 , n10318 , n10319 , n10320 , n10321 , n10322 , n10323 , n10324 , n10325 , n10326 , n10327 , n10328 , n10329 , n10330 , n10331 , n10332 , n10333 , n10334 , n10335 , n10336 , n10337 , n10338 , n10339 , n10340 , n10341 , n10342 , n10343 , n10344 , n10345 , n10346 , n10347 , n10348 , n10349 , n10350 , n10351 , n10352 , n10353 , n10354 , n10355 , n10356 , n10357 , n10358 , n10359 , n10360 , n10361 , n10362 , n10363 , n10364 , n10365 , n10366 , n10367 , n10368 , n10369 , n10370 , n10371 , n10372 , n10373 , n10374 , n10375 , n10376 , n10377 , n10378 , n10379 , n10380 , n10381 , n10382 , n10383 , n10384 , n10385 , n10386 , n10387 , n10388 , n10389 , n10390 , n10391 , n10392 , n10393 , n10394 , n10395 , n10396 , n10397 , n10398 , n10399 , n10400 , n10401 , n10402 , n10403 , n10404 , n10405 , n10406 , n10407 , n10408 , n10409 , n10410 , n10411 , n10412 , n10413 , n10414 , n10415 , n10416 , n10417 , n10418 , n10419 , n10420 , n10421 , n10422 , n10423 , n10424 , n10425 , n10426 , n10427 , n10428 , n10429 , n10430 , n10431 , n10432 , n10433 , n10434 , n10435 , n10436 , n10437 , n10438 , n10439 , n10440 , n10441 , n10442 , n10443 , n10444 , n10445 , n10446 , n10447 , n10448 , n10449 , n10450 , n10451 , n10452 , n10453 , n10454 , n10455 , n10456 , n10457 , n10458 , n10459 , n10460 , n10461 , n10462 , n10463 , n10464 , n10465 , n10466 , n10467 , n10468 , n10469 , n10470 , n10471 , n10472 , n10473 , n10474 , n10475 , n10476 , n10477 , n10478 , n10479 , n10480 , n10481 , n10482 , n10483 , n10484 , n10485 , n10486 , n10487 , n10488 , n10489 , n10490 , n10491 , n10492 , n10493 , n10494 , n10495 , n10496 , n10497 , n10498 , n10499 , n10500 , n10501 , n10502 , n10503 , n10504 , n10505 , n10506 , n10507 , n10508 , n10509 , n10510 , n10511 , n10512 , n10513 , n10514 , n10515 , n10516 , n10517 , n10518 , n10519 , n10520 , n10521 , n10522 , n10523 , n10524 , n10525 , n10526 , n10527 , n10528 , n10529 , n10530 , n10531 , n10532 , n10533 , n10534 , n10535 , n10536 , n10537 , n10538 , n10539 , n10540 , n10541 , n10542 , n10543 , n10544 , n10545 , n10546 , n10547 , n10548 , n10549 , n10550 , n10551 , n10552 , n10553 , n10554 , n10555 , n10556 , n10557 , n10558 , n10559 , n10560 , n10561 , n10562 , n10563 , n10564 , n10565 , n10566 , n10567 , n10568 , n10569 , n10570 , n10571 , n10572 , n10573 , n10574 , n10575 , n10576 , n10577 , n10578 , n10579 , n10580 , n10581 , n10582 , n10583 , n10584 , n10585 , n10586 , n10587 , n10588 , n10589 , n10590 , n10591 , n10592 , n10593 , n10594 , n10595 , n10596 , n10597 , n10598 , n10599 , n10600 , n10601 , n10602 , n10603 , n10604 , n10605 , n10606 , n10607 , n10608 , n10609 , n10610 , n10611 , n10612 , n10613 , n10614 , n10615 , n10616 , n10617 , n10618 , n10619 , n10620 , n10621 , n10622 , n10623 , n10624 , n10625 , n10626 , n10627 , n10628 , n10629 , n10630 , n10631 , n10632 , n10633 , n10634 , n10635 , n10636 , n10637 , n10638 , n10639 , n10640 , n10641 , n10642 , n10643 , n10644 , n10645 , n10646 , n10647 , n10648 , n10649 , n10650 , n10651 , n10652 , n10653 , n10654 , n10655 , n10656 , n10657 , n10658 , n10659 , n10660 , n10661 , n10662 , n10663 , n10664 , n10665 , n10666 , n10667 , n10668 , n10669 , n10670 , n10671 , n10672 , n10673 , n10674 , n10675 , n10676 , n10677 , n10678 , n10679 , n10680 , n10681 , n10682 , n10683 , n10684 , n10685 , n10686 , n10687 , n10688 , n10689 , n10690 , n10691 , n10692 , n10693 , n10694 , n10695 , n10696 , n10697 , n10698 , n10699 , n10700 , n10701 , n10702 , n10703 , n10704 , n10705 , n10706 , n10707 , n10708 , n10709 , n10710 , n10711 , n10712 , n10713 , n10714 , n10715 , n10716 , n10717 , n10718 , n10719 , n10720 , n10721 , n10722 , n10723 , n10724 , n10725 , n10726 , n10727 , n10728 , n10729 , n10730 , n10731 , n10732 , n10733 , n10734 , n10735 , n10736 , n10737 , n10738 , n10739 , n10740 , n10741 , n10742 , n10743 , n10744 , n10745 , n10746 , n10747 , n10748 , n10749 , n10750 , n10751 , n10752 , n10753 , n10754 , n10755 , n10756 , n10757 , n10758 , n10759 , n10760 , n10761 , n10762 , n10763 , n10764 , n10765 , n10766 , n10767 , n10768 , n10769 , n10770 , n10771 , n10772 , n10773 , n10774 , n10775 , n10776 , n10777 , n10778 , n10779 , n10780 , n10781 , n10782 , n10783 , n10784 , n10785 , n10786 , n10787 , n10788 , n10789 , n10790 , n10791 , n10792 , n10793 , n10794 , n10795 , n10796 , n10797 , n10798 , n10799 , n10800 , n10801 , n10802 , n10803 , n10804 , n10805 , n10806 , n10807 , n10808 , n10809 , n10810 , n10811 , n10812 , n10813 , n10814 , n10815 , n10816 , n10817 , n10818 , n10819 , n10820 , n10821 , n10822 , n10823 , n10824 , n10825 , n10826 , n10827 , n10828 , n10829 , n10830 , n10831 , n10832 , n10833 , n10834 , n10835 , n10836 , n10837 , n10838 , n10839 , n10840 , n10841 , n10842 , n10843 , n10844 , n10845 , n10846 , n10847 , n10848 , n10849 , n10850 , n10851 , n10852 , n10853 , n10854 , n10855 , n10856 , n10857 , n10858 , n10859 , n10860 , n10861 , n10862 , n10863 , n10864 , n10865 , n10866 , n10867 , n10868 , n10869 , n10870 , n10871 , n10872 , n10873 , n10874 , n10875 , n10876 , n10877 , n10878 , n10879 , n10880 , n10881 , n10882 , n10883 , n10884 , n10885 , n10886 , n10887 , n10888 , n10889 , n10890 , n10891 , n10892 , n10893 , n10894 , n10895 , n10896 , n10897 , n10898 , n10899 , n10900 , n10901 , n10902 , n10903 , n10904 , n10905 , n10906 , n10907 , n10908 , n10909 , n10910 , n10911 , n10912 , n10913 , n10914 , n10915 , n10916 , n10917 , n10918 , n10919 , n10920 , n10921 , n10922 , n10923 , n10924 , n10925 , n10926 , n10927 , n10928 , n10929 , n10930 , n10931 , n10932 , n10933 , n10934 , n10935 , n10936 , n10937 , n10938 , n10939 , n10940 , n10941 , n10942 , n10943 , n10944 , n10945 , n10946 , n10947 , n10948 , n10949 , n10950 , n10951 , n10952 , n10953 , n10954 , n10955 , n10956 , n10957 , n10958 , n10959 , n10960 , n10961 , n10962 , n10963 , n10964 , n10965 , n10966 , n10967 , n10968 , n10969 , n10970 , n10971 , n10972 , n10973 , n10974 , n10975 , n10976 , n10977 , n10978 , n10979 , n10980 , n10981 , n10982 , n10983 , n10984 , n10985 , n10986 , n10987 , n10988 , n10989 , n10990 , n10991 , n10992 , n10993 , n10994 , n10995 , n10996 , n10997 , n10998 , n10999 , n11000 , n11001 , n11002 , n11003 , n11004 , n11005 , n11006 , n11007 , n11008 , n11009 , n11010 , n11011 , n11012 , n11013 , n11014 , n11015 , n11016 , n11017 , n11018 , n11019 , n11020 , n11021 , n11022 , n11023 , n11024 , n11025 , n11026 , n11027 , n11028 , n11029 , n11030 , n11031 , n11032 , n11033 , n11034 , n11035 , n11036 , n11037 , n11038 , n11039 , n11040 , n11041 , n11042 , n11043 , n11044 , n11045 , n11046 , n11047 , n11048 , n11049 , n11050 , n11051 , n11052 , n11053 , n11054 , n11055 , n11056 , n11057 , n11058 , n11059 , n11060 , n11061 , n11062 , n11063 , n11064 , n11065 , n11066 , n11067 , n11068 , n11069 , n11070 , n11071 , n11072 , n11073 , n11074 , n11075 , n11076 , n11077 , n11078 , n11079 , n11080 , n11081 , n11082 , n11083 , n11084 , n11085 , n11086 , n11087 , n11088 , n11089 , n11090 , n11091 , n11092 , n11093 , n11094 , n11095 , n11096 , n11097 , n11098 , n11099 , n11100 , n11101 , n11102 , n11103 , n11104 , n11105 , n11106 , n11107 , n11108 , n11109 , n11110 , n11111 , n11112 , n11113 , n11114 , n11115 , n11116 , n11117 , n11118 , n11119 , n11120 , n11121 , n11122 , n11123 , n11124 , n11125 , n11126 , n11127 , n11128 , n11129 , n11130 , n11131 , n11132 , n11133 , n11134 , n11135 , n11136 , n11137 , n11138 , n11139 , n11140 , n11141 , n11142 , n11143 , n11144 , n11145 , n11146 , n11147 , n11148 , n11149 , n11150 , n11151 , n11152 , n11153 , n11154 , n11155 , n11156 , n11157 , n11158 , n11159 , n11160 , n11161 , n11162 , n11163 , n11164 , n11165 , n11166 , n11167 , n11168 , n11169 , n11170 , n11171 , n11172 , n11173 , n11174 , n11175 , n11176 , n11177 , n11178 , n11179 , n11180 , n11181 , n11182 , n11183 , n11184 , n11185 , n11186 , n11187 , n11188 , n11189 , n11190 , n11191 , n11192 , n11193 , n11194 , n11195 , n11196 , n11197 , n11198 , n11199 , n11200 , n11201 , n11202 , n11203 , n11204 , n11205 , n11206 , n11207 , n11208 , n11209 , n11210 , n11211 , n11212 , n11213 , n11214 , n11215 , n11216 , n11217 , n11218 , n11219 , n11220 , n11221 , n11222 , n11223 , n11224 , n11225 , n11226 , n11227 , n11228 , n11229 , n11230 , n11231 , n11232 , n11233 , n11234 , n11235 , n11236 , n11237 , n11238 , n11239 , n11240 , n11241 , n11242 , n11243 , n11244 , n11245 , n11246 , n11247 , n11248 , n11249 , n11250 , n11251 , n11252 , n11253 , n11254 , n11255 , n11256 , n11257 , n11258 , n11259 , n11260 , n11261 , n11262 , n11263 , n11264 , n11265 , n11266 , n11267 , n11268 , n11269 , n11270 , n11271 , n11272 , n11273 , n11274 , n11275 , n11276 , n11277 , n11278 , n11279 , n11280 , n11281 , n11282 , n11283 , n11284 , n11285 , n11286 , n11287 , n11288 , n11289 , n11290 , n11291 , n11292 , n11293 , n11294 , n11295 , n11296 , n11297 , n11298 , n11299 , n11300 , n11301 , n11302 , n11303 , n11304 , n11305 , n11306 , n11307 , n11308 , n11309 , n11310 , n11311 , n11312 , n11313 , n11314 , n11315 , n11316 , n11317 , n11318 , n11319 , n11320 , n11321 , n11322 , n11323 , n11324 , n11325 , n11326 , n11327 , n11328 , n11329 , n11330 , n11331 , n11332 , n11333 , n11334 , n11335 , n11336 , n11337 , n11338 , n11339 , n11340 , n11341 , n11342 , n11343 , n11344 , n11345 , n11346 , n11347 , n11348 , n11349 , n11350 , n11351 , n11352 , n11353 , n11354 , n11355 , n11356 , n11357 , n11358 , n11359 , n11360 , n11361 , n11362 , n11363 , n11364 , n11365 , n11366 , n11367 , n11368 , n11369 , n11370 , n11371 , n11372 , n11373 , n11374 , n11375 , n11376 , n11377 , n11378 , n11379 , n11380 , n11381 , n11382 , n11383 , n11384 , n11385 , n11386 , n11387 , n11388 , n11389 , n11390 , n11391 , n11392 , n11393 , n11394 , n11395 , n11396 , n11397 , n11398 , n11399 , n11400 , n11401 , n11402 , n11403 , n11404 , n11405 , n11406 , n11407 , n11408 , n11409 , n11410 , n11411 , n11412 , n11413 , n11414 , n11415 , n11416 , n11417 , n11418 , n11419 , n11420 , n11421 , n11422 , n11423 , n11424 , n11425 , n11426 , n11427 , n11428 , n11429 , n11430 , n11431 , n11432 , n11433 , n11434 , n11435 , n11436 , n11437 , n11438 , n11439 , n11440 , n11441 , n11442 , n11443 , n11444 , n11445 , n11446 , n11447 , n11448 , n11449 , n11450 , n11451 , n11452 , n11453 , n11454 , n11455 , n11456 , n11457 , n11458 , n11459 , n11460 , n11461 , n11462 , n11463 , n11464 , n11465 , n11466 , n11467 , n11468 , n11469 , n11470 , n11471 , n11472 , n11473 , n11474 , n11475 , n11476 , n11477 , n11478 , n11479 , n11480 , n11481 , n11482 , n11483 , n11484 , n11485 , n11486 , n11487 , n11488 , n11489 , n11490 , n11491 , n11492 , n11493 , n11494 , n11495 , n11496 , n11497 , n11498 , n11499 , n11500 , n11501 , n11502 , n11503 , n11504 , n11505 , n11506 , n11507 , n11508 , n11509 , n11510 , n11511 , n11512 , n11513 , n11514 , n11515 , n11516 , n11517 , n11518 , n11519 , n11520 , n11521 , n11522 , n11523 , n11524 , n11525 , n11526 , n11527 , n11528 , n11529 , n11530 , n11531 , n11532 , n11533 , n11534 , n11535 , n11536 , n11537 , n11538 , n11539 , n11540 , n11541 , n11542 , n11543 , n11544 , n11545 , n11546 , n11547 , n11548 , n11549 , n11550 , n11551 , n11552 , n11553 , n11554 , n11555 , n11556 , n11557 , n11558 , n11559 , n11560 , n11561 , n11562 , n11563 , n11564 , n11565 , n11566 , n11567 , n11568 , n11569 , n11570 , n11571 , n11572 , n11573 , n11574 , n11575 , n11576 , n11577 , n11578 , n11579 , n11580 , n11581 , n11582 , n11583 , n11584 , n11585 , n11586 , n11587 , n11588 , n11589 , n11590 , n11591 , n11592 , n11593 , n11594 , n11595 , n11596 , n11597 , n11598 , n11599 , n11600 , n11601 , n11602 , n11603 , n11604 , n11605 , n11606 , n11607 , n11608 , n11609 , n11610 , n11611 , n11612 , n11613 , n11614 , n11615 , n11616 , n11617 , n11618 , n11619 , n11620 , n11621 , n11622 , n11623 , n11624 , n11625 , n11626 , n11627 , n11628 , n11629 , n11630 , n11631 , n11632 , n11633 , n11634 , n11635 , n11636 , n11637 , n11638 , n11639 , n11640 , n11641 , n11642 , n11643 , n11644 , n11645 , n11646 , n11647 , n11648 , n11649 , n11650 , n11651 , n11652 , n11653 , n11654 , n11655 , n11656 , n11657 , n11658 , n11659 , n11660 , n11661 , n11662 , n11663 , n11664 , n11665 , n11666 , n11667 , n11668 , n11669 , n11670 , n11671 , n11672 , n11673 , n11674 , n11675 , n11676 , n11677 , n11678 , n11679 , n11680 , n11681 , n11682 , n11683 , n11684 , n11685 , n11686 , n11687 , n11688 , n11689 , n11690 , n11691 , n11692 , n11693 , n11694 , n11695 , n11696 , n11697 , n11698 , n11699 , n11700 , n11701 , n11702 , n11703 , n11704 , n11705 , n11706 , n11707 , n11708 , n11709 , n11710 , n11711 , n11712 , n11713 , n11714 , n11715 , n11716 , n11717 , n11718 , n11719 , n11720 , n11721 , n11722 , n11723 , n11724 , n11725 , n11726 , n11727 , n11728 , n11729 , n11730 , n11731 , n11732 , n11733 , n11734 , n11735 , n11736 , n11737 , n11738 , n11739 , n11740 , n11741 , n11742 , n11743 , n11744 , n11745 , n11746 , n11747 , n11748 , n11749 , n11750 , n11751 , n11752 , n11753 , n11754 , n11755 , n11756 , n11757 , n11758 , n11759 , n11760 , n11761 , n11762 , n11763 , n11764 , n11765 , n11766 , n11767 , n11768 , n11769 , n11770 , n11771 , n11772 , n11773 , n11774 , n11775 , n11776 , n11777 , n11778 , n11779 , n11780 , n11781 , n11782 , n11783 , n11784 , n11785 , n11786 , n11787 , n11788 , n11789 , n11790 , n11791 , n11792 , n11793 , n11794 , n11795 , n11796 , n11797 , n11798 , n11799 , n11800 , n11801 , n11802 , n11803 , n11804 , n11805 , n11806 , n11807 , n11808 , n11809 , n11810 , n11811 , n11812 , n11813 , n11814 , n11815 , n11816 , n11817 , n11818 , n11819 , n11820 , n11821 , n11822 , n11823 , n11824 , n11825 , n11826 , n11827 , n11828 , n11829 , n11830 , n11831 , n11832 , n11833 , n11834 , n11835 , n11836 , n11837 , n11838 , n11839 , n11840 , n11841 , n11842 , n11843 , n11844 , n11845 , n11846 , n11847 , n11848 , n11849 , n11850 , n11851 , n11852 , n11853 , n11854 , n11855 , n11856 , n11857 , n11858 , n11859 , n11860 , n11861 , n11862 , n11863 , n11864 , n11865 , n11866 , n11867 , n11868 , n11869 , n11870 , n11871 , n11872 , n11873 , n11874 , n11875 , n11876 , n11877 , n11878 , n11879 , n11880 , n11881 , n11882 , n11883 , n11884 , n11885 , n11886 , n11887 , n11888 , n11889 , n11890 , n11891 , n11892 , n11893 , n11894 , n11895 , n11896 , n11897 , n11898 , n11899 , n11900 , n11901 , n11902 , n11903 , n11904 , n11905 , n11906 , n11907 , n11908 , n11909 , n11910 , n11911 , n11912 , n11913 , n11914 , n11915 , n11916 , n11917 , n11918 , n11919 , n11920 , n11921 , n11922 , n11923 , n11924 , n11925 , n11926 , n11927 , n11928 , n11929 , n11930 , n11931 , n11932 , n11933 , n11934 , n11935 , n11936 , n11937 , n11938 , n11939 , n11940 , n11941 , n11942 , n11943 , n11944 , n11945 , n11946 , n11947 , n11948 , n11949 , n11950 , n11951 , n11952 , n11953 , n11954 , n11955 , n11956 , n11957 , n11958 , n11959 , n11960 , n11961 , n11962 , n11963 , n11964 , n11965 , n11966 , n11967 , n11968 , n11969 , n11970 , n11971 , n11972 , n11973 , n11974 , n11975 , n11976 , n11977 , n11978 , n11979 , n11980 , n11981 , n11982 , n11983 , n11984 , n11985 , n11986 , n11987 , n11988 , n11989 , n11990 , n11991 , n11992 , n11993 , n11994 , n11995 , n11996 , n11997 , n11998 , n11999 , n12000 , n12001 , n12002 , n12003 , n12004 , n12005 , n12006 , n12007 , n12008 , n12009 , n12010 , n12011 , n12012 , n12013 , n12014 , n12015 , n12016 , n12017 , n12018 , n12019 , n12020 , n12021 , n12022 , n12023 , n12024 , n12025 , n12026 , n12027 , n12028 , n12029 , n12030 , n12031 , n12032 , n12033 , n12034 , n12035 , n12036 , n12037 , n12038 , n12039 , n12040 , n12041 , n12042 , n12043 , n12044 , n12045 , n12046 , n12047 , n12048 , n12049 , n12050 , n12051 , n12052 , n12053 , n12054 , n12055 , n12056 , n12057 , n12058 , n12059 , n12060 , n12061 , n12062 , n12063 , n12064 , n12065 , n12066 , n12067 , n12068 , n12069 , n12070 , n12071 , n12072 , n12073 , n12074 , n12075 , n12076 , n12077 , n12078 , n12079 , n12080 , n12081 , n12082 , n12083 , n12084 , n12085 , n12086 , n12087 , n12088 , n12089 , n12090 , n12091 , n12092 , n12093 , n12094 , n12095 , n12096 , n12097 , n12098 , n12099 , n12100 , n12101 , n12102 , n12103 , n12104 , n12105 , n12106 , n12107 , n12108 , n12109 , n12110 , n12111 , n12112 , n12113 , n12114 , n12115 , n12116 , n12117 , n12118 , n12119 , n12120 , n12121 , n12122 , n12123 , n12124 , n12125 , n12126 , n12127 , n12128 , n12129 , n12130 , n12131 , n12132 , n12133 , n12134 , n12135 , n12136 , n12137 , n12138 , n12139 , n12140 , n12141 , n12142 , n12143 , n12144 , n12145 , n12146 , n12147 , n12148 , n12149 , n12150 , n12151 , n12152 , n12153 , n12154 , n12155 , n12156 , n12157 , n12158 , n12159 , n12160 , n12161 , n12162 , n12163 , n12164 , n12165 , n12166 , n12167 , n12168 , n12169 , n12170 , n12171 , n12172 , n12173 , n12174 , n12175 , n12176 , n12177 , n12178 , n12179 , n12180 , n12181 , n12182 , n12183 , n12184 , n12185 , n12186 , n12187 , n12188 , n12189 , n12190 , n12191 , n12192 , n12193 , n12194 , n12195 , n12196 , n12197 , n12198 , n12199 , n12200 , n12201 , n12202 , n12203 , n12204 , n12205 , n12206 , n12207 , n12208 , n12209 , n12210 , n12211 , n12212 , n12213 , n12214 , n12215 , n12216 , n12217 , n12218 , n12219 , n12220 , n12221 , n12222 , n12223 , n12224 , n12225 , n12226 , n12227 , n12228 , n12229 , n12230 , n12231 , n12232 , n12233 , n12234 , n12235 , n12236 , n12237 , n12238 , n12239 , n12240 , n12241 , n12242 , n12243 , n12244 , n12245 , n12246 , n12247 , n12248 , n12249 , n12250 , n12251 , n12252 , n12253 , n12254 , n12255 , n12256 , n12257 , n12258 , n12259 , n12260 , n12261 , n12262 , n12263 , n12264 , n12265 , n12266 , n12267 , n12268 , n12269 , n12270 , n12271 , n12272 , n12273 , n12274 , n12275 , n12276 , n12277 , n12278 , n12279 , n12280 , n12281 , n12282 , n12283 , n12284 , n12285 , n12286 , n12287 , n12288 , n12289 , n12290 , n12291 , n12292 , n12293 , n12294 , n12295 , n12296 , n12297 , n12298 , n12299 , n12300 , n12301 , n12302 , n12303 , n12304 , n12305 , n12306 , n12307 , n12308 , n12309 , n12310 , n12311 , n12312 , n12313 , n12314 , n12315 , n12316 , n12317 , n12318 , n12319 , n12320 , n12321 , n12322 , n12323 , n12324 , n12325 , n12326 , n12327 , n12328 , n12329 , n12330 , n12331 , n12332 , n12333 , n12334 , n12335 , n12336 , n12337 , n12338 , n12339 , n12340 , n12341 , n12342 , n12343 , n12344 , n12345 , n12346 , n12347 , n12348 , n12349 , n12350 , n12351 , n12352 , n12353 , n12354 , n12355 , n12356 , n12357 , n12358 , n12359 , n12360 , n12361 , n12362 , n12363 , n12364 , n12365 , n12366 , n12367 , n12368 , n12369 , n12370 , n12371 , n12372 , n12373 , n12374 , n12375 , n12376 , n12377 , n12378 , n12379 , n12380 , n12381 , n12382 , n12383 , n12384 , n12385 , n12386 , n12387 , n12388 , n12389 , n12390 , n12391 , n12392 , n12393 , n12394 , n12395 , n12396 , n12397 , n12398 , n12399 , n12400 , n12401 , n12402 , n12403 , n12404 , n12405 , n12406 , n12407 , n12408 , n12409 , n12410 , n12411 , n12412 , n12413 , n12414 , n12415 , n12416 , n12417 , n12418 , n12419 , n12420 , n12421 , n12422 , n12423 , n12424 , n12425 , n12426 , n12427 , n12428 , n12429 , n12430 , n12431 , n12432 , n12433 , n12434 , n12435 , n12436 , n12437 , n12438 , n12439 , n12440 , n12441 , n12442 , n12443 , n12444 , n12445 , n12446 , n12447 , n12448 , n12449 , n12450 , n12451 , n12452 , n12453 , n12454 , n12455 , n12456 , n12457 , n12458 , n12459 , n12460 , n12461 , n12462 , n12463 , n12464 , n12465 , n12466 , n12467 , n12468 , n12469 , n12470 , n12471 , n12472 , n12473 , n12474 , n12475 , n12476 , n12477 , n12478 , n12479 , n12480 , n12481 , n12482 , n12483 , n12484 , n12485 , n12486 , n12487 , n12488 , n12489 , n12490 , n12491 , n12492 , n12493 , n12494 , n12495 , n12496 , n12497 , n12498 , n12499 , n12500 , n12501 , n12502 , n12503 , n12504 , n12505 , n12506 , n12507 , n12508 , n12509 , n12510 , n12511 , n12512 , n12513 , n12514 , n12515 , n12516 , n12517 , n12518 , n12519 , n12520 , n12521 , n12522 , n12523 , n12524 , n12525 , n12526 , n12527 , n12528 , n12529 , n12530 , n12531 , n12532 , n12533 , n12534 , n12535 , n12536 , n12537 , n12538 , n12539 , n12540 , n12541 , n12542 , n12543 , n12544 , n12545 , n12546 , n12547 , n12548 , n12549 , n12550 , n12551 , n12552 , n12553 , n12554 , n12555 , n12556 , n12557 , n12558 , n12559 , n12560 , n12561 , n12562 , n12563 , n12564 , n12565 , n12566 , n12567 , n12568 , n12569 , n12570 , n12571 , n12572 , n12573 , n12574 , n12575 , n12576 , n12577 , n12578 , n12579 , n12580 , n12581 , n12582 , n12583 , n12584 , n12585 , n12586 , n12587 , n12588 , n12589 , n12590 , n12591 , n12592 , n12593 , n12594 , n12595 , n12596 , n12597 , n12598 , n12599 , n12600 , n12601 , n12602 , n12603 , n12604 , n12605 , n12606 , n12607 , n12608 , n12609 , n12610 , n12611 , n12612 , n12613 , n12614 , n12615 , n12616 , n12617 , n12618 , n12619 , n12620 , n12621 , n12622 , n12623 , n12624 , n12625 , n12626 , n12627 , n12628 , n12629 , n12630 , n12631 , n12632 , n12633 , n12634 , n12635 , n12636 , n12637 , n12638 , n12639 , n12640 , n12641 , n12642 , n12643 , n12644 , n12645 , n12646 , n12647 , n12648 , n12649 , n12650 , n12651 , n12652 , n12653 , n12654 , n12655 , n12656 , n12657 , n12658 , n12659 , n12660 , n12661 , n12662 , n12663 , n12664 , n12665 , n12666 , n12667 , n12668 , n12669 , n12670 , n12671 , n12672 , n12673 , n12674 , n12675 , n12676 , n12677 , n12678 , n12679 , n12680 , n12681 , n12682 , n12683 , n12684 , n12685 , n12686 , n12687 , n12688 , n12689 , n12690 , n12691 , n12692 , n12693 , n12694 , n12695 , n12696 , n12697 , n12698 , n12699 , n12700 , n12701 , n12702 , n12703 , n12704 , n12705 , n12706 , n12707 , n12708 , n12709 , n12710 , n12711 , n12712 , n12713 , n12714 , n12715 , n12716 , n12717 , n12718 , n12719 , n12720 , n12721 , n12722 , n12723 , n12724 , n12725 , n12726 , n12727 , n12728 , n12729 , n12730 , n12731 , n12732 , n12733 , n12734 , n12735 , n12736 , n12737 , n12738 , n12739 , n12740 , n12741 , n12742 , n12743 , n12744 , n12745 , n12746 , n12747 , n12748 , n12749 , n12750 , n12751 , n12752 , n12753 , n12754 , n12755 , n12756 , n12757 , n12758 , n12759 , n12760 , n12761 , n12762 , n12763 , n12764 , n12765 , n12766 , n12767 , n12768 , n12769 , n12770 , n12771 , n12772 , n12773 , n12774 , n12775 , n12776 , n12777 , n12778 , n12779 , n12780 , n12781 , n12782 , n12783 , n12784 , n12785 , n12786 , n12787 , n12788 , n12789 , n12790 , n12791 , n12792 , n12793 , n12794 , n12795 , n12796 , n12797 , n12798 , n12799 , n12800 , n12801 , n12802 , n12803 , n12804 , n12805 , n12806 , n12807 , n12808 , n12809 , n12810 , n12811 , n12812 , n12813 , n12814 , n12815 , n12816 , n12817 , n12818 , n12819 , n12820 , n12821 , n12822 , n12823 , n12824 , n12825 , n12826 , n12827 , n12828 , n12829 ;
  assign n476 = ~\P1_IR_reg[17]/NET0131  & ~\P1_IR_reg[18]/NET0131  ;
  assign n477 = ~\P1_IR_reg[19]/NET0131  & n476 ;
  assign n478 = ~\P1_IR_reg[16]/NET0131  & n477 ;
  assign n462 = ~\P1_IR_reg[6]/NET0131  & ~\P1_IR_reg[7]/NET0131  ;
  assign n463 = ~\P1_IR_reg[0]/NET0131  & ~\P1_IR_reg[1]/NET0131  ;
  assign n464 = ~\P1_IR_reg[2]/NET0131  & n463 ;
  assign n465 = ~\P1_IR_reg[3]/NET0131  & ~\P1_IR_reg[4]/NET0131  ;
  assign n466 = ~\P1_IR_reg[5]/NET0131  & n465 ;
  assign n467 = n464 & n466 ;
  assign n468 = n462 & n467 ;
  assign n469 = ~\P1_IR_reg[10]/NET0131  & ~\P1_IR_reg[9]/NET0131  ;
  assign n470 = ~\P1_IR_reg[11]/NET0131  & n469 ;
  assign n471 = ~\P1_IR_reg[12]/NET0131  & n470 ;
  assign n472 = ~\P1_IR_reg[13]/NET0131  & ~\P1_IR_reg[8]/NET0131  ;
  assign n473 = n471 & n472 ;
  assign n474 = n468 & n473 ;
  assign n475 = ~\P1_IR_reg[14]/NET0131  & ~\P1_IR_reg[15]/NET0131  ;
  assign n514 = n474 & n475 ;
  assign n515 = n478 & n514 ;
  assign n516 = \P1_IR_reg[31]/NET0131  & ~n515 ;
  assign n517 = \P1_IR_reg[20]/NET0131  & n516 ;
  assign n518 = ~\P1_IR_reg[20]/NET0131  & ~n516 ;
  assign n519 = ~n517 & ~n518 ;
  assign n503 = ~\P1_IR_reg[14]/NET0131  & n474 ;
  assign n504 = ~\P1_IR_reg[15]/NET0131  & ~\P1_IR_reg[16]/NET0131  ;
  assign n505 = n476 & n504 ;
  assign n506 = n503 & n505 ;
  assign n479 = ~\P1_IR_reg[20]/NET0131  & ~\P1_IR_reg[21]/NET0131  ;
  assign n502 = ~\P1_IR_reg[22]/NET0131  & n479 ;
  assign n507 = ~\P1_IR_reg[19]/NET0131  & n502 ;
  assign n508 = n506 & n507 ;
  assign n520 = ~\P1_IR_reg[23]/NET0131  & ~\P1_IR_reg[24]/NET0131  ;
  assign n521 = ~\P1_IR_reg[25]/NET0131  & ~\P1_IR_reg[26]/NET0131  ;
  assign n522 = n520 & n521 ;
  assign n523 = n508 & n522 ;
  assign n524 = \P1_IR_reg[31]/NET0131  & ~n523 ;
  assign n525 = \P1_IR_reg[27]/NET0131  & n524 ;
  assign n526 = ~\P1_IR_reg[27]/NET0131  & ~n524 ;
  assign n527 = ~n525 & ~n526 ;
  assign n528 = ~\P1_IR_reg[23]/NET0131  & n502 ;
  assign n529 = n515 & n528 ;
  assign n530 = \P1_IR_reg[31]/NET0131  & ~n529 ;
  assign n531 = ~\P1_IR_reg[24]/NET0131  & ~\P1_IR_reg[27]/NET0131  ;
  assign n532 = n521 & n531 ;
  assign n533 = \P1_IR_reg[31]/NET0131  & ~n532 ;
  assign n534 = ~n530 & ~n533 ;
  assign n535 = \P1_IR_reg[28]/NET0131  & ~n534 ;
  assign n536 = ~\P1_IR_reg[28]/NET0131  & n534 ;
  assign n537 = ~n535 & ~n536 ;
  assign n538 = ~n527 & ~n537 ;
  assign n544 = ~\P2_datao_reg[22]/NET0131  & ~\si[22]_pad  ;
  assign n545 = \P2_datao_reg[22]/NET0131  & \si[22]_pad  ;
  assign n546 = \P2_datao_reg[21]/NET0131  & \si[21]_pad  ;
  assign n547 = ~n545 & ~n546 ;
  assign n548 = ~n544 & ~n547 ;
  assign n549 = ~\P2_datao_reg[21]/NET0131  & ~\si[21]_pad  ;
  assign n550 = ~n544 & ~n549 ;
  assign n551 = ~\P2_datao_reg[20]/NET0131  & ~\si[20]_pad  ;
  assign n552 = \P2_datao_reg[20]/NET0131  & \si[20]_pad  ;
  assign n553 = \P2_datao_reg[19]/NET0131  & \si[19]_pad  ;
  assign n554 = ~n552 & ~n553 ;
  assign n555 = ~n551 & ~n554 ;
  assign n556 = n550 & n555 ;
  assign n557 = ~n548 & ~n556 ;
  assign n558 = ~\P2_datao_reg[19]/NET0131  & ~\si[19]_pad  ;
  assign n559 = ~n551 & ~n558 ;
  assign n560 = n550 & n559 ;
  assign n561 = ~\P2_datao_reg[18]/NET0131  & ~\si[18]_pad  ;
  assign n562 = \P2_datao_reg[18]/NET0131  & \si[18]_pad  ;
  assign n563 = \P2_datao_reg[17]/NET0131  & \si[17]_pad  ;
  assign n564 = ~n562 & ~n563 ;
  assign n565 = ~n561 & ~n564 ;
  assign n566 = ~\P2_datao_reg[17]/NET0131  & ~\si[17]_pad  ;
  assign n567 = ~n561 & ~n566 ;
  assign n568 = ~\P2_datao_reg[16]/NET0131  & ~\si[16]_pad  ;
  assign n569 = \P2_datao_reg[15]/NET0131  & \si[15]_pad  ;
  assign n570 = \P2_datao_reg[16]/NET0131  & \si[16]_pad  ;
  assign n571 = ~n569 & ~n570 ;
  assign n572 = ~n568 & ~n571 ;
  assign n573 = n567 & n572 ;
  assign n574 = ~n565 & ~n573 ;
  assign n575 = ~\P2_datao_reg[14]/NET0131  & ~\si[14]_pad  ;
  assign n576 = \P2_datao_reg[14]/NET0131  & \si[14]_pad  ;
  assign n577 = \P2_datao_reg[13]/NET0131  & \si[13]_pad  ;
  assign n578 = ~n576 & ~n577 ;
  assign n579 = ~n575 & ~n578 ;
  assign n580 = ~\P2_datao_reg[13]/NET0131  & ~\si[13]_pad  ;
  assign n581 = ~n575 & ~n580 ;
  assign n582 = ~\P2_datao_reg[12]/NET0131  & ~\si[12]_pad  ;
  assign n583 = \P2_datao_reg[12]/NET0131  & \si[12]_pad  ;
  assign n584 = \P2_datao_reg[11]/NET0131  & \si[11]_pad  ;
  assign n585 = ~n583 & ~n584 ;
  assign n586 = ~n582 & ~n585 ;
  assign n587 = n581 & n586 ;
  assign n588 = ~n579 & ~n587 ;
  assign n602 = ~\P2_datao_reg[6]/NET0131  & ~\si[6]_pad  ;
  assign n603 = \P2_datao_reg[5]/NET0131  & \si[5]_pad  ;
  assign n604 = \P2_datao_reg[6]/NET0131  & \si[6]_pad  ;
  assign n605 = ~n603 & ~n604 ;
  assign n606 = ~n602 & ~n605 ;
  assign n607 = \P2_datao_reg[4]/NET0131  & \si[4]_pad  ;
  assign n608 = \P2_datao_reg[3]/NET0131  & \si[3]_pad  ;
  assign n609 = ~\P2_datao_reg[3]/NET0131  & ~\si[3]_pad  ;
  assign n610 = ~\P2_datao_reg[2]/NET0131  & ~\si[2]_pad  ;
  assign n611 = ~n609 & ~n610 ;
  assign n612 = \P2_datao_reg[0]/NET0131  & \si[0]_pad  ;
  assign n613 = ~\P2_datao_reg[1]/NET0131  & ~\si[1]_pad  ;
  assign n614 = n612 & ~n613 ;
  assign n615 = \P2_datao_reg[1]/NET0131  & \si[1]_pad  ;
  assign n616 = \P2_datao_reg[2]/NET0131  & \si[2]_pad  ;
  assign n617 = ~n615 & ~n616 ;
  assign n618 = ~n614 & n617 ;
  assign n619 = n611 & ~n618 ;
  assign n620 = ~n608 & ~n619 ;
  assign n621 = ~n607 & n620 ;
  assign n622 = ~\P2_datao_reg[5]/NET0131  & ~\si[5]_pad  ;
  assign n623 = ~\P2_datao_reg[4]/NET0131  & ~\si[4]_pad  ;
  assign n624 = ~n622 & ~n623 ;
  assign n625 = ~n602 & n624 ;
  assign n626 = ~n621 & n625 ;
  assign n627 = ~n606 & ~n626 ;
  assign n592 = ~\P2_datao_reg[9]/NET0131  & ~\si[9]_pad  ;
  assign n593 = ~\P2_datao_reg[10]/NET0131  & ~\si[10]_pad  ;
  assign n594 = ~n592 & ~n593 ;
  assign n595 = ~\P2_datao_reg[8]/NET0131  & ~\si[8]_pad  ;
  assign n628 = ~\P2_datao_reg[7]/NET0131  & ~\si[7]_pad  ;
  assign n629 = ~n595 & ~n628 ;
  assign n630 = n594 & n629 ;
  assign n631 = ~n627 & n630 ;
  assign n589 = \P2_datao_reg[8]/NET0131  & \si[8]_pad  ;
  assign n590 = \P2_datao_reg[7]/NET0131  & \si[7]_pad  ;
  assign n591 = ~n589 & ~n590 ;
  assign n596 = n594 & ~n595 ;
  assign n597 = ~n591 & n596 ;
  assign n598 = \P2_datao_reg[9]/NET0131  & \si[9]_pad  ;
  assign n599 = \P2_datao_reg[10]/NET0131  & \si[10]_pad  ;
  assign n600 = ~n598 & ~n599 ;
  assign n601 = ~n593 & ~n600 ;
  assign n632 = ~n597 & ~n601 ;
  assign n633 = ~n631 & n632 ;
  assign n634 = ~\P2_datao_reg[11]/NET0131  & ~\si[11]_pad  ;
  assign n635 = ~n582 & ~n634 ;
  assign n636 = n581 & n635 ;
  assign n637 = ~n633 & n636 ;
  assign n638 = n588 & ~n637 ;
  assign n639 = ~\P2_datao_reg[15]/NET0131  & ~\si[15]_pad  ;
  assign n640 = ~n568 & ~n639 ;
  assign n641 = n567 & n640 ;
  assign n642 = ~n638 & n641 ;
  assign n643 = n574 & ~n642 ;
  assign n644 = n560 & ~n643 ;
  assign n645 = n557 & ~n644 ;
  assign n646 = ~\P2_datao_reg[30]/NET0131  & ~\si[30]_pad  ;
  assign n647 = ~\P2_datao_reg[29]/NET0131  & ~\si[29]_pad  ;
  assign n648 = ~\P2_datao_reg[27]/NET0131  & ~\si[27]_pad  ;
  assign n649 = ~\P2_datao_reg[28]/NET0131  & ~\si[28]_pad  ;
  assign n650 = ~n648 & ~n649 ;
  assign n651 = ~n647 & n650 ;
  assign n652 = ~n646 & n651 ;
  assign n653 = ~\P2_datao_reg[26]/NET0131  & ~\si[26]_pad  ;
  assign n654 = ~\P2_datao_reg[25]/NET0131  & ~\si[25]_pad  ;
  assign n655 = ~n653 & ~n654 ;
  assign n656 = ~\P2_datao_reg[24]/NET0131  & ~\si[24]_pad  ;
  assign n657 = ~\P2_datao_reg[23]/NET0131  & ~\si[23]_pad  ;
  assign n658 = ~n656 & ~n657 ;
  assign n659 = n655 & n658 ;
  assign n660 = n652 & n659 ;
  assign n661 = ~n645 & n660 ;
  assign n670 = \P2_datao_reg[26]/NET0131  & \si[26]_pad  ;
  assign n671 = \P2_datao_reg[25]/NET0131  & \si[25]_pad  ;
  assign n672 = ~n670 & ~n671 ;
  assign n673 = ~n653 & ~n672 ;
  assign n674 = \P2_datao_reg[24]/NET0131  & \si[24]_pad  ;
  assign n675 = \P2_datao_reg[23]/NET0131  & \si[23]_pad  ;
  assign n676 = ~n674 & ~n675 ;
  assign n677 = ~n656 & ~n676 ;
  assign n678 = n655 & n677 ;
  assign n679 = ~n673 & ~n678 ;
  assign n680 = n652 & ~n679 ;
  assign n662 = \P2_datao_reg[29]/NET0131  & \si[29]_pad  ;
  assign n663 = \P2_datao_reg[27]/NET0131  & \si[27]_pad  ;
  assign n664 = \P2_datao_reg[28]/NET0131  & \si[28]_pad  ;
  assign n665 = ~n663 & ~n664 ;
  assign n666 = ~n647 & ~n649 ;
  assign n667 = ~n665 & n666 ;
  assign n668 = ~n662 & ~n667 ;
  assign n669 = ~n646 & ~n668 ;
  assign n681 = \P2_datao_reg[30]/NET0131  & \si[30]_pad  ;
  assign n682 = ~n669 & ~n681 ;
  assign n683 = ~n680 & n682 ;
  assign n684 = ~n661 & n683 ;
  assign n686 = ~\si[31]_pad  & n684 ;
  assign n539 = ~\P1_addr_reg[19]/NET0131  & ~\P2_addr_reg[19]/NET0131  ;
  assign n540 = ~\P1_rd_reg/NET0131  & n539 ;
  assign n541 = \P1_addr_reg[19]/NET0131  & \P2_addr_reg[19]/NET0131  ;
  assign n542 = ~\P2_rd_reg/NET0131  & n541 ;
  assign n543 = ~n540 & ~n542 ;
  assign n685 = \si[31]_pad  & ~n684 ;
  assign n687 = ~n543 & ~n685 ;
  assign n688 = ~n686 & n687 ;
  assign n689 = \P2_datao_reg[31]/NET0131  & n688 ;
  assign n690 = ~\P2_datao_reg[31]/NET0131  & ~n688 ;
  assign n691 = ~n689 & ~n690 ;
  assign n692 = ~n538 & n691 ;
  assign n480 = n475 & n479 ;
  assign n481 = n478 & n480 ;
  assign n482 = n474 & n481 ;
  assign n693 = ~\P1_IR_reg[22]/NET0131  & ~\P1_IR_reg[25]/NET0131  ;
  assign n694 = n520 & n693 ;
  assign n695 = n482 & n694 ;
  assign n696 = \P1_IR_reg[31]/NET0131  & ~n695 ;
  assign n697 = ~\P1_IR_reg[27]/NET0131  & ~\P1_IR_reg[28]/NET0131  ;
  assign n698 = ~\P1_IR_reg[29]/NET0131  & n697 ;
  assign n699 = ~\P1_IR_reg[26]/NET0131  & n698 ;
  assign n700 = \P1_IR_reg[31]/NET0131  & ~n699 ;
  assign n701 = ~n696 & ~n700 ;
  assign n702 = \P1_IR_reg[30]/NET0131  & ~n701 ;
  assign n703 = ~\P1_IR_reg[30]/NET0131  & n701 ;
  assign n704 = ~n702 & ~n703 ;
  assign n487 = ~\P1_IR_reg[3]/NET0131  & n464 ;
  assign n488 = ~\P1_IR_reg[4]/NET0131  & n487 ;
  assign n489 = ~\P1_IR_reg[8]/NET0131  & n462 ;
  assign n490 = ~\P1_IR_reg[5]/NET0131  & n489 ;
  assign n491 = n488 & n490 ;
  assign n492 = ~\P1_IR_reg[13]/NET0131  & ~\P1_IR_reg[16]/NET0131  ;
  assign n493 = n475 & n492 ;
  assign n494 = n471 & n493 ;
  assign n495 = n491 & n494 ;
  assign n705 = ~\P1_IR_reg[24]/NET0131  & n477 ;
  assign n706 = n528 & n705 ;
  assign n707 = n495 & n706 ;
  assign n708 = \P1_IR_reg[31]/NET0131  & ~n707 ;
  assign n709 = n521 & n697 ;
  assign n710 = \P1_IR_reg[31]/NET0131  & ~n709 ;
  assign n711 = ~n708 & ~n710 ;
  assign n712 = \P1_IR_reg[29]/NET0131  & ~n711 ;
  assign n713 = ~\P1_IR_reg[29]/NET0131  & n711 ;
  assign n714 = ~n712 & ~n713 ;
  assign n715 = n704 & n714 ;
  assign n716 = \P1_reg3_reg[3]/NET0131  & \P1_reg3_reg[4]/NET0131  ;
  assign n717 = \P1_reg3_reg[5]/NET0131  & n716 ;
  assign n718 = \P1_reg3_reg[6]/NET0131  & n717 ;
  assign n719 = \P1_reg3_reg[7]/NET0131  & n718 ;
  assign n720 = \P1_reg3_reg[8]/NET0131  & n719 ;
  assign n721 = \P1_reg3_reg[9]/NET0131  & n720 ;
  assign n722 = \P1_reg3_reg[10]/NET0131  & n721 ;
  assign n723 = \P1_reg3_reg[11]/NET0131  & n722 ;
  assign n724 = \P1_reg3_reg[12]/NET0131  & \P1_reg3_reg[13]/NET0131  ;
  assign n725 = n723 & n724 ;
  assign n726 = \P1_reg3_reg[14]/NET0131  & \P1_reg3_reg[15]/NET0131  ;
  assign n727 = \P1_reg3_reg[16]/NET0131  & n726 ;
  assign n728 = n725 & n727 ;
  assign n731 = \P1_reg3_reg[19]/NET0131  & \P1_reg3_reg[22]/NET0131  ;
  assign n732 = \P1_reg3_reg[23]/NET0131  & \P1_reg3_reg[24]/NET0131  ;
  assign n733 = n731 & n732 ;
  assign n729 = \P1_reg3_reg[20]/NET0131  & \P1_reg3_reg[21]/NET0131  ;
  assign n730 = \P1_reg3_reg[17]/NET0131  & \P1_reg3_reg[18]/NET0131  ;
  assign n734 = n729 & n730 ;
  assign n735 = n733 & n734 ;
  assign n736 = n728 & n735 ;
  assign n737 = \P1_reg3_reg[25]/NET0131  & \P1_reg3_reg[26]/NET0131  ;
  assign n738 = \P1_reg3_reg[27]/NET0131  & \P1_reg3_reg[28]/NET0131  ;
  assign n739 = n737 & n738 ;
  assign n740 = n736 & n739 ;
  assign n741 = n715 & n740 ;
  assign n742 = n704 & ~n714 ;
  assign n743 = \P1_reg2_reg[31]/NET0131  & n742 ;
  assign n748 = ~n741 & ~n743 ;
  assign n744 = ~n704 & ~n714 ;
  assign n745 = \P1_reg0_reg[31]/NET0131  & n744 ;
  assign n746 = ~n704 & n714 ;
  assign n747 = \P1_reg1_reg[31]/NET0131  & n746 ;
  assign n749 = ~n745 & ~n747 ;
  assign n750 = n748 & n749 ;
  assign n751 = \P2_datao_reg[30]/NET0131  & n543 ;
  assign n752 = ~n646 & ~n681 ;
  assign n767 = ~n546 & ~n552 ;
  assign n768 = ~n549 & ~n767 ;
  assign n769 = ~n549 & ~n551 ;
  assign n770 = ~n553 & ~n562 ;
  assign n771 = ~n558 & ~n770 ;
  assign n772 = n769 & n771 ;
  assign n773 = ~n768 & ~n772 ;
  assign n774 = ~n577 & ~n583 ;
  assign n775 = ~n584 & ~n599 ;
  assign n776 = n635 & ~n775 ;
  assign n777 = n774 & ~n776 ;
  assign n778 = ~n580 & ~n777 ;
  assign n779 = ~n614 & ~n615 ;
  assign n780 = n611 & ~n779 ;
  assign n781 = ~n609 & n616 ;
  assign n782 = ~n608 & ~n781 ;
  assign n783 = ~n780 & n782 ;
  assign n784 = n624 & ~n783 ;
  assign n785 = ~n603 & ~n607 ;
  assign n786 = ~n622 & ~n785 ;
  assign n787 = ~n784 & ~n786 ;
  assign n788 = ~n592 & n629 ;
  assign n789 = ~n602 & n788 ;
  assign n790 = ~n787 & n789 ;
  assign n791 = ~n589 & ~n598 ;
  assign n792 = ~n592 & ~n791 ;
  assign n793 = ~n590 & ~n604 ;
  assign n794 = n788 & ~n793 ;
  assign n795 = ~n792 & ~n794 ;
  assign n796 = ~n790 & n795 ;
  assign n797 = ~n580 & ~n593 ;
  assign n798 = n635 & n797 ;
  assign n799 = ~n796 & n798 ;
  assign n800 = ~n778 & ~n799 ;
  assign n801 = ~n566 & ~n575 ;
  assign n802 = n640 & n801 ;
  assign n803 = ~n800 & n802 ;
  assign n804 = ~n563 & ~n570 ;
  assign n805 = ~n569 & ~n576 ;
  assign n806 = n640 & ~n805 ;
  assign n807 = n804 & ~n806 ;
  assign n808 = ~n566 & ~n807 ;
  assign n809 = ~n803 & ~n808 ;
  assign n810 = ~n558 & ~n561 ;
  assign n811 = n769 & n810 ;
  assign n812 = ~n809 & n811 ;
  assign n813 = n773 & ~n812 ;
  assign n754 = n651 & ~n653 ;
  assign n757 = ~n654 & ~n656 ;
  assign n765 = ~n544 & ~n657 ;
  assign n766 = n757 & n765 ;
  assign n814 = n754 & n766 ;
  assign n815 = ~n813 & n814 ;
  assign n755 = ~n671 & ~n674 ;
  assign n756 = ~n654 & ~n755 ;
  assign n758 = ~n545 & ~n675 ;
  assign n759 = ~n657 & ~n758 ;
  assign n760 = n757 & n759 ;
  assign n761 = ~n756 & ~n760 ;
  assign n762 = n754 & ~n761 ;
  assign n763 = ~n663 & ~n670 ;
  assign n764 = n651 & ~n763 ;
  assign n753 = ~n647 & n664 ;
  assign n816 = ~n662 & ~n753 ;
  assign n817 = ~n764 & n816 ;
  assign n818 = ~n762 & n817 ;
  assign n819 = ~n815 & n818 ;
  assign n821 = ~n752 & n819 ;
  assign n820 = n752 & ~n819 ;
  assign n822 = ~n543 & ~n820 ;
  assign n823 = ~n821 & n822 ;
  assign n824 = ~n751 & ~n823 ;
  assign n825 = ~n538 & ~n824 ;
  assign n826 = \P1_reg2_reg[30]/NET0131  & n742 ;
  assign n829 = ~n741 & ~n826 ;
  assign n827 = \P1_reg0_reg[30]/NET0131  & n744 ;
  assign n828 = \P1_reg1_reg[30]/NET0131  & n746 ;
  assign n830 = ~n827 & ~n828 ;
  assign n831 = n829 & n830 ;
  assign n832 = ~n825 & ~n831 ;
  assign n833 = ~n750 & ~n832 ;
  assign n834 = n692 & ~n833 ;
  assign n838 = \P2_datao_reg[29]/NET0131  & n543 ;
  assign n839 = ~n647 & ~n662 ;
  assign n840 = n548 & n658 ;
  assign n841 = ~n677 & ~n840 ;
  assign n842 = n655 & ~n841 ;
  assign n843 = ~n673 & ~n842 ;
  assign n844 = ~n648 & ~n843 ;
  assign n845 = n665 & ~n844 ;
  assign n846 = ~n649 & ~n845 ;
  assign n847 = n559 & n565 ;
  assign n848 = ~n555 & ~n847 ;
  assign n849 = n579 & n640 ;
  assign n850 = ~n572 & ~n849 ;
  assign n853 = ~n620 & ~n623 ;
  assign n854 = ~n607 & ~n853 ;
  assign n855 = ~n602 & ~n628 ;
  assign n856 = ~n595 & ~n622 ;
  assign n857 = n855 & n856 ;
  assign n858 = ~n854 & n857 ;
  assign n851 = ~n590 & ~n606 ;
  assign n852 = n629 & ~n851 ;
  assign n859 = ~n589 & ~n852 ;
  assign n860 = ~n858 & n859 ;
  assign n861 = n594 & n635 ;
  assign n862 = ~n860 & n861 ;
  assign n863 = n601 & n635 ;
  assign n864 = ~n586 & ~n863 ;
  assign n865 = ~n862 & n864 ;
  assign n866 = n581 & n640 ;
  assign n867 = ~n865 & n866 ;
  assign n868 = n850 & ~n867 ;
  assign n869 = n559 & n567 ;
  assign n870 = ~n868 & n869 ;
  assign n871 = n848 & ~n870 ;
  assign n872 = n550 & n659 ;
  assign n873 = n650 & n872 ;
  assign n874 = ~n871 & n873 ;
  assign n875 = ~n846 & ~n874 ;
  assign n877 = ~n839 & n875 ;
  assign n876 = n839 & ~n875 ;
  assign n878 = ~n543 & ~n876 ;
  assign n879 = ~n877 & n878 ;
  assign n880 = ~n838 & ~n879 ;
  assign n881 = ~n538 & ~n880 ;
  assign n882 = \P1_reg1_reg[29]/NET0131  & n746 ;
  assign n885 = ~n741 & ~n882 ;
  assign n883 = \P1_reg0_reg[29]/NET0131  & n744 ;
  assign n884 = \P1_reg2_reg[29]/NET0131  & n742 ;
  assign n886 = ~n883 & ~n884 ;
  assign n887 = n885 & n886 ;
  assign n888 = n881 & n887 ;
  assign n889 = \P2_datao_reg[28]/NET0131  & n543 ;
  assign n890 = ~n649 & ~n664 ;
  assign n891 = ~n653 & n756 ;
  assign n892 = n763 & ~n891 ;
  assign n893 = ~n648 & ~n892 ;
  assign n894 = ~n599 & ~n792 ;
  assign n895 = ~n593 & ~n634 ;
  assign n896 = ~n894 & n895 ;
  assign n897 = ~n584 & ~n896 ;
  assign n898 = ~n582 & ~n897 ;
  assign n899 = n774 & ~n898 ;
  assign n900 = n581 & ~n899 ;
  assign n901 = n805 & ~n900 ;
  assign n902 = ~n639 & ~n901 ;
  assign n903 = ~n604 & ~n786 ;
  assign n904 = ~n784 & n903 ;
  assign n905 = n855 & ~n904 ;
  assign n906 = ~n590 & ~n905 ;
  assign n907 = n596 & ~n634 ;
  assign n908 = ~n906 & n907 ;
  assign n909 = ~n582 & ~n639 ;
  assign n910 = n581 & n909 ;
  assign n911 = n908 & n910 ;
  assign n912 = ~n902 & ~n911 ;
  assign n913 = ~n558 & n567 ;
  assign n914 = ~n568 & n913 ;
  assign n915 = ~n912 & n914 ;
  assign n916 = ~n804 & n913 ;
  assign n917 = ~n771 & ~n916 ;
  assign n918 = ~n915 & n917 ;
  assign n919 = n765 & n769 ;
  assign n920 = ~n918 & n919 ;
  assign n921 = n765 & n768 ;
  assign n922 = ~n759 & ~n921 ;
  assign n923 = ~n920 & n922 ;
  assign n924 = ~n648 & ~n656 ;
  assign n925 = n655 & n924 ;
  assign n926 = ~n923 & n925 ;
  assign n927 = ~n893 & ~n926 ;
  assign n929 = ~n890 & n927 ;
  assign n928 = n890 & ~n927 ;
  assign n930 = ~n543 & ~n928 ;
  assign n931 = ~n929 & n930 ;
  assign n932 = ~n889 & ~n931 ;
  assign n933 = ~n538 & ~n932 ;
  assign n937 = \P1_reg3_reg[25]/NET0131  & n736 ;
  assign n938 = \P1_reg3_reg[26]/NET0131  & n937 ;
  assign n939 = \P1_reg3_reg[27]/NET0131  & n938 ;
  assign n940 = ~\P1_reg3_reg[28]/NET0131  & ~n939 ;
  assign n941 = ~n740 & ~n940 ;
  assign n942 = n715 & n941 ;
  assign n936 = \P1_reg2_reg[28]/NET0131  & n742 ;
  assign n934 = \P1_reg0_reg[28]/NET0131  & n744 ;
  assign n935 = \P1_reg1_reg[28]/NET0131  & n746 ;
  assign n943 = ~n934 & ~n935 ;
  assign n944 = ~n936 & n943 ;
  assign n945 = ~n942 & n944 ;
  assign n946 = ~n933 & ~n945 ;
  assign n947 = ~n881 & ~n887 ;
  assign n948 = ~n946 & ~n947 ;
  assign n949 = ~n888 & ~n948 ;
  assign n950 = n933 & n945 ;
  assign n951 = ~n888 & ~n950 ;
  assign n1302 = \P2_datao_reg[22]/NET0131  & n543 ;
  assign n1303 = ~n544 & ~n545 ;
  assign n1305 = n813 & ~n1303 ;
  assign n1304 = ~n813 & n1303 ;
  assign n1306 = ~n543 & ~n1304 ;
  assign n1307 = ~n1305 & n1306 ;
  assign n1308 = ~n1302 & ~n1307 ;
  assign n1309 = ~n538 & ~n1308 ;
  assign n1051 = \P1_reg3_reg[17]/NET0131  & n728 ;
  assign n1052 = \P1_reg3_reg[18]/NET0131  & n1051 ;
  assign n1053 = \P1_reg3_reg[19]/NET0131  & n1052 ;
  assign n1054 = n729 & n1053 ;
  assign n1055 = \P1_reg3_reg[22]/NET0131  & n1054 ;
  assign n1313 = ~\P1_reg3_reg[22]/NET0131  & ~n1054 ;
  assign n1314 = ~n1055 & ~n1313 ;
  assign n1315 = n715 & n1314 ;
  assign n1312 = \P1_reg0_reg[22]/NET0131  & n744 ;
  assign n1310 = \P1_reg2_reg[22]/NET0131  & n742 ;
  assign n1311 = \P1_reg1_reg[22]/NET0131  & n746 ;
  assign n1316 = ~n1310 & ~n1311 ;
  assign n1317 = ~n1312 & n1316 ;
  assign n1318 = ~n1315 & n1317 ;
  assign n1319 = n1309 & n1318 ;
  assign n1320 = \P2_datao_reg[23]/NET0131  & n543 ;
  assign n1321 = ~n657 & ~n675 ;
  assign n1323 = n645 & ~n1321 ;
  assign n1322 = ~n645 & n1321 ;
  assign n1324 = ~n543 & ~n1322 ;
  assign n1325 = ~n1323 & n1324 ;
  assign n1326 = ~n1320 & ~n1325 ;
  assign n1327 = ~n538 & ~n1326 ;
  assign n1056 = \P1_reg3_reg[23]/NET0131  & n1055 ;
  assign n1329 = ~\P1_reg3_reg[23]/NET0131  & ~n1055 ;
  assign n1330 = ~n1056 & ~n1329 ;
  assign n1331 = n715 & n1330 ;
  assign n1333 = \P1_reg2_reg[23]/NET0131  & n742 ;
  assign n1328 = \P1_reg0_reg[23]/NET0131  & n744 ;
  assign n1332 = \P1_reg1_reg[23]/NET0131  & n746 ;
  assign n1334 = ~n1328 & ~n1332 ;
  assign n1335 = ~n1333 & n1334 ;
  assign n1336 = ~n1331 & n1335 ;
  assign n1337 = n1327 & n1336 ;
  assign n1338 = ~n1319 & ~n1337 ;
  assign n1339 = \P2_datao_reg[21]/NET0131  & n543 ;
  assign n1340 = ~n546 & ~n549 ;
  assign n1342 = n871 & ~n1340 ;
  assign n1341 = ~n871 & n1340 ;
  assign n1343 = ~n543 & ~n1341 ;
  assign n1344 = ~n1342 & n1343 ;
  assign n1345 = ~n1339 & ~n1344 ;
  assign n1346 = ~n538 & ~n1345 ;
  assign n1350 = \P1_reg3_reg[20]/NET0131  & n1053 ;
  assign n1351 = ~\P1_reg3_reg[21]/NET0131  & ~n1350 ;
  assign n1352 = ~n1054 & ~n1351 ;
  assign n1353 = n715 & n1352 ;
  assign n1349 = \P1_reg1_reg[21]/NET0131  & n746 ;
  assign n1347 = \P1_reg0_reg[21]/NET0131  & n744 ;
  assign n1348 = \P1_reg2_reg[21]/NET0131  & n742 ;
  assign n1354 = ~n1347 & ~n1348 ;
  assign n1355 = ~n1349 & n1354 ;
  assign n1356 = ~n1353 & n1355 ;
  assign n1357 = n1346 & n1356 ;
  assign n1698 = ~n1346 & ~n1356 ;
  assign n1358 = \P2_datao_reg[20]/NET0131  & n543 ;
  assign n1359 = ~n551 & ~n552 ;
  assign n1361 = n918 & ~n1359 ;
  assign n1360 = ~n918 & n1359 ;
  assign n1362 = ~n543 & ~n1360 ;
  assign n1363 = ~n1361 & n1362 ;
  assign n1364 = ~n1358 & ~n1363 ;
  assign n1365 = ~n538 & ~n1364 ;
  assign n1369 = ~\P1_reg3_reg[20]/NET0131  & ~n1053 ;
  assign n1370 = ~n1350 & ~n1369 ;
  assign n1371 = n715 & n1370 ;
  assign n1368 = \P1_reg1_reg[20]/NET0131  & n746 ;
  assign n1366 = \P1_reg0_reg[20]/NET0131  & n744 ;
  assign n1367 = \P1_reg2_reg[20]/NET0131  & n742 ;
  assign n1372 = ~n1366 & ~n1367 ;
  assign n1373 = ~n1368 & n1372 ;
  assign n1374 = ~n1371 & n1373 ;
  assign n1704 = ~n1365 & ~n1374 ;
  assign n1705 = ~n1698 & ~n1704 ;
  assign n1706 = ~n1357 & ~n1705 ;
  assign n1707 = n1338 & n1706 ;
  assign n1697 = ~n1327 & ~n1336 ;
  assign n1699 = ~n1309 & ~n1318 ;
  assign n1708 = ~n1697 & ~n1699 ;
  assign n1709 = ~n1337 & ~n1708 ;
  assign n1710 = ~n1707 & ~n1709 ;
  assign n1378 = \P1_IR_reg[31]/NET0131  & ~n514 ;
  assign n1379 = ~\P1_IR_reg[16]/NET0131  & ~\P1_IR_reg[17]/NET0131  ;
  assign n1380 = \P1_IR_reg[31]/NET0131  & ~n1379 ;
  assign n1381 = ~n1378 & ~n1380 ;
  assign n1382 = \P1_IR_reg[18]/NET0131  & ~n1381 ;
  assign n1383 = ~\P1_IR_reg[18]/NET0131  & n1381 ;
  assign n1384 = ~n1382 & ~n1383 ;
  assign n1385 = n538 & ~n1384 ;
  assign n1386 = \P2_datao_reg[18]/NET0131  & n543 ;
  assign n1387 = ~n561 & ~n562 ;
  assign n1389 = n809 & ~n1387 ;
  assign n1388 = ~n809 & n1387 ;
  assign n1390 = ~n543 & ~n1388 ;
  assign n1391 = ~n1389 & n1390 ;
  assign n1392 = ~n1386 & ~n1391 ;
  assign n1393 = ~n538 & n1392 ;
  assign n1394 = ~n1385 & ~n1393 ;
  assign n1398 = ~\P1_reg3_reg[18]/NET0131  & ~n1051 ;
  assign n1399 = ~n1052 & ~n1398 ;
  assign n1400 = n715 & n1399 ;
  assign n1397 = \P1_reg2_reg[18]/NET0131  & n742 ;
  assign n1395 = \P1_reg1_reg[18]/NET0131  & n746 ;
  assign n1396 = \P1_reg0_reg[18]/NET0131  & n744 ;
  assign n1401 = ~n1395 & ~n1396 ;
  assign n1402 = ~n1397 & n1401 ;
  assign n1403 = ~n1400 & n1402 ;
  assign n1404 = n1394 & n1403 ;
  assign n1405 = \P1_IR_reg[31]/NET0131  & ~n506 ;
  assign n1406 = ~\P1_IR_reg[19]/NET0131  & ~n1405 ;
  assign n1407 = \P1_IR_reg[19]/NET0131  & n1405 ;
  assign n1408 = ~n1406 & ~n1407 ;
  assign n1409 = n538 & ~n1408 ;
  assign n1410 = \P2_datao_reg[19]/NET0131  & n543 ;
  assign n1411 = ~n553 & ~n558 ;
  assign n1413 = n643 & ~n1411 ;
  assign n1412 = ~n643 & n1411 ;
  assign n1414 = ~n543 & ~n1412 ;
  assign n1415 = ~n1413 & n1414 ;
  assign n1416 = ~n1410 & ~n1415 ;
  assign n1417 = ~n538 & n1416 ;
  assign n1418 = ~n1409 & ~n1417 ;
  assign n1422 = ~\P1_reg3_reg[19]/NET0131  & ~n1052 ;
  assign n1423 = ~n1053 & ~n1422 ;
  assign n1424 = n715 & n1423 ;
  assign n1421 = \P1_reg1_reg[19]/NET0131  & n746 ;
  assign n1419 = \P1_reg0_reg[19]/NET0131  & n744 ;
  assign n1420 = \P1_reg2_reg[19]/NET0131  & n742 ;
  assign n1425 = ~n1419 & ~n1420 ;
  assign n1426 = ~n1421 & n1425 ;
  assign n1427 = ~n1424 & n1426 ;
  assign n1428 = n1418 & n1427 ;
  assign n1429 = ~n1404 & ~n1428 ;
  assign n1430 = \P1_IR_reg[31]/NET0131  & ~n495 ;
  assign n1431 = \P1_IR_reg[17]/NET0131  & ~n1430 ;
  assign n1432 = ~\P1_IR_reg[17]/NET0131  & n1430 ;
  assign n1433 = ~n1431 & ~n1432 ;
  assign n1434 = n538 & n1433 ;
  assign n1435 = \P2_datao_reg[17]/NET0131  & n543 ;
  assign n1436 = ~n563 & ~n566 ;
  assign n1438 = n868 & ~n1436 ;
  assign n1437 = ~n868 & n1436 ;
  assign n1439 = ~n543 & ~n1437 ;
  assign n1440 = ~n1438 & n1439 ;
  assign n1441 = ~n1435 & ~n1440 ;
  assign n1442 = ~n538 & n1441 ;
  assign n1443 = ~n1434 & ~n1442 ;
  assign n1444 = \P1_reg0_reg[17]/NET0131  & n744 ;
  assign n1445 = \P1_reg1_reg[17]/NET0131  & n746 ;
  assign n1450 = ~n1444 & ~n1445 ;
  assign n1446 = ~\P1_reg3_reg[17]/NET0131  & ~n728 ;
  assign n1447 = ~n1051 & ~n1446 ;
  assign n1448 = n715 & n1447 ;
  assign n1449 = \P1_reg2_reg[17]/NET0131  & n742 ;
  assign n1451 = ~n1448 & ~n1449 ;
  assign n1452 = n1450 & n1451 ;
  assign n1453 = n1443 & n1452 ;
  assign n1711 = ~n1443 & ~n1452 ;
  assign n1454 = ~\P1_IR_reg[16]/NET0131  & ~n1378 ;
  assign n1455 = \P1_IR_reg[16]/NET0131  & n1378 ;
  assign n1456 = ~n1454 & ~n1455 ;
  assign n1457 = n538 & ~n1456 ;
  assign n1458 = \P2_datao_reg[16]/NET0131  & n543 ;
  assign n1459 = ~n568 & ~n570 ;
  assign n1461 = n912 & ~n1459 ;
  assign n1460 = ~n912 & n1459 ;
  assign n1462 = ~n543 & ~n1460 ;
  assign n1463 = ~n1461 & n1462 ;
  assign n1464 = ~n1458 & ~n1463 ;
  assign n1465 = ~n538 & n1464 ;
  assign n1466 = ~n1457 & ~n1465 ;
  assign n1085 = \P1_reg3_reg[14]/NET0131  & n725 ;
  assign n1086 = \P1_reg3_reg[15]/NET0131  & n1085 ;
  assign n1470 = ~\P1_reg3_reg[16]/NET0131  & ~n1086 ;
  assign n1471 = ~n728 & ~n1470 ;
  assign n1472 = n715 & n1471 ;
  assign n1469 = \P1_reg1_reg[16]/NET0131  & n746 ;
  assign n1467 = \P1_reg0_reg[16]/NET0131  & n744 ;
  assign n1468 = \P1_reg2_reg[16]/NET0131  & n742 ;
  assign n1473 = ~n1467 & ~n1468 ;
  assign n1474 = ~n1469 & n1473 ;
  assign n1475 = ~n1472 & n1474 ;
  assign n1712 = ~n1466 & ~n1475 ;
  assign n1713 = ~n1711 & ~n1712 ;
  assign n1714 = ~n1453 & ~n1713 ;
  assign n1715 = n1429 & n1714 ;
  assign n1716 = ~n1418 & ~n1427 ;
  assign n1717 = ~n1394 & ~n1403 ;
  assign n1718 = ~n1716 & ~n1717 ;
  assign n1719 = ~n1428 & ~n1718 ;
  assign n1720 = ~n1715 & ~n1719 ;
  assign n1721 = n1710 & n1720 ;
  assign n952 = \P2_datao_reg[27]/NET0131  & n543 ;
  assign n953 = ~n648 & ~n663 ;
  assign n959 = n559 & n641 ;
  assign n960 = n872 & n959 ;
  assign n961 = n637 & n960 ;
  assign n954 = ~n588 & n641 ;
  assign n955 = n574 & ~n954 ;
  assign n956 = n560 & ~n955 ;
  assign n957 = n557 & ~n956 ;
  assign n958 = n659 & ~n957 ;
  assign n962 = n679 & ~n958 ;
  assign n963 = ~n961 & n962 ;
  assign n965 = ~n953 & n963 ;
  assign n964 = n953 & ~n963 ;
  assign n966 = ~n543 & ~n964 ;
  assign n967 = ~n965 & n966 ;
  assign n968 = ~n952 & ~n967 ;
  assign n969 = ~n538 & ~n968 ;
  assign n973 = ~\P1_reg3_reg[27]/NET0131  & ~n938 ;
  assign n974 = ~n939 & ~n973 ;
  assign n975 = n715 & n974 ;
  assign n972 = \P1_reg1_reg[27]/NET0131  & n746 ;
  assign n970 = \P1_reg0_reg[27]/NET0131  & n744 ;
  assign n971 = \P1_reg2_reg[27]/NET0131  & n742 ;
  assign n976 = ~n970 & ~n971 ;
  assign n977 = ~n972 & n976 ;
  assign n978 = ~n975 & n977 ;
  assign n979 = n969 & n978 ;
  assign n980 = \P2_datao_reg[26]/NET0131  & n543 ;
  assign n981 = ~n653 & ~n670 ;
  assign n987 = n766 & n802 ;
  assign n988 = n811 & n987 ;
  assign n989 = n799 & n988 ;
  assign n982 = n778 & n802 ;
  assign n983 = ~n808 & ~n982 ;
  assign n984 = n811 & ~n983 ;
  assign n985 = n773 & ~n984 ;
  assign n986 = n766 & ~n985 ;
  assign n990 = n761 & ~n986 ;
  assign n991 = ~n989 & n990 ;
  assign n993 = ~n981 & n991 ;
  assign n992 = n981 & ~n991 ;
  assign n994 = ~n543 & ~n992 ;
  assign n995 = ~n993 & n994 ;
  assign n996 = ~n980 & ~n995 ;
  assign n997 = ~n538 & ~n996 ;
  assign n1001 = ~\P1_reg3_reg[26]/NET0131  & ~n937 ;
  assign n1002 = ~n938 & ~n1001 ;
  assign n1003 = n715 & n1002 ;
  assign n1000 = \P1_reg0_reg[26]/NET0131  & n744 ;
  assign n998 = \P1_reg1_reg[26]/NET0131  & n746 ;
  assign n999 = \P1_reg2_reg[26]/NET0131  & n742 ;
  assign n1004 = ~n998 & ~n999 ;
  assign n1005 = ~n1000 & n1004 ;
  assign n1006 = ~n1003 & n1005 ;
  assign n1010 = n997 & n1006 ;
  assign n1298 = ~n979 & ~n1010 ;
  assign n1011 = \P2_datao_reg[25]/NET0131  & n543 ;
  assign n1012 = ~n654 & ~n671 ;
  assign n1013 = n550 & n658 ;
  assign n1019 = n866 & n869 ;
  assign n1020 = n1013 & n1019 ;
  assign n1021 = n862 & n1020 ;
  assign n1014 = ~n864 & n866 ;
  assign n1015 = n850 & ~n1014 ;
  assign n1016 = n869 & ~n1015 ;
  assign n1017 = n848 & ~n1016 ;
  assign n1018 = n1013 & ~n1017 ;
  assign n1022 = n841 & ~n1018 ;
  assign n1023 = ~n1021 & n1022 ;
  assign n1025 = ~n1012 & n1023 ;
  assign n1024 = n1012 & ~n1023 ;
  assign n1026 = ~n543 & ~n1024 ;
  assign n1027 = ~n1025 & n1026 ;
  assign n1028 = ~n1011 & ~n1027 ;
  assign n1029 = ~n538 & ~n1028 ;
  assign n1033 = ~\P1_reg3_reg[25]/NET0131  & ~n736 ;
  assign n1034 = ~n937 & ~n1033 ;
  assign n1035 = n715 & n1034 ;
  assign n1032 = \P1_reg0_reg[25]/NET0131  & n744 ;
  assign n1030 = \P1_reg2_reg[25]/NET0131  & n742 ;
  assign n1031 = \P1_reg1_reg[25]/NET0131  & n746 ;
  assign n1036 = ~n1030 & ~n1031 ;
  assign n1037 = ~n1032 & n1036 ;
  assign n1038 = ~n1035 & n1037 ;
  assign n1039 = n1029 & n1038 ;
  assign n1040 = \P2_datao_reg[24]/NET0131  & n543 ;
  assign n1041 = ~n656 & ~n674 ;
  assign n1043 = n923 & ~n1041 ;
  assign n1042 = ~n923 & n1041 ;
  assign n1044 = ~n543 & ~n1042 ;
  assign n1045 = ~n1043 & n1044 ;
  assign n1046 = ~n1040 & ~n1045 ;
  assign n1047 = ~n538 & ~n1046 ;
  assign n1057 = ~\P1_reg3_reg[24]/NET0131  & ~n1056 ;
  assign n1058 = ~n736 & ~n1057 ;
  assign n1059 = n715 & n1058 ;
  assign n1050 = \P1_reg1_reg[24]/NET0131  & n746 ;
  assign n1048 = \P1_reg2_reg[24]/NET0131  & n742 ;
  assign n1049 = \P1_reg0_reg[24]/NET0131  & n744 ;
  assign n1060 = ~n1048 & ~n1049 ;
  assign n1061 = ~n1050 & n1060 ;
  assign n1062 = ~n1059 & n1061 ;
  assign n1299 = n1047 & n1062 ;
  assign n1300 = ~n1039 & ~n1299 ;
  assign n1301 = n1298 & n1300 ;
  assign n1375 = n1365 & n1374 ;
  assign n1376 = ~n1357 & ~n1375 ;
  assign n1700 = ~n1698 & ~n1699 ;
  assign n1701 = ~n1376 & n1700 ;
  assign n1702 = n1338 & ~n1701 ;
  assign n1703 = ~n1697 & ~n1702 ;
  assign n1722 = n1301 & ~n1703 ;
  assign n1723 = ~n1721 & n1722 ;
  assign n1007 = ~n997 & ~n1006 ;
  assign n1008 = ~n969 & ~n978 ;
  assign n1009 = ~n1007 & ~n1008 ;
  assign n1063 = ~n1047 & ~n1062 ;
  assign n1064 = ~n1029 & ~n1038 ;
  assign n1065 = ~n1063 & ~n1064 ;
  assign n1066 = ~n1039 & ~n1065 ;
  assign n1067 = ~n1010 & n1066 ;
  assign n1068 = n1009 & ~n1067 ;
  assign n1069 = ~n979 & ~n1068 ;
  assign n1490 = ~\P1_reg3_reg[7]/NET0131  & ~n718 ;
  assign n1491 = ~n719 & ~n1490 ;
  assign n1492 = n715 & n1491 ;
  assign n1493 = \P1_reg2_reg[7]/NET0131  & n742 ;
  assign n1496 = ~n1492 & ~n1493 ;
  assign n1494 = \P1_reg1_reg[7]/NET0131  & n746 ;
  assign n1495 = \P1_reg0_reg[7]/NET0131  & n744 ;
  assign n1497 = ~n1494 & ~n1495 ;
  assign n1498 = n1496 & n1497 ;
  assign n1499 = \P2_datao_reg[7]/NET0131  & n543 ;
  assign n1500 = ~n590 & ~n628 ;
  assign n1502 = n627 & ~n1500 ;
  assign n1501 = ~n627 & n1500 ;
  assign n1503 = ~n543 & ~n1501 ;
  assign n1504 = ~n1502 & n1503 ;
  assign n1505 = ~n1499 & ~n1504 ;
  assign n1506 = ~n538 & ~n1505 ;
  assign n1507 = \P1_IR_reg[31]/NET0131  & ~n467 ;
  assign n1508 = \P1_IR_reg[31]/NET0131  & \P1_IR_reg[6]/NET0131  ;
  assign n1509 = ~n1507 & ~n1508 ;
  assign n1510 = \P1_IR_reg[7]/NET0131  & ~n1509 ;
  assign n1511 = ~\P1_IR_reg[7]/NET0131  & n1509 ;
  assign n1512 = ~n1510 & ~n1511 ;
  assign n1513 = n538 & n1512 ;
  assign n1514 = ~n1506 & ~n1513 ;
  assign n1515 = n1498 & ~n1514 ;
  assign n1516 = \P1_reg0_reg[6]/NET0131  & n744 ;
  assign n1517 = ~\P1_reg3_reg[6]/NET0131  & ~n717 ;
  assign n1518 = ~n718 & ~n1517 ;
  assign n1519 = n715 & n1518 ;
  assign n1522 = ~n1516 & ~n1519 ;
  assign n1520 = \P1_reg1_reg[6]/NET0131  & n746 ;
  assign n1521 = \P1_reg2_reg[6]/NET0131  & n742 ;
  assign n1523 = ~n1520 & ~n1521 ;
  assign n1524 = n1522 & n1523 ;
  assign n1525 = \P2_datao_reg[6]/NET0131  & n543 ;
  assign n1526 = ~n602 & ~n604 ;
  assign n1528 = n787 & ~n1526 ;
  assign n1527 = ~n787 & n1526 ;
  assign n1529 = ~n543 & ~n1527 ;
  assign n1530 = ~n1528 & n1529 ;
  assign n1531 = ~n1525 & ~n1530 ;
  assign n1532 = ~n538 & ~n1531 ;
  assign n1533 = \P1_IR_reg[6]/NET0131  & ~n1507 ;
  assign n1534 = ~\P1_IR_reg[6]/NET0131  & n1507 ;
  assign n1535 = ~n1533 & ~n1534 ;
  assign n1536 = n538 & ~n1535 ;
  assign n1537 = ~n1532 & ~n1536 ;
  assign n1538 = n1524 & ~n1537 ;
  assign n1539 = ~n1515 & ~n1538 ;
  assign n1540 = \P1_reg0_reg[5]/NET0131  & n744 ;
  assign n1541 = \P1_reg1_reg[5]/NET0131  & n746 ;
  assign n1546 = ~n1540 & ~n1541 ;
  assign n1542 = ~\P1_reg3_reg[5]/NET0131  & ~n716 ;
  assign n1543 = ~n717 & ~n1542 ;
  assign n1544 = n715 & n1543 ;
  assign n1545 = \P1_reg2_reg[5]/NET0131  & n742 ;
  assign n1547 = ~n1544 & ~n1545 ;
  assign n1548 = n1546 & n1547 ;
  assign n1549 = \P2_datao_reg[5]/NET0131  & n543 ;
  assign n1550 = ~n603 & ~n622 ;
  assign n1552 = n854 & ~n1550 ;
  assign n1551 = ~n854 & n1550 ;
  assign n1553 = ~n543 & ~n1551 ;
  assign n1554 = ~n1552 & n1553 ;
  assign n1555 = ~n1549 & ~n1554 ;
  assign n1556 = ~n538 & ~n1555 ;
  assign n1557 = \P1_IR_reg[31]/NET0131  & ~n488 ;
  assign n1558 = ~\P1_IR_reg[5]/NET0131  & n1557 ;
  assign n1559 = \P1_IR_reg[5]/NET0131  & ~n1557 ;
  assign n1560 = ~n1558 & ~n1559 ;
  assign n1561 = n538 & ~n1560 ;
  assign n1562 = ~n1556 & ~n1561 ;
  assign n1563 = n1548 & ~n1562 ;
  assign n1564 = \P1_reg1_reg[4]/NET0131  & n746 ;
  assign n1565 = \P1_reg2_reg[4]/NET0131  & n742 ;
  assign n1570 = ~n1564 & ~n1565 ;
  assign n1566 = \P1_reg0_reg[4]/NET0131  & n744 ;
  assign n1567 = ~\P1_reg3_reg[3]/NET0131  & ~\P1_reg3_reg[4]/NET0131  ;
  assign n1568 = ~n716 & ~n1567 ;
  assign n1569 = n715 & n1568 ;
  assign n1571 = ~n1566 & ~n1569 ;
  assign n1572 = n1570 & n1571 ;
  assign n1573 = \P2_datao_reg[4]/NET0131  & n543 ;
  assign n1574 = ~n607 & ~n623 ;
  assign n1576 = n783 & ~n1574 ;
  assign n1575 = ~n783 & n1574 ;
  assign n1577 = ~n543 & ~n1575 ;
  assign n1578 = ~n1576 & n1577 ;
  assign n1579 = ~n1573 & ~n1578 ;
  assign n1580 = ~n538 & ~n1579 ;
  assign n1581 = \P1_IR_reg[31]/NET0131  & ~n487 ;
  assign n1582 = \P1_IR_reg[4]/NET0131  & ~n1581 ;
  assign n1583 = ~\P1_IR_reg[4]/NET0131  & n1581 ;
  assign n1584 = ~n1582 & ~n1583 ;
  assign n1585 = n538 & ~n1584 ;
  assign n1586 = ~n1580 & ~n1585 ;
  assign n1587 = n1572 & ~n1586 ;
  assign n1588 = ~n1563 & ~n1587 ;
  assign n1589 = \P1_reg0_reg[2]/NET0131  & n744 ;
  assign n1590 = \P1_reg1_reg[2]/NET0131  & n746 ;
  assign n1593 = ~n1589 & ~n1590 ;
  assign n1591 = \P1_reg2_reg[2]/NET0131  & n742 ;
  assign n1592 = \P1_reg3_reg[2]/NET0131  & n715 ;
  assign n1594 = ~n1591 & ~n1592 ;
  assign n1595 = n1593 & n1594 ;
  assign n1596 = \P2_datao_reg[2]/NET0131  & n543 ;
  assign n1597 = ~n610 & ~n616 ;
  assign n1599 = n779 & ~n1597 ;
  assign n1598 = ~n779 & n1597 ;
  assign n1600 = ~n543 & ~n1598 ;
  assign n1601 = ~n1599 & n1600 ;
  assign n1602 = ~n1596 & ~n1601 ;
  assign n1603 = ~n538 & ~n1602 ;
  assign n1604 = \P1_IR_reg[31]/NET0131  & ~n463 ;
  assign n1605 = \P1_IR_reg[2]/NET0131  & n1604 ;
  assign n1606 = ~\P1_IR_reg[2]/NET0131  & ~n1604 ;
  assign n1607 = ~n1605 & ~n1606 ;
  assign n1608 = n538 & n1607 ;
  assign n1609 = ~n1603 & ~n1608 ;
  assign n1610 = n1595 & ~n1609 ;
  assign n1611 = \P1_reg1_reg[3]/NET0131  & n746 ;
  assign n1612 = \P1_reg2_reg[3]/NET0131  & n742 ;
  assign n1615 = ~n1611 & ~n1612 ;
  assign n1613 = \P1_reg0_reg[3]/NET0131  & n744 ;
  assign n1614 = ~\P1_reg3_reg[3]/NET0131  & n715 ;
  assign n1616 = ~n1613 & ~n1614 ;
  assign n1617 = n1615 & n1616 ;
  assign n1618 = \P1_IR_reg[31]/NET0131  & ~n464 ;
  assign n1619 = \P1_IR_reg[3]/NET0131  & ~n1618 ;
  assign n1620 = ~\P1_IR_reg[3]/NET0131  & n1618 ;
  assign n1621 = ~n1619 & ~n1620 ;
  assign n1622 = n538 & ~n1621 ;
  assign n1623 = ~\P2_datao_reg[3]/NET0131  & n543 ;
  assign n1624 = ~n610 & ~n618 ;
  assign n1625 = ~n608 & ~n609 ;
  assign n1627 = ~n1624 & n1625 ;
  assign n1626 = n1624 & ~n1625 ;
  assign n1628 = ~n543 & ~n1626 ;
  assign n1629 = ~n1627 & n1628 ;
  assign n1630 = ~n1623 & ~n1629 ;
  assign n1631 = ~n538 & n1630 ;
  assign n1632 = ~n1622 & ~n1631 ;
  assign n1633 = n1617 & ~n1632 ;
  assign n1634 = ~n1610 & ~n1633 ;
  assign n1635 = \P1_reg1_reg[1]/NET0131  & n746 ;
  assign n1636 = \P1_reg0_reg[1]/NET0131  & n744 ;
  assign n1639 = ~n1635 & ~n1636 ;
  assign n1637 = \P1_reg3_reg[1]/NET0131  & n715 ;
  assign n1638 = \P1_reg2_reg[1]/NET0131  & n742 ;
  assign n1640 = ~n1637 & ~n1638 ;
  assign n1641 = n1639 & n1640 ;
  assign n1642 = \P1_IR_reg[0]/NET0131  & \P1_IR_reg[31]/NET0131  ;
  assign n1643 = ~\P1_IR_reg[1]/NET0131  & ~n1642 ;
  assign n1644 = \P1_IR_reg[1]/NET0131  & n1642 ;
  assign n1645 = ~n1643 & ~n1644 ;
  assign n1646 = n538 & n1645 ;
  assign n1647 = ~\P2_datao_reg[1]/NET0131  & n543 ;
  assign n1648 = ~n613 & ~n615 ;
  assign n1650 = n612 & ~n1648 ;
  assign n1649 = ~n612 & n1648 ;
  assign n1651 = ~n543 & ~n1649 ;
  assign n1652 = ~n1650 & n1651 ;
  assign n1653 = ~n1647 & ~n1652 ;
  assign n1654 = ~n538 & n1653 ;
  assign n1655 = ~n1646 & ~n1654 ;
  assign n1656 = ~n1641 & n1655 ;
  assign n1657 = n1641 & ~n1655 ;
  assign n1658 = \P1_reg3_reg[0]/NET0131  & n715 ;
  assign n1659 = \P1_reg2_reg[0]/NET0131  & n742 ;
  assign n1662 = ~n1658 & ~n1659 ;
  assign n1660 = \P1_reg0_reg[0]/NET0131  & n744 ;
  assign n1661 = \P1_reg1_reg[0]/NET0131  & n746 ;
  assign n1663 = ~n1660 & ~n1661 ;
  assign n1664 = n1662 & n1663 ;
  assign n1665 = \si[0]_pad  & ~n543 ;
  assign n1666 = ~\P2_datao_reg[0]/NET0131  & ~n1665 ;
  assign n1667 = ~n543 & n612 ;
  assign n1668 = ~n1666 & ~n1667 ;
  assign n1669 = ~n538 & n1668 ;
  assign n1670 = \P1_IR_reg[0]/NET0131  & n538 ;
  assign n1671 = ~n1669 & ~n1670 ;
  assign n1672 = n1664 & ~n1671 ;
  assign n1673 = ~n1657 & ~n1672 ;
  assign n1674 = ~n1656 & ~n1673 ;
  assign n1675 = n1634 & ~n1674 ;
  assign n1676 = ~n1617 & n1632 ;
  assign n1677 = ~n1595 & n1609 ;
  assign n1678 = ~n1676 & ~n1677 ;
  assign n1679 = ~n1633 & ~n1678 ;
  assign n1680 = ~n1675 & ~n1679 ;
  assign n1681 = n1588 & ~n1680 ;
  assign n1682 = ~n1548 & n1562 ;
  assign n1683 = ~n1572 & n1586 ;
  assign n1684 = ~n1563 & n1683 ;
  assign n1685 = ~n1682 & ~n1684 ;
  assign n1686 = ~n1681 & n1685 ;
  assign n1687 = n1539 & ~n1686 ;
  assign n1070 = \P1_IR_reg[31]/NET0131  & ~n503 ;
  assign n1071 = ~\P1_IR_reg[15]/NET0131  & ~n1070 ;
  assign n1072 = \P1_IR_reg[15]/NET0131  & n1070 ;
  assign n1073 = ~n1071 & ~n1072 ;
  assign n1074 = n538 & ~n1073 ;
  assign n1075 = \P2_datao_reg[15]/NET0131  & n543 ;
  assign n1076 = ~n569 & ~n639 ;
  assign n1078 = n638 & ~n1076 ;
  assign n1077 = ~n638 & n1076 ;
  assign n1079 = ~n543 & ~n1077 ;
  assign n1080 = ~n1078 & n1079 ;
  assign n1081 = ~n1075 & ~n1080 ;
  assign n1082 = ~n538 & n1081 ;
  assign n1083 = ~n1074 & ~n1082 ;
  assign n1084 = \P1_reg1_reg[15]/NET0131  & n746 ;
  assign n1087 = ~\P1_reg3_reg[15]/NET0131  & ~n1085 ;
  assign n1088 = ~n1086 & ~n1087 ;
  assign n1089 = n715 & n1088 ;
  assign n1092 = ~n1084 & ~n1089 ;
  assign n1090 = \P1_reg0_reg[15]/NET0131  & n744 ;
  assign n1091 = \P1_reg2_reg[15]/NET0131  & n742 ;
  assign n1093 = ~n1090 & ~n1091 ;
  assign n1094 = n1092 & n1093 ;
  assign n1095 = n1083 & n1094 ;
  assign n1096 = \P1_IR_reg[31]/NET0131  & ~n474 ;
  assign n1097 = \P1_IR_reg[14]/NET0131  & n1096 ;
  assign n1098 = ~\P1_IR_reg[14]/NET0131  & ~n1096 ;
  assign n1099 = ~n1097 & ~n1098 ;
  assign n1100 = n538 & ~n1099 ;
  assign n1101 = \P2_datao_reg[14]/NET0131  & n543 ;
  assign n1102 = ~n575 & ~n576 ;
  assign n1104 = n800 & ~n1102 ;
  assign n1103 = ~n800 & n1102 ;
  assign n1105 = ~n543 & ~n1103 ;
  assign n1106 = ~n1104 & n1105 ;
  assign n1107 = ~n1101 & ~n1106 ;
  assign n1108 = ~n538 & n1107 ;
  assign n1109 = ~n1100 & ~n1108 ;
  assign n1110 = \P1_reg0_reg[14]/NET0131  & n744 ;
  assign n1111 = \P1_reg1_reg[14]/NET0131  & n746 ;
  assign n1116 = ~n1110 & ~n1111 ;
  assign n1112 = ~\P1_reg3_reg[14]/NET0131  & ~n725 ;
  assign n1113 = ~n1085 & ~n1112 ;
  assign n1114 = n715 & n1113 ;
  assign n1115 = \P1_reg2_reg[14]/NET0131  & n742 ;
  assign n1117 = ~n1114 & ~n1115 ;
  assign n1118 = n1116 & n1117 ;
  assign n1119 = n1109 & n1118 ;
  assign n1120 = ~n1095 & ~n1119 ;
  assign n1121 = \P1_IR_reg[31]/NET0131  & ~n491 ;
  assign n1122 = \P1_IR_reg[31]/NET0131  & ~n471 ;
  assign n1123 = ~n1121 & ~n1122 ;
  assign n1124 = \P1_IR_reg[13]/NET0131  & ~n1123 ;
  assign n1125 = ~\P1_IR_reg[13]/NET0131  & n1123 ;
  assign n1126 = ~n1124 & ~n1125 ;
  assign n1127 = n538 & ~n1126 ;
  assign n1128 = \P2_datao_reg[13]/NET0131  & n543 ;
  assign n1129 = ~n577 & ~n580 ;
  assign n1131 = n865 & ~n1129 ;
  assign n1130 = ~n865 & n1129 ;
  assign n1132 = ~n543 & ~n1130 ;
  assign n1133 = ~n1131 & n1132 ;
  assign n1134 = ~n1128 & ~n1133 ;
  assign n1135 = ~n538 & n1134 ;
  assign n1136 = ~n1127 & ~n1135 ;
  assign n1137 = \P1_reg2_reg[13]/NET0131  & n742 ;
  assign n1138 = \P1_reg3_reg[12]/NET0131  & n723 ;
  assign n1139 = ~\P1_reg3_reg[13]/NET0131  & ~n1138 ;
  assign n1140 = ~n725 & ~n1139 ;
  assign n1141 = n715 & n1140 ;
  assign n1144 = ~n1137 & ~n1141 ;
  assign n1142 = \P1_reg0_reg[13]/NET0131  & n744 ;
  assign n1143 = \P1_reg1_reg[13]/NET0131  & n746 ;
  assign n1145 = ~n1142 & ~n1143 ;
  assign n1146 = n1144 & n1145 ;
  assign n1147 = n1136 & n1146 ;
  assign n1148 = ~n1136 & ~n1146 ;
  assign n1149 = n467 & n489 ;
  assign n1150 = n470 & n1149 ;
  assign n1151 = \P1_IR_reg[31]/NET0131  & ~n1150 ;
  assign n1152 = \P1_IR_reg[12]/NET0131  & n1151 ;
  assign n1153 = ~\P1_IR_reg[12]/NET0131  & ~n1151 ;
  assign n1154 = ~n1152 & ~n1153 ;
  assign n1155 = n538 & ~n1154 ;
  assign n1156 = \P2_datao_reg[12]/NET0131  & n543 ;
  assign n1157 = ~n582 & ~n583 ;
  assign n1158 = n897 & ~n908 ;
  assign n1160 = ~n1157 & n1158 ;
  assign n1159 = n1157 & ~n1158 ;
  assign n1161 = ~n543 & ~n1159 ;
  assign n1162 = ~n1160 & n1161 ;
  assign n1163 = ~n1156 & ~n1162 ;
  assign n1164 = ~n538 & n1163 ;
  assign n1165 = ~n1155 & ~n1164 ;
  assign n1166 = \P1_reg2_reg[12]/NET0131  & n742 ;
  assign n1167 = \P1_reg0_reg[12]/NET0131  & n744 ;
  assign n1172 = ~n1166 & ~n1167 ;
  assign n1168 = \P1_reg1_reg[12]/NET0131  & n746 ;
  assign n1169 = ~\P1_reg3_reg[12]/NET0131  & ~n723 ;
  assign n1170 = ~n1138 & ~n1169 ;
  assign n1171 = n715 & n1170 ;
  assign n1173 = ~n1168 & ~n1171 ;
  assign n1174 = n1172 & n1173 ;
  assign n1175 = ~n1165 & ~n1174 ;
  assign n1176 = ~n1148 & ~n1175 ;
  assign n1177 = ~n1147 & ~n1176 ;
  assign n1178 = n1120 & n1177 ;
  assign n1179 = ~n1109 & ~n1118 ;
  assign n1180 = ~n1083 & ~n1094 ;
  assign n1181 = ~n1179 & ~n1180 ;
  assign n1182 = ~n1095 & ~n1181 ;
  assign n1183 = ~n1178 & ~n1182 ;
  assign n1290 = n1165 & n1174 ;
  assign n1291 = ~n1147 & ~n1290 ;
  assign n1480 = n1120 & n1291 ;
  assign n1184 = n469 & n1149 ;
  assign n1185 = \P1_IR_reg[31]/NET0131  & ~n1184 ;
  assign n1186 = ~\P1_IR_reg[11]/NET0131  & ~n1185 ;
  assign n1187 = \P1_IR_reg[11]/NET0131  & n1185 ;
  assign n1188 = ~n1186 & ~n1187 ;
  assign n1189 = n538 & ~n1188 ;
  assign n1190 = \P2_datao_reg[11]/NET0131  & n543 ;
  assign n1191 = ~n584 & ~n634 ;
  assign n1193 = n633 & ~n1191 ;
  assign n1192 = ~n633 & n1191 ;
  assign n1194 = ~n543 & ~n1192 ;
  assign n1195 = ~n1193 & n1194 ;
  assign n1196 = ~n1190 & ~n1195 ;
  assign n1197 = ~n538 & n1196 ;
  assign n1198 = ~n1189 & ~n1197 ;
  assign n1199 = \P1_reg2_reg[11]/NET0131  & n742 ;
  assign n1200 = \P1_reg1_reg[11]/NET0131  & n746 ;
  assign n1205 = ~n1199 & ~n1200 ;
  assign n1201 = \P1_reg0_reg[11]/NET0131  & n744 ;
  assign n1202 = ~\P1_reg3_reg[11]/NET0131  & ~n722 ;
  assign n1203 = ~n723 & ~n1202 ;
  assign n1204 = n715 & n1203 ;
  assign n1206 = ~n1201 & ~n1204 ;
  assign n1207 = n1205 & n1206 ;
  assign n1209 = n1198 & n1207 ;
  assign n1210 = \P1_reg1_reg[10]/NET0131  & n746 ;
  assign n1211 = \P1_reg2_reg[10]/NET0131  & n742 ;
  assign n1216 = ~n1210 & ~n1211 ;
  assign n1212 = \P1_reg0_reg[10]/NET0131  & n744 ;
  assign n1213 = ~\P1_reg3_reg[10]/NET0131  & ~n721 ;
  assign n1214 = ~n722 & ~n1213 ;
  assign n1215 = n715 & n1214 ;
  assign n1217 = ~n1212 & ~n1215 ;
  assign n1218 = n1216 & n1217 ;
  assign n1219 = ~\P1_IR_reg[9]/NET0131  & n1149 ;
  assign n1220 = \P1_IR_reg[31]/NET0131  & ~n1219 ;
  assign n1221 = \P1_IR_reg[10]/NET0131  & n1220 ;
  assign n1222 = ~\P1_IR_reg[10]/NET0131  & ~n1220 ;
  assign n1223 = ~n1221 & ~n1222 ;
  assign n1224 = n538 & ~n1223 ;
  assign n1225 = \P2_datao_reg[10]/NET0131  & n543 ;
  assign n1226 = ~n593 & ~n599 ;
  assign n1228 = n796 & ~n1226 ;
  assign n1227 = ~n796 & n1226 ;
  assign n1229 = ~n543 & ~n1227 ;
  assign n1230 = ~n1228 & n1229 ;
  assign n1231 = ~n1225 & ~n1230 ;
  assign n1232 = ~n538 & n1231 ;
  assign n1233 = ~n1224 & ~n1232 ;
  assign n1234 = n1218 & n1233 ;
  assign n1235 = ~n1209 & ~n1234 ;
  assign n1236 = \P1_reg2_reg[9]/NET0131  & n742 ;
  assign n1237 = \P1_reg0_reg[9]/NET0131  & n744 ;
  assign n1242 = ~n1236 & ~n1237 ;
  assign n1238 = ~\P1_reg3_reg[9]/NET0131  & ~n720 ;
  assign n1239 = ~n721 & ~n1238 ;
  assign n1240 = n715 & n1239 ;
  assign n1241 = \P1_reg1_reg[9]/NET0131  & n746 ;
  assign n1243 = ~n1240 & ~n1241 ;
  assign n1244 = n1242 & n1243 ;
  assign n1245 = ~\P1_IR_reg[9]/NET0131  & ~n1121 ;
  assign n1246 = \P1_IR_reg[9]/NET0131  & n1121 ;
  assign n1247 = ~n1245 & ~n1246 ;
  assign n1248 = n538 & ~n1247 ;
  assign n1249 = \P2_datao_reg[9]/NET0131  & n543 ;
  assign n1250 = ~n592 & ~n598 ;
  assign n1252 = n860 & ~n1250 ;
  assign n1251 = ~n860 & n1250 ;
  assign n1253 = ~n543 & ~n1251 ;
  assign n1254 = ~n1252 & n1253 ;
  assign n1255 = ~n1249 & ~n1254 ;
  assign n1256 = ~n538 & n1255 ;
  assign n1257 = ~n1248 & ~n1256 ;
  assign n1258 = n1244 & n1257 ;
  assign n1284 = ~n1244 & ~n1257 ;
  assign n1259 = \P1_reg1_reg[8]/NET0131  & n746 ;
  assign n1260 = \P1_reg2_reg[8]/NET0131  & n742 ;
  assign n1265 = ~n1259 & ~n1260 ;
  assign n1261 = ~\P1_reg3_reg[8]/NET0131  & ~n719 ;
  assign n1262 = ~n720 & ~n1261 ;
  assign n1263 = n715 & n1262 ;
  assign n1264 = \P1_reg0_reg[8]/NET0131  & n744 ;
  assign n1266 = ~n1263 & ~n1264 ;
  assign n1267 = n1265 & n1266 ;
  assign n1268 = \P1_IR_reg[31]/NET0131  & ~n468 ;
  assign n1269 = ~\P1_IR_reg[8]/NET0131  & ~n1268 ;
  assign n1270 = \P1_IR_reg[8]/NET0131  & n1268 ;
  assign n1271 = ~n1269 & ~n1270 ;
  assign n1272 = n538 & ~n1271 ;
  assign n1273 = \P2_datao_reg[8]/NET0131  & n543 ;
  assign n1274 = ~n589 & ~n595 ;
  assign n1276 = n906 & ~n1274 ;
  assign n1275 = ~n906 & n1274 ;
  assign n1277 = ~n543 & ~n1275 ;
  assign n1278 = ~n1276 & n1277 ;
  assign n1279 = ~n1273 & ~n1278 ;
  assign n1280 = ~n538 & n1279 ;
  assign n1281 = ~n1272 & ~n1280 ;
  assign n1481 = ~n1267 & ~n1281 ;
  assign n1482 = ~n1284 & ~n1481 ;
  assign n1483 = ~n1258 & ~n1482 ;
  assign n1484 = n1235 & n1483 ;
  assign n1208 = ~n1198 & ~n1207 ;
  assign n1285 = ~n1218 & ~n1233 ;
  assign n1485 = ~n1208 & ~n1285 ;
  assign n1486 = ~n1209 & ~n1485 ;
  assign n1487 = ~n1484 & ~n1486 ;
  assign n1488 = n1480 & ~n1487 ;
  assign n1489 = n1183 & ~n1488 ;
  assign n1688 = ~n1498 & n1514 ;
  assign n1689 = ~n1524 & n1537 ;
  assign n1690 = ~n1515 & n1689 ;
  assign n1691 = ~n1688 & ~n1690 ;
  assign n1692 = n1489 & n1691 ;
  assign n1693 = ~n1687 & n1692 ;
  assign n1377 = n1338 & n1376 ;
  assign n1476 = n1466 & n1475 ;
  assign n1477 = ~n1453 & ~n1476 ;
  assign n1478 = n1429 & n1477 ;
  assign n1479 = n1377 & n1478 ;
  assign n1282 = n1267 & n1281 ;
  assign n1283 = ~n1258 & ~n1282 ;
  assign n1286 = ~n1284 & ~n1285 ;
  assign n1287 = ~n1283 & n1286 ;
  assign n1288 = n1235 & ~n1287 ;
  assign n1289 = ~n1208 & ~n1288 ;
  assign n1292 = ~n1148 & ~n1179 ;
  assign n1293 = ~n1291 & n1292 ;
  assign n1294 = n1120 & ~n1293 ;
  assign n1295 = ~n1180 & ~n1294 ;
  assign n1296 = ~n1289 & ~n1295 ;
  assign n1297 = n1183 & ~n1296 ;
  assign n1694 = ~n1297 & n1301 ;
  assign n1695 = n1479 & n1694 ;
  assign n1696 = ~n1693 & n1695 ;
  assign n1724 = ~n1069 & ~n1696 ;
  assign n1725 = ~n1723 & n1724 ;
  assign n1726 = n951 & ~n1725 ;
  assign n1727 = ~n949 & ~n1726 ;
  assign n835 = ~n692 & ~n750 ;
  assign n836 = ~n750 & ~n831 ;
  assign n837 = n825 & ~n836 ;
  assign n1728 = ~n835 & ~n837 ;
  assign n1729 = ~n1727 & n1728 ;
  assign n1730 = ~n834 & ~n1729 ;
  assign n1732 = n519 & ~n1730 ;
  assign n509 = \P1_IR_reg[31]/NET0131  & ~n508 ;
  assign n510 = ~\P1_IR_reg[23]/NET0131  & n509 ;
  assign n511 = \P1_IR_reg[23]/NET0131  & ~n509 ;
  assign n512 = ~n510 & ~n511 ;
  assign n513 = \P1_B_reg/NET0131  & ~n512 ;
  assign n1731 = ~n519 & n1730 ;
  assign n1733 = ~n513 & ~n1731 ;
  assign n1734 = ~n1732 & n1733 ;
  assign n483 = \P1_IR_reg[31]/NET0131  & ~n482 ;
  assign n484 = \P1_IR_reg[22]/NET0131  & n483 ;
  assign n485 = ~\P1_IR_reg[22]/NET0131  & ~n483 ;
  assign n486 = ~n484 & ~n485 ;
  assign n496 = ~\P1_IR_reg[20]/NET0131  & n477 ;
  assign n497 = n495 & n496 ;
  assign n498 = \P1_IR_reg[31]/NET0131  & ~n497 ;
  assign n499 = \P1_IR_reg[21]/NET0131  & n498 ;
  assign n500 = ~\P1_IR_reg[21]/NET0131  & ~n498 ;
  assign n501 = ~n499 & ~n500 ;
  assign n1735 = n486 & n501 ;
  assign n1736 = ~n1734 & n1735 ;
  assign n1737 = n692 & n750 ;
  assign n1738 = ~n832 & ~n1737 ;
  assign n1739 = n825 & n831 ;
  assign n1740 = n949 & ~n1739 ;
  assign n1741 = n1738 & ~n1740 ;
  assign n1742 = ~n835 & ~n1741 ;
  assign n1743 = n1539 & n1681 ;
  assign n1744 = n1539 & ~n1685 ;
  assign n1745 = n1691 & ~n1744 ;
  assign n1746 = ~n1743 & n1745 ;
  assign n1747 = n1235 & n1283 ;
  assign n1748 = ~n1746 & n1747 ;
  assign n1749 = n1480 & n1748 ;
  assign n1750 = n1489 & ~n1749 ;
  assign n1751 = n1479 & ~n1750 ;
  assign n1752 = n1377 & ~n1720 ;
  assign n1753 = n1710 & ~n1752 ;
  assign n1754 = ~n1751 & n1753 ;
  assign n1755 = n1301 & ~n1754 ;
  assign n1756 = ~n1069 & ~n1755 ;
  assign n1757 = ~n835 & ~n1739 ;
  assign n1758 = n951 & n1757 ;
  assign n1759 = ~n1756 & n1758 ;
  assign n1760 = ~n1742 & ~n1759 ;
  assign n1941 = ~\P1_B_reg/NET0131  & n1760 ;
  assign n1761 = ~n501 & n519 ;
  assign n1765 = ~n486 & ~n512 ;
  assign n1942 = n1761 & n1765 ;
  assign n1943 = ~n1941 & n1942 ;
  assign n1889 = ~n1007 & ~n1064 ;
  assign n1890 = ~n1300 & n1889 ;
  assign n1891 = n1298 & ~n1890 ;
  assign n1892 = ~n946 & ~n1008 ;
  assign n1893 = ~n1891 & n1892 ;
  assign n1894 = n951 & ~n1893 ;
  assign n1895 = ~n947 & ~n1894 ;
  assign n1896 = ~n1682 & ~n1689 ;
  assign n1897 = ~n1676 & ~n1683 ;
  assign n1803 = ~n1664 & n1671 ;
  assign n1898 = ~n1657 & n1803 ;
  assign n1899 = ~n1656 & ~n1677 ;
  assign n1900 = ~n1898 & n1899 ;
  assign n1901 = n1634 & ~n1900 ;
  assign n1902 = n1897 & ~n1901 ;
  assign n1903 = n1588 & ~n1902 ;
  assign n1904 = n1896 & ~n1903 ;
  assign n1905 = n1539 & ~n1904 ;
  assign n1906 = n1482 & ~n1688 ;
  assign n1907 = n1485 & n1906 ;
  assign n1908 = n1176 & n1907 ;
  assign n1909 = n1181 & n1908 ;
  assign n1910 = ~n1905 & n1909 ;
  assign n1911 = ~n1297 & ~n1910 ;
  assign n1912 = n1705 & n1708 ;
  assign n1913 = n1713 & n1718 ;
  assign n1914 = n1912 & n1913 ;
  assign n1915 = ~n1911 & n1914 ;
  assign n1916 = ~n1711 & ~n1717 ;
  assign n1917 = ~n1477 & n1916 ;
  assign n1918 = n1429 & ~n1917 ;
  assign n1919 = ~n1716 & ~n1918 ;
  assign n1920 = n1912 & n1919 ;
  assign n1921 = ~n1703 & ~n1920 ;
  assign n1922 = ~n1915 & n1921 ;
  assign n1923 = n1009 & n1065 ;
  assign n1924 = n948 & n1923 ;
  assign n1925 = ~n1922 & n1924 ;
  assign n1926 = ~n1895 & ~n1925 ;
  assign n1927 = ~n832 & ~n1926 ;
  assign n1928 = n1757 & ~n1927 ;
  assign n1929 = ~n1737 & ~n1928 ;
  assign n1934 = ~\P1_B_reg/NET0131  & ~n1929 ;
  assign n1885 = ~n501 & ~n519 ;
  assign n1935 = n486 & ~n512 ;
  assign n1936 = n1885 & n1935 ;
  assign n1937 = ~n1934 & n1936 ;
  assign n1938 = ~\P1_B_reg/NET0131  & n1929 ;
  assign n1939 = n1761 & n1935 ;
  assign n1940 = ~n1938 & n1939 ;
  assign n1948 = ~n1937 & ~n1940 ;
  assign n1949 = ~n1943 & n1948 ;
  assign n1931 = ~n1885 & n1929 ;
  assign n1888 = n486 & n512 ;
  assign n1930 = ~n1761 & ~n1929 ;
  assign n1932 = n1888 & ~n1930 ;
  assign n1933 = ~n1931 & n1932 ;
  assign n1886 = ~n486 & n1885 ;
  assign n1887 = n1760 & n1886 ;
  assign n1762 = ~n486 & n512 ;
  assign n1763 = n1761 & n1762 ;
  assign n1764 = ~n1760 & n1763 ;
  assign n1829 = ~n933 & n945 ;
  assign n1830 = n933 & ~n945 ;
  assign n1831 = ~n1829 & ~n1830 ;
  assign n1826 = ~n1365 & n1374 ;
  assign n1827 = n1365 & ~n1374 ;
  assign n1828 = ~n1826 & ~n1827 ;
  assign n1822 = ~n1394 & n1403 ;
  assign n1823 = n1394 & ~n1403 ;
  assign n1824 = ~n1822 & ~n1823 ;
  assign n1825 = ~n1453 & ~n1711 ;
  assign n1860 = ~n1824 & n1825 ;
  assign n1861 = ~n1828 & n1860 ;
  assign n1767 = ~n969 & n978 ;
  assign n1768 = n969 & ~n978 ;
  assign n1769 = ~n1767 & ~n1768 ;
  assign n1770 = ~n1198 & n1207 ;
  assign n1771 = n1198 & ~n1207 ;
  assign n1772 = ~n1770 & ~n1771 ;
  assign n1773 = ~n1633 & ~n1676 ;
  assign n1774 = n1498 & n1514 ;
  assign n1775 = ~n1498 & ~n1514 ;
  assign n1776 = ~n1774 & ~n1775 ;
  assign n1842 = n1773 & ~n1776 ;
  assign n1777 = ~n1595 & ~n1609 ;
  assign n1778 = n1595 & n1609 ;
  assign n1779 = ~n1777 & ~n1778 ;
  assign n1780 = ~n1244 & n1257 ;
  assign n1781 = n1244 & ~n1257 ;
  assign n1782 = ~n1780 & ~n1781 ;
  assign n1843 = ~n1779 & ~n1782 ;
  assign n1849 = n1842 & n1843 ;
  assign n1850 = ~n1772 & n1849 ;
  assign n1856 = ~n1769 & n1850 ;
  assign n1783 = ~n1466 & n1475 ;
  assign n1784 = n1466 & ~n1475 ;
  assign n1785 = ~n1783 & ~n1784 ;
  assign n1786 = ~n1083 & n1094 ;
  assign n1787 = n1083 & ~n1094 ;
  assign n1788 = ~n1786 & ~n1787 ;
  assign n1857 = ~n1785 & ~n1788 ;
  assign n1858 = n1856 & n1857 ;
  assign n1813 = ~n1109 & n1118 ;
  assign n1814 = n1109 & ~n1118 ;
  assign n1815 = ~n1813 & ~n1814 ;
  assign n1807 = n997 & ~n1006 ;
  assign n1808 = ~n997 & n1006 ;
  assign n1809 = ~n1807 & ~n1808 ;
  assign n1810 = ~n1029 & n1038 ;
  assign n1811 = n1029 & ~n1038 ;
  assign n1812 = ~n1810 & ~n1811 ;
  assign n1853 = ~n1809 & ~n1812 ;
  assign n1854 = ~n1815 & n1853 ;
  assign n1806 = ~n1587 & ~n1683 ;
  assign n1804 = ~n1672 & ~n1803 ;
  assign n1805 = ~n1563 & ~n1682 ;
  assign n1846 = n1804 & n1805 ;
  assign n1847 = n1806 & n1846 ;
  assign n1789 = ~n1218 & n1233 ;
  assign n1790 = n1218 & ~n1233 ;
  assign n1791 = ~n1789 & ~n1790 ;
  assign n1792 = ~n1656 & ~n1657 ;
  assign n1844 = ~n1791 & n1792 ;
  assign n1793 = ~n1538 & ~n1689 ;
  assign n1800 = n1267 & ~n1281 ;
  assign n1801 = ~n1267 & n1281 ;
  assign n1802 = ~n1800 & ~n1801 ;
  assign n1845 = n1793 & ~n1802 ;
  assign n1848 = n1844 & n1845 ;
  assign n1851 = n1847 & n1848 ;
  assign n1794 = ~n1165 & n1174 ;
  assign n1795 = n1165 & ~n1174 ;
  assign n1796 = ~n1794 & ~n1795 ;
  assign n1797 = ~n1136 & n1146 ;
  assign n1798 = n1136 & ~n1146 ;
  assign n1799 = ~n1797 & ~n1798 ;
  assign n1852 = ~n1796 & ~n1799 ;
  assign n1855 = n1851 & n1852 ;
  assign n1859 = n1854 & n1855 ;
  assign n1862 = n1858 & n1859 ;
  assign n1865 = n1861 & n1862 ;
  assign n1816 = ~n1047 & n1062 ;
  assign n1817 = n1047 & ~n1062 ;
  assign n1818 = ~n1816 & ~n1817 ;
  assign n1819 = n1327 & ~n1336 ;
  assign n1820 = ~n1327 & n1336 ;
  assign n1821 = ~n1819 & ~n1820 ;
  assign n1866 = ~n1818 & ~n1821 ;
  assign n1867 = n1865 & n1866 ;
  assign n1832 = ~n888 & ~n947 ;
  assign n1839 = ~n1346 & n1356 ;
  assign n1840 = n1346 & ~n1356 ;
  assign n1841 = ~n1839 & ~n1840 ;
  assign n1833 = ~n1418 & n1427 ;
  assign n1834 = n1418 & ~n1427 ;
  assign n1835 = ~n1833 & ~n1834 ;
  assign n1836 = ~n1309 & n1318 ;
  assign n1837 = n1309 & ~n1318 ;
  assign n1838 = ~n1836 & ~n1837 ;
  assign n1863 = ~n1835 & ~n1838 ;
  assign n1864 = ~n1841 & n1863 ;
  assign n1868 = n1832 & n1864 ;
  assign n1869 = n1867 & n1868 ;
  assign n1870 = ~n1831 & n1869 ;
  assign n1871 = n1738 & n1757 ;
  assign n1872 = n1870 & n1871 ;
  assign n1882 = n519 & n1872 ;
  assign n1880 = n501 & n1762 ;
  assign n1881 = ~n519 & ~n1872 ;
  assign n1883 = n1880 & ~n1881 ;
  assign n1884 = ~n1882 & n1883 ;
  assign n1766 = ~n519 & n1765 ;
  assign n1873 = n501 & n1872 ;
  assign n1874 = ~\P1_B_reg/NET0131  & ~n1873 ;
  assign n1875 = n1766 & ~n1874 ;
  assign n1876 = ~\P1_B_reg/NET0131  & n1872 ;
  assign n1877 = n519 & n1765 ;
  assign n1878 = n501 & n1877 ;
  assign n1879 = ~n1876 & n1878 ;
  assign n1944 = ~n1875 & ~n1879 ;
  assign n1945 = ~n1884 & n1944 ;
  assign n1946 = ~n1764 & n1945 ;
  assign n1947 = ~n1887 & n1946 ;
  assign n1950 = ~n1933 & n1947 ;
  assign n1951 = n1949 & n1950 ;
  assign n1952 = ~n1736 & n1951 ;
  assign n1953 = \P1_state_reg[0]/NET0131  & ~n512 ;
  assign n1954 = ~n1952 & n1953 ;
  assign n1955 = \P1_B_reg/NET0131  & ~n1953 ;
  assign n1956 = ~n1954 & ~n1955 ;
  assign n1961 = ~\P2_IR_reg[0]/NET0131  & ~\P2_IR_reg[1]/NET0131  ;
  assign n1962 = ~\P2_IR_reg[2]/NET0131  & n1961 ;
  assign n1963 = ~\P2_IR_reg[3]/NET0131  & ~\P2_IR_reg[4]/NET0131  ;
  assign n1964 = n1962 & n1963 ;
  assign n1965 = ~\P2_IR_reg[5]/NET0131  & ~\P2_IR_reg[6]/NET0131  ;
  assign n1966 = ~\P2_IR_reg[7]/NET0131  & n1965 ;
  assign n1967 = ~\P2_IR_reg[8]/NET0131  & ~\P2_IR_reg[9]/NET0131  ;
  assign n1968 = n1966 & n1967 ;
  assign n1969 = n1964 & n1968 ;
  assign n1959 = ~\P2_IR_reg[10]/NET0131  & ~\P2_IR_reg[11]/NET0131  ;
  assign n1960 = ~\P2_IR_reg[12]/NET0131  & n1959 ;
  assign n1970 = ~\P2_IR_reg[13]/NET0131  & n1960 ;
  assign n1971 = n1969 & n1970 ;
  assign n1972 = ~\P2_IR_reg[14]/NET0131  & n1971 ;
  assign n1973 = ~\P2_IR_reg[15]/NET0131  & n1972 ;
  assign n1974 = ~\P2_IR_reg[16]/NET0131  & ~\P2_IR_reg[17]/NET0131  ;
  assign n1975 = ~\P2_IR_reg[18]/NET0131  & n1974 ;
  assign n1976 = n1973 & n1975 ;
  assign n1957 = ~\P2_IR_reg[20]/NET0131  & ~\P2_IR_reg[21]/NET0131  ;
  assign n1958 = ~\P2_IR_reg[22]/NET0131  & n1957 ;
  assign n1977 = ~\P2_IR_reg[19]/NET0131  & n1958 ;
  assign n1978 = n1976 & n1977 ;
  assign n1979 = \P2_IR_reg[31]/NET0131  & ~n1978 ;
  assign n1980 = ~\P2_IR_reg[23]/NET0131  & ~n1979 ;
  assign n1981 = \P2_IR_reg[23]/NET0131  & n1979 ;
  assign n1982 = ~n1980 & ~n1981 ;
  assign n1983 = \P1_state_reg[0]/NET0131  & ~n1982 ;
  assign n1984 = \P2_reg0_reg[29]/NET0131  & ~n1983 ;
  assign n1987 = ~\P2_IR_reg[13]/NET0131  & ~\P2_IR_reg[14]/NET0131  ;
  assign n1988 = ~\P2_IR_reg[15]/NET0131  & ~\P2_IR_reg[16]/NET0131  ;
  assign n1989 = n1987 & n1988 ;
  assign n1990 = ~\P2_IR_reg[17]/NET0131  & n1989 ;
  assign n1991 = n1960 & n1990 ;
  assign n1992 = n1969 & n1991 ;
  assign n1993 = ~\P2_IR_reg[18]/NET0131  & ~\P2_IR_reg[19]/NET0131  ;
  assign n1994 = n1957 & n1993 ;
  assign n1995 = n1992 & n1994 ;
  assign n1985 = ~\P2_IR_reg[23]/NET0131  & ~\P2_IR_reg[24]/NET0131  ;
  assign n1986 = ~\P2_IR_reg[22]/NET0131  & n1985 ;
  assign n1996 = ~\P2_IR_reg[25]/NET0131  & n1986 ;
  assign n1997 = n1995 & n1996 ;
  assign n1998 = \P2_IR_reg[31]/NET0131  & ~n1997 ;
  assign n1999 = \P2_IR_reg[26]/NET0131  & n1998 ;
  assign n2000 = ~\P2_IR_reg[26]/NET0131  & ~n1998 ;
  assign n2001 = ~n1999 & ~n2000 ;
  assign n2002 = n1992 & n1993 ;
  assign n2003 = ~\P2_IR_reg[23]/NET0131  & n1958 ;
  assign n2004 = n2002 & n2003 ;
  assign n2005 = \P2_IR_reg[31]/NET0131  & ~n2004 ;
  assign n2006 = ~\P2_IR_reg[24]/NET0131  & ~n2005 ;
  assign n2007 = \P2_IR_reg[24]/NET0131  & n2005 ;
  assign n2008 = ~n2006 & ~n2007 ;
  assign n2009 = n2001 & n2008 ;
  assign n2010 = ~\P2_IR_reg[8]/NET0131  & n1966 ;
  assign n2011 = n1964 & n2010 ;
  assign n2012 = ~\P2_IR_reg[9]/NET0131  & n1960 ;
  assign n2013 = n2011 & n2012 ;
  assign n2014 = ~\P2_IR_reg[20]/NET0131  & n1993 ;
  assign n2015 = n1990 & n2014 ;
  assign n2016 = n2013 & n2015 ;
  assign n2017 = ~\P2_IR_reg[21]/NET0131  & n1986 ;
  assign n2018 = n2016 & n2017 ;
  assign n2019 = \P2_IR_reg[31]/NET0131  & ~n2018 ;
  assign n2020 = \P2_IR_reg[25]/NET0131  & n2019 ;
  assign n2021 = ~\P2_IR_reg[25]/NET0131  & ~n2019 ;
  assign n2022 = ~n2020 & ~n2021 ;
  assign n2023 = n2009 & n2022 ;
  assign n2024 = ~n1982 & n2023 ;
  assign n2025 = \P2_reg0_reg[29]/NET0131  & n2024 ;
  assign n2026 = ~n1982 & ~n2023 ;
  assign n2027 = \P2_B_reg/NET0131  & ~n2008 ;
  assign n2028 = ~n2022 & n2027 ;
  assign n2029 = ~\P2_d_reg[1]/NET0131  & ~n2028 ;
  assign n2030 = n2001 & ~n2029 ;
  assign n2031 = ~\P2_B_reg/NET0131  & ~n2022 ;
  assign n2032 = n2001 & ~n2031 ;
  assign n2033 = ~n2009 & ~n2022 ;
  assign n2034 = ~n2032 & ~n2033 ;
  assign n2035 = ~n2030 & ~n2034 ;
  assign n2036 = ~\P2_d_reg[0]/NET0131  & ~n2028 ;
  assign n2037 = n2001 & ~n2036 ;
  assign n2038 = n2008 & ~n2032 ;
  assign n2039 = ~n2037 & ~n2038 ;
  assign n2040 = n2035 & n2039 ;
  assign n2041 = \P2_reg0_reg[29]/NET0131  & ~n2040 ;
  assign n2042 = \P2_IR_reg[31]/NET0131  & ~n2002 ;
  assign n2043 = ~\P2_IR_reg[25]/NET0131  & ~\P2_IR_reg[26]/NET0131  ;
  assign n2044 = n1985 & n2043 ;
  assign n2045 = ~\P2_IR_reg[22]/NET0131  & n2044 ;
  assign n2046 = n1957 & n2045 ;
  assign n2047 = \P2_IR_reg[31]/NET0131  & ~n2046 ;
  assign n2048 = ~n2042 & ~n2047 ;
  assign n2049 = \P2_IR_reg[27]/NET0131  & ~n2048 ;
  assign n2050 = ~\P2_IR_reg[27]/NET0131  & n2048 ;
  assign n2051 = ~n2049 & ~n2050 ;
  assign n2052 = ~\P2_IR_reg[24]/NET0131  & ~\P2_IR_reg[27]/NET0131  ;
  assign n2053 = n2043 & n2052 ;
  assign n2054 = \P2_IR_reg[31]/NET0131  & ~n2053 ;
  assign n2055 = ~n2005 & ~n2054 ;
  assign n2056 = \P2_IR_reg[28]/NET0131  & ~n2055 ;
  assign n2057 = ~\P2_IR_reg[28]/NET0131  & n2055 ;
  assign n2058 = ~n2056 & ~n2057 ;
  assign n2059 = ~n2051 & ~n2058 ;
  assign n2060 = \P1_datao_reg[29]/NET0131  & ~n543 ;
  assign n2061 = \P1_datao_reg[29]/NET0131  & \si[29]_pad  ;
  assign n2062 = ~\P1_datao_reg[29]/NET0131  & ~\si[29]_pad  ;
  assign n2063 = ~n2061 & ~n2062 ;
  assign n2064 = ~\P1_datao_reg[28]/NET0131  & ~\si[28]_pad  ;
  assign n2119 = ~\P1_datao_reg[4]/NET0131  & ~\si[4]_pad  ;
  assign n2120 = ~\P1_datao_reg[3]/NET0131  & ~\si[3]_pad  ;
  assign n2121 = \P1_datao_reg[2]/NET0131  & \si[2]_pad  ;
  assign n2122 = ~\P1_datao_reg[2]/NET0131  & ~\si[2]_pad  ;
  assign n2123 = ~\P1_datao_reg[1]/NET0131  & ~\si[1]_pad  ;
  assign n2124 = \P1_datao_reg[1]/NET0131  & \si[1]_pad  ;
  assign n2125 = \P1_datao_reg[0]/NET0131  & \si[0]_pad  ;
  assign n2126 = ~n2124 & ~n2125 ;
  assign n2127 = ~n2123 & ~n2126 ;
  assign n2128 = ~n2122 & n2127 ;
  assign n2129 = ~n2121 & ~n2128 ;
  assign n2130 = ~n2120 & ~n2129 ;
  assign n2131 = \P1_datao_reg[4]/NET0131  & \si[4]_pad  ;
  assign n2132 = \P1_datao_reg[3]/NET0131  & \si[3]_pad  ;
  assign n2133 = ~n2131 & ~n2132 ;
  assign n2134 = ~n2130 & n2133 ;
  assign n2135 = ~n2119 & ~n2134 ;
  assign n2108 = ~\P1_datao_reg[7]/NET0131  & ~\si[7]_pad  ;
  assign n2109 = ~\P1_datao_reg[8]/NET0131  & ~\si[8]_pad  ;
  assign n2110 = ~n2108 & ~n2109 ;
  assign n2112 = ~\P1_datao_reg[6]/NET0131  & ~\si[6]_pad  ;
  assign n2136 = ~\P1_datao_reg[5]/NET0131  & ~\si[5]_pad  ;
  assign n2137 = ~n2112 & ~n2136 ;
  assign n2138 = n2110 & n2137 ;
  assign n2139 = n2135 & n2138 ;
  assign n2107 = \P1_datao_reg[8]/NET0131  & \si[8]_pad  ;
  assign n2111 = \P1_datao_reg[7]/NET0131  & \si[7]_pad  ;
  assign n2113 = \P1_datao_reg[5]/NET0131  & \si[5]_pad  ;
  assign n2114 = \P1_datao_reg[6]/NET0131  & \si[6]_pad  ;
  assign n2115 = ~n2113 & ~n2114 ;
  assign n2116 = ~n2112 & ~n2115 ;
  assign n2117 = ~n2111 & ~n2116 ;
  assign n2118 = n2110 & ~n2117 ;
  assign n2140 = ~n2107 & ~n2118 ;
  assign n2141 = ~n2139 & n2140 ;
  assign n2143 = ~\P1_datao_reg[11]/NET0131  & ~\si[11]_pad  ;
  assign n2144 = ~\P1_datao_reg[10]/NET0131  & ~\si[10]_pad  ;
  assign n2145 = ~n2143 & ~n2144 ;
  assign n2142 = ~\P1_datao_reg[12]/NET0131  & ~\si[12]_pad  ;
  assign n2146 = ~\P1_datao_reg[9]/NET0131  & ~\si[9]_pad  ;
  assign n2147 = ~n2142 & ~n2146 ;
  assign n2148 = n2145 & n2147 ;
  assign n2149 = ~n2141 & n2148 ;
  assign n2150 = \P1_datao_reg[12]/NET0131  & \si[12]_pad  ;
  assign n2151 = \P1_datao_reg[11]/NET0131  & \si[11]_pad  ;
  assign n2152 = \P1_datao_reg[10]/NET0131  & \si[10]_pad  ;
  assign n2153 = \P1_datao_reg[9]/NET0131  & \si[9]_pad  ;
  assign n2154 = ~n2152 & ~n2153 ;
  assign n2155 = ~n2144 & ~n2154 ;
  assign n2156 = ~n2151 & ~n2155 ;
  assign n2157 = ~n2142 & ~n2143 ;
  assign n2158 = ~n2156 & n2157 ;
  assign n2159 = ~n2150 & ~n2158 ;
  assign n2160 = ~n2149 & n2159 ;
  assign n2077 = ~\P1_datao_reg[17]/NET0131  & ~\si[17]_pad  ;
  assign n2078 = ~\P1_datao_reg[20]/NET0131  & ~\si[20]_pad  ;
  assign n2079 = ~\P1_datao_reg[18]/NET0131  & ~\si[18]_pad  ;
  assign n2080 = ~\P1_datao_reg[19]/NET0131  & ~\si[19]_pad  ;
  assign n2081 = ~n2079 & ~n2080 ;
  assign n2082 = ~n2078 & n2081 ;
  assign n2083 = ~n2077 & n2082 ;
  assign n2088 = ~\P1_datao_reg[14]/NET0131  & ~\si[14]_pad  ;
  assign n2089 = ~\P1_datao_reg[15]/NET0131  & ~\si[15]_pad  ;
  assign n2090 = ~n2088 & ~n2089 ;
  assign n2084 = ~\P1_datao_reg[16]/NET0131  & ~\si[16]_pad  ;
  assign n2161 = ~\P1_datao_reg[13]/NET0131  & ~\si[13]_pad  ;
  assign n2162 = ~n2084 & ~n2161 ;
  assign n2163 = n2090 & n2162 ;
  assign n2164 = n2083 & n2163 ;
  assign n2165 = ~n2160 & n2164 ;
  assign n2085 = \P1_datao_reg[15]/NET0131  & \si[15]_pad  ;
  assign n2086 = \P1_datao_reg[16]/NET0131  & \si[16]_pad  ;
  assign n2087 = ~n2085 & ~n2086 ;
  assign n2091 = \P1_datao_reg[13]/NET0131  & \si[13]_pad  ;
  assign n2092 = \P1_datao_reg[14]/NET0131  & \si[14]_pad  ;
  assign n2093 = ~n2091 & ~n2092 ;
  assign n2094 = n2090 & ~n2093 ;
  assign n2095 = n2087 & ~n2094 ;
  assign n2096 = ~n2084 & ~n2095 ;
  assign n2097 = n2083 & n2096 ;
  assign n2098 = \P1_datao_reg[19]/NET0131  & \si[19]_pad  ;
  assign n2099 = \P1_datao_reg[20]/NET0131  & \si[20]_pad  ;
  assign n2100 = ~n2098 & ~n2099 ;
  assign n2101 = ~n2078 & ~n2100 ;
  assign n2102 = \P1_datao_reg[17]/NET0131  & \si[17]_pad  ;
  assign n2103 = \P1_datao_reg[18]/NET0131  & \si[18]_pad  ;
  assign n2104 = ~n2102 & ~n2103 ;
  assign n2105 = n2082 & ~n2104 ;
  assign n2106 = ~n2101 & ~n2105 ;
  assign n2166 = ~n2097 & n2106 ;
  assign n2167 = ~n2165 & n2166 ;
  assign n2065 = ~\P1_datao_reg[23]/NET0131  & ~\si[23]_pad  ;
  assign n2066 = ~\P1_datao_reg[24]/NET0131  & ~\si[24]_pad  ;
  assign n2067 = ~n2065 & ~n2066 ;
  assign n2068 = ~\P1_datao_reg[22]/NET0131  & ~\si[22]_pad  ;
  assign n2069 = ~\P1_datao_reg[21]/NET0131  & ~\si[21]_pad  ;
  assign n2070 = ~n2068 & ~n2069 ;
  assign n2071 = n2067 & n2070 ;
  assign n2072 = ~\P1_datao_reg[27]/NET0131  & ~\si[27]_pad  ;
  assign n2073 = ~\P1_datao_reg[26]/NET0131  & ~\si[26]_pad  ;
  assign n2074 = ~\P1_datao_reg[25]/NET0131  & ~\si[25]_pad  ;
  assign n2075 = ~n2073 & ~n2074 ;
  assign n2076 = ~n2072 & n2075 ;
  assign n2168 = n2071 & n2076 ;
  assign n2169 = ~n2167 & n2168 ;
  assign n2170 = \P1_datao_reg[27]/NET0131  & \si[27]_pad  ;
  assign n2171 = \P1_datao_reg[28]/NET0131  & \si[28]_pad  ;
  assign n2172 = ~n2170 & ~n2171 ;
  assign n2173 = \P1_datao_reg[26]/NET0131  & \si[26]_pad  ;
  assign n2174 = \P1_datao_reg[25]/NET0131  & \si[25]_pad  ;
  assign n2175 = ~n2173 & ~n2174 ;
  assign n2176 = ~n2073 & ~n2175 ;
  assign n2177 = \P1_datao_reg[22]/NET0131  & \si[22]_pad  ;
  assign n2178 = \P1_datao_reg[21]/NET0131  & \si[21]_pad  ;
  assign n2179 = ~n2177 & ~n2178 ;
  assign n2180 = ~n2068 & ~n2179 ;
  assign n2181 = n2067 & n2180 ;
  assign n2182 = \P1_datao_reg[23]/NET0131  & \si[23]_pad  ;
  assign n2183 = \P1_datao_reg[24]/NET0131  & \si[24]_pad  ;
  assign n2184 = ~n2182 & ~n2183 ;
  assign n2185 = ~n2066 & ~n2184 ;
  assign n2186 = ~n2181 & ~n2185 ;
  assign n2187 = n2075 & ~n2186 ;
  assign n2188 = ~n2176 & ~n2187 ;
  assign n2189 = ~n2072 & ~n2188 ;
  assign n2190 = n2172 & ~n2189 ;
  assign n2191 = ~n2169 & n2190 ;
  assign n2192 = ~n2064 & ~n2191 ;
  assign n2194 = n2063 & n2192 ;
  assign n2193 = ~n2063 & ~n2192 ;
  assign n2195 = n543 & ~n2193 ;
  assign n2196 = ~n2194 & n2195 ;
  assign n2197 = ~n2060 & ~n2196 ;
  assign n2198 = ~n2059 & ~n2197 ;
  assign n2199 = \P2_IR_reg[31]/NET0131  & ~n1995 ;
  assign n2200 = ~\P2_IR_reg[27]/NET0131  & ~\P2_IR_reg[28]/NET0131  ;
  assign n2201 = ~\P2_IR_reg[29]/NET0131  & n2200 ;
  assign n2202 = n2045 & n2201 ;
  assign n2203 = \P2_IR_reg[31]/NET0131  & ~n2202 ;
  assign n2204 = ~n2199 & ~n2203 ;
  assign n2205 = \P2_IR_reg[30]/NET0131  & ~n2204 ;
  assign n2206 = ~\P2_IR_reg[30]/NET0131  & n2204 ;
  assign n2207 = ~n2205 & ~n2206 ;
  assign n2208 = \P2_IR_reg[31]/NET0131  & ~n2016 ;
  assign n2209 = ~\P2_IR_reg[21]/NET0131  & n2200 ;
  assign n2210 = n2045 & n2209 ;
  assign n2211 = \P2_IR_reg[31]/NET0131  & ~n2210 ;
  assign n2212 = ~n2208 & ~n2211 ;
  assign n2213 = \P2_IR_reg[29]/NET0131  & ~n2212 ;
  assign n2214 = ~\P2_IR_reg[29]/NET0131  & n2212 ;
  assign n2215 = ~n2213 & ~n2214 ;
  assign n2216 = n2207 & n2215 ;
  assign n2217 = \P2_reg3_reg[3]/NET0131  & \P2_reg3_reg[4]/NET0131  ;
  assign n2218 = \P2_reg3_reg[5]/NET0131  & n2217 ;
  assign n2219 = \P2_reg3_reg[6]/NET0131  & n2218 ;
  assign n2220 = \P2_reg3_reg[7]/NET0131  & n2219 ;
  assign n2221 = \P2_reg3_reg[8]/NET0131  & n2220 ;
  assign n2222 = \P2_reg3_reg[9]/NET0131  & n2221 ;
  assign n2223 = \P2_reg3_reg[10]/NET0131  & n2222 ;
  assign n2224 = \P2_reg3_reg[11]/NET0131  & \P2_reg3_reg[12]/NET0131  ;
  assign n2225 = \P2_reg3_reg[13]/NET0131  & \P2_reg3_reg[14]/NET0131  ;
  assign n2226 = n2224 & n2225 ;
  assign n2227 = n2223 & n2226 ;
  assign n2228 = \P2_reg3_reg[15]/NET0131  & \P2_reg3_reg[16]/NET0131  ;
  assign n2229 = n2227 & n2228 ;
  assign n2230 = \P2_reg3_reg[20]/NET0131  & \P2_reg3_reg[21]/NET0131  ;
  assign n2231 = \P2_reg3_reg[22]/NET0131  & n2230 ;
  assign n2232 = \P2_reg3_reg[17]/NET0131  & \P2_reg3_reg[18]/NET0131  ;
  assign n2233 = \P2_reg3_reg[19]/NET0131  & \P2_reg3_reg[23]/NET0131  ;
  assign n2234 = \P2_reg3_reg[24]/NET0131  & n2233 ;
  assign n2235 = n2232 & n2234 ;
  assign n2236 = n2231 & n2235 ;
  assign n2237 = n2229 & n2236 ;
  assign n2238 = \P2_reg3_reg[25]/NET0131  & \P2_reg3_reg[26]/NET0131  ;
  assign n2239 = \P2_reg3_reg[27]/NET0131  & \P2_reg3_reg[28]/NET0131  ;
  assign n2240 = n2238 & n2239 ;
  assign n2241 = n2237 & n2240 ;
  assign n2242 = n2216 & n2241 ;
  assign n2243 = n2207 & ~n2215 ;
  assign n2244 = \P2_reg2_reg[29]/NET0131  & n2243 ;
  assign n2249 = ~n2242 & ~n2244 ;
  assign n2245 = ~n2207 & ~n2215 ;
  assign n2246 = \P2_reg0_reg[29]/NET0131  & n2245 ;
  assign n2247 = ~n2207 & n2215 ;
  assign n2248 = \P2_reg1_reg[29]/NET0131  & n2247 ;
  assign n2250 = ~n2246 & ~n2248 ;
  assign n2251 = n2249 & n2250 ;
  assign n2252 = n2198 & n2251 ;
  assign n2253 = ~n2198 & ~n2251 ;
  assign n2254 = ~n2252 & ~n2253 ;
  assign n2255 = \P2_IR_reg[31]/NET0131  & ~n1976 ;
  assign n2256 = ~\P2_IR_reg[19]/NET0131  & ~n2255 ;
  assign n2257 = \P2_IR_reg[19]/NET0131  & n2255 ;
  assign n2258 = ~n2256 & ~n2257 ;
  assign n2259 = n2059 & ~n2258 ;
  assign n2260 = \P1_datao_reg[19]/NET0131  & ~n543 ;
  assign n2261 = ~n2077 & ~n2084 ;
  assign n2262 = ~n2079 & n2261 ;
  assign n2263 = ~n2089 & n2262 ;
  assign n2264 = ~n2119 & ~n2136 ;
  assign n2265 = ~n2112 & n2264 ;
  assign n2266 = ~n2134 & n2265 ;
  assign n2267 = ~n2116 & ~n2266 ;
  assign n2268 = ~n2109 & ~n2146 ;
  assign n2269 = ~n2108 & n2268 ;
  assign n2270 = ~n2144 & n2269 ;
  assign n2271 = ~n2267 & n2270 ;
  assign n2272 = ~n2107 & ~n2111 ;
  assign n2273 = ~n2144 & n2268 ;
  assign n2274 = ~n2272 & n2273 ;
  assign n2275 = ~n2155 & ~n2274 ;
  assign n2276 = ~n2271 & n2275 ;
  assign n2277 = n2157 & ~n2161 ;
  assign n2278 = ~n2088 & n2277 ;
  assign n2279 = ~n2276 & n2278 ;
  assign n2280 = n2263 & n2279 ;
  assign n2281 = ~n2142 & ~n2161 ;
  assign n2282 = ~n2150 & ~n2151 ;
  assign n2283 = n2281 & ~n2282 ;
  assign n2284 = n2093 & ~n2283 ;
  assign n2285 = ~n2088 & ~n2284 ;
  assign n2286 = n2263 & n2285 ;
  assign n2287 = ~n2087 & n2261 ;
  assign n2288 = n2104 & ~n2287 ;
  assign n2289 = ~n2079 & ~n2288 ;
  assign n2290 = ~n2286 & ~n2289 ;
  assign n2291 = ~n2280 & n2290 ;
  assign n2292 = ~n2080 & ~n2098 ;
  assign n2294 = ~n2291 & n2292 ;
  assign n2293 = n2291 & ~n2292 ;
  assign n2295 = n543 & ~n2293 ;
  assign n2296 = ~n2294 & n2295 ;
  assign n2297 = ~n2260 & ~n2296 ;
  assign n2298 = ~n2059 & n2297 ;
  assign n2299 = ~n2259 & ~n2298 ;
  assign n2303 = \P2_reg3_reg[17]/NET0131  & n2229 ;
  assign n2304 = \P2_reg3_reg[18]/NET0131  & n2303 ;
  assign n2305 = ~\P2_reg3_reg[19]/NET0131  & ~n2304 ;
  assign n2306 = \P2_reg3_reg[19]/NET0131  & n2304 ;
  assign n2307 = ~n2305 & ~n2306 ;
  assign n2308 = n2216 & n2307 ;
  assign n2302 = \P2_reg1_reg[19]/NET0131  & n2247 ;
  assign n2300 = \P2_reg0_reg[19]/NET0131  & n2245 ;
  assign n2301 = \P2_reg2_reg[19]/NET0131  & n2243 ;
  assign n2309 = ~n2300 & ~n2301 ;
  assign n2310 = ~n2302 & n2309 ;
  assign n2311 = ~n2308 & n2310 ;
  assign n2312 = ~n2299 & n2311 ;
  assign n2313 = \P1_datao_reg[20]/NET0131  & ~n543 ;
  assign n2319 = n2090 & n2281 ;
  assign n2320 = ~n2121 & ~n2132 ;
  assign n2321 = ~n2128 & n2320 ;
  assign n2322 = ~n2120 & ~n2321 ;
  assign n2323 = n2265 & n2322 ;
  assign n2324 = ~n2111 & ~n2114 ;
  assign n2325 = ~n2113 & ~n2131 ;
  assign n2326 = ~n2136 & ~n2325 ;
  assign n2327 = ~n2112 & n2326 ;
  assign n2328 = n2324 & ~n2327 ;
  assign n2329 = ~n2323 & n2328 ;
  assign n2330 = ~n2108 & ~n2329 ;
  assign n2331 = n2145 & n2268 ;
  assign n2332 = n2330 & n2331 ;
  assign n2333 = n2319 & n2332 ;
  assign n2337 = ~n2107 & ~n2153 ;
  assign n2338 = ~n2146 & ~n2337 ;
  assign n2339 = ~n2152 & ~n2338 ;
  assign n2340 = n2145 & ~n2339 ;
  assign n2341 = ~n2151 & ~n2340 ;
  assign n2342 = n2319 & ~n2341 ;
  assign n2334 = ~n2091 & ~n2150 ;
  assign n2335 = ~n2161 & ~n2334 ;
  assign n2336 = n2090 & n2335 ;
  assign n2343 = ~n2085 & ~n2092 ;
  assign n2344 = ~n2089 & ~n2343 ;
  assign n2345 = ~n2336 & ~n2344 ;
  assign n2346 = ~n2342 & n2345 ;
  assign n2347 = ~n2333 & n2346 ;
  assign n2348 = ~n2080 & n2262 ;
  assign n2349 = ~n2347 & n2348 ;
  assign n2314 = ~n2098 & ~n2103 ;
  assign n2315 = ~n2080 & ~n2314 ;
  assign n2316 = ~n2086 & ~n2102 ;
  assign n2317 = ~n2077 & ~n2316 ;
  assign n2318 = n2081 & n2317 ;
  assign n2350 = ~n2315 & ~n2318 ;
  assign n2351 = ~n2349 & n2350 ;
  assign n2352 = ~n2078 & ~n2099 ;
  assign n2354 = ~n2351 & n2352 ;
  assign n2353 = n2351 & ~n2352 ;
  assign n2355 = n543 & ~n2353 ;
  assign n2356 = ~n2354 & n2355 ;
  assign n2357 = ~n2313 & ~n2356 ;
  assign n2358 = ~n2059 & ~n2357 ;
  assign n2362 = \P2_reg3_reg[20]/NET0131  & n2306 ;
  assign n2363 = ~\P2_reg3_reg[20]/NET0131  & ~n2306 ;
  assign n2364 = ~n2362 & ~n2363 ;
  assign n2365 = n2216 & n2364 ;
  assign n2361 = \P2_reg2_reg[20]/NET0131  & n2243 ;
  assign n2359 = \P2_reg1_reg[20]/NET0131  & n2247 ;
  assign n2360 = \P2_reg0_reg[20]/NET0131  & n2245 ;
  assign n2366 = ~n2359 & ~n2360 ;
  assign n2367 = ~n2361 & n2366 ;
  assign n2368 = ~n2365 & n2367 ;
  assign n2369 = ~n2358 & n2368 ;
  assign n2370 = ~n2312 & ~n2369 ;
  assign n2371 = \P2_reg1_reg[17]/NET0131  & n2247 ;
  assign n2372 = ~\P2_reg3_reg[17]/NET0131  & ~n2229 ;
  assign n2373 = ~n2303 & ~n2372 ;
  assign n2374 = n2216 & n2373 ;
  assign n2377 = ~n2371 & ~n2374 ;
  assign n2375 = \P2_reg2_reg[17]/NET0131  & n2243 ;
  assign n2376 = \P2_reg0_reg[17]/NET0131  & n2245 ;
  assign n2378 = ~n2375 & ~n2376 ;
  assign n2379 = n2377 & n2378 ;
  assign n2380 = \P2_IR_reg[31]/NET0131  & ~n2013 ;
  assign n2381 = \P2_IR_reg[31]/NET0131  & ~n1989 ;
  assign n2382 = ~n2380 & ~n2381 ;
  assign n2383 = \P2_IR_reg[17]/NET0131  & ~n2382 ;
  assign n2384 = ~\P2_IR_reg[17]/NET0131  & n2382 ;
  assign n2385 = ~n2383 & ~n2384 ;
  assign n2386 = n2059 & ~n2385 ;
  assign n2387 = \P1_datao_reg[17]/NET0131  & ~n543 ;
  assign n2388 = n2149 & n2163 ;
  assign n2389 = ~n2159 & n2163 ;
  assign n2390 = ~n2096 & ~n2389 ;
  assign n2391 = ~n2388 & n2390 ;
  assign n2392 = ~n2077 & ~n2102 ;
  assign n2394 = ~n2391 & n2392 ;
  assign n2393 = n2391 & ~n2392 ;
  assign n2395 = n543 & ~n2393 ;
  assign n2396 = ~n2394 & n2395 ;
  assign n2397 = ~n2387 & ~n2396 ;
  assign n2398 = ~n2059 & n2397 ;
  assign n2399 = ~n2386 & ~n2398 ;
  assign n2400 = n2379 & ~n2399 ;
  assign n2401 = \P2_IR_reg[31]/NET0131  & ~n1992 ;
  assign n2402 = ~\P2_IR_reg[18]/NET0131  & ~n2401 ;
  assign n2403 = \P2_IR_reg[18]/NET0131  & n2401 ;
  assign n2404 = ~n2402 & ~n2403 ;
  assign n2405 = n2059 & ~n2404 ;
  assign n2406 = \P1_datao_reg[18]/NET0131  & ~n543 ;
  assign n2407 = ~n2079 & ~n2103 ;
  assign n2408 = n2264 & n2322 ;
  assign n2409 = ~n2326 & ~n2408 ;
  assign n2410 = ~n2112 & n2269 ;
  assign n2411 = ~n2409 & n2410 ;
  assign n2412 = n2269 & ~n2324 ;
  assign n2413 = ~n2338 & ~n2412 ;
  assign n2414 = ~n2411 & n2413 ;
  assign n2415 = ~n2144 & n2277 ;
  assign n2416 = ~n2414 & n2415 ;
  assign n2417 = n2090 & n2261 ;
  assign n2418 = n2416 & n2417 ;
  assign n2419 = n2261 & n2344 ;
  assign n2420 = ~n2317 & ~n2419 ;
  assign n2421 = ~n2151 & ~n2152 ;
  assign n2422 = n2277 & ~n2421 ;
  assign n2423 = ~n2335 & ~n2422 ;
  assign n2424 = n2417 & ~n2423 ;
  assign n2425 = n2420 & ~n2424 ;
  assign n2426 = ~n2418 & n2425 ;
  assign n2428 = ~n2407 & n2426 ;
  assign n2427 = n2407 & ~n2426 ;
  assign n2429 = n543 & ~n2427 ;
  assign n2430 = ~n2428 & n2429 ;
  assign n2431 = ~n2406 & ~n2430 ;
  assign n2432 = ~n2059 & n2431 ;
  assign n2433 = ~n2405 & ~n2432 ;
  assign n2437 = ~\P2_reg3_reg[18]/NET0131  & ~n2303 ;
  assign n2438 = ~n2304 & ~n2437 ;
  assign n2439 = n2216 & n2438 ;
  assign n2436 = \P2_reg1_reg[18]/NET0131  & n2247 ;
  assign n2434 = \P2_reg2_reg[18]/NET0131  & n2243 ;
  assign n2435 = \P2_reg0_reg[18]/NET0131  & n2245 ;
  assign n2440 = ~n2434 & ~n2435 ;
  assign n2441 = ~n2436 & n2440 ;
  assign n2442 = ~n2439 & n2441 ;
  assign n2443 = ~n2433 & n2442 ;
  assign n2444 = ~n2400 & ~n2443 ;
  assign n2445 = n2370 & n2444 ;
  assign n2446 = ~\P2_reg3_reg[8]/NET0131  & ~n2220 ;
  assign n2447 = ~n2221 & ~n2446 ;
  assign n2448 = n2216 & n2447 ;
  assign n2449 = \P2_reg1_reg[8]/NET0131  & n2247 ;
  assign n2452 = ~n2448 & ~n2449 ;
  assign n2450 = \P2_reg0_reg[8]/NET0131  & n2245 ;
  assign n2451 = \P2_reg2_reg[8]/NET0131  & n2243 ;
  assign n2453 = ~n2450 & ~n2451 ;
  assign n2454 = n2452 & n2453 ;
  assign n2455 = \P2_IR_reg[31]/NET0131  & ~n1964 ;
  assign n2456 = \P2_IR_reg[31]/NET0131  & ~n1966 ;
  assign n2457 = ~n2455 & ~n2456 ;
  assign n2458 = \P2_IR_reg[8]/NET0131  & ~n2457 ;
  assign n2459 = ~\P2_IR_reg[8]/NET0131  & n2457 ;
  assign n2460 = ~n2458 & ~n2459 ;
  assign n2461 = n2059 & ~n2460 ;
  assign n2462 = \P1_datao_reg[8]/NET0131  & ~n543 ;
  assign n2463 = ~n2107 & ~n2109 ;
  assign n2465 = n2330 & n2463 ;
  assign n2464 = ~n2330 & ~n2463 ;
  assign n2466 = n543 & ~n2464 ;
  assign n2467 = ~n2465 & n2466 ;
  assign n2468 = ~n2462 & ~n2467 ;
  assign n2469 = ~n2059 & n2468 ;
  assign n2470 = ~n2461 & ~n2469 ;
  assign n2471 = n2454 & ~n2470 ;
  assign n2472 = \P2_reg2_reg[7]/NET0131  & n2243 ;
  assign n2473 = \P2_reg1_reg[7]/NET0131  & n2247 ;
  assign n2478 = ~n2472 & ~n2473 ;
  assign n2474 = \P2_reg0_reg[7]/NET0131  & n2245 ;
  assign n2475 = ~\P2_reg3_reg[7]/NET0131  & ~n2219 ;
  assign n2476 = ~n2220 & ~n2475 ;
  assign n2477 = n2216 & n2476 ;
  assign n2479 = ~n2474 & ~n2477 ;
  assign n2480 = n2478 & n2479 ;
  assign n2481 = \P2_IR_reg[31]/NET0131  & ~n1965 ;
  assign n2482 = ~n2455 & ~n2481 ;
  assign n2483 = \P2_IR_reg[7]/NET0131  & ~n2482 ;
  assign n2484 = ~\P2_IR_reg[7]/NET0131  & n2482 ;
  assign n2485 = ~n2483 & ~n2484 ;
  assign n2486 = n2059 & ~n2485 ;
  assign n2487 = \P1_datao_reg[7]/NET0131  & ~n543 ;
  assign n2488 = ~n2108 & ~n2111 ;
  assign n2490 = n2267 & ~n2488 ;
  assign n2489 = ~n2267 & n2488 ;
  assign n2491 = n543 & ~n2489 ;
  assign n2492 = ~n2490 & n2491 ;
  assign n2493 = ~n2487 & ~n2492 ;
  assign n2494 = ~n2059 & n2493 ;
  assign n2495 = ~n2486 & ~n2494 ;
  assign n2496 = n2480 & ~n2495 ;
  assign n2497 = ~n2471 & ~n2496 ;
  assign n2546 = \P2_reg0_reg[2]/NET0131  & n2245 ;
  assign n2547 = \P2_reg1_reg[2]/NET0131  & n2247 ;
  assign n2550 = ~n2546 & ~n2547 ;
  assign n2548 = \P2_reg2_reg[2]/NET0131  & n2243 ;
  assign n2549 = \P2_reg3_reg[2]/NET0131  & n2216 ;
  assign n2551 = ~n2548 & ~n2549 ;
  assign n2552 = n2550 & n2551 ;
  assign n2553 = \P1_datao_reg[2]/NET0131  & ~n543 ;
  assign n2554 = ~n2121 & ~n2122 ;
  assign n2556 = n2127 & n2554 ;
  assign n2555 = ~n2127 & ~n2554 ;
  assign n2557 = n543 & ~n2555 ;
  assign n2558 = ~n2556 & n2557 ;
  assign n2559 = ~n2553 & ~n2558 ;
  assign n2560 = ~n2059 & ~n2559 ;
  assign n2561 = \P2_IR_reg[31]/NET0131  & ~n1961 ;
  assign n2562 = \P2_IR_reg[2]/NET0131  & n2561 ;
  assign n2563 = ~\P2_IR_reg[2]/NET0131  & ~n2561 ;
  assign n2564 = ~n2562 & ~n2563 ;
  assign n2565 = n2059 & n2564 ;
  assign n2566 = ~n2560 & ~n2565 ;
  assign n2567 = ~n2552 & ~n2566 ;
  assign n2568 = \P2_reg3_reg[1]/NET0131  & n2216 ;
  assign n2569 = \P2_reg0_reg[1]/NET0131  & n2245 ;
  assign n2572 = ~n2568 & ~n2569 ;
  assign n2570 = \P2_reg2_reg[1]/NET0131  & n2243 ;
  assign n2571 = \P2_reg1_reg[1]/NET0131  & n2247 ;
  assign n2573 = ~n2570 & ~n2571 ;
  assign n2574 = n2572 & n2573 ;
  assign n2575 = \P2_IR_reg[0]/NET0131  & \P2_IR_reg[31]/NET0131  ;
  assign n2576 = ~\P2_IR_reg[1]/NET0131  & ~n2575 ;
  assign n2577 = \P2_IR_reg[1]/NET0131  & n2575 ;
  assign n2578 = ~n2576 & ~n2577 ;
  assign n2579 = n2059 & n2578 ;
  assign n2580 = ~\P1_datao_reg[1]/NET0131  & ~n543 ;
  assign n2581 = ~n2123 & ~n2124 ;
  assign n2583 = n2125 & ~n2581 ;
  assign n2582 = ~n2125 & n2581 ;
  assign n2584 = n543 & ~n2582 ;
  assign n2585 = ~n2583 & n2584 ;
  assign n2586 = ~n2580 & ~n2585 ;
  assign n2587 = ~n2059 & n2586 ;
  assign n2588 = ~n2579 & ~n2587 ;
  assign n2589 = n2574 & n2588 ;
  assign n2590 = ~n2574 & ~n2588 ;
  assign n2591 = \P2_reg2_reg[0]/NET0131  & n2243 ;
  assign n2592 = \P2_reg0_reg[0]/NET0131  & n2245 ;
  assign n2595 = ~n2591 & ~n2592 ;
  assign n2593 = \P2_reg1_reg[0]/NET0131  & n2247 ;
  assign n2594 = \P2_reg3_reg[0]/NET0131  & n2216 ;
  assign n2596 = ~n2593 & ~n2594 ;
  assign n2597 = n2595 & n2596 ;
  assign n2598 = \si[0]_pad  & n543 ;
  assign n2599 = ~\P1_datao_reg[0]/NET0131  & ~n2598 ;
  assign n2600 = \P1_datao_reg[0]/NET0131  & n2598 ;
  assign n2601 = ~n2599 & ~n2600 ;
  assign n2602 = ~n2059 & n2601 ;
  assign n2603 = \P2_IR_reg[0]/NET0131  & n2059 ;
  assign n2604 = ~n2602 & ~n2603 ;
  assign n2605 = ~n2597 & ~n2604 ;
  assign n2606 = ~n2590 & ~n2605 ;
  assign n2607 = ~n2589 & ~n2606 ;
  assign n2608 = ~n2567 & ~n2607 ;
  assign n2609 = n2552 & n2566 ;
  assign n2610 = \P2_reg1_reg[3]/NET0131  & n2247 ;
  assign n2611 = \P2_reg2_reg[3]/NET0131  & n2243 ;
  assign n2614 = ~n2610 & ~n2611 ;
  assign n2612 = \P2_reg0_reg[3]/NET0131  & n2245 ;
  assign n2613 = ~\P2_reg3_reg[3]/NET0131  & n2216 ;
  assign n2615 = ~n2612 & ~n2613 ;
  assign n2616 = n2614 & n2615 ;
  assign n2617 = \P1_datao_reg[3]/NET0131  & ~n543 ;
  assign n2618 = ~n2120 & ~n2132 ;
  assign n2620 = ~n2129 & n2618 ;
  assign n2619 = n2129 & ~n2618 ;
  assign n2621 = n543 & ~n2619 ;
  assign n2622 = ~n2620 & n2621 ;
  assign n2623 = ~n2617 & ~n2622 ;
  assign n2624 = ~n2059 & ~n2623 ;
  assign n2625 = \P2_IR_reg[31]/NET0131  & ~n1962 ;
  assign n2626 = ~\P2_IR_reg[3]/NET0131  & ~n2625 ;
  assign n2627 = \P2_IR_reg[31]/NET0131  & \P2_IR_reg[3]/NET0131  ;
  assign n2628 = ~n1962 & n2627 ;
  assign n2629 = ~n2626 & ~n2628 ;
  assign n2630 = n2059 & n2629 ;
  assign n2631 = ~n2624 & ~n2630 ;
  assign n2632 = n2616 & n2631 ;
  assign n2633 = ~n2609 & ~n2632 ;
  assign n2634 = ~\P2_reg3_reg[3]/NET0131  & ~\P2_reg3_reg[4]/NET0131  ;
  assign n2635 = ~n2217 & ~n2634 ;
  assign n2636 = n2216 & n2635 ;
  assign n2637 = \P2_reg2_reg[4]/NET0131  & n2243 ;
  assign n2640 = ~n2636 & ~n2637 ;
  assign n2638 = \P2_reg1_reg[4]/NET0131  & n2247 ;
  assign n2639 = \P2_reg0_reg[4]/NET0131  & n2245 ;
  assign n2641 = ~n2638 & ~n2639 ;
  assign n2642 = n2640 & n2641 ;
  assign n2643 = ~n2625 & ~n2627 ;
  assign n2644 = \P2_IR_reg[4]/NET0131  & ~n2643 ;
  assign n2645 = ~\P2_IR_reg[4]/NET0131  & n2643 ;
  assign n2646 = ~n2644 & ~n2645 ;
  assign n2647 = n2059 & n2646 ;
  assign n2648 = ~\P1_datao_reg[4]/NET0131  & ~n543 ;
  assign n2649 = ~n2119 & ~n2131 ;
  assign n2651 = n2322 & ~n2649 ;
  assign n2650 = ~n2322 & n2649 ;
  assign n2652 = n543 & ~n2650 ;
  assign n2653 = ~n2651 & n2652 ;
  assign n2654 = ~n2648 & ~n2653 ;
  assign n2655 = ~n2059 & n2654 ;
  assign n2656 = ~n2647 & ~n2655 ;
  assign n2657 = n2642 & n2656 ;
  assign n2658 = n2633 & ~n2657 ;
  assign n2659 = ~n2608 & n2658 ;
  assign n2660 = ~n2642 & ~n2656 ;
  assign n2661 = ~n2616 & ~n2631 ;
  assign n2662 = ~n2660 & ~n2661 ;
  assign n2663 = ~n2657 & ~n2662 ;
  assign n2664 = ~n2659 & ~n2663 ;
  assign n2498 = ~\P2_reg3_reg[6]/NET0131  & ~n2218 ;
  assign n2499 = ~n2219 & ~n2498 ;
  assign n2500 = n2216 & n2499 ;
  assign n2501 = \P2_reg0_reg[6]/NET0131  & n2245 ;
  assign n2504 = ~n2500 & ~n2501 ;
  assign n2502 = \P2_reg1_reg[6]/NET0131  & n2247 ;
  assign n2503 = \P2_reg2_reg[6]/NET0131  & n2243 ;
  assign n2505 = ~n2502 & ~n2503 ;
  assign n2506 = n2504 & n2505 ;
  assign n2507 = \P1_datao_reg[6]/NET0131  & ~n543 ;
  assign n2508 = ~n2112 & ~n2114 ;
  assign n2510 = n2409 & ~n2508 ;
  assign n2509 = ~n2409 & n2508 ;
  assign n2511 = n543 & ~n2509 ;
  assign n2512 = ~n2510 & n2511 ;
  assign n2513 = ~n2507 & ~n2512 ;
  assign n2514 = ~n2059 & ~n2513 ;
  assign n2515 = \P2_IR_reg[31]/NET0131  & \P2_IR_reg[5]/NET0131  ;
  assign n2516 = ~n2455 & ~n2515 ;
  assign n2517 = \P2_IR_reg[6]/NET0131  & ~n2516 ;
  assign n2518 = ~\P2_IR_reg[6]/NET0131  & n2516 ;
  assign n2519 = ~n2517 & ~n2518 ;
  assign n2520 = n2059 & n2519 ;
  assign n2521 = ~n2514 & ~n2520 ;
  assign n2522 = n2506 & n2521 ;
  assign n2523 = \P2_reg0_reg[5]/NET0131  & n2245 ;
  assign n2524 = \P2_reg2_reg[5]/NET0131  & n2243 ;
  assign n2529 = ~n2523 & ~n2524 ;
  assign n2525 = ~\P2_reg3_reg[5]/NET0131  & ~n2217 ;
  assign n2526 = ~n2218 & ~n2525 ;
  assign n2527 = n2216 & n2526 ;
  assign n2528 = \P2_reg1_reg[5]/NET0131  & n2247 ;
  assign n2530 = ~n2527 & ~n2528 ;
  assign n2531 = n2529 & n2530 ;
  assign n2532 = \P1_datao_reg[5]/NET0131  & ~n543 ;
  assign n2533 = ~n2113 & ~n2136 ;
  assign n2535 = n2135 & n2533 ;
  assign n2534 = ~n2135 & ~n2533 ;
  assign n2536 = n543 & ~n2534 ;
  assign n2537 = ~n2535 & n2536 ;
  assign n2538 = ~n2532 & ~n2537 ;
  assign n2539 = ~n2059 & ~n2538 ;
  assign n2540 = \P2_IR_reg[5]/NET0131  & ~n2455 ;
  assign n2541 = ~\P2_IR_reg[5]/NET0131  & n2455 ;
  assign n2542 = ~n2540 & ~n2541 ;
  assign n2543 = n2059 & ~n2542 ;
  assign n2544 = ~n2539 & ~n2543 ;
  assign n2545 = n2531 & n2544 ;
  assign n2665 = ~n2522 & ~n2545 ;
  assign n2666 = ~n2664 & n2665 ;
  assign n2667 = n2497 & n2666 ;
  assign n2668 = ~n2506 & ~n2521 ;
  assign n2669 = ~n2531 & ~n2544 ;
  assign n2670 = ~n2522 & n2669 ;
  assign n2671 = ~n2668 & ~n2670 ;
  assign n2672 = n2497 & ~n2671 ;
  assign n2673 = ~n2454 & n2470 ;
  assign n2674 = ~n2480 & n2495 ;
  assign n2675 = ~n2673 & ~n2674 ;
  assign n2676 = ~n2471 & ~n2675 ;
  assign n2677 = ~n2672 & ~n2676 ;
  assign n2678 = ~n2667 & n2677 ;
  assign n2679 = \P2_reg3_reg[11]/NET0131  & n2223 ;
  assign n2680 = ~\P2_reg3_reg[11]/NET0131  & ~n2223 ;
  assign n2681 = ~n2679 & ~n2680 ;
  assign n2682 = n2216 & n2681 ;
  assign n2683 = \P2_reg0_reg[11]/NET0131  & n2245 ;
  assign n2686 = ~n2682 & ~n2683 ;
  assign n2684 = \P2_reg1_reg[11]/NET0131  & n2247 ;
  assign n2685 = \P2_reg2_reg[11]/NET0131  & n2243 ;
  assign n2687 = ~n2684 & ~n2685 ;
  assign n2688 = n2686 & n2687 ;
  assign n2689 = \P2_IR_reg[31]/NET0131  & ~n1969 ;
  assign n2690 = \P2_IR_reg[10]/NET0131  & \P2_IR_reg[31]/NET0131  ;
  assign n2691 = ~n2689 & ~n2690 ;
  assign n2692 = \P2_IR_reg[11]/NET0131  & ~n2691 ;
  assign n2693 = ~\P2_IR_reg[11]/NET0131  & n2691 ;
  assign n2694 = ~n2692 & ~n2693 ;
  assign n2695 = n2059 & ~n2694 ;
  assign n2696 = \P1_datao_reg[11]/NET0131  & ~n543 ;
  assign n2697 = ~n2143 & ~n2151 ;
  assign n2699 = n2276 & ~n2697 ;
  assign n2698 = ~n2276 & n2697 ;
  assign n2700 = n543 & ~n2698 ;
  assign n2701 = ~n2699 & n2700 ;
  assign n2702 = ~n2696 & ~n2701 ;
  assign n2703 = ~n2059 & n2702 ;
  assign n2704 = ~n2695 & ~n2703 ;
  assign n2705 = n2688 & ~n2704 ;
  assign n2706 = \P2_reg1_reg[12]/NET0131  & n2247 ;
  assign n2707 = \P2_reg3_reg[12]/NET0131  & n2679 ;
  assign n2708 = ~\P2_reg3_reg[12]/NET0131  & ~n2679 ;
  assign n2709 = ~n2707 & ~n2708 ;
  assign n2710 = n2216 & n2709 ;
  assign n2713 = ~n2706 & ~n2710 ;
  assign n2711 = \P2_reg2_reg[12]/NET0131  & n2243 ;
  assign n2712 = \P2_reg0_reg[12]/NET0131  & n2245 ;
  assign n2714 = ~n2711 & ~n2712 ;
  assign n2715 = n2713 & n2714 ;
  assign n2716 = \P2_IR_reg[31]/NET0131  & ~n1959 ;
  assign n2717 = ~n2689 & ~n2716 ;
  assign n2718 = \P2_IR_reg[12]/NET0131  & ~n2717 ;
  assign n2719 = ~\P2_IR_reg[12]/NET0131  & n2717 ;
  assign n2720 = ~n2718 & ~n2719 ;
  assign n2721 = n2059 & ~n2720 ;
  assign n2722 = \P1_datao_reg[12]/NET0131  & ~n543 ;
  assign n2723 = ~n2142 & ~n2150 ;
  assign n2724 = ~n2332 & n2341 ;
  assign n2726 = ~n2723 & n2724 ;
  assign n2725 = n2723 & ~n2724 ;
  assign n2727 = n543 & ~n2725 ;
  assign n2728 = ~n2726 & n2727 ;
  assign n2729 = ~n2722 & ~n2728 ;
  assign n2730 = ~n2059 & n2729 ;
  assign n2731 = ~n2721 & ~n2730 ;
  assign n2732 = n2715 & ~n2731 ;
  assign n2733 = ~n2705 & ~n2732 ;
  assign n2734 = ~\P2_reg3_reg[10]/NET0131  & ~n2222 ;
  assign n2735 = ~n2223 & ~n2734 ;
  assign n2736 = n2216 & n2735 ;
  assign n2737 = \P2_reg1_reg[10]/NET0131  & n2247 ;
  assign n2740 = ~n2736 & ~n2737 ;
  assign n2738 = \P2_reg0_reg[10]/NET0131  & n2245 ;
  assign n2739 = \P2_reg2_reg[10]/NET0131  & n2243 ;
  assign n2741 = ~n2738 & ~n2739 ;
  assign n2742 = n2740 & n2741 ;
  assign n2743 = ~\P2_IR_reg[10]/NET0131  & n2689 ;
  assign n2744 = \P2_IR_reg[10]/NET0131  & ~n2689 ;
  assign n2745 = ~n2743 & ~n2744 ;
  assign n2746 = n2059 & n2745 ;
  assign n2747 = \P1_datao_reg[10]/NET0131  & ~n543 ;
  assign n2748 = ~n2144 & ~n2152 ;
  assign n2750 = n2414 & ~n2748 ;
  assign n2749 = ~n2414 & n2748 ;
  assign n2751 = n543 & ~n2749 ;
  assign n2752 = ~n2750 & n2751 ;
  assign n2753 = ~n2747 & ~n2752 ;
  assign n2754 = ~n2059 & n2753 ;
  assign n2755 = ~n2746 & ~n2754 ;
  assign n2756 = n2742 & ~n2755 ;
  assign n2757 = \P2_reg2_reg[9]/NET0131  & n2243 ;
  assign n2758 = \P2_reg1_reg[9]/NET0131  & n2247 ;
  assign n2763 = ~n2757 & ~n2758 ;
  assign n2759 = ~\P2_reg3_reg[9]/NET0131  & ~n2221 ;
  assign n2760 = ~n2222 & ~n2759 ;
  assign n2761 = n2216 & n2760 ;
  assign n2762 = \P2_reg0_reg[9]/NET0131  & n2245 ;
  assign n2764 = ~n2761 & ~n2762 ;
  assign n2765 = n2763 & n2764 ;
  assign n2766 = \P2_IR_reg[31]/NET0131  & ~n2011 ;
  assign n2767 = ~\P2_IR_reg[9]/NET0131  & n2766 ;
  assign n2768 = \P2_IR_reg[9]/NET0131  & ~n2766 ;
  assign n2769 = ~n2767 & ~n2768 ;
  assign n2770 = n2059 & n2769 ;
  assign n2771 = \P1_datao_reg[9]/NET0131  & ~n543 ;
  assign n2772 = ~n2146 & ~n2153 ;
  assign n2774 = n2141 & ~n2772 ;
  assign n2773 = ~n2141 & n2772 ;
  assign n2775 = n543 & ~n2773 ;
  assign n2776 = ~n2774 & n2775 ;
  assign n2777 = ~n2771 & ~n2776 ;
  assign n2778 = ~n2059 & n2777 ;
  assign n2779 = ~n2770 & ~n2778 ;
  assign n2780 = n2765 & ~n2779 ;
  assign n2781 = ~n2756 & ~n2780 ;
  assign n2782 = n2733 & n2781 ;
  assign n2783 = ~n2678 & n2782 ;
  assign n2784 = ~n2742 & n2755 ;
  assign n2785 = ~n2765 & n2779 ;
  assign n2786 = ~n2756 & n2785 ;
  assign n2787 = ~n2784 & ~n2786 ;
  assign n2788 = n2733 & ~n2787 ;
  assign n2789 = ~n2715 & n2731 ;
  assign n2790 = ~n2688 & n2704 ;
  assign n2791 = ~n2789 & ~n2790 ;
  assign n2792 = ~n2732 & ~n2791 ;
  assign n2793 = ~n2788 & ~n2792 ;
  assign n2794 = ~n2783 & n2793 ;
  assign n2795 = \P2_reg3_reg[15]/NET0131  & n2227 ;
  assign n2796 = ~\P2_reg3_reg[16]/NET0131  & ~n2795 ;
  assign n2797 = ~n2229 & ~n2796 ;
  assign n2798 = n2216 & n2797 ;
  assign n2799 = \P2_reg0_reg[16]/NET0131  & n2245 ;
  assign n2802 = ~n2798 & ~n2799 ;
  assign n2800 = \P2_reg2_reg[16]/NET0131  & n2243 ;
  assign n2801 = \P2_reg1_reg[16]/NET0131  & n2247 ;
  assign n2803 = ~n2800 & ~n2801 ;
  assign n2804 = n2802 & n2803 ;
  assign n2805 = \P2_IR_reg[31]/NET0131  & ~n1973 ;
  assign n2806 = \P2_IR_reg[16]/NET0131  & n2805 ;
  assign n2807 = ~\P2_IR_reg[16]/NET0131  & ~n2805 ;
  assign n2808 = ~n2806 & ~n2807 ;
  assign n2809 = n2059 & ~n2808 ;
  assign n2810 = \P1_datao_reg[16]/NET0131  & ~n543 ;
  assign n2811 = ~n2084 & ~n2086 ;
  assign n2813 = n2347 & ~n2811 ;
  assign n2812 = ~n2347 & n2811 ;
  assign n2814 = n543 & ~n2812 ;
  assign n2815 = ~n2813 & n2814 ;
  assign n2816 = ~n2810 & ~n2815 ;
  assign n2817 = ~n2059 & n2816 ;
  assign n2818 = ~n2809 & ~n2817 ;
  assign n2819 = n2804 & ~n2818 ;
  assign n2820 = \P2_reg2_reg[15]/NET0131  & n2243 ;
  assign n2821 = ~\P2_reg3_reg[15]/NET0131  & ~n2227 ;
  assign n2822 = ~n2795 & ~n2821 ;
  assign n2823 = n2216 & n2822 ;
  assign n2826 = ~n2820 & ~n2823 ;
  assign n2824 = \P2_reg1_reg[15]/NET0131  & n2247 ;
  assign n2825 = \P2_reg0_reg[15]/NET0131  & n2245 ;
  assign n2827 = ~n2824 & ~n2825 ;
  assign n2828 = n2826 & n2827 ;
  assign n2829 = \P2_IR_reg[31]/NET0131  & ~n1972 ;
  assign n2830 = \P2_IR_reg[15]/NET0131  & n2829 ;
  assign n2831 = ~\P2_IR_reg[15]/NET0131  & ~n2829 ;
  assign n2832 = ~n2830 & ~n2831 ;
  assign n2833 = n2059 & ~n2832 ;
  assign n2834 = \P1_datao_reg[15]/NET0131  & ~n543 ;
  assign n2835 = ~n2279 & ~n2285 ;
  assign n2836 = ~n2085 & ~n2089 ;
  assign n2838 = ~n2835 & n2836 ;
  assign n2837 = n2835 & ~n2836 ;
  assign n2839 = n543 & ~n2837 ;
  assign n2840 = ~n2838 & n2839 ;
  assign n2841 = ~n2834 & ~n2840 ;
  assign n2842 = ~n2059 & n2841 ;
  assign n2843 = ~n2833 & ~n2842 ;
  assign n2844 = n2828 & ~n2843 ;
  assign n2845 = ~n2819 & ~n2844 ;
  assign n2846 = \P2_IR_reg[31]/NET0131  & ~n1971 ;
  assign n2847 = \P2_IR_reg[14]/NET0131  & n2846 ;
  assign n2848 = ~\P2_IR_reg[14]/NET0131  & ~n2846 ;
  assign n2849 = ~n2847 & ~n2848 ;
  assign n2850 = n2059 & ~n2849 ;
  assign n2851 = \P1_datao_reg[14]/NET0131  & ~n543 ;
  assign n2852 = ~n2416 & n2423 ;
  assign n2853 = ~n2088 & ~n2092 ;
  assign n2855 = ~n2852 & n2853 ;
  assign n2854 = n2852 & ~n2853 ;
  assign n2856 = n543 & ~n2854 ;
  assign n2857 = ~n2855 & n2856 ;
  assign n2858 = ~n2851 & ~n2857 ;
  assign n2859 = ~n2059 & n2858 ;
  assign n2860 = ~n2850 & ~n2859 ;
  assign n2864 = \P2_reg3_reg[13]/NET0131  & n2707 ;
  assign n2865 = ~\P2_reg3_reg[14]/NET0131  & ~n2864 ;
  assign n2866 = ~n2227 & ~n2865 ;
  assign n2867 = n2216 & n2866 ;
  assign n2863 = \P2_reg0_reg[14]/NET0131  & n2245 ;
  assign n2861 = \P2_reg2_reg[14]/NET0131  & n2243 ;
  assign n2862 = \P2_reg1_reg[14]/NET0131  & n2247 ;
  assign n2868 = ~n2861 & ~n2862 ;
  assign n2869 = ~n2863 & n2868 ;
  assign n2870 = ~n2867 & n2869 ;
  assign n2871 = ~n2860 & n2870 ;
  assign n2872 = \P2_reg2_reg[13]/NET0131  & n2243 ;
  assign n2873 = ~\P2_reg3_reg[13]/NET0131  & ~n2707 ;
  assign n2874 = ~n2864 & ~n2873 ;
  assign n2875 = n2216 & n2874 ;
  assign n2878 = ~n2872 & ~n2875 ;
  assign n2876 = \P2_reg1_reg[13]/NET0131  & n2247 ;
  assign n2877 = \P2_reg0_reg[13]/NET0131  & n2245 ;
  assign n2879 = ~n2876 & ~n2877 ;
  assign n2880 = n2878 & n2879 ;
  assign n2881 = \P2_IR_reg[13]/NET0131  & ~n2380 ;
  assign n2882 = ~\P2_IR_reg[13]/NET0131  & n2380 ;
  assign n2883 = ~n2881 & ~n2882 ;
  assign n2884 = n2059 & n2883 ;
  assign n2885 = \P1_datao_reg[13]/NET0131  & ~n543 ;
  assign n2886 = ~n2091 & ~n2161 ;
  assign n2888 = n2160 & ~n2886 ;
  assign n2887 = ~n2160 & n2886 ;
  assign n2889 = n543 & ~n2887 ;
  assign n2890 = ~n2888 & n2889 ;
  assign n2891 = ~n2885 & ~n2890 ;
  assign n2892 = ~n2059 & n2891 ;
  assign n2893 = ~n2884 & ~n2892 ;
  assign n2894 = n2880 & ~n2893 ;
  assign n2895 = ~n2871 & ~n2894 ;
  assign n2896 = n2845 & n2895 ;
  assign n2897 = ~n2794 & n2896 ;
  assign n2898 = n2445 & n2897 ;
  assign n2899 = n2860 & ~n2870 ;
  assign n2900 = ~n2880 & n2893 ;
  assign n2901 = ~n2871 & n2900 ;
  assign n2902 = ~n2899 & ~n2901 ;
  assign n2903 = n2845 & ~n2902 ;
  assign n2904 = ~n2804 & n2818 ;
  assign n2905 = ~n2828 & n2843 ;
  assign n2906 = ~n2819 & n2905 ;
  assign n2907 = ~n2904 & ~n2906 ;
  assign n2908 = ~n2903 & n2907 ;
  assign n2909 = n2445 & ~n2908 ;
  assign n2910 = n2433 & ~n2442 ;
  assign n2911 = ~n2379 & n2399 ;
  assign n2912 = ~n2910 & ~n2911 ;
  assign n2913 = ~n2443 & ~n2912 ;
  assign n2914 = n2370 & n2913 ;
  assign n2915 = n2358 & ~n2368 ;
  assign n2916 = n2299 & ~n2311 ;
  assign n2917 = ~n2369 & n2916 ;
  assign n2918 = ~n2915 & ~n2917 ;
  assign n2919 = ~n2914 & n2918 ;
  assign n2920 = ~n2909 & n2919 ;
  assign n2921 = ~n2898 & n2920 ;
  assign n2922 = \P1_datao_reg[28]/NET0131  & ~n543 ;
  assign n2923 = ~n2064 & ~n2171 ;
  assign n2924 = ~n2170 & ~n2173 ;
  assign n2925 = ~n2174 & ~n2183 ;
  assign n2926 = ~n2074 & ~n2925 ;
  assign n2927 = ~n2073 & n2926 ;
  assign n2928 = n2924 & ~n2927 ;
  assign n2929 = ~n2072 & ~n2928 ;
  assign n2930 = ~n2065 & ~n2068 ;
  assign n2931 = ~n2069 & ~n2078 ;
  assign n2932 = n2930 & n2931 ;
  assign n2933 = ~n2351 & n2932 ;
  assign n2934 = ~n2177 & ~n2182 ;
  assign n2935 = ~n2065 & ~n2934 ;
  assign n2936 = ~n2099 & ~n2178 ;
  assign n2937 = ~n2069 & ~n2936 ;
  assign n2938 = n2930 & n2937 ;
  assign n2939 = ~n2935 & ~n2938 ;
  assign n2940 = ~n2933 & n2939 ;
  assign n2941 = ~n2066 & n2076 ;
  assign n2942 = ~n2940 & n2941 ;
  assign n2943 = ~n2929 & ~n2942 ;
  assign n2945 = ~n2923 & n2943 ;
  assign n2944 = n2923 & ~n2943 ;
  assign n2946 = n543 & ~n2944 ;
  assign n2947 = ~n2945 & n2946 ;
  assign n2948 = ~n2922 & ~n2947 ;
  assign n2949 = ~n2059 & ~n2948 ;
  assign n2953 = \P2_reg3_reg[25]/NET0131  & n2237 ;
  assign n2954 = \P2_reg3_reg[26]/NET0131  & n2953 ;
  assign n2955 = \P2_reg3_reg[27]/NET0131  & n2954 ;
  assign n2956 = \P2_reg3_reg[28]/NET0131  & ~n2955 ;
  assign n2957 = ~\P2_reg3_reg[28]/NET0131  & n2955 ;
  assign n2958 = ~n2956 & ~n2957 ;
  assign n2959 = n2216 & ~n2958 ;
  assign n2952 = \P2_reg1_reg[28]/NET0131  & n2247 ;
  assign n2950 = \P2_reg0_reg[28]/NET0131  & n2245 ;
  assign n2951 = \P2_reg2_reg[28]/NET0131  & n2243 ;
  assign n2960 = ~n2950 & ~n2951 ;
  assign n2961 = ~n2952 & n2960 ;
  assign n2962 = ~n2959 & n2961 ;
  assign n2963 = ~n2949 & n2962 ;
  assign n2964 = \P1_datao_reg[27]/NET0131  & ~n543 ;
  assign n2965 = ~n2072 & ~n2170 ;
  assign n2966 = n2075 & n2185 ;
  assign n2967 = ~n2176 & ~n2966 ;
  assign n2968 = n2067 & n2075 ;
  assign n2969 = n2070 & n2101 ;
  assign n2970 = ~n2180 & ~n2969 ;
  assign n2971 = ~n2068 & ~n2080 ;
  assign n2972 = n2931 & n2971 ;
  assign n2973 = ~n2291 & n2972 ;
  assign n2974 = n2970 & ~n2973 ;
  assign n2975 = n2968 & ~n2974 ;
  assign n2976 = n2967 & ~n2975 ;
  assign n2978 = ~n2965 & n2976 ;
  assign n2977 = n2965 & ~n2976 ;
  assign n2979 = n543 & ~n2977 ;
  assign n2980 = ~n2978 & n2979 ;
  assign n2981 = ~n2964 & ~n2980 ;
  assign n2982 = ~n2059 & ~n2981 ;
  assign n2986 = ~\P2_reg3_reg[27]/NET0131  & ~n2954 ;
  assign n2987 = ~n2955 & ~n2986 ;
  assign n2988 = n2216 & n2987 ;
  assign n2985 = \P2_reg2_reg[27]/NET0131  & n2243 ;
  assign n2983 = \P2_reg0_reg[27]/NET0131  & n2245 ;
  assign n2984 = \P2_reg1_reg[27]/NET0131  & n2247 ;
  assign n2989 = ~n2983 & ~n2984 ;
  assign n2990 = ~n2985 & n2989 ;
  assign n2991 = ~n2988 & n2990 ;
  assign n2992 = ~n2982 & n2991 ;
  assign n2993 = ~n2963 & ~n2992 ;
  assign n2994 = \P1_datao_reg[26]/NET0131  & ~n543 ;
  assign n2995 = ~n2073 & ~n2173 ;
  assign n2996 = ~n2066 & ~n2074 ;
  assign n2997 = n2935 & n2996 ;
  assign n2998 = ~n2926 & ~n2997 ;
  assign n2999 = n2930 & n2996 ;
  assign n3000 = ~n2069 & n2082 ;
  assign n3001 = ~n2426 & n3000 ;
  assign n3002 = n2315 & n2931 ;
  assign n3003 = ~n2937 & ~n3002 ;
  assign n3004 = ~n3001 & n3003 ;
  assign n3005 = n2999 & ~n3004 ;
  assign n3006 = n2998 & ~n3005 ;
  assign n3008 = ~n2995 & n3006 ;
  assign n3007 = n2995 & ~n3006 ;
  assign n3009 = n543 & ~n3007 ;
  assign n3010 = ~n3008 & n3009 ;
  assign n3011 = ~n2994 & ~n3010 ;
  assign n3012 = ~n2059 & ~n3011 ;
  assign n3016 = ~\P2_reg3_reg[26]/NET0131  & ~n2953 ;
  assign n3017 = ~n2954 & ~n3016 ;
  assign n3018 = n2216 & n3017 ;
  assign n3015 = \P2_reg2_reg[26]/NET0131  & n2243 ;
  assign n3013 = \P2_reg0_reg[26]/NET0131  & n2245 ;
  assign n3014 = \P2_reg1_reg[26]/NET0131  & n2247 ;
  assign n3019 = ~n3013 & ~n3014 ;
  assign n3020 = ~n3015 & n3019 ;
  assign n3021 = ~n3018 & n3020 ;
  assign n3022 = ~n3012 & n3021 ;
  assign n3023 = \P1_datao_reg[25]/NET0131  & ~n543 ;
  assign n3024 = ~n2074 & ~n2174 ;
  assign n3025 = n2083 & ~n2391 ;
  assign n3026 = n2106 & ~n3025 ;
  assign n3027 = n2071 & ~n3026 ;
  assign n3028 = n2186 & ~n3027 ;
  assign n3030 = ~n3024 & n3028 ;
  assign n3029 = n3024 & ~n3028 ;
  assign n3031 = n543 & ~n3029 ;
  assign n3032 = ~n3030 & n3031 ;
  assign n3033 = ~n3023 & ~n3032 ;
  assign n3034 = ~n2059 & ~n3033 ;
  assign n3038 = ~\P2_reg3_reg[25]/NET0131  & ~n2237 ;
  assign n3039 = ~n2953 & ~n3038 ;
  assign n3040 = n2216 & n3039 ;
  assign n3037 = \P2_reg2_reg[25]/NET0131  & n2243 ;
  assign n3035 = \P2_reg0_reg[25]/NET0131  & n2245 ;
  assign n3036 = \P2_reg1_reg[25]/NET0131  & n2247 ;
  assign n3041 = ~n3035 & ~n3036 ;
  assign n3042 = ~n3037 & n3041 ;
  assign n3043 = ~n3040 & n3042 ;
  assign n3044 = ~n3034 & n3043 ;
  assign n3045 = ~n3022 & ~n3044 ;
  assign n3046 = n2993 & n3045 ;
  assign n3047 = \P1_datao_reg[24]/NET0131  & ~n543 ;
  assign n3048 = ~n2066 & ~n2183 ;
  assign n3050 = n2940 & ~n3048 ;
  assign n3049 = ~n2940 & n3048 ;
  assign n3051 = n543 & ~n3049 ;
  assign n3052 = ~n3050 & n3051 ;
  assign n3053 = ~n3047 & ~n3052 ;
  assign n3054 = ~n2059 & ~n3053 ;
  assign n3055 = n2231 & n2306 ;
  assign n3056 = \P2_reg3_reg[23]/NET0131  & n3055 ;
  assign n3057 = ~\P2_reg3_reg[24]/NET0131  & ~n3056 ;
  assign n3058 = ~n2237 & ~n3057 ;
  assign n3059 = n2216 & n3058 ;
  assign n3062 = \P2_reg0_reg[24]/NET0131  & n2245 ;
  assign n3060 = \P2_reg1_reg[24]/NET0131  & n2247 ;
  assign n3061 = \P2_reg2_reg[24]/NET0131  & n2243 ;
  assign n3063 = ~n3060 & ~n3061 ;
  assign n3064 = ~n3062 & n3063 ;
  assign n3065 = ~n3059 & n3064 ;
  assign n3066 = ~n3054 & n3065 ;
  assign n3067 = \P1_datao_reg[23]/NET0131  & ~n543 ;
  assign n3068 = ~n2065 & ~n2182 ;
  assign n3070 = n2263 & n2972 ;
  assign n3071 = ~n2835 & n3070 ;
  assign n3069 = n2289 & n2972 ;
  assign n3072 = n2970 & ~n3069 ;
  assign n3073 = ~n3071 & n3072 ;
  assign n3075 = ~n3068 & n3073 ;
  assign n3074 = n3068 & ~n3073 ;
  assign n3076 = n543 & ~n3074 ;
  assign n3077 = ~n3075 & n3076 ;
  assign n3078 = ~n3067 & ~n3077 ;
  assign n3079 = ~n2059 & ~n3078 ;
  assign n3083 = ~\P2_reg3_reg[23]/NET0131  & ~n3055 ;
  assign n3084 = ~n3056 & ~n3083 ;
  assign n3085 = n2216 & n3084 ;
  assign n3082 = \P2_reg1_reg[23]/NET0131  & n2247 ;
  assign n3080 = \P2_reg0_reg[23]/NET0131  & n2245 ;
  assign n3081 = \P2_reg2_reg[23]/NET0131  & n2243 ;
  assign n3086 = ~n3080 & ~n3081 ;
  assign n3087 = ~n3082 & n3086 ;
  assign n3088 = ~n3085 & n3087 ;
  assign n3089 = ~n3079 & n3088 ;
  assign n3090 = ~n3066 & ~n3089 ;
  assign n3091 = \P1_datao_reg[22]/NET0131  & ~n543 ;
  assign n3092 = ~n2068 & ~n2177 ;
  assign n3093 = n2417 & ~n2852 ;
  assign n3094 = n2420 & ~n3093 ;
  assign n3095 = n3000 & ~n3094 ;
  assign n3096 = n3003 & ~n3095 ;
  assign n3098 = ~n3092 & n3096 ;
  assign n3097 = n3092 & ~n3096 ;
  assign n3099 = n543 & ~n3097 ;
  assign n3100 = ~n3098 & n3099 ;
  assign n3101 = ~n3091 & ~n3100 ;
  assign n3102 = ~n2059 & ~n3101 ;
  assign n3106 = n2230 & n2306 ;
  assign n3107 = ~\P2_reg3_reg[22]/NET0131  & ~n3106 ;
  assign n3108 = ~n3055 & ~n3107 ;
  assign n3109 = n2216 & n3108 ;
  assign n3105 = \P2_reg2_reg[22]/NET0131  & n2243 ;
  assign n3103 = \P2_reg0_reg[22]/NET0131  & n2245 ;
  assign n3104 = \P2_reg1_reg[22]/NET0131  & n2247 ;
  assign n3110 = ~n3103 & ~n3104 ;
  assign n3111 = ~n3105 & n3110 ;
  assign n3112 = ~n3109 & n3111 ;
  assign n3113 = ~n3102 & n3112 ;
  assign n3114 = \P1_datao_reg[21]/NET0131  & ~n543 ;
  assign n3115 = ~n2069 & ~n2178 ;
  assign n3117 = n2167 & ~n3115 ;
  assign n3116 = ~n2167 & n3115 ;
  assign n3118 = n543 & ~n3116 ;
  assign n3119 = ~n3117 & n3118 ;
  assign n3120 = ~n3114 & ~n3119 ;
  assign n3121 = ~n2059 & ~n3120 ;
  assign n3125 = ~\P2_reg3_reg[21]/NET0131  & ~n2362 ;
  assign n3126 = ~n3106 & ~n3125 ;
  assign n3127 = n2216 & n3126 ;
  assign n3124 = \P2_reg1_reg[21]/NET0131  & n2247 ;
  assign n3122 = \P2_reg2_reg[21]/NET0131  & n2243 ;
  assign n3123 = \P2_reg0_reg[21]/NET0131  & n2245 ;
  assign n3128 = ~n3122 & ~n3123 ;
  assign n3129 = ~n3124 & n3128 ;
  assign n3130 = ~n3127 & n3129 ;
  assign n3131 = ~n3121 & n3130 ;
  assign n3132 = ~n3113 & ~n3131 ;
  assign n3133 = n3090 & n3132 ;
  assign n3134 = n3046 & n3133 ;
  assign n3135 = ~n2921 & n3134 ;
  assign n3138 = n3102 & ~n3112 ;
  assign n3139 = n3121 & ~n3130 ;
  assign n3140 = ~n3113 & n3139 ;
  assign n3141 = ~n3138 & ~n3140 ;
  assign n3142 = n3090 & ~n3141 ;
  assign n3143 = n3054 & ~n3065 ;
  assign n3144 = n3079 & ~n3088 ;
  assign n3145 = ~n3066 & n3144 ;
  assign n3146 = ~n3143 & ~n3145 ;
  assign n3147 = ~n3142 & n3146 ;
  assign n3148 = n3046 & ~n3147 ;
  assign n3149 = n3012 & ~n3021 ;
  assign n3150 = n3034 & ~n3043 ;
  assign n3151 = ~n3022 & n3150 ;
  assign n3152 = ~n3149 & ~n3151 ;
  assign n3153 = n2993 & ~n3152 ;
  assign n3136 = n2982 & ~n2991 ;
  assign n3137 = ~n2963 & n3136 ;
  assign n3154 = n2949 & ~n2962 ;
  assign n3155 = ~n3137 & ~n3154 ;
  assign n3156 = ~n3153 & n3155 ;
  assign n3157 = ~n3148 & n3156 ;
  assign n3158 = ~n3135 & n3157 ;
  assign n3159 = n2254 & ~n3158 ;
  assign n3160 = ~n2254 & n3158 ;
  assign n3161 = ~n3159 & ~n3160 ;
  assign n3162 = n2040 & ~n3161 ;
  assign n3163 = ~n2041 & ~n3162 ;
  assign n3164 = ~\P2_IR_reg[22]/NET0131  & ~n2199 ;
  assign n3165 = \P2_IR_reg[22]/NET0131  & n2199 ;
  assign n3166 = ~n3164 & ~n3165 ;
  assign n3167 = ~n1982 & n3166 ;
  assign n3168 = \P2_IR_reg[21]/NET0131  & ~n2208 ;
  assign n3169 = ~\P2_IR_reg[21]/NET0131  & n2208 ;
  assign n3170 = ~n3168 & ~n3169 ;
  assign n3171 = n3167 & n3170 ;
  assign n3172 = n1982 & ~n3166 ;
  assign n3173 = \P2_IR_reg[20]/NET0131  & ~n2042 ;
  assign n3174 = ~\P2_IR_reg[20]/NET0131  & n2042 ;
  assign n3175 = ~n3173 & ~n3174 ;
  assign n3176 = n3172 & n3175 ;
  assign n3177 = ~n3171 & ~n3176 ;
  assign n3178 = ~n3163 & ~n3177 ;
  assign n3210 = n2299 & n2311 ;
  assign n3211 = n2358 & n2368 ;
  assign n3212 = ~n3210 & ~n3211 ;
  assign n3213 = n2379 & n2399 ;
  assign n3214 = n2433 & n2442 ;
  assign n3215 = ~n3213 & ~n3214 ;
  assign n3216 = n3212 & n3215 ;
  assign n3217 = n2804 & n2818 ;
  assign n3218 = n2828 & n2843 ;
  assign n3219 = ~n3217 & ~n3218 ;
  assign n3220 = n2860 & n2870 ;
  assign n3221 = n2880 & n2893 ;
  assign n3222 = ~n3220 & ~n3221 ;
  assign n3223 = n3219 & n3222 ;
  assign n3224 = n3216 & n3223 ;
  assign n3225 = n2688 & n2704 ;
  assign n3226 = n2715 & n2731 ;
  assign n3227 = ~n3225 & ~n3226 ;
  assign n3228 = ~n2742 & ~n2755 ;
  assign n3229 = n2742 & n2755 ;
  assign n3230 = ~n2765 & ~n2779 ;
  assign n3231 = ~n3229 & n3230 ;
  assign n3232 = ~n3228 & ~n3231 ;
  assign n3233 = n3227 & ~n3232 ;
  assign n3234 = ~n2715 & ~n2731 ;
  assign n3235 = ~n2688 & ~n2704 ;
  assign n3236 = ~n3226 & n3235 ;
  assign n3237 = ~n3234 & ~n3236 ;
  assign n3238 = ~n3233 & n3237 ;
  assign n3254 = ~n2552 & n2566 ;
  assign n3255 = ~n2574 & n2588 ;
  assign n3256 = ~n3254 & ~n3255 ;
  assign n3257 = n2574 & ~n2588 ;
  assign n3258 = n2597 & ~n2604 ;
  assign n3259 = ~n3257 & ~n3258 ;
  assign n3260 = n3256 & ~n3259 ;
  assign n3261 = n2552 & ~n2566 ;
  assign n3262 = n2616 & ~n2631 ;
  assign n3263 = ~n3261 & ~n3262 ;
  assign n3264 = n2642 & ~n2656 ;
  assign n3265 = n3263 & ~n3264 ;
  assign n3266 = ~n3260 & n3265 ;
  assign n3267 = ~n2642 & n2656 ;
  assign n3268 = ~n2616 & n2631 ;
  assign n3269 = ~n3267 & ~n3268 ;
  assign n3270 = ~n3264 & ~n3269 ;
  assign n3271 = ~n3266 & ~n3270 ;
  assign n3241 = n2480 & n2495 ;
  assign n3242 = n2454 & n2470 ;
  assign n3243 = ~n3241 & ~n3242 ;
  assign n3244 = n2506 & ~n2521 ;
  assign n3272 = n2531 & ~n2544 ;
  assign n3273 = ~n3244 & ~n3272 ;
  assign n3274 = n3243 & n3273 ;
  assign n3275 = ~n3271 & n3274 ;
  assign n3245 = ~n2506 & n2521 ;
  assign n3246 = ~n2531 & n2544 ;
  assign n3247 = ~n3245 & ~n3246 ;
  assign n3248 = ~n3244 & ~n3247 ;
  assign n3249 = n3243 & n3248 ;
  assign n3250 = ~n2454 & ~n2470 ;
  assign n3251 = ~n2480 & ~n2495 ;
  assign n3252 = ~n3242 & n3251 ;
  assign n3253 = ~n3250 & ~n3252 ;
  assign n3276 = ~n3249 & n3253 ;
  assign n3277 = ~n3275 & n3276 ;
  assign n3239 = n2765 & n2779 ;
  assign n3240 = ~n3229 & ~n3239 ;
  assign n3278 = n3227 & n3240 ;
  assign n3279 = ~n3277 & n3278 ;
  assign n3280 = n3238 & ~n3279 ;
  assign n3281 = n3224 & ~n3280 ;
  assign n3282 = ~n2860 & ~n2870 ;
  assign n3283 = ~n2880 & ~n2893 ;
  assign n3284 = ~n3282 & ~n3283 ;
  assign n3285 = ~n3220 & ~n3284 ;
  assign n3286 = n3219 & n3285 ;
  assign n3287 = ~n2804 & ~n2818 ;
  assign n3288 = ~n2828 & ~n2843 ;
  assign n3289 = ~n3287 & ~n3288 ;
  assign n3290 = ~n3217 & ~n3289 ;
  assign n3291 = ~n3286 & ~n3290 ;
  assign n3292 = n3216 & ~n3291 ;
  assign n3293 = ~n2433 & ~n2442 ;
  assign n3294 = ~n2379 & ~n2399 ;
  assign n3295 = ~n3293 & ~n3294 ;
  assign n3296 = ~n3214 & ~n3295 ;
  assign n3297 = n3212 & n3296 ;
  assign n3298 = ~n2358 & ~n2368 ;
  assign n3299 = ~n2299 & ~n2311 ;
  assign n3300 = ~n3298 & ~n3299 ;
  assign n3301 = ~n3211 & ~n3300 ;
  assign n3302 = ~n3297 & ~n3301 ;
  assign n3303 = ~n3292 & n3302 ;
  assign n3304 = ~n3281 & n3303 ;
  assign n3179 = n2949 & n2962 ;
  assign n3180 = n2982 & n2991 ;
  assign n3181 = ~n3179 & ~n3180 ;
  assign n3182 = n3012 & n3021 ;
  assign n3183 = n3034 & n3043 ;
  assign n3184 = ~n3182 & ~n3183 ;
  assign n3185 = n3181 & n3184 ;
  assign n3186 = n3079 & n3088 ;
  assign n3187 = n3054 & n3065 ;
  assign n3188 = ~n3186 & ~n3187 ;
  assign n3189 = n3102 & n3112 ;
  assign n3305 = n3121 & n3130 ;
  assign n3306 = ~n3189 & ~n3305 ;
  assign n3307 = n3188 & n3306 ;
  assign n3308 = n3185 & n3307 ;
  assign n3309 = ~n3304 & n3308 ;
  assign n3190 = ~n3102 & ~n3112 ;
  assign n3191 = ~n3121 & ~n3130 ;
  assign n3192 = ~n3190 & ~n3191 ;
  assign n3193 = ~n3189 & ~n3192 ;
  assign n3194 = n3188 & n3193 ;
  assign n3195 = ~n3054 & ~n3065 ;
  assign n3196 = ~n3079 & ~n3088 ;
  assign n3197 = ~n3187 & n3196 ;
  assign n3198 = ~n3195 & ~n3197 ;
  assign n3199 = ~n3194 & n3198 ;
  assign n3200 = n3185 & ~n3199 ;
  assign n3201 = ~n3012 & ~n3021 ;
  assign n3202 = ~n3034 & ~n3043 ;
  assign n3203 = ~n3201 & ~n3202 ;
  assign n3204 = ~n3182 & ~n3203 ;
  assign n3205 = n3181 & n3204 ;
  assign n3206 = ~n2949 & ~n2962 ;
  assign n3207 = ~n2982 & ~n2991 ;
  assign n3208 = ~n3206 & ~n3207 ;
  assign n3209 = ~n3179 & ~n3208 ;
  assign n3310 = ~n3205 & ~n3209 ;
  assign n3311 = ~n3200 & n3310 ;
  assign n3312 = ~n3309 & n3311 ;
  assign n3313 = n2254 & ~n3312 ;
  assign n3314 = ~n2254 & n3312 ;
  assign n3315 = ~n3313 & ~n3314 ;
  assign n3316 = n2040 & n3315 ;
  assign n3317 = ~n2041 & ~n3316 ;
  assign n3318 = n3172 & ~n3175 ;
  assign n3319 = n3167 & ~n3170 ;
  assign n3320 = ~n3318 & ~n3319 ;
  assign n3321 = ~n3317 & ~n3320 ;
  assign n3326 = n2588 & n2604 ;
  assign n3327 = n2566 & n3326 ;
  assign n3328 = n2631 & n3327 ;
  assign n3329 = n2656 & n3328 ;
  assign n3330 = n2544 & n3329 ;
  assign n3331 = n2521 & n3330 ;
  assign n3332 = ~n2495 & n3331 ;
  assign n3333 = ~n2470 & ~n2779 ;
  assign n3334 = n3332 & n3333 ;
  assign n3335 = ~n2704 & ~n2755 ;
  assign n3336 = n3334 & n3335 ;
  assign n3337 = ~n2731 & n3336 ;
  assign n3338 = ~n2860 & ~n2893 ;
  assign n3339 = n3337 & n3338 ;
  assign n3340 = ~n2399 & ~n2818 ;
  assign n3341 = ~n2433 & ~n2843 ;
  assign n3342 = n3340 & n3341 ;
  assign n3343 = n3339 & n3342 ;
  assign n3322 = ~n2299 & ~n2358 ;
  assign n3323 = ~n3079 & ~n3121 ;
  assign n3324 = ~n3102 & n3323 ;
  assign n3325 = n3322 & n3324 ;
  assign n3344 = ~n3034 & ~n3054 ;
  assign n3345 = n3325 & n3344 ;
  assign n3346 = n3343 & n3345 ;
  assign n3347 = ~n2982 & ~n3012 ;
  assign n3348 = ~n2949 & n3347 ;
  assign n3349 = n3346 & n3348 ;
  assign n3350 = ~n2198 & n3349 ;
  assign n3351 = n2198 & ~n3349 ;
  assign n3352 = ~n3350 & ~n3351 ;
  assign n3353 = n3170 & n3175 ;
  assign n3354 = ~n3166 & n3353 ;
  assign n3355 = ~n1982 & n3354 ;
  assign n3356 = n3352 & n3355 ;
  assign n3357 = ~n1982 & ~n3166 ;
  assign n3358 = ~n3170 & n3357 ;
  assign n3359 = n2198 & n3358 ;
  assign n3360 = n2058 & ~n2962 ;
  assign n3367 = \P2_reg2_reg[31]/NET0131  & n2243 ;
  assign n3370 = ~n2242 & ~n3367 ;
  assign n3368 = \P2_reg0_reg[31]/NET0131  & n2245 ;
  assign n3369 = \P2_reg1_reg[31]/NET0131  & n2247 ;
  assign n3371 = ~n3368 & ~n3369 ;
  assign n3372 = n3370 & n3371 ;
  assign n3373 = ~n2597 & ~n3372 ;
  assign n3374 = ~n2574 & n3373 ;
  assign n3375 = ~n2552 & n3374 ;
  assign n3376 = ~n2616 & n3375 ;
  assign n3377 = ~n2531 & ~n2642 ;
  assign n3378 = n3376 & n3377 ;
  assign n3379 = ~n2506 & n3378 ;
  assign n3380 = ~n2480 & n3379 ;
  assign n3381 = ~n2454 & ~n2742 ;
  assign n3382 = ~n2765 & n3381 ;
  assign n3383 = n3380 & n3382 ;
  assign n3384 = ~n2688 & ~n2715 ;
  assign n3385 = ~n2880 & n3384 ;
  assign n3386 = ~n2870 & n3385 ;
  assign n3387 = n3383 & n3386 ;
  assign n3388 = ~n2379 & ~n2804 ;
  assign n3389 = ~n2828 & n3388 ;
  assign n3390 = ~n2442 & n3389 ;
  assign n3391 = ~n2311 & ~n2368 ;
  assign n3392 = ~n3130 & n3391 ;
  assign n3393 = n3390 & n3392 ;
  assign n3394 = n3387 & n3393 ;
  assign n3362 = ~n3088 & ~n3112 ;
  assign n3363 = ~n3065 & n3362 ;
  assign n3361 = ~n3021 & ~n3043 ;
  assign n3364 = ~n2991 & n3361 ;
  assign n3365 = n3363 & n3364 ;
  assign n3366 = ~n2962 & n3365 ;
  assign n3395 = ~n2251 & n3366 ;
  assign n3396 = n3394 & n3395 ;
  assign n3397 = \P2_reg2_reg[30]/NET0131  & n2243 ;
  assign n3400 = ~n2242 & ~n3397 ;
  assign n3398 = \P2_reg0_reg[30]/NET0131  & n2245 ;
  assign n3399 = \P2_reg1_reg[30]/NET0131  & n2247 ;
  assign n3401 = ~n3398 & ~n3399 ;
  assign n3402 = n3400 & n3401 ;
  assign n3403 = ~n3396 & n3402 ;
  assign n3404 = n3396 & ~n3402 ;
  assign n3405 = \P2_B_reg/NET0131  & n2051 ;
  assign n3406 = ~n2058 & ~n3405 ;
  assign n3407 = ~n3404 & n3406 ;
  assign n3408 = ~n3403 & n3407 ;
  assign n3409 = ~n3360 & ~n3408 ;
  assign n3410 = n1982 & n3166 ;
  assign n3411 = n3353 & n3410 ;
  assign n3412 = ~n3409 & n3411 ;
  assign n3413 = ~n3359 & ~n3412 ;
  assign n3414 = ~n3356 & n3413 ;
  assign n3415 = n2040 & ~n3414 ;
  assign n3416 = ~n2040 & n3411 ;
  assign n3417 = ~n3353 & n3410 ;
  assign n3418 = n3170 & ~n3175 ;
  assign n3419 = ~n3166 & n3418 ;
  assign n3420 = ~n1982 & n3419 ;
  assign n3421 = ~n3417 & ~n3420 ;
  assign n3422 = ~n2040 & n3358 ;
  assign n3423 = n3421 & ~n3422 ;
  assign n3424 = ~n2040 & n3355 ;
  assign n3425 = n3423 & ~n3424 ;
  assign n3426 = ~n3416 & n3425 ;
  assign n3427 = \P2_reg0_reg[29]/NET0131  & ~n3426 ;
  assign n3428 = ~n3415 & ~n3427 ;
  assign n3429 = ~n3321 & n3428 ;
  assign n3430 = ~n3178 & n3429 ;
  assign n3431 = n2026 & ~n3430 ;
  assign n3432 = ~n2025 & ~n3431 ;
  assign n3433 = \P1_state_reg[0]/NET0131  & ~n3432 ;
  assign n3434 = ~n1984 & ~n3433 ;
  assign n3435 = \P1_state_reg[0]/NET0131  & n512 ;
  assign n3436 = \P1_reg2_reg[29]/NET0131  & ~n3435 ;
  assign n3443 = ~\P1_IR_reg[24]/NET0131  & ~n530 ;
  assign n3444 = \P1_IR_reg[24]/NET0131  & n530 ;
  assign n3445 = ~n3443 & ~n3444 ;
  assign n3437 = \P1_IR_reg[25]/NET0131  & ~n708 ;
  assign n3438 = ~\P1_IR_reg[25]/NET0131  & n708 ;
  assign n3439 = ~n3437 & ~n3438 ;
  assign n3440 = \P1_IR_reg[26]/NET0131  & ~n696 ;
  assign n3441 = ~\P1_IR_reg[26]/NET0131  & n696 ;
  assign n3442 = ~n3440 & ~n3441 ;
  assign n3446 = ~n3439 & ~n3442 ;
  assign n3447 = n3445 & n3446 ;
  assign n3448 = n512 & n3447 ;
  assign n3449 = \P1_reg2_reg[29]/NET0131  & n3448 ;
  assign n3450 = n512 & ~n3447 ;
  assign n3451 = n3439 & ~n3442 ;
  assign n3452 = ~\P1_B_reg/NET0131  & n3445 ;
  assign n3453 = n3451 & n3452 ;
  assign n3454 = ~\P1_d_reg[0]/NET0131  & ~n3453 ;
  assign n3455 = ~n3442 & ~n3454 ;
  assign n3456 = \P1_B_reg/NET0131  & ~n3445 ;
  assign n3457 = n3451 & n3456 ;
  assign n3458 = n3442 & n3445 ;
  assign n3459 = ~n3457 & ~n3458 ;
  assign n3460 = ~n3455 & n3459 ;
  assign n3461 = \P1_d_reg[1]/NET0131  & ~n3442 ;
  assign n3462 = ~n3439 & n3442 ;
  assign n3463 = ~n3461 & ~n3462 ;
  assign n3464 = ~n3453 & n3463 ;
  assign n3465 = ~n3457 & n3464 ;
  assign n3466 = n3460 & ~n3465 ;
  assign n3467 = \P1_reg2_reg[29]/NET0131  & ~n3466 ;
  assign n3468 = ~n1816 & ~n1820 ;
  assign n3469 = ~n1836 & n1840 ;
  assign n3470 = ~n1837 & ~n3469 ;
  assign n3471 = n3468 & ~n3470 ;
  assign n3472 = ~n1816 & n1819 ;
  assign n3473 = ~n1817 & ~n3472 ;
  assign n3474 = ~n3471 & n3473 ;
  assign n3475 = ~n1767 & ~n1808 ;
  assign n3476 = ~n1810 & n3475 ;
  assign n3477 = ~n3474 & n3476 ;
  assign n3478 = ~n1807 & ~n1811 ;
  assign n3479 = n3475 & ~n3478 ;
  assign n3480 = ~n1768 & ~n3479 ;
  assign n3481 = ~n1830 & n3480 ;
  assign n3482 = ~n3477 & n3481 ;
  assign n3483 = ~n1829 & ~n3482 ;
  assign n3484 = ~n1826 & ~n1833 ;
  assign n3485 = ~n1443 & n1452 ;
  assign n3486 = ~n1822 & ~n3485 ;
  assign n3487 = n3484 & n3486 ;
  assign n3488 = ~n1797 & ~n1813 ;
  assign n3489 = ~n1783 & ~n1786 ;
  assign n3490 = n3488 & n3489 ;
  assign n3491 = n3487 & n3490 ;
  assign n3492 = ~n1770 & ~n1794 ;
  assign n3493 = n1780 & ~n1790 ;
  assign n3494 = ~n1789 & ~n3493 ;
  assign n3495 = n3492 & ~n3494 ;
  assign n3496 = n1771 & ~n1794 ;
  assign n3497 = ~n1795 & ~n3496 ;
  assign n3498 = ~n3495 & n3497 ;
  assign n3503 = n1641 & n1655 ;
  assign n3504 = ~n1641 & ~n1655 ;
  assign n3505 = ~n1664 & ~n1671 ;
  assign n3506 = ~n3504 & ~n3505 ;
  assign n3507 = ~n3503 & ~n3506 ;
  assign n3508 = ~n1777 & ~n3507 ;
  assign n3509 = n1617 & n1632 ;
  assign n3510 = ~n1778 & ~n3509 ;
  assign n3511 = n1572 & n1586 ;
  assign n3512 = n3510 & ~n3511 ;
  assign n3513 = ~n3508 & n3512 ;
  assign n3514 = ~n1572 & ~n1586 ;
  assign n3515 = ~n1617 & ~n1632 ;
  assign n3516 = ~n3511 & n3515 ;
  assign n3517 = ~n3514 & ~n3516 ;
  assign n3518 = ~n3513 & n3517 ;
  assign n3499 = n1524 & n1537 ;
  assign n3500 = n1548 & n1562 ;
  assign n3501 = ~n3499 & ~n3500 ;
  assign n3502 = ~n1774 & ~n1800 ;
  assign n3519 = n3501 & n3502 ;
  assign n3520 = ~n3518 & n3519 ;
  assign n3521 = ~n1524 & ~n1537 ;
  assign n3522 = ~n1548 & ~n1562 ;
  assign n3523 = ~n3499 & n3522 ;
  assign n3524 = ~n3521 & ~n3523 ;
  assign n3525 = n3502 & ~n3524 ;
  assign n3526 = n1775 & ~n1800 ;
  assign n3527 = ~n1801 & ~n3526 ;
  assign n3528 = ~n3525 & n3527 ;
  assign n3529 = ~n3520 & n3528 ;
  assign n3530 = ~n1781 & ~n1790 ;
  assign n3531 = n3492 & n3530 ;
  assign n3532 = ~n3529 & n3531 ;
  assign n3533 = n3498 & ~n3532 ;
  assign n3534 = n3491 & ~n3533 ;
  assign n3535 = n1798 & ~n1813 ;
  assign n3536 = ~n1814 & ~n3535 ;
  assign n3537 = n3489 & ~n3536 ;
  assign n3538 = ~n1784 & ~n1787 ;
  assign n3539 = ~n1783 & ~n3538 ;
  assign n3540 = ~n3537 & ~n3539 ;
  assign n3541 = n3487 & ~n3540 ;
  assign n3542 = n1443 & ~n1452 ;
  assign n3543 = ~n1822 & n3542 ;
  assign n3544 = ~n1823 & ~n3543 ;
  assign n3545 = n3484 & ~n3544 ;
  assign n3546 = ~n1826 & n1834 ;
  assign n3547 = ~n1827 & ~n3546 ;
  assign n3548 = ~n3545 & n3547 ;
  assign n3549 = ~n3541 & n3548 ;
  assign n3550 = ~n3534 & n3549 ;
  assign n3551 = ~n1836 & ~n1839 ;
  assign n3552 = n3468 & n3551 ;
  assign n3553 = ~n1829 & n3476 ;
  assign n3554 = n3552 & n3553 ;
  assign n3555 = ~n3550 & n3554 ;
  assign n3556 = ~n3483 & ~n3555 ;
  assign n3557 = n1832 & ~n3556 ;
  assign n3558 = ~n1832 & n3556 ;
  assign n3559 = ~n3557 & ~n3558 ;
  assign n3560 = n3466 & ~n3559 ;
  assign n3561 = ~n3467 & ~n3560 ;
  assign n3562 = ~n501 & n1888 ;
  assign n3563 = ~n1766 & ~n3562 ;
  assign n3564 = ~n3561 & ~n3563 ;
  assign n3679 = n1655 & n1671 ;
  assign n3680 = n1609 & n3679 ;
  assign n3681 = n1632 & n3680 ;
  assign n3682 = n1586 & n3681 ;
  assign n3683 = n1562 & n3682 ;
  assign n3684 = n1537 & n3683 ;
  assign n3685 = ~n1281 & n1514 ;
  assign n3686 = ~n1257 & n3685 ;
  assign n3687 = n3684 & n3686 ;
  assign n3688 = ~n1198 & ~n1233 ;
  assign n3689 = ~n1165 & n3688 ;
  assign n3690 = n3687 & n3689 ;
  assign n3692 = ~n1136 & ~n1466 ;
  assign n3693 = ~n1394 & n3692 ;
  assign n3691 = ~n1083 & ~n1109 ;
  assign n3694 = ~n1443 & n3691 ;
  assign n3695 = n3693 & n3694 ;
  assign n3696 = n3690 & n3695 ;
  assign n3697 = ~n1365 & ~n1418 ;
  assign n3698 = n3696 & n3697 ;
  assign n3699 = ~n1309 & ~n1346 ;
  assign n3700 = n3698 & n3699 ;
  assign n3701 = ~n1047 & ~n1327 ;
  assign n3702 = ~n997 & ~n1029 ;
  assign n3703 = n3701 & n3702 ;
  assign n3704 = n3700 & n3703 ;
  assign n3705 = ~n933 & ~n969 ;
  assign n3706 = n3704 & n3705 ;
  assign n3707 = n881 & ~n3706 ;
  assign n3708 = ~n881 & n3706 ;
  assign n3709 = ~n3707 & ~n3708 ;
  assign n3710 = n3466 & n3709 ;
  assign n3711 = ~n3467 & ~n3710 ;
  assign n3712 = n512 & n1886 ;
  assign n3713 = ~n3711 & n3712 ;
  assign n3714 = n881 & n1880 ;
  assign n3715 = n3466 & n3714 ;
  assign n3716 = ~n1885 & n1935 ;
  assign n3717 = n1880 & ~n3466 ;
  assign n3718 = ~n3716 & ~n3717 ;
  assign n3719 = \P1_reg2_reg[29]/NET0131  & ~n3718 ;
  assign n3720 = n740 & n1763 ;
  assign n3721 = ~n3719 & ~n3720 ;
  assign n3722 = ~n3715 & n3721 ;
  assign n3723 = ~n3713 & n3722 ;
  assign n3724 = ~n3564 & n3723 ;
  assign n3565 = n537 & ~n945 ;
  assign n3570 = ~n750 & ~n1664 ;
  assign n3571 = ~n1641 & n3570 ;
  assign n3572 = ~n1595 & n3571 ;
  assign n3573 = ~n1617 & n3572 ;
  assign n3574 = ~n1548 & ~n1572 ;
  assign n3575 = n3573 & n3574 ;
  assign n3576 = ~n1498 & ~n1524 ;
  assign n3577 = n3575 & n3576 ;
  assign n3578 = ~n1218 & ~n1244 ;
  assign n3579 = ~n1267 & n3578 ;
  assign n3580 = n3577 & n3579 ;
  assign n3581 = ~n1146 & ~n1174 ;
  assign n3582 = ~n1207 & n3581 ;
  assign n3583 = n3580 & n3582 ;
  assign n3568 = ~n1452 & ~n1475 ;
  assign n3569 = ~n1094 & ~n1118 ;
  assign n3584 = n3568 & n3569 ;
  assign n3585 = n3583 & n3584 ;
  assign n3586 = ~n1318 & ~n1336 ;
  assign n3587 = ~n1374 & ~n1427 ;
  assign n3588 = ~n1356 & ~n1403 ;
  assign n3589 = n3587 & n3588 ;
  assign n3590 = n3586 & n3589 ;
  assign n3591 = ~n1062 & n3590 ;
  assign n3592 = ~n1038 & n3591 ;
  assign n3593 = n3585 & n3592 ;
  assign n3594 = ~n1006 & n3593 ;
  assign n3595 = ~n945 & ~n978 ;
  assign n3596 = ~n887 & n3595 ;
  assign n3597 = n3594 & n3596 ;
  assign n3599 = ~n831 & n3597 ;
  assign n3566 = ~\P1_B_reg/NET0131  & ~n537 ;
  assign n3567 = ~n538 & ~n3566 ;
  assign n3598 = n831 & ~n3597 ;
  assign n3600 = ~n3567 & ~n3598 ;
  assign n3601 = ~n3599 & n3600 ;
  assign n3602 = ~n3565 & ~n3601 ;
  assign n3603 = n3466 & ~n3602 ;
  assign n3604 = ~n3467 & ~n3603 ;
  assign n3605 = n1936 & ~n3604 ;
  assign n3606 = ~n1299 & ~n1337 ;
  assign n3607 = ~n1319 & ~n1700 ;
  assign n3608 = n3606 & n3607 ;
  assign n3609 = ~n1063 & ~n1697 ;
  assign n3610 = ~n1299 & ~n3609 ;
  assign n3611 = ~n3608 & ~n3610 ;
  assign n3612 = ~n1010 & ~n1039 ;
  assign n3613 = ~n979 & n3612 ;
  assign n3614 = ~n3611 & n3613 ;
  assign n3615 = ~n1010 & ~n1889 ;
  assign n3616 = ~n979 & n3615 ;
  assign n3617 = n1892 & ~n3616 ;
  assign n3618 = ~n3614 & n3617 ;
  assign n3619 = ~n950 & ~n3618 ;
  assign n3620 = ~n1375 & ~n1428 ;
  assign n3621 = ~n1404 & ~n1453 ;
  assign n3622 = n3620 & n3621 ;
  assign n3623 = ~n1095 & ~n1476 ;
  assign n3624 = ~n1119 & ~n1147 ;
  assign n3625 = n3623 & n3624 ;
  assign n3626 = n3622 & n3625 ;
  assign n3627 = ~n1209 & ~n1290 ;
  assign n3628 = ~n1234 & ~n1286 ;
  assign n3629 = n3627 & n3628 ;
  assign n3630 = ~n1175 & ~n1208 ;
  assign n3631 = ~n1290 & ~n3630 ;
  assign n3632 = ~n3629 & ~n3631 ;
  assign n3633 = ~n1673 & n1899 ;
  assign n3634 = n1634 & ~n3633 ;
  assign n3635 = n1897 & ~n3634 ;
  assign n3636 = ~n1587 & ~n3635 ;
  assign n3637 = ~n1538 & ~n1563 ;
  assign n3638 = ~n1282 & ~n1515 ;
  assign n3639 = n3637 & n3638 ;
  assign n3640 = n3636 & n3639 ;
  assign n3641 = ~n1538 & ~n1896 ;
  assign n3642 = n3638 & n3641 ;
  assign n3643 = ~n1481 & ~n1688 ;
  assign n3644 = ~n1282 & ~n3643 ;
  assign n3645 = ~n3642 & ~n3644 ;
  assign n3646 = ~n3640 & n3645 ;
  assign n3647 = ~n1234 & ~n1258 ;
  assign n3648 = n3627 & n3647 ;
  assign n3649 = ~n3646 & n3648 ;
  assign n3650 = n3632 & ~n3649 ;
  assign n3651 = n3626 & ~n3650 ;
  assign n3652 = ~n1119 & ~n1292 ;
  assign n3653 = n3623 & n3652 ;
  assign n3654 = ~n1180 & ~n1712 ;
  assign n3655 = ~n1476 & ~n3654 ;
  assign n3656 = ~n3653 & ~n3655 ;
  assign n3657 = n3622 & ~n3656 ;
  assign n3658 = ~n1404 & ~n1916 ;
  assign n3659 = n3620 & n3658 ;
  assign n3660 = ~n1375 & n1716 ;
  assign n3661 = ~n1704 & ~n3660 ;
  assign n3662 = ~n3659 & n3661 ;
  assign n3663 = ~n3657 & n3662 ;
  assign n3664 = ~n3651 & n3663 ;
  assign n3665 = ~n1319 & ~n1357 ;
  assign n3666 = n3606 & n3665 ;
  assign n3667 = ~n950 & n3613 ;
  assign n3668 = n3666 & n3667 ;
  assign n3669 = ~n3664 & n3668 ;
  assign n3670 = ~n3619 & ~n3669 ;
  assign n3671 = ~n1832 & n3670 ;
  assign n3672 = n1832 & ~n3670 ;
  assign n3673 = ~n3671 & ~n3672 ;
  assign n3674 = n3466 & n3673 ;
  assign n3675 = ~n3467 & ~n3674 ;
  assign n3676 = n501 & n1888 ;
  assign n3677 = ~n1877 & ~n3676 ;
  assign n3678 = ~n3675 & ~n3677 ;
  assign n3725 = ~n3605 & ~n3678 ;
  assign n3726 = n3724 & n3725 ;
  assign n3727 = n3450 & ~n3726 ;
  assign n3728 = ~n3449 & ~n3727 ;
  assign n3729 = \P1_state_reg[0]/NET0131  & ~n3728 ;
  assign n3730 = ~n3436 & ~n3729 ;
  assign n3731 = \P2_reg1_reg[29]/NET0131  & ~n1983 ;
  assign n3732 = \P2_reg1_reg[29]/NET0131  & n2024 ;
  assign n3733 = n2035 & ~n2039 ;
  assign n3734 = \P2_reg1_reg[29]/NET0131  & ~n3733 ;
  assign n3735 = ~n3161 & n3733 ;
  assign n3736 = ~n3734 & ~n3735 ;
  assign n3737 = ~n3177 & ~n3736 ;
  assign n3738 = n3315 & n3733 ;
  assign n3739 = ~n3734 & ~n3738 ;
  assign n3740 = ~n3320 & ~n3739 ;
  assign n3741 = ~n3414 & n3733 ;
  assign n3742 = n3358 & ~n3733 ;
  assign n3743 = n3421 & ~n3742 ;
  assign n3744 = ~n3167 & ~n3172 ;
  assign n3745 = n3353 & n3744 ;
  assign n3746 = ~n3733 & n3745 ;
  assign n3747 = n3743 & ~n3746 ;
  assign n3748 = \P2_reg1_reg[29]/NET0131  & ~n3747 ;
  assign n3749 = ~n3741 & ~n3748 ;
  assign n3750 = ~n3740 & n3749 ;
  assign n3751 = ~n3737 & n3750 ;
  assign n3752 = n2026 & ~n3751 ;
  assign n3753 = ~n3732 & ~n3752 ;
  assign n3754 = \P1_state_reg[0]/NET0131  & ~n3753 ;
  assign n3755 = ~n3731 & ~n3754 ;
  assign n3756 = \P2_reg2_reg[29]/NET0131  & ~n1983 ;
  assign n3757 = \P2_reg2_reg[29]/NET0131  & n2024 ;
  assign n3758 = ~n2035 & n2039 ;
  assign n3759 = \P2_reg2_reg[29]/NET0131  & ~n3758 ;
  assign n3760 = ~n3161 & n3758 ;
  assign n3761 = ~n3759 & ~n3760 ;
  assign n3762 = ~n3177 & ~n3761 ;
  assign n3763 = n3315 & n3758 ;
  assign n3764 = ~n3759 & ~n3763 ;
  assign n3765 = ~n3320 & ~n3764 ;
  assign n3766 = n3352 & n3758 ;
  assign n3767 = ~n3759 & ~n3766 ;
  assign n3768 = n3355 & ~n3767 ;
  assign n3769 = ~n3409 & n3758 ;
  assign n3770 = ~n3759 & ~n3769 ;
  assign n3771 = n3411 & ~n3770 ;
  assign n3772 = n3359 & n3758 ;
  assign n3773 = n3358 & ~n3758 ;
  assign n3774 = ~n3417 & ~n3773 ;
  assign n3775 = \P2_reg2_reg[29]/NET0131  & ~n3774 ;
  assign n3776 = n2241 & n3420 ;
  assign n3777 = ~n3775 & ~n3776 ;
  assign n3778 = ~n3772 & n3777 ;
  assign n3779 = ~n3771 & n3778 ;
  assign n3780 = ~n3768 & n3779 ;
  assign n3781 = ~n3765 & n3780 ;
  assign n3782 = ~n3762 & n3781 ;
  assign n3783 = n2026 & ~n3782 ;
  assign n3784 = ~n3757 & ~n3783 ;
  assign n3785 = \P1_state_reg[0]/NET0131  & ~n3784 ;
  assign n3786 = ~n3756 & ~n3785 ;
  assign n3787 = n2024 & ~n2958 ;
  assign n3788 = ~n2035 & ~n2039 ;
  assign n3789 = ~n2958 & ~n3788 ;
  assign n3854 = ~n3201 & ~n3207 ;
  assign n3855 = ~n3195 & ~n3202 ;
  assign n3856 = ~n3183 & ~n3855 ;
  assign n3857 = ~n3182 & n3856 ;
  assign n3858 = n3854 & ~n3857 ;
  assign n3859 = ~n3180 & ~n3858 ;
  assign n3790 = ~n3183 & ~n3187 ;
  assign n3791 = ~n3180 & ~n3182 ;
  assign n3792 = n3790 & n3791 ;
  assign n3793 = ~n3186 & ~n3189 ;
  assign n3794 = ~n3211 & ~n3305 ;
  assign n3795 = n3793 & n3794 ;
  assign n3796 = n3792 & n3795 ;
  assign n3814 = ~n3239 & ~n3242 ;
  assign n3815 = ~n3225 & ~n3229 ;
  assign n3816 = n3814 & n3815 ;
  assign n3817 = ~n3241 & ~n3244 ;
  assign n3818 = ~n3264 & ~n3272 ;
  assign n3819 = ~n3255 & ~n3259 ;
  assign n3820 = n3263 & ~n3819 ;
  assign n3821 = ~n3254 & ~n3268 ;
  assign n3822 = ~n3262 & ~n3821 ;
  assign n3823 = ~n3820 & ~n3822 ;
  assign n3824 = n3818 & ~n3823 ;
  assign n3825 = n3267 & ~n3272 ;
  assign n3826 = ~n3246 & ~n3825 ;
  assign n3827 = ~n3824 & n3826 ;
  assign n3828 = n3817 & ~n3827 ;
  assign n3829 = ~n3245 & ~n3251 ;
  assign n3830 = ~n3241 & ~n3829 ;
  assign n3831 = ~n3828 & ~n3830 ;
  assign n3832 = n3816 & ~n3831 ;
  assign n3833 = ~n3230 & ~n3250 ;
  assign n3834 = ~n3239 & ~n3833 ;
  assign n3835 = n3815 & n3834 ;
  assign n3836 = ~n3228 & ~n3235 ;
  assign n3837 = ~n3225 & ~n3836 ;
  assign n3838 = ~n3835 & ~n3837 ;
  assign n3839 = ~n3832 & n3838 ;
  assign n3797 = ~n3210 & ~n3214 ;
  assign n3798 = ~n3213 & ~n3217 ;
  assign n3799 = n3797 & n3798 ;
  assign n3800 = ~n3218 & ~n3220 ;
  assign n3840 = ~n3221 & ~n3226 ;
  assign n3841 = n3800 & n3840 ;
  assign n3842 = n3799 & n3841 ;
  assign n3843 = ~n3839 & n3842 ;
  assign n3801 = ~n3234 & ~n3283 ;
  assign n3802 = ~n3221 & ~n3801 ;
  assign n3803 = n3800 & n3802 ;
  assign n3804 = ~n3282 & ~n3288 ;
  assign n3805 = ~n3218 & ~n3804 ;
  assign n3806 = ~n3803 & ~n3805 ;
  assign n3807 = n3799 & ~n3806 ;
  assign n3808 = ~n3213 & n3287 ;
  assign n3809 = ~n3294 & ~n3808 ;
  assign n3810 = n3797 & ~n3809 ;
  assign n3811 = ~n3210 & n3293 ;
  assign n3812 = ~n3299 & ~n3811 ;
  assign n3813 = ~n3810 & n3812 ;
  assign n3844 = ~n3807 & n3813 ;
  assign n3845 = ~n3843 & n3844 ;
  assign n3846 = n3796 & ~n3845 ;
  assign n3847 = n3298 & ~n3305 ;
  assign n3848 = ~n3191 & ~n3847 ;
  assign n3849 = n3793 & ~n3848 ;
  assign n3850 = ~n3190 & ~n3196 ;
  assign n3851 = ~n3186 & ~n3850 ;
  assign n3852 = ~n3849 & ~n3851 ;
  assign n3853 = n3792 & ~n3852 ;
  assign n3860 = ~n3846 & ~n3853 ;
  assign n3861 = ~n3859 & n3860 ;
  assign n3862 = ~n2963 & ~n3154 ;
  assign n3863 = ~n3861 & n3862 ;
  assign n3864 = n3861 & ~n3862 ;
  assign n3865 = ~n3863 & ~n3864 ;
  assign n3866 = n3788 & ~n3865 ;
  assign n3867 = ~n3789 & ~n3866 ;
  assign n3868 = ~n3320 & ~n3867 ;
  assign n3869 = ~n2705 & ~n2756 ;
  assign n3870 = n2673 & ~n2780 ;
  assign n3871 = ~n2785 & ~n3870 ;
  assign n3872 = n3869 & ~n3871 ;
  assign n3873 = ~n2705 & n2784 ;
  assign n3874 = ~n2790 & ~n3873 ;
  assign n3875 = ~n3872 & n3874 ;
  assign n3876 = ~n2496 & ~n2522 ;
  assign n3877 = n2607 & n2633 ;
  assign n3878 = ~n2567 & ~n2661 ;
  assign n3879 = ~n2632 & ~n3878 ;
  assign n3880 = ~n3877 & ~n3879 ;
  assign n3881 = ~n2545 & ~n2657 ;
  assign n3882 = ~n3880 & n3881 ;
  assign n3883 = ~n2660 & ~n2669 ;
  assign n3884 = ~n2545 & ~n3883 ;
  assign n3885 = ~n3882 & ~n3884 ;
  assign n3886 = n3876 & ~n3885 ;
  assign n3887 = ~n2668 & ~n2674 ;
  assign n3888 = ~n2496 & ~n3887 ;
  assign n3889 = ~n3886 & ~n3888 ;
  assign n3890 = ~n2471 & ~n2780 ;
  assign n3891 = n3869 & n3890 ;
  assign n3892 = ~n3889 & n3891 ;
  assign n3893 = n3875 & ~n3892 ;
  assign n3894 = ~n2844 & ~n2871 ;
  assign n3895 = ~n2732 & ~n2894 ;
  assign n3896 = n3894 & n3895 ;
  assign n3897 = ~n2400 & ~n2819 ;
  assign n3898 = ~n2312 & ~n2443 ;
  assign n3899 = n3897 & n3898 ;
  assign n3900 = n3896 & n3899 ;
  assign n3901 = ~n3893 & n3900 ;
  assign n3902 = ~n2789 & ~n2900 ;
  assign n3903 = ~n2894 & ~n3902 ;
  assign n3904 = n3894 & n3903 ;
  assign n3905 = ~n2899 & ~n2905 ;
  assign n3906 = ~n2844 & ~n3905 ;
  assign n3907 = ~n3904 & ~n3906 ;
  assign n3908 = n3899 & ~n3907 ;
  assign n3909 = ~n2904 & ~n2911 ;
  assign n3910 = ~n2400 & ~n3909 ;
  assign n3911 = n3898 & n3910 ;
  assign n3912 = ~n2312 & n2910 ;
  assign n3913 = ~n2916 & ~n3912 ;
  assign n3914 = ~n3911 & n3913 ;
  assign n3915 = ~n3908 & n3914 ;
  assign n3916 = ~n3901 & n3915 ;
  assign n3917 = ~n3044 & ~n3066 ;
  assign n3918 = ~n2992 & ~n3022 ;
  assign n3919 = n3917 & n3918 ;
  assign n3920 = ~n3089 & ~n3113 ;
  assign n3921 = ~n2369 & ~n3131 ;
  assign n3922 = n3920 & n3921 ;
  assign n3923 = n3919 & n3922 ;
  assign n3924 = ~n3916 & n3923 ;
  assign n3925 = n2915 & ~n3131 ;
  assign n3926 = ~n3139 & ~n3925 ;
  assign n3927 = n3920 & ~n3926 ;
  assign n3928 = ~n3089 & n3138 ;
  assign n3929 = ~n3144 & ~n3928 ;
  assign n3930 = ~n3927 & n3929 ;
  assign n3931 = n3919 & ~n3930 ;
  assign n3932 = ~n3044 & n3143 ;
  assign n3933 = ~n3150 & ~n3932 ;
  assign n3934 = n3918 & ~n3933 ;
  assign n3935 = ~n2992 & n3149 ;
  assign n3936 = ~n3136 & ~n3935 ;
  assign n3937 = ~n3934 & n3936 ;
  assign n3938 = ~n3931 & n3937 ;
  assign n3939 = ~n3924 & n3938 ;
  assign n3940 = n3862 & n3939 ;
  assign n3941 = ~n3862 & ~n3939 ;
  assign n3942 = ~n3940 & ~n3941 ;
  assign n3943 = n3788 & ~n3942 ;
  assign n3944 = ~n3789 & ~n3943 ;
  assign n3945 = ~n3177 & ~n3944 ;
  assign n3946 = n3346 & n3347 ;
  assign n3947 = n2949 & ~n3946 ;
  assign n3948 = ~n3349 & ~n3947 ;
  assign n3949 = n3788 & n3948 ;
  assign n3950 = ~n3789 & ~n3949 ;
  assign n3951 = n3355 & ~n3950 ;
  assign n3952 = n3366 & n3394 ;
  assign n3953 = n2251 & ~n3952 ;
  assign n3954 = ~n3396 & ~n3953 ;
  assign n3955 = ~n2058 & ~n3954 ;
  assign n3956 = n2058 & n2991 ;
  assign n3957 = ~n3955 & ~n3956 ;
  assign n3958 = n3788 & n3957 ;
  assign n3959 = ~n3789 & ~n3958 ;
  assign n3960 = n3411 & ~n3959 ;
  assign n3961 = n3358 & ~n3788 ;
  assign n3962 = ~n3417 & ~n3961 ;
  assign n3963 = ~n2958 & ~n3962 ;
  assign n3964 = n3358 & n3788 ;
  assign n3965 = ~n3420 & ~n3964 ;
  assign n3966 = n2949 & ~n3965 ;
  assign n3967 = ~n3963 & ~n3966 ;
  assign n3968 = ~n3960 & n3967 ;
  assign n3969 = ~n3951 & n3968 ;
  assign n3970 = ~n3945 & n3969 ;
  assign n3971 = ~n3868 & n3970 ;
  assign n3972 = n2026 & ~n3971 ;
  assign n3973 = ~n3787 & ~n3972 ;
  assign n3974 = \P1_state_reg[0]/NET0131  & ~n3973 ;
  assign n3975 = ~\P1_state_reg[0]/NET0131  & \P2_reg3_reg[28]/NET0131  ;
  assign n3976 = \P1_state_reg[0]/NET0131  & n1982 ;
  assign n3977 = ~n2958 & n3976 ;
  assign n3978 = ~n3975 & ~n3977 ;
  assign n3979 = ~n3974 & n3978 ;
  assign n3980 = ~n3460 & ~n3465 ;
  assign n3981 = n941 & ~n3980 ;
  assign n3982 = ~n1774 & ~n3499 ;
  assign n3983 = n3507 & n3510 ;
  assign n3984 = ~n1777 & ~n3515 ;
  assign n3985 = ~n3509 & ~n3984 ;
  assign n3986 = ~n3983 & ~n3985 ;
  assign n3987 = ~n3500 & ~n3511 ;
  assign n3988 = ~n3986 & n3987 ;
  assign n3989 = n3982 & n3988 ;
  assign n3990 = ~n3500 & n3514 ;
  assign n3991 = ~n3522 & ~n3990 ;
  assign n3992 = n3982 & ~n3991 ;
  assign n3993 = ~n1774 & n3521 ;
  assign n3994 = ~n1775 & ~n3993 ;
  assign n3995 = ~n3992 & n3994 ;
  assign n3996 = ~n3989 & n3995 ;
  assign n3997 = ~n1781 & ~n1800 ;
  assign n3998 = ~n1770 & ~n1790 ;
  assign n3999 = n3997 & n3998 ;
  assign n4000 = ~n3996 & n3999 ;
  assign n4001 = ~n1781 & n1801 ;
  assign n4002 = ~n1780 & ~n4001 ;
  assign n4003 = n3998 & ~n4002 ;
  assign n4004 = ~n1771 & ~n1789 ;
  assign n4005 = ~n1770 & ~n4004 ;
  assign n4006 = ~n4003 & ~n4005 ;
  assign n4007 = ~n4000 & n4006 ;
  assign n4008 = ~n1794 & ~n1797 ;
  assign n4009 = ~n1786 & ~n1813 ;
  assign n4010 = n4008 & n4009 ;
  assign n4011 = ~n1783 & ~n3485 ;
  assign n4012 = ~n1822 & ~n1833 ;
  assign n4013 = n4011 & n4012 ;
  assign n4014 = n4010 & n4013 ;
  assign n4015 = ~n4007 & n4014 ;
  assign n4016 = n1795 & ~n1797 ;
  assign n4017 = ~n1798 & ~n4016 ;
  assign n4018 = n4009 & ~n4017 ;
  assign n4019 = ~n1786 & n1814 ;
  assign n4020 = ~n1787 & ~n4019 ;
  assign n4021 = ~n4018 & n4020 ;
  assign n4022 = n4013 & ~n4021 ;
  assign n4023 = ~n1784 & ~n3542 ;
  assign n4024 = ~n3485 & ~n4023 ;
  assign n4025 = n4012 & n4024 ;
  assign n4026 = ~n1823 & ~n1834 ;
  assign n4027 = ~n1833 & ~n4026 ;
  assign n4028 = ~n4025 & ~n4027 ;
  assign n4029 = ~n4022 & n4028 ;
  assign n4030 = ~n4015 & n4029 ;
  assign n4031 = ~n1820 & ~n1836 ;
  assign n4032 = ~n1826 & ~n1839 ;
  assign n4033 = n4031 & n4032 ;
  assign n4034 = ~n1816 & n3476 ;
  assign n4035 = n4033 & n4034 ;
  assign n4036 = ~n4030 & n4035 ;
  assign n4038 = n1827 & ~n1839 ;
  assign n4039 = ~n1840 & ~n4038 ;
  assign n4040 = n4031 & ~n4039 ;
  assign n4041 = ~n1820 & n1837 ;
  assign n4042 = ~n1819 & ~n4041 ;
  assign n4043 = ~n4040 & n4042 ;
  assign n4044 = n4034 & ~n4043 ;
  assign n4045 = ~n1811 & ~n1817 ;
  assign n4046 = n3476 & ~n4045 ;
  assign n4037 = ~n1767 & n1807 ;
  assign n4047 = ~n1768 & ~n4037 ;
  assign n4048 = ~n4046 & n4047 ;
  assign n4049 = ~n4044 & n4048 ;
  assign n4050 = ~n4036 & n4049 ;
  assign n4051 = n1831 & n4050 ;
  assign n4052 = ~n1831 & ~n4050 ;
  assign n4053 = ~n4051 & ~n4052 ;
  assign n4054 = n3980 & ~n4053 ;
  assign n4055 = ~n3981 & ~n4054 ;
  assign n4056 = ~n3563 & ~n4055 ;
  assign n4057 = ~n969 & n3704 ;
  assign n4058 = n933 & ~n4057 ;
  assign n4059 = ~n3706 & ~n4058 ;
  assign n4060 = n3980 & n4059 ;
  assign n4061 = ~n3981 & ~n4060 ;
  assign n4062 = n3712 & ~n4061 ;
  assign n4063 = n1880 & ~n3980 ;
  assign n4064 = ~n3716 & ~n4063 ;
  assign n4065 = n941 & ~n4064 ;
  assign n4066 = n1880 & n3980 ;
  assign n4067 = ~n1763 & ~n4066 ;
  assign n4068 = n933 & ~n4067 ;
  assign n4105 = ~n4065 & ~n4068 ;
  assign n4106 = ~n4062 & n4105 ;
  assign n4107 = ~n4056 & n4106 ;
  assign n4069 = ~n1207 & n3580 ;
  assign n4070 = ~n1174 & n4069 ;
  assign n4071 = ~n1146 & n3569 ;
  assign n4072 = ~n1475 & n4071 ;
  assign n4073 = n4070 & n4072 ;
  assign n4074 = ~n1452 & n3591 ;
  assign n4075 = n4073 & n4074 ;
  assign n4076 = ~n1006 & ~n1038 ;
  assign n4077 = n3595 & n4076 ;
  assign n4078 = n4075 & n4077 ;
  assign n4079 = ~n887 & ~n4078 ;
  assign n4080 = n887 & n4078 ;
  assign n4081 = ~n4079 & ~n4080 ;
  assign n4082 = ~n537 & ~n4081 ;
  assign n4083 = n537 & ~n978 ;
  assign n4084 = ~n4082 & ~n4083 ;
  assign n4085 = n3980 & ~n4084 ;
  assign n4086 = ~n3981 & ~n4085 ;
  assign n4087 = n1936 & ~n4086 ;
  assign n4088 = n1487 & ~n1748 ;
  assign n4089 = n1478 & n1480 ;
  assign n4090 = ~n4088 & n4089 ;
  assign n4091 = ~n1183 & n1478 ;
  assign n4092 = n1720 & ~n4091 ;
  assign n4093 = ~n4090 & n4092 ;
  assign n4094 = n1301 & n1377 ;
  assign n4095 = ~n4093 & n4094 ;
  assign n4096 = n1301 & ~n1710 ;
  assign n4097 = ~n1069 & ~n4096 ;
  assign n4098 = ~n4095 & n4097 ;
  assign n4099 = n1831 & ~n4098 ;
  assign n4100 = ~n1831 & n4098 ;
  assign n4101 = ~n4099 & ~n4100 ;
  assign n4102 = n3980 & ~n4101 ;
  assign n4103 = ~n3981 & ~n4102 ;
  assign n4104 = ~n3677 & ~n4103 ;
  assign n4108 = ~n4087 & ~n4104 ;
  assign n4109 = n4107 & n4108 ;
  assign n4110 = n3450 & ~n4109 ;
  assign n4111 = n941 & n3448 ;
  assign n4112 = ~n4110 & ~n4111 ;
  assign n4113 = \P1_state_reg[0]/NET0131  & ~n4112 ;
  assign n4114 = \P1_reg3_reg[28]/NET0131  & ~\P1_state_reg[0]/NET0131  ;
  assign n4115 = n941 & n1953 ;
  assign n4116 = ~n4114 & ~n4115 ;
  assign n4117 = ~n4113 & n4116 ;
  assign n4118 = ~n3419 & n3976 ;
  assign n4119 = \P2_B_reg/NET0131  & ~n4118 ;
  assign n4120 = ~\P1_datao_reg[30]/NET0131  & ~\si[30]_pad  ;
  assign n4121 = ~n2062 & ~n2064 ;
  assign n4122 = ~n2072 & n4121 ;
  assign n4123 = ~n4120 & n4122 ;
  assign n4124 = n2968 & n4123 ;
  assign n4125 = ~n3073 & n4124 ;
  assign n4129 = ~n2967 & n4123 ;
  assign n4126 = ~n2172 & n4121 ;
  assign n4127 = ~n2061 & ~n4126 ;
  assign n4128 = ~n4120 & ~n4127 ;
  assign n4130 = \P1_datao_reg[30]/NET0131  & \si[30]_pad  ;
  assign n4131 = ~n4128 & ~n4130 ;
  assign n4132 = ~n4129 & n4131 ;
  assign n4133 = ~n4125 & n4132 ;
  assign n4135 = ~\si[31]_pad  & n4133 ;
  assign n4134 = \si[31]_pad  & ~n4133 ;
  assign n4136 = n543 & ~n4134 ;
  assign n4137 = ~n4135 & n4136 ;
  assign n4138 = \P1_datao_reg[31]/NET0131  & n4137 ;
  assign n4139 = ~\P1_datao_reg[31]/NET0131  & ~n4137 ;
  assign n4140 = ~n4138 & ~n4139 ;
  assign n4141 = ~n2059 & n4140 ;
  assign n4142 = \P1_datao_reg[30]/NET0131  & ~n543 ;
  assign n4143 = ~n4120 & ~n4130 ;
  assign n4145 = ~n2073 & n4122 ;
  assign n4148 = n2999 & n4145 ;
  assign n4149 = ~n3096 & n4148 ;
  assign n4146 = ~n2998 & n4145 ;
  assign n4147 = ~n2924 & n4122 ;
  assign n4144 = ~n2062 & n2171 ;
  assign n4150 = ~n2061 & ~n4144 ;
  assign n4151 = ~n4147 & n4150 ;
  assign n4152 = ~n4146 & n4151 ;
  assign n4153 = ~n4149 & n4152 ;
  assign n4155 = ~n4143 & n4153 ;
  assign n4154 = n4143 & ~n4153 ;
  assign n4156 = n543 & ~n4154 ;
  assign n4157 = ~n4155 & n4156 ;
  assign n4158 = ~n4142 & ~n4157 ;
  assign n4159 = ~n2059 & ~n4158 ;
  assign n4160 = ~n3402 & ~n4159 ;
  assign n4161 = ~n3372 & ~n4160 ;
  assign n4162 = n4141 & ~n4161 ;
  assign n4163 = ~n2253 & ~n3206 ;
  assign n4164 = ~n2252 & ~n4163 ;
  assign n4165 = ~n2252 & ~n3179 ;
  assign n4166 = ~n3838 & n3841 ;
  assign n4167 = n3806 & ~n4166 ;
  assign n4168 = n3832 & n3841 ;
  assign n4169 = n4167 & ~n4168 ;
  assign n4170 = n3799 & ~n4169 ;
  assign n4171 = n3796 & n4170 ;
  assign n4172 = n3795 & ~n3813 ;
  assign n4173 = n3852 & ~n4172 ;
  assign n4174 = n3792 & ~n4173 ;
  assign n4175 = ~n3859 & ~n4174 ;
  assign n4176 = ~n4171 & n4175 ;
  assign n4177 = n4165 & ~n4176 ;
  assign n4178 = ~n4164 & ~n4177 ;
  assign n4179 = ~n3372 & ~n4141 ;
  assign n4180 = ~n3372 & ~n3402 ;
  assign n4181 = n4159 & ~n4180 ;
  assign n4182 = ~n4179 & ~n4181 ;
  assign n4183 = ~n4178 & n4182 ;
  assign n4184 = ~n4162 & ~n4183 ;
  assign n4186 = n3175 & ~n4184 ;
  assign n4185 = ~n3175 & n4184 ;
  assign n4187 = n3166 & ~n3170 ;
  assign n4188 = ~n4185 & n4187 ;
  assign n4189 = ~n4186 & n4188 ;
  assign n4222 = n3372 & n4141 ;
  assign n4220 = n3402 & n4159 ;
  assign n4221 = ~n4179 & ~n4220 ;
  assign n4261 = ~n2253 & ~n4160 ;
  assign n4262 = ~n4165 & n4261 ;
  assign n4263 = n4221 & ~n4262 ;
  assign n4264 = ~n4222 & ~n4263 ;
  assign n4223 = ~n4160 & ~n4222 ;
  assign n4265 = n4163 & n4223 ;
  assign n4266 = n3854 & n3855 ;
  assign n4267 = n4265 & n4266 ;
  assign n4268 = n3816 & n3841 ;
  assign n4269 = n4167 & ~n4268 ;
  assign n4203 = ~n2597 & n2604 ;
  assign n4270 = ~n3257 & n4203 ;
  assign n4271 = n3256 & ~n4270 ;
  assign n4272 = n3263 & ~n4271 ;
  assign n4273 = n3269 & ~n4272 ;
  assign n4274 = n3818 & ~n4273 ;
  assign n4275 = n3247 & ~n4274 ;
  assign n4276 = n3817 & ~n4275 ;
  assign n4277 = ~n3251 & n3833 ;
  assign n4278 = n3836 & n4277 ;
  assign n4279 = n3801 & n4278 ;
  assign n4280 = n3804 & n4279 ;
  assign n4281 = ~n4276 & n4280 ;
  assign n4282 = ~n4269 & ~n4281 ;
  assign n4283 = ~n3191 & n3300 ;
  assign n4284 = n3850 & n4283 ;
  assign n4285 = ~n3287 & n3295 ;
  assign n4286 = n4284 & n4285 ;
  assign n4287 = ~n4282 & n4286 ;
  assign n4288 = n4267 & n4287 ;
  assign n4301 = ~n4264 & ~n4288 ;
  assign n4289 = n3192 & ~n3794 ;
  assign n4290 = n3793 & ~n4289 ;
  assign n4291 = ~n3196 & ~n4290 ;
  assign n4292 = n3295 & ~n3798 ;
  assign n4293 = n3797 & ~n4292 ;
  assign n4294 = n4284 & ~n4293 ;
  assign n4295 = ~n4291 & ~n4294 ;
  assign n4296 = n4267 & ~n4295 ;
  assign n4297 = n3203 & ~n3790 ;
  assign n4298 = n3791 & ~n4297 ;
  assign n4299 = ~n3207 & n4265 ;
  assign n4300 = ~n4298 & n4299 ;
  assign n4302 = ~n4296 & ~n4300 ;
  assign n4303 = n4301 & n4302 ;
  assign n4311 = n3175 & n4303 ;
  assign n4310 = ~n3175 & ~n4303 ;
  assign n4312 = n3171 & ~n4310 ;
  assign n4313 = ~n4311 & n4312 ;
  assign n4190 = \P2_B_reg/NET0131  & n1982 ;
  assign n4219 = ~n2992 & ~n3136 ;
  assign n4251 = ~n4219 & n4221 ;
  assign n4252 = n4223 & n4251 ;
  assign n4192 = ~n2894 & ~n2900 ;
  assign n4198 = ~n3230 & ~n3239 ;
  assign n4195 = ~n3228 & ~n3229 ;
  assign n4206 = ~n2657 & ~n2660 ;
  assign n4204 = ~n3258 & ~n4203 ;
  assign n4205 = ~n2522 & ~n2668 ;
  assign n4226 = n4204 & ~n4205 ;
  assign n4227 = ~n4206 & n4226 ;
  assign n4231 = n4195 & n4227 ;
  assign n4232 = n4198 & n4231 ;
  assign n4235 = ~n4192 & n4232 ;
  assign n4210 = ~n2871 & ~n2899 ;
  assign n4211 = ~n2819 & ~n2904 ;
  assign n4236 = ~n4210 & ~n4211 ;
  assign n4237 = n4235 & n4236 ;
  assign n4191 = ~n2400 & ~n2911 ;
  assign n4212 = ~n2732 & ~n2789 ;
  assign n4201 = ~n2705 & ~n2790 ;
  assign n4193 = ~n3262 & ~n3268 ;
  assign n4194 = ~n3246 & ~n3272 ;
  assign n4224 = n4193 & n4194 ;
  assign n4199 = ~n3255 & ~n3257 ;
  assign n4202 = ~n2567 & ~n2609 ;
  assign n4225 = n4199 & ~n4202 ;
  assign n4228 = n4224 & n4225 ;
  assign n4207 = ~n2496 & ~n2674 ;
  assign n4208 = ~n2471 & ~n2673 ;
  assign n4229 = ~n4207 & ~n4208 ;
  assign n4230 = n4228 & n4229 ;
  assign n4233 = ~n4201 & n4230 ;
  assign n4234 = ~n4212 & n4233 ;
  assign n4238 = ~n4191 & n4234 ;
  assign n4242 = n4237 & n4238 ;
  assign n4196 = ~n3089 & ~n3144 ;
  assign n4197 = ~n2312 & ~n2916 ;
  assign n4243 = ~n4196 & ~n4197 ;
  assign n4244 = n4242 & n4243 ;
  assign n4247 = n2254 & n4244 ;
  assign n4213 = ~n3044 & ~n3150 ;
  assign n4214 = ~n3022 & ~n3149 ;
  assign n4248 = ~n4213 & ~n4214 ;
  assign n4249 = n4247 & n4248 ;
  assign n4209 = ~n3113 & ~n3138 ;
  assign n4200 = ~n3066 & ~n3143 ;
  assign n4215 = ~n2844 & ~n2905 ;
  assign n4216 = ~n3131 & ~n3139 ;
  assign n4239 = ~n4215 & ~n4216 ;
  assign n4217 = ~n2369 & ~n2915 ;
  assign n4218 = ~n2443 & ~n2910 ;
  assign n4240 = ~n4217 & ~n4218 ;
  assign n4241 = n4239 & n4240 ;
  assign n4245 = ~n4200 & n4241 ;
  assign n4246 = ~n4209 & n4245 ;
  assign n4250 = ~n3862 & n4246 ;
  assign n4253 = n4249 & n4250 ;
  assign n4254 = n4252 & n4253 ;
  assign n4256 = n3175 & ~n4254 ;
  assign n4255 = ~n3175 & n4254 ;
  assign n4257 = ~n3166 & ~n4255 ;
  assign n4258 = ~n4256 & n4257 ;
  assign n4259 = ~n4190 & ~n4258 ;
  assign n4260 = ~n3170 & ~n4259 ;
  assign n4304 = ~\P2_B_reg/NET0131  & ~n4303 ;
  assign n4305 = n3410 & n3418 ;
  assign n4306 = ~n4304 & n4305 ;
  assign n4307 = n3411 & ~n4303 ;
  assign n4308 = ~n3176 & ~n3411 ;
  assign n4309 = \P2_B_reg/NET0131  & ~n4308 ;
  assign n4319 = ~n4307 & ~n4309 ;
  assign n4320 = ~n4306 & n4319 ;
  assign n4321 = ~n4260 & n4320 ;
  assign n4322 = ~n4313 & n4321 ;
  assign n4314 = ~n4264 & ~n4265 ;
  assign n4315 = n4177 & n4221 ;
  assign n4316 = ~n4314 & ~n4315 ;
  assign n4317 = n3354 & n4316 ;
  assign n4318 = n3419 & ~n4316 ;
  assign n4323 = ~n4317 & ~n4318 ;
  assign n4324 = n4322 & n4323 ;
  assign n4325 = ~n4189 & n4324 ;
  assign n4326 = n3976 & ~n4325 ;
  assign n4327 = ~n4119 & ~n4326 ;
  assign n4328 = \P2_reg0_reg[28]/NET0131  & ~n1983 ;
  assign n4329 = \P2_reg0_reg[28]/NET0131  & n2024 ;
  assign n4330 = \P2_reg0_reg[28]/NET0131  & ~n2040 ;
  assign n4331 = n2040 & ~n3865 ;
  assign n4332 = ~n4330 & ~n4331 ;
  assign n4333 = ~n3320 & ~n4332 ;
  assign n4334 = n2040 & ~n3942 ;
  assign n4335 = ~n4330 & ~n4334 ;
  assign n4336 = ~n3177 & ~n4335 ;
  assign n4337 = n3355 & n3948 ;
  assign n4338 = n2949 & n3358 ;
  assign n4339 = n3411 & n3957 ;
  assign n4340 = ~n4338 & ~n4339 ;
  assign n4341 = ~n4337 & n4340 ;
  assign n4342 = n2040 & ~n4341 ;
  assign n4343 = \P2_reg0_reg[28]/NET0131  & ~n3426 ;
  assign n4344 = ~n4342 & ~n4343 ;
  assign n4345 = ~n4336 & n4344 ;
  assign n4346 = ~n4333 & n4345 ;
  assign n4347 = n2026 & ~n4346 ;
  assign n4348 = ~n4329 & ~n4347 ;
  assign n4349 = \P1_state_reg[0]/NET0131  & ~n4348 ;
  assign n4350 = ~n4328 & ~n4349 ;
  assign n4351 = \P2_reg1_reg[28]/NET0131  & ~n1983 ;
  assign n4352 = \P2_reg1_reg[28]/NET0131  & n2024 ;
  assign n4353 = \P2_reg1_reg[28]/NET0131  & ~n3733 ;
  assign n4354 = n3733 & ~n3865 ;
  assign n4355 = ~n4353 & ~n4354 ;
  assign n4356 = ~n3320 & ~n4355 ;
  assign n4357 = n3733 & ~n3942 ;
  assign n4358 = ~n4353 & ~n4357 ;
  assign n4359 = ~n3177 & ~n4358 ;
  assign n4360 = n3733 & ~n4341 ;
  assign n4361 = \P2_reg1_reg[28]/NET0131  & ~n3747 ;
  assign n4362 = ~n4360 & ~n4361 ;
  assign n4363 = ~n4359 & n4362 ;
  assign n4364 = ~n4356 & n4363 ;
  assign n4365 = n2026 & ~n4364 ;
  assign n4366 = ~n4352 & ~n4365 ;
  assign n4367 = \P1_state_reg[0]/NET0131  & ~n4366 ;
  assign n4368 = ~n4351 & ~n4367 ;
  assign n4369 = \P2_reg2_reg[28]/NET0131  & ~n1983 ;
  assign n4370 = \P2_reg2_reg[28]/NET0131  & n2024 ;
  assign n4371 = \P2_reg2_reg[28]/NET0131  & ~n3758 ;
  assign n4372 = n3758 & ~n3865 ;
  assign n4373 = ~n4371 & ~n4372 ;
  assign n4374 = ~n3320 & ~n4373 ;
  assign n4375 = n3758 & ~n3942 ;
  assign n4376 = ~n4371 & ~n4375 ;
  assign n4377 = ~n3177 & ~n4376 ;
  assign n4378 = n3758 & ~n4341 ;
  assign n4379 = ~n2958 & n3420 ;
  assign n4380 = n3411 & ~n3758 ;
  assign n4381 = n3354 & ~n3758 ;
  assign n4382 = ~n1982 & n4381 ;
  assign n4383 = n3774 & ~n4382 ;
  assign n4384 = ~n4380 & n4383 ;
  assign n4385 = \P2_reg2_reg[28]/NET0131  & ~n4384 ;
  assign n4386 = ~n4379 & ~n4385 ;
  assign n4387 = ~n4378 & n4386 ;
  assign n4388 = ~n4377 & n4387 ;
  assign n4389 = ~n4374 & n4388 ;
  assign n4390 = n2026 & ~n4389 ;
  assign n4391 = ~n4370 & ~n4390 ;
  assign n4392 = \P1_state_reg[0]/NET0131  & ~n4391 ;
  assign n4393 = ~n4369 & ~n4392 ;
  assign n4394 = \P1_reg0_reg[27]/NET0131  & ~n3435 ;
  assign n4395 = \P1_reg0_reg[27]/NET0131  & n3448 ;
  assign n4396 = n3460 & n3465 ;
  assign n4397 = \P1_reg0_reg[27]/NET0131  & ~n4396 ;
  assign n4398 = n3636 & n3637 ;
  assign n4399 = ~n3641 & ~n4398 ;
  assign n4400 = n3638 & n3647 ;
  assign n4401 = ~n4399 & n4400 ;
  assign n4402 = n3644 & n3647 ;
  assign n4403 = ~n3628 & ~n4402 ;
  assign n4404 = ~n4401 & n4403 ;
  assign n4405 = n3621 & n3623 ;
  assign n4406 = n3624 & n3627 ;
  assign n4407 = n4405 & n4406 ;
  assign n4408 = ~n4404 & n4407 ;
  assign n4409 = n3624 & n3631 ;
  assign n4410 = ~n3652 & ~n4409 ;
  assign n4411 = n4405 & ~n4410 ;
  assign n4412 = n3621 & n3655 ;
  assign n4413 = ~n3658 & ~n4412 ;
  assign n4414 = ~n4411 & n4413 ;
  assign n4415 = ~n4408 & n4414 ;
  assign n4416 = n3606 & n3612 ;
  assign n4417 = n3620 & n3665 ;
  assign n4418 = n4416 & n4417 ;
  assign n4419 = ~n4415 & n4418 ;
  assign n4421 = ~n3661 & n3665 ;
  assign n4422 = ~n3607 & ~n4421 ;
  assign n4423 = n4416 & ~n4422 ;
  assign n4420 = n3610 & n3612 ;
  assign n4424 = ~n3615 & ~n4420 ;
  assign n4425 = ~n4423 & n4424 ;
  assign n4426 = ~n4419 & n4425 ;
  assign n4427 = n1769 & ~n4426 ;
  assign n4428 = ~n1769 & n4426 ;
  assign n4429 = ~n4427 & ~n4428 ;
  assign n4430 = n4396 & ~n4429 ;
  assign n4431 = ~n4397 & ~n4430 ;
  assign n4432 = ~n3677 & ~n4431 ;
  assign n4484 = n969 & ~n3704 ;
  assign n4485 = ~n4057 & ~n4484 ;
  assign n4486 = n3712 & n4485 ;
  assign n4487 = n969 & n1880 ;
  assign n4488 = ~n4486 & ~n4487 ;
  assign n4489 = n4396 & ~n4488 ;
  assign n4490 = n3712 & ~n4396 ;
  assign n4491 = ~n1763 & ~n3716 ;
  assign n4492 = n1880 & ~n4396 ;
  assign n4493 = n4491 & ~n4492 ;
  assign n4494 = ~n4490 & n4493 ;
  assign n4495 = \P1_reg0_reg[27]/NET0131  & ~n4494 ;
  assign n4496 = ~n4489 & ~n4495 ;
  assign n4497 = ~n4432 & n4496 ;
  assign n4433 = ~n1810 & n3468 ;
  assign n4434 = ~n3547 & n3551 ;
  assign n4435 = n3470 & ~n4434 ;
  assign n4436 = n4433 & ~n4435 ;
  assign n4437 = ~n1810 & ~n3473 ;
  assign n4438 = n3478 & ~n4437 ;
  assign n4439 = ~n4436 & n4438 ;
  assign n4440 = ~n1808 & ~n4439 ;
  assign n4441 = n3501 & ~n3518 ;
  assign n4442 = n3524 & ~n4441 ;
  assign n4443 = n3502 & n3530 ;
  assign n4444 = ~n4442 & n4443 ;
  assign n4445 = ~n3527 & n3530 ;
  assign n4446 = n3494 & ~n4445 ;
  assign n4447 = ~n4444 & n4446 ;
  assign n4448 = n3488 & n3492 ;
  assign n4449 = n3486 & n3489 ;
  assign n4450 = n4448 & n4449 ;
  assign n4451 = ~n4447 & n4450 ;
  assign n4452 = n3488 & ~n3497 ;
  assign n4453 = n3536 & ~n4452 ;
  assign n4454 = n4449 & ~n4453 ;
  assign n4455 = n3486 & n3539 ;
  assign n4456 = n3544 & ~n4455 ;
  assign n4457 = ~n4454 & n4456 ;
  assign n4458 = ~n4451 & n4457 ;
  assign n4459 = n3484 & n3551 ;
  assign n4460 = ~n1808 & n4459 ;
  assign n4461 = n4433 & n4460 ;
  assign n4462 = ~n4458 & n4461 ;
  assign n4463 = ~n4440 & ~n4462 ;
  assign n4464 = n1769 & n4463 ;
  assign n4465 = ~n1769 & ~n4463 ;
  assign n4466 = ~n4464 & ~n4465 ;
  assign n4467 = n4396 & ~n4466 ;
  assign n4468 = ~n4397 & ~n4467 ;
  assign n4469 = ~n3563 & ~n4468 ;
  assign n4470 = n4070 & n4071 ;
  assign n4471 = n3568 & n3590 ;
  assign n4472 = n4470 & n4471 ;
  assign n4473 = ~n1062 & n4076 ;
  assign n4474 = ~n978 & n4473 ;
  assign n4475 = n4472 & n4474 ;
  assign n4476 = n945 & ~n4475 ;
  assign n4477 = ~n4078 & ~n4476 ;
  assign n4478 = ~n537 & ~n4477 ;
  assign n4479 = n537 & n1006 ;
  assign n4480 = ~n4478 & ~n4479 ;
  assign n4481 = n4396 & n4480 ;
  assign n4482 = ~n4397 & ~n4481 ;
  assign n4483 = n1936 & ~n4482 ;
  assign n4498 = ~n4469 & ~n4483 ;
  assign n4499 = n4497 & n4498 ;
  assign n4500 = n3450 & ~n4499 ;
  assign n4501 = ~n4395 & ~n4500 ;
  assign n4502 = \P1_state_reg[0]/NET0131  & ~n4501 ;
  assign n4503 = ~n4394 & ~n4502 ;
  assign n4504 = \P1_reg0_reg[29]/NET0131  & ~n3435 ;
  assign n4505 = \P1_reg0_reg[29]/NET0131  & n3448 ;
  assign n4506 = \P1_reg0_reg[29]/NET0131  & ~n4396 ;
  assign n4507 = ~n3559 & n4396 ;
  assign n4508 = ~n4506 & ~n4507 ;
  assign n4509 = ~n3563 & ~n4508 ;
  assign n4510 = n3709 & n4396 ;
  assign n4511 = ~n4506 & ~n4510 ;
  assign n4512 = n3712 & ~n4511 ;
  assign n4513 = \P1_reg0_reg[29]/NET0131  & ~n4493 ;
  assign n4514 = n3714 & n4396 ;
  assign n4521 = ~n4513 & ~n4514 ;
  assign n4522 = ~n4512 & n4521 ;
  assign n4523 = ~n4509 & n4522 ;
  assign n4515 = ~n3602 & n4396 ;
  assign n4516 = ~n4506 & ~n4515 ;
  assign n4517 = n1936 & ~n4516 ;
  assign n4518 = n3673 & n4396 ;
  assign n4519 = ~n4506 & ~n4518 ;
  assign n4520 = ~n3677 & ~n4519 ;
  assign n4524 = ~n4517 & ~n4520 ;
  assign n4525 = n4523 & n4524 ;
  assign n4526 = n3450 & ~n4525 ;
  assign n4527 = ~n4505 & ~n4526 ;
  assign n4528 = \P1_state_reg[0]/NET0131  & ~n4527 ;
  assign n4529 = ~n4504 & ~n4528 ;
  assign n4530 = \P1_reg1_reg[29]/NET0131  & ~n3435 ;
  assign n4531 = \P1_reg1_reg[29]/NET0131  & n3448 ;
  assign n4532 = ~n3460 & n3465 ;
  assign n4533 = \P1_reg1_reg[29]/NET0131  & ~n4532 ;
  assign n4534 = ~n3559 & n4532 ;
  assign n4535 = ~n4533 & ~n4534 ;
  assign n4536 = ~n3563 & ~n4535 ;
  assign n4537 = n3709 & n4532 ;
  assign n4538 = ~n4533 & ~n4537 ;
  assign n4539 = n3712 & ~n4538 ;
  assign n4540 = n1880 & ~n4532 ;
  assign n4541 = n4491 & ~n4540 ;
  assign n4542 = \P1_reg1_reg[29]/NET0131  & ~n4541 ;
  assign n4543 = n3714 & n4532 ;
  assign n4550 = ~n4542 & ~n4543 ;
  assign n4551 = ~n4539 & n4550 ;
  assign n4552 = ~n4536 & n4551 ;
  assign n4544 = ~n3602 & n4532 ;
  assign n4545 = ~n4533 & ~n4544 ;
  assign n4546 = n1936 & ~n4545 ;
  assign n4547 = n3673 & n4532 ;
  assign n4548 = ~n4533 & ~n4547 ;
  assign n4549 = ~n3677 & ~n4548 ;
  assign n4553 = ~n4546 & ~n4549 ;
  assign n4554 = n4552 & n4553 ;
  assign n4555 = n3450 & ~n4554 ;
  assign n4556 = ~n4531 & ~n4555 ;
  assign n4557 = \P1_state_reg[0]/NET0131  & ~n4556 ;
  assign n4558 = ~n4530 & ~n4557 ;
  assign n4559 = \P1_reg1_reg[27]/NET0131  & ~n3435 ;
  assign n4560 = \P1_reg1_reg[27]/NET0131  & n3448 ;
  assign n4561 = \P1_reg1_reg[27]/NET0131  & ~n4532 ;
  assign n4562 = ~n4429 & n4532 ;
  assign n4563 = ~n4561 & ~n4562 ;
  assign n4564 = ~n3677 & ~n4563 ;
  assign n4571 = ~n4488 & n4532 ;
  assign n4572 = n3712 & ~n4532 ;
  assign n4573 = n4541 & ~n4572 ;
  assign n4574 = \P1_reg1_reg[27]/NET0131  & ~n4573 ;
  assign n4575 = ~n4571 & ~n4574 ;
  assign n4576 = ~n4564 & n4575 ;
  assign n4565 = ~n4466 & n4532 ;
  assign n4566 = ~n4561 & ~n4565 ;
  assign n4567 = ~n3563 & ~n4566 ;
  assign n4568 = n4480 & n4532 ;
  assign n4569 = ~n4561 & ~n4568 ;
  assign n4570 = n1936 & ~n4569 ;
  assign n4577 = ~n4567 & ~n4570 ;
  assign n4578 = n4576 & n4577 ;
  assign n4579 = n3450 & ~n4578 ;
  assign n4580 = ~n4560 & ~n4579 ;
  assign n4581 = \P1_state_reg[0]/NET0131  & ~n4580 ;
  assign n4582 = ~n4559 & ~n4581 ;
  assign n4585 = n2024 & n3039 ;
  assign n4586 = n3039 & ~n3788 ;
  assign n4602 = n3224 & n3279 ;
  assign n4599 = n3223 & ~n3238 ;
  assign n4600 = n3291 & ~n4599 ;
  assign n4601 = n3216 & ~n4600 ;
  assign n4603 = n3302 & ~n4601 ;
  assign n4604 = ~n4602 & n4603 ;
  assign n4605 = n3307 & ~n4604 ;
  assign n4606 = n3199 & ~n4605 ;
  assign n4607 = n4213 & ~n4606 ;
  assign n4608 = ~n4213 & n4606 ;
  assign n4609 = ~n4607 & ~n4608 ;
  assign n4610 = n3788 & ~n4609 ;
  assign n4611 = ~n4586 & ~n4610 ;
  assign n4612 = ~n3320 & ~n4611 ;
  assign n4587 = ~n2897 & n2908 ;
  assign n4588 = n2445 & n3133 ;
  assign n4589 = ~n4587 & n4588 ;
  assign n4590 = ~n2919 & n3133 ;
  assign n4591 = n3147 & ~n4590 ;
  assign n4592 = ~n4589 & n4591 ;
  assign n4593 = n4213 & n4592 ;
  assign n4594 = ~n4213 & ~n4592 ;
  assign n4595 = ~n4593 & ~n4594 ;
  assign n4596 = n3788 & ~n4595 ;
  assign n4597 = ~n4586 & ~n4596 ;
  assign n4598 = ~n3177 & ~n4597 ;
  assign n4614 = n3325 & n3343 ;
  assign n4615 = ~n3054 & n4614 ;
  assign n4616 = n3034 & ~n4615 ;
  assign n4617 = ~n3346 & ~n4616 ;
  assign n4618 = n3788 & n4617 ;
  assign n4619 = ~n4586 & ~n4618 ;
  assign n4620 = n3355 & ~n4619 ;
  assign n4622 = n3363 & n3394 ;
  assign n4623 = ~n3043 & n4622 ;
  assign n4624 = n3021 & ~n4623 ;
  assign n4625 = n3361 & n4622 ;
  assign n4626 = ~n4624 & ~n4625 ;
  assign n4627 = ~n2058 & ~n4626 ;
  assign n4621 = n2058 & n3065 ;
  assign n4628 = n3411 & ~n4621 ;
  assign n4629 = ~n4627 & n4628 ;
  assign n4630 = n3788 & n4629 ;
  assign n4613 = n3034 & ~n3965 ;
  assign n4631 = n3411 & ~n3788 ;
  assign n4632 = n3962 & ~n4631 ;
  assign n4633 = n3039 & ~n4632 ;
  assign n4634 = ~n4613 & ~n4633 ;
  assign n4635 = ~n4630 & n4634 ;
  assign n4636 = ~n4620 & n4635 ;
  assign n4637 = ~n4598 & n4636 ;
  assign n4638 = ~n4612 & n4637 ;
  assign n4639 = n2026 & ~n4638 ;
  assign n4640 = ~n4585 & ~n4639 ;
  assign n4641 = \P1_state_reg[0]/NET0131  & ~n4640 ;
  assign n4583 = ~\P1_state_reg[0]/NET0131  & \P2_reg3_reg[25]/NET0131  ;
  assign n4584 = n3039 & n3976 ;
  assign n4642 = ~n4583 & ~n4584 ;
  assign n4643 = ~n4641 & n4642 ;
  assign n4646 = n1034 & n3448 ;
  assign n4647 = n1034 & ~n3980 ;
  assign n4686 = n3700 & n3701 ;
  assign n4687 = n1029 & ~n4686 ;
  assign n4688 = ~n1029 & n4686 ;
  assign n4689 = ~n4687 & ~n4688 ;
  assign n4690 = n3980 & n4689 ;
  assign n4691 = ~n4647 & ~n4690 ;
  assign n4692 = n3712 & ~n4691 ;
  assign n4678 = n1006 & ~n3593 ;
  assign n4679 = ~n3594 & ~n4678 ;
  assign n4680 = ~n537 & ~n4679 ;
  assign n4681 = n537 & n1062 ;
  assign n4682 = ~n4680 & ~n4681 ;
  assign n4683 = n3980 & n4682 ;
  assign n4684 = ~n4647 & ~n4683 ;
  assign n4685 = n1936 & ~n4684 ;
  assign n4676 = n1029 & ~n4067 ;
  assign n4677 = n1034 & ~n4064 ;
  assign n4693 = ~n4676 & ~n4677 ;
  assign n4694 = ~n4685 & n4693 ;
  assign n4695 = ~n4692 & n4694 ;
  assign n4648 = n3626 & n3649 ;
  assign n4649 = n3625 & ~n3632 ;
  assign n4650 = n3656 & ~n4649 ;
  assign n4651 = n3622 & ~n4650 ;
  assign n4652 = n3662 & ~n4651 ;
  assign n4653 = ~n4648 & n4652 ;
  assign n4654 = n3666 & ~n4653 ;
  assign n4655 = n3611 & ~n4654 ;
  assign n4656 = n1812 & ~n4655 ;
  assign n4657 = ~n1812 & n4655 ;
  assign n4658 = ~n4656 & ~n4657 ;
  assign n4659 = n3980 & ~n4658 ;
  assign n4660 = ~n4647 & ~n4659 ;
  assign n4661 = ~n3677 & ~n4660 ;
  assign n4662 = n3491 & n3532 ;
  assign n4663 = n3490 & ~n3498 ;
  assign n4664 = n3540 & ~n4663 ;
  assign n4665 = n3487 & ~n4664 ;
  assign n4666 = n3548 & ~n4665 ;
  assign n4667 = ~n4662 & n4666 ;
  assign n4668 = n3552 & ~n4667 ;
  assign n4669 = n3474 & ~n4668 ;
  assign n4670 = n1812 & n4669 ;
  assign n4671 = ~n1812 & ~n4669 ;
  assign n4672 = ~n4670 & ~n4671 ;
  assign n4673 = n3980 & ~n4672 ;
  assign n4674 = ~n4647 & ~n4673 ;
  assign n4675 = ~n3563 & ~n4674 ;
  assign n4696 = ~n4661 & ~n4675 ;
  assign n4697 = n4695 & n4696 ;
  assign n4698 = n3450 & ~n4697 ;
  assign n4699 = ~n4646 & ~n4698 ;
  assign n4700 = \P1_state_reg[0]/NET0131  & ~n4699 ;
  assign n4644 = \P1_reg3_reg[25]/NET0131  & ~\P1_state_reg[0]/NET0131  ;
  assign n4645 = n1034 & n1953 ;
  assign n4701 = ~n4644 & ~n4645 ;
  assign n4702 = ~n4700 & n4701 ;
  assign n4703 = n3017 & ~n3788 ;
  assign n4704 = n3790 & n3793 ;
  assign n4705 = n3814 & n3817 ;
  assign n4706 = ~n3827 & n4705 ;
  assign n4707 = n3814 & n3830 ;
  assign n4708 = ~n3834 & ~n4707 ;
  assign n4709 = ~n4706 & n4708 ;
  assign n4710 = n3815 & n3840 ;
  assign n4711 = ~n4709 & n4710 ;
  assign n4712 = n3837 & n3840 ;
  assign n4713 = ~n3802 & ~n4712 ;
  assign n4714 = ~n4711 & n4713 ;
  assign n4715 = n3798 & n3800 ;
  assign n4716 = ~n4714 & n4715 ;
  assign n4717 = n3798 & n3805 ;
  assign n4718 = n3809 & ~n4717 ;
  assign n4719 = ~n4716 & n4718 ;
  assign n4720 = n3794 & n3797 ;
  assign n4721 = ~n4719 & n4720 ;
  assign n4722 = n4704 & n4721 ;
  assign n4724 = n3794 & ~n3812 ;
  assign n4725 = n3848 & ~n4724 ;
  assign n4726 = n4704 & ~n4725 ;
  assign n4723 = n3790 & n3851 ;
  assign n4727 = ~n3856 & ~n4723 ;
  assign n4728 = ~n4726 & n4727 ;
  assign n4729 = ~n4722 & n4728 ;
  assign n4730 = n4214 & ~n4729 ;
  assign n4731 = ~n4214 & n4729 ;
  assign n4732 = ~n4730 & ~n4731 ;
  assign n4733 = n3788 & ~n4732 ;
  assign n4734 = ~n4703 & ~n4733 ;
  assign n4735 = ~n3320 & ~n4734 ;
  assign n4736 = n3876 & n3890 ;
  assign n4737 = ~n3885 & n4736 ;
  assign n4738 = n3888 & n3890 ;
  assign n4739 = n3871 & ~n4738 ;
  assign n4740 = ~n4737 & n4739 ;
  assign n4741 = n3869 & n3895 ;
  assign n4742 = ~n4740 & n4741 ;
  assign n4743 = ~n3874 & n3895 ;
  assign n4744 = ~n3903 & ~n4743 ;
  assign n4745 = ~n4742 & n4744 ;
  assign n4746 = n3894 & n3897 ;
  assign n4747 = ~n4745 & n4746 ;
  assign n4748 = n3897 & n3906 ;
  assign n4749 = ~n3910 & ~n4748 ;
  assign n4750 = ~n4747 & n4749 ;
  assign n4751 = n3917 & n3920 ;
  assign n4752 = n3898 & n3921 ;
  assign n4753 = n4751 & n4752 ;
  assign n4754 = ~n4750 & n4753 ;
  assign n4756 = ~n3913 & n3921 ;
  assign n4757 = n3926 & ~n4756 ;
  assign n4758 = n4751 & ~n4757 ;
  assign n4755 = n3917 & ~n3929 ;
  assign n4759 = n3933 & ~n4755 ;
  assign n4760 = ~n4758 & n4759 ;
  assign n4761 = ~n4754 & n4760 ;
  assign n4762 = n4214 & n4761 ;
  assign n4763 = ~n4214 & ~n4761 ;
  assign n4764 = ~n4762 & ~n4763 ;
  assign n4765 = n3788 & ~n4764 ;
  assign n4766 = ~n4703 & ~n4765 ;
  assign n4767 = ~n3177 & ~n4766 ;
  assign n4768 = n2991 & ~n4625 ;
  assign n4769 = n3365 & n3394 ;
  assign n4770 = ~n4768 & ~n4769 ;
  assign n4771 = ~n2058 & ~n4770 ;
  assign n4772 = n2058 & n3043 ;
  assign n4773 = ~n4771 & ~n4772 ;
  assign n4774 = n3788 & n4773 ;
  assign n4775 = ~n4703 & ~n4774 ;
  assign n4776 = n3411 & ~n4775 ;
  assign n4777 = n3012 & ~n3346 ;
  assign n4778 = ~n3012 & n3346 ;
  assign n4779 = ~n4777 & ~n4778 ;
  assign n4780 = n3788 & n4779 ;
  assign n4781 = ~n4703 & ~n4780 ;
  assign n4782 = n3355 & ~n4781 ;
  assign n4783 = n3017 & ~n3962 ;
  assign n4784 = n3012 & ~n3965 ;
  assign n4785 = ~n4783 & ~n4784 ;
  assign n4786 = ~n4782 & n4785 ;
  assign n4787 = ~n4776 & n4786 ;
  assign n4788 = ~n4767 & n4787 ;
  assign n4789 = ~n4735 & n4788 ;
  assign n4790 = n2026 & ~n4789 ;
  assign n4791 = n2024 & n3017 ;
  assign n4792 = ~n4790 & ~n4791 ;
  assign n4793 = \P1_state_reg[0]/NET0131  & ~n4792 ;
  assign n4794 = n3017 & n3976 ;
  assign n4795 = ~\P1_state_reg[0]/NET0131  & \P2_reg3_reg[26]/NET0131  ;
  assign n4796 = ~n4794 & ~n4795 ;
  assign n4797 = ~n4793 & n4796 ;
  assign n4798 = n2987 & ~n3788 ;
  assign n4799 = ~n2666 & n2671 ;
  assign n4800 = n2497 & n2781 ;
  assign n4801 = ~n4799 & n4800 ;
  assign n4802 = n2676 & n2781 ;
  assign n4803 = n2787 & ~n4802 ;
  assign n4804 = ~n4801 & n4803 ;
  assign n4805 = n2733 & n2895 ;
  assign n4806 = ~n4804 & n4805 ;
  assign n4807 = n2792 & n2895 ;
  assign n4808 = n2902 & ~n4807 ;
  assign n4809 = ~n4806 & n4808 ;
  assign n4810 = n2444 & n2845 ;
  assign n4811 = ~n4809 & n4810 ;
  assign n4812 = n2444 & ~n2907 ;
  assign n4813 = ~n2913 & ~n4812 ;
  assign n4814 = ~n4811 & n4813 ;
  assign n4815 = n3045 & n3090 ;
  assign n4816 = n2370 & n3132 ;
  assign n4817 = n4815 & n4816 ;
  assign n4818 = ~n4814 & n4817 ;
  assign n4820 = ~n2918 & n3132 ;
  assign n4821 = n3141 & ~n4820 ;
  assign n4822 = n4815 & ~n4821 ;
  assign n4819 = n3045 & ~n3146 ;
  assign n4823 = n3152 & ~n4819 ;
  assign n4824 = ~n4822 & n4823 ;
  assign n4825 = ~n4818 & n4824 ;
  assign n4826 = n4219 & ~n4825 ;
  assign n4827 = ~n4219 & n4825 ;
  assign n4828 = ~n4826 & ~n4827 ;
  assign n4829 = n3788 & n4828 ;
  assign n4830 = ~n4798 & ~n4829 ;
  assign n4831 = ~n3177 & ~n4830 ;
  assign n4868 = n2982 & ~n4778 ;
  assign n4869 = ~n3946 & ~n4868 ;
  assign n4870 = n3788 & n4869 ;
  assign n4871 = ~n4798 & ~n4870 ;
  assign n4872 = n3355 & ~n4871 ;
  assign n4832 = n3266 & n3273 ;
  assign n4833 = n3270 & n3273 ;
  assign n4834 = ~n3248 & ~n4833 ;
  assign n4835 = ~n4832 & n4834 ;
  assign n4836 = n3240 & n3243 ;
  assign n4837 = ~n4835 & n4836 ;
  assign n4838 = n3240 & ~n3253 ;
  assign n4839 = n3232 & ~n4838 ;
  assign n4840 = ~n4837 & n4839 ;
  assign n4841 = n3222 & n3227 ;
  assign n4842 = ~n4840 & n4841 ;
  assign n4843 = n3222 & ~n3237 ;
  assign n4844 = ~n3285 & ~n4843 ;
  assign n4845 = ~n4842 & n4844 ;
  assign n4846 = n3215 & n3219 ;
  assign n4847 = ~n4845 & n4846 ;
  assign n4848 = n3215 & n3290 ;
  assign n4849 = ~n3296 & ~n4848 ;
  assign n4850 = ~n4847 & n4849 ;
  assign n4851 = n3212 & n3306 ;
  assign n4852 = n3184 & n3188 ;
  assign n4853 = n4851 & n4852 ;
  assign n4854 = ~n4850 & n4853 ;
  assign n4855 = n3301 & n3306 ;
  assign n4856 = ~n3193 & ~n4855 ;
  assign n4857 = n4852 & ~n4856 ;
  assign n4858 = n3184 & ~n3198 ;
  assign n4859 = ~n3204 & ~n4858 ;
  assign n4860 = ~n4857 & n4859 ;
  assign n4861 = ~n4854 & n4860 ;
  assign n4862 = n4219 & ~n4861 ;
  assign n4863 = ~n4219 & n4861 ;
  assign n4864 = ~n4862 & ~n4863 ;
  assign n4865 = n3788 & ~n4864 ;
  assign n4866 = ~n4798 & ~n4865 ;
  assign n4867 = ~n3320 & ~n4866 ;
  assign n4873 = n2962 & ~n4769 ;
  assign n4874 = ~n3952 & ~n4873 ;
  assign n4875 = ~n2058 & ~n4874 ;
  assign n4876 = n2058 & n3021 ;
  assign n4877 = ~n4875 & ~n4876 ;
  assign n4878 = n3788 & n4877 ;
  assign n4879 = ~n4798 & ~n4878 ;
  assign n4880 = n3411 & ~n4879 ;
  assign n4881 = n2982 & ~n3965 ;
  assign n4882 = n2987 & ~n3962 ;
  assign n4883 = ~n4881 & ~n4882 ;
  assign n4884 = ~n4880 & n4883 ;
  assign n4885 = ~n4867 & n4884 ;
  assign n4886 = ~n4872 & n4885 ;
  assign n4887 = ~n4831 & n4886 ;
  assign n4888 = n2026 & ~n4887 ;
  assign n4889 = n2024 & n2987 ;
  assign n4890 = ~n4888 & ~n4889 ;
  assign n4891 = \P1_state_reg[0]/NET0131  & ~n4890 ;
  assign n4892 = ~\P1_state_reg[0]/NET0131  & \P2_reg3_reg[27]/NET0131  ;
  assign n4893 = n2987 & n3976 ;
  assign n4894 = ~n4892 & ~n4893 ;
  assign n4895 = ~n4891 & n4894 ;
  assign n4898 = n974 & n3448 ;
  assign n4899 = n974 & ~n3980 ;
  assign n4900 = n3980 & ~n4429 ;
  assign n4901 = ~n4899 & ~n4900 ;
  assign n4902 = ~n3677 & ~n4901 ;
  assign n4912 = n3980 & n4486 ;
  assign n4909 = n3712 & ~n3980 ;
  assign n4910 = n4064 & ~n4909 ;
  assign n4911 = n974 & ~n4910 ;
  assign n4913 = n969 & ~n4067 ;
  assign n4914 = ~n4911 & ~n4913 ;
  assign n4915 = ~n4912 & n4914 ;
  assign n4916 = ~n4902 & n4915 ;
  assign n4903 = n3980 & n4480 ;
  assign n4904 = ~n4899 & ~n4903 ;
  assign n4905 = n1936 & ~n4904 ;
  assign n4906 = n3980 & ~n4466 ;
  assign n4907 = ~n4899 & ~n4906 ;
  assign n4908 = ~n3563 & ~n4907 ;
  assign n4917 = ~n4905 & ~n4908 ;
  assign n4918 = n4916 & n4917 ;
  assign n4919 = n3450 & ~n4918 ;
  assign n4920 = ~n4898 & ~n4919 ;
  assign n4921 = \P1_state_reg[0]/NET0131  & ~n4920 ;
  assign n4896 = \P1_reg3_reg[27]/NET0131  & ~\P1_state_reg[0]/NET0131  ;
  assign n4897 = n974 & n1953 ;
  assign n4922 = ~n4896 & ~n4897 ;
  assign n4923 = ~n4921 & n4922 ;
  assign n4924 = \P2_reg2_reg[25]/NET0131  & ~n1983 ;
  assign n4925 = \P2_reg2_reg[25]/NET0131  & n2024 ;
  assign n4935 = \P2_reg2_reg[25]/NET0131  & ~n3758 ;
  assign n4939 = n3758 & ~n4609 ;
  assign n4940 = ~n4935 & ~n4939 ;
  assign n4941 = ~n3320 & ~n4940 ;
  assign n4936 = n3758 & ~n4595 ;
  assign n4937 = ~n4935 & ~n4936 ;
  assign n4938 = ~n3177 & ~n4937 ;
  assign n4926 = n3355 & n4617 ;
  assign n4927 = n3034 & n3358 ;
  assign n4928 = ~n4629 & ~n4927 ;
  assign n4929 = ~n4926 & n4928 ;
  assign n4930 = n3758 & ~n4929 ;
  assign n4931 = n3039 & n3420 ;
  assign n4932 = n3745 & ~n3758 ;
  assign n4933 = n3774 & ~n4932 ;
  assign n4934 = \P2_reg2_reg[25]/NET0131  & ~n4933 ;
  assign n4942 = ~n4931 & ~n4934 ;
  assign n4943 = ~n4930 & n4942 ;
  assign n4944 = ~n4938 & n4943 ;
  assign n4945 = ~n4941 & n4944 ;
  assign n4946 = n2026 & ~n4945 ;
  assign n4947 = ~n4925 & ~n4946 ;
  assign n4948 = \P1_state_reg[0]/NET0131  & ~n4947 ;
  assign n4949 = ~n4924 & ~n4948 ;
  assign n4950 = \P2_reg2_reg[26]/NET0131  & n2024 ;
  assign n4951 = \P2_reg2_reg[26]/NET0131  & ~n3758 ;
  assign n4952 = n3758 & ~n4732 ;
  assign n4953 = ~n4951 & ~n4952 ;
  assign n4954 = ~n3320 & ~n4953 ;
  assign n4955 = n3758 & ~n4764 ;
  assign n4956 = ~n4951 & ~n4955 ;
  assign n4957 = ~n3177 & ~n4956 ;
  assign n4958 = n3411 & n4773 ;
  assign n4959 = n3012 & n3358 ;
  assign n4960 = n3355 & n4779 ;
  assign n4961 = ~n4959 & ~n4960 ;
  assign n4962 = ~n4958 & n4961 ;
  assign n4963 = n3758 & ~n4962 ;
  assign n4964 = n3017 & n3420 ;
  assign n4965 = \P2_reg2_reg[26]/NET0131  & ~n4384 ;
  assign n4966 = ~n4964 & ~n4965 ;
  assign n4967 = ~n4963 & n4966 ;
  assign n4968 = ~n4957 & n4967 ;
  assign n4969 = ~n4954 & n4968 ;
  assign n4970 = n2026 & ~n4969 ;
  assign n4971 = ~n4950 & ~n4970 ;
  assign n4972 = \P1_state_reg[0]/NET0131  & ~n4971 ;
  assign n4973 = \P2_reg2_reg[26]/NET0131  & ~n1983 ;
  assign n4974 = ~n4972 & ~n4973 ;
  assign n4975 = \P2_reg0_reg[24]/NET0131  & ~n1983 ;
  assign n4976 = \P2_reg0_reg[24]/NET0131  & n2024 ;
  assign n4977 = \P2_reg0_reg[24]/NET0131  & ~n2040 ;
  assign n4978 = n3813 & ~n4170 ;
  assign n4979 = n3795 & ~n4978 ;
  assign n4980 = n3852 & ~n4979 ;
  assign n4981 = n4200 & ~n4980 ;
  assign n4982 = ~n4200 & n4980 ;
  assign n4983 = ~n4981 & ~n4982 ;
  assign n4984 = n2040 & ~n4983 ;
  assign n4985 = ~n4977 & ~n4984 ;
  assign n4986 = ~n3320 & ~n4985 ;
  assign n4990 = n3892 & n3900 ;
  assign n4987 = ~n3875 & n3896 ;
  assign n4988 = n3907 & ~n4987 ;
  assign n4989 = n3899 & ~n4988 ;
  assign n4991 = n3914 & ~n4989 ;
  assign n4992 = ~n4990 & n4991 ;
  assign n4993 = n3922 & ~n4992 ;
  assign n4994 = n3930 & ~n4993 ;
  assign n4995 = n4200 & n4994 ;
  assign n4996 = ~n4200 & ~n4994 ;
  assign n4997 = ~n4995 & ~n4996 ;
  assign n4998 = n2040 & ~n4997 ;
  assign n4999 = ~n4977 & ~n4998 ;
  assign n5000 = ~n3177 & ~n4999 ;
  assign n5004 = n3043 & ~n4622 ;
  assign n5005 = ~n4623 & ~n5004 ;
  assign n5006 = ~n2058 & ~n5005 ;
  assign n5007 = n2058 & n3088 ;
  assign n5008 = ~n5006 & ~n5007 ;
  assign n5009 = n3411 & n5008 ;
  assign n5001 = n3054 & ~n4614 ;
  assign n5002 = ~n4615 & ~n5001 ;
  assign n5003 = n3355 & n5002 ;
  assign n5010 = n3054 & n3358 ;
  assign n5011 = ~n5003 & ~n5010 ;
  assign n5012 = ~n5009 & n5011 ;
  assign n5013 = n2040 & ~n5012 ;
  assign n5014 = \P2_reg0_reg[24]/NET0131  & ~n3426 ;
  assign n5015 = ~n5013 & ~n5014 ;
  assign n5016 = ~n5000 & n5015 ;
  assign n5017 = ~n4986 & n5016 ;
  assign n5018 = n2026 & ~n5017 ;
  assign n5019 = ~n4976 & ~n5018 ;
  assign n5020 = \P1_state_reg[0]/NET0131  & ~n5019 ;
  assign n5021 = ~n4975 & ~n5020 ;
  assign n5022 = \P2_reg0_reg[27]/NET0131  & n2024 ;
  assign n5023 = \P2_reg0_reg[27]/NET0131  & ~n2040 ;
  assign n5024 = n2040 & n4828 ;
  assign n5025 = ~n5023 & ~n5024 ;
  assign n5026 = ~n3177 & ~n5025 ;
  assign n5030 = n2040 & ~n4864 ;
  assign n5031 = ~n5023 & ~n5030 ;
  assign n5032 = ~n3320 & ~n5031 ;
  assign n5027 = n2040 & n4869 ;
  assign n5028 = ~n5023 & ~n5027 ;
  assign n5029 = n3355 & ~n5028 ;
  assign n5033 = n2040 & n4877 ;
  assign n5034 = ~n5023 & ~n5033 ;
  assign n5035 = n3411 & ~n5034 ;
  assign n5036 = n2982 & n3358 ;
  assign n5037 = n2040 & n5036 ;
  assign n5038 = \P2_reg0_reg[27]/NET0131  & ~n3423 ;
  assign n5039 = ~n5037 & ~n5038 ;
  assign n5040 = ~n5035 & n5039 ;
  assign n5041 = ~n5029 & n5040 ;
  assign n5042 = ~n5032 & n5041 ;
  assign n5043 = ~n5026 & n5042 ;
  assign n5044 = n2026 & ~n5043 ;
  assign n5045 = ~n5022 & ~n5044 ;
  assign n5046 = \P1_state_reg[0]/NET0131  & ~n5045 ;
  assign n5047 = \P2_reg0_reg[27]/NET0131  & ~n1983 ;
  assign n5048 = ~n5046 & ~n5047 ;
  assign n5049 = \P1_reg2_reg[27]/NET0131  & ~n3435 ;
  assign n5050 = \P1_reg2_reg[27]/NET0131  & n3448 ;
  assign n5051 = \P1_reg2_reg[27]/NET0131  & ~n3466 ;
  assign n5052 = n3466 & ~n4429 ;
  assign n5053 = ~n5051 & ~n5052 ;
  assign n5054 = ~n3677 & ~n5053 ;
  assign n5062 = n3466 & n4485 ;
  assign n5063 = ~n5051 & ~n5062 ;
  assign n5064 = n3712 & ~n5063 ;
  assign n5065 = n969 & n3466 ;
  assign n5066 = ~n5051 & ~n5065 ;
  assign n5067 = n1880 & ~n5066 ;
  assign n5061 = n974 & n1763 ;
  assign n5068 = \P1_reg2_reg[27]/NET0131  & n3716 ;
  assign n5069 = ~n5061 & ~n5068 ;
  assign n5070 = ~n5067 & n5069 ;
  assign n5071 = ~n5064 & n5070 ;
  assign n5072 = ~n5054 & n5071 ;
  assign n5055 = n3466 & n4480 ;
  assign n5056 = ~n5051 & ~n5055 ;
  assign n5057 = n1936 & ~n5056 ;
  assign n5058 = n3466 & ~n4466 ;
  assign n5059 = ~n5051 & ~n5058 ;
  assign n5060 = ~n3563 & ~n5059 ;
  assign n5073 = ~n5057 & ~n5060 ;
  assign n5074 = n5072 & n5073 ;
  assign n5075 = n3450 & ~n5074 ;
  assign n5076 = ~n5050 & ~n5075 ;
  assign n5077 = \P1_state_reg[0]/NET0131  & ~n5076 ;
  assign n5078 = ~n5049 & ~n5077 ;
  assign n5079 = \P2_reg1_reg[24]/NET0131  & ~n1983 ;
  assign n5080 = \P2_reg1_reg[24]/NET0131  & n2024 ;
  assign n5081 = \P2_reg1_reg[24]/NET0131  & ~n3733 ;
  assign n5082 = n3733 & ~n4983 ;
  assign n5083 = ~n5081 & ~n5082 ;
  assign n5084 = ~n3320 & ~n5083 ;
  assign n5085 = n3733 & ~n4997 ;
  assign n5086 = ~n5081 & ~n5085 ;
  assign n5087 = ~n3177 & ~n5086 ;
  assign n5088 = n3733 & ~n5012 ;
  assign n5089 = \P2_reg1_reg[24]/NET0131  & ~n3747 ;
  assign n5090 = ~n5088 & ~n5089 ;
  assign n5091 = ~n5087 & n5090 ;
  assign n5092 = ~n5084 & n5091 ;
  assign n5093 = n2026 & ~n5092 ;
  assign n5094 = ~n5080 & ~n5093 ;
  assign n5095 = \P1_state_reg[0]/NET0131  & ~n5094 ;
  assign n5096 = ~n5079 & ~n5095 ;
  assign n5097 = \P2_reg1_reg[25]/NET0131  & ~n1983 ;
  assign n5098 = \P2_reg1_reg[25]/NET0131  & n2024 ;
  assign n5101 = \P2_reg1_reg[25]/NET0131  & ~n3733 ;
  assign n5105 = n3733 & ~n4609 ;
  assign n5106 = ~n5101 & ~n5105 ;
  assign n5107 = ~n3320 & ~n5106 ;
  assign n5102 = n3733 & ~n4595 ;
  assign n5103 = ~n5101 & ~n5102 ;
  assign n5104 = ~n3177 & ~n5103 ;
  assign n5099 = \P2_reg1_reg[25]/NET0131  & ~n3747 ;
  assign n5100 = n3733 & ~n4929 ;
  assign n5108 = ~n5099 & ~n5100 ;
  assign n5109 = ~n5104 & n5108 ;
  assign n5110 = ~n5107 & n5109 ;
  assign n5111 = n2026 & ~n5110 ;
  assign n5112 = ~n5098 & ~n5111 ;
  assign n5113 = \P1_state_reg[0]/NET0131  & ~n5112 ;
  assign n5114 = ~n5097 & ~n5113 ;
  assign n5115 = \P2_reg1_reg[26]/NET0131  & ~n1983 ;
  assign n5116 = \P2_reg1_reg[26]/NET0131  & ~n3733 ;
  assign n5117 = n3733 & ~n4732 ;
  assign n5118 = ~n5116 & ~n5117 ;
  assign n5119 = ~n3320 & ~n5118 ;
  assign n5120 = n3733 & ~n4764 ;
  assign n5121 = ~n5116 & ~n5120 ;
  assign n5122 = ~n3177 & ~n5121 ;
  assign n5123 = n3733 & ~n4962 ;
  assign n5124 = \P2_reg1_reg[26]/NET0131  & ~n3747 ;
  assign n5125 = ~n5123 & ~n5124 ;
  assign n5126 = ~n5122 & n5125 ;
  assign n5127 = ~n5119 & n5126 ;
  assign n5128 = n2026 & ~n5127 ;
  assign n5129 = \P2_reg1_reg[26]/NET0131  & n2024 ;
  assign n5130 = ~n5128 & ~n5129 ;
  assign n5131 = \P1_state_reg[0]/NET0131  & ~n5130 ;
  assign n5132 = ~n5115 & ~n5131 ;
  assign n5133 = \P2_reg1_reg[27]/NET0131  & ~n3733 ;
  assign n5134 = n3733 & n4828 ;
  assign n5135 = ~n5133 & ~n5134 ;
  assign n5136 = ~n3177 & ~n5135 ;
  assign n5140 = n3733 & n4869 ;
  assign n5141 = ~n5133 & ~n5140 ;
  assign n5142 = n3355 & ~n5141 ;
  assign n5137 = n3733 & ~n4864 ;
  assign n5138 = ~n5133 & ~n5137 ;
  assign n5139 = ~n3320 & ~n5138 ;
  assign n5143 = n3733 & n4877 ;
  assign n5144 = ~n5133 & ~n5143 ;
  assign n5145 = n3411 & ~n5144 ;
  assign n5146 = n3733 & n5036 ;
  assign n5147 = \P2_reg1_reg[27]/NET0131  & ~n3743 ;
  assign n5148 = ~n5146 & ~n5147 ;
  assign n5149 = ~n5145 & n5148 ;
  assign n5150 = ~n5139 & n5149 ;
  assign n5151 = ~n5142 & n5150 ;
  assign n5152 = ~n5136 & n5151 ;
  assign n5153 = n2026 & ~n5152 ;
  assign n5154 = \P2_reg1_reg[27]/NET0131  & n2024 ;
  assign n5155 = ~n5153 & ~n5154 ;
  assign n5156 = \P1_state_reg[0]/NET0131  & ~n5155 ;
  assign n5157 = \P2_reg1_reg[27]/NET0131  & ~n1983 ;
  assign n5158 = ~n5156 & ~n5157 ;
  assign n5159 = \P1_reg2_reg[24]/NET0131  & ~n3435 ;
  assign n5160 = \P1_reg2_reg[24]/NET0131  & n3448 ;
  assign n5161 = \P1_reg2_reg[24]/NET0131  & ~n3466 ;
  assign n5162 = n4000 & n4014 ;
  assign n5163 = ~n4006 & n4010 ;
  assign n5164 = n4021 & ~n5163 ;
  assign n5165 = n4013 & ~n5164 ;
  assign n5166 = n4028 & ~n5165 ;
  assign n5167 = ~n5162 & n5166 ;
  assign n5168 = n4033 & ~n5167 ;
  assign n5169 = n4043 & ~n5168 ;
  assign n5170 = n1818 & n5169 ;
  assign n5171 = ~n1818 & ~n5169 ;
  assign n5172 = ~n5170 & ~n5171 ;
  assign n5173 = n3466 & ~n5172 ;
  assign n5174 = ~n5161 & ~n5173 ;
  assign n5175 = ~n3563 & ~n5174 ;
  assign n5188 = ~n1327 & n3700 ;
  assign n5189 = n1047 & ~n5188 ;
  assign n5190 = ~n4686 & ~n5189 ;
  assign n5191 = n3466 & n5190 ;
  assign n5192 = ~n5161 & ~n5191 ;
  assign n5193 = n3712 & ~n5192 ;
  assign n5206 = n1047 & n1880 ;
  assign n5207 = n3466 & n5206 ;
  assign n5204 = \P1_reg2_reg[24]/NET0131  & ~n3718 ;
  assign n5205 = n1058 & n1763 ;
  assign n5208 = ~n5204 & ~n5205 ;
  assign n5209 = ~n5207 & n5208 ;
  assign n5210 = ~n5193 & n5209 ;
  assign n5211 = ~n5175 & n5210 ;
  assign n5177 = n1478 & ~n1489 ;
  assign n5178 = n1720 & ~n5177 ;
  assign n5179 = n1377 & ~n5178 ;
  assign n5176 = n1479 & n1749 ;
  assign n5180 = n1710 & ~n5176 ;
  assign n5181 = ~n5179 & n5180 ;
  assign n5182 = n1818 & ~n5181 ;
  assign n5183 = ~n1818 & n5181 ;
  assign n5184 = ~n5182 & ~n5183 ;
  assign n5185 = n3466 & ~n5184 ;
  assign n5186 = ~n5161 & ~n5185 ;
  assign n5187 = ~n3677 & ~n5186 ;
  assign n5194 = n1038 & ~n4075 ;
  assign n5195 = n3568 & n4470 ;
  assign n5196 = n3592 & n5195 ;
  assign n5197 = ~n5194 & ~n5196 ;
  assign n5198 = ~n537 & ~n5197 ;
  assign n5199 = n537 & n1336 ;
  assign n5200 = ~n5198 & ~n5199 ;
  assign n5201 = n3466 & n5200 ;
  assign n5202 = ~n5161 & ~n5201 ;
  assign n5203 = n1936 & ~n5202 ;
  assign n5212 = ~n5187 & ~n5203 ;
  assign n5213 = n5211 & n5212 ;
  assign n5214 = n3450 & ~n5213 ;
  assign n5215 = ~n5160 & ~n5214 ;
  assign n5216 = \P1_state_reg[0]/NET0131  & ~n5215 ;
  assign n5217 = ~n5159 & ~n5216 ;
  assign n5218 = \P1_reg2_reg[28]/NET0131  & ~n3435 ;
  assign n5219 = \P1_reg2_reg[28]/NET0131  & n3448 ;
  assign n5220 = \P1_reg2_reg[28]/NET0131  & ~n3466 ;
  assign n5221 = n3466 & ~n4101 ;
  assign n5222 = ~n5220 & ~n5221 ;
  assign n5223 = ~n3677 & ~n5222 ;
  assign n5224 = n3466 & n4059 ;
  assign n5225 = ~n5220 & ~n5224 ;
  assign n5226 = n3712 & ~n5225 ;
  assign n5229 = n933 & n1880 ;
  assign n5230 = n3466 & n5229 ;
  assign n5227 = \P1_reg2_reg[28]/NET0131  & ~n3718 ;
  assign n5228 = n941 & n1763 ;
  assign n5237 = ~n5227 & ~n5228 ;
  assign n5238 = ~n5230 & n5237 ;
  assign n5239 = ~n5226 & n5238 ;
  assign n5240 = ~n5223 & n5239 ;
  assign n5231 = n3466 & ~n4084 ;
  assign n5232 = ~n5220 & ~n5231 ;
  assign n5233 = n1936 & ~n5232 ;
  assign n5234 = n3466 & ~n4053 ;
  assign n5235 = ~n5220 & ~n5234 ;
  assign n5236 = ~n3563 & ~n5235 ;
  assign n5241 = ~n5233 & ~n5236 ;
  assign n5242 = n5240 & n5241 ;
  assign n5243 = n3450 & ~n5242 ;
  assign n5244 = ~n5219 & ~n5243 ;
  assign n5245 = \P1_state_reg[0]/NET0131  & ~n5244 ;
  assign n5246 = ~n5218 & ~n5245 ;
  assign n5247 = \P2_reg2_reg[27]/NET0131  & ~n3758 ;
  assign n5248 = n3758 & n4828 ;
  assign n5249 = ~n5247 & ~n5248 ;
  assign n5250 = ~n3177 & ~n5249 ;
  assign n5254 = n3758 & ~n4864 ;
  assign n5255 = ~n5247 & ~n5254 ;
  assign n5256 = ~n3320 & ~n5255 ;
  assign n5251 = n3758 & n4869 ;
  assign n5252 = ~n5247 & ~n5251 ;
  assign n5253 = n3355 & ~n5252 ;
  assign n5257 = n3758 & n4877 ;
  assign n5258 = ~n5247 & ~n5257 ;
  assign n5259 = n3411 & ~n5258 ;
  assign n5260 = n3758 & n5036 ;
  assign n5261 = n2987 & n3420 ;
  assign n5262 = \P2_reg2_reg[27]/NET0131  & ~n3774 ;
  assign n5263 = ~n5261 & ~n5262 ;
  assign n5264 = ~n5260 & n5263 ;
  assign n5265 = ~n5259 & n5264 ;
  assign n5266 = ~n5253 & n5265 ;
  assign n5267 = ~n5256 & n5266 ;
  assign n5268 = ~n5250 & n5267 ;
  assign n5269 = n2026 & ~n5268 ;
  assign n5270 = \P2_reg2_reg[27]/NET0131  & n2024 ;
  assign n5271 = ~n5269 & ~n5270 ;
  assign n5272 = \P1_state_reg[0]/NET0131  & ~n5271 ;
  assign n5273 = \P2_reg2_reg[27]/NET0131  & ~n1983 ;
  assign n5274 = ~n5272 & ~n5273 ;
  assign n5275 = n3358 & n4141 ;
  assign n5276 = ~n3372 & n3411 ;
  assign n5277 = n3407 & n5276 ;
  assign n5278 = ~n5275 & ~n5277 ;
  assign n5279 = n3350 & ~n4159 ;
  assign n5280 = n4141 & ~n5279 ;
  assign n5281 = ~n4141 & n5279 ;
  assign n5282 = ~n5280 & ~n5281 ;
  assign n5283 = n3354 & n5282 ;
  assign n5284 = n5278 & ~n5283 ;
  assign n5285 = n3758 & ~n5284 ;
  assign n5286 = ~n3776 & ~n5285 ;
  assign n5287 = n1983 & ~n2023 ;
  assign n5288 = ~n5286 & n5287 ;
  assign n5289 = ~n3357 & ~n3758 ;
  assign n5290 = n3774 & ~n5289 ;
  assign n5291 = ~n4381 & n5287 ;
  assign n5292 = n5290 & n5291 ;
  assign n5293 = \P2_reg2_reg[31]/NET0131  & ~n5292 ;
  assign n5294 = ~n5288 & ~n5293 ;
  assign n5295 = \P1_reg0_reg[25]/NET0131  & ~n3435 ;
  assign n5296 = \P1_reg0_reg[25]/NET0131  & n3448 ;
  assign n5297 = \P1_reg0_reg[25]/NET0131  & ~n4396 ;
  assign n5310 = n4396 & n4689 ;
  assign n5311 = ~n5297 & ~n5310 ;
  assign n5312 = n3712 & ~n5311 ;
  assign n5307 = n4396 & n4682 ;
  assign n5308 = ~n5297 & ~n5307 ;
  assign n5309 = n1936 & ~n5308 ;
  assign n5304 = n1029 & n1880 ;
  assign n5305 = n4396 & n5304 ;
  assign n5306 = \P1_reg0_reg[25]/NET0131  & ~n4493 ;
  assign n5313 = ~n5305 & ~n5306 ;
  assign n5314 = ~n5309 & n5313 ;
  assign n5315 = ~n5312 & n5314 ;
  assign n5298 = n4396 & ~n4658 ;
  assign n5299 = ~n5297 & ~n5298 ;
  assign n5300 = ~n3677 & ~n5299 ;
  assign n5301 = n4396 & ~n4672 ;
  assign n5302 = ~n5297 & ~n5301 ;
  assign n5303 = ~n3563 & ~n5302 ;
  assign n5316 = ~n5300 & ~n5303 ;
  assign n5317 = n5315 & n5316 ;
  assign n5318 = n3450 & ~n5317 ;
  assign n5319 = ~n5296 & ~n5318 ;
  assign n5320 = \P1_state_reg[0]/NET0131  & ~n5319 ;
  assign n5321 = ~n5295 & ~n5320 ;
  assign n5322 = \P1_reg0_reg[28]/NET0131  & n3448 ;
  assign n5323 = \P1_reg0_reg[28]/NET0131  & ~n4396 ;
  assign n5324 = ~n4101 & n4396 ;
  assign n5325 = ~n5323 & ~n5324 ;
  assign n5326 = ~n3677 & ~n5325 ;
  assign n5327 = n4059 & n4396 ;
  assign n5328 = ~n5323 & ~n5327 ;
  assign n5329 = n3712 & ~n5328 ;
  assign n5330 = \P1_reg0_reg[28]/NET0131  & ~n4493 ;
  assign n5331 = n4396 & n5229 ;
  assign n5338 = ~n5330 & ~n5331 ;
  assign n5339 = ~n5329 & n5338 ;
  assign n5340 = ~n5326 & n5339 ;
  assign n5332 = ~n4084 & n4396 ;
  assign n5333 = ~n5323 & ~n5332 ;
  assign n5334 = n1936 & ~n5333 ;
  assign n5335 = ~n4053 & n4396 ;
  assign n5336 = ~n5323 & ~n5335 ;
  assign n5337 = ~n3563 & ~n5336 ;
  assign n5341 = ~n5334 & ~n5337 ;
  assign n5342 = n5340 & n5341 ;
  assign n5343 = n3450 & ~n5342 ;
  assign n5344 = ~n5322 & ~n5343 ;
  assign n5345 = \P1_state_reg[0]/NET0131  & ~n5344 ;
  assign n5346 = \P1_reg0_reg[28]/NET0131  & ~n3435 ;
  assign n5347 = ~n5345 & ~n5346 ;
  assign n5348 = \P1_reg1_reg[24]/NET0131  & ~n3435 ;
  assign n5349 = \P1_reg1_reg[24]/NET0131  & n3448 ;
  assign n5350 = \P1_reg1_reg[24]/NET0131  & ~n4532 ;
  assign n5351 = n4532 & ~n5172 ;
  assign n5352 = ~n5350 & ~n5351 ;
  assign n5353 = ~n3563 & ~n5352 ;
  assign n5359 = n4532 & n5190 ;
  assign n5360 = ~n5350 & ~n5359 ;
  assign n5361 = n3712 & ~n5360 ;
  assign n5357 = \P1_reg1_reg[24]/NET0131  & ~n4541 ;
  assign n5358 = n4532 & n5206 ;
  assign n5365 = ~n5357 & ~n5358 ;
  assign n5366 = ~n5361 & n5365 ;
  assign n5367 = ~n5353 & n5366 ;
  assign n5354 = n4532 & n5200 ;
  assign n5355 = ~n5350 & ~n5354 ;
  assign n5356 = n1936 & ~n5355 ;
  assign n5362 = n4532 & ~n5184 ;
  assign n5363 = ~n5350 & ~n5362 ;
  assign n5364 = ~n3677 & ~n5363 ;
  assign n5368 = ~n5356 & ~n5364 ;
  assign n5369 = n5367 & n5368 ;
  assign n5370 = n3450 & ~n5369 ;
  assign n5371 = ~n5349 & ~n5370 ;
  assign n5372 = \P1_state_reg[0]/NET0131  & ~n5371 ;
  assign n5373 = ~n5348 & ~n5372 ;
  assign n5374 = \P1_reg1_reg[25]/NET0131  & ~n3435 ;
  assign n5375 = \P1_reg1_reg[25]/NET0131  & n3448 ;
  assign n5376 = \P1_reg1_reg[25]/NET0131  & ~n4532 ;
  assign n5388 = n4532 & n4689 ;
  assign n5389 = ~n5376 & ~n5388 ;
  assign n5390 = n3712 & ~n5389 ;
  assign n5385 = n4532 & n4682 ;
  assign n5386 = ~n5376 & ~n5385 ;
  assign n5387 = n1936 & ~n5386 ;
  assign n5383 = n4532 & n5304 ;
  assign n5384 = \P1_reg1_reg[25]/NET0131  & ~n4541 ;
  assign n5391 = ~n5383 & ~n5384 ;
  assign n5392 = ~n5387 & n5391 ;
  assign n5393 = ~n5390 & n5392 ;
  assign n5377 = n4532 & ~n4658 ;
  assign n5378 = ~n5376 & ~n5377 ;
  assign n5379 = ~n3677 & ~n5378 ;
  assign n5380 = n4532 & ~n4672 ;
  assign n5381 = ~n5376 & ~n5380 ;
  assign n5382 = ~n3563 & ~n5381 ;
  assign n5394 = ~n5379 & ~n5382 ;
  assign n5395 = n5393 & n5394 ;
  assign n5396 = n3450 & ~n5395 ;
  assign n5397 = ~n5375 & ~n5396 ;
  assign n5398 = \P1_state_reg[0]/NET0131  & ~n5397 ;
  assign n5399 = ~n5374 & ~n5398 ;
  assign n5400 = \P1_reg1_reg[28]/NET0131  & n3448 ;
  assign n5401 = \P1_reg1_reg[28]/NET0131  & ~n4532 ;
  assign n5402 = ~n4101 & n4532 ;
  assign n5403 = ~n5401 & ~n5402 ;
  assign n5404 = ~n3677 & ~n5403 ;
  assign n5405 = n4059 & n4532 ;
  assign n5406 = ~n5401 & ~n5405 ;
  assign n5407 = n3712 & ~n5406 ;
  assign n5408 = \P1_reg1_reg[28]/NET0131  & ~n4541 ;
  assign n5409 = n4532 & n5229 ;
  assign n5416 = ~n5408 & ~n5409 ;
  assign n5417 = ~n5407 & n5416 ;
  assign n5418 = ~n5404 & n5417 ;
  assign n5410 = ~n4084 & n4532 ;
  assign n5411 = ~n5401 & ~n5410 ;
  assign n5412 = n1936 & ~n5411 ;
  assign n5413 = ~n4053 & n4532 ;
  assign n5414 = ~n5401 & ~n5413 ;
  assign n5415 = ~n3563 & ~n5414 ;
  assign n5419 = ~n5412 & ~n5415 ;
  assign n5420 = n5418 & n5419 ;
  assign n5421 = n3450 & ~n5420 ;
  assign n5422 = ~n5400 & ~n5421 ;
  assign n5423 = \P1_state_reg[0]/NET0131  & ~n5422 ;
  assign n5424 = \P1_reg1_reg[28]/NET0131  & ~n3435 ;
  assign n5425 = ~n5423 & ~n5424 ;
  assign n5428 = n1447 & n3448 ;
  assign n5431 = n1447 & ~n3980 ;
  assign n5457 = n1403 & ~n3585 ;
  assign n5458 = ~n1403 & n3585 ;
  assign n5459 = ~n5457 & ~n5458 ;
  assign n5460 = ~n537 & ~n5459 ;
  assign n5461 = n537 & n1475 ;
  assign n5462 = ~n5460 & ~n5461 ;
  assign n5463 = n3980 & n5462 ;
  assign n5464 = ~n5431 & ~n5463 ;
  assign n5465 = n1936 & ~n5464 ;
  assign n5440 = ~n1136 & n3690 ;
  assign n5441 = n3691 & n5440 ;
  assign n5442 = ~n1466 & n5441 ;
  assign n5443 = n1443 & ~n5442 ;
  assign n5444 = ~n1443 & n5442 ;
  assign n5445 = ~n5443 & ~n5444 ;
  assign n5446 = n3980 & n5445 ;
  assign n5447 = ~n5431 & ~n5446 ;
  assign n5448 = n3712 & ~n5447 ;
  assign n5429 = n1447 & ~n4064 ;
  assign n5430 = n1443 & ~n4067 ;
  assign n5466 = ~n5429 & ~n5430 ;
  assign n5467 = ~n5448 & n5466 ;
  assign n5468 = ~n5465 & n5467 ;
  assign n5432 = n3625 & ~n3650 ;
  assign n5433 = n3656 & ~n5432 ;
  assign n5434 = n1825 & ~n5433 ;
  assign n5435 = ~n1825 & n5433 ;
  assign n5436 = ~n5434 & ~n5435 ;
  assign n5437 = n3980 & n5436 ;
  assign n5438 = ~n5431 & ~n5437 ;
  assign n5439 = ~n3677 & ~n5438 ;
  assign n5449 = n3490 & ~n3533 ;
  assign n5450 = n3540 & ~n5449 ;
  assign n5451 = n1825 & ~n5450 ;
  assign n5452 = ~n1825 & n5450 ;
  assign n5453 = ~n5451 & ~n5452 ;
  assign n5454 = n3980 & ~n5453 ;
  assign n5455 = ~n5431 & ~n5454 ;
  assign n5456 = ~n3563 & ~n5455 ;
  assign n5469 = ~n5439 & ~n5456 ;
  assign n5470 = n5468 & n5469 ;
  assign n5471 = n3450 & ~n5470 ;
  assign n5472 = ~n5428 & ~n5471 ;
  assign n5473 = \P1_state_reg[0]/NET0131  & ~n5472 ;
  assign n5426 = \P1_reg3_reg[17]/NET0131  & ~\P1_state_reg[0]/NET0131  ;
  assign n5427 = n1447 & n1953 ;
  assign n5474 = ~n5426 & ~n5427 ;
  assign n5475 = ~n5473 & n5474 ;
  assign n5478 = n1399 & n3448 ;
  assign n5480 = n1399 & ~n3980 ;
  assign n5481 = n1394 & ~n5444 ;
  assign n5482 = ~n3696 & ~n5481 ;
  assign n5483 = n3980 & n5482 ;
  assign n5484 = ~n5480 & ~n5483 ;
  assign n5485 = n3712 & ~n5484 ;
  assign n5479 = n1399 & ~n4064 ;
  assign n5540 = n1394 & ~n4067 ;
  assign n5541 = ~n5479 & ~n5540 ;
  assign n5542 = ~n5485 & n5541 ;
  assign n5531 = ~n1427 & ~n5458 ;
  assign n5532 = n1427 & n5458 ;
  assign n5533 = ~n5531 & ~n5532 ;
  assign n5534 = ~n537 & ~n5533 ;
  assign n5535 = n537 & ~n1452 ;
  assign n5536 = ~n5534 & ~n5535 ;
  assign n5537 = n3980 & ~n5536 ;
  assign n5538 = ~n5480 & ~n5537 ;
  assign n5539 = n1936 & ~n5538 ;
  assign n5486 = n1120 & n1477 ;
  assign n5487 = n1283 & n1539 ;
  assign n5488 = ~n1686 & n5487 ;
  assign n5489 = n1283 & ~n1691 ;
  assign n5490 = ~n1483 & ~n5489 ;
  assign n5491 = ~n5488 & n5490 ;
  assign n5492 = n1235 & n1291 ;
  assign n5493 = ~n5491 & n5492 ;
  assign n5494 = n5486 & n5493 ;
  assign n5495 = n1291 & n1486 ;
  assign n5496 = ~n1177 & ~n5495 ;
  assign n5497 = n5486 & ~n5496 ;
  assign n5498 = n1182 & n1477 ;
  assign n5499 = ~n1714 & ~n5498 ;
  assign n5500 = ~n5497 & n5499 ;
  assign n5501 = ~n5494 & n5500 ;
  assign n5502 = n1824 & ~n5501 ;
  assign n5503 = ~n1824 & n5501 ;
  assign n5504 = ~n5502 & ~n5503 ;
  assign n5505 = n3980 & ~n5504 ;
  assign n5506 = ~n5480 & ~n5505 ;
  assign n5507 = ~n3677 & ~n5506 ;
  assign n5508 = n4009 & n4011 ;
  assign n5509 = ~n3988 & n3991 ;
  assign n5510 = n3982 & n3997 ;
  assign n5511 = ~n5509 & n5510 ;
  assign n5512 = ~n3994 & n3997 ;
  assign n5513 = n4002 & ~n5512 ;
  assign n5514 = ~n5511 & n5513 ;
  assign n5515 = n3998 & n4008 ;
  assign n5516 = ~n5514 & n5515 ;
  assign n5517 = n5508 & n5516 ;
  assign n5518 = n4005 & n4008 ;
  assign n5519 = n4017 & ~n5518 ;
  assign n5520 = n5508 & ~n5519 ;
  assign n5521 = n4011 & ~n4020 ;
  assign n5522 = ~n4024 & ~n5521 ;
  assign n5523 = ~n5520 & n5522 ;
  assign n5524 = ~n5517 & n5523 ;
  assign n5525 = n1824 & ~n5524 ;
  assign n5526 = ~n1824 & n5524 ;
  assign n5527 = ~n5525 & ~n5526 ;
  assign n5528 = n3980 & n5527 ;
  assign n5529 = ~n5480 & ~n5528 ;
  assign n5530 = ~n3563 & ~n5529 ;
  assign n5543 = ~n5507 & ~n5530 ;
  assign n5544 = ~n5539 & n5543 ;
  assign n5545 = n5542 & n5544 ;
  assign n5546 = n3450 & ~n5545 ;
  assign n5547 = ~n5478 & ~n5546 ;
  assign n5548 = \P1_state_reg[0]/NET0131  & ~n5547 ;
  assign n5476 = n1399 & n1953 ;
  assign n5477 = \P1_reg3_reg[18]/NET0131  & ~\P1_state_reg[0]/NET0131  ;
  assign n5549 = ~n5476 & ~n5477 ;
  assign n5550 = ~n5548 & n5549 ;
  assign n5553 = n2024 & n2373 ;
  assign n5555 = n2373 & ~n3788 ;
  assign n5556 = n4191 & ~n4587 ;
  assign n5557 = ~n4191 & n4587 ;
  assign n5558 = ~n5556 & ~n5557 ;
  assign n5559 = n3788 & n5558 ;
  assign n5560 = ~n5555 & ~n5559 ;
  assign n5561 = ~n3177 & ~n5560 ;
  assign n5582 = n3223 & ~n3280 ;
  assign n5583 = n3291 & ~n5582 ;
  assign n5584 = n4191 & n5583 ;
  assign n5585 = ~n4191 & ~n5583 ;
  assign n5586 = ~n5584 & ~n5585 ;
  assign n5587 = n3788 & n5586 ;
  assign n5588 = ~n5555 & ~n5587 ;
  assign n5589 = ~n3320 & ~n5588 ;
  assign n5554 = n2399 & ~n3965 ;
  assign n5590 = n2373 & ~n3962 ;
  assign n5591 = ~n5554 & ~n5590 ;
  assign n5592 = ~n5589 & n5591 ;
  assign n5593 = ~n5561 & n5592 ;
  assign n5562 = n2058 & ~n2804 ;
  assign n5564 = ~n2828 & n3387 ;
  assign n5565 = ~n2804 & n5564 ;
  assign n5566 = ~n2379 & n5565 ;
  assign n5567 = n2442 & ~n5566 ;
  assign n5563 = n3387 & n3390 ;
  assign n5568 = ~n2058 & ~n5563 ;
  assign n5569 = ~n5567 & n5568 ;
  assign n5570 = ~n5562 & ~n5569 ;
  assign n5571 = n3788 & ~n5570 ;
  assign n5572 = ~n5555 & ~n5571 ;
  assign n5573 = n3411 & ~n5572 ;
  assign n5574 = ~n2843 & n3339 ;
  assign n5575 = ~n2818 & n5574 ;
  assign n5576 = n2399 & ~n5575 ;
  assign n5577 = ~n2399 & n5575 ;
  assign n5578 = ~n5576 & ~n5577 ;
  assign n5579 = n3788 & n5578 ;
  assign n5580 = ~n5555 & ~n5579 ;
  assign n5581 = n3355 & ~n5580 ;
  assign n5594 = ~n5573 & ~n5581 ;
  assign n5595 = n5593 & n5594 ;
  assign n5596 = n2026 & ~n5595 ;
  assign n5597 = ~n5553 & ~n5596 ;
  assign n5598 = \P1_state_reg[0]/NET0131  & ~n5597 ;
  assign n5551 = ~\P1_state_reg[0]/NET0131  & \P2_reg3_reg[17]/NET0131  ;
  assign n5552 = n2373 & n3976 ;
  assign n5599 = ~n5551 & ~n5552 ;
  assign n5600 = ~n5598 & n5599 ;
  assign n5603 = n2024 & n2307 ;
  assign n5605 = n2307 & ~n3788 ;
  assign n5606 = n4197 & ~n4814 ;
  assign n5607 = ~n4197 & n4814 ;
  assign n5608 = ~n5606 & ~n5607 ;
  assign n5609 = n3788 & n5608 ;
  assign n5610 = ~n5605 & ~n5609 ;
  assign n5611 = ~n3177 & ~n5610 ;
  assign n5618 = ~n2311 & n5563 ;
  assign n5619 = n2368 & ~n5618 ;
  assign n5620 = ~n2368 & n5618 ;
  assign n5621 = ~n5619 & ~n5620 ;
  assign n5622 = ~n2058 & ~n5621 ;
  assign n5623 = n2058 & n2442 ;
  assign n5624 = ~n5622 & ~n5623 ;
  assign n5625 = n3788 & n5624 ;
  assign n5626 = ~n5605 & ~n5625 ;
  assign n5627 = n3411 & ~n5626 ;
  assign n5628 = n2299 & ~n3343 ;
  assign n5629 = ~n2299 & n3343 ;
  assign n5630 = ~n5628 & ~n5629 ;
  assign n5631 = n3788 & n5630 ;
  assign n5632 = ~n5605 & ~n5631 ;
  assign n5633 = n3355 & ~n5632 ;
  assign n5612 = n4197 & ~n4850 ;
  assign n5613 = ~n4197 & n4850 ;
  assign n5614 = ~n5612 & ~n5613 ;
  assign n5615 = n3788 & ~n5614 ;
  assign n5616 = ~n5605 & ~n5615 ;
  assign n5617 = ~n3320 & ~n5616 ;
  assign n5604 = n2307 & ~n3962 ;
  assign n5634 = n2299 & ~n3965 ;
  assign n5635 = ~n5604 & ~n5634 ;
  assign n5636 = ~n5617 & n5635 ;
  assign n5637 = ~n5633 & n5636 ;
  assign n5638 = ~n5627 & n5637 ;
  assign n5639 = ~n5611 & n5638 ;
  assign n5640 = n2026 & ~n5639 ;
  assign n5641 = ~n5603 & ~n5640 ;
  assign n5642 = \P1_state_reg[0]/NET0131  & ~n5641 ;
  assign n5601 = n2307 & n3976 ;
  assign n5602 = ~\P1_state_reg[0]/NET0131  & \P2_reg3_reg[19]/NET0131  ;
  assign n5643 = ~n5601 & ~n5602 ;
  assign n5644 = ~n5642 & n5643 ;
  assign n5645 = n1423 & n3448 ;
  assign n5646 = n1423 & ~n3980 ;
  assign n5647 = n537 & ~n1403 ;
  assign n5648 = ~n1403 & n5195 ;
  assign n5650 = ~n1427 & n5648 ;
  assign n5651 = n1374 & ~n5650 ;
  assign n5649 = n3587 & n5648 ;
  assign n5652 = ~n537 & ~n5649 ;
  assign n5653 = ~n5651 & n5652 ;
  assign n5654 = ~n5647 & ~n5653 ;
  assign n5655 = n3980 & ~n5654 ;
  assign n5656 = ~n5646 & ~n5655 ;
  assign n5657 = n1936 & ~n5656 ;
  assign n5665 = n1835 & ~n4415 ;
  assign n5666 = ~n1835 & n4415 ;
  assign n5667 = ~n5665 & ~n5666 ;
  assign n5668 = n3980 & ~n5667 ;
  assign n5669 = ~n5646 & ~n5668 ;
  assign n5670 = ~n3677 & ~n5669 ;
  assign n5659 = n1835 & ~n4458 ;
  assign n5660 = ~n1835 & n4458 ;
  assign n5661 = ~n5659 & ~n5660 ;
  assign n5662 = n3980 & n5661 ;
  assign n5663 = ~n5646 & ~n5662 ;
  assign n5664 = ~n3563 & ~n5663 ;
  assign n5671 = ~n1418 & n3696 ;
  assign n5672 = n1418 & ~n3696 ;
  assign n5673 = ~n5671 & ~n5672 ;
  assign n5674 = n3712 & n5673 ;
  assign n5675 = n3980 & n5674 ;
  assign n5658 = n1423 & ~n4910 ;
  assign n5676 = n1418 & ~n4067 ;
  assign n5677 = ~n5658 & ~n5676 ;
  assign n5678 = ~n5675 & n5677 ;
  assign n5679 = ~n5664 & n5678 ;
  assign n5680 = ~n5670 & n5679 ;
  assign n5681 = ~n5657 & n5680 ;
  assign n5682 = n3450 & ~n5681 ;
  assign n5683 = ~n5645 & ~n5682 ;
  assign n5684 = \P1_state_reg[0]/NET0131  & ~n5683 ;
  assign n5685 = \P1_reg3_reg[19]/NET0131  & ~\P1_state_reg[0]/NET0131  ;
  assign n5686 = n1423 & n1953 ;
  assign n5687 = ~n5685 & ~n5686 ;
  assign n5688 = ~n5684 & n5687 ;
  assign n5689 = n2024 & n3058 ;
  assign n5690 = n3058 & ~n3788 ;
  assign n5691 = n3788 & ~n4983 ;
  assign n5692 = ~n5690 & ~n5691 ;
  assign n5693 = ~n3320 & ~n5692 ;
  assign n5694 = n3788 & ~n4997 ;
  assign n5695 = ~n5690 & ~n5694 ;
  assign n5696 = ~n3177 & ~n5695 ;
  assign n5700 = n3788 & n5008 ;
  assign n5701 = ~n5690 & ~n5700 ;
  assign n5702 = n3411 & ~n5701 ;
  assign n5703 = n3788 & n5003 ;
  assign n5697 = n3355 & ~n3788 ;
  assign n5698 = n3962 & ~n5697 ;
  assign n5699 = n3058 & ~n5698 ;
  assign n5704 = n3054 & ~n3965 ;
  assign n5705 = ~n5699 & ~n5704 ;
  assign n5706 = ~n5703 & n5705 ;
  assign n5707 = ~n5702 & n5706 ;
  assign n5708 = ~n5696 & n5707 ;
  assign n5709 = ~n5693 & n5708 ;
  assign n5710 = n2026 & ~n5709 ;
  assign n5711 = ~n5689 & ~n5710 ;
  assign n5712 = \P1_state_reg[0]/NET0131  & ~n5711 ;
  assign n5713 = ~\P1_state_reg[0]/NET0131  & \P2_reg3_reg[24]/NET0131  ;
  assign n5714 = n3058 & n3976 ;
  assign n5715 = ~n5713 & ~n5714 ;
  assign n5716 = ~n5712 & n5715 ;
  assign n5719 = n1058 & n3448 ;
  assign n5720 = n1058 & ~n3980 ;
  assign n5721 = n3980 & ~n5172 ;
  assign n5722 = ~n5720 & ~n5721 ;
  assign n5723 = ~n3563 & ~n5722 ;
  assign n5729 = n3980 & n5190 ;
  assign n5730 = ~n5720 & ~n5729 ;
  assign n5731 = n3712 & ~n5730 ;
  assign n5727 = n1058 & ~n4064 ;
  assign n5728 = n1047 & ~n4067 ;
  assign n5735 = ~n5727 & ~n5728 ;
  assign n5736 = ~n5731 & n5735 ;
  assign n5737 = ~n5723 & n5736 ;
  assign n5724 = n3980 & ~n5184 ;
  assign n5725 = ~n5720 & ~n5724 ;
  assign n5726 = ~n3677 & ~n5725 ;
  assign n5732 = n3980 & n5200 ;
  assign n5733 = ~n5720 & ~n5732 ;
  assign n5734 = n1936 & ~n5733 ;
  assign n5738 = ~n5726 & ~n5734 ;
  assign n5739 = n5737 & n5738 ;
  assign n5740 = n3450 & ~n5739 ;
  assign n5741 = ~n5719 & ~n5740 ;
  assign n5742 = \P1_state_reg[0]/NET0131  & ~n5741 ;
  assign n5717 = \P1_reg3_reg[24]/NET0131  & ~\P1_state_reg[0]/NET0131  ;
  assign n5718 = n1058 & n1953 ;
  assign n5743 = ~n5717 & ~n5718 ;
  assign n5744 = ~n5742 & n5743 ;
  assign n5747 = n2024 & n3108 ;
  assign n5748 = n3108 & ~n3788 ;
  assign n5757 = ~n4721 & n4725 ;
  assign n5758 = n4209 & n5757 ;
  assign n5759 = ~n4209 & ~n5757 ;
  assign n5760 = ~n5758 & ~n5759 ;
  assign n5761 = n3788 & n5760 ;
  assign n5762 = ~n5748 & ~n5761 ;
  assign n5763 = ~n3320 & ~n5762 ;
  assign n5749 = ~n4750 & n4752 ;
  assign n5750 = n4757 & ~n5749 ;
  assign n5751 = n4209 & n5750 ;
  assign n5752 = ~n4209 & ~n5750 ;
  assign n5753 = ~n5751 & ~n5752 ;
  assign n5754 = n3788 & ~n5753 ;
  assign n5755 = ~n5748 & ~n5754 ;
  assign n5756 = ~n3177 & ~n5755 ;
  assign n5765 = n3322 & n3343 ;
  assign n5766 = ~n3121 & n5765 ;
  assign n5767 = n3102 & ~n5766 ;
  assign n5768 = ~n3102 & n5766 ;
  assign n5769 = ~n5767 & ~n5768 ;
  assign n5770 = n3788 & n5769 ;
  assign n5771 = ~n5748 & ~n5770 ;
  assign n5772 = n3355 & ~n5771 ;
  assign n5773 = ~n3112 & n3394 ;
  assign n5774 = n3088 & ~n5773 ;
  assign n5775 = ~n3088 & n5773 ;
  assign n5776 = ~n5774 & ~n5775 ;
  assign n5777 = ~n2058 & ~n5776 ;
  assign n5778 = n2058 & n3130 ;
  assign n5779 = ~n5777 & ~n5778 ;
  assign n5780 = n3788 & n5779 ;
  assign n5781 = ~n5748 & ~n5780 ;
  assign n5782 = n3411 & ~n5781 ;
  assign n5764 = n3108 & ~n3962 ;
  assign n5783 = n3102 & ~n3965 ;
  assign n5784 = ~n5764 & ~n5783 ;
  assign n5785 = ~n5782 & n5784 ;
  assign n5786 = ~n5772 & n5785 ;
  assign n5787 = ~n5756 & n5786 ;
  assign n5788 = ~n5763 & n5787 ;
  assign n5789 = n2026 & ~n5788 ;
  assign n5790 = ~n5747 & ~n5789 ;
  assign n5791 = \P1_state_reg[0]/NET0131  & ~n5790 ;
  assign n5745 = ~\P1_state_reg[0]/NET0131  & \P2_reg3_reg[22]/NET0131  ;
  assign n5746 = n3108 & n3976 ;
  assign n5792 = ~n5745 & ~n5746 ;
  assign n5793 = ~n5791 & n5792 ;
  assign n5803 = ~n825 & n3708 ;
  assign n5805 = ~n692 & n5803 ;
  assign n5804 = n692 & ~n5803 ;
  assign n5806 = n3712 & ~n5804 ;
  assign n5807 = ~n5805 & n5806 ;
  assign n5794 = n692 & n1880 ;
  assign n5795 = n3585 & n3589 ;
  assign n5796 = n3586 & n5795 ;
  assign n5797 = n4473 & n5796 ;
  assign n5798 = ~n831 & n3596 ;
  assign n5799 = n5797 & n5798 ;
  assign n5800 = n1936 & ~n3567 ;
  assign n5801 = ~n750 & n5800 ;
  assign n5802 = ~n5799 & n5801 ;
  assign n5808 = ~n5794 & ~n5802 ;
  assign n5809 = ~n5807 & n5808 ;
  assign n5810 = n3466 & ~n5809 ;
  assign n5811 = ~n3720 & ~n5810 ;
  assign n5812 = n3435 & ~n3447 ;
  assign n5813 = ~n5811 & n5812 ;
  assign n5814 = ~n1763 & ~n3466 ;
  assign n5815 = ~n3716 & n5812 ;
  assign n5816 = ~n5814 & n5815 ;
  assign n5817 = \P1_reg2_reg[31]/NET0131  & ~n5816 ;
  assign n5818 = ~n5813 & ~n5817 ;
  assign n5819 = \P2_reg0_reg[25]/NET0131  & ~n1983 ;
  assign n5820 = \P2_reg0_reg[25]/NET0131  & n2024 ;
  assign n5821 = \P2_reg0_reg[25]/NET0131  & ~n2040 ;
  assign n5825 = n2040 & ~n4609 ;
  assign n5826 = ~n5821 & ~n5825 ;
  assign n5827 = ~n3320 & ~n5826 ;
  assign n5822 = n2040 & ~n4595 ;
  assign n5823 = ~n5821 & ~n5822 ;
  assign n5824 = ~n3177 & ~n5823 ;
  assign n5829 = n2040 & n4617 ;
  assign n5830 = ~n5821 & ~n5829 ;
  assign n5831 = n3355 & ~n5830 ;
  assign n5828 = n2040 & ~n4928 ;
  assign n5832 = ~n3416 & n3423 ;
  assign n5833 = \P2_reg0_reg[25]/NET0131  & ~n5832 ;
  assign n5834 = ~n5828 & ~n5833 ;
  assign n5835 = ~n5831 & n5834 ;
  assign n5836 = ~n5824 & n5835 ;
  assign n5837 = ~n5827 & n5836 ;
  assign n5838 = n2026 & ~n5837 ;
  assign n5839 = ~n5820 & ~n5838 ;
  assign n5840 = \P1_state_reg[0]/NET0131  & ~n5839 ;
  assign n5841 = ~n5819 & ~n5840 ;
  assign n5842 = \P2_reg0_reg[26]/NET0131  & ~n1983 ;
  assign n5843 = \P2_reg0_reg[26]/NET0131  & ~n2040 ;
  assign n5844 = n2040 & ~n4732 ;
  assign n5845 = ~n5843 & ~n5844 ;
  assign n5846 = ~n3320 & ~n5845 ;
  assign n5847 = n2040 & ~n4764 ;
  assign n5848 = ~n5843 & ~n5847 ;
  assign n5849 = ~n3177 & ~n5848 ;
  assign n5850 = n2040 & ~n4962 ;
  assign n5851 = \P2_reg0_reg[26]/NET0131  & ~n3426 ;
  assign n5852 = ~n5850 & ~n5851 ;
  assign n5853 = ~n5849 & n5852 ;
  assign n5854 = ~n5846 & n5853 ;
  assign n5855 = n2026 & ~n5854 ;
  assign n5856 = \P2_reg0_reg[26]/NET0131  & n2024 ;
  assign n5857 = ~n5855 & ~n5856 ;
  assign n5858 = \P1_state_reg[0]/NET0131  & ~n5857 ;
  assign n5859 = ~n5842 & ~n5858 ;
  assign n5860 = n2040 & n5287 ;
  assign n5861 = n3421 & n5860 ;
  assign n5862 = \P2_reg0_reg[31]/NET0131  & ~n5861 ;
  assign n5863 = n3355 & n5282 ;
  assign n5864 = n5278 & ~n5863 ;
  assign n5865 = n5860 & ~n5864 ;
  assign n5866 = ~n5862 & ~n5865 ;
  assign n5867 = \P1_reg2_reg[25]/NET0131  & ~n3435 ;
  assign n5868 = \P1_reg2_reg[25]/NET0131  & n3448 ;
  assign n5869 = \P1_reg2_reg[25]/NET0131  & ~n3466 ;
  assign n5880 = n3466 & n4689 ;
  assign n5881 = ~n5869 & ~n5880 ;
  assign n5882 = n3712 & ~n5881 ;
  assign n5877 = n3466 & n4682 ;
  assign n5878 = ~n5869 & ~n5877 ;
  assign n5879 = n1936 & ~n5878 ;
  assign n5884 = \P1_reg2_reg[25]/NET0131  & ~n3718 ;
  assign n5876 = n3466 & n5304 ;
  assign n5883 = n1034 & n1763 ;
  assign n5885 = ~n5876 & ~n5883 ;
  assign n5886 = ~n5884 & n5885 ;
  assign n5887 = ~n5879 & n5886 ;
  assign n5888 = ~n5882 & n5887 ;
  assign n5870 = n3466 & ~n4658 ;
  assign n5871 = ~n5869 & ~n5870 ;
  assign n5872 = ~n3677 & ~n5871 ;
  assign n5873 = n3466 & ~n4672 ;
  assign n5874 = ~n5869 & ~n5873 ;
  assign n5875 = ~n3563 & ~n5874 ;
  assign n5889 = ~n5872 & ~n5875 ;
  assign n5890 = n5888 & n5889 ;
  assign n5891 = n3450 & ~n5890 ;
  assign n5892 = ~n5868 & ~n5891 ;
  assign n5893 = \P1_state_reg[0]/NET0131  & ~n5892 ;
  assign n5894 = ~n5867 & ~n5893 ;
  assign n5895 = \P1_reg2_reg[26]/NET0131  & ~n3435 ;
  assign n5896 = \P1_reg2_reg[26]/NET0131  & n3448 ;
  assign n5897 = \P1_reg2_reg[26]/NET0131  & ~n3466 ;
  assign n5898 = ~n978 & ~n5797 ;
  assign n5899 = n978 & n5797 ;
  assign n5900 = ~n5898 & ~n5899 ;
  assign n5901 = ~n537 & ~n5900 ;
  assign n5902 = n537 & ~n1038 ;
  assign n5903 = ~n5901 & ~n5902 ;
  assign n5904 = n3466 & ~n5903 ;
  assign n5905 = ~n5897 & ~n5904 ;
  assign n5906 = n1936 & ~n5905 ;
  assign n5907 = n997 & ~n4688 ;
  assign n5908 = ~n3704 & ~n5907 ;
  assign n5909 = n3712 & n5908 ;
  assign n5910 = n997 & n1880 ;
  assign n5911 = ~n5909 & ~n5910 ;
  assign n5912 = n3466 & ~n5911 ;
  assign n5913 = ~n3466 & n3712 ;
  assign n5914 = n3718 & ~n5913 ;
  assign n5915 = \P1_reg2_reg[26]/NET0131  & ~n5914 ;
  assign n5916 = n1002 & n1763 ;
  assign n5952 = ~n5915 & ~n5916 ;
  assign n5953 = ~n5912 & n5952 ;
  assign n5954 = ~n5906 & n5953 ;
  assign n5917 = n1300 & n1338 ;
  assign n5918 = n1376 & n1429 ;
  assign n5919 = n5917 & n5918 ;
  assign n5920 = ~n5501 & n5919 ;
  assign n5922 = n1376 & n1719 ;
  assign n5923 = ~n1706 & ~n5922 ;
  assign n5924 = n5917 & ~n5923 ;
  assign n5921 = n1300 & n1709 ;
  assign n5925 = ~n1066 & ~n5921 ;
  assign n5926 = ~n5924 & n5925 ;
  assign n5927 = ~n5920 & n5926 ;
  assign n5928 = n1809 & ~n5927 ;
  assign n5929 = ~n1809 & n5927 ;
  assign n5930 = ~n5928 & ~n5929 ;
  assign n5931 = n3466 & ~n5930 ;
  assign n5932 = ~n5897 & ~n5931 ;
  assign n5933 = ~n3677 & ~n5932 ;
  assign n5934 = n4012 & n4032 ;
  assign n5935 = ~n1836 & n4433 ;
  assign n5936 = n5934 & n5935 ;
  assign n5937 = ~n5524 & n5936 ;
  assign n5938 = n4027 & n4032 ;
  assign n5939 = n4039 & ~n5938 ;
  assign n5940 = n5935 & ~n5939 ;
  assign n5941 = ~n1816 & ~n4042 ;
  assign n5942 = n4045 & ~n5941 ;
  assign n5943 = ~n1810 & ~n5942 ;
  assign n5944 = ~n5940 & ~n5943 ;
  assign n5945 = ~n5937 & n5944 ;
  assign n5946 = n1809 & n5945 ;
  assign n5947 = ~n1809 & ~n5945 ;
  assign n5948 = ~n5946 & ~n5947 ;
  assign n5949 = n3466 & ~n5948 ;
  assign n5950 = ~n5897 & ~n5949 ;
  assign n5951 = ~n3563 & ~n5950 ;
  assign n5955 = ~n5933 & ~n5951 ;
  assign n5956 = n5954 & n5955 ;
  assign n5957 = n3450 & ~n5956 ;
  assign n5958 = ~n5896 & ~n5957 ;
  assign n5959 = \P1_state_reg[0]/NET0131  & ~n5958 ;
  assign n5960 = ~n5895 & ~n5959 ;
  assign n5961 = n3421 & n5287 ;
  assign n5962 = n3733 & n5961 ;
  assign n5963 = \P2_reg1_reg[31]/NET0131  & ~n5962 ;
  assign n5964 = n3733 & n5287 ;
  assign n5965 = ~n5864 & n5964 ;
  assign n5966 = ~n5963 & ~n5965 ;
  assign n5967 = \P1_reg0_reg[24]/NET0131  & ~n3435 ;
  assign n5968 = \P1_reg0_reg[24]/NET0131  & n3448 ;
  assign n5969 = \P1_reg0_reg[24]/NET0131  & ~n4396 ;
  assign n5970 = n4396 & ~n5172 ;
  assign n5971 = ~n5969 & ~n5970 ;
  assign n5972 = ~n3563 & ~n5971 ;
  assign n5978 = n4396 & n5190 ;
  assign n5979 = ~n5969 & ~n5978 ;
  assign n5980 = n3712 & ~n5979 ;
  assign n5976 = \P1_reg0_reg[24]/NET0131  & ~n4493 ;
  assign n5977 = n4396 & n5206 ;
  assign n5984 = ~n5976 & ~n5977 ;
  assign n5985 = ~n5980 & n5984 ;
  assign n5986 = ~n5972 & n5985 ;
  assign n5973 = n4396 & n5200 ;
  assign n5974 = ~n5969 & ~n5973 ;
  assign n5975 = n1936 & ~n5974 ;
  assign n5981 = n4396 & ~n5184 ;
  assign n5982 = ~n5969 & ~n5981 ;
  assign n5983 = ~n3677 & ~n5982 ;
  assign n5987 = ~n5975 & ~n5983 ;
  assign n5988 = n5986 & n5987 ;
  assign n5989 = n3450 & ~n5988 ;
  assign n5990 = ~n5968 & ~n5989 ;
  assign n5991 = \P1_state_reg[0]/NET0131  & ~n5990 ;
  assign n5992 = ~n5967 & ~n5991 ;
  assign n5993 = \P1_reg0_reg[26]/NET0131  & ~n3435 ;
  assign n5994 = \P1_reg0_reg[26]/NET0131  & n3448 ;
  assign n5995 = \P1_reg0_reg[26]/NET0131  & ~n4396 ;
  assign n5996 = n4396 & ~n5903 ;
  assign n5997 = ~n5995 & ~n5996 ;
  assign n5998 = n1936 & ~n5997 ;
  assign n5999 = \P1_reg0_reg[26]/NET0131  & ~n4494 ;
  assign n6000 = n4396 & ~n5911 ;
  assign n6007 = ~n5999 & ~n6000 ;
  assign n6008 = ~n5998 & n6007 ;
  assign n6001 = n4396 & ~n5948 ;
  assign n6002 = ~n5995 & ~n6001 ;
  assign n6003 = ~n3563 & ~n6002 ;
  assign n6004 = n4396 & ~n5930 ;
  assign n6005 = ~n5995 & ~n6004 ;
  assign n6006 = ~n3677 & ~n6005 ;
  assign n6009 = ~n6003 & ~n6006 ;
  assign n6010 = n6008 & n6009 ;
  assign n6011 = n3450 & ~n6010 ;
  assign n6012 = ~n5994 & ~n6011 ;
  assign n6013 = \P1_state_reg[0]/NET0131  & ~n6012 ;
  assign n6014 = ~n5993 & ~n6013 ;
  assign n6015 = \P1_reg1_reg[22]/NET0131  & ~n3435 ;
  assign n6016 = \P1_reg1_reg[22]/NET0131  & n3448 ;
  assign n6017 = \P1_reg1_reg[22]/NET0131  & ~n4532 ;
  assign n6031 = ~n5516 & n5519 ;
  assign n6032 = n5508 & n5934 ;
  assign n6033 = ~n6031 & n6032 ;
  assign n6030 = ~n5522 & n5934 ;
  assign n6034 = n5939 & ~n6030 ;
  assign n6035 = ~n6033 & n6034 ;
  assign n6036 = n1838 & n6035 ;
  assign n6037 = ~n1838 & ~n6035 ;
  assign n6038 = ~n6036 & ~n6037 ;
  assign n6039 = n4532 & ~n6038 ;
  assign n6040 = ~n6017 & ~n6039 ;
  assign n6041 = ~n3563 & ~n6040 ;
  assign n6019 = ~n5493 & n5496 ;
  assign n6020 = n5486 & n5918 ;
  assign n6021 = ~n6019 & n6020 ;
  assign n6018 = ~n5499 & n5918 ;
  assign n6022 = n5923 & ~n6018 ;
  assign n6023 = ~n6021 & n6022 ;
  assign n6024 = n1838 & n6023 ;
  assign n6025 = ~n1838 & ~n6023 ;
  assign n6026 = ~n6024 & ~n6025 ;
  assign n6027 = n4532 & n6026 ;
  assign n6028 = ~n6017 & ~n6027 ;
  assign n6029 = ~n3677 & ~n6028 ;
  assign n6043 = n537 & ~n1356 ;
  assign n6044 = ~n1318 & n5795 ;
  assign n6045 = n1336 & ~n6044 ;
  assign n6046 = ~n537 & ~n5796 ;
  assign n6047 = ~n6045 & n6046 ;
  assign n6048 = ~n6043 & ~n6047 ;
  assign n6049 = n4532 & ~n6048 ;
  assign n6050 = ~n6017 & ~n6049 ;
  assign n6051 = n1936 & ~n6050 ;
  assign n6042 = \P1_reg1_reg[22]/NET0131  & ~n4573 ;
  assign n6052 = ~n1346 & n3698 ;
  assign n6053 = n1309 & ~n6052 ;
  assign n6054 = ~n3700 & ~n6053 ;
  assign n6055 = n3712 & n6054 ;
  assign n6056 = n1309 & n1880 ;
  assign n6057 = ~n6055 & ~n6056 ;
  assign n6058 = n4532 & ~n6057 ;
  assign n6059 = ~n6042 & ~n6058 ;
  assign n6060 = ~n6051 & n6059 ;
  assign n6061 = ~n6029 & n6060 ;
  assign n6062 = ~n6041 & n6061 ;
  assign n6063 = n3450 & ~n6062 ;
  assign n6064 = ~n6016 & ~n6063 ;
  assign n6065 = \P1_state_reg[0]/NET0131  & ~n6064 ;
  assign n6066 = ~n6015 & ~n6065 ;
  assign n6067 = \P1_reg1_reg[26]/NET0131  & ~n3435 ;
  assign n6068 = \P1_reg1_reg[26]/NET0131  & n3448 ;
  assign n6069 = \P1_reg1_reg[26]/NET0131  & ~n4532 ;
  assign n6070 = n4532 & ~n5903 ;
  assign n6071 = ~n6069 & ~n6070 ;
  assign n6072 = n1936 & ~n6071 ;
  assign n6073 = \P1_reg1_reg[26]/NET0131  & ~n4573 ;
  assign n6074 = n4532 & ~n5911 ;
  assign n6081 = ~n6073 & ~n6074 ;
  assign n6082 = ~n6072 & n6081 ;
  assign n6075 = n4532 & ~n5948 ;
  assign n6076 = ~n6069 & ~n6075 ;
  assign n6077 = ~n3563 & ~n6076 ;
  assign n6078 = n4532 & ~n5930 ;
  assign n6079 = ~n6069 & ~n6078 ;
  assign n6080 = ~n3677 & ~n6079 ;
  assign n6083 = ~n6077 & ~n6080 ;
  assign n6084 = n6082 & n6083 ;
  assign n6085 = n3450 & ~n6084 ;
  assign n6086 = ~n6068 & ~n6085 ;
  assign n6087 = \P1_state_reg[0]/NET0131  & ~n6086 ;
  assign n6088 = ~n6067 & ~n6087 ;
  assign n6091 = n1170 & n3448 ;
  assign n6093 = n1170 & ~n3980 ;
  assign n6094 = n1146 & ~n4070 ;
  assign n6095 = ~n3583 & ~n6094 ;
  assign n6096 = ~n537 & ~n6095 ;
  assign n6097 = n537 & n1207 ;
  assign n6098 = ~n6096 & ~n6097 ;
  assign n6099 = n3980 & n6098 ;
  assign n6100 = ~n6093 & ~n6099 ;
  assign n6101 = n1936 & ~n6100 ;
  assign n6108 = n1796 & ~n4088 ;
  assign n6109 = ~n1796 & n4088 ;
  assign n6110 = ~n6108 & ~n6109 ;
  assign n6111 = n3980 & ~n6110 ;
  assign n6112 = ~n6093 & ~n6111 ;
  assign n6113 = ~n3677 & ~n6112 ;
  assign n6102 = n1796 & ~n4007 ;
  assign n6103 = ~n1796 & n4007 ;
  assign n6104 = ~n6102 & ~n6103 ;
  assign n6105 = n3980 & n6104 ;
  assign n6106 = ~n6093 & ~n6105 ;
  assign n6107 = ~n3563 & ~n6106 ;
  assign n6114 = ~n1233 & n3687 ;
  assign n6115 = ~n1198 & n6114 ;
  assign n6116 = n1165 & ~n6115 ;
  assign n6117 = ~n3690 & ~n6116 ;
  assign n6118 = n3980 & n6117 ;
  assign n6119 = ~n6093 & ~n6118 ;
  assign n6120 = n3712 & ~n6119 ;
  assign n6092 = n1165 & ~n4067 ;
  assign n6121 = n1170 & ~n4064 ;
  assign n6122 = ~n6092 & ~n6121 ;
  assign n6123 = ~n6120 & n6122 ;
  assign n6124 = ~n6107 & n6123 ;
  assign n6125 = ~n6113 & n6124 ;
  assign n6126 = ~n6101 & n6125 ;
  assign n6127 = n3450 & ~n6126 ;
  assign n6128 = ~n6091 & ~n6127 ;
  assign n6129 = \P1_state_reg[0]/NET0131  & ~n6128 ;
  assign n6089 = \P1_reg3_reg[12]/NET0131  & ~\P1_state_reg[0]/NET0131  ;
  assign n6090 = n1170 & n1953 ;
  assign n6130 = ~n6089 & ~n6090 ;
  assign n6131 = ~n6129 & n6130 ;
  assign n6134 = n1471 & n3448 ;
  assign n6136 = n1471 & ~n3980 ;
  assign n6145 = n1452 & ~n4073 ;
  assign n6146 = ~n5195 & ~n6145 ;
  assign n6147 = ~n537 & ~n6146 ;
  assign n6148 = n537 & n1094 ;
  assign n6149 = ~n6147 & ~n6148 ;
  assign n6150 = n3980 & n6149 ;
  assign n6151 = ~n6136 & ~n6150 ;
  assign n6152 = n1936 & ~n6151 ;
  assign n6137 = ~n4007 & n4010 ;
  assign n6138 = n4021 & ~n6137 ;
  assign n6139 = n1785 & n6138 ;
  assign n6140 = ~n1785 & ~n6138 ;
  assign n6141 = ~n6139 & ~n6140 ;
  assign n6142 = n3980 & ~n6141 ;
  assign n6143 = ~n6136 & ~n6142 ;
  assign n6144 = ~n3563 & ~n6143 ;
  assign n6153 = ~n1750 & n1785 ;
  assign n6154 = n1750 & ~n1785 ;
  assign n6155 = ~n6153 & ~n6154 ;
  assign n6156 = n3980 & ~n6155 ;
  assign n6157 = ~n6136 & ~n6156 ;
  assign n6158 = ~n3677 & ~n6157 ;
  assign n6159 = n1466 & ~n5441 ;
  assign n6160 = ~n5442 & ~n6159 ;
  assign n6161 = n3712 & n6160 ;
  assign n6162 = n3980 & n6161 ;
  assign n6135 = n1471 & ~n4910 ;
  assign n6163 = n1466 & ~n4067 ;
  assign n6164 = ~n6135 & ~n6163 ;
  assign n6165 = ~n6162 & n6164 ;
  assign n6166 = ~n6158 & n6165 ;
  assign n6167 = ~n6144 & n6166 ;
  assign n6168 = ~n6152 & n6167 ;
  assign n6169 = n3450 & ~n6168 ;
  assign n6170 = ~n6134 & ~n6169 ;
  assign n6171 = \P1_state_reg[0]/NET0131  & ~n6170 ;
  assign n6132 = \P1_reg3_reg[16]/NET0131  & ~\P1_state_reg[0]/NET0131  ;
  assign n6133 = n1471 & n1953 ;
  assign n6172 = ~n6132 & ~n6133 ;
  assign n6173 = ~n6171 & n6172 ;
  assign n6176 = n2024 & n2709 ;
  assign n6178 = n2709 & ~n3788 ;
  assign n6179 = ~n2688 & n3383 ;
  assign n6180 = ~n2715 & n6179 ;
  assign n6181 = n2880 & ~n6180 ;
  assign n6182 = ~n2880 & n6180 ;
  assign n6183 = ~n6181 & ~n6182 ;
  assign n6184 = ~n2058 & ~n6183 ;
  assign n6185 = n2058 & n2688 ;
  assign n6186 = ~n6184 & ~n6185 ;
  assign n6187 = n3788 & n6186 ;
  assign n6188 = ~n6178 & ~n6187 ;
  assign n6189 = n3411 & ~n6188 ;
  assign n6196 = ~n3839 & n4212 ;
  assign n6197 = n3839 & ~n4212 ;
  assign n6198 = ~n6196 & ~n6197 ;
  assign n6199 = n3788 & ~n6198 ;
  assign n6200 = ~n6178 & ~n6199 ;
  assign n6201 = ~n3320 & ~n6200 ;
  assign n6190 = ~n3893 & n4212 ;
  assign n6191 = n3893 & ~n4212 ;
  assign n6192 = ~n6190 & ~n6191 ;
  assign n6193 = n3788 & n6192 ;
  assign n6194 = ~n6178 & ~n6193 ;
  assign n6195 = ~n3177 & ~n6194 ;
  assign n6202 = n2731 & ~n3336 ;
  assign n6203 = ~n3337 & ~n6202 ;
  assign n6204 = n3355 & n6203 ;
  assign n6205 = n3788 & n6204 ;
  assign n6177 = n2709 & ~n5698 ;
  assign n6206 = n2731 & ~n3965 ;
  assign n6207 = ~n6177 & ~n6206 ;
  assign n6208 = ~n6205 & n6207 ;
  assign n6209 = ~n6195 & n6208 ;
  assign n6210 = ~n6201 & n6209 ;
  assign n6211 = ~n6189 & n6210 ;
  assign n6212 = n2026 & ~n6211 ;
  assign n6213 = ~n6176 & ~n6212 ;
  assign n6214 = \P1_state_reg[0]/NET0131  & ~n6213 ;
  assign n6174 = ~\P1_state_reg[0]/NET0131  & \P2_reg3_reg[12]/NET0131  ;
  assign n6175 = n2709 & n3976 ;
  assign n6215 = ~n6174 & ~n6175 ;
  assign n6216 = ~n6214 & n6215 ;
  assign n6219 = n2024 & n2797 ;
  assign n6221 = n2797 & ~n3788 ;
  assign n6244 = ~n4169 & n4211 ;
  assign n6245 = n4169 & ~n4211 ;
  assign n6246 = ~n6244 & ~n6245 ;
  assign n6247 = n3788 & ~n6246 ;
  assign n6248 = ~n6221 & ~n6247 ;
  assign n6249 = ~n3320 & ~n6248 ;
  assign n6239 = n2818 & ~n5574 ;
  assign n6240 = ~n5575 & ~n6239 ;
  assign n6241 = n3788 & n6240 ;
  assign n6242 = ~n6221 & ~n6241 ;
  assign n6243 = n3355 & ~n6242 ;
  assign n6220 = n2797 & ~n3962 ;
  assign n6238 = n2818 & ~n3965 ;
  assign n6250 = ~n6220 & ~n6238 ;
  assign n6251 = ~n6243 & n6250 ;
  assign n6252 = ~n6249 & n6251 ;
  assign n6222 = ~n3893 & n3896 ;
  assign n6223 = n3907 & ~n6222 ;
  assign n6224 = n4211 & n6223 ;
  assign n6225 = ~n4211 & ~n6223 ;
  assign n6226 = ~n6224 & ~n6225 ;
  assign n6227 = n3788 & ~n6226 ;
  assign n6228 = ~n6221 & ~n6227 ;
  assign n6229 = ~n3177 & ~n6228 ;
  assign n6230 = n2379 & ~n5565 ;
  assign n6231 = ~n5566 & ~n6230 ;
  assign n6232 = ~n2058 & ~n6231 ;
  assign n6233 = n2058 & n2828 ;
  assign n6234 = ~n6232 & ~n6233 ;
  assign n6235 = n3788 & n6234 ;
  assign n6236 = ~n6221 & ~n6235 ;
  assign n6237 = n3411 & ~n6236 ;
  assign n6253 = ~n6229 & ~n6237 ;
  assign n6254 = n6252 & n6253 ;
  assign n6255 = n2026 & ~n6254 ;
  assign n6256 = ~n6219 & ~n6255 ;
  assign n6257 = \P1_state_reg[0]/NET0131  & ~n6256 ;
  assign n6217 = n2797 & n3976 ;
  assign n6218 = ~\P1_state_reg[0]/NET0131  & \P2_reg3_reg[16]/NET0131  ;
  assign n6258 = ~n6217 & ~n6218 ;
  assign n6259 = ~n6257 & n6258 ;
  assign n6262 = n1314 & n3448 ;
  assign n6263 = n1314 & ~n3980 ;
  assign n6267 = n3980 & n6026 ;
  assign n6268 = ~n6263 & ~n6267 ;
  assign n6269 = ~n3677 & ~n6268 ;
  assign n6264 = n3980 & ~n6038 ;
  assign n6265 = ~n6263 & ~n6264 ;
  assign n6266 = ~n3563 & ~n6265 ;
  assign n6271 = n3980 & ~n6048 ;
  assign n6272 = ~n6263 & ~n6271 ;
  assign n6273 = n1936 & ~n6272 ;
  assign n6274 = n3980 & n6055 ;
  assign n6270 = n1314 & ~n4910 ;
  assign n6275 = n1309 & ~n4067 ;
  assign n6276 = ~n6270 & ~n6275 ;
  assign n6277 = ~n6274 & n6276 ;
  assign n6278 = ~n6273 & n6277 ;
  assign n6279 = ~n6266 & n6278 ;
  assign n6280 = ~n6269 & n6279 ;
  assign n6281 = n3450 & ~n6280 ;
  assign n6282 = ~n6262 & ~n6281 ;
  assign n6283 = \P1_state_reg[0]/NET0131  & ~n6282 ;
  assign n6260 = \P1_reg3_reg[22]/NET0131  & ~\P1_state_reg[0]/NET0131  ;
  assign n6261 = n1314 & n1953 ;
  assign n6284 = ~n6260 & ~n6261 ;
  assign n6285 = ~n6283 & n6284 ;
  assign n6286 = n2024 & n3126 ;
  assign n6301 = n3121 & ~n5765 ;
  assign n6302 = n3355 & ~n5766 ;
  assign n6303 = ~n6301 & n6302 ;
  assign n6296 = n3112 & ~n3394 ;
  assign n6297 = ~n5773 & ~n6296 ;
  assign n6298 = ~n2058 & ~n6297 ;
  assign n6295 = n2058 & n2368 ;
  assign n6299 = n3411 & ~n6295 ;
  assign n6300 = ~n6298 & n6299 ;
  assign n6305 = n3304 & n4216 ;
  assign n6304 = ~n3304 & ~n4216 ;
  assign n6306 = ~n3320 & ~n6304 ;
  assign n6307 = ~n6305 & n6306 ;
  assign n6308 = ~n6300 & ~n6307 ;
  assign n6309 = ~n6303 & n6308 ;
  assign n6310 = n3788 & ~n6309 ;
  assign n6288 = n2921 & n4216 ;
  assign n6289 = ~n2921 & ~n4216 ;
  assign n6290 = ~n6288 & ~n6289 ;
  assign n6291 = n3788 & n6290 ;
  assign n6292 = ~n3126 & ~n3788 ;
  assign n6293 = ~n3177 & ~n6292 ;
  assign n6294 = ~n6291 & n6293 ;
  assign n6287 = n3121 & ~n3965 ;
  assign n6311 = ~n3320 & ~n3788 ;
  assign n6312 = n3962 & ~n6311 ;
  assign n6313 = n3745 & ~n3788 ;
  assign n6314 = n6312 & ~n6313 ;
  assign n6315 = n3126 & ~n6314 ;
  assign n6316 = ~n6287 & ~n6315 ;
  assign n6317 = ~n6294 & n6316 ;
  assign n6318 = ~n6310 & n6317 ;
  assign n6319 = n2026 & ~n6318 ;
  assign n6320 = ~n6286 & ~n6319 ;
  assign n6321 = \P1_state_reg[0]/NET0131  & ~n6320 ;
  assign n6322 = n3126 & n3976 ;
  assign n6323 = ~\P1_state_reg[0]/NET0131  & \P2_reg3_reg[21]/NET0131  ;
  assign n6324 = ~n6322 & ~n6323 ;
  assign n6325 = ~n6321 & n6324 ;
  assign n6326 = \P2_reg2_reg[18]/NET0131  & ~n1983 ;
  assign n6327 = \P2_reg2_reg[18]/NET0131  & n2024 ;
  assign n6329 = \P2_reg2_reg[18]/NET0131  & ~n3758 ;
  assign n6330 = n2433 & ~n5577 ;
  assign n6331 = ~n3343 & ~n6330 ;
  assign n6332 = n3758 & n6331 ;
  assign n6333 = ~n6329 & ~n6332 ;
  assign n6334 = n3355 & ~n6333 ;
  assign n6341 = n4218 & ~n4719 ;
  assign n6342 = ~n4218 & n4719 ;
  assign n6343 = ~n6341 & ~n6342 ;
  assign n6344 = n3758 & ~n6343 ;
  assign n6345 = ~n6329 & ~n6344 ;
  assign n6346 = ~n3320 & ~n6345 ;
  assign n6335 = n4218 & ~n4750 ;
  assign n6336 = ~n4218 & n4750 ;
  assign n6337 = ~n6335 & ~n6336 ;
  assign n6338 = n3758 & n6337 ;
  assign n6339 = ~n6329 & ~n6338 ;
  assign n6340 = ~n3177 & ~n6339 ;
  assign n6347 = n2311 & ~n5563 ;
  assign n6348 = ~n5618 & ~n6347 ;
  assign n6349 = ~n2058 & ~n6348 ;
  assign n6350 = n2058 & n2379 ;
  assign n6351 = ~n6349 & ~n6350 ;
  assign n6352 = n3758 & n6351 ;
  assign n6353 = ~n6329 & ~n6352 ;
  assign n6354 = n3411 & ~n6353 ;
  assign n6356 = n2433 & n3358 ;
  assign n6357 = n3758 & n6356 ;
  assign n6328 = \P2_reg2_reg[18]/NET0131  & ~n3774 ;
  assign n6355 = n2438 & n3420 ;
  assign n6358 = ~n6328 & ~n6355 ;
  assign n6359 = ~n6357 & n6358 ;
  assign n6360 = ~n6354 & n6359 ;
  assign n6361 = ~n6340 & n6360 ;
  assign n6362 = ~n6346 & n6361 ;
  assign n6363 = ~n6334 & n6362 ;
  assign n6364 = n2026 & ~n6363 ;
  assign n6365 = ~n6327 & ~n6364 ;
  assign n6366 = \P1_state_reg[0]/NET0131  & ~n6365 ;
  assign n6367 = ~n6326 & ~n6366 ;
  assign n6368 = n4532 & n5812 ;
  assign n6369 = ~n5809 & n6368 ;
  assign n6370 = n4491 & n6368 ;
  assign n6371 = \P1_reg1_reg[31]/NET0131  & ~n6370 ;
  assign n6372 = ~n6369 & ~n6371 ;
  assign n6373 = \P2_reg0_reg[22]/NET0131  & ~n1983 ;
  assign n6374 = \P2_reg0_reg[22]/NET0131  & n2024 ;
  assign n6382 = \P2_reg0_reg[22]/NET0131  & ~n2040 ;
  assign n6386 = n2040 & n5760 ;
  assign n6387 = ~n6382 & ~n6386 ;
  assign n6388 = ~n3320 & ~n6387 ;
  assign n6383 = n2040 & ~n5753 ;
  assign n6384 = ~n6382 & ~n6383 ;
  assign n6385 = ~n3177 & ~n6384 ;
  assign n6376 = n3355 & n5769 ;
  assign n6375 = n3411 & n5779 ;
  assign n6377 = n3102 & n3358 ;
  assign n6378 = ~n6375 & ~n6377 ;
  assign n6379 = ~n6376 & n6378 ;
  assign n6380 = n2040 & ~n6379 ;
  assign n6381 = \P2_reg0_reg[22]/NET0131  & ~n3426 ;
  assign n6389 = ~n6380 & ~n6381 ;
  assign n6390 = ~n6385 & n6389 ;
  assign n6391 = ~n6388 & n6390 ;
  assign n6392 = n2026 & ~n6391 ;
  assign n6393 = ~n6374 & ~n6392 ;
  assign n6394 = \P1_state_reg[0]/NET0131  & ~n6393 ;
  assign n6395 = ~n6373 & ~n6394 ;
  assign n6396 = \P1_reg2_reg[18]/NET0131  & ~n3435 ;
  assign n6397 = \P1_reg2_reg[18]/NET0131  & n3448 ;
  assign n6399 = \P1_reg2_reg[18]/NET0131  & ~n3466 ;
  assign n6400 = n3466 & n5482 ;
  assign n6401 = ~n6399 & ~n6400 ;
  assign n6402 = n3712 & ~n6401 ;
  assign n6413 = n1394 & n1880 ;
  assign n6414 = n3466 & n6413 ;
  assign n6398 = \P1_reg2_reg[18]/NET0131  & ~n3718 ;
  assign n6412 = n1399 & n1763 ;
  assign n6415 = ~n6398 & ~n6412 ;
  assign n6416 = ~n6414 & n6415 ;
  assign n6417 = ~n6402 & n6416 ;
  assign n6409 = n3466 & ~n5536 ;
  assign n6410 = ~n6399 & ~n6409 ;
  assign n6411 = n1936 & ~n6410 ;
  assign n6403 = n3466 & ~n5504 ;
  assign n6404 = ~n6399 & ~n6403 ;
  assign n6405 = ~n3677 & ~n6404 ;
  assign n6406 = n3466 & n5527 ;
  assign n6407 = ~n6399 & ~n6406 ;
  assign n6408 = ~n3563 & ~n6407 ;
  assign n6418 = ~n6405 & ~n6408 ;
  assign n6419 = ~n6411 & n6418 ;
  assign n6420 = n6417 & n6419 ;
  assign n6421 = n3450 & ~n6420 ;
  assign n6422 = ~n6397 & ~n6421 ;
  assign n6423 = \P1_state_reg[0]/NET0131  & ~n6422 ;
  assign n6424 = ~n6396 & ~n6423 ;
  assign n6425 = \P1_reg2_reg[17]/NET0131  & ~n3435 ;
  assign n6426 = \P1_reg2_reg[17]/NET0131  & n3448 ;
  assign n6427 = \P1_reg2_reg[17]/NET0131  & ~n3466 ;
  assign n6437 = n3466 & n5462 ;
  assign n6438 = ~n6427 & ~n6437 ;
  assign n6439 = n1936 & ~n6438 ;
  assign n6431 = n3466 & n5445 ;
  assign n6432 = ~n6427 & ~n6431 ;
  assign n6433 = n3712 & ~n6432 ;
  assign n6442 = n1443 & n1880 ;
  assign n6443 = n3466 & n6442 ;
  assign n6440 = \P1_reg2_reg[17]/NET0131  & ~n3718 ;
  assign n6441 = n1447 & n1763 ;
  assign n6444 = ~n6440 & ~n6441 ;
  assign n6445 = ~n6443 & n6444 ;
  assign n6446 = ~n6433 & n6445 ;
  assign n6447 = ~n6439 & n6446 ;
  assign n6428 = n3466 & ~n5453 ;
  assign n6429 = ~n6427 & ~n6428 ;
  assign n6430 = ~n3563 & ~n6429 ;
  assign n6434 = n3466 & n5436 ;
  assign n6435 = ~n6427 & ~n6434 ;
  assign n6436 = ~n3677 & ~n6435 ;
  assign n6448 = ~n6430 & ~n6436 ;
  assign n6449 = n6447 & n6448 ;
  assign n6450 = n3450 & ~n6449 ;
  assign n6451 = ~n6426 & ~n6450 ;
  assign n6452 = \P1_state_reg[0]/NET0131  & ~n6451 ;
  assign n6453 = ~n6425 & ~n6452 ;
  assign n6454 = \P1_reg2_reg[19]/NET0131  & n3448 ;
  assign n6455 = \P1_reg2_reg[19]/NET0131  & ~n3466 ;
  assign n6456 = n3466 & ~n5654 ;
  assign n6457 = ~n6455 & ~n6456 ;
  assign n6458 = n1936 & ~n6457 ;
  assign n6463 = n3466 & ~n5667 ;
  assign n6464 = ~n6455 & ~n6463 ;
  assign n6465 = ~n3677 & ~n6464 ;
  assign n6460 = n3466 & n5661 ;
  assign n6461 = ~n6455 & ~n6460 ;
  assign n6462 = ~n3563 & ~n6461 ;
  assign n6466 = n3466 & n5673 ;
  assign n6467 = ~n6455 & ~n6466 ;
  assign n6468 = n3712 & ~n6467 ;
  assign n6469 = n1418 & n3466 ;
  assign n6470 = ~n6455 & ~n6469 ;
  assign n6471 = n1880 & ~n6470 ;
  assign n6459 = n1423 & n1763 ;
  assign n6472 = \P1_reg2_reg[19]/NET0131  & n3716 ;
  assign n6473 = ~n6459 & ~n6472 ;
  assign n6474 = ~n6471 & n6473 ;
  assign n6475 = ~n6468 & n6474 ;
  assign n6476 = ~n6462 & n6475 ;
  assign n6477 = ~n6465 & n6476 ;
  assign n6478 = ~n6458 & n6477 ;
  assign n6479 = n3450 & ~n6478 ;
  assign n6480 = ~n6454 & ~n6479 ;
  assign n6481 = \P1_state_reg[0]/NET0131  & ~n6480 ;
  assign n6482 = \P1_reg2_reg[19]/NET0131  & ~n3435 ;
  assign n6483 = ~n6481 & ~n6482 ;
  assign n6484 = \P1_reg2_reg[20]/NET0131  & ~n3435 ;
  assign n6485 = \P1_reg2_reg[20]/NET0131  & n3448 ;
  assign n6486 = \P1_reg2_reg[20]/NET0131  & ~n3466 ;
  assign n6487 = n1356 & ~n5649 ;
  assign n6488 = n3589 & n5195 ;
  assign n6489 = ~n6487 & ~n6488 ;
  assign n6490 = ~n537 & ~n6489 ;
  assign n6491 = n537 & n1427 ;
  assign n6492 = ~n6490 & ~n6491 ;
  assign n6493 = n3466 & n6492 ;
  assign n6494 = ~n6486 & ~n6493 ;
  assign n6495 = n1936 & ~n6494 ;
  assign n6503 = n1828 & n4030 ;
  assign n6504 = ~n1828 & ~n4030 ;
  assign n6505 = ~n6503 & ~n6504 ;
  assign n6506 = n3466 & ~n6505 ;
  assign n6507 = ~n6486 & ~n6506 ;
  assign n6508 = ~n3563 & ~n6507 ;
  assign n6497 = n1828 & ~n4093 ;
  assign n6498 = ~n1828 & n4093 ;
  assign n6499 = ~n6497 & ~n6498 ;
  assign n6500 = n3466 & ~n6499 ;
  assign n6501 = ~n6486 & ~n6500 ;
  assign n6502 = ~n3677 & ~n6501 ;
  assign n6509 = n1365 & ~n5671 ;
  assign n6510 = ~n3698 & ~n6509 ;
  assign n6511 = n3466 & n6510 ;
  assign n6512 = ~n6486 & ~n6511 ;
  assign n6513 = n3712 & ~n6512 ;
  assign n6515 = n1365 & n1880 ;
  assign n6516 = n3466 & n6515 ;
  assign n6496 = \P1_reg2_reg[20]/NET0131  & ~n3718 ;
  assign n6514 = n1370 & n1763 ;
  assign n6517 = ~n6496 & ~n6514 ;
  assign n6518 = ~n6516 & n6517 ;
  assign n6519 = ~n6513 & n6518 ;
  assign n6520 = ~n6502 & n6519 ;
  assign n6521 = ~n6508 & n6520 ;
  assign n6522 = ~n6495 & n6521 ;
  assign n6523 = n3450 & ~n6522 ;
  assign n6524 = ~n6485 & ~n6523 ;
  assign n6525 = \P1_state_reg[0]/NET0131  & ~n6524 ;
  assign n6526 = ~n6484 & ~n6525 ;
  assign n6527 = \P2_reg1_reg[17]/NET0131  & ~n1983 ;
  assign n6528 = \P2_reg1_reg[17]/NET0131  & n2024 ;
  assign n6531 = \P2_reg1_reg[17]/NET0131  & ~n3733 ;
  assign n6532 = n3733 & n5558 ;
  assign n6533 = ~n6531 & ~n6532 ;
  assign n6534 = ~n3177 & ~n6533 ;
  assign n6541 = n3733 & n5586 ;
  assign n6542 = ~n6531 & ~n6541 ;
  assign n6543 = ~n3320 & ~n6542 ;
  assign n6529 = n2399 & n3358 ;
  assign n6530 = n3733 & n6529 ;
  assign n6544 = \P2_reg1_reg[17]/NET0131  & ~n3743 ;
  assign n6545 = ~n6530 & ~n6544 ;
  assign n6546 = ~n6543 & n6545 ;
  assign n6547 = ~n6534 & n6546 ;
  assign n6535 = n3733 & ~n5570 ;
  assign n6536 = ~n6531 & ~n6535 ;
  assign n6537 = n3411 & ~n6536 ;
  assign n6538 = n3733 & n5578 ;
  assign n6539 = ~n6531 & ~n6538 ;
  assign n6540 = n3355 & ~n6539 ;
  assign n6548 = ~n6537 & ~n6540 ;
  assign n6549 = n6547 & n6548 ;
  assign n6550 = n2026 & ~n6549 ;
  assign n6551 = ~n6528 & ~n6550 ;
  assign n6552 = \P1_state_reg[0]/NET0131  & ~n6551 ;
  assign n6553 = ~n6527 & ~n6552 ;
  assign n6554 = \P1_reg2_reg[22]/NET0131  & ~n3435 ;
  assign n6555 = \P1_reg2_reg[22]/NET0131  & n3448 ;
  assign n6556 = \P1_reg2_reg[22]/NET0131  & ~n3466 ;
  assign n6560 = n3466 & ~n6038 ;
  assign n6561 = ~n6556 & ~n6560 ;
  assign n6562 = ~n3563 & ~n6561 ;
  assign n6557 = n3466 & n6026 ;
  assign n6558 = ~n6556 & ~n6557 ;
  assign n6559 = ~n3677 & ~n6558 ;
  assign n6564 = n3466 & ~n6048 ;
  assign n6565 = ~n6556 & ~n6564 ;
  assign n6566 = n1936 & ~n6565 ;
  assign n6567 = n3466 & n6054 ;
  assign n6568 = ~n6556 & ~n6567 ;
  assign n6569 = n3712 & ~n6568 ;
  assign n6570 = n1309 & n3466 ;
  assign n6571 = ~n6556 & ~n6570 ;
  assign n6572 = n1880 & ~n6571 ;
  assign n6563 = \P1_reg2_reg[22]/NET0131  & n3716 ;
  assign n6573 = n1314 & n1763 ;
  assign n6574 = ~n6563 & ~n6573 ;
  assign n6575 = ~n6572 & n6574 ;
  assign n6576 = ~n6569 & n6575 ;
  assign n6577 = ~n6566 & n6576 ;
  assign n6578 = ~n6559 & n6577 ;
  assign n6579 = ~n6562 & n6578 ;
  assign n6580 = n3450 & ~n6579 ;
  assign n6581 = ~n6555 & ~n6580 ;
  assign n6582 = \P1_state_reg[0]/NET0131  & ~n6581 ;
  assign n6583 = ~n6554 & ~n6582 ;
  assign n6584 = \P2_reg1_reg[18]/NET0131  & ~n1983 ;
  assign n6585 = \P2_reg1_reg[18]/NET0131  & n2024 ;
  assign n6587 = \P2_reg1_reg[18]/NET0131  & ~n3733 ;
  assign n6588 = n3733 & n6331 ;
  assign n6589 = ~n6587 & ~n6588 ;
  assign n6590 = n3355 & ~n6589 ;
  assign n6594 = n3733 & ~n6343 ;
  assign n6595 = ~n6587 & ~n6594 ;
  assign n6596 = ~n3320 & ~n6595 ;
  assign n6591 = n3733 & n6337 ;
  assign n6592 = ~n6587 & ~n6591 ;
  assign n6593 = ~n3177 & ~n6592 ;
  assign n6597 = n3733 & n6351 ;
  assign n6598 = ~n6587 & ~n6597 ;
  assign n6599 = n3411 & ~n6598 ;
  assign n6586 = \P2_reg1_reg[18]/NET0131  & ~n3743 ;
  assign n6600 = n3733 & n6356 ;
  assign n6601 = ~n6586 & ~n6600 ;
  assign n6602 = ~n6599 & n6601 ;
  assign n6603 = ~n6593 & n6602 ;
  assign n6604 = ~n6596 & n6603 ;
  assign n6605 = ~n6590 & n6604 ;
  assign n6606 = n2026 & ~n6605 ;
  assign n6607 = ~n6585 & ~n6606 ;
  assign n6608 = \P1_state_reg[0]/NET0131  & ~n6607 ;
  assign n6609 = ~n6584 & ~n6608 ;
  assign n6610 = \P2_reg1_reg[19]/NET0131  & ~n1983 ;
  assign n6611 = \P2_reg1_reg[19]/NET0131  & n2024 ;
  assign n6613 = \P2_reg1_reg[19]/NET0131  & ~n3733 ;
  assign n6614 = n3733 & n5608 ;
  assign n6615 = ~n6613 & ~n6614 ;
  assign n6616 = ~n3177 & ~n6615 ;
  assign n6620 = n3733 & n5624 ;
  assign n6621 = ~n6613 & ~n6620 ;
  assign n6622 = n3411 & ~n6621 ;
  assign n6623 = n3733 & n5630 ;
  assign n6624 = ~n6613 & ~n6623 ;
  assign n6625 = n3355 & ~n6624 ;
  assign n6617 = n3733 & ~n5614 ;
  assign n6618 = ~n6613 & ~n6617 ;
  assign n6619 = ~n3320 & ~n6618 ;
  assign n6612 = \P2_reg1_reg[19]/NET0131  & ~n3743 ;
  assign n6626 = n2299 & n3358 ;
  assign n6627 = n3733 & n6626 ;
  assign n6628 = ~n6612 & ~n6627 ;
  assign n6629 = ~n6619 & n6628 ;
  assign n6630 = ~n6625 & n6629 ;
  assign n6631 = ~n6622 & n6630 ;
  assign n6632 = ~n6616 & n6631 ;
  assign n6633 = n2026 & ~n6632 ;
  assign n6634 = ~n6611 & ~n6633 ;
  assign n6635 = \P1_state_reg[0]/NET0131  & ~n6634 ;
  assign n6636 = ~n6610 & ~n6635 ;
  assign n6637 = \P2_reg1_reg[21]/NET0131  & ~n1983 ;
  assign n6638 = \P2_reg1_reg[21]/NET0131  & n2024 ;
  assign n6639 = n3320 & ~n3358 ;
  assign n6640 = n3177 & ~n3745 ;
  assign n6641 = n6639 & n6640 ;
  assign n6642 = ~n3733 & ~n6641 ;
  assign n6643 = n3421 & ~n6642 ;
  assign n6644 = \P2_reg1_reg[21]/NET0131  & ~n6643 ;
  assign n6646 = ~n3177 & ~n6290 ;
  assign n6645 = n3121 & n3358 ;
  assign n6647 = n6309 & ~n6645 ;
  assign n6648 = ~n6646 & n6647 ;
  assign n6649 = n3733 & ~n6648 ;
  assign n6650 = ~n6644 & ~n6649 ;
  assign n6651 = n2026 & ~n6650 ;
  assign n6652 = ~n6638 & ~n6651 ;
  assign n6653 = \P1_state_reg[0]/NET0131  & ~n6652 ;
  assign n6654 = ~n6637 & ~n6653 ;
  assign n6655 = \P2_reg1_reg[22]/NET0131  & ~n1983 ;
  assign n6656 = \P2_reg1_reg[22]/NET0131  & n2024 ;
  assign n6659 = \P2_reg1_reg[22]/NET0131  & ~n3733 ;
  assign n6663 = n3733 & n5760 ;
  assign n6664 = ~n6659 & ~n6663 ;
  assign n6665 = ~n3320 & ~n6664 ;
  assign n6660 = n3733 & ~n5753 ;
  assign n6661 = ~n6659 & ~n6660 ;
  assign n6662 = ~n3177 & ~n6661 ;
  assign n6657 = n3733 & ~n6379 ;
  assign n6658 = \P2_reg1_reg[22]/NET0131  & ~n3747 ;
  assign n6666 = ~n6657 & ~n6658 ;
  assign n6667 = ~n6662 & n6666 ;
  assign n6668 = ~n6665 & n6667 ;
  assign n6669 = n2026 & ~n6668 ;
  assign n6670 = ~n6656 & ~n6669 ;
  assign n6671 = \P1_state_reg[0]/NET0131  & ~n6670 ;
  assign n6672 = ~n6655 & ~n6671 ;
  assign n6673 = \P2_reg2_reg[17]/NET0131  & ~n1983 ;
  assign n6674 = \P2_reg2_reg[17]/NET0131  & n2024 ;
  assign n6676 = \P2_reg2_reg[17]/NET0131  & ~n3758 ;
  assign n6677 = n3758 & n5558 ;
  assign n6678 = ~n6676 & ~n6677 ;
  assign n6679 = ~n3177 & ~n6678 ;
  assign n6686 = n3758 & n5586 ;
  assign n6687 = ~n6676 & ~n6686 ;
  assign n6688 = ~n3320 & ~n6687 ;
  assign n6690 = n3758 & n6529 ;
  assign n6675 = \P2_reg2_reg[17]/NET0131  & ~n3774 ;
  assign n6689 = n2373 & n3420 ;
  assign n6691 = ~n6675 & ~n6689 ;
  assign n6692 = ~n6690 & n6691 ;
  assign n6693 = ~n6688 & n6692 ;
  assign n6694 = ~n6679 & n6693 ;
  assign n6680 = n3758 & ~n5570 ;
  assign n6681 = ~n6676 & ~n6680 ;
  assign n6682 = n3411 & ~n6681 ;
  assign n6683 = n3758 & n5578 ;
  assign n6684 = ~n6676 & ~n6683 ;
  assign n6685 = n3355 & ~n6684 ;
  assign n6695 = ~n6682 & ~n6685 ;
  assign n6696 = n6694 & n6695 ;
  assign n6697 = n2026 & ~n6696 ;
  assign n6698 = ~n6674 & ~n6697 ;
  assign n6699 = \P1_state_reg[0]/NET0131  & ~n6698 ;
  assign n6700 = ~n6673 & ~n6699 ;
  assign n6701 = \P2_reg2_reg[19]/NET0131  & ~n1983 ;
  assign n6702 = \P2_reg2_reg[19]/NET0131  & n2024 ;
  assign n6704 = \P2_reg2_reg[19]/NET0131  & ~n3758 ;
  assign n6705 = n3758 & n5608 ;
  assign n6706 = ~n6704 & ~n6705 ;
  assign n6707 = ~n3177 & ~n6706 ;
  assign n6711 = n3758 & n5624 ;
  assign n6712 = ~n6704 & ~n6711 ;
  assign n6713 = n3411 & ~n6712 ;
  assign n6714 = n3758 & n5630 ;
  assign n6715 = ~n6704 & ~n6714 ;
  assign n6716 = n3355 & ~n6715 ;
  assign n6708 = n3758 & ~n5614 ;
  assign n6709 = ~n6704 & ~n6708 ;
  assign n6710 = ~n3320 & ~n6709 ;
  assign n6703 = n3758 & n6626 ;
  assign n6717 = n2307 & n3420 ;
  assign n6718 = \P2_reg2_reg[19]/NET0131  & ~n3774 ;
  assign n6719 = ~n6717 & ~n6718 ;
  assign n6720 = ~n6703 & n6719 ;
  assign n6721 = ~n6710 & n6720 ;
  assign n6722 = ~n6716 & n6721 ;
  assign n6723 = ~n6713 & n6722 ;
  assign n6724 = ~n6707 & n6723 ;
  assign n6725 = n2026 & ~n6724 ;
  assign n6726 = ~n6702 & ~n6725 ;
  assign n6727 = \P1_state_reg[0]/NET0131  & ~n6726 ;
  assign n6728 = ~n6701 & ~n6727 ;
  assign n6729 = \P2_reg2_reg[20]/NET0131  & ~n1983 ;
  assign n6730 = \P2_reg2_reg[20]/NET0131  & n2024 ;
  assign n6732 = \P2_reg2_reg[20]/NET0131  & ~n3758 ;
  assign n6733 = n3130 & ~n5620 ;
  assign n6734 = ~n3394 & ~n6733 ;
  assign n6735 = ~n2058 & ~n6734 ;
  assign n6736 = n2058 & n2311 ;
  assign n6737 = ~n6735 & ~n6736 ;
  assign n6738 = n3758 & n6737 ;
  assign n6739 = ~n6732 & ~n6738 ;
  assign n6740 = n3411 & ~n6739 ;
  assign n6741 = n3916 & n4217 ;
  assign n6742 = ~n3916 & ~n4217 ;
  assign n6743 = ~n6741 & ~n6742 ;
  assign n6744 = n3758 & ~n6743 ;
  assign n6745 = ~n6732 & ~n6744 ;
  assign n6746 = ~n3177 & ~n6745 ;
  assign n6759 = n2358 & n3358 ;
  assign n6760 = n3758 & n6759 ;
  assign n6731 = \P2_reg2_reg[20]/NET0131  & ~n3774 ;
  assign n6758 = n2364 & n3420 ;
  assign n6761 = ~n6731 & ~n6758 ;
  assign n6762 = ~n6760 & n6761 ;
  assign n6763 = ~n6746 & n6762 ;
  assign n6747 = ~n3845 & n4217 ;
  assign n6748 = n3845 & ~n4217 ;
  assign n6749 = ~n6747 & ~n6748 ;
  assign n6750 = n3758 & ~n6749 ;
  assign n6751 = ~n6732 & ~n6750 ;
  assign n6752 = ~n3320 & ~n6751 ;
  assign n6753 = n2358 & ~n5629 ;
  assign n6754 = ~n5765 & ~n6753 ;
  assign n6755 = n3758 & n6754 ;
  assign n6756 = ~n6732 & ~n6755 ;
  assign n6757 = n3355 & ~n6756 ;
  assign n6764 = ~n6752 & ~n6757 ;
  assign n6765 = n6763 & n6764 ;
  assign n6766 = ~n6740 & n6765 ;
  assign n6767 = n2026 & ~n6766 ;
  assign n6768 = ~n6730 & ~n6767 ;
  assign n6769 = \P1_state_reg[0]/NET0131  & ~n6768 ;
  assign n6770 = ~n6729 & ~n6769 ;
  assign n6771 = \P2_reg2_reg[22]/NET0131  & ~n1983 ;
  assign n6772 = \P2_reg2_reg[22]/NET0131  & n2024 ;
  assign n6776 = \P2_reg2_reg[22]/NET0131  & ~n3758 ;
  assign n6780 = n3758 & n5760 ;
  assign n6781 = ~n6776 & ~n6780 ;
  assign n6782 = ~n3320 & ~n6781 ;
  assign n6777 = n3758 & ~n5753 ;
  assign n6778 = ~n6776 & ~n6777 ;
  assign n6779 = ~n3177 & ~n6778 ;
  assign n6773 = n3758 & ~n6379 ;
  assign n6774 = \P2_reg2_reg[22]/NET0131  & ~n4933 ;
  assign n6775 = n3108 & n3420 ;
  assign n6783 = ~n6774 & ~n6775 ;
  assign n6784 = ~n6773 & n6783 ;
  assign n6785 = ~n6779 & n6784 ;
  assign n6786 = ~n6782 & n6785 ;
  assign n6787 = n2026 & ~n6786 ;
  assign n6788 = ~n6772 & ~n6787 ;
  assign n6789 = \P1_state_reg[0]/NET0131  & ~n6788 ;
  assign n6790 = ~n6771 & ~n6789 ;
  assign n6791 = \P1_reg0_reg[17]/NET0131  & ~n3435 ;
  assign n6792 = \P1_reg0_reg[17]/NET0131  & n3448 ;
  assign n6795 = \P1_reg0_reg[17]/NET0131  & ~n4396 ;
  assign n6805 = n4396 & n5462 ;
  assign n6806 = ~n6795 & ~n6805 ;
  assign n6807 = n1936 & ~n6806 ;
  assign n6799 = n4396 & n5445 ;
  assign n6800 = ~n6795 & ~n6799 ;
  assign n6801 = n3712 & ~n6800 ;
  assign n6793 = \P1_reg0_reg[17]/NET0131  & ~n4493 ;
  assign n6794 = n4396 & n6442 ;
  assign n6808 = ~n6793 & ~n6794 ;
  assign n6809 = ~n6801 & n6808 ;
  assign n6810 = ~n6807 & n6809 ;
  assign n6796 = n4396 & n5436 ;
  assign n6797 = ~n6795 & ~n6796 ;
  assign n6798 = ~n3677 & ~n6797 ;
  assign n6802 = n4396 & ~n5453 ;
  assign n6803 = ~n6795 & ~n6802 ;
  assign n6804 = ~n3563 & ~n6803 ;
  assign n6811 = ~n6798 & ~n6804 ;
  assign n6812 = n6810 & n6811 ;
  assign n6813 = n3450 & ~n6812 ;
  assign n6814 = ~n6792 & ~n6813 ;
  assign n6815 = \P1_state_reg[0]/NET0131  & ~n6814 ;
  assign n6816 = ~n6791 & ~n6815 ;
  assign n6817 = \P1_reg0_reg[18]/NET0131  & ~n3435 ;
  assign n6818 = \P1_reg0_reg[18]/NET0131  & n3448 ;
  assign n6820 = \P1_reg0_reg[18]/NET0131  & ~n4396 ;
  assign n6821 = n4396 & n5482 ;
  assign n6822 = ~n6820 & ~n6821 ;
  assign n6823 = n3712 & ~n6822 ;
  assign n6819 = n4396 & n6413 ;
  assign n6833 = \P1_reg0_reg[18]/NET0131  & ~n4493 ;
  assign n6834 = ~n6819 & ~n6833 ;
  assign n6835 = ~n6823 & n6834 ;
  assign n6830 = n4396 & ~n5536 ;
  assign n6831 = ~n6820 & ~n6830 ;
  assign n6832 = n1936 & ~n6831 ;
  assign n6824 = n4396 & ~n5504 ;
  assign n6825 = ~n6820 & ~n6824 ;
  assign n6826 = ~n3677 & ~n6825 ;
  assign n6827 = n4396 & n5527 ;
  assign n6828 = ~n6820 & ~n6827 ;
  assign n6829 = ~n3563 & ~n6828 ;
  assign n6836 = ~n6826 & ~n6829 ;
  assign n6837 = ~n6832 & n6836 ;
  assign n6838 = n6835 & n6837 ;
  assign n6839 = n3450 & ~n6838 ;
  assign n6840 = ~n6818 & ~n6839 ;
  assign n6841 = \P1_state_reg[0]/NET0131  & ~n6840 ;
  assign n6842 = ~n6817 & ~n6841 ;
  assign n6843 = \P1_reg0_reg[19]/NET0131  & ~n3435 ;
  assign n6844 = \P1_reg0_reg[19]/NET0131  & n3448 ;
  assign n6845 = ~n1936 & n3563 ;
  assign n6846 = n3677 & n6845 ;
  assign n6847 = ~n4396 & ~n6846 ;
  assign n6848 = n4494 & ~n6847 ;
  assign n6849 = \P1_reg0_reg[19]/NET0131  & ~n6848 ;
  assign n6850 = n1936 & ~n5654 ;
  assign n6853 = ~n3677 & ~n5667 ;
  assign n6852 = ~n3563 & n5661 ;
  assign n6851 = n1418 & n1880 ;
  assign n6854 = ~n5674 & ~n6851 ;
  assign n6855 = ~n6852 & n6854 ;
  assign n6856 = ~n6853 & n6855 ;
  assign n6857 = ~n6850 & n6856 ;
  assign n6858 = n4396 & ~n6857 ;
  assign n6859 = ~n6849 & ~n6858 ;
  assign n6860 = n3450 & ~n6859 ;
  assign n6861 = ~n6844 & ~n6860 ;
  assign n6862 = \P1_state_reg[0]/NET0131  & ~n6861 ;
  assign n6863 = ~n6843 & ~n6862 ;
  assign n6864 = \P1_reg0_reg[22]/NET0131  & ~n3435 ;
  assign n6865 = \P1_reg0_reg[22]/NET0131  & n3448 ;
  assign n6866 = \P1_reg0_reg[22]/NET0131  & ~n4396 ;
  assign n6870 = n4396 & n6026 ;
  assign n6871 = ~n6866 & ~n6870 ;
  assign n6872 = ~n3677 & ~n6871 ;
  assign n6867 = n4396 & ~n6038 ;
  assign n6868 = ~n6866 & ~n6867 ;
  assign n6869 = ~n3563 & ~n6868 ;
  assign n6874 = n4396 & ~n6048 ;
  assign n6875 = ~n6866 & ~n6874 ;
  assign n6876 = n1936 & ~n6875 ;
  assign n6873 = \P1_reg0_reg[22]/NET0131  & ~n4494 ;
  assign n6877 = n4396 & ~n6057 ;
  assign n6878 = ~n6873 & ~n6877 ;
  assign n6879 = ~n6876 & n6878 ;
  assign n6880 = ~n6869 & n6879 ;
  assign n6881 = ~n6872 & n6880 ;
  assign n6882 = n3450 & ~n6881 ;
  assign n6883 = ~n6865 & ~n6882 ;
  assign n6884 = \P1_state_reg[0]/NET0131  & ~n6883 ;
  assign n6885 = ~n6864 & ~n6884 ;
  assign n6886 = n4396 & n5812 ;
  assign n6887 = n4491 & n6886 ;
  assign n6888 = \P1_reg0_reg[31]/NET0131  & ~n6887 ;
  assign n6889 = ~n5809 & n6886 ;
  assign n6890 = ~n6888 & ~n6889 ;
  assign n6891 = \P1_reg1_reg[17]/NET0131  & ~n3435 ;
  assign n6892 = \P1_reg1_reg[17]/NET0131  & n3448 ;
  assign n6895 = \P1_reg1_reg[17]/NET0131  & ~n4532 ;
  assign n6905 = n4532 & n5462 ;
  assign n6906 = ~n6895 & ~n6905 ;
  assign n6907 = n1936 & ~n6906 ;
  assign n6899 = n4532 & n5445 ;
  assign n6900 = ~n6895 & ~n6899 ;
  assign n6901 = n3712 & ~n6900 ;
  assign n6893 = \P1_reg1_reg[17]/NET0131  & ~n4541 ;
  assign n6894 = n4532 & n6442 ;
  assign n6908 = ~n6893 & ~n6894 ;
  assign n6909 = ~n6901 & n6908 ;
  assign n6910 = ~n6907 & n6909 ;
  assign n6896 = n4532 & n5436 ;
  assign n6897 = ~n6895 & ~n6896 ;
  assign n6898 = ~n3677 & ~n6897 ;
  assign n6902 = n4532 & ~n5453 ;
  assign n6903 = ~n6895 & ~n6902 ;
  assign n6904 = ~n3563 & ~n6903 ;
  assign n6911 = ~n6898 & ~n6904 ;
  assign n6912 = n6910 & n6911 ;
  assign n6913 = n3450 & ~n6912 ;
  assign n6914 = ~n6892 & ~n6913 ;
  assign n6915 = \P1_state_reg[0]/NET0131  & ~n6914 ;
  assign n6916 = ~n6891 & ~n6915 ;
  assign n6917 = \P1_reg1_reg[18]/NET0131  & ~n3435 ;
  assign n6918 = \P1_reg1_reg[18]/NET0131  & n3448 ;
  assign n6920 = \P1_reg1_reg[18]/NET0131  & ~n4532 ;
  assign n6921 = n4532 & n5482 ;
  assign n6922 = ~n6920 & ~n6921 ;
  assign n6923 = n3712 & ~n6922 ;
  assign n6919 = n4532 & n6413 ;
  assign n6933 = \P1_reg1_reg[18]/NET0131  & ~n4541 ;
  assign n6934 = ~n6919 & ~n6933 ;
  assign n6935 = ~n6923 & n6934 ;
  assign n6930 = n4532 & ~n5536 ;
  assign n6931 = ~n6920 & ~n6930 ;
  assign n6932 = n1936 & ~n6931 ;
  assign n6924 = n4532 & ~n5504 ;
  assign n6925 = ~n6920 & ~n6924 ;
  assign n6926 = ~n3677 & ~n6925 ;
  assign n6927 = n4532 & n5527 ;
  assign n6928 = ~n6920 & ~n6927 ;
  assign n6929 = ~n3563 & ~n6928 ;
  assign n6936 = ~n6926 & ~n6929 ;
  assign n6937 = ~n6932 & n6936 ;
  assign n6938 = n6935 & n6937 ;
  assign n6939 = n3450 & ~n6938 ;
  assign n6940 = ~n6918 & ~n6939 ;
  assign n6941 = \P1_state_reg[0]/NET0131  & ~n6940 ;
  assign n6942 = ~n6917 & ~n6941 ;
  assign n6943 = \P1_reg1_reg[19]/NET0131  & ~n3435 ;
  assign n6944 = \P1_reg1_reg[19]/NET0131  & n3448 ;
  assign n6945 = n4491 & n4532 ;
  assign n6946 = \P1_reg1_reg[19]/NET0131  & ~n6945 ;
  assign n6947 = n4532 & ~n6857 ;
  assign n6948 = ~n6946 & ~n6947 ;
  assign n6949 = n3450 & ~n6948 ;
  assign n6950 = ~n6944 & ~n6949 ;
  assign n6951 = \P1_state_reg[0]/NET0131  & ~n6950 ;
  assign n6952 = ~n6943 & ~n6951 ;
  assign n6953 = \P1_reg1_reg[21]/NET0131  & ~n3435 ;
  assign n6954 = \P1_reg1_reg[21]/NET0131  & n3448 ;
  assign n6957 = \P1_reg1_reg[21]/NET0131  & ~n4532 ;
  assign n6958 = n1318 & ~n5795 ;
  assign n6959 = ~n6044 & ~n6958 ;
  assign n6960 = ~n537 & ~n6959 ;
  assign n6961 = n537 & n1374 ;
  assign n6962 = ~n6960 & ~n6961 ;
  assign n6963 = n4532 & n6962 ;
  assign n6964 = ~n6957 & ~n6963 ;
  assign n6965 = n1936 & ~n6964 ;
  assign n6978 = n1346 & ~n3698 ;
  assign n6979 = ~n6052 & ~n6978 ;
  assign n6980 = n4532 & n6979 ;
  assign n6981 = ~n6957 & ~n6980 ;
  assign n6982 = n3712 & ~n6981 ;
  assign n6955 = n1346 & n1880 ;
  assign n6956 = n4532 & n6955 ;
  assign n6983 = \P1_reg1_reg[21]/NET0131  & ~n4541 ;
  assign n6984 = ~n6956 & ~n6983 ;
  assign n6985 = ~n6982 & n6984 ;
  assign n6986 = ~n6965 & n6985 ;
  assign n6966 = n1841 & n3550 ;
  assign n6967 = ~n1841 & ~n3550 ;
  assign n6968 = ~n6966 & ~n6967 ;
  assign n6969 = n4532 & ~n6968 ;
  assign n6970 = ~n6957 & ~n6969 ;
  assign n6971 = ~n3563 & ~n6970 ;
  assign n6972 = n1841 & n3664 ;
  assign n6973 = ~n1841 & ~n3664 ;
  assign n6974 = ~n6972 & ~n6973 ;
  assign n6975 = n4532 & n6974 ;
  assign n6976 = ~n6957 & ~n6975 ;
  assign n6977 = ~n3677 & ~n6976 ;
  assign n6987 = ~n6971 & ~n6977 ;
  assign n6988 = n6986 & n6987 ;
  assign n6989 = n3450 & ~n6988 ;
  assign n6990 = ~n6954 & ~n6989 ;
  assign n6991 = \P1_state_reg[0]/NET0131  & ~n6990 ;
  assign n6992 = ~n6953 & ~n6991 ;
  assign n6993 = \P2_reg0_reg[17]/NET0131  & ~n1983 ;
  assign n6994 = \P2_reg0_reg[17]/NET0131  & n2024 ;
  assign n6996 = \P2_reg0_reg[17]/NET0131  & ~n2040 ;
  assign n6997 = n2040 & n5558 ;
  assign n6998 = ~n6996 & ~n6997 ;
  assign n6999 = ~n3177 & ~n6998 ;
  assign n7006 = n2040 & n5586 ;
  assign n7007 = ~n6996 & ~n7006 ;
  assign n7008 = ~n3320 & ~n7007 ;
  assign n6995 = \P2_reg0_reg[17]/NET0131  & ~n3423 ;
  assign n7009 = n2040 & n6529 ;
  assign n7010 = ~n6995 & ~n7009 ;
  assign n7011 = ~n7008 & n7010 ;
  assign n7012 = ~n6999 & n7011 ;
  assign n7000 = n2040 & ~n5570 ;
  assign n7001 = ~n6996 & ~n7000 ;
  assign n7002 = n3411 & ~n7001 ;
  assign n7003 = n2040 & n5578 ;
  assign n7004 = ~n6996 & ~n7003 ;
  assign n7005 = n3355 & ~n7004 ;
  assign n7013 = ~n7002 & ~n7005 ;
  assign n7014 = n7012 & n7013 ;
  assign n7015 = n2026 & ~n7014 ;
  assign n7016 = ~n6994 & ~n7015 ;
  assign n7017 = \P1_state_reg[0]/NET0131  & ~n7016 ;
  assign n7018 = ~n6993 & ~n7017 ;
  assign n7019 = \P2_reg0_reg[18]/NET0131  & ~n1983 ;
  assign n7020 = \P2_reg0_reg[18]/NET0131  & n2024 ;
  assign n7022 = \P2_reg0_reg[18]/NET0131  & ~n2040 ;
  assign n7023 = n2040 & n6331 ;
  assign n7024 = ~n7022 & ~n7023 ;
  assign n7025 = n3355 & ~n7024 ;
  assign n7029 = n2040 & ~n6343 ;
  assign n7030 = ~n7022 & ~n7029 ;
  assign n7031 = ~n3320 & ~n7030 ;
  assign n7026 = n2040 & n6337 ;
  assign n7027 = ~n7022 & ~n7026 ;
  assign n7028 = ~n3177 & ~n7027 ;
  assign n7032 = n2040 & n6351 ;
  assign n7033 = ~n7022 & ~n7032 ;
  assign n7034 = n3411 & ~n7033 ;
  assign n7021 = n2040 & n6356 ;
  assign n7035 = \P2_reg0_reg[18]/NET0131  & ~n3423 ;
  assign n7036 = ~n7021 & ~n7035 ;
  assign n7037 = ~n7034 & n7036 ;
  assign n7038 = ~n7028 & n7037 ;
  assign n7039 = ~n7031 & n7038 ;
  assign n7040 = ~n7025 & n7039 ;
  assign n7041 = n2026 & ~n7040 ;
  assign n7042 = ~n7020 & ~n7041 ;
  assign n7043 = \P1_state_reg[0]/NET0131  & ~n7042 ;
  assign n7044 = ~n7019 & ~n7043 ;
  assign n7045 = \P2_reg0_reg[19]/NET0131  & ~n1983 ;
  assign n7046 = \P2_reg0_reg[19]/NET0131  & n2024 ;
  assign n7048 = \P2_reg0_reg[19]/NET0131  & ~n2040 ;
  assign n7049 = n2040 & n5608 ;
  assign n7050 = ~n7048 & ~n7049 ;
  assign n7051 = ~n3177 & ~n7050 ;
  assign n7055 = n2040 & n5624 ;
  assign n7056 = ~n7048 & ~n7055 ;
  assign n7057 = n3411 & ~n7056 ;
  assign n7058 = n2040 & n5630 ;
  assign n7059 = ~n7048 & ~n7058 ;
  assign n7060 = n3355 & ~n7059 ;
  assign n7052 = n2040 & ~n5614 ;
  assign n7053 = ~n7048 & ~n7052 ;
  assign n7054 = ~n3320 & ~n7053 ;
  assign n7047 = n2040 & n6626 ;
  assign n7061 = \P2_reg0_reg[19]/NET0131  & ~n3423 ;
  assign n7062 = ~n7047 & ~n7061 ;
  assign n7063 = ~n7054 & n7062 ;
  assign n7064 = ~n7060 & n7063 ;
  assign n7065 = ~n7057 & n7064 ;
  assign n7066 = ~n7051 & n7065 ;
  assign n7067 = n2026 & ~n7066 ;
  assign n7068 = ~n7046 & ~n7067 ;
  assign n7069 = \P1_state_reg[0]/NET0131  & ~n7068 ;
  assign n7070 = ~n7045 & ~n7069 ;
  assign n7073 = n1214 & n3448 ;
  assign n7075 = n1214 & ~n3980 ;
  assign n7076 = n1791 & ~n5491 ;
  assign n7077 = ~n1791 & n5491 ;
  assign n7078 = ~n7076 & ~n7077 ;
  assign n7079 = n3980 & ~n7078 ;
  assign n7080 = ~n7075 & ~n7079 ;
  assign n7081 = ~n3677 & ~n7080 ;
  assign n7096 = n1233 & ~n3687 ;
  assign n7097 = ~n6114 & ~n7096 ;
  assign n7098 = n3980 & n7097 ;
  assign n7099 = ~n7075 & ~n7098 ;
  assign n7100 = n3712 & ~n7099 ;
  assign n7074 = n1233 & ~n4067 ;
  assign n7101 = n1214 & ~n4064 ;
  assign n7102 = ~n7074 & ~n7101 ;
  assign n7103 = ~n7100 & n7102 ;
  assign n7104 = ~n7081 & n7103 ;
  assign n7082 = n1207 & ~n3580 ;
  assign n7083 = ~n4069 & ~n7082 ;
  assign n7084 = ~n537 & ~n7083 ;
  assign n7085 = n537 & n1244 ;
  assign n7086 = ~n7084 & ~n7085 ;
  assign n7087 = n3980 & n7086 ;
  assign n7088 = ~n7075 & ~n7087 ;
  assign n7089 = n1936 & ~n7088 ;
  assign n7090 = n1791 & ~n5514 ;
  assign n7091 = ~n1791 & n5514 ;
  assign n7092 = ~n7090 & ~n7091 ;
  assign n7093 = n3980 & n7092 ;
  assign n7094 = ~n7075 & ~n7093 ;
  assign n7095 = ~n3563 & ~n7094 ;
  assign n7105 = ~n7089 & ~n7095 ;
  assign n7106 = n7104 & n7105 ;
  assign n7107 = n3450 & ~n7106 ;
  assign n7108 = ~n7073 & ~n7107 ;
  assign n7109 = \P1_state_reg[0]/NET0131  & ~n7108 ;
  assign n7071 = \P1_reg3_reg[10]/NET0131  & ~\P1_state_reg[0]/NET0131  ;
  assign n7072 = n1214 & n1953 ;
  assign n7110 = ~n7071 & ~n7072 ;
  assign n7111 = ~n7109 & n7110 ;
  assign n7114 = n1140 & n3448 ;
  assign n7116 = n1140 & ~n3980 ;
  assign n7117 = n1799 & ~n3650 ;
  assign n7118 = ~n1799 & n3650 ;
  assign n7119 = ~n7117 & ~n7118 ;
  assign n7120 = n3980 & ~n7119 ;
  assign n7121 = ~n7116 & ~n7120 ;
  assign n7122 = ~n3677 & ~n7121 ;
  assign n7138 = n1136 & ~n3690 ;
  assign n7139 = ~n5440 & ~n7138 ;
  assign n7140 = n3980 & n7139 ;
  assign n7141 = ~n7116 & ~n7140 ;
  assign n7142 = n3712 & ~n7141 ;
  assign n7115 = n1136 & ~n4067 ;
  assign n7143 = n1140 & ~n4064 ;
  assign n7144 = ~n7115 & ~n7143 ;
  assign n7145 = ~n7142 & n7144 ;
  assign n7146 = ~n7122 & n7145 ;
  assign n7123 = n1799 & ~n3533 ;
  assign n7124 = ~n1799 & n3533 ;
  assign n7125 = ~n7123 & ~n7124 ;
  assign n7126 = n3980 & n7125 ;
  assign n7127 = ~n7116 & ~n7126 ;
  assign n7128 = ~n3563 & ~n7127 ;
  assign n7129 = n1118 & ~n3583 ;
  assign n7130 = ~n1118 & n3583 ;
  assign n7131 = ~n7129 & ~n7130 ;
  assign n7132 = ~n537 & ~n7131 ;
  assign n7133 = n537 & n1174 ;
  assign n7134 = ~n7132 & ~n7133 ;
  assign n7135 = n3980 & n7134 ;
  assign n7136 = ~n7116 & ~n7135 ;
  assign n7137 = n1936 & ~n7136 ;
  assign n7147 = ~n7128 & ~n7137 ;
  assign n7148 = n7146 & n7147 ;
  assign n7149 = n3450 & ~n7148 ;
  assign n7150 = ~n7114 & ~n7149 ;
  assign n7151 = \P1_state_reg[0]/NET0131  & ~n7150 ;
  assign n7112 = n1140 & n1953 ;
  assign n7113 = \P1_reg3_reg[13]/NET0131  & ~\P1_state_reg[0]/NET0131  ;
  assign n7152 = ~n7112 & ~n7113 ;
  assign n7153 = ~n7151 & n7152 ;
  assign n7156 = n2024 & n2735 ;
  assign n7158 = n2735 & ~n3788 ;
  assign n7159 = n2688 & ~n3383 ;
  assign n7160 = ~n6179 & ~n7159 ;
  assign n7161 = ~n2058 & ~n7160 ;
  assign n7162 = n2058 & n2765 ;
  assign n7163 = ~n7161 & ~n7162 ;
  assign n7164 = n3788 & n7163 ;
  assign n7165 = ~n7158 & ~n7164 ;
  assign n7166 = n3411 & ~n7165 ;
  assign n7173 = n4195 & ~n4709 ;
  assign n7174 = ~n4195 & n4709 ;
  assign n7175 = ~n7173 & ~n7174 ;
  assign n7176 = n3788 & n7175 ;
  assign n7177 = ~n7158 & ~n7176 ;
  assign n7178 = ~n3320 & ~n7177 ;
  assign n7167 = n4195 & ~n4740 ;
  assign n7168 = ~n4195 & n4740 ;
  assign n7169 = ~n7167 & ~n7168 ;
  assign n7170 = n3788 & ~n7169 ;
  assign n7171 = ~n7158 & ~n7170 ;
  assign n7172 = ~n3177 & ~n7171 ;
  assign n7179 = ~n2755 & n3334 ;
  assign n7180 = n2755 & ~n3334 ;
  assign n7181 = ~n7179 & ~n7180 ;
  assign n7182 = n3788 & n7181 ;
  assign n7183 = ~n7158 & ~n7182 ;
  assign n7184 = n3355 & ~n7183 ;
  assign n7157 = n2755 & ~n3965 ;
  assign n7185 = n2735 & ~n3962 ;
  assign n7186 = ~n7157 & ~n7185 ;
  assign n7187 = ~n7184 & n7186 ;
  assign n7188 = ~n7172 & n7187 ;
  assign n7189 = ~n7178 & n7188 ;
  assign n7190 = ~n7166 & n7189 ;
  assign n7191 = n2026 & ~n7190 ;
  assign n7192 = ~n7156 & ~n7191 ;
  assign n7193 = \P1_state_reg[0]/NET0131  & ~n7192 ;
  assign n7154 = ~\P1_state_reg[0]/NET0131  & \P2_reg3_reg[10]/NET0131  ;
  assign n7155 = n2735 & n3976 ;
  assign n7194 = ~n7154 & ~n7155 ;
  assign n7195 = ~n7193 & n7194 ;
  assign n7198 = n2024 & n2874 ;
  assign n7200 = n2874 & ~n3788 ;
  assign n7201 = n2058 & ~n2715 ;
  assign n7202 = n2870 & ~n6182 ;
  assign n7203 = ~n2058 & ~n3387 ;
  assign n7204 = ~n7202 & n7203 ;
  assign n7205 = ~n7201 & ~n7204 ;
  assign n7206 = n3788 & ~n7205 ;
  assign n7207 = ~n7200 & ~n7206 ;
  assign n7208 = n3411 & ~n7207 ;
  assign n7209 = ~n2794 & n4192 ;
  assign n7210 = n2794 & ~n4192 ;
  assign n7211 = ~n7209 & ~n7210 ;
  assign n7212 = n3788 & n7211 ;
  assign n7213 = ~n7200 & ~n7212 ;
  assign n7214 = ~n3177 & ~n7213 ;
  assign n7215 = ~n2893 & n3337 ;
  assign n7216 = n2893 & ~n3337 ;
  assign n7217 = ~n7215 & ~n7216 ;
  assign n7218 = n3788 & n7217 ;
  assign n7219 = ~n7200 & ~n7218 ;
  assign n7220 = n3355 & ~n7219 ;
  assign n7221 = ~n3280 & n4192 ;
  assign n7222 = n3280 & ~n4192 ;
  assign n7223 = ~n7221 & ~n7222 ;
  assign n7224 = n3788 & ~n7223 ;
  assign n7225 = ~n7200 & ~n7224 ;
  assign n7226 = ~n3320 & ~n7225 ;
  assign n7199 = n2893 & ~n3965 ;
  assign n7227 = n2874 & ~n3962 ;
  assign n7228 = ~n7199 & ~n7227 ;
  assign n7229 = ~n7226 & n7228 ;
  assign n7230 = ~n7220 & n7229 ;
  assign n7231 = ~n7214 & n7230 ;
  assign n7232 = ~n7208 & n7231 ;
  assign n7233 = n2026 & ~n7232 ;
  assign n7234 = ~n7198 & ~n7233 ;
  assign n7235 = \P1_state_reg[0]/NET0131  & ~n7234 ;
  assign n7196 = n2874 & n3976 ;
  assign n7197 = ~\P1_state_reg[0]/NET0131  & \P2_reg3_reg[13]/NET0131  ;
  assign n7236 = ~n7196 & ~n7197 ;
  assign n7237 = ~n7235 & n7236 ;
  assign n7239 = n2024 & n2760 ;
  assign n7241 = n2760 & ~n3788 ;
  assign n7242 = ~n2454 & n3380 ;
  assign n7243 = ~n2765 & n7242 ;
  assign n7244 = n2742 & ~n7243 ;
  assign n7245 = ~n3383 & ~n7244 ;
  assign n7246 = ~n2058 & ~n7245 ;
  assign n7247 = n2058 & n2454 ;
  assign n7248 = ~n7246 & ~n7247 ;
  assign n7249 = n3788 & n7248 ;
  assign n7250 = ~n7241 & ~n7249 ;
  assign n7251 = n3411 & ~n7250 ;
  assign n7252 = n2678 & ~n4198 ;
  assign n7253 = ~n2678 & n4198 ;
  assign n7254 = ~n7252 & ~n7253 ;
  assign n7255 = n3788 & ~n7254 ;
  assign n7256 = ~n7241 & ~n7255 ;
  assign n7257 = ~n3177 & ~n7256 ;
  assign n7258 = ~n2470 & n3332 ;
  assign n7259 = n2779 & ~n7258 ;
  assign n7260 = ~n3334 & ~n7259 ;
  assign n7261 = n3788 & n7260 ;
  assign n7262 = ~n7241 & ~n7261 ;
  assign n7263 = n3355 & ~n7262 ;
  assign n7264 = n3277 & ~n4198 ;
  assign n7265 = ~n3277 & n4198 ;
  assign n7266 = ~n7264 & ~n7265 ;
  assign n7267 = ~n3320 & n7266 ;
  assign n7268 = n3788 & n7267 ;
  assign n7240 = n2760 & ~n6312 ;
  assign n7269 = n2779 & ~n3965 ;
  assign n7270 = ~n7240 & ~n7269 ;
  assign n7271 = ~n7268 & n7270 ;
  assign n7272 = ~n7263 & n7271 ;
  assign n7273 = ~n7257 & n7272 ;
  assign n7274 = ~n7251 & n7273 ;
  assign n7275 = n2026 & ~n7274 ;
  assign n7276 = ~n7239 & ~n7275 ;
  assign n7277 = \P1_state_reg[0]/NET0131  & ~n7276 ;
  assign n7238 = ~\P1_state_reg[0]/NET0131  & \P2_reg3_reg[9]/NET0131  ;
  assign n7278 = n2760 & n3976 ;
  assign n7279 = ~n7238 & ~n7278 ;
  assign n7280 = ~n7277 & n7279 ;
  assign n7283 = n1239 & n3448 ;
  assign n7285 = n1239 & ~n3980 ;
  assign n7304 = n537 & ~n1267 ;
  assign n7305 = ~n1267 & n3577 ;
  assign n7306 = ~n1244 & n7305 ;
  assign n7307 = n1218 & ~n7306 ;
  assign n7308 = ~n537 & ~n3580 ;
  assign n7309 = ~n7307 & n7308 ;
  assign n7310 = ~n7304 & ~n7309 ;
  assign n7311 = n3980 & ~n7310 ;
  assign n7312 = ~n7285 & ~n7311 ;
  assign n7313 = n1936 & ~n7312 ;
  assign n7292 = n1782 & ~n3529 ;
  assign n7293 = ~n1782 & n3529 ;
  assign n7294 = ~n7292 & ~n7293 ;
  assign n7295 = n3980 & n7294 ;
  assign n7296 = ~n7285 & ~n7295 ;
  assign n7297 = ~n3563 & ~n7296 ;
  assign n7286 = n1782 & ~n3646 ;
  assign n7287 = ~n1782 & n3646 ;
  assign n7288 = ~n7286 & ~n7287 ;
  assign n7289 = n3980 & ~n7288 ;
  assign n7290 = ~n7285 & ~n7289 ;
  assign n7291 = ~n3677 & ~n7290 ;
  assign n7298 = n3684 & n3685 ;
  assign n7299 = n1257 & ~n7298 ;
  assign n7300 = ~n3687 & ~n7299 ;
  assign n7301 = n3980 & n7300 ;
  assign n7302 = ~n7285 & ~n7301 ;
  assign n7303 = n3712 & ~n7302 ;
  assign n7284 = n1257 & ~n4067 ;
  assign n7314 = n1239 & ~n4064 ;
  assign n7315 = ~n7284 & ~n7314 ;
  assign n7316 = ~n7303 & n7315 ;
  assign n7317 = ~n7291 & n7316 ;
  assign n7318 = ~n7297 & n7317 ;
  assign n7319 = ~n7313 & n7318 ;
  assign n7320 = n3450 & ~n7319 ;
  assign n7321 = ~n7283 & ~n7320 ;
  assign n7322 = \P1_state_reg[0]/NET0131  & ~n7321 ;
  assign n7281 = \P1_reg3_reg[9]/NET0131  & ~\P1_state_reg[0]/NET0131  ;
  assign n7282 = n1239 & n1953 ;
  assign n7323 = ~n7281 & ~n7282 ;
  assign n7324 = ~n7322 & n7323 ;
  assign n7327 = n2024 & n2364 ;
  assign n7329 = n2364 & ~n3788 ;
  assign n7330 = n3788 & n6737 ;
  assign n7331 = ~n7329 & ~n7330 ;
  assign n7332 = n3411 & ~n7331 ;
  assign n7333 = n3788 & ~n6743 ;
  assign n7334 = ~n7329 & ~n7333 ;
  assign n7335 = ~n3177 & ~n7334 ;
  assign n7328 = n2364 & ~n3962 ;
  assign n7342 = n2358 & ~n3965 ;
  assign n7343 = ~n7328 & ~n7342 ;
  assign n7344 = ~n7335 & n7343 ;
  assign n7336 = n3788 & ~n6749 ;
  assign n7337 = ~n7329 & ~n7336 ;
  assign n7338 = ~n3320 & ~n7337 ;
  assign n7339 = n3788 & n6754 ;
  assign n7340 = ~n7329 & ~n7339 ;
  assign n7341 = n3355 & ~n7340 ;
  assign n7345 = ~n7338 & ~n7341 ;
  assign n7346 = n7344 & n7345 ;
  assign n7347 = ~n7332 & n7346 ;
  assign n7348 = n2026 & ~n7347 ;
  assign n7349 = ~n7327 & ~n7348 ;
  assign n7350 = \P1_state_reg[0]/NET0131  & ~n7349 ;
  assign n7325 = n2364 & n3976 ;
  assign n7326 = ~\P1_state_reg[0]/NET0131  & \P2_reg3_reg[20]/NET0131  ;
  assign n7351 = ~n7325 & ~n7326 ;
  assign n7352 = ~n7350 & n7351 ;
  assign n7355 = n1370 & n3448 ;
  assign n7356 = n1370 & ~n3980 ;
  assign n7357 = n3980 & n6492 ;
  assign n7358 = ~n7356 & ~n7357 ;
  assign n7359 = n1936 & ~n7358 ;
  assign n7364 = n3980 & ~n6499 ;
  assign n7365 = ~n7356 & ~n7364 ;
  assign n7366 = ~n3677 & ~n7365 ;
  assign n7361 = n3980 & ~n6505 ;
  assign n7362 = ~n7356 & ~n7361 ;
  assign n7363 = ~n3563 & ~n7362 ;
  assign n7367 = n3980 & n6510 ;
  assign n7368 = ~n7356 & ~n7367 ;
  assign n7369 = n3712 & ~n7368 ;
  assign n7360 = n1365 & ~n4067 ;
  assign n7370 = n1370 & ~n4064 ;
  assign n7371 = ~n7360 & ~n7370 ;
  assign n7372 = ~n7369 & n7371 ;
  assign n7373 = ~n7363 & n7372 ;
  assign n7374 = ~n7366 & n7373 ;
  assign n7375 = ~n7359 & n7374 ;
  assign n7376 = n3450 & ~n7375 ;
  assign n7377 = ~n7355 & ~n7376 ;
  assign n7378 = \P1_state_reg[0]/NET0131  & ~n7377 ;
  assign n7353 = \P1_reg3_reg[20]/NET0131  & ~\P1_state_reg[0]/NET0131  ;
  assign n7354 = n1370 & n1953 ;
  assign n7379 = ~n7353 & ~n7354 ;
  assign n7380 = ~n7378 & n7379 ;
  assign n7383 = n1352 & n3448 ;
  assign n7385 = n1352 & ~n3980 ;
  assign n7386 = n3980 & n6962 ;
  assign n7387 = ~n7385 & ~n7386 ;
  assign n7388 = n1936 & ~n7387 ;
  assign n7395 = n3980 & n6979 ;
  assign n7396 = ~n7385 & ~n7395 ;
  assign n7397 = n3712 & ~n7396 ;
  assign n7384 = n1346 & ~n4067 ;
  assign n7398 = n1352 & ~n4064 ;
  assign n7399 = ~n7384 & ~n7398 ;
  assign n7400 = ~n7397 & n7399 ;
  assign n7401 = ~n7388 & n7400 ;
  assign n7389 = n3980 & ~n6968 ;
  assign n7390 = ~n7385 & ~n7389 ;
  assign n7391 = ~n3563 & ~n7390 ;
  assign n7392 = n3980 & n6974 ;
  assign n7393 = ~n7385 & ~n7392 ;
  assign n7394 = ~n3677 & ~n7393 ;
  assign n7402 = ~n7391 & ~n7394 ;
  assign n7403 = n7401 & n7402 ;
  assign n7404 = n3450 & ~n7403 ;
  assign n7405 = ~n7383 & ~n7404 ;
  assign n7406 = \P1_state_reg[0]/NET0131  & ~n7405 ;
  assign n7381 = n1352 & n1953 ;
  assign n7382 = \P1_reg3_reg[21]/NET0131  & ~\P1_state_reg[0]/NET0131  ;
  assign n7407 = ~n7381 & ~n7382 ;
  assign n7408 = ~n7406 & n7407 ;
  assign n7411 = n1330 & n3448 ;
  assign n7412 = n1330 & ~n3980 ;
  assign n7426 = ~n4447 & n4448 ;
  assign n7427 = n4453 & ~n7426 ;
  assign n7428 = n4449 & n4459 ;
  assign n7429 = ~n7427 & n7428 ;
  assign n7430 = ~n4456 & n4459 ;
  assign n7431 = n4435 & ~n7430 ;
  assign n7432 = ~n7429 & n7431 ;
  assign n7433 = n1821 & n7432 ;
  assign n7434 = ~n1821 & ~n7432 ;
  assign n7435 = ~n7433 & ~n7434 ;
  assign n7436 = n3980 & ~n7435 ;
  assign n7437 = ~n7412 & ~n7436 ;
  assign n7438 = ~n3563 & ~n7437 ;
  assign n7413 = ~n4404 & n4406 ;
  assign n7414 = n4410 & ~n7413 ;
  assign n7415 = n4405 & n4417 ;
  assign n7416 = ~n7414 & n7415 ;
  assign n7417 = ~n4413 & n4417 ;
  assign n7418 = n4422 & ~n7417 ;
  assign n7419 = ~n7416 & n7418 ;
  assign n7420 = n1821 & ~n7419 ;
  assign n7421 = ~n1821 & n7419 ;
  assign n7422 = ~n7420 & ~n7421 ;
  assign n7423 = n3980 & ~n7422 ;
  assign n7424 = ~n7412 & ~n7423 ;
  assign n7425 = ~n3677 & ~n7424 ;
  assign n7440 = n1062 & ~n4472 ;
  assign n7441 = ~n4075 & ~n7440 ;
  assign n7442 = ~n537 & ~n7441 ;
  assign n7443 = n537 & n1318 ;
  assign n7444 = ~n7442 & ~n7443 ;
  assign n7445 = n3980 & n7444 ;
  assign n7446 = ~n7412 & ~n7445 ;
  assign n7447 = n1936 & ~n7446 ;
  assign n7448 = n1327 & ~n3700 ;
  assign n7449 = ~n5188 & ~n7448 ;
  assign n7450 = n3712 & n7449 ;
  assign n7451 = n3980 & n7450 ;
  assign n7439 = n1330 & ~n4910 ;
  assign n7452 = n1327 & ~n4067 ;
  assign n7453 = ~n7439 & ~n7452 ;
  assign n7454 = ~n7451 & n7453 ;
  assign n7455 = ~n7447 & n7454 ;
  assign n7456 = ~n7425 & n7455 ;
  assign n7457 = ~n7438 & n7456 ;
  assign n7458 = n3450 & ~n7457 ;
  assign n7459 = ~n7411 & ~n7458 ;
  assign n7460 = \P1_state_reg[0]/NET0131  & ~n7459 ;
  assign n7409 = \P1_reg3_reg[23]/NET0131  & ~\P1_state_reg[0]/NET0131  ;
  assign n7410 = n1330 & n1953 ;
  assign n7461 = ~n7409 & ~n7410 ;
  assign n7462 = ~n7460 & n7461 ;
  assign n7463 = \P2_reg0_reg[20]/NET0131  & ~n1983 ;
  assign n7464 = \P2_reg0_reg[20]/NET0131  & n2024 ;
  assign n7466 = \P2_reg0_reg[20]/NET0131  & ~n2040 ;
  assign n7467 = n2040 & n6737 ;
  assign n7468 = ~n7466 & ~n7467 ;
  assign n7469 = n3411 & ~n7468 ;
  assign n7470 = n2040 & ~n6743 ;
  assign n7471 = ~n7466 & ~n7470 ;
  assign n7472 = ~n3177 & ~n7471 ;
  assign n7465 = \P2_reg0_reg[20]/NET0131  & ~n3423 ;
  assign n7479 = n2040 & n6759 ;
  assign n7480 = ~n7465 & ~n7479 ;
  assign n7481 = ~n7472 & n7480 ;
  assign n7473 = n2040 & ~n6749 ;
  assign n7474 = ~n7466 & ~n7473 ;
  assign n7475 = ~n3320 & ~n7474 ;
  assign n7476 = n2040 & n6754 ;
  assign n7477 = ~n7466 & ~n7476 ;
  assign n7478 = n3355 & ~n7477 ;
  assign n7482 = ~n7475 & ~n7478 ;
  assign n7483 = n7481 & n7482 ;
  assign n7484 = ~n7469 & n7483 ;
  assign n7485 = n2026 & ~n7484 ;
  assign n7486 = ~n7464 & ~n7485 ;
  assign n7487 = \P1_state_reg[0]/NET0131  & ~n7486 ;
  assign n7488 = ~n7463 & ~n7487 ;
  assign n7489 = n825 & n1880 ;
  assign n7490 = ~n5802 & ~n7489 ;
  assign n7491 = n825 & ~n3708 ;
  assign n7492 = ~n5803 & ~n7491 ;
  assign n7493 = n3712 & n7492 ;
  assign n7494 = n7490 & ~n7493 ;
  assign n7495 = n4532 & ~n7494 ;
  assign n7496 = \P1_reg1_reg[30]/NET0131  & ~n6945 ;
  assign n7497 = ~n7495 & ~n7496 ;
  assign n7498 = n3450 & ~n7497 ;
  assign n7499 = \P1_reg1_reg[30]/NET0131  & n3448 ;
  assign n7500 = ~n7498 & ~n7499 ;
  assign n7501 = \P1_state_reg[0]/NET0131  & ~n7500 ;
  assign n7502 = \P1_reg1_reg[30]/NET0131  & ~n3435 ;
  assign n7503 = ~n7501 & ~n7502 ;
  assign n7504 = n5860 & ~n6648 ;
  assign n7508 = ~n3171 & n4308 ;
  assign n7509 = ~n2040 & ~n7508 ;
  assign n7510 = n5287 & ~n7509 ;
  assign n7505 = ~n2040 & ~n6639 ;
  assign n7506 = n3421 & ~n7505 ;
  assign n7507 = ~n2040 & n3354 ;
  assign n7511 = n7506 & ~n7507 ;
  assign n7512 = n7510 & n7511 ;
  assign n7513 = \P2_reg0_reg[21]/NET0131  & ~n7512 ;
  assign n7514 = ~n7504 & ~n7513 ;
  assign n7515 = \P1_reg2_reg[12]/NET0131  & ~n3435 ;
  assign n7516 = \P1_reg2_reg[12]/NET0131  & n3448 ;
  assign n7518 = \P1_reg2_reg[12]/NET0131  & ~n3466 ;
  assign n7519 = n3466 & n6098 ;
  assign n7520 = ~n7518 & ~n7519 ;
  assign n7521 = n1936 & ~n7520 ;
  assign n7525 = n3466 & ~n6110 ;
  assign n7526 = ~n7518 & ~n7525 ;
  assign n7527 = ~n3677 & ~n7526 ;
  assign n7522 = n3466 & n6104 ;
  assign n7523 = ~n7518 & ~n7522 ;
  assign n7524 = ~n3563 & ~n7523 ;
  assign n7528 = n3466 & n6117 ;
  assign n7529 = ~n7518 & ~n7528 ;
  assign n7530 = n3712 & ~n7529 ;
  assign n7517 = \P1_reg2_reg[12]/NET0131  & ~n3718 ;
  assign n7531 = n1170 & n1763 ;
  assign n7532 = n1165 & n1880 ;
  assign n7533 = n3466 & n7532 ;
  assign n7534 = ~n7531 & ~n7533 ;
  assign n7535 = ~n7517 & n7534 ;
  assign n7536 = ~n7530 & n7535 ;
  assign n7537 = ~n7524 & n7536 ;
  assign n7538 = ~n7527 & n7537 ;
  assign n7539 = ~n7521 & n7538 ;
  assign n7540 = n3450 & ~n7539 ;
  assign n7541 = ~n7516 & ~n7540 ;
  assign n7542 = \P1_state_reg[0]/NET0131  & ~n7541 ;
  assign n7543 = ~n7515 & ~n7542 ;
  assign n7544 = \P2_reg0_reg[30]/NET0131  & ~n5861 ;
  assign n7545 = n3358 & n4159 ;
  assign n7546 = ~n5277 & ~n7545 ;
  assign n7547 = ~n3350 & n4159 ;
  assign n7548 = ~n5279 & ~n7547 ;
  assign n7549 = n3355 & n7548 ;
  assign n7550 = n7546 & ~n7549 ;
  assign n7551 = n5860 & ~n7550 ;
  assign n7552 = ~n7544 & ~n7551 ;
  assign n7553 = \P1_reg2_reg[16]/NET0131  & ~n3435 ;
  assign n7554 = \P1_reg2_reg[16]/NET0131  & n3448 ;
  assign n7556 = \P1_reg2_reg[16]/NET0131  & ~n3466 ;
  assign n7560 = n3466 & n6149 ;
  assign n7561 = ~n7556 & ~n7560 ;
  assign n7562 = n1936 & ~n7561 ;
  assign n7557 = n3466 & ~n6141 ;
  assign n7558 = ~n7556 & ~n7557 ;
  assign n7559 = ~n3563 & ~n7558 ;
  assign n7566 = n3466 & ~n6155 ;
  assign n7567 = ~n7556 & ~n7566 ;
  assign n7568 = ~n3677 & ~n7567 ;
  assign n7563 = n3466 & n6160 ;
  assign n7564 = ~n7556 & ~n7563 ;
  assign n7565 = n3712 & ~n7564 ;
  assign n7570 = n1466 & n1880 ;
  assign n7571 = n3466 & n7570 ;
  assign n7555 = \P1_reg2_reg[16]/NET0131  & ~n3718 ;
  assign n7569 = n1471 & n1763 ;
  assign n7572 = ~n7555 & ~n7569 ;
  assign n7573 = ~n7571 & n7572 ;
  assign n7574 = ~n7565 & n7573 ;
  assign n7575 = ~n7568 & n7574 ;
  assign n7576 = ~n7559 & n7575 ;
  assign n7577 = ~n7562 & n7576 ;
  assign n7578 = n3450 & ~n7577 ;
  assign n7579 = ~n7554 & ~n7578 ;
  assign n7580 = \P1_state_reg[0]/NET0131  & ~n7579 ;
  assign n7581 = ~n7553 & ~n7580 ;
  assign n7582 = \P2_reg1_reg[12]/NET0131  & ~n1983 ;
  assign n7583 = \P2_reg1_reg[12]/NET0131  & n2024 ;
  assign n7587 = \P2_reg1_reg[12]/NET0131  & ~n3733 ;
  assign n7588 = n3733 & n6186 ;
  assign n7589 = ~n7587 & ~n7588 ;
  assign n7590 = n3411 & ~n7589 ;
  assign n7594 = n3733 & ~n6198 ;
  assign n7595 = ~n7587 & ~n7594 ;
  assign n7596 = ~n3320 & ~n7595 ;
  assign n7591 = n3733 & n6192 ;
  assign n7592 = ~n7587 & ~n7591 ;
  assign n7593 = ~n3177 & ~n7592 ;
  assign n7584 = n2731 & n3358 ;
  assign n7585 = ~n6204 & ~n7584 ;
  assign n7586 = n3733 & ~n7585 ;
  assign n7597 = n3355 & ~n3733 ;
  assign n7598 = n3743 & ~n7597 ;
  assign n7599 = \P2_reg1_reg[12]/NET0131  & ~n7598 ;
  assign n7600 = ~n7586 & ~n7599 ;
  assign n7601 = ~n7593 & n7600 ;
  assign n7602 = ~n7596 & n7601 ;
  assign n7603 = ~n7590 & n7602 ;
  assign n7604 = n2026 & ~n7603 ;
  assign n7605 = ~n7583 & ~n7604 ;
  assign n7606 = \P1_state_reg[0]/NET0131  & ~n7605 ;
  assign n7607 = ~n7582 & ~n7606 ;
  assign n7608 = \P1_reg2_reg[21]/NET0131  & ~n3435 ;
  assign n7609 = \P1_reg2_reg[21]/NET0131  & n3448 ;
  assign n7611 = \P1_reg2_reg[21]/NET0131  & ~n3466 ;
  assign n7612 = n3466 & n6962 ;
  assign n7613 = ~n7611 & ~n7612 ;
  assign n7614 = n1936 & ~n7613 ;
  assign n7621 = n3466 & n6979 ;
  assign n7622 = ~n7611 & ~n7621 ;
  assign n7623 = n3712 & ~n7622 ;
  assign n7625 = n3466 & n6955 ;
  assign n7610 = \P1_reg2_reg[21]/NET0131  & ~n3718 ;
  assign n7624 = n1352 & n1763 ;
  assign n7626 = ~n7610 & ~n7624 ;
  assign n7627 = ~n7625 & n7626 ;
  assign n7628 = ~n7623 & n7627 ;
  assign n7629 = ~n7614 & n7628 ;
  assign n7615 = n3466 & ~n6968 ;
  assign n7616 = ~n7611 & ~n7615 ;
  assign n7617 = ~n3563 & ~n7616 ;
  assign n7618 = n3466 & n6974 ;
  assign n7619 = ~n7611 & ~n7618 ;
  assign n7620 = ~n3677 & ~n7619 ;
  assign n7630 = ~n7617 & ~n7620 ;
  assign n7631 = n7629 & n7630 ;
  assign n7632 = n3450 & ~n7631 ;
  assign n7633 = ~n7609 & ~n7632 ;
  assign n7634 = \P1_state_reg[0]/NET0131  & ~n7633 ;
  assign n7635 = ~n7608 & ~n7634 ;
  assign n7636 = \P1_reg2_reg[23]/NET0131  & ~n3435 ;
  assign n7637 = \P1_reg2_reg[23]/NET0131  & n3448 ;
  assign n7638 = \P1_reg2_reg[23]/NET0131  & ~n3466 ;
  assign n7642 = n3466 & ~n7435 ;
  assign n7643 = ~n7638 & ~n7642 ;
  assign n7644 = ~n3563 & ~n7643 ;
  assign n7639 = n3466 & ~n7422 ;
  assign n7640 = ~n7638 & ~n7639 ;
  assign n7641 = ~n3677 & ~n7640 ;
  assign n7646 = n3466 & n7444 ;
  assign n7647 = ~n7638 & ~n7646 ;
  assign n7648 = n1936 & ~n7647 ;
  assign n7649 = n3466 & n7449 ;
  assign n7650 = ~n7638 & ~n7649 ;
  assign n7651 = n3712 & ~n7650 ;
  assign n7653 = n1327 & n1880 ;
  assign n7654 = n3466 & n7653 ;
  assign n7645 = \P1_reg2_reg[23]/NET0131  & ~n3718 ;
  assign n7652 = n1330 & n1763 ;
  assign n7655 = ~n7645 & ~n7652 ;
  assign n7656 = ~n7654 & n7655 ;
  assign n7657 = ~n7651 & n7656 ;
  assign n7658 = ~n7648 & n7657 ;
  assign n7659 = ~n7641 & n7658 ;
  assign n7660 = ~n7644 & n7659 ;
  assign n7661 = n3450 & ~n7660 ;
  assign n7662 = ~n7637 & ~n7661 ;
  assign n7663 = \P1_state_reg[0]/NET0131  & ~n7662 ;
  assign n7664 = ~n7636 & ~n7663 ;
  assign n7665 = \P2_reg1_reg[20]/NET0131  & ~n1983 ;
  assign n7666 = \P2_reg1_reg[20]/NET0131  & n2024 ;
  assign n7668 = \P2_reg1_reg[20]/NET0131  & ~n3733 ;
  assign n7669 = n3733 & n6737 ;
  assign n7670 = ~n7668 & ~n7669 ;
  assign n7671 = n3411 & ~n7670 ;
  assign n7672 = n3733 & ~n6743 ;
  assign n7673 = ~n7668 & ~n7672 ;
  assign n7674 = ~n3177 & ~n7673 ;
  assign n7667 = \P2_reg1_reg[20]/NET0131  & ~n3743 ;
  assign n7681 = n3733 & n6759 ;
  assign n7682 = ~n7667 & ~n7681 ;
  assign n7683 = ~n7674 & n7682 ;
  assign n7675 = n3733 & ~n6749 ;
  assign n7676 = ~n7668 & ~n7675 ;
  assign n7677 = ~n3320 & ~n7676 ;
  assign n7678 = n3733 & n6754 ;
  assign n7679 = ~n7668 & ~n7678 ;
  assign n7680 = n3355 & ~n7679 ;
  assign n7684 = ~n7677 & ~n7680 ;
  assign n7685 = n7683 & n7684 ;
  assign n7686 = ~n7671 & n7685 ;
  assign n7687 = n2026 & ~n7686 ;
  assign n7688 = ~n7666 & ~n7687 ;
  assign n7689 = \P1_state_reg[0]/NET0131  & ~n7688 ;
  assign n7690 = ~n7665 & ~n7689 ;
  assign n7691 = \P2_reg1_reg[30]/NET0131  & ~n5962 ;
  assign n7692 = n5964 & ~n7550 ;
  assign n7693 = ~n7691 & ~n7692 ;
  assign n7694 = \P1_reg2_reg[30]/NET0131  & ~n3466 ;
  assign n7695 = n3466 & n5812 ;
  assign n7696 = n7492 & n7695 ;
  assign n7697 = ~n7694 & ~n7696 ;
  assign n7698 = n3712 & ~n7697 ;
  assign n7699 = n3466 & ~n7490 ;
  assign n7700 = ~n3720 & ~n7699 ;
  assign n7701 = n5812 & ~n7700 ;
  assign n7702 = ~n501 & n1762 ;
  assign n7703 = ~n3466 & ~n7702 ;
  assign n7704 = n5815 & ~n7703 ;
  assign n7705 = \P1_reg2_reg[30]/NET0131  & ~n7704 ;
  assign n7706 = ~n7701 & ~n7705 ;
  assign n7707 = ~n7698 & n7706 ;
  assign n7708 = \P2_reg2_reg[12]/NET0131  & ~n1983 ;
  assign n7709 = \P2_reg2_reg[12]/NET0131  & n2024 ;
  assign n7711 = \P2_reg2_reg[12]/NET0131  & ~n3758 ;
  assign n7712 = n3758 & n6186 ;
  assign n7713 = ~n7711 & ~n7712 ;
  assign n7714 = n3411 & ~n7713 ;
  assign n7718 = n3758 & ~n6198 ;
  assign n7719 = ~n7711 & ~n7718 ;
  assign n7720 = ~n3320 & ~n7719 ;
  assign n7715 = n3758 & n6192 ;
  assign n7716 = ~n7711 & ~n7715 ;
  assign n7717 = ~n3177 & ~n7716 ;
  assign n7721 = n3758 & n6203 ;
  assign n7722 = ~n7711 & ~n7721 ;
  assign n7723 = n3355 & ~n7722 ;
  assign n7725 = n3758 & n7584 ;
  assign n7710 = \P2_reg2_reg[12]/NET0131  & ~n3774 ;
  assign n7724 = n2709 & n3420 ;
  assign n7726 = ~n7710 & ~n7724 ;
  assign n7727 = ~n7725 & n7726 ;
  assign n7728 = ~n7723 & n7727 ;
  assign n7729 = ~n7717 & n7728 ;
  assign n7730 = ~n7720 & n7729 ;
  assign n7731 = ~n7714 & n7730 ;
  assign n7732 = n2026 & ~n7731 ;
  assign n7733 = ~n7709 & ~n7732 ;
  assign n7734 = \P1_state_reg[0]/NET0131  & ~n7733 ;
  assign n7735 = ~n7708 & ~n7734 ;
  assign n7736 = \P2_reg2_reg[16]/NET0131  & ~n1983 ;
  assign n7737 = \P2_reg2_reg[16]/NET0131  & n2024 ;
  assign n7739 = \P2_reg2_reg[16]/NET0131  & ~n3758 ;
  assign n7749 = n3758 & ~n6246 ;
  assign n7750 = ~n7739 & ~n7749 ;
  assign n7751 = ~n3320 & ~n7750 ;
  assign n7746 = n3758 & n6240 ;
  assign n7747 = ~n7739 & ~n7746 ;
  assign n7748 = n3355 & ~n7747 ;
  assign n7752 = n2818 & n3358 ;
  assign n7753 = n3758 & n7752 ;
  assign n7738 = \P2_reg2_reg[16]/NET0131  & ~n3774 ;
  assign n7754 = n2797 & n3420 ;
  assign n7755 = ~n7738 & ~n7754 ;
  assign n7756 = ~n7753 & n7755 ;
  assign n7757 = ~n7748 & n7756 ;
  assign n7758 = ~n7751 & n7757 ;
  assign n7740 = n3758 & ~n6226 ;
  assign n7741 = ~n7739 & ~n7740 ;
  assign n7742 = ~n3177 & ~n7741 ;
  assign n7743 = n3758 & n6234 ;
  assign n7744 = ~n7739 & ~n7743 ;
  assign n7745 = n3411 & ~n7744 ;
  assign n7759 = ~n7742 & ~n7745 ;
  assign n7760 = n7758 & n7759 ;
  assign n7761 = n2026 & ~n7760 ;
  assign n7762 = ~n7737 & ~n7761 ;
  assign n7763 = \P1_state_reg[0]/NET0131  & ~n7762 ;
  assign n7764 = ~n7736 & ~n7763 ;
  assign n7765 = n3758 & ~n6648 ;
  assign n7766 = n3126 & n3419 ;
  assign n7767 = ~n7765 & ~n7766 ;
  assign n7768 = n5287 & ~n7767 ;
  assign n7769 = ~n3320 & ~n3758 ;
  assign n7770 = n3774 & ~n7769 ;
  assign n7771 = ~n3758 & ~n6640 ;
  assign n7772 = n5287 & ~n7771 ;
  assign n7773 = n7770 & n7772 ;
  assign n7774 = \P2_reg2_reg[21]/NET0131  & ~n7773 ;
  assign n7775 = ~n7768 & ~n7774 ;
  assign n7776 = \P2_reg2_reg[30]/NET0131  & ~n1983 ;
  assign n7777 = \P2_reg2_reg[30]/NET0131  & n2024 ;
  assign n7779 = n3758 & ~n7548 ;
  assign n7780 = ~\P2_reg2_reg[30]/NET0131  & ~n3758 ;
  assign n7781 = n3355 & ~n7780 ;
  assign n7782 = ~n7779 & n7781 ;
  assign n7783 = n3758 & ~n7546 ;
  assign n7778 = \P2_reg2_reg[30]/NET0131  & ~n5290 ;
  assign n7784 = ~n3776 & ~n7778 ;
  assign n7785 = ~n7783 & n7784 ;
  assign n7786 = ~n7782 & n7785 ;
  assign n7787 = n2026 & ~n7786 ;
  assign n7788 = ~n7777 & ~n7787 ;
  assign n7789 = \P1_state_reg[0]/NET0131  & ~n7788 ;
  assign n7790 = ~n7776 & ~n7789 ;
  assign n7791 = \P1_reg0_reg[12]/NET0131  & ~n3435 ;
  assign n7792 = \P1_reg0_reg[12]/NET0131  & n3448 ;
  assign n7794 = \P1_reg0_reg[12]/NET0131  & ~n4396 ;
  assign n7795 = n4396 & n6098 ;
  assign n7796 = ~n7794 & ~n7795 ;
  assign n7797 = n1936 & ~n7796 ;
  assign n7801 = n4396 & ~n6110 ;
  assign n7802 = ~n7794 & ~n7801 ;
  assign n7803 = ~n3677 & ~n7802 ;
  assign n7798 = n4396 & n6104 ;
  assign n7799 = ~n7794 & ~n7798 ;
  assign n7800 = ~n3563 & ~n7799 ;
  assign n7804 = n4396 & n6117 ;
  assign n7805 = ~n7794 & ~n7804 ;
  assign n7806 = n3712 & ~n7805 ;
  assign n7793 = n4396 & n7532 ;
  assign n7807 = \P1_reg0_reg[12]/NET0131  & ~n4493 ;
  assign n7808 = ~n7793 & ~n7807 ;
  assign n7809 = ~n7806 & n7808 ;
  assign n7810 = ~n7800 & n7809 ;
  assign n7811 = ~n7803 & n7810 ;
  assign n7812 = ~n7797 & n7811 ;
  assign n7813 = n3450 & ~n7812 ;
  assign n7814 = ~n7792 & ~n7813 ;
  assign n7815 = \P1_state_reg[0]/NET0131  & ~n7814 ;
  assign n7816 = ~n7791 & ~n7815 ;
  assign n7817 = \P1_reg0_reg[16]/NET0131  & ~n3435 ;
  assign n7818 = \P1_reg0_reg[16]/NET0131  & n3448 ;
  assign n7819 = \P1_reg0_reg[16]/NET0131  & ~n6848 ;
  assign n7822 = ~n3563 & ~n6141 ;
  assign n7820 = n1936 & n6149 ;
  assign n7821 = ~n3677 & ~n6155 ;
  assign n7823 = ~n6161 & ~n7570 ;
  assign n7824 = ~n7821 & n7823 ;
  assign n7825 = ~n7820 & n7824 ;
  assign n7826 = ~n7822 & n7825 ;
  assign n7827 = n4396 & ~n7826 ;
  assign n7828 = ~n7819 & ~n7827 ;
  assign n7829 = n3450 & ~n7828 ;
  assign n7830 = ~n7818 & ~n7829 ;
  assign n7831 = \P1_state_reg[0]/NET0131  & ~n7830 ;
  assign n7832 = ~n7817 & ~n7831 ;
  assign n7833 = \P1_reg0_reg[20]/NET0131  & ~n3435 ;
  assign n7834 = \P1_reg0_reg[20]/NET0131  & n3448 ;
  assign n7835 = \P1_reg0_reg[20]/NET0131  & ~n4396 ;
  assign n7836 = n4396 & n6492 ;
  assign n7837 = ~n7835 & ~n7836 ;
  assign n7838 = n1936 & ~n7837 ;
  assign n7843 = n4396 & ~n6505 ;
  assign n7844 = ~n7835 & ~n7843 ;
  assign n7845 = ~n3563 & ~n7844 ;
  assign n7840 = n4396 & ~n6499 ;
  assign n7841 = ~n7835 & ~n7840 ;
  assign n7842 = ~n3677 & ~n7841 ;
  assign n7846 = n4396 & n6510 ;
  assign n7847 = ~n7835 & ~n7846 ;
  assign n7848 = n3712 & ~n7847 ;
  assign n7839 = n4396 & n6515 ;
  assign n7849 = \P1_reg0_reg[20]/NET0131  & ~n4493 ;
  assign n7850 = ~n7839 & ~n7849 ;
  assign n7851 = ~n7848 & n7850 ;
  assign n7852 = ~n7842 & n7851 ;
  assign n7853 = ~n7845 & n7852 ;
  assign n7854 = ~n7838 & n7853 ;
  assign n7855 = n3450 & ~n7854 ;
  assign n7856 = ~n7834 & ~n7855 ;
  assign n7857 = \P1_state_reg[0]/NET0131  & ~n7856 ;
  assign n7858 = ~n7833 & ~n7857 ;
  assign n7859 = \P1_reg0_reg[21]/NET0131  & ~n3435 ;
  assign n7860 = \P1_reg0_reg[21]/NET0131  & n3448 ;
  assign n7862 = \P1_reg0_reg[21]/NET0131  & ~n4396 ;
  assign n7863 = n4396 & n6962 ;
  assign n7864 = ~n7862 & ~n7863 ;
  assign n7865 = n1936 & ~n7864 ;
  assign n7872 = n4396 & n6979 ;
  assign n7873 = ~n7862 & ~n7872 ;
  assign n7874 = n3712 & ~n7873 ;
  assign n7861 = n4396 & n6955 ;
  assign n7875 = \P1_reg0_reg[21]/NET0131  & ~n4493 ;
  assign n7876 = ~n7861 & ~n7875 ;
  assign n7877 = ~n7874 & n7876 ;
  assign n7878 = ~n7865 & n7877 ;
  assign n7866 = n4396 & ~n6968 ;
  assign n7867 = ~n7862 & ~n7866 ;
  assign n7868 = ~n3563 & ~n7867 ;
  assign n7869 = n4396 & n6974 ;
  assign n7870 = ~n7862 & ~n7869 ;
  assign n7871 = ~n3677 & ~n7870 ;
  assign n7879 = ~n7868 & ~n7871 ;
  assign n7880 = n7878 & n7879 ;
  assign n7881 = n3450 & ~n7880 ;
  assign n7882 = ~n7860 & ~n7881 ;
  assign n7883 = \P1_state_reg[0]/NET0131  & ~n7882 ;
  assign n7884 = ~n7859 & ~n7883 ;
  assign n7885 = \P1_reg0_reg[30]/NET0131  & ~n6887 ;
  assign n7886 = n6886 & ~n7494 ;
  assign n7887 = ~n7885 & ~n7886 ;
  assign n7888 = \P1_reg1_reg[12]/NET0131  & ~n3435 ;
  assign n7889 = \P1_reg1_reg[12]/NET0131  & n3448 ;
  assign n7891 = \P1_reg1_reg[12]/NET0131  & ~n4532 ;
  assign n7892 = n4532 & n6098 ;
  assign n7893 = ~n7891 & ~n7892 ;
  assign n7894 = n1936 & ~n7893 ;
  assign n7898 = n4532 & ~n6110 ;
  assign n7899 = ~n7891 & ~n7898 ;
  assign n7900 = ~n3677 & ~n7899 ;
  assign n7895 = n4532 & n6104 ;
  assign n7896 = ~n7891 & ~n7895 ;
  assign n7897 = ~n3563 & ~n7896 ;
  assign n7901 = n4532 & n6117 ;
  assign n7902 = ~n7891 & ~n7901 ;
  assign n7903 = n3712 & ~n7902 ;
  assign n7890 = n4532 & n7532 ;
  assign n7904 = \P1_reg1_reg[12]/NET0131  & ~n4541 ;
  assign n7905 = ~n7890 & ~n7904 ;
  assign n7906 = ~n7903 & n7905 ;
  assign n7907 = ~n7897 & n7906 ;
  assign n7908 = ~n7900 & n7907 ;
  assign n7909 = ~n7894 & n7908 ;
  assign n7910 = n3450 & ~n7909 ;
  assign n7911 = ~n7889 & ~n7910 ;
  assign n7912 = \P1_state_reg[0]/NET0131  & ~n7911 ;
  assign n7913 = ~n7888 & ~n7912 ;
  assign n7914 = \P1_reg1_reg[16]/NET0131  & ~n3435 ;
  assign n7915 = \P1_reg1_reg[16]/NET0131  & n3448 ;
  assign n7916 = n4532 & ~n7826 ;
  assign n7917 = ~n4532 & ~n6846 ;
  assign n7918 = n4573 & ~n7917 ;
  assign n7919 = \P1_reg1_reg[16]/NET0131  & ~n7918 ;
  assign n7920 = ~n7916 & ~n7919 ;
  assign n7921 = n3450 & ~n7920 ;
  assign n7922 = ~n7915 & ~n7921 ;
  assign n7923 = \P1_state_reg[0]/NET0131  & ~n7922 ;
  assign n7924 = ~n7914 & ~n7923 ;
  assign n7925 = \P1_reg1_reg[20]/NET0131  & ~n3435 ;
  assign n7926 = \P1_reg1_reg[20]/NET0131  & n3448 ;
  assign n7927 = \P1_reg1_reg[20]/NET0131  & ~n4532 ;
  assign n7928 = n4532 & n6492 ;
  assign n7929 = ~n7927 & ~n7928 ;
  assign n7930 = n1936 & ~n7929 ;
  assign n7935 = n4532 & ~n6505 ;
  assign n7936 = ~n7927 & ~n7935 ;
  assign n7937 = ~n3563 & ~n7936 ;
  assign n7932 = n4532 & ~n6499 ;
  assign n7933 = ~n7927 & ~n7932 ;
  assign n7934 = ~n3677 & ~n7933 ;
  assign n7938 = n4532 & n6510 ;
  assign n7939 = ~n7927 & ~n7938 ;
  assign n7940 = n3712 & ~n7939 ;
  assign n7931 = n4532 & n6515 ;
  assign n7941 = \P1_reg1_reg[20]/NET0131  & ~n4541 ;
  assign n7942 = ~n7931 & ~n7941 ;
  assign n7943 = ~n7940 & n7942 ;
  assign n7944 = ~n7934 & n7943 ;
  assign n7945 = ~n7937 & n7944 ;
  assign n7946 = ~n7930 & n7945 ;
  assign n7947 = n3450 & ~n7946 ;
  assign n7948 = ~n7926 & ~n7947 ;
  assign n7949 = \P1_state_reg[0]/NET0131  & ~n7948 ;
  assign n7950 = ~n7925 & ~n7949 ;
  assign n7951 = \P2_reg0_reg[12]/NET0131  & ~n1983 ;
  assign n7952 = \P2_reg0_reg[12]/NET0131  & n2024 ;
  assign n7954 = \P2_reg0_reg[12]/NET0131  & ~n2040 ;
  assign n7955 = n2040 & n6186 ;
  assign n7956 = ~n7954 & ~n7955 ;
  assign n7957 = n3411 & ~n7956 ;
  assign n7961 = n2040 & ~n6198 ;
  assign n7962 = ~n7954 & ~n7961 ;
  assign n7963 = ~n3320 & ~n7962 ;
  assign n7958 = n2040 & n6192 ;
  assign n7959 = ~n7954 & ~n7958 ;
  assign n7960 = ~n3177 & ~n7959 ;
  assign n7953 = n2040 & ~n7585 ;
  assign n7964 = \P2_reg0_reg[12]/NET0131  & ~n3425 ;
  assign n7965 = ~n7953 & ~n7964 ;
  assign n7966 = ~n7960 & n7965 ;
  assign n7967 = ~n7963 & n7966 ;
  assign n7968 = ~n7957 & n7967 ;
  assign n7969 = n2026 & ~n7968 ;
  assign n7970 = ~n7952 & ~n7969 ;
  assign n7971 = \P1_state_reg[0]/NET0131  & ~n7970 ;
  assign n7972 = ~n7951 & ~n7971 ;
  assign n7973 = \P2_reg0_reg[16]/NET0131  & ~n1983 ;
  assign n7974 = \P2_reg0_reg[16]/NET0131  & n2024 ;
  assign n7982 = ~n3320 & ~n6246 ;
  assign n7983 = ~n7752 & ~n7982 ;
  assign n7984 = n2040 & ~n7983 ;
  assign n7975 = \P2_reg0_reg[16]/NET0131  & ~n2040 ;
  assign n7979 = n2040 & n6240 ;
  assign n7980 = ~n7975 & ~n7979 ;
  assign n7981 = n3355 & ~n7980 ;
  assign n7985 = \P2_reg0_reg[16]/NET0131  & ~n7506 ;
  assign n7989 = ~n7981 & ~n7985 ;
  assign n7990 = ~n7984 & n7989 ;
  assign n7976 = n2040 & ~n6226 ;
  assign n7977 = ~n7975 & ~n7976 ;
  assign n7978 = ~n3177 & ~n7977 ;
  assign n7986 = n2040 & n6234 ;
  assign n7987 = ~n7975 & ~n7986 ;
  assign n7988 = n3411 & ~n7987 ;
  assign n7991 = ~n7978 & ~n7988 ;
  assign n7992 = n7990 & n7991 ;
  assign n7993 = n2026 & ~n7992 ;
  assign n7994 = ~n7974 & ~n7993 ;
  assign n7995 = \P1_state_reg[0]/NET0131  & ~n7994 ;
  assign n7996 = ~n7973 & ~n7995 ;
  assign n7999 = n1203 & n3448 ;
  assign n8001 = n1203 & ~n3980 ;
  assign n8002 = n1772 & ~n4404 ;
  assign n8003 = ~n1772 & n4404 ;
  assign n8004 = ~n8002 & ~n8003 ;
  assign n8005 = n3980 & ~n8004 ;
  assign n8006 = ~n8001 & ~n8005 ;
  assign n8007 = ~n3677 & ~n8006 ;
  assign n8022 = n1198 & ~n6114 ;
  assign n8023 = ~n6115 & ~n8022 ;
  assign n8024 = n3712 & n8023 ;
  assign n8025 = n3980 & n8024 ;
  assign n8000 = n1203 & ~n4910 ;
  assign n8026 = n1198 & ~n4067 ;
  assign n8027 = ~n8000 & ~n8026 ;
  assign n8028 = ~n8025 & n8027 ;
  assign n8029 = ~n8007 & n8028 ;
  assign n8008 = n1772 & ~n4447 ;
  assign n8009 = ~n1772 & n4447 ;
  assign n8010 = ~n8008 & ~n8009 ;
  assign n8011 = n3980 & n8010 ;
  assign n8012 = ~n8001 & ~n8011 ;
  assign n8013 = ~n3563 & ~n8012 ;
  assign n8014 = n1174 & ~n4069 ;
  assign n8015 = ~n4070 & ~n8014 ;
  assign n8016 = ~n537 & ~n8015 ;
  assign n8017 = n537 & n1218 ;
  assign n8018 = ~n8016 & ~n8017 ;
  assign n8019 = n3980 & n8018 ;
  assign n8020 = ~n8001 & ~n8019 ;
  assign n8021 = n1936 & ~n8020 ;
  assign n8030 = ~n8013 & ~n8021 ;
  assign n8031 = n8029 & n8030 ;
  assign n8032 = n3450 & ~n8031 ;
  assign n8033 = ~n7999 & ~n8032 ;
  assign n8034 = \P1_state_reg[0]/NET0131  & ~n8033 ;
  assign n7997 = \P1_reg3_reg[11]/NET0131  & ~\P1_state_reg[0]/NET0131  ;
  assign n7998 = n1203 & n1953 ;
  assign n8035 = ~n7997 & ~n7998 ;
  assign n8036 = ~n8034 & n8035 ;
  assign n8039 = n1113 & n3448 ;
  assign n8041 = n1113 & ~n3980 ;
  assign n8051 = ~n1815 & ~n6031 ;
  assign n8052 = n1815 & n6031 ;
  assign n8053 = ~n8051 & ~n8052 ;
  assign n8054 = ~n3563 & ~n8053 ;
  assign n8055 = n1815 & ~n6019 ;
  assign n8056 = ~n1815 & n6019 ;
  assign n8057 = ~n8055 & ~n8056 ;
  assign n8058 = ~n8054 & n8057 ;
  assign n8059 = n3980 & ~n8058 ;
  assign n8060 = ~n8041 & ~n8059 ;
  assign n8061 = ~n3563 & ~n3980 ;
  assign n8062 = n3677 & ~n8054 ;
  assign n8063 = ~n8061 & n8062 ;
  assign n8064 = ~n8060 & ~n8063 ;
  assign n8042 = ~n1094 & ~n7130 ;
  assign n8043 = n1094 & n7130 ;
  assign n8044 = ~n8042 & ~n8043 ;
  assign n8045 = ~n537 & ~n8044 ;
  assign n8046 = n537 & ~n1146 ;
  assign n8047 = ~n8045 & ~n8046 ;
  assign n8048 = n3980 & ~n8047 ;
  assign n8049 = ~n8041 & ~n8048 ;
  assign n8050 = n1936 & ~n8049 ;
  assign n8065 = ~n1109 & n5440 ;
  assign n8066 = n1109 & ~n5440 ;
  assign n8067 = ~n8065 & ~n8066 ;
  assign n8068 = n3980 & n8067 ;
  assign n8069 = ~n8041 & ~n8068 ;
  assign n8070 = n3712 & ~n8069 ;
  assign n8040 = n1113 & ~n4064 ;
  assign n8071 = n1109 & ~n4067 ;
  assign n8072 = ~n8040 & ~n8071 ;
  assign n8073 = ~n8070 & n8072 ;
  assign n8074 = ~n8050 & n8073 ;
  assign n8075 = ~n8064 & n8074 ;
  assign n8076 = n3450 & ~n8075 ;
  assign n8077 = ~n8039 & ~n8076 ;
  assign n8078 = \P1_state_reg[0]/NET0131  & ~n8077 ;
  assign n8037 = n1113 & n1953 ;
  assign n8038 = \P1_reg3_reg[14]/NET0131  & ~\P1_state_reg[0]/NET0131  ;
  assign n8079 = ~n8037 & ~n8038 ;
  assign n8080 = ~n8078 & n8079 ;
  assign n8083 = n1088 & n3448 ;
  assign n8085 = n1088 & ~n3980 ;
  assign n8086 = n1788 & ~n7414 ;
  assign n8087 = ~n1788 & n7414 ;
  assign n8088 = ~n8086 & ~n8087 ;
  assign n8089 = n3980 & ~n8088 ;
  assign n8090 = ~n8085 & ~n8089 ;
  assign n8091 = ~n3677 & ~n8090 ;
  assign n8106 = n1083 & ~n8065 ;
  assign n8107 = ~n5441 & ~n8106 ;
  assign n8108 = n3712 & n8107 ;
  assign n8109 = n3980 & n8108 ;
  assign n8084 = n1088 & ~n4910 ;
  assign n8110 = n1083 & ~n4067 ;
  assign n8111 = ~n8084 & ~n8110 ;
  assign n8112 = ~n8109 & n8111 ;
  assign n8113 = ~n8091 & n8112 ;
  assign n8092 = n1788 & ~n7427 ;
  assign n8093 = ~n1788 & n7427 ;
  assign n8094 = ~n8092 & ~n8093 ;
  assign n8095 = n3980 & n8094 ;
  assign n8096 = ~n8085 & ~n8095 ;
  assign n8097 = ~n3563 & ~n8096 ;
  assign n8098 = n1475 & ~n4470 ;
  assign n8099 = ~n4073 & ~n8098 ;
  assign n8100 = ~n537 & ~n8099 ;
  assign n8101 = n537 & n1118 ;
  assign n8102 = ~n8100 & ~n8101 ;
  assign n8103 = n3980 & n8102 ;
  assign n8104 = ~n8085 & ~n8103 ;
  assign n8105 = n1936 & ~n8104 ;
  assign n8114 = ~n8097 & ~n8105 ;
  assign n8115 = n8113 & n8114 ;
  assign n8116 = n3450 & ~n8115 ;
  assign n8117 = ~n8083 & ~n8116 ;
  assign n8118 = \P1_state_reg[0]/NET0131  & ~n8117 ;
  assign n8081 = n1088 & n1953 ;
  assign n8082 = \P1_reg3_reg[15]/NET0131  & ~\P1_state_reg[0]/NET0131  ;
  assign n8119 = ~n8081 & ~n8082 ;
  assign n8120 = ~n8118 & n8119 ;
  assign n8122 = n2024 & n2681 ;
  assign n8124 = n2681 & ~n3788 ;
  assign n8125 = n2715 & ~n6179 ;
  assign n8126 = ~n6180 & ~n8125 ;
  assign n8127 = ~n2058 & ~n8126 ;
  assign n8128 = n2058 & n2742 ;
  assign n8129 = ~n8127 & ~n8128 ;
  assign n8130 = n3788 & n8129 ;
  assign n8131 = ~n8124 & ~n8130 ;
  assign n8132 = n3411 & ~n8131 ;
  assign n8133 = n4201 & ~n4804 ;
  assign n8134 = ~n4201 & n4804 ;
  assign n8135 = ~n8133 & ~n8134 ;
  assign n8136 = n3788 & n8135 ;
  assign n8137 = ~n8124 & ~n8136 ;
  assign n8138 = ~n3177 & ~n8137 ;
  assign n8139 = n2704 & ~n7179 ;
  assign n8140 = ~n3336 & ~n8139 ;
  assign n8141 = n3788 & n8140 ;
  assign n8142 = ~n8124 & ~n8141 ;
  assign n8143 = n3355 & ~n8142 ;
  assign n8144 = n4201 & ~n4840 ;
  assign n8145 = ~n4201 & n4840 ;
  assign n8146 = ~n8144 & ~n8145 ;
  assign n8147 = ~n3320 & ~n8146 ;
  assign n8148 = n3788 & n8147 ;
  assign n8123 = n2681 & ~n6312 ;
  assign n8149 = n2704 & ~n3965 ;
  assign n8150 = ~n8123 & ~n8149 ;
  assign n8151 = ~n8148 & n8150 ;
  assign n8152 = ~n8143 & n8151 ;
  assign n8153 = ~n8138 & n8152 ;
  assign n8154 = ~n8132 & n8153 ;
  assign n8155 = n2026 & ~n8154 ;
  assign n8156 = ~n8122 & ~n8155 ;
  assign n8157 = \P1_state_reg[0]/NET0131  & ~n8156 ;
  assign n8121 = ~\P1_state_reg[0]/NET0131  & \P2_reg3_reg[11]/NET0131  ;
  assign n8158 = n2681 & n3976 ;
  assign n8159 = ~n8121 & ~n8158 ;
  assign n8160 = ~n8157 & n8159 ;
  assign n8163 = n2024 & n2866 ;
  assign n8166 = n2866 & ~n3788 ;
  assign n8167 = n2828 & ~n3387 ;
  assign n8168 = ~n5564 & ~n8167 ;
  assign n8169 = ~n2058 & ~n8168 ;
  assign n8170 = n2058 & n2880 ;
  assign n8171 = ~n8169 & ~n8170 ;
  assign n8172 = n3788 & n8171 ;
  assign n8173 = ~n8166 & ~n8172 ;
  assign n8174 = n3411 & ~n8173 ;
  assign n8164 = n2860 & ~n3965 ;
  assign n8165 = n2866 & ~n3962 ;
  assign n8192 = ~n8164 & ~n8165 ;
  assign n8193 = ~n8174 & n8192 ;
  assign n8186 = n4210 & ~n4714 ;
  assign n8187 = ~n4210 & n4714 ;
  assign n8188 = ~n8186 & ~n8187 ;
  assign n8189 = n3788 & ~n8188 ;
  assign n8190 = ~n8166 & ~n8189 ;
  assign n8191 = ~n3320 & ~n8190 ;
  assign n8175 = n2860 & ~n7215 ;
  assign n8176 = ~n3339 & ~n8175 ;
  assign n8177 = n3788 & n8176 ;
  assign n8178 = ~n8166 & ~n8177 ;
  assign n8179 = n3355 & ~n8178 ;
  assign n8180 = n4210 & ~n4745 ;
  assign n8181 = ~n4210 & n4745 ;
  assign n8182 = ~n8180 & ~n8181 ;
  assign n8183 = n3788 & n8182 ;
  assign n8184 = ~n8166 & ~n8183 ;
  assign n8185 = ~n3177 & ~n8184 ;
  assign n8194 = ~n8179 & ~n8185 ;
  assign n8195 = ~n8191 & n8194 ;
  assign n8196 = n8193 & n8195 ;
  assign n8197 = n2026 & ~n8196 ;
  assign n8198 = ~n8163 & ~n8197 ;
  assign n8199 = \P1_state_reg[0]/NET0131  & ~n8198 ;
  assign n8161 = n2866 & n3976 ;
  assign n8162 = ~\P1_state_reg[0]/NET0131  & \P2_reg3_reg[14]/NET0131  ;
  assign n8200 = ~n8161 & ~n8162 ;
  assign n8201 = ~n8199 & n8200 ;
  assign n8204 = n2024 & n2822 ;
  assign n8206 = n2822 & ~n3788 ;
  assign n8215 = n4215 & ~n4809 ;
  assign n8216 = ~n4215 & n4809 ;
  assign n8217 = ~n8215 & ~n8216 ;
  assign n8218 = n3788 & n8217 ;
  assign n8219 = ~n8206 & ~n8218 ;
  assign n8220 = ~n3177 & ~n8219 ;
  assign n8207 = n2804 & ~n5564 ;
  assign n8208 = ~n5565 & ~n8207 ;
  assign n8209 = ~n2058 & ~n8208 ;
  assign n8210 = n2058 & n2870 ;
  assign n8211 = ~n8209 & ~n8210 ;
  assign n8212 = n3788 & n8211 ;
  assign n8213 = ~n8206 & ~n8212 ;
  assign n8214 = n3411 & ~n8213 ;
  assign n8221 = n2843 & ~n3339 ;
  assign n8222 = ~n5574 & ~n8221 ;
  assign n8223 = n3788 & n8222 ;
  assign n8224 = ~n8206 & ~n8223 ;
  assign n8225 = n3355 & ~n8224 ;
  assign n8226 = n4215 & ~n4845 ;
  assign n8227 = ~n4215 & n4845 ;
  assign n8228 = ~n8226 & ~n8227 ;
  assign n8229 = n3788 & ~n8228 ;
  assign n8230 = ~n8206 & ~n8229 ;
  assign n8231 = ~n3320 & ~n8230 ;
  assign n8205 = n2843 & ~n3965 ;
  assign n8232 = n2822 & ~n3962 ;
  assign n8233 = ~n8205 & ~n8232 ;
  assign n8234 = ~n8231 & n8233 ;
  assign n8235 = ~n8225 & n8234 ;
  assign n8236 = ~n8214 & n8235 ;
  assign n8237 = ~n8220 & n8236 ;
  assign n8238 = n2026 & ~n8237 ;
  assign n8239 = ~n8204 & ~n8238 ;
  assign n8240 = \P1_state_reg[0]/NET0131  & ~n8239 ;
  assign n8202 = n2822 & n3976 ;
  assign n8203 = ~\P1_state_reg[0]/NET0131  & \P2_reg3_reg[15]/NET0131  ;
  assign n8241 = ~n8202 & ~n8203 ;
  assign n8242 = ~n8240 & n8241 ;
  assign n8245 = n2024 & n2447 ;
  assign n8247 = n2447 & ~n3788 ;
  assign n8248 = n2765 & ~n7242 ;
  assign n8249 = ~n7243 & ~n8248 ;
  assign n8250 = ~n2058 & ~n8249 ;
  assign n8251 = n2058 & n2480 ;
  assign n8252 = ~n8250 & ~n8251 ;
  assign n8253 = n3788 & n8252 ;
  assign n8254 = ~n8247 & ~n8253 ;
  assign n8255 = n3411 & ~n8254 ;
  assign n8262 = ~n3831 & n4208 ;
  assign n8263 = n3831 & ~n4208 ;
  assign n8264 = ~n8262 & ~n8263 ;
  assign n8265 = n3788 & ~n8264 ;
  assign n8266 = ~n8247 & ~n8265 ;
  assign n8267 = ~n3320 & ~n8266 ;
  assign n8256 = ~n3889 & n4208 ;
  assign n8257 = n3889 & ~n4208 ;
  assign n8258 = ~n8256 & ~n8257 ;
  assign n8259 = n3788 & n8258 ;
  assign n8260 = ~n8247 & ~n8259 ;
  assign n8261 = ~n3177 & ~n8260 ;
  assign n8268 = n2470 & ~n3332 ;
  assign n8269 = ~n7258 & ~n8268 ;
  assign n8270 = n3355 & n8269 ;
  assign n8271 = n3788 & n8270 ;
  assign n8246 = n2447 & ~n5698 ;
  assign n8272 = n2470 & ~n3965 ;
  assign n8273 = ~n8246 & ~n8272 ;
  assign n8274 = ~n8271 & n8273 ;
  assign n8275 = ~n8261 & n8274 ;
  assign n8276 = ~n8267 & n8275 ;
  assign n8277 = ~n8255 & n8276 ;
  assign n8278 = n2026 & ~n8277 ;
  assign n8279 = ~n8245 & ~n8278 ;
  assign n8280 = \P1_state_reg[0]/NET0131  & ~n8279 ;
  assign n8243 = ~\P1_state_reg[0]/NET0131  & \P2_reg3_reg[8]/NET0131  ;
  assign n8244 = n2447 & n3976 ;
  assign n8281 = ~n8243 & ~n8244 ;
  assign n8282 = ~n8280 & n8281 ;
  assign n8285 = n1262 & n3448 ;
  assign n8287 = n1262 & ~n3980 ;
  assign n8288 = n1244 & ~n7305 ;
  assign n8289 = ~n7306 & ~n8288 ;
  assign n8290 = ~n537 & ~n8289 ;
  assign n8291 = n537 & n1498 ;
  assign n8292 = ~n8290 & ~n8291 ;
  assign n8293 = n3980 & n8292 ;
  assign n8294 = ~n8287 & ~n8293 ;
  assign n8295 = n1936 & ~n8294 ;
  assign n8302 = ~n1746 & n1802 ;
  assign n8303 = n1746 & ~n1802 ;
  assign n8304 = ~n8302 & ~n8303 ;
  assign n8305 = n3980 & ~n8304 ;
  assign n8306 = ~n8287 & ~n8305 ;
  assign n8307 = ~n3677 & ~n8306 ;
  assign n8296 = n1802 & ~n3996 ;
  assign n8297 = ~n1802 & n3996 ;
  assign n8298 = ~n8296 & ~n8297 ;
  assign n8299 = n3980 & n8298 ;
  assign n8300 = ~n8287 & ~n8299 ;
  assign n8301 = ~n3563 & ~n8300 ;
  assign n8308 = n1514 & n3684 ;
  assign n8309 = n1281 & ~n8308 ;
  assign n8310 = ~n7298 & ~n8309 ;
  assign n8311 = n3980 & n8310 ;
  assign n8312 = ~n8287 & ~n8311 ;
  assign n8313 = n3712 & ~n8312 ;
  assign n8286 = n1281 & ~n4067 ;
  assign n8314 = n1262 & ~n4064 ;
  assign n8315 = ~n8286 & ~n8314 ;
  assign n8316 = ~n8313 & n8315 ;
  assign n8317 = ~n8301 & n8316 ;
  assign n8318 = ~n8307 & n8317 ;
  assign n8319 = ~n8295 & n8318 ;
  assign n8320 = n3450 & ~n8319 ;
  assign n8321 = ~n8285 & ~n8320 ;
  assign n8322 = \P1_state_reg[0]/NET0131  & ~n8321 ;
  assign n8283 = \P1_reg3_reg[8]/NET0131  & ~\P1_state_reg[0]/NET0131  ;
  assign n8284 = n1262 & n1953 ;
  assign n8323 = ~n8283 & ~n8284 ;
  assign n8324 = ~n8322 & n8323 ;
  assign n8325 = n2024 & n3084 ;
  assign n8326 = n3084 & ~n3788 ;
  assign n8327 = ~n4814 & n4816 ;
  assign n8328 = n4821 & ~n8327 ;
  assign n8329 = n4196 & ~n8328 ;
  assign n8330 = ~n4196 & n8328 ;
  assign n8331 = ~n8329 & ~n8330 ;
  assign n8332 = n3788 & n8331 ;
  assign n8333 = ~n8326 & ~n8332 ;
  assign n8334 = ~n3177 & ~n8333 ;
  assign n8335 = n3079 & ~n5768 ;
  assign n8336 = ~n4614 & ~n8335 ;
  assign n8337 = n3788 & n8336 ;
  assign n8338 = ~n8326 & ~n8337 ;
  assign n8339 = n3355 & ~n8338 ;
  assign n8340 = ~n4850 & n4851 ;
  assign n8341 = n4856 & ~n8340 ;
  assign n8342 = n4196 & ~n8341 ;
  assign n8343 = ~n4196 & n8341 ;
  assign n8344 = ~n8342 & ~n8343 ;
  assign n8345 = n3788 & ~n8344 ;
  assign n8346 = ~n8326 & ~n8345 ;
  assign n8347 = ~n3320 & ~n8346 ;
  assign n8348 = n2058 & ~n3112 ;
  assign n8349 = n3065 & ~n5775 ;
  assign n8350 = ~n2058 & ~n4622 ;
  assign n8351 = ~n8349 & n8350 ;
  assign n8352 = ~n8348 & ~n8351 ;
  assign n8353 = n3788 & ~n8352 ;
  assign n8354 = ~n8326 & ~n8353 ;
  assign n8355 = n3411 & ~n8354 ;
  assign n8356 = n3084 & ~n3962 ;
  assign n8357 = n3079 & ~n3965 ;
  assign n8358 = ~n8356 & ~n8357 ;
  assign n8359 = ~n8355 & n8358 ;
  assign n8360 = ~n8347 & n8359 ;
  assign n8361 = ~n8339 & n8360 ;
  assign n8362 = ~n8334 & n8361 ;
  assign n8363 = n2026 & ~n8362 ;
  assign n8364 = ~n8325 & ~n8363 ;
  assign n8365 = \P1_state_reg[0]/NET0131  & ~n8364 ;
  assign n8366 = ~\P1_state_reg[0]/NET0131  & \P2_reg3_reg[23]/NET0131  ;
  assign n8367 = n3084 & n3976 ;
  assign n8368 = ~n8366 & ~n8367 ;
  assign n8369 = ~n8365 & n8368 ;
  assign n8370 = \P2_reg0_reg[23]/NET0131  & ~n1983 ;
  assign n8371 = \P2_reg0_reg[23]/NET0131  & n2024 ;
  assign n8372 = \P2_reg0_reg[23]/NET0131  & ~n2040 ;
  assign n8373 = n2040 & n8331 ;
  assign n8374 = ~n8372 & ~n8373 ;
  assign n8375 = ~n3177 & ~n8374 ;
  assign n8376 = n3355 & n8336 ;
  assign n8377 = n3079 & n3358 ;
  assign n8378 = ~n3320 & ~n8344 ;
  assign n8379 = ~n8377 & ~n8378 ;
  assign n8380 = ~n8376 & n8379 ;
  assign n8381 = n2040 & ~n8380 ;
  assign n8382 = n2040 & ~n8352 ;
  assign n8383 = ~n8372 & ~n8382 ;
  assign n8384 = n3411 & ~n8383 ;
  assign n8385 = ~n3424 & n7506 ;
  assign n8386 = \P2_reg0_reg[23]/NET0131  & ~n8385 ;
  assign n8387 = ~n8384 & ~n8386 ;
  assign n8388 = ~n8381 & n8387 ;
  assign n8389 = ~n8375 & n8388 ;
  assign n8390 = n2026 & ~n8389 ;
  assign n8391 = ~n8371 & ~n8390 ;
  assign n8392 = \P1_state_reg[0]/NET0131  & ~n8391 ;
  assign n8393 = ~n8370 & ~n8392 ;
  assign n8394 = \P1_reg1_reg[9]/NET0131  & ~n3435 ;
  assign n8395 = \P1_reg1_reg[9]/NET0131  & n3448 ;
  assign n8398 = \P1_reg1_reg[9]/NET0131  & ~n4532 ;
  assign n8408 = n4532 & ~n7310 ;
  assign n8409 = ~n8398 & ~n8408 ;
  assign n8410 = n1936 & ~n8409 ;
  assign n8402 = n4532 & ~n7288 ;
  assign n8403 = ~n8398 & ~n8402 ;
  assign n8404 = ~n3677 & ~n8403 ;
  assign n8399 = n4532 & n7294 ;
  assign n8400 = ~n8398 & ~n8399 ;
  assign n8401 = ~n3563 & ~n8400 ;
  assign n8405 = n4532 & n7300 ;
  assign n8406 = ~n8398 & ~n8405 ;
  assign n8407 = n3712 & ~n8406 ;
  assign n8396 = n1257 & n1880 ;
  assign n8397 = n4532 & n8396 ;
  assign n8411 = \P1_reg1_reg[9]/NET0131  & ~n4541 ;
  assign n8412 = ~n8397 & ~n8411 ;
  assign n8413 = ~n8407 & n8412 ;
  assign n8414 = ~n8401 & n8413 ;
  assign n8415 = ~n8404 & n8414 ;
  assign n8416 = ~n8410 & n8415 ;
  assign n8417 = n3450 & ~n8416 ;
  assign n8418 = ~n8395 & ~n8417 ;
  assign n8419 = \P1_state_reg[0]/NET0131  & ~n8418 ;
  assign n8420 = ~n8394 & ~n8419 ;
  assign n8421 = \P1_reg2_reg[10]/NET0131  & ~n3435 ;
  assign n8422 = \P1_reg2_reg[10]/NET0131  & n3448 ;
  assign n8425 = \P1_reg2_reg[10]/NET0131  & ~n3466 ;
  assign n8426 = n3466 & n7086 ;
  assign n8427 = ~n8425 & ~n8426 ;
  assign n8428 = n1936 & ~n8427 ;
  assign n8435 = n3466 & n7097 ;
  assign n8436 = ~n8425 & ~n8435 ;
  assign n8437 = n3712 & ~n8436 ;
  assign n8439 = \P1_reg2_reg[10]/NET0131  & ~n3718 ;
  assign n8423 = n1233 & n1880 ;
  assign n8424 = n3466 & n8423 ;
  assign n8438 = n1214 & n1763 ;
  assign n8440 = ~n8424 & ~n8438 ;
  assign n8441 = ~n8439 & n8440 ;
  assign n8442 = ~n8437 & n8441 ;
  assign n8443 = ~n8428 & n8442 ;
  assign n8429 = n3466 & n7092 ;
  assign n8430 = ~n8425 & ~n8429 ;
  assign n8431 = ~n3563 & ~n8430 ;
  assign n8432 = n3466 & ~n7078 ;
  assign n8433 = ~n8425 & ~n8432 ;
  assign n8434 = ~n3677 & ~n8433 ;
  assign n8444 = ~n8431 & ~n8434 ;
  assign n8445 = n8443 & n8444 ;
  assign n8446 = n3450 & ~n8445 ;
  assign n8447 = ~n8422 & ~n8446 ;
  assign n8448 = \P1_state_reg[0]/NET0131  & ~n8447 ;
  assign n8449 = ~n8421 & ~n8448 ;
  assign n8450 = \P1_reg2_reg[13]/NET0131  & ~n3435 ;
  assign n8451 = \P1_reg2_reg[13]/NET0131  & n3448 ;
  assign n8453 = \P1_reg2_reg[13]/NET0131  & ~n3466 ;
  assign n8454 = n3466 & n7125 ;
  assign n8455 = ~n8453 & ~n8454 ;
  assign n8456 = ~n3563 & ~n8455 ;
  assign n8463 = n3466 & n7139 ;
  assign n8464 = ~n8453 & ~n8463 ;
  assign n8465 = n3712 & ~n8464 ;
  assign n8452 = \P1_reg2_reg[13]/NET0131  & ~n3718 ;
  assign n8466 = n1140 & n1763 ;
  assign n8467 = n1136 & n1880 ;
  assign n8468 = n3466 & n8467 ;
  assign n8469 = ~n8466 & ~n8468 ;
  assign n8470 = ~n8452 & n8469 ;
  assign n8471 = ~n8465 & n8470 ;
  assign n8472 = ~n8456 & n8471 ;
  assign n8457 = n3466 & n7134 ;
  assign n8458 = ~n8453 & ~n8457 ;
  assign n8459 = n1936 & ~n8458 ;
  assign n8460 = n3466 & ~n7119 ;
  assign n8461 = ~n8453 & ~n8460 ;
  assign n8462 = ~n3677 & ~n8461 ;
  assign n8473 = ~n8459 & ~n8462 ;
  assign n8474 = n8472 & n8473 ;
  assign n8475 = n3450 & ~n8474 ;
  assign n8476 = ~n8451 & ~n8475 ;
  assign n8477 = \P1_state_reg[0]/NET0131  & ~n8476 ;
  assign n8478 = ~n8450 & ~n8477 ;
  assign n8479 = \P2_reg0_reg[9]/NET0131  & ~n1983 ;
  assign n8480 = \P2_reg0_reg[9]/NET0131  & n2024 ;
  assign n8482 = \P2_reg0_reg[9]/NET0131  & ~n2040 ;
  assign n8483 = n2040 & n7248 ;
  assign n8484 = ~n8482 & ~n8483 ;
  assign n8485 = n3411 & ~n8484 ;
  assign n8486 = n2040 & ~n7254 ;
  assign n8487 = ~n8482 & ~n8486 ;
  assign n8488 = ~n3177 & ~n8487 ;
  assign n8481 = \P2_reg0_reg[9]/NET0131  & ~n8385 ;
  assign n8490 = n3355 & n7260 ;
  assign n8489 = n2779 & n3358 ;
  assign n8491 = ~n7267 & ~n8489 ;
  assign n8492 = ~n8490 & n8491 ;
  assign n8493 = n2040 & ~n8492 ;
  assign n8494 = ~n8481 & ~n8493 ;
  assign n8495 = ~n8488 & n8494 ;
  assign n8496 = ~n8485 & n8495 ;
  assign n8497 = n2026 & ~n8496 ;
  assign n8498 = ~n8480 & ~n8497 ;
  assign n8499 = \P1_state_reg[0]/NET0131  & ~n8498 ;
  assign n8500 = ~n8479 & ~n8499 ;
  assign n8501 = \P2_reg1_reg[10]/NET0131  & ~n1983 ;
  assign n8502 = \P2_reg1_reg[10]/NET0131  & n2024 ;
  assign n8505 = \P2_reg1_reg[10]/NET0131  & ~n3733 ;
  assign n8506 = n3733 & n7163 ;
  assign n8507 = ~n8505 & ~n8506 ;
  assign n8508 = n3411 & ~n8507 ;
  assign n8512 = n3733 & n7175 ;
  assign n8513 = ~n8505 & ~n8512 ;
  assign n8514 = ~n3320 & ~n8513 ;
  assign n8509 = n3733 & ~n7169 ;
  assign n8510 = ~n8505 & ~n8509 ;
  assign n8511 = ~n3177 & ~n8510 ;
  assign n8515 = n3733 & n7181 ;
  assign n8516 = ~n8505 & ~n8515 ;
  assign n8517 = n3355 & ~n8516 ;
  assign n8503 = n2755 & n3358 ;
  assign n8504 = n3733 & n8503 ;
  assign n8518 = \P2_reg1_reg[10]/NET0131  & ~n3743 ;
  assign n8519 = ~n8504 & ~n8518 ;
  assign n8520 = ~n8517 & n8519 ;
  assign n8521 = ~n8511 & n8520 ;
  assign n8522 = ~n8514 & n8521 ;
  assign n8523 = ~n8508 & n8522 ;
  assign n8524 = n2026 & ~n8523 ;
  assign n8525 = ~n8502 & ~n8524 ;
  assign n8526 = \P1_state_reg[0]/NET0131  & ~n8525 ;
  assign n8527 = ~n8501 & ~n8526 ;
  assign n8528 = \P2_reg1_reg[13]/NET0131  & ~n1983 ;
  assign n8529 = \P2_reg1_reg[13]/NET0131  & n2024 ;
  assign n8530 = ~n3733 & ~n6639 ;
  assign n8531 = n3421 & ~n8530 ;
  assign n8532 = ~n7597 & n8531 ;
  assign n8533 = ~n3733 & ~n7508 ;
  assign n8534 = n8532 & ~n8533 ;
  assign n8535 = \P2_reg1_reg[13]/NET0131  & ~n8534 ;
  assign n8541 = n3411 & ~n7205 ;
  assign n8536 = n2893 & n3358 ;
  assign n8537 = ~n3320 & ~n7223 ;
  assign n8538 = ~n8536 & ~n8537 ;
  assign n8539 = n3355 & n7217 ;
  assign n8540 = n8538 & ~n8539 ;
  assign n8542 = ~n3177 & n7211 ;
  assign n8543 = n8540 & ~n8542 ;
  assign n8544 = ~n8541 & n8543 ;
  assign n8545 = n3733 & ~n8544 ;
  assign n8546 = ~n8535 & ~n8545 ;
  assign n8547 = n2026 & ~n8546 ;
  assign n8548 = ~n8529 & ~n8547 ;
  assign n8549 = \P1_state_reg[0]/NET0131  & ~n8548 ;
  assign n8550 = ~n8528 & ~n8549 ;
  assign n8551 = \P2_reg1_reg[23]/NET0131  & ~n1983 ;
  assign n8552 = \P2_reg1_reg[23]/NET0131  & n2024 ;
  assign n8553 = \P2_reg1_reg[23]/NET0131  & ~n3733 ;
  assign n8554 = n3733 & n8331 ;
  assign n8555 = ~n8553 & ~n8554 ;
  assign n8556 = ~n3177 & ~n8555 ;
  assign n8557 = n3733 & ~n8380 ;
  assign n8558 = n3733 & ~n8352 ;
  assign n8559 = ~n8553 & ~n8558 ;
  assign n8560 = n3411 & ~n8559 ;
  assign n8561 = \P2_reg1_reg[23]/NET0131  & ~n8532 ;
  assign n8562 = ~n8560 & ~n8561 ;
  assign n8563 = ~n8557 & n8562 ;
  assign n8564 = ~n8556 & n8563 ;
  assign n8565 = n2026 & ~n8564 ;
  assign n8566 = ~n8552 & ~n8565 ;
  assign n8567 = \P1_state_reg[0]/NET0131  & ~n8566 ;
  assign n8568 = ~n8551 & ~n8567 ;
  assign n8569 = \P1_reg0_reg[10]/NET0131  & ~n3435 ;
  assign n8570 = \P1_reg0_reg[10]/NET0131  & n3448 ;
  assign n8572 = \P1_reg0_reg[10]/NET0131  & ~n4396 ;
  assign n8573 = n4396 & n7092 ;
  assign n8574 = ~n8572 & ~n8573 ;
  assign n8575 = ~n3563 & ~n8574 ;
  assign n8582 = n4396 & n7097 ;
  assign n8583 = ~n8572 & ~n8582 ;
  assign n8584 = n3712 & ~n8583 ;
  assign n8571 = n4396 & n8423 ;
  assign n8585 = \P1_reg0_reg[10]/NET0131  & ~n4493 ;
  assign n8586 = ~n8571 & ~n8585 ;
  assign n8587 = ~n8584 & n8586 ;
  assign n8588 = ~n8575 & n8587 ;
  assign n8576 = n4396 & n7086 ;
  assign n8577 = ~n8572 & ~n8576 ;
  assign n8578 = n1936 & ~n8577 ;
  assign n8579 = n4396 & ~n7078 ;
  assign n8580 = ~n8572 & ~n8579 ;
  assign n8581 = ~n3677 & ~n8580 ;
  assign n8589 = ~n8578 & ~n8581 ;
  assign n8590 = n8588 & n8589 ;
  assign n8591 = n3450 & ~n8590 ;
  assign n8592 = ~n8570 & ~n8591 ;
  assign n8593 = \P1_state_reg[0]/NET0131  & ~n8592 ;
  assign n8594 = ~n8569 & ~n8593 ;
  assign n8595 = \P2_reg1_reg[9]/NET0131  & ~n1983 ;
  assign n8596 = \P2_reg1_reg[9]/NET0131  & n2024 ;
  assign n8598 = \P2_reg1_reg[9]/NET0131  & ~n3733 ;
  assign n8599 = n3733 & n7248 ;
  assign n8600 = ~n8598 & ~n8599 ;
  assign n8601 = n3411 & ~n8600 ;
  assign n8602 = n3733 & ~n7254 ;
  assign n8603 = ~n8598 & ~n8602 ;
  assign n8604 = ~n3177 & ~n8603 ;
  assign n8597 = \P2_reg1_reg[9]/NET0131  & ~n8532 ;
  assign n8605 = n3733 & ~n8492 ;
  assign n8606 = ~n8597 & ~n8605 ;
  assign n8607 = ~n8604 & n8606 ;
  assign n8608 = ~n8601 & n8607 ;
  assign n8609 = n2026 & ~n8608 ;
  assign n8610 = ~n8596 & ~n8609 ;
  assign n8611 = \P1_state_reg[0]/NET0131  & ~n8610 ;
  assign n8612 = ~n8595 & ~n8611 ;
  assign n8613 = \P2_reg2_reg[10]/NET0131  & ~n1983 ;
  assign n8614 = \P2_reg2_reg[10]/NET0131  & n2024 ;
  assign n8616 = \P2_reg2_reg[10]/NET0131  & ~n3758 ;
  assign n8617 = n3758 & n7163 ;
  assign n8618 = ~n8616 & ~n8617 ;
  assign n8619 = n3411 & ~n8618 ;
  assign n8623 = n3758 & n7175 ;
  assign n8624 = ~n8616 & ~n8623 ;
  assign n8625 = ~n3320 & ~n8624 ;
  assign n8620 = n3758 & ~n7169 ;
  assign n8621 = ~n8616 & ~n8620 ;
  assign n8622 = ~n3177 & ~n8621 ;
  assign n8626 = n3758 & n7181 ;
  assign n8627 = ~n8616 & ~n8626 ;
  assign n8628 = n3355 & ~n8627 ;
  assign n8630 = \P2_reg2_reg[10]/NET0131  & ~n3774 ;
  assign n8615 = n3758 & n8503 ;
  assign n8629 = n2735 & n3420 ;
  assign n8631 = ~n8615 & ~n8629 ;
  assign n8632 = ~n8630 & n8631 ;
  assign n8633 = ~n8628 & n8632 ;
  assign n8634 = ~n8622 & n8633 ;
  assign n8635 = ~n8625 & n8634 ;
  assign n8636 = ~n8619 & n8635 ;
  assign n8637 = n2026 & ~n8636 ;
  assign n8638 = ~n8614 & ~n8637 ;
  assign n8639 = \P1_state_reg[0]/NET0131  & ~n8638 ;
  assign n8640 = ~n8613 & ~n8639 ;
  assign n8641 = \P2_reg2_reg[13]/NET0131  & ~n1983 ;
  assign n8642 = \P2_reg2_reg[13]/NET0131  & n2024 ;
  assign n8644 = \P2_reg2_reg[13]/NET0131  & ~n3758 ;
  assign n8645 = n3758 & ~n7205 ;
  assign n8646 = ~n8644 & ~n8645 ;
  assign n8647 = n3411 & ~n8646 ;
  assign n8648 = n3758 & n7211 ;
  assign n8649 = ~n8644 & ~n8648 ;
  assign n8650 = ~n3177 & ~n8649 ;
  assign n8651 = n3758 & n7217 ;
  assign n8652 = ~n8644 & ~n8651 ;
  assign n8653 = n3355 & ~n8652 ;
  assign n8654 = n3758 & ~n8538 ;
  assign n8643 = \P2_reg2_reg[13]/NET0131  & ~n7770 ;
  assign n8655 = n2874 & n3420 ;
  assign n8656 = ~n8643 & ~n8655 ;
  assign n8657 = ~n8654 & n8656 ;
  assign n8658 = ~n8653 & n8657 ;
  assign n8659 = ~n8650 & n8658 ;
  assign n8660 = ~n8647 & n8659 ;
  assign n8661 = n2026 & ~n8660 ;
  assign n8662 = ~n8642 & ~n8661 ;
  assign n8663 = \P1_state_reg[0]/NET0131  & ~n8662 ;
  assign n8664 = ~n8641 & ~n8663 ;
  assign n8665 = \P1_reg2_reg[9]/NET0131  & ~n3435 ;
  assign n8666 = \P1_reg2_reg[9]/NET0131  & n3448 ;
  assign n8668 = \P1_reg2_reg[9]/NET0131  & ~n3466 ;
  assign n8678 = n3466 & ~n7310 ;
  assign n8679 = ~n8668 & ~n8678 ;
  assign n8680 = n1936 & ~n8679 ;
  assign n8672 = n3466 & ~n7288 ;
  assign n8673 = ~n8668 & ~n8672 ;
  assign n8674 = ~n3677 & ~n8673 ;
  assign n8669 = n3466 & n7294 ;
  assign n8670 = ~n8668 & ~n8669 ;
  assign n8671 = ~n3563 & ~n8670 ;
  assign n8675 = n3466 & n7300 ;
  assign n8676 = ~n8668 & ~n8675 ;
  assign n8677 = n3712 & ~n8676 ;
  assign n8682 = \P1_reg2_reg[9]/NET0131  & ~n3718 ;
  assign n8667 = n3466 & n8396 ;
  assign n8681 = n1239 & n1763 ;
  assign n8683 = ~n8667 & ~n8681 ;
  assign n8684 = ~n8682 & n8683 ;
  assign n8685 = ~n8677 & n8684 ;
  assign n8686 = ~n8671 & n8685 ;
  assign n8687 = ~n8674 & n8686 ;
  assign n8688 = ~n8680 & n8687 ;
  assign n8689 = n3450 & ~n8688 ;
  assign n8690 = ~n8666 & ~n8689 ;
  assign n8691 = \P1_state_reg[0]/NET0131  & ~n8690 ;
  assign n8692 = ~n8665 & ~n8691 ;
  assign n8693 = \P2_reg2_reg[23]/NET0131  & ~n1983 ;
  assign n8694 = \P2_reg2_reg[23]/NET0131  & n2024 ;
  assign n8695 = \P2_reg2_reg[23]/NET0131  & ~n3758 ;
  assign n8696 = n3758 & n8331 ;
  assign n8697 = ~n8695 & ~n8696 ;
  assign n8698 = ~n3177 & ~n8697 ;
  assign n8699 = n3758 & ~n8380 ;
  assign n8701 = n3758 & ~n8352 ;
  assign n8702 = ~n8695 & ~n8701 ;
  assign n8703 = n3411 & ~n8702 ;
  assign n8700 = n3084 & n3420 ;
  assign n8704 = ~n4382 & n7770 ;
  assign n8705 = \P2_reg2_reg[23]/NET0131  & ~n8704 ;
  assign n8706 = ~n8700 & ~n8705 ;
  assign n8707 = ~n8703 & n8706 ;
  assign n8708 = ~n8699 & n8707 ;
  assign n8709 = ~n8698 & n8708 ;
  assign n8710 = n2026 & ~n8709 ;
  assign n8711 = ~n8694 & ~n8710 ;
  assign n8712 = \P1_state_reg[0]/NET0131  & ~n8711 ;
  assign n8713 = ~n8693 & ~n8712 ;
  assign n8714 = \P2_reg2_reg[9]/NET0131  & ~n1983 ;
  assign n8715 = \P2_reg2_reg[9]/NET0131  & n2024 ;
  assign n8717 = \P2_reg2_reg[9]/NET0131  & ~n3758 ;
  assign n8718 = n3758 & n7248 ;
  assign n8719 = ~n8717 & ~n8718 ;
  assign n8720 = n3411 & ~n8719 ;
  assign n8721 = n3758 & ~n7254 ;
  assign n8722 = ~n8717 & ~n8721 ;
  assign n8723 = ~n3177 & ~n8722 ;
  assign n8724 = n3758 & n7260 ;
  assign n8725 = ~n8717 & ~n8724 ;
  assign n8726 = n3355 & ~n8725 ;
  assign n8727 = n3758 & n7266 ;
  assign n8728 = ~n8717 & ~n8727 ;
  assign n8729 = ~n3320 & ~n8728 ;
  assign n8731 = \P2_reg2_reg[9]/NET0131  & ~n3774 ;
  assign n8716 = n3758 & n8489 ;
  assign n8730 = n2760 & n3420 ;
  assign n8732 = ~n8716 & ~n8730 ;
  assign n8733 = ~n8731 & n8732 ;
  assign n8734 = ~n8729 & n8733 ;
  assign n8735 = ~n8726 & n8734 ;
  assign n8736 = ~n8723 & n8735 ;
  assign n8737 = ~n8720 & n8736 ;
  assign n8738 = n2026 & ~n8737 ;
  assign n8739 = ~n8715 & ~n8738 ;
  assign n8740 = \P1_state_reg[0]/NET0131  & ~n8739 ;
  assign n8741 = ~n8714 & ~n8740 ;
  assign n8742 = \P1_reg0_reg[13]/NET0131  & ~n3435 ;
  assign n8743 = \P1_reg0_reg[13]/NET0131  & n3448 ;
  assign n8745 = \P1_reg0_reg[13]/NET0131  & ~n4396 ;
  assign n8746 = n4396 & ~n7119 ;
  assign n8747 = ~n8745 & ~n8746 ;
  assign n8748 = ~n3677 & ~n8747 ;
  assign n8755 = n4396 & n7139 ;
  assign n8756 = ~n8745 & ~n8755 ;
  assign n8757 = n3712 & ~n8756 ;
  assign n8744 = n4396 & n8467 ;
  assign n8758 = \P1_reg0_reg[13]/NET0131  & ~n4493 ;
  assign n8759 = ~n8744 & ~n8758 ;
  assign n8760 = ~n8757 & n8759 ;
  assign n8761 = ~n8748 & n8760 ;
  assign n8749 = n4396 & n7125 ;
  assign n8750 = ~n8745 & ~n8749 ;
  assign n8751 = ~n3563 & ~n8750 ;
  assign n8752 = n4396 & n7134 ;
  assign n8753 = ~n8745 & ~n8752 ;
  assign n8754 = n1936 & ~n8753 ;
  assign n8762 = ~n8751 & ~n8754 ;
  assign n8763 = n8761 & n8762 ;
  assign n8764 = n3450 & ~n8763 ;
  assign n8765 = ~n8743 & ~n8764 ;
  assign n8766 = \P1_state_reg[0]/NET0131  & ~n8765 ;
  assign n8767 = ~n8742 & ~n8766 ;
  assign n8768 = \P1_reg0_reg[23]/NET0131  & ~n3435 ;
  assign n8769 = \P1_reg0_reg[23]/NET0131  & n3448 ;
  assign n8770 = \P1_reg0_reg[23]/NET0131  & ~n4396 ;
  assign n8774 = n4396 & ~n7435 ;
  assign n8775 = ~n8770 & ~n8774 ;
  assign n8776 = ~n3563 & ~n8775 ;
  assign n8771 = n4396 & ~n7422 ;
  assign n8772 = ~n8770 & ~n8771 ;
  assign n8773 = ~n3677 & ~n8772 ;
  assign n8779 = n4396 & n7444 ;
  assign n8780 = ~n8770 & ~n8779 ;
  assign n8781 = n1936 & ~n8780 ;
  assign n8777 = ~n7450 & ~n7653 ;
  assign n8778 = n4396 & ~n8777 ;
  assign n8782 = \P1_reg0_reg[23]/NET0131  & ~n4494 ;
  assign n8783 = ~n8778 & ~n8782 ;
  assign n8784 = ~n8781 & n8783 ;
  assign n8785 = ~n8773 & n8784 ;
  assign n8786 = ~n8776 & n8785 ;
  assign n8787 = n3450 & ~n8786 ;
  assign n8788 = ~n8769 & ~n8787 ;
  assign n8789 = \P1_state_reg[0]/NET0131  & ~n8788 ;
  assign n8790 = ~n8768 & ~n8789 ;
  assign n8791 = \P1_reg0_reg[9]/NET0131  & ~n3435 ;
  assign n8792 = \P1_reg0_reg[9]/NET0131  & n3448 ;
  assign n8794 = \P1_reg0_reg[9]/NET0131  & ~n4396 ;
  assign n8804 = n4396 & ~n7310 ;
  assign n8805 = ~n8794 & ~n8804 ;
  assign n8806 = n1936 & ~n8805 ;
  assign n8798 = n4396 & ~n7288 ;
  assign n8799 = ~n8794 & ~n8798 ;
  assign n8800 = ~n3677 & ~n8799 ;
  assign n8795 = n4396 & n7294 ;
  assign n8796 = ~n8794 & ~n8795 ;
  assign n8797 = ~n3563 & ~n8796 ;
  assign n8801 = n4396 & n7300 ;
  assign n8802 = ~n8794 & ~n8801 ;
  assign n8803 = n3712 & ~n8802 ;
  assign n8793 = n4396 & n8396 ;
  assign n8807 = \P1_reg0_reg[9]/NET0131  & ~n4493 ;
  assign n8808 = ~n8793 & ~n8807 ;
  assign n8809 = ~n8803 & n8808 ;
  assign n8810 = ~n8797 & n8809 ;
  assign n8811 = ~n8800 & n8810 ;
  assign n8812 = ~n8806 & n8811 ;
  assign n8813 = n3450 & ~n8812 ;
  assign n8814 = ~n8792 & ~n8813 ;
  assign n8815 = \P1_state_reg[0]/NET0131  & ~n8814 ;
  assign n8816 = ~n8791 & ~n8815 ;
  assign n8817 = \P1_reg1_reg[10]/NET0131  & ~n3435 ;
  assign n8818 = \P1_reg1_reg[10]/NET0131  & n3448 ;
  assign n8820 = \P1_reg1_reg[10]/NET0131  & ~n4532 ;
  assign n8821 = n4532 & n7092 ;
  assign n8822 = ~n8820 & ~n8821 ;
  assign n8823 = ~n3563 & ~n8822 ;
  assign n8830 = n4532 & n7097 ;
  assign n8831 = ~n8820 & ~n8830 ;
  assign n8832 = n3712 & ~n8831 ;
  assign n8819 = n4532 & n8423 ;
  assign n8833 = \P1_reg1_reg[10]/NET0131  & ~n4541 ;
  assign n8834 = ~n8819 & ~n8833 ;
  assign n8835 = ~n8832 & n8834 ;
  assign n8836 = ~n8823 & n8835 ;
  assign n8824 = n4532 & n7086 ;
  assign n8825 = ~n8820 & ~n8824 ;
  assign n8826 = n1936 & ~n8825 ;
  assign n8827 = n4532 & ~n7078 ;
  assign n8828 = ~n8820 & ~n8827 ;
  assign n8829 = ~n3677 & ~n8828 ;
  assign n8837 = ~n8826 & ~n8829 ;
  assign n8838 = n8836 & n8837 ;
  assign n8839 = n3450 & ~n8838 ;
  assign n8840 = ~n8818 & ~n8839 ;
  assign n8841 = \P1_state_reg[0]/NET0131  & ~n8840 ;
  assign n8842 = ~n8817 & ~n8841 ;
  assign n8843 = \P1_reg1_reg[13]/NET0131  & ~n3435 ;
  assign n8844 = \P1_reg1_reg[13]/NET0131  & n3448 ;
  assign n8846 = \P1_reg1_reg[13]/NET0131  & ~n4532 ;
  assign n8847 = n4532 & ~n7119 ;
  assign n8848 = ~n8846 & ~n8847 ;
  assign n8849 = ~n3677 & ~n8848 ;
  assign n8856 = n4532 & n7139 ;
  assign n8857 = ~n8846 & ~n8856 ;
  assign n8858 = n3712 & ~n8857 ;
  assign n8845 = n4532 & n8467 ;
  assign n8859 = \P1_reg1_reg[13]/NET0131  & ~n4541 ;
  assign n8860 = ~n8845 & ~n8859 ;
  assign n8861 = ~n8858 & n8860 ;
  assign n8862 = ~n8849 & n8861 ;
  assign n8850 = n4532 & n7125 ;
  assign n8851 = ~n8846 & ~n8850 ;
  assign n8852 = ~n3563 & ~n8851 ;
  assign n8853 = n4532 & n7134 ;
  assign n8854 = ~n8846 & ~n8853 ;
  assign n8855 = n1936 & ~n8854 ;
  assign n8863 = ~n8852 & ~n8855 ;
  assign n8864 = n8862 & n8863 ;
  assign n8865 = n3450 & ~n8864 ;
  assign n8866 = ~n8844 & ~n8865 ;
  assign n8867 = \P1_state_reg[0]/NET0131  & ~n8866 ;
  assign n8868 = ~n8843 & ~n8867 ;
  assign n8869 = \P2_reg0_reg[10]/NET0131  & ~n1983 ;
  assign n8870 = \P2_reg0_reg[10]/NET0131  & n2024 ;
  assign n8872 = \P2_reg0_reg[10]/NET0131  & ~n2040 ;
  assign n8873 = n2040 & n7163 ;
  assign n8874 = ~n8872 & ~n8873 ;
  assign n8875 = n3411 & ~n8874 ;
  assign n8879 = n2040 & n7175 ;
  assign n8880 = ~n8872 & ~n8879 ;
  assign n8881 = ~n3320 & ~n8880 ;
  assign n8876 = n2040 & ~n7169 ;
  assign n8877 = ~n8872 & ~n8876 ;
  assign n8878 = ~n3177 & ~n8877 ;
  assign n8882 = n2040 & n7181 ;
  assign n8883 = ~n8872 & ~n8882 ;
  assign n8884 = n3355 & ~n8883 ;
  assign n8871 = \P2_reg0_reg[10]/NET0131  & ~n3423 ;
  assign n8885 = n2040 & n8503 ;
  assign n8886 = ~n8871 & ~n8885 ;
  assign n8887 = ~n8884 & n8886 ;
  assign n8888 = ~n8878 & n8887 ;
  assign n8889 = ~n8881 & n8888 ;
  assign n8890 = ~n8875 & n8889 ;
  assign n8891 = n2026 & ~n8890 ;
  assign n8892 = ~n8870 & ~n8891 ;
  assign n8893 = \P1_state_reg[0]/NET0131  & ~n8892 ;
  assign n8894 = ~n8869 & ~n8893 ;
  assign n8895 = \P2_reg0_reg[13]/NET0131  & ~n1983 ;
  assign n8896 = \P2_reg0_reg[13]/NET0131  & n2024 ;
  assign n8898 = \P2_reg0_reg[13]/NET0131  & ~n2040 ;
  assign n8899 = n2040 & ~n7205 ;
  assign n8900 = ~n8898 & ~n8899 ;
  assign n8901 = n3411 & ~n8900 ;
  assign n8903 = n2040 & n7211 ;
  assign n8904 = ~n8898 & ~n8903 ;
  assign n8905 = ~n3177 & ~n8904 ;
  assign n8897 = n2040 & ~n8540 ;
  assign n8902 = \P2_reg0_reg[13]/NET0131  & ~n8385 ;
  assign n8906 = ~n8897 & ~n8902 ;
  assign n8907 = ~n8905 & n8906 ;
  assign n8908 = ~n8901 & n8907 ;
  assign n8909 = n2026 & ~n8908 ;
  assign n8910 = ~n8896 & ~n8909 ;
  assign n8911 = \P1_state_reg[0]/NET0131  & ~n8910 ;
  assign n8912 = ~n8895 & ~n8911 ;
  assign n8913 = \P1_reg1_reg[23]/NET0131  & ~n3435 ;
  assign n8914 = \P1_reg1_reg[23]/NET0131  & n3448 ;
  assign n8915 = \P1_reg1_reg[23]/NET0131  & ~n4532 ;
  assign n8919 = n4532 & ~n7435 ;
  assign n8920 = ~n8915 & ~n8919 ;
  assign n8921 = ~n3563 & ~n8920 ;
  assign n8916 = n4532 & ~n7422 ;
  assign n8917 = ~n8915 & ~n8916 ;
  assign n8918 = ~n3677 & ~n8917 ;
  assign n8923 = n4532 & n7444 ;
  assign n8924 = ~n8915 & ~n8923 ;
  assign n8925 = n1936 & ~n8924 ;
  assign n8922 = n4532 & ~n8777 ;
  assign n8926 = \P1_reg1_reg[23]/NET0131  & ~n4573 ;
  assign n8927 = ~n8922 & ~n8926 ;
  assign n8928 = ~n8925 & n8927 ;
  assign n8929 = ~n8918 & n8928 ;
  assign n8930 = ~n8921 & n8929 ;
  assign n8931 = n3450 & ~n8930 ;
  assign n8932 = ~n8914 & ~n8931 ;
  assign n8933 = \P1_state_reg[0]/NET0131  & ~n8932 ;
  assign n8934 = ~n8913 & ~n8933 ;
  assign n8937 = n2024 & n2635 ;
  assign n8939 = n2635 & ~n3788 ;
  assign n8940 = n2058 & ~n2616 ;
  assign n8941 = ~n2642 & n3376 ;
  assign n8942 = n2531 & ~n8941 ;
  assign n8943 = ~n2058 & ~n3378 ;
  assign n8944 = ~n8942 & n8943 ;
  assign n8945 = ~n8940 & ~n8944 ;
  assign n8946 = n3788 & ~n8945 ;
  assign n8947 = ~n8939 & ~n8946 ;
  assign n8948 = n3411 & ~n8947 ;
  assign n8955 = n3823 & ~n4206 ;
  assign n8956 = ~n3823 & n4206 ;
  assign n8957 = ~n8955 & ~n8956 ;
  assign n8958 = n3788 & ~n8957 ;
  assign n8959 = ~n8939 & ~n8958 ;
  assign n8960 = ~n3320 & ~n8959 ;
  assign n8949 = n3880 & ~n4206 ;
  assign n8950 = ~n3880 & n4206 ;
  assign n8951 = ~n8949 & ~n8950 ;
  assign n8952 = n3788 & n8951 ;
  assign n8953 = ~n8939 & ~n8952 ;
  assign n8954 = ~n3177 & ~n8953 ;
  assign n8961 = ~n2656 & ~n3328 ;
  assign n8962 = ~n3329 & ~n8961 ;
  assign n8963 = n3788 & n8962 ;
  assign n8964 = ~n8939 & ~n8963 ;
  assign n8965 = n3355 & ~n8964 ;
  assign n8938 = ~n2656 & ~n3965 ;
  assign n8966 = n2635 & ~n3962 ;
  assign n8967 = ~n8938 & ~n8966 ;
  assign n8968 = ~n8965 & n8967 ;
  assign n8969 = ~n8954 & n8968 ;
  assign n8970 = ~n8960 & n8969 ;
  assign n8971 = ~n8948 & n8970 ;
  assign n8972 = n2026 & ~n8971 ;
  assign n8973 = ~n8937 & ~n8972 ;
  assign n8974 = \P1_state_reg[0]/NET0131  & ~n8973 ;
  assign n8935 = ~\P1_state_reg[0]/NET0131  & \P2_reg3_reg[4]/NET0131  ;
  assign n8936 = n2635 & n3976 ;
  assign n8975 = ~n8935 & ~n8936 ;
  assign n8976 = ~n8974 & n8975 ;
  assign n8978 = n2024 & n2526 ;
  assign n8980 = n2526 & ~n3788 ;
  assign n8981 = n2506 & ~n3378 ;
  assign n8982 = ~n3379 & ~n8981 ;
  assign n8983 = ~n2058 & ~n8982 ;
  assign n8984 = n2058 & n2642 ;
  assign n8985 = ~n8983 & ~n8984 ;
  assign n8986 = n3788 & n8985 ;
  assign n8987 = ~n8980 & ~n8986 ;
  assign n8988 = n3411 & ~n8987 ;
  assign n8989 = ~n2664 & n4194 ;
  assign n8990 = n2664 & ~n4194 ;
  assign n8991 = ~n8989 & ~n8990 ;
  assign n8992 = n3788 & ~n8991 ;
  assign n8993 = ~n8980 & ~n8992 ;
  assign n8994 = ~n3177 & ~n8993 ;
  assign n8995 = ~n2544 & ~n3329 ;
  assign n8996 = ~n3330 & n3355 ;
  assign n8997 = ~n8995 & n8996 ;
  assign n8999 = ~n3271 & n4194 ;
  assign n8998 = n3271 & ~n4194 ;
  assign n9000 = ~n3320 & ~n8998 ;
  assign n9001 = ~n8999 & n9000 ;
  assign n9002 = ~n8997 & ~n9001 ;
  assign n9003 = n3788 & ~n9002 ;
  assign n8979 = ~n2544 & ~n3965 ;
  assign n9004 = n5698 & ~n6311 ;
  assign n9005 = n2526 & ~n9004 ;
  assign n9006 = ~n8979 & ~n9005 ;
  assign n9007 = ~n9003 & n9006 ;
  assign n9008 = ~n8994 & n9007 ;
  assign n9009 = ~n8988 & n9008 ;
  assign n9010 = n2026 & ~n9009 ;
  assign n9011 = ~n8978 & ~n9010 ;
  assign n9012 = \P1_state_reg[0]/NET0131  & ~n9011 ;
  assign n8977 = ~\P1_state_reg[0]/NET0131  & \P2_reg3_reg[5]/NET0131  ;
  assign n9013 = n2526 & n3976 ;
  assign n9014 = ~n8977 & ~n9013 ;
  assign n9015 = ~n9012 & n9014 ;
  assign n9018 = n1568 & n3448 ;
  assign n9020 = n1568 & ~n3980 ;
  assign n9021 = n537 & ~n1617 ;
  assign n9022 = ~n1572 & n3573 ;
  assign n9023 = n1548 & ~n9022 ;
  assign n9024 = ~n537 & ~n3575 ;
  assign n9025 = ~n9023 & n9024 ;
  assign n9026 = ~n9021 & ~n9025 ;
  assign n9027 = n3980 & ~n9026 ;
  assign n9028 = ~n9020 & ~n9027 ;
  assign n9029 = n1936 & ~n9028 ;
  assign n9036 = ~n1680 & n1806 ;
  assign n9037 = n1680 & ~n1806 ;
  assign n9038 = ~n9036 & ~n9037 ;
  assign n9039 = n3980 & n9038 ;
  assign n9040 = ~n9020 & ~n9039 ;
  assign n9041 = ~n3677 & ~n9040 ;
  assign n9030 = n1806 & ~n3986 ;
  assign n9031 = ~n1806 & n3986 ;
  assign n9032 = ~n9030 & ~n9031 ;
  assign n9033 = n3980 & ~n9032 ;
  assign n9034 = ~n9020 & ~n9033 ;
  assign n9035 = ~n3563 & ~n9034 ;
  assign n9042 = ~n1586 & ~n3681 ;
  assign n9043 = ~n3682 & ~n9042 ;
  assign n9044 = n3980 & n9043 ;
  assign n9045 = ~n9020 & ~n9044 ;
  assign n9046 = n3712 & ~n9045 ;
  assign n9019 = ~n1586 & ~n4067 ;
  assign n9047 = n1568 & ~n4064 ;
  assign n9048 = ~n9019 & ~n9047 ;
  assign n9049 = ~n9046 & n9048 ;
  assign n9050 = ~n9035 & n9049 ;
  assign n9051 = ~n9041 & n9050 ;
  assign n9052 = ~n9029 & n9051 ;
  assign n9053 = n3450 & ~n9052 ;
  assign n9054 = ~n9018 & ~n9053 ;
  assign n9055 = \P1_state_reg[0]/NET0131  & ~n9054 ;
  assign n9016 = \P1_reg3_reg[4]/NET0131  & ~\P1_state_reg[0]/NET0131  ;
  assign n9017 = n1568 & n1953 ;
  assign n9056 = ~n9016 & ~n9017 ;
  assign n9057 = ~n9055 & n9056 ;
  assign n9060 = n1543 & n3448 ;
  assign n9067 = n1543 & ~n3980 ;
  assign n9068 = n1524 & ~n3575 ;
  assign n9069 = ~n1524 & n3575 ;
  assign n9070 = ~n9068 & ~n9069 ;
  assign n9071 = ~n537 & ~n9070 ;
  assign n9072 = n537 & n1572 ;
  assign n9073 = ~n9071 & ~n9072 ;
  assign n9074 = n3980 & n9073 ;
  assign n9075 = ~n9067 & ~n9074 ;
  assign n9076 = n1936 & ~n9075 ;
  assign n9083 = n1805 & ~n3636 ;
  assign n9084 = ~n1805 & n3636 ;
  assign n9085 = ~n9083 & ~n9084 ;
  assign n9086 = n3980 & ~n9085 ;
  assign n9087 = ~n9067 & ~n9086 ;
  assign n9088 = ~n3677 & ~n9087 ;
  assign n9077 = n1805 & ~n3518 ;
  assign n9078 = ~n1805 & n3518 ;
  assign n9079 = ~n9077 & ~n9078 ;
  assign n9080 = n3980 & ~n9079 ;
  assign n9081 = ~n9067 & ~n9080 ;
  assign n9082 = ~n3563 & ~n9081 ;
  assign n9061 = ~n1562 & n1880 ;
  assign n9062 = ~n1562 & ~n3682 ;
  assign n9063 = ~n3683 & ~n9062 ;
  assign n9064 = n3712 & n9063 ;
  assign n9065 = ~n9061 & ~n9064 ;
  assign n9066 = n3980 & ~n9065 ;
  assign n9089 = ~n1562 & n1763 ;
  assign n9090 = ~n1761 & n1762 ;
  assign n9091 = ~n3980 & n9090 ;
  assign n9092 = ~n3716 & ~n9091 ;
  assign n9093 = n1543 & ~n9092 ;
  assign n9094 = ~n9089 & ~n9093 ;
  assign n9095 = ~n9066 & n9094 ;
  assign n9096 = ~n9082 & n9095 ;
  assign n9097 = ~n9088 & n9096 ;
  assign n9098 = ~n9076 & n9097 ;
  assign n9099 = n3450 & ~n9098 ;
  assign n9100 = ~n9060 & ~n9099 ;
  assign n9101 = \P1_state_reg[0]/NET0131  & ~n9100 ;
  assign n9058 = \P1_reg3_reg[5]/NET0131  & ~\P1_state_reg[0]/NET0131  ;
  assign n9059 = n1543 & n1953 ;
  assign n9102 = ~n9058 & ~n9059 ;
  assign n9103 = ~n9101 & n9102 ;
  assign n9104 = \P1_reg1_reg[4]/NET0131  & ~n3435 ;
  assign n9105 = \P1_reg1_reg[4]/NET0131  & n3448 ;
  assign n9108 = \P1_reg1_reg[4]/NET0131  & ~n4532 ;
  assign n9109 = n4532 & ~n9026 ;
  assign n9110 = ~n9108 & ~n9109 ;
  assign n9111 = n1936 & ~n9110 ;
  assign n9115 = n4532 & n9038 ;
  assign n9116 = ~n9108 & ~n9115 ;
  assign n9117 = ~n3677 & ~n9116 ;
  assign n9112 = n4532 & ~n9032 ;
  assign n9113 = ~n9108 & ~n9112 ;
  assign n9114 = ~n3563 & ~n9113 ;
  assign n9118 = n4532 & n9043 ;
  assign n9119 = ~n9108 & ~n9118 ;
  assign n9120 = n3712 & ~n9119 ;
  assign n9106 = ~n1586 & n1880 ;
  assign n9107 = n4532 & n9106 ;
  assign n9121 = \P1_reg1_reg[4]/NET0131  & ~n4541 ;
  assign n9122 = ~n9107 & ~n9121 ;
  assign n9123 = ~n9120 & n9122 ;
  assign n9124 = ~n9114 & n9123 ;
  assign n9125 = ~n9117 & n9124 ;
  assign n9126 = ~n9111 & n9125 ;
  assign n9127 = n3450 & ~n9126 ;
  assign n9128 = ~n9105 & ~n9127 ;
  assign n9129 = \P1_state_reg[0]/NET0131  & ~n9128 ;
  assign n9130 = ~n9104 & ~n9129 ;
  assign n9131 = \P1_reg0_reg[4]/NET0131  & ~n3435 ;
  assign n9132 = \P1_reg0_reg[4]/NET0131  & n3448 ;
  assign n9134 = \P1_reg0_reg[4]/NET0131  & ~n4396 ;
  assign n9135 = n4396 & ~n9026 ;
  assign n9136 = ~n9134 & ~n9135 ;
  assign n9137 = n1936 & ~n9136 ;
  assign n9141 = n4396 & n9038 ;
  assign n9142 = ~n9134 & ~n9141 ;
  assign n9143 = ~n3677 & ~n9142 ;
  assign n9138 = n4396 & ~n9032 ;
  assign n9139 = ~n9134 & ~n9138 ;
  assign n9140 = ~n3563 & ~n9139 ;
  assign n9144 = n4396 & n9043 ;
  assign n9145 = ~n9134 & ~n9144 ;
  assign n9146 = n3712 & ~n9145 ;
  assign n9133 = n4396 & n9106 ;
  assign n9147 = \P1_reg0_reg[4]/NET0131  & ~n4493 ;
  assign n9148 = ~n9133 & ~n9147 ;
  assign n9149 = ~n9146 & n9148 ;
  assign n9150 = ~n9140 & n9149 ;
  assign n9151 = ~n9143 & n9150 ;
  assign n9152 = ~n9137 & n9151 ;
  assign n9153 = n3450 & ~n9152 ;
  assign n9154 = ~n9132 & ~n9153 ;
  assign n9155 = \P1_state_reg[0]/NET0131  & ~n9154 ;
  assign n9156 = ~n9131 & ~n9155 ;
  assign n9157 = \P2_reg0_reg[4]/NET0131  & ~n1983 ;
  assign n9158 = \P2_reg0_reg[4]/NET0131  & n2024 ;
  assign n9161 = \P2_reg0_reg[4]/NET0131  & ~n2040 ;
  assign n9162 = n2040 & ~n8945 ;
  assign n9163 = ~n9161 & ~n9162 ;
  assign n9164 = n3411 & ~n9163 ;
  assign n9168 = n2040 & n8951 ;
  assign n9169 = ~n9161 & ~n9168 ;
  assign n9170 = ~n3177 & ~n9169 ;
  assign n9165 = n2040 & ~n8957 ;
  assign n9166 = ~n9161 & ~n9165 ;
  assign n9167 = ~n3320 & ~n9166 ;
  assign n9171 = n2040 & n8962 ;
  assign n9172 = ~n9161 & ~n9171 ;
  assign n9173 = n3355 & ~n9172 ;
  assign n9159 = ~n2656 & n3358 ;
  assign n9160 = n2040 & n9159 ;
  assign n9174 = \P2_reg0_reg[4]/NET0131  & ~n3423 ;
  assign n9175 = ~n9160 & ~n9174 ;
  assign n9176 = ~n9173 & n9175 ;
  assign n9177 = ~n9167 & n9176 ;
  assign n9178 = ~n9170 & n9177 ;
  assign n9179 = ~n9164 & n9178 ;
  assign n9180 = n2026 & ~n9179 ;
  assign n9181 = ~n9158 & ~n9180 ;
  assign n9182 = \P1_state_reg[0]/NET0131  & ~n9181 ;
  assign n9183 = ~n9157 & ~n9182 ;
  assign n9184 = \P2_reg1_reg[4]/NET0131  & ~n1983 ;
  assign n9185 = \P2_reg1_reg[4]/NET0131  & n2024 ;
  assign n9187 = \P2_reg1_reg[4]/NET0131  & ~n3733 ;
  assign n9188 = n3733 & ~n8945 ;
  assign n9189 = ~n9187 & ~n9188 ;
  assign n9190 = n3411 & ~n9189 ;
  assign n9194 = n3733 & ~n8957 ;
  assign n9195 = ~n9187 & ~n9194 ;
  assign n9196 = ~n3320 & ~n9195 ;
  assign n9191 = n3733 & n8951 ;
  assign n9192 = ~n9187 & ~n9191 ;
  assign n9193 = ~n3177 & ~n9192 ;
  assign n9197 = n3733 & n8962 ;
  assign n9198 = ~n9187 & ~n9197 ;
  assign n9199 = n3355 & ~n9198 ;
  assign n9186 = n3733 & n9159 ;
  assign n9200 = \P2_reg1_reg[4]/NET0131  & ~n3743 ;
  assign n9201 = ~n9186 & ~n9200 ;
  assign n9202 = ~n9199 & n9201 ;
  assign n9203 = ~n9193 & n9202 ;
  assign n9204 = ~n9196 & n9203 ;
  assign n9205 = ~n9190 & n9204 ;
  assign n9206 = n2026 & ~n9205 ;
  assign n9207 = ~n9185 & ~n9206 ;
  assign n9208 = \P1_state_reg[0]/NET0131  & ~n9207 ;
  assign n9209 = ~n9184 & ~n9208 ;
  assign n9210 = \P1_reg2_reg[8]/NET0131  & ~n3435 ;
  assign n9211 = \P1_reg2_reg[8]/NET0131  & n3448 ;
  assign n9214 = \P1_reg2_reg[8]/NET0131  & ~n3466 ;
  assign n9215 = n3466 & n8292 ;
  assign n9216 = ~n9214 & ~n9215 ;
  assign n9217 = n1936 & ~n9216 ;
  assign n9221 = n3466 & ~n8304 ;
  assign n9222 = ~n9214 & ~n9221 ;
  assign n9223 = ~n3677 & ~n9222 ;
  assign n9218 = n3466 & n8298 ;
  assign n9219 = ~n9214 & ~n9218 ;
  assign n9220 = ~n3563 & ~n9219 ;
  assign n9224 = n3466 & n8310 ;
  assign n9225 = ~n9214 & ~n9224 ;
  assign n9226 = n3712 & ~n9225 ;
  assign n9228 = \P1_reg2_reg[8]/NET0131  & ~n3718 ;
  assign n9212 = n1281 & n1880 ;
  assign n9213 = n3466 & n9212 ;
  assign n9227 = n1262 & n1763 ;
  assign n9229 = ~n9213 & ~n9227 ;
  assign n9230 = ~n9228 & n9229 ;
  assign n9231 = ~n9226 & n9230 ;
  assign n9232 = ~n9220 & n9231 ;
  assign n9233 = ~n9223 & n9232 ;
  assign n9234 = ~n9217 & n9233 ;
  assign n9235 = n3450 & ~n9234 ;
  assign n9236 = ~n9211 & ~n9235 ;
  assign n9237 = \P1_state_reg[0]/NET0131  & ~n9236 ;
  assign n9238 = ~n9210 & ~n9237 ;
  assign n9239 = \P1_reg1_reg[8]/NET0131  & ~n3435 ;
  assign n9240 = \P1_reg1_reg[8]/NET0131  & n3448 ;
  assign n9242 = \P1_reg1_reg[8]/NET0131  & ~n4532 ;
  assign n9243 = n4532 & n8292 ;
  assign n9244 = ~n9242 & ~n9243 ;
  assign n9245 = n1936 & ~n9244 ;
  assign n9249 = n4532 & n8298 ;
  assign n9250 = ~n9242 & ~n9249 ;
  assign n9251 = ~n3563 & ~n9250 ;
  assign n9246 = n4532 & ~n8304 ;
  assign n9247 = ~n9242 & ~n9246 ;
  assign n9248 = ~n3677 & ~n9247 ;
  assign n9252 = n4532 & n8310 ;
  assign n9253 = ~n9242 & ~n9252 ;
  assign n9254 = n3712 & ~n9253 ;
  assign n9241 = n4532 & n9212 ;
  assign n9255 = \P1_reg1_reg[8]/NET0131  & ~n4541 ;
  assign n9256 = ~n9241 & ~n9255 ;
  assign n9257 = ~n9254 & n9256 ;
  assign n9258 = ~n9248 & n9257 ;
  assign n9259 = ~n9251 & n9258 ;
  assign n9260 = ~n9245 & n9259 ;
  assign n9261 = n3450 & ~n9260 ;
  assign n9262 = ~n9240 & ~n9261 ;
  assign n9263 = \P1_state_reg[0]/NET0131  & ~n9262 ;
  assign n9264 = ~n9239 & ~n9263 ;
  assign n9265 = \P1_reg2_reg[11]/NET0131  & ~n3435 ;
  assign n9266 = \P1_reg2_reg[11]/NET0131  & n3448 ;
  assign n9268 = \P1_reg2_reg[11]/NET0131  & ~n3466 ;
  assign n9269 = n3466 & n8010 ;
  assign n9270 = ~n9268 & ~n9269 ;
  assign n9271 = ~n3563 & ~n9270 ;
  assign n9278 = n1198 & n1880 ;
  assign n9279 = ~n8024 & ~n9278 ;
  assign n9280 = n3466 & ~n9279 ;
  assign n9267 = \P1_reg2_reg[11]/NET0131  & ~n5914 ;
  assign n9281 = n1203 & n1763 ;
  assign n9282 = ~n9267 & ~n9281 ;
  assign n9283 = ~n9280 & n9282 ;
  assign n9284 = ~n9271 & n9283 ;
  assign n9272 = n3466 & n8018 ;
  assign n9273 = ~n9268 & ~n9272 ;
  assign n9274 = n1936 & ~n9273 ;
  assign n9275 = n3466 & ~n8004 ;
  assign n9276 = ~n9268 & ~n9275 ;
  assign n9277 = ~n3677 & ~n9276 ;
  assign n9285 = ~n9274 & ~n9277 ;
  assign n9286 = n9284 & n9285 ;
  assign n9287 = n3450 & ~n9286 ;
  assign n9288 = ~n9266 & ~n9287 ;
  assign n9289 = \P1_state_reg[0]/NET0131  & ~n9288 ;
  assign n9290 = ~n9265 & ~n9289 ;
  assign n9291 = \P1_reg2_reg[14]/NET0131  & ~n3435 ;
  assign n9292 = \P1_reg2_reg[14]/NET0131  & n3448 ;
  assign n9294 = \P1_reg2_reg[14]/NET0131  & ~n3466 ;
  assign n9298 = n3466 & ~n8058 ;
  assign n9299 = ~n9294 & ~n9298 ;
  assign n9300 = ~n3466 & ~n3563 ;
  assign n9301 = n8062 & ~n9300 ;
  assign n9302 = ~n9299 & ~n9301 ;
  assign n9295 = n3466 & ~n8047 ;
  assign n9296 = ~n9294 & ~n9295 ;
  assign n9297 = n1936 & ~n9296 ;
  assign n9303 = n3466 & n8067 ;
  assign n9304 = ~n9294 & ~n9303 ;
  assign n9305 = n3712 & ~n9304 ;
  assign n9293 = \P1_reg2_reg[14]/NET0131  & ~n3718 ;
  assign n9306 = n1113 & n1763 ;
  assign n9307 = n1109 & n1880 ;
  assign n9308 = n3466 & n9307 ;
  assign n9309 = ~n9306 & ~n9308 ;
  assign n9310 = ~n9293 & n9309 ;
  assign n9311 = ~n9305 & n9310 ;
  assign n9312 = ~n9297 & n9311 ;
  assign n9313 = ~n9302 & n9312 ;
  assign n9314 = n3450 & ~n9313 ;
  assign n9315 = ~n9292 & ~n9314 ;
  assign n9316 = \P1_state_reg[0]/NET0131  & ~n9315 ;
  assign n9317 = ~n9291 & ~n9316 ;
  assign n9318 = \P1_reg2_reg[15]/NET0131  & ~n3435 ;
  assign n9319 = \P1_reg2_reg[15]/NET0131  & n3448 ;
  assign n9321 = \P1_reg2_reg[15]/NET0131  & ~n3466 ;
  assign n9322 = n3466 & n8094 ;
  assign n9323 = ~n9321 & ~n9322 ;
  assign n9324 = ~n3563 & ~n9323 ;
  assign n9331 = n1083 & n1880 ;
  assign n9332 = ~n8108 & ~n9331 ;
  assign n9333 = n3466 & ~n9332 ;
  assign n9320 = \P1_reg2_reg[15]/NET0131  & ~n5914 ;
  assign n9334 = n1088 & n1763 ;
  assign n9335 = ~n9320 & ~n9334 ;
  assign n9336 = ~n9333 & n9335 ;
  assign n9337 = ~n9324 & n9336 ;
  assign n9325 = n3466 & n8102 ;
  assign n9326 = ~n9321 & ~n9325 ;
  assign n9327 = n1936 & ~n9326 ;
  assign n9328 = n3466 & ~n8088 ;
  assign n9329 = ~n9321 & ~n9328 ;
  assign n9330 = ~n3677 & ~n9329 ;
  assign n9338 = ~n9327 & ~n9330 ;
  assign n9339 = n9337 & n9338 ;
  assign n9340 = n3450 & ~n9339 ;
  assign n9341 = ~n9319 & ~n9340 ;
  assign n9342 = \P1_state_reg[0]/NET0131  & ~n9341 ;
  assign n9343 = ~n9318 & ~n9342 ;
  assign n9344 = n3411 & n8252 ;
  assign n9347 = ~n3177 & n8258 ;
  assign n9346 = ~n3320 & ~n8264 ;
  assign n9345 = n2470 & n3358 ;
  assign n9348 = ~n8270 & ~n9345 ;
  assign n9349 = ~n9346 & n9348 ;
  assign n9350 = ~n9347 & n9349 ;
  assign n9351 = ~n9344 & n9350 ;
  assign n9352 = n5860 & ~n9351 ;
  assign n9353 = n7510 & n8385 ;
  assign n9354 = ~n9344 & n9353 ;
  assign n9355 = \P2_reg0_reg[8]/NET0131  & ~n9354 ;
  assign n9356 = ~n9352 & ~n9355 ;
  assign n9357 = \P2_reg1_reg[15]/NET0131  & ~n1983 ;
  assign n9358 = \P2_reg1_reg[15]/NET0131  & n2024 ;
  assign n9363 = \P2_reg1_reg[15]/NET0131  & ~n3733 ;
  assign n9367 = n3733 & n8217 ;
  assign n9368 = ~n9363 & ~n9367 ;
  assign n9369 = ~n3177 & ~n9368 ;
  assign n9364 = n3733 & n8211 ;
  assign n9365 = ~n9363 & ~n9364 ;
  assign n9366 = n3411 & ~n9365 ;
  assign n9370 = n3733 & n8222 ;
  assign n9371 = ~n9363 & ~n9370 ;
  assign n9372 = n3355 & ~n9371 ;
  assign n9359 = n2843 & n3358 ;
  assign n9360 = ~n3320 & ~n8228 ;
  assign n9361 = ~n9359 & ~n9360 ;
  assign n9362 = n3733 & ~n9361 ;
  assign n9373 = \P2_reg1_reg[15]/NET0131  & ~n8531 ;
  assign n9374 = ~n9362 & ~n9373 ;
  assign n9375 = ~n9372 & n9374 ;
  assign n9376 = ~n9366 & n9375 ;
  assign n9377 = ~n9369 & n9376 ;
  assign n9378 = n2026 & ~n9377 ;
  assign n9379 = ~n9358 & ~n9378 ;
  assign n9380 = \P1_state_reg[0]/NET0131  & ~n9379 ;
  assign n9381 = ~n9357 & ~n9380 ;
  assign n9382 = \P2_reg1_reg[8]/NET0131  & ~n1983 ;
  assign n9383 = \P2_reg1_reg[8]/NET0131  & n2024 ;
  assign n9384 = \P2_reg1_reg[8]/NET0131  & ~n8534 ;
  assign n9385 = n3733 & ~n9351 ;
  assign n9386 = ~n9384 & ~n9385 ;
  assign n9387 = n2026 & ~n9386 ;
  assign n9388 = ~n9383 & ~n9387 ;
  assign n9389 = \P1_state_reg[0]/NET0131  & ~n9388 ;
  assign n9390 = ~n9382 & ~n9389 ;
  assign n9391 = \P2_reg2_reg[11]/NET0131  & ~n1983 ;
  assign n9392 = \P2_reg2_reg[11]/NET0131  & n2024 ;
  assign n9394 = \P2_reg2_reg[11]/NET0131  & ~n3758 ;
  assign n9395 = n3758 & n8129 ;
  assign n9396 = ~n9394 & ~n9395 ;
  assign n9397 = n3411 & ~n9396 ;
  assign n9398 = n3758 & n8135 ;
  assign n9399 = ~n9394 & ~n9398 ;
  assign n9400 = ~n3177 & ~n9399 ;
  assign n9401 = n3758 & n8140 ;
  assign n9402 = ~n9394 & ~n9401 ;
  assign n9403 = n3355 & ~n9402 ;
  assign n9404 = n3758 & ~n8146 ;
  assign n9405 = ~n9394 & ~n9404 ;
  assign n9406 = ~n3320 & ~n9405 ;
  assign n9408 = n2704 & n3358 ;
  assign n9409 = n3758 & n9408 ;
  assign n9393 = \P2_reg2_reg[11]/NET0131  & ~n3774 ;
  assign n9407 = n2681 & n3420 ;
  assign n9410 = ~n9393 & ~n9407 ;
  assign n9411 = ~n9409 & n9410 ;
  assign n9412 = ~n9406 & n9411 ;
  assign n9413 = ~n9403 & n9412 ;
  assign n9414 = ~n9400 & n9413 ;
  assign n9415 = ~n9397 & n9414 ;
  assign n9416 = n2026 & ~n9415 ;
  assign n9417 = ~n9392 & ~n9416 ;
  assign n9418 = \P1_state_reg[0]/NET0131  & ~n9417 ;
  assign n9419 = ~n9391 & ~n9418 ;
  assign n9420 = \P2_reg2_reg[14]/NET0131  & ~n1983 ;
  assign n9421 = \P2_reg2_reg[14]/NET0131  & n2024 ;
  assign n9423 = \P2_reg2_reg[14]/NET0131  & ~n3758 ;
  assign n9424 = n3758 & n8171 ;
  assign n9425 = ~n9423 & ~n9424 ;
  assign n9426 = n3411 & ~n9425 ;
  assign n9437 = n2860 & n3358 ;
  assign n9438 = n3758 & n9437 ;
  assign n9422 = \P2_reg2_reg[14]/NET0131  & ~n3774 ;
  assign n9436 = n2866 & n3420 ;
  assign n9439 = ~n9422 & ~n9436 ;
  assign n9440 = ~n9438 & n9439 ;
  assign n9441 = ~n9426 & n9440 ;
  assign n9433 = n3758 & ~n8188 ;
  assign n9434 = ~n9423 & ~n9433 ;
  assign n9435 = ~n3320 & ~n9434 ;
  assign n9427 = n3758 & n8176 ;
  assign n9428 = ~n9423 & ~n9427 ;
  assign n9429 = n3355 & ~n9428 ;
  assign n9430 = n3758 & n8182 ;
  assign n9431 = ~n9423 & ~n9430 ;
  assign n9432 = ~n3177 & ~n9431 ;
  assign n9442 = ~n9429 & ~n9432 ;
  assign n9443 = ~n9435 & n9442 ;
  assign n9444 = n9441 & n9443 ;
  assign n9445 = n2026 & ~n9444 ;
  assign n9446 = ~n9421 & ~n9445 ;
  assign n9447 = \P1_state_reg[0]/NET0131  & ~n9446 ;
  assign n9448 = ~n9420 & ~n9447 ;
  assign n9449 = \P2_reg2_reg[8]/NET0131  & ~n1983 ;
  assign n9450 = \P2_reg2_reg[8]/NET0131  & n2024 ;
  assign n9452 = \P2_reg2_reg[8]/NET0131  & ~n3758 ;
  assign n9453 = n3758 & n8252 ;
  assign n9454 = ~n9452 & ~n9453 ;
  assign n9455 = n3411 & ~n9454 ;
  assign n9459 = n3758 & ~n8264 ;
  assign n9460 = ~n9452 & ~n9459 ;
  assign n9461 = ~n3320 & ~n9460 ;
  assign n9456 = n3758 & n8258 ;
  assign n9457 = ~n9452 & ~n9456 ;
  assign n9458 = ~n3177 & ~n9457 ;
  assign n9462 = n3758 & n8269 ;
  assign n9463 = ~n9452 & ~n9462 ;
  assign n9464 = n3355 & ~n9463 ;
  assign n9466 = \P2_reg2_reg[8]/NET0131  & ~n3774 ;
  assign n9451 = n3758 & n9345 ;
  assign n9465 = n2447 & n3420 ;
  assign n9467 = ~n9451 & ~n9465 ;
  assign n9468 = ~n9466 & n9467 ;
  assign n9469 = ~n9464 & n9468 ;
  assign n9470 = ~n9458 & n9469 ;
  assign n9471 = ~n9461 & n9470 ;
  assign n9472 = ~n9455 & n9471 ;
  assign n9473 = n2026 & ~n9472 ;
  assign n9474 = ~n9450 & ~n9473 ;
  assign n9475 = \P1_state_reg[0]/NET0131  & ~n9474 ;
  assign n9476 = ~n9449 & ~n9475 ;
  assign n9477 = \P1_reg0_reg[15]/NET0131  & ~n3435 ;
  assign n9478 = \P1_reg0_reg[15]/NET0131  & n3448 ;
  assign n9480 = \P1_reg0_reg[15]/NET0131  & ~n4396 ;
  assign n9481 = n4396 & n8094 ;
  assign n9482 = ~n9480 & ~n9481 ;
  assign n9483 = ~n3563 & ~n9482 ;
  assign n9479 = \P1_reg0_reg[15]/NET0131  & ~n4494 ;
  assign n9490 = n4396 & ~n9332 ;
  assign n9491 = ~n9479 & ~n9490 ;
  assign n9492 = ~n9483 & n9491 ;
  assign n9484 = n4396 & n8102 ;
  assign n9485 = ~n9480 & ~n9484 ;
  assign n9486 = n1936 & ~n9485 ;
  assign n9487 = n4396 & ~n8088 ;
  assign n9488 = ~n9480 & ~n9487 ;
  assign n9489 = ~n3677 & ~n9488 ;
  assign n9493 = ~n9486 & ~n9489 ;
  assign n9494 = n9492 & n9493 ;
  assign n9495 = n3450 & ~n9494 ;
  assign n9496 = ~n9478 & ~n9495 ;
  assign n9497 = \P1_state_reg[0]/NET0131  & ~n9496 ;
  assign n9498 = ~n9477 & ~n9497 ;
  assign n9499 = \P1_reg0_reg[8]/NET0131  & ~n3435 ;
  assign n9500 = \P1_reg0_reg[8]/NET0131  & n3448 ;
  assign n9502 = \P1_reg0_reg[8]/NET0131  & ~n4396 ;
  assign n9503 = n4396 & n8292 ;
  assign n9504 = ~n9502 & ~n9503 ;
  assign n9505 = n1936 & ~n9504 ;
  assign n9509 = n4396 & ~n8304 ;
  assign n9510 = ~n9502 & ~n9509 ;
  assign n9511 = ~n3677 & ~n9510 ;
  assign n9506 = n4396 & n8298 ;
  assign n9507 = ~n9502 & ~n9506 ;
  assign n9508 = ~n3563 & ~n9507 ;
  assign n9512 = n4396 & n8310 ;
  assign n9513 = ~n9502 & ~n9512 ;
  assign n9514 = n3712 & ~n9513 ;
  assign n9501 = n4396 & n9212 ;
  assign n9515 = \P1_reg0_reg[8]/NET0131  & ~n4493 ;
  assign n9516 = ~n9501 & ~n9515 ;
  assign n9517 = ~n9514 & n9516 ;
  assign n9518 = ~n9508 & n9517 ;
  assign n9519 = ~n9511 & n9518 ;
  assign n9520 = ~n9505 & n9519 ;
  assign n9521 = n3450 & ~n9520 ;
  assign n9522 = ~n9500 & ~n9521 ;
  assign n9523 = \P1_state_reg[0]/NET0131  & ~n9522 ;
  assign n9524 = ~n9499 & ~n9523 ;
  assign n9525 = \P1_reg1_reg[15]/NET0131  & ~n3435 ;
  assign n9526 = \P1_reg1_reg[15]/NET0131  & n3448 ;
  assign n9528 = \P1_reg1_reg[15]/NET0131  & ~n4532 ;
  assign n9529 = n4532 & n8094 ;
  assign n9530 = ~n9528 & ~n9529 ;
  assign n9531 = ~n3563 & ~n9530 ;
  assign n9538 = n4532 & n8107 ;
  assign n9539 = ~n9528 & ~n9538 ;
  assign n9540 = n3712 & ~n9539 ;
  assign n9527 = \P1_reg1_reg[15]/NET0131  & ~n4491 ;
  assign n9541 = n1083 & n4532 ;
  assign n9542 = ~n9528 & ~n9541 ;
  assign n9543 = n1880 & ~n9542 ;
  assign n9544 = ~n9527 & ~n9543 ;
  assign n9545 = ~n9540 & n9544 ;
  assign n9546 = ~n9531 & n9545 ;
  assign n9532 = n4532 & n8102 ;
  assign n9533 = ~n9528 & ~n9532 ;
  assign n9534 = n1936 & ~n9533 ;
  assign n9535 = n4532 & ~n8088 ;
  assign n9536 = ~n9528 & ~n9535 ;
  assign n9537 = ~n3677 & ~n9536 ;
  assign n9547 = ~n9534 & ~n9537 ;
  assign n9548 = n9546 & n9547 ;
  assign n9549 = n3450 & ~n9548 ;
  assign n9550 = ~n9526 & ~n9549 ;
  assign n9551 = \P1_state_reg[0]/NET0131  & ~n9550 ;
  assign n9552 = ~n9525 & ~n9551 ;
  assign n9553 = \P2_reg0_reg[15]/NET0131  & ~n1983 ;
  assign n9554 = \P2_reg0_reg[15]/NET0131  & n2024 ;
  assign n9556 = \P2_reg0_reg[15]/NET0131  & ~n2040 ;
  assign n9560 = n2040 & n8217 ;
  assign n9561 = ~n9556 & ~n9560 ;
  assign n9562 = ~n3177 & ~n9561 ;
  assign n9557 = n2040 & n8211 ;
  assign n9558 = ~n9556 & ~n9557 ;
  assign n9559 = n3411 & ~n9558 ;
  assign n9563 = n2040 & n8222 ;
  assign n9564 = ~n9556 & ~n9563 ;
  assign n9565 = n3355 & ~n9564 ;
  assign n9555 = n2040 & ~n9361 ;
  assign n9566 = \P2_reg0_reg[15]/NET0131  & ~n7506 ;
  assign n9567 = ~n9555 & ~n9566 ;
  assign n9568 = ~n9565 & n9567 ;
  assign n9569 = ~n9559 & n9568 ;
  assign n9570 = ~n9562 & n9569 ;
  assign n9571 = n2026 & ~n9570 ;
  assign n9572 = ~n9554 & ~n9571 ;
  assign n9573 = \P1_state_reg[0]/NET0131  & ~n9572 ;
  assign n9574 = ~n9553 & ~n9573 ;
  assign n9576 = ~\P2_reg3_reg[3]/NET0131  & n2024 ;
  assign n9593 = n2642 & ~n3376 ;
  assign n9594 = ~n8941 & ~n9593 ;
  assign n9595 = ~n2058 & ~n9594 ;
  assign n9596 = n2058 & n2552 ;
  assign n9597 = ~n9595 & ~n9596 ;
  assign n9598 = n3411 & n9597 ;
  assign n9578 = ~n3260 & ~n3261 ;
  assign n9579 = ~n4193 & n9578 ;
  assign n9580 = n4193 & ~n9578 ;
  assign n9581 = ~n9579 & ~n9580 ;
  assign n9582 = ~n3320 & ~n9581 ;
  assign n9577 = ~n2631 & n3358 ;
  assign n9583 = ~n2631 & ~n3327 ;
  assign n9584 = ~n3328 & n3355 ;
  assign n9585 = ~n9583 & n9584 ;
  assign n9586 = ~n9577 & ~n9585 ;
  assign n9587 = ~n9582 & n9586 ;
  assign n9588 = ~n2608 & ~n2609 ;
  assign n9589 = n4193 & n9588 ;
  assign n9590 = ~n4193 & ~n9588 ;
  assign n9591 = ~n9589 & ~n9590 ;
  assign n9592 = ~n3177 & ~n9591 ;
  assign n9599 = n9587 & ~n9592 ;
  assign n9600 = ~n9598 & n9599 ;
  assign n9601 = n3788 & ~n9600 ;
  assign n9604 = ~\P2_reg3_reg[3]/NET0131  & ~n3788 ;
  assign n9605 = ~n6641 & n9604 ;
  assign n9602 = ~\P2_reg3_reg[3]/NET0131  & n3417 ;
  assign n9603 = ~n2631 & n3420 ;
  assign n9606 = ~n9602 & ~n9603 ;
  assign n9607 = ~n9605 & n9606 ;
  assign n9608 = ~n9601 & n9607 ;
  assign n9609 = n2026 & ~n9608 ;
  assign n9610 = ~n9576 & ~n9609 ;
  assign n9611 = \P1_state_reg[0]/NET0131  & ~n9610 ;
  assign n9575 = ~\P1_state_reg[0]/NET0131  & \P2_reg3_reg[3]/NET0131  ;
  assign n9612 = ~\P2_reg3_reg[3]/NET0131  & n3976 ;
  assign n9613 = ~n9575 & ~n9612 ;
  assign n9614 = ~n9611 & n9613 ;
  assign n9617 = n2024 & n2499 ;
  assign n9619 = n2499 & ~n3788 ;
  assign n9620 = n2480 & ~n3379 ;
  assign n9621 = ~n3380 & ~n9620 ;
  assign n9622 = ~n2058 & ~n9621 ;
  assign n9623 = n2058 & n2531 ;
  assign n9624 = ~n9622 & ~n9623 ;
  assign n9625 = n3788 & n9624 ;
  assign n9626 = ~n9619 & ~n9625 ;
  assign n9627 = n3411 & ~n9626 ;
  assign n9634 = n3885 & ~n4205 ;
  assign n9635 = ~n3885 & n4205 ;
  assign n9636 = ~n9634 & ~n9635 ;
  assign n9637 = n3788 & n9636 ;
  assign n9638 = ~n9619 & ~n9637 ;
  assign n9639 = ~n3177 & ~n9638 ;
  assign n9628 = n3827 & ~n4205 ;
  assign n9629 = ~n3827 & n4205 ;
  assign n9630 = ~n9628 & ~n9629 ;
  assign n9631 = n3788 & ~n9630 ;
  assign n9632 = ~n9619 & ~n9631 ;
  assign n9633 = ~n3320 & ~n9632 ;
  assign n9640 = ~n2521 & ~n3330 ;
  assign n9641 = ~n3331 & ~n9640 ;
  assign n9642 = n3788 & n9641 ;
  assign n9643 = ~n9619 & ~n9642 ;
  assign n9644 = n3355 & ~n9643 ;
  assign n9618 = ~n2521 & ~n3965 ;
  assign n9645 = n2499 & ~n3962 ;
  assign n9646 = ~n9618 & ~n9645 ;
  assign n9647 = ~n9644 & n9646 ;
  assign n9648 = ~n9633 & n9647 ;
  assign n9649 = ~n9639 & n9648 ;
  assign n9650 = ~n9627 & n9649 ;
  assign n9651 = n2026 & ~n9650 ;
  assign n9652 = ~n9617 & ~n9651 ;
  assign n9653 = \P1_state_reg[0]/NET0131  & ~n9652 ;
  assign n9615 = ~\P1_state_reg[0]/NET0131  & \P2_reg3_reg[6]/NET0131  ;
  assign n9616 = n2499 & n3976 ;
  assign n9654 = ~n9615 & ~n9616 ;
  assign n9655 = ~n9653 & n9654 ;
  assign n9657 = n2024 & n2476 ;
  assign n9659 = n2476 & ~n3788 ;
  assign n9660 = n2454 & ~n3380 ;
  assign n9661 = ~n7242 & ~n9660 ;
  assign n9662 = ~n2058 & ~n9661 ;
  assign n9663 = n2058 & n2506 ;
  assign n9664 = ~n9662 & ~n9663 ;
  assign n9665 = n3788 & n9664 ;
  assign n9666 = ~n9659 & ~n9665 ;
  assign n9667 = n3411 & ~n9666 ;
  assign n9668 = n4207 & ~n4799 ;
  assign n9669 = ~n4207 & n4799 ;
  assign n9670 = ~n9668 & ~n9669 ;
  assign n9671 = n3788 & n9670 ;
  assign n9672 = ~n9659 & ~n9671 ;
  assign n9673 = ~n3177 & ~n9672 ;
  assign n9674 = n4207 & ~n4835 ;
  assign n9675 = ~n4207 & n4835 ;
  assign n9676 = ~n9674 & ~n9675 ;
  assign n9677 = n3788 & ~n9676 ;
  assign n9678 = ~n9659 & ~n9677 ;
  assign n9679 = ~n3320 & ~n9678 ;
  assign n9680 = n2495 & ~n3331 ;
  assign n9681 = ~n3332 & ~n9680 ;
  assign n9682 = n3355 & n9681 ;
  assign n9683 = n3788 & n9682 ;
  assign n9658 = n2476 & ~n5698 ;
  assign n9684 = n2495 & ~n3965 ;
  assign n9685 = ~n9658 & ~n9684 ;
  assign n9686 = ~n9683 & n9685 ;
  assign n9687 = ~n9679 & n9686 ;
  assign n9688 = ~n9673 & n9687 ;
  assign n9689 = ~n9667 & n9688 ;
  assign n9690 = n2026 & ~n9689 ;
  assign n9691 = ~n9657 & ~n9690 ;
  assign n9692 = \P1_state_reg[0]/NET0131  & ~n9691 ;
  assign n9656 = ~\P1_state_reg[0]/NET0131  & \P2_reg3_reg[7]/NET0131  ;
  assign n9693 = n2476 & n3976 ;
  assign n9694 = ~n9656 & ~n9693 ;
  assign n9695 = ~n9692 & n9694 ;
  assign n9697 = ~\P1_reg3_reg[3]/NET0131  & n3448 ;
  assign n9704 = ~\P1_reg3_reg[3]/NET0131  & ~n3980 ;
  assign n9705 = n1572 & ~n3573 ;
  assign n9706 = ~n9022 & ~n9705 ;
  assign n9707 = ~n537 & ~n9706 ;
  assign n9708 = n537 & n1595 ;
  assign n9709 = ~n9707 & ~n9708 ;
  assign n9710 = n3980 & n9709 ;
  assign n9711 = ~n9704 & ~n9710 ;
  assign n9712 = n1936 & ~n9711 ;
  assign n9713 = ~n1778 & ~n3508 ;
  assign n9714 = n1773 & n9713 ;
  assign n9715 = ~n1773 & ~n9713 ;
  assign n9716 = ~n9714 & ~n9715 ;
  assign n9717 = n3980 & ~n9716 ;
  assign n9718 = ~n9704 & ~n9717 ;
  assign n9719 = ~n3563 & ~n9718 ;
  assign n9720 = ~n1610 & ~n3633 ;
  assign n9721 = n1773 & n9720 ;
  assign n9722 = ~n1773 & ~n9720 ;
  assign n9723 = ~n9721 & ~n9722 ;
  assign n9724 = n3980 & n9723 ;
  assign n9725 = ~n9704 & ~n9724 ;
  assign n9726 = ~n3677 & ~n9725 ;
  assign n9698 = ~n1632 & n1880 ;
  assign n9699 = ~n1632 & ~n3680 ;
  assign n9700 = ~n3681 & n3712 ;
  assign n9701 = ~n9699 & n9700 ;
  assign n9702 = ~n9698 & ~n9701 ;
  assign n9703 = n3980 & ~n9702 ;
  assign n9727 = ~n1632 & n1763 ;
  assign n9728 = ~\P1_reg3_reg[3]/NET0131  & ~n9092 ;
  assign n9729 = ~n9727 & ~n9728 ;
  assign n9730 = ~n9703 & n9729 ;
  assign n9731 = ~n9726 & n9730 ;
  assign n9732 = ~n9719 & n9731 ;
  assign n9733 = ~n9712 & n9732 ;
  assign n9734 = n3450 & ~n9733 ;
  assign n9735 = ~n9697 & ~n9734 ;
  assign n9736 = \P1_state_reg[0]/NET0131  & ~n9735 ;
  assign n9696 = \P1_reg3_reg[3]/NET0131  & ~\P1_state_reg[0]/NET0131  ;
  assign n9737 = ~\P1_reg3_reg[3]/NET0131  & n1953 ;
  assign n9738 = ~n9696 & ~n9737 ;
  assign n9739 = ~n9736 & n9738 ;
  assign n9742 = n1518 & n3448 ;
  assign n9744 = n1518 & ~n3980 ;
  assign n9745 = n537 & ~n1548 ;
  assign n9746 = n1498 & ~n9069 ;
  assign n9747 = ~n537 & ~n3577 ;
  assign n9748 = ~n9746 & n9747 ;
  assign n9749 = ~n9745 & ~n9748 ;
  assign n9750 = n3980 & ~n9749 ;
  assign n9751 = ~n9744 & ~n9750 ;
  assign n9752 = n1936 & ~n9751 ;
  assign n9765 = ~n1537 & ~n3683 ;
  assign n9766 = ~n3684 & ~n9765 ;
  assign n9767 = n3980 & n9766 ;
  assign n9768 = ~n9744 & ~n9767 ;
  assign n9769 = n3712 & ~n9768 ;
  assign n9743 = ~n1537 & ~n4067 ;
  assign n9770 = n1518 & ~n4064 ;
  assign n9771 = ~n9743 & ~n9770 ;
  assign n9772 = ~n9769 & n9771 ;
  assign n9773 = ~n9752 & n9772 ;
  assign n9753 = ~n1686 & n1793 ;
  assign n9754 = n1686 & ~n1793 ;
  assign n9755 = ~n9753 & ~n9754 ;
  assign n9756 = n3980 & n9755 ;
  assign n9757 = ~n9744 & ~n9756 ;
  assign n9758 = ~n3677 & ~n9757 ;
  assign n9759 = n1793 & ~n5509 ;
  assign n9760 = ~n1793 & n5509 ;
  assign n9761 = ~n9759 & ~n9760 ;
  assign n9762 = n3980 & ~n9761 ;
  assign n9763 = ~n9744 & ~n9762 ;
  assign n9764 = ~n3563 & ~n9763 ;
  assign n9774 = ~n9758 & ~n9764 ;
  assign n9775 = n9773 & n9774 ;
  assign n9776 = n3450 & ~n9775 ;
  assign n9777 = ~n9742 & ~n9776 ;
  assign n9778 = \P1_state_reg[0]/NET0131  & ~n9777 ;
  assign n9740 = \P1_reg3_reg[6]/NET0131  & ~\P1_state_reg[0]/NET0131  ;
  assign n9741 = n1518 & n1953 ;
  assign n9779 = ~n9740 & ~n9741 ;
  assign n9780 = ~n9778 & n9779 ;
  assign n9783 = n1491 & n3448 ;
  assign n9785 = n1491 & ~n3980 ;
  assign n9786 = n1776 & ~n4399 ;
  assign n9787 = ~n1776 & n4399 ;
  assign n9788 = ~n9786 & ~n9787 ;
  assign n9789 = n3980 & ~n9788 ;
  assign n9790 = ~n9785 & ~n9789 ;
  assign n9791 = ~n3677 & ~n9790 ;
  assign n9806 = ~n1514 & ~n3684 ;
  assign n9807 = ~n8308 & ~n9806 ;
  assign n9808 = n3712 & n9807 ;
  assign n9809 = n3980 & n9808 ;
  assign n9784 = n1491 & ~n4910 ;
  assign n9810 = ~n1514 & ~n4067 ;
  assign n9811 = ~n9784 & ~n9810 ;
  assign n9812 = ~n9809 & n9811 ;
  assign n9813 = ~n9791 & n9812 ;
  assign n9792 = n1776 & ~n4442 ;
  assign n9793 = ~n1776 & n4442 ;
  assign n9794 = ~n9792 & ~n9793 ;
  assign n9795 = n3980 & n9794 ;
  assign n9796 = ~n9785 & ~n9795 ;
  assign n9797 = ~n3563 & ~n9796 ;
  assign n9798 = n1267 & ~n3577 ;
  assign n9799 = ~n7305 & ~n9798 ;
  assign n9800 = ~n537 & ~n9799 ;
  assign n9801 = n537 & n1524 ;
  assign n9802 = ~n9800 & ~n9801 ;
  assign n9803 = n3980 & n9802 ;
  assign n9804 = ~n9785 & ~n9803 ;
  assign n9805 = n1936 & ~n9804 ;
  assign n9814 = ~n9797 & ~n9805 ;
  assign n9815 = n9813 & n9814 ;
  assign n9816 = n3450 & ~n9815 ;
  assign n9817 = ~n9783 & ~n9816 ;
  assign n9818 = \P1_state_reg[0]/NET0131  & ~n9817 ;
  assign n9781 = \P1_reg3_reg[7]/NET0131  & ~\P1_state_reg[0]/NET0131  ;
  assign n9782 = n1491 & n1953 ;
  assign n9819 = ~n9781 & ~n9782 ;
  assign n9820 = ~n9818 & n9819 ;
  assign n9821 = \P1_reg1_reg[5]/NET0131  & ~n3435 ;
  assign n9822 = \P1_reg1_reg[5]/NET0131  & n3448 ;
  assign n9824 = \P1_reg1_reg[5]/NET0131  & ~n4532 ;
  assign n9825 = n4532 & n9073 ;
  assign n9826 = ~n9824 & ~n9825 ;
  assign n9827 = n1936 & ~n9826 ;
  assign n9831 = n4532 & ~n9085 ;
  assign n9832 = ~n9824 & ~n9831 ;
  assign n9833 = ~n3677 & ~n9832 ;
  assign n9828 = n4532 & ~n9079 ;
  assign n9829 = ~n9824 & ~n9828 ;
  assign n9830 = ~n3563 & ~n9829 ;
  assign n9823 = n4532 & ~n9065 ;
  assign n9834 = ~n4532 & n9090 ;
  assign n9835 = n4491 & ~n9834 ;
  assign n9836 = \P1_reg1_reg[5]/NET0131  & ~n9835 ;
  assign n9837 = ~n9823 & ~n9836 ;
  assign n9838 = ~n9830 & n9837 ;
  assign n9839 = ~n9833 & n9838 ;
  assign n9840 = ~n9827 & n9839 ;
  assign n9841 = n3450 & ~n9840 ;
  assign n9842 = ~n9822 & ~n9841 ;
  assign n9843 = \P1_state_reg[0]/NET0131  & ~n9842 ;
  assign n9844 = ~n9821 & ~n9843 ;
  assign n9845 = n3411 & n8985 ;
  assign n9846 = n9353 & ~n9845 ;
  assign n9847 = \P2_reg0_reg[5]/NET0131  & ~n9846 ;
  assign n9849 = ~n3177 & ~n8991 ;
  assign n9848 = ~n2544 & n3358 ;
  assign n9850 = n9002 & ~n9848 ;
  assign n9851 = ~n9849 & n9850 ;
  assign n9852 = ~n9845 & n9851 ;
  assign n9853 = n5860 & ~n9852 ;
  assign n9854 = ~n9847 & ~n9853 ;
  assign n9855 = \P2_reg1_reg[11]/NET0131  & ~n1983 ;
  assign n9856 = \P2_reg1_reg[11]/NET0131  & n2024 ;
  assign n9858 = \P2_reg1_reg[11]/NET0131  & ~n3733 ;
  assign n9859 = n3733 & n8129 ;
  assign n9860 = ~n9858 & ~n9859 ;
  assign n9861 = n3411 & ~n9860 ;
  assign n9862 = n3733 & n8135 ;
  assign n9863 = ~n9858 & ~n9862 ;
  assign n9864 = ~n3177 & ~n9863 ;
  assign n9857 = \P2_reg1_reg[11]/NET0131  & ~n8532 ;
  assign n9865 = n3355 & n8140 ;
  assign n9866 = ~n8147 & ~n9408 ;
  assign n9867 = ~n9865 & n9866 ;
  assign n9868 = n3733 & ~n9867 ;
  assign n9869 = ~n9857 & ~n9868 ;
  assign n9870 = ~n9864 & n9869 ;
  assign n9871 = ~n9861 & n9870 ;
  assign n9872 = n2026 & ~n9871 ;
  assign n9873 = ~n9856 & ~n9872 ;
  assign n9874 = \P1_state_reg[0]/NET0131  & ~n9873 ;
  assign n9875 = ~n9855 & ~n9874 ;
  assign n9876 = \P2_reg1_reg[14]/NET0131  & ~n1983 ;
  assign n9877 = \P2_reg1_reg[14]/NET0131  & n2024 ;
  assign n9880 = \P2_reg1_reg[14]/NET0131  & ~n3733 ;
  assign n9881 = n3733 & n8176 ;
  assign n9882 = ~n9880 & ~n9881 ;
  assign n9883 = n3355 & ~n9882 ;
  assign n9878 = n3733 & n9437 ;
  assign n9879 = \P2_reg1_reg[14]/NET0131  & ~n3743 ;
  assign n9893 = ~n9878 & ~n9879 ;
  assign n9894 = ~n9883 & n9893 ;
  assign n9890 = n3733 & n8171 ;
  assign n9891 = ~n9880 & ~n9890 ;
  assign n9892 = n3411 & ~n9891 ;
  assign n9884 = n3733 & n8182 ;
  assign n9885 = ~n9880 & ~n9884 ;
  assign n9886 = ~n3177 & ~n9885 ;
  assign n9887 = n3733 & ~n8188 ;
  assign n9888 = ~n9880 & ~n9887 ;
  assign n9889 = ~n3320 & ~n9888 ;
  assign n9895 = ~n9886 & ~n9889 ;
  assign n9896 = ~n9892 & n9895 ;
  assign n9897 = n9894 & n9896 ;
  assign n9898 = n2026 & ~n9897 ;
  assign n9899 = ~n9877 & ~n9898 ;
  assign n9900 = \P1_state_reg[0]/NET0131  & ~n9899 ;
  assign n9901 = ~n9876 & ~n9900 ;
  assign n9902 = n5964 & ~n9852 ;
  assign n9903 = n3357 & ~n3418 ;
  assign n9904 = n3320 & ~n9903 ;
  assign n9905 = ~n3733 & ~n9904 ;
  assign n9906 = n3421 & ~n9905 ;
  assign n9907 = n5287 & ~n8533 ;
  assign n9908 = n9906 & n9907 ;
  assign n9909 = \P2_reg1_reg[5]/NET0131  & ~n9908 ;
  assign n9910 = ~n9902 & ~n9909 ;
  assign n9911 = \P1_reg2_reg[4]/NET0131  & ~n3435 ;
  assign n9912 = \P1_reg2_reg[4]/NET0131  & n3448 ;
  assign n9914 = \P1_reg2_reg[4]/NET0131  & ~n3466 ;
  assign n9915 = n3466 & ~n9026 ;
  assign n9916 = ~n9914 & ~n9915 ;
  assign n9917 = n1936 & ~n9916 ;
  assign n9921 = n3466 & n9038 ;
  assign n9922 = ~n9914 & ~n9921 ;
  assign n9923 = ~n3677 & ~n9922 ;
  assign n9918 = n3466 & ~n9032 ;
  assign n9919 = ~n9914 & ~n9918 ;
  assign n9920 = ~n3563 & ~n9919 ;
  assign n9924 = n3466 & n9043 ;
  assign n9925 = ~n9914 & ~n9924 ;
  assign n9926 = n3712 & ~n9925 ;
  assign n9928 = \P1_reg2_reg[4]/NET0131  & ~n3718 ;
  assign n9913 = n3466 & n9106 ;
  assign n9927 = n1568 & n1763 ;
  assign n9929 = ~n9913 & ~n9927 ;
  assign n9930 = ~n9928 & n9929 ;
  assign n9931 = ~n9926 & n9930 ;
  assign n9932 = ~n9920 & n9931 ;
  assign n9933 = ~n9923 & n9932 ;
  assign n9934 = ~n9917 & n9933 ;
  assign n9935 = n3450 & ~n9934 ;
  assign n9936 = ~n9912 & ~n9935 ;
  assign n9937 = \P1_state_reg[0]/NET0131  & ~n9936 ;
  assign n9938 = ~n9911 & ~n9937 ;
  assign n9939 = \P1_reg2_reg[5]/NET0131  & ~n3435 ;
  assign n9940 = \P1_reg2_reg[5]/NET0131  & n3448 ;
  assign n9942 = \P1_reg2_reg[5]/NET0131  & ~n3466 ;
  assign n9943 = n3466 & n9073 ;
  assign n9944 = ~n9942 & ~n9943 ;
  assign n9945 = n1936 & ~n9944 ;
  assign n9949 = n3466 & ~n9085 ;
  assign n9950 = ~n9942 & ~n9949 ;
  assign n9951 = ~n3677 & ~n9950 ;
  assign n9946 = n3466 & ~n9079 ;
  assign n9947 = ~n9942 & ~n9946 ;
  assign n9948 = ~n3563 & ~n9947 ;
  assign n9941 = n3466 & ~n9065 ;
  assign n9952 = n1543 & n1763 ;
  assign n9953 = ~n3466 & n9090 ;
  assign n9954 = ~n3716 & ~n9953 ;
  assign n9955 = \P1_reg2_reg[5]/NET0131  & ~n9954 ;
  assign n9956 = ~n9952 & ~n9955 ;
  assign n9957 = ~n9941 & n9956 ;
  assign n9958 = ~n9948 & n9957 ;
  assign n9959 = ~n9951 & n9958 ;
  assign n9960 = ~n9945 & n9959 ;
  assign n9961 = n3450 & ~n9960 ;
  assign n9962 = ~n9940 & ~n9961 ;
  assign n9963 = \P1_state_reg[0]/NET0131  & ~n9962 ;
  assign n9964 = ~n9939 & ~n9963 ;
  assign n9965 = \P1_reg0_reg[11]/NET0131  & ~n3435 ;
  assign n9966 = \P1_reg0_reg[11]/NET0131  & n3448 ;
  assign n9968 = \P1_reg0_reg[11]/NET0131  & ~n4396 ;
  assign n9969 = n4396 & n8010 ;
  assign n9970 = ~n9968 & ~n9969 ;
  assign n9971 = ~n3563 & ~n9970 ;
  assign n9967 = \P1_reg0_reg[11]/NET0131  & ~n4494 ;
  assign n9978 = n4396 & ~n9279 ;
  assign n9979 = ~n9967 & ~n9978 ;
  assign n9980 = ~n9971 & n9979 ;
  assign n9972 = n4396 & n8018 ;
  assign n9973 = ~n9968 & ~n9972 ;
  assign n9974 = n1936 & ~n9973 ;
  assign n9975 = n4396 & ~n8004 ;
  assign n9976 = ~n9968 & ~n9975 ;
  assign n9977 = ~n3677 & ~n9976 ;
  assign n9981 = ~n9974 & ~n9977 ;
  assign n9982 = n9980 & n9981 ;
  assign n9983 = n3450 & ~n9982 ;
  assign n9984 = ~n9966 & ~n9983 ;
  assign n9985 = \P1_state_reg[0]/NET0131  & ~n9984 ;
  assign n9986 = ~n9965 & ~n9985 ;
  assign n9987 = \P2_reg2_reg[4]/NET0131  & ~n1983 ;
  assign n9988 = \P2_reg2_reg[4]/NET0131  & n2024 ;
  assign n9990 = \P2_reg2_reg[4]/NET0131  & ~n3758 ;
  assign n9991 = n3758 & ~n8945 ;
  assign n9992 = ~n9990 & ~n9991 ;
  assign n9993 = n3411 & ~n9992 ;
  assign n9997 = n3758 & ~n8957 ;
  assign n9998 = ~n9990 & ~n9997 ;
  assign n9999 = ~n3320 & ~n9998 ;
  assign n9994 = n3758 & n8951 ;
  assign n9995 = ~n9990 & ~n9994 ;
  assign n9996 = ~n3177 & ~n9995 ;
  assign n10000 = n3758 & n8962 ;
  assign n10001 = ~n9990 & ~n10000 ;
  assign n10002 = n3355 & ~n10001 ;
  assign n10004 = \P2_reg2_reg[4]/NET0131  & ~n3774 ;
  assign n9989 = n3758 & n9159 ;
  assign n10003 = n2635 & n3420 ;
  assign n10005 = ~n9989 & ~n10003 ;
  assign n10006 = ~n10004 & n10005 ;
  assign n10007 = ~n10002 & n10006 ;
  assign n10008 = ~n9996 & n10007 ;
  assign n10009 = ~n9999 & n10008 ;
  assign n10010 = ~n9993 & n10009 ;
  assign n10011 = n2026 & ~n10010 ;
  assign n10012 = ~n9988 & ~n10011 ;
  assign n10013 = \P1_state_reg[0]/NET0131  & ~n10012 ;
  assign n10014 = ~n9987 & ~n10013 ;
  assign n10015 = ~n3758 & n9903 ;
  assign n10016 = ~n3417 & ~n10015 ;
  assign n10017 = n5287 & ~n5289 ;
  assign n10018 = n10016 & n10017 ;
  assign n10019 = \P2_reg2_reg[5]/NET0131  & ~n10018 ;
  assign n10020 = n2526 & n3420 ;
  assign n10021 = n3758 & ~n9852 ;
  assign n10022 = ~n10020 & ~n10021 ;
  assign n10023 = n5287 & ~n10022 ;
  assign n10024 = ~n10019 & ~n10023 ;
  assign n10025 = \P1_reg0_reg[14]/NET0131  & ~n3435 ;
  assign n10026 = \P1_reg0_reg[14]/NET0131  & n3448 ;
  assign n10028 = \P1_reg0_reg[14]/NET0131  & ~n4396 ;
  assign n10032 = n4396 & ~n8058 ;
  assign n10033 = ~n10028 & ~n10032 ;
  assign n10034 = ~n3563 & ~n4396 ;
  assign n10035 = n8062 & ~n10034 ;
  assign n10036 = ~n10033 & ~n10035 ;
  assign n10029 = n4396 & ~n8047 ;
  assign n10030 = ~n10028 & ~n10029 ;
  assign n10031 = n1936 & ~n10030 ;
  assign n10037 = n4396 & n8067 ;
  assign n10038 = ~n10028 & ~n10037 ;
  assign n10039 = n3712 & ~n10038 ;
  assign n10027 = n4396 & n9307 ;
  assign n10040 = \P1_reg0_reg[14]/NET0131  & ~n4493 ;
  assign n10041 = ~n10027 & ~n10040 ;
  assign n10042 = ~n10039 & n10041 ;
  assign n10043 = ~n10031 & n10042 ;
  assign n10044 = ~n10036 & n10043 ;
  assign n10045 = n3450 & ~n10044 ;
  assign n10046 = ~n10026 & ~n10045 ;
  assign n10047 = \P1_state_reg[0]/NET0131  & ~n10046 ;
  assign n10048 = ~n10025 & ~n10047 ;
  assign n10049 = \P1_reg0_reg[5]/NET0131  & ~n3435 ;
  assign n10050 = \P1_reg0_reg[5]/NET0131  & n3448 ;
  assign n10052 = \P1_reg0_reg[5]/NET0131  & ~n4396 ;
  assign n10053 = n4396 & n9073 ;
  assign n10054 = ~n10052 & ~n10053 ;
  assign n10055 = n1936 & ~n10054 ;
  assign n10059 = n4396 & ~n9085 ;
  assign n10060 = ~n10052 & ~n10059 ;
  assign n10061 = ~n3677 & ~n10060 ;
  assign n10056 = n4396 & ~n9079 ;
  assign n10057 = ~n10052 & ~n10056 ;
  assign n10058 = ~n3563 & ~n10057 ;
  assign n10062 = n4396 & n9063 ;
  assign n10063 = ~n10052 & ~n10062 ;
  assign n10064 = n3712 & ~n10063 ;
  assign n10051 = \P1_reg0_reg[5]/NET0131  & ~n4491 ;
  assign n10065 = ~n1562 & n4396 ;
  assign n10066 = ~n10052 & ~n10065 ;
  assign n10067 = n1880 & ~n10066 ;
  assign n10068 = ~n10051 & ~n10067 ;
  assign n10069 = ~n10064 & n10068 ;
  assign n10070 = ~n10058 & n10069 ;
  assign n10071 = ~n10061 & n10070 ;
  assign n10072 = ~n10055 & n10071 ;
  assign n10073 = n3450 & ~n10072 ;
  assign n10074 = ~n10050 & ~n10073 ;
  assign n10075 = \P1_state_reg[0]/NET0131  & ~n10074 ;
  assign n10076 = ~n10049 & ~n10075 ;
  assign n10077 = \P1_reg1_reg[11]/NET0131  & ~n3435 ;
  assign n10078 = \P1_reg1_reg[11]/NET0131  & n3448 ;
  assign n10080 = \P1_reg1_reg[11]/NET0131  & ~n4532 ;
  assign n10081 = n4532 & n8010 ;
  assign n10082 = ~n10080 & ~n10081 ;
  assign n10083 = ~n3563 & ~n10082 ;
  assign n10090 = n4532 & n8023 ;
  assign n10091 = ~n10080 & ~n10090 ;
  assign n10092 = n3712 & ~n10091 ;
  assign n10079 = \P1_reg1_reg[11]/NET0131  & ~n4491 ;
  assign n10093 = n1198 & n4532 ;
  assign n10094 = ~n10080 & ~n10093 ;
  assign n10095 = n1880 & ~n10094 ;
  assign n10096 = ~n10079 & ~n10095 ;
  assign n10097 = ~n10092 & n10096 ;
  assign n10098 = ~n10083 & n10097 ;
  assign n10084 = n4532 & n8018 ;
  assign n10085 = ~n10080 & ~n10084 ;
  assign n10086 = n1936 & ~n10085 ;
  assign n10087 = n4532 & ~n8004 ;
  assign n10088 = ~n10080 & ~n10087 ;
  assign n10089 = ~n3677 & ~n10088 ;
  assign n10099 = ~n10086 & ~n10089 ;
  assign n10100 = n10098 & n10099 ;
  assign n10101 = n3450 & ~n10100 ;
  assign n10102 = ~n10078 & ~n10101 ;
  assign n10103 = \P1_state_reg[0]/NET0131  & ~n10102 ;
  assign n10104 = ~n10077 & ~n10103 ;
  assign n10105 = \P1_reg1_reg[14]/NET0131  & ~n3435 ;
  assign n10106 = \P1_reg1_reg[14]/NET0131  & n3448 ;
  assign n10108 = \P1_reg1_reg[14]/NET0131  & ~n4532 ;
  assign n10112 = n4532 & ~n8058 ;
  assign n10113 = ~n10108 & ~n10112 ;
  assign n10114 = ~n3563 & ~n4532 ;
  assign n10115 = n8062 & ~n10114 ;
  assign n10116 = ~n10113 & ~n10115 ;
  assign n10109 = n4532 & ~n8047 ;
  assign n10110 = ~n10108 & ~n10109 ;
  assign n10111 = n1936 & ~n10110 ;
  assign n10117 = n4532 & n8067 ;
  assign n10118 = ~n10108 & ~n10117 ;
  assign n10119 = n3712 & ~n10118 ;
  assign n10107 = n4532 & n9307 ;
  assign n10120 = \P1_reg1_reg[14]/NET0131  & ~n4541 ;
  assign n10121 = ~n10107 & ~n10120 ;
  assign n10122 = ~n10119 & n10121 ;
  assign n10123 = ~n10111 & n10122 ;
  assign n10124 = ~n10116 & n10123 ;
  assign n10125 = n3450 & ~n10124 ;
  assign n10126 = ~n10106 & ~n10125 ;
  assign n10127 = \P1_state_reg[0]/NET0131  & ~n10126 ;
  assign n10128 = ~n10105 & ~n10127 ;
  assign n10129 = \P2_reg0_reg[11]/NET0131  & ~n1983 ;
  assign n10130 = \P2_reg0_reg[11]/NET0131  & n2024 ;
  assign n10132 = \P2_reg0_reg[11]/NET0131  & ~n2040 ;
  assign n10133 = n2040 & n8129 ;
  assign n10134 = ~n10132 & ~n10133 ;
  assign n10135 = n3411 & ~n10134 ;
  assign n10136 = n2040 & n8135 ;
  assign n10137 = ~n10132 & ~n10136 ;
  assign n10138 = ~n3177 & ~n10137 ;
  assign n10131 = \P2_reg0_reg[11]/NET0131  & ~n8385 ;
  assign n10139 = n2040 & ~n9867 ;
  assign n10140 = ~n10131 & ~n10139 ;
  assign n10141 = ~n10138 & n10140 ;
  assign n10142 = ~n10135 & n10141 ;
  assign n10143 = n2026 & ~n10142 ;
  assign n10144 = ~n10130 & ~n10143 ;
  assign n10145 = \P1_state_reg[0]/NET0131  & ~n10144 ;
  assign n10146 = ~n10129 & ~n10145 ;
  assign n10147 = \P2_reg0_reg[14]/NET0131  & ~n1983 ;
  assign n10148 = \P2_reg0_reg[14]/NET0131  & n2024 ;
  assign n10151 = \P2_reg0_reg[14]/NET0131  & ~n2040 ;
  assign n10152 = n2040 & n8176 ;
  assign n10153 = ~n10151 & ~n10152 ;
  assign n10154 = n3355 & ~n10153 ;
  assign n10149 = \P2_reg0_reg[14]/NET0131  & ~n3423 ;
  assign n10150 = n2040 & n9437 ;
  assign n10164 = ~n10149 & ~n10150 ;
  assign n10165 = ~n10154 & n10164 ;
  assign n10161 = n2040 & n8171 ;
  assign n10162 = ~n10151 & ~n10161 ;
  assign n10163 = n3411 & ~n10162 ;
  assign n10155 = n2040 & n8182 ;
  assign n10156 = ~n10151 & ~n10155 ;
  assign n10157 = ~n3177 & ~n10156 ;
  assign n10158 = n2040 & ~n8188 ;
  assign n10159 = ~n10151 & ~n10158 ;
  assign n10160 = ~n3320 & ~n10159 ;
  assign n10166 = ~n10157 & ~n10160 ;
  assign n10167 = ~n10163 & n10166 ;
  assign n10168 = n10165 & n10167 ;
  assign n10169 = n2026 & ~n10168 ;
  assign n10170 = ~n10148 & ~n10169 ;
  assign n10171 = \P1_state_reg[0]/NET0131  & ~n10170 ;
  assign n10172 = ~n10147 & ~n10171 ;
  assign n10173 = \P1_reg1_reg[3]/NET0131  & ~n3435 ;
  assign n10174 = \P1_reg1_reg[3]/NET0131  & n3448 ;
  assign n10178 = \P1_reg1_reg[3]/NET0131  & ~n4532 ;
  assign n10179 = n4532 & n9709 ;
  assign n10180 = ~n10178 & ~n10179 ;
  assign n10181 = n1936 & ~n10180 ;
  assign n10182 = n4532 & ~n9716 ;
  assign n10183 = ~n10178 & ~n10182 ;
  assign n10184 = ~n3563 & ~n10183 ;
  assign n10175 = ~n3677 & n9723 ;
  assign n10176 = n9702 & ~n10175 ;
  assign n10177 = n4532 & ~n10176 ;
  assign n10185 = ~n3677 & ~n4532 ;
  assign n10186 = n9835 & ~n10185 ;
  assign n10187 = \P1_reg1_reg[3]/NET0131  & ~n10186 ;
  assign n10188 = ~n10177 & ~n10187 ;
  assign n10189 = ~n10184 & n10188 ;
  assign n10190 = ~n10181 & n10189 ;
  assign n10191 = n3450 & ~n10190 ;
  assign n10192 = ~n10174 & ~n10191 ;
  assign n10193 = \P1_state_reg[0]/NET0131  & ~n10192 ;
  assign n10194 = ~n10173 & ~n10193 ;
  assign n10195 = \P1_reg1_reg[7]/NET0131  & ~n3435 ;
  assign n10196 = \P1_reg1_reg[7]/NET0131  & n3448 ;
  assign n10198 = \P1_reg1_reg[7]/NET0131  & ~n4532 ;
  assign n10199 = n4532 & n9794 ;
  assign n10200 = ~n10198 & ~n10199 ;
  assign n10201 = ~n3563 & ~n10200 ;
  assign n10197 = \P1_reg1_reg[7]/NET0131  & ~n4573 ;
  assign n10208 = ~n1514 & n1880 ;
  assign n10209 = ~n9808 & ~n10208 ;
  assign n10210 = n4532 & ~n10209 ;
  assign n10211 = ~n10197 & ~n10210 ;
  assign n10212 = ~n10201 & n10211 ;
  assign n10202 = n4532 & n9802 ;
  assign n10203 = ~n10198 & ~n10202 ;
  assign n10204 = n1936 & ~n10203 ;
  assign n10205 = n4532 & ~n9788 ;
  assign n10206 = ~n10198 & ~n10205 ;
  assign n10207 = ~n3677 & ~n10206 ;
  assign n10213 = ~n10204 & ~n10207 ;
  assign n10214 = n10212 & n10213 ;
  assign n10215 = n3450 & ~n10214 ;
  assign n10216 = ~n10196 & ~n10215 ;
  assign n10217 = \P1_state_reg[0]/NET0131  & ~n10216 ;
  assign n10218 = ~n10195 & ~n10217 ;
  assign n10219 = \P2_reg0_reg[3]/NET0131  & ~n1983 ;
  assign n10220 = \P2_reg0_reg[3]/NET0131  & n2024 ;
  assign n10222 = \P2_reg0_reg[3]/NET0131  & ~n2040 ;
  assign n10223 = n2040 & n9597 ;
  assign n10224 = ~n10222 & ~n10223 ;
  assign n10225 = n3411 & ~n10224 ;
  assign n10226 = n2040 & ~n9591 ;
  assign n10227 = ~n10222 & ~n10226 ;
  assign n10228 = ~n3177 & ~n10227 ;
  assign n10221 = n2040 & ~n9587 ;
  assign n10229 = ~n2040 & ~n9904 ;
  assign n10230 = n3421 & ~n10229 ;
  assign n10231 = \P2_reg0_reg[3]/NET0131  & ~n10230 ;
  assign n10232 = ~n10221 & ~n10231 ;
  assign n10233 = ~n10228 & n10232 ;
  assign n10234 = ~n10225 & n10233 ;
  assign n10235 = n2026 & ~n10234 ;
  assign n10236 = ~n10220 & ~n10235 ;
  assign n10237 = \P1_state_reg[0]/NET0131  & ~n10236 ;
  assign n10238 = ~n10219 & ~n10237 ;
  assign n10239 = \P2_reg0_reg[7]/NET0131  & ~n1983 ;
  assign n10240 = \P2_reg0_reg[7]/NET0131  & n2024 ;
  assign n10242 = \P2_reg0_reg[7]/NET0131  & ~n2040 ;
  assign n10243 = n2040 & n9664 ;
  assign n10244 = ~n10242 & ~n10243 ;
  assign n10245 = n3411 & ~n10244 ;
  assign n10246 = n2040 & n9670 ;
  assign n10247 = ~n10242 & ~n10246 ;
  assign n10248 = ~n3177 & ~n10247 ;
  assign n10241 = \P2_reg0_reg[7]/NET0131  & ~n8385 ;
  assign n10250 = ~n3320 & ~n9676 ;
  assign n10249 = n2495 & n3358 ;
  assign n10251 = ~n9682 & ~n10249 ;
  assign n10252 = ~n10250 & n10251 ;
  assign n10253 = n2040 & ~n10252 ;
  assign n10254 = ~n10241 & ~n10253 ;
  assign n10255 = ~n10248 & n10254 ;
  assign n10256 = ~n10245 & n10255 ;
  assign n10257 = n2026 & ~n10256 ;
  assign n10258 = ~n10240 & ~n10257 ;
  assign n10259 = \P1_state_reg[0]/NET0131  & ~n10258 ;
  assign n10260 = ~n10239 & ~n10259 ;
  assign n10261 = \P2_reg1_reg[3]/NET0131  & ~n1983 ;
  assign n10262 = \P2_reg1_reg[3]/NET0131  & n2024 ;
  assign n10264 = \P2_reg1_reg[3]/NET0131  & ~n3733 ;
  assign n10265 = n3733 & n9597 ;
  assign n10266 = ~n10264 & ~n10265 ;
  assign n10267 = n3411 & ~n10266 ;
  assign n10268 = n3733 & ~n9591 ;
  assign n10269 = ~n10264 & ~n10268 ;
  assign n10270 = ~n3177 & ~n10269 ;
  assign n10263 = \P2_reg1_reg[3]/NET0131  & ~n9906 ;
  assign n10271 = n3733 & ~n9587 ;
  assign n10272 = ~n10263 & ~n10271 ;
  assign n10273 = ~n10270 & n10272 ;
  assign n10274 = ~n10267 & n10273 ;
  assign n10275 = n2026 & ~n10274 ;
  assign n10276 = ~n10262 & ~n10275 ;
  assign n10277 = \P1_state_reg[0]/NET0131  & ~n10276 ;
  assign n10278 = ~n10261 & ~n10277 ;
  assign n10279 = \P2_reg1_reg[7]/NET0131  & ~n1983 ;
  assign n10280 = \P2_reg1_reg[7]/NET0131  & n2024 ;
  assign n10282 = \P2_reg1_reg[7]/NET0131  & ~n3733 ;
  assign n10283 = n3733 & n9664 ;
  assign n10284 = ~n10282 & ~n10283 ;
  assign n10285 = n3411 & ~n10284 ;
  assign n10286 = n3733 & n9670 ;
  assign n10287 = ~n10282 & ~n10286 ;
  assign n10288 = ~n3177 & ~n10287 ;
  assign n10281 = \P2_reg1_reg[7]/NET0131  & ~n8532 ;
  assign n10289 = n3733 & ~n10252 ;
  assign n10290 = ~n10281 & ~n10289 ;
  assign n10291 = ~n10288 & n10290 ;
  assign n10292 = ~n10285 & n10291 ;
  assign n10293 = n2026 & ~n10292 ;
  assign n10294 = ~n10280 & ~n10293 ;
  assign n10295 = \P1_state_reg[0]/NET0131  & ~n10294 ;
  assign n10296 = ~n10279 & ~n10295 ;
  assign n10297 = \P1_reg2_reg[3]/NET0131  & ~n3435 ;
  assign n10298 = \P1_reg2_reg[3]/NET0131  & n3448 ;
  assign n10300 = \P1_reg2_reg[3]/NET0131  & ~n3466 ;
  assign n10301 = n3466 & n9709 ;
  assign n10302 = ~n10300 & ~n10301 ;
  assign n10303 = n1936 & ~n10302 ;
  assign n10304 = n3466 & ~n9716 ;
  assign n10305 = ~n10300 & ~n10304 ;
  assign n10306 = ~n3563 & ~n10305 ;
  assign n10307 = n3466 & n9723 ;
  assign n10308 = ~n10300 & ~n10307 ;
  assign n10309 = ~n3677 & ~n10308 ;
  assign n10299 = n3466 & ~n9702 ;
  assign n10310 = ~\P1_reg3_reg[3]/NET0131  & n1763 ;
  assign n10311 = \P1_reg2_reg[3]/NET0131  & ~n9954 ;
  assign n10312 = ~n10310 & ~n10311 ;
  assign n10313 = ~n10299 & n10312 ;
  assign n10314 = ~n10309 & n10313 ;
  assign n10315 = ~n10306 & n10314 ;
  assign n10316 = ~n10303 & n10315 ;
  assign n10317 = n3450 & ~n10316 ;
  assign n10318 = ~n10298 & ~n10317 ;
  assign n10319 = \P1_state_reg[0]/NET0131  & ~n10318 ;
  assign n10320 = ~n10297 & ~n10319 ;
  assign n10321 = \P1_reg2_reg[6]/NET0131  & ~n3435 ;
  assign n10322 = \P1_reg2_reg[6]/NET0131  & n3448 ;
  assign n10325 = \P1_reg2_reg[6]/NET0131  & ~n3466 ;
  assign n10326 = n3466 & n9755 ;
  assign n10327 = ~n10325 & ~n10326 ;
  assign n10328 = ~n3677 & ~n10327 ;
  assign n10335 = n3466 & n9766 ;
  assign n10336 = ~n10325 & ~n10335 ;
  assign n10337 = n3712 & ~n10336 ;
  assign n10339 = \P1_reg2_reg[6]/NET0131  & ~n3718 ;
  assign n10323 = ~n1537 & n1880 ;
  assign n10324 = n3466 & n10323 ;
  assign n10338 = n1518 & n1763 ;
  assign n10340 = ~n10324 & ~n10338 ;
  assign n10341 = ~n10339 & n10340 ;
  assign n10342 = ~n10337 & n10341 ;
  assign n10343 = ~n10328 & n10342 ;
  assign n10329 = n3466 & ~n9761 ;
  assign n10330 = ~n10325 & ~n10329 ;
  assign n10331 = ~n3563 & ~n10330 ;
  assign n10332 = n3466 & ~n9749 ;
  assign n10333 = ~n10325 & ~n10332 ;
  assign n10334 = n1936 & ~n10333 ;
  assign n10344 = ~n10331 & ~n10334 ;
  assign n10345 = n10343 & n10344 ;
  assign n10346 = n3450 & ~n10345 ;
  assign n10347 = ~n10322 & ~n10346 ;
  assign n10348 = \P1_state_reg[0]/NET0131  & ~n10347 ;
  assign n10349 = ~n10321 & ~n10348 ;
  assign n10350 = \P1_reg2_reg[7]/NET0131  & ~n3435 ;
  assign n10351 = \P1_reg2_reg[7]/NET0131  & n3448 ;
  assign n10353 = \P1_reg2_reg[7]/NET0131  & ~n3466 ;
  assign n10354 = n3466 & n9794 ;
  assign n10355 = ~n10353 & ~n10354 ;
  assign n10356 = ~n3563 & ~n10355 ;
  assign n10363 = n3466 & ~n10209 ;
  assign n10352 = \P1_reg2_reg[7]/NET0131  & ~n5914 ;
  assign n10364 = n1491 & n1763 ;
  assign n10365 = ~n10352 & ~n10364 ;
  assign n10366 = ~n10363 & n10365 ;
  assign n10367 = ~n10356 & n10366 ;
  assign n10357 = n3466 & n9802 ;
  assign n10358 = ~n10353 & ~n10357 ;
  assign n10359 = n1936 & ~n10358 ;
  assign n10360 = n3466 & ~n9788 ;
  assign n10361 = ~n10353 & ~n10360 ;
  assign n10362 = ~n3677 & ~n10361 ;
  assign n10368 = ~n10359 & ~n10362 ;
  assign n10369 = n10367 & n10368 ;
  assign n10370 = n3450 & ~n10369 ;
  assign n10371 = ~n10351 & ~n10370 ;
  assign n10372 = \P1_state_reg[0]/NET0131  & ~n10371 ;
  assign n10373 = ~n10350 & ~n10372 ;
  assign n10374 = \P2_reg2_reg[3]/NET0131  & ~n1983 ;
  assign n10375 = \P2_reg2_reg[3]/NET0131  & n2024 ;
  assign n10377 = \P2_reg2_reg[3]/NET0131  & ~n3758 ;
  assign n10378 = n3758 & n9597 ;
  assign n10379 = ~n10377 & ~n10378 ;
  assign n10380 = n3411 & ~n10379 ;
  assign n10381 = n3758 & ~n9591 ;
  assign n10382 = ~n10377 & ~n10381 ;
  assign n10383 = ~n3177 & ~n10382 ;
  assign n10384 = n3758 & ~n9587 ;
  assign n10376 = ~\P2_reg3_reg[3]/NET0131  & n3420 ;
  assign n10385 = ~n7769 & n10016 ;
  assign n10386 = \P2_reg2_reg[3]/NET0131  & ~n10385 ;
  assign n10387 = ~n10376 & ~n10386 ;
  assign n10388 = ~n10384 & n10387 ;
  assign n10389 = ~n10383 & n10388 ;
  assign n10390 = ~n10380 & n10389 ;
  assign n10391 = n2026 & ~n10390 ;
  assign n10392 = ~n10375 & ~n10391 ;
  assign n10393 = \P1_state_reg[0]/NET0131  & ~n10392 ;
  assign n10394 = ~n10374 & ~n10393 ;
  assign n10395 = \P2_reg2_reg[6]/NET0131  & ~n1983 ;
  assign n10396 = \P2_reg2_reg[6]/NET0131  & n2024 ;
  assign n10399 = \P2_reg2_reg[6]/NET0131  & ~n3758 ;
  assign n10400 = n3758 & n9624 ;
  assign n10401 = ~n10399 & ~n10400 ;
  assign n10402 = n3411 & ~n10401 ;
  assign n10406 = n3758 & n9636 ;
  assign n10407 = ~n10399 & ~n10406 ;
  assign n10408 = ~n3177 & ~n10407 ;
  assign n10403 = n3758 & ~n9630 ;
  assign n10404 = ~n10399 & ~n10403 ;
  assign n10405 = ~n3320 & ~n10404 ;
  assign n10409 = n3758 & n9641 ;
  assign n10410 = ~n10399 & ~n10409 ;
  assign n10411 = n3355 & ~n10410 ;
  assign n10413 = \P2_reg2_reg[6]/NET0131  & ~n3774 ;
  assign n10397 = ~n2521 & n3358 ;
  assign n10398 = n3758 & n10397 ;
  assign n10412 = n2499 & n3420 ;
  assign n10414 = ~n10398 & ~n10412 ;
  assign n10415 = ~n10413 & n10414 ;
  assign n10416 = ~n10411 & n10415 ;
  assign n10417 = ~n10405 & n10416 ;
  assign n10418 = ~n10408 & n10417 ;
  assign n10419 = ~n10402 & n10418 ;
  assign n10420 = n2026 & ~n10419 ;
  assign n10421 = ~n10396 & ~n10420 ;
  assign n10422 = \P1_state_reg[0]/NET0131  & ~n10421 ;
  assign n10423 = ~n10395 & ~n10422 ;
  assign n10424 = \P2_reg2_reg[7]/NET0131  & n2024 ;
  assign n10426 = \P2_reg2_reg[7]/NET0131  & ~n3758 ;
  assign n10427 = n3758 & n9664 ;
  assign n10428 = ~n10426 & ~n10427 ;
  assign n10429 = n3411 & ~n10428 ;
  assign n10430 = n3758 & n9670 ;
  assign n10431 = ~n10426 & ~n10430 ;
  assign n10432 = ~n3177 & ~n10431 ;
  assign n10436 = n3758 & n9681 ;
  assign n10437 = ~n10426 & ~n10436 ;
  assign n10438 = n3355 & ~n10437 ;
  assign n10433 = n3758 & ~n9676 ;
  assign n10434 = ~n10426 & ~n10433 ;
  assign n10435 = ~n3320 & ~n10434 ;
  assign n10425 = \P2_reg2_reg[7]/NET0131  & ~n3774 ;
  assign n10439 = n2476 & n3420 ;
  assign n10440 = n3758 & n10249 ;
  assign n10441 = ~n10439 & ~n10440 ;
  assign n10442 = ~n10425 & n10441 ;
  assign n10443 = ~n10435 & n10442 ;
  assign n10444 = ~n10438 & n10443 ;
  assign n10445 = ~n10432 & n10444 ;
  assign n10446 = ~n10429 & n10445 ;
  assign n10447 = n2026 & ~n10446 ;
  assign n10448 = ~n10424 & ~n10447 ;
  assign n10449 = \P1_state_reg[0]/NET0131  & ~n10448 ;
  assign n10450 = \P2_reg2_reg[7]/NET0131  & ~n1983 ;
  assign n10451 = ~n10449 & ~n10450 ;
  assign n10452 = \P1_reg0_reg[3]/NET0131  & ~n3435 ;
  assign n10453 = \P1_reg0_reg[3]/NET0131  & n3448 ;
  assign n10455 = \P1_reg0_reg[3]/NET0131  & ~n4396 ;
  assign n10456 = n4396 & n9709 ;
  assign n10457 = ~n10455 & ~n10456 ;
  assign n10458 = n1936 & ~n10457 ;
  assign n10459 = n4396 & ~n9716 ;
  assign n10460 = ~n10455 & ~n10459 ;
  assign n10461 = ~n3563 & ~n10460 ;
  assign n10454 = n4396 & ~n10176 ;
  assign n10462 = ~n3677 & ~n4396 ;
  assign n10463 = n4494 & ~n10462 ;
  assign n10464 = \P1_reg0_reg[3]/NET0131  & ~n10463 ;
  assign n10465 = ~n10454 & ~n10464 ;
  assign n10466 = ~n10461 & n10465 ;
  assign n10467 = ~n10458 & n10466 ;
  assign n10468 = n3450 & ~n10467 ;
  assign n10469 = ~n10453 & ~n10468 ;
  assign n10470 = \P1_state_reg[0]/NET0131  & ~n10469 ;
  assign n10471 = ~n10452 & ~n10470 ;
  assign n10472 = \P1_reg0_reg[7]/NET0131  & ~n3435 ;
  assign n10473 = \P1_reg0_reg[7]/NET0131  & n3448 ;
  assign n10475 = \P1_reg0_reg[7]/NET0131  & ~n4396 ;
  assign n10476 = n4396 & n9794 ;
  assign n10477 = ~n10475 & ~n10476 ;
  assign n10478 = ~n3563 & ~n10477 ;
  assign n10485 = n4396 & n9807 ;
  assign n10486 = ~n10475 & ~n10485 ;
  assign n10487 = n3712 & ~n10486 ;
  assign n10474 = \P1_reg0_reg[7]/NET0131  & ~n4491 ;
  assign n10488 = ~n1514 & n4396 ;
  assign n10489 = ~n10475 & ~n10488 ;
  assign n10490 = n1880 & ~n10489 ;
  assign n10491 = ~n10474 & ~n10490 ;
  assign n10492 = ~n10487 & n10491 ;
  assign n10493 = ~n10478 & n10492 ;
  assign n10479 = n4396 & n9802 ;
  assign n10480 = ~n10475 & ~n10479 ;
  assign n10481 = n1936 & ~n10480 ;
  assign n10482 = n4396 & ~n9788 ;
  assign n10483 = ~n10475 & ~n10482 ;
  assign n10484 = ~n3677 & ~n10483 ;
  assign n10494 = ~n10481 & ~n10484 ;
  assign n10495 = n10493 & n10494 ;
  assign n10496 = n3450 & ~n10495 ;
  assign n10497 = ~n10473 & ~n10496 ;
  assign n10498 = \P1_state_reg[0]/NET0131  & ~n10497 ;
  assign n10499 = ~n10472 & ~n10498 ;
  assign n10500 = \P1_reg1_reg[6]/NET0131  & ~n3435 ;
  assign n10501 = \P1_reg1_reg[6]/NET0131  & n3448 ;
  assign n10503 = \P1_reg1_reg[6]/NET0131  & ~n4532 ;
  assign n10504 = n4532 & ~n9749 ;
  assign n10505 = ~n10503 & ~n10504 ;
  assign n10506 = n1936 & ~n10505 ;
  assign n10513 = n4532 & n9766 ;
  assign n10514 = ~n10503 & ~n10513 ;
  assign n10515 = n3712 & ~n10514 ;
  assign n10502 = n4532 & n10323 ;
  assign n10516 = \P1_reg1_reg[6]/NET0131  & ~n4541 ;
  assign n10517 = ~n10502 & ~n10516 ;
  assign n10518 = ~n10515 & n10517 ;
  assign n10519 = ~n10506 & n10518 ;
  assign n10507 = n4532 & ~n9761 ;
  assign n10508 = ~n10503 & ~n10507 ;
  assign n10509 = ~n3563 & ~n10508 ;
  assign n10510 = n4532 & n9755 ;
  assign n10511 = ~n10503 & ~n10510 ;
  assign n10512 = ~n3677 & ~n10511 ;
  assign n10520 = ~n10509 & ~n10512 ;
  assign n10521 = n10519 & n10520 ;
  assign n10522 = n3450 & ~n10521 ;
  assign n10523 = ~n10501 & ~n10522 ;
  assign n10524 = \P1_state_reg[0]/NET0131  & ~n10523 ;
  assign n10525 = ~n10500 & ~n10524 ;
  assign n10526 = \P2_reg0_reg[6]/NET0131  & ~n1983 ;
  assign n10527 = \P2_reg0_reg[6]/NET0131  & n2024 ;
  assign n10529 = \P2_reg0_reg[6]/NET0131  & ~n2040 ;
  assign n10530 = n2040 & n9624 ;
  assign n10531 = ~n10529 & ~n10530 ;
  assign n10532 = n3411 & ~n10531 ;
  assign n10536 = n2040 & ~n9630 ;
  assign n10537 = ~n10529 & ~n10536 ;
  assign n10538 = ~n3320 & ~n10537 ;
  assign n10533 = n2040 & n9636 ;
  assign n10534 = ~n10529 & ~n10533 ;
  assign n10535 = ~n3177 & ~n10534 ;
  assign n10539 = n2040 & n9641 ;
  assign n10540 = ~n10529 & ~n10539 ;
  assign n10541 = n3355 & ~n10540 ;
  assign n10528 = \P2_reg0_reg[6]/NET0131  & ~n3423 ;
  assign n10542 = n2040 & n10397 ;
  assign n10543 = ~n10528 & ~n10542 ;
  assign n10544 = ~n10541 & n10543 ;
  assign n10545 = ~n10535 & n10544 ;
  assign n10546 = ~n10538 & n10545 ;
  assign n10547 = ~n10532 & n10546 ;
  assign n10548 = n2026 & ~n10547 ;
  assign n10549 = ~n10527 & ~n10548 ;
  assign n10550 = \P1_state_reg[0]/NET0131  & ~n10549 ;
  assign n10551 = ~n10526 & ~n10550 ;
  assign n10552 = \P2_reg1_reg[6]/NET0131  & ~n1983 ;
  assign n10553 = \P2_reg1_reg[6]/NET0131  & n2024 ;
  assign n10555 = \P2_reg1_reg[6]/NET0131  & ~n3733 ;
  assign n10556 = n3733 & n9624 ;
  assign n10557 = ~n10555 & ~n10556 ;
  assign n10558 = n3411 & ~n10557 ;
  assign n10562 = n3733 & ~n9630 ;
  assign n10563 = ~n10555 & ~n10562 ;
  assign n10564 = ~n3320 & ~n10563 ;
  assign n10559 = n3733 & n9636 ;
  assign n10560 = ~n10555 & ~n10559 ;
  assign n10561 = ~n3177 & ~n10560 ;
  assign n10565 = n3733 & n9641 ;
  assign n10566 = ~n10555 & ~n10565 ;
  assign n10567 = n3355 & ~n10566 ;
  assign n10554 = n3733 & n10397 ;
  assign n10568 = \P2_reg1_reg[6]/NET0131  & ~n3743 ;
  assign n10569 = ~n10554 & ~n10568 ;
  assign n10570 = ~n10567 & n10569 ;
  assign n10571 = ~n10561 & n10570 ;
  assign n10572 = ~n10564 & n10571 ;
  assign n10573 = ~n10558 & n10572 ;
  assign n10574 = n2026 & ~n10573 ;
  assign n10575 = ~n10553 & ~n10574 ;
  assign n10576 = \P1_state_reg[0]/NET0131  & ~n10575 ;
  assign n10577 = ~n10552 & ~n10576 ;
  assign n10578 = \P1_reg0_reg[6]/NET0131  & ~n3435 ;
  assign n10579 = \P1_reg0_reg[6]/NET0131  & n3448 ;
  assign n10581 = \P1_reg0_reg[6]/NET0131  & ~n4396 ;
  assign n10582 = n4396 & ~n9761 ;
  assign n10583 = ~n10581 & ~n10582 ;
  assign n10584 = ~n3563 & ~n10583 ;
  assign n10591 = n4396 & n9766 ;
  assign n10592 = ~n10581 & ~n10591 ;
  assign n10593 = n3712 & ~n10592 ;
  assign n10580 = n4396 & n10323 ;
  assign n10594 = \P1_reg0_reg[6]/NET0131  & ~n4493 ;
  assign n10595 = ~n10580 & ~n10594 ;
  assign n10596 = ~n10593 & n10595 ;
  assign n10597 = ~n10584 & n10596 ;
  assign n10585 = n4396 & ~n9749 ;
  assign n10586 = ~n10581 & ~n10585 ;
  assign n10587 = n1936 & ~n10586 ;
  assign n10588 = n4396 & n9755 ;
  assign n10589 = ~n10581 & ~n10588 ;
  assign n10590 = ~n3677 & ~n10589 ;
  assign n10598 = ~n10587 & ~n10590 ;
  assign n10599 = n10597 & n10598 ;
  assign n10600 = n3450 & ~n10599 ;
  assign n10601 = ~n10579 & ~n10600 ;
  assign n10602 = \P1_state_reg[0]/NET0131  & ~n10601 ;
  assign n10603 = ~n10578 & ~n10602 ;
  assign n10604 = \P2_reg3_reg[2]/NET0131  & ~n1983 ;
  assign n10605 = \P2_reg3_reg[2]/NET0131  & n2024 ;
  assign n10607 = \P2_reg3_reg[2]/NET0131  & ~n3788 ;
  assign n10620 = n2616 & ~n3375 ;
  assign n10621 = ~n3376 & ~n10620 ;
  assign n10622 = ~n2058 & ~n10621 ;
  assign n10623 = n2058 & n2574 ;
  assign n10624 = ~n10622 & ~n10623 ;
  assign n10625 = n3788 & n10624 ;
  assign n10626 = ~n10607 & ~n10625 ;
  assign n10627 = n3411 & ~n10626 ;
  assign n10614 = n3819 & ~n4202 ;
  assign n10615 = ~n3819 & n4202 ;
  assign n10616 = ~n10614 & ~n10615 ;
  assign n10617 = n3788 & ~n10616 ;
  assign n10618 = ~n10607 & ~n10617 ;
  assign n10619 = ~n3320 & ~n10618 ;
  assign n10608 = ~n2607 & n4202 ;
  assign n10609 = n2607 & ~n4202 ;
  assign n10610 = ~n10608 & ~n10609 ;
  assign n10611 = n3788 & ~n10610 ;
  assign n10612 = ~n10607 & ~n10611 ;
  assign n10613 = ~n3177 & ~n10612 ;
  assign n10628 = ~n2566 & ~n3326 ;
  assign n10629 = ~n3327 & ~n10628 ;
  assign n10630 = n3788 & n10629 ;
  assign n10631 = ~n10607 & ~n10630 ;
  assign n10632 = n3355 & ~n10631 ;
  assign n10606 = ~n2566 & ~n3965 ;
  assign n10633 = \P2_reg3_reg[2]/NET0131  & ~n3962 ;
  assign n10634 = ~n10606 & ~n10633 ;
  assign n10635 = ~n10632 & n10634 ;
  assign n10636 = ~n10613 & n10635 ;
  assign n10637 = ~n10619 & n10636 ;
  assign n10638 = ~n10627 & n10637 ;
  assign n10639 = n2026 & ~n10638 ;
  assign n10640 = ~n10605 & ~n10639 ;
  assign n10641 = \P1_state_reg[0]/NET0131  & ~n10640 ;
  assign n10642 = ~n10604 & ~n10641 ;
  assign n10643 = \P1_reg3_reg[2]/NET0131  & ~n3435 ;
  assign n10644 = \P1_reg3_reg[2]/NET0131  & n3448 ;
  assign n10646 = \P1_reg3_reg[2]/NET0131  & ~n3980 ;
  assign n10659 = n1617 & ~n3572 ;
  assign n10660 = ~n3573 & ~n10659 ;
  assign n10661 = ~n537 & ~n10660 ;
  assign n10662 = n537 & n1641 ;
  assign n10663 = ~n10661 & ~n10662 ;
  assign n10664 = n3980 & n10663 ;
  assign n10665 = ~n10646 & ~n10664 ;
  assign n10666 = n1936 & ~n10665 ;
  assign n10653 = n1674 & ~n1779 ;
  assign n10654 = ~n1674 & n1779 ;
  assign n10655 = ~n10653 & ~n10654 ;
  assign n10656 = n3980 & ~n10655 ;
  assign n10657 = ~n10646 & ~n10656 ;
  assign n10658 = ~n3677 & ~n10657 ;
  assign n10647 = n1779 & ~n3507 ;
  assign n10648 = ~n1779 & n3507 ;
  assign n10649 = ~n10647 & ~n10648 ;
  assign n10650 = n3980 & ~n10649 ;
  assign n10651 = ~n10646 & ~n10650 ;
  assign n10652 = ~n3563 & ~n10651 ;
  assign n10667 = ~n1609 & ~n3679 ;
  assign n10668 = ~n3680 & ~n10667 ;
  assign n10669 = n3980 & n10668 ;
  assign n10670 = ~n10646 & ~n10669 ;
  assign n10671 = n3712 & ~n10670 ;
  assign n10645 = ~n1609 & ~n4067 ;
  assign n10672 = \P1_reg3_reg[2]/NET0131  & ~n4064 ;
  assign n10673 = ~n10645 & ~n10672 ;
  assign n10674 = ~n10671 & n10673 ;
  assign n10675 = ~n10652 & n10674 ;
  assign n10676 = ~n10658 & n10675 ;
  assign n10677 = ~n10666 & n10676 ;
  assign n10678 = n3450 & ~n10677 ;
  assign n10679 = ~n10644 & ~n10678 ;
  assign n10680 = \P1_state_reg[0]/NET0131  & ~n10679 ;
  assign n10681 = ~n10643 & ~n10680 ;
  assign n10682 = \P2_reg0_reg[2]/NET0131  & ~n1983 ;
  assign n10683 = \P2_reg0_reg[2]/NET0131  & n2024 ;
  assign n10686 = \P2_reg0_reg[2]/NET0131  & ~n2040 ;
  assign n10693 = n2040 & n10624 ;
  assign n10694 = ~n10686 & ~n10693 ;
  assign n10695 = n3411 & ~n10694 ;
  assign n10690 = n2040 & ~n10616 ;
  assign n10691 = ~n10686 & ~n10690 ;
  assign n10692 = ~n3320 & ~n10691 ;
  assign n10687 = n2040 & ~n10610 ;
  assign n10688 = ~n10686 & ~n10687 ;
  assign n10689 = ~n3177 & ~n10688 ;
  assign n10696 = n2040 & n10629 ;
  assign n10697 = ~n10686 & ~n10696 ;
  assign n10698 = n3355 & ~n10697 ;
  assign n10684 = ~n2566 & n3358 ;
  assign n10685 = n2040 & n10684 ;
  assign n10699 = \P2_reg0_reg[2]/NET0131  & ~n3423 ;
  assign n10700 = ~n10685 & ~n10699 ;
  assign n10701 = ~n10698 & n10700 ;
  assign n10702 = ~n10689 & n10701 ;
  assign n10703 = ~n10692 & n10702 ;
  assign n10704 = ~n10695 & n10703 ;
  assign n10705 = n2026 & ~n10704 ;
  assign n10706 = ~n10683 & ~n10705 ;
  assign n10707 = \P1_state_reg[0]/NET0131  & ~n10706 ;
  assign n10708 = ~n10682 & ~n10707 ;
  assign n10709 = \P2_reg1_reg[2]/NET0131  & ~n1983 ;
  assign n10710 = \P2_reg1_reg[2]/NET0131  & n2024 ;
  assign n10712 = \P2_reg1_reg[2]/NET0131  & ~n3733 ;
  assign n10719 = n3733 & n10624 ;
  assign n10720 = ~n10712 & ~n10719 ;
  assign n10721 = n3411 & ~n10720 ;
  assign n10716 = n3733 & ~n10610 ;
  assign n10717 = ~n10712 & ~n10716 ;
  assign n10718 = ~n3177 & ~n10717 ;
  assign n10713 = n3733 & ~n10616 ;
  assign n10714 = ~n10712 & ~n10713 ;
  assign n10715 = ~n3320 & ~n10714 ;
  assign n10722 = n3733 & n10629 ;
  assign n10723 = ~n10712 & ~n10722 ;
  assign n10724 = n3355 & ~n10723 ;
  assign n10711 = n3733 & n10684 ;
  assign n10725 = \P2_reg1_reg[2]/NET0131  & ~n3743 ;
  assign n10726 = ~n10711 & ~n10725 ;
  assign n10727 = ~n10724 & n10726 ;
  assign n10728 = ~n10715 & n10727 ;
  assign n10729 = ~n10718 & n10728 ;
  assign n10730 = ~n10721 & n10729 ;
  assign n10731 = n2026 & ~n10730 ;
  assign n10732 = ~n10710 & ~n10731 ;
  assign n10733 = \P1_state_reg[0]/NET0131  & ~n10732 ;
  assign n10734 = ~n10709 & ~n10733 ;
  assign n10735 = \P1_reg2_reg[2]/NET0131  & ~n3435 ;
  assign n10736 = \P1_reg2_reg[2]/NET0131  & n3448 ;
  assign n10739 = \P1_reg2_reg[2]/NET0131  & ~n3466 ;
  assign n10746 = n3466 & n10663 ;
  assign n10747 = ~n10739 & ~n10746 ;
  assign n10748 = n1936 & ~n10747 ;
  assign n10743 = n3466 & ~n10649 ;
  assign n10744 = ~n10739 & ~n10743 ;
  assign n10745 = ~n3563 & ~n10744 ;
  assign n10740 = n3466 & ~n10655 ;
  assign n10741 = ~n10739 & ~n10740 ;
  assign n10742 = ~n3677 & ~n10741 ;
  assign n10749 = n3466 & n10668 ;
  assign n10750 = ~n10739 & ~n10749 ;
  assign n10751 = n3712 & ~n10750 ;
  assign n10753 = \P1_reg2_reg[2]/NET0131  & ~n3718 ;
  assign n10737 = ~n1609 & n1880 ;
  assign n10738 = n3466 & n10737 ;
  assign n10752 = \P1_reg3_reg[2]/NET0131  & n1763 ;
  assign n10754 = ~n10738 & ~n10752 ;
  assign n10755 = ~n10753 & n10754 ;
  assign n10756 = ~n10751 & n10755 ;
  assign n10757 = ~n10742 & n10756 ;
  assign n10758 = ~n10745 & n10757 ;
  assign n10759 = ~n10748 & n10758 ;
  assign n10760 = n3450 & ~n10759 ;
  assign n10761 = ~n10736 & ~n10760 ;
  assign n10762 = \P1_state_reg[0]/NET0131  & ~n10761 ;
  assign n10763 = ~n10735 & ~n10762 ;
  assign n10764 = \P1_reg0_reg[2]/NET0131  & ~n3435 ;
  assign n10765 = \P1_reg0_reg[2]/NET0131  & n3448 ;
  assign n10767 = \P1_reg0_reg[2]/NET0131  & ~n4396 ;
  assign n10774 = n4396 & n10663 ;
  assign n10775 = ~n10767 & ~n10774 ;
  assign n10776 = n1936 & ~n10775 ;
  assign n10771 = n4396 & ~n10649 ;
  assign n10772 = ~n10767 & ~n10771 ;
  assign n10773 = ~n3563 & ~n10772 ;
  assign n10768 = n4396 & ~n10655 ;
  assign n10769 = ~n10767 & ~n10768 ;
  assign n10770 = ~n3677 & ~n10769 ;
  assign n10777 = n4396 & n10668 ;
  assign n10778 = ~n10767 & ~n10777 ;
  assign n10779 = n3712 & ~n10778 ;
  assign n10766 = n4396 & n10737 ;
  assign n10780 = \P1_reg0_reg[2]/NET0131  & ~n4493 ;
  assign n10781 = ~n10766 & ~n10780 ;
  assign n10782 = ~n10779 & n10781 ;
  assign n10783 = ~n10770 & n10782 ;
  assign n10784 = ~n10773 & n10783 ;
  assign n10785 = ~n10776 & n10784 ;
  assign n10786 = n3450 & ~n10785 ;
  assign n10787 = ~n10765 & ~n10786 ;
  assign n10788 = \P1_state_reg[0]/NET0131  & ~n10787 ;
  assign n10789 = ~n10764 & ~n10788 ;
  assign n10790 = \P1_reg1_reg[2]/NET0131  & ~n3435 ;
  assign n10791 = \P1_reg1_reg[2]/NET0131  & n3448 ;
  assign n10793 = \P1_reg1_reg[2]/NET0131  & ~n4532 ;
  assign n10800 = n4532 & n10663 ;
  assign n10801 = ~n10793 & ~n10800 ;
  assign n10802 = n1936 & ~n10801 ;
  assign n10797 = n4532 & ~n10649 ;
  assign n10798 = ~n10793 & ~n10797 ;
  assign n10799 = ~n3563 & ~n10798 ;
  assign n10794 = n4532 & ~n10655 ;
  assign n10795 = ~n10793 & ~n10794 ;
  assign n10796 = ~n3677 & ~n10795 ;
  assign n10803 = n4532 & n10668 ;
  assign n10804 = ~n10793 & ~n10803 ;
  assign n10805 = n3712 & ~n10804 ;
  assign n10792 = n4532 & n10737 ;
  assign n10806 = \P1_reg1_reg[2]/NET0131  & ~n4541 ;
  assign n10807 = ~n10792 & ~n10806 ;
  assign n10808 = ~n10805 & n10807 ;
  assign n10809 = ~n10796 & n10808 ;
  assign n10810 = ~n10799 & n10809 ;
  assign n10811 = ~n10802 & n10810 ;
  assign n10812 = n3450 & ~n10811 ;
  assign n10813 = ~n10791 & ~n10812 ;
  assign n10814 = \P1_state_reg[0]/NET0131  & ~n10813 ;
  assign n10815 = ~n10790 & ~n10814 ;
  assign n10816 = \P1_reg3_reg[1]/NET0131  & ~n3435 ;
  assign n10817 = \P1_reg3_reg[1]/NET0131  & n3448 ;
  assign n10822 = \P1_reg3_reg[1]/NET0131  & ~n3980 ;
  assign n10832 = n1595 & ~n3571 ;
  assign n10833 = ~n3572 & ~n10832 ;
  assign n10834 = ~n537 & ~n10833 ;
  assign n10835 = n537 & n1664 ;
  assign n10836 = ~n10834 & ~n10835 ;
  assign n10837 = n3980 & n10836 ;
  assign n10838 = ~n10822 & ~n10837 ;
  assign n10839 = n1936 & ~n10838 ;
  assign n10823 = n1792 & n3505 ;
  assign n10824 = ~n1792 & ~n3505 ;
  assign n10825 = ~n10823 & ~n10824 ;
  assign n10826 = ~n1671 & n10825 ;
  assign n10827 = n1671 & ~n1792 ;
  assign n10828 = ~n10826 & ~n10827 ;
  assign n10829 = n3980 & ~n10828 ;
  assign n10830 = ~n10822 & ~n10829 ;
  assign n10831 = ~n3677 & ~n10830 ;
  assign n10840 = n3980 & ~n10825 ;
  assign n10841 = ~n10822 & ~n10840 ;
  assign n10842 = ~n3563 & ~n10841 ;
  assign n10844 = \P1_reg3_reg[1]/NET0131  & ~n4910 ;
  assign n10818 = ~n1655 & ~n1671 ;
  assign n10819 = ~n3679 & ~n10818 ;
  assign n10820 = n3712 & n10819 ;
  assign n10821 = n3980 & n10820 ;
  assign n10843 = ~n1655 & ~n4067 ;
  assign n10845 = ~n10821 & ~n10843 ;
  assign n10846 = ~n10844 & n10845 ;
  assign n10847 = ~n10842 & n10846 ;
  assign n10848 = ~n10831 & n10847 ;
  assign n10849 = ~n10839 & n10848 ;
  assign n10850 = n3450 & ~n10849 ;
  assign n10851 = ~n10817 & ~n10850 ;
  assign n10852 = \P1_state_reg[0]/NET0131  & ~n10851 ;
  assign n10853 = ~n10816 & ~n10852 ;
  assign n10854 = \P2_reg3_reg[1]/NET0131  & ~n1983 ;
  assign n10855 = \P2_reg3_reg[1]/NET0131  & n2024 ;
  assign n10857 = \P2_reg3_reg[1]/NET0131  & ~n3788 ;
  assign n10867 = n2552 & ~n3374 ;
  assign n10868 = ~n3375 & ~n10867 ;
  assign n10869 = ~n2058 & ~n10868 ;
  assign n10870 = n2058 & n2597 ;
  assign n10871 = ~n10869 & ~n10870 ;
  assign n10872 = n3788 & n10871 ;
  assign n10873 = ~n10857 & ~n10872 ;
  assign n10874 = n3411 & ~n10873 ;
  assign n10858 = ~n2605 & n4199 ;
  assign n10859 = n2605 & ~n4199 ;
  assign n10860 = ~n10858 & ~n10859 ;
  assign n10861 = ~n2604 & ~n10860 ;
  assign n10862 = n2604 & ~n4199 ;
  assign n10863 = ~n10861 & ~n10862 ;
  assign n10864 = n3788 & ~n10863 ;
  assign n10865 = ~n10857 & ~n10864 ;
  assign n10866 = ~n3320 & ~n10865 ;
  assign n10875 = n3788 & n10860 ;
  assign n10876 = ~n10857 & ~n10875 ;
  assign n10877 = ~n3177 & ~n10876 ;
  assign n10856 = \P2_reg3_reg[1]/NET0131  & ~n5698 ;
  assign n10878 = ~n2588 & ~n3965 ;
  assign n10879 = ~n2588 & ~n2604 ;
  assign n10880 = ~n3326 & n3355 ;
  assign n10881 = ~n10879 & n10880 ;
  assign n10882 = n3788 & n10881 ;
  assign n10883 = ~n10878 & ~n10882 ;
  assign n10884 = ~n10856 & n10883 ;
  assign n10885 = ~n10877 & n10884 ;
  assign n10886 = ~n10866 & n10885 ;
  assign n10887 = ~n10874 & n10886 ;
  assign n10888 = n2026 & ~n10887 ;
  assign n10889 = ~n10855 & ~n10888 ;
  assign n10890 = \P1_state_reg[0]/NET0131  & ~n10889 ;
  assign n10891 = ~n10854 & ~n10890 ;
  assign n10892 = \P2_reg0_reg[1]/NET0131  & ~n1983 ;
  assign n10893 = \P2_reg0_reg[1]/NET0131  & n2024 ;
  assign n10897 = \P2_reg0_reg[1]/NET0131  & ~n2040 ;
  assign n10901 = n2040 & n10871 ;
  assign n10902 = ~n10897 & ~n10901 ;
  assign n10903 = n3411 & ~n10902 ;
  assign n10898 = n2040 & ~n10863 ;
  assign n10899 = ~n10897 & ~n10898 ;
  assign n10900 = ~n3320 & ~n10899 ;
  assign n10904 = n2040 & n10860 ;
  assign n10905 = ~n10897 & ~n10904 ;
  assign n10906 = ~n3177 & ~n10905 ;
  assign n10894 = ~n2588 & n3358 ;
  assign n10895 = ~n10881 & ~n10894 ;
  assign n10896 = n2040 & ~n10895 ;
  assign n10907 = \P2_reg0_reg[1]/NET0131  & ~n3425 ;
  assign n10908 = ~n10896 & ~n10907 ;
  assign n10909 = ~n10906 & n10908 ;
  assign n10910 = ~n10900 & n10909 ;
  assign n10911 = ~n10903 & n10910 ;
  assign n10912 = n2026 & ~n10911 ;
  assign n10913 = ~n10893 & ~n10912 ;
  assign n10914 = \P1_state_reg[0]/NET0131  & ~n10913 ;
  assign n10915 = ~n10892 & ~n10914 ;
  assign n10916 = \P2_reg1_reg[1]/NET0131  & ~n1983 ;
  assign n10917 = \P2_reg1_reg[1]/NET0131  & n2024 ;
  assign n10919 = \P2_reg1_reg[1]/NET0131  & ~n3733 ;
  assign n10923 = n3733 & n10871 ;
  assign n10924 = ~n10919 & ~n10923 ;
  assign n10925 = n3411 & ~n10924 ;
  assign n10920 = n3733 & ~n10863 ;
  assign n10921 = ~n10919 & ~n10920 ;
  assign n10922 = ~n3320 & ~n10921 ;
  assign n10926 = n3733 & n10860 ;
  assign n10927 = ~n10919 & ~n10926 ;
  assign n10928 = ~n3177 & ~n10927 ;
  assign n10918 = n3733 & ~n10895 ;
  assign n10929 = \P2_reg1_reg[1]/NET0131  & ~n7598 ;
  assign n10930 = ~n10918 & ~n10929 ;
  assign n10931 = ~n10928 & n10930 ;
  assign n10932 = ~n10922 & n10931 ;
  assign n10933 = ~n10925 & n10932 ;
  assign n10934 = n2026 & ~n10933 ;
  assign n10935 = ~n10917 & ~n10934 ;
  assign n10936 = \P1_state_reg[0]/NET0131  & ~n10935 ;
  assign n10937 = ~n10916 & ~n10936 ;
  assign n10938 = \P2_reg2_reg[2]/NET0131  & ~n1983 ;
  assign n10939 = \P2_reg2_reg[2]/NET0131  & n2024 ;
  assign n10941 = \P2_reg2_reg[2]/NET0131  & ~n3758 ;
  assign n10948 = n3758 & n10624 ;
  assign n10949 = ~n10941 & ~n10948 ;
  assign n10950 = n3411 & ~n10949 ;
  assign n10945 = n3758 & ~n10610 ;
  assign n10946 = ~n10941 & ~n10945 ;
  assign n10947 = ~n3177 & ~n10946 ;
  assign n10942 = n3758 & ~n10616 ;
  assign n10943 = ~n10941 & ~n10942 ;
  assign n10944 = ~n3320 & ~n10943 ;
  assign n10951 = n3758 & n10629 ;
  assign n10952 = ~n10941 & ~n10951 ;
  assign n10953 = n3355 & ~n10952 ;
  assign n10955 = \P2_reg2_reg[2]/NET0131  & ~n3774 ;
  assign n10940 = n3758 & n10684 ;
  assign n10954 = \P2_reg3_reg[2]/NET0131  & n3420 ;
  assign n10956 = ~n10940 & ~n10954 ;
  assign n10957 = ~n10955 & n10956 ;
  assign n10958 = ~n10953 & n10957 ;
  assign n10959 = ~n10944 & n10958 ;
  assign n10960 = ~n10947 & n10959 ;
  assign n10961 = ~n10950 & n10960 ;
  assign n10962 = n2026 & ~n10961 ;
  assign n10963 = ~n10939 & ~n10962 ;
  assign n10964 = \P1_state_reg[0]/NET0131  & ~n10963 ;
  assign n10965 = ~n10938 & ~n10964 ;
  assign n10966 = \P1_reg0_reg[1]/NET0131  & ~n3435 ;
  assign n10967 = \P1_reg0_reg[1]/NET0131  & n3448 ;
  assign n10969 = \P1_reg0_reg[1]/NET0131  & ~n4396 ;
  assign n10973 = n4396 & n10836 ;
  assign n10974 = ~n10969 & ~n10973 ;
  assign n10975 = n1936 & ~n10974 ;
  assign n10970 = n4396 & ~n10828 ;
  assign n10971 = ~n10969 & ~n10970 ;
  assign n10972 = ~n3677 & ~n10971 ;
  assign n10976 = n4396 & ~n10825 ;
  assign n10977 = ~n10969 & ~n10976 ;
  assign n10978 = ~n3563 & ~n10977 ;
  assign n10968 = \P1_reg0_reg[1]/NET0131  & ~n4494 ;
  assign n10979 = ~n1655 & n1880 ;
  assign n10980 = ~n10820 & ~n10979 ;
  assign n10981 = n4396 & ~n10980 ;
  assign n10982 = ~n10968 & ~n10981 ;
  assign n10983 = ~n10978 & n10982 ;
  assign n10984 = ~n10972 & n10983 ;
  assign n10985 = ~n10975 & n10984 ;
  assign n10986 = n3450 & ~n10985 ;
  assign n10987 = ~n10967 & ~n10986 ;
  assign n10988 = \P1_state_reg[0]/NET0131  & ~n10987 ;
  assign n10989 = ~n10966 & ~n10988 ;
  assign n10990 = \P1_reg1_reg[1]/NET0131  & ~n3435 ;
  assign n10991 = \P1_reg1_reg[1]/NET0131  & n3448 ;
  assign n10993 = \P1_reg1_reg[1]/NET0131  & ~n4532 ;
  assign n10997 = n4532 & n10836 ;
  assign n10998 = ~n10993 & ~n10997 ;
  assign n10999 = n1936 & ~n10998 ;
  assign n10994 = n4532 & ~n10828 ;
  assign n10995 = ~n10993 & ~n10994 ;
  assign n10996 = ~n3677 & ~n10995 ;
  assign n11000 = n4532 & ~n10825 ;
  assign n11001 = ~n10993 & ~n11000 ;
  assign n11002 = ~n3563 & ~n11001 ;
  assign n10992 = \P1_reg1_reg[1]/NET0131  & ~n4573 ;
  assign n11003 = n4532 & ~n10980 ;
  assign n11004 = ~n10992 & ~n11003 ;
  assign n11005 = ~n11002 & n11004 ;
  assign n11006 = ~n10996 & n11005 ;
  assign n11007 = ~n10999 & n11006 ;
  assign n11008 = n3450 & ~n11007 ;
  assign n11009 = ~n10991 & ~n11008 ;
  assign n11010 = \P1_state_reg[0]/NET0131  & ~n11009 ;
  assign n11011 = ~n10990 & ~n11010 ;
  assign n11012 = \P1_reg2_reg[1]/NET0131  & ~n3435 ;
  assign n11013 = \P1_reg2_reg[1]/NET0131  & n3448 ;
  assign n11015 = \P1_reg2_reg[1]/NET0131  & ~n3466 ;
  assign n11019 = n3466 & n10836 ;
  assign n11020 = ~n11015 & ~n11019 ;
  assign n11021 = n1936 & ~n11020 ;
  assign n11016 = n3466 & ~n10828 ;
  assign n11017 = ~n11015 & ~n11016 ;
  assign n11018 = ~n3677 & ~n11017 ;
  assign n11022 = n3466 & ~n10825 ;
  assign n11023 = ~n11015 & ~n11022 ;
  assign n11024 = ~n3563 & ~n11023 ;
  assign n11028 = n3466 & n10819 ;
  assign n11029 = ~n11015 & ~n11028 ;
  assign n11030 = n3712 & ~n11029 ;
  assign n11025 = ~n1655 & n3466 ;
  assign n11026 = ~n11015 & ~n11025 ;
  assign n11027 = n1880 & ~n11026 ;
  assign n11014 = \P1_reg3_reg[1]/NET0131  & n1763 ;
  assign n11031 = \P1_reg2_reg[1]/NET0131  & n3716 ;
  assign n11032 = ~n11014 & ~n11031 ;
  assign n11033 = ~n11027 & n11032 ;
  assign n11034 = ~n11030 & n11033 ;
  assign n11035 = ~n11024 & n11034 ;
  assign n11036 = ~n11018 & n11035 ;
  assign n11037 = ~n11021 & n11036 ;
  assign n11038 = n3450 & ~n11037 ;
  assign n11039 = ~n11013 & ~n11038 ;
  assign n11040 = \P1_state_reg[0]/NET0131  & ~n11039 ;
  assign n11041 = ~n11012 & ~n11040 ;
  assign n11042 = \P2_reg2_reg[1]/NET0131  & ~n1983 ;
  assign n11043 = \P2_reg2_reg[1]/NET0131  & n2024 ;
  assign n11045 = \P2_reg2_reg[1]/NET0131  & ~n3758 ;
  assign n11049 = n3758 & n10871 ;
  assign n11050 = ~n11045 & ~n11049 ;
  assign n11051 = n3411 & ~n11050 ;
  assign n11046 = n3758 & ~n10863 ;
  assign n11047 = ~n11045 & ~n11046 ;
  assign n11048 = ~n3320 & ~n11047 ;
  assign n11052 = n3758 & n10860 ;
  assign n11053 = ~n11045 & ~n11052 ;
  assign n11054 = ~n3177 & ~n11053 ;
  assign n11055 = \P2_reg2_reg[1]/NET0131  & ~n4383 ;
  assign n11044 = \P2_reg3_reg[1]/NET0131  & n3420 ;
  assign n11056 = n3758 & ~n10895 ;
  assign n11057 = ~n11044 & ~n11056 ;
  assign n11058 = ~n11055 & n11057 ;
  assign n11059 = ~n11054 & n11058 ;
  assign n11060 = ~n11048 & n11059 ;
  assign n11061 = ~n11051 & n11060 ;
  assign n11062 = n2026 & ~n11061 ;
  assign n11063 = ~n11043 & ~n11062 ;
  assign n11064 = \P1_state_reg[0]/NET0131  & ~n11063 ;
  assign n11065 = ~n11042 & ~n11064 ;
  assign n11066 = \P1_reg3_reg[0]/NET0131  & ~n3435 ;
  assign n11067 = \P1_reg3_reg[0]/NET0131  & n3448 ;
  assign n11069 = \P1_reg3_reg[0]/NET0131  & ~n3980 ;
  assign n11077 = n1641 & ~n3570 ;
  assign n11078 = ~n537 & ~n3571 ;
  assign n11079 = ~n11077 & n11078 ;
  assign n11080 = n3980 & n11079 ;
  assign n11081 = ~n11069 & ~n11080 ;
  assign n11082 = n1936 & ~n11081 ;
  assign n11076 = \P1_reg3_reg[0]/NET0131  & ~n9092 ;
  assign n11068 = ~n1765 & ~n1888 ;
  assign n11070 = ~n1804 & n3980 ;
  assign n11071 = ~n11069 & ~n11070 ;
  assign n11072 = ~n11068 & ~n11071 ;
  assign n11073 = ~n1761 & ~n3980 ;
  assign n11074 = ~n1671 & n1762 ;
  assign n11075 = ~n11073 & n11074 ;
  assign n11083 = ~n11072 & ~n11075 ;
  assign n11084 = ~n11076 & n11083 ;
  assign n11085 = ~n11082 & n11084 ;
  assign n11086 = n3450 & ~n11085 ;
  assign n11087 = ~n11067 & ~n11086 ;
  assign n11088 = \P1_state_reg[0]/NET0131  & ~n11087 ;
  assign n11089 = ~n11066 & ~n11088 ;
  assign n11090 = \P2_reg3_reg[0]/NET0131  & ~n1983 ;
  assign n11091 = \P2_reg3_reg[0]/NET0131  & n2024 ;
  assign n11093 = \P2_reg3_reg[0]/NET0131  & ~n3788 ;
  assign n11100 = n2574 & ~n3373 ;
  assign n11101 = ~n2058 & ~n3374 ;
  assign n11102 = ~n11100 & n11101 ;
  assign n11103 = n3788 & n11102 ;
  assign n11104 = ~n11093 & ~n11103 ;
  assign n11105 = n3411 & ~n11104 ;
  assign n11097 = ~n2604 & n3788 ;
  assign n11098 = ~n11093 & ~n11097 ;
  assign n11099 = n9903 & ~n11098 ;
  assign n11094 = n3788 & ~n4204 ;
  assign n11095 = ~n11093 & ~n11094 ;
  assign n11096 = ~n3744 & ~n11095 ;
  assign n11092 = \P2_reg3_reg[0]/NET0131  & n3417 ;
  assign n11106 = ~n2604 & n3420 ;
  assign n11107 = ~n11092 & ~n11106 ;
  assign n11108 = ~n11096 & n11107 ;
  assign n11109 = ~n11099 & n11108 ;
  assign n11110 = ~n11105 & n11109 ;
  assign n11111 = n2026 & ~n11110 ;
  assign n11112 = ~n11091 & ~n11111 ;
  assign n11113 = \P1_state_reg[0]/NET0131  & ~n11112 ;
  assign n11114 = ~n11090 & ~n11113 ;
  assign n11115 = ~\P1_reg2_reg[0]/NET0131  & ~n5812 ;
  assign n11117 = n1936 & n11079 ;
  assign n11118 = ~n1671 & n9090 ;
  assign n11119 = ~n1804 & ~n11068 ;
  assign n11120 = ~n11118 & ~n11119 ;
  assign n11121 = ~n11117 & n11120 ;
  assign n11122 = n3466 & ~n11121 ;
  assign n11116 = \P1_reg3_reg[0]/NET0131  & n1763 ;
  assign n11123 = ~n1936 & n11068 ;
  assign n11124 = ~n3466 & ~n11123 ;
  assign n11125 = n5815 & ~n9953 ;
  assign n11126 = ~n11124 & n11125 ;
  assign n11127 = \P1_reg2_reg[0]/NET0131  & ~n11126 ;
  assign n11128 = ~n11116 & ~n11127 ;
  assign n11129 = ~n11122 & n11128 ;
  assign n11130 = ~n11115 & ~n11129 ;
  assign n11131 = \P2_reg1_reg[0]/NET0131  & ~n1983 ;
  assign n11132 = \P2_reg1_reg[0]/NET0131  & n2024 ;
  assign n11133 = \P2_reg1_reg[0]/NET0131  & ~n3733 ;
  assign n11141 = n3733 & n11102 ;
  assign n11142 = ~n11133 & ~n11141 ;
  assign n11143 = n3411 & ~n11142 ;
  assign n11137 = n3733 & ~n4204 ;
  assign n11138 = ~n11133 & ~n11137 ;
  assign n11139 = ~n3744 & ~n11138 ;
  assign n11134 = ~n2604 & n3733 ;
  assign n11135 = ~n11133 & ~n11134 ;
  assign n11136 = n9903 & ~n11135 ;
  assign n11140 = \P2_reg1_reg[0]/NET0131  & ~n3421 ;
  assign n11144 = ~n11136 & ~n11140 ;
  assign n11145 = ~n11139 & n11144 ;
  assign n11146 = ~n11143 & n11145 ;
  assign n11147 = n2026 & ~n11146 ;
  assign n11148 = ~n11132 & ~n11147 ;
  assign n11149 = \P1_state_reg[0]/NET0131  & ~n11148 ;
  assign n11150 = ~n11131 & ~n11149 ;
  assign n11151 = \P2_reg3_reg[0]/NET0131  & n3420 ;
  assign n11154 = n3411 & n11102 ;
  assign n11152 = ~n3744 & ~n4204 ;
  assign n11153 = ~n2604 & n9903 ;
  assign n11155 = ~n11152 & ~n11153 ;
  assign n11156 = ~n11154 & n11155 ;
  assign n11157 = n3758 & ~n11156 ;
  assign n11158 = ~n11151 & ~n11157 ;
  assign n11159 = n5287 & ~n11158 ;
  assign n11160 = \P2_reg2_reg[0]/NET0131  & ~n10018 ;
  assign n11161 = ~n11159 & ~n11160 ;
  assign n11162 = \P1_reg0_reg[0]/NET0131  & ~n3435 ;
  assign n11163 = \P1_reg0_reg[0]/NET0131  & n3448 ;
  assign n11164 = \P1_reg0_reg[0]/NET0131  & ~n4396 ;
  assign n11172 = n4396 & n11079 ;
  assign n11173 = ~n11164 & ~n11172 ;
  assign n11174 = n1936 & ~n11173 ;
  assign n11168 = ~n1671 & n4396 ;
  assign n11169 = ~n11164 & ~n11168 ;
  assign n11170 = n9090 & ~n11169 ;
  assign n11165 = ~n1804 & n4396 ;
  assign n11166 = ~n11164 & ~n11165 ;
  assign n11167 = ~n11068 & ~n11166 ;
  assign n11171 = \P1_reg0_reg[0]/NET0131  & ~n4491 ;
  assign n11175 = ~n11167 & ~n11171 ;
  assign n11176 = ~n11170 & n11175 ;
  assign n11177 = ~n11174 & n11176 ;
  assign n11178 = n3450 & ~n11177 ;
  assign n11179 = ~n11163 & ~n11178 ;
  assign n11180 = \P1_state_reg[0]/NET0131  & ~n11179 ;
  assign n11181 = ~n11162 & ~n11180 ;
  assign n11182 = n6368 & ~n11121 ;
  assign n11183 = ~n4532 & ~n11123 ;
  assign n11184 = n5812 & ~n11183 ;
  assign n11185 = n9835 & n11184 ;
  assign n11186 = \P1_reg1_reg[0]/NET0131  & ~n11185 ;
  assign n11187 = ~n11182 & ~n11186 ;
  assign n11188 = \P2_reg0_reg[0]/NET0131  & ~n1983 ;
  assign n11189 = \P2_reg0_reg[0]/NET0131  & n2024 ;
  assign n11190 = \P2_reg0_reg[0]/NET0131  & ~n2040 ;
  assign n11198 = n2040 & n11102 ;
  assign n11199 = ~n11190 & ~n11198 ;
  assign n11200 = n3411 & ~n11199 ;
  assign n11194 = n2040 & ~n4204 ;
  assign n11195 = ~n11190 & ~n11194 ;
  assign n11196 = ~n3744 & ~n11195 ;
  assign n11191 = n2040 & ~n2604 ;
  assign n11192 = ~n11190 & ~n11191 ;
  assign n11193 = n9903 & ~n11192 ;
  assign n11197 = \P2_reg0_reg[0]/NET0131  & ~n3421 ;
  assign n11201 = ~n11193 & ~n11197 ;
  assign n11202 = ~n11196 & n11201 ;
  assign n11203 = ~n11200 & n11202 ;
  assign n11204 = n2026 & ~n11203 ;
  assign n11205 = ~n11189 & ~n11204 ;
  assign n11206 = \P1_state_reg[0]/NET0131  & ~n11205 ;
  assign n11207 = ~n11188 & ~n11206 ;
  assign n11208 = ~\P1_state_reg[0]/NET0131  & ~n1028 ;
  assign n11209 = \P1_state_reg[0]/NET0131  & ~n3439 ;
  assign n11210 = ~n11208 & ~n11209 ;
  assign n11211 = ~\P1_state_reg[0]/NET0131  & ~n996 ;
  assign n11212 = \P1_state_reg[0]/NET0131  & ~n3442 ;
  assign n11213 = ~n11211 & ~n11212 ;
  assign n11214 = ~\P1_state_reg[0]/NET0131  & ~n968 ;
  assign n11215 = \P1_state_reg[0]/NET0131  & n527 ;
  assign n11216 = ~n11214 & ~n11215 ;
  assign n11217 = ~\P1_state_reg[0]/NET0131  & ~n3033 ;
  assign n11218 = \P1_state_reg[0]/NET0131  & n2022 ;
  assign n11219 = ~n11217 & ~n11218 ;
  assign n11220 = ~\P1_state_reg[0]/NET0131  & ~n3011 ;
  assign n11221 = \P1_state_reg[0]/NET0131  & n2001 ;
  assign n11222 = ~n11220 & ~n11221 ;
  assign n11223 = ~\P1_state_reg[0]/NET0131  & ~n2981 ;
  assign n11224 = \P1_state_reg[0]/NET0131  & n2051 ;
  assign n11225 = ~n11223 & ~n11224 ;
  assign n11226 = ~\P1_state_reg[0]/NET0131  & ~n2753 ;
  assign n11227 = \P1_state_reg[0]/NET0131  & ~n2745 ;
  assign n11228 = ~n11226 & ~n11227 ;
  assign n11229 = \P1_state_reg[0]/NET0131  & ~n2694 ;
  assign n11230 = ~\P1_state_reg[0]/NET0131  & n2702 ;
  assign n11231 = ~n11229 & ~n11230 ;
  assign n11232 = \P1_state_reg[0]/NET0131  & ~n2720 ;
  assign n11233 = ~\P1_state_reg[0]/NET0131  & n2729 ;
  assign n11234 = ~n11232 & ~n11233 ;
  assign n11235 = ~\P1_state_reg[0]/NET0131  & ~n2891 ;
  assign n11236 = \P1_state_reg[0]/NET0131  & ~n2883 ;
  assign n11237 = ~n11235 & ~n11236 ;
  assign n11238 = \P1_state_reg[0]/NET0131  & ~n2849 ;
  assign n11239 = ~\P1_state_reg[0]/NET0131  & n2858 ;
  assign n11240 = ~n11238 & ~n11239 ;
  assign n11241 = ~\P1_state_reg[0]/NET0131  & ~n2841 ;
  assign n11242 = \P1_state_reg[0]/NET0131  & n2832 ;
  assign n11243 = ~n11241 & ~n11242 ;
  assign n11244 = \P1_state_reg[0]/NET0131  & ~n2808 ;
  assign n11245 = ~\P1_state_reg[0]/NET0131  & n2816 ;
  assign n11246 = ~n11244 & ~n11245 ;
  assign n11247 = \P1_state_reg[0]/NET0131  & ~n2385 ;
  assign n11248 = ~\P1_state_reg[0]/NET0131  & n2397 ;
  assign n11249 = ~n11247 & ~n11248 ;
  assign n11250 = \P1_state_reg[0]/NET0131  & ~n2404 ;
  assign n11251 = ~\P1_state_reg[0]/NET0131  & n2431 ;
  assign n11252 = ~n11250 & ~n11251 ;
  assign n11253 = ~\P1_state_reg[0]/NET0131  & ~n2297 ;
  assign n11254 = \P1_state_reg[0]/NET0131  & n2258 ;
  assign n11255 = ~n11253 & ~n11254 ;
  assign n11256 = \P1_state_reg[0]/NET0131  & n2578 ;
  assign n11257 = ~\P1_state_reg[0]/NET0131  & n2586 ;
  assign n11258 = ~n11256 & ~n11257 ;
  assign n11259 = ~\P1_state_reg[0]/NET0131  & ~n2357 ;
  assign n11260 = \P1_state_reg[0]/NET0131  & ~n3175 ;
  assign n11261 = ~n11259 & ~n11260 ;
  assign n11262 = ~\P1_state_reg[0]/NET0131  & ~n3120 ;
  assign n11263 = \P1_state_reg[0]/NET0131  & ~n3170 ;
  assign n11264 = ~n11262 & ~n11263 ;
  assign n11265 = ~\P1_state_reg[0]/NET0131  & ~n3101 ;
  assign n11266 = \P1_state_reg[0]/NET0131  & n3166 ;
  assign n11267 = ~n11265 & ~n11266 ;
  assign n11268 = ~\P1_state_reg[0]/NET0131  & ~n3078 ;
  assign n11269 = ~n3976 & ~n11268 ;
  assign n11270 = ~\P1_state_reg[0]/NET0131  & ~n3053 ;
  assign n11271 = \P1_state_reg[0]/NET0131  & n2008 ;
  assign n11272 = ~n11270 & ~n11271 ;
  assign n11273 = \P1_state_reg[0]/NET0131  & ~n2215 ;
  assign n11274 = ~\P1_state_reg[0]/NET0131  & n2197 ;
  assign n11275 = ~n11273 & ~n11274 ;
  assign n11276 = ~\P1_state_reg[0]/NET0131  & ~n2559 ;
  assign n11277 = \P1_state_reg[0]/NET0131  & n2564 ;
  assign n11278 = ~n11276 & ~n11277 ;
  assign n11279 = ~\P1_state_reg[0]/NET0131  & ~n4158 ;
  assign n11280 = \P1_state_reg[0]/NET0131  & n2207 ;
  assign n11281 = ~n11279 & ~n11280 ;
  assign n11282 = \P1_state_reg[0]/NET0131  & ~n2629 ;
  assign n11283 = ~\P1_state_reg[0]/NET0131  & n2623 ;
  assign n11284 = ~n11282 & ~n11283 ;
  assign n11285 = \P1_state_reg[0]/NET0131  & n2646 ;
  assign n11286 = ~\P1_state_reg[0]/NET0131  & n2654 ;
  assign n11287 = ~n11285 & ~n11286 ;
  assign n11288 = ~\P1_state_reg[0]/NET0131  & ~n2538 ;
  assign n11289 = \P1_state_reg[0]/NET0131  & ~n2542 ;
  assign n11290 = ~n11288 & ~n11289 ;
  assign n11291 = ~\P1_state_reg[0]/NET0131  & ~n2513 ;
  assign n11292 = \P1_state_reg[0]/NET0131  & n2519 ;
  assign n11293 = ~n11291 & ~n11292 ;
  assign n11294 = \P1_state_reg[0]/NET0131  & ~n2485 ;
  assign n11295 = ~\P1_state_reg[0]/NET0131  & n2493 ;
  assign n11296 = ~n11294 & ~n11295 ;
  assign n11297 = \P1_state_reg[0]/NET0131  & ~n2460 ;
  assign n11298 = ~\P1_state_reg[0]/NET0131  & n2468 ;
  assign n11299 = ~n11297 & ~n11298 ;
  assign n11300 = ~\P1_state_reg[0]/NET0131  & ~n2777 ;
  assign n11301 = \P1_state_reg[0]/NET0131  & ~n2769 ;
  assign n11302 = ~n11300 & ~n11301 ;
  assign n11303 = ~\P1_state_reg[0]/NET0131  & ~n2948 ;
  assign n11304 = \P1_state_reg[0]/NET0131  & n2058 ;
  assign n11305 = ~n11303 & ~n11304 ;
  assign n11306 = \P1_state_reg[0]/NET0131  & ~n1223 ;
  assign n11307 = ~\P1_state_reg[0]/NET0131  & n1231 ;
  assign n11308 = ~n11306 & ~n11307 ;
  assign n11309 = ~\P1_state_reg[0]/NET0131  & ~n1196 ;
  assign n11310 = \P1_state_reg[0]/NET0131  & n1188 ;
  assign n11311 = ~n11309 & ~n11310 ;
  assign n11312 = \P1_state_reg[0]/NET0131  & ~n1154 ;
  assign n11313 = ~\P1_state_reg[0]/NET0131  & n1163 ;
  assign n11314 = ~n11312 & ~n11313 ;
  assign n11315 = \P1_state_reg[0]/NET0131  & ~n1126 ;
  assign n11316 = ~\P1_state_reg[0]/NET0131  & n1134 ;
  assign n11317 = ~n11315 & ~n11316 ;
  assign n11318 = ~\P1_state_reg[0]/NET0131  & ~n1107 ;
  assign n11319 = \P1_state_reg[0]/NET0131  & n1099 ;
  assign n11320 = ~n11318 & ~n11319 ;
  assign n11321 = ~\P1_state_reg[0]/NET0131  & ~n1081 ;
  assign n11322 = \P1_state_reg[0]/NET0131  & n1073 ;
  assign n11323 = ~n11321 & ~n11322 ;
  assign n11324 = ~\P1_state_reg[0]/NET0131  & ~n1464 ;
  assign n11325 = \P1_state_reg[0]/NET0131  & n1456 ;
  assign n11326 = ~n11324 & ~n11325 ;
  assign n11327 = ~\P1_state_reg[0]/NET0131  & ~n1441 ;
  assign n11328 = \P1_state_reg[0]/NET0131  & ~n1433 ;
  assign n11329 = ~n11327 & ~n11328 ;
  assign n11330 = \P1_state_reg[0]/NET0131  & ~n1384 ;
  assign n11331 = ~\P1_state_reg[0]/NET0131  & n1392 ;
  assign n11332 = ~n11330 & ~n11331 ;
  assign n11333 = ~\P1_state_reg[0]/NET0131  & ~n1416 ;
  assign n11334 = \P1_state_reg[0]/NET0131  & n1408 ;
  assign n11335 = ~n11333 & ~n11334 ;
  assign n11336 = \P1_state_reg[0]/NET0131  & n1645 ;
  assign n11337 = ~\P1_state_reg[0]/NET0131  & n1653 ;
  assign n11338 = ~n11336 & ~n11337 ;
  assign n11339 = \P1_state_reg[0]/NET0131  & ~n519 ;
  assign n11340 = ~\P1_state_reg[0]/NET0131  & n1364 ;
  assign n11341 = ~n11339 & ~n11340 ;
  assign n11342 = ~\P1_state_reg[0]/NET0131  & ~n1345 ;
  assign n11343 = \P1_state_reg[0]/NET0131  & n501 ;
  assign n11344 = ~n11342 & ~n11343 ;
  assign n11345 = ~\P1_state_reg[0]/NET0131  & ~n1326 ;
  assign n11346 = ~n1953 & ~n11345 ;
  assign n11347 = ~\P1_state_reg[0]/NET0131  & ~n1046 ;
  assign n11348 = \P1_state_reg[0]/NET0131  & n3445 ;
  assign n11349 = ~n11347 & ~n11348 ;
  assign n11350 = ~\P1_state_reg[0]/NET0131  & ~n1308 ;
  assign n11351 = \P1_state_reg[0]/NET0131  & n486 ;
  assign n11352 = ~n11350 & ~n11351 ;
  assign n11353 = ~\P1_state_reg[0]/NET0131  & ~n932 ;
  assign n11354 = \P1_state_reg[0]/NET0131  & n537 ;
  assign n11355 = ~n11353 & ~n11354 ;
  assign n11356 = ~\P1_state_reg[0]/NET0131  & ~n880 ;
  assign n11357 = \P1_state_reg[0]/NET0131  & n714 ;
  assign n11358 = ~n11356 & ~n11357 ;
  assign n11359 = ~\P1_state_reg[0]/NET0131  & ~n1602 ;
  assign n11360 = \P1_state_reg[0]/NET0131  & n1607 ;
  assign n11361 = ~n11359 & ~n11360 ;
  assign n11362 = ~\P1_state_reg[0]/NET0131  & ~n824 ;
  assign n11363 = \P1_state_reg[0]/NET0131  & n704 ;
  assign n11364 = ~n11362 & ~n11363 ;
  assign n11365 = ~\P1_state_reg[0]/NET0131  & n691 ;
  assign n11366 = ~\P1_IR_reg[30]/NET0131  & \P1_IR_reg[31]/NET0131  ;
  assign n11367 = \P1_state_reg[0]/NET0131  & n11366 ;
  assign n11368 = n698 & n11367 ;
  assign n11369 = n523 & n11368 ;
  assign n11370 = ~n11365 & ~n11369 ;
  assign n11371 = \P1_state_reg[0]/NET0131  & ~n1621 ;
  assign n11372 = ~\P1_state_reg[0]/NET0131  & n1630 ;
  assign n11373 = ~n11371 & ~n11372 ;
  assign n11374 = ~\P1_state_reg[0]/NET0131  & ~n1579 ;
  assign n11375 = \P1_state_reg[0]/NET0131  & ~n1584 ;
  assign n11376 = ~n11374 & ~n11375 ;
  assign n11377 = ~\P1_state_reg[0]/NET0131  & ~n1555 ;
  assign n11378 = \P1_state_reg[0]/NET0131  & ~n1560 ;
  assign n11379 = ~n11377 & ~n11378 ;
  assign n11380 = ~\P1_state_reg[0]/NET0131  & ~n1531 ;
  assign n11381 = \P1_state_reg[0]/NET0131  & ~n1535 ;
  assign n11382 = ~n11380 & ~n11381 ;
  assign n11383 = ~\P1_state_reg[0]/NET0131  & ~n1505 ;
  assign n11384 = \P1_state_reg[0]/NET0131  & n1512 ;
  assign n11385 = ~n11383 & ~n11384 ;
  assign n11386 = ~\P1_state_reg[0]/NET0131  & ~n1279 ;
  assign n11387 = \P1_state_reg[0]/NET0131  & n1271 ;
  assign n11388 = ~n11386 & ~n11387 ;
  assign n11389 = ~\P1_state_reg[0]/NET0131  & ~n1255 ;
  assign n11390 = \P1_state_reg[0]/NET0131  & n1247 ;
  assign n11391 = ~n11389 & ~n11390 ;
  assign n11392 = ~\P1_state_reg[0]/NET0131  & n4140 ;
  assign n11393 = \P1_state_reg[0]/NET0131  & ~\P2_IR_reg[30]/NET0131  ;
  assign n11394 = \P2_IR_reg[31]/NET0131  & n11393 ;
  assign n11395 = n2044 & n11394 ;
  assign n11396 = n2201 & n11395 ;
  assign n11397 = n1978 & n11396 ;
  assign n11398 = ~n11392 & ~n11397 ;
  assign n11438 = \P1_reg2_reg[7]/NET0131  & n1512 ;
  assign n11439 = ~\P1_reg2_reg[7]/NET0131  & ~n1512 ;
  assign n11440 = ~n11438 & ~n11439 ;
  assign n11441 = \P1_reg2_reg[6]/NET0131  & ~n1535 ;
  assign n11442 = ~\P1_reg2_reg[6]/NET0131  & n1535 ;
  assign n11443 = \P1_reg2_reg[5]/NET0131  & ~n1560 ;
  assign n11444 = \P1_reg2_reg[4]/NET0131  & ~n1584 ;
  assign n11445 = ~\P1_reg2_reg[3]/NET0131  & n1621 ;
  assign n11446 = \P1_reg2_reg[3]/NET0131  & ~n1621 ;
  assign n11447 = ~\P1_reg2_reg[2]/NET0131  & ~n1607 ;
  assign n11448 = \P1_reg2_reg[2]/NET0131  & n1607 ;
  assign n11449 = ~\P1_reg2_reg[1]/NET0131  & ~n1645 ;
  assign n11450 = \P1_reg2_reg[1]/NET0131  & n1645 ;
  assign n11451 = \P1_IR_reg[0]/NET0131  & \P1_reg2_reg[0]/NET0131  ;
  assign n11452 = ~n11450 & ~n11451 ;
  assign n11453 = ~n11449 & ~n11452 ;
  assign n11454 = ~n11448 & ~n11453 ;
  assign n11455 = ~n11447 & ~n11454 ;
  assign n11456 = ~n11446 & ~n11455 ;
  assign n11457 = ~n11445 & ~n11456 ;
  assign n11458 = ~n11444 & ~n11457 ;
  assign n11459 = ~\P1_reg2_reg[5]/NET0131  & n1560 ;
  assign n11460 = ~\P1_reg2_reg[4]/NET0131  & n1584 ;
  assign n11461 = ~n11459 & ~n11460 ;
  assign n11462 = ~n11458 & n11461 ;
  assign n11463 = ~n11443 & ~n11462 ;
  assign n11464 = ~n11442 & ~n11463 ;
  assign n11465 = ~n11441 & ~n11464 ;
  assign n11467 = n11440 & ~n11465 ;
  assign n11437 = n527 & n537 ;
  assign n11466 = ~n11440 & n11465 ;
  assign n11468 = n11437 & ~n11466 ;
  assign n11469 = ~n11467 & n11468 ;
  assign n11399 = ~n527 & ~n3448 ;
  assign n11401 = ~n1512 & ~n11399 ;
  assign n11400 = ~\P1_addr_reg[7]/NET0131  & n11399 ;
  assign n11402 = ~n537 & ~n11400 ;
  assign n11403 = ~n11401 & n11402 ;
  assign n11405 = \P1_reg1_reg[7]/NET0131  & n1512 ;
  assign n11406 = ~\P1_reg1_reg[7]/NET0131  & ~n1512 ;
  assign n11407 = ~n11405 & ~n11406 ;
  assign n11408 = \P1_reg1_reg[6]/NET0131  & ~n1535 ;
  assign n11409 = ~\P1_reg1_reg[6]/NET0131  & n1535 ;
  assign n11410 = \P1_reg1_reg[5]/NET0131  & ~n1560 ;
  assign n11411 = \P1_reg1_reg[4]/NET0131  & ~n1584 ;
  assign n11412 = ~\P1_reg1_reg[3]/NET0131  & n1621 ;
  assign n11413 = \P1_reg1_reg[3]/NET0131  & ~n1621 ;
  assign n11414 = ~\P1_reg1_reg[2]/NET0131  & ~n1607 ;
  assign n11415 = \P1_reg1_reg[2]/NET0131  & n1607 ;
  assign n11416 = ~\P1_reg1_reg[1]/NET0131  & ~n1645 ;
  assign n11417 = \P1_reg1_reg[1]/NET0131  & n1645 ;
  assign n11418 = \P1_IR_reg[0]/NET0131  & \P1_reg1_reg[0]/NET0131  ;
  assign n11419 = ~n11417 & ~n11418 ;
  assign n11420 = ~n11416 & ~n11419 ;
  assign n11421 = ~n11415 & ~n11420 ;
  assign n11422 = ~n11414 & ~n11421 ;
  assign n11423 = ~n11413 & ~n11422 ;
  assign n11424 = ~n11412 & ~n11423 ;
  assign n11425 = ~n11411 & ~n11424 ;
  assign n11426 = ~\P1_reg1_reg[5]/NET0131  & n1560 ;
  assign n11427 = ~\P1_reg1_reg[4]/NET0131  & n1584 ;
  assign n11428 = ~n11426 & ~n11427 ;
  assign n11429 = ~n11425 & n11428 ;
  assign n11430 = ~n11410 & ~n11429 ;
  assign n11431 = ~n11409 & ~n11430 ;
  assign n11432 = ~n11408 & ~n11431 ;
  assign n11434 = n11407 & ~n11432 ;
  assign n11404 = ~n527 & n537 ;
  assign n11433 = ~n11407 & n11432 ;
  assign n11435 = n11404 & ~n11433 ;
  assign n11436 = ~n11434 & n11435 ;
  assign n11470 = ~n11403 & ~n11436 ;
  assign n11471 = ~n11469 & n11470 ;
  assign n11472 = \P1_state_reg[0]/NET0131  & ~n11471 ;
  assign n11473 = ~n9781 & ~n11472 ;
  assign n11491 = ~\P1_reg2_reg[9]/NET0131  & ~n1247 ;
  assign n11492 = \P1_reg2_reg[9]/NET0131  & n1247 ;
  assign n11493 = ~n11491 & ~n11492 ;
  assign n11494 = ~\P1_reg2_reg[8]/NET0131  & ~n1271 ;
  assign n11495 = ~n11439 & ~n11465 ;
  assign n11496 = \P1_reg2_reg[8]/NET0131  & n1271 ;
  assign n11497 = ~n11438 & ~n11496 ;
  assign n11498 = ~n11495 & n11497 ;
  assign n11499 = ~n11494 & ~n11498 ;
  assign n11501 = n11493 & n11499 ;
  assign n11500 = ~n11493 & ~n11499 ;
  assign n11502 = n11437 & ~n11500 ;
  assign n11503 = ~n11501 & n11502 ;
  assign n11475 = ~n1247 & ~n11399 ;
  assign n11474 = ~\P1_addr_reg[9]/NET0131  & n11399 ;
  assign n11476 = ~n537 & ~n11474 ;
  assign n11477 = ~n11475 & n11476 ;
  assign n11478 = ~\P1_reg1_reg[8]/NET0131  & ~n1271 ;
  assign n11479 = ~n11406 & ~n11432 ;
  assign n11480 = \P1_reg1_reg[8]/NET0131  & n1271 ;
  assign n11481 = ~n11405 & ~n11480 ;
  assign n11482 = ~n11479 & n11481 ;
  assign n11483 = ~n11478 & ~n11482 ;
  assign n11484 = \P1_reg1_reg[9]/NET0131  & n1247 ;
  assign n11485 = ~\P1_reg1_reg[9]/NET0131  & ~n1247 ;
  assign n11486 = ~n11484 & ~n11485 ;
  assign n11488 = n11483 & n11486 ;
  assign n11487 = ~n11483 & ~n11486 ;
  assign n11489 = n11404 & ~n11487 ;
  assign n11490 = ~n11488 & n11489 ;
  assign n11504 = ~n11477 & ~n11490 ;
  assign n11505 = ~n11503 & n11504 ;
  assign n11506 = \P1_state_reg[0]/NET0131  & ~n11505 ;
  assign n11507 = ~n7281 & ~n11506 ;
  assign n11519 = n1535 & ~n11399 ;
  assign n11518 = ~\P1_addr_reg[6]/NET0131  & n11399 ;
  assign n11520 = ~n537 & ~n11518 ;
  assign n11521 = ~n11519 & n11520 ;
  assign n11508 = ~n11408 & ~n11409 ;
  assign n11510 = ~n11430 & n11508 ;
  assign n11509 = n11430 & ~n11508 ;
  assign n11511 = n11404 & ~n11509 ;
  assign n11512 = ~n11510 & n11511 ;
  assign n11513 = ~n11441 & ~n11442 ;
  assign n11515 = ~n11463 & n11513 ;
  assign n11514 = n11463 & ~n11513 ;
  assign n11516 = n11437 & ~n11514 ;
  assign n11517 = ~n11515 & n11516 ;
  assign n11522 = ~n11512 & ~n11517 ;
  assign n11523 = ~n11521 & n11522 ;
  assign n11524 = \P1_state_reg[0]/NET0131  & ~n11523 ;
  assign n11525 = ~n9740 & ~n11524 ;
  assign n11526 = \P1_reg3_reg[2]/NET0131  & ~\P1_state_reg[0]/NET0131  ;
  assign n11530 = ~n1607 & n3448 ;
  assign n11529 = ~\P1_addr_reg[2]/NET0131  & ~n3448 ;
  assign n11531 = n538 & ~n11529 ;
  assign n11532 = ~n11530 & n11531 ;
  assign n11538 = ~n11414 & ~n11415 ;
  assign n11539 = ~n11420 & ~n11538 ;
  assign n11540 = n11420 & n11538 ;
  assign n11541 = ~n11539 & ~n11540 ;
  assign n11542 = n11404 & n11541 ;
  assign n11527 = n527 & ~n537 ;
  assign n11528 = n1607 & n11527 ;
  assign n11533 = ~n11447 & ~n11448 ;
  assign n11534 = ~n11453 & ~n11533 ;
  assign n11535 = n11453 & n11533 ;
  assign n11536 = ~n11534 & ~n11535 ;
  assign n11537 = n11437 & n11536 ;
  assign n11543 = ~n11528 & ~n11537 ;
  assign n11544 = ~n11542 & n11543 ;
  assign n11545 = ~n11532 & n11544 ;
  assign n11546 = \P1_state_reg[0]/NET0131  & ~n11545 ;
  assign n11547 = ~n11526 & ~n11546 ;
  assign n11550 = n1621 & n3448 ;
  assign n11549 = ~\P1_addr_reg[3]/NET0131  & ~n3448 ;
  assign n11551 = n538 & ~n11549 ;
  assign n11552 = ~n11550 & n11551 ;
  assign n11558 = ~n11445 & ~n11446 ;
  assign n11559 = ~n11455 & ~n11558 ;
  assign n11560 = n11455 & n11558 ;
  assign n11561 = ~n11559 & ~n11560 ;
  assign n11562 = n11437 & n11561 ;
  assign n11548 = ~n1621 & n11527 ;
  assign n11553 = ~n11412 & ~n11413 ;
  assign n11554 = ~n11422 & ~n11553 ;
  assign n11555 = n11422 & n11553 ;
  assign n11556 = ~n11554 & ~n11555 ;
  assign n11557 = n11404 & n11556 ;
  assign n11563 = ~n11548 & ~n11557 ;
  assign n11564 = ~n11562 & n11563 ;
  assign n11565 = ~n11552 & n11564 ;
  assign n11566 = \P1_state_reg[0]/NET0131  & ~n11565 ;
  assign n11567 = ~n9696 & ~n11566 ;
  assign n11593 = \P1_reg1_reg[13]/NET0131  & n1126 ;
  assign n11594 = ~\P1_reg1_reg[13]/NET0131  & ~n1126 ;
  assign n11595 = ~n11593 & ~n11594 ;
  assign n11596 = ~\P1_reg1_reg[12]/NET0131  & ~n1154 ;
  assign n11597 = ~\P1_reg1_reg[11]/NET0131  & ~n1188 ;
  assign n11598 = ~\P1_reg1_reg[10]/NET0131  & ~n1223 ;
  assign n11599 = n11483 & ~n11485 ;
  assign n11600 = \P1_reg1_reg[10]/NET0131  & n1223 ;
  assign n11601 = ~n11484 & ~n11600 ;
  assign n11602 = ~n11599 & n11601 ;
  assign n11603 = ~n11598 & ~n11602 ;
  assign n11604 = ~n11597 & n11603 ;
  assign n11605 = \P1_reg1_reg[12]/NET0131  & n1154 ;
  assign n11606 = \P1_reg1_reg[11]/NET0131  & n1188 ;
  assign n11607 = ~n11605 & ~n11606 ;
  assign n11608 = ~n11604 & n11607 ;
  assign n11609 = ~n11596 & ~n11608 ;
  assign n11611 = n11595 & n11609 ;
  assign n11610 = ~n11595 & ~n11609 ;
  assign n11612 = n11404 & ~n11610 ;
  assign n11613 = ~n11611 & n11612 ;
  assign n11568 = \P1_reg2_reg[13]/NET0131  & n1126 ;
  assign n11569 = ~\P1_reg2_reg[13]/NET0131  & ~n1126 ;
  assign n11570 = ~n11568 & ~n11569 ;
  assign n11571 = ~\P1_reg2_reg[12]/NET0131  & ~n1154 ;
  assign n11572 = ~\P1_reg2_reg[11]/NET0131  & ~n1188 ;
  assign n11573 = ~\P1_reg2_reg[10]/NET0131  & ~n1223 ;
  assign n11574 = ~n11491 & n11499 ;
  assign n11575 = \P1_reg2_reg[10]/NET0131  & n1223 ;
  assign n11576 = ~n11492 & ~n11575 ;
  assign n11577 = ~n11574 & n11576 ;
  assign n11578 = ~n11573 & ~n11577 ;
  assign n11579 = ~n11572 & n11578 ;
  assign n11580 = \P1_reg2_reg[12]/NET0131  & n1154 ;
  assign n11581 = \P1_reg2_reg[11]/NET0131  & n1188 ;
  assign n11582 = ~n11580 & ~n11581 ;
  assign n11583 = ~n11579 & n11582 ;
  assign n11584 = ~n11571 & ~n11583 ;
  assign n11586 = n11570 & n11584 ;
  assign n11585 = ~n11570 & ~n11584 ;
  assign n11587 = n11437 & ~n11585 ;
  assign n11588 = ~n11586 & n11587 ;
  assign n11590 = ~n1126 & ~n11399 ;
  assign n11589 = ~\P1_addr_reg[13]/NET0131  & n11399 ;
  assign n11591 = ~n537 & ~n11589 ;
  assign n11592 = ~n11590 & n11591 ;
  assign n11614 = ~n11588 & ~n11592 ;
  assign n11615 = ~n11613 & n11614 ;
  assign n11616 = \P1_state_reg[0]/NET0131  & ~n11615 ;
  assign n11617 = ~n7113 & ~n11616 ;
  assign n11618 = ~\P1_state_reg[0]/NET0131  & \P2_reg3_reg[0]/NET0131  ;
  assign n11622 = ~\P2_IR_reg[0]/NET0131  & n2024 ;
  assign n11621 = ~\P2_addr_reg[0]/NET0131  & ~n2024 ;
  assign n11623 = n2059 & ~n11621 ;
  assign n11624 = ~n11622 & n11623 ;
  assign n11630 = n2051 & n2058 ;
  assign n11631 = ~\P2_IR_reg[0]/NET0131  & ~\P2_reg2_reg[0]/NET0131  ;
  assign n11632 = \P2_IR_reg[0]/NET0131  & \P2_reg2_reg[0]/NET0131  ;
  assign n11633 = ~n11631 & ~n11632 ;
  assign n11634 = n11630 & n11633 ;
  assign n11619 = n2051 & ~n2058 ;
  assign n11620 = \P2_IR_reg[0]/NET0131  & n11619 ;
  assign n11626 = ~n2051 & n2058 ;
  assign n11625 = ~\P2_IR_reg[0]/NET0131  & ~\P2_reg1_reg[0]/NET0131  ;
  assign n11627 = \P2_IR_reg[0]/NET0131  & \P2_reg1_reg[0]/NET0131  ;
  assign n11628 = ~n11625 & ~n11627 ;
  assign n11629 = n11626 & n11628 ;
  assign n11635 = ~n11620 & ~n11629 ;
  assign n11636 = ~n11634 & n11635 ;
  assign n11637 = ~n11624 & n11636 ;
  assign n11638 = \P1_state_reg[0]/NET0131  & ~n11637 ;
  assign n11639 = ~n11618 & ~n11638 ;
  assign n11640 = \P1_reg3_reg[0]/NET0131  & ~\P1_state_reg[0]/NET0131  ;
  assign n11643 = ~\P1_IR_reg[0]/NET0131  & n3448 ;
  assign n11642 = ~\P1_addr_reg[0]/NET0131  & ~n3448 ;
  assign n11644 = n538 & ~n11642 ;
  assign n11645 = ~n11643 & n11644 ;
  assign n11649 = ~\P1_IR_reg[0]/NET0131  & ~\P1_reg2_reg[0]/NET0131  ;
  assign n11650 = ~n11451 & ~n11649 ;
  assign n11651 = n11437 & n11650 ;
  assign n11641 = \P1_IR_reg[0]/NET0131  & n11527 ;
  assign n11646 = ~\P1_IR_reg[0]/NET0131  & ~\P1_reg1_reg[0]/NET0131  ;
  assign n11647 = ~n11418 & ~n11646 ;
  assign n11648 = n11404 & n11647 ;
  assign n11652 = ~n11641 & ~n11648 ;
  assign n11653 = ~n11651 & n11652 ;
  assign n11654 = ~n11645 & n11653 ;
  assign n11655 = \P1_state_reg[0]/NET0131  & ~n11654 ;
  assign n11656 = ~n11640 & ~n11655 ;
  assign n11671 = ~n11573 & ~n11575 ;
  assign n11672 = ~n11438 & ~n11495 ;
  assign n11673 = ~n11494 & ~n11672 ;
  assign n11674 = ~n11492 & ~n11496 ;
  assign n11675 = ~n11673 & n11674 ;
  assign n11676 = ~n11491 & ~n11675 ;
  assign n11678 = n11671 & n11676 ;
  assign n11677 = ~n11671 & ~n11676 ;
  assign n11679 = n11437 & ~n11677 ;
  assign n11680 = ~n11678 & n11679 ;
  assign n11658 = ~n1223 & ~n11399 ;
  assign n11657 = ~\P1_addr_reg[10]/NET0131  & n11399 ;
  assign n11659 = ~n537 & ~n11657 ;
  assign n11660 = ~n11658 & n11659 ;
  assign n11661 = ~n11598 & ~n11600 ;
  assign n11662 = ~n11405 & ~n11479 ;
  assign n11663 = ~n11478 & ~n11662 ;
  assign n11664 = ~n11480 & ~n11484 ;
  assign n11665 = ~n11663 & n11664 ;
  assign n11666 = ~n11485 & ~n11665 ;
  assign n11668 = n11661 & n11666 ;
  assign n11667 = ~n11661 & ~n11666 ;
  assign n11669 = n11404 & ~n11667 ;
  assign n11670 = ~n11668 & n11669 ;
  assign n11681 = ~n11660 & ~n11670 ;
  assign n11682 = ~n11680 & n11681 ;
  assign n11683 = \P1_state_reg[0]/NET0131  & ~n11682 ;
  assign n11684 = ~n7071 & ~n11683 ;
  assign n11694 = ~n11572 & ~n11581 ;
  assign n11696 = n11578 & n11694 ;
  assign n11695 = ~n11578 & ~n11694 ;
  assign n11697 = n11437 & ~n11695 ;
  assign n11698 = ~n11696 & n11697 ;
  assign n11686 = ~n1188 & ~n11399 ;
  assign n11685 = ~\P1_addr_reg[11]/NET0131  & n11399 ;
  assign n11687 = ~n537 & ~n11685 ;
  assign n11688 = ~n11686 & n11687 ;
  assign n11689 = ~n11597 & ~n11606 ;
  assign n11691 = n11603 & n11689 ;
  assign n11690 = ~n11603 & ~n11689 ;
  assign n11692 = n11404 & ~n11690 ;
  assign n11693 = ~n11691 & n11692 ;
  assign n11699 = ~n11688 & ~n11693 ;
  assign n11700 = ~n11698 & n11699 ;
  assign n11701 = \P1_state_reg[0]/NET0131  & ~n11700 ;
  assign n11702 = ~n7997 & ~n11701 ;
  assign n11716 = ~n11571 & ~n11580 ;
  assign n11717 = ~n11573 & n11676 ;
  assign n11718 = ~n11575 & ~n11581 ;
  assign n11719 = ~n11717 & n11718 ;
  assign n11720 = ~n11572 & ~n11719 ;
  assign n11722 = n11716 & n11720 ;
  assign n11721 = ~n11716 & ~n11720 ;
  assign n11723 = n11437 & ~n11721 ;
  assign n11724 = ~n11722 & n11723 ;
  assign n11704 = ~n1154 & ~n11399 ;
  assign n11703 = ~\P1_addr_reg[12]/NET0131  & n11399 ;
  assign n11705 = ~n537 & ~n11703 ;
  assign n11706 = ~n11704 & n11705 ;
  assign n11707 = ~n11596 & ~n11605 ;
  assign n11708 = ~n11598 & n11666 ;
  assign n11709 = ~n11600 & ~n11606 ;
  assign n11710 = ~n11708 & n11709 ;
  assign n11711 = ~n11597 & ~n11710 ;
  assign n11713 = n11707 & n11711 ;
  assign n11712 = ~n11707 & ~n11711 ;
  assign n11714 = n11404 & ~n11712 ;
  assign n11715 = ~n11713 & n11714 ;
  assign n11725 = ~n11706 & ~n11715 ;
  assign n11726 = ~n11724 & n11725 ;
  assign n11727 = \P1_state_reg[0]/NET0131  & ~n11726 ;
  assign n11728 = ~n6089 & ~n11727 ;
  assign n11777 = \P2_reg2_reg[10]/NET0131  & ~n2745 ;
  assign n11778 = ~\P2_reg2_reg[10]/NET0131  & n2745 ;
  assign n11779 = ~n11777 & ~n11778 ;
  assign n11780 = \P2_reg2_reg[9]/NET0131  & ~n2769 ;
  assign n11781 = ~\P2_reg2_reg[9]/NET0131  & n2769 ;
  assign n11782 = ~\P2_reg2_reg[8]/NET0131  & ~n2460 ;
  assign n11783 = ~n11781 & ~n11782 ;
  assign n11784 = \P2_reg2_reg[8]/NET0131  & n2460 ;
  assign n11785 = ~\P2_reg2_reg[7]/NET0131  & ~n2485 ;
  assign n11787 = ~\P2_reg2_reg[6]/NET0131  & ~n2519 ;
  assign n11788 = \P2_reg2_reg[5]/NET0131  & ~n2542 ;
  assign n11789 = ~\P2_reg2_reg[5]/NET0131  & n2542 ;
  assign n11790 = ~\P2_reg2_reg[4]/NET0131  & ~n2646 ;
  assign n11791 = \P2_reg2_reg[4]/NET0131  & n2646 ;
  assign n11792 = ~\P2_reg2_reg[3]/NET0131  & ~n2629 ;
  assign n11793 = \P2_reg2_reg[3]/NET0131  & n2629 ;
  assign n11794 = ~\P2_reg2_reg[2]/NET0131  & ~n2564 ;
  assign n11795 = \P2_reg2_reg[2]/NET0131  & n2564 ;
  assign n11796 = ~\P2_reg2_reg[1]/NET0131  & ~n2578 ;
  assign n11797 = \P2_reg2_reg[1]/NET0131  & n2578 ;
  assign n11798 = ~n11632 & ~n11797 ;
  assign n11799 = ~n11796 & ~n11798 ;
  assign n11800 = ~n11795 & ~n11799 ;
  assign n11801 = ~n11794 & ~n11800 ;
  assign n11802 = ~n11793 & ~n11801 ;
  assign n11803 = ~n11792 & ~n11802 ;
  assign n11804 = ~n11791 & ~n11803 ;
  assign n11805 = ~n11790 & ~n11804 ;
  assign n11806 = ~n11789 & n11805 ;
  assign n11807 = ~n11788 & ~n11806 ;
  assign n11808 = ~n11787 & ~n11807 ;
  assign n11786 = \P2_reg2_reg[6]/NET0131  & n2519 ;
  assign n11809 = \P2_reg2_reg[7]/NET0131  & n2485 ;
  assign n11810 = ~n11786 & ~n11809 ;
  assign n11811 = ~n11808 & n11810 ;
  assign n11812 = ~n11785 & ~n11811 ;
  assign n11813 = ~n11784 & ~n11812 ;
  assign n11814 = n11783 & ~n11813 ;
  assign n11815 = ~n11780 & ~n11814 ;
  assign n11817 = n11779 & ~n11815 ;
  assign n11816 = ~n11779 & n11815 ;
  assign n11818 = n11630 & ~n11816 ;
  assign n11819 = ~n11817 & n11818 ;
  assign n11729 = ~n2024 & ~n2051 ;
  assign n11731 = n2745 & ~n11729 ;
  assign n11730 = ~\P2_addr_reg[10]/NET0131  & n11729 ;
  assign n11732 = ~n2058 & ~n11730 ;
  assign n11733 = ~n11731 & n11732 ;
  assign n11734 = \P2_reg1_reg[10]/NET0131  & ~n2745 ;
  assign n11735 = ~\P2_reg1_reg[10]/NET0131  & n2745 ;
  assign n11736 = ~n11734 & ~n11735 ;
  assign n11737 = \P2_reg1_reg[9]/NET0131  & ~n2769 ;
  assign n11738 = ~\P2_reg1_reg[9]/NET0131  & n2769 ;
  assign n11739 = ~\P2_reg1_reg[8]/NET0131  & ~n2460 ;
  assign n11740 = ~n11738 & ~n11739 ;
  assign n11741 = \P2_reg1_reg[8]/NET0131  & n2460 ;
  assign n11742 = ~\P2_reg1_reg[7]/NET0131  & ~n2485 ;
  assign n11744 = ~\P2_reg1_reg[6]/NET0131  & ~n2519 ;
  assign n11745 = \P2_reg1_reg[5]/NET0131  & ~n2542 ;
  assign n11746 = ~\P2_reg1_reg[5]/NET0131  & n2542 ;
  assign n11747 = ~\P2_reg1_reg[4]/NET0131  & ~n2646 ;
  assign n11748 = ~\P2_reg1_reg[3]/NET0131  & ~n2629 ;
  assign n11749 = ~\P2_reg1_reg[2]/NET0131  & ~n2564 ;
  assign n11750 = \P2_reg1_reg[2]/NET0131  & n2564 ;
  assign n11751 = ~\P2_reg1_reg[1]/NET0131  & ~n2578 ;
  assign n11752 = \P2_reg1_reg[1]/NET0131  & n2578 ;
  assign n11753 = ~n11627 & ~n11752 ;
  assign n11754 = ~n11751 & ~n11753 ;
  assign n11755 = ~n11750 & ~n11754 ;
  assign n11756 = ~n11749 & ~n11755 ;
  assign n11757 = ~n11748 & n11756 ;
  assign n11758 = \P2_reg1_reg[4]/NET0131  & n2646 ;
  assign n11759 = \P2_reg1_reg[3]/NET0131  & n2629 ;
  assign n11760 = ~n11758 & ~n11759 ;
  assign n11761 = ~n11757 & n11760 ;
  assign n11762 = ~n11747 & ~n11761 ;
  assign n11763 = ~n11746 & n11762 ;
  assign n11764 = ~n11745 & ~n11763 ;
  assign n11765 = ~n11744 & ~n11764 ;
  assign n11743 = \P2_reg1_reg[6]/NET0131  & n2519 ;
  assign n11766 = \P2_reg1_reg[7]/NET0131  & n2485 ;
  assign n11767 = ~n11743 & ~n11766 ;
  assign n11768 = ~n11765 & n11767 ;
  assign n11769 = ~n11742 & ~n11768 ;
  assign n11770 = ~n11741 & ~n11769 ;
  assign n11771 = n11740 & ~n11770 ;
  assign n11772 = ~n11737 & ~n11771 ;
  assign n11774 = n11736 & ~n11772 ;
  assign n11773 = ~n11736 & n11772 ;
  assign n11775 = n11626 & ~n11773 ;
  assign n11776 = ~n11774 & n11775 ;
  assign n11820 = ~n11733 & ~n11776 ;
  assign n11821 = ~n11819 & n11820 ;
  assign n11822 = \P1_state_reg[0]/NET0131  & ~n11821 ;
  assign n11823 = ~n7154 & ~n11822 ;
  assign n11839 = \P1_reg2_reg[14]/NET0131  & n1099 ;
  assign n11840 = ~\P1_reg2_reg[14]/NET0131  & ~n1099 ;
  assign n11841 = ~n11839 & ~n11840 ;
  assign n11842 = ~n11571 & n11720 ;
  assign n11843 = ~n11568 & ~n11580 ;
  assign n11844 = ~n11842 & n11843 ;
  assign n11845 = ~n11569 & ~n11844 ;
  assign n11847 = n11841 & n11845 ;
  assign n11846 = ~n11841 & ~n11845 ;
  assign n11848 = n11437 & ~n11846 ;
  assign n11849 = ~n11847 & n11848 ;
  assign n11825 = ~n1099 & ~n11399 ;
  assign n11824 = ~\P1_addr_reg[14]/NET0131  & n11399 ;
  assign n11826 = ~n537 & ~n11824 ;
  assign n11827 = ~n11825 & n11826 ;
  assign n11828 = \P1_reg1_reg[14]/NET0131  & n1099 ;
  assign n11829 = ~\P1_reg1_reg[14]/NET0131  & ~n1099 ;
  assign n11830 = ~n11828 & ~n11829 ;
  assign n11831 = ~n11596 & n11711 ;
  assign n11832 = ~n11593 & ~n11605 ;
  assign n11833 = ~n11831 & n11832 ;
  assign n11834 = ~n11594 & ~n11833 ;
  assign n11836 = n11830 & n11834 ;
  assign n11835 = ~n11830 & ~n11834 ;
  assign n11837 = n11404 & ~n11835 ;
  assign n11838 = ~n11836 & n11837 ;
  assign n11850 = ~n11827 & ~n11838 ;
  assign n11851 = ~n11849 & n11850 ;
  assign n11852 = \P1_state_reg[0]/NET0131  & ~n11851 ;
  assign n11853 = ~n8038 & ~n11852 ;
  assign n11875 = ~\P2_reg2_reg[11]/NET0131  & ~n2694 ;
  assign n11876 = \P2_reg2_reg[11]/NET0131  & n2694 ;
  assign n11877 = ~n11875 & ~n11876 ;
  assign n11878 = ~n11786 & ~n11788 ;
  assign n11879 = ~n11806 & n11878 ;
  assign n11880 = ~n11787 & ~n11879 ;
  assign n11881 = ~n11785 & n11880 ;
  assign n11882 = ~n11784 & ~n11809 ;
  assign n11883 = ~n11881 & n11882 ;
  assign n11884 = n11783 & ~n11883 ;
  assign n11885 = ~n11777 & ~n11780 ;
  assign n11886 = ~n11884 & n11885 ;
  assign n11887 = ~n11778 & ~n11886 ;
  assign n11889 = n11877 & n11887 ;
  assign n11888 = ~n11877 & ~n11887 ;
  assign n11890 = n11630 & ~n11888 ;
  assign n11891 = ~n11889 & n11890 ;
  assign n11855 = ~n2694 & ~n11729 ;
  assign n11854 = ~\P2_addr_reg[11]/NET0131  & n11729 ;
  assign n11856 = ~n2058 & ~n11854 ;
  assign n11857 = ~n11855 & n11856 ;
  assign n11858 = ~\P2_reg1_reg[11]/NET0131  & ~n2694 ;
  assign n11859 = \P2_reg1_reg[11]/NET0131  & n2694 ;
  assign n11860 = ~n11858 & ~n11859 ;
  assign n11861 = ~n11743 & ~n11745 ;
  assign n11862 = ~n11763 & n11861 ;
  assign n11863 = ~n11744 & ~n11862 ;
  assign n11864 = ~n11742 & n11863 ;
  assign n11865 = ~n11741 & ~n11766 ;
  assign n11866 = ~n11864 & n11865 ;
  assign n11867 = n11740 & ~n11866 ;
  assign n11868 = ~n11734 & ~n11737 ;
  assign n11869 = ~n11867 & n11868 ;
  assign n11870 = ~n11735 & ~n11869 ;
  assign n11872 = n11860 & n11870 ;
  assign n11871 = ~n11860 & ~n11870 ;
  assign n11873 = n11626 & ~n11871 ;
  assign n11874 = ~n11872 & n11873 ;
  assign n11892 = ~n11857 & ~n11874 ;
  assign n11893 = ~n11891 & n11892 ;
  assign n11894 = \P1_state_reg[0]/NET0131  & ~n11893 ;
  assign n11895 = ~n8121 & ~n11894 ;
  assign n11911 = \P2_reg2_reg[12]/NET0131  & n2720 ;
  assign n11912 = ~\P2_reg2_reg[12]/NET0131  & ~n2720 ;
  assign n11913 = ~n11911 & ~n11912 ;
  assign n11914 = ~n11778 & ~n11815 ;
  assign n11915 = ~n11777 & ~n11876 ;
  assign n11916 = ~n11914 & n11915 ;
  assign n11917 = ~n11875 & ~n11916 ;
  assign n11919 = n11913 & n11917 ;
  assign n11918 = ~n11913 & ~n11917 ;
  assign n11920 = n11630 & ~n11918 ;
  assign n11921 = ~n11919 & n11920 ;
  assign n11897 = ~n2720 & ~n11729 ;
  assign n11896 = ~\P2_addr_reg[12]/NET0131  & n11729 ;
  assign n11898 = ~n2058 & ~n11896 ;
  assign n11899 = ~n11897 & n11898 ;
  assign n11900 = \P2_reg1_reg[12]/NET0131  & n2720 ;
  assign n11901 = ~\P2_reg1_reg[12]/NET0131  & ~n2720 ;
  assign n11902 = ~n11900 & ~n11901 ;
  assign n11903 = ~n11735 & ~n11772 ;
  assign n11904 = ~n11734 & ~n11859 ;
  assign n11905 = ~n11903 & n11904 ;
  assign n11906 = ~n11858 & ~n11905 ;
  assign n11908 = n11902 & n11906 ;
  assign n11907 = ~n11902 & ~n11906 ;
  assign n11909 = n11626 & ~n11907 ;
  assign n11910 = ~n11908 & n11909 ;
  assign n11922 = ~n11899 & ~n11910 ;
  assign n11923 = ~n11921 & n11922 ;
  assign n11924 = \P1_state_reg[0]/NET0131  & ~n11923 ;
  assign n11925 = ~n6174 & ~n11924 ;
  assign n11941 = \P2_reg2_reg[13]/NET0131  & ~n2883 ;
  assign n11942 = ~\P2_reg2_reg[13]/NET0131  & n2883 ;
  assign n11943 = ~n11941 & ~n11942 ;
  assign n11944 = ~n11875 & n11887 ;
  assign n11945 = ~n11876 & ~n11911 ;
  assign n11946 = ~n11944 & n11945 ;
  assign n11947 = ~n11912 & ~n11946 ;
  assign n11949 = n11943 & n11947 ;
  assign n11948 = ~n11943 & ~n11947 ;
  assign n11950 = n11630 & ~n11948 ;
  assign n11951 = ~n11949 & n11950 ;
  assign n11927 = n2883 & ~n11729 ;
  assign n11926 = ~\P2_addr_reg[13]/NET0131  & n11729 ;
  assign n11928 = ~n2058 & ~n11926 ;
  assign n11929 = ~n11927 & n11928 ;
  assign n11930 = \P2_reg1_reg[13]/NET0131  & ~n2883 ;
  assign n11931 = ~\P2_reg1_reg[13]/NET0131  & n2883 ;
  assign n11932 = ~n11930 & ~n11931 ;
  assign n11933 = ~n11858 & n11870 ;
  assign n11934 = ~n11859 & ~n11900 ;
  assign n11935 = ~n11933 & n11934 ;
  assign n11936 = ~n11901 & ~n11935 ;
  assign n11938 = n11932 & n11936 ;
  assign n11937 = ~n11932 & ~n11936 ;
  assign n11939 = n11626 & ~n11937 ;
  assign n11940 = ~n11938 & n11939 ;
  assign n11952 = ~n11929 & ~n11940 ;
  assign n11953 = ~n11951 & n11952 ;
  assign n11954 = \P1_state_reg[0]/NET0131  & ~n11953 ;
  assign n11955 = ~n7197 & ~n11954 ;
  assign n11972 = ~\P1_reg1_reg[15]/NET0131  & ~n1073 ;
  assign n11973 = \P1_reg1_reg[15]/NET0131  & n1073 ;
  assign n11974 = ~n11972 & ~n11973 ;
  assign n11975 = ~n11594 & n11609 ;
  assign n11976 = ~n11593 & ~n11828 ;
  assign n11977 = ~n11975 & n11976 ;
  assign n11978 = ~n11829 & ~n11977 ;
  assign n11980 = n11974 & n11978 ;
  assign n11979 = ~n11974 & ~n11978 ;
  assign n11981 = n11404 & ~n11979 ;
  assign n11982 = ~n11980 & n11981 ;
  assign n11957 = ~n1073 & ~n11399 ;
  assign n11956 = ~\P1_addr_reg[15]/NET0131  & n11399 ;
  assign n11958 = ~n537 & ~n11956 ;
  assign n11959 = ~n11957 & n11958 ;
  assign n11960 = ~\P1_reg2_reg[15]/NET0131  & ~n1073 ;
  assign n11961 = \P1_reg2_reg[15]/NET0131  & n1073 ;
  assign n11962 = ~n11960 & ~n11961 ;
  assign n11963 = ~n11569 & ~n11840 ;
  assign n11964 = n11584 & n11963 ;
  assign n11965 = n11568 & ~n11840 ;
  assign n11966 = ~n11839 & ~n11965 ;
  assign n11967 = ~n11964 & n11966 ;
  assign n11969 = n11962 & ~n11967 ;
  assign n11968 = ~n11962 & n11967 ;
  assign n11970 = n11437 & ~n11968 ;
  assign n11971 = ~n11969 & n11970 ;
  assign n11983 = ~n11959 & ~n11971 ;
  assign n11984 = ~n11982 & n11983 ;
  assign n11985 = \P1_state_reg[0]/NET0131  & ~n11984 ;
  assign n11986 = ~n8082 & ~n11985 ;
  assign n12002 = \P2_reg2_reg[14]/NET0131  & n2849 ;
  assign n12003 = ~\P2_reg2_reg[14]/NET0131  & ~n2849 ;
  assign n12004 = ~n12002 & ~n12003 ;
  assign n12005 = ~n11912 & n11917 ;
  assign n12006 = ~n11911 & ~n11941 ;
  assign n12007 = ~n12005 & n12006 ;
  assign n12008 = ~n11942 & ~n12007 ;
  assign n12010 = n12004 & n12008 ;
  assign n12009 = ~n12004 & ~n12008 ;
  assign n12011 = n11630 & ~n12009 ;
  assign n12012 = ~n12010 & n12011 ;
  assign n11988 = ~n2849 & ~n11729 ;
  assign n11987 = ~\P2_addr_reg[14]/NET0131  & n11729 ;
  assign n11989 = ~n2058 & ~n11987 ;
  assign n11990 = ~n11988 & n11989 ;
  assign n11991 = \P2_reg1_reg[14]/NET0131  & n2849 ;
  assign n11992 = ~\P2_reg1_reg[14]/NET0131  & ~n2849 ;
  assign n11993 = ~n11991 & ~n11992 ;
  assign n11994 = ~n11901 & n11906 ;
  assign n11995 = ~n11900 & ~n11930 ;
  assign n11996 = ~n11994 & n11995 ;
  assign n11997 = ~n11931 & ~n11996 ;
  assign n11999 = n11993 & n11997 ;
  assign n11998 = ~n11993 & ~n11997 ;
  assign n12000 = n11626 & ~n11998 ;
  assign n12001 = ~n11999 & n12000 ;
  assign n12013 = ~n11990 & ~n12001 ;
  assign n12014 = ~n12012 & n12013 ;
  assign n12015 = \P1_state_reg[0]/NET0131  & ~n12014 ;
  assign n12016 = ~n8162 & ~n12015 ;
  assign n12032 = ~\P2_reg2_reg[15]/NET0131  & ~n2832 ;
  assign n12033 = \P2_reg2_reg[15]/NET0131  & n2832 ;
  assign n12034 = ~n12032 & ~n12033 ;
  assign n12035 = ~n11942 & n11947 ;
  assign n12036 = ~n11941 & ~n12002 ;
  assign n12037 = ~n12035 & n12036 ;
  assign n12038 = ~n12003 & ~n12037 ;
  assign n12040 = n12034 & n12038 ;
  assign n12039 = ~n12034 & ~n12038 ;
  assign n12041 = n11630 & ~n12039 ;
  assign n12042 = ~n12040 & n12041 ;
  assign n12018 = ~n2832 & ~n11729 ;
  assign n12017 = ~\P2_addr_reg[15]/NET0131  & n11729 ;
  assign n12019 = ~n2058 & ~n12017 ;
  assign n12020 = ~n12018 & n12019 ;
  assign n12021 = ~\P2_reg1_reg[15]/NET0131  & ~n2832 ;
  assign n12022 = \P2_reg1_reg[15]/NET0131  & n2832 ;
  assign n12023 = ~n12021 & ~n12022 ;
  assign n12024 = ~n11931 & n11936 ;
  assign n12025 = ~n11930 & ~n11991 ;
  assign n12026 = ~n12024 & n12025 ;
  assign n12027 = ~n11992 & ~n12026 ;
  assign n12029 = n12023 & n12027 ;
  assign n12028 = ~n12023 & ~n12027 ;
  assign n12030 = n11626 & ~n12028 ;
  assign n12031 = ~n12029 & n12030 ;
  assign n12043 = ~n12020 & ~n12031 ;
  assign n12044 = ~n12042 & n12043 ;
  assign n12045 = \P1_state_reg[0]/NET0131  & ~n12044 ;
  assign n12046 = ~n8203 & ~n12045 ;
  assign n12062 = \P2_reg2_reg[16]/NET0131  & n2808 ;
  assign n12063 = ~\P2_reg2_reg[16]/NET0131  & ~n2808 ;
  assign n12064 = ~n12062 & ~n12063 ;
  assign n12065 = ~n12003 & n12008 ;
  assign n12066 = ~n12002 & ~n12033 ;
  assign n12067 = ~n12065 & n12066 ;
  assign n12068 = ~n12032 & ~n12067 ;
  assign n12070 = n12064 & n12068 ;
  assign n12069 = ~n12064 & ~n12068 ;
  assign n12071 = n11630 & ~n12069 ;
  assign n12072 = ~n12070 & n12071 ;
  assign n12048 = ~n2808 & ~n11729 ;
  assign n12047 = ~\P2_addr_reg[16]/NET0131  & n11729 ;
  assign n12049 = ~n2058 & ~n12047 ;
  assign n12050 = ~n12048 & n12049 ;
  assign n12051 = \P2_reg1_reg[16]/NET0131  & n2808 ;
  assign n12052 = ~\P2_reg1_reg[16]/NET0131  & ~n2808 ;
  assign n12053 = ~n12051 & ~n12052 ;
  assign n12054 = ~n11992 & n11997 ;
  assign n12055 = ~n11991 & ~n12022 ;
  assign n12056 = ~n12054 & n12055 ;
  assign n12057 = ~n12021 & ~n12056 ;
  assign n12059 = n12053 & n12057 ;
  assign n12058 = ~n12053 & ~n12057 ;
  assign n12060 = n11626 & ~n12058 ;
  assign n12061 = ~n12059 & n12060 ;
  assign n12073 = ~n12050 & ~n12061 ;
  assign n12074 = ~n12072 & n12073 ;
  assign n12075 = \P1_state_reg[0]/NET0131  & ~n12074 ;
  assign n12076 = ~n6218 & ~n12075 ;
  assign n12092 = ~\P2_reg2_reg[17]/NET0131  & ~n2385 ;
  assign n12093 = \P2_reg2_reg[17]/NET0131  & n2385 ;
  assign n12094 = ~n12092 & ~n12093 ;
  assign n12095 = ~n12032 & n12038 ;
  assign n12096 = ~n12033 & ~n12062 ;
  assign n12097 = ~n12095 & n12096 ;
  assign n12098 = ~n12063 & ~n12097 ;
  assign n12100 = n12094 & n12098 ;
  assign n12099 = ~n12094 & ~n12098 ;
  assign n12101 = n11630 & ~n12099 ;
  assign n12102 = ~n12100 & n12101 ;
  assign n12078 = ~n2385 & ~n11729 ;
  assign n12077 = ~\P2_addr_reg[17]/NET0131  & n11729 ;
  assign n12079 = ~n2058 & ~n12077 ;
  assign n12080 = ~n12078 & n12079 ;
  assign n12081 = ~\P2_reg1_reg[17]/NET0131  & ~n2385 ;
  assign n12082 = \P2_reg1_reg[17]/NET0131  & n2385 ;
  assign n12083 = ~n12081 & ~n12082 ;
  assign n12084 = ~n12021 & n12027 ;
  assign n12085 = ~n12022 & ~n12051 ;
  assign n12086 = ~n12084 & n12085 ;
  assign n12087 = ~n12052 & ~n12086 ;
  assign n12089 = n12083 & n12087 ;
  assign n12088 = ~n12083 & ~n12087 ;
  assign n12090 = n11626 & ~n12088 ;
  assign n12091 = ~n12089 & n12090 ;
  assign n12103 = ~n12080 & ~n12091 ;
  assign n12104 = ~n12102 & n12103 ;
  assign n12105 = \P1_state_reg[0]/NET0131  & ~n12104 ;
  assign n12106 = ~n5551 & ~n12105 ;
  assign n12122 = \P1_reg2_reg[16]/NET0131  & n1456 ;
  assign n12123 = ~\P1_reg2_reg[16]/NET0131  & ~n1456 ;
  assign n12124 = ~n12122 & ~n12123 ;
  assign n12125 = ~n11840 & n11845 ;
  assign n12126 = ~n11839 & ~n11961 ;
  assign n12127 = ~n12125 & n12126 ;
  assign n12128 = ~n11960 & ~n12127 ;
  assign n12130 = n12124 & n12128 ;
  assign n12129 = ~n12124 & ~n12128 ;
  assign n12131 = n11437 & ~n12129 ;
  assign n12132 = ~n12130 & n12131 ;
  assign n12108 = ~n1456 & ~n11399 ;
  assign n12107 = ~\P1_addr_reg[16]/NET0131  & n11399 ;
  assign n12109 = ~n537 & ~n12107 ;
  assign n12110 = ~n12108 & n12109 ;
  assign n12111 = \P1_reg1_reg[16]/NET0131  & n1456 ;
  assign n12112 = ~\P1_reg1_reg[16]/NET0131  & ~n1456 ;
  assign n12113 = ~n12111 & ~n12112 ;
  assign n12114 = ~n11829 & n11834 ;
  assign n12115 = ~n11828 & ~n11973 ;
  assign n12116 = ~n12114 & n12115 ;
  assign n12117 = ~n11972 & ~n12116 ;
  assign n12119 = n12113 & n12117 ;
  assign n12118 = ~n12113 & ~n12117 ;
  assign n12120 = n11404 & ~n12118 ;
  assign n12121 = ~n12119 & n12120 ;
  assign n12133 = ~n12110 & ~n12121 ;
  assign n12134 = ~n12132 & n12133 ;
  assign n12135 = \P1_state_reg[0]/NET0131  & ~n12134 ;
  assign n12136 = ~n6132 & ~n12135 ;
  assign n12137 = ~\P1_state_reg[0]/NET0131  & \P2_reg3_reg[1]/NET0131  ;
  assign n12140 = n2024 & ~n2578 ;
  assign n12139 = ~\P2_addr_reg[1]/NET0131  & ~n2024 ;
  assign n12141 = n2059 & ~n12139 ;
  assign n12142 = ~n12140 & n12141 ;
  assign n12148 = ~n11751 & ~n11752 ;
  assign n12149 = ~n11627 & ~n12148 ;
  assign n12150 = n11627 & n12148 ;
  assign n12151 = ~n12149 & ~n12150 ;
  assign n12152 = n11626 & n12151 ;
  assign n12138 = n2578 & n11619 ;
  assign n12143 = ~n11796 & ~n11797 ;
  assign n12144 = ~n11632 & ~n12143 ;
  assign n12145 = n11632 & n12143 ;
  assign n12146 = ~n12144 & ~n12145 ;
  assign n12147 = n11630 & n12146 ;
  assign n12153 = ~n12138 & ~n12147 ;
  assign n12154 = ~n12152 & n12153 ;
  assign n12155 = ~n12142 & n12154 ;
  assign n12156 = \P1_state_reg[0]/NET0131  & ~n12155 ;
  assign n12157 = ~n12137 & ~n12156 ;
  assign n12173 = ~\P1_reg1_reg[17]/NET0131  & n1433 ;
  assign n12174 = \P1_reg1_reg[17]/NET0131  & ~n1433 ;
  assign n12175 = ~n12173 & ~n12174 ;
  assign n12176 = ~n11972 & n11978 ;
  assign n12177 = ~n11973 & ~n12111 ;
  assign n12178 = ~n12176 & n12177 ;
  assign n12179 = ~n12112 & ~n12178 ;
  assign n12181 = n12175 & n12179 ;
  assign n12180 = ~n12175 & ~n12179 ;
  assign n12182 = n11404 & ~n12180 ;
  assign n12183 = ~n12181 & n12182 ;
  assign n12159 = n1433 & ~n11399 ;
  assign n12158 = ~\P1_addr_reg[17]/NET0131  & n11399 ;
  assign n12160 = ~n537 & ~n12158 ;
  assign n12161 = ~n12159 & n12160 ;
  assign n12162 = ~\P1_reg2_reg[17]/NET0131  & n1433 ;
  assign n12163 = \P1_reg2_reg[17]/NET0131  & ~n1433 ;
  assign n12164 = ~n12162 & ~n12163 ;
  assign n12165 = ~n11960 & ~n11967 ;
  assign n12166 = ~n11961 & ~n12122 ;
  assign n12167 = ~n12165 & n12166 ;
  assign n12168 = ~n12123 & ~n12167 ;
  assign n12170 = n12164 & n12168 ;
  assign n12169 = ~n12164 & ~n12168 ;
  assign n12171 = n11437 & ~n12169 ;
  assign n12172 = ~n12170 & n12171 ;
  assign n12184 = ~n12161 & ~n12172 ;
  assign n12185 = ~n12183 & n12184 ;
  assign n12186 = \P1_state_reg[0]/NET0131  & ~n12185 ;
  assign n12187 = ~n5426 & ~n12186 ;
  assign n12188 = ~\P1_state_reg[0]/NET0131  & \P2_reg3_reg[2]/NET0131  ;
  assign n12191 = n2024 & ~n2564 ;
  assign n12190 = ~\P2_addr_reg[2]/NET0131  & ~n2024 ;
  assign n12192 = n2059 & ~n12190 ;
  assign n12193 = ~n12191 & n12192 ;
  assign n12199 = ~n11749 & ~n11750 ;
  assign n12200 = ~n11754 & ~n12199 ;
  assign n12201 = n11754 & n12199 ;
  assign n12202 = ~n12200 & ~n12201 ;
  assign n12203 = n11626 & n12202 ;
  assign n12189 = n2564 & n11619 ;
  assign n12194 = ~n11794 & ~n11795 ;
  assign n12195 = ~n11799 & ~n12194 ;
  assign n12196 = n11799 & n12194 ;
  assign n12197 = ~n12195 & ~n12196 ;
  assign n12198 = n11630 & n12197 ;
  assign n12204 = ~n12189 & ~n12198 ;
  assign n12205 = ~n12203 & n12204 ;
  assign n12206 = ~n12193 & n12205 ;
  assign n12207 = \P1_state_reg[0]/NET0131  & ~n12206 ;
  assign n12208 = ~n12188 & ~n12207 ;
  assign n12211 = n2024 & ~n2629 ;
  assign n12210 = ~\P2_addr_reg[3]/NET0131  & ~n2024 ;
  assign n12212 = n2059 & ~n12210 ;
  assign n12213 = ~n12211 & n12212 ;
  assign n12219 = ~n11792 & ~n11793 ;
  assign n12220 = ~n11801 & ~n12219 ;
  assign n12221 = n11801 & n12219 ;
  assign n12222 = ~n12220 & ~n12221 ;
  assign n12223 = n11630 & n12222 ;
  assign n12209 = n2629 & n11619 ;
  assign n12214 = ~n11748 & ~n11759 ;
  assign n12215 = ~n11756 & ~n12214 ;
  assign n12216 = n11756 & n12214 ;
  assign n12217 = ~n12215 & ~n12216 ;
  assign n12218 = n11626 & n12217 ;
  assign n12224 = ~n12209 & ~n12218 ;
  assign n12225 = ~n12223 & n12224 ;
  assign n12226 = ~n12213 & n12225 ;
  assign n12227 = \P1_state_reg[0]/NET0131  & ~n12226 ;
  assign n12228 = ~n9575 & ~n12227 ;
  assign n12231 = n2024 & ~n2646 ;
  assign n12230 = ~\P2_addr_reg[4]/NET0131  & ~n2024 ;
  assign n12232 = n2059 & ~n12230 ;
  assign n12233 = ~n12231 & n12232 ;
  assign n12239 = ~n11757 & ~n11759 ;
  assign n12240 = ~n11747 & ~n11758 ;
  assign n12241 = n12239 & ~n12240 ;
  assign n12242 = ~n12239 & n12240 ;
  assign n12243 = ~n12241 & ~n12242 ;
  assign n12244 = n11626 & n12243 ;
  assign n12229 = n2646 & n11619 ;
  assign n12234 = ~n11790 & ~n11791 ;
  assign n12235 = ~n11803 & ~n12234 ;
  assign n12236 = n11803 & n12234 ;
  assign n12237 = ~n12235 & ~n12236 ;
  assign n12238 = n11630 & n12237 ;
  assign n12245 = ~n12229 & ~n12238 ;
  assign n12246 = ~n12244 & n12245 ;
  assign n12247 = ~n12233 & n12246 ;
  assign n12248 = \P1_state_reg[0]/NET0131  & ~n12247 ;
  assign n12249 = ~n8935 & ~n12248 ;
  assign n12252 = n2024 & n2542 ;
  assign n12251 = ~\P2_addr_reg[5]/NET0131  & ~n2024 ;
  assign n12253 = n2059 & ~n12251 ;
  assign n12254 = ~n12252 & n12253 ;
  assign n12260 = ~n11788 & ~n11789 ;
  assign n12262 = n11805 & n12260 ;
  assign n12261 = ~n11805 & ~n12260 ;
  assign n12263 = n11630 & ~n12261 ;
  assign n12264 = ~n12262 & n12263 ;
  assign n12250 = ~n2542 & n11619 ;
  assign n12257 = ~n11745 & n11763 ;
  assign n12255 = ~n11745 & ~n11746 ;
  assign n12256 = ~n11762 & ~n12255 ;
  assign n12258 = n11626 & ~n12256 ;
  assign n12259 = ~n12257 & n12258 ;
  assign n12265 = ~n12250 & ~n12259 ;
  assign n12266 = ~n12264 & n12265 ;
  assign n12267 = ~n12254 & n12266 ;
  assign n12268 = \P1_state_reg[0]/NET0131  & ~n12267 ;
  assign n12269 = ~n8977 & ~n12268 ;
  assign n12279 = ~n11786 & ~n11787 ;
  assign n12281 = ~n11807 & n12279 ;
  assign n12280 = n11807 & ~n12279 ;
  assign n12282 = n11630 & ~n12280 ;
  assign n12283 = ~n12281 & n12282 ;
  assign n12271 = ~n2519 & ~n11729 ;
  assign n12270 = ~\P2_addr_reg[6]/NET0131  & n11729 ;
  assign n12272 = ~n2058 & ~n12270 ;
  assign n12273 = ~n12271 & n12272 ;
  assign n12274 = ~n11743 & ~n11744 ;
  assign n12276 = ~n11764 & n12274 ;
  assign n12275 = n11764 & ~n12274 ;
  assign n12277 = n11626 & ~n12275 ;
  assign n12278 = ~n12276 & n12277 ;
  assign n12284 = ~n12273 & ~n12278 ;
  assign n12285 = ~n12283 & n12284 ;
  assign n12286 = \P1_state_reg[0]/NET0131  & ~n12285 ;
  assign n12287 = ~n9615 & ~n12286 ;
  assign n12299 = ~n11809 & n11881 ;
  assign n12297 = ~n11785 & ~n11809 ;
  assign n12298 = ~n11880 & ~n12297 ;
  assign n12300 = n11630 & ~n12298 ;
  assign n12301 = ~n12299 & n12300 ;
  assign n12290 = ~n11766 & n11864 ;
  assign n12288 = ~n11742 & ~n11766 ;
  assign n12289 = ~n11863 & ~n12288 ;
  assign n12291 = n11626 & ~n12289 ;
  assign n12292 = ~n12290 & n12291 ;
  assign n12294 = ~n2485 & ~n11729 ;
  assign n12293 = ~\P2_addr_reg[7]/NET0131  & n11729 ;
  assign n12295 = ~n2058 & ~n12293 ;
  assign n12296 = ~n12294 & n12295 ;
  assign n12302 = ~n12292 & ~n12296 ;
  assign n12303 = ~n12301 & n12302 ;
  assign n12304 = \P1_state_reg[0]/NET0131  & ~n12303 ;
  assign n12305 = ~n9656 & ~n12304 ;
  assign n12315 = ~n11782 & ~n11784 ;
  assign n12317 = n11812 & n12315 ;
  assign n12316 = ~n11812 & ~n12315 ;
  assign n12318 = n11630 & ~n12316 ;
  assign n12319 = ~n12317 & n12318 ;
  assign n12306 = ~n11739 & ~n11741 ;
  assign n12308 = n11769 & n12306 ;
  assign n12307 = ~n11769 & ~n12306 ;
  assign n12309 = n11626 & ~n12307 ;
  assign n12310 = ~n12308 & n12309 ;
  assign n12312 = ~n2460 & ~n11729 ;
  assign n12311 = ~\P2_addr_reg[8]/NET0131  & n11729 ;
  assign n12313 = ~n2058 & ~n12311 ;
  assign n12314 = ~n12312 & n12313 ;
  assign n12320 = ~n12310 & ~n12314 ;
  assign n12321 = ~n12319 & n12320 ;
  assign n12322 = \P1_state_reg[0]/NET0131  & ~n12321 ;
  assign n12323 = ~n8243 & ~n12322 ;
  assign n12337 = ~n11780 & n11884 ;
  assign n12334 = ~n11780 & ~n11781 ;
  assign n12335 = ~n11782 & ~n11883 ;
  assign n12336 = ~n12334 & ~n12335 ;
  assign n12338 = n11630 & ~n12336 ;
  assign n12339 = ~n12337 & n12338 ;
  assign n12327 = ~n11737 & n11867 ;
  assign n12324 = ~n11737 & ~n11738 ;
  assign n12325 = ~n11739 & ~n11866 ;
  assign n12326 = ~n12324 & ~n12325 ;
  assign n12328 = n11626 & ~n12326 ;
  assign n12329 = ~n12327 & n12328 ;
  assign n12331 = n2769 & ~n11729 ;
  assign n12330 = ~\P2_addr_reg[9]/NET0131  & n11729 ;
  assign n12332 = ~n2058 & ~n12330 ;
  assign n12333 = ~n12331 & n12332 ;
  assign n12340 = ~n12329 & ~n12333 ;
  assign n12341 = ~n12339 & n12340 ;
  assign n12342 = \P1_state_reg[0]/NET0131  & ~n12341 ;
  assign n12343 = ~n7238 & ~n12342 ;
  assign n12353 = ~n11478 & ~n11480 ;
  assign n12355 = ~n11662 & n12353 ;
  assign n12354 = n11662 & ~n12353 ;
  assign n12356 = n11404 & ~n12354 ;
  assign n12357 = ~n12355 & n12356 ;
  assign n12345 = ~n1271 & ~n11399 ;
  assign n12344 = ~\P1_addr_reg[8]/NET0131  & n11399 ;
  assign n12346 = ~n537 & ~n12344 ;
  assign n12347 = ~n12345 & n12346 ;
  assign n12348 = ~n11494 & ~n11496 ;
  assign n12350 = ~n11672 & n12348 ;
  assign n12349 = n11672 & ~n12348 ;
  assign n12351 = n11437 & ~n12349 ;
  assign n12352 = ~n12350 & n12351 ;
  assign n12358 = ~n12347 & ~n12352 ;
  assign n12359 = ~n12357 & n12358 ;
  assign n12360 = \P1_state_reg[0]/NET0131  & ~n12359 ;
  assign n12361 = ~n8283 & ~n12360 ;
  assign n12362 = \P1_reg3_reg[1]/NET0131  & ~\P1_state_reg[0]/NET0131  ;
  assign n12365 = ~n1645 & n3448 ;
  assign n12364 = ~\P1_addr_reg[1]/NET0131  & ~n3448 ;
  assign n12366 = n538 & ~n12364 ;
  assign n12367 = ~n12365 & n12366 ;
  assign n12373 = ~n11449 & ~n11450 ;
  assign n12374 = ~n11451 & ~n12373 ;
  assign n12375 = n11451 & n12373 ;
  assign n12376 = ~n12374 & ~n12375 ;
  assign n12377 = n11437 & n12376 ;
  assign n12363 = n1645 & n11527 ;
  assign n12368 = ~n11416 & ~n11417 ;
  assign n12369 = ~n11418 & ~n12368 ;
  assign n12370 = n11418 & n12368 ;
  assign n12371 = ~n12369 & ~n12370 ;
  assign n12372 = n11404 & n12371 ;
  assign n12378 = ~n12363 & ~n12372 ;
  assign n12379 = ~n12377 & n12378 ;
  assign n12380 = ~n12367 & n12379 ;
  assign n12381 = \P1_state_reg[0]/NET0131  & ~n12380 ;
  assign n12382 = ~n12362 & ~n12381 ;
  assign n12385 = n1584 & n3448 ;
  assign n12384 = ~\P1_addr_reg[4]/NET0131  & ~n3448 ;
  assign n12386 = n538 & ~n12384 ;
  assign n12387 = ~n12385 & n12386 ;
  assign n12393 = ~n11411 & ~n11427 ;
  assign n12394 = ~n11424 & ~n12393 ;
  assign n12395 = n11424 & n12393 ;
  assign n12396 = ~n12394 & ~n12395 ;
  assign n12397 = n11404 & n12396 ;
  assign n12383 = ~n1584 & n11527 ;
  assign n12388 = ~n11444 & ~n11460 ;
  assign n12389 = ~n11457 & ~n12388 ;
  assign n12390 = n11457 & n12388 ;
  assign n12391 = ~n12389 & ~n12390 ;
  assign n12392 = n11437 & n12391 ;
  assign n12398 = ~n12383 & ~n12392 ;
  assign n12399 = ~n12397 & n12398 ;
  assign n12400 = ~n12387 & n12399 ;
  assign n12401 = \P1_state_reg[0]/NET0131  & ~n12400 ;
  assign n12402 = ~n9016 & ~n12401 ;
  assign n12416 = n1560 & ~n11399 ;
  assign n12415 = ~\P1_addr_reg[5]/NET0131  & n11399 ;
  assign n12417 = ~n537 & ~n12415 ;
  assign n12418 = ~n12416 & n12417 ;
  assign n12406 = ~n11410 & n11429 ;
  assign n12403 = ~n11425 & ~n11427 ;
  assign n12404 = ~n11410 & ~n11426 ;
  assign n12405 = ~n12403 & ~n12404 ;
  assign n12407 = n11404 & ~n12405 ;
  assign n12408 = ~n12406 & n12407 ;
  assign n12412 = ~n11443 & n11462 ;
  assign n12409 = ~n11458 & ~n11460 ;
  assign n12410 = ~n11443 & ~n11459 ;
  assign n12411 = ~n12409 & ~n12410 ;
  assign n12413 = n11437 & ~n12411 ;
  assign n12414 = ~n12412 & n12413 ;
  assign n12419 = ~n12408 & ~n12414 ;
  assign n12420 = ~n12418 & n12419 ;
  assign n12421 = \P1_state_reg[0]/NET0131  & ~n12420 ;
  assign n12422 = ~n9058 & ~n12421 ;
  assign n12423 = ~\P1_state_reg[0]/NET0131  & \P2_reg3_reg[18]/NET0131  ;
  assign n12439 = \P2_reg2_reg[18]/NET0131  & n2404 ;
  assign n12440 = ~\P2_reg2_reg[18]/NET0131  & ~n2404 ;
  assign n12441 = ~n12439 & ~n12440 ;
  assign n12442 = ~n12063 & n12068 ;
  assign n12443 = ~n12062 & ~n12093 ;
  assign n12444 = ~n12442 & n12443 ;
  assign n12445 = ~n12092 & ~n12444 ;
  assign n12447 = n12441 & n12445 ;
  assign n12446 = ~n12441 & ~n12445 ;
  assign n12448 = n11630 & ~n12446 ;
  assign n12449 = ~n12447 & n12448 ;
  assign n12424 = \P2_reg1_reg[18]/NET0131  & n2404 ;
  assign n12425 = ~\P2_reg1_reg[18]/NET0131  & ~n2404 ;
  assign n12426 = ~n12424 & ~n12425 ;
  assign n12427 = ~n12052 & n12057 ;
  assign n12428 = ~n12051 & ~n12082 ;
  assign n12429 = ~n12427 & n12428 ;
  assign n12430 = ~n12081 & ~n12429 ;
  assign n12432 = n12426 & n12430 ;
  assign n12431 = ~n12426 & ~n12430 ;
  assign n12433 = n11626 & ~n12431 ;
  assign n12434 = ~n12432 & n12433 ;
  assign n12436 = ~n2404 & ~n11729 ;
  assign n12435 = ~\P2_addr_reg[18]/NET0131  & n11729 ;
  assign n12437 = ~n2058 & ~n12435 ;
  assign n12438 = ~n12436 & n12437 ;
  assign n12450 = ~n12434 & ~n12438 ;
  assign n12451 = ~n12449 & n12450 ;
  assign n12452 = \P1_state_reg[0]/NET0131  & ~n12451 ;
  assign n12453 = ~n12423 & ~n12452 ;
  assign n12469 = ~n12092 & n12098 ;
  assign n12470 = ~n12093 & ~n12439 ;
  assign n12471 = ~n12469 & n12470 ;
  assign n12472 = ~n12440 & ~n12471 ;
  assign n12473 = \P2_reg2_reg[19]/NET0131  & n12472 ;
  assign n12474 = ~\P2_reg2_reg[19]/NET0131  & ~n12472 ;
  assign n12475 = ~n12473 & ~n12474 ;
  assign n12477 = ~n2258 & ~n12475 ;
  assign n12476 = n2258 & n12475 ;
  assign n12478 = n11630 & ~n12476 ;
  assign n12479 = ~n12477 & n12478 ;
  assign n12454 = ~n12081 & n12087 ;
  assign n12455 = ~n12082 & ~n12424 ;
  assign n12456 = ~n12454 & n12455 ;
  assign n12457 = ~n12425 & ~n12456 ;
  assign n12458 = \P2_reg1_reg[19]/NET0131  & ~n12457 ;
  assign n12459 = ~\P2_reg1_reg[19]/NET0131  & n12457 ;
  assign n12460 = ~n12458 & ~n12459 ;
  assign n12462 = ~n2258 & n12460 ;
  assign n12461 = n2258 & ~n12460 ;
  assign n12463 = n11626 & ~n12461 ;
  assign n12464 = ~n12462 & n12463 ;
  assign n12466 = ~n2258 & ~n11729 ;
  assign n12465 = ~\P2_addr_reg[19]/NET0131  & n11729 ;
  assign n12467 = ~n2058 & ~n12465 ;
  assign n12468 = ~n12466 & n12467 ;
  assign n12480 = ~n12464 & ~n12468 ;
  assign n12481 = ~n12479 & n12480 ;
  assign n12482 = \P1_state_reg[0]/NET0131  & ~n12481 ;
  assign n12483 = ~n5602 & ~n12482 ;
  assign n12499 = \P1_reg2_reg[18]/NET0131  & n1384 ;
  assign n12500 = ~\P1_reg2_reg[18]/NET0131  & ~n1384 ;
  assign n12501 = ~n12499 & ~n12500 ;
  assign n12502 = ~n12123 & n12128 ;
  assign n12503 = ~n12122 & ~n12163 ;
  assign n12504 = ~n12502 & n12503 ;
  assign n12505 = ~n12162 & ~n12504 ;
  assign n12507 = n12501 & n12505 ;
  assign n12506 = ~n12501 & ~n12505 ;
  assign n12508 = n11437 & ~n12506 ;
  assign n12509 = ~n12507 & n12508 ;
  assign n12484 = \P1_reg1_reg[18]/NET0131  & n1384 ;
  assign n12485 = ~\P1_reg1_reg[18]/NET0131  & ~n1384 ;
  assign n12486 = ~n12484 & ~n12485 ;
  assign n12487 = ~n12112 & n12117 ;
  assign n12488 = ~n12111 & ~n12174 ;
  assign n12489 = ~n12487 & n12488 ;
  assign n12490 = ~n12173 & ~n12489 ;
  assign n12492 = n12486 & n12490 ;
  assign n12491 = ~n12486 & ~n12490 ;
  assign n12493 = n11404 & ~n12491 ;
  assign n12494 = ~n12492 & n12493 ;
  assign n12496 = ~n1384 & ~n11399 ;
  assign n12495 = ~\P1_addr_reg[18]/NET0131  & n11399 ;
  assign n12497 = ~n537 & ~n12495 ;
  assign n12498 = ~n12496 & n12497 ;
  assign n12510 = ~n12494 & ~n12498 ;
  assign n12511 = ~n12509 & n12510 ;
  assign n12512 = \P1_state_reg[0]/NET0131  & ~n12511 ;
  assign n12513 = ~n5477 & ~n12512 ;
  assign n12529 = ~n12162 & n12168 ;
  assign n12530 = ~n12163 & ~n12499 ;
  assign n12531 = ~n12529 & n12530 ;
  assign n12532 = ~n12500 & ~n12531 ;
  assign n12533 = \P1_reg2_reg[19]/NET0131  & n12532 ;
  assign n12534 = ~\P1_reg2_reg[19]/NET0131  & ~n12532 ;
  assign n12535 = ~n12533 & ~n12534 ;
  assign n12537 = ~n1408 & ~n12535 ;
  assign n12536 = n1408 & n12535 ;
  assign n12538 = n11437 & ~n12536 ;
  assign n12539 = ~n12537 & n12538 ;
  assign n12514 = ~n12173 & n12179 ;
  assign n12515 = ~n12174 & ~n12484 ;
  assign n12516 = ~n12514 & n12515 ;
  assign n12517 = ~n12485 & ~n12516 ;
  assign n12518 = ~\P1_reg1_reg[19]/NET0131  & ~n1408 ;
  assign n12519 = \P1_reg1_reg[19]/NET0131  & n1408 ;
  assign n12520 = ~n12518 & ~n12519 ;
  assign n12522 = n12517 & n12520 ;
  assign n12521 = ~n12517 & ~n12520 ;
  assign n12523 = n11404 & ~n12521 ;
  assign n12524 = ~n12522 & n12523 ;
  assign n12526 = ~n1408 & ~n11399 ;
  assign n12525 = ~\P1_addr_reg[19]/NET0131  & n11399 ;
  assign n12527 = ~n537 & ~n12525 ;
  assign n12528 = ~n12526 & n12527 ;
  assign n12540 = ~n12524 & ~n12528 ;
  assign n12541 = ~n12539 & n12540 ;
  assign n12542 = \P1_state_reg[0]/NET0131  & ~n12541 ;
  assign n12543 = ~n5685 & ~n12542 ;
  assign n12544 = ~n538 & ~n3448 ;
  assign n12545 = \P1_state_reg[0]/NET0131  & ~n12544 ;
  assign n12546 = ~n2024 & ~n2059 ;
  assign n12547 = \P1_state_reg[0]/NET0131  & ~n12546 ;
  assign n12548 = \P1_state_reg[0]/NET0131  & n3448 ;
  assign n12549 = \P1_state_reg[0]/NET0131  & n2024 ;
  assign n12550 = n2023 & ~n3043 ;
  assign n12551 = \P2_datao_reg[25]/NET0131  & ~n2023 ;
  assign n12552 = ~n12550 & ~n12551 ;
  assign n12553 = ~n1038 & n3447 ;
  assign n12554 = \P1_datao_reg[25]/NET0131  & ~n3447 ;
  assign n12555 = ~n12553 & ~n12554 ;
  assign n12556 = \P2_reg1_reg[16]/NET0131  & ~n5961 ;
  assign n12557 = \P2_reg1_reg[16]/NET0131  & n6642 ;
  assign n12558 = n3355 & n6240 ;
  assign n12561 = n7983 & ~n12558 ;
  assign n12559 = ~n3177 & ~n6226 ;
  assign n12560 = n3411 & n6234 ;
  assign n12562 = ~n12559 & ~n12560 ;
  assign n12563 = n12561 & n12562 ;
  assign n12564 = n3733 & ~n12563 ;
  assign n12565 = ~n12557 & ~n12564 ;
  assign n12566 = n5287 & ~n12565 ;
  assign n12567 = ~n12556 & ~n12566 ;
  assign n12569 = n2024 & n2438 ;
  assign n12571 = n2438 & ~n3788 ;
  assign n12572 = n3788 & n6331 ;
  assign n12573 = ~n12571 & ~n12572 ;
  assign n12574 = n3355 & ~n12573 ;
  assign n12578 = n3788 & ~n6343 ;
  assign n12579 = ~n12571 & ~n12578 ;
  assign n12580 = ~n3320 & ~n12579 ;
  assign n12575 = n3788 & n6337 ;
  assign n12576 = ~n12571 & ~n12575 ;
  assign n12577 = ~n3177 & ~n12576 ;
  assign n12581 = n3788 & n6351 ;
  assign n12582 = ~n12571 & ~n12581 ;
  assign n12583 = n3411 & ~n12582 ;
  assign n12570 = n2438 & ~n3962 ;
  assign n12584 = n2433 & ~n3965 ;
  assign n12585 = ~n12570 & ~n12584 ;
  assign n12586 = ~n12583 & n12585 ;
  assign n12587 = ~n12577 & n12586 ;
  assign n12588 = ~n12580 & n12587 ;
  assign n12589 = ~n12574 & n12588 ;
  assign n12590 = n2026 & ~n12589 ;
  assign n12591 = ~n12569 & ~n12590 ;
  assign n12592 = \P1_state_reg[0]/NET0131  & ~n12591 ;
  assign n12568 = n2438 & n3976 ;
  assign n12593 = ~n12423 & ~n12568 ;
  assign n12594 = ~n12592 & n12593 ;
  assign n12596 = n1002 & ~n3980 ;
  assign n12597 = n3980 & ~n5948 ;
  assign n12598 = ~n12596 & ~n12597 ;
  assign n12599 = ~n3563 & ~n12598 ;
  assign n12606 = n3980 & n5908 ;
  assign n12607 = ~n12596 & ~n12606 ;
  assign n12608 = n3712 & ~n12607 ;
  assign n12595 = n997 & ~n4067 ;
  assign n12609 = n1002 & ~n4064 ;
  assign n12610 = ~n12595 & ~n12609 ;
  assign n12611 = ~n12608 & n12610 ;
  assign n12612 = ~n12599 & n12611 ;
  assign n12600 = n3980 & ~n5930 ;
  assign n12601 = ~n12596 & ~n12600 ;
  assign n12602 = ~n3677 & ~n12601 ;
  assign n12603 = n3980 & ~n5903 ;
  assign n12604 = ~n12596 & ~n12603 ;
  assign n12605 = n1936 & ~n12604 ;
  assign n12613 = ~n12602 & ~n12605 ;
  assign n12614 = n12612 & n12613 ;
  assign n12615 = n5812 & ~n12614 ;
  assign n12616 = \P1_reg3_reg[26]/NET0131  & ~\P1_state_reg[0]/NET0131  ;
  assign n12617 = \P1_state_reg[0]/NET0131  & ~n3450 ;
  assign n12618 = n1002 & n12617 ;
  assign n12619 = ~n12616 & ~n12618 ;
  assign n12620 = ~n12615 & n12619 ;
  assign n12621 = \P2_reg2_reg[15]/NET0131  & ~n1983 ;
  assign n12622 = \P2_reg2_reg[15]/NET0131  & n2024 ;
  assign n12624 = \P2_reg2_reg[15]/NET0131  & ~n3758 ;
  assign n12628 = n3758 & n8217 ;
  assign n12629 = ~n12624 & ~n12628 ;
  assign n12630 = ~n3177 & ~n12629 ;
  assign n12625 = n3758 & n8211 ;
  assign n12626 = ~n12624 & ~n12625 ;
  assign n12627 = n3411 & ~n12626 ;
  assign n12633 = n3758 & n8222 ;
  assign n12634 = ~n12624 & ~n12633 ;
  assign n12635 = n3355 & ~n12634 ;
  assign n12632 = n3758 & ~n9361 ;
  assign n12623 = n2822 & n3420 ;
  assign n12631 = \P2_reg2_reg[15]/NET0131  & ~n7770 ;
  assign n12636 = ~n12623 & ~n12631 ;
  assign n12637 = ~n12632 & n12636 ;
  assign n12638 = ~n12635 & n12637 ;
  assign n12639 = ~n12627 & n12638 ;
  assign n12640 = ~n12630 & n12639 ;
  assign n12641 = n2026 & ~n12640 ;
  assign n12642 = ~n12622 & ~n12641 ;
  assign n12643 = \P1_state_reg[0]/NET0131  & ~n12642 ;
  assign n12644 = ~n12621 & ~n12643 ;
  assign n12645 = \P2_reg2_reg[24]/NET0131  & ~n1983 ;
  assign n12646 = \P2_reg2_reg[24]/NET0131  & n2024 ;
  assign n12647 = \P2_reg2_reg[24]/NET0131  & ~n3758 ;
  assign n12648 = n3758 & ~n4983 ;
  assign n12649 = ~n12647 & ~n12648 ;
  assign n12650 = ~n3320 & ~n12649 ;
  assign n12651 = n3758 & ~n4997 ;
  assign n12652 = ~n12647 & ~n12651 ;
  assign n12653 = ~n3177 & ~n12652 ;
  assign n12657 = n3758 & n5008 ;
  assign n12658 = ~n12647 & ~n12657 ;
  assign n12659 = n3411 & ~n12658 ;
  assign n12654 = n3758 & n5002 ;
  assign n12655 = ~n12647 & ~n12654 ;
  assign n12656 = n3355 & ~n12655 ;
  assign n12660 = n3758 & n5010 ;
  assign n12661 = n3058 & n3420 ;
  assign n12662 = \P2_reg2_reg[24]/NET0131  & ~n3774 ;
  assign n12663 = ~n12661 & ~n12662 ;
  assign n12664 = ~n12660 & n12663 ;
  assign n12665 = ~n12656 & n12664 ;
  assign n12666 = ~n12659 & n12665 ;
  assign n12667 = ~n12653 & n12666 ;
  assign n12668 = ~n12650 & n12667 ;
  assign n12669 = n2026 & ~n12668 ;
  assign n12670 = ~n12646 & ~n12669 ;
  assign n12671 = \P1_state_reg[0]/NET0131  & ~n12670 ;
  assign n12672 = ~n12645 & ~n12671 ;
  assign n12673 = ~\P1_rd_reg/NET0131  & ~\P2_rd_reg/NET0131  ;
  assign n12674 = \P1_rd_reg/NET0131  & \P2_rd_reg/NET0131  ;
  assign n12675 = ~n12673 & ~n12674 ;
  assign n12676 = \P1_addr_reg[0]/NET0131  & \P2_addr_reg[0]/NET0131  ;
  assign n12677 = ~\P1_addr_reg[0]/NET0131  & ~\P2_addr_reg[0]/NET0131  ;
  assign n12678 = ~n12676 & ~n12677 ;
  assign n12679 = \P1_addr_reg[10]/NET0131  & \P2_addr_reg[10]/NET0131  ;
  assign n12680 = ~\P1_addr_reg[10]/NET0131  & ~\P2_addr_reg[10]/NET0131  ;
  assign n12681 = ~n12679 & ~n12680 ;
  assign n12682 = ~\P1_addr_reg[9]/NET0131  & ~\P2_addr_reg[9]/NET0131  ;
  assign n12683 = \P1_addr_reg[9]/NET0131  & \P2_addr_reg[9]/NET0131  ;
  assign n12684 = ~\P1_addr_reg[8]/NET0131  & ~\P2_addr_reg[8]/NET0131  ;
  assign n12685 = \P1_addr_reg[8]/NET0131  & \P2_addr_reg[8]/NET0131  ;
  assign n12686 = ~\P1_addr_reg[7]/NET0131  & ~\P2_addr_reg[7]/NET0131  ;
  assign n12687 = \P1_addr_reg[7]/NET0131  & \P2_addr_reg[7]/NET0131  ;
  assign n12688 = ~\P1_addr_reg[6]/NET0131  & ~\P2_addr_reg[6]/NET0131  ;
  assign n12689 = \P1_addr_reg[6]/NET0131  & \P2_addr_reg[6]/NET0131  ;
  assign n12690 = ~\P1_addr_reg[5]/NET0131  & ~\P2_addr_reg[5]/NET0131  ;
  assign n12691 = \P1_addr_reg[5]/NET0131  & \P2_addr_reg[5]/NET0131  ;
  assign n12692 = ~\P1_addr_reg[4]/NET0131  & ~\P2_addr_reg[4]/NET0131  ;
  assign n12693 = \P1_addr_reg[4]/NET0131  & \P2_addr_reg[4]/NET0131  ;
  assign n12694 = ~\P1_addr_reg[3]/NET0131  & ~\P2_addr_reg[3]/NET0131  ;
  assign n12695 = \P1_addr_reg[3]/NET0131  & \P2_addr_reg[3]/NET0131  ;
  assign n12696 = ~\P1_addr_reg[2]/NET0131  & ~\P2_addr_reg[2]/NET0131  ;
  assign n12697 = \P1_addr_reg[2]/NET0131  & \P2_addr_reg[2]/NET0131  ;
  assign n12698 = ~\P1_addr_reg[1]/NET0131  & ~\P2_addr_reg[1]/NET0131  ;
  assign n12699 = \P1_addr_reg[1]/NET0131  & \P2_addr_reg[1]/NET0131  ;
  assign n12700 = ~n12676 & ~n12699 ;
  assign n12701 = ~n12698 & ~n12700 ;
  assign n12702 = ~n12697 & ~n12701 ;
  assign n12703 = ~n12696 & ~n12702 ;
  assign n12704 = ~n12695 & ~n12703 ;
  assign n12705 = ~n12694 & ~n12704 ;
  assign n12706 = ~n12693 & ~n12705 ;
  assign n12707 = ~n12692 & ~n12706 ;
  assign n12708 = ~n12691 & ~n12707 ;
  assign n12709 = ~n12690 & ~n12708 ;
  assign n12710 = ~n12689 & ~n12709 ;
  assign n12711 = ~n12688 & ~n12710 ;
  assign n12712 = ~n12687 & ~n12711 ;
  assign n12713 = ~n12686 & ~n12712 ;
  assign n12714 = ~n12685 & ~n12713 ;
  assign n12715 = ~n12684 & ~n12714 ;
  assign n12716 = ~n12683 & ~n12715 ;
  assign n12717 = ~n12682 & ~n12716 ;
  assign n12718 = ~n12681 & n12717 ;
  assign n12719 = n12681 & ~n12717 ;
  assign n12720 = ~n12718 & ~n12719 ;
  assign n12721 = \P1_addr_reg[11]/NET0131  & \P2_addr_reg[11]/NET0131  ;
  assign n12722 = ~\P1_addr_reg[11]/NET0131  & ~\P2_addr_reg[11]/NET0131  ;
  assign n12723 = ~n12721 & ~n12722 ;
  assign n12724 = ~n12679 & ~n12717 ;
  assign n12725 = ~n12680 & ~n12724 ;
  assign n12726 = ~n12723 & n12725 ;
  assign n12727 = n12723 & ~n12725 ;
  assign n12728 = ~n12726 & ~n12727 ;
  assign n12729 = \P1_addr_reg[12]/NET0131  & \P2_addr_reg[12]/NET0131  ;
  assign n12730 = ~\P1_addr_reg[12]/NET0131  & ~\P2_addr_reg[12]/NET0131  ;
  assign n12731 = ~n12729 & ~n12730 ;
  assign n12732 = ~n12721 & ~n12725 ;
  assign n12733 = ~n12722 & ~n12732 ;
  assign n12734 = ~n12731 & n12733 ;
  assign n12735 = n12731 & ~n12733 ;
  assign n12736 = ~n12734 & ~n12735 ;
  assign n12737 = \P1_addr_reg[13]/NET0131  & \P2_addr_reg[13]/NET0131  ;
  assign n12738 = ~\P1_addr_reg[13]/NET0131  & ~\P2_addr_reg[13]/NET0131  ;
  assign n12739 = ~n12737 & ~n12738 ;
  assign n12740 = ~n12729 & ~n12733 ;
  assign n12741 = ~n12730 & ~n12740 ;
  assign n12742 = ~n12739 & n12741 ;
  assign n12743 = n12739 & ~n12741 ;
  assign n12744 = ~n12742 & ~n12743 ;
  assign n12745 = \P1_addr_reg[14]/NET0131  & \P2_addr_reg[14]/NET0131  ;
  assign n12746 = ~\P1_addr_reg[14]/NET0131  & ~\P2_addr_reg[14]/NET0131  ;
  assign n12747 = ~n12745 & ~n12746 ;
  assign n12748 = ~n12737 & ~n12741 ;
  assign n12749 = ~n12738 & ~n12748 ;
  assign n12750 = ~n12747 & n12749 ;
  assign n12751 = n12747 & ~n12749 ;
  assign n12752 = ~n12750 & ~n12751 ;
  assign n12753 = \P1_addr_reg[15]/NET0131  & \P2_addr_reg[15]/NET0131  ;
  assign n12754 = ~\P1_addr_reg[15]/NET0131  & ~\P2_addr_reg[15]/NET0131  ;
  assign n12755 = ~n12753 & ~n12754 ;
  assign n12756 = ~n12745 & ~n12749 ;
  assign n12757 = ~n12746 & ~n12756 ;
  assign n12758 = ~n12755 & n12757 ;
  assign n12759 = n12755 & ~n12757 ;
  assign n12760 = ~n12758 & ~n12759 ;
  assign n12761 = \P1_addr_reg[16]/NET0131  & \P2_addr_reg[16]/NET0131  ;
  assign n12762 = ~\P1_addr_reg[16]/NET0131  & ~\P2_addr_reg[16]/NET0131  ;
  assign n12763 = ~n12761 & ~n12762 ;
  assign n12764 = ~n12753 & ~n12757 ;
  assign n12765 = ~n12754 & ~n12764 ;
  assign n12766 = ~n12763 & n12765 ;
  assign n12767 = n12763 & ~n12765 ;
  assign n12768 = ~n12766 & ~n12767 ;
  assign n12769 = \P1_addr_reg[17]/NET0131  & \P2_addr_reg[17]/NET0131  ;
  assign n12770 = ~\P1_addr_reg[17]/NET0131  & ~\P2_addr_reg[17]/NET0131  ;
  assign n12771 = ~n12769 & ~n12770 ;
  assign n12772 = ~n12761 & ~n12765 ;
  assign n12773 = ~n12762 & ~n12772 ;
  assign n12774 = ~n12771 & n12773 ;
  assign n12775 = n12771 & ~n12773 ;
  assign n12776 = ~n12774 & ~n12775 ;
  assign n12777 = \P1_addr_reg[18]/NET0131  & \P2_addr_reg[18]/NET0131  ;
  assign n12778 = ~\P1_addr_reg[18]/NET0131  & ~\P2_addr_reg[18]/NET0131  ;
  assign n12779 = ~n12777 & ~n12778 ;
  assign n12780 = ~n12769 & ~n12773 ;
  assign n12781 = ~n12770 & ~n12780 ;
  assign n12782 = ~n12779 & n12781 ;
  assign n12783 = n12779 & ~n12781 ;
  assign n12784 = ~n12782 & ~n12783 ;
  assign n12785 = ~n539 & ~n541 ;
  assign n12786 = ~n12777 & ~n12781 ;
  assign n12787 = ~n12778 & ~n12786 ;
  assign n12788 = n12785 & ~n12787 ;
  assign n12789 = ~n12785 & n12787 ;
  assign n12790 = ~n12788 & ~n12789 ;
  assign n12791 = ~n12698 & ~n12699 ;
  assign n12792 = n12676 & ~n12791 ;
  assign n12793 = ~n12676 & n12791 ;
  assign n12794 = ~n12792 & ~n12793 ;
  assign n12795 = ~n12696 & ~n12697 ;
  assign n12796 = n12701 & ~n12795 ;
  assign n12797 = ~n12701 & n12795 ;
  assign n12798 = ~n12796 & ~n12797 ;
  assign n12799 = ~n12694 & ~n12695 ;
  assign n12800 = n12703 & ~n12799 ;
  assign n12801 = ~n12703 & n12799 ;
  assign n12802 = ~n12800 & ~n12801 ;
  assign n12803 = ~n12692 & ~n12693 ;
  assign n12804 = n12705 & ~n12803 ;
  assign n12805 = ~n12705 & n12803 ;
  assign n12806 = ~n12804 & ~n12805 ;
  assign n12807 = ~n12690 & ~n12691 ;
  assign n12808 = n12707 & ~n12807 ;
  assign n12809 = ~n12707 & n12807 ;
  assign n12810 = ~n12808 & ~n12809 ;
  assign n12811 = ~n12688 & ~n12689 ;
  assign n12812 = n12709 & ~n12811 ;
  assign n12813 = ~n12709 & n12811 ;
  assign n12814 = ~n12812 & ~n12813 ;
  assign n12815 = ~n12686 & ~n12687 ;
  assign n12816 = n12711 & ~n12815 ;
  assign n12817 = ~n12711 & n12815 ;
  assign n12818 = ~n12816 & ~n12817 ;
  assign n12819 = ~n12684 & ~n12685 ;
  assign n12820 = n12713 & ~n12819 ;
  assign n12821 = ~n12713 & n12819 ;
  assign n12822 = ~n12820 & ~n12821 ;
  assign n12823 = ~n12682 & ~n12683 ;
  assign n12824 = n12715 & ~n12823 ;
  assign n12825 = ~n12715 & n12823 ;
  assign n12826 = ~n12824 & ~n12825 ;
  assign n12827 = ~\P1_wr_reg/NET0131  & ~\P2_wr_reg/NET0131  ;
  assign n12828 = \P1_wr_reg/NET0131  & \P2_wr_reg/NET0131  ;
  assign n12829 = ~n12827 & ~n12828 ;
  assign \P1_state_reg[0]/NET0131_syn_2  = ~\P1_state_reg[0]/NET0131  ;
  assign \_al_n0  = 1'b0 ;
  assign \_al_n1  = ~1'b0 ;
  assign \g73521/_0_  = ~n1956 ;
  assign \g73537/_0_  = ~n3434 ;
  assign \g73538/_0_  = ~n3730 ;
  assign \g73539/_0_  = ~n3755 ;
  assign \g73540/_0_  = ~n3786 ;
  assign \g73570/_0_  = ~n3979 ;
  assign \g73571/_0_  = ~n4117 ;
  assign \g73572/_0_  = ~n4327 ;
  assign \g73573/_0_  = ~n4350 ;
  assign \g73574/_0_  = ~n4368 ;
  assign \g73575/_0_  = ~n4393 ;
  assign \g73576/_0_  = ~n4503 ;
  assign \g73577/_0_  = ~n4529 ;
  assign \g73578/_0_  = ~n4558 ;
  assign \g73579/_0_  = ~n4582 ;
  assign \g73609/_0_  = ~n4643 ;
  assign \g73610/_0_  = ~n4702 ;
  assign \g73611/_0_  = ~n4797 ;
  assign \g73613/_0_  = ~n4895 ;
  assign \g73614/_0_  = ~n4923 ;
  assign \g73615/_0_  = ~n4949 ;
  assign \g73617/_0_  = ~n4974 ;
  assign \g73618/_0_  = ~n5021 ;
  assign \g73619/_0_  = ~n5048 ;
  assign \g73620/_0_  = ~n5078 ;
  assign \g73621/_0_  = ~n5096 ;
  assign \g73622/_0_  = ~n5114 ;
  assign \g73623/_0_  = ~n5132 ;
  assign \g73624/_0_  = ~n5158 ;
  assign \g73625/_0_  = ~n5217 ;
  assign \g73626/_0_  = ~n5246 ;
  assign \g73627/_0_  = ~n5274 ;
  assign \g73628/_0_  = ~n5294 ;
  assign \g73629/_0_  = ~n5321 ;
  assign \g73630/_0_  = ~n5347 ;
  assign \g73631/_0_  = ~n5373 ;
  assign \g73632/_0_  = ~n5399 ;
  assign \g73633/_0_  = ~n5425 ;
  assign \g73692/_0_  = ~n5475 ;
  assign \g73693/_0_  = ~n5550 ;
  assign \g73694/_0_  = ~n5600 ;
  assign \g73696/_0_  = ~n5644 ;
  assign \g73697/_0_  = ~n5688 ;
  assign \g73703/_0_  = ~n5716 ;
  assign \g73704/_0_  = ~n5744 ;
  assign \g73709/_0_  = ~n5793 ;
  assign \g73710/_0_  = ~n5818 ;
  assign \g73711/_0_  = ~n5841 ;
  assign \g73712/_0_  = ~n5859 ;
  assign \g73713/_0_  = ~n5866 ;
  assign \g73714/_0_  = ~n5894 ;
  assign \g73715/_0_  = ~n5960 ;
  assign \g73716/_0_  = ~n5966 ;
  assign \g73717/_0_  = ~n5992 ;
  assign \g73718/_0_  = ~n6014 ;
  assign \g73719/_0_  = ~n6066 ;
  assign \g73720/_0_  = ~n6088 ;
  assign \g73774/_0_  = ~n6131 ;
  assign \g73775/_0_  = ~n6173 ;
  assign \g73776/_0_  = ~n6216 ;
  assign \g73777/_0_  = ~n6259 ;
  assign \g73806/_0_  = ~n6285 ;
  assign \g73807/_0_  = ~n6325 ;
  assign \g73808/_0_  = ~n6367 ;
  assign \g73809/_0_  = ~n6372 ;
  assign \g73810/_0_  = ~n6395 ;
  assign \g73811/_0_  = ~n6424 ;
  assign \g73812/_0_  = ~n6453 ;
  assign \g73813/_0_  = ~n6483 ;
  assign \g73814/_0_  = ~n6526 ;
  assign \g73815/_0_  = ~n6553 ;
  assign \g73816/_0_  = ~n6583 ;
  assign \g73817/_0_  = ~n6609 ;
  assign \g73818/_0_  = ~n6636 ;
  assign \g73819/_0_  = ~n6654 ;
  assign \g73820/_0_  = ~n6672 ;
  assign \g73821/_0_  = ~n6700 ;
  assign \g73822/_0_  = ~n6728 ;
  assign \g73823/_0_  = ~n6770 ;
  assign \g73824/_0_  = ~n6790 ;
  assign \g73825/_0_  = ~n6816 ;
  assign \g73826/_0_  = ~n6842 ;
  assign \g73827/_0_  = ~n6863 ;
  assign \g73828/_0_  = ~n6885 ;
  assign \g73829/_0_  = ~n6890 ;
  assign \g73830/_0_  = ~n6916 ;
  assign \g73831/_0_  = ~n6942 ;
  assign \g73832/_0_  = ~n6952 ;
  assign \g73833/_0_  = ~n6992 ;
  assign \g73834/_0_  = ~n7018 ;
  assign \g73835/_0_  = ~n7044 ;
  assign \g73836/_0_  = ~n7070 ;
  assign \g73908/_0_  = ~n7111 ;
  assign \g73909/_0_  = ~n7153 ;
  assign \g73911/_0_  = ~n7195 ;
  assign \g73912/_0_  = ~n7237 ;
  assign \g73915/_0_  = ~n7280 ;
  assign \g73916/_0_  = ~n7324 ;
  assign \g73946/_0_  = ~n7352 ;
  assign \g73950/_0_  = ~n7380 ;
  assign \g73957/_0_  = ~n7408 ;
  assign \g73958/_0_  = ~n7462 ;
  assign \g73959/_0_  = ~n7488 ;
  assign \g73960/_0_  = ~n7503 ;
  assign \g73961/_0_  = ~n7514 ;
  assign \g73962/_0_  = ~n7543 ;
  assign \g73963/_0_  = ~n7552 ;
  assign \g73964/_0_  = ~n7581 ;
  assign \g73965/_0_  = ~n7607 ;
  assign \g73966/_0_  = ~n7635 ;
  assign \g73968/_0_  = ~n7664 ;
  assign \g73969/_0_  = ~n7690 ;
  assign \g73970/_0_  = ~n7693 ;
  assign \g73971/_0_  = ~n7707 ;
  assign \g73972/_0_  = ~n7735 ;
  assign \g73973/_0_  = ~n7764 ;
  assign \g73974/_0_  = ~n7775 ;
  assign \g73975/_0_  = ~n7790 ;
  assign \g73976/_0_  = ~n7816 ;
  assign \g73977/_0_  = ~n7832 ;
  assign \g73978/_0_  = ~n7858 ;
  assign \g73979/_0_  = ~n7884 ;
  assign \g73980/_0_  = ~n7887 ;
  assign \g73981/_0_  = ~n7913 ;
  assign \g73982/_0_  = ~n7924 ;
  assign \g73983/_0_  = ~n7950 ;
  assign \g73984/_0_  = ~n7972 ;
  assign \g73985/_0_  = ~n7996 ;
  assign \g74044/_0_  = ~n8036 ;
  assign \g74045/_0_  = ~n8080 ;
  assign \g74046/_0_  = ~n8120 ;
  assign \g74047/_0_  = ~n8160 ;
  assign \g74048/_0_  = ~n8201 ;
  assign \g74049/_0_  = ~n8242 ;
  assign \g74051/_0_  = ~n8282 ;
  assign \g74052/_0_  = ~n8324 ;
  assign \g74099/_0_  = ~n8369 ;
  assign \g74100/_0_  = ~n8393 ;
  assign \g74101/_0_  = ~n8420 ;
  assign \g74102/_0_  = ~n8449 ;
  assign \g74103/_0_  = ~n8478 ;
  assign \g74104/_0_  = ~n8500 ;
  assign \g74105/_0_  = ~n8527 ;
  assign \g74106/_0_  = ~n8550 ;
  assign \g74107/_0_  = ~n8568 ;
  assign \g74108/_0_  = ~n8594 ;
  assign \g74109/_0_  = ~n8612 ;
  assign \g74110/_0_  = ~n8640 ;
  assign \g74111/_0_  = ~n8664 ;
  assign \g74112/_0_  = ~n8692 ;
  assign \g74113/_0_  = ~n8713 ;
  assign \g74114/_0_  = ~n8741 ;
  assign \g74115/_0_  = ~n8767 ;
  assign \g74116/_0_  = ~n8790 ;
  assign \g74117/_0_  = ~n8816 ;
  assign \g74118/_0_  = ~n8842 ;
  assign \g74119/_0_  = ~n8868 ;
  assign \g74120/_0_  = ~n8894 ;
  assign \g74121/_0_  = ~n8912 ;
  assign \g74122/_0_  = ~n8934 ;
  assign \g74199/_0_  = ~n8976 ;
  assign \g74200/_0_  = ~n9015 ;
  assign \g74201/_0_  = ~n9057 ;
  assign \g74202/_0_  = ~n9103 ;
  assign \g74279/_0_  = ~n9130 ;
  assign \g74280/_0_  = ~n9156 ;
  assign \g74284/_0_  = ~n9183 ;
  assign \g74285/_0_  = ~n9209 ;
  assign \g74287/_0_  = ~n9238 ;
  assign \g74288/_0_  = ~n9264 ;
  assign \g74289/_0_  = ~n9290 ;
  assign \g74290/_0_  = ~n9317 ;
  assign \g74291/_0_  = ~n9343 ;
  assign \g74292/_0_  = ~n9356 ;
  assign \g74293/_0_  = ~n9381 ;
  assign \g74294/_0_  = ~n9390 ;
  assign \g74295/_0_  = ~n9419 ;
  assign \g74296/_0_  = ~n9448 ;
  assign \g74298/_0_  = ~n9476 ;
  assign \g74299/_0_  = ~n9498 ;
  assign \g74300/_0_  = ~n9524 ;
  assign \g74301/_0_  = ~n9552 ;
  assign \g74302/_0_  = ~n9574 ;
  assign \g74382/_0_  = ~n9614 ;
  assign \g74383/_0_  = ~n9655 ;
  assign \g74384/_0_  = ~n9695 ;
  assign \g74385/_0_  = ~n9739 ;
  assign \g74386/_0_  = ~n9780 ;
  assign \g74387/_0_  = ~n9820 ;
  assign \g74456/_0_  = ~n9844 ;
  assign \g74457/_0_  = ~n9854 ;
  assign \g74458/_0_  = ~n9875 ;
  assign \g74459/_0_  = ~n9901 ;
  assign \g74460/_0_  = ~n9910 ;
  assign \g74461/_0_  = ~n9938 ;
  assign \g74462/_0_  = ~n9964 ;
  assign \g74463/_0_  = ~n9986 ;
  assign \g74464/_0_  = ~n10014 ;
  assign \g74465/_0_  = ~n10024 ;
  assign \g74466/_0_  = ~n10048 ;
  assign \g74467/_0_  = ~n10076 ;
  assign \g74468/_0_  = ~n10104 ;
  assign \g74469/_0_  = ~n10128 ;
  assign \g74470/_0_  = ~n10146 ;
  assign \g74471/_0_  = ~n10172 ;
  assign \g74661/_0_  = ~n10194 ;
  assign \g74662/_0_  = ~n10218 ;
  assign \g74663/_0_  = ~n10238 ;
  assign \g74664/_0_  = ~n10260 ;
  assign \g74665/_0_  = ~n10278 ;
  assign \g74666/_0_  = ~n10296 ;
  assign \g74667/_0_  = ~n10320 ;
  assign \g74668/_0_  = ~n10349 ;
  assign \g74669/_0_  = ~n10373 ;
  assign \g74670/_0_  = ~n10394 ;
  assign \g74671/_0_  = ~n10423 ;
  assign \g74672/_0_  = ~n10451 ;
  assign \g74673/_0_  = ~n10471 ;
  assign \g74674/_0_  = ~n10499 ;
  assign \g74899/_0_  = ~n10525 ;
  assign \g74900/_0_  = ~n10551 ;
  assign \g74901/_0_  = ~n10577 ;
  assign \g74902/_0_  = ~n10603 ;
  assign \g75002/_0_  = ~n10642 ;
  assign \g75005/_0_  = ~n10681 ;
  assign \g75191/_0_  = ~n10708 ;
  assign \g75192/_0_  = ~n10734 ;
  assign \g75193/_0_  = ~n10763 ;
  assign \g75194/_0_  = ~n10789 ;
  assign \g75195/_0_  = ~n10815 ;
  assign \g75392/_0_  = ~n10853 ;
  assign \g75399/_0_  = ~n10891 ;
  assign \g75606/_0_  = ~n10915 ;
  assign \g75607/_0_  = ~n10937 ;
  assign \g75608/_0_  = ~n10965 ;
  assign \g75609/_0_  = ~n10989 ;
  assign \g75610/_0_  = ~n11011 ;
  assign \g76007/_0_  = ~n11041 ;
  assign \g76008/_0_  = ~n11065 ;
  assign \g76685/_0_  = ~n11089 ;
  assign \g76696/_0_  = ~n11114 ;
  assign \g77574/_0_  = n11130 ;
  assign \g77575/_0_  = ~n11150 ;
  assign \g77576/_0_  = ~n11161 ;
  assign \g77577/_0_  = ~n11181 ;
  assign \g77578/_0_  = ~n11187 ;
  assign \g77579/_0_  = ~n11207 ;
  assign \g82699/_3_  = ~n11210 ;
  assign \g82700/_3_  = ~n11213 ;
  assign \g82701/_3_  = ~n11216 ;
  assign \g82702/_3_  = ~n11219 ;
  assign \g82703/_3_  = ~n11222 ;
  assign \g82704/_3_  = ~n11225 ;
  assign \g83319/_0_  = ~n11228 ;
  assign \g83320/_0_  = n11231 ;
  assign \g83321/_0_  = n11234 ;
  assign \g83322/_0_  = ~n11237 ;
  assign \g83323/_3_  = n11240 ;
  assign \g83324/_0_  = ~n11243 ;
  assign \g83325/_0_  = n11246 ;
  assign \g83326/_0_  = n11249 ;
  assign \g83327/_0_  = n11252 ;
  assign \g83328/_0_  = ~n11255 ;
  assign \g83329/_0_  = ~n11258 ;
  assign \g83330/_0_  = ~n11261 ;
  assign \g83331/_0_  = ~n11264 ;
  assign \g83332/_0_  = ~n11267 ;
  assign \g83333/_0_  = ~n11269 ;
  assign \g83334/_0_  = ~n11272 ;
  assign \g83335/_0_  = n11275 ;
  assign \g83336/_3_  = ~n11278 ;
  assign \g83337/_0_  = ~n11281 ;
  assign \g83338/_0_  = n11284 ;
  assign \g83339/_0_  = ~n11287 ;
  assign \g83340/_0_  = ~n11290 ;
  assign \g83341/_0_  = ~n11293 ;
  assign \g83342/_0_  = n11296 ;
  assign \g83343/_0_  = n11299 ;
  assign \g83344/_0_  = ~n11302 ;
  assign \g83345/_0_  = ~n11305 ;
  assign \g83347/_3_  = n11308 ;
  assign \g83348/_3_  = ~n11311 ;
  assign \g83349/_3_  = n11314 ;
  assign \g83350/_3_  = n11317 ;
  assign \g83351/_3_  = ~n11320 ;
  assign \g83352/_3_  = ~n11323 ;
  assign \g83353/_3_  = ~n11326 ;
  assign \g83354/_3_  = ~n11329 ;
  assign \g83355/_3_  = n11332 ;
  assign \g83356/_3_  = ~n11335 ;
  assign \g83357/_0_  = ~n11338 ;
  assign \g83358/_3_  = n11341 ;
  assign \g83359/_3_  = ~n11344 ;
  assign \g83360/_3_  = ~n11346 ;
  assign \g83361/_3_  = ~n11349 ;
  assign \g83362/_3_  = ~n11352 ;
  assign \g83363/_3_  = ~n11355 ;
  assign \g83364/_3_  = ~n11358 ;
  assign \g83365/_0_  = ~n11361 ;
  assign \g83366/_3_  = ~n11364 ;
  assign \g83367/_0_  = ~n11370 ;
  assign \g83368/_3_  = ~n11373 ;
  assign \g83369/_3_  = ~n11376 ;
  assign \g83370/_0_  = ~n11379 ;
  assign \g83371/_3_  = ~n11382 ;
  assign \g83372/_3_  = ~n11385 ;
  assign \g83373/_3_  = ~n11388 ;
  assign \g83374/_3_  = ~n11391 ;
  assign \g83376/_0_  = ~n11398 ;
  assign \g83778/_0_  = n1668 ;
  assign \g83784/_0_  = n2601 ;
  assign \g84388/_0_  = ~n11473 ;
  assign \g84389/_0_  = ~n11507 ;
  assign \g84391/_0_  = ~n11525 ;
  assign \g84395/_0_  = ~n11547 ;
  assign \g84397/_0_  = ~n11567 ;
  assign \g84398/_0_  = ~n11617 ;
  assign \g84399/_0_  = ~n11639 ;
  assign \g84400/_0_  = ~n11656 ;
  assign \g84401/_0_  = ~n11684 ;
  assign \g84402/_0_  = ~n11702 ;
  assign \g84403/_0_  = ~n11728 ;
  assign \g84405/_0_  = ~n11823 ;
  assign \g84406/_0_  = ~n11853 ;
  assign \g84407/_0_  = ~n11895 ;
  assign \g84408/_0_  = ~n11925 ;
  assign \g84409/_0_  = ~n11955 ;
  assign \g84410/_0_  = ~n11986 ;
  assign \g84411/_0_  = ~n12016 ;
  assign \g84412/_0_  = ~n12046 ;
  assign \g84413/_0_  = ~n12076 ;
  assign \g84414/_0_  = ~n12106 ;
  assign \g84415/_0_  = ~n12136 ;
  assign \g84416/_0_  = ~n12157 ;
  assign \g84417/_0_  = ~n12187 ;
  assign \g84418/_0_  = ~n12208 ;
  assign \g84419/_0_  = ~n12228 ;
  assign \g84420/_0_  = ~n12249 ;
  assign \g84421/_0_  = ~n12269 ;
  assign \g84422/_0_  = ~n12287 ;
  assign \g84423/_0_  = ~n12305 ;
  assign \g84424/_0_  = ~n12323 ;
  assign \g84425/_0_  = ~n12343 ;
  assign \g84426/_0_  = ~n12361 ;
  assign \g84427/_0_  = ~n12382 ;
  assign \g84429/_0_  = ~n12402 ;
  assign \g84430/_0_  = ~n12422 ;
  assign \g84442/_0_  = ~n12453 ;
  assign \g84443/_0_  = ~n12483 ;
  assign \g84444/_0_  = ~n12513 ;
  assign \g84445/_0_  = ~n12543 ;
  assign \g84908/_0_  = ~n12545 ;
  assign \g84961/_0_  = ~n12547 ;
  assign \g84984/u3_syn_4  = n5812 ;
  assign \g84985/u3_syn_4  = n5287 ;
  assign \g85802/_0_  = ~n3460 ;
  assign \g86055/_1_  = ~n2035 ;
  assign \g86073/_0_  = ~n3465 ;
  assign \g86298/u3_syn_4  = n12548 ;
  assign \g86300/u3_syn_4  = n12549 ;
  assign \g87397/_0_  = ~n12552 ;
  assign \g87409/_0_  = ~n12555 ;
  assign \g87480/_0_  = ~n887 ;
  assign \g87494/_0_  = ~n831 ;
  assign \g87544/_0_  = ~n750 ;
  assign \g87555/_0_  = ~n2251 ;
  assign \g87567/_0_  = ~n3372 ;
  assign \g87576/_0_  = ~n3402 ;
  assign \g87894/_0_  = ~n1475 ;
  assign \g87905/_0_  = ~n3021 ;
  assign \g87914/_0_  = ~n978 ;
  assign \g87955/_1_  = ~n1062 ;
  assign \g88030/_0_  = ~n1524 ;
  assign \g88039/_0_  = ~n1244 ;
  assign \g88054/_0_  = ~n1267 ;
  assign \g88079/_0_  = ~n2828 ;
  assign \g88094/_0_  = ~n945 ;
  assign \g88111/_0_  = ~n1498 ;
  assign \g88122/_0_  = ~n1664 ;
  assign \g88129/_0_  = ~n1427 ;
  assign \g88162/_0_  = ~n1174 ;
  assign \g88185/_0_  = ~n2715 ;
  assign \g88196/_0_  = ~n2880 ;
  assign \g88204/_0_  = ~n1118 ;
  assign \g88220/_0_  = ~n1218 ;
  assign \g88226/_0_  = ~n2597 ;
  assign \g88243/_0_  = ~n1548 ;
  assign \g88252/_0_  = ~n2531 ;
  assign \g88261/_0_  = ~n2506 ;
  assign \g88269/_0_  = ~n2742 ;
  assign \g88288/_0_  = ~n2379 ;
  assign \g88299/_0_  = ~n2442 ;
  assign \g88310/_0_  = ~n2962 ;
  assign \g88321/_0_  = ~n3130 ;
  assign \g88328/_0_  = ~n3112 ;
  assign \g88335/_0_  = ~n3088 ;
  assign \g88356/_0_  = ~n2454 ;
  assign \g88366/_0_  = ~n2688 ;
  assign \g88372/_0_  = ~n2552 ;
  assign \g88380/_0_  = ~n2311 ;
  assign \g88395_dup/_0_  = ~n2574 ;
  assign \g88403/_0_  = ~n2991 ;
  assign \g88414/_0_  = ~n2368 ;
  assign \g88425/_0_  = ~n1146 ;
  assign \g88443/_0_  = ~n1374 ;
  assign \g88453/_0_  = ~n1318 ;
  assign \g88471/_0_  = ~n1336 ;
  assign \g88524/_0_  = ~n1356 ;
  assign \g88546/_0_  = ~n1006 ;
  assign \g88556/_0_  = ~n2765 ;
  assign \g88563/_0_  = ~n1207 ;
  assign \g89966/_1_  = n3435 ;
  assign \g89999/_1_  = n1983 ;
  assign \g95209/_0_  = ~n12567 ;
  assign \g95269/_0_  = ~n2642 ;
  assign \g95319/_0_  = ~n12594 ;
  assign \g95354/_0_  = ~n2804 ;
  assign \g95786/_0_  = ~n2616 ;
  assign \g95909/_0_  = ~n1595 ;
  assign \g95914/_0_  = ~n1572 ;
  assign \g95918/_0_  = ~n1617 ;
  assign \g95984/_0_  = ~n2870 ;
  assign \g96009/_0_  = ~n3065 ;
  assign \g96124/_0_  = ~n1094 ;
  assign \g96218/_0_  = ~n1452 ;
  assign \g96286/_0_  = ~n1641 ;
  assign \g96335/_0_  = ~n2480 ;
  assign \g96465/_0_  = ~n2039 ;
  assign \g96694/_0_  = ~n12620 ;
  assign \g96713/_0_  = ~n1403 ;
  assign \g96830/_0_  = ~n12644 ;
  assign \g96875/_0_  = ~n12672 ;
  assign rd_pad = ~n12675 ;
  assign \so[0]_pad  = n12678 ;
  assign \so[10]_pad  = ~n12720 ;
  assign \so[11]_pad  = ~n12728 ;
  assign \so[12]_pad  = ~n12736 ;
  assign \so[13]_pad  = ~n12744 ;
  assign \so[14]_pad  = ~n12752 ;
  assign \so[15]_pad  = ~n12760 ;
  assign \so[16]_pad  = ~n12768 ;
  assign \so[17]_pad  = ~n12776 ;
  assign \so[18]_pad  = ~n12784 ;
  assign \so[19]_pad  = ~n12790 ;
  assign \so[1]_pad  = ~n12794 ;
  assign \so[2]_pad  = ~n12798 ;
  assign \so[3]_pad  = ~n12802 ;
  assign \so[4]_pad  = ~n12806 ;
  assign \so[5]_pad  = ~n12810 ;
  assign \so[6]_pad  = ~n12814 ;
  assign \so[7]_pad  = ~n12818 ;
  assign \so[8]_pad  = ~n12822 ;
  assign \so[9]_pad  = ~n12826 ;
  assign wr_pad = ~n12829 ;
endmodule
