module top( \a[0]  , \a[1]  , \a[2]  , \a[3]  , \a[4]  , \a[5]  , \a[6]  , \a[7]  , \a[8]  , \a[9]  , \a[10]  , \a[11]  , \a[12]  , \a[13]  , \a[14]  , \a[15]  , \a[16]  , \a[17]  , \a[18]  , \a[19]  , \a[20]  , \a[21]  , \a[22]  , \a[23]  , \a[24]  , \a[25]  , \a[26]  , \a[27]  , \a[28]  , \a[29]  , \a[30]  , \a[31]  , \a[32]  , \a[33]  , \a[34]  , \a[35]  , \a[36]  , \a[37]  , \a[38]  , \a[39]  , \a[40]  , \a[41]  , \a[42]  , \a[43]  , \a[44]  , \a[45]  , \a[46]  , \a[47]  , \a[48]  , \a[49]  , \a[50]  , \a[51]  , \a[52]  , \a[53]  , \a[54]  , \a[55]  , \a[56]  , \a[57]  , \a[58]  , \a[59]  , \a[60]  , \a[61]  , \a[62]  , \a[63]  , \a[64]  , \a[65]  , \a[66]  , \a[67]  , \a[68]  , \a[69]  , \a[70]  , \a[71]  , \a[72]  , \a[73]  , \a[74]  , \a[75]  , \a[76]  , \a[77]  , \a[78]  , \a[79]  , \a[80]  , \a[81]  , \a[82]  , \a[83]  , \a[84]  , \a[85]  , \a[86]  , \a[87]  , \a[88]  , \a[89]  , \a[90]  , \a[91]  , \a[92]  , \a[93]  , \a[94]  , \a[95]  , \a[96]  , \a[97]  , \a[98]  , \a[99]  , \a[100]  , \a[101]  , \a[102]  , \a[103]  , \a[104]  , \a[105]  , \a[106]  , \a[107]  , \a[108]  , \a[109]  , \a[110]  , \a[111]  , \a[112]  , \a[113]  , \a[114]  , \a[115]  , \a[116]  , \a[117]  , \a[118]  , \a[119]  , \a[120]  , \a[121]  , \a[122]  , \a[123]  , \a[124]  , \a[125]  , \a[126]  , \a[127]  , \shift[0]  , \shift[1]  , \shift[2]  , \shift[3]  , \shift[4]  , \shift[5]  , \shift[6]  , \result[0]  , \result[1]  , \result[2]  , \result[3]  , \result[4]  , \result[5]  , \result[6]  , \result[7]  , \result[8]  , \result[9]  , \result[10]  , \result[11]  , \result[12]  , \result[13]  , \result[14]  , \result[15]  , \result[16]  , \result[17]  , \result[18]  , \result[19]  , \result[20]  , \result[21]  , \result[22]  , \result[23]  , \result[24]  , \result[25]  , \result[26]  , \result[27]  , \result[28]  , \result[29]  , \result[30]  , \result[31]  , \result[32]  , \result[33]  , \result[34]  , \result[35]  , \result[36]  , \result[37]  , \result[38]  , \result[39]  , \result[40]  , \result[41]  , \result[42]  , \result[43]  , \result[44]  , \result[45]  , \result[46]  , \result[47]  , \result[48]  , \result[49]  , \result[50]  , \result[51]  , \result[52]  , \result[53]  , \result[54]  , \result[55]  , \result[56]  , \result[57]  , \result[58]  , \result[59]  , \result[60]  , \result[61]  , \result[62]  , \result[63]  , \result[64]  , \result[65]  , \result[66]  , \result[67]  , \result[68]  , \result[69]  , \result[70]  , \result[71]  , \result[72]  , \result[73]  , \result[74]  , \result[75]  , \result[76]  , \result[77]  , \result[78]  , \result[79]  , \result[80]  , \result[81]  , \result[82]  , \result[83]  , \result[84]  , \result[85]  , \result[86]  , \result[87]  , \result[88]  , \result[89]  , \result[90]  , \result[91]  , \result[92]  , \result[93]  , \result[94]  , \result[95]  , \result[96]  , \result[97]  , \result[98]  , \result[99]  , \result[100]  , \result[101]  , \result[102]  , \result[103]  , \result[104]  , \result[105]  , \result[106]  , \result[107]  , \result[108]  , \result[109]  , \result[110]  , \result[111]  , \result[112]  , \result[113]  , \result[114]  , \result[115]  , \result[116]  , \result[117]  , \result[118]  , \result[119]  , \result[120]  , \result[121]  , \result[122]  , \result[123]  , \result[124]  , \result[125]  , \result[126]  , \result[127]  );
  input \a[0]  ;
  input \a[1]  ;
  input \a[2]  ;
  input \a[3]  ;
  input \a[4]  ;
  input \a[5]  ;
  input \a[6]  ;
  input \a[7]  ;
  input \a[8]  ;
  input \a[9]  ;
  input \a[10]  ;
  input \a[11]  ;
  input \a[12]  ;
  input \a[13]  ;
  input \a[14]  ;
  input \a[15]  ;
  input \a[16]  ;
  input \a[17]  ;
  input \a[18]  ;
  input \a[19]  ;
  input \a[20]  ;
  input \a[21]  ;
  input \a[22]  ;
  input \a[23]  ;
  input \a[24]  ;
  input \a[25]  ;
  input \a[26]  ;
  input \a[27]  ;
  input \a[28]  ;
  input \a[29]  ;
  input \a[30]  ;
  input \a[31]  ;
  input \a[32]  ;
  input \a[33]  ;
  input \a[34]  ;
  input \a[35]  ;
  input \a[36]  ;
  input \a[37]  ;
  input \a[38]  ;
  input \a[39]  ;
  input \a[40]  ;
  input \a[41]  ;
  input \a[42]  ;
  input \a[43]  ;
  input \a[44]  ;
  input \a[45]  ;
  input \a[46]  ;
  input \a[47]  ;
  input \a[48]  ;
  input \a[49]  ;
  input \a[50]  ;
  input \a[51]  ;
  input \a[52]  ;
  input \a[53]  ;
  input \a[54]  ;
  input \a[55]  ;
  input \a[56]  ;
  input \a[57]  ;
  input \a[58]  ;
  input \a[59]  ;
  input \a[60]  ;
  input \a[61]  ;
  input \a[62]  ;
  input \a[63]  ;
  input \a[64]  ;
  input \a[65]  ;
  input \a[66]  ;
  input \a[67]  ;
  input \a[68]  ;
  input \a[69]  ;
  input \a[70]  ;
  input \a[71]  ;
  input \a[72]  ;
  input \a[73]  ;
  input \a[74]  ;
  input \a[75]  ;
  input \a[76]  ;
  input \a[77]  ;
  input \a[78]  ;
  input \a[79]  ;
  input \a[80]  ;
  input \a[81]  ;
  input \a[82]  ;
  input \a[83]  ;
  input \a[84]  ;
  input \a[85]  ;
  input \a[86]  ;
  input \a[87]  ;
  input \a[88]  ;
  input \a[89]  ;
  input \a[90]  ;
  input \a[91]  ;
  input \a[92]  ;
  input \a[93]  ;
  input \a[94]  ;
  input \a[95]  ;
  input \a[96]  ;
  input \a[97]  ;
  input \a[98]  ;
  input \a[99]  ;
  input \a[100]  ;
  input \a[101]  ;
  input \a[102]  ;
  input \a[103]  ;
  input \a[104]  ;
  input \a[105]  ;
  input \a[106]  ;
  input \a[107]  ;
  input \a[108]  ;
  input \a[109]  ;
  input \a[110]  ;
  input \a[111]  ;
  input \a[112]  ;
  input \a[113]  ;
  input \a[114]  ;
  input \a[115]  ;
  input \a[116]  ;
  input \a[117]  ;
  input \a[118]  ;
  input \a[119]  ;
  input \a[120]  ;
  input \a[121]  ;
  input \a[122]  ;
  input \a[123]  ;
  input \a[124]  ;
  input \a[125]  ;
  input \a[126]  ;
  input \a[127]  ;
  input \shift[0]  ;
  input \shift[1]  ;
  input \shift[2]  ;
  input \shift[3]  ;
  input \shift[4]  ;
  input \shift[5]  ;
  input \shift[6]  ;
  output \result[0]  ;
  output \result[1]  ;
  output \result[2]  ;
  output \result[3]  ;
  output \result[4]  ;
  output \result[5]  ;
  output \result[6]  ;
  output \result[7]  ;
  output \result[8]  ;
  output \result[9]  ;
  output \result[10]  ;
  output \result[11]  ;
  output \result[12]  ;
  output \result[13]  ;
  output \result[14]  ;
  output \result[15]  ;
  output \result[16]  ;
  output \result[17]  ;
  output \result[18]  ;
  output \result[19]  ;
  output \result[20]  ;
  output \result[21]  ;
  output \result[22]  ;
  output \result[23]  ;
  output \result[24]  ;
  output \result[25]  ;
  output \result[26]  ;
  output \result[27]  ;
  output \result[28]  ;
  output \result[29]  ;
  output \result[30]  ;
  output \result[31]  ;
  output \result[32]  ;
  output \result[33]  ;
  output \result[34]  ;
  output \result[35]  ;
  output \result[36]  ;
  output \result[37]  ;
  output \result[38]  ;
  output \result[39]  ;
  output \result[40]  ;
  output \result[41]  ;
  output \result[42]  ;
  output \result[43]  ;
  output \result[44]  ;
  output \result[45]  ;
  output \result[46]  ;
  output \result[47]  ;
  output \result[48]  ;
  output \result[49]  ;
  output \result[50]  ;
  output \result[51]  ;
  output \result[52]  ;
  output \result[53]  ;
  output \result[54]  ;
  output \result[55]  ;
  output \result[56]  ;
  output \result[57]  ;
  output \result[58]  ;
  output \result[59]  ;
  output \result[60]  ;
  output \result[61]  ;
  output \result[62]  ;
  output \result[63]  ;
  output \result[64]  ;
  output \result[65]  ;
  output \result[66]  ;
  output \result[67]  ;
  output \result[68]  ;
  output \result[69]  ;
  output \result[70]  ;
  output \result[71]  ;
  output \result[72]  ;
  output \result[73]  ;
  output \result[74]  ;
  output \result[75]  ;
  output \result[76]  ;
  output \result[77]  ;
  output \result[78]  ;
  output \result[79]  ;
  output \result[80]  ;
  output \result[81]  ;
  output \result[82]  ;
  output \result[83]  ;
  output \result[84]  ;
  output \result[85]  ;
  output \result[86]  ;
  output \result[87]  ;
  output \result[88]  ;
  output \result[89]  ;
  output \result[90]  ;
  output \result[91]  ;
  output \result[92]  ;
  output \result[93]  ;
  output \result[94]  ;
  output \result[95]  ;
  output \result[96]  ;
  output \result[97]  ;
  output \result[98]  ;
  output \result[99]  ;
  output \result[100]  ;
  output \result[101]  ;
  output \result[102]  ;
  output \result[103]  ;
  output \result[104]  ;
  output \result[105]  ;
  output \result[106]  ;
  output \result[107]  ;
  output \result[108]  ;
  output \result[109]  ;
  output \result[110]  ;
  output \result[111]  ;
  output \result[112]  ;
  output \result[113]  ;
  output \result[114]  ;
  output \result[115]  ;
  output \result[116]  ;
  output \result[117]  ;
  output \result[118]  ;
  output \result[119]  ;
  output \result[120]  ;
  output \result[121]  ;
  output \result[122]  ;
  output \result[123]  ;
  output \result[124]  ;
  output \result[125]  ;
  output \result[126]  ;
  output \result[127]  ;
  wire n136 , n137 , n138 , n139 , n140 , n141 , n142 , n143 , n144 , n145 , n146 , n147 , n148 , n149 , n150 , n151 , n152 , n153 , n154 , n155 , n156 , n157 , n158 , n159 , n160 , n161 , n162 , n163 , n164 , n165 , n166 , n167 , n168 , n169 , n170 , n171 , n172 , n173 , n174 , n175 , n176 , n177 , n178 , n179 , n180 , n181 , n182 , n183 , n184 , n185 , n186 , n187 , n188 , n189 , n190 , n191 , n192 , n193 , n194 , n195 , n196 , n197 , n198 , n199 , n200 , n201 , n202 , n203 , n204 , n205 , n206 , n207 , n208 , n209 , n210 , n211 , n212 , n213 , n214 , n215 , n216 , n217 , n218 , n219 , n220 , n221 , n222 , n223 , n224 , n225 , n226 , n227 , n228 , n229 , n230 , n231 , n232 , n233 , n234 , n235 , n236 , n237 , n238 , n239 , n240 , n241 , n242 , n243 , n244 , n245 , n246 , n247 , n248 , n249 , n250 , n251 , n252 , n253 , n254 , n255 , n256 , n257 , n258 , n259 , n260 , n261 , n262 , n263 , n264 , n265 , n266 , n267 , n268 , n269 , n270 , n271 , n272 , n273 , n274 , n275 , n276 , n277 , n278 , n279 , n280 , n281 , n282 , n283 , n284 , n285 , n286 , n287 , n288 , n289 , n290 , n291 , n292 , n293 , n294 , n295 , n296 , n297 , n298 , n299 , n300 , n301 , n302 , n303 , n304 , n305 , n306 , n307 , n308 , n309 , n310 , n311 , n312 , n313 , n314 , n315 , n316 , n317 , n318 , n319 , n320 , n321 , n322 , n323 , n324 , n325 , n326 , n327 , n328 , n329 , n330 , n331 , n332 , n333 , n334 , n335 , n336 , n337 , n338 , n339 , n340 , n341 , n342 , n343 , n344 , n345 , n346 , n347 , n348 , n349 , n350 , n351 , n352 , n353 , n354 , n355 , n356 , n357 , n358 , n359 , n360 , n361 , n362 , n363 , n364 , n365 , n366 , n367 , n368 , n369 , n370 , n371 , n372 , n373 , n374 , n375 , n376 , n377 , n378 , n379 , n380 , n381 , n382 , n383 , n384 , n385 , n386 , n387 , n388 , n389 , n390 , n391 , n392 , n393 , n394 , n395 , n396 , n397 , n398 , n399 , n400 , n401 , n402 , n403 , n404 , n405 , n406 , n407 , n408 , n409 , n410 , n411 , n412 , n413 , n414 , n415 , n416 , n417 , n418 , n419 , n420 , n421 , n422 , n423 , n424 , n425 , n426 , n427 , n428 , n429 , n430 , n431 , n432 , n433 , n434 , n435 , n436 , n437 , n438 , n439 , n440 , n441 , n442 , n443 , n444 , n445 , n446 , n447 , n448 , n449 , n450 , n451 , n452 , n453 , n454 , n455 , n456 , n457 , n458 , n459 , n460 , n461 , n462 , n463 , n464 , n465 , n466 , n467 , n468 , n469 , n470 , n471 , n472 , n473 , n474 , n475 , n476 , n477 , n478 , n479 , n480 , n481 , n482 , n483 , n484 , n485 , n486 , n487 , n488 , n489 , n490 , n491 , n492 , n493 , n494 , n495 , n496 , n497 , n498 , n499 , n500 , n501 , n502 , n503 , n504 , n505 , n506 , n507 , n508 , n509 , n510 , n511 , n512 , n513 , n514 , n515 , n516 , n517 , n518 , n519 , n520 , n521 , n522 , n523 , n524 , n525 , n526 , n527 , n528 , n529 , n530 , n531 , n532 , n533 , n534 , n535 , n536 , n537 , n538 , n539 , n540 , n541 , n542 , n543 , n544 , n545 , n546 , n547 , n548 , n549 , n550 , n551 , n552 , n553 , n554 , n555 , n556 , n557 , n558 , n559 , n560 , n561 , n562 , n563 , n564 , n565 , n566 , n567 , n568 , n569 , n570 , n571 , n572 , n573 , n574 , n575 , n576 , n577 , n578 , n579 , n580 , n581 , n582 , n583 , n584 , n585 , n586 , n587 , n588 , n589 , n590 , n591 , n592 , n593 , n594 , n595 , n596 , n597 , n598 , n599 , n600 , n601 , n602 , n603 , n604 , n605 , n606 , n607 , n608 , n609 , n610 , n611 , n612 , n613 , n614 , n615 , n616 , n617 , n618 , n619 , n620 , n621 , n622 , n623 , n624 , n625 , n626 , n627 , n628 , n629 , n630 , n631 , n632 , n633 , n634 , n635 , n636 , n637 , n638 , n639 , n640 , n641 , n642 , n643 , n644 , n645 , n646 , n647 , n648 , n649 , n650 , n651 , n652 , n653 , n654 , n655 , n656 , n657 , n658 , n659 , n660 , n661 , n662 , n663 , n664 , n665 , n666 , n667 , n668 , n669 , n670 , n671 , n672 , n673 , n674 , n675 , n676 , n677 , n678 , n679 , n680 , n681 , n682 , n683 , n684 , n685 , n686 , n687 , n688 , n689 , n690 , n691 , n692 , n693 , n694 , n695 , n696 , n697 , n698 , n699 , n700 , n701 , n702 , n703 , n704 , n705 , n706 , n707 , n708 , n709 , n710 , n711 , n712 , n713 , n714 , n715 , n716 , n717 , n718 , n719 , n720 , n721 , n722 , n723 , n724 , n725 , n726 , n727 , n728 , n729 , n730 , n731 , n732 , n733 , n734 , n735 , n736 , n737 , n738 , n739 , n740 , n741 , n742 , n743 , n744 , n745 , n746 , n747 , n748 , n749 , n750 , n751 , n752 , n753 , n754 , n755 , n756 , n757 , n758 , n759 , n760 , n761 , n762 , n763 , n764 , n765 , n766 , n767 , n768 , n769 , n770 , n771 , n772 , n773 , n774 , n775 , n776 , n777 , n778 , n779 , n780 , n781 , n782 , n783 , n784 , n785 , n786 , n787 , n788 , n789 , n790 , n791 , n792 , n793 , n794 , n795 , n796 , n797 , n798 , n799 , n800 , n801 , n802 , n803 , n804 , n805 , n806 , n807 , n808 , n809 , n810 , n811 , n812 , n813 , n814 , n815 , n816 , n817 , n818 , n819 , n820 , n821 , n822 , n823 , n824 , n825 , n826 , n827 , n828 , n829 , n830 , n831 , n832 , n833 , n834 , n835 , n836 , n837 , n838 , n839 , n840 , n841 , n842 , n843 , n844 , n845 , n846 , n847 , n848 , n849 , n850 , n851 , n852 , n853 , n854 , n855 , n856 , n857 , n858 , n859 , n860 , n861 , n862 , n863 , n864 , n865 , n866 , n867 , n868 , n869 , n870 , n871 , n872 , n873 , n874 , n875 , n876 , n877 , n878 , n879 , n880 , n881 , n882 , n883 , n884 , n885 , n886 , n887 , n888 , n889 , n890 , n891 , n892 , n893 , n894 , n895 , n896 , n897 , n898 , n899 , n900 , n901 , n902 , n903 , n904 , n905 , n906 , n907 , n908 , n909 , n910 , n911 , n912 , n913 , n914 , n915 , n916 , n917 , n918 , n919 , n920 , n921 , n922 , n923 , n924 , n925 , n926 , n927 , n928 , n929 , n930 , n931 , n932 , n933 , n934 , n935 , n936 , n937 , n938 , n939 , n940 , n941 , n942 , n943 , n944 , n945 , n946 , n947 , n948 , n949 , n950 , n951 , n952 , n953 , n954 , n955 , n956 , n957 , n958 , n959 , n960 , n961 , n962 , n963 , n964 , n965 , n966 , n967 , n968 , n969 , n970 , n971 , n972 , n973 , n974 , n975 , n976 , n977 , n978 , n979 , n980 , n981 , n982 , n983 , n984 , n985 , n986 , n987 , n988 , n989 , n990 , n991 , n992 , n993 , n994 , n995 , n996 , n997 , n998 , n999 , n1000 , n1001 , n1002 , n1003 , n1004 , n1005 , n1006 , n1007 , n1008 , n1009 , n1010 , n1011 , n1012 , n1013 , n1014 , n1015 , n1016 , n1017 , n1018 , n1019 , n1020 , n1021 , n1022 , n1023 , n1024 , n1025 , n1026 , n1027 , n1028 , n1029 , n1030 , n1031 , n1032 , n1033 , n1034 , n1035 , n1036 , n1037 , n1038 , n1039 , n1040 , n1041 , n1042 , n1043 , n1044 , n1045 , n1046 , n1047 , n1048 , n1049 , n1050 , n1051 , n1052 , n1053 , n1054 , n1055 , n1056 , n1057 , n1058 , n1059 , n1060 , n1061 , n1062 , n1063 , n1064 , n1065 , n1066 , n1067 , n1068 , n1069 , n1070 , n1071 , n1072 , n1073 , n1074 , n1075 , n1076 , n1077 , n1078 , n1079 , n1080 , n1081 , n1082 , n1083 , n1084 , n1085 , n1086 , n1087 , n1088 , n1089 , n1090 , n1091 , n1092 , n1093 , n1094 , n1095 , n1096 , n1097 , n1098 , n1099 , n1100 , n1101 , n1102 , n1103 , n1104 , n1105 , n1106 , n1107 , n1108 , n1109 , n1110 , n1111 , n1112 , n1113 , n1114 , n1115 , n1116 , n1117 , n1118 , n1119 , n1120 , n1121 , n1122 , n1123 , n1124 , n1125 , n1126 , n1127 , n1128 , n1129 , n1130 , n1131 , n1132 , n1133 , n1134 , n1135 , n1136 , n1137 , n1138 , n1139 , n1140 , n1141 , n1142 , n1143 , n1144 , n1145 , n1146 , n1147 , n1148 , n1149 , n1150 , n1151 , n1152 , n1153 , n1154 , n1155 , n1156 , n1157 , n1158 , n1159 , n1160 , n1161 , n1162 , n1163 , n1164 , n1165 , n1166 , n1167 , n1168 , n1169 , n1170 , n1171 , n1172 , n1173 , n1174 , n1175 , n1176 , n1177 , n1178 , n1179 , n1180 , n1181 , n1182 , n1183 , n1184 , n1185 , n1186 , n1187 , n1188 , n1189 , n1190 , n1191 , n1192 , n1193 , n1194 , n1195 , n1196 , n1197 , n1198 , n1199 , n1200 , n1201 , n1202 , n1203 , n1204 , n1205 , n1206 , n1207 , n1208 , n1209 , n1210 , n1211 , n1212 , n1213 , n1214 , n1215 , n1216 , n1217 , n1218 , n1219 , n1220 , n1221 , n1222 , n1223 , n1224 , n1225 , n1226 , n1227 , n1228 , n1229 , n1230 , n1231 , n1232 , n1233 , n1234 , n1235 , n1236 , n1237 , n1238 , n1239 , n1240 , n1241 , n1242 , n1243 , n1244 , n1245 , n1246 , n1247 , n1248 , n1249 , n1250 , n1251 , n1252 , n1253 , n1254 , n1255 , n1256 , n1257 , n1258 , n1259 , n1260 , n1261 , n1262 , n1263 , n1264 , n1265 , n1266 , n1267 , n1268 , n1269 , n1270 , n1271 , n1272 , n1273 , n1274 , n1275 , n1276 , n1277 , n1278 , n1279 , n1280 , n1281 , n1282 , n1283 , n1284 , n1285 , n1286 , n1287 , n1288 , n1289 , n1290 , n1291 , n1292 , n1293 , n1294 , n1295 , n1296 , n1297 , n1298 , n1299 , n1300 , n1301 , n1302 , n1303 , n1304 , n1305 , n1306 , n1307 , n1308 , n1309 , n1310 , n1311 , n1312 , n1313 , n1314 , n1315 , n1316 , n1317 , n1318 , n1319 , n1320 , n1321 , n1322 , n1323 , n1324 , n1325 , n1326 , n1327 , n1328 , n1329 , n1330 , n1331 , n1332 , n1333 , n1334 , n1335 , n1336 , n1337 , n1338 , n1339 , n1340 , n1341 , n1342 , n1343 , n1344 , n1345 , n1346 , n1347 , n1348 , n1349 , n1350 , n1351 , n1352 , n1353 , n1354 , n1355 , n1356 , n1357 , n1358 , n1359 , n1360 , n1361 , n1362 , n1363 , n1364 , n1365 , n1366 , n1367 , n1368 , n1369 , n1370 , n1371 , n1372 , n1373 , n1374 , n1375 , n1376 , n1377 , n1378 , n1379 , n1380 , n1381 , n1382 , n1383 , n1384 , n1385 , n1386 , n1387 , n1388 , n1389 , n1390 , n1391 , n1392 , n1393 , n1394 , n1395 , n1396 , n1397 , n1398 , n1399 , n1400 , n1401 , n1402 , n1403 , n1404 , n1405 , n1406 , n1407 , n1408 , n1409 , n1410 , n1411 , n1412 , n1413 , n1414 , n1415 , n1416 , n1417 , n1418 , n1419 , n1420 , n1421 , n1422 , n1423 , n1424 , n1425 , n1426 , n1427 , n1428 , n1429 , n1430 , n1431 , n1432 , n1433 , n1434 , n1435 , n1436 , n1437 , n1438 , n1439 , n1440 , n1441 , n1442 , n1443 , n1444 , n1445 , n1446 , n1447 , n1448 , n1449 , n1450 , n1451 , n1452 , n1453 , n1454 , n1455 , n1456 , n1457 , n1458 , n1459 , n1460 , n1461 , n1462 , n1463 , n1464 , n1465 , n1466 , n1467 , n1468 , n1469 , n1470 , n1471 , n1472 , n1473 , n1474 , n1475 , n1476 , n1477 , n1478 , n1479 , n1480 , n1481 , n1482 , n1483 , n1484 , n1485 , n1486 , n1487 , n1488 , n1489 , n1490 , n1491 , n1492 , n1493 , n1494 , n1495 , n1496 , n1497 , n1498 , n1499 , n1500 , n1501 , n1502 , n1503 , n1504 , n1505 , n1506 , n1507 , n1508 , n1509 , n1510 , n1511 , n1512 , n1513 , n1514 , n1515 , n1516 , n1517 , n1518 , n1519 , n1520 , n1521 , n1522 , n1523 , n1524 , n1525 , n1526 , n1527 , n1528 , n1529 , n1530 , n1531 , n1532 , n1533 , n1534 , n1535 , n1536 , n1537 , n1538 , n1539 , n1540 , n1541 , n1542 , n1543 , n1544 , n1545 , n1546 , n1547 , n1548 , n1549 , n1550 , n1551 , n1552 , n1553 , n1554 , n1555 , n1556 , n1557 , n1558 , n1559 , n1560 , n1561 , n1562 , n1563 , n1564 , n1565 , n1566 , n1567 , n1568 , n1569 , n1570 , n1571 , n1572 , n1573 , n1574 , n1575 , n1576 , n1577 , n1578 , n1579 , n1580 , n1581 , n1582 , n1583 , n1584 , n1585 , n1586 , n1587 , n1588 , n1589 , n1590 , n1591 , n1592 , n1593 , n1594 , n1595 , n1596 , n1597 , n1598 , n1599 , n1600 , n1601 , n1602 , n1603 , n1604 , n1605 , n1606 , n1607 , n1608 , n1609 , n1610 , n1611 , n1612 , n1613 , n1614 , n1615 , n1616 , n1617 , n1618 , n1619 , n1620 , n1621 , n1622 , n1623 , n1624 , n1625 , n1626 , n1627 , n1628 , n1629 , n1630 , n1631 , n1632 , n1633 , n1634 , n1635 , n1636 , n1637 , n1638 , n1639 , n1640 , n1641 , n1642 , n1643 , n1644 , n1645 , n1646 , n1647 , n1648 , n1649 , n1650 , n1651 , n1652 , n1653 , n1654 , n1655 , n1656 , n1657 , n1658 , n1659 , n1660 , n1661 , n1662 , n1663 , n1664 , n1665 , n1666 , n1667 , n1668 , n1669 , n1670 , n1671 , n1672 , n1673 , n1674 , n1675 , n1676 , n1677 , n1678 , n1679 , n1680 , n1681 , n1682 , n1683 , n1684 , n1685 , n1686 , n1687 , n1688 , n1689 , n1690 , n1691 , n1692 , n1693 , n1694 , n1695 , n1696 , n1697 , n1698 , n1699 , n1700 , n1701 , n1702 , n1703 , n1704 , n1705 , n1706 , n1707 , n1708 , n1709 , n1710 , n1711 , n1712 , n1713 , n1714 , n1715 , n1716 , n1717 , n1718 , n1719 , n1720 , n1721 , n1722 , n1723 , n1724 , n1725 , n1726 , n1727 , n1728 , n1729 , n1730 , n1731 , n1732 , n1733 , n1734 , n1735 , n1736 , n1737 , n1738 , n1739 , n1740 , n1741 , n1742 , n1743 , n1744 , n1745 , n1746 , n1747 , n1748 , n1749 , n1750 , n1751 , n1752 , n1753 , n1754 , n1755 , n1756 , n1757 , n1758 , n1759 , n1760 , n1761 , n1762 , n1763 , n1764 , n1765 , n1766 , n1767 , n1768 , n1769 , n1770 , n1771 , n1772 , n1773 , n1774 , n1775 , n1776 , n1777 , n1778 , n1779 , n1780 , n1781 , n1782 , n1783 , n1784 , n1785 , n1786 , n1787 , n1788 , n1789 , n1790 , n1791 , n1792 , n1793 , n1794 , n1795 , n1796 , n1797 , n1798 , n1799 , n1800 , n1801 , n1802 , n1803 , n1804 , n1805 , n1806 , n1807 , n1808 , n1809 , n1810 , n1811 , n1812 , n1813 , n1814 , n1815 , n1816 , n1817 , n1818 , n1819 , n1820 , n1821 , n1822 , n1823 , n1824 , n1825 , n1826 , n1827 , n1828 , n1829 , n1830 , n1831 , n1832 , n1833 , n1834 , n1835 , n1836 , n1837 , n1838 , n1839 , n1840 , n1841 , n1842 , n1843 , n1844 , n1845 , n1846 , n1847 , n1848 , n1849 , n1850 , n1851 , n1852 , n1853 , n1854 , n1855 , n1856 , n1857 , n1858 , n1859 , n1860 , n1861 , n1862 , n1863 , n1864 , n1865 , n1866 , n1867 , n1868 , n1869 , n1870 , n1871 , n1872 , n1873 , n1874 , n1875 , n1876 , n1877 , n1878 , n1879 , n1880 , n1881 , n1882 , n1883 , n1884 , n1885 , n1886 , n1887 , n1888 , n1889 , n1890 , n1891 , n1892 , n1893 , n1894 , n1895 , n1896 , n1897 , n1898 , n1899 , n1900 , n1901 , n1902 , n1903 , n1904 , n1905 , n1906 , n1907 , n1908 , n1909 , n1910 , n1911 , n1912 , n1913 , n1914 , n1915 , n1916 , n1917 , n1918 , n1919 , n1920 , n1921 , n1922 , n1923 , n1924 , n1925 , n1926 , n1927 , n1928 , n1929 , n1930 , n1931 , n1932 , n1933 , n1934 , n1935 , n1936 , n1937 , n1938 , n1939 , n1940 , n1941 , n1942 , n1943 , n1944 , n1945 , n1946 , n1947 , n1948 , n1949 , n1950 , n1951 , n1952 , n1953 , n1954 , n1955 , n1956 , n1957 , n1958 , n1959 , n1960 , n1961 , n1962 , n1963 , n1964 , n1965 , n1966 , n1967 , n1968 , n1969 , n1970 , n1971 , n1972 , n1973 , n1974 , n1975 , n1976 , n1977 , n1978 , n1979 , n1980 , n1981 , n1982 , n1983 , n1984 , n1985 , n1986 , n1987 , n1988 , n1989 , n1990 , n1991 , n1992 , n1993 , n1994 , n1995 , n1996 , n1997 , n1998 , n1999 , n2000 , n2001 , n2002 , n2003 , n2004 , n2005 , n2006 , n2007 , n2008 , n2009 , n2010 , n2011 , n2012 , n2013 , n2014 , n2015 , n2016 , n2017 , n2018 , n2019 , n2020 , n2021 , n2022 , n2023 , n2024 , n2025 , n2026 , n2027 , n2028 , n2029 , n2030 , n2031 , n2032 , n2033 , n2034 , n2035 , n2036 , n2037 , n2038 , n2039 , n2040 , n2041 , n2042 , n2043 , n2044 , n2045 , n2046 , n2047 , n2048 , n2049 , n2050 , n2051 , n2052 , n2053 , n2054 , n2055 , n2056 , n2057 , n2058 , n2059 , n2060 , n2061 , n2062 , n2063 , n2064 , n2065 , n2066 , n2067 , n2068 , n2069 , n2070 , n2071 , n2072 , n2073 , n2074 , n2075 , n2076 , n2077 , n2078 , n2079 , n2080 , n2081 , n2082 , n2083 , n2084 , n2085 , n2086 , n2087 , n2088 , n2089 , n2090 , n2091 , n2092 , n2093 , n2094 , n2095 , n2096 , n2097 , n2098 , n2099 , n2100 , n2101 , n2102 , n2103 , n2104 , n2105 , n2106 , n2107 , n2108 , n2109 , n2110 , n2111 , n2112 , n2113 , n2114 , n2115 , n2116 , n2117 , n2118 , n2119 , n2120 , n2121 , n2122 , n2123 , n2124 , n2125 , n2126 , n2127 , n2128 , n2129 , n2130 , n2131 , n2132 , n2133 , n2134 , n2135 , n2136 , n2137 , n2138 , n2139 , n2140 , n2141 , n2142 , n2143 , n2144 , n2145 , n2146 , n2147 , n2148 , n2149 , n2150 , n2151 , n2152 , n2153 , n2154 , n2155 , n2156 , n2157 , n2158 , n2159 , n2160 , n2161 , n2162 , n2163 , n2164 , n2165 , n2166 , n2167 , n2168 , n2169 , n2170 , n2171 , n2172 , n2173 , n2174 , n2175 , n2176 , n2177 , n2178 , n2179 , n2180 , n2181 , n2182 , n2183 , n2184 , n2185 , n2186 , n2187 , n2188 , n2189 , n2190 , n2191 , n2192 , n2193 , n2194 , n2195 , n2196 , n2197 , n2198 , n2199 , n2200 , n2201 , n2202 , n2203 , n2204 , n2205 , n2206 , n2207 , n2208 , n2209 , n2210 , n2211 , n2212 , n2213 , n2214 , n2215 , n2216 , n2217 , n2218 , n2219 , n2220 , n2221 , n2222 , n2223 , n2224 , n2225 , n2226 , n2227 , n2228 , n2229 , n2230 , n2231 , n2232 , n2233 , n2234 , n2235 , n2236 , n2237 , n2238 , n2239 , n2240 , n2241 , n2242 , n2243 , n2244 , n2245 , n2246 , n2247 , n2248 , n2249 , n2250 , n2251 , n2252 , n2253 , n2254 , n2255 , n2256 , n2257 , n2258 , n2259 , n2260 , n2261 , n2262 , n2263 , n2264 , n2265 , n2266 , n2267 , n2268 , n2269 , n2270 , n2271 , n2272 , n2273 , n2274 , n2275 , n2276 , n2277 , n2278 , n2279 , n2280 , n2281 , n2282 , n2283 , n2284 , n2285 , n2286 , n2287 , n2288 , n2289 , n2290 , n2291 , n2292 , n2293 , n2294 , n2295 , n2296 , n2297 , n2298 , n2299 , n2300 , n2301 , n2302 , n2303 , n2304 , n2305 , n2306 , n2307 , n2308 , n2309 , n2310 , n2311 , n2312 , n2313 , n2314 , n2315 , n2316 , n2317 , n2318 , n2319 , n2320 , n2321 , n2322 , n2323 , n2324 , n2325 , n2326 , n2327 , n2328 , n2329 , n2330 , n2331 , n2332 , n2333 , n2334 , n2335 , n2336 , n2337 , n2338 , n2339 , n2340 , n2341 , n2342 , n2343 , n2344 , n2345 , n2346 , n2347 , n2348 , n2349 , n2350 , n2351 , n2352 , n2353 , n2354 , n2355 , n2356 , n2357 , n2358 , n2359 , n2360 , n2361 , n2362 , n2363 , n2364 , n2365 , n2366 , n2367 , n2368 , n2369 , n2370 , n2371 , n2372 , n2373 , n2374 , n2375 , n2376 , n2377 , n2378 , n2379 , n2380 , n2381 , n2382 , n2383 , n2384 , n2385 , n2386 , n2387 , n2388 , n2389 , n2390 , n2391 , n2392 , n2393 , n2394 , n2395 , n2396 , n2397 , n2398 , n2399 , n2400 , n2401 , n2402 , n2403 , n2404 , n2405 , n2406 , n2407 , n2408 , n2409 , n2410 , n2411 , n2412 , n2413 , n2414 , n2415 , n2416 , n2417 , n2418 , n2419 , n2420 , n2421 , n2422 , n2423 , n2424 , n2425 , n2426 , n2427 , n2428 , n2429 , n2430 , n2431 , n2432 , n2433 , n2434 , n2435 , n2436 , n2437 , n2438 , n2439 , n2440 , n2441 , n2442 , n2443 , n2444 , n2445 , n2446 , n2447 , n2448 , n2449 , n2450 , n2451 , n2452 , n2453 , n2454 , n2455 , n2456 , n2457 , n2458 , n2459 , n2460 , n2461 , n2462 , n2463 , n2464 , n2465 , n2466 , n2467 , n2468 , n2469 , n2470 , n2471 , n2472 , n2473 , n2474 , n2475 , n2476 , n2477 , n2478 , n2479 , n2480 , n2481 , n2482 , n2483 , n2484 , n2485 , n2486 , n2487 , n2488 , n2489 , n2490 , n2491 , n2492 , n2493 , n2494 , n2495 , n2496 , n2497 , n2498 , n2499 , n2500 , n2501 , n2502 , n2503 , n2504 , n2505 , n2506 , n2507 , n2508 , n2509 , n2510 , n2511 , n2512 , n2513 , n2514 , n2515 , n2516 , n2517 , n2518 , n2519 , n2520 , n2521 , n2522 , n2523 , n2524 , n2525 , n2526 , n2527 , n2528 , n2529 , n2530 , n2531 , n2532 , n2533 , n2534 , n2535 , n2536 , n2537 , n2538 , n2539 , n2540 , n2541 , n2542 , n2543 , n2544 , n2545 , n2546 , n2547 , n2548 , n2549 , n2550 , n2551 , n2552 , n2553 , n2554 , n2555 , n2556 , n2557 , n2558 , n2559 , n2560 , n2561 , n2562 , n2563 , n2564 , n2565 , n2566 , n2567 , n2568 , n2569 , n2570 , n2571 , n2572 , n2573 , n2574 , n2575 , n2576 , n2577 , n2578 , n2579 , n2580 , n2581 , n2582 , n2583 , n2584 , n2585 , n2586 , n2587 , n2588 , n2589 , n2590 , n2591 , n2592 , n2593 , n2594 , n2595 , n2596 , n2597 , n2598 , n2599 , n2600 , n2601 , n2602 , n2603 , n2604 , n2605 , n2606 , n2607 , n2608 , n2609 , n2610 , n2611 , n2612 , n2613 , n2614 , n2615 , n2616 , n2617 , n2618 , n2619 , n2620 , n2621 , n2622 , n2623 , n2624 , n2625 , n2626 , n2627 , n2628 , n2629 , n2630 , n2631 , n2632 , n2633 , n2634 , n2635 , n2636 , n2637 , n2638 , n2639 , n2640 , n2641 , n2642 , n2643 , n2644 , n2645 , n2646 , n2647 , n2648 , n2649 , n2650 , n2651 , n2652 , n2653 , n2654 , n2655 , n2656 , n2657 , n2658 , n2659 , n2660 , n2661 , n2662 , n2663 , n2664 , n2665 , n2666 , n2667 , n2668 , n2669 , n2670 , n2671 , n2672 , n2673 , n2674 , n2675 , n2676 , n2677 , n2678 , n2679 , n2680 , n2681 , n2682 , n2683 , n2684 , n2685 , n2686 , n2687 , n2688 , n2689 , n2690 , n2691 , n2692 , n2693 , n2694 , n2695 , n2696 , n2697 , n2698 , n2699 , n2700 , n2701 , n2702 , n2703 , n2704 , n2705 , n2706 , n2707 , n2708 , n2709 , n2710 , n2711 , n2712 , n2713 , n2714 , n2715 , n2716 , n2717 , n2718 , n2719 , n2720 , n2721 , n2722 , n2723 , n2724 , n2725 , n2726 , n2727 , n2728 , n2729 , n2730 , n2731 , n2732 , n2733 , n2734 , n2735 , n2736 , n2737 , n2738 , n2739 , n2740 , n2741 , n2742 , n2743 , n2744 , n2745 , n2746 , n2747 , n2748 , n2749 , n2750 , n2751 , n2752 , n2753 , n2754 , n2755 , n2756 , n2757 , n2758 , n2759 , n2760 , n2761 , n2762 , n2763 , n2764 , n2765 , n2766 , n2767 , n2768 , n2769 , n2770 , n2771 , n2772 , n2773 , n2774 , n2775 , n2776 , n2777 , n2778 , n2779 , n2780 , n2781 , n2782 , n2783 , n2784 , n2785 , n2786 , n2787 , n2788 , n2789 , n2790 , n2791 , n2792 , n2793 , n2794 , n2795 , n2796 , n2797 , n2798 , n2799 , n2800 , n2801 , n2802 , n2803 , n2804 , n2805 , n2806 , n2807 , n2808 , n2809 , n2810 , n2811 , n2812 , n2813 , n2814 , n2815 , n2816 , n2817 , n2818 , n2819 , n2820 , n2821 , n2822 , n2823 , n2824 , n2825 , n2826 , n2827 , n2828 , n2829 , n2830 , n2831 , n2832 , n2833 , n2834 , n2835 , n2836 , n2837 , n2838 , n2839 , n2840 , n2841 , n2842 , n2843 , n2844 , n2845 , n2846 , n2847 , n2848 , n2849 , n2850 , n2851 , n2852 , n2853 , n2854 , n2855 , n2856 , n2857 , n2858 , n2859 , n2860 , n2861 , n2862 , n2863 , n2864 , n2865 , n2866 , n2867 , n2868 , n2869 , n2870 , n2871 , n2872 , n2873 , n2874 , n2875 , n2876 , n2877 , n2878 , n2879 , n2880 , n2881 , n2882 , n2883 , n2884 , n2885 , n2886 , n2887 , n2888 , n2889 , n2890 , n2891 , n2892 , n2893 , n2894 , n2895 , n2896 , n2897 , n2898 , n2899 , n2900 , n2901 , n2902 , n2903 , n2904 , n2905 , n2906 , n2907 , n2908 , n2909 , n2910 , n2911 , n2912 , n2913 , n2914 , n2915 , n2916 , n2917 , n2918 , n2919 , n2920 , n2921 , n2922 , n2923 , n2924 , n2925 , n2926 , n2927 , n2928 , n2929 , n2930 , n2931 , n2932 , n2933 , n2934 , n2935 , n2936 , n2937 , n2938 , n2939 , n2940 , n2941 , n2942 , n2943 , n2944 , n2945 , n2946 , n2947 , n2948 , n2949 , n2950 , n2951 , n2952 , n2953 , n2954 , n2955 , n2956 , n2957 , n2958 , n2959 , n2960 , n2961 , n2962 , n2963 , n2964 , n2965 , n2966 , n2967 , n2968 , n2969 , n2970 , n2971 , n2972 , n2973 , n2974 , n2975 , n2976 , n2977 , n2978 , n2979 , n2980 , n2981 , n2982 , n2983 , n2984 , n2985 , n2986 , n2987 , n2988 , n2989 , n2990 , n2991 , n2992 , n2993 , n2994 , n2995 , n2996 , n2997 , n2998 , n2999 , n3000 , n3001 , n3002 , n3003 , n3004 , n3005 , n3006 , n3007 , n3008 , n3009 , n3010 , n3011 , n3012 , n3013 , n3014 , n3015 , n3016 , n3017 , n3018 , n3019 , n3020 , n3021 , n3022 , n3023 , n3024 , n3025 , n3026 , n3027 , n3028 , n3029 , n3030 , n3031 , n3032 , n3033 , n3034 , n3035 , n3036 , n3037 , n3038 , n3039 , n3040 , n3041 , n3042 , n3043 , n3044 , n3045 , n3046 , n3047 , n3048 , n3049 , n3050 , n3051 , n3052 , n3053 , n3054 , n3055 , n3056 , n3057 , n3058 , n3059 , n3060 , n3061 , n3062 , n3063 , n3064 , n3065 , n3066 , n3067 , n3068 , n3069 , n3070 , n3071 , n3072 , n3073 , n3074 , n3075 , n3076 , n3077 , n3078 , n3079 , n3080 , n3081 , n3082 , n3083 , n3084 , n3085 , n3086 , n3087 , n3088 , n3089 , n3090 , n3091 , n3092 , n3093 , n3094 , n3095 , n3096 , n3097 , n3098 , n3099 , n3100 , n3101 , n3102 , n3103 , n3104 , n3105 , n3106 , n3107 , n3108 , n3109 , n3110 , n3111 , n3112 , n3113 , n3114 , n3115 , n3116 , n3117 , n3118 , n3119 , n3120 , n3121 , n3122 , n3123 , n3124 , n3125 , n3126 , n3127 , n3128 , n3129 , n3130 , n3131 , n3132 , n3133 , n3134 , n3135 , n3136 , n3137 , n3138 , n3139 , n3140 , n3141 , n3142 , n3143 , n3144 , n3145 , n3146 , n3147 , n3148 , n3149 , n3150 , n3151 , n3152 , n3153 , n3154 , n3155 , n3156 , n3157 , n3158 , n3159 , n3160 , n3161 , n3162 , n3163 , n3164 , n3165 , n3166 , n3167 , n3168 , n3169 , n3170 , n3171 , n3172 , n3173 , n3174 , n3175 , n3176 , n3177 , n3178 , n3179 , n3180 , n3181 , n3182 , n3183 , n3184 , n3185 , n3186 , n3187 , n3188 , n3189 , n3190 , n3191 , n3192 , n3193 , n3194 , n3195 , n3196 , n3197 , n3198 , n3199 , n3200 , n3201 , n3202 , n3203 , n3204 , n3205 , n3206 , n3207 , n3208 , n3209 , n3210 , n3211 , n3212 , n3213 , n3214 , n3215 , n3216 , n3217 , n3218 , n3219 , n3220 , n3221 , n3222 , n3223 , n3224 , n3225 , n3226 , n3227 , n3228 , n3229 , n3230 , n3231 , n3232 , n3233 , n3234 , n3235 , n3236 , n3237 , n3238 , n3239 , n3240 , n3241 , n3242 , n3243 , n3244 , n3245 , n3246 , n3247 , n3248 , n3249 , n3250 , n3251 , n3252 , n3253 , n3254 , n3255 , n3256 , n3257 , n3258 , n3259 , n3260 , n3261 , n3262 , n3263 , n3264 , n3265 , n3266 , n3267 , n3268 , n3269 , n3270 , n3271 , n3272 , n3273 , n3274 , n3275 , n3276 ;
  assign n136 = ~\shift[2]  & ~\shift[3]  ;
  assign n137 = \a[77]  & \shift[0]  ;
  assign n138 = \a[78]  & ~\shift[0]  ;
  assign n139 = ~n137 & ~n138 ;
  assign n140 = \shift[1]  & ~n139 ;
  assign n141 = \a[80]  & ~\shift[0]  ;
  assign n142 = \a[79]  & \shift[0]  ;
  assign n143 = ~n141 & ~n142 ;
  assign n144 = ~\shift[1]  & ~n143 ;
  assign n145 = ~n140 & ~n144 ;
  assign n146 = n136 & ~n145 ;
  assign n147 = \shift[2]  & ~\shift[3]  ;
  assign n148 = \a[73]  & \shift[0]  ;
  assign n149 = \a[74]  & ~\shift[0]  ;
  assign n150 = ~n148 & ~n149 ;
  assign n151 = \shift[1]  & ~n150 ;
  assign n152 = \a[76]  & ~\shift[0]  ;
  assign n153 = \a[75]  & \shift[0]  ;
  assign n154 = ~n152 & ~n153 ;
  assign n155 = ~\shift[1]  & ~n154 ;
  assign n156 = ~n151 & ~n155 ;
  assign n157 = n147 & ~n156 ;
  assign n180 = ~n146 & ~n157 ;
  assign n158 = \shift[2]  & \shift[3]  ;
  assign n159 = \a[65]  & \shift[0]  ;
  assign n160 = \a[66]  & ~\shift[0]  ;
  assign n161 = ~n159 & ~n160 ;
  assign n162 = \shift[1]  & ~n161 ;
  assign n163 = \a[68]  & ~\shift[0]  ;
  assign n164 = \a[67]  & \shift[0]  ;
  assign n165 = ~n163 & ~n164 ;
  assign n166 = ~\shift[1]  & ~n165 ;
  assign n167 = ~n162 & ~n166 ;
  assign n168 = n158 & ~n167 ;
  assign n169 = ~\shift[2]  & \shift[3]  ;
  assign n170 = \a[69]  & \shift[0]  ;
  assign n171 = \a[70]  & ~\shift[0]  ;
  assign n172 = ~n170 & ~n171 ;
  assign n173 = \shift[1]  & ~n172 ;
  assign n174 = \a[72]  & ~\shift[0]  ;
  assign n175 = \a[71]  & \shift[0]  ;
  assign n176 = ~n174 & ~n175 ;
  assign n177 = ~\shift[1]  & ~n176 ;
  assign n178 = ~n173 & ~n177 ;
  assign n179 = n169 & ~n178 ;
  assign n181 = ~n168 & ~n179 ;
  assign n182 = n180 & n181 ;
  assign n183 = \shift[4]  & \shift[5]  ;
  assign n184 = ~n182 & n183 ;
  assign n185 = \a[93]  & \shift[0]  ;
  assign n186 = \a[94]  & ~\shift[0]  ;
  assign n187 = ~n185 & ~n186 ;
  assign n188 = \shift[1]  & ~n187 ;
  assign n189 = \a[96]  & ~\shift[0]  ;
  assign n190 = \a[95]  & \shift[0]  ;
  assign n191 = ~n189 & ~n190 ;
  assign n192 = ~\shift[1]  & ~n191 ;
  assign n193 = ~n188 & ~n192 ;
  assign n194 = n136 & ~n193 ;
  assign n195 = \a[89]  & \shift[0]  ;
  assign n196 = \a[90]  & ~\shift[0]  ;
  assign n197 = ~n195 & ~n196 ;
  assign n198 = \shift[1]  & ~n197 ;
  assign n199 = \a[92]  & ~\shift[0]  ;
  assign n200 = \a[91]  & \shift[0]  ;
  assign n201 = ~n199 & ~n200 ;
  assign n202 = ~\shift[1]  & ~n201 ;
  assign n203 = ~n198 & ~n202 ;
  assign n204 = n147 & ~n203 ;
  assign n225 = ~n194 & ~n204 ;
  assign n205 = \a[81]  & \shift[0]  ;
  assign n206 = \a[82]  & ~\shift[0]  ;
  assign n207 = ~n205 & ~n206 ;
  assign n208 = \shift[1]  & ~n207 ;
  assign n209 = \a[84]  & ~\shift[0]  ;
  assign n210 = \a[83]  & \shift[0]  ;
  assign n211 = ~n209 & ~n210 ;
  assign n212 = ~\shift[1]  & ~n211 ;
  assign n213 = ~n208 & ~n212 ;
  assign n214 = n158 & ~n213 ;
  assign n215 = \a[85]  & \shift[0]  ;
  assign n216 = \a[86]  & ~\shift[0]  ;
  assign n217 = ~n215 & ~n216 ;
  assign n218 = \shift[1]  & ~n217 ;
  assign n219 = \a[88]  & ~\shift[0]  ;
  assign n220 = \a[87]  & \shift[0]  ;
  assign n221 = ~n219 & ~n220 ;
  assign n222 = ~\shift[1]  & ~n221 ;
  assign n223 = ~n218 & ~n222 ;
  assign n224 = n169 & ~n223 ;
  assign n226 = ~n214 & ~n224 ;
  assign n227 = n225 & n226 ;
  assign n228 = ~\shift[4]  & \shift[5]  ;
  assign n229 = ~n227 & n228 ;
  assign n320 = ~n184 & ~n229 ;
  assign n230 = \a[125]  & \shift[0]  ;
  assign n231 = \a[126]  & ~\shift[0]  ;
  assign n232 = ~n230 & ~n231 ;
  assign n233 = \shift[1]  & ~n232 ;
  assign n234 = \a[0]  & ~\shift[0]  ;
  assign n235 = \a[127]  & \shift[0]  ;
  assign n236 = ~n234 & ~n235 ;
  assign n237 = ~\shift[1]  & ~n236 ;
  assign n238 = ~n233 & ~n237 ;
  assign n239 = n136 & ~n238 ;
  assign n240 = \a[121]  & \shift[0]  ;
  assign n241 = \a[122]  & ~\shift[0]  ;
  assign n242 = ~n240 & ~n241 ;
  assign n243 = \shift[1]  & ~n242 ;
  assign n244 = \a[124]  & ~\shift[0]  ;
  assign n245 = \a[123]  & \shift[0]  ;
  assign n246 = ~n244 & ~n245 ;
  assign n247 = ~\shift[1]  & ~n246 ;
  assign n248 = ~n243 & ~n247 ;
  assign n249 = n147 & ~n248 ;
  assign n270 = ~n239 & ~n249 ;
  assign n250 = \a[113]  & \shift[0]  ;
  assign n251 = \a[114]  & ~\shift[0]  ;
  assign n252 = ~n250 & ~n251 ;
  assign n253 = \shift[1]  & ~n252 ;
  assign n254 = \a[116]  & ~\shift[0]  ;
  assign n255 = \a[115]  & \shift[0]  ;
  assign n256 = ~n254 & ~n255 ;
  assign n257 = ~\shift[1]  & ~n256 ;
  assign n258 = ~n253 & ~n257 ;
  assign n259 = n158 & ~n258 ;
  assign n260 = \a[117]  & \shift[0]  ;
  assign n261 = \a[118]  & ~\shift[0]  ;
  assign n262 = ~n260 & ~n261 ;
  assign n263 = \shift[1]  & ~n262 ;
  assign n264 = \a[120]  & ~\shift[0]  ;
  assign n265 = \a[119]  & \shift[0]  ;
  assign n266 = ~n264 & ~n265 ;
  assign n267 = ~\shift[1]  & ~n266 ;
  assign n268 = ~n263 & ~n267 ;
  assign n269 = n169 & ~n268 ;
  assign n271 = ~n259 & ~n269 ;
  assign n272 = n270 & n271 ;
  assign n273 = ~\shift[4]  & ~\shift[5]  ;
  assign n274 = ~n272 & n273 ;
  assign n275 = \a[109]  & \shift[0]  ;
  assign n276 = \a[110]  & ~\shift[0]  ;
  assign n277 = ~n275 & ~n276 ;
  assign n278 = \shift[1]  & ~n277 ;
  assign n279 = \a[112]  & ~\shift[0]  ;
  assign n280 = \a[111]  & \shift[0]  ;
  assign n281 = ~n279 & ~n280 ;
  assign n282 = ~\shift[1]  & ~n281 ;
  assign n283 = ~n278 & ~n282 ;
  assign n284 = n136 & ~n283 ;
  assign n285 = \a[105]  & \shift[0]  ;
  assign n286 = \a[106]  & ~\shift[0]  ;
  assign n287 = ~n285 & ~n286 ;
  assign n288 = \shift[1]  & ~n287 ;
  assign n289 = \a[108]  & ~\shift[0]  ;
  assign n290 = \a[107]  & \shift[0]  ;
  assign n291 = ~n289 & ~n290 ;
  assign n292 = ~\shift[1]  & ~n291 ;
  assign n293 = ~n288 & ~n292 ;
  assign n294 = n147 & ~n293 ;
  assign n315 = ~n284 & ~n294 ;
  assign n295 = \a[97]  & \shift[0]  ;
  assign n296 = \a[98]  & ~\shift[0]  ;
  assign n297 = ~n295 & ~n296 ;
  assign n298 = \shift[1]  & ~n297 ;
  assign n299 = \a[100]  & ~\shift[0]  ;
  assign n300 = \a[99]  & \shift[0]  ;
  assign n301 = ~n299 & ~n300 ;
  assign n302 = ~\shift[1]  & ~n301 ;
  assign n303 = ~n298 & ~n302 ;
  assign n304 = n158 & ~n303 ;
  assign n305 = \a[101]  & \shift[0]  ;
  assign n306 = \a[102]  & ~\shift[0]  ;
  assign n307 = ~n305 & ~n306 ;
  assign n308 = \shift[1]  & ~n307 ;
  assign n309 = \a[104]  & ~\shift[0]  ;
  assign n310 = \a[103]  & \shift[0]  ;
  assign n311 = ~n309 & ~n310 ;
  assign n312 = ~\shift[1]  & ~n311 ;
  assign n313 = ~n308 & ~n312 ;
  assign n314 = n169 & ~n313 ;
  assign n316 = ~n304 & ~n314 ;
  assign n317 = n315 & n316 ;
  assign n318 = \shift[4]  & ~\shift[5]  ;
  assign n319 = ~n317 & n318 ;
  assign n321 = ~n274 & ~n319 ;
  assign n322 = n320 & n321 ;
  assign n323 = ~\shift[6]  & ~n322 ;
  assign n324 = \a[13]  & \shift[0]  ;
  assign n325 = \a[14]  & ~\shift[0]  ;
  assign n326 = ~n324 & ~n325 ;
  assign n327 = \shift[1]  & ~n326 ;
  assign n328 = \a[16]  & ~\shift[0]  ;
  assign n329 = \a[15]  & \shift[0]  ;
  assign n330 = ~n328 & ~n329 ;
  assign n331 = ~\shift[1]  & ~n330 ;
  assign n332 = ~n327 & ~n331 ;
  assign n333 = n136 & ~n332 ;
  assign n334 = \a[9]  & \shift[0]  ;
  assign n335 = \a[10]  & ~\shift[0]  ;
  assign n336 = ~n334 & ~n335 ;
  assign n337 = \shift[1]  & ~n336 ;
  assign n338 = \a[12]  & ~\shift[0]  ;
  assign n339 = \a[11]  & \shift[0]  ;
  assign n340 = ~n338 & ~n339 ;
  assign n341 = ~\shift[1]  & ~n340 ;
  assign n342 = ~n337 & ~n341 ;
  assign n343 = n147 & ~n342 ;
  assign n364 = ~n333 & ~n343 ;
  assign n344 = \a[1]  & \shift[0]  ;
  assign n345 = \a[2]  & ~\shift[0]  ;
  assign n346 = ~n344 & ~n345 ;
  assign n347 = \shift[1]  & ~n346 ;
  assign n348 = \a[4]  & ~\shift[0]  ;
  assign n349 = \a[3]  & \shift[0]  ;
  assign n350 = ~n348 & ~n349 ;
  assign n351 = ~\shift[1]  & ~n350 ;
  assign n352 = ~n347 & ~n351 ;
  assign n353 = n158 & ~n352 ;
  assign n354 = \a[5]  & \shift[0]  ;
  assign n355 = \a[6]  & ~\shift[0]  ;
  assign n356 = ~n354 & ~n355 ;
  assign n357 = \shift[1]  & ~n356 ;
  assign n358 = \a[8]  & ~\shift[0]  ;
  assign n359 = \a[7]  & \shift[0]  ;
  assign n360 = ~n358 & ~n359 ;
  assign n361 = ~\shift[1]  & ~n360 ;
  assign n362 = ~n357 & ~n361 ;
  assign n363 = n169 & ~n362 ;
  assign n365 = ~n353 & ~n363 ;
  assign n366 = n364 & n365 ;
  assign n367 = n183 & ~n366 ;
  assign n368 = \a[29]  & \shift[0]  ;
  assign n369 = \a[30]  & ~\shift[0]  ;
  assign n370 = ~n368 & ~n369 ;
  assign n371 = \shift[1]  & ~n370 ;
  assign n372 = \a[32]  & ~\shift[0]  ;
  assign n373 = \a[31]  & \shift[0]  ;
  assign n374 = ~n372 & ~n373 ;
  assign n375 = ~\shift[1]  & ~n374 ;
  assign n376 = ~n371 & ~n375 ;
  assign n377 = n136 & ~n376 ;
  assign n378 = \a[25]  & \shift[0]  ;
  assign n379 = \a[26]  & ~\shift[0]  ;
  assign n380 = ~n378 & ~n379 ;
  assign n381 = \shift[1]  & ~n380 ;
  assign n382 = \a[28]  & ~\shift[0]  ;
  assign n383 = \a[27]  & \shift[0]  ;
  assign n384 = ~n382 & ~n383 ;
  assign n385 = ~\shift[1]  & ~n384 ;
  assign n386 = ~n381 & ~n385 ;
  assign n387 = n147 & ~n386 ;
  assign n408 = ~n377 & ~n387 ;
  assign n388 = \a[17]  & \shift[0]  ;
  assign n389 = \a[18]  & ~\shift[0]  ;
  assign n390 = ~n388 & ~n389 ;
  assign n391 = \shift[1]  & ~n390 ;
  assign n392 = \a[20]  & ~\shift[0]  ;
  assign n393 = \a[19]  & \shift[0]  ;
  assign n394 = ~n392 & ~n393 ;
  assign n395 = ~\shift[1]  & ~n394 ;
  assign n396 = ~n391 & ~n395 ;
  assign n397 = n158 & ~n396 ;
  assign n398 = \a[21]  & \shift[0]  ;
  assign n399 = \a[22]  & ~\shift[0]  ;
  assign n400 = ~n398 & ~n399 ;
  assign n401 = \shift[1]  & ~n400 ;
  assign n402 = \a[24]  & ~\shift[0]  ;
  assign n403 = \a[23]  & \shift[0]  ;
  assign n404 = ~n402 & ~n403 ;
  assign n405 = ~\shift[1]  & ~n404 ;
  assign n406 = ~n401 & ~n405 ;
  assign n407 = n169 & ~n406 ;
  assign n409 = ~n397 & ~n407 ;
  assign n410 = n408 & n409 ;
  assign n411 = n228 & ~n410 ;
  assign n502 = ~n367 & ~n411 ;
  assign n412 = \a[61]  & \shift[0]  ;
  assign n413 = \a[62]  & ~\shift[0]  ;
  assign n414 = ~n412 & ~n413 ;
  assign n415 = \shift[1]  & ~n414 ;
  assign n416 = \a[64]  & ~\shift[0]  ;
  assign n417 = \a[63]  & \shift[0]  ;
  assign n418 = ~n416 & ~n417 ;
  assign n419 = ~\shift[1]  & ~n418 ;
  assign n420 = ~n415 & ~n419 ;
  assign n421 = n136 & ~n420 ;
  assign n422 = \a[57]  & \shift[0]  ;
  assign n423 = \a[58]  & ~\shift[0]  ;
  assign n424 = ~n422 & ~n423 ;
  assign n425 = \shift[1]  & ~n424 ;
  assign n426 = \a[60]  & ~\shift[0]  ;
  assign n427 = \a[59]  & \shift[0]  ;
  assign n428 = ~n426 & ~n427 ;
  assign n429 = ~\shift[1]  & ~n428 ;
  assign n430 = ~n425 & ~n429 ;
  assign n431 = n147 & ~n430 ;
  assign n452 = ~n421 & ~n431 ;
  assign n432 = \a[49]  & \shift[0]  ;
  assign n433 = \a[50]  & ~\shift[0]  ;
  assign n434 = ~n432 & ~n433 ;
  assign n435 = \shift[1]  & ~n434 ;
  assign n436 = \a[52]  & ~\shift[0]  ;
  assign n437 = \a[51]  & \shift[0]  ;
  assign n438 = ~n436 & ~n437 ;
  assign n439 = ~\shift[1]  & ~n438 ;
  assign n440 = ~n435 & ~n439 ;
  assign n441 = n158 & ~n440 ;
  assign n442 = \a[53]  & \shift[0]  ;
  assign n443 = \a[54]  & ~\shift[0]  ;
  assign n444 = ~n442 & ~n443 ;
  assign n445 = \shift[1]  & ~n444 ;
  assign n446 = \a[56]  & ~\shift[0]  ;
  assign n447 = \a[55]  & \shift[0]  ;
  assign n448 = ~n446 & ~n447 ;
  assign n449 = ~\shift[1]  & ~n448 ;
  assign n450 = ~n445 & ~n449 ;
  assign n451 = n169 & ~n450 ;
  assign n453 = ~n441 & ~n451 ;
  assign n454 = n452 & n453 ;
  assign n455 = n273 & ~n454 ;
  assign n456 = \a[45]  & \shift[0]  ;
  assign n457 = \a[46]  & ~\shift[0]  ;
  assign n458 = ~n456 & ~n457 ;
  assign n459 = \shift[1]  & ~n458 ;
  assign n460 = \a[48]  & ~\shift[0]  ;
  assign n461 = \a[47]  & \shift[0]  ;
  assign n462 = ~n460 & ~n461 ;
  assign n463 = ~\shift[1]  & ~n462 ;
  assign n464 = ~n459 & ~n463 ;
  assign n465 = n136 & ~n464 ;
  assign n466 = \a[41]  & \shift[0]  ;
  assign n467 = \a[42]  & ~\shift[0]  ;
  assign n468 = ~n466 & ~n467 ;
  assign n469 = \shift[1]  & ~n468 ;
  assign n470 = \a[44]  & ~\shift[0]  ;
  assign n471 = \a[43]  & \shift[0]  ;
  assign n472 = ~n470 & ~n471 ;
  assign n473 = ~\shift[1]  & ~n472 ;
  assign n474 = ~n469 & ~n473 ;
  assign n475 = n147 & ~n474 ;
  assign n498 = ~n465 & ~n475 ;
  assign n476 = \a[33]  & \shift[0]  ;
  assign n477 = \a[34]  & ~\shift[0]  ;
  assign n478 = ~n476 & ~n477 ;
  assign n479 = \shift[1]  & ~n478 ;
  assign n480 = \a[36]  & ~\shift[0]  ;
  assign n481 = \a[35]  & \shift[0]  ;
  assign n482 = ~n480 & ~n481 ;
  assign n483 = ~\shift[1]  & ~n482 ;
  assign n484 = ~n479 & ~n483 ;
  assign n485 = n158 & ~n484 ;
  assign n486 = \a[40]  & ~\shift[0]  ;
  assign n487 = ~\shift[1]  & ~n486 ;
  assign n488 = \a[37]  & \shift[0]  ;
  assign n489 = \shift[1]  & ~n488 ;
  assign n490 = ~n487 & ~n489 ;
  assign n491 = \a[38]  & ~\shift[0]  ;
  assign n492 = \shift[1]  & n491 ;
  assign n493 = \a[39]  & \shift[0]  ;
  assign n494 = ~\shift[1]  & n493 ;
  assign n495 = ~n492 & ~n494 ;
  assign n496 = ~n490 & n495 ;
  assign n497 = n169 & ~n496 ;
  assign n499 = ~n485 & ~n497 ;
  assign n500 = n498 & n499 ;
  assign n501 = n318 & ~n500 ;
  assign n503 = ~n455 & ~n501 ;
  assign n504 = n502 & n503 ;
  assign n505 = \shift[6]  & ~n504 ;
  assign n506 = ~n323 & ~n505 ;
  assign n507 = \a[81]  & ~\shift[0]  ;
  assign n508 = ~\shift[1]  & ~n507 ;
  assign n509 = \a[78]  & \shift[0]  ;
  assign n510 = \shift[1]  & ~n509 ;
  assign n511 = ~n508 & ~n510 ;
  assign n512 = \a[79]  & ~\shift[0]  ;
  assign n513 = \shift[1]  & n512 ;
  assign n514 = \a[80]  & \shift[0]  ;
  assign n515 = ~\shift[1]  & n514 ;
  assign n516 = ~n513 & ~n515 ;
  assign n517 = ~n511 & n516 ;
  assign n518 = n136 & ~n517 ;
  assign n519 = \a[77]  & ~\shift[0]  ;
  assign n520 = ~\shift[1]  & ~n519 ;
  assign n521 = \a[74]  & \shift[0]  ;
  assign n522 = \shift[1]  & ~n521 ;
  assign n523 = ~n520 & ~n522 ;
  assign n524 = \a[75]  & ~\shift[0]  ;
  assign n525 = \shift[1]  & n524 ;
  assign n526 = \a[76]  & \shift[0]  ;
  assign n527 = ~\shift[1]  & n526 ;
  assign n528 = ~n525 & ~n527 ;
  assign n529 = ~n523 & n528 ;
  assign n530 = n147 & ~n529 ;
  assign n555 = ~n518 & ~n530 ;
  assign n531 = \a[69]  & ~\shift[0]  ;
  assign n532 = ~\shift[1]  & ~n531 ;
  assign n533 = \a[66]  & \shift[0]  ;
  assign n534 = \shift[1]  & ~n533 ;
  assign n535 = ~n532 & ~n534 ;
  assign n536 = \a[67]  & ~\shift[0]  ;
  assign n537 = \shift[1]  & n536 ;
  assign n538 = \a[68]  & \shift[0]  ;
  assign n539 = ~\shift[1]  & n538 ;
  assign n540 = ~n537 & ~n539 ;
  assign n541 = ~n535 & n540 ;
  assign n542 = n158 & ~n541 ;
  assign n543 = \a[73]  & ~\shift[0]  ;
  assign n544 = ~\shift[1]  & ~n543 ;
  assign n545 = \a[70]  & \shift[0]  ;
  assign n546 = \shift[1]  & ~n545 ;
  assign n547 = ~n544 & ~n546 ;
  assign n548 = \a[71]  & ~\shift[0]  ;
  assign n549 = \shift[1]  & n548 ;
  assign n550 = \a[72]  & \shift[0]  ;
  assign n551 = ~\shift[1]  & n550 ;
  assign n552 = ~n549 & ~n551 ;
  assign n553 = ~n547 & n552 ;
  assign n554 = n169 & ~n553 ;
  assign n556 = ~n542 & ~n554 ;
  assign n557 = n555 & n556 ;
  assign n558 = n183 & ~n557 ;
  assign n559 = \a[97]  & ~\shift[0]  ;
  assign n560 = ~\shift[1]  & ~n559 ;
  assign n561 = \a[94]  & \shift[0]  ;
  assign n562 = \shift[1]  & ~n561 ;
  assign n563 = ~n560 & ~n562 ;
  assign n564 = \a[95]  & ~\shift[0]  ;
  assign n565 = \shift[1]  & n564 ;
  assign n566 = \a[96]  & \shift[0]  ;
  assign n567 = ~\shift[1]  & n566 ;
  assign n568 = ~n565 & ~n567 ;
  assign n569 = ~n563 & n568 ;
  assign n570 = n136 & ~n569 ;
  assign n571 = \a[93]  & ~\shift[0]  ;
  assign n572 = ~\shift[1]  & ~n571 ;
  assign n573 = \a[90]  & \shift[0]  ;
  assign n574 = \shift[1]  & ~n573 ;
  assign n575 = ~n572 & ~n574 ;
  assign n576 = \a[91]  & ~\shift[0]  ;
  assign n577 = \shift[1]  & n576 ;
  assign n578 = \a[92]  & \shift[0]  ;
  assign n579 = ~\shift[1]  & n578 ;
  assign n580 = ~n577 & ~n579 ;
  assign n581 = ~n575 & n580 ;
  assign n582 = n147 & ~n581 ;
  assign n607 = ~n570 & ~n582 ;
  assign n583 = \a[85]  & ~\shift[0]  ;
  assign n584 = ~\shift[1]  & ~n583 ;
  assign n585 = \a[82]  & \shift[0]  ;
  assign n586 = \shift[1]  & ~n585 ;
  assign n587 = ~n584 & ~n586 ;
  assign n588 = \a[83]  & ~\shift[0]  ;
  assign n589 = \shift[1]  & n588 ;
  assign n590 = \a[84]  & \shift[0]  ;
  assign n591 = ~\shift[1]  & n590 ;
  assign n592 = ~n589 & ~n591 ;
  assign n593 = ~n587 & n592 ;
  assign n594 = n158 & ~n593 ;
  assign n595 = \a[89]  & ~\shift[0]  ;
  assign n596 = ~\shift[1]  & ~n595 ;
  assign n597 = \a[86]  & \shift[0]  ;
  assign n598 = \shift[1]  & ~n597 ;
  assign n599 = ~n596 & ~n598 ;
  assign n600 = \a[87]  & ~\shift[0]  ;
  assign n601 = \shift[1]  & n600 ;
  assign n602 = \a[88]  & \shift[0]  ;
  assign n603 = ~\shift[1]  & n602 ;
  assign n604 = ~n601 & ~n603 ;
  assign n605 = ~n599 & n604 ;
  assign n606 = n169 & ~n605 ;
  assign n608 = ~n594 & ~n606 ;
  assign n609 = n607 & n608 ;
  assign n610 = n228 & ~n609 ;
  assign n715 = ~n558 & ~n610 ;
  assign n611 = \a[1]  & ~\shift[0]  ;
  assign n612 = ~\shift[1]  & ~n611 ;
  assign n613 = \a[126]  & \shift[0]  ;
  assign n614 = \shift[1]  & ~n613 ;
  assign n615 = ~n612 & ~n614 ;
  assign n616 = \a[127]  & ~\shift[0]  ;
  assign n617 = \shift[1]  & n616 ;
  assign n618 = \a[0]  & \shift[0]  ;
  assign n619 = ~\shift[1]  & n618 ;
  assign n620 = ~n617 & ~n619 ;
  assign n621 = ~n615 & n620 ;
  assign n622 = n136 & ~n621 ;
  assign n623 = \a[125]  & ~\shift[0]  ;
  assign n624 = ~\shift[1]  & ~n623 ;
  assign n625 = \a[122]  & \shift[0]  ;
  assign n626 = \shift[1]  & ~n625 ;
  assign n627 = ~n624 & ~n626 ;
  assign n628 = \a[123]  & ~\shift[0]  ;
  assign n629 = \shift[1]  & n628 ;
  assign n630 = \a[124]  & \shift[0]  ;
  assign n631 = ~\shift[1]  & n630 ;
  assign n632 = ~n629 & ~n631 ;
  assign n633 = ~n627 & n632 ;
  assign n634 = n147 & ~n633 ;
  assign n659 = ~n622 & ~n634 ;
  assign n635 = \a[117]  & ~\shift[0]  ;
  assign n636 = ~\shift[1]  & ~n635 ;
  assign n637 = \a[114]  & \shift[0]  ;
  assign n638 = \shift[1]  & ~n637 ;
  assign n639 = ~n636 & ~n638 ;
  assign n640 = \a[115]  & ~\shift[0]  ;
  assign n641 = \shift[1]  & n640 ;
  assign n642 = \a[116]  & \shift[0]  ;
  assign n643 = ~\shift[1]  & n642 ;
  assign n644 = ~n641 & ~n643 ;
  assign n645 = ~n639 & n644 ;
  assign n646 = n158 & ~n645 ;
  assign n647 = \a[121]  & ~\shift[0]  ;
  assign n648 = ~\shift[1]  & ~n647 ;
  assign n649 = \a[118]  & \shift[0]  ;
  assign n650 = \shift[1]  & ~n649 ;
  assign n651 = ~n648 & ~n650 ;
  assign n652 = \a[119]  & ~\shift[0]  ;
  assign n653 = \shift[1]  & n652 ;
  assign n654 = \a[120]  & \shift[0]  ;
  assign n655 = ~\shift[1]  & n654 ;
  assign n656 = ~n653 & ~n655 ;
  assign n657 = ~n651 & n656 ;
  assign n658 = n169 & ~n657 ;
  assign n660 = ~n646 & ~n658 ;
  assign n661 = n659 & n660 ;
  assign n662 = n273 & ~n661 ;
  assign n663 = \a[113]  & ~\shift[0]  ;
  assign n664 = ~\shift[1]  & ~n663 ;
  assign n665 = \a[110]  & \shift[0]  ;
  assign n666 = \shift[1]  & ~n665 ;
  assign n667 = ~n664 & ~n666 ;
  assign n668 = \a[111]  & ~\shift[0]  ;
  assign n669 = \shift[1]  & n668 ;
  assign n670 = \a[112]  & \shift[0]  ;
  assign n671 = ~\shift[1]  & n670 ;
  assign n672 = ~n669 & ~n671 ;
  assign n673 = ~n667 & n672 ;
  assign n674 = n136 & ~n673 ;
  assign n675 = \a[109]  & ~\shift[0]  ;
  assign n676 = ~\shift[1]  & ~n675 ;
  assign n677 = \a[106]  & \shift[0]  ;
  assign n678 = \shift[1]  & ~n677 ;
  assign n679 = ~n676 & ~n678 ;
  assign n680 = \a[107]  & ~\shift[0]  ;
  assign n681 = \shift[1]  & n680 ;
  assign n682 = \a[108]  & \shift[0]  ;
  assign n683 = ~\shift[1]  & n682 ;
  assign n684 = ~n681 & ~n683 ;
  assign n685 = ~n679 & n684 ;
  assign n686 = n147 & ~n685 ;
  assign n711 = ~n674 & ~n686 ;
  assign n687 = \a[101]  & ~\shift[0]  ;
  assign n688 = ~\shift[1]  & ~n687 ;
  assign n689 = \a[98]  & \shift[0]  ;
  assign n690 = \shift[1]  & ~n689 ;
  assign n691 = ~n688 & ~n690 ;
  assign n692 = \a[99]  & ~\shift[0]  ;
  assign n693 = \shift[1]  & n692 ;
  assign n694 = \a[100]  & \shift[0]  ;
  assign n695 = ~\shift[1]  & n694 ;
  assign n696 = ~n693 & ~n695 ;
  assign n697 = ~n691 & n696 ;
  assign n698 = n158 & ~n697 ;
  assign n699 = \a[105]  & ~\shift[0]  ;
  assign n700 = ~\shift[1]  & ~n699 ;
  assign n701 = \a[102]  & \shift[0]  ;
  assign n702 = \shift[1]  & ~n701 ;
  assign n703 = ~n700 & ~n702 ;
  assign n704 = \a[103]  & ~\shift[0]  ;
  assign n705 = \shift[1]  & n704 ;
  assign n706 = \a[104]  & \shift[0]  ;
  assign n707 = ~\shift[1]  & n706 ;
  assign n708 = ~n705 & ~n707 ;
  assign n709 = ~n703 & n708 ;
  assign n710 = n169 & ~n709 ;
  assign n712 = ~n698 & ~n710 ;
  assign n713 = n711 & n712 ;
  assign n714 = n318 & ~n713 ;
  assign n716 = ~n662 & ~n714 ;
  assign n717 = n715 & n716 ;
  assign n718 = ~\shift[6]  & ~n717 ;
  assign n719 = \a[65]  & ~\shift[0]  ;
  assign n720 = ~\shift[1]  & ~n719 ;
  assign n721 = \a[62]  & \shift[0]  ;
  assign n722 = \shift[1]  & ~n721 ;
  assign n723 = ~n720 & ~n722 ;
  assign n724 = \a[63]  & ~\shift[0]  ;
  assign n725 = \shift[1]  & n724 ;
  assign n726 = \a[64]  & \shift[0]  ;
  assign n727 = ~\shift[1]  & n726 ;
  assign n728 = ~n725 & ~n727 ;
  assign n729 = ~n723 & n728 ;
  assign n730 = n136 & ~n729 ;
  assign n731 = \a[61]  & ~\shift[0]  ;
  assign n732 = ~\shift[1]  & ~n731 ;
  assign n733 = \a[58]  & \shift[0]  ;
  assign n734 = \shift[1]  & ~n733 ;
  assign n735 = ~n732 & ~n734 ;
  assign n736 = \a[59]  & ~\shift[0]  ;
  assign n737 = \shift[1]  & n736 ;
  assign n738 = \a[60]  & \shift[0]  ;
  assign n739 = ~\shift[1]  & n738 ;
  assign n740 = ~n737 & ~n739 ;
  assign n741 = ~n735 & n740 ;
  assign n742 = n147 & ~n741 ;
  assign n767 = ~n730 & ~n742 ;
  assign n743 = \a[53]  & ~\shift[0]  ;
  assign n744 = ~\shift[1]  & ~n743 ;
  assign n745 = \a[50]  & \shift[0]  ;
  assign n746 = \shift[1]  & ~n745 ;
  assign n747 = ~n744 & ~n746 ;
  assign n748 = \a[51]  & ~\shift[0]  ;
  assign n749 = \shift[1]  & n748 ;
  assign n750 = \a[52]  & \shift[0]  ;
  assign n751 = ~\shift[1]  & n750 ;
  assign n752 = ~n749 & ~n751 ;
  assign n753 = ~n747 & n752 ;
  assign n754 = n158 & ~n753 ;
  assign n755 = \a[57]  & ~\shift[0]  ;
  assign n756 = ~\shift[1]  & ~n755 ;
  assign n757 = \a[54]  & \shift[0]  ;
  assign n758 = \shift[1]  & ~n757 ;
  assign n759 = ~n756 & ~n758 ;
  assign n760 = \a[55]  & ~\shift[0]  ;
  assign n761 = \shift[1]  & n760 ;
  assign n762 = \a[56]  & \shift[0]  ;
  assign n763 = ~\shift[1]  & n762 ;
  assign n764 = ~n761 & ~n763 ;
  assign n765 = ~n759 & n764 ;
  assign n766 = n169 & ~n765 ;
  assign n768 = ~n754 & ~n766 ;
  assign n769 = n767 & n768 ;
  assign n770 = n273 & ~n769 ;
  assign n771 = \a[17]  & ~\shift[0]  ;
  assign n772 = ~\shift[1]  & ~n771 ;
  assign n773 = \a[14]  & \shift[0]  ;
  assign n774 = \shift[1]  & ~n773 ;
  assign n775 = ~n772 & ~n774 ;
  assign n776 = \a[15]  & ~\shift[0]  ;
  assign n777 = \shift[1]  & n776 ;
  assign n778 = \a[16]  & \shift[0]  ;
  assign n779 = ~\shift[1]  & n778 ;
  assign n780 = ~n777 & ~n779 ;
  assign n781 = ~n775 & n780 ;
  assign n782 = n136 & ~n781 ;
  assign n783 = \a[13]  & ~\shift[0]  ;
  assign n784 = ~\shift[1]  & ~n783 ;
  assign n785 = \a[10]  & \shift[0]  ;
  assign n786 = \shift[1]  & ~n785 ;
  assign n787 = ~n784 & ~n786 ;
  assign n788 = \a[11]  & ~\shift[0]  ;
  assign n789 = \shift[1]  & n788 ;
  assign n790 = \a[12]  & \shift[0]  ;
  assign n791 = ~\shift[1]  & n790 ;
  assign n792 = ~n789 & ~n791 ;
  assign n793 = ~n787 & n792 ;
  assign n794 = n147 & ~n793 ;
  assign n819 = ~n782 & ~n794 ;
  assign n795 = \a[5]  & ~\shift[0]  ;
  assign n796 = ~\shift[1]  & ~n795 ;
  assign n797 = \a[2]  & \shift[0]  ;
  assign n798 = \shift[1]  & ~n797 ;
  assign n799 = ~n796 & ~n798 ;
  assign n800 = \a[3]  & ~\shift[0]  ;
  assign n801 = \shift[1]  & n800 ;
  assign n802 = \a[4]  & \shift[0]  ;
  assign n803 = ~\shift[1]  & n802 ;
  assign n804 = ~n801 & ~n803 ;
  assign n805 = ~n799 & n804 ;
  assign n806 = n158 & ~n805 ;
  assign n807 = \a[9]  & ~\shift[0]  ;
  assign n808 = ~\shift[1]  & ~n807 ;
  assign n809 = \a[6]  & \shift[0]  ;
  assign n810 = \shift[1]  & ~n809 ;
  assign n811 = ~n808 & ~n810 ;
  assign n812 = \a[7]  & ~\shift[0]  ;
  assign n813 = \shift[1]  & n812 ;
  assign n814 = \a[8]  & \shift[0]  ;
  assign n815 = ~\shift[1]  & n814 ;
  assign n816 = ~n813 & ~n815 ;
  assign n817 = ~n811 & n816 ;
  assign n818 = n169 & ~n817 ;
  assign n820 = ~n806 & ~n818 ;
  assign n821 = n819 & n820 ;
  assign n822 = n183 & ~n821 ;
  assign n923 = ~n770 & ~n822 ;
  assign n823 = \a[49]  & ~\shift[0]  ;
  assign n824 = ~\shift[1]  & ~n823 ;
  assign n825 = \a[46]  & \shift[0]  ;
  assign n826 = \shift[1]  & ~n825 ;
  assign n827 = ~n824 & ~n826 ;
  assign n828 = \a[47]  & ~\shift[0]  ;
  assign n829 = \shift[1]  & n828 ;
  assign n830 = \a[48]  & \shift[0]  ;
  assign n831 = ~\shift[1]  & n830 ;
  assign n832 = ~n829 & ~n831 ;
  assign n833 = ~n827 & n832 ;
  assign n834 = n136 & ~n833 ;
  assign n835 = \a[42]  & \shift[0]  ;
  assign n836 = \a[43]  & ~\shift[0]  ;
  assign n837 = ~n835 & ~n836 ;
  assign n838 = \shift[1]  & ~n837 ;
  assign n839 = \a[45]  & ~\shift[0]  ;
  assign n840 = \a[44]  & \shift[0]  ;
  assign n841 = ~n839 & ~n840 ;
  assign n842 = ~\shift[1]  & ~n841 ;
  assign n843 = ~n838 & ~n842 ;
  assign n844 = n147 & ~n843 ;
  assign n867 = ~n834 & ~n844 ;
  assign n845 = \a[37]  & ~\shift[0]  ;
  assign n846 = ~\shift[1]  & ~n845 ;
  assign n847 = \a[34]  & \shift[0]  ;
  assign n848 = \shift[1]  & ~n847 ;
  assign n849 = ~n846 & ~n848 ;
  assign n850 = \a[35]  & ~\shift[0]  ;
  assign n851 = \shift[1]  & n850 ;
  assign n852 = \a[36]  & \shift[0]  ;
  assign n853 = ~\shift[1]  & n852 ;
  assign n854 = ~n851 & ~n853 ;
  assign n855 = ~n849 & n854 ;
  assign n856 = n158 & ~n855 ;
  assign n857 = \a[41]  & ~\shift[0]  ;
  assign n858 = \a[40]  & \shift[0]  ;
  assign n859 = ~n857 & ~n858 ;
  assign n860 = ~\shift[1]  & ~n859 ;
  assign n861 = \a[39]  & ~\shift[0]  ;
  assign n862 = \a[38]  & \shift[0]  ;
  assign n863 = ~n861 & ~n862 ;
  assign n864 = \shift[1]  & ~n863 ;
  assign n865 = ~n860 & ~n864 ;
  assign n866 = n169 & ~n865 ;
  assign n868 = ~n856 & ~n866 ;
  assign n869 = n867 & n868 ;
  assign n870 = n318 & ~n869 ;
  assign n871 = \a[33]  & ~\shift[0]  ;
  assign n872 = ~\shift[1]  & ~n871 ;
  assign n873 = \a[30]  & \shift[0]  ;
  assign n874 = \shift[1]  & ~n873 ;
  assign n875 = ~n872 & ~n874 ;
  assign n876 = \a[31]  & ~\shift[0]  ;
  assign n877 = \shift[1]  & n876 ;
  assign n878 = \a[32]  & \shift[0]  ;
  assign n879 = ~\shift[1]  & n878 ;
  assign n880 = ~n877 & ~n879 ;
  assign n881 = ~n875 & n880 ;
  assign n882 = n136 & ~n881 ;
  assign n883 = \a[29]  & ~\shift[0]  ;
  assign n884 = ~\shift[1]  & ~n883 ;
  assign n885 = \a[26]  & \shift[0]  ;
  assign n886 = \shift[1]  & ~n885 ;
  assign n887 = ~n884 & ~n886 ;
  assign n888 = \a[27]  & ~\shift[0]  ;
  assign n889 = \shift[1]  & n888 ;
  assign n890 = \a[28]  & \shift[0]  ;
  assign n891 = ~\shift[1]  & n890 ;
  assign n892 = ~n889 & ~n891 ;
  assign n893 = ~n887 & n892 ;
  assign n894 = n147 & ~n893 ;
  assign n919 = ~n882 & ~n894 ;
  assign n895 = \a[21]  & ~\shift[0]  ;
  assign n896 = ~\shift[1]  & ~n895 ;
  assign n897 = \a[18]  & \shift[0]  ;
  assign n898 = \shift[1]  & ~n897 ;
  assign n899 = ~n896 & ~n898 ;
  assign n900 = \a[19]  & ~\shift[0]  ;
  assign n901 = \shift[1]  & n900 ;
  assign n902 = \a[20]  & \shift[0]  ;
  assign n903 = ~\shift[1]  & n902 ;
  assign n904 = ~n901 & ~n903 ;
  assign n905 = ~n899 & n904 ;
  assign n906 = n158 & ~n905 ;
  assign n907 = \a[25]  & ~\shift[0]  ;
  assign n908 = ~\shift[1]  & ~n907 ;
  assign n909 = \a[22]  & \shift[0]  ;
  assign n910 = \shift[1]  & ~n909 ;
  assign n911 = ~n908 & ~n910 ;
  assign n912 = \a[23]  & ~\shift[0]  ;
  assign n913 = \shift[1]  & n912 ;
  assign n914 = \a[24]  & \shift[0]  ;
  assign n915 = ~\shift[1]  & n914 ;
  assign n916 = ~n913 & ~n915 ;
  assign n917 = ~n911 & n916 ;
  assign n918 = n169 & ~n917 ;
  assign n920 = ~n906 & ~n918 ;
  assign n921 = n919 & n920 ;
  assign n922 = n228 & ~n921 ;
  assign n924 = ~n870 & ~n922 ;
  assign n925 = n923 & n924 ;
  assign n926 = \shift[6]  & ~n925 ;
  assign n927 = ~n718 & ~n926 ;
  assign n928 = \shift[1]  & ~n143 ;
  assign n929 = ~\shift[1]  & ~n207 ;
  assign n930 = ~n928 & ~n929 ;
  assign n931 = n136 & ~n930 ;
  assign n932 = \shift[1]  & ~n154 ;
  assign n933 = ~\shift[1]  & ~n139 ;
  assign n934 = ~n932 & ~n933 ;
  assign n935 = n147 & ~n934 ;
  assign n944 = ~n931 & ~n935 ;
  assign n936 = \shift[1]  & ~n165 ;
  assign n937 = ~\shift[1]  & ~n172 ;
  assign n938 = ~n936 & ~n937 ;
  assign n939 = n158 & ~n938 ;
  assign n940 = \shift[1]  & ~n176 ;
  assign n941 = ~\shift[1]  & ~n150 ;
  assign n942 = ~n940 & ~n941 ;
  assign n943 = n169 & ~n942 ;
  assign n945 = ~n939 & ~n943 ;
  assign n946 = n944 & n945 ;
  assign n947 = n183 & ~n946 ;
  assign n948 = \shift[1]  & ~n191 ;
  assign n949 = ~\shift[1]  & ~n297 ;
  assign n950 = ~n948 & ~n949 ;
  assign n951 = n136 & ~n950 ;
  assign n952 = \shift[1]  & ~n201 ;
  assign n953 = ~\shift[1]  & ~n187 ;
  assign n954 = ~n952 & ~n953 ;
  assign n955 = n147 & ~n954 ;
  assign n964 = ~n951 & ~n955 ;
  assign n956 = \shift[1]  & ~n211 ;
  assign n957 = ~\shift[1]  & ~n217 ;
  assign n958 = ~n956 & ~n957 ;
  assign n959 = n158 & ~n958 ;
  assign n960 = \shift[1]  & ~n221 ;
  assign n961 = ~\shift[1]  & ~n197 ;
  assign n962 = ~n960 & ~n961 ;
  assign n963 = n169 & ~n962 ;
  assign n965 = ~n959 & ~n963 ;
  assign n966 = n964 & n965 ;
  assign n967 = n228 & ~n966 ;
  assign n1008 = ~n947 & ~n967 ;
  assign n968 = \shift[1]  & ~n236 ;
  assign n969 = ~\shift[1]  & ~n346 ;
  assign n970 = ~n968 & ~n969 ;
  assign n971 = n136 & ~n970 ;
  assign n972 = \shift[1]  & ~n246 ;
  assign n973 = ~\shift[1]  & ~n232 ;
  assign n974 = ~n972 & ~n973 ;
  assign n975 = n147 & ~n974 ;
  assign n984 = ~n971 & ~n975 ;
  assign n976 = \shift[1]  & ~n256 ;
  assign n977 = ~\shift[1]  & ~n262 ;
  assign n978 = ~n976 & ~n977 ;
  assign n979 = n158 & ~n978 ;
  assign n980 = \shift[1]  & ~n266 ;
  assign n981 = ~\shift[1]  & ~n242 ;
  assign n982 = ~n980 & ~n981 ;
  assign n983 = n169 & ~n982 ;
  assign n985 = ~n979 & ~n983 ;
  assign n986 = n984 & n985 ;
  assign n987 = n273 & ~n986 ;
  assign n988 = \shift[1]  & ~n281 ;
  assign n989 = ~\shift[1]  & ~n252 ;
  assign n990 = ~n988 & ~n989 ;
  assign n991 = n136 & ~n990 ;
  assign n992 = \shift[1]  & ~n291 ;
  assign n993 = ~\shift[1]  & ~n277 ;
  assign n994 = ~n992 & ~n993 ;
  assign n995 = n147 & ~n994 ;
  assign n1004 = ~n991 & ~n995 ;
  assign n996 = \shift[1]  & ~n301 ;
  assign n997 = ~\shift[1]  & ~n307 ;
  assign n998 = ~n996 & ~n997 ;
  assign n999 = n158 & ~n998 ;
  assign n1000 = \shift[1]  & ~n311 ;
  assign n1001 = ~\shift[1]  & ~n287 ;
  assign n1002 = ~n1000 & ~n1001 ;
  assign n1003 = n169 & ~n1002 ;
  assign n1005 = ~n999 & ~n1003 ;
  assign n1006 = n1004 & n1005 ;
  assign n1007 = n318 & ~n1006 ;
  assign n1009 = ~n987 & ~n1007 ;
  assign n1010 = n1008 & n1009 ;
  assign n1011 = ~\shift[6]  & ~n1010 ;
  assign n1012 = \shift[1]  & ~n418 ;
  assign n1013 = ~\shift[1]  & ~n161 ;
  assign n1014 = ~n1012 & ~n1013 ;
  assign n1015 = n136 & ~n1014 ;
  assign n1016 = \shift[1]  & ~n428 ;
  assign n1017 = ~\shift[1]  & ~n414 ;
  assign n1018 = ~n1016 & ~n1017 ;
  assign n1019 = n147 & ~n1018 ;
  assign n1028 = ~n1015 & ~n1019 ;
  assign n1020 = \shift[1]  & ~n438 ;
  assign n1021 = ~\shift[1]  & ~n444 ;
  assign n1022 = ~n1020 & ~n1021 ;
  assign n1023 = n158 & ~n1022 ;
  assign n1024 = \shift[1]  & ~n448 ;
  assign n1025 = ~\shift[1]  & ~n424 ;
  assign n1026 = ~n1024 & ~n1025 ;
  assign n1027 = n169 & ~n1026 ;
  assign n1029 = ~n1023 & ~n1027 ;
  assign n1030 = n1028 & n1029 ;
  assign n1031 = n273 & ~n1030 ;
  assign n1032 = \shift[1]  & ~n330 ;
  assign n1033 = ~\shift[1]  & ~n390 ;
  assign n1034 = ~n1032 & ~n1033 ;
  assign n1035 = n136 & ~n1034 ;
  assign n1036 = \shift[1]  & ~n340 ;
  assign n1037 = ~\shift[1]  & ~n326 ;
  assign n1038 = ~n1036 & ~n1037 ;
  assign n1039 = n147 & ~n1038 ;
  assign n1048 = ~n1035 & ~n1039 ;
  assign n1040 = \shift[1]  & ~n350 ;
  assign n1041 = ~\shift[1]  & ~n356 ;
  assign n1042 = ~n1040 & ~n1041 ;
  assign n1043 = n158 & ~n1042 ;
  assign n1044 = \shift[1]  & ~n360 ;
  assign n1045 = ~\shift[1]  & ~n336 ;
  assign n1046 = ~n1044 & ~n1045 ;
  assign n1047 = n169 & ~n1046 ;
  assign n1049 = ~n1043 & ~n1047 ;
  assign n1050 = n1048 & n1049 ;
  assign n1051 = n183 & ~n1050 ;
  assign n1094 = ~n1031 & ~n1051 ;
  assign n1052 = \shift[1]  & ~n462 ;
  assign n1053 = ~\shift[1]  & ~n434 ;
  assign n1054 = ~n1052 & ~n1053 ;
  assign n1055 = n136 & ~n1054 ;
  assign n1056 = \shift[1]  & ~n472 ;
  assign n1057 = ~\shift[1]  & ~n458 ;
  assign n1058 = ~n1056 & ~n1057 ;
  assign n1059 = n147 & ~n1058 ;
  assign n1070 = ~n1055 & ~n1059 ;
  assign n1060 = ~n488 & ~n491 ;
  assign n1061 = ~\shift[1]  & ~n1060 ;
  assign n1062 = \shift[1]  & ~n482 ;
  assign n1063 = ~n1061 & ~n1062 ;
  assign n1064 = n158 & ~n1063 ;
  assign n1065 = ~\shift[1]  & ~n468 ;
  assign n1066 = ~n486 & ~n493 ;
  assign n1067 = \shift[1]  & ~n1066 ;
  assign n1068 = ~n1065 & ~n1067 ;
  assign n1069 = n169 & ~n1068 ;
  assign n1071 = ~n1064 & ~n1069 ;
  assign n1072 = n1070 & n1071 ;
  assign n1073 = n318 & ~n1072 ;
  assign n1074 = \shift[1]  & ~n374 ;
  assign n1075 = ~\shift[1]  & ~n478 ;
  assign n1076 = ~n1074 & ~n1075 ;
  assign n1077 = n136 & ~n1076 ;
  assign n1078 = \shift[1]  & ~n384 ;
  assign n1079 = ~\shift[1]  & ~n370 ;
  assign n1080 = ~n1078 & ~n1079 ;
  assign n1081 = n147 & ~n1080 ;
  assign n1090 = ~n1077 & ~n1081 ;
  assign n1082 = \shift[1]  & ~n394 ;
  assign n1083 = ~\shift[1]  & ~n400 ;
  assign n1084 = ~n1082 & ~n1083 ;
  assign n1085 = n158 & ~n1084 ;
  assign n1086 = \shift[1]  & ~n404 ;
  assign n1087 = ~\shift[1]  & ~n380 ;
  assign n1088 = ~n1086 & ~n1087 ;
  assign n1089 = n169 & ~n1088 ;
  assign n1091 = ~n1085 & ~n1089 ;
  assign n1092 = n1090 & n1091 ;
  assign n1093 = n228 & ~n1092 ;
  assign n1095 = ~n1073 & ~n1093 ;
  assign n1096 = n1094 & n1095 ;
  assign n1097 = \shift[6]  & ~n1096 ;
  assign n1098 = ~n1011 & ~n1097 ;
  assign n1099 = ~\shift[1]  & ~n637 ;
  assign n1100 = \shift[1]  & ~n663 ;
  assign n1101 = ~n1099 & ~n1100 ;
  assign n1102 = \shift[1]  & n670 ;
  assign n1103 = ~\shift[1]  & n640 ;
  assign n1104 = ~n1102 & ~n1103 ;
  assign n1105 = ~n1101 & n1104 ;
  assign n1106 = n136 & ~n1105 ;
  assign n1107 = ~\shift[1]  & ~n665 ;
  assign n1108 = \shift[1]  & ~n675 ;
  assign n1109 = ~n1107 & ~n1108 ;
  assign n1110 = \shift[1]  & n682 ;
  assign n1111 = ~\shift[1]  & n668 ;
  assign n1112 = ~n1110 & ~n1111 ;
  assign n1113 = ~n1109 & n1112 ;
  assign n1114 = n147 & ~n1113 ;
  assign n1131 = ~n1106 & ~n1114 ;
  assign n1115 = ~\shift[1]  & ~n701 ;
  assign n1116 = \shift[1]  & ~n687 ;
  assign n1117 = ~n1115 & ~n1116 ;
  assign n1118 = \shift[1]  & n694 ;
  assign n1119 = ~\shift[1]  & n704 ;
  assign n1120 = ~n1118 & ~n1119 ;
  assign n1121 = ~n1117 & n1120 ;
  assign n1122 = n158 & ~n1121 ;
  assign n1123 = ~\shift[1]  & ~n677 ;
  assign n1124 = \shift[1]  & ~n699 ;
  assign n1125 = ~n1123 & ~n1124 ;
  assign n1126 = \shift[1]  & n706 ;
  assign n1127 = ~\shift[1]  & n680 ;
  assign n1128 = ~n1126 & ~n1127 ;
  assign n1129 = ~n1125 & n1128 ;
  assign n1130 = n169 & ~n1129 ;
  assign n1132 = ~n1122 & ~n1130 ;
  assign n1133 = n1131 & n1132 ;
  assign n1134 = n318 & ~n1133 ;
  assign n1135 = ~\shift[1]  & ~n689 ;
  assign n1136 = \shift[1]  & ~n559 ;
  assign n1137 = ~n1135 & ~n1136 ;
  assign n1138 = \shift[1]  & n566 ;
  assign n1139 = ~\shift[1]  & n692 ;
  assign n1140 = ~n1138 & ~n1139 ;
  assign n1141 = ~n1137 & n1140 ;
  assign n1142 = n136 & ~n1141 ;
  assign n1143 = ~\shift[1]  & ~n561 ;
  assign n1144 = \shift[1]  & ~n571 ;
  assign n1145 = ~n1143 & ~n1144 ;
  assign n1146 = \shift[1]  & n578 ;
  assign n1147 = ~\shift[1]  & n564 ;
  assign n1148 = ~n1146 & ~n1147 ;
  assign n1149 = ~n1145 & n1148 ;
  assign n1150 = n147 & ~n1149 ;
  assign n1167 = ~n1142 & ~n1150 ;
  assign n1151 = ~\shift[1]  & ~n597 ;
  assign n1152 = \shift[1]  & ~n583 ;
  assign n1153 = ~n1151 & ~n1152 ;
  assign n1154 = \shift[1]  & n590 ;
  assign n1155 = ~\shift[1]  & n600 ;
  assign n1156 = ~n1154 & ~n1155 ;
  assign n1157 = ~n1153 & n1156 ;
  assign n1158 = n158 & ~n1157 ;
  assign n1159 = ~\shift[1]  & ~n573 ;
  assign n1160 = \shift[1]  & ~n595 ;
  assign n1161 = ~n1159 & ~n1160 ;
  assign n1162 = \shift[1]  & n602 ;
  assign n1163 = ~\shift[1]  & n576 ;
  assign n1164 = ~n1162 & ~n1163 ;
  assign n1165 = ~n1161 & n1164 ;
  assign n1166 = n169 & ~n1165 ;
  assign n1168 = ~n1158 & ~n1166 ;
  assign n1169 = n1167 & n1168 ;
  assign n1170 = n228 & ~n1169 ;
  assign n1243 = ~n1134 & ~n1170 ;
  assign n1171 = ~\shift[1]  & ~n797 ;
  assign n1172 = \shift[1]  & ~n611 ;
  assign n1173 = ~n1171 & ~n1172 ;
  assign n1174 = \shift[1]  & n618 ;
  assign n1175 = ~\shift[1]  & n800 ;
  assign n1176 = ~n1174 & ~n1175 ;
  assign n1177 = ~n1173 & n1176 ;
  assign n1178 = n136 & ~n1177 ;
  assign n1179 = ~\shift[1]  & ~n613 ;
  assign n1180 = \shift[1]  & ~n623 ;
  assign n1181 = ~n1179 & ~n1180 ;
  assign n1182 = \shift[1]  & n630 ;
  assign n1183 = ~\shift[1]  & n616 ;
  assign n1184 = ~n1182 & ~n1183 ;
  assign n1185 = ~n1181 & n1184 ;
  assign n1186 = n147 & ~n1185 ;
  assign n1203 = ~n1178 & ~n1186 ;
  assign n1187 = ~\shift[1]  & ~n649 ;
  assign n1188 = \shift[1]  & ~n635 ;
  assign n1189 = ~n1187 & ~n1188 ;
  assign n1190 = \shift[1]  & n642 ;
  assign n1191 = ~\shift[1]  & n652 ;
  assign n1192 = ~n1190 & ~n1191 ;
  assign n1193 = ~n1189 & n1192 ;
  assign n1194 = n158 & ~n1193 ;
  assign n1195 = ~\shift[1]  & ~n625 ;
  assign n1196 = \shift[1]  & ~n647 ;
  assign n1197 = ~n1195 & ~n1196 ;
  assign n1198 = \shift[1]  & n654 ;
  assign n1199 = ~\shift[1]  & n628 ;
  assign n1200 = ~n1198 & ~n1199 ;
  assign n1201 = ~n1197 & n1200 ;
  assign n1202 = n169 & ~n1201 ;
  assign n1204 = ~n1194 & ~n1202 ;
  assign n1205 = n1203 & n1204 ;
  assign n1206 = n273 & ~n1205 ;
  assign n1207 = ~\shift[1]  & ~n585 ;
  assign n1208 = \shift[1]  & ~n507 ;
  assign n1209 = ~n1207 & ~n1208 ;
  assign n1210 = \shift[1]  & n514 ;
  assign n1211 = ~\shift[1]  & n588 ;
  assign n1212 = ~n1210 & ~n1211 ;
  assign n1213 = ~n1209 & n1212 ;
  assign n1214 = n136 & ~n1213 ;
  assign n1215 = ~\shift[1]  & ~n509 ;
  assign n1216 = \shift[1]  & ~n519 ;
  assign n1217 = ~n1215 & ~n1216 ;
  assign n1218 = \shift[1]  & n526 ;
  assign n1219 = ~\shift[1]  & n512 ;
  assign n1220 = ~n1218 & ~n1219 ;
  assign n1221 = ~n1217 & n1220 ;
  assign n1222 = n147 & ~n1221 ;
  assign n1239 = ~n1214 & ~n1222 ;
  assign n1223 = ~\shift[1]  & ~n545 ;
  assign n1224 = \shift[1]  & ~n531 ;
  assign n1225 = ~n1223 & ~n1224 ;
  assign n1226 = \shift[1]  & n538 ;
  assign n1227 = ~\shift[1]  & n548 ;
  assign n1228 = ~n1226 & ~n1227 ;
  assign n1229 = ~n1225 & n1228 ;
  assign n1230 = n158 & ~n1229 ;
  assign n1231 = ~\shift[1]  & ~n521 ;
  assign n1232 = \shift[1]  & ~n543 ;
  assign n1233 = ~n1231 & ~n1232 ;
  assign n1234 = \shift[1]  & n550 ;
  assign n1235 = ~\shift[1]  & n524 ;
  assign n1236 = ~n1234 & ~n1235 ;
  assign n1237 = ~n1233 & n1236 ;
  assign n1238 = n169 & ~n1237 ;
  assign n1240 = ~n1230 & ~n1238 ;
  assign n1241 = n1239 & n1240 ;
  assign n1242 = n183 & ~n1241 ;
  assign n1244 = ~n1206 & ~n1242 ;
  assign n1245 = n1243 & n1244 ;
  assign n1246 = ~\shift[6]  & ~n1245 ;
  assign n1247 = ~\shift[1]  & ~n533 ;
  assign n1248 = \shift[1]  & ~n719 ;
  assign n1249 = ~n1247 & ~n1248 ;
  assign n1250 = \shift[1]  & n726 ;
  assign n1251 = ~\shift[1]  & n536 ;
  assign n1252 = ~n1250 & ~n1251 ;
  assign n1253 = ~n1249 & n1252 ;
  assign n1254 = n136 & ~n1253 ;
  assign n1255 = ~\shift[1]  & ~n721 ;
  assign n1256 = \shift[1]  & ~n731 ;
  assign n1257 = ~n1255 & ~n1256 ;
  assign n1258 = \shift[1]  & n738 ;
  assign n1259 = ~\shift[1]  & n724 ;
  assign n1260 = ~n1258 & ~n1259 ;
  assign n1261 = ~n1257 & n1260 ;
  assign n1262 = n147 & ~n1261 ;
  assign n1279 = ~n1254 & ~n1262 ;
  assign n1263 = ~\shift[1]  & ~n757 ;
  assign n1264 = \shift[1]  & ~n743 ;
  assign n1265 = ~n1263 & ~n1264 ;
  assign n1266 = \shift[1]  & n750 ;
  assign n1267 = ~\shift[1]  & n760 ;
  assign n1268 = ~n1266 & ~n1267 ;
  assign n1269 = ~n1265 & n1268 ;
  assign n1270 = n158 & ~n1269 ;
  assign n1271 = ~\shift[1]  & ~n733 ;
  assign n1272 = \shift[1]  & ~n755 ;
  assign n1273 = ~n1271 & ~n1272 ;
  assign n1274 = \shift[1]  & n762 ;
  assign n1275 = ~\shift[1]  & n736 ;
  assign n1276 = ~n1274 & ~n1275 ;
  assign n1277 = ~n1273 & n1276 ;
  assign n1278 = n169 & ~n1277 ;
  assign n1280 = ~n1270 & ~n1278 ;
  assign n1281 = n1279 & n1280 ;
  assign n1282 = n273 & ~n1281 ;
  assign n1283 = ~\shift[1]  & ~n745 ;
  assign n1284 = \shift[1]  & ~n823 ;
  assign n1285 = ~n1283 & ~n1284 ;
  assign n1286 = \shift[1]  & n830 ;
  assign n1287 = ~\shift[1]  & n748 ;
  assign n1288 = ~n1286 & ~n1287 ;
  assign n1289 = ~n1285 & n1288 ;
  assign n1290 = n136 & ~n1289 ;
  assign n1291 = \shift[1]  & ~n841 ;
  assign n1292 = ~n825 & ~n828 ;
  assign n1293 = ~\shift[1]  & ~n1292 ;
  assign n1294 = ~n1291 & ~n1293 ;
  assign n1295 = n147 & ~n1294 ;
  assign n1312 = ~n1290 & ~n1295 ;
  assign n1296 = ~\shift[1]  & ~n862 ;
  assign n1297 = \shift[1]  & ~n845 ;
  assign n1298 = ~n1296 & ~n1297 ;
  assign n1299 = \shift[1]  & n852 ;
  assign n1300 = ~\shift[1]  & n861 ;
  assign n1301 = ~n1299 & ~n1300 ;
  assign n1302 = ~n1298 & n1301 ;
  assign n1303 = n158 & ~n1302 ;
  assign n1304 = ~\shift[1]  & ~n835 ;
  assign n1305 = \shift[1]  & ~n857 ;
  assign n1306 = ~n1304 & ~n1305 ;
  assign n1307 = \shift[1]  & n858 ;
  assign n1308 = ~\shift[1]  & n836 ;
  assign n1309 = ~n1307 & ~n1308 ;
  assign n1310 = ~n1306 & n1309 ;
  assign n1311 = n169 & ~n1310 ;
  assign n1313 = ~n1303 & ~n1311 ;
  assign n1314 = n1312 & n1313 ;
  assign n1315 = n318 & ~n1314 ;
  assign n1388 = ~n1282 & ~n1315 ;
  assign n1316 = ~\shift[1]  & ~n897 ;
  assign n1317 = \shift[1]  & ~n771 ;
  assign n1318 = ~n1316 & ~n1317 ;
  assign n1319 = \shift[1]  & n778 ;
  assign n1320 = ~\shift[1]  & n900 ;
  assign n1321 = ~n1319 & ~n1320 ;
  assign n1322 = ~n1318 & n1321 ;
  assign n1323 = n136 & ~n1322 ;
  assign n1324 = ~\shift[1]  & ~n773 ;
  assign n1325 = \shift[1]  & ~n783 ;
  assign n1326 = ~n1324 & ~n1325 ;
  assign n1327 = \shift[1]  & n790 ;
  assign n1328 = ~\shift[1]  & n776 ;
  assign n1329 = ~n1327 & ~n1328 ;
  assign n1330 = ~n1326 & n1329 ;
  assign n1331 = n147 & ~n1330 ;
  assign n1348 = ~n1323 & ~n1331 ;
  assign n1332 = ~\shift[1]  & ~n809 ;
  assign n1333 = \shift[1]  & ~n795 ;
  assign n1334 = ~n1332 & ~n1333 ;
  assign n1335 = \shift[1]  & n802 ;
  assign n1336 = ~\shift[1]  & n812 ;
  assign n1337 = ~n1335 & ~n1336 ;
  assign n1338 = ~n1334 & n1337 ;
  assign n1339 = n158 & ~n1338 ;
  assign n1340 = ~\shift[1]  & ~n785 ;
  assign n1341 = \shift[1]  & ~n807 ;
  assign n1342 = ~n1340 & ~n1341 ;
  assign n1343 = \shift[1]  & n814 ;
  assign n1344 = ~\shift[1]  & n788 ;
  assign n1345 = ~n1343 & ~n1344 ;
  assign n1346 = ~n1342 & n1345 ;
  assign n1347 = n169 & ~n1346 ;
  assign n1349 = ~n1339 & ~n1347 ;
  assign n1350 = n1348 & n1349 ;
  assign n1351 = n183 & ~n1350 ;
  assign n1352 = ~\shift[1]  & ~n847 ;
  assign n1353 = \shift[1]  & ~n871 ;
  assign n1354 = ~n1352 & ~n1353 ;
  assign n1355 = \shift[1]  & n878 ;
  assign n1356 = ~\shift[1]  & n850 ;
  assign n1357 = ~n1355 & ~n1356 ;
  assign n1358 = ~n1354 & n1357 ;
  assign n1359 = n136 & ~n1358 ;
  assign n1360 = ~\shift[1]  & ~n873 ;
  assign n1361 = \shift[1]  & ~n883 ;
  assign n1362 = ~n1360 & ~n1361 ;
  assign n1363 = \shift[1]  & n890 ;
  assign n1364 = ~\shift[1]  & n876 ;
  assign n1365 = ~n1363 & ~n1364 ;
  assign n1366 = ~n1362 & n1365 ;
  assign n1367 = n147 & ~n1366 ;
  assign n1384 = ~n1359 & ~n1367 ;
  assign n1368 = ~\shift[1]  & ~n909 ;
  assign n1369 = \shift[1]  & ~n895 ;
  assign n1370 = ~n1368 & ~n1369 ;
  assign n1371 = \shift[1]  & n902 ;
  assign n1372 = ~\shift[1]  & n912 ;
  assign n1373 = ~n1371 & ~n1372 ;
  assign n1374 = ~n1370 & n1373 ;
  assign n1375 = n158 & ~n1374 ;
  assign n1376 = ~\shift[1]  & ~n885 ;
  assign n1377 = \shift[1]  & ~n907 ;
  assign n1378 = ~n1376 & ~n1377 ;
  assign n1379 = \shift[1]  & n914 ;
  assign n1380 = ~\shift[1]  & n888 ;
  assign n1381 = ~n1379 & ~n1380 ;
  assign n1382 = ~n1378 & n1381 ;
  assign n1383 = n169 & ~n1382 ;
  assign n1385 = ~n1375 & ~n1383 ;
  assign n1386 = n1384 & n1385 ;
  assign n1387 = n228 & ~n1386 ;
  assign n1389 = ~n1351 & ~n1387 ;
  assign n1390 = n1388 & n1389 ;
  assign n1391 = \shift[6]  & ~n1390 ;
  assign n1392 = ~n1246 & ~n1391 ;
  assign n1393 = n136 & ~n213 ;
  assign n1394 = ~n145 & n147 ;
  assign n1397 = ~n1393 & ~n1394 ;
  assign n1395 = n158 & ~n178 ;
  assign n1396 = ~n156 & n169 ;
  assign n1398 = ~n1395 & ~n1396 ;
  assign n1399 = n1397 & n1398 ;
  assign n1400 = n183 & ~n1399 ;
  assign n1401 = n136 & ~n303 ;
  assign n1402 = n147 & ~n193 ;
  assign n1405 = ~n1401 & ~n1402 ;
  assign n1403 = n158 & ~n223 ;
  assign n1404 = n169 & ~n203 ;
  assign n1406 = ~n1403 & ~n1404 ;
  assign n1407 = n1405 & n1406 ;
  assign n1408 = n228 & ~n1407 ;
  assign n1425 = ~n1400 & ~n1408 ;
  assign n1409 = n136 & ~n352 ;
  assign n1410 = n147 & ~n238 ;
  assign n1413 = ~n1409 & ~n1410 ;
  assign n1411 = n158 & ~n268 ;
  assign n1412 = n169 & ~n248 ;
  assign n1414 = ~n1411 & ~n1412 ;
  assign n1415 = n1413 & n1414 ;
  assign n1416 = n273 & ~n1415 ;
  assign n1417 = n136 & ~n258 ;
  assign n1418 = n147 & ~n283 ;
  assign n1421 = ~n1417 & ~n1418 ;
  assign n1419 = n158 & ~n313 ;
  assign n1420 = n169 & ~n293 ;
  assign n1422 = ~n1419 & ~n1420 ;
  assign n1423 = n1421 & n1422 ;
  assign n1424 = n318 & ~n1423 ;
  assign n1426 = ~n1416 & ~n1424 ;
  assign n1427 = n1425 & n1426 ;
  assign n1428 = ~\shift[6]  & ~n1427 ;
  assign n1429 = n136 & ~n440 ;
  assign n1430 = n147 & ~n464 ;
  assign n1433 = ~n1429 & ~n1430 ;
  assign n1431 = n158 & ~n496 ;
  assign n1432 = n169 & ~n474 ;
  assign n1434 = ~n1431 & ~n1432 ;
  assign n1435 = n1433 & n1434 ;
  assign n1436 = n318 & ~n1435 ;
  assign n1437 = n136 & ~n167 ;
  assign n1438 = n147 & ~n420 ;
  assign n1441 = ~n1437 & ~n1438 ;
  assign n1439 = n158 & ~n450 ;
  assign n1440 = n169 & ~n430 ;
  assign n1442 = ~n1439 & ~n1440 ;
  assign n1443 = n1441 & n1442 ;
  assign n1444 = n273 & ~n1443 ;
  assign n1461 = ~n1436 & ~n1444 ;
  assign n1445 = n136 & ~n484 ;
  assign n1446 = n147 & ~n376 ;
  assign n1449 = ~n1445 & ~n1446 ;
  assign n1447 = n158 & ~n406 ;
  assign n1448 = n169 & ~n386 ;
  assign n1450 = ~n1447 & ~n1448 ;
  assign n1451 = n1449 & n1450 ;
  assign n1452 = n228 & ~n1451 ;
  assign n1453 = n136 & ~n396 ;
  assign n1454 = n147 & ~n332 ;
  assign n1457 = ~n1453 & ~n1454 ;
  assign n1455 = n158 & ~n362 ;
  assign n1456 = n169 & ~n342 ;
  assign n1458 = ~n1455 & ~n1456 ;
  assign n1459 = n1457 & n1458 ;
  assign n1460 = n183 & ~n1459 ;
  assign n1462 = ~n1452 & ~n1460 ;
  assign n1463 = n1461 & n1462 ;
  assign n1464 = \shift[6]  & ~n1463 ;
  assign n1465 = ~n1428 & ~n1464 ;
  assign n1466 = n136 & ~n593 ;
  assign n1467 = n147 & ~n517 ;
  assign n1470 = ~n1466 & ~n1467 ;
  assign n1468 = n158 & ~n553 ;
  assign n1469 = n169 & ~n529 ;
  assign n1471 = ~n1468 & ~n1469 ;
  assign n1472 = n1470 & n1471 ;
  assign n1473 = n183 & ~n1472 ;
  assign n1474 = n136 & ~n697 ;
  assign n1475 = n147 & ~n569 ;
  assign n1478 = ~n1474 & ~n1475 ;
  assign n1476 = n158 & ~n605 ;
  assign n1477 = n169 & ~n581 ;
  assign n1479 = ~n1476 & ~n1477 ;
  assign n1480 = n1478 & n1479 ;
  assign n1481 = n228 & ~n1480 ;
  assign n1498 = ~n1473 & ~n1481 ;
  assign n1482 = n136 & ~n805 ;
  assign n1483 = n147 & ~n621 ;
  assign n1486 = ~n1482 & ~n1483 ;
  assign n1484 = n158 & ~n657 ;
  assign n1485 = n169 & ~n633 ;
  assign n1487 = ~n1484 & ~n1485 ;
  assign n1488 = n1486 & n1487 ;
  assign n1489 = n273 & ~n1488 ;
  assign n1490 = n136 & ~n645 ;
  assign n1491 = n147 & ~n673 ;
  assign n1494 = ~n1490 & ~n1491 ;
  assign n1492 = n158 & ~n709 ;
  assign n1493 = n169 & ~n685 ;
  assign n1495 = ~n1492 & ~n1493 ;
  assign n1496 = n1494 & n1495 ;
  assign n1497 = n318 & ~n1496 ;
  assign n1499 = ~n1489 & ~n1497 ;
  assign n1500 = n1498 & n1499 ;
  assign n1501 = ~\shift[6]  & ~n1500 ;
  assign n1502 = n136 & ~n753 ;
  assign n1503 = n147 & ~n833 ;
  assign n1506 = ~n1502 & ~n1503 ;
  assign n1504 = n158 & ~n865 ;
  assign n1505 = n169 & ~n843 ;
  assign n1507 = ~n1504 & ~n1505 ;
  assign n1508 = n1506 & n1507 ;
  assign n1509 = n318 & ~n1508 ;
  assign n1510 = n136 & ~n541 ;
  assign n1511 = n147 & ~n729 ;
  assign n1514 = ~n1510 & ~n1511 ;
  assign n1512 = n158 & ~n765 ;
  assign n1513 = n169 & ~n741 ;
  assign n1515 = ~n1512 & ~n1513 ;
  assign n1516 = n1514 & n1515 ;
  assign n1517 = n273 & ~n1516 ;
  assign n1534 = ~n1509 & ~n1517 ;
  assign n1518 = n136 & ~n855 ;
  assign n1519 = n147 & ~n881 ;
  assign n1522 = ~n1518 & ~n1519 ;
  assign n1520 = n158 & ~n917 ;
  assign n1521 = n169 & ~n893 ;
  assign n1523 = ~n1520 & ~n1521 ;
  assign n1524 = n1522 & n1523 ;
  assign n1525 = n228 & ~n1524 ;
  assign n1526 = n136 & ~n905 ;
  assign n1527 = n147 & ~n781 ;
  assign n1530 = ~n1526 & ~n1527 ;
  assign n1528 = n158 & ~n817 ;
  assign n1529 = n169 & ~n793 ;
  assign n1531 = ~n1528 & ~n1529 ;
  assign n1532 = n1530 & n1531 ;
  assign n1533 = n183 & ~n1532 ;
  assign n1535 = ~n1525 & ~n1533 ;
  assign n1536 = n1534 & n1535 ;
  assign n1537 = \shift[6]  & ~n1536 ;
  assign n1538 = ~n1501 & ~n1537 ;
  assign n1539 = n136 & ~n958 ;
  assign n1540 = n147 & ~n930 ;
  assign n1543 = ~n1539 & ~n1540 ;
  assign n1541 = n158 & ~n942 ;
  assign n1542 = n169 & ~n934 ;
  assign n1544 = ~n1541 & ~n1542 ;
  assign n1545 = n1543 & n1544 ;
  assign n1546 = n183 & ~n1545 ;
  assign n1547 = n136 & ~n998 ;
  assign n1548 = n147 & ~n950 ;
  assign n1551 = ~n1547 & ~n1548 ;
  assign n1549 = n158 & ~n962 ;
  assign n1550 = n169 & ~n954 ;
  assign n1552 = ~n1549 & ~n1550 ;
  assign n1553 = n1551 & n1552 ;
  assign n1554 = n228 & ~n1553 ;
  assign n1571 = ~n1546 & ~n1554 ;
  assign n1555 = n136 & ~n1042 ;
  assign n1556 = n147 & ~n970 ;
  assign n1559 = ~n1555 & ~n1556 ;
  assign n1557 = n158 & ~n982 ;
  assign n1558 = n169 & ~n974 ;
  assign n1560 = ~n1557 & ~n1558 ;
  assign n1561 = n1559 & n1560 ;
  assign n1562 = n273 & ~n1561 ;
  assign n1563 = n136 & ~n978 ;
  assign n1564 = n147 & ~n990 ;
  assign n1567 = ~n1563 & ~n1564 ;
  assign n1565 = n158 & ~n1002 ;
  assign n1566 = n169 & ~n994 ;
  assign n1568 = ~n1565 & ~n1566 ;
  assign n1569 = n1567 & n1568 ;
  assign n1570 = n318 & ~n1569 ;
  assign n1572 = ~n1562 & ~n1570 ;
  assign n1573 = n1571 & n1572 ;
  assign n1574 = ~\shift[6]  & ~n1573 ;
  assign n1575 = n136 & ~n1022 ;
  assign n1576 = n147 & ~n1054 ;
  assign n1579 = ~n1575 & ~n1576 ;
  assign n1577 = n158 & ~n1068 ;
  assign n1578 = n169 & ~n1058 ;
  assign n1580 = ~n1577 & ~n1578 ;
  assign n1581 = n1579 & n1580 ;
  assign n1582 = n318 & ~n1581 ;
  assign n1583 = n136 & ~n938 ;
  assign n1584 = n147 & ~n1014 ;
  assign n1587 = ~n1583 & ~n1584 ;
  assign n1585 = n158 & ~n1026 ;
  assign n1586 = n169 & ~n1018 ;
  assign n1588 = ~n1585 & ~n1586 ;
  assign n1589 = n1587 & n1588 ;
  assign n1590 = n273 & ~n1589 ;
  assign n1607 = ~n1582 & ~n1590 ;
  assign n1591 = n136 & ~n1063 ;
  assign n1592 = n147 & ~n1076 ;
  assign n1595 = ~n1591 & ~n1592 ;
  assign n1593 = n158 & ~n1088 ;
  assign n1594 = n169 & ~n1080 ;
  assign n1596 = ~n1593 & ~n1594 ;
  assign n1597 = n1595 & n1596 ;
  assign n1598 = n228 & ~n1597 ;
  assign n1599 = n136 & ~n1084 ;
  assign n1600 = n147 & ~n1034 ;
  assign n1603 = ~n1599 & ~n1600 ;
  assign n1601 = n158 & ~n1046 ;
  assign n1602 = n169 & ~n1038 ;
  assign n1604 = ~n1601 & ~n1602 ;
  assign n1605 = n1603 & n1604 ;
  assign n1606 = n183 & ~n1605 ;
  assign n1608 = ~n1598 & ~n1606 ;
  assign n1609 = n1607 & n1608 ;
  assign n1610 = \shift[6]  & ~n1609 ;
  assign n1611 = ~n1574 & ~n1610 ;
  assign n1612 = n136 & ~n1157 ;
  assign n1613 = n147 & ~n1213 ;
  assign n1616 = ~n1612 & ~n1613 ;
  assign n1614 = n158 & ~n1237 ;
  assign n1615 = n169 & ~n1221 ;
  assign n1617 = ~n1614 & ~n1615 ;
  assign n1618 = n1616 & n1617 ;
  assign n1619 = n183 & ~n1618 ;
  assign n1620 = n136 & ~n1121 ;
  assign n1621 = n147 & ~n1141 ;
  assign n1624 = ~n1620 & ~n1621 ;
  assign n1622 = n158 & ~n1165 ;
  assign n1623 = n169 & ~n1149 ;
  assign n1625 = ~n1622 & ~n1623 ;
  assign n1626 = n1624 & n1625 ;
  assign n1627 = n228 & ~n1626 ;
  assign n1644 = ~n1619 & ~n1627 ;
  assign n1628 = n136 & ~n1338 ;
  assign n1629 = n147 & ~n1177 ;
  assign n1632 = ~n1628 & ~n1629 ;
  assign n1630 = n158 & ~n1201 ;
  assign n1631 = n169 & ~n1185 ;
  assign n1633 = ~n1630 & ~n1631 ;
  assign n1634 = n1632 & n1633 ;
  assign n1635 = n273 & ~n1634 ;
  assign n1636 = n136 & ~n1193 ;
  assign n1637 = n147 & ~n1105 ;
  assign n1640 = ~n1636 & ~n1637 ;
  assign n1638 = n158 & ~n1129 ;
  assign n1639 = n169 & ~n1113 ;
  assign n1641 = ~n1638 & ~n1639 ;
  assign n1642 = n1640 & n1641 ;
  assign n1643 = n318 & ~n1642 ;
  assign n1645 = ~n1635 & ~n1643 ;
  assign n1646 = n1644 & n1645 ;
  assign n1647 = ~\shift[6]  & ~n1646 ;
  assign n1648 = n147 & ~n1289 ;
  assign n1649 = n169 & ~n1294 ;
  assign n1652 = ~n1648 & ~n1649 ;
  assign n1650 = n158 & ~n1310 ;
  assign n1651 = n136 & ~n1269 ;
  assign n1653 = ~n1650 & ~n1651 ;
  assign n1654 = n1652 & n1653 ;
  assign n1655 = n318 & ~n1654 ;
  assign n1656 = n136 & ~n1229 ;
  assign n1657 = n147 & ~n1253 ;
  assign n1660 = ~n1656 & ~n1657 ;
  assign n1658 = n158 & ~n1277 ;
  assign n1659 = n169 & ~n1261 ;
  assign n1661 = ~n1658 & ~n1659 ;
  assign n1662 = n1660 & n1661 ;
  assign n1663 = n273 & ~n1662 ;
  assign n1680 = ~n1655 & ~n1663 ;
  assign n1664 = n136 & ~n1302 ;
  assign n1665 = n147 & ~n1358 ;
  assign n1668 = ~n1664 & ~n1665 ;
  assign n1666 = n158 & ~n1382 ;
  assign n1667 = n169 & ~n1366 ;
  assign n1669 = ~n1666 & ~n1667 ;
  assign n1670 = n1668 & n1669 ;
  assign n1671 = n228 & ~n1670 ;
  assign n1672 = n136 & ~n1374 ;
  assign n1673 = n147 & ~n1322 ;
  assign n1676 = ~n1672 & ~n1673 ;
  assign n1674 = n158 & ~n1346 ;
  assign n1675 = n169 & ~n1330 ;
  assign n1677 = ~n1674 & ~n1675 ;
  assign n1678 = n1676 & n1677 ;
  assign n1679 = n183 & ~n1678 ;
  assign n1681 = ~n1671 & ~n1679 ;
  assign n1682 = n1680 & n1681 ;
  assign n1683 = \shift[6]  & ~n1682 ;
  assign n1684 = ~n1647 & ~n1683 ;
  assign n1685 = n136 & ~n223 ;
  assign n1686 = n147 & ~n213 ;
  assign n1689 = ~n1685 & ~n1686 ;
  assign n1687 = ~n156 & n158 ;
  assign n1688 = ~n145 & n169 ;
  assign n1690 = ~n1687 & ~n1688 ;
  assign n1691 = n1689 & n1690 ;
  assign n1692 = n183 & ~n1691 ;
  assign n1693 = n136 & ~n313 ;
  assign n1694 = n147 & ~n303 ;
  assign n1697 = ~n1693 & ~n1694 ;
  assign n1695 = n158 & ~n203 ;
  assign n1696 = n169 & ~n193 ;
  assign n1698 = ~n1695 & ~n1696 ;
  assign n1699 = n1697 & n1698 ;
  assign n1700 = n228 & ~n1699 ;
  assign n1717 = ~n1692 & ~n1700 ;
  assign n1701 = n136 & ~n362 ;
  assign n1702 = n147 & ~n352 ;
  assign n1705 = ~n1701 & ~n1702 ;
  assign n1703 = n158 & ~n248 ;
  assign n1704 = n169 & ~n238 ;
  assign n1706 = ~n1703 & ~n1704 ;
  assign n1707 = n1705 & n1706 ;
  assign n1708 = n273 & ~n1707 ;
  assign n1709 = n136 & ~n268 ;
  assign n1710 = n147 & ~n258 ;
  assign n1713 = ~n1709 & ~n1710 ;
  assign n1711 = n158 & ~n293 ;
  assign n1712 = n169 & ~n283 ;
  assign n1714 = ~n1711 & ~n1712 ;
  assign n1715 = n1713 & n1714 ;
  assign n1716 = n318 & ~n1715 ;
  assign n1718 = ~n1708 & ~n1716 ;
  assign n1719 = n1717 & n1718 ;
  assign n1720 = ~\shift[6]  & ~n1719 ;
  assign n1721 = n136 & ~n450 ;
  assign n1722 = n147 & ~n440 ;
  assign n1725 = ~n1721 & ~n1722 ;
  assign n1723 = n158 & ~n474 ;
  assign n1724 = n169 & ~n464 ;
  assign n1726 = ~n1723 & ~n1724 ;
  assign n1727 = n1725 & n1726 ;
  assign n1728 = n318 & ~n1727 ;
  assign n1729 = n136 & ~n178 ;
  assign n1730 = n147 & ~n167 ;
  assign n1733 = ~n1729 & ~n1730 ;
  assign n1731 = n158 & ~n430 ;
  assign n1732 = n169 & ~n420 ;
  assign n1734 = ~n1731 & ~n1732 ;
  assign n1735 = n1733 & n1734 ;
  assign n1736 = n273 & ~n1735 ;
  assign n1753 = ~n1728 & ~n1736 ;
  assign n1737 = n136 & ~n496 ;
  assign n1738 = n147 & ~n484 ;
  assign n1741 = ~n1737 & ~n1738 ;
  assign n1739 = n158 & ~n386 ;
  assign n1740 = n169 & ~n376 ;
  assign n1742 = ~n1739 & ~n1740 ;
  assign n1743 = n1741 & n1742 ;
  assign n1744 = n228 & ~n1743 ;
  assign n1745 = n136 & ~n406 ;
  assign n1746 = n147 & ~n396 ;
  assign n1749 = ~n1745 & ~n1746 ;
  assign n1747 = n158 & ~n342 ;
  assign n1748 = n169 & ~n332 ;
  assign n1750 = ~n1747 & ~n1748 ;
  assign n1751 = n1749 & n1750 ;
  assign n1752 = n183 & ~n1751 ;
  assign n1754 = ~n1744 & ~n1752 ;
  assign n1755 = n1753 & n1754 ;
  assign n1756 = \shift[6]  & ~n1755 ;
  assign n1757 = ~n1720 & ~n1756 ;
  assign n1758 = n136 & ~n605 ;
  assign n1759 = n147 & ~n593 ;
  assign n1762 = ~n1758 & ~n1759 ;
  assign n1760 = n158 & ~n529 ;
  assign n1761 = n169 & ~n517 ;
  assign n1763 = ~n1760 & ~n1761 ;
  assign n1764 = n1762 & n1763 ;
  assign n1765 = n183 & ~n1764 ;
  assign n1766 = n136 & ~n709 ;
  assign n1767 = n147 & ~n697 ;
  assign n1770 = ~n1766 & ~n1767 ;
  assign n1768 = n158 & ~n581 ;
  assign n1769 = n169 & ~n569 ;
  assign n1771 = ~n1768 & ~n1769 ;
  assign n1772 = n1770 & n1771 ;
  assign n1773 = n228 & ~n1772 ;
  assign n1790 = ~n1765 & ~n1773 ;
  assign n1774 = n136 & ~n817 ;
  assign n1775 = n147 & ~n805 ;
  assign n1778 = ~n1774 & ~n1775 ;
  assign n1776 = n158 & ~n633 ;
  assign n1777 = n169 & ~n621 ;
  assign n1779 = ~n1776 & ~n1777 ;
  assign n1780 = n1778 & n1779 ;
  assign n1781 = n273 & ~n1780 ;
  assign n1782 = n136 & ~n657 ;
  assign n1783 = n147 & ~n645 ;
  assign n1786 = ~n1782 & ~n1783 ;
  assign n1784 = n158 & ~n685 ;
  assign n1785 = n169 & ~n673 ;
  assign n1787 = ~n1784 & ~n1785 ;
  assign n1788 = n1786 & n1787 ;
  assign n1789 = n318 & ~n1788 ;
  assign n1791 = ~n1781 & ~n1789 ;
  assign n1792 = n1790 & n1791 ;
  assign n1793 = ~\shift[6]  & ~n1792 ;
  assign n1794 = n136 & ~n765 ;
  assign n1795 = n147 & ~n753 ;
  assign n1798 = ~n1794 & ~n1795 ;
  assign n1796 = n158 & ~n843 ;
  assign n1797 = n169 & ~n833 ;
  assign n1799 = ~n1796 & ~n1797 ;
  assign n1800 = n1798 & n1799 ;
  assign n1801 = n318 & ~n1800 ;
  assign n1802 = n136 & ~n553 ;
  assign n1803 = n147 & ~n541 ;
  assign n1806 = ~n1802 & ~n1803 ;
  assign n1804 = n158 & ~n741 ;
  assign n1805 = n169 & ~n729 ;
  assign n1807 = ~n1804 & ~n1805 ;
  assign n1808 = n1806 & n1807 ;
  assign n1809 = n273 & ~n1808 ;
  assign n1826 = ~n1801 & ~n1809 ;
  assign n1810 = n136 & ~n865 ;
  assign n1811 = n147 & ~n855 ;
  assign n1814 = ~n1810 & ~n1811 ;
  assign n1812 = n158 & ~n893 ;
  assign n1813 = n169 & ~n881 ;
  assign n1815 = ~n1812 & ~n1813 ;
  assign n1816 = n1814 & n1815 ;
  assign n1817 = n228 & ~n1816 ;
  assign n1818 = n136 & ~n917 ;
  assign n1819 = n147 & ~n905 ;
  assign n1822 = ~n1818 & ~n1819 ;
  assign n1820 = n158 & ~n793 ;
  assign n1821 = n169 & ~n781 ;
  assign n1823 = ~n1820 & ~n1821 ;
  assign n1824 = n1822 & n1823 ;
  assign n1825 = n183 & ~n1824 ;
  assign n1827 = ~n1817 & ~n1825 ;
  assign n1828 = n1826 & n1827 ;
  assign n1829 = \shift[6]  & ~n1828 ;
  assign n1830 = ~n1793 & ~n1829 ;
  assign n1831 = n136 & ~n962 ;
  assign n1832 = n147 & ~n958 ;
  assign n1835 = ~n1831 & ~n1832 ;
  assign n1833 = n158 & ~n934 ;
  assign n1834 = n169 & ~n930 ;
  assign n1836 = ~n1833 & ~n1834 ;
  assign n1837 = n1835 & n1836 ;
  assign n1838 = n183 & ~n1837 ;
  assign n1839 = n136 & ~n1002 ;
  assign n1840 = n147 & ~n998 ;
  assign n1843 = ~n1839 & ~n1840 ;
  assign n1841 = n158 & ~n954 ;
  assign n1842 = n169 & ~n950 ;
  assign n1844 = ~n1841 & ~n1842 ;
  assign n1845 = n1843 & n1844 ;
  assign n1846 = n228 & ~n1845 ;
  assign n1863 = ~n1838 & ~n1846 ;
  assign n1847 = n136 & ~n1046 ;
  assign n1848 = n147 & ~n1042 ;
  assign n1851 = ~n1847 & ~n1848 ;
  assign n1849 = n158 & ~n974 ;
  assign n1850 = n169 & ~n970 ;
  assign n1852 = ~n1849 & ~n1850 ;
  assign n1853 = n1851 & n1852 ;
  assign n1854 = n273 & ~n1853 ;
  assign n1855 = n136 & ~n982 ;
  assign n1856 = n147 & ~n978 ;
  assign n1859 = ~n1855 & ~n1856 ;
  assign n1857 = n158 & ~n994 ;
  assign n1858 = n169 & ~n990 ;
  assign n1860 = ~n1857 & ~n1858 ;
  assign n1861 = n1859 & n1860 ;
  assign n1862 = n318 & ~n1861 ;
  assign n1864 = ~n1854 & ~n1862 ;
  assign n1865 = n1863 & n1864 ;
  assign n1866 = ~\shift[6]  & ~n1865 ;
  assign n1867 = n136 & ~n1026 ;
  assign n1868 = n147 & ~n1022 ;
  assign n1871 = ~n1867 & ~n1868 ;
  assign n1869 = n158 & ~n1058 ;
  assign n1870 = n169 & ~n1054 ;
  assign n1872 = ~n1869 & ~n1870 ;
  assign n1873 = n1871 & n1872 ;
  assign n1874 = n318 & ~n1873 ;
  assign n1875 = n136 & ~n942 ;
  assign n1876 = n147 & ~n938 ;
  assign n1879 = ~n1875 & ~n1876 ;
  assign n1877 = n158 & ~n1018 ;
  assign n1878 = n169 & ~n1014 ;
  assign n1880 = ~n1877 & ~n1878 ;
  assign n1881 = n1879 & n1880 ;
  assign n1882 = n273 & ~n1881 ;
  assign n1899 = ~n1874 & ~n1882 ;
  assign n1883 = n136 & ~n1068 ;
  assign n1884 = n147 & ~n1063 ;
  assign n1887 = ~n1883 & ~n1884 ;
  assign n1885 = n158 & ~n1080 ;
  assign n1886 = n169 & ~n1076 ;
  assign n1888 = ~n1885 & ~n1886 ;
  assign n1889 = n1887 & n1888 ;
  assign n1890 = n228 & ~n1889 ;
  assign n1891 = n136 & ~n1088 ;
  assign n1892 = n147 & ~n1084 ;
  assign n1895 = ~n1891 & ~n1892 ;
  assign n1893 = n158 & ~n1038 ;
  assign n1894 = n169 & ~n1034 ;
  assign n1896 = ~n1893 & ~n1894 ;
  assign n1897 = n1895 & n1896 ;
  assign n1898 = n183 & ~n1897 ;
  assign n1900 = ~n1890 & ~n1898 ;
  assign n1901 = n1899 & n1900 ;
  assign n1902 = \shift[6]  & ~n1901 ;
  assign n1903 = ~n1866 & ~n1902 ;
  assign n1904 = n136 & ~n1165 ;
  assign n1905 = n147 & ~n1157 ;
  assign n1908 = ~n1904 & ~n1905 ;
  assign n1906 = n158 & ~n1221 ;
  assign n1907 = n169 & ~n1213 ;
  assign n1909 = ~n1906 & ~n1907 ;
  assign n1910 = n1908 & n1909 ;
  assign n1911 = n183 & ~n1910 ;
  assign n1912 = n136 & ~n1129 ;
  assign n1913 = n147 & ~n1121 ;
  assign n1916 = ~n1912 & ~n1913 ;
  assign n1914 = n158 & ~n1149 ;
  assign n1915 = n169 & ~n1141 ;
  assign n1917 = ~n1914 & ~n1915 ;
  assign n1918 = n1916 & n1917 ;
  assign n1919 = n228 & ~n1918 ;
  assign n1936 = ~n1911 & ~n1919 ;
  assign n1920 = n136 & ~n1346 ;
  assign n1921 = n147 & ~n1338 ;
  assign n1924 = ~n1920 & ~n1921 ;
  assign n1922 = n158 & ~n1185 ;
  assign n1923 = n169 & ~n1177 ;
  assign n1925 = ~n1922 & ~n1923 ;
  assign n1926 = n1924 & n1925 ;
  assign n1927 = n273 & ~n1926 ;
  assign n1928 = n136 & ~n1201 ;
  assign n1929 = n147 & ~n1193 ;
  assign n1932 = ~n1928 & ~n1929 ;
  assign n1930 = n158 & ~n1113 ;
  assign n1931 = n169 & ~n1105 ;
  assign n1933 = ~n1930 & ~n1931 ;
  assign n1934 = n1932 & n1933 ;
  assign n1935 = n318 & ~n1934 ;
  assign n1937 = ~n1927 & ~n1935 ;
  assign n1938 = n1936 & n1937 ;
  assign n1939 = ~\shift[6]  & ~n1938 ;
  assign n1940 = n136 & ~n1277 ;
  assign n1941 = n169 & ~n1289 ;
  assign n1944 = ~n1940 & ~n1941 ;
  assign n1942 = n158 & ~n1294 ;
  assign n1943 = n147 & ~n1269 ;
  assign n1945 = ~n1942 & ~n1943 ;
  assign n1946 = n1944 & n1945 ;
  assign n1947 = n318 & ~n1946 ;
  assign n1948 = n136 & ~n1237 ;
  assign n1949 = n147 & ~n1229 ;
  assign n1952 = ~n1948 & ~n1949 ;
  assign n1950 = n158 & ~n1261 ;
  assign n1951 = n169 & ~n1253 ;
  assign n1953 = ~n1950 & ~n1951 ;
  assign n1954 = n1952 & n1953 ;
  assign n1955 = n273 & ~n1954 ;
  assign n1972 = ~n1947 & ~n1955 ;
  assign n1956 = n136 & ~n1310 ;
  assign n1957 = n147 & ~n1302 ;
  assign n1960 = ~n1956 & ~n1957 ;
  assign n1958 = n158 & ~n1366 ;
  assign n1959 = n169 & ~n1358 ;
  assign n1961 = ~n1958 & ~n1959 ;
  assign n1962 = n1960 & n1961 ;
  assign n1963 = n228 & ~n1962 ;
  assign n1964 = n136 & ~n1382 ;
  assign n1965 = n147 & ~n1374 ;
  assign n1968 = ~n1964 & ~n1965 ;
  assign n1966 = n158 & ~n1330 ;
  assign n1967 = n169 & ~n1322 ;
  assign n1969 = ~n1966 & ~n1967 ;
  assign n1970 = n1968 & n1969 ;
  assign n1971 = n183 & ~n1970 ;
  assign n1973 = ~n1963 & ~n1971 ;
  assign n1974 = n1972 & n1973 ;
  assign n1975 = \shift[6]  & ~n1974 ;
  assign n1976 = ~n1939 & ~n1975 ;
  assign n1977 = n136 & ~n203 ;
  assign n1978 = n147 & ~n223 ;
  assign n1981 = ~n1977 & ~n1978 ;
  assign n1979 = ~n145 & n158 ;
  assign n1980 = n169 & ~n213 ;
  assign n1982 = ~n1979 & ~n1980 ;
  assign n1983 = n1981 & n1982 ;
  assign n1984 = n183 & ~n1983 ;
  assign n1985 = n136 & ~n293 ;
  assign n1986 = n147 & ~n313 ;
  assign n1989 = ~n1985 & ~n1986 ;
  assign n1987 = n158 & ~n193 ;
  assign n1988 = n169 & ~n303 ;
  assign n1990 = ~n1987 & ~n1988 ;
  assign n1991 = n1989 & n1990 ;
  assign n1992 = n228 & ~n1991 ;
  assign n2009 = ~n1984 & ~n1992 ;
  assign n1993 = n136 & ~n342 ;
  assign n1994 = n147 & ~n362 ;
  assign n1997 = ~n1993 & ~n1994 ;
  assign n1995 = n158 & ~n238 ;
  assign n1996 = n169 & ~n352 ;
  assign n1998 = ~n1995 & ~n1996 ;
  assign n1999 = n1997 & n1998 ;
  assign n2000 = n273 & ~n1999 ;
  assign n2001 = n136 & ~n248 ;
  assign n2002 = n147 & ~n268 ;
  assign n2005 = ~n2001 & ~n2002 ;
  assign n2003 = n158 & ~n283 ;
  assign n2004 = n169 & ~n258 ;
  assign n2006 = ~n2003 & ~n2004 ;
  assign n2007 = n2005 & n2006 ;
  assign n2008 = n318 & ~n2007 ;
  assign n2010 = ~n2000 & ~n2008 ;
  assign n2011 = n2009 & n2010 ;
  assign n2012 = ~\shift[6]  & ~n2011 ;
  assign n2013 = n136 & ~n430 ;
  assign n2014 = n147 & ~n450 ;
  assign n2017 = ~n2013 & ~n2014 ;
  assign n2015 = n158 & ~n464 ;
  assign n2016 = n169 & ~n440 ;
  assign n2018 = ~n2015 & ~n2016 ;
  assign n2019 = n2017 & n2018 ;
  assign n2020 = n318 & ~n2019 ;
  assign n2021 = n136 & ~n156 ;
  assign n2022 = n147 & ~n178 ;
  assign n2025 = ~n2021 & ~n2022 ;
  assign n2023 = n158 & ~n420 ;
  assign n2024 = ~n167 & n169 ;
  assign n2026 = ~n2023 & ~n2024 ;
  assign n2027 = n2025 & n2026 ;
  assign n2028 = n273 & ~n2027 ;
  assign n2045 = ~n2020 & ~n2028 ;
  assign n2029 = n136 & ~n474 ;
  assign n2030 = n147 & ~n496 ;
  assign n2033 = ~n2029 & ~n2030 ;
  assign n2031 = n158 & ~n376 ;
  assign n2032 = n169 & ~n484 ;
  assign n2034 = ~n2031 & ~n2032 ;
  assign n2035 = n2033 & n2034 ;
  assign n2036 = n228 & ~n2035 ;
  assign n2037 = n136 & ~n386 ;
  assign n2038 = n147 & ~n406 ;
  assign n2041 = ~n2037 & ~n2038 ;
  assign n2039 = n158 & ~n332 ;
  assign n2040 = n169 & ~n396 ;
  assign n2042 = ~n2039 & ~n2040 ;
  assign n2043 = n2041 & n2042 ;
  assign n2044 = n183 & ~n2043 ;
  assign n2046 = ~n2036 & ~n2044 ;
  assign n2047 = n2045 & n2046 ;
  assign n2048 = \shift[6]  & ~n2047 ;
  assign n2049 = ~n2012 & ~n2048 ;
  assign n2050 = n136 & ~n581 ;
  assign n2051 = n147 & ~n605 ;
  assign n2054 = ~n2050 & ~n2051 ;
  assign n2052 = n158 & ~n517 ;
  assign n2053 = n169 & ~n593 ;
  assign n2055 = ~n2052 & ~n2053 ;
  assign n2056 = n2054 & n2055 ;
  assign n2057 = n183 & ~n2056 ;
  assign n2058 = n136 & ~n685 ;
  assign n2059 = n147 & ~n709 ;
  assign n2062 = ~n2058 & ~n2059 ;
  assign n2060 = n158 & ~n569 ;
  assign n2061 = n169 & ~n697 ;
  assign n2063 = ~n2060 & ~n2061 ;
  assign n2064 = n2062 & n2063 ;
  assign n2065 = n228 & ~n2064 ;
  assign n2082 = ~n2057 & ~n2065 ;
  assign n2066 = n136 & ~n793 ;
  assign n2067 = n147 & ~n817 ;
  assign n2070 = ~n2066 & ~n2067 ;
  assign n2068 = n158 & ~n621 ;
  assign n2069 = n169 & ~n805 ;
  assign n2071 = ~n2068 & ~n2069 ;
  assign n2072 = n2070 & n2071 ;
  assign n2073 = n273 & ~n2072 ;
  assign n2074 = n136 & ~n633 ;
  assign n2075 = n147 & ~n657 ;
  assign n2078 = ~n2074 & ~n2075 ;
  assign n2076 = n158 & ~n673 ;
  assign n2077 = n169 & ~n645 ;
  assign n2079 = ~n2076 & ~n2077 ;
  assign n2080 = n2078 & n2079 ;
  assign n2081 = n318 & ~n2080 ;
  assign n2083 = ~n2073 & ~n2081 ;
  assign n2084 = n2082 & n2083 ;
  assign n2085 = ~\shift[6]  & ~n2084 ;
  assign n2086 = n136 & ~n741 ;
  assign n2087 = n147 & ~n765 ;
  assign n2090 = ~n2086 & ~n2087 ;
  assign n2088 = n158 & ~n833 ;
  assign n2089 = n169 & ~n753 ;
  assign n2091 = ~n2088 & ~n2089 ;
  assign n2092 = n2090 & n2091 ;
  assign n2093 = n318 & ~n2092 ;
  assign n2094 = n136 & ~n529 ;
  assign n2095 = n147 & ~n553 ;
  assign n2098 = ~n2094 & ~n2095 ;
  assign n2096 = n158 & ~n729 ;
  assign n2097 = n169 & ~n541 ;
  assign n2099 = ~n2096 & ~n2097 ;
  assign n2100 = n2098 & n2099 ;
  assign n2101 = n273 & ~n2100 ;
  assign n2118 = ~n2093 & ~n2101 ;
  assign n2102 = n136 & ~n843 ;
  assign n2103 = n147 & ~n865 ;
  assign n2106 = ~n2102 & ~n2103 ;
  assign n2104 = n158 & ~n881 ;
  assign n2105 = n169 & ~n855 ;
  assign n2107 = ~n2104 & ~n2105 ;
  assign n2108 = n2106 & n2107 ;
  assign n2109 = n228 & ~n2108 ;
  assign n2110 = n136 & ~n893 ;
  assign n2111 = n147 & ~n917 ;
  assign n2114 = ~n2110 & ~n2111 ;
  assign n2112 = n158 & ~n781 ;
  assign n2113 = n169 & ~n905 ;
  assign n2115 = ~n2112 & ~n2113 ;
  assign n2116 = n2114 & n2115 ;
  assign n2117 = n183 & ~n2116 ;
  assign n2119 = ~n2109 & ~n2117 ;
  assign n2120 = n2118 & n2119 ;
  assign n2121 = \shift[6]  & ~n2120 ;
  assign n2122 = ~n2085 & ~n2121 ;
  assign n2123 = n136 & ~n954 ;
  assign n2124 = n147 & ~n962 ;
  assign n2127 = ~n2123 & ~n2124 ;
  assign n2125 = n158 & ~n930 ;
  assign n2126 = n169 & ~n958 ;
  assign n2128 = ~n2125 & ~n2126 ;
  assign n2129 = n2127 & n2128 ;
  assign n2130 = n183 & ~n2129 ;
  assign n2131 = n136 & ~n994 ;
  assign n2132 = n147 & ~n1002 ;
  assign n2135 = ~n2131 & ~n2132 ;
  assign n2133 = n158 & ~n950 ;
  assign n2134 = n169 & ~n998 ;
  assign n2136 = ~n2133 & ~n2134 ;
  assign n2137 = n2135 & n2136 ;
  assign n2138 = n228 & ~n2137 ;
  assign n2155 = ~n2130 & ~n2138 ;
  assign n2139 = n136 & ~n1038 ;
  assign n2140 = n147 & ~n1046 ;
  assign n2143 = ~n2139 & ~n2140 ;
  assign n2141 = n158 & ~n970 ;
  assign n2142 = n169 & ~n1042 ;
  assign n2144 = ~n2141 & ~n2142 ;
  assign n2145 = n2143 & n2144 ;
  assign n2146 = n273 & ~n2145 ;
  assign n2147 = n136 & ~n974 ;
  assign n2148 = n147 & ~n982 ;
  assign n2151 = ~n2147 & ~n2148 ;
  assign n2149 = n158 & ~n990 ;
  assign n2150 = n169 & ~n978 ;
  assign n2152 = ~n2149 & ~n2150 ;
  assign n2153 = n2151 & n2152 ;
  assign n2154 = n318 & ~n2153 ;
  assign n2156 = ~n2146 & ~n2154 ;
  assign n2157 = n2155 & n2156 ;
  assign n2158 = ~\shift[6]  & ~n2157 ;
  assign n2159 = n136 & ~n1018 ;
  assign n2160 = n147 & ~n1026 ;
  assign n2163 = ~n2159 & ~n2160 ;
  assign n2161 = n158 & ~n1054 ;
  assign n2162 = n169 & ~n1022 ;
  assign n2164 = ~n2161 & ~n2162 ;
  assign n2165 = n2163 & n2164 ;
  assign n2166 = n318 & ~n2165 ;
  assign n2167 = n136 & ~n934 ;
  assign n2168 = n147 & ~n942 ;
  assign n2171 = ~n2167 & ~n2168 ;
  assign n2169 = n158 & ~n1014 ;
  assign n2170 = n169 & ~n938 ;
  assign n2172 = ~n2169 & ~n2170 ;
  assign n2173 = n2171 & n2172 ;
  assign n2174 = n273 & ~n2173 ;
  assign n2191 = ~n2166 & ~n2174 ;
  assign n2175 = n136 & ~n1058 ;
  assign n2176 = n147 & ~n1068 ;
  assign n2179 = ~n2175 & ~n2176 ;
  assign n2177 = n158 & ~n1076 ;
  assign n2178 = n169 & ~n1063 ;
  assign n2180 = ~n2177 & ~n2178 ;
  assign n2181 = n2179 & n2180 ;
  assign n2182 = n228 & ~n2181 ;
  assign n2183 = n136 & ~n1080 ;
  assign n2184 = n147 & ~n1088 ;
  assign n2187 = ~n2183 & ~n2184 ;
  assign n2185 = n158 & ~n1034 ;
  assign n2186 = n169 & ~n1084 ;
  assign n2188 = ~n2185 & ~n2186 ;
  assign n2189 = n2187 & n2188 ;
  assign n2190 = n183 & ~n2189 ;
  assign n2192 = ~n2182 & ~n2190 ;
  assign n2193 = n2191 & n2192 ;
  assign n2194 = \shift[6]  & ~n2193 ;
  assign n2195 = ~n2158 & ~n2194 ;
  assign n2196 = n136 & ~n1149 ;
  assign n2197 = n147 & ~n1165 ;
  assign n2200 = ~n2196 & ~n2197 ;
  assign n2198 = n158 & ~n1213 ;
  assign n2199 = n169 & ~n1157 ;
  assign n2201 = ~n2198 & ~n2199 ;
  assign n2202 = n2200 & n2201 ;
  assign n2203 = n183 & ~n2202 ;
  assign n2204 = n136 & ~n1113 ;
  assign n2205 = n147 & ~n1129 ;
  assign n2208 = ~n2204 & ~n2205 ;
  assign n2206 = n158 & ~n1141 ;
  assign n2207 = n169 & ~n1121 ;
  assign n2209 = ~n2206 & ~n2207 ;
  assign n2210 = n2208 & n2209 ;
  assign n2211 = n228 & ~n2210 ;
  assign n2228 = ~n2203 & ~n2211 ;
  assign n2212 = n136 & ~n1330 ;
  assign n2213 = n147 & ~n1346 ;
  assign n2216 = ~n2212 & ~n2213 ;
  assign n2214 = n158 & ~n1177 ;
  assign n2215 = n169 & ~n1338 ;
  assign n2217 = ~n2214 & ~n2215 ;
  assign n2218 = n2216 & n2217 ;
  assign n2219 = n273 & ~n2218 ;
  assign n2220 = n136 & ~n1185 ;
  assign n2221 = n147 & ~n1201 ;
  assign n2224 = ~n2220 & ~n2221 ;
  assign n2222 = n158 & ~n1105 ;
  assign n2223 = n169 & ~n1193 ;
  assign n2225 = ~n2222 & ~n2223 ;
  assign n2226 = n2224 & n2225 ;
  assign n2227 = n318 & ~n2226 ;
  assign n2229 = ~n2219 & ~n2227 ;
  assign n2230 = n2228 & n2229 ;
  assign n2231 = ~\shift[6]  & ~n2230 ;
  assign n2232 = n136 & ~n1261 ;
  assign n2233 = n147 & ~n1277 ;
  assign n2236 = ~n2232 & ~n2233 ;
  assign n2234 = n158 & ~n1289 ;
  assign n2235 = n169 & ~n1269 ;
  assign n2237 = ~n2234 & ~n2235 ;
  assign n2238 = n2236 & n2237 ;
  assign n2239 = n318 & ~n2238 ;
  assign n2240 = n136 & ~n1221 ;
  assign n2241 = n147 & ~n1237 ;
  assign n2244 = ~n2240 & ~n2241 ;
  assign n2242 = n158 & ~n1253 ;
  assign n2243 = n169 & ~n1229 ;
  assign n2245 = ~n2242 & ~n2243 ;
  assign n2246 = n2244 & n2245 ;
  assign n2247 = n273 & ~n2246 ;
  assign n2264 = ~n2239 & ~n2247 ;
  assign n2248 = n136 & ~n1294 ;
  assign n2249 = n147 & ~n1310 ;
  assign n2252 = ~n2248 & ~n2249 ;
  assign n2250 = n158 & ~n1358 ;
  assign n2251 = n169 & ~n1302 ;
  assign n2253 = ~n2250 & ~n2251 ;
  assign n2254 = n2252 & n2253 ;
  assign n2255 = n228 & ~n2254 ;
  assign n2256 = n136 & ~n1366 ;
  assign n2257 = n147 & ~n1382 ;
  assign n2260 = ~n2256 & ~n2257 ;
  assign n2258 = n158 & ~n1322 ;
  assign n2259 = n169 & ~n1374 ;
  assign n2261 = ~n2258 & ~n2259 ;
  assign n2262 = n2260 & n2261 ;
  assign n2263 = n183 & ~n2262 ;
  assign n2265 = ~n2255 & ~n2263 ;
  assign n2266 = n2264 & n2265 ;
  assign n2267 = \shift[6]  & ~n2266 ;
  assign n2268 = ~n2231 & ~n2267 ;
  assign n2269 = n183 & ~n227 ;
  assign n2270 = n228 & ~n317 ;
  assign n2273 = ~n2269 & ~n2270 ;
  assign n2271 = n273 & ~n366 ;
  assign n2272 = ~n272 & n318 ;
  assign n2274 = ~n2271 & ~n2272 ;
  assign n2275 = n2273 & n2274 ;
  assign n2276 = ~\shift[6]  & ~n2275 ;
  assign n2277 = ~n182 & n273 ;
  assign n2278 = n183 & ~n410 ;
  assign n2281 = ~n2277 & ~n2278 ;
  assign n2279 = n318 & ~n454 ;
  assign n2280 = n228 & ~n500 ;
  assign n2282 = ~n2279 & ~n2280 ;
  assign n2283 = n2281 & n2282 ;
  assign n2284 = \shift[6]  & ~n2283 ;
  assign n2285 = ~n2276 & ~n2284 ;
  assign n2286 = n183 & ~n609 ;
  assign n2287 = n228 & ~n713 ;
  assign n2290 = ~n2286 & ~n2287 ;
  assign n2288 = n273 & ~n821 ;
  assign n2289 = n318 & ~n661 ;
  assign n2291 = ~n2288 & ~n2289 ;
  assign n2292 = n2290 & n2291 ;
  assign n2293 = ~\shift[6]  & ~n2292 ;
  assign n2294 = n318 & ~n769 ;
  assign n2295 = n273 & ~n557 ;
  assign n2298 = ~n2294 & ~n2295 ;
  assign n2296 = n228 & ~n869 ;
  assign n2297 = n183 & ~n921 ;
  assign n2299 = ~n2296 & ~n2297 ;
  assign n2300 = n2298 & n2299 ;
  assign n2301 = \shift[6]  & ~n2300 ;
  assign n2302 = ~n2293 & ~n2301 ;
  assign n2303 = n183 & ~n966 ;
  assign n2304 = n228 & ~n1006 ;
  assign n2307 = ~n2303 & ~n2304 ;
  assign n2305 = n273 & ~n1050 ;
  assign n2306 = n318 & ~n986 ;
  assign n2308 = ~n2305 & ~n2306 ;
  assign n2309 = n2307 & n2308 ;
  assign n2310 = ~\shift[6]  & ~n2309 ;
  assign n2311 = n318 & ~n1030 ;
  assign n2312 = n273 & ~n946 ;
  assign n2315 = ~n2311 & ~n2312 ;
  assign n2313 = n228 & ~n1072 ;
  assign n2314 = n183 & ~n1092 ;
  assign n2316 = ~n2313 & ~n2314 ;
  assign n2317 = n2315 & n2316 ;
  assign n2318 = \shift[6]  & ~n2317 ;
  assign n2319 = ~n2310 & ~n2318 ;
  assign n2320 = n228 & ~n1133 ;
  assign n2321 = n183 & ~n1169 ;
  assign n2324 = ~n2320 & ~n2321 ;
  assign n2322 = n318 & ~n1205 ;
  assign n2323 = n273 & ~n1350 ;
  assign n2325 = ~n2322 & ~n2323 ;
  assign n2326 = n2324 & n2325 ;
  assign n2327 = ~\shift[6]  & ~n2326 ;
  assign n2328 = n318 & ~n1281 ;
  assign n2329 = n273 & ~n1241 ;
  assign n2332 = ~n2328 & ~n2329 ;
  assign n2330 = n183 & ~n1386 ;
  assign n2331 = n228 & ~n1314 ;
  assign n2333 = ~n2330 & ~n2331 ;
  assign n2334 = n2332 & n2333 ;
  assign n2335 = \shift[6]  & ~n2334 ;
  assign n2336 = ~n2327 & ~n2335 ;
  assign n2337 = n183 & ~n1407 ;
  assign n2338 = n228 & ~n1423 ;
  assign n2341 = ~n2337 & ~n2338 ;
  assign n2339 = n273 & ~n1459 ;
  assign n2340 = n318 & ~n1415 ;
  assign n2342 = ~n2339 & ~n2340 ;
  assign n2343 = n2341 & n2342 ;
  assign n2344 = ~\shift[6]  & ~n2343 ;
  assign n2345 = n273 & ~n1399 ;
  assign n2346 = n228 & ~n1435 ;
  assign n2349 = ~n2345 & ~n2346 ;
  assign n2347 = n183 & ~n1451 ;
  assign n2348 = n318 & ~n1443 ;
  assign n2350 = ~n2347 & ~n2348 ;
  assign n2351 = n2349 & n2350 ;
  assign n2352 = \shift[6]  & ~n2351 ;
  assign n2353 = ~n2344 & ~n2352 ;
  assign n2354 = n183 & ~n1480 ;
  assign n2355 = n228 & ~n1496 ;
  assign n2358 = ~n2354 & ~n2355 ;
  assign n2356 = n273 & ~n1532 ;
  assign n2357 = n318 & ~n1488 ;
  assign n2359 = ~n2356 & ~n2357 ;
  assign n2360 = n2358 & n2359 ;
  assign n2361 = ~\shift[6]  & ~n2360 ;
  assign n2362 = n273 & ~n1472 ;
  assign n2363 = n228 & ~n1508 ;
  assign n2366 = ~n2362 & ~n2363 ;
  assign n2364 = n183 & ~n1524 ;
  assign n2365 = n318 & ~n1516 ;
  assign n2367 = ~n2364 & ~n2365 ;
  assign n2368 = n2366 & n2367 ;
  assign n2369 = \shift[6]  & ~n2368 ;
  assign n2370 = ~n2361 & ~n2369 ;
  assign n2371 = n183 & ~n1553 ;
  assign n2372 = n228 & ~n1569 ;
  assign n2375 = ~n2371 & ~n2372 ;
  assign n2373 = n273 & ~n1605 ;
  assign n2374 = n318 & ~n1561 ;
  assign n2376 = ~n2373 & ~n2374 ;
  assign n2377 = n2375 & n2376 ;
  assign n2378 = ~\shift[6]  & ~n2377 ;
  assign n2379 = n273 & ~n1545 ;
  assign n2380 = n228 & ~n1581 ;
  assign n2383 = ~n2379 & ~n2380 ;
  assign n2381 = n183 & ~n1597 ;
  assign n2382 = n318 & ~n1589 ;
  assign n2384 = ~n2381 & ~n2382 ;
  assign n2385 = n2383 & n2384 ;
  assign n2386 = \shift[6]  & ~n2385 ;
  assign n2387 = ~n2378 & ~n2386 ;
  assign n2388 = n183 & ~n1626 ;
  assign n2389 = n273 & ~n1678 ;
  assign n2392 = ~n2388 & ~n2389 ;
  assign n2390 = n318 & ~n1634 ;
  assign n2391 = n228 & ~n1642 ;
  assign n2393 = ~n2390 & ~n2391 ;
  assign n2394 = n2392 & n2393 ;
  assign n2395 = ~\shift[6]  & ~n2394 ;
  assign n2396 = n228 & ~n1654 ;
  assign n2397 = n318 & ~n1662 ;
  assign n2400 = ~n2396 & ~n2397 ;
  assign n2398 = n183 & ~n1670 ;
  assign n2399 = n273 & ~n1618 ;
  assign n2401 = ~n2398 & ~n2399 ;
  assign n2402 = n2400 & n2401 ;
  assign n2403 = \shift[6]  & ~n2402 ;
  assign n2404 = ~n2395 & ~n2403 ;
  assign n2405 = n183 & ~n1699 ;
  assign n2406 = n273 & ~n1751 ;
  assign n2409 = ~n2405 & ~n2406 ;
  assign n2407 = n318 & ~n1707 ;
  assign n2408 = n228 & ~n1715 ;
  assign n2410 = ~n2407 & ~n2408 ;
  assign n2411 = n2409 & n2410 ;
  assign n2412 = ~\shift[6]  & ~n2411 ;
  assign n2413 = n228 & ~n1727 ;
  assign n2414 = n318 & ~n1735 ;
  assign n2417 = ~n2413 & ~n2414 ;
  assign n2415 = n183 & ~n1743 ;
  assign n2416 = n273 & ~n1691 ;
  assign n2418 = ~n2415 & ~n2416 ;
  assign n2419 = n2417 & n2418 ;
  assign n2420 = \shift[6]  & ~n2419 ;
  assign n2421 = ~n2412 & ~n2420 ;
  assign n2422 = n183 & ~n1772 ;
  assign n2423 = n273 & ~n1824 ;
  assign n2426 = ~n2422 & ~n2423 ;
  assign n2424 = n318 & ~n1780 ;
  assign n2425 = n228 & ~n1788 ;
  assign n2427 = ~n2424 & ~n2425 ;
  assign n2428 = n2426 & n2427 ;
  assign n2429 = ~\shift[6]  & ~n2428 ;
  assign n2430 = n228 & ~n1800 ;
  assign n2431 = n318 & ~n1808 ;
  assign n2434 = ~n2430 & ~n2431 ;
  assign n2432 = n183 & ~n1816 ;
  assign n2433 = n273 & ~n1764 ;
  assign n2435 = ~n2432 & ~n2433 ;
  assign n2436 = n2434 & n2435 ;
  assign n2437 = \shift[6]  & ~n2436 ;
  assign n2438 = ~n2429 & ~n2437 ;
  assign n2439 = n183 & ~n1845 ;
  assign n2440 = n228 & ~n1861 ;
  assign n2443 = ~n2439 & ~n2440 ;
  assign n2441 = n273 & ~n1897 ;
  assign n2442 = n318 & ~n1853 ;
  assign n2444 = ~n2441 & ~n2442 ;
  assign n2445 = n2443 & n2444 ;
  assign n2446 = ~\shift[6]  & ~n2445 ;
  assign n2447 = n228 & ~n1873 ;
  assign n2448 = n318 & ~n1881 ;
  assign n2451 = ~n2447 & ~n2448 ;
  assign n2449 = n183 & ~n1889 ;
  assign n2450 = n273 & ~n1837 ;
  assign n2452 = ~n2449 & ~n2450 ;
  assign n2453 = n2451 & n2452 ;
  assign n2454 = \shift[6]  & ~n2453 ;
  assign n2455 = ~n2446 & ~n2454 ;
  assign n2456 = n183 & ~n1918 ;
  assign n2457 = n228 & ~n1934 ;
  assign n2460 = ~n2456 & ~n2457 ;
  assign n2458 = n273 & ~n1970 ;
  assign n2459 = n318 & ~n1926 ;
  assign n2461 = ~n2458 & ~n2459 ;
  assign n2462 = n2460 & n2461 ;
  assign n2463 = ~\shift[6]  & ~n2462 ;
  assign n2464 = n228 & ~n1946 ;
  assign n2465 = n318 & ~n1954 ;
  assign n2468 = ~n2464 & ~n2465 ;
  assign n2466 = n183 & ~n1962 ;
  assign n2467 = n273 & ~n1910 ;
  assign n2469 = ~n2466 & ~n2467 ;
  assign n2470 = n2468 & n2469 ;
  assign n2471 = \shift[6]  & ~n2470 ;
  assign n2472 = ~n2463 & ~n2471 ;
  assign n2473 = n183 & ~n1991 ;
  assign n2474 = n228 & ~n2007 ;
  assign n2477 = ~n2473 & ~n2474 ;
  assign n2475 = n273 & ~n2043 ;
  assign n2476 = n318 & ~n1999 ;
  assign n2478 = ~n2475 & ~n2476 ;
  assign n2479 = n2477 & n2478 ;
  assign n2480 = ~\shift[6]  & ~n2479 ;
  assign n2481 = n228 & ~n2019 ;
  assign n2482 = n318 & ~n2027 ;
  assign n2485 = ~n2481 & ~n2482 ;
  assign n2483 = n183 & ~n2035 ;
  assign n2484 = n273 & ~n1983 ;
  assign n2486 = ~n2483 & ~n2484 ;
  assign n2487 = n2485 & n2486 ;
  assign n2488 = \shift[6]  & ~n2487 ;
  assign n2489 = ~n2480 & ~n2488 ;
  assign n2490 = n183 & ~n2064 ;
  assign n2491 = n228 & ~n2080 ;
  assign n2494 = ~n2490 & ~n2491 ;
  assign n2492 = n273 & ~n2116 ;
  assign n2493 = n318 & ~n2072 ;
  assign n2495 = ~n2492 & ~n2493 ;
  assign n2496 = n2494 & n2495 ;
  assign n2497 = ~\shift[6]  & ~n2496 ;
  assign n2498 = n228 & ~n2092 ;
  assign n2499 = n318 & ~n2100 ;
  assign n2502 = ~n2498 & ~n2499 ;
  assign n2500 = n183 & ~n2108 ;
  assign n2501 = n273 & ~n2056 ;
  assign n2503 = ~n2500 & ~n2501 ;
  assign n2504 = n2502 & n2503 ;
  assign n2505 = \shift[6]  & ~n2504 ;
  assign n2506 = ~n2497 & ~n2505 ;
  assign n2507 = n183 & ~n2137 ;
  assign n2508 = n228 & ~n2153 ;
  assign n2511 = ~n2507 & ~n2508 ;
  assign n2509 = n273 & ~n2189 ;
  assign n2510 = n318 & ~n2145 ;
  assign n2512 = ~n2509 & ~n2510 ;
  assign n2513 = n2511 & n2512 ;
  assign n2514 = ~\shift[6]  & ~n2513 ;
  assign n2515 = n228 & ~n2165 ;
  assign n2516 = n318 & ~n2173 ;
  assign n2519 = ~n2515 & ~n2516 ;
  assign n2517 = n183 & ~n2181 ;
  assign n2518 = n273 & ~n2129 ;
  assign n2520 = ~n2517 & ~n2518 ;
  assign n2521 = n2519 & n2520 ;
  assign n2522 = \shift[6]  & ~n2521 ;
  assign n2523 = ~n2514 & ~n2522 ;
  assign n2524 = n183 & ~n2210 ;
  assign n2525 = n228 & ~n2226 ;
  assign n2528 = ~n2524 & ~n2525 ;
  assign n2526 = n273 & ~n2262 ;
  assign n2527 = n318 & ~n2218 ;
  assign n2529 = ~n2526 & ~n2527 ;
  assign n2530 = n2528 & n2529 ;
  assign n2531 = ~\shift[6]  & ~n2530 ;
  assign n2532 = n228 & ~n2238 ;
  assign n2533 = n318 & ~n2246 ;
  assign n2536 = ~n2532 & ~n2533 ;
  assign n2534 = n183 & ~n2254 ;
  assign n2535 = n273 & ~n2202 ;
  assign n2537 = ~n2534 & ~n2535 ;
  assign n2538 = n2536 & n2537 ;
  assign n2539 = \shift[6]  & ~n2538 ;
  assign n2540 = ~n2531 & ~n2539 ;
  assign n2541 = n183 & ~n317 ;
  assign n2542 = n228 & ~n272 ;
  assign n2545 = ~n2541 & ~n2542 ;
  assign n2543 = n273 & ~n410 ;
  assign n2544 = n318 & ~n366 ;
  assign n2546 = ~n2543 & ~n2544 ;
  assign n2547 = n2545 & n2546 ;
  assign n2548 = ~\shift[6]  & ~n2547 ;
  assign n2549 = ~n182 & n318 ;
  assign n2550 = ~n227 & n273 ;
  assign n2553 = ~n2549 & ~n2550 ;
  assign n2551 = n228 & ~n454 ;
  assign n2552 = n183 & ~n500 ;
  assign n2554 = ~n2551 & ~n2552 ;
  assign n2555 = n2553 & n2554 ;
  assign n2556 = \shift[6]  & ~n2555 ;
  assign n2557 = ~n2548 & ~n2556 ;
  assign n2558 = n183 & ~n713 ;
  assign n2559 = n228 & ~n661 ;
  assign n2562 = ~n2558 & ~n2559 ;
  assign n2560 = n273 & ~n921 ;
  assign n2561 = n318 & ~n821 ;
  assign n2563 = ~n2560 & ~n2561 ;
  assign n2564 = n2562 & n2563 ;
  assign n2565 = ~\shift[6]  & ~n2564 ;
  assign n2566 = n228 & ~n769 ;
  assign n2567 = n318 & ~n557 ;
  assign n2570 = ~n2566 & ~n2567 ;
  assign n2568 = n183 & ~n869 ;
  assign n2569 = n273 & ~n609 ;
  assign n2571 = ~n2568 & ~n2569 ;
  assign n2572 = n2570 & n2571 ;
  assign n2573 = \shift[6]  & ~n2572 ;
  assign n2574 = ~n2565 & ~n2573 ;
  assign n2575 = n183 & ~n1006 ;
  assign n2576 = n228 & ~n986 ;
  assign n2579 = ~n2575 & ~n2576 ;
  assign n2577 = n273 & ~n1092 ;
  assign n2578 = n318 & ~n1050 ;
  assign n2580 = ~n2577 & ~n2578 ;
  assign n2581 = n2579 & n2580 ;
  assign n2582 = ~\shift[6]  & ~n2581 ;
  assign n2583 = n228 & ~n1030 ;
  assign n2584 = n318 & ~n946 ;
  assign n2587 = ~n2583 & ~n2584 ;
  assign n2585 = n183 & ~n1072 ;
  assign n2586 = n273 & ~n966 ;
  assign n2588 = ~n2585 & ~n2586 ;
  assign n2589 = n2587 & n2588 ;
  assign n2590 = \shift[6]  & ~n2589 ;
  assign n2591 = ~n2582 & ~n2590 ;
  assign n2592 = n183 & ~n1133 ;
  assign n2593 = n273 & ~n1386 ;
  assign n2596 = ~n2592 & ~n2593 ;
  assign n2594 = n228 & ~n1205 ;
  assign n2595 = n318 & ~n1350 ;
  assign n2597 = ~n2594 & ~n2595 ;
  assign n2598 = n2596 & n2597 ;
  assign n2599 = ~\shift[6]  & ~n2598 ;
  assign n2600 = n228 & ~n1281 ;
  assign n2601 = n273 & ~n1169 ;
  assign n2604 = ~n2600 & ~n2601 ;
  assign n2602 = n183 & ~n1314 ;
  assign n2603 = n318 & ~n1241 ;
  assign n2605 = ~n2602 & ~n2603 ;
  assign n2606 = n2604 & n2605 ;
  assign n2607 = \shift[6]  & ~n2606 ;
  assign n2608 = ~n2599 & ~n2607 ;
  assign n2609 = n183 & ~n1423 ;
  assign n2610 = n228 & ~n1415 ;
  assign n2613 = ~n2609 & ~n2610 ;
  assign n2611 = n273 & ~n1451 ;
  assign n2612 = n318 & ~n1459 ;
  assign n2614 = ~n2611 & ~n2612 ;
  assign n2615 = n2613 & n2614 ;
  assign n2616 = ~\shift[6]  & ~n2615 ;
  assign n2617 = n318 & ~n1399 ;
  assign n2618 = n273 & ~n1407 ;
  assign n2621 = ~n2617 & ~n2618 ;
  assign n2619 = n228 & ~n1443 ;
  assign n2620 = n183 & ~n1435 ;
  assign n2622 = ~n2619 & ~n2620 ;
  assign n2623 = n2621 & n2622 ;
  assign n2624 = \shift[6]  & ~n2623 ;
  assign n2625 = ~n2616 & ~n2624 ;
  assign n2626 = n183 & ~n1496 ;
  assign n2627 = n228 & ~n1488 ;
  assign n2630 = ~n2626 & ~n2627 ;
  assign n2628 = n273 & ~n1524 ;
  assign n2629 = n318 & ~n1532 ;
  assign n2631 = ~n2628 & ~n2629 ;
  assign n2632 = n2630 & n2631 ;
  assign n2633 = ~\shift[6]  & ~n2632 ;
  assign n2634 = n318 & ~n1472 ;
  assign n2635 = n273 & ~n1480 ;
  assign n2638 = ~n2634 & ~n2635 ;
  assign n2636 = n228 & ~n1516 ;
  assign n2637 = n183 & ~n1508 ;
  assign n2639 = ~n2636 & ~n2637 ;
  assign n2640 = n2638 & n2639 ;
  assign n2641 = \shift[6]  & ~n2640 ;
  assign n2642 = ~n2633 & ~n2641 ;
  assign n2643 = n183 & ~n1569 ;
  assign n2644 = n228 & ~n1561 ;
  assign n2647 = ~n2643 & ~n2644 ;
  assign n2645 = n273 & ~n1597 ;
  assign n2646 = n318 & ~n1605 ;
  assign n2648 = ~n2645 & ~n2646 ;
  assign n2649 = n2647 & n2648 ;
  assign n2650 = ~\shift[6]  & ~n2649 ;
  assign n2651 = n318 & ~n1545 ;
  assign n2652 = n273 & ~n1553 ;
  assign n2655 = ~n2651 & ~n2652 ;
  assign n2653 = n228 & ~n1589 ;
  assign n2654 = n183 & ~n1581 ;
  assign n2656 = ~n2653 & ~n2654 ;
  assign n2657 = n2655 & n2656 ;
  assign n2658 = \shift[6]  & ~n2657 ;
  assign n2659 = ~n2650 & ~n2658 ;
  assign n2660 = n318 & ~n1678 ;
  assign n2661 = n273 & ~n1670 ;
  assign n2664 = ~n2660 & ~n2661 ;
  assign n2662 = n228 & ~n1634 ;
  assign n2663 = n183 & ~n1642 ;
  assign n2665 = ~n2662 & ~n2663 ;
  assign n2666 = n2664 & n2665 ;
  assign n2667 = ~\shift[6]  & ~n2666 ;
  assign n2668 = n183 & ~n1654 ;
  assign n2669 = n228 & ~n1662 ;
  assign n2672 = ~n2668 & ~n2669 ;
  assign n2670 = n273 & ~n1626 ;
  assign n2671 = n318 & ~n1618 ;
  assign n2673 = ~n2670 & ~n2671 ;
  assign n2674 = n2672 & n2673 ;
  assign n2675 = \shift[6]  & ~n2674 ;
  assign n2676 = ~n2667 & ~n2675 ;
  assign n2677 = n318 & ~n1751 ;
  assign n2678 = n273 & ~n1743 ;
  assign n2681 = ~n2677 & ~n2678 ;
  assign n2679 = n228 & ~n1707 ;
  assign n2680 = n183 & ~n1715 ;
  assign n2682 = ~n2679 & ~n2680 ;
  assign n2683 = n2681 & n2682 ;
  assign n2684 = ~\shift[6]  & ~n2683 ;
  assign n2685 = n183 & ~n1727 ;
  assign n2686 = n228 & ~n1735 ;
  assign n2689 = ~n2685 & ~n2686 ;
  assign n2687 = n273 & ~n1699 ;
  assign n2688 = n318 & ~n1691 ;
  assign n2690 = ~n2687 & ~n2688 ;
  assign n2691 = n2689 & n2690 ;
  assign n2692 = \shift[6]  & ~n2691 ;
  assign n2693 = ~n2684 & ~n2692 ;
  assign n2694 = n318 & ~n1824 ;
  assign n2695 = n273 & ~n1816 ;
  assign n2698 = ~n2694 & ~n2695 ;
  assign n2696 = n228 & ~n1780 ;
  assign n2697 = n183 & ~n1788 ;
  assign n2699 = ~n2696 & ~n2697 ;
  assign n2700 = n2698 & n2699 ;
  assign n2701 = ~\shift[6]  & ~n2700 ;
  assign n2702 = n183 & ~n1800 ;
  assign n2703 = n228 & ~n1808 ;
  assign n2706 = ~n2702 & ~n2703 ;
  assign n2704 = n273 & ~n1772 ;
  assign n2705 = n318 & ~n1764 ;
  assign n2707 = ~n2704 & ~n2705 ;
  assign n2708 = n2706 & n2707 ;
  assign n2709 = \shift[6]  & ~n2708 ;
  assign n2710 = ~n2701 & ~n2709 ;
  assign n2711 = n183 & ~n1861 ;
  assign n2712 = n228 & ~n1853 ;
  assign n2715 = ~n2711 & ~n2712 ;
  assign n2713 = n273 & ~n1889 ;
  assign n2714 = n318 & ~n1897 ;
  assign n2716 = ~n2713 & ~n2714 ;
  assign n2717 = n2715 & n2716 ;
  assign n2718 = ~\shift[6]  & ~n2717 ;
  assign n2719 = n183 & ~n1873 ;
  assign n2720 = n228 & ~n1881 ;
  assign n2723 = ~n2719 & ~n2720 ;
  assign n2721 = n273 & ~n1845 ;
  assign n2722 = n318 & ~n1837 ;
  assign n2724 = ~n2721 & ~n2722 ;
  assign n2725 = n2723 & n2724 ;
  assign n2726 = \shift[6]  & ~n2725 ;
  assign n2727 = ~n2718 & ~n2726 ;
  assign n2728 = n183 & ~n1934 ;
  assign n2729 = n228 & ~n1926 ;
  assign n2732 = ~n2728 & ~n2729 ;
  assign n2730 = n273 & ~n1962 ;
  assign n2731 = n318 & ~n1970 ;
  assign n2733 = ~n2730 & ~n2731 ;
  assign n2734 = n2732 & n2733 ;
  assign n2735 = ~\shift[6]  & ~n2734 ;
  assign n2736 = n183 & ~n1946 ;
  assign n2737 = n228 & ~n1954 ;
  assign n2740 = ~n2736 & ~n2737 ;
  assign n2738 = n273 & ~n1918 ;
  assign n2739 = n318 & ~n1910 ;
  assign n2741 = ~n2738 & ~n2739 ;
  assign n2742 = n2740 & n2741 ;
  assign n2743 = \shift[6]  & ~n2742 ;
  assign n2744 = ~n2735 & ~n2743 ;
  assign n2745 = n183 & ~n2007 ;
  assign n2746 = n228 & ~n1999 ;
  assign n2749 = ~n2745 & ~n2746 ;
  assign n2747 = n273 & ~n2035 ;
  assign n2748 = n318 & ~n2043 ;
  assign n2750 = ~n2747 & ~n2748 ;
  assign n2751 = n2749 & n2750 ;
  assign n2752 = ~\shift[6]  & ~n2751 ;
  assign n2753 = n183 & ~n2019 ;
  assign n2754 = n228 & ~n2027 ;
  assign n2757 = ~n2753 & ~n2754 ;
  assign n2755 = n273 & ~n1991 ;
  assign n2756 = n318 & ~n1983 ;
  assign n2758 = ~n2755 & ~n2756 ;
  assign n2759 = n2757 & n2758 ;
  assign n2760 = \shift[6]  & ~n2759 ;
  assign n2761 = ~n2752 & ~n2760 ;
  assign n2762 = n183 & ~n2080 ;
  assign n2763 = n228 & ~n2072 ;
  assign n2766 = ~n2762 & ~n2763 ;
  assign n2764 = n273 & ~n2108 ;
  assign n2765 = n318 & ~n2116 ;
  assign n2767 = ~n2764 & ~n2765 ;
  assign n2768 = n2766 & n2767 ;
  assign n2769 = ~\shift[6]  & ~n2768 ;
  assign n2770 = n183 & ~n2092 ;
  assign n2771 = n228 & ~n2100 ;
  assign n2774 = ~n2770 & ~n2771 ;
  assign n2772 = n273 & ~n2064 ;
  assign n2773 = n318 & ~n2056 ;
  assign n2775 = ~n2772 & ~n2773 ;
  assign n2776 = n2774 & n2775 ;
  assign n2777 = \shift[6]  & ~n2776 ;
  assign n2778 = ~n2769 & ~n2777 ;
  assign n2779 = n183 & ~n2153 ;
  assign n2780 = n228 & ~n2145 ;
  assign n2783 = ~n2779 & ~n2780 ;
  assign n2781 = n273 & ~n2181 ;
  assign n2782 = n318 & ~n2189 ;
  assign n2784 = ~n2781 & ~n2782 ;
  assign n2785 = n2783 & n2784 ;
  assign n2786 = ~\shift[6]  & ~n2785 ;
  assign n2787 = n183 & ~n2165 ;
  assign n2788 = n228 & ~n2173 ;
  assign n2791 = ~n2787 & ~n2788 ;
  assign n2789 = n273 & ~n2137 ;
  assign n2790 = n318 & ~n2129 ;
  assign n2792 = ~n2789 & ~n2790 ;
  assign n2793 = n2791 & n2792 ;
  assign n2794 = \shift[6]  & ~n2793 ;
  assign n2795 = ~n2786 & ~n2794 ;
  assign n2796 = n183 & ~n2226 ;
  assign n2797 = n228 & ~n2218 ;
  assign n2800 = ~n2796 & ~n2797 ;
  assign n2798 = n273 & ~n2254 ;
  assign n2799 = n318 & ~n2262 ;
  assign n2801 = ~n2798 & ~n2799 ;
  assign n2802 = n2800 & n2801 ;
  assign n2803 = ~\shift[6]  & ~n2802 ;
  assign n2804 = n183 & ~n2238 ;
  assign n2805 = n228 & ~n2246 ;
  assign n2808 = ~n2804 & ~n2805 ;
  assign n2806 = n273 & ~n2210 ;
  assign n2807 = n318 & ~n2202 ;
  assign n2809 = ~n2806 & ~n2807 ;
  assign n2810 = n2808 & n2809 ;
  assign n2811 = \shift[6]  & ~n2810 ;
  assign n2812 = ~n2803 & ~n2811 ;
  assign n2813 = n183 & ~n272 ;
  assign n2814 = n228 & ~n366 ;
  assign n2817 = ~n2813 & ~n2814 ;
  assign n2815 = n273 & ~n500 ;
  assign n2816 = n318 & ~n410 ;
  assign n2818 = ~n2815 & ~n2816 ;
  assign n2819 = n2817 & n2818 ;
  assign n2820 = ~\shift[6]  & ~n2819 ;
  assign n2821 = ~n182 & n228 ;
  assign n2822 = ~n227 & n318 ;
  assign n2825 = ~n2821 & ~n2822 ;
  assign n2823 = n183 & ~n454 ;
  assign n2824 = n273 & ~n317 ;
  assign n2826 = ~n2823 & ~n2824 ;
  assign n2827 = n2825 & n2826 ;
  assign n2828 = \shift[6]  & ~n2827 ;
  assign n2829 = ~n2820 & ~n2828 ;
  assign n2830 = n183 & ~n661 ;
  assign n2831 = n228 & ~n821 ;
  assign n2834 = ~n2830 & ~n2831 ;
  assign n2832 = n273 & ~n869 ;
  assign n2833 = n318 & ~n921 ;
  assign n2835 = ~n2832 & ~n2833 ;
  assign n2836 = n2834 & n2835 ;
  assign n2837 = ~\shift[6]  & ~n2836 ;
  assign n2838 = n183 & ~n769 ;
  assign n2839 = n228 & ~n557 ;
  assign n2842 = ~n2838 & ~n2839 ;
  assign n2840 = n273 & ~n713 ;
  assign n2841 = n318 & ~n609 ;
  assign n2843 = ~n2840 & ~n2841 ;
  assign n2844 = n2842 & n2843 ;
  assign n2845 = \shift[6]  & ~n2844 ;
  assign n2846 = ~n2837 & ~n2845 ;
  assign n2847 = n183 & ~n986 ;
  assign n2848 = n228 & ~n1050 ;
  assign n2851 = ~n2847 & ~n2848 ;
  assign n2849 = n273 & ~n1072 ;
  assign n2850 = n318 & ~n1092 ;
  assign n2852 = ~n2849 & ~n2850 ;
  assign n2853 = n2851 & n2852 ;
  assign n2854 = ~\shift[6]  & ~n2853 ;
  assign n2855 = n183 & ~n1030 ;
  assign n2856 = n228 & ~n946 ;
  assign n2859 = ~n2855 & ~n2856 ;
  assign n2857 = n273 & ~n1006 ;
  assign n2858 = n318 & ~n966 ;
  assign n2860 = ~n2857 & ~n2858 ;
  assign n2861 = n2859 & n2860 ;
  assign n2862 = \shift[6]  & ~n2861 ;
  assign n2863 = ~n2854 & ~n2862 ;
  assign n2864 = n273 & ~n1314 ;
  assign n2865 = n318 & ~n1386 ;
  assign n2868 = ~n2864 & ~n2865 ;
  assign n2866 = n183 & ~n1205 ;
  assign n2867 = n228 & ~n1350 ;
  assign n2869 = ~n2866 & ~n2867 ;
  assign n2870 = n2868 & n2869 ;
  assign n2871 = ~\shift[6]  & ~n2870 ;
  assign n2872 = n183 & ~n1281 ;
  assign n2873 = n273 & ~n1133 ;
  assign n2876 = ~n2872 & ~n2873 ;
  assign n2874 = n228 & ~n1241 ;
  assign n2875 = n318 & ~n1169 ;
  assign n2877 = ~n2874 & ~n2875 ;
  assign n2878 = n2876 & n2877 ;
  assign n2879 = \shift[6]  & ~n2878 ;
  assign n2880 = ~n2871 & ~n2879 ;
  assign n2881 = n273 & ~n1435 ;
  assign n2882 = n183 & ~n1415 ;
  assign n2885 = ~n2881 & ~n2882 ;
  assign n2883 = n318 & ~n1451 ;
  assign n2884 = n228 & ~n1459 ;
  assign n2886 = ~n2883 & ~n2884 ;
  assign n2887 = n2885 & n2886 ;
  assign n2888 = ~\shift[6]  & ~n2887 ;
  assign n2889 = n228 & ~n1399 ;
  assign n2890 = n318 & ~n1407 ;
  assign n2893 = ~n2889 & ~n2890 ;
  assign n2891 = n273 & ~n1423 ;
  assign n2892 = n183 & ~n1443 ;
  assign n2894 = ~n2891 & ~n2892 ;
  assign n2895 = n2893 & n2894 ;
  assign n2896 = \shift[6]  & ~n2895 ;
  assign n2897 = ~n2888 & ~n2896 ;
  assign n2898 = n273 & ~n1508 ;
  assign n2899 = n183 & ~n1488 ;
  assign n2902 = ~n2898 & ~n2899 ;
  assign n2900 = n318 & ~n1524 ;
  assign n2901 = n228 & ~n1532 ;
  assign n2903 = ~n2900 & ~n2901 ;
  assign n2904 = n2902 & n2903 ;
  assign n2905 = ~\shift[6]  & ~n2904 ;
  assign n2906 = n228 & ~n1472 ;
  assign n2907 = n318 & ~n1480 ;
  assign n2910 = ~n2906 & ~n2907 ;
  assign n2908 = n273 & ~n1496 ;
  assign n2909 = n183 & ~n1516 ;
  assign n2911 = ~n2908 & ~n2909 ;
  assign n2912 = n2910 & n2911 ;
  assign n2913 = \shift[6]  & ~n2912 ;
  assign n2914 = ~n2905 & ~n2913 ;
  assign n2915 = n273 & ~n1581 ;
  assign n2916 = n183 & ~n1561 ;
  assign n2919 = ~n2915 & ~n2916 ;
  assign n2917 = n318 & ~n1597 ;
  assign n2918 = n228 & ~n1605 ;
  assign n2920 = ~n2917 & ~n2918 ;
  assign n2921 = n2919 & n2920 ;
  assign n2922 = ~\shift[6]  & ~n2921 ;
  assign n2923 = n228 & ~n1545 ;
  assign n2924 = n318 & ~n1553 ;
  assign n2927 = ~n2923 & ~n2924 ;
  assign n2925 = n273 & ~n1569 ;
  assign n2926 = n183 & ~n1589 ;
  assign n2928 = ~n2925 & ~n2926 ;
  assign n2929 = n2927 & n2928 ;
  assign n2930 = \shift[6]  & ~n2929 ;
  assign n2931 = ~n2922 & ~n2930 ;
  assign n2932 = n273 & ~n1654 ;
  assign n2933 = n228 & ~n1678 ;
  assign n2936 = ~n2932 & ~n2933 ;
  assign n2934 = n183 & ~n1634 ;
  assign n2935 = n318 & ~n1670 ;
  assign n2937 = ~n2934 & ~n2935 ;
  assign n2938 = n2936 & n2937 ;
  assign n2939 = ~\shift[6]  & ~n2938 ;
  assign n2940 = n183 & ~n1662 ;
  assign n2941 = n228 & ~n1618 ;
  assign n2944 = ~n2940 & ~n2941 ;
  assign n2942 = n273 & ~n1642 ;
  assign n2943 = n318 & ~n1626 ;
  assign n2945 = ~n2942 & ~n2943 ;
  assign n2946 = n2944 & n2945 ;
  assign n2947 = \shift[6]  & ~n2946 ;
  assign n2948 = ~n2939 & ~n2947 ;
  assign n2949 = n273 & ~n1727 ;
  assign n2950 = n228 & ~n1751 ;
  assign n2953 = ~n2949 & ~n2950 ;
  assign n2951 = n183 & ~n1707 ;
  assign n2952 = n318 & ~n1743 ;
  assign n2954 = ~n2951 & ~n2952 ;
  assign n2955 = n2953 & n2954 ;
  assign n2956 = ~\shift[6]  & ~n2955 ;
  assign n2957 = n183 & ~n1735 ;
  assign n2958 = n228 & ~n1691 ;
  assign n2961 = ~n2957 & ~n2958 ;
  assign n2959 = n273 & ~n1715 ;
  assign n2960 = n318 & ~n1699 ;
  assign n2962 = ~n2959 & ~n2960 ;
  assign n2963 = n2961 & n2962 ;
  assign n2964 = \shift[6]  & ~n2963 ;
  assign n2965 = ~n2956 & ~n2964 ;
  assign n2966 = n273 & ~n1800 ;
  assign n2967 = n228 & ~n1824 ;
  assign n2970 = ~n2966 & ~n2967 ;
  assign n2968 = n183 & ~n1780 ;
  assign n2969 = n318 & ~n1816 ;
  assign n2971 = ~n2968 & ~n2969 ;
  assign n2972 = n2970 & n2971 ;
  assign n2973 = ~\shift[6]  & ~n2972 ;
  assign n2974 = n183 & ~n1808 ;
  assign n2975 = n228 & ~n1764 ;
  assign n2978 = ~n2974 & ~n2975 ;
  assign n2976 = n273 & ~n1788 ;
  assign n2977 = n318 & ~n1772 ;
  assign n2979 = ~n2976 & ~n2977 ;
  assign n2980 = n2978 & n2979 ;
  assign n2981 = \shift[6]  & ~n2980 ;
  assign n2982 = ~n2973 & ~n2981 ;
  assign n2983 = n273 & ~n1873 ;
  assign n2984 = n183 & ~n1853 ;
  assign n2987 = ~n2983 & ~n2984 ;
  assign n2985 = n318 & ~n1889 ;
  assign n2986 = n228 & ~n1897 ;
  assign n2988 = ~n2985 & ~n2986 ;
  assign n2989 = n2987 & n2988 ;
  assign n2990 = ~\shift[6]  & ~n2989 ;
  assign n2991 = n183 & ~n1881 ;
  assign n2992 = n228 & ~n1837 ;
  assign n2995 = ~n2991 & ~n2992 ;
  assign n2993 = n273 & ~n1861 ;
  assign n2994 = n318 & ~n1845 ;
  assign n2996 = ~n2993 & ~n2994 ;
  assign n2997 = n2995 & n2996 ;
  assign n2998 = \shift[6]  & ~n2997 ;
  assign n2999 = ~n2990 & ~n2998 ;
  assign n3000 = n273 & ~n1946 ;
  assign n3001 = n183 & ~n1926 ;
  assign n3004 = ~n3000 & ~n3001 ;
  assign n3002 = n318 & ~n1962 ;
  assign n3003 = n228 & ~n1970 ;
  assign n3005 = ~n3002 & ~n3003 ;
  assign n3006 = n3004 & n3005 ;
  assign n3007 = ~\shift[6]  & ~n3006 ;
  assign n3008 = n183 & ~n1954 ;
  assign n3009 = n228 & ~n1910 ;
  assign n3012 = ~n3008 & ~n3009 ;
  assign n3010 = n273 & ~n1934 ;
  assign n3011 = n318 & ~n1918 ;
  assign n3013 = ~n3010 & ~n3011 ;
  assign n3014 = n3012 & n3013 ;
  assign n3015 = \shift[6]  & ~n3014 ;
  assign n3016 = ~n3007 & ~n3015 ;
  assign n3017 = n273 & ~n2019 ;
  assign n3018 = n183 & ~n1999 ;
  assign n3021 = ~n3017 & ~n3018 ;
  assign n3019 = n318 & ~n2035 ;
  assign n3020 = n228 & ~n2043 ;
  assign n3022 = ~n3019 & ~n3020 ;
  assign n3023 = n3021 & n3022 ;
  assign n3024 = ~\shift[6]  & ~n3023 ;
  assign n3025 = n183 & ~n2027 ;
  assign n3026 = n228 & ~n1983 ;
  assign n3029 = ~n3025 & ~n3026 ;
  assign n3027 = n273 & ~n2007 ;
  assign n3028 = n318 & ~n1991 ;
  assign n3030 = ~n3027 & ~n3028 ;
  assign n3031 = n3029 & n3030 ;
  assign n3032 = \shift[6]  & ~n3031 ;
  assign n3033 = ~n3024 & ~n3032 ;
  assign n3034 = n273 & ~n2092 ;
  assign n3035 = n183 & ~n2072 ;
  assign n3038 = ~n3034 & ~n3035 ;
  assign n3036 = n318 & ~n2108 ;
  assign n3037 = n228 & ~n2116 ;
  assign n3039 = ~n3036 & ~n3037 ;
  assign n3040 = n3038 & n3039 ;
  assign n3041 = ~\shift[6]  & ~n3040 ;
  assign n3042 = n183 & ~n2100 ;
  assign n3043 = n228 & ~n2056 ;
  assign n3046 = ~n3042 & ~n3043 ;
  assign n3044 = n273 & ~n2080 ;
  assign n3045 = n318 & ~n2064 ;
  assign n3047 = ~n3044 & ~n3045 ;
  assign n3048 = n3046 & n3047 ;
  assign n3049 = \shift[6]  & ~n3048 ;
  assign n3050 = ~n3041 & ~n3049 ;
  assign n3051 = n273 & ~n2165 ;
  assign n3052 = n183 & ~n2145 ;
  assign n3055 = ~n3051 & ~n3052 ;
  assign n3053 = n318 & ~n2181 ;
  assign n3054 = n228 & ~n2189 ;
  assign n3056 = ~n3053 & ~n3054 ;
  assign n3057 = n3055 & n3056 ;
  assign n3058 = ~\shift[6]  & ~n3057 ;
  assign n3059 = n183 & ~n2173 ;
  assign n3060 = n228 & ~n2129 ;
  assign n3063 = ~n3059 & ~n3060 ;
  assign n3061 = n273 & ~n2153 ;
  assign n3062 = n318 & ~n2137 ;
  assign n3064 = ~n3061 & ~n3062 ;
  assign n3065 = n3063 & n3064 ;
  assign n3066 = \shift[6]  & ~n3065 ;
  assign n3067 = ~n3058 & ~n3066 ;
  assign n3068 = n273 & ~n2238 ;
  assign n3069 = n183 & ~n2218 ;
  assign n3072 = ~n3068 & ~n3069 ;
  assign n3070 = n318 & ~n2254 ;
  assign n3071 = n228 & ~n2262 ;
  assign n3073 = ~n3070 & ~n3071 ;
  assign n3074 = n3072 & n3073 ;
  assign n3075 = ~\shift[6]  & ~n3074 ;
  assign n3076 = n183 & ~n2246 ;
  assign n3077 = n228 & ~n2202 ;
  assign n3080 = ~n3076 & ~n3077 ;
  assign n3078 = n273 & ~n2226 ;
  assign n3079 = n318 & ~n2210 ;
  assign n3081 = ~n3078 & ~n3079 ;
  assign n3082 = n3080 & n3081 ;
  assign n3083 = \shift[6]  & ~n3082 ;
  assign n3084 = ~n3075 & ~n3083 ;
  assign n3085 = ~\shift[6]  & ~n504 ;
  assign n3086 = \shift[6]  & ~n322 ;
  assign n3087 = ~n3085 & ~n3086 ;
  assign n3088 = ~\shift[6]  & ~n925 ;
  assign n3089 = \shift[6]  & ~n717 ;
  assign n3090 = ~n3088 & ~n3089 ;
  assign n3091 = ~\shift[6]  & ~n1096 ;
  assign n3092 = \shift[6]  & ~n1010 ;
  assign n3093 = ~n3091 & ~n3092 ;
  assign n3094 = ~\shift[6]  & ~n1390 ;
  assign n3095 = \shift[6]  & ~n1245 ;
  assign n3096 = ~n3094 & ~n3095 ;
  assign n3097 = ~\shift[6]  & ~n1463 ;
  assign n3098 = \shift[6]  & ~n1427 ;
  assign n3099 = ~n3097 & ~n3098 ;
  assign n3100 = ~\shift[6]  & ~n1536 ;
  assign n3101 = \shift[6]  & ~n1500 ;
  assign n3102 = ~n3100 & ~n3101 ;
  assign n3103 = ~\shift[6]  & ~n1609 ;
  assign n3104 = \shift[6]  & ~n1573 ;
  assign n3105 = ~n3103 & ~n3104 ;
  assign n3106 = ~\shift[6]  & ~n1682 ;
  assign n3107 = \shift[6]  & ~n1646 ;
  assign n3108 = ~n3106 & ~n3107 ;
  assign n3109 = ~\shift[6]  & ~n1755 ;
  assign n3110 = \shift[6]  & ~n1719 ;
  assign n3111 = ~n3109 & ~n3110 ;
  assign n3112 = ~\shift[6]  & ~n1828 ;
  assign n3113 = \shift[6]  & ~n1792 ;
  assign n3114 = ~n3112 & ~n3113 ;
  assign n3115 = ~\shift[6]  & ~n1901 ;
  assign n3116 = \shift[6]  & ~n1865 ;
  assign n3117 = ~n3115 & ~n3116 ;
  assign n3118 = ~\shift[6]  & ~n1974 ;
  assign n3119 = \shift[6]  & ~n1938 ;
  assign n3120 = ~n3118 & ~n3119 ;
  assign n3121 = ~\shift[6]  & ~n2047 ;
  assign n3122 = \shift[6]  & ~n2011 ;
  assign n3123 = ~n3121 & ~n3122 ;
  assign n3124 = ~\shift[6]  & ~n2120 ;
  assign n3125 = \shift[6]  & ~n2084 ;
  assign n3126 = ~n3124 & ~n3125 ;
  assign n3127 = ~\shift[6]  & ~n2193 ;
  assign n3128 = \shift[6]  & ~n2157 ;
  assign n3129 = ~n3127 & ~n3128 ;
  assign n3130 = ~\shift[6]  & ~n2266 ;
  assign n3131 = \shift[6]  & ~n2230 ;
  assign n3132 = ~n3130 & ~n3131 ;
  assign n3133 = ~\shift[6]  & ~n2283 ;
  assign n3134 = \shift[6]  & ~n2275 ;
  assign n3135 = ~n3133 & ~n3134 ;
  assign n3136 = ~\shift[6]  & ~n2300 ;
  assign n3137 = \shift[6]  & ~n2292 ;
  assign n3138 = ~n3136 & ~n3137 ;
  assign n3139 = ~\shift[6]  & ~n2317 ;
  assign n3140 = \shift[6]  & ~n2309 ;
  assign n3141 = ~n3139 & ~n3140 ;
  assign n3142 = ~\shift[6]  & ~n2334 ;
  assign n3143 = \shift[6]  & ~n2326 ;
  assign n3144 = ~n3142 & ~n3143 ;
  assign n3145 = ~\shift[6]  & ~n2351 ;
  assign n3146 = \shift[6]  & ~n2343 ;
  assign n3147 = ~n3145 & ~n3146 ;
  assign n3148 = ~\shift[6]  & ~n2368 ;
  assign n3149 = \shift[6]  & ~n2360 ;
  assign n3150 = ~n3148 & ~n3149 ;
  assign n3151 = ~\shift[6]  & ~n2385 ;
  assign n3152 = \shift[6]  & ~n2377 ;
  assign n3153 = ~n3151 & ~n3152 ;
  assign n3154 = ~\shift[6]  & ~n2402 ;
  assign n3155 = \shift[6]  & ~n2394 ;
  assign n3156 = ~n3154 & ~n3155 ;
  assign n3157 = ~\shift[6]  & ~n2419 ;
  assign n3158 = \shift[6]  & ~n2411 ;
  assign n3159 = ~n3157 & ~n3158 ;
  assign n3160 = ~\shift[6]  & ~n2436 ;
  assign n3161 = \shift[6]  & ~n2428 ;
  assign n3162 = ~n3160 & ~n3161 ;
  assign n3163 = ~\shift[6]  & ~n2453 ;
  assign n3164 = \shift[6]  & ~n2445 ;
  assign n3165 = ~n3163 & ~n3164 ;
  assign n3166 = ~\shift[6]  & ~n2470 ;
  assign n3167 = \shift[6]  & ~n2462 ;
  assign n3168 = ~n3166 & ~n3167 ;
  assign n3169 = ~\shift[6]  & ~n2487 ;
  assign n3170 = \shift[6]  & ~n2479 ;
  assign n3171 = ~n3169 & ~n3170 ;
  assign n3172 = ~\shift[6]  & ~n2504 ;
  assign n3173 = \shift[6]  & ~n2496 ;
  assign n3174 = ~n3172 & ~n3173 ;
  assign n3175 = ~\shift[6]  & ~n2521 ;
  assign n3176 = \shift[6]  & ~n2513 ;
  assign n3177 = ~n3175 & ~n3176 ;
  assign n3178 = ~\shift[6]  & ~n2538 ;
  assign n3179 = \shift[6]  & ~n2530 ;
  assign n3180 = ~n3178 & ~n3179 ;
  assign n3181 = ~\shift[6]  & ~n2555 ;
  assign n3182 = \shift[6]  & ~n2547 ;
  assign n3183 = ~n3181 & ~n3182 ;
  assign n3184 = ~\shift[6]  & ~n2572 ;
  assign n3185 = \shift[6]  & ~n2564 ;
  assign n3186 = ~n3184 & ~n3185 ;
  assign n3187 = ~\shift[6]  & ~n2589 ;
  assign n3188 = \shift[6]  & ~n2581 ;
  assign n3189 = ~n3187 & ~n3188 ;
  assign n3190 = ~\shift[6]  & ~n2606 ;
  assign n3191 = \shift[6]  & ~n2598 ;
  assign n3192 = ~n3190 & ~n3191 ;
  assign n3193 = ~\shift[6]  & ~n2623 ;
  assign n3194 = \shift[6]  & ~n2615 ;
  assign n3195 = ~n3193 & ~n3194 ;
  assign n3196 = ~\shift[6]  & ~n2640 ;
  assign n3197 = \shift[6]  & ~n2632 ;
  assign n3198 = ~n3196 & ~n3197 ;
  assign n3199 = ~\shift[6]  & ~n2657 ;
  assign n3200 = \shift[6]  & ~n2649 ;
  assign n3201 = ~n3199 & ~n3200 ;
  assign n3202 = ~\shift[6]  & ~n2674 ;
  assign n3203 = \shift[6]  & ~n2666 ;
  assign n3204 = ~n3202 & ~n3203 ;
  assign n3205 = ~\shift[6]  & ~n2691 ;
  assign n3206 = \shift[6]  & ~n2683 ;
  assign n3207 = ~n3205 & ~n3206 ;
  assign n3208 = ~\shift[6]  & ~n2708 ;
  assign n3209 = \shift[6]  & ~n2700 ;
  assign n3210 = ~n3208 & ~n3209 ;
  assign n3211 = ~\shift[6]  & ~n2725 ;
  assign n3212 = \shift[6]  & ~n2717 ;
  assign n3213 = ~n3211 & ~n3212 ;
  assign n3214 = ~\shift[6]  & ~n2742 ;
  assign n3215 = \shift[6]  & ~n2734 ;
  assign n3216 = ~n3214 & ~n3215 ;
  assign n3217 = ~\shift[6]  & ~n2759 ;
  assign n3218 = \shift[6]  & ~n2751 ;
  assign n3219 = ~n3217 & ~n3218 ;
  assign n3220 = ~\shift[6]  & ~n2776 ;
  assign n3221 = \shift[6]  & ~n2768 ;
  assign n3222 = ~n3220 & ~n3221 ;
  assign n3223 = ~\shift[6]  & ~n2793 ;
  assign n3224 = \shift[6]  & ~n2785 ;
  assign n3225 = ~n3223 & ~n3224 ;
  assign n3226 = ~\shift[6]  & ~n2810 ;
  assign n3227 = \shift[6]  & ~n2802 ;
  assign n3228 = ~n3226 & ~n3227 ;
  assign n3229 = ~\shift[6]  & ~n2827 ;
  assign n3230 = \shift[6]  & ~n2819 ;
  assign n3231 = ~n3229 & ~n3230 ;
  assign n3232 = ~\shift[6]  & ~n2844 ;
  assign n3233 = \shift[6]  & ~n2836 ;
  assign n3234 = ~n3232 & ~n3233 ;
  assign n3235 = ~\shift[6]  & ~n2861 ;
  assign n3236 = \shift[6]  & ~n2853 ;
  assign n3237 = ~n3235 & ~n3236 ;
  assign n3238 = ~\shift[6]  & ~n2878 ;
  assign n3239 = \shift[6]  & ~n2870 ;
  assign n3240 = ~n3238 & ~n3239 ;
  assign n3241 = ~\shift[6]  & ~n2895 ;
  assign n3242 = \shift[6]  & ~n2887 ;
  assign n3243 = ~n3241 & ~n3242 ;
  assign n3244 = ~\shift[6]  & ~n2912 ;
  assign n3245 = \shift[6]  & ~n2904 ;
  assign n3246 = ~n3244 & ~n3245 ;
  assign n3247 = ~\shift[6]  & ~n2929 ;
  assign n3248 = \shift[6]  & ~n2921 ;
  assign n3249 = ~n3247 & ~n3248 ;
  assign n3250 = ~\shift[6]  & ~n2946 ;
  assign n3251 = \shift[6]  & ~n2938 ;
  assign n3252 = ~n3250 & ~n3251 ;
  assign n3253 = ~\shift[6]  & ~n2963 ;
  assign n3254 = \shift[6]  & ~n2955 ;
  assign n3255 = ~n3253 & ~n3254 ;
  assign n3256 = ~\shift[6]  & ~n2980 ;
  assign n3257 = \shift[6]  & ~n2972 ;
  assign n3258 = ~n3256 & ~n3257 ;
  assign n3259 = ~\shift[6]  & ~n2997 ;
  assign n3260 = \shift[6]  & ~n2989 ;
  assign n3261 = ~n3259 & ~n3260 ;
  assign n3262 = ~\shift[6]  & ~n3014 ;
  assign n3263 = \shift[6]  & ~n3006 ;
  assign n3264 = ~n3262 & ~n3263 ;
  assign n3265 = ~\shift[6]  & ~n3031 ;
  assign n3266 = \shift[6]  & ~n3023 ;
  assign n3267 = ~n3265 & ~n3266 ;
  assign n3268 = ~\shift[6]  & ~n3048 ;
  assign n3269 = \shift[6]  & ~n3040 ;
  assign n3270 = ~n3268 & ~n3269 ;
  assign n3271 = ~\shift[6]  & ~n3065 ;
  assign n3272 = \shift[6]  & ~n3057 ;
  assign n3273 = ~n3271 & ~n3272 ;
  assign n3274 = ~\shift[6]  & ~n3082 ;
  assign n3275 = \shift[6]  & ~n3074 ;
  assign n3276 = ~n3274 & ~n3275 ;
  assign \result[0]  = ~n506 ;
  assign \result[1]  = ~n927 ;
  assign \result[2]  = ~n1098 ;
  assign \result[3]  = ~n1392 ;
  assign \result[4]  = ~n1465 ;
  assign \result[5]  = ~n1538 ;
  assign \result[6]  = ~n1611 ;
  assign \result[7]  = ~n1684 ;
  assign \result[8]  = ~n1757 ;
  assign \result[9]  = ~n1830 ;
  assign \result[10]  = ~n1903 ;
  assign \result[11]  = ~n1976 ;
  assign \result[12]  = ~n2049 ;
  assign \result[13]  = ~n2122 ;
  assign \result[14]  = ~n2195 ;
  assign \result[15]  = ~n2268 ;
  assign \result[16]  = ~n2285 ;
  assign \result[17]  = ~n2302 ;
  assign \result[18]  = ~n2319 ;
  assign \result[19]  = ~n2336 ;
  assign \result[20]  = ~n2353 ;
  assign \result[21]  = ~n2370 ;
  assign \result[22]  = ~n2387 ;
  assign \result[23]  = ~n2404 ;
  assign \result[24]  = ~n2421 ;
  assign \result[25]  = ~n2438 ;
  assign \result[26]  = ~n2455 ;
  assign \result[27]  = ~n2472 ;
  assign \result[28]  = ~n2489 ;
  assign \result[29]  = ~n2506 ;
  assign \result[30]  = ~n2523 ;
  assign \result[31]  = ~n2540 ;
  assign \result[32]  = ~n2557 ;
  assign \result[33]  = ~n2574 ;
  assign \result[34]  = ~n2591 ;
  assign \result[35]  = ~n2608 ;
  assign \result[36]  = ~n2625 ;
  assign \result[37]  = ~n2642 ;
  assign \result[38]  = ~n2659 ;
  assign \result[39]  = ~n2676 ;
  assign \result[40]  = ~n2693 ;
  assign \result[41]  = ~n2710 ;
  assign \result[42]  = ~n2727 ;
  assign \result[43]  = ~n2744 ;
  assign \result[44]  = ~n2761 ;
  assign \result[45]  = ~n2778 ;
  assign \result[46]  = ~n2795 ;
  assign \result[47]  = ~n2812 ;
  assign \result[48]  = ~n2829 ;
  assign \result[49]  = ~n2846 ;
  assign \result[50]  = ~n2863 ;
  assign \result[51]  = ~n2880 ;
  assign \result[52]  = ~n2897 ;
  assign \result[53]  = ~n2914 ;
  assign \result[54]  = ~n2931 ;
  assign \result[55]  = ~n2948 ;
  assign \result[56]  = ~n2965 ;
  assign \result[57]  = ~n2982 ;
  assign \result[58]  = ~n2999 ;
  assign \result[59]  = ~n3016 ;
  assign \result[60]  = ~n3033 ;
  assign \result[61]  = ~n3050 ;
  assign \result[62]  = ~n3067 ;
  assign \result[63]  = ~n3084 ;
  assign \result[64]  = ~n3087 ;
  assign \result[65]  = ~n3090 ;
  assign \result[66]  = ~n3093 ;
  assign \result[67]  = ~n3096 ;
  assign \result[68]  = ~n3099 ;
  assign \result[69]  = ~n3102 ;
  assign \result[70]  = ~n3105 ;
  assign \result[71]  = ~n3108 ;
  assign \result[72]  = ~n3111 ;
  assign \result[73]  = ~n3114 ;
  assign \result[74]  = ~n3117 ;
  assign \result[75]  = ~n3120 ;
  assign \result[76]  = ~n3123 ;
  assign \result[77]  = ~n3126 ;
  assign \result[78]  = ~n3129 ;
  assign \result[79]  = ~n3132 ;
  assign \result[80]  = ~n3135 ;
  assign \result[81]  = ~n3138 ;
  assign \result[82]  = ~n3141 ;
  assign \result[83]  = ~n3144 ;
  assign \result[84]  = ~n3147 ;
  assign \result[85]  = ~n3150 ;
  assign \result[86]  = ~n3153 ;
  assign \result[87]  = ~n3156 ;
  assign \result[88]  = ~n3159 ;
  assign \result[89]  = ~n3162 ;
  assign \result[90]  = ~n3165 ;
  assign \result[91]  = ~n3168 ;
  assign \result[92]  = ~n3171 ;
  assign \result[93]  = ~n3174 ;
  assign \result[94]  = ~n3177 ;
  assign \result[95]  = ~n3180 ;
  assign \result[96]  = ~n3183 ;
  assign \result[97]  = ~n3186 ;
  assign \result[98]  = ~n3189 ;
  assign \result[99]  = ~n3192 ;
  assign \result[100]  = ~n3195 ;
  assign \result[101]  = ~n3198 ;
  assign \result[102]  = ~n3201 ;
  assign \result[103]  = ~n3204 ;
  assign \result[104]  = ~n3207 ;
  assign \result[105]  = ~n3210 ;
  assign \result[106]  = ~n3213 ;
  assign \result[107]  = ~n3216 ;
  assign \result[108]  = ~n3219 ;
  assign \result[109]  = ~n3222 ;
  assign \result[110]  = ~n3225 ;
  assign \result[111]  = ~n3228 ;
  assign \result[112]  = ~n3231 ;
  assign \result[113]  = ~n3234 ;
  assign \result[114]  = ~n3237 ;
  assign \result[115]  = ~n3240 ;
  assign \result[116]  = ~n3243 ;
  assign \result[117]  = ~n3246 ;
  assign \result[118]  = ~n3249 ;
  assign \result[119]  = ~n3252 ;
  assign \result[120]  = ~n3255 ;
  assign \result[121]  = ~n3258 ;
  assign \result[122]  = ~n3261 ;
  assign \result[123]  = ~n3264 ;
  assign \result[124]  = ~n3267 ;
  assign \result[125]  = ~n3270 ;
  assign \result[126]  = ~n3273 ;
  assign \result[127]  = ~n3276 ;
endmodule
