module top (\g100_reg/NET0131 , \g1037_reg/NET0131 , \g103_reg/NET0131 , \g1041_reg/NET0131 , \g1045_reg/NET0131 , \g1049_reg/NET0131 , \g104_reg/NET0131 , \g1053_reg/NET0131 , \g1057_reg/NET0131 , \g1061_reg/NET0131 , \g1065_reg/NET0131 , \g1069_reg/NET0131 , \g1073_reg/NET0131 , \g1077_reg/NET0131 , \g1080_pad , \g1087_reg/NET0131 , \g1092_reg/NET0131 , \g1097_reg/NET0131 , \g1098_reg/NET0131 , \g1102_reg/NET0131 , \g1106_reg/NET0131 , \g1110_reg/NET0131 , \g1114_reg/NET0131 , \g1118_reg/NET0131 , \g1122_reg/NET0131 , \g1126_reg/NET0131 , \g1130_reg/NET0131 , \g1134_reg/NET0131 , \g1138_reg/NET0131 , \g1142_reg/NET0131 , \g1148_reg/NET0131 , \g1149_reg/NET0131 , \g1158_reg/NET0131 , \g1166_reg/NET0131 , \g1176_reg/NET0131 , \g1179_reg/NET0131 , \g1189_reg/NET0131 , \g1207_reg/NET0131 , \g1211_reg/NET0131 , \g1214_reg/NET0131 , \g1217_reg/NET0131 , \g1220_reg/NET0131 , \g1223_reg/NET0131 , \g1224_reg/NET0131 , \g1225_reg/NET0131 , \g1226_reg/NET0131 , \g1227_reg/NET0131 , \g1228_reg/NET0131 , \g1229_reg/NET0131 , \g1230_reg/NET0131 , \g1231_reg/NET0131 , \g1247_reg/NET0131 , \g1251_reg/NET0131 , \g1252_reg/NET0131 , \g1253_reg/NET0131 , \g1257_reg/NET0131 , \g1260_reg/NET0131 , \g1263_reg/NET0131 , \g1266_reg/NET0131 , \g1268_reg/NET0131 , \g1269_reg/NET0131 , \g1272_reg/NET0131 , \g1276_reg/NET0131 , \g1280_reg/NET0131 , \g1284_reg/NET0131 , \g1288_reg/NET0131 , \g1292_reg/NET0131 , \g1296_reg/NET0131 , \g1300_reg/NET0131 , \g1304_reg/NET0131 , \g1307_reg/NET0131 , \g1313_reg/NET0131 , \g1317_reg/NET0131 , \g1318_reg/NET0131 , \g1319_reg/NET0131 , \g1320_reg/NET0131 , \g1321_reg/NET0131 , \g1322_reg/NET0131 , \g1323_reg/NET0131 , \g1324_reg/NET0131 , \g1325_reg/NET0131 , \g1326_reg/NET0131 , \g1327_reg/NET0131 , \g1328_reg/NET0131 , \g1329_reg/NET0131 , \g1330_reg/NET0131 , \g1333_reg/NET0131 , \g1336_reg/NET0131 , \g1339_reg/NET0131 , \g1342_reg/NET0131 , \g1345_reg/NET0131 , \g1348_reg/NET0131 , \g1351_reg/NET0131 , \g1354_reg/NET0131 , \g1357_reg/NET0131 , \g1360_reg/NET0131 , \g1363_reg/NET0131 , \g1364_reg/NET0131 , \g1365_reg/NET0131 , \g1366_reg/NET0131 , \g1367_reg/NET0131 , \g1368_reg/NET0131 , \g1369_reg/NET0131 , \g1370_reg/NET0131 , \g1371_reg/NET0131 , \g1372_reg/NET0131 , \g1373_reg/NET0131 , \g1374_reg/NET0131 , \g1375_reg/NET0131 , \g1405_reg/NET0131 , \g1408_reg/NET0131 , \g1412_reg/NET0131 , \g1415_reg/NET0131 , \g1416_reg/NET0131 , \g1421_reg/NET0131 , \g1428_reg/NET0131 , \g1430_reg/NET0131 , \g1432_reg/NET0131 , \g1435_reg/NET0131 , \g1439_reg/NET0131 , \g1444_reg/NET0131 , \g1450_reg/NET0131 , \g1454_reg/NET0131 , \g1462_reg/NET0131 , \g1467_reg/NET0131 , \g1472_reg/NET0131 , \g1481_reg/NET0131 , \g1486_reg/NET0131 , \g1489_reg/NET0131 , \g1494_reg/NET0131 , \g1499_reg/NET0131 , \g1504_reg/NET0131 , \g1509_reg/NET0131 , \g1514_reg/NET0131 , \g1519_reg/NET0131 , \g1944_pad , \g2662_pad , \g2888_pad , \g2_reg/NET0131 , \g4370_pad , \g4371_pad , \g4372_pad , \g4373_pad , \g43_pad , \g652_reg/NET0131 , \g7423_pad , \g7424_pad , \g7425_pad , \g7504_pad , \g7505_pad , \g7507_pad , \g7508_pad , \g785_pad , \g866_reg/NET0131 , \g871_reg/NET0131 , \g889_reg/NET0131 , \g929_reg/NET0131 , \g933_reg/NET0131 , \g936_reg/NET0131 , \g940_reg/NET0131 , \g942_reg/NET0131 , \g943_reg/NET0131 , \g944_reg/NET0131 , \g950_reg/NET0131 , \g951_reg/NET0131 , \g952_reg/NET0131 , \g953_reg/NET0131 , \g954_reg/NET0131 , \g962_pad , \g1006_pad , \g1158_reg/P0001 , \g1252_reg/P0001 , \g1260_reg/P0001 , \g1416_reg/NET0131_syn_2 , \g17/_0_ , \g19189/_0_ , \g19252/_0_ , \g19253/_0_ , \g19273/_3_ , \g19284/_0_ , \g19285/_0_ , \g19295/_3_ , \g19302/_0_ , \g19303/_0_ , \g19304/_0_ , \g19308/_0_ , \g19309/_0_ , \g19310/_0_ , \g19321/_0_ , \g19326/_3_ , \g19331/_0_ , \g19341/_0_ , \g19366/_0_ , \g19372/_3_ , \g19385/_0_ , \g19386/_0_ , \g19387/_0_ , \g19388/_0_ , \g19389/_0_ , \g19390/_0_ , \g19392/_0_ , \g19393/_0_ , \g19394/_0_ , \g19398/_0_ , \g19399/_0_ , \g19400/_0_ , \g19401/_0_ , \g19403/_0_ , \g19405/_0_ , \g19406/_0_ , \g19437/_0_ , \g19438/_0_ , \g19445/_0_ , \g19446/_0_ , \g19450/_3_ , \g19472/_0_ , \g19473/_0_ , \g19474/_0_ , \g19476/_0_ , \g19484/_0_ , \g19485/_0_ , \g19492/_0_ , \g19493/_0_ , \g19499/_0_ , \g19500/_0_ , \g19501/_0_ , \g19502/_0_ , \g19503/_0_ , \g19504/_0_ , \g19507/_3_ , \g19508/_3_ , \g19512/_3_ , \g19513/_3_ , \g19514/_3_ , \g19528/_0_ , \g19529/_0_ , \g19534/_0_ , \g19535/_0_ , \g19536/_0_ , \g19538/_0_ , \g19542/_0_ , \g19560/_0_ , \g19563/_0_ , \g19565/_0_ , \g19567/_0_ , \g19569/_1_ , \g19572/_0_ , \g19574/_3_ , \g19614/_0_ , \g19615/_0_ , \g19620/_0_ , \g19626/_0_ , \g19629/_0_ , \g19631/_0_ , \g19666/_0_ , \g19667/_0_ , \g19669/_0_ , \g19677/_0_ , \g19690/_3_ , \g19721/_0_ , \g19723/_0_ , \g19723/_1_ , \g19725/_2_ , \g19751/_0_ , \g19752/_0_ , \g19753/_0_ , \g19755/_0_ , \g19815/_0_ , \g19821/_0_ , \g19822/_0_ , \g19833/_0_ , \g19877/_0_ , \g19898/_0_ , \g19899/_0_ , \g19900/_0_ , \g19901/_0_ , \g19908/_0_ , \g19927/_0_ , \g19928/_0_ , \g19930/_0_ , \g19931/_0_ , \g19932/_0_ , \g19934/_0_ , \g19992/_0_ , \g19993/_0_ , \g20002/_0_ , \g20008/_0_ , \g20010/_0_ , \g20016/_0_ , \g20110/_0_ , \g20117/_0_ , \g20118/_0_ , \g20131/_0_ , \g20246/_0_ , \g20704/_0_ , \g20722/_0_ , \g20731/_0_ , \g20732/_2_ , \g20870/_0_ , \g20883/_0_ , \g20931/_0_ , \g20951/_0_ , \g20969/_0_ , \g20989/_0_ , \g21/_2_ , \g21070/_0_ , \g21108/_0_ , \g21122/_0_ , \g21152/_0_ , \g21191/_0_ , \g21279/_0_ , \g21316/_0_ , \g21323/_0_ , \g21349/_3_ , \g21352/_3_ , \g21464/_0_ , \g21472/_0_ , \g21484/_0_ , \g21510/_0_ , \g21517/_0_ , \g21608/_0_ , \g21625/_0_ , \g21644/_1_ , \g4655_pad , \g6850_pad , \g6895_pad , \g7048_pad , \g7103_pad , \g7731_pad , \g7732_pad , \g8219_pad , \g8663_pad );
	input \g100_reg/NET0131  ;
	input \g1037_reg/NET0131  ;
	input \g103_reg/NET0131  ;
	input \g1041_reg/NET0131  ;
	input \g1045_reg/NET0131  ;
	input \g1049_reg/NET0131  ;
	input \g104_reg/NET0131  ;
	input \g1053_reg/NET0131  ;
	input \g1057_reg/NET0131  ;
	input \g1061_reg/NET0131  ;
	input \g1065_reg/NET0131  ;
	input \g1069_reg/NET0131  ;
	input \g1073_reg/NET0131  ;
	input \g1077_reg/NET0131  ;
	input \g1080_pad  ;
	input \g1087_reg/NET0131  ;
	input \g1092_reg/NET0131  ;
	input \g1097_reg/NET0131  ;
	input \g1098_reg/NET0131  ;
	input \g1102_reg/NET0131  ;
	input \g1106_reg/NET0131  ;
	input \g1110_reg/NET0131  ;
	input \g1114_reg/NET0131  ;
	input \g1118_reg/NET0131  ;
	input \g1122_reg/NET0131  ;
	input \g1126_reg/NET0131  ;
	input \g1130_reg/NET0131  ;
	input \g1134_reg/NET0131  ;
	input \g1138_reg/NET0131  ;
	input \g1142_reg/NET0131  ;
	input \g1148_reg/NET0131  ;
	input \g1149_reg/NET0131  ;
	input \g1158_reg/NET0131  ;
	input \g1166_reg/NET0131  ;
	input \g1176_reg/NET0131  ;
	input \g1179_reg/NET0131  ;
	input \g1189_reg/NET0131  ;
	input \g1207_reg/NET0131  ;
	input \g1211_reg/NET0131  ;
	input \g1214_reg/NET0131  ;
	input \g1217_reg/NET0131  ;
	input \g1220_reg/NET0131  ;
	input \g1223_reg/NET0131  ;
	input \g1224_reg/NET0131  ;
	input \g1225_reg/NET0131  ;
	input \g1226_reg/NET0131  ;
	input \g1227_reg/NET0131  ;
	input \g1228_reg/NET0131  ;
	input \g1229_reg/NET0131  ;
	input \g1230_reg/NET0131  ;
	input \g1231_reg/NET0131  ;
	input \g1247_reg/NET0131  ;
	input \g1251_reg/NET0131  ;
	input \g1252_reg/NET0131  ;
	input \g1253_reg/NET0131  ;
	input \g1257_reg/NET0131  ;
	input \g1260_reg/NET0131  ;
	input \g1263_reg/NET0131  ;
	input \g1266_reg/NET0131  ;
	input \g1268_reg/NET0131  ;
	input \g1269_reg/NET0131  ;
	input \g1272_reg/NET0131  ;
	input \g1276_reg/NET0131  ;
	input \g1280_reg/NET0131  ;
	input \g1284_reg/NET0131  ;
	input \g1288_reg/NET0131  ;
	input \g1292_reg/NET0131  ;
	input \g1296_reg/NET0131  ;
	input \g1300_reg/NET0131  ;
	input \g1304_reg/NET0131  ;
	input \g1307_reg/NET0131  ;
	input \g1313_reg/NET0131  ;
	input \g1317_reg/NET0131  ;
	input \g1318_reg/NET0131  ;
	input \g1319_reg/NET0131  ;
	input \g1320_reg/NET0131  ;
	input \g1321_reg/NET0131  ;
	input \g1322_reg/NET0131  ;
	input \g1323_reg/NET0131  ;
	input \g1324_reg/NET0131  ;
	input \g1325_reg/NET0131  ;
	input \g1326_reg/NET0131  ;
	input \g1327_reg/NET0131  ;
	input \g1328_reg/NET0131  ;
	input \g1329_reg/NET0131  ;
	input \g1330_reg/NET0131  ;
	input \g1333_reg/NET0131  ;
	input \g1336_reg/NET0131  ;
	input \g1339_reg/NET0131  ;
	input \g1342_reg/NET0131  ;
	input \g1345_reg/NET0131  ;
	input \g1348_reg/NET0131  ;
	input \g1351_reg/NET0131  ;
	input \g1354_reg/NET0131  ;
	input \g1357_reg/NET0131  ;
	input \g1360_reg/NET0131  ;
	input \g1363_reg/NET0131  ;
	input \g1364_reg/NET0131  ;
	input \g1365_reg/NET0131  ;
	input \g1366_reg/NET0131  ;
	input \g1367_reg/NET0131  ;
	input \g1368_reg/NET0131  ;
	input \g1369_reg/NET0131  ;
	input \g1370_reg/NET0131  ;
	input \g1371_reg/NET0131  ;
	input \g1372_reg/NET0131  ;
	input \g1373_reg/NET0131  ;
	input \g1374_reg/NET0131  ;
	input \g1375_reg/NET0131  ;
	input \g1405_reg/NET0131  ;
	input \g1408_reg/NET0131  ;
	input \g1412_reg/NET0131  ;
	input \g1415_reg/NET0131  ;
	input \g1416_reg/NET0131  ;
	input \g1421_reg/NET0131  ;
	input \g1428_reg/NET0131  ;
	input \g1430_reg/NET0131  ;
	input \g1432_reg/NET0131  ;
	input \g1435_reg/NET0131  ;
	input \g1439_reg/NET0131  ;
	input \g1444_reg/NET0131  ;
	input \g1450_reg/NET0131  ;
	input \g1454_reg/NET0131  ;
	input \g1462_reg/NET0131  ;
	input \g1467_reg/NET0131  ;
	input \g1472_reg/NET0131  ;
	input \g1481_reg/NET0131  ;
	input \g1486_reg/NET0131  ;
	input \g1489_reg/NET0131  ;
	input \g1494_reg/NET0131  ;
	input \g1499_reg/NET0131  ;
	input \g1504_reg/NET0131  ;
	input \g1509_reg/NET0131  ;
	input \g1514_reg/NET0131  ;
	input \g1519_reg/NET0131  ;
	input \g1944_pad  ;
	input \g2662_pad  ;
	input \g2888_pad  ;
	input \g2_reg/NET0131  ;
	input \g4370_pad  ;
	input \g4371_pad  ;
	input \g4372_pad  ;
	input \g4373_pad  ;
	input \g43_pad  ;
	input \g652_reg/NET0131  ;
	input \g7423_pad  ;
	input \g7424_pad  ;
	input \g7425_pad  ;
	input \g7504_pad  ;
	input \g7505_pad  ;
	input \g7507_pad  ;
	input \g7508_pad  ;
	input \g785_pad  ;
	input \g866_reg/NET0131  ;
	input \g871_reg/NET0131  ;
	input \g889_reg/NET0131  ;
	input \g929_reg/NET0131  ;
	input \g933_reg/NET0131  ;
	input \g936_reg/NET0131  ;
	input \g940_reg/NET0131  ;
	input \g942_reg/NET0131  ;
	input \g943_reg/NET0131  ;
	input \g944_reg/NET0131  ;
	input \g950_reg/NET0131  ;
	input \g951_reg/NET0131  ;
	input \g952_reg/NET0131  ;
	input \g953_reg/NET0131  ;
	input \g954_reg/NET0131  ;
	input \g962_pad  ;
	output \g1006_pad  ;
	output \g1158_reg/P0001  ;
	output \g1252_reg/P0001  ;
	output \g1260_reg/P0001  ;
	output \g1416_reg/NET0131_syn_2  ;
	output \g17/_0_  ;
	output \g19189/_0_  ;
	output \g19252/_0_  ;
	output \g19253/_0_  ;
	output \g19273/_3_  ;
	output \g19284/_0_  ;
	output \g19285/_0_  ;
	output \g19295/_3_  ;
	output \g19302/_0_  ;
	output \g19303/_0_  ;
	output \g19304/_0_  ;
	output \g19308/_0_  ;
	output \g19309/_0_  ;
	output \g19310/_0_  ;
	output \g19321/_0_  ;
	output \g19326/_3_  ;
	output \g19331/_0_  ;
	output \g19341/_0_  ;
	output \g19366/_0_  ;
	output \g19372/_3_  ;
	output \g19385/_0_  ;
	output \g19386/_0_  ;
	output \g19387/_0_  ;
	output \g19388/_0_  ;
	output \g19389/_0_  ;
	output \g19390/_0_  ;
	output \g19392/_0_  ;
	output \g19393/_0_  ;
	output \g19394/_0_  ;
	output \g19398/_0_  ;
	output \g19399/_0_  ;
	output \g19400/_0_  ;
	output \g19401/_0_  ;
	output \g19403/_0_  ;
	output \g19405/_0_  ;
	output \g19406/_0_  ;
	output \g19437/_0_  ;
	output \g19438/_0_  ;
	output \g19445/_0_  ;
	output \g19446/_0_  ;
	output \g19450/_3_  ;
	output \g19472/_0_  ;
	output \g19473/_0_  ;
	output \g19474/_0_  ;
	output \g19476/_0_  ;
	output \g19484/_0_  ;
	output \g19485/_0_  ;
	output \g19492/_0_  ;
	output \g19493/_0_  ;
	output \g19499/_0_  ;
	output \g19500/_0_  ;
	output \g19501/_0_  ;
	output \g19502/_0_  ;
	output \g19503/_0_  ;
	output \g19504/_0_  ;
	output \g19507/_3_  ;
	output \g19508/_3_  ;
	output \g19512/_3_  ;
	output \g19513/_3_  ;
	output \g19514/_3_  ;
	output \g19528/_0_  ;
	output \g19529/_0_  ;
	output \g19534/_0_  ;
	output \g19535/_0_  ;
	output \g19536/_0_  ;
	output \g19538/_0_  ;
	output \g19542/_0_  ;
	output \g19560/_0_  ;
	output \g19563/_0_  ;
	output \g19565/_0_  ;
	output \g19567/_0_  ;
	output \g19569/_1_  ;
	output \g19572/_0_  ;
	output \g19574/_3_  ;
	output \g19614/_0_  ;
	output \g19615/_0_  ;
	output \g19620/_0_  ;
	output \g19626/_0_  ;
	output \g19629/_0_  ;
	output \g19631/_0_  ;
	output \g19666/_0_  ;
	output \g19667/_0_  ;
	output \g19669/_0_  ;
	output \g19677/_0_  ;
	output \g19690/_3_  ;
	output \g19721/_0_  ;
	output \g19723/_0_  ;
	output \g19723/_1_  ;
	output \g19725/_2_  ;
	output \g19751/_0_  ;
	output \g19752/_0_  ;
	output \g19753/_0_  ;
	output \g19755/_0_  ;
	output \g19815/_0_  ;
	output \g19821/_0_  ;
	output \g19822/_0_  ;
	output \g19833/_0_  ;
	output \g19877/_0_  ;
	output \g19898/_0_  ;
	output \g19899/_0_  ;
	output \g19900/_0_  ;
	output \g19901/_0_  ;
	output \g19908/_0_  ;
	output \g19927/_0_  ;
	output \g19928/_0_  ;
	output \g19930/_0_  ;
	output \g19931/_0_  ;
	output \g19932/_0_  ;
	output \g19934/_0_  ;
	output \g19992/_0_  ;
	output \g19993/_0_  ;
	output \g20002/_0_  ;
	output \g20008/_0_  ;
	output \g20010/_0_  ;
	output \g20016/_0_  ;
	output \g20110/_0_  ;
	output \g20117/_0_  ;
	output \g20118/_0_  ;
	output \g20131/_0_  ;
	output \g20246/_0_  ;
	output \g20704/_0_  ;
	output \g20722/_0_  ;
	output \g20731/_0_  ;
	output \g20732/_2_  ;
	output \g20870/_0_  ;
	output \g20883/_0_  ;
	output \g20931/_0_  ;
	output \g20951/_0_  ;
	output \g20969/_0_  ;
	output \g20989/_0_  ;
	output \g21/_2_  ;
	output \g21070/_0_  ;
	output \g21108/_0_  ;
	output \g21122/_0_  ;
	output \g21152/_0_  ;
	output \g21191/_0_  ;
	output \g21279/_0_  ;
	output \g21316/_0_  ;
	output \g21323/_0_  ;
	output \g21349/_3_  ;
	output \g21352/_3_  ;
	output \g21464/_0_  ;
	output \g21472/_0_  ;
	output \g21484/_0_  ;
	output \g21510/_0_  ;
	output \g21517/_0_  ;
	output \g21608/_0_  ;
	output \g21625/_0_  ;
	output \g21644/_1_  ;
	output \g4655_pad  ;
	output \g6850_pad  ;
	output \g6895_pad  ;
	output \g7048_pad  ;
	output \g7103_pad  ;
	output \g7731_pad  ;
	output \g7732_pad  ;
	output \g8219_pad  ;
	output \g8663_pad  ;
	wire _w792_ ;
	wire _w791_ ;
	wire _w790_ ;
	wire _w789_ ;
	wire _w788_ ;
	wire _w787_ ;
	wire _w786_ ;
	wire _w785_ ;
	wire _w784_ ;
	wire _w783_ ;
	wire _w782_ ;
	wire _w781_ ;
	wire _w780_ ;
	wire _w779_ ;
	wire _w778_ ;
	wire _w777_ ;
	wire _w776_ ;
	wire _w775_ ;
	wire _w774_ ;
	wire _w773_ ;
	wire _w772_ ;
	wire _w771_ ;
	wire _w770_ ;
	wire _w769_ ;
	wire _w768_ ;
	wire _w767_ ;
	wire _w766_ ;
	wire _w765_ ;
	wire _w764_ ;
	wire _w763_ ;
	wire _w762_ ;
	wire _w761_ ;
	wire _w760_ ;
	wire _w759_ ;
	wire _w758_ ;
	wire _w757_ ;
	wire _w756_ ;
	wire _w755_ ;
	wire _w754_ ;
	wire _w753_ ;
	wire _w752_ ;
	wire _w751_ ;
	wire _w750_ ;
	wire _w749_ ;
	wire _w748_ ;
	wire _w747_ ;
	wire _w746_ ;
	wire _w745_ ;
	wire _w744_ ;
	wire _w743_ ;
	wire _w742_ ;
	wire _w741_ ;
	wire _w740_ ;
	wire _w739_ ;
	wire _w738_ ;
	wire _w737_ ;
	wire _w736_ ;
	wire _w735_ ;
	wire _w734_ ;
	wire _w733_ ;
	wire _w732_ ;
	wire _w731_ ;
	wire _w730_ ;
	wire _w729_ ;
	wire _w728_ ;
	wire _w727_ ;
	wire _w726_ ;
	wire _w725_ ;
	wire _w724_ ;
	wire _w723_ ;
	wire _w722_ ;
	wire _w721_ ;
	wire _w720_ ;
	wire _w719_ ;
	wire _w718_ ;
	wire _w717_ ;
	wire _w716_ ;
	wire _w715_ ;
	wire _w714_ ;
	wire _w713_ ;
	wire _w712_ ;
	wire _w711_ ;
	wire _w426_ ;
	wire _w425_ ;
	wire _w424_ ;
	wire _w423_ ;
	wire _w422_ ;
	wire _w421_ ;
	wire _w420_ ;
	wire _w419_ ;
	wire _w418_ ;
	wire _w417_ ;
	wire _w416_ ;
	wire _w415_ ;
	wire _w414_ ;
	wire _w413_ ;
	wire _w412_ ;
	wire _w411_ ;
	wire _w410_ ;
	wire _w409_ ;
	wire _w408_ ;
	wire _w407_ ;
	wire _w406_ ;
	wire _w405_ ;
	wire _w404_ ;
	wire _w403_ ;
	wire _w402_ ;
	wire _w401_ ;
	wire _w400_ ;
	wire _w399_ ;
	wire _w398_ ;
	wire _w397_ ;
	wire _w396_ ;
	wire _w395_ ;
	wire _w394_ ;
	wire _w393_ ;
	wire _w392_ ;
	wire _w391_ ;
	wire _w390_ ;
	wire _w389_ ;
	wire _w388_ ;
	wire _w387_ ;
	wire _w386_ ;
	wire _w385_ ;
	wire _w384_ ;
	wire _w383_ ;
	wire _w382_ ;
	wire _w381_ ;
	wire _w380_ ;
	wire _w379_ ;
	wire _w378_ ;
	wire _w377_ ;
	wire _w376_ ;
	wire _w375_ ;
	wire _w374_ ;
	wire _w373_ ;
	wire _w372_ ;
	wire _w371_ ;
	wire _w370_ ;
	wire _w369_ ;
	wire _w368_ ;
	wire _w367_ ;
	wire _w366_ ;
	wire _w365_ ;
	wire _w364_ ;
	wire _w363_ ;
	wire _w362_ ;
	wire _w361_ ;
	wire _w360_ ;
	wire _w359_ ;
	wire _w358_ ;
	wire _w357_ ;
	wire _w356_ ;
	wire _w355_ ;
	wire _w354_ ;
	wire _w353_ ;
	wire _w352_ ;
	wire _w351_ ;
	wire _w350_ ;
	wire _w349_ ;
	wire _w348_ ;
	wire _w347_ ;
	wire _w346_ ;
	wire _w345_ ;
	wire _w344_ ;
	wire _w343_ ;
	wire _w342_ ;
	wire _w341_ ;
	wire _w340_ ;
	wire _w339_ ;
	wire _w338_ ;
	wire _w337_ ;
	wire _w336_ ;
	wire _w335_ ;
	wire _w334_ ;
	wire _w333_ ;
	wire _w332_ ;
	wire _w331_ ;
	wire _w330_ ;
	wire _w329_ ;
	wire _w328_ ;
	wire _w327_ ;
	wire _w326_ ;
	wire _w325_ ;
	wire _w324_ ;
	wire _w323_ ;
	wire _w322_ ;
	wire _w321_ ;
	wire _w320_ ;
	wire _w319_ ;
	wire _w318_ ;
	wire _w317_ ;
	wire _w316_ ;
	wire _w315_ ;
	wire _w314_ ;
	wire _w313_ ;
	wire _w312_ ;
	wire _w311_ ;
	wire _w310_ ;
	wire _w309_ ;
	wire _w308_ ;
	wire _w307_ ;
	wire _w306_ ;
	wire _w305_ ;
	wire _w304_ ;
	wire _w303_ ;
	wire _w302_ ;
	wire _w301_ ;
	wire _w300_ ;
	wire _w299_ ;
	wire _w298_ ;
	wire _w297_ ;
	wire _w228_ ;
	wire _w227_ ;
	wire _w226_ ;
	wire _w225_ ;
	wire _w224_ ;
	wire _w223_ ;
	wire _w222_ ;
	wire _w221_ ;
	wire _w220_ ;
	wire _w219_ ;
	wire _w218_ ;
	wire _w217_ ;
	wire _w216_ ;
	wire _w215_ ;
	wire _w214_ ;
	wire _w213_ ;
	wire _w212_ ;
	wire _w211_ ;
	wire _w210_ ;
	wire _w209_ ;
	wire _w208_ ;
	wire _w207_ ;
	wire _w206_ ;
	wire _w205_ ;
	wire _w204_ ;
	wire _w203_ ;
	wire _w202_ ;
	wire _w201_ ;
	wire _w200_ ;
	wire _w199_ ;
	wire _w182_ ;
	wire _w181_ ;
	wire _w180_ ;
	wire _w179_ ;
	wire _w178_ ;
	wire _w177_ ;
	wire _w176_ ;
	wire _w175_ ;
	wire _w174_ ;
	wire _w173_ ;
	wire _w172_ ;
	wire _w171_ ;
	wire _w170_ ;
	wire _w183_ ;
	wire _w184_ ;
	wire _w185_ ;
	wire _w186_ ;
	wire _w187_ ;
	wire _w188_ ;
	wire _w189_ ;
	wire _w190_ ;
	wire _w191_ ;
	wire _w192_ ;
	wire _w193_ ;
	wire _w194_ ;
	wire _w195_ ;
	wire _w196_ ;
	wire _w197_ ;
	wire _w198_ ;
	wire _w229_ ;
	wire _w230_ ;
	wire _w231_ ;
	wire _w232_ ;
	wire _w233_ ;
	wire _w234_ ;
	wire _w235_ ;
	wire _w236_ ;
	wire _w237_ ;
	wire _w238_ ;
	wire _w239_ ;
	wire _w240_ ;
	wire _w241_ ;
	wire _w242_ ;
	wire _w243_ ;
	wire _w244_ ;
	wire _w245_ ;
	wire _w246_ ;
	wire _w247_ ;
	wire _w248_ ;
	wire _w249_ ;
	wire _w250_ ;
	wire _w251_ ;
	wire _w252_ ;
	wire _w253_ ;
	wire _w254_ ;
	wire _w255_ ;
	wire _w256_ ;
	wire _w257_ ;
	wire _w258_ ;
	wire _w259_ ;
	wire _w260_ ;
	wire _w261_ ;
	wire _w262_ ;
	wire _w263_ ;
	wire _w264_ ;
	wire _w265_ ;
	wire _w266_ ;
	wire _w267_ ;
	wire _w268_ ;
	wire _w269_ ;
	wire _w270_ ;
	wire _w271_ ;
	wire _w272_ ;
	wire _w273_ ;
	wire _w274_ ;
	wire _w275_ ;
	wire _w276_ ;
	wire _w277_ ;
	wire _w278_ ;
	wire _w279_ ;
	wire _w280_ ;
	wire _w281_ ;
	wire _w282_ ;
	wire _w283_ ;
	wire _w284_ ;
	wire _w285_ ;
	wire _w286_ ;
	wire _w287_ ;
	wire _w288_ ;
	wire _w289_ ;
	wire _w290_ ;
	wire _w291_ ;
	wire _w292_ ;
	wire _w293_ ;
	wire _w294_ ;
	wire _w295_ ;
	wire _w296_ ;
	wire _w427_ ;
	wire _w428_ ;
	wire _w429_ ;
	wire _w430_ ;
	wire _w431_ ;
	wire _w432_ ;
	wire _w433_ ;
	wire _w434_ ;
	wire _w435_ ;
	wire _w436_ ;
	wire _w437_ ;
	wire _w438_ ;
	wire _w439_ ;
	wire _w440_ ;
	wire _w441_ ;
	wire _w442_ ;
	wire _w443_ ;
	wire _w444_ ;
	wire _w445_ ;
	wire _w446_ ;
	wire _w447_ ;
	wire _w448_ ;
	wire _w449_ ;
	wire _w450_ ;
	wire _w451_ ;
	wire _w452_ ;
	wire _w453_ ;
	wire _w454_ ;
	wire _w455_ ;
	wire _w456_ ;
	wire _w457_ ;
	wire _w458_ ;
	wire _w459_ ;
	wire _w460_ ;
	wire _w461_ ;
	wire _w462_ ;
	wire _w463_ ;
	wire _w464_ ;
	wire _w465_ ;
	wire _w466_ ;
	wire _w467_ ;
	wire _w468_ ;
	wire _w469_ ;
	wire _w470_ ;
	wire _w471_ ;
	wire _w472_ ;
	wire _w473_ ;
	wire _w474_ ;
	wire _w475_ ;
	wire _w476_ ;
	wire _w477_ ;
	wire _w478_ ;
	wire _w479_ ;
	wire _w480_ ;
	wire _w481_ ;
	wire _w482_ ;
	wire _w483_ ;
	wire _w484_ ;
	wire _w485_ ;
	wire _w486_ ;
	wire _w487_ ;
	wire _w488_ ;
	wire _w489_ ;
	wire _w490_ ;
	wire _w491_ ;
	wire _w492_ ;
	wire _w493_ ;
	wire _w494_ ;
	wire _w495_ ;
	wire _w496_ ;
	wire _w497_ ;
	wire _w498_ ;
	wire _w499_ ;
	wire _w500_ ;
	wire _w501_ ;
	wire _w502_ ;
	wire _w503_ ;
	wire _w504_ ;
	wire _w505_ ;
	wire _w506_ ;
	wire _w507_ ;
	wire _w508_ ;
	wire _w509_ ;
	wire _w510_ ;
	wire _w511_ ;
	wire _w512_ ;
	wire _w513_ ;
	wire _w514_ ;
	wire _w515_ ;
	wire _w516_ ;
	wire _w517_ ;
	wire _w518_ ;
	wire _w519_ ;
	wire _w520_ ;
	wire _w521_ ;
	wire _w522_ ;
	wire _w523_ ;
	wire _w524_ ;
	wire _w525_ ;
	wire _w526_ ;
	wire _w527_ ;
	wire _w528_ ;
	wire _w529_ ;
	wire _w530_ ;
	wire _w531_ ;
	wire _w532_ ;
	wire _w533_ ;
	wire _w534_ ;
	wire _w535_ ;
	wire _w536_ ;
	wire _w537_ ;
	wire _w538_ ;
	wire _w539_ ;
	wire _w540_ ;
	wire _w541_ ;
	wire _w542_ ;
	wire _w543_ ;
	wire _w544_ ;
	wire _w545_ ;
	wire _w546_ ;
	wire _w547_ ;
	wire _w548_ ;
	wire _w549_ ;
	wire _w550_ ;
	wire _w551_ ;
	wire _w552_ ;
	wire _w553_ ;
	wire _w554_ ;
	wire _w555_ ;
	wire _w556_ ;
	wire _w557_ ;
	wire _w558_ ;
	wire _w559_ ;
	wire _w560_ ;
	wire _w561_ ;
	wire _w562_ ;
	wire _w563_ ;
	wire _w564_ ;
	wire _w565_ ;
	wire _w566_ ;
	wire _w567_ ;
	wire _w568_ ;
	wire _w569_ ;
	wire _w570_ ;
	wire _w571_ ;
	wire _w572_ ;
	wire _w573_ ;
	wire _w574_ ;
	wire _w575_ ;
	wire _w576_ ;
	wire _w577_ ;
	wire _w578_ ;
	wire _w579_ ;
	wire _w580_ ;
	wire _w581_ ;
	wire _w582_ ;
	wire _w583_ ;
	wire _w584_ ;
	wire _w585_ ;
	wire _w586_ ;
	wire _w587_ ;
	wire _w588_ ;
	wire _w589_ ;
	wire _w590_ ;
	wire _w591_ ;
	wire _w592_ ;
	wire _w593_ ;
	wire _w594_ ;
	wire _w595_ ;
	wire _w596_ ;
	wire _w597_ ;
	wire _w598_ ;
	wire _w599_ ;
	wire _w600_ ;
	wire _w601_ ;
	wire _w602_ ;
	wire _w603_ ;
	wire _w604_ ;
	wire _w605_ ;
	wire _w606_ ;
	wire _w607_ ;
	wire _w608_ ;
	wire _w609_ ;
	wire _w610_ ;
	wire _w611_ ;
	wire _w612_ ;
	wire _w613_ ;
	wire _w614_ ;
	wire _w615_ ;
	wire _w616_ ;
	wire _w617_ ;
	wire _w618_ ;
	wire _w619_ ;
	wire _w620_ ;
	wire _w621_ ;
	wire _w622_ ;
	wire _w623_ ;
	wire _w624_ ;
	wire _w625_ ;
	wire _w626_ ;
	wire _w627_ ;
	wire _w628_ ;
	wire _w629_ ;
	wire _w630_ ;
	wire _w631_ ;
	wire _w632_ ;
	wire _w633_ ;
	wire _w634_ ;
	wire _w635_ ;
	wire _w636_ ;
	wire _w637_ ;
	wire _w638_ ;
	wire _w639_ ;
	wire _w640_ ;
	wire _w641_ ;
	wire _w642_ ;
	wire _w643_ ;
	wire _w644_ ;
	wire _w645_ ;
	wire _w646_ ;
	wire _w647_ ;
	wire _w648_ ;
	wire _w649_ ;
	wire _w650_ ;
	wire _w651_ ;
	wire _w652_ ;
	wire _w653_ ;
	wire _w654_ ;
	wire _w655_ ;
	wire _w656_ ;
	wire _w657_ ;
	wire _w658_ ;
	wire _w659_ ;
	wire _w660_ ;
	wire _w661_ ;
	wire _w662_ ;
	wire _w663_ ;
	wire _w664_ ;
	wire _w665_ ;
	wire _w666_ ;
	wire _w667_ ;
	wire _w668_ ;
	wire _w669_ ;
	wire _w670_ ;
	wire _w671_ ;
	wire _w672_ ;
	wire _w673_ ;
	wire _w674_ ;
	wire _w675_ ;
	wire _w676_ ;
	wire _w677_ ;
	wire _w678_ ;
	wire _w679_ ;
	wire _w680_ ;
	wire _w681_ ;
	wire _w682_ ;
	wire _w683_ ;
	wire _w684_ ;
	wire _w685_ ;
	wire _w686_ ;
	wire _w687_ ;
	wire _w688_ ;
	wire _w689_ ;
	wire _w690_ ;
	wire _w691_ ;
	wire _w692_ ;
	wire _w693_ ;
	wire _w694_ ;
	wire _w695_ ;
	wire _w696_ ;
	wire _w697_ ;
	wire _w698_ ;
	wire _w699_ ;
	wire _w700_ ;
	wire _w701_ ;
	wire _w702_ ;
	wire _w703_ ;
	wire _w704_ ;
	wire _w705_ ;
	wire _w706_ ;
	wire _w707_ ;
	wire _w708_ ;
	wire _w709_ ;
	wire _w710_ ;
	LUT2 #(
		.INIT('h8)
	) name0 (
		\g1330_reg/NET0131 ,
		\g1333_reg/NET0131 ,
		_w170_
	);
	LUT2 #(
		.INIT('h8)
	) name1 (
		\g1336_reg/NET0131 ,
		_w170_,
		_w171_
	);
	LUT2 #(
		.INIT('h8)
	) name2 (
		\g1339_reg/NET0131 ,
		_w171_,
		_w172_
	);
	LUT2 #(
		.INIT('h8)
	) name3 (
		\g1342_reg/NET0131 ,
		_w172_,
		_w173_
	);
	LUT2 #(
		.INIT('h8)
	) name4 (
		\g1345_reg/NET0131 ,
		_w173_,
		_w174_
	);
	LUT2 #(
		.INIT('h1)
	) name5 (
		\g1348_reg/NET0131 ,
		_w174_,
		_w175_
	);
	LUT2 #(
		.INIT('h8)
	) name6 (
		\g1348_reg/NET0131 ,
		_w174_,
		_w176_
	);
	LUT2 #(
		.INIT('h2)
	) name7 (
		\g1247_reg/NET0131 ,
		_w175_,
		_w177_
	);
	LUT2 #(
		.INIT('h4)
	) name8 (
		_w176_,
		_w177_,
		_w178_
	);
	LUT2 #(
		.INIT('h2)
	) name9 (
		\g1073_reg/NET0131 ,
		\g1158_reg/NET0131 ,
		_w179_
	);
	LUT2 #(
		.INIT('h4)
	) name10 (
		\g1073_reg/NET0131 ,
		\g1158_reg/NET0131 ,
		_w180_
	);
	LUT2 #(
		.INIT('h4)
	) name11 (
		\g1251_reg/NET0131 ,
		_w180_,
		_w181_
	);
	LUT2 #(
		.INIT('h8)
	) name12 (
		\g1092_reg/NET0131 ,
		\g1130_reg/NET0131 ,
		_w182_
	);
	LUT2 #(
		.INIT('h8)
	) name13 (
		\g1134_reg/NET0131 ,
		_w182_,
		_w183_
	);
	LUT2 #(
		.INIT('h8)
	) name14 (
		\g1138_reg/NET0131 ,
		_w183_,
		_w184_
	);
	LUT2 #(
		.INIT('h8)
	) name15 (
		\g1149_reg/NET0131 ,
		_w184_,
		_w185_
	);
	LUT2 #(
		.INIT('h8)
	) name16 (
		\g1037_reg/NET0131 ,
		\g1041_reg/NET0131 ,
		_w186_
	);
	LUT2 #(
		.INIT('h8)
	) name17 (
		\g1045_reg/NET0131 ,
		_w186_,
		_w187_
	);
	LUT2 #(
		.INIT('h8)
	) name18 (
		_w185_,
		_w187_,
		_w188_
	);
	LUT2 #(
		.INIT('h8)
	) name19 (
		\g1049_reg/NET0131 ,
		\g1053_reg/NET0131 ,
		_w189_
	);
	LUT2 #(
		.INIT('h8)
	) name20 (
		\g1057_reg/NET0131 ,
		\g1061_reg/NET0131 ,
		_w190_
	);
	LUT2 #(
		.INIT('h8)
	) name21 (
		_w189_,
		_w190_,
		_w191_
	);
	LUT2 #(
		.INIT('h8)
	) name22 (
		_w188_,
		_w191_,
		_w192_
	);
	LUT2 #(
		.INIT('h8)
	) name23 (
		\g1065_reg/NET0131 ,
		_w192_,
		_w193_
	);
	LUT2 #(
		.INIT('h8)
	) name24 (
		_w181_,
		_w193_,
		_w194_
	);
	LUT2 #(
		.INIT('h8)
	) name25 (
		\g1069_reg/NET0131 ,
		_w194_,
		_w195_
	);
	LUT2 #(
		.INIT('h1)
	) name26 (
		_w179_,
		_w195_,
		_w196_
	);
	LUT2 #(
		.INIT('h2)
	) name27 (
		\g936_reg/NET0131 ,
		\g940_reg/NET0131 ,
		_w197_
	);
	LUT2 #(
		.INIT('h4)
	) name28 (
		\g936_reg/NET0131 ,
		\g940_reg/NET0131 ,
		_w198_
	);
	LUT2 #(
		.INIT('h4)
	) name29 (
		\g943_reg/NET0131 ,
		_w198_,
		_w199_
	);
	LUT2 #(
		.INIT('h1)
	) name30 (
		_w197_,
		_w199_,
		_w200_
	);
	LUT2 #(
		.INIT('h2)
	) name31 (
		\g1158_reg/NET0131 ,
		\g1251_reg/NET0131 ,
		_w201_
	);
	LUT2 #(
		.INIT('h8)
	) name32 (
		\g1073_reg/NET0131 ,
		\g1158_reg/NET0131 ,
		_w202_
	);
	LUT2 #(
		.INIT('h1)
	) name33 (
		_w201_,
		_w202_,
		_w203_
	);
	LUT2 #(
		.INIT('h8)
	) name34 (
		\g1049_reg/NET0131 ,
		_w203_,
		_w204_
	);
	LUT2 #(
		.INIT('h1)
	) name35 (
		\g1049_reg/NET0131 ,
		_w188_,
		_w205_
	);
	LUT2 #(
		.INIT('h8)
	) name36 (
		\g1049_reg/NET0131 ,
		_w188_,
		_w206_
	);
	LUT2 #(
		.INIT('h2)
	) name37 (
		_w181_,
		_w205_,
		_w207_
	);
	LUT2 #(
		.INIT('h4)
	) name38 (
		_w206_,
		_w207_,
		_w208_
	);
	LUT2 #(
		.INIT('h1)
	) name39 (
		_w204_,
		_w208_,
		_w209_
	);
	LUT2 #(
		.INIT('h2)
	) name40 (
		\g954_reg/NET0131 ,
		_w197_,
		_w210_
	);
	LUT2 #(
		.INIT('h8)
	) name41 (
		\g2_reg/NET0131 ,
		_w197_,
		_w211_
	);
	LUT2 #(
		.INIT('h1)
	) name42 (
		_w210_,
		_w211_,
		_w212_
	);
	LUT2 #(
		.INIT('h4)
	) name43 (
		\g1251_reg/NET0131 ,
		\g1481_reg/NET0131 ,
		_w213_
	);
	LUT2 #(
		.INIT('h8)
	) name44 (
		\g1489_reg/NET0131 ,
		\g1494_reg/NET0131 ,
		_w214_
	);
	LUT2 #(
		.INIT('h8)
	) name45 (
		_w213_,
		_w214_,
		_w215_
	);
	LUT2 #(
		.INIT('h8)
	) name46 (
		\g1514_reg/NET0131 ,
		\g1519_reg/NET0131 ,
		_w216_
	);
	LUT2 #(
		.INIT('h8)
	) name47 (
		\g1462_reg/NET0131 ,
		\g1467_reg/NET0131 ,
		_w217_
	);
	LUT2 #(
		.INIT('h8)
	) name48 (
		\g1472_reg/NET0131 ,
		\g1499_reg/NET0131 ,
		_w218_
	);
	LUT2 #(
		.INIT('h8)
	) name49 (
		_w217_,
		_w218_,
		_w219_
	);
	LUT2 #(
		.INIT('h8)
	) name50 (
		_w216_,
		_w219_,
		_w220_
	);
	LUT2 #(
		.INIT('h8)
	) name51 (
		_w215_,
		_w220_,
		_w221_
	);
	LUT2 #(
		.INIT('h8)
	) name52 (
		\g1499_reg/NET0131 ,
		\g1504_reg/NET0131 ,
		_w222_
	);
	LUT2 #(
		.INIT('h8)
	) name53 (
		_w215_,
		_w222_,
		_w223_
	);
	LUT2 #(
		.INIT('h8)
	) name54 (
		\g1509_reg/NET0131 ,
		_w223_,
		_w224_
	);
	LUT2 #(
		.INIT('h8)
	) name55 (
		\g1514_reg/NET0131 ,
		_w224_,
		_w225_
	);
	LUT2 #(
		.INIT('h1)
	) name56 (
		\g1514_reg/NET0131 ,
		_w224_,
		_w226_
	);
	LUT2 #(
		.INIT('h1)
	) name57 (
		_w221_,
		_w225_,
		_w227_
	);
	LUT2 #(
		.INIT('h4)
	) name58 (
		_w226_,
		_w227_,
		_w228_
	);
	LUT2 #(
		.INIT('h8)
	) name59 (
		\g1087_reg/NET0131 ,
		\g1098_reg/NET0131 ,
		_w229_
	);
	LUT2 #(
		.INIT('h8)
	) name60 (
		\g1102_reg/NET0131 ,
		_w229_,
		_w230_
	);
	LUT2 #(
		.INIT('h8)
	) name61 (
		\g1106_reg/NET0131 ,
		_w230_,
		_w231_
	);
	LUT2 #(
		.INIT('h8)
	) name62 (
		\g1148_reg/NET0131 ,
		_w231_,
		_w232_
	);
	LUT2 #(
		.INIT('h8)
	) name63 (
		\g1110_reg/NET0131 ,
		_w232_,
		_w233_
	);
	LUT2 #(
		.INIT('h8)
	) name64 (
		\g1114_reg/NET0131 ,
		_w233_,
		_w234_
	);
	LUT2 #(
		.INIT('h1)
	) name65 (
		\g1118_reg/NET0131 ,
		_w234_,
		_w235_
	);
	LUT2 #(
		.INIT('h8)
	) name66 (
		\g1118_reg/NET0131 ,
		_w234_,
		_w236_
	);
	LUT2 #(
		.INIT('h1)
	) name67 (
		_w235_,
		_w236_,
		_w237_
	);
	LUT2 #(
		.INIT('h1)
	) name68 (
		\g1097_reg/NET0131 ,
		_w237_,
		_w238_
	);
	LUT2 #(
		.INIT('h2)
	) name69 (
		\g953_reg/NET0131 ,
		_w197_,
		_w239_
	);
	LUT2 #(
		.INIT('h1)
	) name70 (
		_w211_,
		_w239_,
		_w240_
	);
	LUT2 #(
		.INIT('h8)
	) name71 (
		\g1148_reg/NET0131 ,
		_w230_,
		_w241_
	);
	LUT2 #(
		.INIT('h1)
	) name72 (
		\g1106_reg/NET0131 ,
		_w241_,
		_w242_
	);
	LUT2 #(
		.INIT('h1)
	) name73 (
		_w232_,
		_w242_,
		_w243_
	);
	LUT2 #(
		.INIT('h1)
	) name74 (
		\g1097_reg/NET0131 ,
		_w243_,
		_w244_
	);
	LUT2 #(
		.INIT('h1)
	) name75 (
		\g1110_reg/NET0131 ,
		_w232_,
		_w245_
	);
	LUT2 #(
		.INIT('h1)
	) name76 (
		_w233_,
		_w245_,
		_w246_
	);
	LUT2 #(
		.INIT('h1)
	) name77 (
		\g1097_reg/NET0131 ,
		_w246_,
		_w247_
	);
	LUT2 #(
		.INIT('h1)
	) name78 (
		\g1114_reg/NET0131 ,
		_w233_,
		_w248_
	);
	LUT2 #(
		.INIT('h1)
	) name79 (
		_w234_,
		_w248_,
		_w249_
	);
	LUT2 #(
		.INIT('h1)
	) name80 (
		\g1097_reg/NET0131 ,
		_w249_,
		_w250_
	);
	LUT2 #(
		.INIT('h1)
	) name81 (
		\g1509_reg/NET0131 ,
		_w223_,
		_w251_
	);
	LUT2 #(
		.INIT('h1)
	) name82 (
		_w221_,
		_w224_,
		_w252_
	);
	LUT2 #(
		.INIT('h4)
	) name83 (
		_w251_,
		_w252_,
		_w253_
	);
	LUT2 #(
		.INIT('h1)
	) name84 (
		\g1097_reg/NET0131 ,
		\g1148_reg/NET0131 ,
		_w254_
	);
	LUT2 #(
		.INIT('h8)
	) name85 (
		\g1098_reg/NET0131 ,
		_w254_,
		_w255_
	);
	LUT2 #(
		.INIT('h4)
	) name86 (
		\g1097_reg/NET0131 ,
		\g1148_reg/NET0131 ,
		_w256_
	);
	LUT2 #(
		.INIT('h1)
	) name87 (
		\g1087_reg/NET0131 ,
		\g1098_reg/NET0131 ,
		_w257_
	);
	LUT2 #(
		.INIT('h4)
	) name88 (
		_w229_,
		_w256_,
		_w258_
	);
	LUT2 #(
		.INIT('h4)
	) name89 (
		_w257_,
		_w258_,
		_w259_
	);
	LUT2 #(
		.INIT('h1)
	) name90 (
		_w255_,
		_w259_,
		_w260_
	);
	LUT2 #(
		.INIT('h8)
	) name91 (
		\g1102_reg/NET0131 ,
		_w254_,
		_w261_
	);
	LUT2 #(
		.INIT('h1)
	) name92 (
		\g1102_reg/NET0131 ,
		_w229_,
		_w262_
	);
	LUT2 #(
		.INIT('h4)
	) name93 (
		_w230_,
		_w256_,
		_w263_
	);
	LUT2 #(
		.INIT('h4)
	) name94 (
		_w262_,
		_w263_,
		_w264_
	);
	LUT2 #(
		.INIT('h1)
	) name95 (
		_w261_,
		_w264_,
		_w265_
	);
	LUT2 #(
		.INIT('h8)
	) name96 (
		\g1037_reg/NET0131 ,
		_w203_,
		_w266_
	);
	LUT2 #(
		.INIT('h1)
	) name97 (
		\g1037_reg/NET0131 ,
		_w185_,
		_w267_
	);
	LUT2 #(
		.INIT('h8)
	) name98 (
		\g1037_reg/NET0131 ,
		_w185_,
		_w268_
	);
	LUT2 #(
		.INIT('h2)
	) name99 (
		_w181_,
		_w267_,
		_w269_
	);
	LUT2 #(
		.INIT('h4)
	) name100 (
		_w268_,
		_w269_,
		_w270_
	);
	LUT2 #(
		.INIT('h1)
	) name101 (
		_w266_,
		_w270_,
		_w271_
	);
	LUT2 #(
		.INIT('h2)
	) name102 (
		\g952_reg/NET0131 ,
		_w197_,
		_w272_
	);
	LUT2 #(
		.INIT('h1)
	) name103 (
		_w211_,
		_w272_,
		_w273_
	);
	LUT2 #(
		.INIT('h2)
	) name104 (
		\g1087_reg/NET0131 ,
		\g1148_reg/NET0131 ,
		_w274_
	);
	LUT2 #(
		.INIT('h4)
	) name105 (
		\g1087_reg/NET0131 ,
		\g1148_reg/NET0131 ,
		_w275_
	);
	LUT2 #(
		.INIT('h1)
	) name106 (
		_w274_,
		_w275_,
		_w276_
	);
	LUT2 #(
		.INIT('h1)
	) name107 (
		\g1097_reg/NET0131 ,
		_w276_,
		_w277_
	);
	LUT2 #(
		.INIT('h8)
	) name108 (
		\g1499_reg/NET0131 ,
		_w215_,
		_w278_
	);
	LUT2 #(
		.INIT('h1)
	) name109 (
		\g1504_reg/NET0131 ,
		_w278_,
		_w279_
	);
	LUT2 #(
		.INIT('h1)
	) name110 (
		_w221_,
		_w223_,
		_w280_
	);
	LUT2 #(
		.INIT('h4)
	) name111 (
		_w279_,
		_w280_,
		_w281_
	);
	LUT2 #(
		.INIT('h8)
	) name112 (
		\g1149_reg/NET0131 ,
		_w203_,
		_w282_
	);
	LUT2 #(
		.INIT('h1)
	) name113 (
		\g1149_reg/NET0131 ,
		_w184_,
		_w283_
	);
	LUT2 #(
		.INIT('h2)
	) name114 (
		_w181_,
		_w185_,
		_w284_
	);
	LUT2 #(
		.INIT('h4)
	) name115 (
		_w283_,
		_w284_,
		_w285_
	);
	LUT2 #(
		.INIT('h1)
	) name116 (
		_w282_,
		_w285_,
		_w286_
	);
	LUT2 #(
		.INIT('h2)
	) name117 (
		\g951_reg/NET0131 ,
		_w197_,
		_w287_
	);
	LUT2 #(
		.INIT('h1)
	) name118 (
		_w211_,
		_w287_,
		_w288_
	);
	LUT2 #(
		.INIT('h4)
	) name119 (
		\g1092_reg/NET0131 ,
		_w201_,
		_w289_
	);
	LUT2 #(
		.INIT('h2)
	) name120 (
		\g1092_reg/NET0131 ,
		_w201_,
		_w290_
	);
	LUT2 #(
		.INIT('h1)
	) name121 (
		_w289_,
		_w290_,
		_w291_
	);
	LUT2 #(
		.INIT('h1)
	) name122 (
		_w202_,
		_w291_,
		_w292_
	);
	LUT2 #(
		.INIT('h8)
	) name123 (
		\g100_reg/NET0131 ,
		\g1329_reg/NET0131 ,
		_w293_
	);
	LUT2 #(
		.INIT('h8)
	) name124 (
		\g1313_reg/NET0131 ,
		\g1317_reg/NET0131 ,
		_w294_
	);
	LUT2 #(
		.INIT('h1)
	) name125 (
		\g1318_reg/NET0131 ,
		_w294_,
		_w295_
	);
	LUT2 #(
		.INIT('h8)
	) name126 (
		\g1318_reg/NET0131 ,
		_w294_,
		_w296_
	);
	LUT2 #(
		.INIT('h1)
	) name127 (
		\g1329_reg/NET0131 ,
		_w295_,
		_w297_
	);
	LUT2 #(
		.INIT('h4)
	) name128 (
		_w296_,
		_w297_,
		_w298_
	);
	LUT2 #(
		.INIT('h1)
	) name129 (
		_w293_,
		_w298_,
		_w299_
	);
	LUT2 #(
		.INIT('h2)
	) name130 (
		\g1251_reg/NET0131 ,
		\g1481_reg/NET0131 ,
		_w300_
	);
	LUT2 #(
		.INIT('h1)
	) name131 (
		_w213_,
		_w300_,
		_w301_
	);
	LUT2 #(
		.INIT('h8)
	) name132 (
		\g1489_reg/NET0131 ,
		_w213_,
		_w302_
	);
	LUT2 #(
		.INIT('h1)
	) name133 (
		\g1489_reg/NET0131 ,
		_w213_,
		_w303_
	);
	LUT2 #(
		.INIT('h1)
	) name134 (
		_w302_,
		_w303_,
		_w304_
	);
	LUT2 #(
		.INIT('h8)
	) name135 (
		\g103_reg/NET0131 ,
		\g1329_reg/NET0131 ,
		_w305_
	);
	LUT2 #(
		.INIT('h8)
	) name136 (
		\g1318_reg/NET0131 ,
		\g1319_reg/NET0131 ,
		_w306_
	);
	LUT2 #(
		.INIT('h8)
	) name137 (
		_w294_,
		_w306_,
		_w307_
	);
	LUT2 #(
		.INIT('h8)
	) name138 (
		\g1320_reg/NET0131 ,
		\g1321_reg/NET0131 ,
		_w308_
	);
	LUT2 #(
		.INIT('h8)
	) name139 (
		\g1322_reg/NET0131 ,
		_w308_,
		_w309_
	);
	LUT2 #(
		.INIT('h8)
	) name140 (
		_w307_,
		_w309_,
		_w310_
	);
	LUT2 #(
		.INIT('h8)
	) name141 (
		\g1323_reg/NET0131 ,
		_w310_,
		_w311_
	);
	LUT2 #(
		.INIT('h1)
	) name142 (
		\g1324_reg/NET0131 ,
		_w311_,
		_w312_
	);
	LUT2 #(
		.INIT('h8)
	) name143 (
		\g1324_reg/NET0131 ,
		_w311_,
		_w313_
	);
	LUT2 #(
		.INIT('h1)
	) name144 (
		\g1329_reg/NET0131 ,
		_w312_,
		_w314_
	);
	LUT2 #(
		.INIT('h4)
	) name145 (
		_w313_,
		_w314_,
		_w315_
	);
	LUT2 #(
		.INIT('h1)
	) name146 (
		_w305_,
		_w315_,
		_w316_
	);
	LUT2 #(
		.INIT('h8)
	) name147 (
		\g1342_reg/NET0131 ,
		\g1345_reg/NET0131 ,
		_w317_
	);
	LUT2 #(
		.INIT('h8)
	) name148 (
		\g1348_reg/NET0131 ,
		\g1351_reg/NET0131 ,
		_w318_
	);
	LUT2 #(
		.INIT('h8)
	) name149 (
		_w317_,
		_w318_,
		_w319_
	);
	LUT2 #(
		.INIT('h8)
	) name150 (
		_w172_,
		_w319_,
		_w320_
	);
	LUT2 #(
		.INIT('h1)
	) name151 (
		\g1354_reg/NET0131 ,
		_w320_,
		_w321_
	);
	LUT2 #(
		.INIT('h8)
	) name152 (
		\g1354_reg/NET0131 ,
		_w320_,
		_w322_
	);
	LUT2 #(
		.INIT('h2)
	) name153 (
		\g1247_reg/NET0131 ,
		_w321_,
		_w323_
	);
	LUT2 #(
		.INIT('h4)
	) name154 (
		_w322_,
		_w323_,
		_w324_
	);
	LUT2 #(
		.INIT('h1)
	) name155 (
		\g1363_reg/NET0131 ,
		\g1364_reg/NET0131 ,
		_w325_
	);
	LUT2 #(
		.INIT('h1)
	) name156 (
		\g1365_reg/NET0131 ,
		\g1366_reg/NET0131 ,
		_w326_
	);
	LUT2 #(
		.INIT('h1)
	) name157 (
		\g1367_reg/NET0131 ,
		\g1368_reg/NET0131 ,
		_w327_
	);
	LUT2 #(
		.INIT('h1)
	) name158 (
		\g1369_reg/NET0131 ,
		\g1370_reg/NET0131 ,
		_w328_
	);
	LUT2 #(
		.INIT('h1)
	) name159 (
		\g1371_reg/NET0131 ,
		\g1372_reg/NET0131 ,
		_w329_
	);
	LUT2 #(
		.INIT('h1)
	) name160 (
		\g1373_reg/NET0131 ,
		\g1374_reg/NET0131 ,
		_w330_
	);
	LUT2 #(
		.INIT('h4)
	) name161 (
		\g1375_reg/NET0131 ,
		_w330_,
		_w331_
	);
	LUT2 #(
		.INIT('h8)
	) name162 (
		_w328_,
		_w329_,
		_w332_
	);
	LUT2 #(
		.INIT('h8)
	) name163 (
		_w326_,
		_w327_,
		_w333_
	);
	LUT2 #(
		.INIT('h8)
	) name164 (
		_w325_,
		_w333_,
		_w334_
	);
	LUT2 #(
		.INIT('h8)
	) name165 (
		_w331_,
		_w332_,
		_w335_
	);
	LUT2 #(
		.INIT('h8)
	) name166 (
		_w334_,
		_w335_,
		_w336_
	);
	LUT2 #(
		.INIT('h8)
	) name167 (
		\g1325_reg/NET0131 ,
		\g1326_reg/NET0131 ,
		_w337_
	);
	LUT2 #(
		.INIT('h8)
	) name168 (
		\g1327_reg/NET0131 ,
		_w337_,
		_w338_
	);
	LUT2 #(
		.INIT('h8)
	) name169 (
		_w313_,
		_w338_,
		_w339_
	);
	LUT2 #(
		.INIT('h8)
	) name170 (
		\g1328_reg/NET0131 ,
		_w339_,
		_w340_
	);
	LUT2 #(
		.INIT('h1)
	) name171 (
		\g7504_pad ,
		_w340_,
		_w341_
	);
	LUT2 #(
		.INIT('h1)
	) name172 (
		\g1329_reg/NET0131 ,
		_w341_,
		_w342_
	);
	LUT2 #(
		.INIT('h8)
	) name173 (
		\g929_reg/NET0131 ,
		\g933_reg/NET0131 ,
		_w343_
	);
	LUT2 #(
		.INIT('h8)
	) name174 (
		\g871_reg/NET0131 ,
		_w343_,
		_w344_
	);
	LUT2 #(
		.INIT('h4)
	) name175 (
		\g889_reg/NET0131 ,
		_w344_,
		_w345_
	);
	LUT2 #(
		.INIT('h1)
	) name176 (
		\g785_pad ,
		_w345_,
		_w346_
	);
	LUT2 #(
		.INIT('h8)
	) name177 (
		\g1325_reg/NET0131 ,
		_w313_,
		_w347_
	);
	LUT2 #(
		.INIT('h1)
	) name178 (
		\g1326_reg/NET0131 ,
		\g1329_reg/NET0131 ,
		_w348_
	);
	LUT2 #(
		.INIT('h8)
	) name179 (
		_w347_,
		_w348_,
		_w349_
	);
	LUT2 #(
		.INIT('h1)
	) name180 (
		\g1329_reg/NET0131 ,
		_w347_,
		_w350_
	);
	LUT2 #(
		.INIT('h8)
	) name181 (
		\g1326_reg/NET0131 ,
		_w350_,
		_w351_
	);
	LUT2 #(
		.INIT('h1)
	) name182 (
		_w305_,
		_w349_,
		_w352_
	);
	LUT2 #(
		.INIT('h4)
	) name183 (
		_w351_,
		_w352_,
		_w353_
	);
	LUT2 #(
		.INIT('h8)
	) name184 (
		\g1134_reg/NET0131 ,
		_w203_,
		_w354_
	);
	LUT2 #(
		.INIT('h1)
	) name185 (
		\g1134_reg/NET0131 ,
		_w182_,
		_w355_
	);
	LUT2 #(
		.INIT('h2)
	) name186 (
		_w181_,
		_w183_,
		_w356_
	);
	LUT2 #(
		.INIT('h4)
	) name187 (
		_w355_,
		_w356_,
		_w357_
	);
	LUT2 #(
		.INIT('h1)
	) name188 (
		_w354_,
		_w357_,
		_w358_
	);
	LUT2 #(
		.INIT('h8)
	) name189 (
		\g1320_reg/NET0131 ,
		_w307_,
		_w359_
	);
	LUT2 #(
		.INIT('h1)
	) name190 (
		\g1321_reg/NET0131 ,
		_w359_,
		_w360_
	);
	LUT2 #(
		.INIT('h8)
	) name191 (
		\g1321_reg/NET0131 ,
		_w359_,
		_w361_
	);
	LUT2 #(
		.INIT('h1)
	) name192 (
		\g1329_reg/NET0131 ,
		_w360_,
		_w362_
	);
	LUT2 #(
		.INIT('h4)
	) name193 (
		_w361_,
		_w362_,
		_w363_
	);
	LUT2 #(
		.INIT('h1)
	) name194 (
		_w293_,
		_w363_,
		_w364_
	);
	LUT2 #(
		.INIT('h8)
	) name195 (
		\g1138_reg/NET0131 ,
		_w203_,
		_w365_
	);
	LUT2 #(
		.INIT('h1)
	) name196 (
		\g1138_reg/NET0131 ,
		_w183_,
		_w366_
	);
	LUT2 #(
		.INIT('h2)
	) name197 (
		_w181_,
		_w184_,
		_w367_
	);
	LUT2 #(
		.INIT('h4)
	) name198 (
		_w366_,
		_w367_,
		_w368_
	);
	LUT2 #(
		.INIT('h1)
	) name199 (
		_w365_,
		_w368_,
		_w369_
	);
	LUT2 #(
		.INIT('h8)
	) name200 (
		\g1130_reg/NET0131 ,
		_w203_,
		_w370_
	);
	LUT2 #(
		.INIT('h1)
	) name201 (
		\g1092_reg/NET0131 ,
		\g1130_reg/NET0131 ,
		_w371_
	);
	LUT2 #(
		.INIT('h1)
	) name202 (
		_w182_,
		_w371_,
		_w372_
	);
	LUT2 #(
		.INIT('h8)
	) name203 (
		_w181_,
		_w372_,
		_w373_
	);
	LUT2 #(
		.INIT('h1)
	) name204 (
		_w370_,
		_w373_,
		_w374_
	);
	LUT2 #(
		.INIT('h8)
	) name205 (
		\g1405_reg/NET0131 ,
		\g1408_reg/NET0131 ,
		_w375_
	);
	LUT2 #(
		.INIT('h1)
	) name206 (
		\g1231_reg/NET0131 ,
		\g1428_reg/NET0131 ,
		_w376_
	);
	LUT2 #(
		.INIT('h4)
	) name207 (
		_w375_,
		_w376_,
		_w377_
	);
	LUT2 #(
		.INIT('h8)
	) name208 (
		\g1412_reg/NET0131 ,
		\g1415_reg/NET0131 ,
		_w378_
	);
	LUT2 #(
		.INIT('h1)
	) name209 (
		\g1231_reg/NET0131 ,
		\g1430_reg/NET0131 ,
		_w379_
	);
	LUT2 #(
		.INIT('h4)
	) name210 (
		_w378_,
		_w379_,
		_w380_
	);
	LUT2 #(
		.INIT('h8)
	) name211 (
		\g1272_reg/NET0131 ,
		\g1307_reg/NET0131 ,
		_w381_
	);
	LUT2 #(
		.INIT('h8)
	) name212 (
		\g1276_reg/NET0131 ,
		_w381_,
		_w382_
	);
	LUT2 #(
		.INIT('h8)
	) name213 (
		\g1280_reg/NET0131 ,
		_w382_,
		_w383_
	);
	LUT2 #(
		.INIT('h1)
	) name214 (
		\g1280_reg/NET0131 ,
		_w382_,
		_w384_
	);
	LUT2 #(
		.INIT('h1)
	) name215 (
		\g1304_reg/NET0131 ,
		_w383_,
		_w385_
	);
	LUT2 #(
		.INIT('h4)
	) name216 (
		_w384_,
		_w385_,
		_w386_
	);
	LUT2 #(
		.INIT('h8)
	) name217 (
		\g1272_reg/NET0131 ,
		\g1276_reg/NET0131 ,
		_w387_
	);
	LUT2 #(
		.INIT('h8)
	) name218 (
		\g1280_reg/NET0131 ,
		\g1284_reg/NET0131 ,
		_w388_
	);
	LUT2 #(
		.INIT('h8)
	) name219 (
		_w387_,
		_w388_,
		_w389_
	);
	LUT2 #(
		.INIT('h8)
	) name220 (
		\g1307_reg/NET0131 ,
		_w389_,
		_w390_
	);
	LUT2 #(
		.INIT('h8)
	) name221 (
		\g1288_reg/NET0131 ,
		_w390_,
		_w391_
	);
	LUT2 #(
		.INIT('h1)
	) name222 (
		\g1292_reg/NET0131 ,
		_w391_,
		_w392_
	);
	LUT2 #(
		.INIT('h8)
	) name223 (
		\g1292_reg/NET0131 ,
		_w391_,
		_w393_
	);
	LUT2 #(
		.INIT('h1)
	) name224 (
		\g1304_reg/NET0131 ,
		_w392_,
		_w394_
	);
	LUT2 #(
		.INIT('h4)
	) name225 (
		_w393_,
		_w394_,
		_w395_
	);
	LUT2 #(
		.INIT('h8)
	) name226 (
		\g1300_reg/NET0131 ,
		_w393_,
		_w396_
	);
	LUT2 #(
		.INIT('h1)
	) name227 (
		\g1296_reg/NET0131 ,
		_w396_,
		_w397_
	);
	LUT2 #(
		.INIT('h8)
	) name228 (
		\g1296_reg/NET0131 ,
		_w396_,
		_w398_
	);
	LUT2 #(
		.INIT('h1)
	) name229 (
		\g1304_reg/NET0131 ,
		_w397_,
		_w399_
	);
	LUT2 #(
		.INIT('h4)
	) name230 (
		_w398_,
		_w399_,
		_w400_
	);
	LUT2 #(
		.INIT('h1)
	) name231 (
		\g1300_reg/NET0131 ,
		_w393_,
		_w401_
	);
	LUT2 #(
		.INIT('h1)
	) name232 (
		\g1304_reg/NET0131 ,
		_w396_,
		_w402_
	);
	LUT2 #(
		.INIT('h4)
	) name233 (
		_w401_,
		_w402_,
		_w403_
	);
	LUT2 #(
		.INIT('h1)
	) name234 (
		\g1276_reg/NET0131 ,
		_w381_,
		_w404_
	);
	LUT2 #(
		.INIT('h1)
	) name235 (
		\g1304_reg/NET0131 ,
		_w382_,
		_w405_
	);
	LUT2 #(
		.INIT('h4)
	) name236 (
		_w404_,
		_w405_,
		_w406_
	);
	LUT2 #(
		.INIT('h8)
	) name237 (
		\g1432_reg/NET0131 ,
		\g1439_reg/NET0131 ,
		_w407_
	);
	LUT2 #(
		.INIT('h1)
	) name238 (
		\g1430_reg/NET0131 ,
		_w407_,
		_w408_
	);
	LUT2 #(
		.INIT('h8)
	) name239 (
		\g1435_reg/NET0131 ,
		_w408_,
		_w409_
	);
	LUT2 #(
		.INIT('h8)
	) name240 (
		\g1435_reg/NET0131 ,
		\g1439_reg/NET0131 ,
		_w410_
	);
	LUT2 #(
		.INIT('h1)
	) name241 (
		\g1435_reg/NET0131 ,
		\g1439_reg/NET0131 ,
		_w411_
	);
	LUT2 #(
		.INIT('h1)
	) name242 (
		_w410_,
		_w411_,
		_w412_
	);
	LUT2 #(
		.INIT('h8)
	) name243 (
		_w408_,
		_w412_,
		_w413_
	);
	LUT2 #(
		.INIT('h4)
	) name244 (
		\g7507_pad ,
		_w407_,
		_w414_
	);
	LUT2 #(
		.INIT('h2)
	) name245 (
		\g7507_pad ,
		_w407_,
		_w415_
	);
	LUT2 #(
		.INIT('h1)
	) name246 (
		\g1430_reg/NET0131 ,
		_w414_,
		_w416_
	);
	LUT2 #(
		.INIT('h4)
	) name247 (
		_w415_,
		_w416_,
		_w417_
	);
	LUT2 #(
		.INIT('h1)
	) name248 (
		\g1432_reg/NET0131 ,
		_w410_,
		_w418_
	);
	LUT2 #(
		.INIT('h2)
	) name249 (
		_w408_,
		_w418_,
		_w419_
	);
	LUT2 #(
		.INIT('h1)
	) name250 (
		\g1284_reg/NET0131 ,
		_w383_,
		_w420_
	);
	LUT2 #(
		.INIT('h1)
	) name251 (
		\g1304_reg/NET0131 ,
		_w390_,
		_w421_
	);
	LUT2 #(
		.INIT('h4)
	) name252 (
		_w420_,
		_w421_,
		_w422_
	);
	LUT2 #(
		.INIT('h8)
	) name253 (
		\g1288_reg/NET0131 ,
		\g1292_reg/NET0131 ,
		_w423_
	);
	LUT2 #(
		.INIT('h8)
	) name254 (
		\g1296_reg/NET0131 ,
		\g1300_reg/NET0131 ,
		_w424_
	);
	LUT2 #(
		.INIT('h8)
	) name255 (
		_w423_,
		_w424_,
		_w425_
	);
	LUT2 #(
		.INIT('h1)
	) name256 (
		\g1288_reg/NET0131 ,
		_w390_,
		_w426_
	);
	LUT2 #(
		.INIT('h1)
	) name257 (
		_w391_,
		_w426_,
		_w427_
	);
	LUT2 #(
		.INIT('h1)
	) name258 (
		\g1304_reg/NET0131 ,
		_w425_,
		_w428_
	);
	LUT2 #(
		.INIT('h4)
	) name259 (
		_w427_,
		_w428_,
		_w429_
	);
	LUT2 #(
		.INIT('h8)
	) name260 (
		\g1211_reg/NET0131 ,
		\g1214_reg/NET0131 ,
		_w430_
	);
	LUT2 #(
		.INIT('h8)
	) name261 (
		\g1207_reg/NET0131 ,
		_w430_,
		_w431_
	);
	LUT2 #(
		.INIT('h8)
	) name262 (
		\g1217_reg/NET0131 ,
		_w431_,
		_w432_
	);
	LUT2 #(
		.INIT('h8)
	) name263 (
		\g1220_reg/NET0131 ,
		_w432_,
		_w433_
	);
	LUT2 #(
		.INIT('h1)
	) name264 (
		\g1223_reg/NET0131 ,
		_w433_,
		_w434_
	);
	LUT2 #(
		.INIT('h8)
	) name265 (
		\g1223_reg/NET0131 ,
		_w433_,
		_w435_
	);
	LUT2 #(
		.INIT('h1)
	) name266 (
		_w434_,
		_w435_,
		_w436_
	);
	LUT2 #(
		.INIT('h1)
	) name267 (
		\g1231_reg/NET0131 ,
		_w436_,
		_w437_
	);
	LUT2 #(
		.INIT('h1)
	) name268 (
		\g1272_reg/NET0131 ,
		\g1307_reg/NET0131 ,
		_w438_
	);
	LUT2 #(
		.INIT('h1)
	) name269 (
		\g1304_reg/NET0131 ,
		_w381_,
		_w439_
	);
	LUT2 #(
		.INIT('h4)
	) name270 (
		_w438_,
		_w439_,
		_w440_
	);
	LUT2 #(
		.INIT('h1)
	) name271 (
		\g1313_reg/NET0131 ,
		\g1329_reg/NET0131 ,
		_w441_
	);
	LUT2 #(
		.INIT('h1)
	) name272 (
		_w293_,
		_w441_,
		_w442_
	);
	LUT2 #(
		.INIT('h1)
	) name273 (
		\g1322_reg/NET0131 ,
		_w361_,
		_w443_
	);
	LUT2 #(
		.INIT('h1)
	) name274 (
		\g1329_reg/NET0131 ,
		_w310_,
		_w444_
	);
	LUT2 #(
		.INIT('h4)
	) name275 (
		_w443_,
		_w444_,
		_w445_
	);
	LUT2 #(
		.INIT('h1)
	) name276 (
		_w293_,
		_w445_,
		_w446_
	);
	LUT2 #(
		.INIT('h1)
	) name277 (
		\g1323_reg/NET0131 ,
		_w310_,
		_w447_
	);
	LUT2 #(
		.INIT('h1)
	) name278 (
		\g1329_reg/NET0131 ,
		_w311_,
		_w448_
	);
	LUT2 #(
		.INIT('h4)
	) name279 (
		_w447_,
		_w448_,
		_w449_
	);
	LUT2 #(
		.INIT('h1)
	) name280 (
		_w293_,
		_w449_,
		_w450_
	);
	LUT2 #(
		.INIT('h1)
	) name281 (
		\g1325_reg/NET0131 ,
		_w313_,
		_w451_
	);
	LUT2 #(
		.INIT('h2)
	) name282 (
		_w350_,
		_w451_,
		_w452_
	);
	LUT2 #(
		.INIT('h1)
	) name283 (
		_w305_,
		_w452_,
		_w453_
	);
	LUT2 #(
		.INIT('h1)
	) name284 (
		\g1319_reg/NET0131 ,
		_w296_,
		_w454_
	);
	LUT2 #(
		.INIT('h1)
	) name285 (
		\g1329_reg/NET0131 ,
		_w307_,
		_w455_
	);
	LUT2 #(
		.INIT('h4)
	) name286 (
		_w454_,
		_w455_,
		_w456_
	);
	LUT2 #(
		.INIT('h1)
	) name287 (
		_w293_,
		_w456_,
		_w457_
	);
	LUT2 #(
		.INIT('h8)
	) name288 (
		_w313_,
		_w337_,
		_w458_
	);
	LUT2 #(
		.INIT('h1)
	) name289 (
		\g1327_reg/NET0131 ,
		_w458_,
		_w459_
	);
	LUT2 #(
		.INIT('h1)
	) name290 (
		\g1329_reg/NET0131 ,
		_w339_,
		_w460_
	);
	LUT2 #(
		.INIT('h4)
	) name291 (
		_w459_,
		_w460_,
		_w461_
	);
	LUT2 #(
		.INIT('h1)
	) name292 (
		_w305_,
		_w461_,
		_w462_
	);
	LUT2 #(
		.INIT('h1)
	) name293 (
		\g1494_reg/NET0131 ,
		_w302_,
		_w463_
	);
	LUT2 #(
		.INIT('h1)
	) name294 (
		_w215_,
		_w463_,
		_w464_
	);
	LUT2 #(
		.INIT('h1)
	) name295 (
		\g1499_reg/NET0131 ,
		_w215_,
		_w465_
	);
	LUT2 #(
		.INIT('h1)
	) name296 (
		_w278_,
		_w465_,
		_w466_
	);
	LUT2 #(
		.INIT('h1)
	) name297 (
		\g1313_reg/NET0131 ,
		\g1317_reg/NET0131 ,
		_w467_
	);
	LUT2 #(
		.INIT('h1)
	) name298 (
		\g1329_reg/NET0131 ,
		_w294_,
		_w468_
	);
	LUT2 #(
		.INIT('h4)
	) name299 (
		_w467_,
		_w468_,
		_w469_
	);
	LUT2 #(
		.INIT('h1)
	) name300 (
		_w293_,
		_w469_,
		_w470_
	);
	LUT2 #(
		.INIT('h2)
	) name301 (
		\g950_reg/NET0131 ,
		_w197_,
		_w471_
	);
	LUT2 #(
		.INIT('h1)
	) name302 (
		_w211_,
		_w471_,
		_w472_
	);
	LUT2 #(
		.INIT('h1)
	) name303 (
		\g1320_reg/NET0131 ,
		_w307_,
		_w473_
	);
	LUT2 #(
		.INIT('h1)
	) name304 (
		\g1329_reg/NET0131 ,
		_w359_,
		_w474_
	);
	LUT2 #(
		.INIT('h4)
	) name305 (
		_w473_,
		_w474_,
		_w475_
	);
	LUT2 #(
		.INIT('h1)
	) name306 (
		_w293_,
		_w475_,
		_w476_
	);
	LUT2 #(
		.INIT('h8)
	) name307 (
		\g1450_reg/NET0131 ,
		\g1454_reg/NET0131 ,
		_w477_
	);
	LUT2 #(
		.INIT('h1)
	) name308 (
		\g1307_reg/NET0131 ,
		_w477_,
		_w478_
	);
	LUT2 #(
		.INIT('h8)
	) name309 (
		\g1444_reg/NET0131 ,
		_w478_,
		_w479_
	);
	LUT2 #(
		.INIT('h2)
	) name310 (
		\g1444_reg/NET0131 ,
		\g1450_reg/NET0131 ,
		_w480_
	);
	LUT2 #(
		.INIT('h4)
	) name311 (
		\g1444_reg/NET0131 ,
		\g1450_reg/NET0131 ,
		_w481_
	);
	LUT2 #(
		.INIT('h4)
	) name312 (
		\g1454_reg/NET0131 ,
		_w481_,
		_w482_
	);
	LUT2 #(
		.INIT('h1)
	) name313 (
		_w480_,
		_w482_,
		_w483_
	);
	LUT2 #(
		.INIT('h1)
	) name314 (
		\g1307_reg/NET0131 ,
		_w483_,
		_w484_
	);
	LUT2 #(
		.INIT('h4)
	) name315 (
		\g1405_reg/NET0131 ,
		_w376_,
		_w485_
	);
	LUT2 #(
		.INIT('h4)
	) name316 (
		\g1412_reg/NET0131 ,
		_w379_,
		_w486_
	);
	LUT2 #(
		.INIT('h4)
	) name317 (
		\g1307_reg/NET0131 ,
		\g1416_reg/NET0131 ,
		_w487_
	);
	LUT2 #(
		.INIT('h4)
	) name318 (
		\g1421_reg/NET0131 ,
		_w487_,
		_w488_
	);
	LUT2 #(
		.INIT('h8)
	) name319 (
		\g1444_reg/NET0131 ,
		\g1450_reg/NET0131 ,
		_w489_
	);
	LUT2 #(
		.INIT('h1)
	) name320 (
		\g1454_reg/NET0131 ,
		_w489_,
		_w490_
	);
	LUT2 #(
		.INIT('h2)
	) name321 (
		_w478_,
		_w490_,
		_w491_
	);
	LUT2 #(
		.INIT('h2)
	) name322 (
		\g7508_pad ,
		_w414_,
		_w492_
	);
	LUT2 #(
		.INIT('h4)
	) name323 (
		\g7508_pad ,
		_w414_,
		_w493_
	);
	LUT2 #(
		.INIT('h1)
	) name324 (
		\g1430_reg/NET0131 ,
		_w492_,
		_w494_
	);
	LUT2 #(
		.INIT('h4)
	) name325 (
		_w493_,
		_w494_,
		_w495_
	);
	LUT2 #(
		.INIT('h1)
	) name326 (
		\g104_reg/NET0131 ,
		\g1339_reg/NET0131 ,
		_w496_
	);
	LUT2 #(
		.INIT('h1)
	) name327 (
		_w170_,
		_w496_,
		_w497_
	);
	LUT2 #(
		.INIT('h1)
	) name328 (
		\g1330_reg/NET0131 ,
		\g1333_reg/NET0131 ,
		_w498_
	);
	LUT2 #(
		.INIT('h8)
	) name329 (
		\g104_reg/NET0131 ,
		\g1339_reg/NET0131 ,
		_w499_
	);
	LUT2 #(
		.INIT('h1)
	) name330 (
		_w498_,
		_w499_,
		_w500_
	);
	LUT2 #(
		.INIT('h1)
	) name331 (
		\g104_reg/NET0131 ,
		\g1336_reg/NET0131 ,
		_w501_
	);
	LUT2 #(
		.INIT('h1)
	) name332 (
		\g1342_reg/NET0131 ,
		\g1345_reg/NET0131 ,
		_w502_
	);
	LUT2 #(
		.INIT('h1)
	) name333 (
		\g1348_reg/NET0131 ,
		\g1351_reg/NET0131 ,
		_w503_
	);
	LUT2 #(
		.INIT('h1)
	) name334 (
		\g1354_reg/NET0131 ,
		\g1357_reg/NET0131 ,
		_w504_
	);
	LUT2 #(
		.INIT('h4)
	) name335 (
		\g1360_reg/NET0131 ,
		_w504_,
		_w505_
	);
	LUT2 #(
		.INIT('h8)
	) name336 (
		_w502_,
		_w503_,
		_w506_
	);
	LUT2 #(
		.INIT('h8)
	) name337 (
		_w501_,
		_w506_,
		_w507_
	);
	LUT2 #(
		.INIT('h8)
	) name338 (
		_w505_,
		_w507_,
		_w508_
	);
	LUT2 #(
		.INIT('h8)
	) name339 (
		\g1354_reg/NET0131 ,
		\g1357_reg/NET0131 ,
		_w509_
	);
	LUT2 #(
		.INIT('h8)
	) name340 (
		\g104_reg/NET0131 ,
		\g1336_reg/NET0131 ,
		_w510_
	);
	LUT2 #(
		.INIT('h8)
	) name341 (
		\g1360_reg/NET0131 ,
		_w510_,
		_w511_
	);
	LUT2 #(
		.INIT('h8)
	) name342 (
		_w509_,
		_w511_,
		_w512_
	);
	LUT2 #(
		.INIT('h8)
	) name343 (
		_w319_,
		_w512_,
		_w513_
	);
	LUT2 #(
		.INIT('h1)
	) name344 (
		_w508_,
		_w513_,
		_w514_
	);
	LUT2 #(
		.INIT('h1)
	) name345 (
		_w497_,
		_w500_,
		_w515_
	);
	LUT2 #(
		.INIT('h4)
	) name346 (
		_w514_,
		_w515_,
		_w516_
	);
	LUT2 #(
		.INIT('h8)
	) name347 (
		\g1077_reg/NET0131 ,
		\g2888_pad ,
		_w517_
	);
	LUT2 #(
		.INIT('h8)
	) name348 (
		\g1158_reg/NET0131 ,
		\g652_reg/NET0131 ,
		_w518_
	);
	LUT2 #(
		.INIT('h8)
	) name349 (
		\g1176_reg/NET0131 ,
		_w518_,
		_w519_
	);
	LUT2 #(
		.INIT('h1)
	) name350 (
		_w517_,
		_w519_,
		_w520_
	);
	LUT2 #(
		.INIT('h2)
	) name351 (
		\g1247_reg/NET0131 ,
		_w170_,
		_w521_
	);
	LUT2 #(
		.INIT('h4)
	) name352 (
		_w498_,
		_w521_,
		_w522_
	);
	LUT2 #(
		.INIT('h1)
	) name353 (
		\g1351_reg/NET0131 ,
		_w176_,
		_w523_
	);
	LUT2 #(
		.INIT('h2)
	) name354 (
		\g1247_reg/NET0131 ,
		_w320_,
		_w524_
	);
	LUT2 #(
		.INIT('h4)
	) name355 (
		_w523_,
		_w524_,
		_w525_
	);
	LUT2 #(
		.INIT('h4)
	) name356 (
		\g785_pad ,
		\g866_reg/NET0131 ,
		_w526_
	);
	LUT2 #(
		.INIT('h8)
	) name357 (
		\g889_reg/NET0131 ,
		_w526_,
		_w527_
	);
	LUT2 #(
		.INIT('h8)
	) name358 (
		\g1179_reg/NET0131 ,
		_w518_,
		_w528_
	);
	LUT2 #(
		.INIT('h2)
	) name359 (
		\g2888_pad ,
		_w528_,
		_w529_
	);
	LUT2 #(
		.INIT('h4)
	) name360 (
		\g2888_pad ,
		_w528_,
		_w530_
	);
	LUT2 #(
		.INIT('h1)
	) name361 (
		_w529_,
		_w530_,
		_w531_
	);
	LUT2 #(
		.INIT('h1)
	) name362 (
		_w517_,
		_w531_,
		_w532_
	);
	LUT2 #(
		.INIT('h4)
	) name363 (
		\g1176_reg/NET0131 ,
		\g1944_pad ,
		_w533_
	);
	LUT2 #(
		.INIT('h2)
	) name364 (
		\g1080_pad ,
		\g1944_pad ,
		_w534_
	);
	LUT2 #(
		.INIT('h1)
	) name365 (
		_w533_,
		_w534_,
		_w535_
	);
	LUT2 #(
		.INIT('h1)
	) name366 (
		\g1224_reg/NET0131 ,
		_w435_,
		_w536_
	);
	LUT2 #(
		.INIT('h8)
	) name367 (
		\g1223_reg/NET0131 ,
		\g1224_reg/NET0131 ,
		_w537_
	);
	LUT2 #(
		.INIT('h8)
	) name368 (
		_w433_,
		_w537_,
		_w538_
	);
	LUT2 #(
		.INIT('h1)
	) name369 (
		_w536_,
		_w538_,
		_w539_
	);
	LUT2 #(
		.INIT('h1)
	) name370 (
		\g1231_reg/NET0131 ,
		_w539_,
		_w540_
	);
	LUT2 #(
		.INIT('h1)
	) name371 (
		_w496_,
		_w499_,
		_w541_
	);
	LUT2 #(
		.INIT('h2)
	) name372 (
		_w498_,
		_w541_,
		_w542_
	);
	LUT2 #(
		.INIT('h4)
	) name373 (
		_w514_,
		_w542_,
		_w543_
	);
	LUT2 #(
		.INIT('h1)
	) name374 (
		\g1257_reg/NET0131 ,
		\g1263_reg/NET0131 ,
		_w544_
	);
	LUT2 #(
		.INIT('h8)
	) name375 (
		\g1225_reg/NET0131 ,
		_w537_,
		_w545_
	);
	LUT2 #(
		.INIT('h8)
	) name376 (
		\g1227_reg/NET0131 ,
		\g1228_reg/NET0131 ,
		_w546_
	);
	LUT2 #(
		.INIT('h2)
	) name377 (
		\g1226_reg/NET0131 ,
		\g1229_reg/NET0131 ,
		_w547_
	);
	LUT2 #(
		.INIT('h8)
	) name378 (
		\g1230_reg/NET0131 ,
		_w547_,
		_w548_
	);
	LUT2 #(
		.INIT('h8)
	) name379 (
		_w546_,
		_w548_,
		_w549_
	);
	LUT2 #(
		.INIT('h8)
	) name380 (
		_w545_,
		_w549_,
		_w550_
	);
	LUT2 #(
		.INIT('h4)
	) name381 (
		_w544_,
		_w550_,
		_w551_
	);
	LUT2 #(
		.INIT('h2)
	) name382 (
		\g1247_reg/NET0131 ,
		_w551_,
		_w552_
	);
	LUT2 #(
		.INIT('h2)
	) name383 (
		\g1253_reg/NET0131 ,
		_w552_,
		_w553_
	);
	LUT2 #(
		.INIT('h1)
	) name384 (
		\g1339_reg/NET0131 ,
		_w171_,
		_w554_
	);
	LUT2 #(
		.INIT('h2)
	) name385 (
		\g1247_reg/NET0131 ,
		_w172_,
		_w555_
	);
	LUT2 #(
		.INIT('h4)
	) name386 (
		_w554_,
		_w555_,
		_w556_
	);
	LUT2 #(
		.INIT('h1)
	) name387 (
		\g1220_reg/NET0131 ,
		_w432_,
		_w557_
	);
	LUT2 #(
		.INIT('h1)
	) name388 (
		_w433_,
		_w557_,
		_w558_
	);
	LUT2 #(
		.INIT('h1)
	) name389 (
		\g1231_reg/NET0131 ,
		_w558_,
		_w559_
	);
	LUT2 #(
		.INIT('h1)
	) name390 (
		\g1416_reg/NET0131 ,
		\g1421_reg/NET0131 ,
		_w560_
	);
	LUT2 #(
		.INIT('h1)
	) name391 (
		\g1307_reg/NET0131 ,
		_w560_,
		_w561_
	);
	LUT2 #(
		.INIT('h2)
	) name392 (
		\g1247_reg/NET0131 ,
		\g1330_reg/NET0131 ,
		_w562_
	);
	LUT2 #(
		.INIT('h1)
	) name393 (
		\g1336_reg/NET0131 ,
		_w170_,
		_w563_
	);
	LUT2 #(
		.INIT('h2)
	) name394 (
		\g1247_reg/NET0131 ,
		_w171_,
		_w564_
	);
	LUT2 #(
		.INIT('h4)
	) name395 (
		_w563_,
		_w564_,
		_w565_
	);
	LUT2 #(
		.INIT('h1)
	) name396 (
		\g1342_reg/NET0131 ,
		_w172_,
		_w566_
	);
	LUT2 #(
		.INIT('h2)
	) name397 (
		\g1247_reg/NET0131 ,
		_w173_,
		_w567_
	);
	LUT2 #(
		.INIT('h4)
	) name398 (
		_w566_,
		_w567_,
		_w568_
	);
	LUT2 #(
		.INIT('h8)
	) name399 (
		_w389_,
		_w425_,
		_w569_
	);
	LUT2 #(
		.INIT('h8)
	) name400 (
		\g104_reg/NET0131 ,
		_w569_,
		_w570_
	);
	LUT2 #(
		.INIT('h1)
	) name401 (
		\g104_reg/NET0131 ,
		\g1272_reg/NET0131 ,
		_w571_
	);
	LUT2 #(
		.INIT('h1)
	) name402 (
		\g1276_reg/NET0131 ,
		\g1280_reg/NET0131 ,
		_w572_
	);
	LUT2 #(
		.INIT('h1)
	) name403 (
		\g1284_reg/NET0131 ,
		\g1288_reg/NET0131 ,
		_w573_
	);
	LUT2 #(
		.INIT('h1)
	) name404 (
		\g1292_reg/NET0131 ,
		\g1296_reg/NET0131 ,
		_w574_
	);
	LUT2 #(
		.INIT('h4)
	) name405 (
		\g1300_reg/NET0131 ,
		_w574_,
		_w575_
	);
	LUT2 #(
		.INIT('h8)
	) name406 (
		_w572_,
		_w573_,
		_w576_
	);
	LUT2 #(
		.INIT('h8)
	) name407 (
		_w571_,
		_w576_,
		_w577_
	);
	LUT2 #(
		.INIT('h8)
	) name408 (
		_w575_,
		_w577_,
		_w578_
	);
	LUT2 #(
		.INIT('h1)
	) name409 (
		_w570_,
		_w578_,
		_w579_
	);
	LUT2 #(
		.INIT('h2)
	) name410 (
		\g104_reg/NET0131 ,
		_w197_,
		_w580_
	);
	LUT2 #(
		.INIT('h1)
	) name411 (
		_w211_,
		_w580_,
		_w581_
	);
	LUT2 #(
		.INIT('h1)
	) name412 (
		\g1268_reg/NET0131 ,
		\g1269_reg/NET0131 ,
		_w582_
	);
	LUT2 #(
		.INIT('h1)
	) name413 (
		_w197_,
		_w198_,
		_w583_
	);
	LUT2 #(
		.INIT('h1)
	) name414 (
		_w344_,
		_w583_,
		_w584_
	);
	LUT2 #(
		.INIT('h1)
	) name415 (
		\g1073_reg/NET0131 ,
		\g1179_reg/NET0131 ,
		_w585_
	);
	LUT2 #(
		.INIT('h1)
	) name416 (
		\g4370_pad ,
		\g4371_pad ,
		_w586_
	);
	LUT2 #(
		.INIT('h1)
	) name417 (
		\g4372_pad ,
		\g4373_pad ,
		_w587_
	);
	LUT2 #(
		.INIT('h8)
	) name418 (
		_w586_,
		_w587_,
		_w588_
	);
	LUT2 #(
		.INIT('h8)
	) name419 (
		_w585_,
		_w588_,
		_w589_
	);
	LUT2 #(
		.INIT('h8)
	) name420 (
		\g1263_reg/NET0131 ,
		_w550_,
		_w590_
	);
	LUT2 #(
		.INIT('h8)
	) name421 (
		\g1257_reg/NET0131 ,
		_w550_,
		_w591_
	);
	LUT2 #(
		.INIT('h8)
	) name422 (
		\g1266_reg/NET0131 ,
		_w550_,
		_w592_
	);
	LUT2 #(
		.INIT('h1)
	) name423 (
		\g1217_reg/NET0131 ,
		_w431_,
		_w593_
	);
	LUT2 #(
		.INIT('h1)
	) name424 (
		_w432_,
		_w593_,
		_w594_
	);
	LUT2 #(
		.INIT('h1)
	) name425 (
		\g1231_reg/NET0131 ,
		_w594_,
		_w595_
	);
	LUT2 #(
		.INIT('h1)
	) name426 (
		\g1223_reg/NET0131 ,
		\g1224_reg/NET0131 ,
		_w596_
	);
	LUT2 #(
		.INIT('h1)
	) name427 (
		\g1225_reg/NET0131 ,
		\g1226_reg/NET0131 ,
		_w597_
	);
	LUT2 #(
		.INIT('h1)
	) name428 (
		\g1227_reg/NET0131 ,
		\g1228_reg/NET0131 ,
		_w598_
	);
	LUT2 #(
		.INIT('h1)
	) name429 (
		\g1229_reg/NET0131 ,
		\g1230_reg/NET0131 ,
		_w599_
	);
	LUT2 #(
		.INIT('h8)
	) name430 (
		_w598_,
		_w599_,
		_w600_
	);
	LUT2 #(
		.INIT('h8)
	) name431 (
		_w596_,
		_w597_,
		_w601_
	);
	LUT2 #(
		.INIT('h8)
	) name432 (
		_w600_,
		_w601_,
		_w602_
	);
	LUT2 #(
		.INIT('h8)
	) name433 (
		\g1207_reg/NET0131 ,
		\g1211_reg/NET0131 ,
		_w603_
	);
	LUT2 #(
		.INIT('h1)
	) name434 (
		\g1207_reg/NET0131 ,
		\g1211_reg/NET0131 ,
		_w604_
	);
	LUT2 #(
		.INIT('h1)
	) name435 (
		_w603_,
		_w604_,
		_w605_
	);
	LUT2 #(
		.INIT('h1)
	) name436 (
		\g1231_reg/NET0131 ,
		_w605_,
		_w606_
	);
	LUT2 #(
		.INIT('h4)
	) name437 (
		\g1231_reg/NET0131 ,
		\g2662_pad ,
		_w607_
	);
	LUT2 #(
		.INIT('h1)
	) name438 (
		\g1214_reg/NET0131 ,
		_w603_,
		_w608_
	);
	LUT2 #(
		.INIT('h4)
	) name439 (
		_w431_,
		_w607_,
		_w609_
	);
	LUT2 #(
		.INIT('h4)
	) name440 (
		_w608_,
		_w609_,
		_w610_
	);
	LUT2 #(
		.INIT('h1)
	) name441 (
		\g871_reg/NET0131 ,
		_w343_,
		_w611_
	);
	LUT2 #(
		.INIT('h1)
	) name442 (
		_w344_,
		_w611_,
		_w612_
	);
	LUT2 #(
		.INIT('h2)
	) name443 (
		\g1207_reg/NET0131 ,
		\g1231_reg/NET0131 ,
		_w613_
	);
	LUT2 #(
		.INIT('h2)
	) name444 (
		\g104_reg/NET0131 ,
		\g1211_reg/NET0131 ,
		_w614_
	);
	LUT2 #(
		.INIT('h4)
	) name445 (
		\g104_reg/NET0131 ,
		\g1211_reg/NET0131 ,
		_w615_
	);
	LUT2 #(
		.INIT('h1)
	) name446 (
		_w614_,
		_w615_,
		_w616_
	);
	LUT2 #(
		.INIT('h2)
	) name447 (
		\g104_reg/NET0131 ,
		\g1214_reg/NET0131 ,
		_w617_
	);
	LUT2 #(
		.INIT('h4)
	) name448 (
		\g104_reg/NET0131 ,
		\g1214_reg/NET0131 ,
		_w618_
	);
	LUT2 #(
		.INIT('h1)
	) name449 (
		_w617_,
		_w618_,
		_w619_
	);
	LUT2 #(
		.INIT('h2)
	) name450 (
		\g104_reg/NET0131 ,
		\g1220_reg/NET0131 ,
		_w620_
	);
	LUT2 #(
		.INIT('h4)
	) name451 (
		\g104_reg/NET0131 ,
		\g1220_reg/NET0131 ,
		_w621_
	);
	LUT2 #(
		.INIT('h1)
	) name452 (
		_w620_,
		_w621_,
		_w622_
	);
	LUT2 #(
		.INIT('h2)
	) name453 (
		\g104_reg/NET0131 ,
		\g1207_reg/NET0131 ,
		_w623_
	);
	LUT2 #(
		.INIT('h4)
	) name454 (
		\g104_reg/NET0131 ,
		\g1207_reg/NET0131 ,
		_w624_
	);
	LUT2 #(
		.INIT('h1)
	) name455 (
		_w623_,
		_w624_,
		_w625_
	);
	LUT2 #(
		.INIT('h2)
	) name456 (
		\g104_reg/NET0131 ,
		\g1225_reg/NET0131 ,
		_w626_
	);
	LUT2 #(
		.INIT('h4)
	) name457 (
		\g104_reg/NET0131 ,
		\g1225_reg/NET0131 ,
		_w627_
	);
	LUT2 #(
		.INIT('h1)
	) name458 (
		_w626_,
		_w627_,
		_w628_
	);
	LUT2 #(
		.INIT('h2)
	) name459 (
		\g104_reg/NET0131 ,
		\g1227_reg/NET0131 ,
		_w629_
	);
	LUT2 #(
		.INIT('h4)
	) name460 (
		\g104_reg/NET0131 ,
		\g1227_reg/NET0131 ,
		_w630_
	);
	LUT2 #(
		.INIT('h1)
	) name461 (
		_w629_,
		_w630_,
		_w631_
	);
	LUT2 #(
		.INIT('h2)
	) name462 (
		\g104_reg/NET0131 ,
		\g1228_reg/NET0131 ,
		_w632_
	);
	LUT2 #(
		.INIT('h4)
	) name463 (
		\g104_reg/NET0131 ,
		\g1228_reg/NET0131 ,
		_w633_
	);
	LUT2 #(
		.INIT('h1)
	) name464 (
		_w632_,
		_w633_,
		_w634_
	);
	LUT2 #(
		.INIT('h2)
	) name465 (
		\g104_reg/NET0131 ,
		\g1230_reg/NET0131 ,
		_w635_
	);
	LUT2 #(
		.INIT('h4)
	) name466 (
		\g104_reg/NET0131 ,
		\g1230_reg/NET0131 ,
		_w636_
	);
	LUT2 #(
		.INIT('h1)
	) name467 (
		_w635_,
		_w636_,
		_w637_
	);
	LUT2 #(
		.INIT('h2)
	) name468 (
		\g104_reg/NET0131 ,
		\g1223_reg/NET0131 ,
		_w638_
	);
	LUT2 #(
		.INIT('h4)
	) name469 (
		\g104_reg/NET0131 ,
		\g1223_reg/NET0131 ,
		_w639_
	);
	LUT2 #(
		.INIT('h1)
	) name470 (
		_w638_,
		_w639_,
		_w640_
	);
	LUT2 #(
		.INIT('h2)
	) name471 (
		\g104_reg/NET0131 ,
		\g1224_reg/NET0131 ,
		_w641_
	);
	LUT2 #(
		.INIT('h4)
	) name472 (
		\g104_reg/NET0131 ,
		\g1224_reg/NET0131 ,
		_w642_
	);
	LUT2 #(
		.INIT('h1)
	) name473 (
		_w641_,
		_w642_,
		_w643_
	);
	LUT2 #(
		.INIT('h2)
	) name474 (
		\g104_reg/NET0131 ,
		\g1226_reg/NET0131 ,
		_w644_
	);
	LUT2 #(
		.INIT('h4)
	) name475 (
		\g104_reg/NET0131 ,
		\g1226_reg/NET0131 ,
		_w645_
	);
	LUT2 #(
		.INIT('h1)
	) name476 (
		_w644_,
		_w645_,
		_w646_
	);
	LUT2 #(
		.INIT('h8)
	) name477 (
		\g1217_reg/NET0131 ,
		\g1220_reg/NET0131 ,
		_w647_
	);
	LUT2 #(
		.INIT('h4)
	) name478 (
		\g1211_reg/NET0131 ,
		_w647_,
		_w648_
	);
	LUT2 #(
		.INIT('h8)
	) name479 (
		\g1207_reg/NET0131 ,
		\g1214_reg/NET0131 ,
		_w649_
	);
	LUT2 #(
		.INIT('h8)
	) name480 (
		_w648_,
		_w649_,
		_w650_
	);
	LUT2 #(
		.INIT('h4)
	) name481 (
		\g1207_reg/NET0131 ,
		\g1214_reg/NET0131 ,
		_w651_
	);
	LUT2 #(
		.INIT('h8)
	) name482 (
		_w648_,
		_w651_,
		_w652_
	);
	LUT2 #(
		.INIT('h8)
	) name483 (
		\g1211_reg/NET0131 ,
		_w647_,
		_w653_
	);
	LUT2 #(
		.INIT('h8)
	) name484 (
		_w651_,
		_w653_,
		_w654_
	);
	LUT2 #(
		.INIT('h2)
	) name485 (
		\g104_reg/NET0131 ,
		\g1217_reg/NET0131 ,
		_w655_
	);
	LUT2 #(
		.INIT('h4)
	) name486 (
		\g104_reg/NET0131 ,
		\g1217_reg/NET0131 ,
		_w656_
	);
	LUT2 #(
		.INIT('h1)
	) name487 (
		_w655_,
		_w656_,
		_w657_
	);
	LUT2 #(
		.INIT('h2)
	) name488 (
		\g104_reg/NET0131 ,
		\g1229_reg/NET0131 ,
		_w658_
	);
	LUT2 #(
		.INIT('h4)
	) name489 (
		\g104_reg/NET0131 ,
		\g1229_reg/NET0131 ,
		_w659_
	);
	LUT2 #(
		.INIT('h1)
	) name490 (
		_w658_,
		_w659_,
		_w660_
	);
	LUT2 #(
		.INIT('h1)
	) name491 (
		\g929_reg/NET0131 ,
		\g933_reg/NET0131 ,
		_w661_
	);
	LUT2 #(
		.INIT('h1)
	) name492 (
		_w343_,
		_w661_,
		_w662_
	);
	LUT2 #(
		.INIT('h1)
	) name493 (
		\g1217_reg/NET0131 ,
		\g1220_reg/NET0131 ,
		_w663_
	);
	LUT2 #(
		.INIT('h8)
	) name494 (
		_w430_,
		_w663_,
		_w664_
	);
	LUT2 #(
		.INIT('h8)
	) name495 (
		\g1454_reg/NET0131 ,
		_w480_,
		_w665_
	);
	LUT2 #(
		.INIT('h2)
	) name496 (
		\g942_reg/NET0131 ,
		_w198_,
		_w666_
	);
	LUT2 #(
		.INIT('h1)
	) name497 (
		\g1122_reg/NET0131 ,
		_w236_,
		_w667_
	);
	LUT2 #(
		.INIT('h8)
	) name498 (
		\g1114_reg/NET0131 ,
		\g1118_reg/NET0131 ,
		_w668_
	);
	LUT2 #(
		.INIT('h8)
	) name499 (
		\g1122_reg/NET0131 ,
		_w668_,
		_w669_
	);
	LUT2 #(
		.INIT('h8)
	) name500 (
		_w233_,
		_w669_,
		_w670_
	);
	LUT2 #(
		.INIT('h1)
	) name501 (
		_w667_,
		_w670_,
		_w671_
	);
	LUT2 #(
		.INIT('h1)
	) name502 (
		\g1097_reg/NET0131 ,
		_w671_,
		_w672_
	);
	LUT2 #(
		.INIT('h8)
	) name503 (
		\g1126_reg/NET0131 ,
		_w670_,
		_w673_
	);
	LUT2 #(
		.INIT('h1)
	) name504 (
		\g1126_reg/NET0131 ,
		_w670_,
		_w674_
	);
	LUT2 #(
		.INIT('h1)
	) name505 (
		_w673_,
		_w674_,
		_w675_
	);
	LUT2 #(
		.INIT('h1)
	) name506 (
		\g1097_reg/NET0131 ,
		_w675_,
		_w676_
	);
	LUT2 #(
		.INIT('h8)
	) name507 (
		\g1110_reg/NET0131 ,
		\g1126_reg/NET0131 ,
		_w677_
	);
	LUT2 #(
		.INIT('h8)
	) name508 (
		\g1142_reg/NET0131 ,
		_w677_,
		_w678_
	);
	LUT2 #(
		.INIT('h8)
	) name509 (
		_w669_,
		_w678_,
		_w679_
	);
	LUT2 #(
		.INIT('h8)
	) name510 (
		_w231_,
		_w679_,
		_w680_
	);
	LUT2 #(
		.INIT('h1)
	) name511 (
		\g1166_reg/NET0131 ,
		\g7423_pad ,
		_w681_
	);
	LUT2 #(
		.INIT('h1)
	) name512 (
		\g7424_pad ,
		\g7425_pad ,
		_w682_
	);
	LUT2 #(
		.INIT('h8)
	) name513 (
		_w681_,
		_w682_,
		_w683_
	);
	LUT2 #(
		.INIT('h4)
	) name514 (
		_w680_,
		_w683_,
		_w684_
	);
	LUT2 #(
		.INIT('h8)
	) name515 (
		_w545_,
		_w649_,
		_w685_
	);
	LUT2 #(
		.INIT('h8)
	) name516 (
		_w653_,
		_w685_,
		_w686_
	);
	LUT2 #(
		.INIT('h8)
	) name517 (
		\g1226_reg/NET0131 ,
		_w686_,
		_w687_
	);
	LUT2 #(
		.INIT('h8)
	) name518 (
		\g1227_reg/NET0131 ,
		_w687_,
		_w688_
	);
	LUT2 #(
		.INIT('h1)
	) name519 (
		\g1228_reg/NET0131 ,
		_w688_,
		_w689_
	);
	LUT2 #(
		.INIT('h8)
	) name520 (
		_w546_,
		_w687_,
		_w690_
	);
	LUT2 #(
		.INIT('h1)
	) name521 (
		_w689_,
		_w690_,
		_w691_
	);
	LUT2 #(
		.INIT('h1)
	) name522 (
		\g1231_reg/NET0131 ,
		_w691_,
		_w692_
	);
	LUT2 #(
		.INIT('h8)
	) name523 (
		\g1229_reg/NET0131 ,
		_w546_,
		_w693_
	);
	LUT2 #(
		.INIT('h8)
	) name524 (
		_w687_,
		_w693_,
		_w694_
	);
	LUT2 #(
		.INIT('h1)
	) name525 (
		\g1229_reg/NET0131 ,
		_w690_,
		_w695_
	);
	LUT2 #(
		.INIT('h2)
	) name526 (
		_w607_,
		_w694_,
		_w696_
	);
	LUT2 #(
		.INIT('h4)
	) name527 (
		_w695_,
		_w696_,
		_w697_
	);
	LUT2 #(
		.INIT('h8)
	) name528 (
		_w216_,
		_w224_,
		_w698_
	);
	LUT2 #(
		.INIT('h8)
	) name529 (
		\g1462_reg/NET0131 ,
		_w698_,
		_w699_
	);
	LUT2 #(
		.INIT('h1)
	) name530 (
		\g1467_reg/NET0131 ,
		_w699_,
		_w700_
	);
	LUT2 #(
		.INIT('h8)
	) name531 (
		\g1467_reg/NET0131 ,
		_w699_,
		_w701_
	);
	LUT2 #(
		.INIT('h1)
	) name532 (
		_w221_,
		_w700_,
		_w702_
	);
	LUT2 #(
		.INIT('h4)
	) name533 (
		_w701_,
		_w702_,
		_w703_
	);
	LUT2 #(
		.INIT('h2)
	) name534 (
		\g1486_reg/NET0131 ,
		_w221_,
		_w704_
	);
	LUT2 #(
		.INIT('h4)
	) name535 (
		\g1486_reg/NET0131 ,
		_w221_,
		_w705_
	);
	LUT2 #(
		.INIT('h1)
	) name536 (
		_w704_,
		_w705_,
		_w706_
	);
	LUT2 #(
		.INIT('h1)
	) name537 (
		\g1227_reg/NET0131 ,
		_w687_,
		_w707_
	);
	LUT2 #(
		.INIT('h1)
	) name538 (
		_w688_,
		_w707_,
		_w708_
	);
	LUT2 #(
		.INIT('h1)
	) name539 (
		\g1231_reg/NET0131 ,
		_w708_,
		_w709_
	);
	LUT2 #(
		.INIT('h1)
	) name540 (
		\g1519_reg/NET0131 ,
		_w225_,
		_w710_
	);
	LUT2 #(
		.INIT('h1)
	) name541 (
		_w221_,
		_w698_,
		_w711_
	);
	LUT2 #(
		.INIT('h4)
	) name542 (
		_w710_,
		_w711_,
		_w712_
	);
	LUT2 #(
		.INIT('h1)
	) name543 (
		\g1462_reg/NET0131 ,
		_w698_,
		_w713_
	);
	LUT2 #(
		.INIT('h1)
	) name544 (
		_w221_,
		_w699_,
		_w714_
	);
	LUT2 #(
		.INIT('h4)
	) name545 (
		_w713_,
		_w714_,
		_w715_
	);
	LUT2 #(
		.INIT('h1)
	) name546 (
		\g1226_reg/NET0131 ,
		_w686_,
		_w716_
	);
	LUT2 #(
		.INIT('h1)
	) name547 (
		_w687_,
		_w716_,
		_w717_
	);
	LUT2 #(
		.INIT('h1)
	) name548 (
		\g1231_reg/NET0131 ,
		_w717_,
		_w718_
	);
	LUT2 #(
		.INIT('h2)
	) name549 (
		\g1225_reg/NET0131 ,
		_w538_,
		_w719_
	);
	LUT2 #(
		.INIT('h4)
	) name550 (
		\g1225_reg/NET0131 ,
		_w538_,
		_w720_
	);
	LUT2 #(
		.INIT('h1)
	) name551 (
		\g1231_reg/NET0131 ,
		_w719_,
		_w721_
	);
	LUT2 #(
		.INIT('h4)
	) name552 (
		_w720_,
		_w721_,
		_w722_
	);
	LUT2 #(
		.INIT('h1)
	) name553 (
		\g1230_reg/NET0131 ,
		_w694_,
		_w723_
	);
	LUT2 #(
		.INIT('h8)
	) name554 (
		\g1230_reg/NET0131 ,
		_w694_,
		_w724_
	);
	LUT2 #(
		.INIT('h2)
	) name555 (
		\g2662_pad ,
		_w723_,
		_w725_
	);
	LUT2 #(
		.INIT('h4)
	) name556 (
		_w724_,
		_w725_,
		_w726_
	);
	LUT2 #(
		.INIT('h1)
	) name557 (
		\g1231_reg/NET0131 ,
		_w726_,
		_w727_
	);
	LUT2 #(
		.INIT('h8)
	) name558 (
		_w320_,
		_w509_,
		_w728_
	);
	LUT2 #(
		.INIT('h1)
	) name559 (
		\g1357_reg/NET0131 ,
		_w322_,
		_w729_
	);
	LUT2 #(
		.INIT('h2)
	) name560 (
		\g1247_reg/NET0131 ,
		_w728_,
		_w730_
	);
	LUT2 #(
		.INIT('h4)
	) name561 (
		_w729_,
		_w730_,
		_w731_
	);
	LUT2 #(
		.INIT('h8)
	) name562 (
		\g1041_reg/NET0131 ,
		_w268_,
		_w732_
	);
	LUT2 #(
		.INIT('h2)
	) name563 (
		_w181_,
		_w732_,
		_w733_
	);
	LUT2 #(
		.INIT('h1)
	) name564 (
		_w203_,
		_w733_,
		_w734_
	);
	LUT2 #(
		.INIT('h2)
	) name565 (
		\g1045_reg/NET0131 ,
		_w734_,
		_w735_
	);
	LUT2 #(
		.INIT('h4)
	) name566 (
		\g1045_reg/NET0131 ,
		_w181_,
		_w736_
	);
	LUT2 #(
		.INIT('h8)
	) name567 (
		_w732_,
		_w736_,
		_w737_
	);
	LUT2 #(
		.INIT('h1)
	) name568 (
		_w735_,
		_w737_,
		_w738_
	);
	LUT2 #(
		.INIT('h8)
	) name569 (
		\g1065_reg/NET0131 ,
		_w203_,
		_w739_
	);
	LUT2 #(
		.INIT('h1)
	) name570 (
		\g1065_reg/NET0131 ,
		_w192_,
		_w740_
	);
	LUT2 #(
		.INIT('h2)
	) name571 (
		_w181_,
		_w193_,
		_w741_
	);
	LUT2 #(
		.INIT('h4)
	) name572 (
		_w740_,
		_w741_,
		_w742_
	);
	LUT2 #(
		.INIT('h1)
	) name573 (
		_w739_,
		_w742_,
		_w743_
	);
	LUT2 #(
		.INIT('h8)
	) name574 (
		\g1053_reg/NET0131 ,
		_w203_,
		_w744_
	);
	LUT2 #(
		.INIT('h1)
	) name575 (
		\g1053_reg/NET0131 ,
		_w206_,
		_w745_
	);
	LUT2 #(
		.INIT('h8)
	) name576 (
		\g1053_reg/NET0131 ,
		_w206_,
		_w746_
	);
	LUT2 #(
		.INIT('h2)
	) name577 (
		_w181_,
		_w746_,
		_w747_
	);
	LUT2 #(
		.INIT('h4)
	) name578 (
		_w745_,
		_w747_,
		_w748_
	);
	LUT2 #(
		.INIT('h1)
	) name579 (
		_w744_,
		_w748_,
		_w749_
	);
	LUT2 #(
		.INIT('h1)
	) name580 (
		\g1345_reg/NET0131 ,
		_w173_,
		_w750_
	);
	LUT2 #(
		.INIT('h2)
	) name581 (
		\g1247_reg/NET0131 ,
		_w174_,
		_w751_
	);
	LUT2 #(
		.INIT('h4)
	) name582 (
		_w750_,
		_w751_,
		_w752_
	);
	LUT2 #(
		.INIT('h1)
	) name583 (
		\g1142_reg/NET0131 ,
		_w673_,
		_w753_
	);
	LUT2 #(
		.INIT('h8)
	) name584 (
		\g1142_reg/NET0131 ,
		_w673_,
		_w754_
	);
	LUT2 #(
		.INIT('h1)
	) name585 (
		\g1097_reg/NET0131 ,
		_w753_,
		_w755_
	);
	LUT2 #(
		.INIT('h4)
	) name586 (
		_w754_,
		_w755_,
		_w756_
	);
	LUT2 #(
		.INIT('h1)
	) name587 (
		\g1069_reg/NET0131 ,
		_w194_,
		_w757_
	);
	LUT2 #(
		.INIT('h2)
	) name588 (
		\g1069_reg/NET0131 ,
		_w203_,
		_w758_
	);
	LUT2 #(
		.INIT('h4)
	) name589 (
		_w741_,
		_w758_,
		_w759_
	);
	LUT2 #(
		.INIT('h1)
	) name590 (
		_w757_,
		_w759_,
		_w760_
	);
	LUT2 #(
		.INIT('h8)
	) name591 (
		\g1057_reg/NET0131 ,
		_w746_,
		_w761_
	);
	LUT2 #(
		.INIT('h8)
	) name592 (
		\g1061_reg/NET0131 ,
		_w181_,
		_w762_
	);
	LUT2 #(
		.INIT('h4)
	) name593 (
		_w761_,
		_w762_,
		_w763_
	);
	LUT2 #(
		.INIT('h8)
	) name594 (
		\g1061_reg/NET0131 ,
		_w203_,
		_w764_
	);
	LUT2 #(
		.INIT('h2)
	) name595 (
		\g1057_reg/NET0131 ,
		\g1061_reg/NET0131 ,
		_w765_
	);
	LUT2 #(
		.INIT('h8)
	) name596 (
		_w181_,
		_w765_,
		_w766_
	);
	LUT2 #(
		.INIT('h8)
	) name597 (
		_w746_,
		_w766_,
		_w767_
	);
	LUT2 #(
		.INIT('h1)
	) name598 (
		_w764_,
		_w767_,
		_w768_
	);
	LUT2 #(
		.INIT('h4)
	) name599 (
		_w763_,
		_w768_,
		_w769_
	);
	LUT2 #(
		.INIT('h1)
	) name600 (
		\g1360_reg/NET0131 ,
		_w728_,
		_w770_
	);
	LUT2 #(
		.INIT('h8)
	) name601 (
		\g1360_reg/NET0131 ,
		_w728_,
		_w771_
	);
	LUT2 #(
		.INIT('h2)
	) name602 (
		\g1247_reg/NET0131 ,
		_w770_,
		_w772_
	);
	LUT2 #(
		.INIT('h4)
	) name603 (
		_w771_,
		_w772_,
		_w773_
	);
	LUT2 #(
		.INIT('h8)
	) name604 (
		_w181_,
		_w746_,
		_w774_
	);
	LUT2 #(
		.INIT('h1)
	) name605 (
		\g1057_reg/NET0131 ,
		_w774_,
		_w775_
	);
	LUT2 #(
		.INIT('h2)
	) name606 (
		\g1057_reg/NET0131 ,
		_w203_,
		_w776_
	);
	LUT2 #(
		.INIT('h4)
	) name607 (
		_w747_,
		_w776_,
		_w777_
	);
	LUT2 #(
		.INIT('h1)
	) name608 (
		_w775_,
		_w777_,
		_w778_
	);
	LUT2 #(
		.INIT('h1)
	) name609 (
		\g1328_reg/NET0131 ,
		_w339_,
		_w779_
	);
	LUT2 #(
		.INIT('h1)
	) name610 (
		\g1329_reg/NET0131 ,
		_w340_,
		_w780_
	);
	LUT2 #(
		.INIT('h4)
	) name611 (
		_w779_,
		_w780_,
		_w781_
	);
	LUT2 #(
		.INIT('h1)
	) name612 (
		_w305_,
		_w781_,
		_w782_
	);
	LUT2 #(
		.INIT('h2)
	) name613 (
		\g1041_reg/NET0131 ,
		_w734_,
		_w783_
	);
	LUT2 #(
		.INIT('h8)
	) name614 (
		_w268_,
		_w733_,
		_w784_
	);
	LUT2 #(
		.INIT('h1)
	) name615 (
		_w783_,
		_w784_,
		_w785_
	);
	LUT2 #(
		.INIT('h1)
	) name616 (
		\g1472_reg/NET0131 ,
		_w701_,
		_w786_
	);
	LUT2 #(
		.INIT('h8)
	) name617 (
		\g1472_reg/NET0131 ,
		_w701_,
		_w787_
	);
	LUT2 #(
		.INIT('h1)
	) name618 (
		_w221_,
		_w786_,
		_w788_
	);
	LUT2 #(
		.INIT('h4)
	) name619 (
		_w787_,
		_w788_,
		_w789_
	);
	LUT2 #(
		.INIT('h1)
	) name620 (
		\g2_reg/NET0131 ,
		\g962_pad ,
		_w790_
	);
	LUT2 #(
		.INIT('h1)
	) name621 (
		\g1189_reg/NET0131 ,
		\g7505_pad ,
		_w791_
	);
	LUT2 #(
		.INIT('h8)
	) name622 (
		\g1405_reg/NET0131 ,
		\g1412_reg/NET0131 ,
		_w792_
	);
	assign \g1006_pad  = 1'b0;
	assign \g1158_reg/P0001  = \g1158_reg/NET0131 ;
	assign \g1252_reg/P0001  = \g1252_reg/NET0131 ;
	assign \g1260_reg/P0001  = \g1260_reg/NET0131 ;
	assign \g1416_reg/NET0131_syn_2  = \g1416_reg/NET0131 ;
	assign \g17/_0_  = _w178_ ;
	assign \g19189/_0_  = _w196_ ;
	assign \g19252/_0_  = _w200_ ;
	assign \g19253/_0_  = _w209_ ;
	assign \g19273/_3_  = _w212_ ;
	assign \g19284/_0_  = _w228_ ;
	assign \g19285/_0_  = _w238_ ;
	assign \g19295/_3_  = _w240_ ;
	assign \g19302/_0_  = _w244_ ;
	assign \g19303/_0_  = _w247_ ;
	assign \g19304/_0_  = _w250_ ;
	assign \g19308/_0_  = _w253_ ;
	assign \g19309/_0_  = _w260_ ;
	assign \g19310/_0_  = _w265_ ;
	assign \g19321/_0_  = _w271_ ;
	assign \g19326/_3_  = _w273_ ;
	assign \g19331/_0_  = _w277_ ;
	assign \g19341/_0_  = _w281_ ;
	assign \g19366/_0_  = _w286_ ;
	assign \g19372/_3_  = _w288_ ;
	assign \g19385/_0_  = _w292_ ;
	assign \g19386/_0_  = _w299_ ;
	assign \g19387/_0_  = _w301_ ;
	assign \g19388/_0_  = _w304_ ;
	assign \g19389/_0_  = _w316_ ;
	assign \g19390/_0_  = _w324_ ;
	assign \g19392/_0_  = _w336_ ;
	assign \g19393/_0_  = _w342_ ;
	assign \g19394/_0_  = _w346_ ;
	assign \g19398/_0_  = _w353_ ;
	assign \g19399/_0_  = _w358_ ;
	assign \g19400/_0_  = _w364_ ;
	assign \g19401/_0_  = _w369_ ;
	assign \g19403/_0_  = _w374_ ;
	assign \g19405/_0_  = _w377_ ;
	assign \g19406/_0_  = _w380_ ;
	assign \g19437/_0_  = _w386_ ;
	assign \g19438/_0_  = _w395_ ;
	assign \g19445/_0_  = _w400_ ;
	assign \g19446/_0_  = _w403_ ;
	assign \g19450/_3_  = _w406_ ;
	assign \g19472/_0_  = _w409_ ;
	assign \g19473/_0_  = _w413_ ;
	assign \g19474/_0_  = _w417_ ;
	assign \g19476/_0_  = _w419_ ;
	assign \g19484/_0_  = _w422_ ;
	assign \g19485/_0_  = _w429_ ;
	assign \g19492/_0_  = _w437_ ;
	assign \g19493/_0_  = _w440_ ;
	assign \g19499/_0_  = _w442_ ;
	assign \g19500/_0_  = _w446_ ;
	assign \g19501/_0_  = _w450_ ;
	assign \g19502/_0_  = _w453_ ;
	assign \g19503/_0_  = _w457_ ;
	assign \g19504/_0_  = _w462_ ;
	assign \g19507/_3_  = _w464_ ;
	assign \g19508/_3_  = _w466_ ;
	assign \g19512/_3_  = _w470_ ;
	assign \g19513/_3_  = _w472_ ;
	assign \g19514/_3_  = _w476_ ;
	assign \g19528/_0_  = _w479_ ;
	assign \g19529/_0_  = _w484_ ;
	assign \g19534/_0_  = _w485_ ;
	assign \g19535/_0_  = _w486_ ;
	assign \g19536/_0_  = _w488_ ;
	assign \g19538/_0_  = _w491_ ;
	assign \g19542/_0_  = _w495_ ;
	assign \g19560/_0_  = _w516_ ;
	assign \g19563/_0_  = _w520_ ;
	assign \g19565/_0_  = _w522_ ;
	assign \g19567/_0_  = _w525_ ;
	assign \g19569/_1_  = _w527_ ;
	assign \g19572/_0_  = _w532_ ;
	assign \g19574/_3_  = _w535_ ;
	assign \g19614/_0_  = _w540_ ;
	assign \g19615/_0_  = _w543_ ;
	assign \g19620/_0_  = _w553_ ;
	assign \g19626/_0_  = _w556_ ;
	assign \g19629/_0_  = _w559_ ;
	assign \g19631/_0_  = _w561_ ;
	assign \g19666/_0_  = _w562_ ;
	assign \g19667/_0_  = _w565_ ;
	assign \g19669/_0_  = _w568_ ;
	assign \g19677/_0_  = _w579_ ;
	assign \g19690/_3_  = _w581_ ;
	assign \g19721/_0_  = _w582_ ;
	assign \g19723/_0_  = _w584_ ;
	assign \g19723/_1_  = _w344_ ;
	assign \g19725/_2_  = _w589_ ;
	assign \g19751/_0_  = _w590_ ;
	assign \g19752/_0_  = _w591_ ;
	assign \g19753/_0_  = _w592_ ;
	assign \g19755/_0_  = _w595_ ;
	assign \g19815/_0_  = _w602_ ;
	assign \g19821/_0_  = _w606_ ;
	assign \g19822/_0_  = _w610_ ;
	assign \g19833/_0_  = _w612_ ;
	assign \g19877/_0_  = _w613_ ;
	assign \g19898/_0_  = _w616_ ;
	assign \g19899/_0_  = _w619_ ;
	assign \g19900/_0_  = _w622_ ;
	assign \g19901/_0_  = _w625_ ;
	assign \g19908/_0_  = _w628_ ;
	assign \g19927/_0_  = _w631_ ;
	assign \g19928/_0_  = _w634_ ;
	assign \g19930/_0_  = _w637_ ;
	assign \g19931/_0_  = _w640_ ;
	assign \g19932/_0_  = _w643_ ;
	assign \g19934/_0_  = _w646_ ;
	assign \g19992/_0_  = _w650_ ;
	assign \g19993/_0_  = _w652_ ;
	assign \g20002/_0_  = _w654_ ;
	assign \g20008/_0_  = _w657_ ;
	assign \g20010/_0_  = _w660_ ;
	assign \g20016/_0_  = _w662_ ;
	assign \g20110/_0_  = _w664_ ;
	assign \g20117/_0_  = _w482_ ;
	assign \g20118/_0_  = _w665_ ;
	assign \g20131/_0_  = _w666_ ;
	assign \g20246/_0_  = \g929_reg/NET0131 ;
	assign \g20704/_0_  = _w672_ ;
	assign \g20722/_0_  = _w676_ ;
	assign \g20731/_0_  = _w684_ ;
	assign \g20732/_2_  = _w680_ ;
	assign \g20870/_0_  = _w692_ ;
	assign \g20883/_0_  = _w697_ ;
	assign \g20931/_0_  = _w703_ ;
	assign \g20951/_0_  = _w706_ ;
	assign \g20969/_0_  = _w709_ ;
	assign \g20989/_0_  = _w552_ ;
	assign \g21/_2_  = _w712_ ;
	assign \g21070/_0_  = _w715_ ;
	assign \g21108/_0_  = _w718_ ;
	assign \g21122/_0_  = _w722_ ;
	assign \g21152/_0_  = _w727_ ;
	assign \g21191/_0_  = _w731_ ;
	assign \g21279/_0_  = _w738_ ;
	assign \g21316/_0_  = _w743_ ;
	assign \g21323/_0_  = _w749_ ;
	assign \g21349/_3_  = _w569_ ;
	assign \g21352/_3_  = _w752_ ;
	assign \g21464/_0_  = _w756_ ;
	assign \g21472/_0_  = _w760_ ;
	assign \g21484/_0_  = _w769_ ;
	assign \g21510/_0_  = _w773_ ;
	assign \g21517/_0_  = _w778_ ;
	assign \g21608/_0_  = _w782_ ;
	assign \g21625/_0_  = _w785_ ;
	assign \g21644/_1_  = _w789_ ;
	assign \g4655_pad  = _w583_ ;
	assign \g6850_pad  = \g43_pad ;
	assign \g6895_pad  = 1'b0;
	assign \g7048_pad  = \g944_reg/NET0131 ;
	assign \g7103_pad  = _w790_ ;
	assign \g7731_pad  = _w791_ ;
	assign \g7732_pad  = \g1486_reg/NET0131 ;
	assign \g8219_pad  = \g1432_reg/NET0131 ;
	assign \g8663_pad  = _w792_ ;
endmodule;