module top (\G0_pad , \G10_pad , \G11_pad , \G12_pad , \G13_pad , \G1_pad , \G29_reg/NET0131 , \G2_pad , \G30_reg/NET0131 , \G31_reg/NET0131 , \G32_reg/NET0131 , \G33_reg/NET0131 , \G34_reg/NET0131 , \G35_reg/NET0131 , \G36_reg/NET0131 , \G37_reg/NET0131 , \G38_reg/NET0131 , \G39_reg/NET0131 , \G3_pad , \G40_reg/NET0131 , \G41_reg/NET0131 , \G42_reg/NET0131 , \G43_reg/NET0131 , \G44_reg/NET0131 , \G46_reg/NET0131 , \G4_pad , \G5_pad , \G6_pad , \G7_pad , \G8_pad , \G9_pad , \G532_pad , \G537_pad , \G539_pad , \G542_pad , \G546_pad , \G547_pad , \G548_pad , \G549_pad , \G550_pad , \G551_pad , \G552_pad , \_al_n0 , \_al_n1 , \g1667/_3_ , \g1737/_0_ , \g1744/_0_ , \g1787/_0_ , \g1811/_0_ , \g1830/_0_ , \g1831/_0_ , \g1846/_0_ , \g1852/_0_ , \g1866/_0_ , \g19/_2_ , \g1931/_0_ , \g1945/_0_ , \g2014/_0_ , \g2015/_0_ , \g2643/_0_ , \g2859/_1_ , \g3397/_2_ , \g3546/_0_ , \g3606/_3_ );
	input \G0_pad  ;
	input \G10_pad  ;
	input \G11_pad  ;
	input \G12_pad  ;
	input \G13_pad  ;
	input \G1_pad  ;
	input \G29_reg/NET0131  ;
	input \G2_pad  ;
	input \G30_reg/NET0131  ;
	input \G31_reg/NET0131  ;
	input \G32_reg/NET0131  ;
	input \G33_reg/NET0131  ;
	input \G34_reg/NET0131  ;
	input \G35_reg/NET0131  ;
	input \G36_reg/NET0131  ;
	input \G37_reg/NET0131  ;
	input \G38_reg/NET0131  ;
	input \G39_reg/NET0131  ;
	input \G3_pad  ;
	input \G40_reg/NET0131  ;
	input \G41_reg/NET0131  ;
	input \G42_reg/NET0131  ;
	input \G43_reg/NET0131  ;
	input \G44_reg/NET0131  ;
	input \G46_reg/NET0131  ;
	input \G4_pad  ;
	input \G5_pad  ;
	input \G6_pad  ;
	input \G7_pad  ;
	input \G8_pad  ;
	input \G9_pad  ;
	output \G532_pad  ;
	output \G537_pad  ;
	output \G539_pad  ;
	output \G542_pad  ;
	output \G546_pad  ;
	output \G547_pad  ;
	output \G548_pad  ;
	output \G549_pad  ;
	output \G550_pad  ;
	output \G551_pad  ;
	output \G552_pad  ;
	output \_al_n0  ;
	output \_al_n1  ;
	output \g1667/_3_  ;
	output \g1737/_0_  ;
	output \g1744/_0_  ;
	output \g1787/_0_  ;
	output \g1811/_0_  ;
	output \g1830/_0_  ;
	output \g1831/_0_  ;
	output \g1846/_0_  ;
	output \g1852/_0_  ;
	output \g1866/_0_  ;
	output \g19/_2_  ;
	output \g1931/_0_  ;
	output \g1945/_0_  ;
	output \g2014/_0_  ;
	output \g2015/_0_  ;
	output \g2643/_0_  ;
	output \g2859/_1_  ;
	output \g3397/_2_  ;
	output \g3546/_0_  ;
	output \g3606/_3_  ;
	wire _w311_ ;
	wire _w310_ ;
	wire _w309_ ;
	wire _w308_ ;
	wire _w307_ ;
	wire _w306_ ;
	wire _w305_ ;
	wire _w304_ ;
	wire _w303_ ;
	wire _w302_ ;
	wire _w301_ ;
	wire _w300_ ;
	wire _w299_ ;
	wire _w298_ ;
	wire _w297_ ;
	wire _w296_ ;
	wire _w295_ ;
	wire _w294_ ;
	wire _w293_ ;
	wire _w292_ ;
	wire _w291_ ;
	wire _w290_ ;
	wire _w159_ ;
	wire _w158_ ;
	wire _w157_ ;
	wire _w156_ ;
	wire _w155_ ;
	wire _w154_ ;
	wire _w153_ ;
	wire _w152_ ;
	wire _w151_ ;
	wire _w149_ ;
	wire _w148_ ;
	wire _w147_ ;
	wire _w146_ ;
	wire _w145_ ;
	wire _w144_ ;
	wire _w143_ ;
	wire _w142_ ;
	wire _w141_ ;
	wire _w140_ ;
	wire _w139_ ;
	wire _w138_ ;
	wire _w137_ ;
	wire _w136_ ;
	wire _w135_ ;
	wire _w134_ ;
	wire _w133_ ;
	wire _w132_ ;
	wire _w131_ ;
	wire _w130_ ;
	wire _w129_ ;
	wire _w128_ ;
	wire _w127_ ;
	wire _w126_ ;
	wire _w125_ ;
	wire _w124_ ;
	wire _w123_ ;
	wire _w122_ ;
	wire _w121_ ;
	wire _w120_ ;
	wire _w119_ ;
	wire _w118_ ;
	wire _w117_ ;
	wire _w116_ ;
	wire _w115_ ;
	wire _w114_ ;
	wire _w113_ ;
	wire _w112_ ;
	wire _w111_ ;
	wire _w110_ ;
	wire _w109_ ;
	wire _w108_ ;
	wire _w107_ ;
	wire _w106_ ;
	wire _w105_ ;
	wire _w104_ ;
	wire _w103_ ;
	wire _w102_ ;
	wire _w101_ ;
	wire _w100_ ;
	wire _w99_ ;
	wire _w98_ ;
	wire _w97_ ;
	wire _w96_ ;
	wire _w95_ ;
	wire _w94_ ;
	wire _w93_ ;
	wire _w92_ ;
	wire _w61_ ;
	wire _w60_ ;
	wire _w59_ ;
	wire _w58_ ;
	wire _w57_ ;
	wire _w56_ ;
	wire _w55_ ;
	wire _w54_ ;
	wire _w53_ ;
	wire _w51_ ;
	wire _w50_ ;
	wire _w49_ ;
	wire _w48_ ;
	wire _w47_ ;
	wire _w46_ ;
	wire _w52_ ;
	wire _w150_ ;
	wire _w23_ ;
	wire _w280_ ;
	wire _w82_ ;
	wire _w36_ ;
	wire _w34_ ;
	wire _w35_ ;
	wire _w37_ ;
	wire _w38_ ;
	wire _w39_ ;
	wire _w40_ ;
	wire _w41_ ;
	wire _w42_ ;
	wire _w43_ ;
	wire _w44_ ;
	wire _w45_ ;
	wire _w62_ ;
	wire _w63_ ;
	wire _w64_ ;
	wire _w65_ ;
	wire _w66_ ;
	wire _w67_ ;
	wire _w68_ ;
	wire _w69_ ;
	wire _w70_ ;
	wire _w71_ ;
	wire _w72_ ;
	wire _w73_ ;
	wire _w74_ ;
	wire _w75_ ;
	wire _w76_ ;
	wire _w77_ ;
	wire _w78_ ;
	wire _w79_ ;
	wire _w80_ ;
	wire _w81_ ;
	wire _w83_ ;
	wire _w84_ ;
	wire _w85_ ;
	wire _w86_ ;
	wire _w87_ ;
	wire _w88_ ;
	wire _w89_ ;
	wire _w90_ ;
	wire _w91_ ;
	wire _w160_ ;
	wire _w161_ ;
	wire _w162_ ;
	wire _w163_ ;
	wire _w164_ ;
	wire _w165_ ;
	wire _w166_ ;
	wire _w167_ ;
	wire _w168_ ;
	wire _w169_ ;
	wire _w170_ ;
	wire _w171_ ;
	wire _w172_ ;
	wire _w173_ ;
	wire _w174_ ;
	wire _w175_ ;
	wire _w176_ ;
	wire _w177_ ;
	wire _w178_ ;
	wire _w179_ ;
	wire _w180_ ;
	wire _w181_ ;
	wire _w182_ ;
	wire _w183_ ;
	wire _w184_ ;
	wire _w185_ ;
	wire _w186_ ;
	wire _w187_ ;
	wire _w188_ ;
	wire _w189_ ;
	wire _w190_ ;
	wire _w191_ ;
	wire _w192_ ;
	wire _w193_ ;
	wire _w194_ ;
	wire _w195_ ;
	wire _w196_ ;
	wire _w197_ ;
	wire _w198_ ;
	wire _w199_ ;
	wire _w200_ ;
	wire _w201_ ;
	wire _w202_ ;
	wire _w203_ ;
	wire _w204_ ;
	wire _w205_ ;
	wire _w206_ ;
	wire _w207_ ;
	wire _w208_ ;
	wire _w209_ ;
	wire _w210_ ;
	wire _w211_ ;
	wire _w212_ ;
	wire _w213_ ;
	wire _w214_ ;
	wire _w215_ ;
	wire _w216_ ;
	wire _w217_ ;
	wire _w218_ ;
	wire _w219_ ;
	wire _w220_ ;
	wire _w221_ ;
	wire _w222_ ;
	wire _w223_ ;
	wire _w224_ ;
	wire _w225_ ;
	wire _w226_ ;
	wire _w227_ ;
	wire _w228_ ;
	wire _w229_ ;
	wire _w230_ ;
	wire _w231_ ;
	wire _w232_ ;
	wire _w233_ ;
	wire _w234_ ;
	wire _w235_ ;
	wire _w236_ ;
	wire _w237_ ;
	wire _w238_ ;
	wire _w239_ ;
	wire _w240_ ;
	wire _w241_ ;
	wire _w242_ ;
	wire _w243_ ;
	wire _w244_ ;
	wire _w245_ ;
	wire _w246_ ;
	wire _w247_ ;
	wire _w248_ ;
	wire _w249_ ;
	wire _w250_ ;
	wire _w251_ ;
	wire _w252_ ;
	wire _w253_ ;
	wire _w254_ ;
	wire _w255_ ;
	wire _w256_ ;
	wire _w257_ ;
	wire _w258_ ;
	wire _w259_ ;
	wire _w260_ ;
	wire _w261_ ;
	wire _w262_ ;
	wire _w263_ ;
	wire _w264_ ;
	wire _w265_ ;
	wire _w266_ ;
	wire _w267_ ;
	wire _w268_ ;
	wire _w269_ ;
	wire _w270_ ;
	wire _w271_ ;
	wire _w272_ ;
	wire _w273_ ;
	wire _w274_ ;
	wire _w275_ ;
	wire _w276_ ;
	wire _w277_ ;
	wire _w278_ ;
	wire _w279_ ;
	wire _w281_ ;
	wire _w282_ ;
	wire _w283_ ;
	wire _w284_ ;
	wire _w285_ ;
	wire _w286_ ;
	wire _w287_ ;
	wire _w288_ ;
	wire _w289_ ;
	LUT1 #(
		.INIT('h1)
	) name0 (
		\G41_reg/NET0131 ,
		_w23_
	);
	LUT3 #(
		.INIT('h80)
	) name1 (
		\G11_pad ,
		\G8_pad ,
		\G9_pad ,
		_w34_
	);
	LUT2 #(
		.INIT('h8)
	) name2 (
		\G10_pad ,
		\G7_pad ,
		_w35_
	);
	LUT3 #(
		.INIT('h20)
	) name3 (
		\G30_reg/NET0131 ,
		\G7_pad ,
		\G8_pad ,
		_w36_
	);
	LUT3 #(
		.INIT('h40)
	) name4 (
		\G10_pad ,
		\G7_pad ,
		\G9_pad ,
		_w37_
	);
	LUT4 #(
		.INIT('h0045)
	) name5 (
		_w36_,
		_w34_,
		_w35_,
		_w37_,
		_w38_
	);
	LUT3 #(
		.INIT('h51)
	) name6 (
		\G13_pad ,
		\G32_reg/NET0131 ,
		_w38_,
		_w39_
	);
	LUT4 #(
		.INIT('h0800)
	) name7 (
		\G3_pad ,
		\G4_pad ,
		\G5_pad ,
		\G6_pad ,
		_w40_
	);
	LUT2 #(
		.INIT('h8)
	) name8 (
		\G8_pad ,
		\G9_pad ,
		_w41_
	);
	LUT4 #(
		.INIT('h0240)
	) name9 (
		\G10_pad ,
		\G7_pad ,
		\G8_pad ,
		\G9_pad ,
		_w42_
	);
	LUT3 #(
		.INIT('h10)
	) name10 (
		\G10_pad ,
		\G7_pad ,
		\G9_pad ,
		_w43_
	);
	LUT4 #(
		.INIT('hedbf)
	) name11 (
		\G10_pad ,
		\G7_pad ,
		\G8_pad ,
		\G9_pad ,
		_w44_
	);
	LUT3 #(
		.INIT('h08)
	) name12 (
		\G11_pad ,
		_w40_,
		_w44_,
		_w45_
	);
	LUT2 #(
		.INIT('h2)
	) name13 (
		\G36_reg/NET0131 ,
		\G6_pad ,
		_w46_
	);
	LUT3 #(
		.INIT('h80)
	) name14 (
		\G4_pad ,
		\G5_pad ,
		\G6_pad ,
		_w47_
	);
	LUT4 #(
		.INIT('h8000)
	) name15 (
		\G11_pad ,
		\G4_pad ,
		\G5_pad ,
		\G6_pad ,
		_w48_
	);
	LUT4 #(
		.INIT('h5450)
	) name16 (
		\G3_pad ,
		_w42_,
		_w46_,
		_w48_,
		_w49_
	);
	LUT3 #(
		.INIT('h54)
	) name17 (
		\G2_pad ,
		_w45_,
		_w49_,
		_w50_
	);
	LUT3 #(
		.INIT('h80)
	) name18 (
		\G3_pad ,
		_w39_,
		_w50_,
		_w51_
	);
	LUT2 #(
		.INIT('h4)
	) name19 (
		\G1_pad ,
		\G2_pad ,
		_w52_
	);
	LUT2 #(
		.INIT('h8)
	) name20 (
		\G3_pad ,
		\G5_pad ,
		_w53_
	);
	LUT2 #(
		.INIT('h4)
	) name21 (
		\G2_pad ,
		\G3_pad ,
		_w54_
	);
	LUT4 #(
		.INIT('h8909)
	) name22 (
		\G2_pad ,
		\G3_pad ,
		\G4_pad ,
		\G5_pad ,
		_w55_
	);
	LUT2 #(
		.INIT('h2)
	) name23 (
		\G4_pad ,
		\G5_pad ,
		_w56_
	);
	LUT3 #(
		.INIT('h04)
	) name24 (
		\G3_pad ,
		\G4_pad ,
		\G5_pad ,
		_w57_
	);
	LUT4 #(
		.INIT('haa08)
	) name25 (
		\G1_pad ,
		\G6_pad ,
		_w55_,
		_w57_,
		_w58_
	);
	LUT3 #(
		.INIT('h31)
	) name26 (
		\G1_pad ,
		\G2_pad ,
		\G4_pad ,
		_w59_
	);
	LUT4 #(
		.INIT('h00f8)
	) name27 (
		\G1_pad ,
		\G4_pad ,
		\G5_pad ,
		\G6_pad ,
		_w60_
	);
	LUT2 #(
		.INIT('h4)
	) name28 (
		_w59_,
		_w60_,
		_w61_
	);
	LUT3 #(
		.INIT('h23)
	) name29 (
		\G4_pad ,
		\G5_pad ,
		\G6_pad ,
		_w62_
	);
	LUT2 #(
		.INIT('h8)
	) name30 (
		\G1_pad ,
		\G3_pad ,
		_w63_
	);
	LUT3 #(
		.INIT('h4c)
	) name31 (
		\G4_pad ,
		\G5_pad ,
		\G6_pad ,
		_w64_
	);
	LUT4 #(
		.INIT('h0ddd)
	) name32 (
		_w52_,
		_w62_,
		_w63_,
		_w64_,
		_w65_
	);
	LUT4 #(
		.INIT('h5455)
	) name33 (
		_w38_,
		_w58_,
		_w61_,
		_w65_,
		_w66_
	);
	LUT2 #(
		.INIT('h2)
	) name34 (
		\G11_pad ,
		\G9_pad ,
		_w67_
	);
	LUT3 #(
		.INIT('h40)
	) name35 (
		\G10_pad ,
		\G7_pad ,
		\G8_pad ,
		_w68_
	);
	LUT2 #(
		.INIT('h1)
	) name36 (
		\G7_pad ,
		\G8_pad ,
		_w69_
	);
	LUT3 #(
		.INIT('h80)
	) name37 (
		\G10_pad ,
		\G11_pad ,
		\G9_pad ,
		_w70_
	);
	LUT4 #(
		.INIT('h0777)
	) name38 (
		_w67_,
		_w68_,
		_w69_,
		_w70_,
		_w71_
	);
	LUT4 #(
		.INIT('h4800)
	) name39 (
		\G1_pad ,
		\G3_pad ,
		\G4_pad ,
		\G6_pad ,
		_w72_
	);
	LUT2 #(
		.INIT('h4)
	) name40 (
		\G1_pad ,
		\G3_pad ,
		_w73_
	);
	LUT4 #(
		.INIT('h0040)
	) name41 (
		\G10_pad ,
		\G4_pad ,
		\G6_pad ,
		\G7_pad ,
		_w74_
	);
	LUT3 #(
		.INIT('h04)
	) name42 (
		\G10_pad ,
		\G7_pad ,
		\G8_pad ,
		_w75_
	);
	LUT4 #(
		.INIT('h0002)
	) name43 (
		\G11_pad ,
		\G4_pad ,
		\G6_pad ,
		\G9_pad ,
		_w76_
	);
	LUT4 #(
		.INIT('h0777)
	) name44 (
		_w34_,
		_w74_,
		_w75_,
		_w76_,
		_w77_
	);
	LUT4 #(
		.INIT('hbb0b)
	) name45 (
		_w71_,
		_w72_,
		_w73_,
		_w77_,
		_w78_
	);
	LUT2 #(
		.INIT('h2)
	) name46 (
		\G2_pad ,
		\G5_pad ,
		_w79_
	);
	LUT2 #(
		.INIT('h1)
	) name47 (
		\G10_pad ,
		\G11_pad ,
		_w80_
	);
	LUT4 #(
		.INIT('h0001)
	) name48 (
		\G10_pad ,
		\G11_pad ,
		\G7_pad ,
		\G8_pad ,
		_w81_
	);
	LUT4 #(
		.INIT('h153f)
	) name49 (
		\G9_pad ,
		_w34_,
		_w35_,
		_w81_,
		_w82_
	);
	LUT4 #(
		.INIT('h8000)
	) name50 (
		\G3_pad ,
		\G4_pad ,
		\G5_pad ,
		\G6_pad ,
		_w83_
	);
	LUT2 #(
		.INIT('h8)
	) name51 (
		\G1_pad ,
		\G2_pad ,
		_w84_
	);
	LUT3 #(
		.INIT('h40)
	) name52 (
		_w82_,
		_w83_,
		_w84_,
		_w85_
	);
	LUT3 #(
		.INIT('h0b)
	) name53 (
		_w78_,
		_w79_,
		_w85_,
		_w86_
	);
	LUT4 #(
		.INIT('h5510)
	) name54 (
		_w66_,
		_w78_,
		_w79_,
		_w85_,
		_w87_
	);
	LUT4 #(
		.INIT('h1333)
	) name55 (
		\G13_pad ,
		_w51_,
		_w52_,
		_w87_,
		_w88_
	);
	LUT3 #(
		.INIT('h20)
	) name56 (
		\G4_pad ,
		\G5_pad ,
		\G6_pad ,
		_w89_
	);
	LUT3 #(
		.INIT('h80)
	) name57 (
		_w69_,
		_w70_,
		_w89_,
		_w90_
	);
	LUT2 #(
		.INIT('h1)
	) name58 (
		\G4_pad ,
		\G5_pad ,
		_w91_
	);
	LUT3 #(
		.INIT('h02)
	) name59 (
		\G11_pad ,
		\G4_pad ,
		\G5_pad ,
		_w92_
	);
	LUT2 #(
		.INIT('h8)
	) name60 (
		\G35_reg/NET0131 ,
		\G3_pad ,
		_w93_
	);
	LUT2 #(
		.INIT('h8)
	) name61 (
		_w92_,
		_w93_,
		_w94_
	);
	LUT4 #(
		.INIT('haa20)
	) name62 (
		\G2_pad ,
		_w82_,
		_w83_,
		_w94_,
		_w95_
	);
	LUT3 #(
		.INIT('ha8)
	) name63 (
		_w39_,
		_w50_,
		_w95_,
		_w96_
	);
	LUT2 #(
		.INIT('h8)
	) name64 (
		\G13_pad ,
		\G1_pad ,
		_w97_
	);
	LUT2 #(
		.INIT('h8)
	) name65 (
		\G4_pad ,
		\G5_pad ,
		_w98_
	);
	LUT3 #(
		.INIT('h80)
	) name66 (
		\G9_pad ,
		_w81_,
		_w98_,
		_w99_
	);
	LUT2 #(
		.INIT('h8)
	) name67 (
		_w42_,
		_w92_,
		_w100_
	);
	LUT3 #(
		.INIT('h80)
	) name68 (
		\G2_pad ,
		\G3_pad ,
		\G6_pad ,
		_w101_
	);
	LUT3 #(
		.INIT('he0)
	) name69 (
		_w99_,
		_w100_,
		_w101_,
		_w102_
	);
	LUT4 #(
		.INIT('hec00)
	) name70 (
		_w87_,
		_w96_,
		_w97_,
		_w102_,
		_w103_
	);
	LUT2 #(
		.INIT('h2)
	) name71 (
		\G13_pad ,
		\G43_reg/NET0131 ,
		_w104_
	);
	LUT2 #(
		.INIT('h8)
	) name72 (
		_w66_,
		_w104_,
		_w105_
	);
	LUT3 #(
		.INIT('h02)
	) name73 (
		\G36_reg/NET0131 ,
		\G4_pad ,
		\G6_pad ,
		_w106_
	);
	LUT4 #(
		.INIT('h007f)
	) name74 (
		_w47_,
		_w67_,
		_w68_,
		_w106_,
		_w107_
	);
	LUT2 #(
		.INIT('h1)
	) name75 (
		\G3_pad ,
		_w107_,
		_w108_
	);
	LUT3 #(
		.INIT('h80)
	) name76 (
		_w39_,
		_w50_,
		_w108_,
		_w109_
	);
	LUT2 #(
		.INIT('h1)
	) name77 (
		_w105_,
		_w109_,
		_w110_
	);
	LUT4 #(
		.INIT('h0b00)
	) name78 (
		_w88_,
		_w90_,
		_w103_,
		_w110_,
		_w111_
	);
	LUT2 #(
		.INIT('h2)
	) name79 (
		\G12_pad ,
		\G13_pad ,
		_w112_
	);
	LUT3 #(
		.INIT('h20)
	) name80 (
		\G30_reg/NET0131 ,
		\G6_pad ,
		\G7_pad ,
		_w113_
	);
	LUT4 #(
		.INIT('h5155)
	) name81 (
		\G10_pad ,
		\G30_reg/NET0131 ,
		\G6_pad ,
		\G7_pad ,
		_w114_
	);
	LUT2 #(
		.INIT('h8)
	) name82 (
		\G31_reg/NET0131 ,
		\G8_pad ,
		_w115_
	);
	LUT3 #(
		.INIT('h32)
	) name83 (
		\G10_pad ,
		\G7_pad ,
		\G8_pad ,
		_w116_
	);
	LUT4 #(
		.INIT('h3120)
	) name84 (
		\G9_pad ,
		_w115_,
		_w116_,
		_w114_,
		_w117_
	);
	LUT4 #(
		.INIT('h3133)
	) name85 (
		\G30_reg/NET0131 ,
		\G31_reg/NET0131 ,
		\G6_pad ,
		\G7_pad ,
		_w118_
	);
	LUT4 #(
		.INIT('ha0f3)
	) name86 (
		\G10_pad ,
		\G7_pad ,
		\G8_pad ,
		\G9_pad ,
		_w119_
	);
	LUT3 #(
		.INIT('ha8)
	) name87 (
		\G11_pad ,
		\G30_reg/NET0131 ,
		\G6_pad ,
		_w120_
	);
	LUT4 #(
		.INIT('h2f00)
	) name88 (
		\G8_pad ,
		_w118_,
		_w119_,
		_w120_,
		_w121_
	);
	LUT2 #(
		.INIT('h8)
	) name89 (
		\G0_pad ,
		\G3_pad ,
		_w122_
	);
	LUT3 #(
		.INIT('h23)
	) name90 (
		\G3_pad ,
		\G4_pad ,
		\G5_pad ,
		_w123_
	);
	LUT4 #(
		.INIT('h0407)
	) name91 (
		\G0_pad ,
		\G3_pad ,
		\G4_pad ,
		\G5_pad ,
		_w124_
	);
	LUT2 #(
		.INIT('h2)
	) name92 (
		\G46_reg/NET0131 ,
		_w124_,
		_w125_
	);
	LUT4 #(
		.INIT('hf100)
	) name93 (
		\G11_pad ,
		_w117_,
		_w121_,
		_w125_,
		_w126_
	);
	LUT4 #(
		.INIT('ha2f3)
	) name94 (
		\G2_pad ,
		\G3_pad ,
		\G4_pad ,
		\G5_pad ,
		_w127_
	);
	LUT3 #(
		.INIT('h4c)
	) name95 (
		\G1_pad ,
		\G2_pad ,
		\G3_pad ,
		_w128_
	);
	LUT4 #(
		.INIT('h83b0)
	) name96 (
		\G1_pad ,
		\G2_pad ,
		\G3_pad ,
		\G5_pad ,
		_w129_
	);
	LUT4 #(
		.INIT('hf531)
	) name97 (
		\G1_pad ,
		\G4_pad ,
		_w127_,
		_w129_,
		_w130_
	);
	LUT2 #(
		.INIT('h2)
	) name98 (
		\G0_pad ,
		_w130_,
		_w131_
	);
	LUT3 #(
		.INIT('h80)
	) name99 (
		_w112_,
		_w126_,
		_w131_,
		_w132_
	);
	LUT3 #(
		.INIT('hf1)
	) name100 (
		\G12_pad ,
		_w111_,
		_w132_,
		_w133_
	);
	LUT3 #(
		.INIT('h01)
	) name101 (
		\G4_pad ,
		\G5_pad ,
		\G6_pad ,
		_w134_
	);
	LUT4 #(
		.INIT('h0777)
	) name102 (
		_w47_,
		_w70_,
		_w80_,
		_w134_,
		_w135_
	);
	LUT3 #(
		.INIT('h20)
	) name103 (
		\G10_pad ,
		\G6_pad ,
		\G7_pad ,
		_w136_
	);
	LUT3 #(
		.INIT('h80)
	) name104 (
		_w34_,
		_w56_,
		_w136_,
		_w137_
	);
	LUT4 #(
		.INIT('h5504)
	) name105 (
		\G3_pad ,
		_w69_,
		_w135_,
		_w137_,
		_w138_
	);
	LUT2 #(
		.INIT('h8)
	) name106 (
		_w40_,
		_w42_,
		_w139_
	);
	LUT3 #(
		.INIT('h80)
	) name107 (
		\G11_pad ,
		_w40_,
		_w42_,
		_w140_
	);
	LUT2 #(
		.INIT('h1)
	) name108 (
		_w138_,
		_w140_,
		_w141_
	);
	LUT3 #(
		.INIT('h40)
	) name109 (
		\G12_pad ,
		_w39_,
		_w50_,
		_w142_
	);
	LUT2 #(
		.INIT('h4)
	) name110 (
		_w141_,
		_w142_,
		_w143_
	);
	LUT2 #(
		.INIT('h8)
	) name111 (
		\G11_pad ,
		\G2_pad ,
		_w144_
	);
	LUT2 #(
		.INIT('h8)
	) name112 (
		\G6_pad ,
		\G9_pad ,
		_w145_
	);
	LUT3 #(
		.INIT('h80)
	) name113 (
		\G10_pad ,
		\G4_pad ,
		\G7_pad ,
		_w146_
	);
	LUT3 #(
		.INIT('h80)
	) name114 (
		_w53_,
		_w145_,
		_w146_,
		_w147_
	);
	LUT3 #(
		.INIT('h04)
	) name115 (
		\G10_pad ,
		\G7_pad ,
		\G9_pad ,
		_w148_
	);
	LUT4 #(
		.INIT('h0200)
	) name116 (
		\G3_pad ,
		\G4_pad ,
		\G5_pad ,
		\G6_pad ,
		_w149_
	);
	LUT2 #(
		.INIT('h8)
	) name117 (
		_w148_,
		_w149_,
		_w150_
	);
	LUT3 #(
		.INIT('ha8)
	) name118 (
		\G8_pad ,
		_w147_,
		_w150_,
		_w151_
	);
	LUT4 #(
		.INIT('hec00)
	) name119 (
		_w87_,
		_w96_,
		_w97_,
		_w151_,
		_w152_
	);
	LUT4 #(
		.INIT('h2000)
	) name120 (
		\G13_pad ,
		\G1_pad ,
		_w87_,
		_w139_,
		_w153_
	);
	LUT2 #(
		.INIT('h1)
	) name121 (
		\G0_pad ,
		\G4_pad ,
		_w154_
	);
	LUT4 #(
		.INIT('h0002)
	) name122 (
		\G10_pad ,
		\G3_pad ,
		\G5_pad ,
		\G8_pad ,
		_w155_
	);
	LUT4 #(
		.INIT('h0008)
	) name123 (
		\G11_pad ,
		\G6_pad ,
		\G7_pad ,
		\G9_pad ,
		_w156_
	);
	LUT4 #(
		.INIT('h8000)
	) name124 (
		\G11_pad ,
		\G37_reg/NET0131 ,
		\G3_pad ,
		\G5_pad ,
		_w157_
	);
	LUT4 #(
		.INIT('h153f)
	) name125 (
		_w68_,
		_w155_,
		_w156_,
		_w157_,
		_w158_
	);
	LUT4 #(
		.INIT('h8000)
	) name126 (
		_w34_,
		_w35_,
		_w47_,
		_w122_,
		_w159_
	);
	LUT4 #(
		.INIT('haa08)
	) name127 (
		_w84_,
		_w154_,
		_w158_,
		_w159_,
		_w160_
	);
	LUT3 #(
		.INIT('h20)
	) name128 (
		_w112_,
		_w126_,
		_w160_,
		_w161_
	);
	LUT3 #(
		.INIT('h08)
	) name129 (
		\G38_reg/NET0131 ,
		\G6_pad ,
		\G9_pad ,
		_w162_
	);
	LUT4 #(
		.INIT('h007f)
	) name130 (
		\G0_pad ,
		_w145_,
		_w146_,
		_w162_,
		_w163_
	);
	LUT4 #(
		.INIT('h8000)
	) name131 (
		\G1_pad ,
		\G3_pad ,
		\G5_pad ,
		\G8_pad ,
		_w164_
	);
	LUT2 #(
		.INIT('h4)
	) name132 (
		_w163_,
		_w164_,
		_w165_
	);
	LUT4 #(
		.INIT('h2000)
	) name133 (
		_w112_,
		_w126_,
		_w160_,
		_w165_,
		_w166_
	);
	LUT4 #(
		.INIT('h00ab)
	) name134 (
		\G12_pad ,
		_w152_,
		_w153_,
		_w166_,
		_w167_
	);
	LUT3 #(
		.INIT('hae)
	) name135 (
		_w143_,
		_w144_,
		_w167_,
		_w168_
	);
	LUT4 #(
		.INIT('h1101)
	) name136 (
		\G12_pad ,
		\G13_pad ,
		\G32_reg/NET0131 ,
		_w38_,
		_w169_
	);
	LUT3 #(
		.INIT('h10)
	) name137 (
		_w50_,
		_w95_,
		_w169_,
		_w170_
	);
	LUT3 #(
		.INIT('h02)
	) name138 (
		_w112_,
		_w126_,
		_w160_,
		_w171_
	);
	LUT2 #(
		.INIT('h4)
	) name139 (
		\G12_pad ,
		\G13_pad ,
		_w172_
	);
	LUT2 #(
		.INIT('h4)
	) name140 (
		_w66_,
		_w172_,
		_w173_
	);
	LUT4 #(
		.INIT('hffec)
	) name141 (
		_w86_,
		_w171_,
		_w173_,
		_w170_,
		_w174_
	);
	LUT2 #(
		.INIT('h8)
	) name142 (
		\G34_reg/NET0131 ,
		\G8_pad ,
		_w175_
	);
	LUT4 #(
		.INIT('h007f)
	) name143 (
		\G6_pad ,
		_w112_,
		_w126_,
		_w175_,
		_w176_
	);
	LUT3 #(
		.INIT('h80)
	) name144 (
		\G10_pad ,
		\G34_reg/NET0131 ,
		\G7_pad ,
		_w177_
	);
	LUT2 #(
		.INIT('h4)
	) name145 (
		_w41_,
		_w177_,
		_w178_
	);
	LUT4 #(
		.INIT('h0800)
	) name146 (
		\G10_pad ,
		\G11_pad ,
		\G8_pad ,
		\G9_pad ,
		_w179_
	);
	LUT3 #(
		.INIT('ha2)
	) name147 (
		\G11_pad ,
		\G7_pad ,
		\G8_pad ,
		_w180_
	);
	LUT3 #(
		.INIT('h0e)
	) name148 (
		\G10_pad ,
		\G11_pad ,
		\G9_pad ,
		_w181_
	);
	LUT4 #(
		.INIT('h20a0)
	) name149 (
		\G10_pad ,
		\G7_pad ,
		\G8_pad ,
		\G9_pad ,
		_w182_
	);
	LUT4 #(
		.INIT('h000b)
	) name150 (
		_w180_,
		_w181_,
		_w182_,
		_w179_,
		_w183_
	);
	LUT4 #(
		.INIT('h0080)
	) name151 (
		\G6_pad ,
		_w112_,
		_w126_,
		_w183_,
		_w184_
	);
	LUT4 #(
		.INIT('hffce)
	) name152 (
		_w37_,
		_w178_,
		_w176_,
		_w184_,
		_w185_
	);
	LUT4 #(
		.INIT('h48c0)
	) name153 (
		\G10_pad ,
		\G34_reg/NET0131 ,
		\G7_pad ,
		\G8_pad ,
		_w186_
	);
	LUT4 #(
		.INIT('h007f)
	) name154 (
		_w112_,
		_w126_,
		_w136_,
		_w186_,
		_w187_
	);
	LUT4 #(
		.INIT('h3010)
	) name155 (
		\G10_pad ,
		\G7_pad ,
		\G8_pad ,
		\G9_pad ,
		_w188_
	);
	LUT4 #(
		.INIT('h0d00)
	) name156 (
		\G10_pad ,
		\G11_pad ,
		\G8_pad ,
		\G9_pad ,
		_w189_
	);
	LUT4 #(
		.INIT('h0405)
	) name157 (
		_w37_,
		_w80_,
		_w189_,
		_w188_,
		_w190_
	);
	LUT4 #(
		.INIT('h0080)
	) name158 (
		\G6_pad ,
		_w112_,
		_w126_,
		_w190_,
		_w191_
	);
	LUT3 #(
		.INIT('hf2)
	) name159 (
		\G9_pad ,
		_w187_,
		_w191_,
		_w192_
	);
	LUT4 #(
		.INIT('h8044)
	) name160 (
		\G10_pad ,
		\G7_pad ,
		\G8_pad ,
		\G9_pad ,
		_w193_
	);
	LUT4 #(
		.INIT('h8880)
	) name161 (
		\G11_pad ,
		\G34_reg/NET0131 ,
		\G7_pad ,
		\G8_pad ,
		_w194_
	);
	LUT3 #(
		.INIT('h10)
	) name162 (
		_w43_,
		_w193_,
		_w194_,
		_w195_
	);
	LUT4 #(
		.INIT('hff40)
	) name163 (
		\G42_reg/NET0131 ,
		_w112_,
		_w126_,
		_w195_,
		_w196_
	);
	LUT4 #(
		.INIT('h1d0f)
	) name164 (
		\G2_pad ,
		\G3_pad ,
		\G5_pad ,
		\G6_pad ,
		_w197_
	);
	LUT2 #(
		.INIT('h1)
	) name165 (
		\G4_pad ,
		_w197_,
		_w198_
	);
	LUT3 #(
		.INIT('h40)
	) name166 (
		\G3_pad ,
		\G4_pad ,
		\G6_pad ,
		_w199_
	);
	LUT4 #(
		.INIT('h8bbb)
	) name167 (
		\G2_pad ,
		\G3_pad ,
		\G4_pad ,
		\G6_pad ,
		_w200_
	);
	LUT3 #(
		.INIT('h08)
	) name168 (
		\G2_pad ,
		\G4_pad ,
		\G5_pad ,
		_w201_
	);
	LUT3 #(
		.INIT('h0d)
	) name169 (
		\G5_pad ,
		_w200_,
		_w201_,
		_w202_
	);
	LUT2 #(
		.INIT('h4)
	) name170 (
		_w198_,
		_w202_,
		_w203_
	);
	LUT4 #(
		.INIT('h0080)
	) name171 (
		\G1_pad ,
		_w66_,
		_w172_,
		_w203_,
		_w204_
	);
	LUT4 #(
		.INIT('h4c00)
	) name172 (
		\G0_pad ,
		\G1_pad ,
		\G3_pad ,
		\G4_pad ,
		_w205_
	);
	LUT3 #(
		.INIT('h80)
	) name173 (
		_w112_,
		_w126_,
		_w205_,
		_w206_
	);
	LUT3 #(
		.INIT('h10)
	) name174 (
		\G13_pad ,
		\G33_reg/NET0131 ,
		\G3_pad ,
		_w207_
	);
	LUT4 #(
		.INIT('h0010)
	) name175 (
		\G12_pad ,
		\G13_pad ,
		\G32_reg/NET0131 ,
		_w38_,
		_w208_
	);
	LUT4 #(
		.INIT('h2a00)
	) name176 (
		\G2_pad ,
		\G3_pad ,
		\G4_pad ,
		\G5_pad ,
		_w209_
	);
	LUT3 #(
		.INIT('h15)
	) name177 (
		_w207_,
		_w208_,
		_w209_,
		_w210_
	);
	LUT3 #(
		.INIT('hef)
	) name178 (
		_w204_,
		_w206_,
		_w210_,
		_w211_
	);
	LUT4 #(
		.INIT('h4c80)
	) name179 (
		\G1_pad ,
		\G2_pad ,
		\G4_pad ,
		\G5_pad ,
		_w212_
	);
	LUT3 #(
		.INIT('h80)
	) name180 (
		_w66_,
		_w172_,
		_w212_,
		_w213_
	);
	LUT2 #(
		.INIT('h2)
	) name181 (
		\G0_pad ,
		\G29_reg/NET0131 ,
		_w214_
	);
	LUT4 #(
		.INIT('h4000)
	) name182 (
		\G0_pad ,
		\G1_pad ,
		\G3_pad ,
		\G4_pad ,
		_w215_
	);
	LUT2 #(
		.INIT('h1)
	) name183 (
		_w214_,
		_w215_,
		_w216_
	);
	LUT3 #(
		.INIT('h08)
	) name184 (
		_w112_,
		_w126_,
		_w216_,
		_w217_
	);
	LUT4 #(
		.INIT('h4c00)
	) name185 (
		\G2_pad ,
		\G3_pad ,
		\G4_pad ,
		\G5_pad ,
		_w218_
	);
	LUT3 #(
		.INIT('h15)
	) name186 (
		_w207_,
		_w208_,
		_w218_,
		_w219_
	);
	LUT3 #(
		.INIT('hef)
	) name187 (
		_w217_,
		_w213_,
		_w219_,
		_w220_
	);
	LUT3 #(
		.INIT('h08)
	) name188 (
		\G0_pad ,
		\G2_pad ,
		\G4_pad ,
		_w221_
	);
	LUT4 #(
		.INIT('h00ec)
	) name189 (
		\G0_pad ,
		\G1_pad ,
		\G2_pad ,
		\G3_pad ,
		_w222_
	);
	LUT4 #(
		.INIT('h9b5f)
	) name190 (
		\G0_pad ,
		\G1_pad ,
		\G3_pad ,
		\G4_pad ,
		_w223_
	);
	LUT3 #(
		.INIT('hb0)
	) name191 (
		_w221_,
		_w222_,
		_w223_,
		_w224_
	);
	LUT3 #(
		.INIT('h08)
	) name192 (
		_w112_,
		_w126_,
		_w224_,
		_w225_
	);
	LUT4 #(
		.INIT('h6400)
	) name193 (
		\G1_pad ,
		\G2_pad ,
		\G3_pad ,
		\G4_pad ,
		_w226_
	);
	LUT3 #(
		.INIT('h80)
	) name194 (
		_w66_,
		_w172_,
		_w226_,
		_w227_
	);
	LUT3 #(
		.INIT('ha8)
	) name195 (
		\G5_pad ,
		_w225_,
		_w227_,
		_w228_
	);
	LUT4 #(
		.INIT('h0400)
	) name196 (
		\G2_pad ,
		\G3_pad ,
		\G5_pad ,
		\G6_pad ,
		_w229_
	);
	LUT4 #(
		.INIT('h00b0)
	) name197 (
		\G2_pad ,
		\G3_pad ,
		\G4_pad ,
		\G5_pad ,
		_w230_
	);
	LUT3 #(
		.INIT('h01)
	) name198 (
		_w199_,
		_w230_,
		_w229_,
		_w231_
	);
	LUT4 #(
		.INIT('h0080)
	) name199 (
		\G1_pad ,
		_w66_,
		_w172_,
		_w231_,
		_w232_
	);
	LUT2 #(
		.INIT('h8)
	) name200 (
		\G39_reg/NET0131 ,
		\G4_pad ,
		_w233_
	);
	LUT2 #(
		.INIT('h8)
	) name201 (
		_w208_,
		_w233_,
		_w234_
	);
	LUT2 #(
		.INIT('h1)
	) name202 (
		_w232_,
		_w234_,
		_w235_
	);
	LUT2 #(
		.INIT('hb)
	) name203 (
		_w228_,
		_w235_,
		_w236_
	);
	LUT3 #(
		.INIT('h8c)
	) name204 (
		\G1_pad ,
		\G4_pad ,
		\G5_pad ,
		_w237_
	);
	LUT4 #(
		.INIT('h0800)
	) name205 (
		\G1_pad ,
		\G3_pad ,
		\G4_pad ,
		\G5_pad ,
		_w238_
	);
	LUT3 #(
		.INIT('h0d)
	) name206 (
		_w128_,
		_w237_,
		_w238_,
		_w239_
	);
	LUT3 #(
		.INIT('h08)
	) name207 (
		_w66_,
		_w172_,
		_w239_,
		_w240_
	);
	LUT4 #(
		.INIT('h4404)
	) name208 (
		\G2_pad ,
		\G3_pad ,
		\G4_pad ,
		\G5_pad ,
		_w241_
	);
	LUT3 #(
		.INIT('ha8)
	) name209 (
		\G2_pad ,
		\G4_pad ,
		\G5_pad ,
		_w242_
	);
	LUT4 #(
		.INIT('h915b)
	) name210 (
		\G2_pad ,
		\G3_pad ,
		\G4_pad ,
		\G5_pad ,
		_w243_
	);
	LUT2 #(
		.INIT('h2)
	) name211 (
		_w208_,
		_w243_,
		_w244_
	);
	LUT3 #(
		.INIT('ha8)
	) name212 (
		\G6_pad ,
		_w240_,
		_w244_,
		_w245_
	);
	LUT3 #(
		.INIT('h40)
	) name213 (
		\G40_reg/NET0131 ,
		_w112_,
		_w126_,
		_w246_
	);
	LUT4 #(
		.INIT('h4c00)
	) name214 (
		\G2_pad ,
		\G4_pad ,
		\G5_pad ,
		\G6_pad ,
		_w247_
	);
	LUT4 #(
		.INIT('h8000)
	) name215 (
		\G1_pad ,
		_w66_,
		_w172_,
		_w247_,
		_w248_
	);
	LUT2 #(
		.INIT('h1)
	) name216 (
		_w246_,
		_w248_,
		_w249_
	);
	LUT2 #(
		.INIT('hb)
	) name217 (
		_w245_,
		_w249_,
		_w250_
	);
	LUT4 #(
		.INIT('h4000)
	) name218 (
		\G12_pad ,
		_w39_,
		_w49_,
		_w50_,
		_w251_
	);
	LUT4 #(
		.INIT('h44c4)
	) name219 (
		\G0_pad ,
		\G1_pad ,
		\G3_pad ,
		\G4_pad ,
		_w252_
	);
	LUT4 #(
		.INIT('h8a0f)
	) name220 (
		\G1_pad ,
		\G3_pad ,
		\G4_pad ,
		\G5_pad ,
		_w253_
	);
	LUT4 #(
		.INIT('h4f45)
	) name221 (
		\G0_pad ,
		_w123_,
		_w252_,
		_w253_,
		_w254_
	);
	LUT2 #(
		.INIT('h2)
	) name222 (
		\G2_pad ,
		_w254_,
		_w255_
	);
	LUT3 #(
		.INIT('h80)
	) name223 (
		_w112_,
		_w126_,
		_w255_,
		_w256_
	);
	LUT2 #(
		.INIT('he)
	) name224 (
		_w251_,
		_w256_,
		_w257_
	);
	LUT4 #(
		.INIT('h1143)
	) name225 (
		\G2_pad ,
		\G3_pad ,
		\G4_pad ,
		\G5_pad ,
		_w258_
	);
	LUT3 #(
		.INIT('h31)
	) name226 (
		\G0_pad ,
		\G1_pad ,
		_w258_,
		_w259_
	);
	LUT4 #(
		.INIT('h010f)
	) name227 (
		\G10_pad ,
		\G30_reg/NET0131 ,
		\G6_pad ,
		\G7_pad ,
		_w260_
	);
	LUT4 #(
		.INIT('h4044)
	) name228 (
		\G1_pad ,
		\G3_pad ,
		\G4_pad ,
		\G5_pad ,
		_w261_
	);
	LUT4 #(
		.INIT('ha202)
	) name229 (
		\G0_pad ,
		\G3_pad ,
		\G4_pad ,
		\G5_pad ,
		_w262_
	);
	LUT4 #(
		.INIT('h8880)
	) name230 (
		\G2_pad ,
		_w253_,
		_w261_,
		_w262_,
		_w263_
	);
	LUT3 #(
		.INIT('h01)
	) name231 (
		_w259_,
		_w260_,
		_w263_,
		_w264_
	);
	LUT3 #(
		.INIT('hf8)
	) name232 (
		_w66_,
		_w172_,
		_w208_,
		_w265_
	);
	LUT4 #(
		.INIT('h7400)
	) name233 (
		\G10_pad ,
		\G11_pad ,
		\G7_pad ,
		\G9_pad ,
		_w266_
	);
	LUT4 #(
		.INIT('h0307)
	) name234 (
		\G31_reg/NET0131 ,
		\G6_pad ,
		_w113_,
		_w266_,
		_w267_
	);
	LUT2 #(
		.INIT('hd)
	) name235 (
		\G8_pad ,
		_w267_,
		_w268_
	);
	LUT4 #(
		.INIT('h770f)
	) name236 (
		\G10_pad ,
		\G6_pad ,
		\G7_pad ,
		\G8_pad ,
		_w269_
	);
	LUT4 #(
		.INIT('h93cf)
	) name237 (
		\G10_pad ,
		\G6_pad ,
		\G7_pad ,
		\G9_pad ,
		_w270_
	);
	LUT4 #(
		.INIT('hfd55)
	) name238 (
		\G11_pad ,
		\G9_pad ,
		_w269_,
		_w270_,
		_w271_
	);
	LUT4 #(
		.INIT('h8207)
	) name239 (
		\G2_pad ,
		\G4_pad ,
		\G5_pad ,
		\G6_pad ,
		_w272_
	);
	LUT4 #(
		.INIT('hfb51)
	) name240 (
		\G1_pad ,
		\G2_pad ,
		_w62_,
		_w272_,
		_w273_
	);
	LUT2 #(
		.INIT('hd)
	) name241 (
		\G3_pad ,
		_w273_,
		_w274_
	);
	LUT3 #(
		.INIT('h80)
	) name242 (
		_w47_,
		_w69_,
		_w70_,
		_w275_
	);
	LUT3 #(
		.INIT('h80)
	) name243 (
		_w34_,
		_w35_,
		_w134_,
		_w276_
	);
	LUT3 #(
		.INIT('h01)
	) name244 (
		\G5_pad ,
		\G6_pad ,
		\G9_pad ,
		_w277_
	);
	LUT2 #(
		.INIT('h8)
	) name245 (
		_w81_,
		_w277_,
		_w278_
	);
	LUT3 #(
		.INIT('h01)
	) name246 (
		_w276_,
		_w275_,
		_w278_,
		_w279_
	);
	LUT4 #(
		.INIT('h5540)
	) name247 (
		\G5_pad ,
		_w34_,
		_w35_,
		_w81_,
		_w280_
	);
	LUT4 #(
		.INIT('h2f22)
	) name248 (
		_w54_,
		_w62_,
		_w83_,
		_w242_,
		_w281_
	);
	LUT3 #(
		.INIT('h47)
	) name249 (
		\G3_pad ,
		\G4_pad ,
		\G5_pad ,
		_w282_
	);
	LUT3 #(
		.INIT('h31)
	) name250 (
		_w52_,
		_w241_,
		_w282_,
		_w283_
	);
	LUT4 #(
		.INIT('h0100)
	) name251 (
		\G0_pad ,
		\G10_pad ,
		\G4_pad ,
		\G7_pad ,
		_w284_
	);
	LUT3 #(
		.INIT('h6a)
	) name252 (
		\G2_pad ,
		\G3_pad ,
		\G5_pad ,
		_w285_
	);
	LUT4 #(
		.INIT('h2eae)
	) name253 (
		\G10_pad ,
		\G11_pad ,
		\G7_pad ,
		\G9_pad ,
		_w286_
	);
	LUT3 #(
		.INIT('hae)
	) name254 (
		\G10_pad ,
		\G11_pad ,
		\G9_pad ,
		_w287_
	);
	LUT2 #(
		.INIT('h6)
	) name255 (
		\G6_pad ,
		\G9_pad ,
		_w288_
	);
	LUT4 #(
		.INIT('h5540)
	) name256 (
		\G12_pad ,
		\G13_pad ,
		_w87_,
		_w96_,
		_w289_
	);
	LUT2 #(
		.INIT('he)
	) name257 (
		_w161_,
		_w289_,
		_w290_
	);
	LUT4 #(
		.INIT('h1040)
	) name258 (
		\G10_pad ,
		\G7_pad ,
		\G8_pad ,
		\G9_pad ,
		_w291_
	);
	LUT2 #(
		.INIT('h1)
	) name259 (
		\G3_pad ,
		\G44_reg/NET0131 ,
		_w292_
	);
	LUT4 #(
		.INIT('h007f)
	) name260 (
		\G11_pad ,
		_w40_,
		_w291_,
		_w292_,
		_w293_
	);
	LUT4 #(
		.INIT('h0040)
	) name261 (
		\G12_pad ,
		_w39_,
		_w50_,
		_w293_,
		_w294_
	);
	LUT2 #(
		.INIT('h8)
	) name262 (
		_w42_,
		_w91_,
		_w295_
	);
	LUT4 #(
		.INIT('hec00)
	) name263 (
		_w87_,
		_w96_,
		_w97_,
		_w295_,
		_w296_
	);
	LUT4 #(
		.INIT('h2000)
	) name264 (
		\G13_pad ,
		\G1_pad ,
		_w87_,
		_w291_,
		_w297_
	);
	LUT3 #(
		.INIT('h40)
	) name265 (
		\G12_pad ,
		\G3_pad ,
		\G6_pad ,
		_w298_
	);
	LUT2 #(
		.INIT('h8)
	) name266 (
		\G37_reg/NET0131 ,
		\G38_reg/NET0131 ,
		_w299_
	);
	LUT2 #(
		.INIT('h8)
	) name267 (
		_w164_,
		_w299_,
		_w300_
	);
	LUT4 #(
		.INIT('h2000)
	) name268 (
		_w112_,
		_w126_,
		_w160_,
		_w300_,
		_w301_
	);
	LUT4 #(
		.INIT('h001f)
	) name269 (
		_w296_,
		_w297_,
		_w298_,
		_w301_,
		_w302_
	);
	LUT3 #(
		.INIT('hce)
	) name270 (
		_w144_,
		_w294_,
		_w302_,
		_w303_
	);
	LUT4 #(
		.INIT('h20a0)
	) name271 (
		\G10_pad ,
		\G6_pad ,
		\G7_pad ,
		\G9_pad ,
		_w304_
	);
	LUT2 #(
		.INIT('h8)
	) name272 (
		\G34_reg/NET0131 ,
		_w182_,
		_w305_
	);
	LUT4 #(
		.INIT('h007f)
	) name273 (
		_w112_,
		_w126_,
		_w304_,
		_w305_,
		_w306_
	);
	LUT3 #(
		.INIT('hd0)
	) name274 (
		_w37_,
		_w176_,
		_w306_,
		_w307_
	);
	LUT4 #(
		.INIT('h0400)
	) name275 (
		\G12_pad ,
		\G32_reg/NET0131 ,
		_w38_,
		_w201_,
		_w308_
	);
	LUT4 #(
		.INIT('h0080)
	) name276 (
		\G0_pad ,
		\G12_pad ,
		\G1_pad ,
		\G4_pad ,
		_w309_
	);
	LUT3 #(
		.INIT('h13)
	) name277 (
		_w126_,
		_w308_,
		_w309_,
		_w310_
	);
	LUT4 #(
		.INIT('hb1a0)
	) name278 (
		\G6_pad ,
		\G9_pad ,
		_w42_,
		_w75_,
		_w311_
	);
	assign \G532_pad  = _w133_ ;
	assign \G537_pad  = _w168_ ;
	assign \G539_pad  = _w174_ ;
	assign \G542_pad  = _w185_ ;
	assign \G546_pad  = _w23_ ;
	assign \G547_pad  = _w192_ ;
	assign \G548_pad  = _w196_ ;
	assign \G549_pad  = _w211_ ;
	assign \G550_pad  = _w220_ ;
	assign \G551_pad  = _w236_ ;
	assign \G552_pad  = _w250_ ;
	assign \_al_n0  = 1'b0;
	assign \_al_n1  = 1'b1;
	assign \g1667/_3_  = _w257_ ;
	assign \g1737/_0_  = _w264_ ;
	assign \g1744/_0_  = _w265_ ;
	assign \g1787/_0_  = _w268_ ;
	assign \g1811/_0_  = _w271_ ;
	assign \g1830/_0_  = _w274_ ;
	assign \g1831/_0_  = _w279_ ;
	assign \g1846/_0_  = _w280_ ;
	assign \g1852/_0_  = _w281_ ;
	assign \g1866/_0_  = _w283_ ;
	assign \g19/_2_  = _w284_ ;
	assign \g1931/_0_  = _w285_ ;
	assign \g1945/_0_  = _w286_ ;
	assign \g2014/_0_  = _w287_ ;
	assign \g2015/_0_  = _w288_ ;
	assign \g2643/_0_  = _w290_ ;
	assign \g2859/_1_  = _w303_ ;
	assign \g3397/_2_  = _w307_ ;
	assign \g3546/_0_  = _w310_ ;
	assign \g3606/_3_  = _w311_ ;
endmodule;