module top( \a0_pad  , a_pad , \b0_pad  , b_pad , \c0_pad  , c_pad , \d0_pad  , d_pad , \e0_pad  , e_pad , \f0_pad  , f_pad , \g0_pad  , g_pad , \h0_pad  , h_pad , \i0_pad  , i_pad , \j0_pad  , j_pad , \k0_pad  , k_pad , l_pad , m_pad , n_pad , o_pad , p_pad , q_pad , s_pad , t_pad , u_pad , v_pad , w_pad , x_pad , y_pad , z_pad , \a1_pad  , \l0_pad  , \m0_pad  , \n0_pad  , \o0_pad  , \p0_pad  , \q0_pad  , \r0_pad  , \s0_pad  , \t0_pad  , \u0_pad  , \v0_pad  , \w0_pad  , \x0_pad  , \y0_pad  , \z0_pad  );
  input \a0_pad  ;
  input a_pad ;
  input \b0_pad  ;
  input b_pad ;
  input \c0_pad  ;
  input c_pad ;
  input \d0_pad  ;
  input d_pad ;
  input \e0_pad  ;
  input e_pad ;
  input \f0_pad  ;
  input f_pad ;
  input \g0_pad  ;
  input g_pad ;
  input \h0_pad  ;
  input h_pad ;
  input \i0_pad  ;
  input i_pad ;
  input \j0_pad  ;
  input j_pad ;
  input \k0_pad  ;
  input k_pad ;
  input l_pad ;
  input m_pad ;
  input n_pad ;
  input o_pad ;
  input p_pad ;
  input q_pad ;
  input s_pad ;
  input t_pad ;
  input u_pad ;
  input v_pad ;
  input w_pad ;
  input x_pad ;
  input y_pad ;
  input z_pad ;
  output \a1_pad  ;
  output \l0_pad  ;
  output \m0_pad  ;
  output \n0_pad  ;
  output \o0_pad  ;
  output \p0_pad  ;
  output \q0_pad  ;
  output \r0_pad  ;
  output \s0_pad  ;
  output \t0_pad  ;
  output \u0_pad  ;
  output \v0_pad  ;
  output \w0_pad  ;
  output \x0_pad  ;
  output \y0_pad  ;
  output \z0_pad  ;
  wire n37 , n38 , n39 , n40 , n41 , n42 , n43 , n44 , n45 , n46 , n47 , n48 , n49 , n50 , n51 , n52 , n53 , n54 , n55 , n56 , n57 , n58 , n59 , n60 , n61 , n62 , n63 , n64 , n65 , n66 , n67 , n68 , n69 , n70 , n71 , n72 , n73 , n74 , n75 , n76 , n77 , n78 , n79 , n80 , n81 , n82 , n83 , n84 , n85 , n86 , n87 , n88 , n89 , n90 , n91 , n92 , n93 , n94 , n95 , n96 , n97 , n98 , n99 , n100 , n101 , n102 , n103 , n104 , n105 , n106 , n107 , n108 , n109 , n110 , n111 , n112 , n113 , n114 , n115 , n116 , n117 , n118 , n119 , n120 , n121 , n122 , n123 , n124 , n125 , n126 , n127 , n128 , n129 , n130 , n131 , n132 , n133 ;
  assign n37 = ~\k0_pad  & ~u_pad ;
  assign n40 = \d0_pad  & t_pad ;
  assign n38 = ~s_pad & u_pad ;
  assign n39 = ~m_pad & ~t_pad ;
  assign n41 = n38 & ~n39 ;
  assign n42 = ~n40 & n41 ;
  assign n43 = ~n37 & ~n42 ;
  assign n44 = ~u_pad & ~v_pad ;
  assign n46 = t_pad & w_pad ;
  assign n45 = ~d_pad & ~t_pad ;
  assign n47 = n38 & ~n45 ;
  assign n48 = ~n46 & n47 ;
  assign n49 = ~n44 & ~n48 ;
  assign n50 = ~u_pad & ~w_pad ;
  assign n52 = t_pad & x_pad ;
  assign n51 = ~c_pad & ~t_pad ;
  assign n53 = n38 & ~n51 ;
  assign n54 = ~n52 & n53 ;
  assign n55 = ~n50 & ~n54 ;
  assign n56 = ~u_pad & ~x_pad ;
  assign n58 = t_pad & y_pad ;
  assign n57 = ~b_pad & ~t_pad ;
  assign n59 = n38 & ~n57 ;
  assign n60 = ~n58 & n59 ;
  assign n61 = ~n56 & ~n60 ;
  assign n62 = ~u_pad & ~y_pad ;
  assign n64 = ~q_pad & t_pad ;
  assign n63 = ~a_pad & ~t_pad ;
  assign n65 = n38 & ~n63 ;
  assign n66 = ~n64 & n65 ;
  assign n67 = ~n62 & ~n66 ;
  assign n68 = ~u_pad & ~z_pad ;
  assign n70 = \a0_pad  & t_pad ;
  assign n69 = ~h_pad & ~t_pad ;
  assign n71 = n38 & ~n69 ;
  assign n72 = ~n70 & n71 ;
  assign n73 = ~n68 & ~n72 ;
  assign n74 = ~\a0_pad  & ~u_pad ;
  assign n76 = \b0_pad  & t_pad ;
  assign n75 = ~g_pad & ~t_pad ;
  assign n77 = n38 & ~n75 ;
  assign n78 = ~n76 & n77 ;
  assign n79 = ~n74 & ~n78 ;
  assign n80 = ~\b0_pad  & ~u_pad ;
  assign n82 = \c0_pad  & t_pad ;
  assign n81 = ~f_pad & ~t_pad ;
  assign n83 = n38 & ~n81 ;
  assign n84 = ~n82 & n83 ;
  assign n85 = ~n80 & ~n84 ;
  assign n86 = ~\c0_pad  & ~u_pad ;
  assign n88 = t_pad & v_pad ;
  assign n87 = ~e_pad & ~t_pad ;
  assign n89 = n38 & ~n87 ;
  assign n90 = ~n88 & n89 ;
  assign n91 = ~n86 & ~n90 ;
  assign n92 = ~\d0_pad  & ~u_pad ;
  assign n94 = \e0_pad  & t_pad ;
  assign n93 = ~l_pad & ~t_pad ;
  assign n95 = n38 & ~n93 ;
  assign n96 = ~n94 & n95 ;
  assign n97 = ~n92 & ~n96 ;
  assign n98 = ~\e0_pad  & ~u_pad ;
  assign n100 = \f0_pad  & t_pad ;
  assign n99 = ~k_pad & ~t_pad ;
  assign n101 = n38 & ~n99 ;
  assign n102 = ~n100 & n101 ;
  assign n103 = ~n98 & ~n102 ;
  assign n104 = ~\f0_pad  & ~u_pad ;
  assign n106 = \g0_pad  & t_pad ;
  assign n105 = ~j_pad & ~t_pad ;
  assign n107 = n38 & ~n105 ;
  assign n108 = ~n106 & n107 ;
  assign n109 = ~n104 & ~n108 ;
  assign n110 = ~\g0_pad  & ~u_pad ;
  assign n112 = t_pad & z_pad ;
  assign n111 = ~i_pad & ~t_pad ;
  assign n113 = n38 & ~n111 ;
  assign n114 = ~n112 & n113 ;
  assign n115 = ~n110 & ~n114 ;
  assign n116 = ~\h0_pad  & ~u_pad ;
  assign n118 = \i0_pad  & t_pad ;
  assign n117 = ~p_pad & ~t_pad ;
  assign n119 = n38 & ~n117 ;
  assign n120 = ~n118 & n119 ;
  assign n121 = ~n116 & ~n120 ;
  assign n122 = ~\i0_pad  & ~u_pad ;
  assign n124 = \j0_pad  & t_pad ;
  assign n123 = ~o_pad & ~t_pad ;
  assign n125 = n38 & ~n123 ;
  assign n126 = ~n124 & n125 ;
  assign n127 = ~n122 & ~n126 ;
  assign n128 = ~\j0_pad  & ~u_pad ;
  assign n130 = \k0_pad  & t_pad ;
  assign n129 = ~n_pad & ~t_pad ;
  assign n131 = n38 & ~n129 ;
  assign n132 = ~n130 & n131 ;
  assign n133 = ~n128 & ~n132 ;
  assign \a1_pad  = ~n43 ;
  assign \l0_pad  = ~n49 ;
  assign \m0_pad  = ~n55 ;
  assign \n0_pad  = ~n61 ;
  assign \o0_pad  = ~n67 ;
  assign \p0_pad  = ~n73 ;
  assign \q0_pad  = ~n79 ;
  assign \r0_pad  = ~n85 ;
  assign \s0_pad  = ~n91 ;
  assign \t0_pad  = ~n97 ;
  assign \u0_pad  = ~n103 ;
  assign \v0_pad  = ~n109 ;
  assign \w0_pad  = ~n115 ;
  assign \x0_pad  = ~n121 ;
  assign \y0_pad  = ~n127 ;
  assign \z0_pad  = ~n133 ;
endmodule
