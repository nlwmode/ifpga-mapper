module top( \al_reg/NET0131  , \byte_controller_ack_out_reg/NET0131  , \byte_controller_bit_controller_al_reg/NET0131  , \byte_controller_bit_controller_busy_reg/NET0131  , \byte_controller_bit_controller_c_state_reg[0]/NET0131  , \byte_controller_bit_controller_c_state_reg[10]/NET0131  , \byte_controller_bit_controller_c_state_reg[11]/NET0131  , \byte_controller_bit_controller_c_state_reg[12]/NET0131  , \byte_controller_bit_controller_c_state_reg[13]/NET0131  , \byte_controller_bit_controller_c_state_reg[14]/NET0131  , \byte_controller_bit_controller_c_state_reg[15]/NET0131  , \byte_controller_bit_controller_c_state_reg[16]/NET0131  , \byte_controller_bit_controller_c_state_reg[1]/NET0131  , \byte_controller_bit_controller_c_state_reg[2]/NET0131  , \byte_controller_bit_controller_c_state_reg[3]/NET0131  , \byte_controller_bit_controller_c_state_reg[4]/NET0131  , \byte_controller_bit_controller_c_state_reg[5]/NET0131  , \byte_controller_bit_controller_c_state_reg[6]/NET0131  , \byte_controller_bit_controller_c_state_reg[7]/NET0131  , \byte_controller_bit_controller_c_state_reg[8]/NET0131  , \byte_controller_bit_controller_c_state_reg[9]/NET0131  , \byte_controller_bit_controller_clk_en_reg/NET0131  , \byte_controller_bit_controller_cmd_ack_reg/NET0131  , \byte_controller_bit_controller_cmd_stop_reg/NET0131  , \byte_controller_bit_controller_cnt_reg[0]/NET0131  , \byte_controller_bit_controller_cnt_reg[10]/NET0131  , \byte_controller_bit_controller_cnt_reg[11]/NET0131  , \byte_controller_bit_controller_cnt_reg[12]/NET0131  , \byte_controller_bit_controller_cnt_reg[13]/NET0131  , \byte_controller_bit_controller_cnt_reg[14]/NET0131  , \byte_controller_bit_controller_cnt_reg[15]/NET0131  , \byte_controller_bit_controller_cnt_reg[1]/NET0131  , \byte_controller_bit_controller_cnt_reg[2]/NET0131  , \byte_controller_bit_controller_cnt_reg[3]/NET0131  , \byte_controller_bit_controller_cnt_reg[4]/NET0131  , \byte_controller_bit_controller_cnt_reg[5]/NET0131  , \byte_controller_bit_controller_cnt_reg[6]/NET0131  , \byte_controller_bit_controller_cnt_reg[7]/NET0131  , \byte_controller_bit_controller_cnt_reg[8]/NET0131  , \byte_controller_bit_controller_cnt_reg[9]/NET0131  , \byte_controller_bit_controller_dSCL_reg/NET0131  , \byte_controller_bit_controller_dSDA_reg/NET0131  , \byte_controller_bit_controller_dout_reg/P0001  , \byte_controller_bit_controller_dscl_oen_reg/P0001  , \byte_controller_bit_controller_sSCL_reg/NET0131  , \byte_controller_bit_controller_sSDA_reg/NET0131  , \byte_controller_bit_controller_sda_chk_reg/NET0131  , \byte_controller_bit_controller_sta_condition_reg/NET0131  , \byte_controller_bit_controller_sto_condition_reg/NET0131  , \byte_controller_c_state_reg[0]/NET0131  , \byte_controller_c_state_reg[1]/NET0131  , \byte_controller_c_state_reg[2]/NET0131  , \byte_controller_c_state_reg[3]/NET0131  , \byte_controller_c_state_reg[4]/NET0131  , \byte_controller_cmd_ack_reg/NET0131  , \byte_controller_core_cmd_reg[2]/NET0131  , \byte_controller_core_cmd_reg[3]/NET0131  , \byte_controller_core_txd_reg/NET0131  , \byte_controller_dcnt_reg[0]/NET0131  , \byte_controller_dcnt_reg[1]/NET0131  , \byte_controller_dcnt_reg[2]/NET0131  , \byte_controller_ld_reg/NET0131  , \byte_controller_shift_reg/NET0131  , \byte_controller_sr_reg[0]/NET0131  , \byte_controller_sr_reg[1]/NET0131  , \byte_controller_sr_reg[2]/NET0131  , \byte_controller_sr_reg[3]/NET0131  , \byte_controller_sr_reg[4]/NET0131  , \byte_controller_sr_reg[5]/NET0131  , \byte_controller_sr_reg[6]/NET0131  , \byte_controller_sr_reg[7]/NET0131  , \cr_reg[0]/NET0131  , \cr_reg[1]/NET0131  , \cr_reg[2]/NET0131  , \cr_reg[3]/NET0131  , \cr_reg[4]/NET0131  , \cr_reg[5]/NET0131  , \cr_reg[6]/NET0131  , \cr_reg[7]/NET0131  , \ctr_reg[0]/NET0131  , \ctr_reg[1]/NET0131  , \ctr_reg[2]/NET0131  , \ctr_reg[3]/NET0131  , \ctr_reg[4]/NET0131  , \ctr_reg[5]/NET0131  , \ctr_reg[6]/NET0131  , \ctr_reg[7]/NET0131  , \irq_flag_reg/NET0131  , \prer_reg[0]/NET0131  , \prer_reg[10]/NET0131  , \prer_reg[11]/NET0131  , \prer_reg[12]/NET0131  , \prer_reg[13]/NET0131  , \prer_reg[14]/NET0131  , \prer_reg[15]/NET0131  , \prer_reg[1]/NET0131  , \prer_reg[2]/NET0131  , \prer_reg[3]/NET0131  , \prer_reg[4]/NET0131  , \prer_reg[5]/NET0131  , \prer_reg[6]/NET0131  , \prer_reg[7]/NET0131  , \prer_reg[8]/NET0131  , \prer_reg[9]/NET0131  , \rxack_reg/NET0131  , scl_pad_i_pad , scl_padoen_o_pad , sda_pad_i_pad , sda_padoen_o_pad , \tip_reg/NET0131  , \txr_reg[0]/NET0131  , \txr_reg[1]/NET0131  , \txr_reg[2]/NET0131  , \txr_reg[3]/NET0131  , \txr_reg[4]/NET0131  , \txr_reg[5]/NET0131  , \txr_reg[6]/NET0131  , \txr_reg[7]/NET0131  , wb_ack_o_pad , \wb_adr_i[0]_pad  , \wb_adr_i[1]_pad  , \wb_adr_i[2]_pad  , wb_cyc_i_pad , \wb_dat_i[0]_pad  , \wb_dat_i[1]_pad  , \wb_dat_i[2]_pad  , \wb_dat_i[3]_pad  , \wb_dat_i[4]_pad  , \wb_dat_i[5]_pad  , \wb_dat_i[6]_pad  , \wb_dat_i[7]_pad  , wb_rst_i_pad , wb_stb_i_pad , wb_we_i_pad , \_al_n1  , \byte_controller_bit_controller_dout_reg/P0001_reg_syn_3  , \g3074/_0_  , \g3075/_0_  , \g3102/_0_  , \g3106/_0_  , \g3117/_0_  , \g3120/_0_  , \g3127/_0_  , \g3128/_0_  , \g3129/_0_  , \g3130/_0_  , \g3131/_0_  , \g3132/_0_  , \g3160/_0_  , \g3164/_0_  , \g3166/_0_  , \g3167/_0_  , \g3171/_0_  , \g3174/_3_  , \g3184/_0_  , \g3185/_0_  , \g3188/_0_  , \g3193/_0_  , \g3195/_0_  , \g3198/_0_  , \g3199/_0_  , \g32/_1_  , \g3200/_0_  , \g3201/_0_  , \g3203/_0_  , \g3204/_0_  , \g3205/_0_  , \g3206/_0_  , \g3207/_0_  , \g3208/_0_  , \g3209/_0_  , \g3211/_0_  , \g3246/_0_  , \g3250/_2_  , \g3251/_0_  , \g3255/_0_  , \g3256/_0_  , \g3259/_0_  , \g3262/_0_  , \g3269/_0_  , \g3270/_0_  , \g3271/_0_  , \g3272/_0_  , \g3273/_0_  , \g3274/_0_  , \g3275/_0_  , \g3276/_0_  , \g3277/_0_  , \g3278/_0_  , \g3279/_0_  , \g3280/_0_  , \g3281/_0_  , \g3282/_0_  , \g3283/_0_  , \g3284/_0_  , \g3285/_0_  , \g3286/_0_  , \g3307/_0_  , \g3339/_0_  , \g3392/_0_  , \g3419/_0_  , \g3421/_0_  , \g3422/_0_  , \g3423/_0_  , \g3424/_0_  , \g3425/_0_  , \g3426/_0_  , \g3427/_0_  , \g3428/_0_  , \g3429/_0_  , \g3430/_0_  , \g3431/_0_  , \g3452/_0_  , \g3453/_0_  , \g3454/_0_  , \g3455/_0_  , \g3456/_0_  , \g3457/_0_  , \g3458/_0_  , \g3459/_0_  , \g3460/_0_  , \g3462/_0_  , \g3464/_0_  , \g3465/_0_  , \g3471/_0_  , \g3472/_0_  , \g3476/_0_  , \g3477/_0_  , \g3478/_0_  , \g3479/_0_  , \g3499/_0_  , \g3506/_0_  , \g3507/_0_  , \g3591/_0_  , \g3601/_0_  , \g3602/_0_  , \g3603/_0_  , \g3693/_0_  , \g3694/_0_  , \g3761/_0_  , \g3785/_0_  , \g3798/_0_  , \g3815/_1_  , \g3840/_0_  , \g3874/_0_  , \g3915/_0_  , \g3927/_2_  , \g3978/_0_  , \g4004/_0_  , \g4021/_0_  , \g4582/_0_  , \g4804/_0_  , \g4866/_0_  , \g4876/_0_  , \g4942/_0_  , \g4996/_0_  , \g5146/_0_  , \g5236/_0_  , \g5411/_0_  , \g5433/_0_  , scl_pad_o_pad );
  input \al_reg/NET0131  ;
  input \byte_controller_ack_out_reg/NET0131  ;
  input \byte_controller_bit_controller_al_reg/NET0131  ;
  input \byte_controller_bit_controller_busy_reg/NET0131  ;
  input \byte_controller_bit_controller_c_state_reg[0]/NET0131  ;
  input \byte_controller_bit_controller_c_state_reg[10]/NET0131  ;
  input \byte_controller_bit_controller_c_state_reg[11]/NET0131  ;
  input \byte_controller_bit_controller_c_state_reg[12]/NET0131  ;
  input \byte_controller_bit_controller_c_state_reg[13]/NET0131  ;
  input \byte_controller_bit_controller_c_state_reg[14]/NET0131  ;
  input \byte_controller_bit_controller_c_state_reg[15]/NET0131  ;
  input \byte_controller_bit_controller_c_state_reg[16]/NET0131  ;
  input \byte_controller_bit_controller_c_state_reg[1]/NET0131  ;
  input \byte_controller_bit_controller_c_state_reg[2]/NET0131  ;
  input \byte_controller_bit_controller_c_state_reg[3]/NET0131  ;
  input \byte_controller_bit_controller_c_state_reg[4]/NET0131  ;
  input \byte_controller_bit_controller_c_state_reg[5]/NET0131  ;
  input \byte_controller_bit_controller_c_state_reg[6]/NET0131  ;
  input \byte_controller_bit_controller_c_state_reg[7]/NET0131  ;
  input \byte_controller_bit_controller_c_state_reg[8]/NET0131  ;
  input \byte_controller_bit_controller_c_state_reg[9]/NET0131  ;
  input \byte_controller_bit_controller_clk_en_reg/NET0131  ;
  input \byte_controller_bit_controller_cmd_ack_reg/NET0131  ;
  input \byte_controller_bit_controller_cmd_stop_reg/NET0131  ;
  input \byte_controller_bit_controller_cnt_reg[0]/NET0131  ;
  input \byte_controller_bit_controller_cnt_reg[10]/NET0131  ;
  input \byte_controller_bit_controller_cnt_reg[11]/NET0131  ;
  input \byte_controller_bit_controller_cnt_reg[12]/NET0131  ;
  input \byte_controller_bit_controller_cnt_reg[13]/NET0131  ;
  input \byte_controller_bit_controller_cnt_reg[14]/NET0131  ;
  input \byte_controller_bit_controller_cnt_reg[15]/NET0131  ;
  input \byte_controller_bit_controller_cnt_reg[1]/NET0131  ;
  input \byte_controller_bit_controller_cnt_reg[2]/NET0131  ;
  input \byte_controller_bit_controller_cnt_reg[3]/NET0131  ;
  input \byte_controller_bit_controller_cnt_reg[4]/NET0131  ;
  input \byte_controller_bit_controller_cnt_reg[5]/NET0131  ;
  input \byte_controller_bit_controller_cnt_reg[6]/NET0131  ;
  input \byte_controller_bit_controller_cnt_reg[7]/NET0131  ;
  input \byte_controller_bit_controller_cnt_reg[8]/NET0131  ;
  input \byte_controller_bit_controller_cnt_reg[9]/NET0131  ;
  input \byte_controller_bit_controller_dSCL_reg/NET0131  ;
  input \byte_controller_bit_controller_dSDA_reg/NET0131  ;
  input \byte_controller_bit_controller_dout_reg/P0001  ;
  input \byte_controller_bit_controller_dscl_oen_reg/P0001  ;
  input \byte_controller_bit_controller_sSCL_reg/NET0131  ;
  input \byte_controller_bit_controller_sSDA_reg/NET0131  ;
  input \byte_controller_bit_controller_sda_chk_reg/NET0131  ;
  input \byte_controller_bit_controller_sta_condition_reg/NET0131  ;
  input \byte_controller_bit_controller_sto_condition_reg/NET0131  ;
  input \byte_controller_c_state_reg[0]/NET0131  ;
  input \byte_controller_c_state_reg[1]/NET0131  ;
  input \byte_controller_c_state_reg[2]/NET0131  ;
  input \byte_controller_c_state_reg[3]/NET0131  ;
  input \byte_controller_c_state_reg[4]/NET0131  ;
  input \byte_controller_cmd_ack_reg/NET0131  ;
  input \byte_controller_core_cmd_reg[2]/NET0131  ;
  input \byte_controller_core_cmd_reg[3]/NET0131  ;
  input \byte_controller_core_txd_reg/NET0131  ;
  input \byte_controller_dcnt_reg[0]/NET0131  ;
  input \byte_controller_dcnt_reg[1]/NET0131  ;
  input \byte_controller_dcnt_reg[2]/NET0131  ;
  input \byte_controller_ld_reg/NET0131  ;
  input \byte_controller_shift_reg/NET0131  ;
  input \byte_controller_sr_reg[0]/NET0131  ;
  input \byte_controller_sr_reg[1]/NET0131  ;
  input \byte_controller_sr_reg[2]/NET0131  ;
  input \byte_controller_sr_reg[3]/NET0131  ;
  input \byte_controller_sr_reg[4]/NET0131  ;
  input \byte_controller_sr_reg[5]/NET0131  ;
  input \byte_controller_sr_reg[6]/NET0131  ;
  input \byte_controller_sr_reg[7]/NET0131  ;
  input \cr_reg[0]/NET0131  ;
  input \cr_reg[1]/NET0131  ;
  input \cr_reg[2]/NET0131  ;
  input \cr_reg[3]/NET0131  ;
  input \cr_reg[4]/NET0131  ;
  input \cr_reg[5]/NET0131  ;
  input \cr_reg[6]/NET0131  ;
  input \cr_reg[7]/NET0131  ;
  input \ctr_reg[0]/NET0131  ;
  input \ctr_reg[1]/NET0131  ;
  input \ctr_reg[2]/NET0131  ;
  input \ctr_reg[3]/NET0131  ;
  input \ctr_reg[4]/NET0131  ;
  input \ctr_reg[5]/NET0131  ;
  input \ctr_reg[6]/NET0131  ;
  input \ctr_reg[7]/NET0131  ;
  input \irq_flag_reg/NET0131  ;
  input \prer_reg[0]/NET0131  ;
  input \prer_reg[10]/NET0131  ;
  input \prer_reg[11]/NET0131  ;
  input \prer_reg[12]/NET0131  ;
  input \prer_reg[13]/NET0131  ;
  input \prer_reg[14]/NET0131  ;
  input \prer_reg[15]/NET0131  ;
  input \prer_reg[1]/NET0131  ;
  input \prer_reg[2]/NET0131  ;
  input \prer_reg[3]/NET0131  ;
  input \prer_reg[4]/NET0131  ;
  input \prer_reg[5]/NET0131  ;
  input \prer_reg[6]/NET0131  ;
  input \prer_reg[7]/NET0131  ;
  input \prer_reg[8]/NET0131  ;
  input \prer_reg[9]/NET0131  ;
  input \rxack_reg/NET0131  ;
  input scl_pad_i_pad ;
  input scl_padoen_o_pad ;
  input sda_pad_i_pad ;
  input sda_padoen_o_pad ;
  input \tip_reg/NET0131  ;
  input \txr_reg[0]/NET0131  ;
  input \txr_reg[1]/NET0131  ;
  input \txr_reg[2]/NET0131  ;
  input \txr_reg[3]/NET0131  ;
  input \txr_reg[4]/NET0131  ;
  input \txr_reg[5]/NET0131  ;
  input \txr_reg[6]/NET0131  ;
  input \txr_reg[7]/NET0131  ;
  input wb_ack_o_pad ;
  input \wb_adr_i[0]_pad  ;
  input \wb_adr_i[1]_pad  ;
  input \wb_adr_i[2]_pad  ;
  input wb_cyc_i_pad ;
  input \wb_dat_i[0]_pad  ;
  input \wb_dat_i[1]_pad  ;
  input \wb_dat_i[2]_pad  ;
  input \wb_dat_i[3]_pad  ;
  input \wb_dat_i[4]_pad  ;
  input \wb_dat_i[5]_pad  ;
  input \wb_dat_i[6]_pad  ;
  input \wb_dat_i[7]_pad  ;
  input wb_rst_i_pad ;
  input wb_stb_i_pad ;
  input wb_we_i_pad ;
  output \_al_n1  ;
  output \byte_controller_bit_controller_dout_reg/P0001_reg_syn_3  ;
  output \g3074/_0_  ;
  output \g3075/_0_  ;
  output \g3102/_0_  ;
  output \g3106/_0_  ;
  output \g3117/_0_  ;
  output \g3120/_0_  ;
  output \g3127/_0_  ;
  output \g3128/_0_  ;
  output \g3129/_0_  ;
  output \g3130/_0_  ;
  output \g3131/_0_  ;
  output \g3132/_0_  ;
  output \g3160/_0_  ;
  output \g3164/_0_  ;
  output \g3166/_0_  ;
  output \g3167/_0_  ;
  output \g3171/_0_  ;
  output \g3174/_3_  ;
  output \g3184/_0_  ;
  output \g3185/_0_  ;
  output \g3188/_0_  ;
  output \g3193/_0_  ;
  output \g3195/_0_  ;
  output \g3198/_0_  ;
  output \g3199/_0_  ;
  output \g32/_1_  ;
  output \g3200/_0_  ;
  output \g3201/_0_  ;
  output \g3203/_0_  ;
  output \g3204/_0_  ;
  output \g3205/_0_  ;
  output \g3206/_0_  ;
  output \g3207/_0_  ;
  output \g3208/_0_  ;
  output \g3209/_0_  ;
  output \g3211/_0_  ;
  output \g3246/_0_  ;
  output \g3250/_2_  ;
  output \g3251/_0_  ;
  output \g3255/_0_  ;
  output \g3256/_0_  ;
  output \g3259/_0_  ;
  output \g3262/_0_  ;
  output \g3269/_0_  ;
  output \g3270/_0_  ;
  output \g3271/_0_  ;
  output \g3272/_0_  ;
  output \g3273/_0_  ;
  output \g3274/_0_  ;
  output \g3275/_0_  ;
  output \g3276/_0_  ;
  output \g3277/_0_  ;
  output \g3278/_0_  ;
  output \g3279/_0_  ;
  output \g3280/_0_  ;
  output \g3281/_0_  ;
  output \g3282/_0_  ;
  output \g3283/_0_  ;
  output \g3284/_0_  ;
  output \g3285/_0_  ;
  output \g3286/_0_  ;
  output \g3307/_0_  ;
  output \g3339/_0_  ;
  output \g3392/_0_  ;
  output \g3419/_0_  ;
  output \g3421/_0_  ;
  output \g3422/_0_  ;
  output \g3423/_0_  ;
  output \g3424/_0_  ;
  output \g3425/_0_  ;
  output \g3426/_0_  ;
  output \g3427/_0_  ;
  output \g3428/_0_  ;
  output \g3429/_0_  ;
  output \g3430/_0_  ;
  output \g3431/_0_  ;
  output \g3452/_0_  ;
  output \g3453/_0_  ;
  output \g3454/_0_  ;
  output \g3455/_0_  ;
  output \g3456/_0_  ;
  output \g3457/_0_  ;
  output \g3458/_0_  ;
  output \g3459/_0_  ;
  output \g3460/_0_  ;
  output \g3462/_0_  ;
  output \g3464/_0_  ;
  output \g3465/_0_  ;
  output \g3471/_0_  ;
  output \g3472/_0_  ;
  output \g3476/_0_  ;
  output \g3477/_0_  ;
  output \g3478/_0_  ;
  output \g3479/_0_  ;
  output \g3499/_0_  ;
  output \g3506/_0_  ;
  output \g3507/_0_  ;
  output \g3591/_0_  ;
  output \g3601/_0_  ;
  output \g3602/_0_  ;
  output \g3603/_0_  ;
  output \g3693/_0_  ;
  output \g3694/_0_  ;
  output \g3761/_0_  ;
  output \g3785/_0_  ;
  output \g3798/_0_  ;
  output \g3815/_1_  ;
  output \g3840/_0_  ;
  output \g3874/_0_  ;
  output \g3915/_0_  ;
  output \g3927/_2_  ;
  output \g3978/_0_  ;
  output \g4004/_0_  ;
  output \g4021/_0_  ;
  output \g4582/_0_  ;
  output \g4804/_0_  ;
  output \g4866/_0_  ;
  output \g4876/_0_  ;
  output \g4942/_0_  ;
  output \g4996/_0_  ;
  output \g5146/_0_  ;
  output \g5236/_0_  ;
  output \g5411/_0_  ;
  output \g5433/_0_  ;
  output scl_pad_o_pad ;
  wire n135 , n136 , n137 , n138 , n139 , n140 , n141 , n142 , n143 , n144 , n145 , n146 , n147 , n148 , n149 , n150 , n151 , n152 , n153 , n154 , n155 , n156 , n157 , n158 , n159 , n160 , n161 , n162 , n163 , n164 , n165 , n166 , n167 , n168 , n169 , n170 , n171 , n172 , n173 , n174 , n175 , n176 , n177 , n178 , n179 , n180 , n181 , n182 , n183 , n184 , n185 , n186 , n187 , n188 , n189 , n190 , n191 , n192 , n193 , n194 , n195 , n196 , n197 , n198 , n199 , n200 , n201 , n202 , n203 , n204 , n205 , n206 , n207 , n208 , n209 , n210 , n211 , n212 , n213 , n214 , n215 , n216 , n217 , n218 , n219 , n220 , n221 , n222 , n223 , n224 , n225 , n226 , n227 , n228 , n229 , n230 , n231 , n232 , n233 , n234 , n235 , n236 , n237 , n238 , n239 , n240 , n241 , n242 , n243 , n244 , n245 , n246 , n247 , n248 , n249 , n250 , n251 , n252 , n253 , n254 , n255 , n256 , n257 , n258 , n259 , n260 , n261 , n262 , n263 , n264 , n265 , n266 , n267 , n268 , n269 , n270 , n271 , n272 , n273 , n274 , n275 , n276 , n277 , n278 , n279 , n280 , n281 , n282 , n283 , n284 , n285 , n286 , n287 , n288 , n289 , n290 , n291 , n292 , n293 , n294 , n295 , n296 , n297 , n298 , n299 , n300 , n301 , n302 , n303 , n304 , n305 , n306 , n307 , n308 , n309 , n310 , n311 , n312 , n313 , n314 , n315 , n316 , n317 , n318 , n319 , n320 , n321 , n322 , n323 , n324 , n325 , n326 , n327 , n328 , n329 , n330 , n331 , n332 , n333 , n334 , n335 , n336 , n337 , n338 , n339 , n340 , n341 , n342 , n343 , n344 , n345 , n346 , n347 , n348 , n349 , n350 , n351 , n352 , n353 , n354 , n355 , n356 , n357 , n358 , n359 , n360 , n361 , n362 , n363 , n364 , n365 , n366 , n367 , n368 , n369 , n370 , n371 , n372 , n373 , n374 , n375 , n376 , n377 , n378 , n379 , n380 , n381 , n382 , n383 , n384 , n385 , n386 , n387 , n388 , n389 , n390 , n391 , n392 , n393 , n394 , n395 , n396 , n397 , n398 , n399 , n400 , n401 , n402 , n403 , n404 , n405 , n406 , n407 , n408 , n409 , n410 , n411 , n412 , n413 , n414 , n415 , n416 , n417 , n418 , n419 , n420 , n421 , n422 , n423 , n424 , n425 , n426 , n427 , n428 , n429 , n430 , n431 , n432 , n433 , n434 , n435 , n436 , n437 , n438 , n439 , n440 , n441 , n442 , n443 , n444 , n445 , n446 , n447 , n448 , n449 , n450 , n451 , n452 , n453 , n454 , n455 , n456 , n457 , n458 , n459 , n460 , n461 , n462 , n463 , n464 , n465 , n466 , n467 , n468 , n469 , n470 , n471 , n472 , n473 , n474 , n475 , n476 , n477 , n478 , n479 , n480 , n481 , n482 , n483 , n484 , n485 , n486 , n487 , n488 , n489 , n490 , n491 , n492 , n493 , n494 , n495 , n496 , n497 , n498 , n499 , n500 , n501 , n502 , n503 , n504 , n505 , n506 , n507 , n508 , n509 , n510 , n511 , n512 , n513 , n514 , n515 , n516 , n517 , n518 , n519 , n520 , n521 , n522 , n523 , n524 , n525 , n526 , n527 , n528 , n529 , n530 , n531 , n532 , n533 , n534 , n535 , n536 , n537 , n538 , n539 , n540 , n541 , n542 , n543 , n544 , n545 , n546 , n547 , n548 , n549 , n550 , n551 , n552 , n553 , n554 , n555 , n556 , n557 , n558 , n559 , n560 , n561 , n562 , n563 , n564 , n565 , n566 , n567 , n568 , n569 , n570 , n571 , n572 , n573 , n574 , n575 , n576 , n577 , n578 , n579 , n580 , n581 , n582 , n583 , n584 , n585 , n586 , n587 , n588 , n589 , n590 , n591 , n592 , n593 , n594 , n595 , n596 , n597 , n598 , n599 , n600 , n601 , n602 , n603 , n604 , n605 , n606 , n607 , n608 , n609 , n610 , n611 , n612 , n613 , n614 , n615 , n616 , n617 , n618 , n619 , n620 , n621 , n622 , n623 , n624 , n625 , n626 , n627 , n628 , n629 , n630 , n631 , n632 , n633 , n634 , n635 , n636 , n637 , n638 , n639 , n640 , n641 , n642 , n643 , n644 , n645 , n646 , n647 , n648 , n649 , n650 , n651 , n652 , n653 , n654 , n655 , n656 , n657 , n658 , n659 , n660 , n661 , n662 , n663 , n664 , n665 , n666 , n667 , n668 , n669 , n670 , n671 , n672 , n673 , n674 , n675 , n676 , n677 , n678 , n679 , n680 , n681 , n682 , n683 , n684 , n685 , n686 , n687 , n688 , n689 , n690 , n691 , n692 , n693 , n694 , n695 , n696 , n697 , n698 , n699 , n700 , n701 , n702 , n703 , n704 , n705 , n706 , n707 , n708 , n709 , n710 , n711 , n712 , n713 , n714 , n715 , n716 , n717 , n718 , n719 , n720 , n721 , n722 , n723 , n724 , n725 , n726 , n727 , n728 , n729 , n730 , n731 , n732 , n733 , n734 , n735 , n736 , n737 , n738 , n739 , n740 , n741 , n742 , n743 , n744 , n745 , n746 , n747 , n748 , n749 , n750 , n751 , n752 , n753 , n754 , n755 , n756 , n757 , n758 , n759 , n760 , n761 , n762 , n763 , n764 , n765 , n766 , n767 , n768 , n769 , n770 , n771 , n772 , n773 , n774 , n775 , n776 , n777 , n778 , n779 , n780 , n781 , n782 , n783 , n784 , n785 , n786 , n787 , n788 , n789 , n790 , n791 , n792 , n793 , n794 , n795 , n796 , n797 , n798 , n799 , n800 , n801 , n802 , n803 , n804 , n805 , n806 , n807 , n808 , n809 , n810 , n811 , n812 , n813 , n814 , n815 , n816 , n817 , n818 , n819 , n820 , n821 , n822 , n823 , n824 , n825 , n826 , n827 , n828 , n829 , n830 , n831 , n832 , n833 , n834 , n835 , n836 , n837 , n838 , n839 , n840 , n841 , n842 , n843 , n844 , n845 , n846 , n847 , n848 , n849 , n850 , n851 , n852 , n853 , n854 , n855 , n856 , n857 , n858 , n859 , n860 , n861 , n862 , n863 , n864 , n865 , n866 , n867 , n868 , n869 , n870 , n871 , n872 , n873 , n874 , n875 , n876 , n877 , n878 , n879 , n880 , n881 , n882 , n883 , n884 , n885 , n886 , n887 , n888 , n889 , n890 , n891 , n892 , n893 , n894 , n895 , n896 , n897 , n898 , n899 , n900 , n901 , n902 , n903 , n904 , n905 , n906 , n907 , n908 , n909 , n910 , n911 , n912 , n913 , n914 , n915 , n916 , n917 , n918 , n919 , n920 , n921 , n922 , n923 , n924 , n925 , n926 , n927 , n928 , n929 , n930 , n931 , n932 , n933 , n934 , n935 , n936 , n937 , n938 , n939 , n940 , n941 , n942 , n943 , n944 , n945 , n946 , n947 , n948 , n949 , n950 , n951 , n952 , n953 , n954 , n955 , n956 , n957 , n958 , n959 , n960 , n961 , n962 , n963 , n964 , n965 , n966 , n967 , n968 , n969 , n970 , n971 , n972 , n973 , n974 , n975 , n976 , n977 , n978 , n979 , n980 , n981 , n982 , n983 , n984 , n985 , n986 , n987 , n988 , n989 , n990 , n991 , n992 , n993 , n994 , n995 , n996 , n997 , n998 , n999 , n1000 , n1001 , n1002 , n1003 , n1004 , n1005 , n1006 ;
  assign n135 = ~\byte_controller_bit_controller_dSCL_reg/NET0131  & \byte_controller_bit_controller_sSCL_reg/NET0131  ;
  assign n136 = \byte_controller_bit_controller_dout_reg/P0001  & ~n135 ;
  assign n137 = \byte_controller_bit_controller_sSDA_reg/NET0131  & n135 ;
  assign n138 = ~n136 & ~n137 ;
  assign n139 = ~\byte_controller_bit_controller_al_reg/NET0131  & ~wb_rst_i_pad ;
  assign n140 = ~\byte_controller_bit_controller_clk_en_reg/NET0131  & ~sda_padoen_o_pad ;
  assign n141 = ~\byte_controller_bit_controller_c_state_reg[0]/NET0131  & ~\byte_controller_bit_controller_c_state_reg[1]/NET0131  ;
  assign n142 = ~\byte_controller_bit_controller_c_state_reg[11]/NET0131  & ~\byte_controller_bit_controller_c_state_reg[13]/NET0131  ;
  assign n143 = ~\byte_controller_bit_controller_c_state_reg[10]/NET0131  & ~\byte_controller_bit_controller_c_state_reg[12]/NET0131  ;
  assign n144 = n142 & n143 ;
  assign n145 = ~\byte_controller_bit_controller_c_state_reg[14]/NET0131  & ~\byte_controller_bit_controller_c_state_reg[15]/NET0131  ;
  assign n146 = ~\byte_controller_bit_controller_c_state_reg[16]/NET0131  & n145 ;
  assign n147 = n144 & n146 ;
  assign n148 = ~\byte_controller_bit_controller_c_state_reg[8]/NET0131  & ~\byte_controller_bit_controller_c_state_reg[9]/NET0131  ;
  assign n149 = n147 & n148 ;
  assign n150 = ~\byte_controller_bit_controller_c_state_reg[6]/NET0131  & ~\byte_controller_bit_controller_c_state_reg[7]/NET0131  ;
  assign n151 = n149 & n150 ;
  assign n152 = \byte_controller_bit_controller_c_state_reg[3]/NET0131  & \byte_controller_bit_controller_c_state_reg[4]/NET0131  ;
  assign n153 = ~\byte_controller_bit_controller_c_state_reg[2]/NET0131  & ~\byte_controller_bit_controller_c_state_reg[5]/NET0131  ;
  assign n154 = ~n152 & n153 ;
  assign n155 = n151 & n154 ;
  assign n159 = ~\byte_controller_bit_controller_c_state_reg[5]/NET0131  & ~\byte_controller_bit_controller_c_state_reg[6]/NET0131  ;
  assign n160 = \byte_controller_bit_controller_c_state_reg[7]/NET0131  & ~n159 ;
  assign n156 = ~\byte_controller_bit_controller_c_state_reg[3]/NET0131  & ~\byte_controller_bit_controller_c_state_reg[4]/NET0131  ;
  assign n157 = ~\byte_controller_bit_controller_c_state_reg[2]/NET0131  & n156 ;
  assign n158 = \byte_controller_bit_controller_c_state_reg[5]/NET0131  & \byte_controller_bit_controller_c_state_reg[6]/NET0131  ;
  assign n161 = n157 & ~n158 ;
  assign n162 = ~n160 & n161 ;
  assign n163 = n149 & n162 ;
  assign n164 = ~n155 & ~n163 ;
  assign n165 = n141 & ~n164 ;
  assign n166 = ~\byte_controller_bit_controller_c_state_reg[15]/NET0131  & ~\byte_controller_bit_controller_c_state_reg[16]/NET0131  ;
  assign n167 = ~\byte_controller_bit_controller_c_state_reg[13]/NET0131  & ~\byte_controller_bit_controller_c_state_reg[14]/NET0131  ;
  assign n168 = ~n166 & ~n167 ;
  assign n169 = ~\byte_controller_bit_controller_c_state_reg[5]/NET0131  & ~\byte_controller_bit_controller_c_state_reg[8]/NET0131  ;
  assign n170 = n150 & n169 ;
  assign n171 = n156 & n170 ;
  assign n172 = ~\byte_controller_bit_controller_c_state_reg[9]/NET0131  & n171 ;
  assign n173 = ~\byte_controller_bit_controller_c_state_reg[0]/NET0131  & ~\byte_controller_bit_controller_c_state_reg[12]/NET0131  ;
  assign n174 = n142 & n173 ;
  assign n175 = ~\byte_controller_bit_controller_c_state_reg[1]/NET0131  & ~\byte_controller_bit_controller_c_state_reg[2]/NET0131  ;
  assign n176 = ~\byte_controller_bit_controller_c_state_reg[10]/NET0131  & n175 ;
  assign n177 = n174 & n176 ;
  assign n178 = ~\byte_controller_bit_controller_c_state_reg[15]/NET0131  & n177 ;
  assign n179 = n172 & n178 ;
  assign n180 = n166 & n167 ;
  assign n181 = ~n179 & n180 ;
  assign n182 = ~n168 & ~n181 ;
  assign n183 = ~\byte_controller_bit_controller_c_state_reg[4]/NET0131  & ~\byte_controller_bit_controller_c_state_reg[5]/NET0131  ;
  assign n184 = ~\byte_controller_bit_controller_c_state_reg[7]/NET0131  & n183 ;
  assign n185 = n149 & n184 ;
  assign n186 = ~\byte_controller_bit_controller_c_state_reg[6]/NET0131  & n185 ;
  assign n187 = ~\byte_controller_bit_controller_c_state_reg[3]/NET0131  & n141 ;
  assign n188 = n186 & n187 ;
  assign n189 = ~n182 & ~n188 ;
  assign n190 = ~n165 & n189 ;
  assign n191 = \byte_controller_core_txd_reg/NET0131  & ~n167 ;
  assign n192 = sda_padoen_o_pad & n167 ;
  assign n193 = n179 & n192 ;
  assign n194 = ~n191 & ~n193 ;
  assign n195 = n166 & ~n194 ;
  assign n196 = \byte_controller_core_txd_reg/NET0131  & ~n166 ;
  assign n197 = n167 & n196 ;
  assign n198 = \byte_controller_bit_controller_clk_en_reg/NET0131  & ~n197 ;
  assign n199 = ~n195 & n198 ;
  assign n200 = ~n190 & n199 ;
  assign n201 = ~n140 & ~n200 ;
  assign n202 = n139 & ~n201 ;
  assign n203 = n146 & n177 ;
  assign n204 = n172 & n203 ;
  assign n205 = \byte_controller_bit_controller_clk_en_reg/NET0131  & ~n204 ;
  assign n206 = ~\byte_controller_bit_controller_c_state_reg[0]/NET0131  & n205 ;
  assign n207 = ~scl_padoen_o_pad & ~n206 ;
  assign n208 = n175 & n206 ;
  assign n209 = ~\byte_controller_bit_controller_c_state_reg[3]/NET0131  & n208 ;
  assign n210 = \byte_controller_bit_controller_c_state_reg[4]/NET0131  & \byte_controller_bit_controller_c_state_reg[5]/NET0131  ;
  assign n211 = n151 & ~n210 ;
  assign n214 = \byte_controller_bit_controller_c_state_reg[12]/NET0131  & ~n180 ;
  assign n212 = ~\byte_controller_bit_controller_c_state_reg[10]/NET0131  & ~\byte_controller_bit_controller_c_state_reg[11]/NET0131  ;
  assign n213 = ~\byte_controller_bit_controller_c_state_reg[9]/NET0131  & n212 ;
  assign n215 = \byte_controller_bit_controller_c_state_reg[13]/NET0131  & \byte_controller_bit_controller_c_state_reg[16]/NET0131  ;
  assign n216 = n145 & ~n215 ;
  assign n217 = n213 & n216 ;
  assign n218 = ~n214 & n217 ;
  assign n219 = ~n147 & ~n218 ;
  assign n220 = ~\byte_controller_bit_controller_c_state_reg[4]/NET0131  & n170 ;
  assign n221 = ~n219 & n220 ;
  assign n222 = ~n211 & ~n221 ;
  assign n223 = n209 & ~n222 ;
  assign n224 = ~n207 & ~n223 ;
  assign n225 = n139 & ~n224 ;
  assign n226 = \byte_controller_bit_controller_c_state_reg[9]/NET0131  & ~\byte_controller_bit_controller_clk_en_reg/NET0131  ;
  assign n228 = \byte_controller_bit_controller_clk_en_reg/NET0131  & ~\byte_controller_c_state_reg[0]/NET0131  ;
  assign n227 = ~\byte_controller_c_state_reg[4]/NET0131  & ~\byte_controller_core_cmd_reg[2]/NET0131  ;
  assign n229 = \byte_controller_core_cmd_reg[3]/NET0131  & n227 ;
  assign n230 = n228 & n229 ;
  assign n231 = n204 & n230 ;
  assign n232 = ~n226 & ~n231 ;
  assign n233 = n139 & ~n232 ;
  assign n234 = \byte_controller_bit_controller_c_state_reg[3]/NET0131  & ~\byte_controller_bit_controller_clk_en_reg/NET0131  ;
  assign n235 = n188 & n205 ;
  assign n236 = ~n234 & ~n235 ;
  assign n237 = n139 & ~n236 ;
  assign n238 = ~\byte_controller_core_cmd_reg[3]/NET0131  & n228 ;
  assign n239 = \byte_controller_c_state_reg[4]/NET0131  & ~\byte_controller_core_cmd_reg[2]/NET0131  ;
  assign n240 = n238 & n239 ;
  assign n241 = n204 & n240 ;
  assign n242 = \byte_controller_bit_controller_c_state_reg[5]/NET0131  & ~\byte_controller_bit_controller_clk_en_reg/NET0131  ;
  assign n243 = ~n241 & ~n242 ;
  assign n244 = n139 & ~n243 ;
  assign n245 = ~\byte_controller_bit_controller_cnt_reg[0]/NET0131  & ~\byte_controller_bit_controller_cnt_reg[1]/NET0131  ;
  assign n246 = ~\byte_controller_bit_controller_cnt_reg[2]/NET0131  & ~\byte_controller_bit_controller_cnt_reg[3]/NET0131  ;
  assign n247 = n245 & n246 ;
  assign n248 = ~\byte_controller_bit_controller_cnt_reg[4]/NET0131  & ~\byte_controller_bit_controller_cnt_reg[5]/NET0131  ;
  assign n249 = n247 & n248 ;
  assign n250 = ~\byte_controller_bit_controller_cnt_reg[6]/NET0131  & ~\byte_controller_bit_controller_cnt_reg[7]/NET0131  ;
  assign n251 = n249 & n250 ;
  assign n252 = ~\byte_controller_bit_controller_cnt_reg[8]/NET0131  & ~\byte_controller_bit_controller_cnt_reg[9]/NET0131  ;
  assign n253 = n251 & n252 ;
  assign n254 = ~\byte_controller_bit_controller_cnt_reg[10]/NET0131  & ~\byte_controller_bit_controller_cnt_reg[11]/NET0131  ;
  assign n255 = n253 & n254 ;
  assign n256 = ~\byte_controller_bit_controller_cnt_reg[12]/NET0131  & ~\byte_controller_bit_controller_cnt_reg[13]/NET0131  ;
  assign n257 = ~\byte_controller_bit_controller_cnt_reg[14]/NET0131  & ~\byte_controller_bit_controller_cnt_reg[15]/NET0131  ;
  assign n258 = n256 & n257 ;
  assign n259 = n255 & n258 ;
  assign n260 = \ctr_reg[7]/NET0131  & ~n259 ;
  assign n261 = ~\byte_controller_bit_controller_cnt_reg[6]/NET0131  & n249 ;
  assign n262 = \byte_controller_bit_controller_cnt_reg[7]/NET0131  & ~n261 ;
  assign n263 = ~n251 & ~n262 ;
  assign n264 = n260 & ~n263 ;
  assign n265 = \byte_controller_bit_controller_dscl_oen_reg/P0001  & ~\byte_controller_bit_controller_sSCL_reg/NET0131  ;
  assign n266 = ~\prer_reg[7]/NET0131  & ~n265 ;
  assign n267 = ~\byte_controller_bit_controller_cnt_reg[7]/NET0131  & n265 ;
  assign n268 = ~n266 & ~n267 ;
  assign n269 = ~n260 & n268 ;
  assign n270 = ~n264 & ~n269 ;
  assign n271 = ~wb_rst_i_pad & ~n270 ;
  assign n272 = \byte_controller_bit_controller_c_state_reg[6]/NET0131  & ~\byte_controller_bit_controller_clk_en_reg/NET0131  ;
  assign n273 = n151 & n156 ;
  assign n274 = n208 & n273 ;
  assign n275 = ~n272 & ~n274 ;
  assign n276 = n139 & ~n275 ;
  assign n277 = \byte_controller_bit_controller_c_state_reg[7]/NET0131  & ~\byte_controller_bit_controller_clk_en_reg/NET0131  ;
  assign n278 = n185 & n209 ;
  assign n279 = ~n277 & ~n278 ;
  assign n280 = n139 & ~n279 ;
  assign n281 = \byte_controller_bit_controller_c_state_reg[0]/NET0131  & ~\byte_controller_bit_controller_clk_en_reg/NET0131  ;
  assign n282 = \byte_controller_bit_controller_clk_en_reg/NET0131  & \byte_controller_c_state_reg[0]/NET0131  ;
  assign n283 = ~\byte_controller_core_cmd_reg[3]/NET0131  & n282 ;
  assign n284 = n227 & n283 ;
  assign n285 = n204 & n284 ;
  assign n286 = ~n281 & ~n285 ;
  assign n287 = n139 & ~n286 ;
  assign n288 = ~\byte_controller_bit_controller_clk_en_reg/NET0131  & n139 ;
  assign n289 = \byte_controller_bit_controller_c_state_reg[12]/NET0131  & n288 ;
  assign n290 = \byte_controller_bit_controller_clk_en_reg/NET0131  & n139 ;
  assign n291 = n157 & n290 ;
  assign n292 = ~\byte_controller_bit_controller_c_state_reg[9]/NET0131  & n141 ;
  assign n293 = n170 & n292 ;
  assign n294 = n291 & n293 ;
  assign n295 = n143 & n180 ;
  assign n296 = n294 & n295 ;
  assign n297 = ~n204 & n296 ;
  assign n298 = ~n289 & ~n297 ;
  assign n299 = \byte_controller_bit_controller_c_state_reg[15]/NET0131  & n288 ;
  assign n300 = ~\byte_controller_bit_controller_c_state_reg[16]/NET0131  & n144 ;
  assign n301 = ~\byte_controller_bit_controller_c_state_reg[15]/NET0131  & n300 ;
  assign n302 = n294 & n301 ;
  assign n303 = ~n204 & n302 ;
  assign n304 = ~n299 & ~n303 ;
  assign n305 = \byte_controller_bit_controller_c_state_reg[16]/NET0131  & n288 ;
  assign n307 = ~n204 & n290 ;
  assign n308 = ~\byte_controller_bit_controller_c_state_reg[0]/NET0131  & n307 ;
  assign n306 = n172 & n175 ;
  assign n309 = ~\byte_controller_bit_controller_c_state_reg[14]/NET0131  & n300 ;
  assign n310 = n306 & n309 ;
  assign n311 = n308 & n310 ;
  assign n312 = ~n305 & ~n311 ;
  assign n313 = ~\byte_controller_bit_controller_sSDA_reg/NET0131  & \byte_controller_bit_controller_sda_chk_reg/NET0131  ;
  assign n314 = sda_padoen_o_pad & n313 ;
  assign n315 = ~\byte_controller_bit_controller_c_state_reg[1]/NET0131  & n173 ;
  assign n316 = n170 & n315 ;
  assign n317 = n213 & n316 ;
  assign n318 = n157 & n180 ;
  assign n319 = n317 & n318 ;
  assign n320 = ~\byte_controller_bit_controller_cmd_stop_reg/NET0131  & \byte_controller_bit_controller_sto_condition_reg/NET0131  ;
  assign n321 = ~n319 & n320 ;
  assign n322 = ~n314 & ~n321 ;
  assign n323 = ~wb_rst_i_pad & ~n322 ;
  assign n324 = \byte_controller_bit_controller_c_state_reg[14]/NET0131  & n288 ;
  assign n325 = n146 & n291 ;
  assign n326 = n317 & n325 ;
  assign n327 = ~n204 & n326 ;
  assign n328 = ~n324 & ~n327 ;
  assign n329 = \byte_controller_bit_controller_c_state_reg[10]/NET0131  & n288 ;
  assign n330 = n171 & n203 ;
  assign n331 = n307 & n330 ;
  assign n332 = ~n329 & ~n331 ;
  assign n333 = \byte_controller_bit_controller_c_state_reg[11]/NET0131  & n288 ;
  assign n334 = n146 & n174 ;
  assign n335 = n306 & n334 ;
  assign n336 = n307 & n335 ;
  assign n337 = ~n333 & ~n336 ;
  assign n338 = \byte_controller_bit_controller_c_state_reg[1]/NET0131  & n288 ;
  assign n339 = ~\byte_controller_bit_controller_c_state_reg[2]/NET0131  & ~\byte_controller_bit_controller_c_state_reg[3]/NET0131  ;
  assign n340 = n186 & n339 ;
  assign n341 = ~\byte_controller_bit_controller_c_state_reg[1]/NET0131  & n307 ;
  assign n342 = n340 & n341 ;
  assign n343 = ~n338 & ~n342 ;
  assign n344 = \byte_controller_bit_controller_c_state_reg[2]/NET0131  & n288 ;
  assign n345 = n308 & n340 ;
  assign n346 = ~n344 & ~n345 ;
  assign n347 = ~\byte_controller_bit_controller_cnt_reg[8]/NET0131  & n251 ;
  assign n348 = \byte_controller_bit_controller_cnt_reg[8]/NET0131  & ~n251 ;
  assign n349 = ~n347 & ~n348 ;
  assign n350 = n260 & ~n349 ;
  assign n351 = ~\prer_reg[8]/NET0131  & ~n265 ;
  assign n352 = ~\byte_controller_bit_controller_cnt_reg[8]/NET0131  & n265 ;
  assign n353 = ~n351 & ~n352 ;
  assign n354 = ~n260 & n353 ;
  assign n355 = ~n350 & ~n354 ;
  assign n356 = ~wb_rst_i_pad & ~n355 ;
  assign n357 = \byte_controller_bit_controller_cnt_reg[6]/NET0131  & ~n249 ;
  assign n358 = ~n261 & ~n357 ;
  assign n359 = n260 & ~n358 ;
  assign n360 = ~\prer_reg[6]/NET0131  & ~n265 ;
  assign n361 = ~\byte_controller_bit_controller_cnt_reg[6]/NET0131  & n265 ;
  assign n362 = ~n360 & ~n361 ;
  assign n363 = ~n260 & n362 ;
  assign n364 = ~n359 & ~n363 ;
  assign n365 = ~wb_rst_i_pad & ~n364 ;
  assign n369 = \byte_controller_bit_controller_cnt_reg[9]/NET0131  & n265 ;
  assign n370 = \prer_reg[9]/NET0131  & ~n265 ;
  assign n371 = ~n369 & ~n370 ;
  assign n372 = ~n260 & n371 ;
  assign n366 = \byte_controller_bit_controller_cnt_reg[9]/NET0131  & ~n347 ;
  assign n367 = ~n253 & ~n366 ;
  assign n368 = n260 & n367 ;
  assign n373 = ~wb_rst_i_pad & ~n368 ;
  assign n374 = ~n372 & n373 ;
  assign n378 = ~\byte_controller_c_state_reg[1]/NET0131  & ~\byte_controller_c_state_reg[2]/NET0131  ;
  assign n379 = ~\byte_controller_c_state_reg[3]/NET0131  & ~\byte_controller_c_state_reg[4]/NET0131  ;
  assign n398 = n378 & n379 ;
  assign n399 = \byte_controller_c_state_reg[0]/NET0131  & n398 ;
  assign n400 = \byte_controller_bit_controller_cmd_ack_reg/NET0131  & n399 ;
  assign n401 = ~\cr_reg[5]/NET0131  & n400 ;
  assign n402 = ~\byte_controller_bit_controller_cmd_ack_reg/NET0131  & \byte_controller_core_cmd_reg[2]/NET0131  ;
  assign n403 = ~n401 & ~n402 ;
  assign n380 = ~\byte_controller_c_state_reg[0]/NET0131  & n379 ;
  assign n384 = \byte_controller_c_state_reg[1]/NET0131  & ~\byte_controller_c_state_reg[2]/NET0131  ;
  assign n385 = n380 & n384 ;
  assign n404 = ~\byte_controller_c_state_reg[0]/NET0131  & ~\byte_controller_c_state_reg[1]/NET0131  ;
  assign n405 = ~\byte_controller_c_state_reg[2]/NET0131  & n404 ;
  assign n406 = ~\byte_controller_c_state_reg[3]/NET0131  & n405 ;
  assign n407 = \byte_controller_c_state_reg[4]/NET0131  & n406 ;
  assign n408 = ~n385 & ~n407 ;
  assign n394 = ~\byte_controller_c_state_reg[1]/NET0131  & \byte_controller_c_state_reg[2]/NET0131  ;
  assign n395 = n380 & n394 ;
  assign n409 = ~n395 & ~n399 ;
  assign n410 = \byte_controller_c_state_reg[3]/NET0131  & ~\byte_controller_c_state_reg[4]/NET0131  ;
  assign n411 = n405 & n410 ;
  assign n412 = n409 & ~n411 ;
  assign n413 = n408 & n412 ;
  assign n414 = ~n403 & ~n413 ;
  assign n375 = ~\cr_reg[4]/NET0131  & ~\cr_reg[5]/NET0131  ;
  assign n376 = ~\cr_reg[6]/NET0131  & n375 ;
  assign n377 = ~\byte_controller_cmd_ack_reg/NET0131  & ~n376 ;
  assign n381 = n378 & n380 ;
  assign n390 = n377 & n381 ;
  assign n391 = ~\cr_reg[7]/NET0131  & n390 ;
  assign n392 = \cr_reg[4]/NET0131  & ~\cr_reg[5]/NET0131  ;
  assign n393 = n391 & n392 ;
  assign n382 = ~n377 & n381 ;
  assign n383 = \byte_controller_core_cmd_reg[2]/NET0131  & n382 ;
  assign n386 = ~\byte_controller_dcnt_reg[0]/NET0131  & ~\byte_controller_dcnt_reg[1]/NET0131  ;
  assign n387 = ~\byte_controller_dcnt_reg[2]/NET0131  & n386 ;
  assign n388 = \byte_controller_bit_controller_cmd_ack_reg/NET0131  & n387 ;
  assign n389 = n385 & n388 ;
  assign n396 = \byte_controller_bit_controller_cmd_ack_reg/NET0131  & ~n387 ;
  assign n397 = n395 & n396 ;
  assign n415 = ~n389 & ~n397 ;
  assign n416 = ~n383 & n415 ;
  assign n417 = ~n393 & n416 ;
  assign n418 = ~n414 & n417 ;
  assign n419 = n139 & ~n418 ;
  assign n420 = ~\byte_controller_bit_controller_cmd_ack_reg/NET0131  & ~n413 ;
  assign n421 = ~n382 & ~n420 ;
  assign n422 = \byte_controller_core_cmd_reg[3]/NET0131  & ~n421 ;
  assign n424 = ~n391 & ~n400 ;
  assign n425 = \cr_reg[5]/NET0131  & ~n424 ;
  assign n423 = n388 & n395 ;
  assign n426 = n385 & n396 ;
  assign n427 = ~n423 & ~n426 ;
  assign n428 = ~n425 & n427 ;
  assign n429 = ~n422 & n428 ;
  assign n430 = n139 & ~n429 ;
  assign n432 = ~\byte_controller_shift_reg/NET0131  & ~\byte_controller_sr_reg[0]/NET0131  ;
  assign n433 = ~\byte_controller_bit_controller_dout_reg/P0001  & \byte_controller_shift_reg/NET0131  ;
  assign n434 = ~n432 & ~n433 ;
  assign n435 = ~\byte_controller_ld_reg/NET0131  & ~n434 ;
  assign n431 = \byte_controller_ld_reg/NET0131  & ~\txr_reg[0]/NET0131  ;
  assign n436 = ~wb_rst_i_pad & ~n431 ;
  assign n437 = ~n435 & n436 ;
  assign n439 = ~\byte_controller_shift_reg/NET0131  & ~\byte_controller_sr_reg[1]/NET0131  ;
  assign n440 = \byte_controller_shift_reg/NET0131  & ~\byte_controller_sr_reg[0]/NET0131  ;
  assign n441 = ~n439 & ~n440 ;
  assign n442 = ~\byte_controller_ld_reg/NET0131  & ~n441 ;
  assign n438 = \byte_controller_ld_reg/NET0131  & ~\txr_reg[1]/NET0131  ;
  assign n443 = ~wb_rst_i_pad & ~n438 ;
  assign n444 = ~n442 & n443 ;
  assign n445 = ~n260 & ~n265 ;
  assign n447 = ~\byte_controller_bit_controller_cnt_reg[15]/NET0131  & ~n445 ;
  assign n446 = ~\prer_reg[15]/NET0131  & n445 ;
  assign n448 = n255 & n256 ;
  assign n449 = ~\byte_controller_bit_controller_cnt_reg[14]/NET0131  & n448 ;
  assign n450 = n260 & n449 ;
  assign n451 = ~wb_rst_i_pad & ~n450 ;
  assign n452 = ~n446 & n451 ;
  assign n453 = ~n447 & n452 ;
  assign n455 = ~\byte_controller_shift_reg/NET0131  & ~\byte_controller_sr_reg[2]/NET0131  ;
  assign n456 = \byte_controller_shift_reg/NET0131  & ~\byte_controller_sr_reg[1]/NET0131  ;
  assign n457 = ~n455 & ~n456 ;
  assign n458 = ~\byte_controller_ld_reg/NET0131  & ~n457 ;
  assign n454 = \byte_controller_ld_reg/NET0131  & ~\txr_reg[2]/NET0131  ;
  assign n459 = ~wb_rst_i_pad & ~n454 ;
  assign n460 = ~n458 & n459 ;
  assign n462 = ~\byte_controller_shift_reg/NET0131  & ~\byte_controller_sr_reg[3]/NET0131  ;
  assign n463 = \byte_controller_shift_reg/NET0131  & ~\byte_controller_sr_reg[2]/NET0131  ;
  assign n464 = ~n462 & ~n463 ;
  assign n465 = ~\byte_controller_ld_reg/NET0131  & ~n464 ;
  assign n461 = \byte_controller_ld_reg/NET0131  & ~\txr_reg[3]/NET0131  ;
  assign n466 = ~wb_rst_i_pad & ~n461 ;
  assign n467 = ~n465 & n466 ;
  assign n469 = ~\byte_controller_shift_reg/NET0131  & ~\byte_controller_sr_reg[4]/NET0131  ;
  assign n470 = \byte_controller_shift_reg/NET0131  & ~\byte_controller_sr_reg[3]/NET0131  ;
  assign n471 = ~n469 & ~n470 ;
  assign n472 = ~\byte_controller_ld_reg/NET0131  & ~n471 ;
  assign n468 = \byte_controller_ld_reg/NET0131  & ~\txr_reg[4]/NET0131  ;
  assign n473 = ~wb_rst_i_pad & ~n468 ;
  assign n474 = ~n472 & n473 ;
  assign n475 = \byte_controller_bit_controller_cnt_reg[0]/NET0131  & \byte_controller_bit_controller_cnt_reg[1]/NET0131  ;
  assign n476 = ~n245 & ~n475 ;
  assign n477 = n260 & ~n476 ;
  assign n478 = ~\prer_reg[1]/NET0131  & ~n265 ;
  assign n479 = ~\byte_controller_bit_controller_cnt_reg[1]/NET0131  & n265 ;
  assign n480 = ~n478 & ~n479 ;
  assign n481 = ~n260 & n480 ;
  assign n482 = ~n477 & ~n481 ;
  assign n483 = ~wb_rst_i_pad & ~n482 ;
  assign n485 = ~\byte_controller_shift_reg/NET0131  & ~\byte_controller_sr_reg[5]/NET0131  ;
  assign n486 = \byte_controller_shift_reg/NET0131  & ~\byte_controller_sr_reg[4]/NET0131  ;
  assign n487 = ~n485 & ~n486 ;
  assign n488 = ~\byte_controller_ld_reg/NET0131  & ~n487 ;
  assign n484 = \byte_controller_ld_reg/NET0131  & ~\txr_reg[5]/NET0131  ;
  assign n489 = ~wb_rst_i_pad & ~n484 ;
  assign n490 = ~n488 & n489 ;
  assign n492 = ~\byte_controller_shift_reg/NET0131  & ~\byte_controller_sr_reg[6]/NET0131  ;
  assign n493 = \byte_controller_shift_reg/NET0131  & ~\byte_controller_sr_reg[5]/NET0131  ;
  assign n494 = ~n492 & ~n493 ;
  assign n495 = ~\byte_controller_ld_reg/NET0131  & ~n494 ;
  assign n491 = \byte_controller_ld_reg/NET0131  & ~\txr_reg[6]/NET0131  ;
  assign n496 = ~wb_rst_i_pad & ~n491 ;
  assign n497 = ~n495 & n496 ;
  assign n498 = ~\byte_controller_bit_controller_cnt_reg[2]/NET0131  & n245 ;
  assign n499 = \byte_controller_bit_controller_cnt_reg[2]/NET0131  & ~n245 ;
  assign n500 = ~n498 & ~n499 ;
  assign n501 = n260 & ~n500 ;
  assign n502 = ~\prer_reg[2]/NET0131  & ~n265 ;
  assign n503 = ~\byte_controller_bit_controller_cnt_reg[2]/NET0131  & n265 ;
  assign n504 = ~n502 & ~n503 ;
  assign n505 = ~n260 & n504 ;
  assign n506 = ~n501 & ~n505 ;
  assign n507 = ~wb_rst_i_pad & ~n506 ;
  assign n509 = ~\byte_controller_shift_reg/NET0131  & ~\byte_controller_sr_reg[7]/NET0131  ;
  assign n510 = \byte_controller_shift_reg/NET0131  & ~\byte_controller_sr_reg[6]/NET0131  ;
  assign n511 = ~n509 & ~n510 ;
  assign n512 = ~\byte_controller_ld_reg/NET0131  & ~n511 ;
  assign n508 = \byte_controller_ld_reg/NET0131  & ~\txr_reg[7]/NET0131  ;
  assign n513 = ~wb_rst_i_pad & ~n508 ;
  assign n514 = ~n512 & n513 ;
  assign n515 = \byte_controller_bit_controller_cnt_reg[3]/NET0131  & ~n498 ;
  assign n516 = ~n247 & ~n515 ;
  assign n517 = n260 & ~n516 ;
  assign n518 = ~\prer_reg[3]/NET0131  & ~n265 ;
  assign n519 = ~\byte_controller_bit_controller_cnt_reg[3]/NET0131  & n265 ;
  assign n520 = ~n518 & ~n519 ;
  assign n521 = ~n260 & n520 ;
  assign n522 = ~n517 & ~n521 ;
  assign n523 = ~wb_rst_i_pad & ~n522 ;
  assign n524 = ~\byte_controller_bit_controller_cnt_reg[4]/NET0131  & n247 ;
  assign n525 = \byte_controller_bit_controller_cnt_reg[5]/NET0131  & ~n524 ;
  assign n526 = ~n249 & ~n525 ;
  assign n527 = n260 & ~n526 ;
  assign n528 = ~\prer_reg[5]/NET0131  & ~n265 ;
  assign n529 = ~\byte_controller_bit_controller_cnt_reg[5]/NET0131  & n265 ;
  assign n530 = ~n528 & ~n529 ;
  assign n531 = ~n260 & n530 ;
  assign n532 = ~n527 & ~n531 ;
  assign n533 = ~wb_rst_i_pad & ~n532 ;
  assign n535 = n375 & n391 ;
  assign n534 = ~\byte_controller_bit_controller_cmd_ack_reg/NET0131  & n407 ;
  assign n536 = \byte_controller_bit_controller_cmd_ack_reg/NET0131  & \cr_reg[6]/NET0131  ;
  assign n537 = n411 & n536 ;
  assign n538 = ~n534 & ~n537 ;
  assign n539 = ~n535 & n538 ;
  assign n540 = n139 & ~n539 ;
  assign n541 = ~wb_rst_i_pad & ~n445 ;
  assign n542 = ~n388 & n395 ;
  assign n543 = ~n401 & ~n542 ;
  assign n544 = ~n393 & n543 ;
  assign n545 = n139 & ~n544 ;
  assign n546 = ~\byte_controller_dcnt_reg[0]/NET0131  & \byte_controller_shift_reg/NET0131  ;
  assign n548 = \byte_controller_dcnt_reg[1]/NET0131  & ~n546 ;
  assign n547 = ~\byte_controller_dcnt_reg[1]/NET0131  & n546 ;
  assign n549 = ~\byte_controller_ld_reg/NET0131  & ~n547 ;
  assign n550 = ~n548 & n549 ;
  assign n551 = ~wb_rst_i_pad & ~n550 ;
  assign n553 = ~\byte_controller_dcnt_reg[2]/NET0131  & n547 ;
  assign n552 = \byte_controller_dcnt_reg[2]/NET0131  & ~n547 ;
  assign n554 = ~\byte_controller_ld_reg/NET0131  & ~n552 ;
  assign n555 = ~n553 & n554 ;
  assign n556 = ~wb_rst_i_pad & ~n555 ;
  assign n557 = n385 & ~n388 ;
  assign n558 = ~n425 & ~n557 ;
  assign n559 = n139 & ~n558 ;
  assign n560 = \byte_controller_dcnt_reg[0]/NET0131  & ~\byte_controller_shift_reg/NET0131  ;
  assign n561 = ~\byte_controller_ld_reg/NET0131  & ~n546 ;
  assign n562 = ~n560 & n561 ;
  assign n563 = ~wb_rst_i_pad & ~n562 ;
  assign n564 = ~\wb_adr_i[1]_pad  & ~\wb_adr_i[2]_pad  ;
  assign n565 = ~\wb_adr_i[0]_pad  & n564 ;
  assign n566 = wb_cyc_i_pad & wb_stb_i_pad ;
  assign n567 = wb_we_i_pad & n566 ;
  assign n568 = n565 & n567 ;
  assign n569 = ~\prer_reg[0]/NET0131  & ~n568 ;
  assign n570 = ~\wb_dat_i[0]_pad  & n567 ;
  assign n571 = n565 & n570 ;
  assign n572 = ~n569 & ~n571 ;
  assign n573 = ~wb_rst_i_pad & ~n572 ;
  assign n574 = \wb_adr_i[0]_pad  & n564 ;
  assign n575 = n567 & n574 ;
  assign n576 = ~\prer_reg[10]/NET0131  & ~n575 ;
  assign n577 = ~\wb_dat_i[2]_pad  & n567 ;
  assign n578 = n574 & n577 ;
  assign n579 = ~n576 & ~n578 ;
  assign n580 = ~wb_rst_i_pad & ~n579 ;
  assign n581 = ~\prer_reg[11]/NET0131  & ~n575 ;
  assign n582 = ~\wb_dat_i[3]_pad  & n567 ;
  assign n583 = n574 & n582 ;
  assign n584 = ~n581 & ~n583 ;
  assign n585 = ~wb_rst_i_pad & ~n584 ;
  assign n586 = ~\prer_reg[12]/NET0131  & ~n575 ;
  assign n587 = ~\wb_dat_i[4]_pad  & n567 ;
  assign n588 = n574 & n587 ;
  assign n589 = ~n586 & ~n588 ;
  assign n590 = ~wb_rst_i_pad & ~n589 ;
  assign n591 = ~\prer_reg[13]/NET0131  & ~n575 ;
  assign n592 = ~\wb_dat_i[5]_pad  & n567 ;
  assign n593 = n574 & n592 ;
  assign n594 = ~n591 & ~n593 ;
  assign n595 = ~wb_rst_i_pad & ~n594 ;
  assign n596 = ~\prer_reg[14]/NET0131  & ~n575 ;
  assign n597 = ~\wb_dat_i[6]_pad  & n567 ;
  assign n598 = n574 & n597 ;
  assign n599 = ~n596 & ~n598 ;
  assign n600 = ~wb_rst_i_pad & ~n599 ;
  assign n601 = ~\prer_reg[15]/NET0131  & ~n575 ;
  assign n602 = ~\wb_dat_i[7]_pad  & n567 ;
  assign n603 = n574 & n602 ;
  assign n604 = ~n601 & ~n603 ;
  assign n605 = ~wb_rst_i_pad & ~n604 ;
  assign n606 = ~\prer_reg[1]/NET0131  & ~n568 ;
  assign n607 = ~\wb_dat_i[1]_pad  & n567 ;
  assign n608 = n565 & n607 ;
  assign n609 = ~n606 & ~n608 ;
  assign n610 = ~wb_rst_i_pad & ~n609 ;
  assign n611 = ~\prer_reg[2]/NET0131  & ~n568 ;
  assign n612 = n565 & n577 ;
  assign n613 = ~n611 & ~n612 ;
  assign n614 = ~wb_rst_i_pad & ~n613 ;
  assign n615 = ~\prer_reg[3]/NET0131  & ~n568 ;
  assign n616 = n565 & n582 ;
  assign n617 = ~n615 & ~n616 ;
  assign n618 = ~wb_rst_i_pad & ~n617 ;
  assign n619 = ~\prer_reg[4]/NET0131  & ~n568 ;
  assign n620 = n565 & n587 ;
  assign n621 = ~n619 & ~n620 ;
  assign n622 = ~wb_rst_i_pad & ~n621 ;
  assign n623 = ~\prer_reg[5]/NET0131  & ~n568 ;
  assign n624 = n565 & n592 ;
  assign n625 = ~n623 & ~n624 ;
  assign n626 = ~wb_rst_i_pad & ~n625 ;
  assign n627 = ~\prer_reg[6]/NET0131  & ~n568 ;
  assign n628 = n565 & n597 ;
  assign n629 = ~n627 & ~n628 ;
  assign n630 = ~wb_rst_i_pad & ~n629 ;
  assign n631 = ~\prer_reg[7]/NET0131  & ~n568 ;
  assign n632 = n565 & n602 ;
  assign n633 = ~n631 & ~n632 ;
  assign n634 = ~wb_rst_i_pad & ~n633 ;
  assign n635 = ~\prer_reg[8]/NET0131  & ~n575 ;
  assign n636 = n570 & n574 ;
  assign n637 = ~n635 & ~n636 ;
  assign n638 = ~wb_rst_i_pad & ~n637 ;
  assign n639 = ~\prer_reg[9]/NET0131  & ~n575 ;
  assign n640 = n574 & n607 ;
  assign n641 = ~n639 & ~n640 ;
  assign n642 = ~wb_rst_i_pad & ~n641 ;
  assign n643 = ~\byte_controller_ack_out_reg/NET0131  & ~\byte_controller_bit_controller_cmd_ack_reg/NET0131  ;
  assign n644 = \byte_controller_bit_controller_cmd_ack_reg/NET0131  & ~\byte_controller_bit_controller_dout_reg/P0001  ;
  assign n645 = ~n643 & ~n644 ;
  assign n646 = n411 & n645 ;
  assign n647 = ~n395 & ~n398 ;
  assign n648 = n408 & n647 ;
  assign n649 = \byte_controller_ack_out_reg/NET0131  & ~n648 ;
  assign n650 = ~n646 & ~n649 ;
  assign n651 = n139 & ~n650 ;
  assign n652 = ~n406 & n409 ;
  assign n653 = \byte_controller_sr_reg[7]/NET0131  & ~n652 ;
  assign n654 = ~\byte_controller_bit_controller_cmd_ack_reg/NET0131  & ~\cr_reg[3]/NET0131  ;
  assign n655 = n411 & ~n654 ;
  assign n656 = ~\byte_controller_bit_controller_cmd_ack_reg/NET0131  & ~\byte_controller_sr_reg[7]/NET0131  ;
  assign n657 = \byte_controller_bit_controller_cmd_ack_reg/NET0131  & ~\cr_reg[3]/NET0131  ;
  assign n658 = ~n656 & ~n657 ;
  assign n659 = n385 & n658 ;
  assign n660 = ~n655 & ~n659 ;
  assign n661 = ~n653 & n660 ;
  assign n662 = n139 & ~n661 ;
  assign n663 = ~\byte_controller_bit_controller_busy_reg/NET0131  & ~\byte_controller_bit_controller_sta_condition_reg/NET0131  ;
  assign n664 = ~\byte_controller_bit_controller_sto_condition_reg/NET0131  & ~wb_rst_i_pad ;
  assign n665 = ~n663 & n664 ;
  assign n666 = ~n395 & ~n411 ;
  assign n667 = ~\byte_controller_bit_controller_cmd_ack_reg/NET0131  & \byte_controller_c_state_reg[3]/NET0131  ;
  assign n668 = ~n666 & n667 ;
  assign n669 = ~n389 & ~n423 ;
  assign n670 = ~n668 & n669 ;
  assign n671 = n139 & ~n670 ;
  assign n672 = ~\byte_controller_bit_controller_cmd_ack_reg/NET0131  & n399 ;
  assign n673 = \cr_reg[7]/NET0131  & n390 ;
  assign n674 = ~n672 & ~n673 ;
  assign n675 = n139 & ~n674 ;
  assign n676 = \byte_controller_bit_controller_cmd_ack_reg/NET0131  & \byte_controller_c_state_reg[0]/NET0131  ;
  assign n677 = ~n390 & ~n676 ;
  assign n678 = n139 & ~n677 ;
  assign n679 = ~\wb_adr_i[1]_pad  & \wb_adr_i[2]_pad  ;
  assign n680 = ~\wb_adr_i[0]_pad  & n679 ;
  assign n681 = \ctr_reg[7]/NET0131  & n680 ;
  assign n682 = n567 & n681 ;
  assign n683 = ~\byte_controller_bit_controller_al_reg/NET0131  & ~\byte_controller_cmd_ack_reg/NET0131  ;
  assign n684 = ~n567 & ~n683 ;
  assign n685 = ~n682 & ~n684 ;
  assign n686 = \cr_reg[4]/NET0131  & n685 ;
  assign n687 = \wb_dat_i[4]_pad  & n682 ;
  assign n688 = ~n686 & ~n687 ;
  assign n689 = ~wb_rst_i_pad & ~n688 ;
  assign n690 = \cr_reg[5]/NET0131  & n685 ;
  assign n691 = \wb_dat_i[5]_pad  & n682 ;
  assign n692 = ~n690 & ~n691 ;
  assign n693 = ~wb_rst_i_pad & ~n692 ;
  assign n694 = \cr_reg[6]/NET0131  & n685 ;
  assign n695 = \wb_dat_i[6]_pad  & n682 ;
  assign n696 = ~n694 & ~n695 ;
  assign n697 = ~wb_rst_i_pad & ~n696 ;
  assign n698 = \cr_reg[7]/NET0131  & n685 ;
  assign n699 = \wb_dat_i[7]_pad  & n682 ;
  assign n700 = ~n698 & ~n699 ;
  assign n701 = ~wb_rst_i_pad & ~n700 ;
  assign n702 = \wb_adr_i[1]_pad  & ~\wb_adr_i[2]_pad  ;
  assign n703 = ~\wb_adr_i[0]_pad  & n702 ;
  assign n704 = n567 & n703 ;
  assign n706 = ~\wb_dat_i[1]_pad  & n704 ;
  assign n705 = ~\ctr_reg[1]/NET0131  & ~n704 ;
  assign n707 = ~wb_rst_i_pad & ~n705 ;
  assign n708 = ~n706 & n707 ;
  assign n710 = ~\wb_dat_i[2]_pad  & n704 ;
  assign n709 = ~\ctr_reg[2]/NET0131  & ~n704 ;
  assign n711 = ~wb_rst_i_pad & ~n709 ;
  assign n712 = ~n710 & n711 ;
  assign n714 = ~\wb_dat_i[3]_pad  & n704 ;
  assign n713 = ~\ctr_reg[3]/NET0131  & ~n704 ;
  assign n715 = ~wb_rst_i_pad & ~n713 ;
  assign n716 = ~n714 & n715 ;
  assign n718 = ~\wb_dat_i[4]_pad  & n704 ;
  assign n717 = ~\ctr_reg[4]/NET0131  & ~n704 ;
  assign n719 = ~wb_rst_i_pad & ~n717 ;
  assign n720 = ~n718 & n719 ;
  assign n722 = ~\wb_dat_i[5]_pad  & n704 ;
  assign n721 = ~\ctr_reg[5]/NET0131  & ~n704 ;
  assign n723 = ~wb_rst_i_pad & ~n721 ;
  assign n724 = ~n722 & n723 ;
  assign n726 = ~\wb_dat_i[6]_pad  & n704 ;
  assign n725 = ~\ctr_reg[6]/NET0131  & ~n704 ;
  assign n727 = ~wb_rst_i_pad & ~n725 ;
  assign n728 = ~n726 & n727 ;
  assign n730 = ~\wb_dat_i[7]_pad  & n704 ;
  assign n729 = ~\ctr_reg[7]/NET0131  & ~n704 ;
  assign n731 = ~wb_rst_i_pad & ~n729 ;
  assign n732 = ~n730 & n731 ;
  assign n733 = \wb_adr_i[0]_pad  & n702 ;
  assign n734 = n567 & n733 ;
  assign n736 = ~\wb_dat_i[0]_pad  & n734 ;
  assign n735 = ~\txr_reg[0]/NET0131  & ~n734 ;
  assign n737 = ~wb_rst_i_pad & ~n735 ;
  assign n738 = ~n736 & n737 ;
  assign n740 = ~\wb_dat_i[1]_pad  & n734 ;
  assign n739 = ~\txr_reg[1]/NET0131  & ~n734 ;
  assign n741 = ~wb_rst_i_pad & ~n739 ;
  assign n742 = ~n740 & n741 ;
  assign n744 = ~\wb_dat_i[2]_pad  & n734 ;
  assign n743 = ~\txr_reg[2]/NET0131  & ~n734 ;
  assign n745 = ~wb_rst_i_pad & ~n743 ;
  assign n746 = ~n744 & n745 ;
  assign n748 = ~\wb_dat_i[3]_pad  & n734 ;
  assign n747 = ~\txr_reg[3]/NET0131  & ~n734 ;
  assign n749 = ~wb_rst_i_pad & ~n747 ;
  assign n750 = ~n748 & n749 ;
  assign n752 = ~\wb_dat_i[4]_pad  & n734 ;
  assign n751 = ~\txr_reg[4]/NET0131  & ~n734 ;
  assign n753 = ~wb_rst_i_pad & ~n751 ;
  assign n754 = ~n752 & n753 ;
  assign n756 = ~\wb_dat_i[5]_pad  & n734 ;
  assign n755 = ~\txr_reg[5]/NET0131  & ~n734 ;
  assign n757 = ~wb_rst_i_pad & ~n755 ;
  assign n758 = ~n756 & n757 ;
  assign n760 = ~\wb_dat_i[6]_pad  & n734 ;
  assign n759 = ~\txr_reg[6]/NET0131  & ~n734 ;
  assign n761 = ~wb_rst_i_pad & ~n759 ;
  assign n762 = ~n760 & n761 ;
  assign n764 = ~\wb_dat_i[7]_pad  & n734 ;
  assign n763 = ~\txr_reg[7]/NET0131  & ~n734 ;
  assign n765 = ~wb_rst_i_pad & ~n763 ;
  assign n766 = ~n764 & n765 ;
  assign n776 = \prer_reg[8]/NET0131  & n574 ;
  assign n774 = \ctr_reg[0]/NET0131  & n703 ;
  assign n775 = \prer_reg[0]/NET0131  & n565 ;
  assign n779 = ~n774 & ~n775 ;
  assign n780 = ~n776 & n779 ;
  assign n767 = \irq_flag_reg/NET0131  & n680 ;
  assign n768 = \byte_controller_sr_reg[0]/NET0131  & n733 ;
  assign n777 = ~n767 & ~n768 ;
  assign n769 = \wb_adr_i[0]_pad  & n679 ;
  assign n770 = \txr_reg[0]/NET0131  & n769 ;
  assign n771 = ~\wb_adr_i[0]_pad  & \wb_adr_i[1]_pad  ;
  assign n772 = \wb_adr_i[2]_pad  & n771 ;
  assign n773 = \cr_reg[0]/NET0131  & n772 ;
  assign n778 = ~n770 & ~n773 ;
  assign n781 = n777 & n778 ;
  assign n782 = n780 & n781 ;
  assign n783 = \prer_reg[10]/NET0131  & n574 ;
  assign n784 = \byte_controller_sr_reg[2]/NET0131  & n733 ;
  assign n789 = ~n783 & ~n784 ;
  assign n785 = \prer_reg[2]/NET0131  & n565 ;
  assign n786 = \cr_reg[2]/NET0131  & n772 ;
  assign n790 = ~n785 & ~n786 ;
  assign n787 = \ctr_reg[2]/NET0131  & n703 ;
  assign n788 = \txr_reg[2]/NET0131  & n769 ;
  assign n791 = ~n787 & ~n788 ;
  assign n792 = n790 & n791 ;
  assign n793 = n789 & n792 ;
  assign n794 = \prer_reg[11]/NET0131  & n574 ;
  assign n795 = \byte_controller_sr_reg[3]/NET0131  & n733 ;
  assign n800 = ~n794 & ~n795 ;
  assign n796 = \prer_reg[3]/NET0131  & n565 ;
  assign n797 = \cr_reg[3]/NET0131  & n772 ;
  assign n801 = ~n796 & ~n797 ;
  assign n798 = \ctr_reg[3]/NET0131  & n703 ;
  assign n799 = \txr_reg[3]/NET0131  & n769 ;
  assign n802 = ~n798 & ~n799 ;
  assign n803 = n801 & n802 ;
  assign n804 = n800 & n803 ;
  assign n805 = \prer_reg[12]/NET0131  & n574 ;
  assign n806 = \byte_controller_sr_reg[4]/NET0131  & n733 ;
  assign n811 = ~n805 & ~n806 ;
  assign n807 = \prer_reg[4]/NET0131  & n565 ;
  assign n808 = \cr_reg[4]/NET0131  & n772 ;
  assign n812 = ~n807 & ~n808 ;
  assign n809 = \ctr_reg[4]/NET0131  & n703 ;
  assign n810 = \txr_reg[4]/NET0131  & n769 ;
  assign n813 = ~n809 & ~n810 ;
  assign n814 = n812 & n813 ;
  assign n815 = n811 & n814 ;
  assign n817 = ~\wb_dat_i[3]_pad  & n682 ;
  assign n816 = ~\cr_reg[3]/NET0131  & ~n682 ;
  assign n818 = ~wb_rst_i_pad & ~n816 ;
  assign n819 = ~n817 & n818 ;
  assign n821 = ~\wb_dat_i[0]_pad  & n704 ;
  assign n820 = ~\ctr_reg[0]/NET0131  & ~n704 ;
  assign n822 = ~wb_rst_i_pad & ~n820 ;
  assign n823 = ~n821 & n822 ;
  assign n830 = \tip_reg/NET0131  & n680 ;
  assign n828 = \cr_reg[1]/NET0131  & n772 ;
  assign n829 = \prer_reg[9]/NET0131  & n574 ;
  assign n833 = ~n828 & ~n829 ;
  assign n834 = ~n830 & n833 ;
  assign n824 = \ctr_reg[1]/NET0131  & n703 ;
  assign n825 = \prer_reg[1]/NET0131  & n565 ;
  assign n831 = ~n824 & ~n825 ;
  assign n826 = \txr_reg[1]/NET0131  & n769 ;
  assign n827 = \byte_controller_sr_reg[1]/NET0131  & n733 ;
  assign n832 = ~n826 & ~n827 ;
  assign n835 = n831 & n832 ;
  assign n836 = n834 & n835 ;
  assign n843 = \txr_reg[5]/NET0131  & n769 ;
  assign n841 = \cr_reg[5]/NET0131  & n772 ;
  assign n842 = \byte_controller_sr_reg[5]/NET0131  & n733 ;
  assign n846 = ~n841 & ~n842 ;
  assign n847 = ~n843 & n846 ;
  assign n837 = \al_reg/NET0131  & n680 ;
  assign n838 = \prer_reg[5]/NET0131  & n565 ;
  assign n844 = ~n837 & ~n838 ;
  assign n839 = \prer_reg[13]/NET0131  & n574 ;
  assign n840 = \ctr_reg[5]/NET0131  & n703 ;
  assign n845 = ~n839 & ~n840 ;
  assign n848 = n844 & n845 ;
  assign n849 = n847 & n848 ;
  assign n856 = \txr_reg[6]/NET0131  & n769 ;
  assign n854 = \cr_reg[6]/NET0131  & n772 ;
  assign n855 = \byte_controller_sr_reg[6]/NET0131  & n733 ;
  assign n859 = ~n854 & ~n855 ;
  assign n860 = ~n856 & n859 ;
  assign n850 = \byte_controller_bit_controller_busy_reg/NET0131  & n680 ;
  assign n851 = \ctr_reg[6]/NET0131  & n703 ;
  assign n857 = ~n850 & ~n851 ;
  assign n852 = \prer_reg[6]/NET0131  & n565 ;
  assign n853 = \prer_reg[14]/NET0131  & n574 ;
  assign n858 = ~n852 & ~n853 ;
  assign n861 = n857 & n858 ;
  assign n862 = n860 & n861 ;
  assign n869 = \rxack_reg/NET0131  & n680 ;
  assign n867 = \cr_reg[7]/NET0131  & n772 ;
  assign n868 = \prer_reg[15]/NET0131  & n574 ;
  assign n872 = ~n867 & ~n868 ;
  assign n873 = ~n869 & n872 ;
  assign n863 = \ctr_reg[7]/NET0131  & n703 ;
  assign n864 = \prer_reg[7]/NET0131  & n565 ;
  assign n870 = ~n863 & ~n864 ;
  assign n865 = \txr_reg[7]/NET0131  & n769 ;
  assign n866 = \byte_controller_sr_reg[7]/NET0131  & n733 ;
  assign n871 = ~n865 & ~n866 ;
  assign n874 = n870 & n871 ;
  assign n875 = n873 & n874 ;
  assign n876 = \byte_controller_bit_controller_cmd_ack_reg/NET0131  & n139 ;
  assign n877 = ~n387 & n394 ;
  assign n878 = ~n384 & ~n877 ;
  assign n879 = n876 & ~n878 ;
  assign n880 = ~\byte_controller_bit_controller_sSDA_reg/NET0131  & ~wb_rst_i_pad ;
  assign n881 = \byte_controller_bit_controller_dSDA_reg/NET0131  & \byte_controller_bit_controller_sSCL_reg/NET0131  ;
  assign n882 = n880 & n881 ;
  assign n883 = ~\byte_controller_bit_controller_dSDA_reg/NET0131  & \byte_controller_bit_controller_sSCL_reg/NET0131  ;
  assign n884 = \byte_controller_bit_controller_sSDA_reg/NET0131  & ~wb_rst_i_pad ;
  assign n885 = n883 & n884 ;
  assign n886 = ~\byte_controller_bit_controller_clk_en_reg/NET0131  & \byte_controller_bit_controller_cmd_stop_reg/NET0131  ;
  assign n887 = ~n240 & ~n886 ;
  assign n888 = ~wb_rst_i_pad & ~n887 ;
  assign n891 = ~\wb_dat_i[0]_pad  & n681 ;
  assign n889 = ~wb_rst_i_pad & n567 ;
  assign n890 = ~\cr_reg[0]/NET0131  & ~n681 ;
  assign n892 = n889 & ~n890 ;
  assign n893 = ~n891 & n892 ;
  assign n895 = ~\wb_dat_i[1]_pad  & n681 ;
  assign n894 = ~\cr_reg[1]/NET0131  & ~n681 ;
  assign n896 = n889 & ~n894 ;
  assign n897 = ~n895 & n896 ;
  assign n899 = ~\wb_dat_i[2]_pad  & n681 ;
  assign n898 = ~\cr_reg[2]/NET0131  & ~n681 ;
  assign n900 = n889 & ~n898 ;
  assign n901 = ~n899 & n900 ;
  assign n902 = ~\byte_controller_c_state_reg[4]/NET0131  & ~\cr_reg[6]/NET0131  ;
  assign n903 = \byte_controller_c_state_reg[3]/NET0131  & ~n902 ;
  assign n904 = ~n379 & n876 ;
  assign n905 = ~n903 & n904 ;
  assign n906 = \byte_controller_bit_controller_sda_chk_reg/NET0131  & n288 ;
  assign n907 = ~n145 & n290 ;
  assign n908 = ~n906 & ~n907 ;
  assign n909 = \al_reg/NET0131  & ~\cr_reg[7]/NET0131  ;
  assign n910 = ~\byte_controller_bit_controller_al_reg/NET0131  & ~n909 ;
  assign n911 = ~wb_rst_i_pad & ~n910 ;
  assign n912 = ~\byte_controller_bit_controller_sSCL_reg/NET0131  & ~wb_rst_i_pad ;
  assign n913 = ~\byte_controller_bit_controller_c_state_reg[12]/NET0131  & ~\byte_controller_bit_controller_c_state_reg[16]/NET0131  ;
  assign n914 = ~\byte_controller_bit_controller_c_state_reg[4]/NET0131  & ~\byte_controller_bit_controller_c_state_reg[8]/NET0131  ;
  assign n915 = n913 & n914 ;
  assign n916 = n290 & ~n915 ;
  assign n917 = ~\irq_flag_reg/NET0131  & n683 ;
  assign n918 = ~\cr_reg[0]/NET0131  & ~wb_rst_i_pad ;
  assign n919 = ~n917 & n918 ;
  assign n920 = ~wb_rst_i_pad & ~n375 ;
  assign n921 = \ctr_reg[6]/NET0131  & \irq_flag_reg/NET0131  ;
  assign n922 = ~wb_rst_i_pad & n921 ;
  assign n923 = ~wb_ack_o_pad & wb_cyc_i_pad ;
  assign n924 = wb_stb_i_pad & n923 ;
  assign n925 = \byte_controller_ack_out_reg/NET0131  & ~wb_rst_i_pad ;
  assign n926 = ~scl_pad_i_pad & ~wb_rst_i_pad ;
  assign n927 = ~sda_pad_i_pad & ~wb_rst_i_pad ;
  assign n928 = \byte_controller_bit_controller_c_state_reg[8]/NET0131  & ~\byte_controller_bit_controller_clk_en_reg/NET0131  ;
  assign n929 = n156 & n159 ;
  assign n930 = n149 & n929 ;
  assign n931 = n208 & n930 ;
  assign n932 = ~n928 & ~n931 ;
  assign n933 = n139 & ~n932 ;
  assign n934 = \byte_controller_bit_controller_cnt_reg[14]/NET0131  & ~n448 ;
  assign n935 = ~n449 & ~n934 ;
  assign n936 = n260 & ~n935 ;
  assign n937 = ~\prer_reg[14]/NET0131  & ~n265 ;
  assign n938 = ~\byte_controller_bit_controller_cnt_reg[14]/NET0131  & n265 ;
  assign n939 = ~n937 & ~n938 ;
  assign n940 = ~n260 & n939 ;
  assign n941 = ~n936 & ~n940 ;
  assign n942 = ~wb_rst_i_pad & ~n941 ;
  assign n943 = ~\byte_controller_bit_controller_cnt_reg[10]/NET0131  & n253 ;
  assign n944 = \byte_controller_bit_controller_cnt_reg[10]/NET0131  & ~n253 ;
  assign n945 = ~n943 & ~n944 ;
  assign n946 = n260 & ~n945 ;
  assign n947 = ~\prer_reg[10]/NET0131  & ~n265 ;
  assign n948 = ~\byte_controller_bit_controller_cnt_reg[10]/NET0131  & n265 ;
  assign n949 = ~n947 & ~n948 ;
  assign n950 = ~n260 & n949 ;
  assign n951 = ~n946 & ~n950 ;
  assign n952 = ~wb_rst_i_pad & ~n951 ;
  assign n953 = \byte_controller_bit_controller_c_state_reg[4]/NET0131  & ~\byte_controller_bit_controller_clk_en_reg/NET0131  ;
  assign n954 = n186 & n208 ;
  assign n955 = ~n953 & ~n954 ;
  assign n956 = n139 & ~n955 ;
  assign n957 = ~\byte_controller_bit_controller_cnt_reg[12]/NET0131  & n255 ;
  assign n958 = \byte_controller_bit_controller_cnt_reg[12]/NET0131  & ~n255 ;
  assign n959 = ~n957 & ~n958 ;
  assign n960 = n260 & ~n959 ;
  assign n961 = ~\prer_reg[12]/NET0131  & ~n265 ;
  assign n962 = ~\byte_controller_bit_controller_cnt_reg[12]/NET0131  & n265 ;
  assign n963 = ~n961 & ~n962 ;
  assign n964 = ~n260 & n963 ;
  assign n965 = ~n960 & ~n964 ;
  assign n966 = ~wb_rst_i_pad & ~n965 ;
  assign n967 = \byte_controller_bit_controller_c_state_reg[13]/NET0131  & ~\byte_controller_bit_controller_clk_en_reg/NET0131  ;
  assign n968 = ~\byte_controller_c_state_reg[4]/NET0131  & \byte_controller_core_cmd_reg[2]/NET0131  ;
  assign n969 = n238 & n968 ;
  assign n970 = n204 & n969 ;
  assign n971 = ~n967 & ~n970 ;
  assign n972 = n139 & ~n971 ;
  assign n977 = \byte_controller_bit_controller_cnt_reg[0]/NET0131  & n260 ;
  assign n973 = \prer_reg[0]/NET0131  & ~n265 ;
  assign n974 = \byte_controller_bit_controller_cnt_reg[0]/NET0131  & n265 ;
  assign n975 = ~n973 & ~n974 ;
  assign n976 = ~n260 & n975 ;
  assign n978 = ~wb_rst_i_pad & ~n976 ;
  assign n979 = ~n977 & n978 ;
  assign n980 = \byte_controller_bit_controller_cnt_reg[13]/NET0131  & ~n957 ;
  assign n981 = ~n448 & ~n980 ;
  assign n982 = n260 & ~n981 ;
  assign n983 = ~\prer_reg[13]/NET0131  & ~n265 ;
  assign n984 = ~\byte_controller_bit_controller_cnt_reg[13]/NET0131  & n265 ;
  assign n985 = ~n983 & ~n984 ;
  assign n986 = ~n260 & n985 ;
  assign n987 = ~n982 & ~n986 ;
  assign n988 = ~wb_rst_i_pad & ~n987 ;
  assign n989 = \byte_controller_bit_controller_cnt_reg[4]/NET0131  & ~n247 ;
  assign n990 = ~n524 & ~n989 ;
  assign n991 = n260 & ~n990 ;
  assign n992 = ~\prer_reg[4]/NET0131  & ~n265 ;
  assign n993 = ~\byte_controller_bit_controller_cnt_reg[4]/NET0131  & n265 ;
  assign n994 = ~n992 & ~n993 ;
  assign n995 = ~n260 & n994 ;
  assign n996 = ~n991 & ~n995 ;
  assign n997 = ~wb_rst_i_pad & ~n996 ;
  assign n998 = \byte_controller_bit_controller_cnt_reg[11]/NET0131  & ~n943 ;
  assign n999 = ~n255 & ~n998 ;
  assign n1000 = n260 & ~n999 ;
  assign n1001 = ~\prer_reg[11]/NET0131  & ~n265 ;
  assign n1002 = ~\byte_controller_bit_controller_cnt_reg[11]/NET0131  & n265 ;
  assign n1003 = ~n1001 & ~n1002 ;
  assign n1004 = ~n260 & n1003 ;
  assign n1005 = ~n1000 & ~n1004 ;
  assign n1006 = ~wb_rst_i_pad & ~n1005 ;
  assign \_al_n1  = ~1'b0 ;
  assign \byte_controller_bit_controller_dout_reg/P0001_reg_syn_3  = ~n138 ;
  assign \g3074/_0_  = ~n202 ;
  assign \g3075/_0_  = ~n225 ;
  assign \g3102/_0_  = n233 ;
  assign \g3106/_0_  = n237 ;
  assign \g3117/_0_  = n244 ;
  assign \g3120/_0_  = n271 ;
  assign \g3127/_0_  = n276 ;
  assign \g3128/_0_  = n280 ;
  assign \g3129/_0_  = n287 ;
  assign \g3130/_0_  = ~n298 ;
  assign \g3131/_0_  = ~n304 ;
  assign \g3132/_0_  = ~n312 ;
  assign \g3160/_0_  = n323 ;
  assign \g3164/_0_  = ~n328 ;
  assign \g3166/_0_  = ~n332 ;
  assign \g3167/_0_  = ~n337 ;
  assign \g3171/_0_  = ~n343 ;
  assign \g3174/_3_  = ~n346 ;
  assign \g3184/_0_  = n356 ;
  assign \g3185/_0_  = n365 ;
  assign \g3188/_0_  = n374 ;
  assign \g3193/_0_  = n419 ;
  assign \g3195/_0_  = n430 ;
  assign \g3198/_0_  = n437 ;
  assign \g3199/_0_  = n444 ;
  assign \g32/_1_  = n453 ;
  assign \g3200/_0_  = n460 ;
  assign \g3201/_0_  = n467 ;
  assign \g3203/_0_  = n474 ;
  assign \g3204/_0_  = n483 ;
  assign \g3205/_0_  = n490 ;
  assign \g3206/_0_  = n497 ;
  assign \g3207/_0_  = n507 ;
  assign \g3208/_0_  = n514 ;
  assign \g3209/_0_  = n523 ;
  assign \g3211/_0_  = n533 ;
  assign \g3246/_0_  = n540 ;
  assign \g3250/_2_  = ~n541 ;
  assign \g3251/_0_  = n545 ;
  assign \g3255/_0_  = n551 ;
  assign \g3256/_0_  = n556 ;
  assign \g3259/_0_  = n559 ;
  assign \g3262/_0_  = n563 ;
  assign \g3269/_0_  = ~n573 ;
  assign \g3270/_0_  = ~n580 ;
  assign \g3271/_0_  = ~n585 ;
  assign \g3272/_0_  = ~n590 ;
  assign \g3273/_0_  = ~n595 ;
  assign \g3274/_0_  = ~n600 ;
  assign \g3275/_0_  = ~n605 ;
  assign \g3276/_0_  = ~n610 ;
  assign \g3277/_0_  = ~n614 ;
  assign \g3278/_0_  = ~n618 ;
  assign \g3279/_0_  = ~n622 ;
  assign \g3280/_0_  = ~n626 ;
  assign \g3281/_0_  = ~n630 ;
  assign \g3282/_0_  = ~n634 ;
  assign \g3283/_0_  = ~n638 ;
  assign \g3284/_0_  = ~n642 ;
  assign \g3285/_0_  = n651 ;
  assign \g3286/_0_  = n662 ;
  assign \g3307/_0_  = n665 ;
  assign \g3339/_0_  = n671 ;
  assign \g3392/_0_  = n675 ;
  assign \g3419/_0_  = n678 ;
  assign \g3421/_0_  = n689 ;
  assign \g3422/_0_  = n693 ;
  assign \g3423/_0_  = n697 ;
  assign \g3424/_0_  = n701 ;
  assign \g3425/_0_  = n708 ;
  assign \g3426/_0_  = n712 ;
  assign \g3427/_0_  = n716 ;
  assign \g3428/_0_  = n720 ;
  assign \g3429/_0_  = n724 ;
  assign \g3430/_0_  = n728 ;
  assign \g3431/_0_  = n732 ;
  assign \g3452/_0_  = n738 ;
  assign \g3453/_0_  = n742 ;
  assign \g3454/_0_  = n746 ;
  assign \g3455/_0_  = n750 ;
  assign \g3456/_0_  = n754 ;
  assign \g3457/_0_  = n758 ;
  assign \g3458/_0_  = n762 ;
  assign \g3459/_0_  = n766 ;
  assign \g3460/_0_  = ~n782 ;
  assign \g3462/_0_  = ~n793 ;
  assign \g3464/_0_  = ~n804 ;
  assign \g3465/_0_  = ~n815 ;
  assign \g3471/_0_  = n819 ;
  assign \g3472/_0_  = n823 ;
  assign \g3476/_0_  = ~n836 ;
  assign \g3477/_0_  = ~n849 ;
  assign \g3478/_0_  = ~n862 ;
  assign \g3479/_0_  = ~n875 ;
  assign \g3499/_0_  = n879 ;
  assign \g3506/_0_  = n882 ;
  assign \g3507/_0_  = n885 ;
  assign \g3591/_0_  = n888 ;
  assign \g3601/_0_  = n893 ;
  assign \g3602/_0_  = n897 ;
  assign \g3603/_0_  = n901 ;
  assign \g3693/_0_  = n905 ;
  assign \g3694/_0_  = ~n908 ;
  assign \g3761/_0_  = n911 ;
  assign \g3785/_0_  = ~n912 ;
  assign \g3798/_0_  = n916 ;
  assign \g3815/_1_  = ~n880 ;
  assign \g3840/_0_  = n919 ;
  assign \g3874/_0_  = n920 ;
  assign \g3915/_0_  = n922 ;
  assign \g3927/_2_  = n924 ;
  assign \g3978/_0_  = n925 ;
  assign \g4004/_0_  = ~n926 ;
  assign \g4021/_0_  = ~n927 ;
  assign \g4582/_0_  = n933 ;
  assign \g4804/_0_  = n942 ;
  assign \g4866/_0_  = n952 ;
  assign \g4876/_0_  = n956 ;
  assign \g4942/_0_  = n966 ;
  assign \g4996/_0_  = n972 ;
  assign \g5146/_0_  = n979 ;
  assign \g5236/_0_  = n988 ;
  assign \g5411/_0_  = n997 ;
  assign \g5433/_0_  = n1006 ;
  assign scl_pad_o_pad = 1'b0 ;
endmodule
