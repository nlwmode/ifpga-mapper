module top (\a0_pad , a_pad, b_pad, c_pad, \d0_pad , d_pad, e_pad, f_pad, g_pad, h_pad, j_pad, k_pad, l_pad, m_pad, n_pad, o_pad, p_pad, q_pad, s_pad, t_pad, u_pad, v_pad, w_pad, x_pad, y_pad, z_pad, \b0_pad , \c0_pad , \e0_pad , \f0_pad , \g0_pad , \h0_pad , \i0_pad , \j0_pad , \k0_pad , \l0_pad , \m0_pad , \n0_pad , \o0_pad , \p0_pad , \q0_pad , \r0_pad , \s0_pad , \t0_pad );
	input \a0_pad  ;
	input a_pad ;
	input b_pad ;
	input c_pad ;
	input \d0_pad  ;
	input d_pad ;
	input e_pad ;
	input f_pad ;
	input g_pad ;
	input h_pad ;
	input j_pad ;
	input k_pad ;
	input l_pad ;
	input m_pad ;
	input n_pad ;
	input o_pad ;
	input p_pad ;
	input q_pad ;
	input s_pad ;
	input t_pad ;
	input u_pad ;
	input v_pad ;
	input w_pad ;
	input x_pad ;
	input y_pad ;
	input z_pad ;
	output \b0_pad  ;
	output \c0_pad  ;
	output \e0_pad  ;
	output \f0_pad  ;
	output \g0_pad  ;
	output \h0_pad  ;
	output \i0_pad  ;
	output \j0_pad  ;
	output \k0_pad  ;
	output \l0_pad  ;
	output \m0_pad  ;
	output \n0_pad  ;
	output \o0_pad  ;
	output \p0_pad  ;
	output \q0_pad  ;
	output \r0_pad  ;
	output \s0_pad  ;
	output \t0_pad  ;
	wire _w97_ ;
	wire _w96_ ;
	wire _w95_ ;
	wire _w94_ ;
	wire _w93_ ;
	wire _w92_ ;
	wire _w91_ ;
	wire _w90_ ;
	wire _w89_ ;
	wire _w88_ ;
	wire _w87_ ;
	wire _w86_ ;
	wire _w55_ ;
	wire _w54_ ;
	wire _w53_ ;
	wire _w52_ ;
	wire _w51_ ;
	wire _w50_ ;
	wire _w49_ ;
	wire _w48_ ;
	wire _w47_ ;
	wire _w46_ ;
	wire _w45_ ;
	wire _w44_ ;
	wire _w43_ ;
	wire _w42_ ;
	wire _w41_ ;
	wire _w40_ ;
	wire _w27_ ;
	wire _w28_ ;
	wire _w29_ ;
	wire _w30_ ;
	wire _w31_ ;
	wire _w32_ ;
	wire _w33_ ;
	wire _w34_ ;
	wire _w35_ ;
	wire _w36_ ;
	wire _w37_ ;
	wire _w38_ ;
	wire _w39_ ;
	wire _w56_ ;
	wire _w57_ ;
	wire _w58_ ;
	wire _w59_ ;
	wire _w60_ ;
	wire _w61_ ;
	wire _w62_ ;
	wire _w63_ ;
	wire _w64_ ;
	wire _w65_ ;
	wire _w66_ ;
	wire _w67_ ;
	wire _w68_ ;
	wire _w69_ ;
	wire _w70_ ;
	wire _w71_ ;
	wire _w72_ ;
	wire _w73_ ;
	wire _w74_ ;
	wire _w75_ ;
	wire _w76_ ;
	wire _w77_ ;
	wire _w78_ ;
	wire _w79_ ;
	wire _w80_ ;
	wire _w81_ ;
	wire _w82_ ;
	wire _w83_ ;
	wire _w84_ ;
	wire _w85_ ;
	LUT2 #(
		.INIT('h4)
	) name0 (
		\d0_pad ,
		j_pad,
		_w27_
	);
	LUT2 #(
		.INIT('h1)
	) name1 (
		s_pad,
		t_pad,
		_w28_
	);
	LUT2 #(
		.INIT('h4)
	) name2 (
		u_pad,
		_w28_,
		_w29_
	);
	LUT2 #(
		.INIT('h1)
	) name3 (
		v_pad,
		_w29_,
		_w30_
	);
	LUT2 #(
		.INIT('h8)
	) name4 (
		w_pad,
		x_pad,
		_w31_
	);
	LUT2 #(
		.INIT('h4)
	) name5 (
		_w30_,
		_w31_,
		_w32_
	);
	LUT2 #(
		.INIT('h1)
	) name6 (
		y_pad,
		_w32_,
		_w33_
	);
	LUT2 #(
		.INIT('h4)
	) name7 (
		\a0_pad ,
		_w33_,
		_w34_
	);
	LUT2 #(
		.INIT('h8)
	) name8 (
		e_pad,
		f_pad,
		_w35_
	);
	LUT2 #(
		.INIT('h1)
	) name9 (
		\a0_pad ,
		z_pad,
		_w36_
	);
	LUT2 #(
		.INIT('h1)
	) name10 (
		h_pad,
		_w35_,
		_w37_
	);
	LUT2 #(
		.INIT('h4)
	) name11 (
		_w36_,
		_w37_,
		_w38_
	);
	LUT2 #(
		.INIT('h4)
	) name12 (
		_w34_,
		_w38_,
		_w39_
	);
	LUT2 #(
		.INIT('h2)
	) name13 (
		z_pad,
		_w33_,
		_w40_
	);
	LUT2 #(
		.INIT('h1)
	) name14 (
		\a0_pad ,
		_w40_,
		_w41_
	);
	LUT2 #(
		.INIT('h2)
	) name15 (
		b_pad,
		l_pad,
		_w42_
	);
	LUT2 #(
		.INIT('h4)
	) name16 (
		b_pad,
		l_pad,
		_w43_
	);
	LUT2 #(
		.INIT('h2)
	) name17 (
		c_pad,
		m_pad,
		_w44_
	);
	LUT2 #(
		.INIT('h4)
	) name18 (
		c_pad,
		m_pad,
		_w45_
	);
	LUT2 #(
		.INIT('h1)
	) name19 (
		d_pad,
		n_pad,
		_w46_
	);
	LUT2 #(
		.INIT('h8)
	) name20 (
		d_pad,
		n_pad,
		_w47_
	);
	LUT2 #(
		.INIT('h1)
	) name21 (
		_w46_,
		_w47_,
		_w48_
	);
	LUT2 #(
		.INIT('h2)
	) name22 (
		a_pad,
		k_pad,
		_w49_
	);
	LUT2 #(
		.INIT('h4)
	) name23 (
		a_pad,
		k_pad,
		_w50_
	);
	LUT2 #(
		.INIT('h1)
	) name24 (
		_w42_,
		_w43_,
		_w51_
	);
	LUT2 #(
		.INIT('h1)
	) name25 (
		_w44_,
		_w45_,
		_w52_
	);
	LUT2 #(
		.INIT('h1)
	) name26 (
		_w49_,
		_w50_,
		_w53_
	);
	LUT2 #(
		.INIT('h8)
	) name27 (
		_w52_,
		_w53_,
		_w54_
	);
	LUT2 #(
		.INIT('h4)
	) name28 (
		_w48_,
		_w51_,
		_w55_
	);
	LUT2 #(
		.INIT('h8)
	) name29 (
		_w54_,
		_w55_,
		_w56_
	);
	LUT2 #(
		.INIT('h1)
	) name30 (
		j_pad,
		_w56_,
		_w57_
	);
	LUT2 #(
		.INIT('h1)
	) name31 (
		j_pad,
		o_pad,
		_w58_
	);
	LUT2 #(
		.INIT('h4)
	) name32 (
		j_pad,
		p_pad,
		_w59_
	);
	LUT2 #(
		.INIT('h2)
	) name33 (
		g_pad,
		j_pad,
		_w60_
	);
	LUT2 #(
		.INIT('h1)
	) name34 (
		h_pad,
		q_pad,
		_w61_
	);
	LUT2 #(
		.INIT('h8)
	) name35 (
		_w35_,
		_w61_,
		_w62_
	);
	LUT2 #(
		.INIT('h4)
	) name36 (
		_w35_,
		_w61_,
		_w63_
	);
	LUT2 #(
		.INIT('h4)
	) name37 (
		s_pad,
		_w63_,
		_w64_
	);
	LUT2 #(
		.INIT('h8)
	) name38 (
		s_pad,
		t_pad,
		_w65_
	);
	LUT2 #(
		.INIT('h1)
	) name39 (
		_w28_,
		_w65_,
		_w66_
	);
	LUT2 #(
		.INIT('h8)
	) name40 (
		_w63_,
		_w66_,
		_w67_
	);
	LUT2 #(
		.INIT('h1)
	) name41 (
		u_pad,
		_w65_,
		_w68_
	);
	LUT2 #(
		.INIT('h8)
	) name42 (
		u_pad,
		_w65_,
		_w69_
	);
	LUT2 #(
		.INIT('h2)
	) name43 (
		_w63_,
		_w69_,
		_w70_
	);
	LUT2 #(
		.INIT('h4)
	) name44 (
		_w68_,
		_w70_,
		_w71_
	);
	LUT2 #(
		.INIT('h2)
	) name45 (
		u_pad,
		v_pad,
		_w72_
	);
	LUT2 #(
		.INIT('h8)
	) name46 (
		_w65_,
		_w72_,
		_w73_
	);
	LUT2 #(
		.INIT('h8)
	) name47 (
		v_pad,
		_w70_,
		_w74_
	);
	LUT2 #(
		.INIT('h2)
	) name48 (
		_w63_,
		_w73_,
		_w75_
	);
	LUT2 #(
		.INIT('h4)
	) name49 (
		_w74_,
		_w75_,
		_w76_
	);
	LUT2 #(
		.INIT('h2)
	) name50 (
		w_pad,
		_w73_,
		_w77_
	);
	LUT2 #(
		.INIT('h4)
	) name51 (
		w_pad,
		_w73_,
		_w78_
	);
	LUT2 #(
		.INIT('h2)
	) name52 (
		_w63_,
		_w77_,
		_w79_
	);
	LUT2 #(
		.INIT('h4)
	) name53 (
		_w78_,
		_w79_,
		_w80_
	);
	LUT2 #(
		.INIT('h1)
	) name54 (
		w_pad,
		x_pad,
		_w81_
	);
	LUT2 #(
		.INIT('h8)
	) name55 (
		_w73_,
		_w81_,
		_w82_
	);
	LUT2 #(
		.INIT('h2)
	) name56 (
		x_pad,
		_w78_,
		_w83_
	);
	LUT2 #(
		.INIT('h2)
	) name57 (
		_w63_,
		_w82_,
		_w84_
	);
	LUT2 #(
		.INIT('h4)
	) name58 (
		_w83_,
		_w84_,
		_w85_
	);
	LUT2 #(
		.INIT('h2)
	) name59 (
		y_pad,
		_w82_,
		_w86_
	);
	LUT2 #(
		.INIT('h4)
	) name60 (
		y_pad,
		_w82_,
		_w87_
	);
	LUT2 #(
		.INIT('h2)
	) name61 (
		_w63_,
		_w86_,
		_w88_
	);
	LUT2 #(
		.INIT('h4)
	) name62 (
		_w87_,
		_w88_,
		_w89_
	);
	LUT2 #(
		.INIT('h2)
	) name63 (
		z_pad,
		_w87_,
		_w90_
	);
	LUT2 #(
		.INIT('h4)
	) name64 (
		z_pad,
		_w87_,
		_w91_
	);
	LUT2 #(
		.INIT('h2)
	) name65 (
		_w63_,
		_w90_,
		_w92_
	);
	LUT2 #(
		.INIT('h4)
	) name66 (
		_w91_,
		_w92_,
		_w93_
	);
	LUT2 #(
		.INIT('h2)
	) name67 (
		\a0_pad ,
		_w91_,
		_w94_
	);
	LUT2 #(
		.INIT('h8)
	) name68 (
		_w36_,
		_w87_,
		_w95_
	);
	LUT2 #(
		.INIT('h2)
	) name69 (
		_w63_,
		_w95_,
		_w96_
	);
	LUT2 #(
		.INIT('h4)
	) name70 (
		_w94_,
		_w96_,
		_w97_
	);
	assign \b0_pad  = _w27_ ;
	assign \c0_pad  = _w39_ ;
	assign \e0_pad  = _w41_ ;
	assign \f0_pad  = _w57_ ;
	assign \g0_pad  = _w58_ ;
	assign \h0_pad  = _w59_ ;
	assign \i0_pad  = _w60_ ;
	assign \j0_pad  = _w41_ ;
	assign \k0_pad  = _w62_ ;
	assign \l0_pad  = _w64_ ;
	assign \m0_pad  = _w67_ ;
	assign \n0_pad  = _w71_ ;
	assign \o0_pad  = _w76_ ;
	assign \p0_pad  = _w80_ ;
	assign \q0_pad  = _w85_ ;
	assign \r0_pad  = _w89_ ;
	assign \s0_pad  = _w93_ ;
	assign \t0_pad  = _w97_ ;
endmodule;