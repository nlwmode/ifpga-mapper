module top (\a0_pad , a_pad, \b0_pad , b_pad, \c0_pad , c_pad, \d0_pad , d_pad, \e0_pad , e_pad, \f0_pad , f_pad, \g0_pad , g_pad, \h0_pad , h_pad, \i0_pad , i_pad, \j0_pad , j_pad, \k0_pad , k_pad, l_pad, m_pad, n_pad, o_pad, p_pad, q_pad, s_pad, t_pad, u_pad, v_pad, w_pad, x_pad, y_pad, z_pad, \a1_pad , \l0_pad , \m0_pad , \n0_pad , \o0_pad , \p0_pad , \q0_pad , \r0_pad , \s0_pad , \t0_pad , \u0_pad , \v0_pad , \w0_pad , \x0_pad , \y0_pad , \z0_pad );
	input \a0_pad  ;
	input a_pad ;
	input \b0_pad  ;
	input b_pad ;
	input \c0_pad  ;
	input c_pad ;
	input \d0_pad  ;
	input d_pad ;
	input \e0_pad  ;
	input e_pad ;
	input \f0_pad  ;
	input f_pad ;
	input \g0_pad  ;
	input g_pad ;
	input \h0_pad  ;
	input h_pad ;
	input \i0_pad  ;
	input i_pad ;
	input \j0_pad  ;
	input j_pad ;
	input \k0_pad  ;
	input k_pad ;
	input l_pad ;
	input m_pad ;
	input n_pad ;
	input o_pad ;
	input p_pad ;
	input q_pad ;
	input s_pad ;
	input t_pad ;
	input u_pad ;
	input v_pad ;
	input w_pad ;
	input x_pad ;
	input y_pad ;
	input z_pad ;
	output \a1_pad  ;
	output \l0_pad  ;
	output \m0_pad  ;
	output \n0_pad  ;
	output \o0_pad  ;
	output \p0_pad  ;
	output \q0_pad  ;
	output \r0_pad  ;
	output \s0_pad  ;
	output \t0_pad  ;
	output \u0_pad  ;
	output \v0_pad  ;
	output \w0_pad  ;
	output \x0_pad  ;
	output \y0_pad  ;
	output \z0_pad  ;
	wire _w101_ ;
	wire _w100_ ;
	wire _w99_ ;
	wire _w98_ ;
	wire _w97_ ;
	wire _w66_ ;
	wire _w65_ ;
	wire _w64_ ;
	wire _w63_ ;
	wire _w62_ ;
	wire _w61_ ;
	wire _w60_ ;
	wire _w59_ ;
	wire _w58_ ;
	wire _w57_ ;
	wire _w56_ ;
	wire _w55_ ;
	wire _w54_ ;
	wire _w53_ ;
	wire _w52_ ;
	wire _w51_ ;
	wire _w38_ ;
	wire _w39_ ;
	wire _w40_ ;
	wire _w41_ ;
	wire _w42_ ;
	wire _w43_ ;
	wire _w44_ ;
	wire _w45_ ;
	wire _w46_ ;
	wire _w47_ ;
	wire _w48_ ;
	wire _w49_ ;
	wire _w50_ ;
	wire _w67_ ;
	wire _w68_ ;
	wire _w69_ ;
	wire _w70_ ;
	wire _w71_ ;
	wire _w72_ ;
	wire _w73_ ;
	wire _w74_ ;
	wire _w75_ ;
	wire _w76_ ;
	wire _w77_ ;
	wire _w78_ ;
	wire _w79_ ;
	wire _w80_ ;
	wire _w81_ ;
	wire _w82_ ;
	wire _w83_ ;
	wire _w84_ ;
	wire _w85_ ;
	wire _w86_ ;
	wire _w87_ ;
	wire _w88_ ;
	wire _w89_ ;
	wire _w90_ ;
	wire _w91_ ;
	wire _w92_ ;
	wire _w93_ ;
	wire _w94_ ;
	wire _w95_ ;
	wire _w96_ ;
	LUT2 #(
		.INIT('h1)
	) name0 (
		\k0_pad ,
		u_pad,
		_w38_
	);
	LUT2 #(
		.INIT('h8)
	) name1 (
		\d0_pad ,
		t_pad,
		_w39_
	);
	LUT4 #(
		.INIT('h3200)
	) name2 (
		m_pad,
		s_pad,
		t_pad,
		u_pad,
		_w40_
	);
	LUT3 #(
		.INIT('hba)
	) name3 (
		_w38_,
		_w39_,
		_w40_,
		_w41_
	);
	LUT2 #(
		.INIT('h1)
	) name4 (
		u_pad,
		v_pad,
		_w42_
	);
	LUT2 #(
		.INIT('h8)
	) name5 (
		t_pad,
		w_pad,
		_w43_
	);
	LUT4 #(
		.INIT('h3200)
	) name6 (
		d_pad,
		s_pad,
		t_pad,
		u_pad,
		_w44_
	);
	LUT3 #(
		.INIT('hba)
	) name7 (
		_w42_,
		_w43_,
		_w44_,
		_w45_
	);
	LUT2 #(
		.INIT('h1)
	) name8 (
		u_pad,
		w_pad,
		_w46_
	);
	LUT2 #(
		.INIT('h8)
	) name9 (
		t_pad,
		x_pad,
		_w47_
	);
	LUT4 #(
		.INIT('h3200)
	) name10 (
		c_pad,
		s_pad,
		t_pad,
		u_pad,
		_w48_
	);
	LUT3 #(
		.INIT('hba)
	) name11 (
		_w46_,
		_w47_,
		_w48_,
		_w49_
	);
	LUT2 #(
		.INIT('h1)
	) name12 (
		u_pad,
		x_pad,
		_w50_
	);
	LUT2 #(
		.INIT('h8)
	) name13 (
		t_pad,
		y_pad,
		_w51_
	);
	LUT4 #(
		.INIT('h3200)
	) name14 (
		b_pad,
		s_pad,
		t_pad,
		u_pad,
		_w52_
	);
	LUT3 #(
		.INIT('hba)
	) name15 (
		_w50_,
		_w51_,
		_w52_,
		_w53_
	);
	LUT2 #(
		.INIT('h1)
	) name16 (
		u_pad,
		y_pad,
		_w54_
	);
	LUT2 #(
		.INIT('h4)
	) name17 (
		q_pad,
		t_pad,
		_w55_
	);
	LUT4 #(
		.INIT('h3200)
	) name18 (
		a_pad,
		s_pad,
		t_pad,
		u_pad,
		_w56_
	);
	LUT3 #(
		.INIT('hba)
	) name19 (
		_w54_,
		_w55_,
		_w56_,
		_w57_
	);
	LUT2 #(
		.INIT('h1)
	) name20 (
		u_pad,
		z_pad,
		_w58_
	);
	LUT2 #(
		.INIT('h8)
	) name21 (
		\a0_pad ,
		t_pad,
		_w59_
	);
	LUT4 #(
		.INIT('h3200)
	) name22 (
		h_pad,
		s_pad,
		t_pad,
		u_pad,
		_w60_
	);
	LUT3 #(
		.INIT('hba)
	) name23 (
		_w58_,
		_w59_,
		_w60_,
		_w61_
	);
	LUT2 #(
		.INIT('h1)
	) name24 (
		\a0_pad ,
		u_pad,
		_w62_
	);
	LUT2 #(
		.INIT('h8)
	) name25 (
		\b0_pad ,
		t_pad,
		_w63_
	);
	LUT4 #(
		.INIT('h3200)
	) name26 (
		g_pad,
		s_pad,
		t_pad,
		u_pad,
		_w64_
	);
	LUT3 #(
		.INIT('hba)
	) name27 (
		_w62_,
		_w63_,
		_w64_,
		_w65_
	);
	LUT2 #(
		.INIT('h1)
	) name28 (
		\b0_pad ,
		u_pad,
		_w66_
	);
	LUT2 #(
		.INIT('h8)
	) name29 (
		\c0_pad ,
		t_pad,
		_w67_
	);
	LUT4 #(
		.INIT('h3200)
	) name30 (
		f_pad,
		s_pad,
		t_pad,
		u_pad,
		_w68_
	);
	LUT3 #(
		.INIT('hba)
	) name31 (
		_w66_,
		_w67_,
		_w68_,
		_w69_
	);
	LUT2 #(
		.INIT('h1)
	) name32 (
		\c0_pad ,
		u_pad,
		_w70_
	);
	LUT2 #(
		.INIT('h8)
	) name33 (
		t_pad,
		v_pad,
		_w71_
	);
	LUT4 #(
		.INIT('h3200)
	) name34 (
		e_pad,
		s_pad,
		t_pad,
		u_pad,
		_w72_
	);
	LUT3 #(
		.INIT('hba)
	) name35 (
		_w70_,
		_w71_,
		_w72_,
		_w73_
	);
	LUT2 #(
		.INIT('h1)
	) name36 (
		\d0_pad ,
		u_pad,
		_w74_
	);
	LUT2 #(
		.INIT('h8)
	) name37 (
		\e0_pad ,
		t_pad,
		_w75_
	);
	LUT4 #(
		.INIT('h3200)
	) name38 (
		l_pad,
		s_pad,
		t_pad,
		u_pad,
		_w76_
	);
	LUT3 #(
		.INIT('hba)
	) name39 (
		_w74_,
		_w75_,
		_w76_,
		_w77_
	);
	LUT2 #(
		.INIT('h1)
	) name40 (
		\e0_pad ,
		u_pad,
		_w78_
	);
	LUT2 #(
		.INIT('h8)
	) name41 (
		\f0_pad ,
		t_pad,
		_w79_
	);
	LUT4 #(
		.INIT('h3200)
	) name42 (
		k_pad,
		s_pad,
		t_pad,
		u_pad,
		_w80_
	);
	LUT3 #(
		.INIT('hba)
	) name43 (
		_w78_,
		_w79_,
		_w80_,
		_w81_
	);
	LUT2 #(
		.INIT('h1)
	) name44 (
		\f0_pad ,
		u_pad,
		_w82_
	);
	LUT2 #(
		.INIT('h8)
	) name45 (
		\g0_pad ,
		t_pad,
		_w83_
	);
	LUT4 #(
		.INIT('h3200)
	) name46 (
		j_pad,
		s_pad,
		t_pad,
		u_pad,
		_w84_
	);
	LUT3 #(
		.INIT('hba)
	) name47 (
		_w82_,
		_w83_,
		_w84_,
		_w85_
	);
	LUT2 #(
		.INIT('h1)
	) name48 (
		\g0_pad ,
		u_pad,
		_w86_
	);
	LUT2 #(
		.INIT('h8)
	) name49 (
		t_pad,
		z_pad,
		_w87_
	);
	LUT4 #(
		.INIT('h3200)
	) name50 (
		i_pad,
		s_pad,
		t_pad,
		u_pad,
		_w88_
	);
	LUT3 #(
		.INIT('hba)
	) name51 (
		_w86_,
		_w87_,
		_w88_,
		_w89_
	);
	LUT2 #(
		.INIT('h1)
	) name52 (
		\h0_pad ,
		u_pad,
		_w90_
	);
	LUT2 #(
		.INIT('h8)
	) name53 (
		\i0_pad ,
		t_pad,
		_w91_
	);
	LUT4 #(
		.INIT('h3200)
	) name54 (
		p_pad,
		s_pad,
		t_pad,
		u_pad,
		_w92_
	);
	LUT3 #(
		.INIT('hba)
	) name55 (
		_w90_,
		_w91_,
		_w92_,
		_w93_
	);
	LUT2 #(
		.INIT('h1)
	) name56 (
		\i0_pad ,
		u_pad,
		_w94_
	);
	LUT2 #(
		.INIT('h8)
	) name57 (
		\j0_pad ,
		t_pad,
		_w95_
	);
	LUT4 #(
		.INIT('h3200)
	) name58 (
		o_pad,
		s_pad,
		t_pad,
		u_pad,
		_w96_
	);
	LUT3 #(
		.INIT('hba)
	) name59 (
		_w94_,
		_w95_,
		_w96_,
		_w97_
	);
	LUT2 #(
		.INIT('h1)
	) name60 (
		\j0_pad ,
		u_pad,
		_w98_
	);
	LUT2 #(
		.INIT('h8)
	) name61 (
		\k0_pad ,
		t_pad,
		_w99_
	);
	LUT4 #(
		.INIT('h3200)
	) name62 (
		n_pad,
		s_pad,
		t_pad,
		u_pad,
		_w100_
	);
	LUT3 #(
		.INIT('hba)
	) name63 (
		_w98_,
		_w99_,
		_w100_,
		_w101_
	);
	assign \a1_pad  = _w41_ ;
	assign \l0_pad  = _w45_ ;
	assign \m0_pad  = _w49_ ;
	assign \n0_pad  = _w53_ ;
	assign \o0_pad  = _w57_ ;
	assign \p0_pad  = _w61_ ;
	assign \q0_pad  = _w65_ ;
	assign \r0_pad  = _w69_ ;
	assign \s0_pad  = _w73_ ;
	assign \t0_pad  = _w77_ ;
	assign \u0_pad  = _w81_ ;
	assign \v0_pad  = _w85_ ;
	assign \w0_pad  = _w89_ ;
	assign \x0_pad  = _w93_ ;
	assign \y0_pad  = _w97_ ;
	assign \z0_pad  = _w101_ ;
endmodule;