module top( \coda0_reg[0]/NET0131  , \coda0_reg[1]/NET0131  , \coda0_reg[2]/NET0131  , \coda1_reg[0]/NET0131  , \coda1_reg[1]/NET0131  , \coda1_reg[2]/NET0131  , \coda2_reg[0]/NET0131  , \coda2_reg[1]/NET0131  , \coda2_reg[2]/NET0131  , \coda3_reg[0]/NET0131  , \coda3_reg[1]/NET0131  , \coda3_reg[2]/NET0131  , \fu1_reg/NET0131  , \fu2_reg/NET0131  , \fu3_reg/NET0131  , \fu4_reg/NET0131  , \grant_o[0]_pad  , \grant_o[1]_pad  , \grant_o[2]_pad  , \grant_o[3]_pad  , \grant_reg[0]/NET0131  , \grant_reg[1]/NET0131  , \grant_reg[2]/NET0131  , \grant_reg[3]/NET0131  , \request1_pad  , \request2_pad  , \request3_pad  , \request4_pad  , \ru1_reg/NET0131  , \ru2_reg/NET0131  , \ru3_reg/NET0131  , \ru4_reg/NET0131  , \stato_reg[0]/NET0131  , \stato_reg[1]/NET0131  , \_al_n0  , \_al_n1  , \g1143/_0_  , \g1144/_0_  , \g1145/_0_  , \g1146/_0_  , \g1147/_0_  , \g1148/_0_  , \g1149/_0_  , \g1150/_0_  , \g1151/_0_  , \g1152/_0_  , \g1153/_0_  , \g1154/_0_  , \g1174/_0_  , \g1175/_0_  , \g1176/_0_  , \g1177/_0_  , \g1238/_0_  , \g1239/_0_  , \g1240/_0_  , \g1241/_0_  , \g1242/_0_  , \g1243/_0_  , \g1244/_0_  , \g1245/_0_  , \g1247/_0_  , \g1248/_0_  , \g1249/_0_  , \g1250/_0_  , \g1520/_0_  );
  input \coda0_reg[0]/NET0131  ;
  input \coda0_reg[1]/NET0131  ;
  input \coda0_reg[2]/NET0131  ;
  input \coda1_reg[0]/NET0131  ;
  input \coda1_reg[1]/NET0131  ;
  input \coda1_reg[2]/NET0131  ;
  input \coda2_reg[0]/NET0131  ;
  input \coda2_reg[1]/NET0131  ;
  input \coda2_reg[2]/NET0131  ;
  input \coda3_reg[0]/NET0131  ;
  input \coda3_reg[1]/NET0131  ;
  input \coda3_reg[2]/NET0131  ;
  input \fu1_reg/NET0131  ;
  input \fu2_reg/NET0131  ;
  input \fu3_reg/NET0131  ;
  input \fu4_reg/NET0131  ;
  input \grant_o[0]_pad  ;
  input \grant_o[1]_pad  ;
  input \grant_o[2]_pad  ;
  input \grant_o[3]_pad  ;
  input \grant_reg[0]/NET0131  ;
  input \grant_reg[1]/NET0131  ;
  input \grant_reg[2]/NET0131  ;
  input \grant_reg[3]/NET0131  ;
  input \request1_pad  ;
  input \request2_pad  ;
  input \request3_pad  ;
  input \request4_pad  ;
  input \ru1_reg/NET0131  ;
  input \ru2_reg/NET0131  ;
  input \ru3_reg/NET0131  ;
  input \ru4_reg/NET0131  ;
  input \stato_reg[0]/NET0131  ;
  input \stato_reg[1]/NET0131  ;
  output \_al_n0  ;
  output \_al_n1  ;
  output \g1143/_0_  ;
  output \g1144/_0_  ;
  output \g1145/_0_  ;
  output \g1146/_0_  ;
  output \g1147/_0_  ;
  output \g1148/_0_  ;
  output \g1149/_0_  ;
  output \g1150/_0_  ;
  output \g1151/_0_  ;
  output \g1152/_0_  ;
  output \g1153/_0_  ;
  output \g1154/_0_  ;
  output \g1174/_0_  ;
  output \g1175/_0_  ;
  output \g1176/_0_  ;
  output \g1177/_0_  ;
  output \g1238/_0_  ;
  output \g1239/_0_  ;
  output \g1240/_0_  ;
  output \g1241/_0_  ;
  output \g1242/_0_  ;
  output \g1243/_0_  ;
  output \g1244/_0_  ;
  output \g1245/_0_  ;
  output \g1247/_0_  ;
  output \g1248/_0_  ;
  output \g1249/_0_  ;
  output \g1250/_0_  ;
  output \g1520/_0_  ;
  wire n35 , n36 , n37 , n38 , n39 , n40 , n41 , n42 , n43 , n44 , n45 , n46 , n47 , n48 , n49 , n50 , n51 , n52 , n53 , n54 , n55 , n56 , n57 , n58 , n59 , n60 , n61 , n62 , n63 , n64 , n65 , n66 , n67 , n68 , n69 , n70 , n71 , n72 , n73 , n74 , n75 , n76 , n77 , n78 , n79 , n80 , n81 , n82 , n83 , n84 , n85 , n86 , n87 , n88 , n89 , n90 , n91 , n92 , n93 , n94 , n95 , n96 , n97 , n98 , n99 , n100 , n101 , n102 , n103 , n104 , n105 , n106 , n107 , n108 , n109 , n110 , n111 , n112 , n113 , n114 , n115 , n116 , n117 , n118 , n119 , n120 , n121 , n122 , n123 , n124 , n125 , n126 , n127 , n128 , n129 , n130 , n131 , n132 , n133 , n134 , n135 , n136 , n137 , n138 , n139 , n140 , n141 , n142 , n143 , n144 , n145 , n146 , n147 , n148 , n149 , n150 , n151 , n152 , n153 , n154 , n155 , n156 , n157 , n158 , n159 , n160 , n161 , n162 , n163 , n164 , n165 , n166 , n167 , n168 , n169 , n170 , n171 , n172 , n173 , n174 , n175 , n176 , n177 , n178 , n179 , n180 , n181 , n182 , n183 , n184 , n185 , n186 , n187 , n188 , n189 , n190 , n191 , n192 , n193 , n194 , n195 , n196 , n197 , n198 , n199 , n200 , n201 , n202 , n203 , n204 , n205 , n206 , n207 , n208 , n209 , n210 , n211 , n212 , n213 , n214 , n215 , n216 , n217 , n218 , n219 , n220 , n221 , n222 , n223 , n224 , n225 , n226 , n227 , n228 , n229 , n230 , n231 , n232 , n233 , n234 , n235 , n236 , n237 , n238 , n239 , n240 , n241 , n242 , n243 , n244 , n245 , n246 , n247 , n248 , n249 , n250 , n251 , n252 , n253 , n254 , n255 , n256 , n257 , n258 , n259 , n260 , n261 , n262 , n263 , n264 , n265 , n266 , n267 , n268 , n269 , n270 , n271 , n272 , n273 , n274 , n275 , n276 , n277 , n278 , n279 , n280 , n281 , n282 , n283 , n284 , n285 , n286 , n287 , n288 , n289 , n290 , n291 , n292 , n293 , n294 , n295 , n296 , n297 , n298 , n299 , n300 , n301 , n302 , n303 , n304 , n305 , n306 , n307 , n308 , n309 , n310 , n311 , n312 , n313 , n314 , n315 , n316 , n317 , n318 , n319 , n320 , n321 , n322 , n323 , n324 , n325 , n326 , n327 , n328 , n329 , n330 , n331 , n332 , n333 , n334 , n335 , n336 , n337 , n338 , n339 , n340 , n341 , n342 , n343 , n344 , n345 , n346 , n347 , n348 , n349 , n350 , n351 , n352 , n353 , n354 , n355 , n356 , n357 , n358 , n359 , n360 , n361 , n362 , n363 , n364 , n365 , n366 , n367 , n368 , n369 , n370 , n371 , n372 , n373 , n374 , n375 , n376 , n377 , n378 , n379 , n380 , n381 , n382 , n383 ;
  assign n35 = ~\fu4_reg/NET0131  & ~\ru3_reg/NET0131  ;
  assign n36 = \ru4_reg/NET0131  & n35 ;
  assign n37 = ~\fu3_reg/NET0131  & \ru3_reg/NET0131  ;
  assign n38 = \coda0_reg[2]/NET0131  & ~n37 ;
  assign n39 = ~n36 & ~n38 ;
  assign n40 = ~\ru2_reg/NET0131  & ~n39 ;
  assign n41 = \fu2_reg/NET0131  & \ru2_reg/NET0131  ;
  assign n42 = \coda0_reg[2]/NET0131  & n41 ;
  assign n43 = ~\ru1_reg/NET0131  & ~n42 ;
  assign n44 = ~n40 & n43 ;
  assign n45 = \fu1_reg/NET0131  & \ru1_reg/NET0131  ;
  assign n46 = ~\coda0_reg[2]/NET0131  & n45 ;
  assign n47 = \stato_reg[0]/NET0131  & ~\stato_reg[1]/NET0131  ;
  assign n48 = ~n46 & n47 ;
  assign n49 = ~n44 & n48 ;
  assign n50 = ~\fu1_reg/NET0131  & ~\fu2_reg/NET0131  ;
  assign n51 = ~\fu3_reg/NET0131  & ~\fu4_reg/NET0131  ;
  assign n52 = n50 & n51 ;
  assign n53 = ~\coda1_reg[2]/NET0131  & \stato_reg[1]/NET0131  ;
  assign n54 = ~n52 & n53 ;
  assign n55 = \coda0_reg[2]/NET0131  & ~\stato_reg[0]/NET0131  ;
  assign n56 = ~\stato_reg[0]/NET0131  & \stato_reg[1]/NET0131  ;
  assign n57 = ~n52 & n56 ;
  assign n58 = ~n55 & ~n57 ;
  assign n59 = ~n54 & ~n58 ;
  assign n60 = ~n49 & ~n59 ;
  assign n61 = \coda0_reg[0]/NET0131  & n45 ;
  assign n62 = \ru1_reg/NET0131  & ~n61 ;
  assign n63 = ~\ru2_reg/NET0131  & \ru4_reg/NET0131  ;
  assign n64 = n35 & n63 ;
  assign n65 = ~\ru2_reg/NET0131  & n37 ;
  assign n66 = ~n64 & ~n65 ;
  assign n67 = ~\fu2_reg/NET0131  & \ru2_reg/NET0131  ;
  assign n68 = \coda0_reg[0]/NET0131  & ~n67 ;
  assign n69 = ~n61 & ~n68 ;
  assign n70 = n66 & n69 ;
  assign n71 = ~n62 & ~n70 ;
  assign n72 = n47 & n71 ;
  assign n73 = ~\coda1_reg[0]/NET0131  & \stato_reg[1]/NET0131  ;
  assign n74 = ~n52 & n73 ;
  assign n75 = \coda0_reg[0]/NET0131  & ~\stato_reg[0]/NET0131  ;
  assign n76 = ~n57 & ~n75 ;
  assign n77 = ~n74 & ~n76 ;
  assign n78 = ~n72 & ~n77 ;
  assign n79 = \coda0_reg[1]/NET0131  & n45 ;
  assign n80 = ~\coda0_reg[1]/NET0131  & n41 ;
  assign n81 = ~\ru1_reg/NET0131  & ~n80 ;
  assign n82 = ~n79 & ~n81 ;
  assign n83 = ~\ru2_reg/NET0131  & ~n36 ;
  assign n84 = \coda0_reg[1]/NET0131  & ~n37 ;
  assign n85 = ~n79 & ~n84 ;
  assign n86 = n83 & n85 ;
  assign n87 = ~n82 & ~n86 ;
  assign n88 = n47 & n87 ;
  assign n89 = ~\coda1_reg[1]/NET0131  & \stato_reg[1]/NET0131  ;
  assign n90 = ~n52 & n89 ;
  assign n91 = \coda0_reg[1]/NET0131  & ~\stato_reg[0]/NET0131  ;
  assign n92 = ~n57 & ~n91 ;
  assign n93 = ~n90 & ~n92 ;
  assign n94 = ~n88 & ~n93 ;
  assign n95 = ~\ru1_reg/NET0131  & n47 ;
  assign n96 = ~\coda1_reg[1]/NET0131  & \fu2_reg/NET0131  ;
  assign n97 = ~\coda0_reg[1]/NET0131  & ~\fu2_reg/NET0131  ;
  assign n98 = \ru2_reg/NET0131  & ~n97 ;
  assign n99 = ~n96 & n98 ;
  assign n100 = n95 & n99 ;
  assign n101 = ~\coda1_reg[1]/NET0131  & \fu3_reg/NET0131  ;
  assign n102 = ~\coda0_reg[1]/NET0131  & ~\fu3_reg/NET0131  ;
  assign n103 = \ru3_reg/NET0131  & ~n102 ;
  assign n104 = ~n101 & n103 ;
  assign n105 = ~\fu4_reg/NET0131  & \ru4_reg/NET0131  ;
  assign n106 = \coda1_reg[1]/NET0131  & ~\ru3_reg/NET0131  ;
  assign n107 = ~n105 & n106 ;
  assign n108 = \coda0_reg[1]/NET0131  & ~\ru3_reg/NET0131  ;
  assign n109 = n105 & n108 ;
  assign n110 = ~n107 & ~n109 ;
  assign n111 = ~n104 & n110 ;
  assign n112 = ~\ru2_reg/NET0131  & n95 ;
  assign n113 = ~n111 & n112 ;
  assign n114 = ~n100 & ~n113 ;
  assign n115 = ~\stato_reg[0]/NET0131  & n52 ;
  assign n116 = ~\stato_reg[1]/NET0131  & n45 ;
  assign n117 = ~\stato_reg[0]/NET0131  & ~\stato_reg[1]/NET0131  ;
  assign n118 = ~n116 & ~n117 ;
  assign n119 = ~n115 & n118 ;
  assign n120 = \coda1_reg[1]/NET0131  & ~n119 ;
  assign n121 = \coda2_reg[1]/NET0131  & \stato_reg[1]/NET0131  ;
  assign n122 = ~\stato_reg[0]/NET0131  & n121 ;
  assign n123 = ~n52 & n122 ;
  assign n124 = ~\fu1_reg/NET0131  & \ru1_reg/NET0131  ;
  assign n125 = n47 & n124 ;
  assign n126 = \coda0_reg[1]/NET0131  & n125 ;
  assign n127 = ~n123 & ~n126 ;
  assign n128 = ~n120 & n127 ;
  assign n129 = n114 & n128 ;
  assign n130 = ~\coda2_reg[2]/NET0131  & \fu2_reg/NET0131  ;
  assign n131 = ~\coda1_reg[2]/NET0131  & ~\fu2_reg/NET0131  ;
  assign n132 = \ru2_reg/NET0131  & ~n131 ;
  assign n133 = ~n130 & n132 ;
  assign n134 = n95 & n133 ;
  assign n135 = ~\coda2_reg[2]/NET0131  & \fu3_reg/NET0131  ;
  assign n136 = ~\coda1_reg[2]/NET0131  & ~\fu3_reg/NET0131  ;
  assign n137 = \ru3_reg/NET0131  & ~n136 ;
  assign n138 = ~n135 & n137 ;
  assign n139 = \coda2_reg[2]/NET0131  & ~\ru3_reg/NET0131  ;
  assign n140 = ~n105 & n139 ;
  assign n141 = \coda1_reg[2]/NET0131  & ~\ru3_reg/NET0131  ;
  assign n142 = n105 & n141 ;
  assign n143 = ~n140 & ~n142 ;
  assign n144 = ~n138 & n143 ;
  assign n145 = n112 & ~n144 ;
  assign n146 = ~n134 & ~n145 ;
  assign n147 = \coda2_reg[2]/NET0131  & ~n119 ;
  assign n148 = \coda3_reg[2]/NET0131  & \stato_reg[1]/NET0131  ;
  assign n149 = ~\stato_reg[0]/NET0131  & n148 ;
  assign n150 = ~n52 & n149 ;
  assign n151 = \coda1_reg[2]/NET0131  & n125 ;
  assign n152 = ~n150 & ~n151 ;
  assign n153 = ~n147 & n152 ;
  assign n154 = n146 & n153 ;
  assign n155 = ~\coda1_reg[2]/NET0131  & \fu2_reg/NET0131  ;
  assign n156 = ~\coda0_reg[2]/NET0131  & ~\fu2_reg/NET0131  ;
  assign n157 = \ru2_reg/NET0131  & ~n156 ;
  assign n158 = ~n155 & n157 ;
  assign n159 = n95 & n158 ;
  assign n160 = ~\coda1_reg[2]/NET0131  & \fu3_reg/NET0131  ;
  assign n161 = ~\coda0_reg[2]/NET0131  & ~\fu3_reg/NET0131  ;
  assign n162 = \ru3_reg/NET0131  & ~n161 ;
  assign n163 = ~n160 & n162 ;
  assign n164 = ~n105 & n141 ;
  assign n165 = \coda0_reg[2]/NET0131  & ~\ru3_reg/NET0131  ;
  assign n166 = n105 & n165 ;
  assign n167 = ~n164 & ~n166 ;
  assign n168 = ~n163 & n167 ;
  assign n169 = n112 & ~n168 ;
  assign n170 = ~n159 & ~n169 ;
  assign n171 = \coda1_reg[2]/NET0131  & ~n119 ;
  assign n172 = \coda2_reg[2]/NET0131  & \stato_reg[1]/NET0131  ;
  assign n173 = ~\stato_reg[0]/NET0131  & n172 ;
  assign n174 = ~n52 & n173 ;
  assign n175 = \coda0_reg[2]/NET0131  & n125 ;
  assign n176 = ~n174 & ~n175 ;
  assign n177 = ~n171 & n176 ;
  assign n178 = n170 & n177 ;
  assign n179 = ~\coda1_reg[0]/NET0131  & \fu2_reg/NET0131  ;
  assign n180 = ~\coda0_reg[0]/NET0131  & ~\fu2_reg/NET0131  ;
  assign n181 = \ru2_reg/NET0131  & ~n180 ;
  assign n182 = ~n179 & n181 ;
  assign n183 = n95 & n182 ;
  assign n184 = ~\coda1_reg[0]/NET0131  & \fu3_reg/NET0131  ;
  assign n185 = ~\coda0_reg[0]/NET0131  & ~\fu3_reg/NET0131  ;
  assign n186 = \ru3_reg/NET0131  & ~n185 ;
  assign n187 = ~n184 & n186 ;
  assign n188 = \coda1_reg[0]/NET0131  & ~\ru3_reg/NET0131  ;
  assign n189 = ~n105 & n188 ;
  assign n190 = \coda0_reg[0]/NET0131  & ~\ru3_reg/NET0131  ;
  assign n191 = n105 & n190 ;
  assign n192 = ~n189 & ~n191 ;
  assign n193 = ~n187 & n192 ;
  assign n194 = n112 & ~n193 ;
  assign n195 = ~n183 & ~n194 ;
  assign n196 = \coda1_reg[0]/NET0131  & ~n119 ;
  assign n197 = \coda2_reg[0]/NET0131  & \stato_reg[1]/NET0131  ;
  assign n198 = ~\stato_reg[0]/NET0131  & n197 ;
  assign n199 = ~n52 & n198 ;
  assign n200 = \coda0_reg[0]/NET0131  & n125 ;
  assign n201 = ~n199 & ~n200 ;
  assign n202 = ~n196 & n201 ;
  assign n203 = n195 & n202 ;
  assign n204 = ~\coda2_reg[0]/NET0131  & \fu2_reg/NET0131  ;
  assign n205 = ~\coda1_reg[0]/NET0131  & ~\fu2_reg/NET0131  ;
  assign n206 = \ru2_reg/NET0131  & ~n205 ;
  assign n207 = ~n204 & n206 ;
  assign n208 = n95 & n207 ;
  assign n209 = ~\coda2_reg[0]/NET0131  & \fu3_reg/NET0131  ;
  assign n210 = ~\coda1_reg[0]/NET0131  & ~\fu3_reg/NET0131  ;
  assign n211 = \ru3_reg/NET0131  & ~n210 ;
  assign n212 = ~n209 & n211 ;
  assign n213 = \coda2_reg[0]/NET0131  & ~\ru3_reg/NET0131  ;
  assign n214 = ~n105 & n213 ;
  assign n215 = n105 & n188 ;
  assign n216 = ~n214 & ~n215 ;
  assign n217 = ~n212 & n216 ;
  assign n218 = n112 & ~n217 ;
  assign n219 = ~n208 & ~n218 ;
  assign n220 = \coda2_reg[0]/NET0131  & ~n119 ;
  assign n221 = \coda3_reg[0]/NET0131  & \stato_reg[1]/NET0131  ;
  assign n222 = ~\stato_reg[0]/NET0131  & n221 ;
  assign n223 = ~n52 & n222 ;
  assign n224 = \coda1_reg[0]/NET0131  & n125 ;
  assign n225 = ~n223 & ~n224 ;
  assign n226 = ~n220 & n225 ;
  assign n227 = n219 & n226 ;
  assign n228 = ~\coda2_reg[1]/NET0131  & \fu2_reg/NET0131  ;
  assign n229 = ~\coda1_reg[1]/NET0131  & ~\fu2_reg/NET0131  ;
  assign n230 = \ru2_reg/NET0131  & ~n229 ;
  assign n231 = ~n228 & n230 ;
  assign n232 = n95 & n231 ;
  assign n233 = ~\coda2_reg[1]/NET0131  & \fu3_reg/NET0131  ;
  assign n234 = ~\coda1_reg[1]/NET0131  & ~\fu3_reg/NET0131  ;
  assign n235 = \ru3_reg/NET0131  & ~n234 ;
  assign n236 = ~n233 & n235 ;
  assign n237 = \coda2_reg[1]/NET0131  & ~\ru3_reg/NET0131  ;
  assign n238 = ~n105 & n237 ;
  assign n239 = n105 & n106 ;
  assign n240 = ~n238 & ~n239 ;
  assign n241 = ~n236 & n240 ;
  assign n242 = n112 & ~n241 ;
  assign n243 = ~n232 & ~n242 ;
  assign n244 = \ru1_reg/NET0131  & n47 ;
  assign n245 = ~\coda1_reg[1]/NET0131  & ~\fu1_reg/NET0131  ;
  assign n246 = ~\coda2_reg[1]/NET0131  & \fu1_reg/NET0131  ;
  assign n247 = ~n245 & ~n246 ;
  assign n248 = n244 & n247 ;
  assign n249 = ~\coda3_reg[1]/NET0131  & \stato_reg[1]/NET0131  ;
  assign n250 = ~n52 & n249 ;
  assign n251 = \coda2_reg[1]/NET0131  & ~\stato_reg[0]/NET0131  ;
  assign n252 = ~n57 & ~n251 ;
  assign n253 = ~n250 & ~n252 ;
  assign n254 = ~n248 & ~n253 ;
  assign n255 = n243 & n254 ;
  assign n256 = ~\coda3_reg[0]/NET0131  & \fu2_reg/NET0131  ;
  assign n257 = ~\ru1_reg/NET0131  & \ru2_reg/NET0131  ;
  assign n258 = ~\coda2_reg[0]/NET0131  & ~\fu2_reg/NET0131  ;
  assign n259 = n257 & ~n258 ;
  assign n260 = ~n256 & n259 ;
  assign n261 = n47 & n260 ;
  assign n262 = ~\coda3_reg[0]/NET0131  & \fu3_reg/NET0131  ;
  assign n263 = ~\coda2_reg[0]/NET0131  & ~\fu3_reg/NET0131  ;
  assign n264 = \ru3_reg/NET0131  & ~n263 ;
  assign n265 = ~n262 & n264 ;
  assign n266 = \coda3_reg[0]/NET0131  & ~\ru3_reg/NET0131  ;
  assign n267 = ~n105 & n266 ;
  assign n268 = n105 & n213 ;
  assign n269 = ~n267 & ~n268 ;
  assign n270 = ~n265 & n269 ;
  assign n271 = ~\ru1_reg/NET0131  & ~\ru2_reg/NET0131  ;
  assign n272 = n47 & n271 ;
  assign n273 = ~n270 & n272 ;
  assign n274 = ~n261 & ~n273 ;
  assign n275 = \coda3_reg[0]/NET0131  & ~n119 ;
  assign n276 = \coda2_reg[0]/NET0131  & n125 ;
  assign n277 = ~n275 & ~n276 ;
  assign n278 = n274 & n277 ;
  assign n279 = ~\coda3_reg[1]/NET0131  & \fu2_reg/NET0131  ;
  assign n280 = ~\coda2_reg[1]/NET0131  & ~\fu2_reg/NET0131  ;
  assign n281 = n257 & ~n280 ;
  assign n282 = ~n279 & n281 ;
  assign n283 = n47 & n282 ;
  assign n284 = ~\coda3_reg[1]/NET0131  & \fu3_reg/NET0131  ;
  assign n285 = ~\coda2_reg[1]/NET0131  & ~\fu3_reg/NET0131  ;
  assign n286 = \ru3_reg/NET0131  & ~n285 ;
  assign n287 = ~n284 & n286 ;
  assign n288 = \coda3_reg[1]/NET0131  & ~\ru3_reg/NET0131  ;
  assign n289 = ~n105 & n288 ;
  assign n290 = n105 & n237 ;
  assign n291 = ~n289 & ~n290 ;
  assign n292 = ~n287 & n291 ;
  assign n293 = n272 & ~n292 ;
  assign n294 = ~n283 & ~n293 ;
  assign n295 = \coda2_reg[1]/NET0131  & n125 ;
  assign n296 = \coda3_reg[1]/NET0131  & ~n119 ;
  assign n297 = ~n295 & ~n296 ;
  assign n298 = n294 & n297 ;
  assign n299 = ~\coda3_reg[2]/NET0131  & \fu2_reg/NET0131  ;
  assign n300 = ~\coda2_reg[2]/NET0131  & ~\fu2_reg/NET0131  ;
  assign n301 = n257 & ~n300 ;
  assign n302 = ~n299 & n301 ;
  assign n303 = n47 & n302 ;
  assign n304 = ~\coda3_reg[2]/NET0131  & \fu3_reg/NET0131  ;
  assign n305 = ~\coda2_reg[2]/NET0131  & ~\fu3_reg/NET0131  ;
  assign n306 = \ru3_reg/NET0131  & ~n305 ;
  assign n307 = ~n304 & n306 ;
  assign n308 = \coda3_reg[2]/NET0131  & ~\ru3_reg/NET0131  ;
  assign n309 = ~n105 & n308 ;
  assign n310 = n105 & n139 ;
  assign n311 = ~n309 & ~n310 ;
  assign n312 = ~n307 & n311 ;
  assign n313 = n272 & ~n312 ;
  assign n314 = ~n303 & ~n313 ;
  assign n315 = \coda2_reg[2]/NET0131  & n125 ;
  assign n316 = \coda3_reg[2]/NET0131  & ~n119 ;
  assign n317 = ~n315 & ~n316 ;
  assign n318 = n314 & n317 ;
  assign n319 = \grant_reg[0]/NET0131  & ~\stato_reg[1]/NET0131  ;
  assign n320 = \grant_reg[0]/NET0131  & ~\stato_reg[0]/NET0131  ;
  assign n321 = n52 & n320 ;
  assign n322 = ~n319 & ~n321 ;
  assign n323 = \coda0_reg[1]/NET0131  & \stato_reg[1]/NET0131  ;
  assign n324 = ~\stato_reg[0]/NET0131  & n323 ;
  assign n325 = ~n52 & n324 ;
  assign n326 = \coda0_reg[0]/NET0131  & \coda0_reg[2]/NET0131  ;
  assign n327 = n325 & n326 ;
  assign n328 = n322 & ~n327 ;
  assign n329 = \grant_reg[1]/NET0131  & ~\stato_reg[1]/NET0131  ;
  assign n330 = \grant_reg[1]/NET0131  & ~\stato_reg[0]/NET0131  ;
  assign n331 = n52 & n330 ;
  assign n332 = ~n329 & ~n331 ;
  assign n333 = ~\coda0_reg[1]/NET0131  & \stato_reg[1]/NET0131  ;
  assign n334 = ~\stato_reg[0]/NET0131  & n333 ;
  assign n335 = ~n52 & n334 ;
  assign n336 = \coda0_reg[0]/NET0131  & ~\coda0_reg[2]/NET0131  ;
  assign n337 = n335 & n336 ;
  assign n338 = n332 & ~n337 ;
  assign n339 = \grant_reg[2]/NET0131  & ~\stato_reg[1]/NET0131  ;
  assign n340 = \grant_reg[2]/NET0131  & ~\stato_reg[0]/NET0131  ;
  assign n341 = n52 & n340 ;
  assign n342 = ~n339 & ~n341 ;
  assign n343 = ~\coda0_reg[0]/NET0131  & ~\coda0_reg[2]/NET0131  ;
  assign n344 = n325 & n343 ;
  assign n345 = n342 & ~n344 ;
  assign n346 = \grant_reg[3]/NET0131  & ~\stato_reg[1]/NET0131  ;
  assign n347 = \grant_reg[3]/NET0131  & ~\stato_reg[0]/NET0131  ;
  assign n348 = n52 & n347 ;
  assign n349 = ~n346 & ~n348 ;
  assign n350 = ~\coda0_reg[0]/NET0131  & \coda0_reg[2]/NET0131  ;
  assign n351 = n335 & n350 ;
  assign n352 = n349 & ~n351 ;
  assign n353 = \fu1_reg/NET0131  & ~\stato_reg[0]/NET0131  ;
  assign n354 = ~n244 & ~n353 ;
  assign n355 = \ru2_reg/NET0131  & n47 ;
  assign n356 = \fu2_reg/NET0131  & ~\stato_reg[0]/NET0131  ;
  assign n357 = ~n355 & ~n356 ;
  assign n358 = \ru3_reg/NET0131  & n47 ;
  assign n359 = \fu3_reg/NET0131  & ~\stato_reg[0]/NET0131  ;
  assign n360 = ~n358 & ~n359 ;
  assign n361 = \ru4_reg/NET0131  & n47 ;
  assign n362 = \fu4_reg/NET0131  & ~\stato_reg[0]/NET0131  ;
  assign n363 = ~n361 & ~n362 ;
  assign n364 = \grant_reg[0]/NET0131  & n47 ;
  assign n365 = \grant_o[0]_pad  & ~\stato_reg[0]/NET0131  ;
  assign n366 = ~n364 & ~n365 ;
  assign n367 = \grant_reg[1]/NET0131  & n47 ;
  assign n368 = \grant_o[1]_pad  & ~\stato_reg[0]/NET0131  ;
  assign n369 = ~n367 & ~n368 ;
  assign n370 = \grant_reg[2]/NET0131  & n47 ;
  assign n371 = \grant_o[2]_pad  & ~\stato_reg[0]/NET0131  ;
  assign n372 = ~n370 & ~n371 ;
  assign n373 = \grant_reg[3]/NET0131  & n47 ;
  assign n374 = \grant_o[3]_pad  & ~\stato_reg[0]/NET0131  ;
  assign n375 = ~n373 & ~n374 ;
  assign n376 = \request1_pad  & ~\stato_reg[0]/NET0131  ;
  assign n377 = ~n244 & ~n376 ;
  assign n378 = \request2_pad  & ~\stato_reg[0]/NET0131  ;
  assign n379 = ~n355 & ~n378 ;
  assign n380 = \request3_pad  & ~\stato_reg[0]/NET0131  ;
  assign n381 = ~n358 & ~n380 ;
  assign n382 = \request4_pad  & ~\stato_reg[0]/NET0131  ;
  assign n383 = ~n361 & ~n382 ;
  assign \_al_n0  = 1'b0 ;
  assign \_al_n1  = ~1'b0 ;
  assign \g1143/_0_  = ~n60 ;
  assign \g1144/_0_  = ~n78 ;
  assign \g1145/_0_  = ~n94 ;
  assign \g1146/_0_  = ~n129 ;
  assign \g1147/_0_  = ~n154 ;
  assign \g1148/_0_  = ~n178 ;
  assign \g1149/_0_  = ~n203 ;
  assign \g1150/_0_  = ~n227 ;
  assign \g1151/_0_  = ~n255 ;
  assign \g1152/_0_  = ~n278 ;
  assign \g1153/_0_  = ~n298 ;
  assign \g1154/_0_  = ~n318 ;
  assign \g1174/_0_  = ~n328 ;
  assign \g1175/_0_  = ~n338 ;
  assign \g1176/_0_  = ~n345 ;
  assign \g1177/_0_  = ~n352 ;
  assign \g1238/_0_  = ~n354 ;
  assign \g1239/_0_  = ~n357 ;
  assign \g1240/_0_  = ~n360 ;
  assign \g1241/_0_  = ~n363 ;
  assign \g1242/_0_  = ~n366 ;
  assign \g1243/_0_  = ~n369 ;
  assign \g1244/_0_  = ~n372 ;
  assign \g1245/_0_  = ~n375 ;
  assign \g1247/_0_  = ~n377 ;
  assign \g1248/_0_  = ~n379 ;
  assign \g1249/_0_  = ~n381 ;
  assign \g1250/_0_  = ~n383 ;
  assign \g1520/_0_  = ~\stato_reg[0]/NET0131  ;
endmodule
