module top (\P1_B_reg/NET0131 , \P1_IR_reg[0]/NET0131 , \P1_IR_reg[10]/NET0131 , \P1_IR_reg[11]/NET0131 , \P1_IR_reg[12]/NET0131 , \P1_IR_reg[13]/NET0131 , \P1_IR_reg[14]/NET0131 , \P1_IR_reg[15]/NET0131 , \P1_IR_reg[16]/NET0131 , \P1_IR_reg[17]/NET0131 , \P1_IR_reg[18]/NET0131 , \P1_IR_reg[19]/NET0131 , \P1_IR_reg[1]/NET0131 , \P1_IR_reg[20]/NET0131 , \P1_IR_reg[21]/NET0131 , \P1_IR_reg[22]/NET0131 , \P1_IR_reg[23]/NET0131 , \P1_IR_reg[24]/NET0131 , \P1_IR_reg[25]/NET0131 , \P1_IR_reg[26]/NET0131 , \P1_IR_reg[27]/NET0131 , \P1_IR_reg[28]/NET0131 , \P1_IR_reg[29]/NET0131 , \P1_IR_reg[2]/NET0131 , \P1_IR_reg[30]/NET0131 , \P1_IR_reg[31]/NET0131 , \P1_IR_reg[3]/NET0131 , \P1_IR_reg[4]/NET0131 , \P1_IR_reg[5]/NET0131 , \P1_IR_reg[6]/NET0131 , \P1_IR_reg[7]/NET0131 , \P1_IR_reg[8]/NET0131 , \P1_IR_reg[9]/NET0131 , \P1_addr_reg[0]/NET0131 , \P1_addr_reg[10]/NET0131 , \P1_addr_reg[11]/NET0131 , \P1_addr_reg[12]/NET0131 , \P1_addr_reg[13]/NET0131 , \P1_addr_reg[14]/NET0131 , \P1_addr_reg[15]/NET0131 , \P1_addr_reg[16]/NET0131 , \P1_addr_reg[17]/NET0131 , \P1_addr_reg[18]/NET0131 , \P1_addr_reg[19]/NET0131 , \P1_addr_reg[1]/NET0131 , \P1_addr_reg[2]/NET0131 , \P1_addr_reg[3]/NET0131 , \P1_addr_reg[4]/NET0131 , \P1_addr_reg[5]/NET0131 , \P1_addr_reg[6]/NET0131 , \P1_addr_reg[7]/NET0131 , \P1_addr_reg[8]/NET0131 , \P1_addr_reg[9]/NET0131 , \P1_d_reg[0]/NET0131 , \P1_d_reg[1]/NET0131 , \P1_datao_reg[0]/NET0131 , \P1_datao_reg[10]/NET0131 , \P1_datao_reg[11]/NET0131 , \P1_datao_reg[12]/NET0131 , \P1_datao_reg[13]/NET0131 , \P1_datao_reg[14]/NET0131 , \P1_datao_reg[15]/NET0131 , \P1_datao_reg[16]/NET0131 , \P1_datao_reg[17]/NET0131 , \P1_datao_reg[18]/NET0131 , \P1_datao_reg[19]/NET0131 , \P1_datao_reg[1]/NET0131 , \P1_datao_reg[20]/NET0131 , \P1_datao_reg[21]/NET0131 , \P1_datao_reg[22]/NET0131 , \P1_datao_reg[23]/NET0131 , \P1_datao_reg[24]/NET0131 , \P1_datao_reg[25]/NET0131 , \P1_datao_reg[26]/NET0131 , \P1_datao_reg[27]/NET0131 , \P1_datao_reg[28]/NET0131 , \P1_datao_reg[29]/NET0131 , \P1_datao_reg[2]/NET0131 , \P1_datao_reg[30]/NET0131 , \P1_datao_reg[31]/NET0131 , \P1_datao_reg[3]/NET0131 , \P1_datao_reg[4]/NET0131 , \P1_datao_reg[5]/NET0131 , \P1_datao_reg[6]/NET0131 , \P1_datao_reg[7]/NET0131 , \P1_datao_reg[8]/NET0131 , \P1_datao_reg[9]/NET0131 , \P1_rd_reg/NET0131 , \P1_reg0_reg[0]/NET0131 , \P1_reg0_reg[10]/NET0131 , \P1_reg0_reg[11]/NET0131 , \P1_reg0_reg[12]/NET0131 , \P1_reg0_reg[13]/NET0131 , \P1_reg0_reg[14]/NET0131 , \P1_reg0_reg[15]/NET0131 , \P1_reg0_reg[16]/NET0131 , \P1_reg0_reg[17]/NET0131 , \P1_reg0_reg[18]/NET0131 , \P1_reg0_reg[19]/NET0131 , \P1_reg0_reg[1]/NET0131 , \P1_reg0_reg[20]/NET0131 , \P1_reg0_reg[21]/NET0131 , \P1_reg0_reg[22]/NET0131 , \P1_reg0_reg[23]/NET0131 , \P1_reg0_reg[24]/NET0131 , \P1_reg0_reg[25]/NET0131 , \P1_reg0_reg[26]/NET0131 , \P1_reg0_reg[27]/NET0131 , \P1_reg0_reg[28]/NET0131 , \P1_reg0_reg[29]/NET0131 , \P1_reg0_reg[2]/NET0131 , \P1_reg0_reg[30]/NET0131 , \P1_reg0_reg[31]/NET0131 , \P1_reg0_reg[3]/NET0131 , \P1_reg0_reg[4]/NET0131 , \P1_reg0_reg[5]/NET0131 , \P1_reg0_reg[6]/NET0131 , \P1_reg0_reg[7]/NET0131 , \P1_reg0_reg[8]/NET0131 , \P1_reg0_reg[9]/NET0131 , \P1_reg1_reg[0]/NET0131 , \P1_reg1_reg[10]/NET0131 , \P1_reg1_reg[11]/NET0131 , \P1_reg1_reg[12]/NET0131 , \P1_reg1_reg[13]/NET0131 , \P1_reg1_reg[14]/NET0131 , \P1_reg1_reg[15]/NET0131 , \P1_reg1_reg[16]/NET0131 , \P1_reg1_reg[17]/NET0131 , \P1_reg1_reg[18]/NET0131 , \P1_reg1_reg[19]/NET0131 , \P1_reg1_reg[1]/NET0131 , \P1_reg1_reg[20]/NET0131 , \P1_reg1_reg[21]/NET0131 , \P1_reg1_reg[22]/NET0131 , \P1_reg1_reg[23]/NET0131 , \P1_reg1_reg[24]/NET0131 , \P1_reg1_reg[25]/NET0131 , \P1_reg1_reg[26]/NET0131 , \P1_reg1_reg[27]/NET0131 , \P1_reg1_reg[28]/NET0131 , \P1_reg1_reg[29]/NET0131 , \P1_reg1_reg[2]/NET0131 , \P1_reg1_reg[30]/NET0131 , \P1_reg1_reg[31]/NET0131 , \P1_reg1_reg[3]/NET0131 , \P1_reg1_reg[4]/NET0131 , \P1_reg1_reg[5]/NET0131 , \P1_reg1_reg[6]/NET0131 , \P1_reg1_reg[7]/NET0131 , \P1_reg1_reg[8]/NET0131 , \P1_reg1_reg[9]/NET0131 , \P1_reg2_reg[0]/NET0131 , \P1_reg2_reg[10]/NET0131 , \P1_reg2_reg[11]/NET0131 , \P1_reg2_reg[12]/NET0131 , \P1_reg2_reg[13]/NET0131 , \P1_reg2_reg[14]/NET0131 , \P1_reg2_reg[15]/NET0131 , \P1_reg2_reg[16]/NET0131 , \P1_reg2_reg[17]/NET0131 , \P1_reg2_reg[18]/NET0131 , \P1_reg2_reg[19]/NET0131 , \P1_reg2_reg[1]/NET0131 , \P1_reg2_reg[20]/NET0131 , \P1_reg2_reg[21]/NET0131 , \P1_reg2_reg[22]/NET0131 , \P1_reg2_reg[23]/NET0131 , \P1_reg2_reg[24]/NET0131 , \P1_reg2_reg[25]/NET0131 , \P1_reg2_reg[26]/NET0131 , \P1_reg2_reg[27]/NET0131 , \P1_reg2_reg[28]/NET0131 , \P1_reg2_reg[29]/NET0131 , \P1_reg2_reg[2]/NET0131 , \P1_reg2_reg[30]/NET0131 , \P1_reg2_reg[31]/NET0131 , \P1_reg2_reg[3]/NET0131 , \P1_reg2_reg[4]/NET0131 , \P1_reg2_reg[5]/NET0131 , \P1_reg2_reg[6]/NET0131 , \P1_reg2_reg[7]/NET0131 , \P1_reg2_reg[8]/NET0131 , \P1_reg2_reg[9]/NET0131 , \P1_reg3_reg[0]/NET0131 , \P1_reg3_reg[10]/NET0131 , \P1_reg3_reg[11]/NET0131 , \P1_reg3_reg[12]/NET0131 , \P1_reg3_reg[13]/NET0131 , \P1_reg3_reg[14]/NET0131 , \P1_reg3_reg[15]/NET0131 , \P1_reg3_reg[16]/NET0131 , \P1_reg3_reg[17]/NET0131 , \P1_reg3_reg[18]/NET0131 , \P1_reg3_reg[19]/NET0131 , \P1_reg3_reg[1]/NET0131 , \P1_reg3_reg[20]/NET0131 , \P1_reg3_reg[21]/NET0131 , \P1_reg3_reg[22]/NET0131 , \P1_reg3_reg[23]/NET0131 , \P1_reg3_reg[24]/NET0131 , \P1_reg3_reg[25]/NET0131 , \P1_reg3_reg[26]/NET0131 , \P1_reg3_reg[27]/NET0131 , \P1_reg3_reg[28]/NET0131 , \P1_reg3_reg[2]/NET0131 , \P1_reg3_reg[3]/NET0131 , \P1_reg3_reg[4]/NET0131 , \P1_reg3_reg[5]/NET0131 , \P1_reg3_reg[6]/NET0131 , \P1_reg3_reg[7]/NET0131 , \P1_reg3_reg[8]/NET0131 , \P1_reg3_reg[9]/NET0131 , \P1_state_reg[0]/NET0131 , \P1_wr_reg/NET0131 , \P2_B_reg/NET0131 , \P2_IR_reg[0]/NET0131 , \P2_IR_reg[10]/NET0131 , \P2_IR_reg[11]/NET0131 , \P2_IR_reg[12]/NET0131 , \P2_IR_reg[13]/NET0131 , \P2_IR_reg[14]/NET0131 , \P2_IR_reg[15]/NET0131 , \P2_IR_reg[16]/NET0131 , \P2_IR_reg[17]/NET0131 , \P2_IR_reg[18]/NET0131 , \P2_IR_reg[19]/NET0131 , \P2_IR_reg[1]/NET0131 , \P2_IR_reg[20]/NET0131 , \P2_IR_reg[21]/NET0131 , \P2_IR_reg[22]/NET0131 , \P2_IR_reg[23]/NET0131 , \P2_IR_reg[24]/NET0131 , \P2_IR_reg[25]/NET0131 , \P2_IR_reg[26]/NET0131 , \P2_IR_reg[27]/NET0131 , \P2_IR_reg[28]/NET0131 , \P2_IR_reg[29]/NET0131 , \P2_IR_reg[2]/NET0131 , \P2_IR_reg[30]/NET0131 , \P2_IR_reg[31]/NET0131 , \P2_IR_reg[3]/NET0131 , \P2_IR_reg[4]/NET0131 , \P2_IR_reg[5]/NET0131 , \P2_IR_reg[6]/NET0131 , \P2_IR_reg[7]/NET0131 , \P2_IR_reg[8]/NET0131 , \P2_IR_reg[9]/NET0131 , \P2_addr_reg[0]/NET0131 , \P2_addr_reg[10]/NET0131 , \P2_addr_reg[11]/NET0131 , \P2_addr_reg[12]/NET0131 , \P2_addr_reg[13]/NET0131 , \P2_addr_reg[14]/NET0131 , \P2_addr_reg[15]/NET0131 , \P2_addr_reg[16]/NET0131 , \P2_addr_reg[17]/NET0131 , \P2_addr_reg[18]/NET0131 , \P2_addr_reg[19]/NET0131 , \P2_addr_reg[1]/NET0131 , \P2_addr_reg[2]/NET0131 , \P2_addr_reg[3]/NET0131 , \P2_addr_reg[4]/NET0131 , \P2_addr_reg[5]/NET0131 , \P2_addr_reg[6]/NET0131 , \P2_addr_reg[7]/NET0131 , \P2_addr_reg[8]/NET0131 , \P2_addr_reg[9]/NET0131 , \P2_d_reg[0]/NET0131 , \P2_d_reg[1]/NET0131 , \P2_datao_reg[0]/NET0131 , \P2_datao_reg[10]/NET0131 , \P2_datao_reg[11]/NET0131 , \P2_datao_reg[12]/NET0131 , \P2_datao_reg[13]/NET0131 , \P2_datao_reg[14]/NET0131 , \P2_datao_reg[15]/NET0131 , \P2_datao_reg[16]/NET0131 , \P2_datao_reg[17]/NET0131 , \P2_datao_reg[18]/NET0131 , \P2_datao_reg[19]/NET0131 , \P2_datao_reg[1]/NET0131 , \P2_datao_reg[20]/NET0131 , \P2_datao_reg[21]/NET0131 , \P2_datao_reg[22]/NET0131 , \P2_datao_reg[23]/NET0131 , \P2_datao_reg[24]/NET0131 , \P2_datao_reg[25]/NET0131 , \P2_datao_reg[26]/NET0131 , \P2_datao_reg[27]/NET0131 , \P2_datao_reg[28]/NET0131 , \P2_datao_reg[29]/NET0131 , \P2_datao_reg[2]/NET0131 , \P2_datao_reg[30]/NET0131 , \P2_datao_reg[31]/NET0131 , \P2_datao_reg[3]/NET0131 , \P2_datao_reg[4]/NET0131 , \P2_datao_reg[5]/NET0131 , \P2_datao_reg[6]/NET0131 , \P2_datao_reg[7]/NET0131 , \P2_datao_reg[8]/NET0131 , \P2_datao_reg[9]/NET0131 , \P2_rd_reg/NET0131 , \P2_reg0_reg[0]/NET0131 , \P2_reg0_reg[10]/NET0131 , \P2_reg0_reg[11]/NET0131 , \P2_reg0_reg[12]/NET0131 , \P2_reg0_reg[13]/NET0131 , \P2_reg0_reg[14]/NET0131 , \P2_reg0_reg[15]/NET0131 , \P2_reg0_reg[16]/NET0131 , \P2_reg0_reg[17]/NET0131 , \P2_reg0_reg[18]/NET0131 , \P2_reg0_reg[19]/NET0131 , \P2_reg0_reg[1]/NET0131 , \P2_reg0_reg[20]/NET0131 , \P2_reg0_reg[21]/NET0131 , \P2_reg0_reg[22]/NET0131 , \P2_reg0_reg[23]/NET0131 , \P2_reg0_reg[24]/NET0131 , \P2_reg0_reg[25]/NET0131 , \P2_reg0_reg[26]/NET0131 , \P2_reg0_reg[27]/NET0131 , \P2_reg0_reg[28]/NET0131 , \P2_reg0_reg[29]/NET0131 , \P2_reg0_reg[2]/NET0131 , \P2_reg0_reg[30]/NET0131 , \P2_reg0_reg[31]/NET0131 , \P2_reg0_reg[3]/NET0131 , \P2_reg0_reg[4]/NET0131 , \P2_reg0_reg[5]/NET0131 , \P2_reg0_reg[6]/NET0131 , \P2_reg0_reg[7]/NET0131 , \P2_reg0_reg[8]/NET0131 , \P2_reg0_reg[9]/NET0131 , \P2_reg1_reg[0]/NET0131 , \P2_reg1_reg[10]/NET0131 , \P2_reg1_reg[11]/NET0131 , \P2_reg1_reg[12]/NET0131 , \P2_reg1_reg[13]/NET0131 , \P2_reg1_reg[14]/NET0131 , \P2_reg1_reg[15]/NET0131 , \P2_reg1_reg[16]/NET0131 , \P2_reg1_reg[17]/NET0131 , \P2_reg1_reg[18]/NET0131 , \P2_reg1_reg[19]/NET0131 , \P2_reg1_reg[1]/NET0131 , \P2_reg1_reg[20]/NET0131 , \P2_reg1_reg[21]/NET0131 , \P2_reg1_reg[22]/NET0131 , \P2_reg1_reg[23]/NET0131 , \P2_reg1_reg[24]/NET0131 , \P2_reg1_reg[25]/NET0131 , \P2_reg1_reg[26]/NET0131 , \P2_reg1_reg[27]/NET0131 , \P2_reg1_reg[28]/NET0131 , \P2_reg1_reg[29]/NET0131 , \P2_reg1_reg[2]/NET0131 , \P2_reg1_reg[30]/NET0131 , \P2_reg1_reg[31]/NET0131 , \P2_reg1_reg[3]/NET0131 , \P2_reg1_reg[4]/NET0131 , \P2_reg1_reg[5]/NET0131 , \P2_reg1_reg[6]/NET0131 , \P2_reg1_reg[7]/NET0131 , \P2_reg1_reg[8]/NET0131 , \P2_reg1_reg[9]/NET0131 , \P2_reg2_reg[0]/NET0131 , \P2_reg2_reg[10]/NET0131 , \P2_reg2_reg[11]/NET0131 , \P2_reg2_reg[12]/NET0131 , \P2_reg2_reg[13]/NET0131 , \P2_reg2_reg[14]/NET0131 , \P2_reg2_reg[15]/NET0131 , \P2_reg2_reg[16]/NET0131 , \P2_reg2_reg[17]/NET0131 , \P2_reg2_reg[18]/NET0131 , \P2_reg2_reg[19]/NET0131 , \P2_reg2_reg[1]/NET0131 , \P2_reg2_reg[20]/NET0131 , \P2_reg2_reg[21]/NET0131 , \P2_reg2_reg[22]/NET0131 , \P2_reg2_reg[23]/NET0131 , \P2_reg2_reg[24]/NET0131 , \P2_reg2_reg[25]/NET0131 , \P2_reg2_reg[26]/NET0131 , \P2_reg2_reg[27]/NET0131 , \P2_reg2_reg[28]/NET0131 , \P2_reg2_reg[29]/NET0131 , \P2_reg2_reg[2]/NET0131 , \P2_reg2_reg[30]/NET0131 , \P2_reg2_reg[31]/NET0131 , \P2_reg2_reg[3]/NET0131 , \P2_reg2_reg[4]/NET0131 , \P2_reg2_reg[5]/NET0131 , \P2_reg2_reg[6]/NET0131 , \P2_reg2_reg[7]/NET0131 , \P2_reg2_reg[8]/NET0131 , \P2_reg2_reg[9]/NET0131 , \P2_reg3_reg[0]/NET0131 , \P2_reg3_reg[10]/NET0131 , \P2_reg3_reg[11]/NET0131 , \P2_reg3_reg[12]/NET0131 , \P2_reg3_reg[13]/NET0131 , \P2_reg3_reg[14]/NET0131 , \P2_reg3_reg[15]/NET0131 , \P2_reg3_reg[16]/NET0131 , \P2_reg3_reg[17]/NET0131 , \P2_reg3_reg[18]/NET0131 , \P2_reg3_reg[19]/NET0131 , \P2_reg3_reg[1]/NET0131 , \P2_reg3_reg[20]/NET0131 , \P2_reg3_reg[21]/NET0131 , \P2_reg3_reg[22]/NET0131 , \P2_reg3_reg[23]/NET0131 , \P2_reg3_reg[24]/NET0131 , \P2_reg3_reg[25]/NET0131 , \P2_reg3_reg[26]/NET0131 , \P2_reg3_reg[27]/NET0131 , \P2_reg3_reg[28]/NET0131 , \P2_reg3_reg[2]/NET0131 , \P2_reg3_reg[3]/NET0131 , \P2_reg3_reg[4]/NET0131 , \P2_reg3_reg[5]/NET0131 , \P2_reg3_reg[6]/NET0131 , \P2_reg3_reg[7]/NET0131 , \P2_reg3_reg[8]/NET0131 , \P2_reg3_reg[9]/NET0131 , \P2_wr_reg/NET0131 , \si[0]_pad , \si[10]_pad , \si[11]_pad , \si[12]_pad , \si[13]_pad , \si[14]_pad , \si[15]_pad , \si[16]_pad , \si[17]_pad , \si[18]_pad , \si[19]_pad , \si[1]_pad , \si[20]_pad , \si[21]_pad , \si[22]_pad , \si[23]_pad , \si[24]_pad , \si[25]_pad , \si[26]_pad , \si[27]_pad , \si[28]_pad , \si[29]_pad , \si[2]_pad , \si[30]_pad , \si[31]_pad , \si[3]_pad , \si[4]_pad , \si[5]_pad , \si[6]_pad , \si[7]_pad , \si[8]_pad , \si[9]_pad , \P1_state_reg[0]/NET0131_syn_2 , \_al_n0 , \_al_n1 , \g73521/_0_ , \g73537/_0_ , \g73538/_0_ , \g73539/_0_ , \g73540/_0_ , \g73570/_0_ , \g73571/_0_ , \g73572/_0_ , \g73573/_0_ , \g73574/_0_ , \g73575/_0_ , \g73576/_0_ , \g73577/_0_ , \g73578/_0_ , \g73579/_0_ , \g73609/_0_ , \g73610/_0_ , \g73611/_0_ , \g73613/_0_ , \g73614/_0_ , \g73615/_0_ , \g73617/_0_ , \g73618/_0_ , \g73619/_0_ , \g73620/_0_ , \g73621/_0_ , \g73622/_0_ , \g73623/_0_ , \g73624/_0_ , \g73625/_0_ , \g73626/_0_ , \g73627/_0_ , \g73628/_0_ , \g73629/_0_ , \g73630/_0_ , \g73631/_0_ , \g73632/_0_ , \g73633/_0_ , \g73692/_0_ , \g73693/_0_ , \g73694/_0_ , \g73696/_0_ , \g73697/_0_ , \g73703/_0_ , \g73704/_0_ , \g73709/_0_ , \g73710/_0_ , \g73711/_0_ , \g73712/_0_ , \g73713/_0_ , \g73714/_0_ , \g73715/_0_ , \g73716/_0_ , \g73717/_0_ , \g73718/_0_ , \g73719/_0_ , \g73720/_0_ , \g73774/_0_ , \g73775/_0_ , \g73776/_0_ , \g73777/_0_ , \g73806/_0_ , \g73807/_0_ , \g73808/_0_ , \g73809/_0_ , \g73810/_0_ , \g73811/_0_ , \g73812/_0_ , \g73813/_0_ , \g73814/_0_ , \g73815/_0_ , \g73816/_0_ , \g73817/_0_ , \g73818/_0_ , \g73819/_0_ , \g73820/_0_ , \g73821/_0_ , \g73822/_0_ , \g73823/_0_ , \g73824/_0_ , \g73825/_0_ , \g73826/_0_ , \g73827/_0_ , \g73828/_0_ , \g73829/_0_ , \g73830/_0_ , \g73831/_0_ , \g73832/_0_ , \g73833/_0_ , \g73834/_0_ , \g73835/_0_ , \g73836/_0_ , \g73908/_0_ , \g73909/_0_ , \g73911/_0_ , \g73912/_0_ , \g73915/_0_ , \g73916/_0_ , \g73946/_0_ , \g73950/_0_ , \g73957/_0_ , \g73958/_0_ , \g73959/_0_ , \g73960/_0_ , \g73961/_0_ , \g73962/_0_ , \g73963/_0_ , \g73964/_0_ , \g73965/_0_ , \g73966/_0_ , \g73968/_0_ , \g73969/_0_ , \g73970/_0_ , \g73971/_0_ , \g73972/_0_ , \g73973/_0_ , \g73974/_0_ , \g73975/_0_ , \g73976/_0_ , \g73977/_0_ , \g73978/_0_ , \g73979/_0_ , \g73980/_0_ , \g73981/_0_ , \g73982/_0_ , \g73983/_0_ , \g73984/_0_ , \g73985/_0_ , \g74044/_0_ , \g74045/_0_ , \g74046/_0_ , \g74047/_0_ , \g74048/_0_ , \g74049/_0_ , \g74051/_0_ , \g74052/_0_ , \g74099/_0_ , \g74100/_0_ , \g74101/_0_ , \g74102/_0_ , \g74103/_0_ , \g74104/_0_ , \g74105/_0_ , \g74106/_0_ , \g74107/_0_ , \g74108/_0_ , \g74109/_0_ , \g74110/_0_ , \g74111/_0_ , \g74112/_0_ , \g74113/_0_ , \g74114/_0_ , \g74115/_0_ , \g74116/_0_ , \g74117/_0_ , \g74118/_0_ , \g74119/_0_ , \g74120/_0_ , \g74121/_0_ , \g74122/_0_ , \g74199/_0_ , \g74200/_0_ , \g74201/_0_ , \g74202/_0_ , \g74279/_0_ , \g74280/_0_ , \g74284/_0_ , \g74285/_0_ , \g74287/_0_ , \g74288/_0_ , \g74289/_0_ , \g74290/_0_ , \g74291/_0_ , \g74292/_0_ , \g74293/_0_ , \g74294/_0_ , \g74295/_0_ , \g74296/_0_ , \g74298/_0_ , \g74299/_0_ , \g74300/_0_ , \g74301/_0_ , \g74302/_0_ , \g74382/_0_ , \g74383/_0_ , \g74384/_0_ , \g74385/_0_ , \g74386/_0_ , \g74387/_0_ , \g74456/_0_ , \g74457/_0_ , \g74458/_0_ , \g74459/_0_ , \g74460/_0_ , \g74461/_0_ , \g74462/_0_ , \g74463/_0_ , \g74464/_0_ , \g74465/_0_ , \g74466/_0_ , \g74467/_0_ , \g74468/_0_ , \g74469/_0_ , \g74470/_0_ , \g74471/_0_ , \g74661/_0_ , \g74662/_0_ , \g74663/_0_ , \g74664/_0_ , \g74665/_0_ , \g74666/_0_ , \g74667/_0_ , \g74668/_0_ , \g74669/_0_ , \g74670/_0_ , \g74671/_0_ , \g74672/_0_ , \g74673/_0_ , \g74674/_0_ , \g74899/_0_ , \g74900/_0_ , \g74901/_0_ , \g74902/_0_ , \g75002/_0_ , \g75005/_0_ , \g75191/_0_ , \g75192/_0_ , \g75193/_0_ , \g75194/_0_ , \g75195/_0_ , \g75392/_0_ , \g75399/_0_ , \g75606/_0_ , \g75607/_0_ , \g75608/_0_ , \g75609/_0_ , \g75610/_0_ , \g76007/_0_ , \g76008/_0_ , \g76685/_0_ , \g76696/_0_ , \g77574/_0_ , \g77575/_0_ , \g77576/_0_ , \g77577/_0_ , \g77578/_0_ , \g77579/_0_ , \g82699/_3_ , \g82700/_3_ , \g82701/_3_ , \g82702/_3_ , \g82703/_3_ , \g82704/_3_ , \g83319/_0_ , \g83320/_0_ , \g83321/_0_ , \g83322/_0_ , \g83323/_3_ , \g83324/_0_ , \g83325/_0_ , \g83326/_0_ , \g83327/_0_ , \g83328/_0_ , \g83329/_0_ , \g83330/_0_ , \g83331/_0_ , \g83332/_0_ , \g83333/_0_ , \g83334/_0_ , \g83335/_0_ , \g83336/_3_ , \g83337/_0_ , \g83338/_0_ , \g83339/_0_ , \g83340/_0_ , \g83341/_0_ , \g83342/_0_ , \g83343/_0_ , \g83344/_0_ , \g83345/_0_ , \g83347/_3_ , \g83348/_3_ , \g83349/_3_ , \g83350/_3_ , \g83351/_3_ , \g83352/_3_ , \g83353/_3_ , \g83354/_3_ , \g83355/_3_ , \g83356/_3_ , \g83357/_0_ , \g83358/_3_ , \g83359/_3_ , \g83360/_3_ , \g83361/_3_ , \g83362/_3_ , \g83363/_3_ , \g83364/_3_ , \g83365/_0_ , \g83366/_3_ , \g83367/_0_ , \g83368/_3_ , \g83369/_3_ , \g83370/_0_ , \g83371/_3_ , \g83372/_3_ , \g83373/_3_ , \g83374/_3_ , \g83376/_0_ , \g83778/_0_ , \g83784/_0_ , \g84388/_0_ , \g84389/_0_ , \g84391/_0_ , \g84395/_0_ , \g84397/_0_ , \g84398/_0_ , \g84399/_0_ , \g84400/_0_ , \g84401/_0_ , \g84402/_0_ , \g84403/_0_ , \g84405/_0_ , \g84406/_0_ , \g84407/_0_ , \g84408/_0_ , \g84409/_0_ , \g84410/_0_ , \g84411/_0_ , \g84412/_0_ , \g84413/_0_ , \g84414/_0_ , \g84415/_0_ , \g84416/_0_ , \g84417/_0_ , \g84418/_0_ , \g84419/_0_ , \g84420/_0_ , \g84421/_0_ , \g84422/_0_ , \g84423/_0_ , \g84424/_0_ , \g84425/_0_ , \g84426/_0_ , \g84427/_0_ , \g84429/_0_ , \g84430/_0_ , \g84442/_0_ , \g84443/_0_ , \g84444/_0_ , \g84445/_0_ , \g84908/_0_ , \g84961/_0_ , \g84984/u3_syn_4 , \g84985/u3_syn_4 , \g85802/_0_ , \g86055/_1_ , \g86073/_0_ , \g86298/u3_syn_4 , \g86300/u3_syn_4 , \g87397/_0_ , \g87409/_0_ , \g87480/_0_ , \g87494/_0_ , \g87544/_0_ , \g87555/_0_ , \g87567/_0_ , \g87576/_0_ , \g87894/_0_ , \g87905/_0_ , \g87914/_0_ , \g87955/_1_ , \g88030/_0_ , \g88039/_0_ , \g88054/_0_ , \g88079/_0_ , \g88094/_0_ , \g88111/_0_ , \g88122/_0_ , \g88129/_0_ , \g88162/_0_ , \g88185/_0_ , \g88196/_0_ , \g88204/_0_ , \g88220/_0_ , \g88226/_0_ , \g88243/_0_ , \g88252/_0_ , \g88261/_0_ , \g88269/_0_ , \g88288/_0_ , \g88299/_0_ , \g88310/_0_ , \g88321/_0_ , \g88328/_0_ , \g88335/_0_ , \g88356/_0_ , \g88366/_0_ , \g88372/_0_ , \g88380/_0_ , \g88395_dup/_0_ , \g88403/_0_ , \g88414/_0_ , \g88425/_0_ , \g88443/_0_ , \g88453/_0_ , \g88471/_0_ , \g88524/_0_ , \g88546/_0_ , \g88556/_0_ , \g88563/_0_ , \g89966/_1_ , \g89999/_1_ , \g95209/_0_ , \g95269/_0_ , \g95319/_0_ , \g95354/_0_ , \g95786/_0_ , \g95909/_0_ , \g95914/_0_ , \g95918/_0_ , \g95984/_0_ , \g96009/_0_ , \g96124/_0_ , \g96218/_0_ , \g96286/_0_ , \g96335/_0_ , \g96465/_0_ , \g96694/_0_ , \g96713/_0_ , \g96830/_0_ , \g96875/_0_ , rd_pad, \so[0]_pad , \so[10]_pad , \so[11]_pad , \so[12]_pad , \so[13]_pad , \so[14]_pad , \so[15]_pad , \so[16]_pad , \so[17]_pad , \so[18]_pad , \so[19]_pad , \so[1]_pad , \so[2]_pad , \so[3]_pad , \so[4]_pad , \so[5]_pad , \so[6]_pad , \so[7]_pad , \so[8]_pad , \so[9]_pad , wr_pad);
	input \P1_B_reg/NET0131  ;
	input \P1_IR_reg[0]/NET0131  ;
	input \P1_IR_reg[10]/NET0131  ;
	input \P1_IR_reg[11]/NET0131  ;
	input \P1_IR_reg[12]/NET0131  ;
	input \P1_IR_reg[13]/NET0131  ;
	input \P1_IR_reg[14]/NET0131  ;
	input \P1_IR_reg[15]/NET0131  ;
	input \P1_IR_reg[16]/NET0131  ;
	input \P1_IR_reg[17]/NET0131  ;
	input \P1_IR_reg[18]/NET0131  ;
	input \P1_IR_reg[19]/NET0131  ;
	input \P1_IR_reg[1]/NET0131  ;
	input \P1_IR_reg[20]/NET0131  ;
	input \P1_IR_reg[21]/NET0131  ;
	input \P1_IR_reg[22]/NET0131  ;
	input \P1_IR_reg[23]/NET0131  ;
	input \P1_IR_reg[24]/NET0131  ;
	input \P1_IR_reg[25]/NET0131  ;
	input \P1_IR_reg[26]/NET0131  ;
	input \P1_IR_reg[27]/NET0131  ;
	input \P1_IR_reg[28]/NET0131  ;
	input \P1_IR_reg[29]/NET0131  ;
	input \P1_IR_reg[2]/NET0131  ;
	input \P1_IR_reg[30]/NET0131  ;
	input \P1_IR_reg[31]/NET0131  ;
	input \P1_IR_reg[3]/NET0131  ;
	input \P1_IR_reg[4]/NET0131  ;
	input \P1_IR_reg[5]/NET0131  ;
	input \P1_IR_reg[6]/NET0131  ;
	input \P1_IR_reg[7]/NET0131  ;
	input \P1_IR_reg[8]/NET0131  ;
	input \P1_IR_reg[9]/NET0131  ;
	input \P1_addr_reg[0]/NET0131  ;
	input \P1_addr_reg[10]/NET0131  ;
	input \P1_addr_reg[11]/NET0131  ;
	input \P1_addr_reg[12]/NET0131  ;
	input \P1_addr_reg[13]/NET0131  ;
	input \P1_addr_reg[14]/NET0131  ;
	input \P1_addr_reg[15]/NET0131  ;
	input \P1_addr_reg[16]/NET0131  ;
	input \P1_addr_reg[17]/NET0131  ;
	input \P1_addr_reg[18]/NET0131  ;
	input \P1_addr_reg[19]/NET0131  ;
	input \P1_addr_reg[1]/NET0131  ;
	input \P1_addr_reg[2]/NET0131  ;
	input \P1_addr_reg[3]/NET0131  ;
	input \P1_addr_reg[4]/NET0131  ;
	input \P1_addr_reg[5]/NET0131  ;
	input \P1_addr_reg[6]/NET0131  ;
	input \P1_addr_reg[7]/NET0131  ;
	input \P1_addr_reg[8]/NET0131  ;
	input \P1_addr_reg[9]/NET0131  ;
	input \P1_d_reg[0]/NET0131  ;
	input \P1_d_reg[1]/NET0131  ;
	input \P1_datao_reg[0]/NET0131  ;
	input \P1_datao_reg[10]/NET0131  ;
	input \P1_datao_reg[11]/NET0131  ;
	input \P1_datao_reg[12]/NET0131  ;
	input \P1_datao_reg[13]/NET0131  ;
	input \P1_datao_reg[14]/NET0131  ;
	input \P1_datao_reg[15]/NET0131  ;
	input \P1_datao_reg[16]/NET0131  ;
	input \P1_datao_reg[17]/NET0131  ;
	input \P1_datao_reg[18]/NET0131  ;
	input \P1_datao_reg[19]/NET0131  ;
	input \P1_datao_reg[1]/NET0131  ;
	input \P1_datao_reg[20]/NET0131  ;
	input \P1_datao_reg[21]/NET0131  ;
	input \P1_datao_reg[22]/NET0131  ;
	input \P1_datao_reg[23]/NET0131  ;
	input \P1_datao_reg[24]/NET0131  ;
	input \P1_datao_reg[25]/NET0131  ;
	input \P1_datao_reg[26]/NET0131  ;
	input \P1_datao_reg[27]/NET0131  ;
	input \P1_datao_reg[28]/NET0131  ;
	input \P1_datao_reg[29]/NET0131  ;
	input \P1_datao_reg[2]/NET0131  ;
	input \P1_datao_reg[30]/NET0131  ;
	input \P1_datao_reg[31]/NET0131  ;
	input \P1_datao_reg[3]/NET0131  ;
	input \P1_datao_reg[4]/NET0131  ;
	input \P1_datao_reg[5]/NET0131  ;
	input \P1_datao_reg[6]/NET0131  ;
	input \P1_datao_reg[7]/NET0131  ;
	input \P1_datao_reg[8]/NET0131  ;
	input \P1_datao_reg[9]/NET0131  ;
	input \P1_rd_reg/NET0131  ;
	input \P1_reg0_reg[0]/NET0131  ;
	input \P1_reg0_reg[10]/NET0131  ;
	input \P1_reg0_reg[11]/NET0131  ;
	input \P1_reg0_reg[12]/NET0131  ;
	input \P1_reg0_reg[13]/NET0131  ;
	input \P1_reg0_reg[14]/NET0131  ;
	input \P1_reg0_reg[15]/NET0131  ;
	input \P1_reg0_reg[16]/NET0131  ;
	input \P1_reg0_reg[17]/NET0131  ;
	input \P1_reg0_reg[18]/NET0131  ;
	input \P1_reg0_reg[19]/NET0131  ;
	input \P1_reg0_reg[1]/NET0131  ;
	input \P1_reg0_reg[20]/NET0131  ;
	input \P1_reg0_reg[21]/NET0131  ;
	input \P1_reg0_reg[22]/NET0131  ;
	input \P1_reg0_reg[23]/NET0131  ;
	input \P1_reg0_reg[24]/NET0131  ;
	input \P1_reg0_reg[25]/NET0131  ;
	input \P1_reg0_reg[26]/NET0131  ;
	input \P1_reg0_reg[27]/NET0131  ;
	input \P1_reg0_reg[28]/NET0131  ;
	input \P1_reg0_reg[29]/NET0131  ;
	input \P1_reg0_reg[2]/NET0131  ;
	input \P1_reg0_reg[30]/NET0131  ;
	input \P1_reg0_reg[31]/NET0131  ;
	input \P1_reg0_reg[3]/NET0131  ;
	input \P1_reg0_reg[4]/NET0131  ;
	input \P1_reg0_reg[5]/NET0131  ;
	input \P1_reg0_reg[6]/NET0131  ;
	input \P1_reg0_reg[7]/NET0131  ;
	input \P1_reg0_reg[8]/NET0131  ;
	input \P1_reg0_reg[9]/NET0131  ;
	input \P1_reg1_reg[0]/NET0131  ;
	input \P1_reg1_reg[10]/NET0131  ;
	input \P1_reg1_reg[11]/NET0131  ;
	input \P1_reg1_reg[12]/NET0131  ;
	input \P1_reg1_reg[13]/NET0131  ;
	input \P1_reg1_reg[14]/NET0131  ;
	input \P1_reg1_reg[15]/NET0131  ;
	input \P1_reg1_reg[16]/NET0131  ;
	input \P1_reg1_reg[17]/NET0131  ;
	input \P1_reg1_reg[18]/NET0131  ;
	input \P1_reg1_reg[19]/NET0131  ;
	input \P1_reg1_reg[1]/NET0131  ;
	input \P1_reg1_reg[20]/NET0131  ;
	input \P1_reg1_reg[21]/NET0131  ;
	input \P1_reg1_reg[22]/NET0131  ;
	input \P1_reg1_reg[23]/NET0131  ;
	input \P1_reg1_reg[24]/NET0131  ;
	input \P1_reg1_reg[25]/NET0131  ;
	input \P1_reg1_reg[26]/NET0131  ;
	input \P1_reg1_reg[27]/NET0131  ;
	input \P1_reg1_reg[28]/NET0131  ;
	input \P1_reg1_reg[29]/NET0131  ;
	input \P1_reg1_reg[2]/NET0131  ;
	input \P1_reg1_reg[30]/NET0131  ;
	input \P1_reg1_reg[31]/NET0131  ;
	input \P1_reg1_reg[3]/NET0131  ;
	input \P1_reg1_reg[4]/NET0131  ;
	input \P1_reg1_reg[5]/NET0131  ;
	input \P1_reg1_reg[6]/NET0131  ;
	input \P1_reg1_reg[7]/NET0131  ;
	input \P1_reg1_reg[8]/NET0131  ;
	input \P1_reg1_reg[9]/NET0131  ;
	input \P1_reg2_reg[0]/NET0131  ;
	input \P1_reg2_reg[10]/NET0131  ;
	input \P1_reg2_reg[11]/NET0131  ;
	input \P1_reg2_reg[12]/NET0131  ;
	input \P1_reg2_reg[13]/NET0131  ;
	input \P1_reg2_reg[14]/NET0131  ;
	input \P1_reg2_reg[15]/NET0131  ;
	input \P1_reg2_reg[16]/NET0131  ;
	input \P1_reg2_reg[17]/NET0131  ;
	input \P1_reg2_reg[18]/NET0131  ;
	input \P1_reg2_reg[19]/NET0131  ;
	input \P1_reg2_reg[1]/NET0131  ;
	input \P1_reg2_reg[20]/NET0131  ;
	input \P1_reg2_reg[21]/NET0131  ;
	input \P1_reg2_reg[22]/NET0131  ;
	input \P1_reg2_reg[23]/NET0131  ;
	input \P1_reg2_reg[24]/NET0131  ;
	input \P1_reg2_reg[25]/NET0131  ;
	input \P1_reg2_reg[26]/NET0131  ;
	input \P1_reg2_reg[27]/NET0131  ;
	input \P1_reg2_reg[28]/NET0131  ;
	input \P1_reg2_reg[29]/NET0131  ;
	input \P1_reg2_reg[2]/NET0131  ;
	input \P1_reg2_reg[30]/NET0131  ;
	input \P1_reg2_reg[31]/NET0131  ;
	input \P1_reg2_reg[3]/NET0131  ;
	input \P1_reg2_reg[4]/NET0131  ;
	input \P1_reg2_reg[5]/NET0131  ;
	input \P1_reg2_reg[6]/NET0131  ;
	input \P1_reg2_reg[7]/NET0131  ;
	input \P1_reg2_reg[8]/NET0131  ;
	input \P1_reg2_reg[9]/NET0131  ;
	input \P1_reg3_reg[0]/NET0131  ;
	input \P1_reg3_reg[10]/NET0131  ;
	input \P1_reg3_reg[11]/NET0131  ;
	input \P1_reg3_reg[12]/NET0131  ;
	input \P1_reg3_reg[13]/NET0131  ;
	input \P1_reg3_reg[14]/NET0131  ;
	input \P1_reg3_reg[15]/NET0131  ;
	input \P1_reg3_reg[16]/NET0131  ;
	input \P1_reg3_reg[17]/NET0131  ;
	input \P1_reg3_reg[18]/NET0131  ;
	input \P1_reg3_reg[19]/NET0131  ;
	input \P1_reg3_reg[1]/NET0131  ;
	input \P1_reg3_reg[20]/NET0131  ;
	input \P1_reg3_reg[21]/NET0131  ;
	input \P1_reg3_reg[22]/NET0131  ;
	input \P1_reg3_reg[23]/NET0131  ;
	input \P1_reg3_reg[24]/NET0131  ;
	input \P1_reg3_reg[25]/NET0131  ;
	input \P1_reg3_reg[26]/NET0131  ;
	input \P1_reg3_reg[27]/NET0131  ;
	input \P1_reg3_reg[28]/NET0131  ;
	input \P1_reg3_reg[2]/NET0131  ;
	input \P1_reg3_reg[3]/NET0131  ;
	input \P1_reg3_reg[4]/NET0131  ;
	input \P1_reg3_reg[5]/NET0131  ;
	input \P1_reg3_reg[6]/NET0131  ;
	input \P1_reg3_reg[7]/NET0131  ;
	input \P1_reg3_reg[8]/NET0131  ;
	input \P1_reg3_reg[9]/NET0131  ;
	input \P1_state_reg[0]/NET0131  ;
	input \P1_wr_reg/NET0131  ;
	input \P2_B_reg/NET0131  ;
	input \P2_IR_reg[0]/NET0131  ;
	input \P2_IR_reg[10]/NET0131  ;
	input \P2_IR_reg[11]/NET0131  ;
	input \P2_IR_reg[12]/NET0131  ;
	input \P2_IR_reg[13]/NET0131  ;
	input \P2_IR_reg[14]/NET0131  ;
	input \P2_IR_reg[15]/NET0131  ;
	input \P2_IR_reg[16]/NET0131  ;
	input \P2_IR_reg[17]/NET0131  ;
	input \P2_IR_reg[18]/NET0131  ;
	input \P2_IR_reg[19]/NET0131  ;
	input \P2_IR_reg[1]/NET0131  ;
	input \P2_IR_reg[20]/NET0131  ;
	input \P2_IR_reg[21]/NET0131  ;
	input \P2_IR_reg[22]/NET0131  ;
	input \P2_IR_reg[23]/NET0131  ;
	input \P2_IR_reg[24]/NET0131  ;
	input \P2_IR_reg[25]/NET0131  ;
	input \P2_IR_reg[26]/NET0131  ;
	input \P2_IR_reg[27]/NET0131  ;
	input \P2_IR_reg[28]/NET0131  ;
	input \P2_IR_reg[29]/NET0131  ;
	input \P2_IR_reg[2]/NET0131  ;
	input \P2_IR_reg[30]/NET0131  ;
	input \P2_IR_reg[31]/NET0131  ;
	input \P2_IR_reg[3]/NET0131  ;
	input \P2_IR_reg[4]/NET0131  ;
	input \P2_IR_reg[5]/NET0131  ;
	input \P2_IR_reg[6]/NET0131  ;
	input \P2_IR_reg[7]/NET0131  ;
	input \P2_IR_reg[8]/NET0131  ;
	input \P2_IR_reg[9]/NET0131  ;
	input \P2_addr_reg[0]/NET0131  ;
	input \P2_addr_reg[10]/NET0131  ;
	input \P2_addr_reg[11]/NET0131  ;
	input \P2_addr_reg[12]/NET0131  ;
	input \P2_addr_reg[13]/NET0131  ;
	input \P2_addr_reg[14]/NET0131  ;
	input \P2_addr_reg[15]/NET0131  ;
	input \P2_addr_reg[16]/NET0131  ;
	input \P2_addr_reg[17]/NET0131  ;
	input \P2_addr_reg[18]/NET0131  ;
	input \P2_addr_reg[19]/NET0131  ;
	input \P2_addr_reg[1]/NET0131  ;
	input \P2_addr_reg[2]/NET0131  ;
	input \P2_addr_reg[3]/NET0131  ;
	input \P2_addr_reg[4]/NET0131  ;
	input \P2_addr_reg[5]/NET0131  ;
	input \P2_addr_reg[6]/NET0131  ;
	input \P2_addr_reg[7]/NET0131  ;
	input \P2_addr_reg[8]/NET0131  ;
	input \P2_addr_reg[9]/NET0131  ;
	input \P2_d_reg[0]/NET0131  ;
	input \P2_d_reg[1]/NET0131  ;
	input \P2_datao_reg[0]/NET0131  ;
	input \P2_datao_reg[10]/NET0131  ;
	input \P2_datao_reg[11]/NET0131  ;
	input \P2_datao_reg[12]/NET0131  ;
	input \P2_datao_reg[13]/NET0131  ;
	input \P2_datao_reg[14]/NET0131  ;
	input \P2_datao_reg[15]/NET0131  ;
	input \P2_datao_reg[16]/NET0131  ;
	input \P2_datao_reg[17]/NET0131  ;
	input \P2_datao_reg[18]/NET0131  ;
	input \P2_datao_reg[19]/NET0131  ;
	input \P2_datao_reg[1]/NET0131  ;
	input \P2_datao_reg[20]/NET0131  ;
	input \P2_datao_reg[21]/NET0131  ;
	input \P2_datao_reg[22]/NET0131  ;
	input \P2_datao_reg[23]/NET0131  ;
	input \P2_datao_reg[24]/NET0131  ;
	input \P2_datao_reg[25]/NET0131  ;
	input \P2_datao_reg[26]/NET0131  ;
	input \P2_datao_reg[27]/NET0131  ;
	input \P2_datao_reg[28]/NET0131  ;
	input \P2_datao_reg[29]/NET0131  ;
	input \P2_datao_reg[2]/NET0131  ;
	input \P2_datao_reg[30]/NET0131  ;
	input \P2_datao_reg[31]/NET0131  ;
	input \P2_datao_reg[3]/NET0131  ;
	input \P2_datao_reg[4]/NET0131  ;
	input \P2_datao_reg[5]/NET0131  ;
	input \P2_datao_reg[6]/NET0131  ;
	input \P2_datao_reg[7]/NET0131  ;
	input \P2_datao_reg[8]/NET0131  ;
	input \P2_datao_reg[9]/NET0131  ;
	input \P2_rd_reg/NET0131  ;
	input \P2_reg0_reg[0]/NET0131  ;
	input \P2_reg0_reg[10]/NET0131  ;
	input \P2_reg0_reg[11]/NET0131  ;
	input \P2_reg0_reg[12]/NET0131  ;
	input \P2_reg0_reg[13]/NET0131  ;
	input \P2_reg0_reg[14]/NET0131  ;
	input \P2_reg0_reg[15]/NET0131  ;
	input \P2_reg0_reg[16]/NET0131  ;
	input \P2_reg0_reg[17]/NET0131  ;
	input \P2_reg0_reg[18]/NET0131  ;
	input \P2_reg0_reg[19]/NET0131  ;
	input \P2_reg0_reg[1]/NET0131  ;
	input \P2_reg0_reg[20]/NET0131  ;
	input \P2_reg0_reg[21]/NET0131  ;
	input \P2_reg0_reg[22]/NET0131  ;
	input \P2_reg0_reg[23]/NET0131  ;
	input \P2_reg0_reg[24]/NET0131  ;
	input \P2_reg0_reg[25]/NET0131  ;
	input \P2_reg0_reg[26]/NET0131  ;
	input \P2_reg0_reg[27]/NET0131  ;
	input \P2_reg0_reg[28]/NET0131  ;
	input \P2_reg0_reg[29]/NET0131  ;
	input \P2_reg0_reg[2]/NET0131  ;
	input \P2_reg0_reg[30]/NET0131  ;
	input \P2_reg0_reg[31]/NET0131  ;
	input \P2_reg0_reg[3]/NET0131  ;
	input \P2_reg0_reg[4]/NET0131  ;
	input \P2_reg0_reg[5]/NET0131  ;
	input \P2_reg0_reg[6]/NET0131  ;
	input \P2_reg0_reg[7]/NET0131  ;
	input \P2_reg0_reg[8]/NET0131  ;
	input \P2_reg0_reg[9]/NET0131  ;
	input \P2_reg1_reg[0]/NET0131  ;
	input \P2_reg1_reg[10]/NET0131  ;
	input \P2_reg1_reg[11]/NET0131  ;
	input \P2_reg1_reg[12]/NET0131  ;
	input \P2_reg1_reg[13]/NET0131  ;
	input \P2_reg1_reg[14]/NET0131  ;
	input \P2_reg1_reg[15]/NET0131  ;
	input \P2_reg1_reg[16]/NET0131  ;
	input \P2_reg1_reg[17]/NET0131  ;
	input \P2_reg1_reg[18]/NET0131  ;
	input \P2_reg1_reg[19]/NET0131  ;
	input \P2_reg1_reg[1]/NET0131  ;
	input \P2_reg1_reg[20]/NET0131  ;
	input \P2_reg1_reg[21]/NET0131  ;
	input \P2_reg1_reg[22]/NET0131  ;
	input \P2_reg1_reg[23]/NET0131  ;
	input \P2_reg1_reg[24]/NET0131  ;
	input \P2_reg1_reg[25]/NET0131  ;
	input \P2_reg1_reg[26]/NET0131  ;
	input \P2_reg1_reg[27]/NET0131  ;
	input \P2_reg1_reg[28]/NET0131  ;
	input \P2_reg1_reg[29]/NET0131  ;
	input \P2_reg1_reg[2]/NET0131  ;
	input \P2_reg1_reg[30]/NET0131  ;
	input \P2_reg1_reg[31]/NET0131  ;
	input \P2_reg1_reg[3]/NET0131  ;
	input \P2_reg1_reg[4]/NET0131  ;
	input \P2_reg1_reg[5]/NET0131  ;
	input \P2_reg1_reg[6]/NET0131  ;
	input \P2_reg1_reg[7]/NET0131  ;
	input \P2_reg1_reg[8]/NET0131  ;
	input \P2_reg1_reg[9]/NET0131  ;
	input \P2_reg2_reg[0]/NET0131  ;
	input \P2_reg2_reg[10]/NET0131  ;
	input \P2_reg2_reg[11]/NET0131  ;
	input \P2_reg2_reg[12]/NET0131  ;
	input \P2_reg2_reg[13]/NET0131  ;
	input \P2_reg2_reg[14]/NET0131  ;
	input \P2_reg2_reg[15]/NET0131  ;
	input \P2_reg2_reg[16]/NET0131  ;
	input \P2_reg2_reg[17]/NET0131  ;
	input \P2_reg2_reg[18]/NET0131  ;
	input \P2_reg2_reg[19]/NET0131  ;
	input \P2_reg2_reg[1]/NET0131  ;
	input \P2_reg2_reg[20]/NET0131  ;
	input \P2_reg2_reg[21]/NET0131  ;
	input \P2_reg2_reg[22]/NET0131  ;
	input \P2_reg2_reg[23]/NET0131  ;
	input \P2_reg2_reg[24]/NET0131  ;
	input \P2_reg2_reg[25]/NET0131  ;
	input \P2_reg2_reg[26]/NET0131  ;
	input \P2_reg2_reg[27]/NET0131  ;
	input \P2_reg2_reg[28]/NET0131  ;
	input \P2_reg2_reg[29]/NET0131  ;
	input \P2_reg2_reg[2]/NET0131  ;
	input \P2_reg2_reg[30]/NET0131  ;
	input \P2_reg2_reg[31]/NET0131  ;
	input \P2_reg2_reg[3]/NET0131  ;
	input \P2_reg2_reg[4]/NET0131  ;
	input \P2_reg2_reg[5]/NET0131  ;
	input \P2_reg2_reg[6]/NET0131  ;
	input \P2_reg2_reg[7]/NET0131  ;
	input \P2_reg2_reg[8]/NET0131  ;
	input \P2_reg2_reg[9]/NET0131  ;
	input \P2_reg3_reg[0]/NET0131  ;
	input \P2_reg3_reg[10]/NET0131  ;
	input \P2_reg3_reg[11]/NET0131  ;
	input \P2_reg3_reg[12]/NET0131  ;
	input \P2_reg3_reg[13]/NET0131  ;
	input \P2_reg3_reg[14]/NET0131  ;
	input \P2_reg3_reg[15]/NET0131  ;
	input \P2_reg3_reg[16]/NET0131  ;
	input \P2_reg3_reg[17]/NET0131  ;
	input \P2_reg3_reg[18]/NET0131  ;
	input \P2_reg3_reg[19]/NET0131  ;
	input \P2_reg3_reg[1]/NET0131  ;
	input \P2_reg3_reg[20]/NET0131  ;
	input \P2_reg3_reg[21]/NET0131  ;
	input \P2_reg3_reg[22]/NET0131  ;
	input \P2_reg3_reg[23]/NET0131  ;
	input \P2_reg3_reg[24]/NET0131  ;
	input \P2_reg3_reg[25]/NET0131  ;
	input \P2_reg3_reg[26]/NET0131  ;
	input \P2_reg3_reg[27]/NET0131  ;
	input \P2_reg3_reg[28]/NET0131  ;
	input \P2_reg3_reg[2]/NET0131  ;
	input \P2_reg3_reg[3]/NET0131  ;
	input \P2_reg3_reg[4]/NET0131  ;
	input \P2_reg3_reg[5]/NET0131  ;
	input \P2_reg3_reg[6]/NET0131  ;
	input \P2_reg3_reg[7]/NET0131  ;
	input \P2_reg3_reg[8]/NET0131  ;
	input \P2_reg3_reg[9]/NET0131  ;
	input \P2_wr_reg/NET0131  ;
	input \si[0]_pad  ;
	input \si[10]_pad  ;
	input \si[11]_pad  ;
	input \si[12]_pad  ;
	input \si[13]_pad  ;
	input \si[14]_pad  ;
	input \si[15]_pad  ;
	input \si[16]_pad  ;
	input \si[17]_pad  ;
	input \si[18]_pad  ;
	input \si[19]_pad  ;
	input \si[1]_pad  ;
	input \si[20]_pad  ;
	input \si[21]_pad  ;
	input \si[22]_pad  ;
	input \si[23]_pad  ;
	input \si[24]_pad  ;
	input \si[25]_pad  ;
	input \si[26]_pad  ;
	input \si[27]_pad  ;
	input \si[28]_pad  ;
	input \si[29]_pad  ;
	input \si[2]_pad  ;
	input \si[30]_pad  ;
	input \si[31]_pad  ;
	input \si[3]_pad  ;
	input \si[4]_pad  ;
	input \si[5]_pad  ;
	input \si[6]_pad  ;
	input \si[7]_pad  ;
	input \si[8]_pad  ;
	input \si[9]_pad  ;
	output \P1_state_reg[0]/NET0131_syn_2  ;
	output \_al_n0  ;
	output \_al_n1  ;
	output \g73521/_0_  ;
	output \g73537/_0_  ;
	output \g73538/_0_  ;
	output \g73539/_0_  ;
	output \g73540/_0_  ;
	output \g73570/_0_  ;
	output \g73571/_0_  ;
	output \g73572/_0_  ;
	output \g73573/_0_  ;
	output \g73574/_0_  ;
	output \g73575/_0_  ;
	output \g73576/_0_  ;
	output \g73577/_0_  ;
	output \g73578/_0_  ;
	output \g73579/_0_  ;
	output \g73609/_0_  ;
	output \g73610/_0_  ;
	output \g73611/_0_  ;
	output \g73613/_0_  ;
	output \g73614/_0_  ;
	output \g73615/_0_  ;
	output \g73617/_0_  ;
	output \g73618/_0_  ;
	output \g73619/_0_  ;
	output \g73620/_0_  ;
	output \g73621/_0_  ;
	output \g73622/_0_  ;
	output \g73623/_0_  ;
	output \g73624/_0_  ;
	output \g73625/_0_  ;
	output \g73626/_0_  ;
	output \g73627/_0_  ;
	output \g73628/_0_  ;
	output \g73629/_0_  ;
	output \g73630/_0_  ;
	output \g73631/_0_  ;
	output \g73632/_0_  ;
	output \g73633/_0_  ;
	output \g73692/_0_  ;
	output \g73693/_0_  ;
	output \g73694/_0_  ;
	output \g73696/_0_  ;
	output \g73697/_0_  ;
	output \g73703/_0_  ;
	output \g73704/_0_  ;
	output \g73709/_0_  ;
	output \g73710/_0_  ;
	output \g73711/_0_  ;
	output \g73712/_0_  ;
	output \g73713/_0_  ;
	output \g73714/_0_  ;
	output \g73715/_0_  ;
	output \g73716/_0_  ;
	output \g73717/_0_  ;
	output \g73718/_0_  ;
	output \g73719/_0_  ;
	output \g73720/_0_  ;
	output \g73774/_0_  ;
	output \g73775/_0_  ;
	output \g73776/_0_  ;
	output \g73777/_0_  ;
	output \g73806/_0_  ;
	output \g73807/_0_  ;
	output \g73808/_0_  ;
	output \g73809/_0_  ;
	output \g73810/_0_  ;
	output \g73811/_0_  ;
	output \g73812/_0_  ;
	output \g73813/_0_  ;
	output \g73814/_0_  ;
	output \g73815/_0_  ;
	output \g73816/_0_  ;
	output \g73817/_0_  ;
	output \g73818/_0_  ;
	output \g73819/_0_  ;
	output \g73820/_0_  ;
	output \g73821/_0_  ;
	output \g73822/_0_  ;
	output \g73823/_0_  ;
	output \g73824/_0_  ;
	output \g73825/_0_  ;
	output \g73826/_0_  ;
	output \g73827/_0_  ;
	output \g73828/_0_  ;
	output \g73829/_0_  ;
	output \g73830/_0_  ;
	output \g73831/_0_  ;
	output \g73832/_0_  ;
	output \g73833/_0_  ;
	output \g73834/_0_  ;
	output \g73835/_0_  ;
	output \g73836/_0_  ;
	output \g73908/_0_  ;
	output \g73909/_0_  ;
	output \g73911/_0_  ;
	output \g73912/_0_  ;
	output \g73915/_0_  ;
	output \g73916/_0_  ;
	output \g73946/_0_  ;
	output \g73950/_0_  ;
	output \g73957/_0_  ;
	output \g73958/_0_  ;
	output \g73959/_0_  ;
	output \g73960/_0_  ;
	output \g73961/_0_  ;
	output \g73962/_0_  ;
	output \g73963/_0_  ;
	output \g73964/_0_  ;
	output \g73965/_0_  ;
	output \g73966/_0_  ;
	output \g73968/_0_  ;
	output \g73969/_0_  ;
	output \g73970/_0_  ;
	output \g73971/_0_  ;
	output \g73972/_0_  ;
	output \g73973/_0_  ;
	output \g73974/_0_  ;
	output \g73975/_0_  ;
	output \g73976/_0_  ;
	output \g73977/_0_  ;
	output \g73978/_0_  ;
	output \g73979/_0_  ;
	output \g73980/_0_  ;
	output \g73981/_0_  ;
	output \g73982/_0_  ;
	output \g73983/_0_  ;
	output \g73984/_0_  ;
	output \g73985/_0_  ;
	output \g74044/_0_  ;
	output \g74045/_0_  ;
	output \g74046/_0_  ;
	output \g74047/_0_  ;
	output \g74048/_0_  ;
	output \g74049/_0_  ;
	output \g74051/_0_  ;
	output \g74052/_0_  ;
	output \g74099/_0_  ;
	output \g74100/_0_  ;
	output \g74101/_0_  ;
	output \g74102/_0_  ;
	output \g74103/_0_  ;
	output \g74104/_0_  ;
	output \g74105/_0_  ;
	output \g74106/_0_  ;
	output \g74107/_0_  ;
	output \g74108/_0_  ;
	output \g74109/_0_  ;
	output \g74110/_0_  ;
	output \g74111/_0_  ;
	output \g74112/_0_  ;
	output \g74113/_0_  ;
	output \g74114/_0_  ;
	output \g74115/_0_  ;
	output \g74116/_0_  ;
	output \g74117/_0_  ;
	output \g74118/_0_  ;
	output \g74119/_0_  ;
	output \g74120/_0_  ;
	output \g74121/_0_  ;
	output \g74122/_0_  ;
	output \g74199/_0_  ;
	output \g74200/_0_  ;
	output \g74201/_0_  ;
	output \g74202/_0_  ;
	output \g74279/_0_  ;
	output \g74280/_0_  ;
	output \g74284/_0_  ;
	output \g74285/_0_  ;
	output \g74287/_0_  ;
	output \g74288/_0_  ;
	output \g74289/_0_  ;
	output \g74290/_0_  ;
	output \g74291/_0_  ;
	output \g74292/_0_  ;
	output \g74293/_0_  ;
	output \g74294/_0_  ;
	output \g74295/_0_  ;
	output \g74296/_0_  ;
	output \g74298/_0_  ;
	output \g74299/_0_  ;
	output \g74300/_0_  ;
	output \g74301/_0_  ;
	output \g74302/_0_  ;
	output \g74382/_0_  ;
	output \g74383/_0_  ;
	output \g74384/_0_  ;
	output \g74385/_0_  ;
	output \g74386/_0_  ;
	output \g74387/_0_  ;
	output \g74456/_0_  ;
	output \g74457/_0_  ;
	output \g74458/_0_  ;
	output \g74459/_0_  ;
	output \g74460/_0_  ;
	output \g74461/_0_  ;
	output \g74462/_0_  ;
	output \g74463/_0_  ;
	output \g74464/_0_  ;
	output \g74465/_0_  ;
	output \g74466/_0_  ;
	output \g74467/_0_  ;
	output \g74468/_0_  ;
	output \g74469/_0_  ;
	output \g74470/_0_  ;
	output \g74471/_0_  ;
	output \g74661/_0_  ;
	output \g74662/_0_  ;
	output \g74663/_0_  ;
	output \g74664/_0_  ;
	output \g74665/_0_  ;
	output \g74666/_0_  ;
	output \g74667/_0_  ;
	output \g74668/_0_  ;
	output \g74669/_0_  ;
	output \g74670/_0_  ;
	output \g74671/_0_  ;
	output \g74672/_0_  ;
	output \g74673/_0_  ;
	output \g74674/_0_  ;
	output \g74899/_0_  ;
	output \g74900/_0_  ;
	output \g74901/_0_  ;
	output \g74902/_0_  ;
	output \g75002/_0_  ;
	output \g75005/_0_  ;
	output \g75191/_0_  ;
	output \g75192/_0_  ;
	output \g75193/_0_  ;
	output \g75194/_0_  ;
	output \g75195/_0_  ;
	output \g75392/_0_  ;
	output \g75399/_0_  ;
	output \g75606/_0_  ;
	output \g75607/_0_  ;
	output \g75608/_0_  ;
	output \g75609/_0_  ;
	output \g75610/_0_  ;
	output \g76007/_0_  ;
	output \g76008/_0_  ;
	output \g76685/_0_  ;
	output \g76696/_0_  ;
	output \g77574/_0_  ;
	output \g77575/_0_  ;
	output \g77576/_0_  ;
	output \g77577/_0_  ;
	output \g77578/_0_  ;
	output \g77579/_0_  ;
	output \g82699/_3_  ;
	output \g82700/_3_  ;
	output \g82701/_3_  ;
	output \g82702/_3_  ;
	output \g82703/_3_  ;
	output \g82704/_3_  ;
	output \g83319/_0_  ;
	output \g83320/_0_  ;
	output \g83321/_0_  ;
	output \g83322/_0_  ;
	output \g83323/_3_  ;
	output \g83324/_0_  ;
	output \g83325/_0_  ;
	output \g83326/_0_  ;
	output \g83327/_0_  ;
	output \g83328/_0_  ;
	output \g83329/_0_  ;
	output \g83330/_0_  ;
	output \g83331/_0_  ;
	output \g83332/_0_  ;
	output \g83333/_0_  ;
	output \g83334/_0_  ;
	output \g83335/_0_  ;
	output \g83336/_3_  ;
	output \g83337/_0_  ;
	output \g83338/_0_  ;
	output \g83339/_0_  ;
	output \g83340/_0_  ;
	output \g83341/_0_  ;
	output \g83342/_0_  ;
	output \g83343/_0_  ;
	output \g83344/_0_  ;
	output \g83345/_0_  ;
	output \g83347/_3_  ;
	output \g83348/_3_  ;
	output \g83349/_3_  ;
	output \g83350/_3_  ;
	output \g83351/_3_  ;
	output \g83352/_3_  ;
	output \g83353/_3_  ;
	output \g83354/_3_  ;
	output \g83355/_3_  ;
	output \g83356/_3_  ;
	output \g83357/_0_  ;
	output \g83358/_3_  ;
	output \g83359/_3_  ;
	output \g83360/_3_  ;
	output \g83361/_3_  ;
	output \g83362/_3_  ;
	output \g83363/_3_  ;
	output \g83364/_3_  ;
	output \g83365/_0_  ;
	output \g83366/_3_  ;
	output \g83367/_0_  ;
	output \g83368/_3_  ;
	output \g83369/_3_  ;
	output \g83370/_0_  ;
	output \g83371/_3_  ;
	output \g83372/_3_  ;
	output \g83373/_3_  ;
	output \g83374/_3_  ;
	output \g83376/_0_  ;
	output \g83778/_0_  ;
	output \g83784/_0_  ;
	output \g84388/_0_  ;
	output \g84389/_0_  ;
	output \g84391/_0_  ;
	output \g84395/_0_  ;
	output \g84397/_0_  ;
	output \g84398/_0_  ;
	output \g84399/_0_  ;
	output \g84400/_0_  ;
	output \g84401/_0_  ;
	output \g84402/_0_  ;
	output \g84403/_0_  ;
	output \g84405/_0_  ;
	output \g84406/_0_  ;
	output \g84407/_0_  ;
	output \g84408/_0_  ;
	output \g84409/_0_  ;
	output \g84410/_0_  ;
	output \g84411/_0_  ;
	output \g84412/_0_  ;
	output \g84413/_0_  ;
	output \g84414/_0_  ;
	output \g84415/_0_  ;
	output \g84416/_0_  ;
	output \g84417/_0_  ;
	output \g84418/_0_  ;
	output \g84419/_0_  ;
	output \g84420/_0_  ;
	output \g84421/_0_  ;
	output \g84422/_0_  ;
	output \g84423/_0_  ;
	output \g84424/_0_  ;
	output \g84425/_0_  ;
	output \g84426/_0_  ;
	output \g84427/_0_  ;
	output \g84429/_0_  ;
	output \g84430/_0_  ;
	output \g84442/_0_  ;
	output \g84443/_0_  ;
	output \g84444/_0_  ;
	output \g84445/_0_  ;
	output \g84908/_0_  ;
	output \g84961/_0_  ;
	output \g84984/u3_syn_4  ;
	output \g84985/u3_syn_4  ;
	output \g85802/_0_  ;
	output \g86055/_1_  ;
	output \g86073/_0_  ;
	output \g86298/u3_syn_4  ;
	output \g86300/u3_syn_4  ;
	output \g87397/_0_  ;
	output \g87409/_0_  ;
	output \g87480/_0_  ;
	output \g87494/_0_  ;
	output \g87544/_0_  ;
	output \g87555/_0_  ;
	output \g87567/_0_  ;
	output \g87576/_0_  ;
	output \g87894/_0_  ;
	output \g87905/_0_  ;
	output \g87914/_0_  ;
	output \g87955/_1_  ;
	output \g88030/_0_  ;
	output \g88039/_0_  ;
	output \g88054/_0_  ;
	output \g88079/_0_  ;
	output \g88094/_0_  ;
	output \g88111/_0_  ;
	output \g88122/_0_  ;
	output \g88129/_0_  ;
	output \g88162/_0_  ;
	output \g88185/_0_  ;
	output \g88196/_0_  ;
	output \g88204/_0_  ;
	output \g88220/_0_  ;
	output \g88226/_0_  ;
	output \g88243/_0_  ;
	output \g88252/_0_  ;
	output \g88261/_0_  ;
	output \g88269/_0_  ;
	output \g88288/_0_  ;
	output \g88299/_0_  ;
	output \g88310/_0_  ;
	output \g88321/_0_  ;
	output \g88328/_0_  ;
	output \g88335/_0_  ;
	output \g88356/_0_  ;
	output \g88366/_0_  ;
	output \g88372/_0_  ;
	output \g88380/_0_  ;
	output \g88395_dup/_0_  ;
	output \g88403/_0_  ;
	output \g88414/_0_  ;
	output \g88425/_0_  ;
	output \g88443/_0_  ;
	output \g88453/_0_  ;
	output \g88471/_0_  ;
	output \g88524/_0_  ;
	output \g88546/_0_  ;
	output \g88556/_0_  ;
	output \g88563/_0_  ;
	output \g89966/_1_  ;
	output \g89999/_1_  ;
	output \g95209/_0_  ;
	output \g95269/_0_  ;
	output \g95319/_0_  ;
	output \g95354/_0_  ;
	output \g95786/_0_  ;
	output \g95909/_0_  ;
	output \g95914/_0_  ;
	output \g95918/_0_  ;
	output \g95984/_0_  ;
	output \g96009/_0_  ;
	output \g96124/_0_  ;
	output \g96218/_0_  ;
	output \g96286/_0_  ;
	output \g96335/_0_  ;
	output \g96465/_0_  ;
	output \g96694/_0_  ;
	output \g96713/_0_  ;
	output \g96830/_0_  ;
	output \g96875/_0_  ;
	output rd_pad ;
	output \so[0]_pad  ;
	output \so[10]_pad  ;
	output \so[11]_pad  ;
	output \so[12]_pad  ;
	output \so[13]_pad  ;
	output \so[14]_pad  ;
	output \so[15]_pad  ;
	output \so[16]_pad  ;
	output \so[17]_pad  ;
	output \so[18]_pad  ;
	output \so[19]_pad  ;
	output \so[1]_pad  ;
	output \so[2]_pad  ;
	output \so[3]_pad  ;
	output \so[4]_pad  ;
	output \so[5]_pad  ;
	output \so[6]_pad  ;
	output \so[7]_pad  ;
	output \so[8]_pad  ;
	output \so[9]_pad  ;
	output wr_pad ;
	wire _w12829_ ;
	wire _w12828_ ;
	wire _w12827_ ;
	wire _w12826_ ;
	wire _w12825_ ;
	wire _w12824_ ;
	wire _w12823_ ;
	wire _w12822_ ;
	wire _w12821_ ;
	wire _w12820_ ;
	wire _w12819_ ;
	wire _w12818_ ;
	wire _w12817_ ;
	wire _w12816_ ;
	wire _w12815_ ;
	wire _w12814_ ;
	wire _w12813_ ;
	wire _w12812_ ;
	wire _w12811_ ;
	wire _w12810_ ;
	wire _w12809_ ;
	wire _w12808_ ;
	wire _w12807_ ;
	wire _w12806_ ;
	wire _w12805_ ;
	wire _w12804_ ;
	wire _w12803_ ;
	wire _w12802_ ;
	wire _w12801_ ;
	wire _w12800_ ;
	wire _w12799_ ;
	wire _w12798_ ;
	wire _w12797_ ;
	wire _w12796_ ;
	wire _w12795_ ;
	wire _w12794_ ;
	wire _w12793_ ;
	wire _w12792_ ;
	wire _w12791_ ;
	wire _w12790_ ;
	wire _w12789_ ;
	wire _w12788_ ;
	wire _w12787_ ;
	wire _w12786_ ;
	wire _w12785_ ;
	wire _w12784_ ;
	wire _w12783_ ;
	wire _w12782_ ;
	wire _w12781_ ;
	wire _w12780_ ;
	wire _w12779_ ;
	wire _w12778_ ;
	wire _w12777_ ;
	wire _w12776_ ;
	wire _w12775_ ;
	wire _w12774_ ;
	wire _w12773_ ;
	wire _w12772_ ;
	wire _w12771_ ;
	wire _w12770_ ;
	wire _w12769_ ;
	wire _w12768_ ;
	wire _w12767_ ;
	wire _w12766_ ;
	wire _w12765_ ;
	wire _w12764_ ;
	wire _w12763_ ;
	wire _w12762_ ;
	wire _w12761_ ;
	wire _w12760_ ;
	wire _w12759_ ;
	wire _w12758_ ;
	wire _w12757_ ;
	wire _w12756_ ;
	wire _w12755_ ;
	wire _w12754_ ;
	wire _w12753_ ;
	wire _w12752_ ;
	wire _w12751_ ;
	wire _w12750_ ;
	wire _w12749_ ;
	wire _w12748_ ;
	wire _w12747_ ;
	wire _w12746_ ;
	wire _w12745_ ;
	wire _w12744_ ;
	wire _w12743_ ;
	wire _w12742_ ;
	wire _w12741_ ;
	wire _w12740_ ;
	wire _w12739_ ;
	wire _w12738_ ;
	wire _w12737_ ;
	wire _w12736_ ;
	wire _w12735_ ;
	wire _w12734_ ;
	wire _w12733_ ;
	wire _w12732_ ;
	wire _w12731_ ;
	wire _w12730_ ;
	wire _w12729_ ;
	wire _w12728_ ;
	wire _w12727_ ;
	wire _w12726_ ;
	wire _w12725_ ;
	wire _w12724_ ;
	wire _w12723_ ;
	wire _w12722_ ;
	wire _w12721_ ;
	wire _w12720_ ;
	wire _w12719_ ;
	wire _w12718_ ;
	wire _w12717_ ;
	wire _w12716_ ;
	wire _w12715_ ;
	wire _w12714_ ;
	wire _w12713_ ;
	wire _w12712_ ;
	wire _w12711_ ;
	wire _w12710_ ;
	wire _w12709_ ;
	wire _w12708_ ;
	wire _w12707_ ;
	wire _w12706_ ;
	wire _w12705_ ;
	wire _w12704_ ;
	wire _w12703_ ;
	wire _w12702_ ;
	wire _w12701_ ;
	wire _w12700_ ;
	wire _w12699_ ;
	wire _w12698_ ;
	wire _w12697_ ;
	wire _w12696_ ;
	wire _w12695_ ;
	wire _w12694_ ;
	wire _w12693_ ;
	wire _w12692_ ;
	wire _w12691_ ;
	wire _w12690_ ;
	wire _w12689_ ;
	wire _w12688_ ;
	wire _w12687_ ;
	wire _w12686_ ;
	wire _w12685_ ;
	wire _w12684_ ;
	wire _w12683_ ;
	wire _w12682_ ;
	wire _w12681_ ;
	wire _w12680_ ;
	wire _w12679_ ;
	wire _w12678_ ;
	wire _w12677_ ;
	wire _w12676_ ;
	wire _w12675_ ;
	wire _w12674_ ;
	wire _w12673_ ;
	wire _w12672_ ;
	wire _w12671_ ;
	wire _w12670_ ;
	wire _w12669_ ;
	wire _w12668_ ;
	wire _w12667_ ;
	wire _w12666_ ;
	wire _w12665_ ;
	wire _w12664_ ;
	wire _w12663_ ;
	wire _w12662_ ;
	wire _w12661_ ;
	wire _w12660_ ;
	wire _w12659_ ;
	wire _w12658_ ;
	wire _w12657_ ;
	wire _w12656_ ;
	wire _w12655_ ;
	wire _w12654_ ;
	wire _w12653_ ;
	wire _w12652_ ;
	wire _w12651_ ;
	wire _w12650_ ;
	wire _w12649_ ;
	wire _w12648_ ;
	wire _w12647_ ;
	wire _w12646_ ;
	wire _w12645_ ;
	wire _w12644_ ;
	wire _w12643_ ;
	wire _w12642_ ;
	wire _w12641_ ;
	wire _w12640_ ;
	wire _w12639_ ;
	wire _w12638_ ;
	wire _w12637_ ;
	wire _w12636_ ;
	wire _w12635_ ;
	wire _w12634_ ;
	wire _w12633_ ;
	wire _w12632_ ;
	wire _w12631_ ;
	wire _w12630_ ;
	wire _w12629_ ;
	wire _w12628_ ;
	wire _w12627_ ;
	wire _w12626_ ;
	wire _w12625_ ;
	wire _w12624_ ;
	wire _w12623_ ;
	wire _w12622_ ;
	wire _w12621_ ;
	wire _w12620_ ;
	wire _w12619_ ;
	wire _w12618_ ;
	wire _w12617_ ;
	wire _w12616_ ;
	wire _w12615_ ;
	wire _w12614_ ;
	wire _w12613_ ;
	wire _w12612_ ;
	wire _w12611_ ;
	wire _w12610_ ;
	wire _w12609_ ;
	wire _w12608_ ;
	wire _w12607_ ;
	wire _w12606_ ;
	wire _w12605_ ;
	wire _w12604_ ;
	wire _w12603_ ;
	wire _w12602_ ;
	wire _w12601_ ;
	wire _w12600_ ;
	wire _w12599_ ;
	wire _w12598_ ;
	wire _w12597_ ;
	wire _w12596_ ;
	wire _w12595_ ;
	wire _w12594_ ;
	wire _w12593_ ;
	wire _w12592_ ;
	wire _w12591_ ;
	wire _w12590_ ;
	wire _w12589_ ;
	wire _w12588_ ;
	wire _w12587_ ;
	wire _w12586_ ;
	wire _w12585_ ;
	wire _w12584_ ;
	wire _w12583_ ;
	wire _w12582_ ;
	wire _w12581_ ;
	wire _w12580_ ;
	wire _w12579_ ;
	wire _w12578_ ;
	wire _w12577_ ;
	wire _w12576_ ;
	wire _w12575_ ;
	wire _w12574_ ;
	wire _w12573_ ;
	wire _w12572_ ;
	wire _w12571_ ;
	wire _w12570_ ;
	wire _w12569_ ;
	wire _w12568_ ;
	wire _w12567_ ;
	wire _w12566_ ;
	wire _w12565_ ;
	wire _w12564_ ;
	wire _w12563_ ;
	wire _w12562_ ;
	wire _w12561_ ;
	wire _w12560_ ;
	wire _w12559_ ;
	wire _w12558_ ;
	wire _w12557_ ;
	wire _w12556_ ;
	wire _w12555_ ;
	wire _w12554_ ;
	wire _w12553_ ;
	wire _w12552_ ;
	wire _w12551_ ;
	wire _w12550_ ;
	wire _w12549_ ;
	wire _w12548_ ;
	wire _w12547_ ;
	wire _w12546_ ;
	wire _w12545_ ;
	wire _w12544_ ;
	wire _w12543_ ;
	wire _w12542_ ;
	wire _w12541_ ;
	wire _w12540_ ;
	wire _w12539_ ;
	wire _w12538_ ;
	wire _w12537_ ;
	wire _w12536_ ;
	wire _w12535_ ;
	wire _w12534_ ;
	wire _w12533_ ;
	wire _w12532_ ;
	wire _w12531_ ;
	wire _w12530_ ;
	wire _w12529_ ;
	wire _w12528_ ;
	wire _w12527_ ;
	wire _w12526_ ;
	wire _w12525_ ;
	wire _w12524_ ;
	wire _w12523_ ;
	wire _w12522_ ;
	wire _w12521_ ;
	wire _w12520_ ;
	wire _w12519_ ;
	wire _w12518_ ;
	wire _w12517_ ;
	wire _w12516_ ;
	wire _w12515_ ;
	wire _w12514_ ;
	wire _w12513_ ;
	wire _w12512_ ;
	wire _w12511_ ;
	wire _w12510_ ;
	wire _w12509_ ;
	wire _w12508_ ;
	wire _w12507_ ;
	wire _w12506_ ;
	wire _w12505_ ;
	wire _w12504_ ;
	wire _w12503_ ;
	wire _w12502_ ;
	wire _w12501_ ;
	wire _w12500_ ;
	wire _w12499_ ;
	wire _w12498_ ;
	wire _w12497_ ;
	wire _w12496_ ;
	wire _w12495_ ;
	wire _w12494_ ;
	wire _w12493_ ;
	wire _w12492_ ;
	wire _w12491_ ;
	wire _w12490_ ;
	wire _w12489_ ;
	wire _w12488_ ;
	wire _w12487_ ;
	wire _w12486_ ;
	wire _w12485_ ;
	wire _w12484_ ;
	wire _w12483_ ;
	wire _w12482_ ;
	wire _w12481_ ;
	wire _w12480_ ;
	wire _w12479_ ;
	wire _w12478_ ;
	wire _w12477_ ;
	wire _w12476_ ;
	wire _w12475_ ;
	wire _w12474_ ;
	wire _w12473_ ;
	wire _w12472_ ;
	wire _w12471_ ;
	wire _w12470_ ;
	wire _w12469_ ;
	wire _w12468_ ;
	wire _w12467_ ;
	wire _w12466_ ;
	wire _w12465_ ;
	wire _w12464_ ;
	wire _w12463_ ;
	wire _w12462_ ;
	wire _w12461_ ;
	wire _w12460_ ;
	wire _w12459_ ;
	wire _w12458_ ;
	wire _w12457_ ;
	wire _w12456_ ;
	wire _w12455_ ;
	wire _w12454_ ;
	wire _w12453_ ;
	wire _w12452_ ;
	wire _w12451_ ;
	wire _w12450_ ;
	wire _w12449_ ;
	wire _w12448_ ;
	wire _w12447_ ;
	wire _w12446_ ;
	wire _w12445_ ;
	wire _w12444_ ;
	wire _w12443_ ;
	wire _w12442_ ;
	wire _w12441_ ;
	wire _w12440_ ;
	wire _w12439_ ;
	wire _w12438_ ;
	wire _w12437_ ;
	wire _w12436_ ;
	wire _w12435_ ;
	wire _w12434_ ;
	wire _w12433_ ;
	wire _w12432_ ;
	wire _w12431_ ;
	wire _w12430_ ;
	wire _w12429_ ;
	wire _w12428_ ;
	wire _w12427_ ;
	wire _w12426_ ;
	wire _w12425_ ;
	wire _w12424_ ;
	wire _w12423_ ;
	wire _w12422_ ;
	wire _w12421_ ;
	wire _w12420_ ;
	wire _w12419_ ;
	wire _w12418_ ;
	wire _w12417_ ;
	wire _w12416_ ;
	wire _w12415_ ;
	wire _w12414_ ;
	wire _w12413_ ;
	wire _w12412_ ;
	wire _w12411_ ;
	wire _w12410_ ;
	wire _w12409_ ;
	wire _w12408_ ;
	wire _w12407_ ;
	wire _w12406_ ;
	wire _w12405_ ;
	wire _w12404_ ;
	wire _w12403_ ;
	wire _w12402_ ;
	wire _w12401_ ;
	wire _w12400_ ;
	wire _w12399_ ;
	wire _w12398_ ;
	wire _w12397_ ;
	wire _w12396_ ;
	wire _w12395_ ;
	wire _w12394_ ;
	wire _w12393_ ;
	wire _w12392_ ;
	wire _w12391_ ;
	wire _w12390_ ;
	wire _w12389_ ;
	wire _w12388_ ;
	wire _w12387_ ;
	wire _w12386_ ;
	wire _w12385_ ;
	wire _w12384_ ;
	wire _w12383_ ;
	wire _w12382_ ;
	wire _w12381_ ;
	wire _w12380_ ;
	wire _w12379_ ;
	wire _w12378_ ;
	wire _w12377_ ;
	wire _w12376_ ;
	wire _w12375_ ;
	wire _w12374_ ;
	wire _w12373_ ;
	wire _w12372_ ;
	wire _w12371_ ;
	wire _w12370_ ;
	wire _w12369_ ;
	wire _w12368_ ;
	wire _w12367_ ;
	wire _w12366_ ;
	wire _w12365_ ;
	wire _w12364_ ;
	wire _w12363_ ;
	wire _w12362_ ;
	wire _w12361_ ;
	wire _w12360_ ;
	wire _w12359_ ;
	wire _w12358_ ;
	wire _w12357_ ;
	wire _w12356_ ;
	wire _w12355_ ;
	wire _w12354_ ;
	wire _w12353_ ;
	wire _w12352_ ;
	wire _w12351_ ;
	wire _w12350_ ;
	wire _w12349_ ;
	wire _w12348_ ;
	wire _w12347_ ;
	wire _w12346_ ;
	wire _w12345_ ;
	wire _w12344_ ;
	wire _w12343_ ;
	wire _w12342_ ;
	wire _w12341_ ;
	wire _w12340_ ;
	wire _w12339_ ;
	wire _w12338_ ;
	wire _w12337_ ;
	wire _w12336_ ;
	wire _w12335_ ;
	wire _w12334_ ;
	wire _w12333_ ;
	wire _w12332_ ;
	wire _w12331_ ;
	wire _w12330_ ;
	wire _w12329_ ;
	wire _w12328_ ;
	wire _w12327_ ;
	wire _w12326_ ;
	wire _w12325_ ;
	wire _w12324_ ;
	wire _w12323_ ;
	wire _w12322_ ;
	wire _w12321_ ;
	wire _w12320_ ;
	wire _w12319_ ;
	wire _w12318_ ;
	wire _w12317_ ;
	wire _w12316_ ;
	wire _w12315_ ;
	wire _w12314_ ;
	wire _w12313_ ;
	wire _w12312_ ;
	wire _w12311_ ;
	wire _w12310_ ;
	wire _w12309_ ;
	wire _w12308_ ;
	wire _w12307_ ;
	wire _w12306_ ;
	wire _w12305_ ;
	wire _w12304_ ;
	wire _w12303_ ;
	wire _w12302_ ;
	wire _w12301_ ;
	wire _w12300_ ;
	wire _w12299_ ;
	wire _w12298_ ;
	wire _w12297_ ;
	wire _w12296_ ;
	wire _w12295_ ;
	wire _w12294_ ;
	wire _w12293_ ;
	wire _w12292_ ;
	wire _w12291_ ;
	wire _w12290_ ;
	wire _w12289_ ;
	wire _w12288_ ;
	wire _w12287_ ;
	wire _w12286_ ;
	wire _w12285_ ;
	wire _w12284_ ;
	wire _w12283_ ;
	wire _w12282_ ;
	wire _w12281_ ;
	wire _w12280_ ;
	wire _w12279_ ;
	wire _w12278_ ;
	wire _w12277_ ;
	wire _w12276_ ;
	wire _w12275_ ;
	wire _w12274_ ;
	wire _w12273_ ;
	wire _w12272_ ;
	wire _w12271_ ;
	wire _w12270_ ;
	wire _w12269_ ;
	wire _w12268_ ;
	wire _w12267_ ;
	wire _w12266_ ;
	wire _w12265_ ;
	wire _w12264_ ;
	wire _w12263_ ;
	wire _w12262_ ;
	wire _w12261_ ;
	wire _w12260_ ;
	wire _w12259_ ;
	wire _w12258_ ;
	wire _w12257_ ;
	wire _w12256_ ;
	wire _w12255_ ;
	wire _w12254_ ;
	wire _w12253_ ;
	wire _w12252_ ;
	wire _w12251_ ;
	wire _w12250_ ;
	wire _w12249_ ;
	wire _w12248_ ;
	wire _w12247_ ;
	wire _w12246_ ;
	wire _w12245_ ;
	wire _w12244_ ;
	wire _w12243_ ;
	wire _w12242_ ;
	wire _w12241_ ;
	wire _w12240_ ;
	wire _w12239_ ;
	wire _w12238_ ;
	wire _w12237_ ;
	wire _w12236_ ;
	wire _w12235_ ;
	wire _w12234_ ;
	wire _w12233_ ;
	wire _w12232_ ;
	wire _w12231_ ;
	wire _w12230_ ;
	wire _w12229_ ;
	wire _w12228_ ;
	wire _w12227_ ;
	wire _w12226_ ;
	wire _w12225_ ;
	wire _w12224_ ;
	wire _w12223_ ;
	wire _w12222_ ;
	wire _w12221_ ;
	wire _w12220_ ;
	wire _w12219_ ;
	wire _w12218_ ;
	wire _w12217_ ;
	wire _w12216_ ;
	wire _w12215_ ;
	wire _w12214_ ;
	wire _w12213_ ;
	wire _w12212_ ;
	wire _w12211_ ;
	wire _w12210_ ;
	wire _w12209_ ;
	wire _w12208_ ;
	wire _w12207_ ;
	wire _w12206_ ;
	wire _w12205_ ;
	wire _w12204_ ;
	wire _w12203_ ;
	wire _w12202_ ;
	wire _w12201_ ;
	wire _w12200_ ;
	wire _w12199_ ;
	wire _w12198_ ;
	wire _w12197_ ;
	wire _w12196_ ;
	wire _w12195_ ;
	wire _w12194_ ;
	wire _w12193_ ;
	wire _w12192_ ;
	wire _w12191_ ;
	wire _w12190_ ;
	wire _w12189_ ;
	wire _w12188_ ;
	wire _w12187_ ;
	wire _w12186_ ;
	wire _w12185_ ;
	wire _w12184_ ;
	wire _w12183_ ;
	wire _w12182_ ;
	wire _w12181_ ;
	wire _w12180_ ;
	wire _w12179_ ;
	wire _w12178_ ;
	wire _w12177_ ;
	wire _w12176_ ;
	wire _w12175_ ;
	wire _w12174_ ;
	wire _w12173_ ;
	wire _w12172_ ;
	wire _w12171_ ;
	wire _w12170_ ;
	wire _w12169_ ;
	wire _w12168_ ;
	wire _w12167_ ;
	wire _w12166_ ;
	wire _w12165_ ;
	wire _w12164_ ;
	wire _w12163_ ;
	wire _w12162_ ;
	wire _w12161_ ;
	wire _w12160_ ;
	wire _w12159_ ;
	wire _w12158_ ;
	wire _w12157_ ;
	wire _w12156_ ;
	wire _w12155_ ;
	wire _w12154_ ;
	wire _w12153_ ;
	wire _w12152_ ;
	wire _w12151_ ;
	wire _w12150_ ;
	wire _w12149_ ;
	wire _w12148_ ;
	wire _w12147_ ;
	wire _w12146_ ;
	wire _w12145_ ;
	wire _w12144_ ;
	wire _w12143_ ;
	wire _w12142_ ;
	wire _w12141_ ;
	wire _w12140_ ;
	wire _w12139_ ;
	wire _w12138_ ;
	wire _w12137_ ;
	wire _w12136_ ;
	wire _w12135_ ;
	wire _w12134_ ;
	wire _w12133_ ;
	wire _w12132_ ;
	wire _w12131_ ;
	wire _w12130_ ;
	wire _w12129_ ;
	wire _w12128_ ;
	wire _w12127_ ;
	wire _w12126_ ;
	wire _w12125_ ;
	wire _w12124_ ;
	wire _w12123_ ;
	wire _w12122_ ;
	wire _w12121_ ;
	wire _w12120_ ;
	wire _w12119_ ;
	wire _w12118_ ;
	wire _w12117_ ;
	wire _w12116_ ;
	wire _w12115_ ;
	wire _w12114_ ;
	wire _w12113_ ;
	wire _w12112_ ;
	wire _w12111_ ;
	wire _w12110_ ;
	wire _w12109_ ;
	wire _w12108_ ;
	wire _w12107_ ;
	wire _w12106_ ;
	wire _w12105_ ;
	wire _w12104_ ;
	wire _w12103_ ;
	wire _w12102_ ;
	wire _w12101_ ;
	wire _w12100_ ;
	wire _w12099_ ;
	wire _w12098_ ;
	wire _w12097_ ;
	wire _w12096_ ;
	wire _w12095_ ;
	wire _w12094_ ;
	wire _w12093_ ;
	wire _w12092_ ;
	wire _w12091_ ;
	wire _w12090_ ;
	wire _w12089_ ;
	wire _w12088_ ;
	wire _w12087_ ;
	wire _w12086_ ;
	wire _w12085_ ;
	wire _w12084_ ;
	wire _w12083_ ;
	wire _w12082_ ;
	wire _w12081_ ;
	wire _w12080_ ;
	wire _w12079_ ;
	wire _w12078_ ;
	wire _w12077_ ;
	wire _w12076_ ;
	wire _w12075_ ;
	wire _w12074_ ;
	wire _w12073_ ;
	wire _w12072_ ;
	wire _w12071_ ;
	wire _w12070_ ;
	wire _w12069_ ;
	wire _w12068_ ;
	wire _w12067_ ;
	wire _w12066_ ;
	wire _w12065_ ;
	wire _w12064_ ;
	wire _w12063_ ;
	wire _w12062_ ;
	wire _w12061_ ;
	wire _w12060_ ;
	wire _w12059_ ;
	wire _w12058_ ;
	wire _w12057_ ;
	wire _w12056_ ;
	wire _w12055_ ;
	wire _w12054_ ;
	wire _w12053_ ;
	wire _w12052_ ;
	wire _w12051_ ;
	wire _w12050_ ;
	wire _w12049_ ;
	wire _w12048_ ;
	wire _w12047_ ;
	wire _w12046_ ;
	wire _w12045_ ;
	wire _w12044_ ;
	wire _w12043_ ;
	wire _w12042_ ;
	wire _w12041_ ;
	wire _w12040_ ;
	wire _w12039_ ;
	wire _w12038_ ;
	wire _w12037_ ;
	wire _w12036_ ;
	wire _w12035_ ;
	wire _w12034_ ;
	wire _w12033_ ;
	wire _w12032_ ;
	wire _w12031_ ;
	wire _w12030_ ;
	wire _w12029_ ;
	wire _w12028_ ;
	wire _w12027_ ;
	wire _w12026_ ;
	wire _w12025_ ;
	wire _w12024_ ;
	wire _w12023_ ;
	wire _w12022_ ;
	wire _w12021_ ;
	wire _w12020_ ;
	wire _w12019_ ;
	wire _w12018_ ;
	wire _w12017_ ;
	wire _w12016_ ;
	wire _w12015_ ;
	wire _w12014_ ;
	wire _w12013_ ;
	wire _w12012_ ;
	wire _w12011_ ;
	wire _w12010_ ;
	wire _w12009_ ;
	wire _w12008_ ;
	wire _w12007_ ;
	wire _w12006_ ;
	wire _w12005_ ;
	wire _w12004_ ;
	wire _w12003_ ;
	wire _w12002_ ;
	wire _w12001_ ;
	wire _w12000_ ;
	wire _w11999_ ;
	wire _w11998_ ;
	wire _w11997_ ;
	wire _w11996_ ;
	wire _w11995_ ;
	wire _w11994_ ;
	wire _w11993_ ;
	wire _w11992_ ;
	wire _w11991_ ;
	wire _w11990_ ;
	wire _w11989_ ;
	wire _w11988_ ;
	wire _w11987_ ;
	wire _w11986_ ;
	wire _w11985_ ;
	wire _w11984_ ;
	wire _w11983_ ;
	wire _w11982_ ;
	wire _w11981_ ;
	wire _w11980_ ;
	wire _w11979_ ;
	wire _w11978_ ;
	wire _w11977_ ;
	wire _w11976_ ;
	wire _w11975_ ;
	wire _w11974_ ;
	wire _w11973_ ;
	wire _w11972_ ;
	wire _w11971_ ;
	wire _w11970_ ;
	wire _w11969_ ;
	wire _w11968_ ;
	wire _w11967_ ;
	wire _w11966_ ;
	wire _w11965_ ;
	wire _w11964_ ;
	wire _w11963_ ;
	wire _w11962_ ;
	wire _w11961_ ;
	wire _w11960_ ;
	wire _w11959_ ;
	wire _w11958_ ;
	wire _w11957_ ;
	wire _w11956_ ;
	wire _w11955_ ;
	wire _w11954_ ;
	wire _w11953_ ;
	wire _w11952_ ;
	wire _w11951_ ;
	wire _w11950_ ;
	wire _w11949_ ;
	wire _w11948_ ;
	wire _w11947_ ;
	wire _w11946_ ;
	wire _w11945_ ;
	wire _w11944_ ;
	wire _w11943_ ;
	wire _w11942_ ;
	wire _w11941_ ;
	wire _w11940_ ;
	wire _w11939_ ;
	wire _w11938_ ;
	wire _w11937_ ;
	wire _w11936_ ;
	wire _w11935_ ;
	wire _w11934_ ;
	wire _w11933_ ;
	wire _w11932_ ;
	wire _w11931_ ;
	wire _w11930_ ;
	wire _w11929_ ;
	wire _w11928_ ;
	wire _w11927_ ;
	wire _w11926_ ;
	wire _w11925_ ;
	wire _w11924_ ;
	wire _w11923_ ;
	wire _w11922_ ;
	wire _w11921_ ;
	wire _w11920_ ;
	wire _w11919_ ;
	wire _w11918_ ;
	wire _w11917_ ;
	wire _w11916_ ;
	wire _w11915_ ;
	wire _w11914_ ;
	wire _w11913_ ;
	wire _w11912_ ;
	wire _w11911_ ;
	wire _w11910_ ;
	wire _w11909_ ;
	wire _w11908_ ;
	wire _w11907_ ;
	wire _w11906_ ;
	wire _w11905_ ;
	wire _w11904_ ;
	wire _w11903_ ;
	wire _w11902_ ;
	wire _w11901_ ;
	wire _w11900_ ;
	wire _w11899_ ;
	wire _w11898_ ;
	wire _w11897_ ;
	wire _w11896_ ;
	wire _w11895_ ;
	wire _w11894_ ;
	wire _w11893_ ;
	wire _w11892_ ;
	wire _w11891_ ;
	wire _w11890_ ;
	wire _w11889_ ;
	wire _w11888_ ;
	wire _w11887_ ;
	wire _w11886_ ;
	wire _w11885_ ;
	wire _w11884_ ;
	wire _w11883_ ;
	wire _w11882_ ;
	wire _w11881_ ;
	wire _w11880_ ;
	wire _w11879_ ;
	wire _w11878_ ;
	wire _w11877_ ;
	wire _w11876_ ;
	wire _w11875_ ;
	wire _w11874_ ;
	wire _w11873_ ;
	wire _w11872_ ;
	wire _w11871_ ;
	wire _w11870_ ;
	wire _w11869_ ;
	wire _w11868_ ;
	wire _w11867_ ;
	wire _w11866_ ;
	wire _w11865_ ;
	wire _w11864_ ;
	wire _w11863_ ;
	wire _w11862_ ;
	wire _w11861_ ;
	wire _w11860_ ;
	wire _w11859_ ;
	wire _w11858_ ;
	wire _w11857_ ;
	wire _w11856_ ;
	wire _w11855_ ;
	wire _w11854_ ;
	wire _w11853_ ;
	wire _w11852_ ;
	wire _w11851_ ;
	wire _w11850_ ;
	wire _w11849_ ;
	wire _w11848_ ;
	wire _w11847_ ;
	wire _w11846_ ;
	wire _w11845_ ;
	wire _w11844_ ;
	wire _w11843_ ;
	wire _w11842_ ;
	wire _w11841_ ;
	wire _w11840_ ;
	wire _w11839_ ;
	wire _w11838_ ;
	wire _w11837_ ;
	wire _w11836_ ;
	wire _w11835_ ;
	wire _w11834_ ;
	wire _w11833_ ;
	wire _w11832_ ;
	wire _w11831_ ;
	wire _w11830_ ;
	wire _w11829_ ;
	wire _w11828_ ;
	wire _w11827_ ;
	wire _w11826_ ;
	wire _w11825_ ;
	wire _w11824_ ;
	wire _w11823_ ;
	wire _w11822_ ;
	wire _w11821_ ;
	wire _w11820_ ;
	wire _w11819_ ;
	wire _w11818_ ;
	wire _w11817_ ;
	wire _w11816_ ;
	wire _w11815_ ;
	wire _w11814_ ;
	wire _w11813_ ;
	wire _w11812_ ;
	wire _w11811_ ;
	wire _w11810_ ;
	wire _w11809_ ;
	wire _w11808_ ;
	wire _w11807_ ;
	wire _w11806_ ;
	wire _w11805_ ;
	wire _w11804_ ;
	wire _w11803_ ;
	wire _w11802_ ;
	wire _w11801_ ;
	wire _w11800_ ;
	wire _w11799_ ;
	wire _w11798_ ;
	wire _w11797_ ;
	wire _w11796_ ;
	wire _w11795_ ;
	wire _w11794_ ;
	wire _w11793_ ;
	wire _w11792_ ;
	wire _w11791_ ;
	wire _w11790_ ;
	wire _w11789_ ;
	wire _w11788_ ;
	wire _w11787_ ;
	wire _w11786_ ;
	wire _w11785_ ;
	wire _w11784_ ;
	wire _w11783_ ;
	wire _w11782_ ;
	wire _w11781_ ;
	wire _w11780_ ;
	wire _w11779_ ;
	wire _w11778_ ;
	wire _w11777_ ;
	wire _w11776_ ;
	wire _w11775_ ;
	wire _w11774_ ;
	wire _w11773_ ;
	wire _w11772_ ;
	wire _w11771_ ;
	wire _w11770_ ;
	wire _w11769_ ;
	wire _w11768_ ;
	wire _w11767_ ;
	wire _w11766_ ;
	wire _w11765_ ;
	wire _w11764_ ;
	wire _w11763_ ;
	wire _w11762_ ;
	wire _w11761_ ;
	wire _w11760_ ;
	wire _w11759_ ;
	wire _w11758_ ;
	wire _w11757_ ;
	wire _w11756_ ;
	wire _w11755_ ;
	wire _w11754_ ;
	wire _w11753_ ;
	wire _w11752_ ;
	wire _w11751_ ;
	wire _w11750_ ;
	wire _w11749_ ;
	wire _w11748_ ;
	wire _w11747_ ;
	wire _w11746_ ;
	wire _w11745_ ;
	wire _w11744_ ;
	wire _w11743_ ;
	wire _w11742_ ;
	wire _w11741_ ;
	wire _w11740_ ;
	wire _w11739_ ;
	wire _w11738_ ;
	wire _w11737_ ;
	wire _w11736_ ;
	wire _w11735_ ;
	wire _w11734_ ;
	wire _w11733_ ;
	wire _w11732_ ;
	wire _w11731_ ;
	wire _w11730_ ;
	wire _w11729_ ;
	wire _w11728_ ;
	wire _w11727_ ;
	wire _w11726_ ;
	wire _w11725_ ;
	wire _w11724_ ;
	wire _w11723_ ;
	wire _w11722_ ;
	wire _w11721_ ;
	wire _w11720_ ;
	wire _w11719_ ;
	wire _w11718_ ;
	wire _w11717_ ;
	wire _w11716_ ;
	wire _w11715_ ;
	wire _w11714_ ;
	wire _w11713_ ;
	wire _w11712_ ;
	wire _w11711_ ;
	wire _w11710_ ;
	wire _w11709_ ;
	wire _w11708_ ;
	wire _w11707_ ;
	wire _w11706_ ;
	wire _w11705_ ;
	wire _w11704_ ;
	wire _w11703_ ;
	wire _w11702_ ;
	wire _w11701_ ;
	wire _w11700_ ;
	wire _w11699_ ;
	wire _w11698_ ;
	wire _w11697_ ;
	wire _w11696_ ;
	wire _w11695_ ;
	wire _w11694_ ;
	wire _w11693_ ;
	wire _w11692_ ;
	wire _w11691_ ;
	wire _w11690_ ;
	wire _w11689_ ;
	wire _w11688_ ;
	wire _w11687_ ;
	wire _w11686_ ;
	wire _w11685_ ;
	wire _w11684_ ;
	wire _w11683_ ;
	wire _w11682_ ;
	wire _w11681_ ;
	wire _w11680_ ;
	wire _w11679_ ;
	wire _w11678_ ;
	wire _w11677_ ;
	wire _w11676_ ;
	wire _w11675_ ;
	wire _w11674_ ;
	wire _w11673_ ;
	wire _w11672_ ;
	wire _w11671_ ;
	wire _w11670_ ;
	wire _w11669_ ;
	wire _w11668_ ;
	wire _w11667_ ;
	wire _w11666_ ;
	wire _w11665_ ;
	wire _w11664_ ;
	wire _w11663_ ;
	wire _w11662_ ;
	wire _w11661_ ;
	wire _w11660_ ;
	wire _w11659_ ;
	wire _w11658_ ;
	wire _w11657_ ;
	wire _w11656_ ;
	wire _w11655_ ;
	wire _w11654_ ;
	wire _w11653_ ;
	wire _w11652_ ;
	wire _w11651_ ;
	wire _w11650_ ;
	wire _w11649_ ;
	wire _w11648_ ;
	wire _w11647_ ;
	wire _w11646_ ;
	wire _w11645_ ;
	wire _w11644_ ;
	wire _w11643_ ;
	wire _w11642_ ;
	wire _w11641_ ;
	wire _w11640_ ;
	wire _w11639_ ;
	wire _w11638_ ;
	wire _w11637_ ;
	wire _w11636_ ;
	wire _w11635_ ;
	wire _w11634_ ;
	wire _w11633_ ;
	wire _w11632_ ;
	wire _w11631_ ;
	wire _w11630_ ;
	wire _w11629_ ;
	wire _w11628_ ;
	wire _w11627_ ;
	wire _w11626_ ;
	wire _w11625_ ;
	wire _w11624_ ;
	wire _w11623_ ;
	wire _w11622_ ;
	wire _w11621_ ;
	wire _w11620_ ;
	wire _w11619_ ;
	wire _w11618_ ;
	wire _w11617_ ;
	wire _w11616_ ;
	wire _w11615_ ;
	wire _w11614_ ;
	wire _w11613_ ;
	wire _w11612_ ;
	wire _w11611_ ;
	wire _w11610_ ;
	wire _w11609_ ;
	wire _w11608_ ;
	wire _w11607_ ;
	wire _w11606_ ;
	wire _w11605_ ;
	wire _w11604_ ;
	wire _w11603_ ;
	wire _w11602_ ;
	wire _w11601_ ;
	wire _w11600_ ;
	wire _w11599_ ;
	wire _w11598_ ;
	wire _w11597_ ;
	wire _w11596_ ;
	wire _w11595_ ;
	wire _w11594_ ;
	wire _w11593_ ;
	wire _w11592_ ;
	wire _w11591_ ;
	wire _w11590_ ;
	wire _w11589_ ;
	wire _w11588_ ;
	wire _w11587_ ;
	wire _w11586_ ;
	wire _w11585_ ;
	wire _w11584_ ;
	wire _w11583_ ;
	wire _w11582_ ;
	wire _w11581_ ;
	wire _w11580_ ;
	wire _w11579_ ;
	wire _w11578_ ;
	wire _w11577_ ;
	wire _w11576_ ;
	wire _w11575_ ;
	wire _w11574_ ;
	wire _w11573_ ;
	wire _w11572_ ;
	wire _w11571_ ;
	wire _w11570_ ;
	wire _w11569_ ;
	wire _w11568_ ;
	wire _w11567_ ;
	wire _w11566_ ;
	wire _w11565_ ;
	wire _w11564_ ;
	wire _w11563_ ;
	wire _w11562_ ;
	wire _w11561_ ;
	wire _w11560_ ;
	wire _w11559_ ;
	wire _w11558_ ;
	wire _w11557_ ;
	wire _w11556_ ;
	wire _w11555_ ;
	wire _w11554_ ;
	wire _w11553_ ;
	wire _w11552_ ;
	wire _w11551_ ;
	wire _w11550_ ;
	wire _w11549_ ;
	wire _w11548_ ;
	wire _w11547_ ;
	wire _w11546_ ;
	wire _w11545_ ;
	wire _w11544_ ;
	wire _w11543_ ;
	wire _w11542_ ;
	wire _w11541_ ;
	wire _w11540_ ;
	wire _w11539_ ;
	wire _w11538_ ;
	wire _w11537_ ;
	wire _w11536_ ;
	wire _w11535_ ;
	wire _w11534_ ;
	wire _w11533_ ;
	wire _w11532_ ;
	wire _w11531_ ;
	wire _w11530_ ;
	wire _w11529_ ;
	wire _w11528_ ;
	wire _w11527_ ;
	wire _w11526_ ;
	wire _w11525_ ;
	wire _w11524_ ;
	wire _w11523_ ;
	wire _w11522_ ;
	wire _w11521_ ;
	wire _w11520_ ;
	wire _w11519_ ;
	wire _w11518_ ;
	wire _w11517_ ;
	wire _w11516_ ;
	wire _w11515_ ;
	wire _w11514_ ;
	wire _w11513_ ;
	wire _w11512_ ;
	wire _w11511_ ;
	wire _w11510_ ;
	wire _w11509_ ;
	wire _w11508_ ;
	wire _w11507_ ;
	wire _w11506_ ;
	wire _w11505_ ;
	wire _w11504_ ;
	wire _w11503_ ;
	wire _w11502_ ;
	wire _w11501_ ;
	wire _w11500_ ;
	wire _w11499_ ;
	wire _w11498_ ;
	wire _w11497_ ;
	wire _w11496_ ;
	wire _w11495_ ;
	wire _w11494_ ;
	wire _w11493_ ;
	wire _w11492_ ;
	wire _w11491_ ;
	wire _w11490_ ;
	wire _w11489_ ;
	wire _w11488_ ;
	wire _w11487_ ;
	wire _w11486_ ;
	wire _w11485_ ;
	wire _w11484_ ;
	wire _w11483_ ;
	wire _w11482_ ;
	wire _w11481_ ;
	wire _w11480_ ;
	wire _w11479_ ;
	wire _w11478_ ;
	wire _w11477_ ;
	wire _w11476_ ;
	wire _w11475_ ;
	wire _w11474_ ;
	wire _w11473_ ;
	wire _w11472_ ;
	wire _w11471_ ;
	wire _w11470_ ;
	wire _w11469_ ;
	wire _w11468_ ;
	wire _w11467_ ;
	wire _w11466_ ;
	wire _w11465_ ;
	wire _w11464_ ;
	wire _w11463_ ;
	wire _w11462_ ;
	wire _w11461_ ;
	wire _w11460_ ;
	wire _w11459_ ;
	wire _w11458_ ;
	wire _w11457_ ;
	wire _w11456_ ;
	wire _w11455_ ;
	wire _w11454_ ;
	wire _w11453_ ;
	wire _w11452_ ;
	wire _w11451_ ;
	wire _w11450_ ;
	wire _w11449_ ;
	wire _w11448_ ;
	wire _w11447_ ;
	wire _w11446_ ;
	wire _w11445_ ;
	wire _w11444_ ;
	wire _w11443_ ;
	wire _w11442_ ;
	wire _w11441_ ;
	wire _w11440_ ;
	wire _w11439_ ;
	wire _w11438_ ;
	wire _w11437_ ;
	wire _w11436_ ;
	wire _w11435_ ;
	wire _w11434_ ;
	wire _w11433_ ;
	wire _w11432_ ;
	wire _w11431_ ;
	wire _w11430_ ;
	wire _w11429_ ;
	wire _w11428_ ;
	wire _w11427_ ;
	wire _w11426_ ;
	wire _w11425_ ;
	wire _w11424_ ;
	wire _w11423_ ;
	wire _w11422_ ;
	wire _w11421_ ;
	wire _w11420_ ;
	wire _w11419_ ;
	wire _w11418_ ;
	wire _w11417_ ;
	wire _w11416_ ;
	wire _w11415_ ;
	wire _w11414_ ;
	wire _w11413_ ;
	wire _w11412_ ;
	wire _w11411_ ;
	wire _w11410_ ;
	wire _w11409_ ;
	wire _w11408_ ;
	wire _w11407_ ;
	wire _w11406_ ;
	wire _w11405_ ;
	wire _w11404_ ;
	wire _w11403_ ;
	wire _w11402_ ;
	wire _w11401_ ;
	wire _w11400_ ;
	wire _w11399_ ;
	wire _w11398_ ;
	wire _w11397_ ;
	wire _w11396_ ;
	wire _w11395_ ;
	wire _w11394_ ;
	wire _w11393_ ;
	wire _w11392_ ;
	wire _w11391_ ;
	wire _w11390_ ;
	wire _w11389_ ;
	wire _w11388_ ;
	wire _w11387_ ;
	wire _w11386_ ;
	wire _w11385_ ;
	wire _w11384_ ;
	wire _w11383_ ;
	wire _w11382_ ;
	wire _w11381_ ;
	wire _w11380_ ;
	wire _w11379_ ;
	wire _w11378_ ;
	wire _w11377_ ;
	wire _w11376_ ;
	wire _w11375_ ;
	wire _w11374_ ;
	wire _w11373_ ;
	wire _w11372_ ;
	wire _w11371_ ;
	wire _w11370_ ;
	wire _w11369_ ;
	wire _w11368_ ;
	wire _w11367_ ;
	wire _w11366_ ;
	wire _w11365_ ;
	wire _w11364_ ;
	wire _w11363_ ;
	wire _w11362_ ;
	wire _w11361_ ;
	wire _w11360_ ;
	wire _w11359_ ;
	wire _w11358_ ;
	wire _w11357_ ;
	wire _w11356_ ;
	wire _w11355_ ;
	wire _w11354_ ;
	wire _w11353_ ;
	wire _w11352_ ;
	wire _w11351_ ;
	wire _w11350_ ;
	wire _w11349_ ;
	wire _w11348_ ;
	wire _w11347_ ;
	wire _w11346_ ;
	wire _w11345_ ;
	wire _w11344_ ;
	wire _w11343_ ;
	wire _w11342_ ;
	wire _w11341_ ;
	wire _w11340_ ;
	wire _w11339_ ;
	wire _w11338_ ;
	wire _w11337_ ;
	wire _w11336_ ;
	wire _w11335_ ;
	wire _w11334_ ;
	wire _w11333_ ;
	wire _w11332_ ;
	wire _w11331_ ;
	wire _w11330_ ;
	wire _w11329_ ;
	wire _w11328_ ;
	wire _w11327_ ;
	wire _w11326_ ;
	wire _w11325_ ;
	wire _w11324_ ;
	wire _w11323_ ;
	wire _w11322_ ;
	wire _w11321_ ;
	wire _w11320_ ;
	wire _w11319_ ;
	wire _w11318_ ;
	wire _w11317_ ;
	wire _w11316_ ;
	wire _w11315_ ;
	wire _w11314_ ;
	wire _w11313_ ;
	wire _w11312_ ;
	wire _w11311_ ;
	wire _w11310_ ;
	wire _w11309_ ;
	wire _w11308_ ;
	wire _w11307_ ;
	wire _w11306_ ;
	wire _w11305_ ;
	wire _w11304_ ;
	wire _w11303_ ;
	wire _w11302_ ;
	wire _w11301_ ;
	wire _w11300_ ;
	wire _w11299_ ;
	wire _w11298_ ;
	wire _w11297_ ;
	wire _w11296_ ;
	wire _w11295_ ;
	wire _w11294_ ;
	wire _w11293_ ;
	wire _w11292_ ;
	wire _w11291_ ;
	wire _w11290_ ;
	wire _w11289_ ;
	wire _w11288_ ;
	wire _w11287_ ;
	wire _w11286_ ;
	wire _w11285_ ;
	wire _w11284_ ;
	wire _w11283_ ;
	wire _w11282_ ;
	wire _w11281_ ;
	wire _w11280_ ;
	wire _w11279_ ;
	wire _w11278_ ;
	wire _w11277_ ;
	wire _w11276_ ;
	wire _w11275_ ;
	wire _w11274_ ;
	wire _w11273_ ;
	wire _w11272_ ;
	wire _w11271_ ;
	wire _w11270_ ;
	wire _w11269_ ;
	wire _w11268_ ;
	wire _w11267_ ;
	wire _w11266_ ;
	wire _w11265_ ;
	wire _w11264_ ;
	wire _w11263_ ;
	wire _w11262_ ;
	wire _w11261_ ;
	wire _w11260_ ;
	wire _w11259_ ;
	wire _w11258_ ;
	wire _w11257_ ;
	wire _w11256_ ;
	wire _w11255_ ;
	wire _w11254_ ;
	wire _w11253_ ;
	wire _w11252_ ;
	wire _w11251_ ;
	wire _w11250_ ;
	wire _w11249_ ;
	wire _w11248_ ;
	wire _w11247_ ;
	wire _w11246_ ;
	wire _w11245_ ;
	wire _w11244_ ;
	wire _w11243_ ;
	wire _w11242_ ;
	wire _w11241_ ;
	wire _w11240_ ;
	wire _w11239_ ;
	wire _w11238_ ;
	wire _w11237_ ;
	wire _w11236_ ;
	wire _w11235_ ;
	wire _w11234_ ;
	wire _w11233_ ;
	wire _w11232_ ;
	wire _w11231_ ;
	wire _w11230_ ;
	wire _w11229_ ;
	wire _w11228_ ;
	wire _w11227_ ;
	wire _w11226_ ;
	wire _w11225_ ;
	wire _w11224_ ;
	wire _w11223_ ;
	wire _w11222_ ;
	wire _w11221_ ;
	wire _w11220_ ;
	wire _w11219_ ;
	wire _w11218_ ;
	wire _w11217_ ;
	wire _w11216_ ;
	wire _w11215_ ;
	wire _w11214_ ;
	wire _w11213_ ;
	wire _w11212_ ;
	wire _w11211_ ;
	wire _w11210_ ;
	wire _w11209_ ;
	wire _w11208_ ;
	wire _w11207_ ;
	wire _w11206_ ;
	wire _w11205_ ;
	wire _w11204_ ;
	wire _w11203_ ;
	wire _w11202_ ;
	wire _w11201_ ;
	wire _w11200_ ;
	wire _w11199_ ;
	wire _w11198_ ;
	wire _w11197_ ;
	wire _w11196_ ;
	wire _w11195_ ;
	wire _w11194_ ;
	wire _w11193_ ;
	wire _w11192_ ;
	wire _w11191_ ;
	wire _w11190_ ;
	wire _w11189_ ;
	wire _w11188_ ;
	wire _w11187_ ;
	wire _w11186_ ;
	wire _w11185_ ;
	wire _w11184_ ;
	wire _w11183_ ;
	wire _w11182_ ;
	wire _w11181_ ;
	wire _w11180_ ;
	wire _w11179_ ;
	wire _w11178_ ;
	wire _w11177_ ;
	wire _w11176_ ;
	wire _w11175_ ;
	wire _w11174_ ;
	wire _w11173_ ;
	wire _w11172_ ;
	wire _w11171_ ;
	wire _w11170_ ;
	wire _w11169_ ;
	wire _w11168_ ;
	wire _w11167_ ;
	wire _w11166_ ;
	wire _w11165_ ;
	wire _w11164_ ;
	wire _w11163_ ;
	wire _w11162_ ;
	wire _w11161_ ;
	wire _w11160_ ;
	wire _w11159_ ;
	wire _w11158_ ;
	wire _w11157_ ;
	wire _w11156_ ;
	wire _w11155_ ;
	wire _w11154_ ;
	wire _w11153_ ;
	wire _w11152_ ;
	wire _w11151_ ;
	wire _w11150_ ;
	wire _w11149_ ;
	wire _w11148_ ;
	wire _w11147_ ;
	wire _w11146_ ;
	wire _w11145_ ;
	wire _w11144_ ;
	wire _w11143_ ;
	wire _w11142_ ;
	wire _w11141_ ;
	wire _w11140_ ;
	wire _w11139_ ;
	wire _w11138_ ;
	wire _w11137_ ;
	wire _w11136_ ;
	wire _w11135_ ;
	wire _w11134_ ;
	wire _w11133_ ;
	wire _w11132_ ;
	wire _w11131_ ;
	wire _w11130_ ;
	wire _w11129_ ;
	wire _w11128_ ;
	wire _w11127_ ;
	wire _w11126_ ;
	wire _w11125_ ;
	wire _w11124_ ;
	wire _w11123_ ;
	wire _w11122_ ;
	wire _w11121_ ;
	wire _w11120_ ;
	wire _w11119_ ;
	wire _w11118_ ;
	wire _w11117_ ;
	wire _w11116_ ;
	wire _w11115_ ;
	wire _w11114_ ;
	wire _w11113_ ;
	wire _w11112_ ;
	wire _w11111_ ;
	wire _w11110_ ;
	wire _w11109_ ;
	wire _w11108_ ;
	wire _w11107_ ;
	wire _w11106_ ;
	wire _w11105_ ;
	wire _w11104_ ;
	wire _w11103_ ;
	wire _w11102_ ;
	wire _w11101_ ;
	wire _w11100_ ;
	wire _w11099_ ;
	wire _w11098_ ;
	wire _w11097_ ;
	wire _w11096_ ;
	wire _w11095_ ;
	wire _w11094_ ;
	wire _w11093_ ;
	wire _w11092_ ;
	wire _w11091_ ;
	wire _w11090_ ;
	wire _w11089_ ;
	wire _w11088_ ;
	wire _w11087_ ;
	wire _w11086_ ;
	wire _w11085_ ;
	wire _w11084_ ;
	wire _w11083_ ;
	wire _w11082_ ;
	wire _w11081_ ;
	wire _w11080_ ;
	wire _w11079_ ;
	wire _w11078_ ;
	wire _w11077_ ;
	wire _w11076_ ;
	wire _w11075_ ;
	wire _w11074_ ;
	wire _w11073_ ;
	wire _w11072_ ;
	wire _w11071_ ;
	wire _w11070_ ;
	wire _w11069_ ;
	wire _w11068_ ;
	wire _w11067_ ;
	wire _w11066_ ;
	wire _w11065_ ;
	wire _w11064_ ;
	wire _w11063_ ;
	wire _w11062_ ;
	wire _w11061_ ;
	wire _w11060_ ;
	wire _w11059_ ;
	wire _w11058_ ;
	wire _w11057_ ;
	wire _w11056_ ;
	wire _w11055_ ;
	wire _w11054_ ;
	wire _w11053_ ;
	wire _w11052_ ;
	wire _w11051_ ;
	wire _w11050_ ;
	wire _w11049_ ;
	wire _w11048_ ;
	wire _w11047_ ;
	wire _w11046_ ;
	wire _w11045_ ;
	wire _w11044_ ;
	wire _w11043_ ;
	wire _w11042_ ;
	wire _w11041_ ;
	wire _w11040_ ;
	wire _w11039_ ;
	wire _w11038_ ;
	wire _w11037_ ;
	wire _w11036_ ;
	wire _w11035_ ;
	wire _w11034_ ;
	wire _w11033_ ;
	wire _w11032_ ;
	wire _w11031_ ;
	wire _w11030_ ;
	wire _w11029_ ;
	wire _w11028_ ;
	wire _w11027_ ;
	wire _w11026_ ;
	wire _w11025_ ;
	wire _w11024_ ;
	wire _w11023_ ;
	wire _w11022_ ;
	wire _w11021_ ;
	wire _w11020_ ;
	wire _w11019_ ;
	wire _w11018_ ;
	wire _w11017_ ;
	wire _w11016_ ;
	wire _w11015_ ;
	wire _w11014_ ;
	wire _w11013_ ;
	wire _w11012_ ;
	wire _w11011_ ;
	wire _w11010_ ;
	wire _w11009_ ;
	wire _w11008_ ;
	wire _w11007_ ;
	wire _w11006_ ;
	wire _w11005_ ;
	wire _w11004_ ;
	wire _w11003_ ;
	wire _w11002_ ;
	wire _w11001_ ;
	wire _w11000_ ;
	wire _w10999_ ;
	wire _w10998_ ;
	wire _w10997_ ;
	wire _w10996_ ;
	wire _w10995_ ;
	wire _w10994_ ;
	wire _w10993_ ;
	wire _w10992_ ;
	wire _w10991_ ;
	wire _w10990_ ;
	wire _w10989_ ;
	wire _w10988_ ;
	wire _w10987_ ;
	wire _w10986_ ;
	wire _w10985_ ;
	wire _w10984_ ;
	wire _w10983_ ;
	wire _w10982_ ;
	wire _w10981_ ;
	wire _w10980_ ;
	wire _w10979_ ;
	wire _w10978_ ;
	wire _w10977_ ;
	wire _w10976_ ;
	wire _w10975_ ;
	wire _w10974_ ;
	wire _w10973_ ;
	wire _w10972_ ;
	wire _w10971_ ;
	wire _w10970_ ;
	wire _w10969_ ;
	wire _w10968_ ;
	wire _w10967_ ;
	wire _w10966_ ;
	wire _w10965_ ;
	wire _w10964_ ;
	wire _w10963_ ;
	wire _w10962_ ;
	wire _w10961_ ;
	wire _w10960_ ;
	wire _w10959_ ;
	wire _w10958_ ;
	wire _w10957_ ;
	wire _w10956_ ;
	wire _w10955_ ;
	wire _w10954_ ;
	wire _w10953_ ;
	wire _w10952_ ;
	wire _w10951_ ;
	wire _w10950_ ;
	wire _w10949_ ;
	wire _w10948_ ;
	wire _w10947_ ;
	wire _w10946_ ;
	wire _w10945_ ;
	wire _w10944_ ;
	wire _w10943_ ;
	wire _w10942_ ;
	wire _w10941_ ;
	wire _w10940_ ;
	wire _w10939_ ;
	wire _w10938_ ;
	wire _w10937_ ;
	wire _w10936_ ;
	wire _w10935_ ;
	wire _w10934_ ;
	wire _w10933_ ;
	wire _w10932_ ;
	wire _w10931_ ;
	wire _w10930_ ;
	wire _w10929_ ;
	wire _w10928_ ;
	wire _w10927_ ;
	wire _w10926_ ;
	wire _w10925_ ;
	wire _w10924_ ;
	wire _w10923_ ;
	wire _w10922_ ;
	wire _w10921_ ;
	wire _w10920_ ;
	wire _w10919_ ;
	wire _w10918_ ;
	wire _w10917_ ;
	wire _w10916_ ;
	wire _w10915_ ;
	wire _w10914_ ;
	wire _w10913_ ;
	wire _w10912_ ;
	wire _w10911_ ;
	wire _w10910_ ;
	wire _w10909_ ;
	wire _w10908_ ;
	wire _w10907_ ;
	wire _w10906_ ;
	wire _w10905_ ;
	wire _w10904_ ;
	wire _w10903_ ;
	wire _w10902_ ;
	wire _w10901_ ;
	wire _w10900_ ;
	wire _w10899_ ;
	wire _w10898_ ;
	wire _w10897_ ;
	wire _w10896_ ;
	wire _w10895_ ;
	wire _w10894_ ;
	wire _w10893_ ;
	wire _w10892_ ;
	wire _w10891_ ;
	wire _w10890_ ;
	wire _w10889_ ;
	wire _w10888_ ;
	wire _w10887_ ;
	wire _w10886_ ;
	wire _w10885_ ;
	wire _w10884_ ;
	wire _w10883_ ;
	wire _w10882_ ;
	wire _w10881_ ;
	wire _w10880_ ;
	wire _w10879_ ;
	wire _w10878_ ;
	wire _w10877_ ;
	wire _w10876_ ;
	wire _w10875_ ;
	wire _w10874_ ;
	wire _w10873_ ;
	wire _w10872_ ;
	wire _w10871_ ;
	wire _w10870_ ;
	wire _w10869_ ;
	wire _w10868_ ;
	wire _w10867_ ;
	wire _w10866_ ;
	wire _w10865_ ;
	wire _w10864_ ;
	wire _w10863_ ;
	wire _w10862_ ;
	wire _w10861_ ;
	wire _w10860_ ;
	wire _w10859_ ;
	wire _w10858_ ;
	wire _w10857_ ;
	wire _w10856_ ;
	wire _w10855_ ;
	wire _w10854_ ;
	wire _w10853_ ;
	wire _w10852_ ;
	wire _w10851_ ;
	wire _w10850_ ;
	wire _w10849_ ;
	wire _w10848_ ;
	wire _w10847_ ;
	wire _w10846_ ;
	wire _w10845_ ;
	wire _w10844_ ;
	wire _w10843_ ;
	wire _w10842_ ;
	wire _w10841_ ;
	wire _w10840_ ;
	wire _w10839_ ;
	wire _w10838_ ;
	wire _w10837_ ;
	wire _w10836_ ;
	wire _w10835_ ;
	wire _w10834_ ;
	wire _w10833_ ;
	wire _w10832_ ;
	wire _w10831_ ;
	wire _w10830_ ;
	wire _w10829_ ;
	wire _w10828_ ;
	wire _w10827_ ;
	wire _w10826_ ;
	wire _w10825_ ;
	wire _w10824_ ;
	wire _w10823_ ;
	wire _w10822_ ;
	wire _w10821_ ;
	wire _w10820_ ;
	wire _w10819_ ;
	wire _w10818_ ;
	wire _w10817_ ;
	wire _w10816_ ;
	wire _w10815_ ;
	wire _w10814_ ;
	wire _w10813_ ;
	wire _w10812_ ;
	wire _w10811_ ;
	wire _w10810_ ;
	wire _w10809_ ;
	wire _w10808_ ;
	wire _w10807_ ;
	wire _w10806_ ;
	wire _w10805_ ;
	wire _w10804_ ;
	wire _w10803_ ;
	wire _w10802_ ;
	wire _w10801_ ;
	wire _w10800_ ;
	wire _w10799_ ;
	wire _w10798_ ;
	wire _w10797_ ;
	wire _w10796_ ;
	wire _w10795_ ;
	wire _w10794_ ;
	wire _w10793_ ;
	wire _w10792_ ;
	wire _w10791_ ;
	wire _w10790_ ;
	wire _w10789_ ;
	wire _w10788_ ;
	wire _w10787_ ;
	wire _w10786_ ;
	wire _w10785_ ;
	wire _w10784_ ;
	wire _w10783_ ;
	wire _w10782_ ;
	wire _w10781_ ;
	wire _w10780_ ;
	wire _w10779_ ;
	wire _w10778_ ;
	wire _w10777_ ;
	wire _w10776_ ;
	wire _w10775_ ;
	wire _w10774_ ;
	wire _w10773_ ;
	wire _w10772_ ;
	wire _w10771_ ;
	wire _w10770_ ;
	wire _w10769_ ;
	wire _w10768_ ;
	wire _w10767_ ;
	wire _w10766_ ;
	wire _w10765_ ;
	wire _w10764_ ;
	wire _w10763_ ;
	wire _w10762_ ;
	wire _w10761_ ;
	wire _w10760_ ;
	wire _w10759_ ;
	wire _w10758_ ;
	wire _w10757_ ;
	wire _w10756_ ;
	wire _w10755_ ;
	wire _w10754_ ;
	wire _w10753_ ;
	wire _w10752_ ;
	wire _w10751_ ;
	wire _w10750_ ;
	wire _w10749_ ;
	wire _w10748_ ;
	wire _w10747_ ;
	wire _w10746_ ;
	wire _w10745_ ;
	wire _w10744_ ;
	wire _w10743_ ;
	wire _w10742_ ;
	wire _w10741_ ;
	wire _w10740_ ;
	wire _w10739_ ;
	wire _w10738_ ;
	wire _w10737_ ;
	wire _w10736_ ;
	wire _w10735_ ;
	wire _w5548_ ;
	wire _w5547_ ;
	wire _w5546_ ;
	wire _w5545_ ;
	wire _w5544_ ;
	wire _w5543_ ;
	wire _w5542_ ;
	wire _w5541_ ;
	wire _w5540_ ;
	wire _w5539_ ;
	wire _w5538_ ;
	wire _w5537_ ;
	wire _w5536_ ;
	wire _w5535_ ;
	wire _w5534_ ;
	wire _w5533_ ;
	wire _w5532_ ;
	wire _w5531_ ;
	wire _w5530_ ;
	wire _w5529_ ;
	wire _w5528_ ;
	wire _w5527_ ;
	wire _w5526_ ;
	wire _w5525_ ;
	wire _w5524_ ;
	wire _w5523_ ;
	wire _w5522_ ;
	wire _w5521_ ;
	wire _w5520_ ;
	wire _w5519_ ;
	wire _w5518_ ;
	wire _w5517_ ;
	wire _w5516_ ;
	wire _w5515_ ;
	wire _w5514_ ;
	wire _w5513_ ;
	wire _w5512_ ;
	wire _w5511_ ;
	wire _w5510_ ;
	wire _w5509_ ;
	wire _w5508_ ;
	wire _w5507_ ;
	wire _w5506_ ;
	wire _w5505_ ;
	wire _w5504_ ;
	wire _w5503_ ;
	wire _w5502_ ;
	wire _w5501_ ;
	wire _w5500_ ;
	wire _w5499_ ;
	wire _w5498_ ;
	wire _w5497_ ;
	wire _w5496_ ;
	wire _w5495_ ;
	wire _w5494_ ;
	wire _w5493_ ;
	wire _w5492_ ;
	wire _w5491_ ;
	wire _w5490_ ;
	wire _w5489_ ;
	wire _w5488_ ;
	wire _w5487_ ;
	wire _w5486_ ;
	wire _w5485_ ;
	wire _w5484_ ;
	wire _w5483_ ;
	wire _w5482_ ;
	wire _w5481_ ;
	wire _w5480_ ;
	wire _w5479_ ;
	wire _w5478_ ;
	wire _w5477_ ;
	wire _w5476_ ;
	wire _w5475_ ;
	wire _w5474_ ;
	wire _w5473_ ;
	wire _w5472_ ;
	wire _w5471_ ;
	wire _w5470_ ;
	wire _w5469_ ;
	wire _w5468_ ;
	wire _w5467_ ;
	wire _w5466_ ;
	wire _w5465_ ;
	wire _w5464_ ;
	wire _w5463_ ;
	wire _w5462_ ;
	wire _w5461_ ;
	wire _w5460_ ;
	wire _w5459_ ;
	wire _w5458_ ;
	wire _w5457_ ;
	wire _w5456_ ;
	wire _w5455_ ;
	wire _w5454_ ;
	wire _w5453_ ;
	wire _w5452_ ;
	wire _w5451_ ;
	wire _w5450_ ;
	wire _w5449_ ;
	wire _w5448_ ;
	wire _w5447_ ;
	wire _w5446_ ;
	wire _w5445_ ;
	wire _w5444_ ;
	wire _w5443_ ;
	wire _w5442_ ;
	wire _w5441_ ;
	wire _w5440_ ;
	wire _w5439_ ;
	wire _w5438_ ;
	wire _w5437_ ;
	wire _w5436_ ;
	wire _w5435_ ;
	wire _w5434_ ;
	wire _w5433_ ;
	wire _w5432_ ;
	wire _w5431_ ;
	wire _w5430_ ;
	wire _w5429_ ;
	wire _w5428_ ;
	wire _w5427_ ;
	wire _w5426_ ;
	wire _w5425_ ;
	wire _w5424_ ;
	wire _w5423_ ;
	wire _w5422_ ;
	wire _w5421_ ;
	wire _w5420_ ;
	wire _w5419_ ;
	wire _w5418_ ;
	wire _w5417_ ;
	wire _w5416_ ;
	wire _w5415_ ;
	wire _w5414_ ;
	wire _w5413_ ;
	wire _w5412_ ;
	wire _w5411_ ;
	wire _w5410_ ;
	wire _w5409_ ;
	wire _w5408_ ;
	wire _w5407_ ;
	wire _w5406_ ;
	wire _w5405_ ;
	wire _w5404_ ;
	wire _w5403_ ;
	wire _w5402_ ;
	wire _w5401_ ;
	wire _w5400_ ;
	wire _w5399_ ;
	wire _w5398_ ;
	wire _w5397_ ;
	wire _w5396_ ;
	wire _w5395_ ;
	wire _w5394_ ;
	wire _w5393_ ;
	wire _w5392_ ;
	wire _w5391_ ;
	wire _w5390_ ;
	wire _w5389_ ;
	wire _w5388_ ;
	wire _w5387_ ;
	wire _w5386_ ;
	wire _w5385_ ;
	wire _w5384_ ;
	wire _w5383_ ;
	wire _w5382_ ;
	wire _w5381_ ;
	wire _w5380_ ;
	wire _w5379_ ;
	wire _w5378_ ;
	wire _w5377_ ;
	wire _w5376_ ;
	wire _w5375_ ;
	wire _w5374_ ;
	wire _w5373_ ;
	wire _w5372_ ;
	wire _w5371_ ;
	wire _w5370_ ;
	wire _w5369_ ;
	wire _w5368_ ;
	wire _w5367_ ;
	wire _w5366_ ;
	wire _w5365_ ;
	wire _w5364_ ;
	wire _w5363_ ;
	wire _w5362_ ;
	wire _w5361_ ;
	wire _w5360_ ;
	wire _w5359_ ;
	wire _w5358_ ;
	wire _w5357_ ;
	wire _w5356_ ;
	wire _w5355_ ;
	wire _w5354_ ;
	wire _w5353_ ;
	wire _w5352_ ;
	wire _w5351_ ;
	wire _w5350_ ;
	wire _w5349_ ;
	wire _w5348_ ;
	wire _w5347_ ;
	wire _w5346_ ;
	wire _w5345_ ;
	wire _w5344_ ;
	wire _w5343_ ;
	wire _w5342_ ;
	wire _w5341_ ;
	wire _w5340_ ;
	wire _w5339_ ;
	wire _w5338_ ;
	wire _w5337_ ;
	wire _w5336_ ;
	wire _w5335_ ;
	wire _w5334_ ;
	wire _w5333_ ;
	wire _w5332_ ;
	wire _w5331_ ;
	wire _w5330_ ;
	wire _w5329_ ;
	wire _w5328_ ;
	wire _w5327_ ;
	wire _w5326_ ;
	wire _w5325_ ;
	wire _w5324_ ;
	wire _w5323_ ;
	wire _w5322_ ;
	wire _w5321_ ;
	wire _w5320_ ;
	wire _w5319_ ;
	wire _w5318_ ;
	wire _w5317_ ;
	wire _w5316_ ;
	wire _w5315_ ;
	wire _w5314_ ;
	wire _w5313_ ;
	wire _w5312_ ;
	wire _w5311_ ;
	wire _w5310_ ;
	wire _w5309_ ;
	wire _w5308_ ;
	wire _w5307_ ;
	wire _w5306_ ;
	wire _w5305_ ;
	wire _w5304_ ;
	wire _w5303_ ;
	wire _w5302_ ;
	wire _w5301_ ;
	wire _w5300_ ;
	wire _w5299_ ;
	wire _w5298_ ;
	wire _w5297_ ;
	wire _w5296_ ;
	wire _w5295_ ;
	wire _w5294_ ;
	wire _w5293_ ;
	wire _w5292_ ;
	wire _w5291_ ;
	wire _w5290_ ;
	wire _w5289_ ;
	wire _w5288_ ;
	wire _w5287_ ;
	wire _w5286_ ;
	wire _w5285_ ;
	wire _w5284_ ;
	wire _w5283_ ;
	wire _w5282_ ;
	wire _w5281_ ;
	wire _w5280_ ;
	wire _w5279_ ;
	wire _w5278_ ;
	wire _w5277_ ;
	wire _w5276_ ;
	wire _w5275_ ;
	wire _w5274_ ;
	wire _w5273_ ;
	wire _w5272_ ;
	wire _w5271_ ;
	wire _w5270_ ;
	wire _w5269_ ;
	wire _w5268_ ;
	wire _w5267_ ;
	wire _w5266_ ;
	wire _w5265_ ;
	wire _w5264_ ;
	wire _w5263_ ;
	wire _w5262_ ;
	wire _w5261_ ;
	wire _w5260_ ;
	wire _w5259_ ;
	wire _w5258_ ;
	wire _w5257_ ;
	wire _w5256_ ;
	wire _w5255_ ;
	wire _w5254_ ;
	wire _w5253_ ;
	wire _w5252_ ;
	wire _w5251_ ;
	wire _w5250_ ;
	wire _w5249_ ;
	wire _w5248_ ;
	wire _w5247_ ;
	wire _w5246_ ;
	wire _w5245_ ;
	wire _w5244_ ;
	wire _w5243_ ;
	wire _w5242_ ;
	wire _w5241_ ;
	wire _w5240_ ;
	wire _w5239_ ;
	wire _w5238_ ;
	wire _w5237_ ;
	wire _w5236_ ;
	wire _w5235_ ;
	wire _w5234_ ;
	wire _w5233_ ;
	wire _w5232_ ;
	wire _w5231_ ;
	wire _w5230_ ;
	wire _w5229_ ;
	wire _w5228_ ;
	wire _w5227_ ;
	wire _w5226_ ;
	wire _w5225_ ;
	wire _w5224_ ;
	wire _w5223_ ;
	wire _w5222_ ;
	wire _w5221_ ;
	wire _w5220_ ;
	wire _w5219_ ;
	wire _w5218_ ;
	wire _w5217_ ;
	wire _w5216_ ;
	wire _w5215_ ;
	wire _w5214_ ;
	wire _w5213_ ;
	wire _w5212_ ;
	wire _w5211_ ;
	wire _w5210_ ;
	wire _w5209_ ;
	wire _w5208_ ;
	wire _w5207_ ;
	wire _w5206_ ;
	wire _w5205_ ;
	wire _w5204_ ;
	wire _w5203_ ;
	wire _w5202_ ;
	wire _w5201_ ;
	wire _w5200_ ;
	wire _w5199_ ;
	wire _w5198_ ;
	wire _w5197_ ;
	wire _w5196_ ;
	wire _w5195_ ;
	wire _w5194_ ;
	wire _w5193_ ;
	wire _w5192_ ;
	wire _w5191_ ;
	wire _w5190_ ;
	wire _w5189_ ;
	wire _w5188_ ;
	wire _w5187_ ;
	wire _w5186_ ;
	wire _w5185_ ;
	wire _w5184_ ;
	wire _w5183_ ;
	wire _w5182_ ;
	wire _w5181_ ;
	wire _w5180_ ;
	wire _w5179_ ;
	wire _w5178_ ;
	wire _w5177_ ;
	wire _w5176_ ;
	wire _w5175_ ;
	wire _w5174_ ;
	wire _w5173_ ;
	wire _w5172_ ;
	wire _w5171_ ;
	wire _w5170_ ;
	wire _w5169_ ;
	wire _w5168_ ;
	wire _w5167_ ;
	wire _w5166_ ;
	wire _w5165_ ;
	wire _w5164_ ;
	wire _w5163_ ;
	wire _w5162_ ;
	wire _w5161_ ;
	wire _w5160_ ;
	wire _w5159_ ;
	wire _w5158_ ;
	wire _w5157_ ;
	wire _w5156_ ;
	wire _w5155_ ;
	wire _w5154_ ;
	wire _w5153_ ;
	wire _w5152_ ;
	wire _w5151_ ;
	wire _w5150_ ;
	wire _w5149_ ;
	wire _w5148_ ;
	wire _w5147_ ;
	wire _w5146_ ;
	wire _w5145_ ;
	wire _w5144_ ;
	wire _w5143_ ;
	wire _w5142_ ;
	wire _w5141_ ;
	wire _w5140_ ;
	wire _w5139_ ;
	wire _w5138_ ;
	wire _w5137_ ;
	wire _w5136_ ;
	wire _w5135_ ;
	wire _w5134_ ;
	wire _w5133_ ;
	wire _w5132_ ;
	wire _w5131_ ;
	wire _w5130_ ;
	wire _w5129_ ;
	wire _w5128_ ;
	wire _w5127_ ;
	wire _w5126_ ;
	wire _w5125_ ;
	wire _w5124_ ;
	wire _w5123_ ;
	wire _w5122_ ;
	wire _w5121_ ;
	wire _w5120_ ;
	wire _w5119_ ;
	wire _w5118_ ;
	wire _w5117_ ;
	wire _w5116_ ;
	wire _w5115_ ;
	wire _w5114_ ;
	wire _w5113_ ;
	wire _w5112_ ;
	wire _w5111_ ;
	wire _w5110_ ;
	wire _w5109_ ;
	wire _w5108_ ;
	wire _w5107_ ;
	wire _w5106_ ;
	wire _w5105_ ;
	wire _w5104_ ;
	wire _w5103_ ;
	wire _w5102_ ;
	wire _w5101_ ;
	wire _w5100_ ;
	wire _w5099_ ;
	wire _w5098_ ;
	wire _w5097_ ;
	wire _w5096_ ;
	wire _w5095_ ;
	wire _w5094_ ;
	wire _w5093_ ;
	wire _w5092_ ;
	wire _w5091_ ;
	wire _w5090_ ;
	wire _w5089_ ;
	wire _w5088_ ;
	wire _w5087_ ;
	wire _w5086_ ;
	wire _w5085_ ;
	wire _w5084_ ;
	wire _w5083_ ;
	wire _w5082_ ;
	wire _w5081_ ;
	wire _w5080_ ;
	wire _w5079_ ;
	wire _w5078_ ;
	wire _w5077_ ;
	wire _w5076_ ;
	wire _w5075_ ;
	wire _w5074_ ;
	wire _w5073_ ;
	wire _w5072_ ;
	wire _w5071_ ;
	wire _w5070_ ;
	wire _w5069_ ;
	wire _w5068_ ;
	wire _w5067_ ;
	wire _w5066_ ;
	wire _w5065_ ;
	wire _w5064_ ;
	wire _w5063_ ;
	wire _w5062_ ;
	wire _w5061_ ;
	wire _w5060_ ;
	wire _w5059_ ;
	wire _w5058_ ;
	wire _w5057_ ;
	wire _w5056_ ;
	wire _w5055_ ;
	wire _w5054_ ;
	wire _w5053_ ;
	wire _w5052_ ;
	wire _w5051_ ;
	wire _w5050_ ;
	wire _w5049_ ;
	wire _w5048_ ;
	wire _w5047_ ;
	wire _w5046_ ;
	wire _w5045_ ;
	wire _w5044_ ;
	wire _w5043_ ;
	wire _w5042_ ;
	wire _w5041_ ;
	wire _w5040_ ;
	wire _w5039_ ;
	wire _w5038_ ;
	wire _w5037_ ;
	wire _w5036_ ;
	wire _w5035_ ;
	wire _w5034_ ;
	wire _w5033_ ;
	wire _w5032_ ;
	wire _w5031_ ;
	wire _w5030_ ;
	wire _w5029_ ;
	wire _w5028_ ;
	wire _w5027_ ;
	wire _w5026_ ;
	wire _w5025_ ;
	wire _w5024_ ;
	wire _w5023_ ;
	wire _w5022_ ;
	wire _w5021_ ;
	wire _w5020_ ;
	wire _w5019_ ;
	wire _w5018_ ;
	wire _w5017_ ;
	wire _w5016_ ;
	wire _w5015_ ;
	wire _w5014_ ;
	wire _w5013_ ;
	wire _w5012_ ;
	wire _w5011_ ;
	wire _w5010_ ;
	wire _w5009_ ;
	wire _w5008_ ;
	wire _w5007_ ;
	wire _w5006_ ;
	wire _w5005_ ;
	wire _w5004_ ;
	wire _w5003_ ;
	wire _w5002_ ;
	wire _w5001_ ;
	wire _w5000_ ;
	wire _w4999_ ;
	wire _w4998_ ;
	wire _w4997_ ;
	wire _w4996_ ;
	wire _w4995_ ;
	wire _w4994_ ;
	wire _w4993_ ;
	wire _w4992_ ;
	wire _w4991_ ;
	wire _w4990_ ;
	wire _w4989_ ;
	wire _w4988_ ;
	wire _w4987_ ;
	wire _w4986_ ;
	wire _w4985_ ;
	wire _w4984_ ;
	wire _w4983_ ;
	wire _w4982_ ;
	wire _w4981_ ;
	wire _w4980_ ;
	wire _w4979_ ;
	wire _w4978_ ;
	wire _w4977_ ;
	wire _w4976_ ;
	wire _w4975_ ;
	wire _w4974_ ;
	wire _w4973_ ;
	wire _w4972_ ;
	wire _w4971_ ;
	wire _w4970_ ;
	wire _w4969_ ;
	wire _w4968_ ;
	wire _w4967_ ;
	wire _w4966_ ;
	wire _w4965_ ;
	wire _w4964_ ;
	wire _w4963_ ;
	wire _w4962_ ;
	wire _w4961_ ;
	wire _w4960_ ;
	wire _w4959_ ;
	wire _w4958_ ;
	wire _w4957_ ;
	wire _w4956_ ;
	wire _w4955_ ;
	wire _w4954_ ;
	wire _w4953_ ;
	wire _w4952_ ;
	wire _w4951_ ;
	wire _w4950_ ;
	wire _w4949_ ;
	wire _w4948_ ;
	wire _w4947_ ;
	wire _w4946_ ;
	wire _w4945_ ;
	wire _w4944_ ;
	wire _w4943_ ;
	wire _w4942_ ;
	wire _w4941_ ;
	wire _w4940_ ;
	wire _w4939_ ;
	wire _w4938_ ;
	wire _w4937_ ;
	wire _w4936_ ;
	wire _w4935_ ;
	wire _w4934_ ;
	wire _w4933_ ;
	wire _w4932_ ;
	wire _w4931_ ;
	wire _w4930_ ;
	wire _w4929_ ;
	wire _w4928_ ;
	wire _w4927_ ;
	wire _w4926_ ;
	wire _w4925_ ;
	wire _w4924_ ;
	wire _w4923_ ;
	wire _w4922_ ;
	wire _w4921_ ;
	wire _w4920_ ;
	wire _w4919_ ;
	wire _w4918_ ;
	wire _w4917_ ;
	wire _w4916_ ;
	wire _w4915_ ;
	wire _w4914_ ;
	wire _w4913_ ;
	wire _w4912_ ;
	wire _w4911_ ;
	wire _w4910_ ;
	wire _w4909_ ;
	wire _w4908_ ;
	wire _w4907_ ;
	wire _w4906_ ;
	wire _w4905_ ;
	wire _w4904_ ;
	wire _w4903_ ;
	wire _w4902_ ;
	wire _w4901_ ;
	wire _w4900_ ;
	wire _w4899_ ;
	wire _w4898_ ;
	wire _w4897_ ;
	wire _w4896_ ;
	wire _w4895_ ;
	wire _w4894_ ;
	wire _w4893_ ;
	wire _w4892_ ;
	wire _w4891_ ;
	wire _w4890_ ;
	wire _w4889_ ;
	wire _w4888_ ;
	wire _w4887_ ;
	wire _w4886_ ;
	wire _w4885_ ;
	wire _w4884_ ;
	wire _w4883_ ;
	wire _w4882_ ;
	wire _w4881_ ;
	wire _w4880_ ;
	wire _w4879_ ;
	wire _w4878_ ;
	wire _w4877_ ;
	wire _w4876_ ;
	wire _w4875_ ;
	wire _w4874_ ;
	wire _w4873_ ;
	wire _w4872_ ;
	wire _w4871_ ;
	wire _w4870_ ;
	wire _w4869_ ;
	wire _w4868_ ;
	wire _w4867_ ;
	wire _w4866_ ;
	wire _w4865_ ;
	wire _w4864_ ;
	wire _w4863_ ;
	wire _w4862_ ;
	wire _w4861_ ;
	wire _w4860_ ;
	wire _w4859_ ;
	wire _w4858_ ;
	wire _w4857_ ;
	wire _w4856_ ;
	wire _w4855_ ;
	wire _w4854_ ;
	wire _w4853_ ;
	wire _w4852_ ;
	wire _w4851_ ;
	wire _w4850_ ;
	wire _w4849_ ;
	wire _w4848_ ;
	wire _w4847_ ;
	wire _w4846_ ;
	wire _w4845_ ;
	wire _w4844_ ;
	wire _w4843_ ;
	wire _w4842_ ;
	wire _w4841_ ;
	wire _w4840_ ;
	wire _w4839_ ;
	wire _w4838_ ;
	wire _w4837_ ;
	wire _w4836_ ;
	wire _w4835_ ;
	wire _w4834_ ;
	wire _w4833_ ;
	wire _w4832_ ;
	wire _w4831_ ;
	wire _w4830_ ;
	wire _w4829_ ;
	wire _w4828_ ;
	wire _w4827_ ;
	wire _w4826_ ;
	wire _w4825_ ;
	wire _w4824_ ;
	wire _w4823_ ;
	wire _w4822_ ;
	wire _w4821_ ;
	wire _w4820_ ;
	wire _w4819_ ;
	wire _w4818_ ;
	wire _w4817_ ;
	wire _w4816_ ;
	wire _w4815_ ;
	wire _w4814_ ;
	wire _w4813_ ;
	wire _w4812_ ;
	wire _w4811_ ;
	wire _w4810_ ;
	wire _w4809_ ;
	wire _w4808_ ;
	wire _w4807_ ;
	wire _w4806_ ;
	wire _w4805_ ;
	wire _w4804_ ;
	wire _w4803_ ;
	wire _w4802_ ;
	wire _w4801_ ;
	wire _w4800_ ;
	wire _w4799_ ;
	wire _w4798_ ;
	wire _w4797_ ;
	wire _w4796_ ;
	wire _w4795_ ;
	wire _w4794_ ;
	wire _w4793_ ;
	wire _w4792_ ;
	wire _w4791_ ;
	wire _w4790_ ;
	wire _w4789_ ;
	wire _w4788_ ;
	wire _w4787_ ;
	wire _w4786_ ;
	wire _w4785_ ;
	wire _w4784_ ;
	wire _w4783_ ;
	wire _w4782_ ;
	wire _w4781_ ;
	wire _w4780_ ;
	wire _w4779_ ;
	wire _w4778_ ;
	wire _w4777_ ;
	wire _w4776_ ;
	wire _w4775_ ;
	wire _w4774_ ;
	wire _w4773_ ;
	wire _w4772_ ;
	wire _w4771_ ;
	wire _w4770_ ;
	wire _w4769_ ;
	wire _w4768_ ;
	wire _w4767_ ;
	wire _w4766_ ;
	wire _w4765_ ;
	wire _w4764_ ;
	wire _w4763_ ;
	wire _w4762_ ;
	wire _w4761_ ;
	wire _w4760_ ;
	wire _w4759_ ;
	wire _w4758_ ;
	wire _w4757_ ;
	wire _w4756_ ;
	wire _w4755_ ;
	wire _w4754_ ;
	wire _w4753_ ;
	wire _w4752_ ;
	wire _w4751_ ;
	wire _w4750_ ;
	wire _w4749_ ;
	wire _w4748_ ;
	wire _w4747_ ;
	wire _w4746_ ;
	wire _w4745_ ;
	wire _w4744_ ;
	wire _w4743_ ;
	wire _w4742_ ;
	wire _w4741_ ;
	wire _w4740_ ;
	wire _w4739_ ;
	wire _w4738_ ;
	wire _w4737_ ;
	wire _w4736_ ;
	wire _w4735_ ;
	wire _w4734_ ;
	wire _w4733_ ;
	wire _w4732_ ;
	wire _w4731_ ;
	wire _w4730_ ;
	wire _w4729_ ;
	wire _w4728_ ;
	wire _w4727_ ;
	wire _w4726_ ;
	wire _w4725_ ;
	wire _w4724_ ;
	wire _w4723_ ;
	wire _w4722_ ;
	wire _w4721_ ;
	wire _w4720_ ;
	wire _w4719_ ;
	wire _w4718_ ;
	wire _w4717_ ;
	wire _w4716_ ;
	wire _w4715_ ;
	wire _w4714_ ;
	wire _w4713_ ;
	wire _w4712_ ;
	wire _w4711_ ;
	wire _w4710_ ;
	wire _w4709_ ;
	wire _w4708_ ;
	wire _w4707_ ;
	wire _w4706_ ;
	wire _w4705_ ;
	wire _w4704_ ;
	wire _w4703_ ;
	wire _w4702_ ;
	wire _w4701_ ;
	wire _w4700_ ;
	wire _w4699_ ;
	wire _w4698_ ;
	wire _w4697_ ;
	wire _w4696_ ;
	wire _w4695_ ;
	wire _w4694_ ;
	wire _w4693_ ;
	wire _w4692_ ;
	wire _w4691_ ;
	wire _w4690_ ;
	wire _w4689_ ;
	wire _w4688_ ;
	wire _w4687_ ;
	wire _w4686_ ;
	wire _w4685_ ;
	wire _w4684_ ;
	wire _w4683_ ;
	wire _w4682_ ;
	wire _w4681_ ;
	wire _w4680_ ;
	wire _w4679_ ;
	wire _w4678_ ;
	wire _w4677_ ;
	wire _w4676_ ;
	wire _w4675_ ;
	wire _w4674_ ;
	wire _w4673_ ;
	wire _w4672_ ;
	wire _w4671_ ;
	wire _w4670_ ;
	wire _w4669_ ;
	wire _w4668_ ;
	wire _w4667_ ;
	wire _w4666_ ;
	wire _w4665_ ;
	wire _w4664_ ;
	wire _w4663_ ;
	wire _w4662_ ;
	wire _w4661_ ;
	wire _w4660_ ;
	wire _w4659_ ;
	wire _w4658_ ;
	wire _w4657_ ;
	wire _w4656_ ;
	wire _w4655_ ;
	wire _w4654_ ;
	wire _w4653_ ;
	wire _w4652_ ;
	wire _w4651_ ;
	wire _w4650_ ;
	wire _w4649_ ;
	wire _w4648_ ;
	wire _w4647_ ;
	wire _w4646_ ;
	wire _w4645_ ;
	wire _w4644_ ;
	wire _w4643_ ;
	wire _w4642_ ;
	wire _w4641_ ;
	wire _w4640_ ;
	wire _w4639_ ;
	wire _w4638_ ;
	wire _w4637_ ;
	wire _w4636_ ;
	wire _w4635_ ;
	wire _w4634_ ;
	wire _w4633_ ;
	wire _w4632_ ;
	wire _w4631_ ;
	wire _w4630_ ;
	wire _w4629_ ;
	wire _w4628_ ;
	wire _w4627_ ;
	wire _w4626_ ;
	wire _w4625_ ;
	wire _w4624_ ;
	wire _w4623_ ;
	wire _w4622_ ;
	wire _w4621_ ;
	wire _w4620_ ;
	wire _w4619_ ;
	wire _w4618_ ;
	wire _w4617_ ;
	wire _w4616_ ;
	wire _w4615_ ;
	wire _w4614_ ;
	wire _w4613_ ;
	wire _w4612_ ;
	wire _w4611_ ;
	wire _w4610_ ;
	wire _w4609_ ;
	wire _w4608_ ;
	wire _w4607_ ;
	wire _w4606_ ;
	wire _w4605_ ;
	wire _w4604_ ;
	wire _w4603_ ;
	wire _w4602_ ;
	wire _w4601_ ;
	wire _w4600_ ;
	wire _w4599_ ;
	wire _w4598_ ;
	wire _w4597_ ;
	wire _w4596_ ;
	wire _w4595_ ;
	wire _w4594_ ;
	wire _w4593_ ;
	wire _w4592_ ;
	wire _w4591_ ;
	wire _w4590_ ;
	wire _w4589_ ;
	wire _w4588_ ;
	wire _w4587_ ;
	wire _w4586_ ;
	wire _w4585_ ;
	wire _w4584_ ;
	wire _w4583_ ;
	wire _w4582_ ;
	wire _w4581_ ;
	wire _w4580_ ;
	wire _w4579_ ;
	wire _w4578_ ;
	wire _w4577_ ;
	wire _w4576_ ;
	wire _w4575_ ;
	wire _w4574_ ;
	wire _w4573_ ;
	wire _w4572_ ;
	wire _w4571_ ;
	wire _w4570_ ;
	wire _w4569_ ;
	wire _w4568_ ;
	wire _w4567_ ;
	wire _w4566_ ;
	wire _w4565_ ;
	wire _w4564_ ;
	wire _w4563_ ;
	wire _w4562_ ;
	wire _w4561_ ;
	wire _w4560_ ;
	wire _w4559_ ;
	wire _w4558_ ;
	wire _w4557_ ;
	wire _w4556_ ;
	wire _w4555_ ;
	wire _w4554_ ;
	wire _w4553_ ;
	wire _w4552_ ;
	wire _w4551_ ;
	wire _w4550_ ;
	wire _w4549_ ;
	wire _w4548_ ;
	wire _w4547_ ;
	wire _w4546_ ;
	wire _w4545_ ;
	wire _w4544_ ;
	wire _w4543_ ;
	wire _w4542_ ;
	wire _w4541_ ;
	wire _w4540_ ;
	wire _w4539_ ;
	wire _w4538_ ;
	wire _w4537_ ;
	wire _w4536_ ;
	wire _w4535_ ;
	wire _w4534_ ;
	wire _w4533_ ;
	wire _w4532_ ;
	wire _w4531_ ;
	wire _w4530_ ;
	wire _w4529_ ;
	wire _w4528_ ;
	wire _w4527_ ;
	wire _w4526_ ;
	wire _w4525_ ;
	wire _w4524_ ;
	wire _w4523_ ;
	wire _w4522_ ;
	wire _w4521_ ;
	wire _w4520_ ;
	wire _w4519_ ;
	wire _w4518_ ;
	wire _w4517_ ;
	wire _w4516_ ;
	wire _w4515_ ;
	wire _w4514_ ;
	wire _w4513_ ;
	wire _w4512_ ;
	wire _w4511_ ;
	wire _w4510_ ;
	wire _w4509_ ;
	wire _w4508_ ;
	wire _w4507_ ;
	wire _w4506_ ;
	wire _w4505_ ;
	wire _w4504_ ;
	wire _w4503_ ;
	wire _w4502_ ;
	wire _w4501_ ;
	wire _w4500_ ;
	wire _w4499_ ;
	wire _w4498_ ;
	wire _w4497_ ;
	wire _w4496_ ;
	wire _w4495_ ;
	wire _w4494_ ;
	wire _w4493_ ;
	wire _w4492_ ;
	wire _w4491_ ;
	wire _w4490_ ;
	wire _w4489_ ;
	wire _w4488_ ;
	wire _w4487_ ;
	wire _w4486_ ;
	wire _w4485_ ;
	wire _w4484_ ;
	wire _w4483_ ;
	wire _w4482_ ;
	wire _w4481_ ;
	wire _w4480_ ;
	wire _w4479_ ;
	wire _w4478_ ;
	wire _w4477_ ;
	wire _w4476_ ;
	wire _w4475_ ;
	wire _w4474_ ;
	wire _w4473_ ;
	wire _w4472_ ;
	wire _w4471_ ;
	wire _w4470_ ;
	wire _w4469_ ;
	wire _w4468_ ;
	wire _w4467_ ;
	wire _w4466_ ;
	wire _w4465_ ;
	wire _w4464_ ;
	wire _w4463_ ;
	wire _w4462_ ;
	wire _w4461_ ;
	wire _w4460_ ;
	wire _w4459_ ;
	wire _w4458_ ;
	wire _w4457_ ;
	wire _w4456_ ;
	wire _w4455_ ;
	wire _w4454_ ;
	wire _w4453_ ;
	wire _w4452_ ;
	wire _w4451_ ;
	wire _w4450_ ;
	wire _w4449_ ;
	wire _w4448_ ;
	wire _w4447_ ;
	wire _w4446_ ;
	wire _w4445_ ;
	wire _w4444_ ;
	wire _w4443_ ;
	wire _w4442_ ;
	wire _w4441_ ;
	wire _w4440_ ;
	wire _w4439_ ;
	wire _w4438_ ;
	wire _w4437_ ;
	wire _w4436_ ;
	wire _w4435_ ;
	wire _w4434_ ;
	wire _w4433_ ;
	wire _w4432_ ;
	wire _w4431_ ;
	wire _w4430_ ;
	wire _w4429_ ;
	wire _w4428_ ;
	wire _w4427_ ;
	wire _w4426_ ;
	wire _w4425_ ;
	wire _w4424_ ;
	wire _w4423_ ;
	wire _w4422_ ;
	wire _w4421_ ;
	wire _w4420_ ;
	wire _w4419_ ;
	wire _w4418_ ;
	wire _w4417_ ;
	wire _w4416_ ;
	wire _w4415_ ;
	wire _w4414_ ;
	wire _w4413_ ;
	wire _w4412_ ;
	wire _w4411_ ;
	wire _w4410_ ;
	wire _w4409_ ;
	wire _w4408_ ;
	wire _w4407_ ;
	wire _w4406_ ;
	wire _w4405_ ;
	wire _w4404_ ;
	wire _w4403_ ;
	wire _w4402_ ;
	wire _w4401_ ;
	wire _w4400_ ;
	wire _w4399_ ;
	wire _w4398_ ;
	wire _w4397_ ;
	wire _w4396_ ;
	wire _w4395_ ;
	wire _w4394_ ;
	wire _w4393_ ;
	wire _w4392_ ;
	wire _w4391_ ;
	wire _w4390_ ;
	wire _w4389_ ;
	wire _w4388_ ;
	wire _w4387_ ;
	wire _w4386_ ;
	wire _w4385_ ;
	wire _w4384_ ;
	wire _w4383_ ;
	wire _w4382_ ;
	wire _w4381_ ;
	wire _w4380_ ;
	wire _w4379_ ;
	wire _w4378_ ;
	wire _w4377_ ;
	wire _w4376_ ;
	wire _w4375_ ;
	wire _w4374_ ;
	wire _w4373_ ;
	wire _w4372_ ;
	wire _w4371_ ;
	wire _w4370_ ;
	wire _w4369_ ;
	wire _w4368_ ;
	wire _w4367_ ;
	wire _w4366_ ;
	wire _w4365_ ;
	wire _w4364_ ;
	wire _w4363_ ;
	wire _w4362_ ;
	wire _w4361_ ;
	wire _w4360_ ;
	wire _w4359_ ;
	wire _w4358_ ;
	wire _w4357_ ;
	wire _w4356_ ;
	wire _w4355_ ;
	wire _w4354_ ;
	wire _w4353_ ;
	wire _w4352_ ;
	wire _w4351_ ;
	wire _w4350_ ;
	wire _w4349_ ;
	wire _w4348_ ;
	wire _w4347_ ;
	wire _w4346_ ;
	wire _w4345_ ;
	wire _w4344_ ;
	wire _w4343_ ;
	wire _w4342_ ;
	wire _w4341_ ;
	wire _w4340_ ;
	wire _w4339_ ;
	wire _w4338_ ;
	wire _w4337_ ;
	wire _w4336_ ;
	wire _w4335_ ;
	wire _w4334_ ;
	wire _w4333_ ;
	wire _w4332_ ;
	wire _w4331_ ;
	wire _w4330_ ;
	wire _w4329_ ;
	wire _w4328_ ;
	wire _w4327_ ;
	wire _w4326_ ;
	wire _w4325_ ;
	wire _w4324_ ;
	wire _w4323_ ;
	wire _w4322_ ;
	wire _w4321_ ;
	wire _w4320_ ;
	wire _w4319_ ;
	wire _w4318_ ;
	wire _w4317_ ;
	wire _w4316_ ;
	wire _w4315_ ;
	wire _w4314_ ;
	wire _w4313_ ;
	wire _w4312_ ;
	wire _w4311_ ;
	wire _w4310_ ;
	wire _w4309_ ;
	wire _w4308_ ;
	wire _w4307_ ;
	wire _w4306_ ;
	wire _w4305_ ;
	wire _w4304_ ;
	wire _w4303_ ;
	wire _w4302_ ;
	wire _w4301_ ;
	wire _w4300_ ;
	wire _w4299_ ;
	wire _w4298_ ;
	wire _w4297_ ;
	wire _w4296_ ;
	wire _w4295_ ;
	wire _w4294_ ;
	wire _w4293_ ;
	wire _w4292_ ;
	wire _w4291_ ;
	wire _w4290_ ;
	wire _w4289_ ;
	wire _w4288_ ;
	wire _w4287_ ;
	wire _w4286_ ;
	wire _w4285_ ;
	wire _w4284_ ;
	wire _w4283_ ;
	wire _w4282_ ;
	wire _w4281_ ;
	wire _w4280_ ;
	wire _w4279_ ;
	wire _w4278_ ;
	wire _w4277_ ;
	wire _w4276_ ;
	wire _w4275_ ;
	wire _w4274_ ;
	wire _w4273_ ;
	wire _w4272_ ;
	wire _w4271_ ;
	wire _w4270_ ;
	wire _w4269_ ;
	wire _w4268_ ;
	wire _w4267_ ;
	wire _w4266_ ;
	wire _w4265_ ;
	wire _w4264_ ;
	wire _w4263_ ;
	wire _w4262_ ;
	wire _w4261_ ;
	wire _w4260_ ;
	wire _w4259_ ;
	wire _w4258_ ;
	wire _w4257_ ;
	wire _w4256_ ;
	wire _w4255_ ;
	wire _w4254_ ;
	wire _w4253_ ;
	wire _w4252_ ;
	wire _w4251_ ;
	wire _w4250_ ;
	wire _w4249_ ;
	wire _w4248_ ;
	wire _w4247_ ;
	wire _w4246_ ;
	wire _w4245_ ;
	wire _w4244_ ;
	wire _w4243_ ;
	wire _w4242_ ;
	wire _w4241_ ;
	wire _w4240_ ;
	wire _w4239_ ;
	wire _w4238_ ;
	wire _w4237_ ;
	wire _w4236_ ;
	wire _w4235_ ;
	wire _w4234_ ;
	wire _w4233_ ;
	wire _w4232_ ;
	wire _w4231_ ;
	wire _w4230_ ;
	wire _w4229_ ;
	wire _w4228_ ;
	wire _w4227_ ;
	wire _w4226_ ;
	wire _w4225_ ;
	wire _w4224_ ;
	wire _w4223_ ;
	wire _w4222_ ;
	wire _w4221_ ;
	wire _w4220_ ;
	wire _w4219_ ;
	wire _w4218_ ;
	wire _w4217_ ;
	wire _w4216_ ;
	wire _w4215_ ;
	wire _w4214_ ;
	wire _w4213_ ;
	wire _w4212_ ;
	wire _w4211_ ;
	wire _w4210_ ;
	wire _w4209_ ;
	wire _w4208_ ;
	wire _w4207_ ;
	wire _w4206_ ;
	wire _w4205_ ;
	wire _w4204_ ;
	wire _w4203_ ;
	wire _w4202_ ;
	wire _w4201_ ;
	wire _w4200_ ;
	wire _w4199_ ;
	wire _w4198_ ;
	wire _w4197_ ;
	wire _w4196_ ;
	wire _w4195_ ;
	wire _w4194_ ;
	wire _w4193_ ;
	wire _w4192_ ;
	wire _w4191_ ;
	wire _w4190_ ;
	wire _w4189_ ;
	wire _w4188_ ;
	wire _w4187_ ;
	wire _w4186_ ;
	wire _w4185_ ;
	wire _w4184_ ;
	wire _w4183_ ;
	wire _w4182_ ;
	wire _w4181_ ;
	wire _w4180_ ;
	wire _w4179_ ;
	wire _w4178_ ;
	wire _w4177_ ;
	wire _w4176_ ;
	wire _w4175_ ;
	wire _w4174_ ;
	wire _w4173_ ;
	wire _w4172_ ;
	wire _w4171_ ;
	wire _w4170_ ;
	wire _w4169_ ;
	wire _w4168_ ;
	wire _w4167_ ;
	wire _w4166_ ;
	wire _w4165_ ;
	wire _w4164_ ;
	wire _w4163_ ;
	wire _w4162_ ;
	wire _w4161_ ;
	wire _w4160_ ;
	wire _w4159_ ;
	wire _w4158_ ;
	wire _w4157_ ;
	wire _w4156_ ;
	wire _w4155_ ;
	wire _w4154_ ;
	wire _w4153_ ;
	wire _w4152_ ;
	wire _w4151_ ;
	wire _w4150_ ;
	wire _w4149_ ;
	wire _w4148_ ;
	wire _w4147_ ;
	wire _w4146_ ;
	wire _w4145_ ;
	wire _w4144_ ;
	wire _w4143_ ;
	wire _w4142_ ;
	wire _w4141_ ;
	wire _w4140_ ;
	wire _w4139_ ;
	wire _w4138_ ;
	wire _w4137_ ;
	wire _w4136_ ;
	wire _w4135_ ;
	wire _w4134_ ;
	wire _w4133_ ;
	wire _w4132_ ;
	wire _w4131_ ;
	wire _w4130_ ;
	wire _w4129_ ;
	wire _w4128_ ;
	wire _w4127_ ;
	wire _w4126_ ;
	wire _w4125_ ;
	wire _w4124_ ;
	wire _w4123_ ;
	wire _w4122_ ;
	wire _w4121_ ;
	wire _w4120_ ;
	wire _w4119_ ;
	wire _w4118_ ;
	wire _w4117_ ;
	wire _w4116_ ;
	wire _w4115_ ;
	wire _w4114_ ;
	wire _w4113_ ;
	wire _w4112_ ;
	wire _w4111_ ;
	wire _w4110_ ;
	wire _w4109_ ;
	wire _w4108_ ;
	wire _w4107_ ;
	wire _w4106_ ;
	wire _w4105_ ;
	wire _w4104_ ;
	wire _w4103_ ;
	wire _w4102_ ;
	wire _w4101_ ;
	wire _w4100_ ;
	wire _w4099_ ;
	wire _w4098_ ;
	wire _w4097_ ;
	wire _w4096_ ;
	wire _w4095_ ;
	wire _w4094_ ;
	wire _w4093_ ;
	wire _w4092_ ;
	wire _w4091_ ;
	wire _w4090_ ;
	wire _w4089_ ;
	wire _w4088_ ;
	wire _w4087_ ;
	wire _w4086_ ;
	wire _w4085_ ;
	wire _w4084_ ;
	wire _w4083_ ;
	wire _w4082_ ;
	wire _w4081_ ;
	wire _w4080_ ;
	wire _w4079_ ;
	wire _w4078_ ;
	wire _w4077_ ;
	wire _w4076_ ;
	wire _w4075_ ;
	wire _w4074_ ;
	wire _w4073_ ;
	wire _w4072_ ;
	wire _w4071_ ;
	wire _w4070_ ;
	wire _w4069_ ;
	wire _w4068_ ;
	wire _w4067_ ;
	wire _w4066_ ;
	wire _w4065_ ;
	wire _w4064_ ;
	wire _w4063_ ;
	wire _w4062_ ;
	wire _w4061_ ;
	wire _w4060_ ;
	wire _w4059_ ;
	wire _w4058_ ;
	wire _w4057_ ;
	wire _w4056_ ;
	wire _w4055_ ;
	wire _w4054_ ;
	wire _w4053_ ;
	wire _w4052_ ;
	wire _w4051_ ;
	wire _w4050_ ;
	wire _w4049_ ;
	wire _w4048_ ;
	wire _w4047_ ;
	wire _w4046_ ;
	wire _w4045_ ;
	wire _w4044_ ;
	wire _w4043_ ;
	wire _w4042_ ;
	wire _w4041_ ;
	wire _w4040_ ;
	wire _w4039_ ;
	wire _w4038_ ;
	wire _w4037_ ;
	wire _w4036_ ;
	wire _w4035_ ;
	wire _w4034_ ;
	wire _w4033_ ;
	wire _w4032_ ;
	wire _w4031_ ;
	wire _w4030_ ;
	wire _w4029_ ;
	wire _w4028_ ;
	wire _w4027_ ;
	wire _w4026_ ;
	wire _w4025_ ;
	wire _w4024_ ;
	wire _w4023_ ;
	wire _w4022_ ;
	wire _w4021_ ;
	wire _w4020_ ;
	wire _w4019_ ;
	wire _w4018_ ;
	wire _w4017_ ;
	wire _w4016_ ;
	wire _w4015_ ;
	wire _w4014_ ;
	wire _w4013_ ;
	wire _w4012_ ;
	wire _w4011_ ;
	wire _w4010_ ;
	wire _w4009_ ;
	wire _w4008_ ;
	wire _w4007_ ;
	wire _w4006_ ;
	wire _w4005_ ;
	wire _w4004_ ;
	wire _w4003_ ;
	wire _w4002_ ;
	wire _w4001_ ;
	wire _w4000_ ;
	wire _w3999_ ;
	wire _w3998_ ;
	wire _w3997_ ;
	wire _w3996_ ;
	wire _w3995_ ;
	wire _w3994_ ;
	wire _w3993_ ;
	wire _w3992_ ;
	wire _w3991_ ;
	wire _w3990_ ;
	wire _w3989_ ;
	wire _w3988_ ;
	wire _w3987_ ;
	wire _w3986_ ;
	wire _w3985_ ;
	wire _w3984_ ;
	wire _w3983_ ;
	wire _w3982_ ;
	wire _w3981_ ;
	wire _w3980_ ;
	wire _w3979_ ;
	wire _w3978_ ;
	wire _w3977_ ;
	wire _w3976_ ;
	wire _w3975_ ;
	wire _w3974_ ;
	wire _w3973_ ;
	wire _w3972_ ;
	wire _w3971_ ;
	wire _w3970_ ;
	wire _w3969_ ;
	wire _w3968_ ;
	wire _w3967_ ;
	wire _w3966_ ;
	wire _w3965_ ;
	wire _w3964_ ;
	wire _w3963_ ;
	wire _w3962_ ;
	wire _w3961_ ;
	wire _w3960_ ;
	wire _w3959_ ;
	wire _w3958_ ;
	wire _w3957_ ;
	wire _w3956_ ;
	wire _w3955_ ;
	wire _w3954_ ;
	wire _w3953_ ;
	wire _w3952_ ;
	wire _w3951_ ;
	wire _w3950_ ;
	wire _w3949_ ;
	wire _w3948_ ;
	wire _w3947_ ;
	wire _w3946_ ;
	wire _w3945_ ;
	wire _w3944_ ;
	wire _w3943_ ;
	wire _w3942_ ;
	wire _w3941_ ;
	wire _w3940_ ;
	wire _w3939_ ;
	wire _w3938_ ;
	wire _w3937_ ;
	wire _w3936_ ;
	wire _w3935_ ;
	wire _w3934_ ;
	wire _w3933_ ;
	wire _w3932_ ;
	wire _w3931_ ;
	wire _w3930_ ;
	wire _w3929_ ;
	wire _w3928_ ;
	wire _w3927_ ;
	wire _w3926_ ;
	wire _w3925_ ;
	wire _w3924_ ;
	wire _w3923_ ;
	wire _w3922_ ;
	wire _w3921_ ;
	wire _w3920_ ;
	wire _w3919_ ;
	wire _w3918_ ;
	wire _w3917_ ;
	wire _w3916_ ;
	wire _w3915_ ;
	wire _w3914_ ;
	wire _w3913_ ;
	wire _w3912_ ;
	wire _w3911_ ;
	wire _w3910_ ;
	wire _w3909_ ;
	wire _w3908_ ;
	wire _w3907_ ;
	wire _w3906_ ;
	wire _w3905_ ;
	wire _w3904_ ;
	wire _w3903_ ;
	wire _w3902_ ;
	wire _w3901_ ;
	wire _w3900_ ;
	wire _w3899_ ;
	wire _w3898_ ;
	wire _w3897_ ;
	wire _w3896_ ;
	wire _w3895_ ;
	wire _w3894_ ;
	wire _w3893_ ;
	wire _w3892_ ;
	wire _w3891_ ;
	wire _w3890_ ;
	wire _w3889_ ;
	wire _w3888_ ;
	wire _w3887_ ;
	wire _w3886_ ;
	wire _w3885_ ;
	wire _w3884_ ;
	wire _w3883_ ;
	wire _w3882_ ;
	wire _w3881_ ;
	wire _w3880_ ;
	wire _w3879_ ;
	wire _w3878_ ;
	wire _w3877_ ;
	wire _w3876_ ;
	wire _w3875_ ;
	wire _w3874_ ;
	wire _w3873_ ;
	wire _w3872_ ;
	wire _w3871_ ;
	wire _w3870_ ;
	wire _w3869_ ;
	wire _w3868_ ;
	wire _w3867_ ;
	wire _w3866_ ;
	wire _w3865_ ;
	wire _w3864_ ;
	wire _w3863_ ;
	wire _w3862_ ;
	wire _w3861_ ;
	wire _w3860_ ;
	wire _w3859_ ;
	wire _w3858_ ;
	wire _w3857_ ;
	wire _w3856_ ;
	wire _w3855_ ;
	wire _w3854_ ;
	wire _w3853_ ;
	wire _w3852_ ;
	wire _w3851_ ;
	wire _w3850_ ;
	wire _w3849_ ;
	wire _w3848_ ;
	wire _w3847_ ;
	wire _w3846_ ;
	wire _w3845_ ;
	wire _w3844_ ;
	wire _w3843_ ;
	wire _w3842_ ;
	wire _w3841_ ;
	wire _w3840_ ;
	wire _w3839_ ;
	wire _w3838_ ;
	wire _w3837_ ;
	wire _w3836_ ;
	wire _w3835_ ;
	wire _w3834_ ;
	wire _w3833_ ;
	wire _w3832_ ;
	wire _w3831_ ;
	wire _w3830_ ;
	wire _w3829_ ;
	wire _w3828_ ;
	wire _w3827_ ;
	wire _w3826_ ;
	wire _w3825_ ;
	wire _w3824_ ;
	wire _w3823_ ;
	wire _w3822_ ;
	wire _w3821_ ;
	wire _w3820_ ;
	wire _w3819_ ;
	wire _w3818_ ;
	wire _w3817_ ;
	wire _w3816_ ;
	wire _w3815_ ;
	wire _w3814_ ;
	wire _w3813_ ;
	wire _w3812_ ;
	wire _w3811_ ;
	wire _w3810_ ;
	wire _w3809_ ;
	wire _w3808_ ;
	wire _w3807_ ;
	wire _w3806_ ;
	wire _w3805_ ;
	wire _w3804_ ;
	wire _w3803_ ;
	wire _w3802_ ;
	wire _w3801_ ;
	wire _w3800_ ;
	wire _w3799_ ;
	wire _w3798_ ;
	wire _w3797_ ;
	wire _w3796_ ;
	wire _w3795_ ;
	wire _w3794_ ;
	wire _w3793_ ;
	wire _w3792_ ;
	wire _w3791_ ;
	wire _w3790_ ;
	wire _w3789_ ;
	wire _w3788_ ;
	wire _w3787_ ;
	wire _w3786_ ;
	wire _w3785_ ;
	wire _w3784_ ;
	wire _w3783_ ;
	wire _w3782_ ;
	wire _w3781_ ;
	wire _w3780_ ;
	wire _w3779_ ;
	wire _w3778_ ;
	wire _w3777_ ;
	wire _w3776_ ;
	wire _w3775_ ;
	wire _w3774_ ;
	wire _w3773_ ;
	wire _w3772_ ;
	wire _w3771_ ;
	wire _w3770_ ;
	wire _w3769_ ;
	wire _w3768_ ;
	wire _w3767_ ;
	wire _w3766_ ;
	wire _w3765_ ;
	wire _w3764_ ;
	wire _w3763_ ;
	wire _w3762_ ;
	wire _w3761_ ;
	wire _w3760_ ;
	wire _w3759_ ;
	wire _w3758_ ;
	wire _w3757_ ;
	wire _w3756_ ;
	wire _w3755_ ;
	wire _w3754_ ;
	wire _w3753_ ;
	wire _w3752_ ;
	wire _w3751_ ;
	wire _w3750_ ;
	wire _w3749_ ;
	wire _w3748_ ;
	wire _w3747_ ;
	wire _w3746_ ;
	wire _w3745_ ;
	wire _w3744_ ;
	wire _w3743_ ;
	wire _w3742_ ;
	wire _w3741_ ;
	wire _w3740_ ;
	wire _w3739_ ;
	wire _w3738_ ;
	wire _w3737_ ;
	wire _w3736_ ;
	wire _w3735_ ;
	wire _w3734_ ;
	wire _w3733_ ;
	wire _w3732_ ;
	wire _w3731_ ;
	wire _w3730_ ;
	wire _w3729_ ;
	wire _w3728_ ;
	wire _w3727_ ;
	wire _w3726_ ;
	wire _w3725_ ;
	wire _w3724_ ;
	wire _w3723_ ;
	wire _w3722_ ;
	wire _w3721_ ;
	wire _w3720_ ;
	wire _w3719_ ;
	wire _w3718_ ;
	wire _w3717_ ;
	wire _w3716_ ;
	wire _w3715_ ;
	wire _w3714_ ;
	wire _w3713_ ;
	wire _w3712_ ;
	wire _w3711_ ;
	wire _w3710_ ;
	wire _w3709_ ;
	wire _w3708_ ;
	wire _w3707_ ;
	wire _w3706_ ;
	wire _w3705_ ;
	wire _w3704_ ;
	wire _w3703_ ;
	wire _w3702_ ;
	wire _w3701_ ;
	wire _w3700_ ;
	wire _w3699_ ;
	wire _w3698_ ;
	wire _w3697_ ;
	wire _w3696_ ;
	wire _w3695_ ;
	wire _w3694_ ;
	wire _w3693_ ;
	wire _w3692_ ;
	wire _w3691_ ;
	wire _w3690_ ;
	wire _w3689_ ;
	wire _w3688_ ;
	wire _w3687_ ;
	wire _w3686_ ;
	wire _w3685_ ;
	wire _w3684_ ;
	wire _w3683_ ;
	wire _w3682_ ;
	wire _w3681_ ;
	wire _w3680_ ;
	wire _w3679_ ;
	wire _w3678_ ;
	wire _w3677_ ;
	wire _w3676_ ;
	wire _w3675_ ;
	wire _w3674_ ;
	wire _w3673_ ;
	wire _w3672_ ;
	wire _w3671_ ;
	wire _w3670_ ;
	wire _w3669_ ;
	wire _w3668_ ;
	wire _w3667_ ;
	wire _w3666_ ;
	wire _w3665_ ;
	wire _w3664_ ;
	wire _w3663_ ;
	wire _w3662_ ;
	wire _w3661_ ;
	wire _w3660_ ;
	wire _w3659_ ;
	wire _w3658_ ;
	wire _w3657_ ;
	wire _w3656_ ;
	wire _w3655_ ;
	wire _w3654_ ;
	wire _w3653_ ;
	wire _w3652_ ;
	wire _w3651_ ;
	wire _w3650_ ;
	wire _w3649_ ;
	wire _w3648_ ;
	wire _w3647_ ;
	wire _w3646_ ;
	wire _w3645_ ;
	wire _w3644_ ;
	wire _w3643_ ;
	wire _w3642_ ;
	wire _w3641_ ;
	wire _w3640_ ;
	wire _w3639_ ;
	wire _w3638_ ;
	wire _w3637_ ;
	wire _w3636_ ;
	wire _w3635_ ;
	wire _w3634_ ;
	wire _w3633_ ;
	wire _w3632_ ;
	wire _w3631_ ;
	wire _w3630_ ;
	wire _w3629_ ;
	wire _w3628_ ;
	wire _w3627_ ;
	wire _w3626_ ;
	wire _w3625_ ;
	wire _w3624_ ;
	wire _w3623_ ;
	wire _w3622_ ;
	wire _w3621_ ;
	wire _w3620_ ;
	wire _w3619_ ;
	wire _w3618_ ;
	wire _w3617_ ;
	wire _w3616_ ;
	wire _w3615_ ;
	wire _w3614_ ;
	wire _w3613_ ;
	wire _w3612_ ;
	wire _w3611_ ;
	wire _w3610_ ;
	wire _w3609_ ;
	wire _w3608_ ;
	wire _w3607_ ;
	wire _w3606_ ;
	wire _w3605_ ;
	wire _w3604_ ;
	wire _w3603_ ;
	wire _w3602_ ;
	wire _w3601_ ;
	wire _w3600_ ;
	wire _w3599_ ;
	wire _w3598_ ;
	wire _w3597_ ;
	wire _w3596_ ;
	wire _w3595_ ;
	wire _w3594_ ;
	wire _w3593_ ;
	wire _w3592_ ;
	wire _w3591_ ;
	wire _w3590_ ;
	wire _w3589_ ;
	wire _w3588_ ;
	wire _w3587_ ;
	wire _w3586_ ;
	wire _w3585_ ;
	wire _w3584_ ;
	wire _w3583_ ;
	wire _w3582_ ;
	wire _w3581_ ;
	wire _w3580_ ;
	wire _w3579_ ;
	wire _w3578_ ;
	wire _w3577_ ;
	wire _w3576_ ;
	wire _w3575_ ;
	wire _w3574_ ;
	wire _w3573_ ;
	wire _w3572_ ;
	wire _w3571_ ;
	wire _w3570_ ;
	wire _w3569_ ;
	wire _w3568_ ;
	wire _w3567_ ;
	wire _w3566_ ;
	wire _w3565_ ;
	wire _w3564_ ;
	wire _w3563_ ;
	wire _w3562_ ;
	wire _w3561_ ;
	wire _w3560_ ;
	wire _w3559_ ;
	wire _w3558_ ;
	wire _w3557_ ;
	wire _w3556_ ;
	wire _w3555_ ;
	wire _w3554_ ;
	wire _w3553_ ;
	wire _w3552_ ;
	wire _w3551_ ;
	wire _w3550_ ;
	wire _w3549_ ;
	wire _w3548_ ;
	wire _w3547_ ;
	wire _w3546_ ;
	wire _w3545_ ;
	wire _w3544_ ;
	wire _w3543_ ;
	wire _w3542_ ;
	wire _w3541_ ;
	wire _w3540_ ;
	wire _w3539_ ;
	wire _w3538_ ;
	wire _w3537_ ;
	wire _w3536_ ;
	wire _w3535_ ;
	wire _w3534_ ;
	wire _w3533_ ;
	wire _w3532_ ;
	wire _w3531_ ;
	wire _w3530_ ;
	wire _w3529_ ;
	wire _w3528_ ;
	wire _w3527_ ;
	wire _w3526_ ;
	wire _w3525_ ;
	wire _w3524_ ;
	wire _w3523_ ;
	wire _w3522_ ;
	wire _w3521_ ;
	wire _w3520_ ;
	wire _w3519_ ;
	wire _w3518_ ;
	wire _w3517_ ;
	wire _w3516_ ;
	wire _w3515_ ;
	wire _w3514_ ;
	wire _w3513_ ;
	wire _w3512_ ;
	wire _w3511_ ;
	wire _w3510_ ;
	wire _w3509_ ;
	wire _w3508_ ;
	wire _w3507_ ;
	wire _w3506_ ;
	wire _w3505_ ;
	wire _w3504_ ;
	wire _w3503_ ;
	wire _w3502_ ;
	wire _w3501_ ;
	wire _w3500_ ;
	wire _w3499_ ;
	wire _w3498_ ;
	wire _w3497_ ;
	wire _w3496_ ;
	wire _w3495_ ;
	wire _w3494_ ;
	wire _w3493_ ;
	wire _w3492_ ;
	wire _w3491_ ;
	wire _w3490_ ;
	wire _w3489_ ;
	wire _w3488_ ;
	wire _w3487_ ;
	wire _w3486_ ;
	wire _w3485_ ;
	wire _w3484_ ;
	wire _w3483_ ;
	wire _w3482_ ;
	wire _w3481_ ;
	wire _w3480_ ;
	wire _w3479_ ;
	wire _w3478_ ;
	wire _w3477_ ;
	wire _w3476_ ;
	wire _w3475_ ;
	wire _w3474_ ;
	wire _w3473_ ;
	wire _w3472_ ;
	wire _w3471_ ;
	wire _w3470_ ;
	wire _w3469_ ;
	wire _w3468_ ;
	wire _w3467_ ;
	wire _w3466_ ;
	wire _w3465_ ;
	wire _w3464_ ;
	wire _w3463_ ;
	wire _w3462_ ;
	wire _w3461_ ;
	wire _w3460_ ;
	wire _w3459_ ;
	wire _w3458_ ;
	wire _w3457_ ;
	wire _w3456_ ;
	wire _w3455_ ;
	wire _w3454_ ;
	wire _w3453_ ;
	wire _w3452_ ;
	wire _w3451_ ;
	wire _w3450_ ;
	wire _w3449_ ;
	wire _w3448_ ;
	wire _w3447_ ;
	wire _w3446_ ;
	wire _w3445_ ;
	wire _w3444_ ;
	wire _w3443_ ;
	wire _w3442_ ;
	wire _w3441_ ;
	wire _w3440_ ;
	wire _w3439_ ;
	wire _w3438_ ;
	wire _w3437_ ;
	wire _w3436_ ;
	wire _w3435_ ;
	wire _w3434_ ;
	wire _w3433_ ;
	wire _w3432_ ;
	wire _w3431_ ;
	wire _w3430_ ;
	wire _w3429_ ;
	wire _w3428_ ;
	wire _w3427_ ;
	wire _w3426_ ;
	wire _w3425_ ;
	wire _w3424_ ;
	wire _w3423_ ;
	wire _w3422_ ;
	wire _w3421_ ;
	wire _w3420_ ;
	wire _w3419_ ;
	wire _w3418_ ;
	wire _w3417_ ;
	wire _w3416_ ;
	wire _w3415_ ;
	wire _w3414_ ;
	wire _w3413_ ;
	wire _w3412_ ;
	wire _w3411_ ;
	wire _w3410_ ;
	wire _w3409_ ;
	wire _w3408_ ;
	wire _w3407_ ;
	wire _w3406_ ;
	wire _w3405_ ;
	wire _w3404_ ;
	wire _w3403_ ;
	wire _w3402_ ;
	wire _w3401_ ;
	wire _w3400_ ;
	wire _w3399_ ;
	wire _w3398_ ;
	wire _w3397_ ;
	wire _w3396_ ;
	wire _w3395_ ;
	wire _w3394_ ;
	wire _w3393_ ;
	wire _w3392_ ;
	wire _w3391_ ;
	wire _w3390_ ;
	wire _w3389_ ;
	wire _w3388_ ;
	wire _w3387_ ;
	wire _w3386_ ;
	wire _w3385_ ;
	wire _w3384_ ;
	wire _w3383_ ;
	wire _w3382_ ;
	wire _w3381_ ;
	wire _w3380_ ;
	wire _w3379_ ;
	wire _w3378_ ;
	wire _w3377_ ;
	wire _w3376_ ;
	wire _w3375_ ;
	wire _w3374_ ;
	wire _w3373_ ;
	wire _w3372_ ;
	wire _w3371_ ;
	wire _w3370_ ;
	wire _w3369_ ;
	wire _w3368_ ;
	wire _w3367_ ;
	wire _w3366_ ;
	wire _w3365_ ;
	wire _w3364_ ;
	wire _w3363_ ;
	wire _w3362_ ;
	wire _w3361_ ;
	wire _w3360_ ;
	wire _w3359_ ;
	wire _w3358_ ;
	wire _w3357_ ;
	wire _w3356_ ;
	wire _w3355_ ;
	wire _w3354_ ;
	wire _w3353_ ;
	wire _w3352_ ;
	wire _w3351_ ;
	wire _w3350_ ;
	wire _w3349_ ;
	wire _w3348_ ;
	wire _w3347_ ;
	wire _w3346_ ;
	wire _w3345_ ;
	wire _w3344_ ;
	wire _w3343_ ;
	wire _w3342_ ;
	wire _w3341_ ;
	wire _w3340_ ;
	wire _w3339_ ;
	wire _w3338_ ;
	wire _w3337_ ;
	wire _w3336_ ;
	wire _w3335_ ;
	wire _w3334_ ;
	wire _w3333_ ;
	wire _w3332_ ;
	wire _w3331_ ;
	wire _w3330_ ;
	wire _w3329_ ;
	wire _w3328_ ;
	wire _w3327_ ;
	wire _w3326_ ;
	wire _w3325_ ;
	wire _w3324_ ;
	wire _w3323_ ;
	wire _w3322_ ;
	wire _w3321_ ;
	wire _w3320_ ;
	wire _w3319_ ;
	wire _w3318_ ;
	wire _w3317_ ;
	wire _w3316_ ;
	wire _w3315_ ;
	wire _w3314_ ;
	wire _w3313_ ;
	wire _w3312_ ;
	wire _w3311_ ;
	wire _w3310_ ;
	wire _w3309_ ;
	wire _w3308_ ;
	wire _w3307_ ;
	wire _w3306_ ;
	wire _w3305_ ;
	wire _w3304_ ;
	wire _w3303_ ;
	wire _w3302_ ;
	wire _w3301_ ;
	wire _w3300_ ;
	wire _w3299_ ;
	wire _w3298_ ;
	wire _w3297_ ;
	wire _w3296_ ;
	wire _w3295_ ;
	wire _w3294_ ;
	wire _w3293_ ;
	wire _w3292_ ;
	wire _w3291_ ;
	wire _w3290_ ;
	wire _w3289_ ;
	wire _w3288_ ;
	wire _w3287_ ;
	wire _w3286_ ;
	wire _w3285_ ;
	wire _w3284_ ;
	wire _w3283_ ;
	wire _w3282_ ;
	wire _w3281_ ;
	wire _w3280_ ;
	wire _w3279_ ;
	wire _w3278_ ;
	wire _w3277_ ;
	wire _w3276_ ;
	wire _w3275_ ;
	wire _w3274_ ;
	wire _w3273_ ;
	wire _w3272_ ;
	wire _w3271_ ;
	wire _w3270_ ;
	wire _w3269_ ;
	wire _w3268_ ;
	wire _w3267_ ;
	wire _w3266_ ;
	wire _w3265_ ;
	wire _w3264_ ;
	wire _w3263_ ;
	wire _w3262_ ;
	wire _w3261_ ;
	wire _w3260_ ;
	wire _w3259_ ;
	wire _w3258_ ;
	wire _w3257_ ;
	wire _w3256_ ;
	wire _w3255_ ;
	wire _w3254_ ;
	wire _w3253_ ;
	wire _w3252_ ;
	wire _w3251_ ;
	wire _w3250_ ;
	wire _w3249_ ;
	wire _w3248_ ;
	wire _w3247_ ;
	wire _w3246_ ;
	wire _w3245_ ;
	wire _w3244_ ;
	wire _w3243_ ;
	wire _w3242_ ;
	wire _w3241_ ;
	wire _w3240_ ;
	wire _w3239_ ;
	wire _w3238_ ;
	wire _w3237_ ;
	wire _w3236_ ;
	wire _w3235_ ;
	wire _w3234_ ;
	wire _w3233_ ;
	wire _w3232_ ;
	wire _w3231_ ;
	wire _w3230_ ;
	wire _w3229_ ;
	wire _w3228_ ;
	wire _w3227_ ;
	wire _w3226_ ;
	wire _w3225_ ;
	wire _w3224_ ;
	wire _w3223_ ;
	wire _w3222_ ;
	wire _w3221_ ;
	wire _w3220_ ;
	wire _w3219_ ;
	wire _w3218_ ;
	wire _w3217_ ;
	wire _w3216_ ;
	wire _w3215_ ;
	wire _w3214_ ;
	wire _w3213_ ;
	wire _w3212_ ;
	wire _w3211_ ;
	wire _w3210_ ;
	wire _w3209_ ;
	wire _w3208_ ;
	wire _w3207_ ;
	wire _w3206_ ;
	wire _w3205_ ;
	wire _w3204_ ;
	wire _w3203_ ;
	wire _w3202_ ;
	wire _w3201_ ;
	wire _w3200_ ;
	wire _w3199_ ;
	wire _w3198_ ;
	wire _w3197_ ;
	wire _w3196_ ;
	wire _w3195_ ;
	wire _w3194_ ;
	wire _w3193_ ;
	wire _w3192_ ;
	wire _w3191_ ;
	wire _w3190_ ;
	wire _w3189_ ;
	wire _w3188_ ;
	wire _w3187_ ;
	wire _w3186_ ;
	wire _w3185_ ;
	wire _w3184_ ;
	wire _w3183_ ;
	wire _w3182_ ;
	wire _w3181_ ;
	wire _w3180_ ;
	wire _w3179_ ;
	wire _w3178_ ;
	wire _w3177_ ;
	wire _w3176_ ;
	wire _w3175_ ;
	wire _w3174_ ;
	wire _w3173_ ;
	wire _w3172_ ;
	wire _w3171_ ;
	wire _w3170_ ;
	wire _w3169_ ;
	wire _w3168_ ;
	wire _w3167_ ;
	wire _w3166_ ;
	wire _w3165_ ;
	wire _w3164_ ;
	wire _w3163_ ;
	wire _w3162_ ;
	wire _w3161_ ;
	wire _w3160_ ;
	wire _w3159_ ;
	wire _w3158_ ;
	wire _w3157_ ;
	wire _w3156_ ;
	wire _w3155_ ;
	wire _w3154_ ;
	wire _w3153_ ;
	wire _w3152_ ;
	wire _w3151_ ;
	wire _w3150_ ;
	wire _w3149_ ;
	wire _w3148_ ;
	wire _w3147_ ;
	wire _w3146_ ;
	wire _w3145_ ;
	wire _w3144_ ;
	wire _w3143_ ;
	wire _w3142_ ;
	wire _w3141_ ;
	wire _w3140_ ;
	wire _w3139_ ;
	wire _w3138_ ;
	wire _w3137_ ;
	wire _w3136_ ;
	wire _w3135_ ;
	wire _w3134_ ;
	wire _w3133_ ;
	wire _w3132_ ;
	wire _w3131_ ;
	wire _w3130_ ;
	wire _w3129_ ;
	wire _w3128_ ;
	wire _w3127_ ;
	wire _w3126_ ;
	wire _w3125_ ;
	wire _w3124_ ;
	wire _w3123_ ;
	wire _w3122_ ;
	wire _w3121_ ;
	wire _w3120_ ;
	wire _w3119_ ;
	wire _w3118_ ;
	wire _w3117_ ;
	wire _w3116_ ;
	wire _w3115_ ;
	wire _w3114_ ;
	wire _w3113_ ;
	wire _w3112_ ;
	wire _w3111_ ;
	wire _w3110_ ;
	wire _w3109_ ;
	wire _w3108_ ;
	wire _w3107_ ;
	wire _w3106_ ;
	wire _w3105_ ;
	wire _w3104_ ;
	wire _w3103_ ;
	wire _w3102_ ;
	wire _w3101_ ;
	wire _w3100_ ;
	wire _w3099_ ;
	wire _w3098_ ;
	wire _w3097_ ;
	wire _w3096_ ;
	wire _w3095_ ;
	wire _w3094_ ;
	wire _w3093_ ;
	wire _w3092_ ;
	wire _w3091_ ;
	wire _w3090_ ;
	wire _w3089_ ;
	wire _w3088_ ;
	wire _w3087_ ;
	wire _w3086_ ;
	wire _w3085_ ;
	wire _w3084_ ;
	wire _w3083_ ;
	wire _w3082_ ;
	wire _w3081_ ;
	wire _w3080_ ;
	wire _w3079_ ;
	wire _w3078_ ;
	wire _w3077_ ;
	wire _w3076_ ;
	wire _w3075_ ;
	wire _w3074_ ;
	wire _w3073_ ;
	wire _w3072_ ;
	wire _w3071_ ;
	wire _w3070_ ;
	wire _w3069_ ;
	wire _w3068_ ;
	wire _w3067_ ;
	wire _w3066_ ;
	wire _w3065_ ;
	wire _w3064_ ;
	wire _w3063_ ;
	wire _w3062_ ;
	wire _w3061_ ;
	wire _w3060_ ;
	wire _w3059_ ;
	wire _w3058_ ;
	wire _w3057_ ;
	wire _w3056_ ;
	wire _w3055_ ;
	wire _w3054_ ;
	wire _w3053_ ;
	wire _w3052_ ;
	wire _w3051_ ;
	wire _w3050_ ;
	wire _w3049_ ;
	wire _w3048_ ;
	wire _w3047_ ;
	wire _w3046_ ;
	wire _w3045_ ;
	wire _w3044_ ;
	wire _w3043_ ;
	wire _w3042_ ;
	wire _w3041_ ;
	wire _w3040_ ;
	wire _w3039_ ;
	wire _w3038_ ;
	wire _w3037_ ;
	wire _w3036_ ;
	wire _w3035_ ;
	wire _w3034_ ;
	wire _w3033_ ;
	wire _w3032_ ;
	wire _w3031_ ;
	wire _w3030_ ;
	wire _w3029_ ;
	wire _w3028_ ;
	wire _w3027_ ;
	wire _w3026_ ;
	wire _w3025_ ;
	wire _w3024_ ;
	wire _w3023_ ;
	wire _w3022_ ;
	wire _w3021_ ;
	wire _w3020_ ;
	wire _w3019_ ;
	wire _w3018_ ;
	wire _w3017_ ;
	wire _w3016_ ;
	wire _w3015_ ;
	wire _w3014_ ;
	wire _w3013_ ;
	wire _w3012_ ;
	wire _w3011_ ;
	wire _w3010_ ;
	wire _w3009_ ;
	wire _w3008_ ;
	wire _w3007_ ;
	wire _w3006_ ;
	wire _w3005_ ;
	wire _w3004_ ;
	wire _w3003_ ;
	wire _w3002_ ;
	wire _w3001_ ;
	wire _w3000_ ;
	wire _w2999_ ;
	wire _w2998_ ;
	wire _w2997_ ;
	wire _w2996_ ;
	wire _w2995_ ;
	wire _w2994_ ;
	wire _w2993_ ;
	wire _w2992_ ;
	wire _w2991_ ;
	wire _w2990_ ;
	wire _w2989_ ;
	wire _w2988_ ;
	wire _w2987_ ;
	wire _w2986_ ;
	wire _w2985_ ;
	wire _w2984_ ;
	wire _w2983_ ;
	wire _w2982_ ;
	wire _w2981_ ;
	wire _w2980_ ;
	wire _w2979_ ;
	wire _w2978_ ;
	wire _w2977_ ;
	wire _w2976_ ;
	wire _w2975_ ;
	wire _w2974_ ;
	wire _w2973_ ;
	wire _w2972_ ;
	wire _w2971_ ;
	wire _w2970_ ;
	wire _w2969_ ;
	wire _w2968_ ;
	wire _w2967_ ;
	wire _w2966_ ;
	wire _w2965_ ;
	wire _w2964_ ;
	wire _w2963_ ;
	wire _w2962_ ;
	wire _w2961_ ;
	wire _w2960_ ;
	wire _w2959_ ;
	wire _w2958_ ;
	wire _w2957_ ;
	wire _w2956_ ;
	wire _w2955_ ;
	wire _w2954_ ;
	wire _w2953_ ;
	wire _w2952_ ;
	wire _w2951_ ;
	wire _w2950_ ;
	wire _w2949_ ;
	wire _w2948_ ;
	wire _w2947_ ;
	wire _w2946_ ;
	wire _w2945_ ;
	wire _w2944_ ;
	wire _w2943_ ;
	wire _w2942_ ;
	wire _w2941_ ;
	wire _w2940_ ;
	wire _w2939_ ;
	wire _w2938_ ;
	wire _w2937_ ;
	wire _w2936_ ;
	wire _w2935_ ;
	wire _w2934_ ;
	wire _w2933_ ;
	wire _w2932_ ;
	wire _w2931_ ;
	wire _w2930_ ;
	wire _w2929_ ;
	wire _w2928_ ;
	wire _w2927_ ;
	wire _w2926_ ;
	wire _w2925_ ;
	wire _w2924_ ;
	wire _w2923_ ;
	wire _w2922_ ;
	wire _w2921_ ;
	wire _w2920_ ;
	wire _w2919_ ;
	wire _w2918_ ;
	wire _w2917_ ;
	wire _w2916_ ;
	wire _w2915_ ;
	wire _w2914_ ;
	wire _w2913_ ;
	wire _w2912_ ;
	wire _w2911_ ;
	wire _w2910_ ;
	wire _w2909_ ;
	wire _w2908_ ;
	wire _w2907_ ;
	wire _w2906_ ;
	wire _w2905_ ;
	wire _w2904_ ;
	wire _w2903_ ;
	wire _w2902_ ;
	wire _w2901_ ;
	wire _w2900_ ;
	wire _w2899_ ;
	wire _w2898_ ;
	wire _w2897_ ;
	wire _w2896_ ;
	wire _w2895_ ;
	wire _w2894_ ;
	wire _w2893_ ;
	wire _w2892_ ;
	wire _w2891_ ;
	wire _w2890_ ;
	wire _w2889_ ;
	wire _w2888_ ;
	wire _w2887_ ;
	wire _w2886_ ;
	wire _w2885_ ;
	wire _w2884_ ;
	wire _w2883_ ;
	wire _w2882_ ;
	wire _w2881_ ;
	wire _w2880_ ;
	wire _w2879_ ;
	wire _w2878_ ;
	wire _w2877_ ;
	wire _w2876_ ;
	wire _w2875_ ;
	wire _w2874_ ;
	wire _w2873_ ;
	wire _w2872_ ;
	wire _w2871_ ;
	wire _w2870_ ;
	wire _w2869_ ;
	wire _w2868_ ;
	wire _w2867_ ;
	wire _w2866_ ;
	wire _w2865_ ;
	wire _w2864_ ;
	wire _w2863_ ;
	wire _w2862_ ;
	wire _w2861_ ;
	wire _w2860_ ;
	wire _w2859_ ;
	wire _w2858_ ;
	wire _w2857_ ;
	wire _w2856_ ;
	wire _w2855_ ;
	wire _w2854_ ;
	wire _w2853_ ;
	wire _w2852_ ;
	wire _w2851_ ;
	wire _w2850_ ;
	wire _w2849_ ;
	wire _w2848_ ;
	wire _w2847_ ;
	wire _w2846_ ;
	wire _w2845_ ;
	wire _w2844_ ;
	wire _w2843_ ;
	wire _w2842_ ;
	wire _w2841_ ;
	wire _w2840_ ;
	wire _w2839_ ;
	wire _w2838_ ;
	wire _w2837_ ;
	wire _w2836_ ;
	wire _w2835_ ;
	wire _w2834_ ;
	wire _w2833_ ;
	wire _w2832_ ;
	wire _w2831_ ;
	wire _w2830_ ;
	wire _w2829_ ;
	wire _w2828_ ;
	wire _w2827_ ;
	wire _w2826_ ;
	wire _w2825_ ;
	wire _w2824_ ;
	wire _w2823_ ;
	wire _w2822_ ;
	wire _w2821_ ;
	wire _w2820_ ;
	wire _w2819_ ;
	wire _w1570_ ;
	wire _w1569_ ;
	wire _w1568_ ;
	wire _w1567_ ;
	wire _w1566_ ;
	wire _w1565_ ;
	wire _w1564_ ;
	wire _w1563_ ;
	wire _w1562_ ;
	wire _w1561_ ;
	wire _w1560_ ;
	wire _w1559_ ;
	wire _w1558_ ;
	wire _w1557_ ;
	wire _w1556_ ;
	wire _w1555_ ;
	wire _w1554_ ;
	wire _w1553_ ;
	wire _w1552_ ;
	wire _w1551_ ;
	wire _w1550_ ;
	wire _w1549_ ;
	wire _w1548_ ;
	wire _w1547_ ;
	wire _w1546_ ;
	wire _w1545_ ;
	wire _w1544_ ;
	wire _w1543_ ;
	wire _w1542_ ;
	wire _w1541_ ;
	wire _w1540_ ;
	wire _w1539_ ;
	wire _w1538_ ;
	wire _w1537_ ;
	wire _w1536_ ;
	wire _w1535_ ;
	wire _w1534_ ;
	wire _w1533_ ;
	wire _w1532_ ;
	wire _w1531_ ;
	wire _w1530_ ;
	wire _w1529_ ;
	wire _w1528_ ;
	wire _w1527_ ;
	wire _w1526_ ;
	wire _w1525_ ;
	wire _w1524_ ;
	wire _w1523_ ;
	wire _w1522_ ;
	wire _w1521_ ;
	wire _w1520_ ;
	wire _w1519_ ;
	wire _w1518_ ;
	wire _w1517_ ;
	wire _w1516_ ;
	wire _w1515_ ;
	wire _w1514_ ;
	wire _w1513_ ;
	wire _w1512_ ;
	wire _w1511_ ;
	wire _w1510_ ;
	wire _w1509_ ;
	wire _w1508_ ;
	wire _w1507_ ;
	wire _w1506_ ;
	wire _w1505_ ;
	wire _w1504_ ;
	wire _w1503_ ;
	wire _w1502_ ;
	wire _w1501_ ;
	wire _w1500_ ;
	wire _w1499_ ;
	wire _w1498_ ;
	wire _w1497_ ;
	wire _w1496_ ;
	wire _w1495_ ;
	wire _w1494_ ;
	wire _w1493_ ;
	wire _w1492_ ;
	wire _w1491_ ;
	wire _w1490_ ;
	wire _w1489_ ;
	wire _w1488_ ;
	wire _w1487_ ;
	wire _w1486_ ;
	wire _w1485_ ;
	wire _w1484_ ;
	wire _w1483_ ;
	wire _w1482_ ;
	wire _w1481_ ;
	wire _w1480_ ;
	wire _w1479_ ;
	wire _w1478_ ;
	wire _w1477_ ;
	wire _w1476_ ;
	wire _w1475_ ;
	wire _w1474_ ;
	wire _w1473_ ;
	wire _w1472_ ;
	wire _w1471_ ;
	wire _w1470_ ;
	wire _w1469_ ;
	wire _w1468_ ;
	wire _w1467_ ;
	wire _w1466_ ;
	wire _w1465_ ;
	wire _w1464_ ;
	wire _w1463_ ;
	wire _w1462_ ;
	wire _w1461_ ;
	wire _w1460_ ;
	wire _w1459_ ;
	wire _w1458_ ;
	wire _w1457_ ;
	wire _w1456_ ;
	wire _w1455_ ;
	wire _w1454_ ;
	wire _w1453_ ;
	wire _w1452_ ;
	wire _w1451_ ;
	wire _w1450_ ;
	wire _w1449_ ;
	wire _w1448_ ;
	wire _w1447_ ;
	wire _w1446_ ;
	wire _w1445_ ;
	wire _w1444_ ;
	wire _w1443_ ;
	wire _w1442_ ;
	wire _w1441_ ;
	wire _w1440_ ;
	wire _w1439_ ;
	wire _w1438_ ;
	wire _w1437_ ;
	wire _w1436_ ;
	wire _w1435_ ;
	wire _w1434_ ;
	wire _w1433_ ;
	wire _w1432_ ;
	wire _w1431_ ;
	wire _w1430_ ;
	wire _w1429_ ;
	wire _w1428_ ;
	wire _w1427_ ;
	wire _w1426_ ;
	wire _w1425_ ;
	wire _w1424_ ;
	wire _w1423_ ;
	wire _w1422_ ;
	wire _w1421_ ;
	wire _w1420_ ;
	wire _w1419_ ;
	wire _w1418_ ;
	wire _w1417_ ;
	wire _w1416_ ;
	wire _w1415_ ;
	wire _w1414_ ;
	wire _w1413_ ;
	wire _w1412_ ;
	wire _w1411_ ;
	wire _w1410_ ;
	wire _w1409_ ;
	wire _w1408_ ;
	wire _w1407_ ;
	wire _w1406_ ;
	wire _w1405_ ;
	wire _w1404_ ;
	wire _w1403_ ;
	wire _w1402_ ;
	wire _w1401_ ;
	wire _w1400_ ;
	wire _w1399_ ;
	wire _w1398_ ;
	wire _w1397_ ;
	wire _w1396_ ;
	wire _w1395_ ;
	wire _w1394_ ;
	wire _w1393_ ;
	wire _w1392_ ;
	wire _w1391_ ;
	wire _w1390_ ;
	wire _w1389_ ;
	wire _w1388_ ;
	wire _w1387_ ;
	wire _w1386_ ;
	wire _w1385_ ;
	wire _w1384_ ;
	wire _w1383_ ;
	wire _w1382_ ;
	wire _w1381_ ;
	wire _w1380_ ;
	wire _w1379_ ;
	wire _w1378_ ;
	wire _w1377_ ;
	wire _w1376_ ;
	wire _w1375_ ;
	wire _w1374_ ;
	wire _w1373_ ;
	wire _w1372_ ;
	wire _w1371_ ;
	wire _w1370_ ;
	wire _w1369_ ;
	wire _w1368_ ;
	wire _w1367_ ;
	wire _w1366_ ;
	wire _w1365_ ;
	wire _w1364_ ;
	wire _w1363_ ;
	wire _w1362_ ;
	wire _w1361_ ;
	wire _w1360_ ;
	wire _w1359_ ;
	wire _w1358_ ;
	wire _w1357_ ;
	wire _w1356_ ;
	wire _w1355_ ;
	wire _w1354_ ;
	wire _w1353_ ;
	wire _w1352_ ;
	wire _w1351_ ;
	wire _w1350_ ;
	wire _w1349_ ;
	wire _w1348_ ;
	wire _w1347_ ;
	wire _w1346_ ;
	wire _w1345_ ;
	wire _w1344_ ;
	wire _w1343_ ;
	wire _w1342_ ;
	wire _w1341_ ;
	wire _w1340_ ;
	wire _w1339_ ;
	wire _w1338_ ;
	wire _w1337_ ;
	wire _w1336_ ;
	wire _w1335_ ;
	wire _w1334_ ;
	wire _w1333_ ;
	wire _w1332_ ;
	wire _w1331_ ;
	wire _w1330_ ;
	wire _w1329_ ;
	wire _w1328_ ;
	wire _w1327_ ;
	wire _w1326_ ;
	wire _w1325_ ;
	wire _w1324_ ;
	wire _w1323_ ;
	wire _w1322_ ;
	wire _w1321_ ;
	wire _w1320_ ;
	wire _w1319_ ;
	wire _w1318_ ;
	wire _w1317_ ;
	wire _w1316_ ;
	wire _w1315_ ;
	wire _w1314_ ;
	wire _w1313_ ;
	wire _w1312_ ;
	wire _w1311_ ;
	wire _w1310_ ;
	wire _w1309_ ;
	wire _w1308_ ;
	wire _w1307_ ;
	wire _w1306_ ;
	wire _w1305_ ;
	wire _w1304_ ;
	wire _w1303_ ;
	wire _w1302_ ;
	wire _w1301_ ;
	wire _w1300_ ;
	wire _w1299_ ;
	wire _w1298_ ;
	wire _w1297_ ;
	wire _w1296_ ;
	wire _w1295_ ;
	wire _w1294_ ;
	wire _w1293_ ;
	wire _w1292_ ;
	wire _w1291_ ;
	wire _w1290_ ;
	wire _w1289_ ;
	wire _w1288_ ;
	wire _w1287_ ;
	wire _w1286_ ;
	wire _w1285_ ;
	wire _w1284_ ;
	wire _w1283_ ;
	wire _w1282_ ;
	wire _w1281_ ;
	wire _w1280_ ;
	wire _w1279_ ;
	wire _w1278_ ;
	wire _w1277_ ;
	wire _w1276_ ;
	wire _w1275_ ;
	wire _w1274_ ;
	wire _w1273_ ;
	wire _w1272_ ;
	wire _w1271_ ;
	wire _w1270_ ;
	wire _w1269_ ;
	wire _w1268_ ;
	wire _w1267_ ;
	wire _w1266_ ;
	wire _w1265_ ;
	wire _w1264_ ;
	wire _w1263_ ;
	wire _w1262_ ;
	wire _w1261_ ;
	wire _w1260_ ;
	wire _w1259_ ;
	wire _w1258_ ;
	wire _w1257_ ;
	wire _w1256_ ;
	wire _w1255_ ;
	wire _w1254_ ;
	wire _w1253_ ;
	wire _w1252_ ;
	wire _w1251_ ;
	wire _w1250_ ;
	wire _w1249_ ;
	wire _w1248_ ;
	wire _w1247_ ;
	wire _w1246_ ;
	wire _w1245_ ;
	wire _w1244_ ;
	wire _w1243_ ;
	wire _w1242_ ;
	wire _w1241_ ;
	wire _w1240_ ;
	wire _w1239_ ;
	wire _w1238_ ;
	wire _w1237_ ;
	wire _w1236_ ;
	wire _w1235_ ;
	wire _w1234_ ;
	wire _w1233_ ;
	wire _w1232_ ;
	wire _w1231_ ;
	wire _w1230_ ;
	wire _w1229_ ;
	wire _w1228_ ;
	wire _w1227_ ;
	wire _w1226_ ;
	wire _w1225_ ;
	wire _w1224_ ;
	wire _w1223_ ;
	wire _w1222_ ;
	wire _w1221_ ;
	wire _w1220_ ;
	wire _w1219_ ;
	wire _w1218_ ;
	wire _w1217_ ;
	wire _w1216_ ;
	wire _w1215_ ;
	wire _w1214_ ;
	wire _w1213_ ;
	wire _w1212_ ;
	wire _w1211_ ;
	wire _w1210_ ;
	wire _w1209_ ;
	wire _w1208_ ;
	wire _w1207_ ;
	wire _w1206_ ;
	wire _w1205_ ;
	wire _w1204_ ;
	wire _w1203_ ;
	wire _w1202_ ;
	wire _w1201_ ;
	wire _w1200_ ;
	wire _w1199_ ;
	wire _w1198_ ;
	wire _w1197_ ;
	wire _w1196_ ;
	wire _w1195_ ;
	wire _w1194_ ;
	wire _w1193_ ;
	wire _w1192_ ;
	wire _w1191_ ;
	wire _w1190_ ;
	wire _w1189_ ;
	wire _w1188_ ;
	wire _w1187_ ;
	wire _w1186_ ;
	wire _w1185_ ;
	wire _w1184_ ;
	wire _w1183_ ;
	wire _w1182_ ;
	wire _w1181_ ;
	wire _w1180_ ;
	wire _w1179_ ;
	wire _w1178_ ;
	wire _w1177_ ;
	wire _w1176_ ;
	wire _w1175_ ;
	wire _w1174_ ;
	wire _w1173_ ;
	wire _w1172_ ;
	wire _w1171_ ;
	wire _w1170_ ;
	wire _w1169_ ;
	wire _w1168_ ;
	wire _w1167_ ;
	wire _w1166_ ;
	wire _w1165_ ;
	wire _w1164_ ;
	wire _w1163_ ;
	wire _w1162_ ;
	wire _w1161_ ;
	wire _w1160_ ;
	wire _w1159_ ;
	wire _w1158_ ;
	wire _w1157_ ;
	wire _w1156_ ;
	wire _w1155_ ;
	wire _w1154_ ;
	wire _w1153_ ;
	wire _w1152_ ;
	wire _w1151_ ;
	wire _w1150_ ;
	wire _w1149_ ;
	wire _w1148_ ;
	wire _w1147_ ;
	wire _w1146_ ;
	wire _w1145_ ;
	wire _w1144_ ;
	wire _w1143_ ;
	wire _w1142_ ;
	wire _w1141_ ;
	wire _w1140_ ;
	wire _w1139_ ;
	wire _w1138_ ;
	wire _w1137_ ;
	wire _w1136_ ;
	wire _w1135_ ;
	wire _w1134_ ;
	wire _w1133_ ;
	wire _w1132_ ;
	wire _w1131_ ;
	wire _w1130_ ;
	wire _w1129_ ;
	wire _w1128_ ;
	wire _w1127_ ;
	wire _w1126_ ;
	wire _w1125_ ;
	wire _w1124_ ;
	wire _w1123_ ;
	wire _w1122_ ;
	wire _w1121_ ;
	wire _w1120_ ;
	wire _w1119_ ;
	wire _w1118_ ;
	wire _w1117_ ;
	wire _w1116_ ;
	wire _w1115_ ;
	wire _w1114_ ;
	wire _w1113_ ;
	wire _w1112_ ;
	wire _w1111_ ;
	wire _w1110_ ;
	wire _w1109_ ;
	wire _w1108_ ;
	wire _w1107_ ;
	wire _w1106_ ;
	wire _w1105_ ;
	wire _w1104_ ;
	wire _w1103_ ;
	wire _w1102_ ;
	wire _w1101_ ;
	wire _w1100_ ;
	wire _w1099_ ;
	wire _w1098_ ;
	wire _w1097_ ;
	wire _w1096_ ;
	wire _w1095_ ;
	wire _w1094_ ;
	wire _w1093_ ;
	wire _w1092_ ;
	wire _w1091_ ;
	wire _w1090_ ;
	wire _w1089_ ;
	wire _w1088_ ;
	wire _w1087_ ;
	wire _w1086_ ;
	wire _w1085_ ;
	wire _w1084_ ;
	wire _w1083_ ;
	wire _w1082_ ;
	wire _w1081_ ;
	wire _w1080_ ;
	wire _w1079_ ;
	wire _w1078_ ;
	wire _w1077_ ;
	wire _w1076_ ;
	wire _w1075_ ;
	wire _w1074_ ;
	wire _w1073_ ;
	wire _w1072_ ;
	wire _w1071_ ;
	wire _w1070_ ;
	wire _w1069_ ;
	wire _w1068_ ;
	wire _w1067_ ;
	wire _w1066_ ;
	wire _w1065_ ;
	wire _w1064_ ;
	wire _w1063_ ;
	wire _w1062_ ;
	wire _w1061_ ;
	wire _w1060_ ;
	wire _w1059_ ;
	wire _w1058_ ;
	wire _w1057_ ;
	wire _w1056_ ;
	wire _w1055_ ;
	wire _w1054_ ;
	wire _w1053_ ;
	wire _w1052_ ;
	wire _w1051_ ;
	wire _w1050_ ;
	wire _w1049_ ;
	wire _w1048_ ;
	wire _w1047_ ;
	wire _w1046_ ;
	wire _w1045_ ;
	wire _w1044_ ;
	wire _w1043_ ;
	wire _w1042_ ;
	wire _w1041_ ;
	wire _w1040_ ;
	wire _w1039_ ;
	wire _w1038_ ;
	wire _w1037_ ;
	wire _w1036_ ;
	wire _w1035_ ;
	wire _w1034_ ;
	wire _w1033_ ;
	wire _w1032_ ;
	wire _w1031_ ;
	wire _w1030_ ;
	wire _w1029_ ;
	wire _w1028_ ;
	wire _w1027_ ;
	wire _w1026_ ;
	wire _w1025_ ;
	wire _w1024_ ;
	wire _w1023_ ;
	wire _w1022_ ;
	wire _w1021_ ;
	wire _w1020_ ;
	wire _w1019_ ;
	wire _w1018_ ;
	wire _w1017_ ;
	wire _w1016_ ;
	wire _w1015_ ;
	wire _w1014_ ;
	wire _w1013_ ;
	wire _w1012_ ;
	wire _w1011_ ;
	wire _w1010_ ;
	wire _w1009_ ;
	wire _w1008_ ;
	wire _w1007_ ;
	wire _w1006_ ;
	wire _w1005_ ;
	wire _w1004_ ;
	wire _w1003_ ;
	wire _w718_ ;
	wire _w717_ ;
	wire _w716_ ;
	wire _w715_ ;
	wire _w714_ ;
	wire _w713_ ;
	wire _w712_ ;
	wire _w711_ ;
	wire _w710_ ;
	wire _w709_ ;
	wire _w708_ ;
	wire _w707_ ;
	wire _w706_ ;
	wire _w705_ ;
	wire _w704_ ;
	wire _w703_ ;
	wire _w702_ ;
	wire _w701_ ;
	wire _w700_ ;
	wire _w699_ ;
	wire _w698_ ;
	wire _w697_ ;
	wire _w696_ ;
	wire _w695_ ;
	wire _w694_ ;
	wire _w693_ ;
	wire _w692_ ;
	wire _w691_ ;
	wire _w690_ ;
	wire _w689_ ;
	wire _w688_ ;
	wire _w687_ ;
	wire _w686_ ;
	wire _w685_ ;
	wire _w684_ ;
	wire _w683_ ;
	wire _w682_ ;
	wire _w681_ ;
	wire _w680_ ;
	wire _w679_ ;
	wire _w678_ ;
	wire _w677_ ;
	wire _w676_ ;
	wire _w675_ ;
	wire _w674_ ;
	wire _w673_ ;
	wire _w672_ ;
	wire _w671_ ;
	wire _w670_ ;
	wire _w669_ ;
	wire _w668_ ;
	wire _w667_ ;
	wire _w666_ ;
	wire _w665_ ;
	wire _w664_ ;
	wire _w663_ ;
	wire _w662_ ;
	wire _w661_ ;
	wire _w660_ ;
	wire _w659_ ;
	wire _w658_ ;
	wire _w657_ ;
	wire _w656_ ;
	wire _w655_ ;
	wire _w654_ ;
	wire _w653_ ;
	wire _w652_ ;
	wire _w651_ ;
	wire _w650_ ;
	wire _w649_ ;
	wire _w648_ ;
	wire _w647_ ;
	wire _w646_ ;
	wire _w645_ ;
	wire _w644_ ;
	wire _w643_ ;
	wire _w642_ ;
	wire _w641_ ;
	wire _w640_ ;
	wire _w639_ ;
	wire _w638_ ;
	wire _w637_ ;
	wire _w636_ ;
	wire _w635_ ;
	wire _w634_ ;
	wire _w633_ ;
	wire _w632_ ;
	wire _w631_ ;
	wire _w630_ ;
	wire _w629_ ;
	wire _w628_ ;
	wire _w627_ ;
	wire _w626_ ;
	wire _w625_ ;
	wire _w624_ ;
	wire _w623_ ;
	wire _w622_ ;
	wire _w621_ ;
	wire _w620_ ;
	wire _w619_ ;
	wire _w618_ ;
	wire _w617_ ;
	wire _w616_ ;
	wire _w615_ ;
	wire _w614_ ;
	wire _w613_ ;
	wire _w612_ ;
	wire _w611_ ;
	wire _w610_ ;
	wire _w609_ ;
	wire _w608_ ;
	wire _w607_ ;
	wire _w606_ ;
	wire _w605_ ;
	wire _w604_ ;
	wire _w603_ ;
	wire _w602_ ;
	wire _w601_ ;
	wire _w600_ ;
	wire _w599_ ;
	wire _w598_ ;
	wire _w597_ ;
	wire _w596_ ;
	wire _w595_ ;
	wire _w594_ ;
	wire _w593_ ;
	wire _w592_ ;
	wire _w591_ ;
	wire _w590_ ;
	wire _w589_ ;
	wire _w520_ ;
	wire _w519_ ;
	wire _w518_ ;
	wire _w517_ ;
	wire _w516_ ;
	wire _w515_ ;
	wire _w514_ ;
	wire _w513_ ;
	wire _w512_ ;
	wire _w511_ ;
	wire _w510_ ;
	wire _w509_ ;
	wire _w508_ ;
	wire _w507_ ;
	wire _w506_ ;
	wire _w505_ ;
	wire _w504_ ;
	wire _w503_ ;
	wire _w502_ ;
	wire _w501_ ;
	wire _w500_ ;
	wire _w499_ ;
	wire _w498_ ;
	wire _w497_ ;
	wire _w496_ ;
	wire _w495_ ;
	wire _w494_ ;
	wire _w493_ ;
	wire _w492_ ;
	wire _w491_ ;
	wire _w474_ ;
	wire _w473_ ;
	wire _w472_ ;
	wire _w471_ ;
	wire _w470_ ;
	wire _w469_ ;
	wire _w468_ ;
	wire _w467_ ;
	wire _w466_ ;
	wire _w465_ ;
	wire _w464_ ;
	wire _w463_ ;
	wire _w462_ ;
	wire _w475_ ;
	wire _w476_ ;
	wire _w477_ ;
	wire _w478_ ;
	wire _w479_ ;
	wire _w480_ ;
	wire _w481_ ;
	wire _w482_ ;
	wire _w483_ ;
	wire _w484_ ;
	wire _w485_ ;
	wire _w486_ ;
	wire _w487_ ;
	wire _w488_ ;
	wire _w489_ ;
	wire _w490_ ;
	wire _w521_ ;
	wire _w522_ ;
	wire _w523_ ;
	wire _w524_ ;
	wire _w525_ ;
	wire _w526_ ;
	wire _w527_ ;
	wire _w528_ ;
	wire _w529_ ;
	wire _w530_ ;
	wire _w531_ ;
	wire _w532_ ;
	wire _w533_ ;
	wire _w534_ ;
	wire _w535_ ;
	wire _w536_ ;
	wire _w537_ ;
	wire _w538_ ;
	wire _w539_ ;
	wire _w540_ ;
	wire _w541_ ;
	wire _w542_ ;
	wire _w543_ ;
	wire _w544_ ;
	wire _w545_ ;
	wire _w546_ ;
	wire _w547_ ;
	wire _w548_ ;
	wire _w549_ ;
	wire _w550_ ;
	wire _w551_ ;
	wire _w552_ ;
	wire _w553_ ;
	wire _w554_ ;
	wire _w555_ ;
	wire _w556_ ;
	wire _w557_ ;
	wire _w558_ ;
	wire _w559_ ;
	wire _w560_ ;
	wire _w561_ ;
	wire _w562_ ;
	wire _w563_ ;
	wire _w564_ ;
	wire _w565_ ;
	wire _w566_ ;
	wire _w567_ ;
	wire _w568_ ;
	wire _w569_ ;
	wire _w570_ ;
	wire _w571_ ;
	wire _w572_ ;
	wire _w573_ ;
	wire _w574_ ;
	wire _w575_ ;
	wire _w576_ ;
	wire _w577_ ;
	wire _w578_ ;
	wire _w579_ ;
	wire _w580_ ;
	wire _w581_ ;
	wire _w582_ ;
	wire _w583_ ;
	wire _w584_ ;
	wire _w585_ ;
	wire _w586_ ;
	wire _w587_ ;
	wire _w588_ ;
	wire _w719_ ;
	wire _w720_ ;
	wire _w721_ ;
	wire _w722_ ;
	wire _w723_ ;
	wire _w724_ ;
	wire _w725_ ;
	wire _w726_ ;
	wire _w727_ ;
	wire _w728_ ;
	wire _w729_ ;
	wire _w730_ ;
	wire _w731_ ;
	wire _w732_ ;
	wire _w733_ ;
	wire _w734_ ;
	wire _w735_ ;
	wire _w736_ ;
	wire _w737_ ;
	wire _w738_ ;
	wire _w739_ ;
	wire _w740_ ;
	wire _w741_ ;
	wire _w742_ ;
	wire _w743_ ;
	wire _w744_ ;
	wire _w745_ ;
	wire _w746_ ;
	wire _w747_ ;
	wire _w748_ ;
	wire _w749_ ;
	wire _w750_ ;
	wire _w751_ ;
	wire _w752_ ;
	wire _w753_ ;
	wire _w754_ ;
	wire _w755_ ;
	wire _w756_ ;
	wire _w757_ ;
	wire _w758_ ;
	wire _w759_ ;
	wire _w760_ ;
	wire _w761_ ;
	wire _w762_ ;
	wire _w763_ ;
	wire _w764_ ;
	wire _w765_ ;
	wire _w766_ ;
	wire _w767_ ;
	wire _w768_ ;
	wire _w769_ ;
	wire _w770_ ;
	wire _w771_ ;
	wire _w772_ ;
	wire _w773_ ;
	wire _w774_ ;
	wire _w775_ ;
	wire _w776_ ;
	wire _w777_ ;
	wire _w778_ ;
	wire _w779_ ;
	wire _w780_ ;
	wire _w781_ ;
	wire _w782_ ;
	wire _w783_ ;
	wire _w784_ ;
	wire _w785_ ;
	wire _w786_ ;
	wire _w787_ ;
	wire _w788_ ;
	wire _w789_ ;
	wire _w790_ ;
	wire _w791_ ;
	wire _w792_ ;
	wire _w793_ ;
	wire _w794_ ;
	wire _w795_ ;
	wire _w796_ ;
	wire _w797_ ;
	wire _w798_ ;
	wire _w799_ ;
	wire _w800_ ;
	wire _w801_ ;
	wire _w802_ ;
	wire _w803_ ;
	wire _w804_ ;
	wire _w805_ ;
	wire _w806_ ;
	wire _w807_ ;
	wire _w808_ ;
	wire _w809_ ;
	wire _w810_ ;
	wire _w811_ ;
	wire _w812_ ;
	wire _w813_ ;
	wire _w814_ ;
	wire _w815_ ;
	wire _w816_ ;
	wire _w817_ ;
	wire _w818_ ;
	wire _w819_ ;
	wire _w820_ ;
	wire _w821_ ;
	wire _w822_ ;
	wire _w823_ ;
	wire _w824_ ;
	wire _w825_ ;
	wire _w826_ ;
	wire _w827_ ;
	wire _w828_ ;
	wire _w829_ ;
	wire _w830_ ;
	wire _w831_ ;
	wire _w832_ ;
	wire _w833_ ;
	wire _w834_ ;
	wire _w835_ ;
	wire _w836_ ;
	wire _w837_ ;
	wire _w838_ ;
	wire _w839_ ;
	wire _w840_ ;
	wire _w841_ ;
	wire _w842_ ;
	wire _w843_ ;
	wire _w844_ ;
	wire _w845_ ;
	wire _w846_ ;
	wire _w847_ ;
	wire _w848_ ;
	wire _w849_ ;
	wire _w850_ ;
	wire _w851_ ;
	wire _w852_ ;
	wire _w853_ ;
	wire _w854_ ;
	wire _w855_ ;
	wire _w856_ ;
	wire _w857_ ;
	wire _w858_ ;
	wire _w859_ ;
	wire _w860_ ;
	wire _w861_ ;
	wire _w862_ ;
	wire _w863_ ;
	wire _w864_ ;
	wire _w865_ ;
	wire _w866_ ;
	wire _w867_ ;
	wire _w868_ ;
	wire _w869_ ;
	wire _w870_ ;
	wire _w871_ ;
	wire _w872_ ;
	wire _w873_ ;
	wire _w874_ ;
	wire _w875_ ;
	wire _w876_ ;
	wire _w877_ ;
	wire _w878_ ;
	wire _w879_ ;
	wire _w880_ ;
	wire _w881_ ;
	wire _w882_ ;
	wire _w883_ ;
	wire _w884_ ;
	wire _w885_ ;
	wire _w886_ ;
	wire _w887_ ;
	wire _w888_ ;
	wire _w889_ ;
	wire _w890_ ;
	wire _w891_ ;
	wire _w892_ ;
	wire _w893_ ;
	wire _w894_ ;
	wire _w895_ ;
	wire _w896_ ;
	wire _w897_ ;
	wire _w898_ ;
	wire _w899_ ;
	wire _w900_ ;
	wire _w901_ ;
	wire _w902_ ;
	wire _w903_ ;
	wire _w904_ ;
	wire _w905_ ;
	wire _w906_ ;
	wire _w907_ ;
	wire _w908_ ;
	wire _w909_ ;
	wire _w910_ ;
	wire _w911_ ;
	wire _w912_ ;
	wire _w913_ ;
	wire _w914_ ;
	wire _w915_ ;
	wire _w916_ ;
	wire _w917_ ;
	wire _w918_ ;
	wire _w919_ ;
	wire _w920_ ;
	wire _w921_ ;
	wire _w922_ ;
	wire _w923_ ;
	wire _w924_ ;
	wire _w925_ ;
	wire _w926_ ;
	wire _w927_ ;
	wire _w928_ ;
	wire _w929_ ;
	wire _w930_ ;
	wire _w931_ ;
	wire _w932_ ;
	wire _w933_ ;
	wire _w934_ ;
	wire _w935_ ;
	wire _w936_ ;
	wire _w937_ ;
	wire _w938_ ;
	wire _w939_ ;
	wire _w940_ ;
	wire _w941_ ;
	wire _w942_ ;
	wire _w943_ ;
	wire _w944_ ;
	wire _w945_ ;
	wire _w946_ ;
	wire _w947_ ;
	wire _w948_ ;
	wire _w949_ ;
	wire _w950_ ;
	wire _w951_ ;
	wire _w952_ ;
	wire _w953_ ;
	wire _w954_ ;
	wire _w955_ ;
	wire _w956_ ;
	wire _w957_ ;
	wire _w958_ ;
	wire _w959_ ;
	wire _w960_ ;
	wire _w961_ ;
	wire _w962_ ;
	wire _w963_ ;
	wire _w964_ ;
	wire _w965_ ;
	wire _w966_ ;
	wire _w967_ ;
	wire _w968_ ;
	wire _w969_ ;
	wire _w970_ ;
	wire _w971_ ;
	wire _w972_ ;
	wire _w973_ ;
	wire _w974_ ;
	wire _w975_ ;
	wire _w976_ ;
	wire _w977_ ;
	wire _w978_ ;
	wire _w979_ ;
	wire _w980_ ;
	wire _w981_ ;
	wire _w982_ ;
	wire _w983_ ;
	wire _w984_ ;
	wire _w985_ ;
	wire _w986_ ;
	wire _w987_ ;
	wire _w988_ ;
	wire _w989_ ;
	wire _w990_ ;
	wire _w991_ ;
	wire _w992_ ;
	wire _w993_ ;
	wire _w994_ ;
	wire _w995_ ;
	wire _w996_ ;
	wire _w997_ ;
	wire _w998_ ;
	wire _w999_ ;
	wire _w1000_ ;
	wire _w1001_ ;
	wire _w1002_ ;
	wire _w1571_ ;
	wire _w1572_ ;
	wire _w1573_ ;
	wire _w1574_ ;
	wire _w1575_ ;
	wire _w1576_ ;
	wire _w1577_ ;
	wire _w1578_ ;
	wire _w1579_ ;
	wire _w1580_ ;
	wire _w1581_ ;
	wire _w1582_ ;
	wire _w1583_ ;
	wire _w1584_ ;
	wire _w1585_ ;
	wire _w1586_ ;
	wire _w1587_ ;
	wire _w1588_ ;
	wire _w1589_ ;
	wire _w1590_ ;
	wire _w1591_ ;
	wire _w1592_ ;
	wire _w1593_ ;
	wire _w1594_ ;
	wire _w1595_ ;
	wire _w1596_ ;
	wire _w1597_ ;
	wire _w1598_ ;
	wire _w1599_ ;
	wire _w1600_ ;
	wire _w1601_ ;
	wire _w1602_ ;
	wire _w1603_ ;
	wire _w1604_ ;
	wire _w1605_ ;
	wire _w1606_ ;
	wire _w1607_ ;
	wire _w1608_ ;
	wire _w1609_ ;
	wire _w1610_ ;
	wire _w1611_ ;
	wire _w1612_ ;
	wire _w1613_ ;
	wire _w1614_ ;
	wire _w1615_ ;
	wire _w1616_ ;
	wire _w1617_ ;
	wire _w1618_ ;
	wire _w1619_ ;
	wire _w1620_ ;
	wire _w1621_ ;
	wire _w1622_ ;
	wire _w1623_ ;
	wire _w1624_ ;
	wire _w1625_ ;
	wire _w1626_ ;
	wire _w1627_ ;
	wire _w1628_ ;
	wire _w1629_ ;
	wire _w1630_ ;
	wire _w1631_ ;
	wire _w1632_ ;
	wire _w1633_ ;
	wire _w1634_ ;
	wire _w1635_ ;
	wire _w1636_ ;
	wire _w1637_ ;
	wire _w1638_ ;
	wire _w1639_ ;
	wire _w1640_ ;
	wire _w1641_ ;
	wire _w1642_ ;
	wire _w1643_ ;
	wire _w1644_ ;
	wire _w1645_ ;
	wire _w1646_ ;
	wire _w1647_ ;
	wire _w1648_ ;
	wire _w1649_ ;
	wire _w1650_ ;
	wire _w1651_ ;
	wire _w1652_ ;
	wire _w1653_ ;
	wire _w1654_ ;
	wire _w1655_ ;
	wire _w1656_ ;
	wire _w1657_ ;
	wire _w1658_ ;
	wire _w1659_ ;
	wire _w1660_ ;
	wire _w1661_ ;
	wire _w1662_ ;
	wire _w1663_ ;
	wire _w1664_ ;
	wire _w1665_ ;
	wire _w1666_ ;
	wire _w1667_ ;
	wire _w1668_ ;
	wire _w1669_ ;
	wire _w1670_ ;
	wire _w1671_ ;
	wire _w1672_ ;
	wire _w1673_ ;
	wire _w1674_ ;
	wire _w1675_ ;
	wire _w1676_ ;
	wire _w1677_ ;
	wire _w1678_ ;
	wire _w1679_ ;
	wire _w1680_ ;
	wire _w1681_ ;
	wire _w1682_ ;
	wire _w1683_ ;
	wire _w1684_ ;
	wire _w1685_ ;
	wire _w1686_ ;
	wire _w1687_ ;
	wire _w1688_ ;
	wire _w1689_ ;
	wire _w1690_ ;
	wire _w1691_ ;
	wire _w1692_ ;
	wire _w1693_ ;
	wire _w1694_ ;
	wire _w1695_ ;
	wire _w1696_ ;
	wire _w1697_ ;
	wire _w1698_ ;
	wire _w1699_ ;
	wire _w1700_ ;
	wire _w1701_ ;
	wire _w1702_ ;
	wire _w1703_ ;
	wire _w1704_ ;
	wire _w1705_ ;
	wire _w1706_ ;
	wire _w1707_ ;
	wire _w1708_ ;
	wire _w1709_ ;
	wire _w1710_ ;
	wire _w1711_ ;
	wire _w1712_ ;
	wire _w1713_ ;
	wire _w1714_ ;
	wire _w1715_ ;
	wire _w1716_ ;
	wire _w1717_ ;
	wire _w1718_ ;
	wire _w1719_ ;
	wire _w1720_ ;
	wire _w1721_ ;
	wire _w1722_ ;
	wire _w1723_ ;
	wire _w1724_ ;
	wire _w1725_ ;
	wire _w1726_ ;
	wire _w1727_ ;
	wire _w1728_ ;
	wire _w1729_ ;
	wire _w1730_ ;
	wire _w1731_ ;
	wire _w1732_ ;
	wire _w1733_ ;
	wire _w1734_ ;
	wire _w1735_ ;
	wire _w1736_ ;
	wire _w1737_ ;
	wire _w1738_ ;
	wire _w1739_ ;
	wire _w1740_ ;
	wire _w1741_ ;
	wire _w1742_ ;
	wire _w1743_ ;
	wire _w1744_ ;
	wire _w1745_ ;
	wire _w1746_ ;
	wire _w1747_ ;
	wire _w1748_ ;
	wire _w1749_ ;
	wire _w1750_ ;
	wire _w1751_ ;
	wire _w1752_ ;
	wire _w1753_ ;
	wire _w1754_ ;
	wire _w1755_ ;
	wire _w1756_ ;
	wire _w1757_ ;
	wire _w1758_ ;
	wire _w1759_ ;
	wire _w1760_ ;
	wire _w1761_ ;
	wire _w1762_ ;
	wire _w1763_ ;
	wire _w1764_ ;
	wire _w1765_ ;
	wire _w1766_ ;
	wire _w1767_ ;
	wire _w1768_ ;
	wire _w1769_ ;
	wire _w1770_ ;
	wire _w1771_ ;
	wire _w1772_ ;
	wire _w1773_ ;
	wire _w1774_ ;
	wire _w1775_ ;
	wire _w1776_ ;
	wire _w1777_ ;
	wire _w1778_ ;
	wire _w1779_ ;
	wire _w1780_ ;
	wire _w1781_ ;
	wire _w1782_ ;
	wire _w1783_ ;
	wire _w1784_ ;
	wire _w1785_ ;
	wire _w1786_ ;
	wire _w1787_ ;
	wire _w1788_ ;
	wire _w1789_ ;
	wire _w1790_ ;
	wire _w1791_ ;
	wire _w1792_ ;
	wire _w1793_ ;
	wire _w1794_ ;
	wire _w1795_ ;
	wire _w1796_ ;
	wire _w1797_ ;
	wire _w1798_ ;
	wire _w1799_ ;
	wire _w1800_ ;
	wire _w1801_ ;
	wire _w1802_ ;
	wire _w1803_ ;
	wire _w1804_ ;
	wire _w1805_ ;
	wire _w1806_ ;
	wire _w1807_ ;
	wire _w1808_ ;
	wire _w1809_ ;
	wire _w1810_ ;
	wire _w1811_ ;
	wire _w1812_ ;
	wire _w1813_ ;
	wire _w1814_ ;
	wire _w1815_ ;
	wire _w1816_ ;
	wire _w1817_ ;
	wire _w1818_ ;
	wire _w1819_ ;
	wire _w1820_ ;
	wire _w1821_ ;
	wire _w1822_ ;
	wire _w1823_ ;
	wire _w1824_ ;
	wire _w1825_ ;
	wire _w1826_ ;
	wire _w1827_ ;
	wire _w1828_ ;
	wire _w1829_ ;
	wire _w1830_ ;
	wire _w1831_ ;
	wire _w1832_ ;
	wire _w1833_ ;
	wire _w1834_ ;
	wire _w1835_ ;
	wire _w1836_ ;
	wire _w1837_ ;
	wire _w1838_ ;
	wire _w1839_ ;
	wire _w1840_ ;
	wire _w1841_ ;
	wire _w1842_ ;
	wire _w1843_ ;
	wire _w1844_ ;
	wire _w1845_ ;
	wire _w1846_ ;
	wire _w1847_ ;
	wire _w1848_ ;
	wire _w1849_ ;
	wire _w1850_ ;
	wire _w1851_ ;
	wire _w1852_ ;
	wire _w1853_ ;
	wire _w1854_ ;
	wire _w1855_ ;
	wire _w1856_ ;
	wire _w1857_ ;
	wire _w1858_ ;
	wire _w1859_ ;
	wire _w1860_ ;
	wire _w1861_ ;
	wire _w1862_ ;
	wire _w1863_ ;
	wire _w1864_ ;
	wire _w1865_ ;
	wire _w1866_ ;
	wire _w1867_ ;
	wire _w1868_ ;
	wire _w1869_ ;
	wire _w1870_ ;
	wire _w1871_ ;
	wire _w1872_ ;
	wire _w1873_ ;
	wire _w1874_ ;
	wire _w1875_ ;
	wire _w1876_ ;
	wire _w1877_ ;
	wire _w1878_ ;
	wire _w1879_ ;
	wire _w1880_ ;
	wire _w1881_ ;
	wire _w1882_ ;
	wire _w1883_ ;
	wire _w1884_ ;
	wire _w1885_ ;
	wire _w1886_ ;
	wire _w1887_ ;
	wire _w1888_ ;
	wire _w1889_ ;
	wire _w1890_ ;
	wire _w1891_ ;
	wire _w1892_ ;
	wire _w1893_ ;
	wire _w1894_ ;
	wire _w1895_ ;
	wire _w1896_ ;
	wire _w1897_ ;
	wire _w1898_ ;
	wire _w1899_ ;
	wire _w1900_ ;
	wire _w1901_ ;
	wire _w1902_ ;
	wire _w1903_ ;
	wire _w1904_ ;
	wire _w1905_ ;
	wire _w1906_ ;
	wire _w1907_ ;
	wire _w1908_ ;
	wire _w1909_ ;
	wire _w1910_ ;
	wire _w1911_ ;
	wire _w1912_ ;
	wire _w1913_ ;
	wire _w1914_ ;
	wire _w1915_ ;
	wire _w1916_ ;
	wire _w1917_ ;
	wire _w1918_ ;
	wire _w1919_ ;
	wire _w1920_ ;
	wire _w1921_ ;
	wire _w1922_ ;
	wire _w1923_ ;
	wire _w1924_ ;
	wire _w1925_ ;
	wire _w1926_ ;
	wire _w1927_ ;
	wire _w1928_ ;
	wire _w1929_ ;
	wire _w1930_ ;
	wire _w1931_ ;
	wire _w1932_ ;
	wire _w1933_ ;
	wire _w1934_ ;
	wire _w1935_ ;
	wire _w1936_ ;
	wire _w1937_ ;
	wire _w1938_ ;
	wire _w1939_ ;
	wire _w1940_ ;
	wire _w1941_ ;
	wire _w1942_ ;
	wire _w1943_ ;
	wire _w1944_ ;
	wire _w1945_ ;
	wire _w1946_ ;
	wire _w1947_ ;
	wire _w1948_ ;
	wire _w1949_ ;
	wire _w1950_ ;
	wire _w1951_ ;
	wire _w1952_ ;
	wire _w1953_ ;
	wire _w1954_ ;
	wire _w1955_ ;
	wire _w1956_ ;
	wire _w1957_ ;
	wire _w1958_ ;
	wire _w1959_ ;
	wire _w1960_ ;
	wire _w1961_ ;
	wire _w1962_ ;
	wire _w1963_ ;
	wire _w1964_ ;
	wire _w1965_ ;
	wire _w1966_ ;
	wire _w1967_ ;
	wire _w1968_ ;
	wire _w1969_ ;
	wire _w1970_ ;
	wire _w1971_ ;
	wire _w1972_ ;
	wire _w1973_ ;
	wire _w1974_ ;
	wire _w1975_ ;
	wire _w1976_ ;
	wire _w1977_ ;
	wire _w1978_ ;
	wire _w1979_ ;
	wire _w1980_ ;
	wire _w1981_ ;
	wire _w1982_ ;
	wire _w1983_ ;
	wire _w1984_ ;
	wire _w1985_ ;
	wire _w1986_ ;
	wire _w1987_ ;
	wire _w1988_ ;
	wire _w1989_ ;
	wire _w1990_ ;
	wire _w1991_ ;
	wire _w1992_ ;
	wire _w1993_ ;
	wire _w1994_ ;
	wire _w1995_ ;
	wire _w1996_ ;
	wire _w1997_ ;
	wire _w1998_ ;
	wire _w1999_ ;
	wire _w2000_ ;
	wire _w2001_ ;
	wire _w2002_ ;
	wire _w2003_ ;
	wire _w2004_ ;
	wire _w2005_ ;
	wire _w2006_ ;
	wire _w2007_ ;
	wire _w2008_ ;
	wire _w2009_ ;
	wire _w2010_ ;
	wire _w2011_ ;
	wire _w2012_ ;
	wire _w2013_ ;
	wire _w2014_ ;
	wire _w2015_ ;
	wire _w2016_ ;
	wire _w2017_ ;
	wire _w2018_ ;
	wire _w2019_ ;
	wire _w2020_ ;
	wire _w2021_ ;
	wire _w2022_ ;
	wire _w2023_ ;
	wire _w2024_ ;
	wire _w2025_ ;
	wire _w2026_ ;
	wire _w2027_ ;
	wire _w2028_ ;
	wire _w2029_ ;
	wire _w2030_ ;
	wire _w2031_ ;
	wire _w2032_ ;
	wire _w2033_ ;
	wire _w2034_ ;
	wire _w2035_ ;
	wire _w2036_ ;
	wire _w2037_ ;
	wire _w2038_ ;
	wire _w2039_ ;
	wire _w2040_ ;
	wire _w2041_ ;
	wire _w2042_ ;
	wire _w2043_ ;
	wire _w2044_ ;
	wire _w2045_ ;
	wire _w2046_ ;
	wire _w2047_ ;
	wire _w2048_ ;
	wire _w2049_ ;
	wire _w2050_ ;
	wire _w2051_ ;
	wire _w2052_ ;
	wire _w2053_ ;
	wire _w2054_ ;
	wire _w2055_ ;
	wire _w2056_ ;
	wire _w2057_ ;
	wire _w2058_ ;
	wire _w2059_ ;
	wire _w2060_ ;
	wire _w2061_ ;
	wire _w2062_ ;
	wire _w2063_ ;
	wire _w2064_ ;
	wire _w2065_ ;
	wire _w2066_ ;
	wire _w2067_ ;
	wire _w2068_ ;
	wire _w2069_ ;
	wire _w2070_ ;
	wire _w2071_ ;
	wire _w2072_ ;
	wire _w2073_ ;
	wire _w2074_ ;
	wire _w2075_ ;
	wire _w2076_ ;
	wire _w2077_ ;
	wire _w2078_ ;
	wire _w2079_ ;
	wire _w2080_ ;
	wire _w2081_ ;
	wire _w2082_ ;
	wire _w2083_ ;
	wire _w2084_ ;
	wire _w2085_ ;
	wire _w2086_ ;
	wire _w2087_ ;
	wire _w2088_ ;
	wire _w2089_ ;
	wire _w2090_ ;
	wire _w2091_ ;
	wire _w2092_ ;
	wire _w2093_ ;
	wire _w2094_ ;
	wire _w2095_ ;
	wire _w2096_ ;
	wire _w2097_ ;
	wire _w2098_ ;
	wire _w2099_ ;
	wire _w2100_ ;
	wire _w2101_ ;
	wire _w2102_ ;
	wire _w2103_ ;
	wire _w2104_ ;
	wire _w2105_ ;
	wire _w2106_ ;
	wire _w2107_ ;
	wire _w2108_ ;
	wire _w2109_ ;
	wire _w2110_ ;
	wire _w2111_ ;
	wire _w2112_ ;
	wire _w2113_ ;
	wire _w2114_ ;
	wire _w2115_ ;
	wire _w2116_ ;
	wire _w2117_ ;
	wire _w2118_ ;
	wire _w2119_ ;
	wire _w2120_ ;
	wire _w2121_ ;
	wire _w2122_ ;
	wire _w2123_ ;
	wire _w2124_ ;
	wire _w2125_ ;
	wire _w2126_ ;
	wire _w2127_ ;
	wire _w2128_ ;
	wire _w2129_ ;
	wire _w2130_ ;
	wire _w2131_ ;
	wire _w2132_ ;
	wire _w2133_ ;
	wire _w2134_ ;
	wire _w2135_ ;
	wire _w2136_ ;
	wire _w2137_ ;
	wire _w2138_ ;
	wire _w2139_ ;
	wire _w2140_ ;
	wire _w2141_ ;
	wire _w2142_ ;
	wire _w2143_ ;
	wire _w2144_ ;
	wire _w2145_ ;
	wire _w2146_ ;
	wire _w2147_ ;
	wire _w2148_ ;
	wire _w2149_ ;
	wire _w2150_ ;
	wire _w2151_ ;
	wire _w2152_ ;
	wire _w2153_ ;
	wire _w2154_ ;
	wire _w2155_ ;
	wire _w2156_ ;
	wire _w2157_ ;
	wire _w2158_ ;
	wire _w2159_ ;
	wire _w2160_ ;
	wire _w2161_ ;
	wire _w2162_ ;
	wire _w2163_ ;
	wire _w2164_ ;
	wire _w2165_ ;
	wire _w2166_ ;
	wire _w2167_ ;
	wire _w2168_ ;
	wire _w2169_ ;
	wire _w2170_ ;
	wire _w2171_ ;
	wire _w2172_ ;
	wire _w2173_ ;
	wire _w2174_ ;
	wire _w2175_ ;
	wire _w2176_ ;
	wire _w2177_ ;
	wire _w2178_ ;
	wire _w2179_ ;
	wire _w2180_ ;
	wire _w2181_ ;
	wire _w2182_ ;
	wire _w2183_ ;
	wire _w2184_ ;
	wire _w2185_ ;
	wire _w2186_ ;
	wire _w2187_ ;
	wire _w2188_ ;
	wire _w2189_ ;
	wire _w2190_ ;
	wire _w2191_ ;
	wire _w2192_ ;
	wire _w2193_ ;
	wire _w2194_ ;
	wire _w2195_ ;
	wire _w2196_ ;
	wire _w2197_ ;
	wire _w2198_ ;
	wire _w2199_ ;
	wire _w2200_ ;
	wire _w2201_ ;
	wire _w2202_ ;
	wire _w2203_ ;
	wire _w2204_ ;
	wire _w2205_ ;
	wire _w2206_ ;
	wire _w2207_ ;
	wire _w2208_ ;
	wire _w2209_ ;
	wire _w2210_ ;
	wire _w2211_ ;
	wire _w2212_ ;
	wire _w2213_ ;
	wire _w2214_ ;
	wire _w2215_ ;
	wire _w2216_ ;
	wire _w2217_ ;
	wire _w2218_ ;
	wire _w2219_ ;
	wire _w2220_ ;
	wire _w2221_ ;
	wire _w2222_ ;
	wire _w2223_ ;
	wire _w2224_ ;
	wire _w2225_ ;
	wire _w2226_ ;
	wire _w2227_ ;
	wire _w2228_ ;
	wire _w2229_ ;
	wire _w2230_ ;
	wire _w2231_ ;
	wire _w2232_ ;
	wire _w2233_ ;
	wire _w2234_ ;
	wire _w2235_ ;
	wire _w2236_ ;
	wire _w2237_ ;
	wire _w2238_ ;
	wire _w2239_ ;
	wire _w2240_ ;
	wire _w2241_ ;
	wire _w2242_ ;
	wire _w2243_ ;
	wire _w2244_ ;
	wire _w2245_ ;
	wire _w2246_ ;
	wire _w2247_ ;
	wire _w2248_ ;
	wire _w2249_ ;
	wire _w2250_ ;
	wire _w2251_ ;
	wire _w2252_ ;
	wire _w2253_ ;
	wire _w2254_ ;
	wire _w2255_ ;
	wire _w2256_ ;
	wire _w2257_ ;
	wire _w2258_ ;
	wire _w2259_ ;
	wire _w2260_ ;
	wire _w2261_ ;
	wire _w2262_ ;
	wire _w2263_ ;
	wire _w2264_ ;
	wire _w2265_ ;
	wire _w2266_ ;
	wire _w2267_ ;
	wire _w2268_ ;
	wire _w2269_ ;
	wire _w2270_ ;
	wire _w2271_ ;
	wire _w2272_ ;
	wire _w2273_ ;
	wire _w2274_ ;
	wire _w2275_ ;
	wire _w2276_ ;
	wire _w2277_ ;
	wire _w2278_ ;
	wire _w2279_ ;
	wire _w2280_ ;
	wire _w2281_ ;
	wire _w2282_ ;
	wire _w2283_ ;
	wire _w2284_ ;
	wire _w2285_ ;
	wire _w2286_ ;
	wire _w2287_ ;
	wire _w2288_ ;
	wire _w2289_ ;
	wire _w2290_ ;
	wire _w2291_ ;
	wire _w2292_ ;
	wire _w2293_ ;
	wire _w2294_ ;
	wire _w2295_ ;
	wire _w2296_ ;
	wire _w2297_ ;
	wire _w2298_ ;
	wire _w2299_ ;
	wire _w2300_ ;
	wire _w2301_ ;
	wire _w2302_ ;
	wire _w2303_ ;
	wire _w2304_ ;
	wire _w2305_ ;
	wire _w2306_ ;
	wire _w2307_ ;
	wire _w2308_ ;
	wire _w2309_ ;
	wire _w2310_ ;
	wire _w2311_ ;
	wire _w2312_ ;
	wire _w2313_ ;
	wire _w2314_ ;
	wire _w2315_ ;
	wire _w2316_ ;
	wire _w2317_ ;
	wire _w2318_ ;
	wire _w2319_ ;
	wire _w2320_ ;
	wire _w2321_ ;
	wire _w2322_ ;
	wire _w2323_ ;
	wire _w2324_ ;
	wire _w2325_ ;
	wire _w2326_ ;
	wire _w2327_ ;
	wire _w2328_ ;
	wire _w2329_ ;
	wire _w2330_ ;
	wire _w2331_ ;
	wire _w2332_ ;
	wire _w2333_ ;
	wire _w2334_ ;
	wire _w2335_ ;
	wire _w2336_ ;
	wire _w2337_ ;
	wire _w2338_ ;
	wire _w2339_ ;
	wire _w2340_ ;
	wire _w2341_ ;
	wire _w2342_ ;
	wire _w2343_ ;
	wire _w2344_ ;
	wire _w2345_ ;
	wire _w2346_ ;
	wire _w2347_ ;
	wire _w2348_ ;
	wire _w2349_ ;
	wire _w2350_ ;
	wire _w2351_ ;
	wire _w2352_ ;
	wire _w2353_ ;
	wire _w2354_ ;
	wire _w2355_ ;
	wire _w2356_ ;
	wire _w2357_ ;
	wire _w2358_ ;
	wire _w2359_ ;
	wire _w2360_ ;
	wire _w2361_ ;
	wire _w2362_ ;
	wire _w2363_ ;
	wire _w2364_ ;
	wire _w2365_ ;
	wire _w2366_ ;
	wire _w2367_ ;
	wire _w2368_ ;
	wire _w2369_ ;
	wire _w2370_ ;
	wire _w2371_ ;
	wire _w2372_ ;
	wire _w2373_ ;
	wire _w2374_ ;
	wire _w2375_ ;
	wire _w2376_ ;
	wire _w2377_ ;
	wire _w2378_ ;
	wire _w2379_ ;
	wire _w2380_ ;
	wire _w2381_ ;
	wire _w2382_ ;
	wire _w2383_ ;
	wire _w2384_ ;
	wire _w2385_ ;
	wire _w2386_ ;
	wire _w2387_ ;
	wire _w2388_ ;
	wire _w2389_ ;
	wire _w2390_ ;
	wire _w2391_ ;
	wire _w2392_ ;
	wire _w2393_ ;
	wire _w2394_ ;
	wire _w2395_ ;
	wire _w2396_ ;
	wire _w2397_ ;
	wire _w2398_ ;
	wire _w2399_ ;
	wire _w2400_ ;
	wire _w2401_ ;
	wire _w2402_ ;
	wire _w2403_ ;
	wire _w2404_ ;
	wire _w2405_ ;
	wire _w2406_ ;
	wire _w2407_ ;
	wire _w2408_ ;
	wire _w2409_ ;
	wire _w2410_ ;
	wire _w2411_ ;
	wire _w2412_ ;
	wire _w2413_ ;
	wire _w2414_ ;
	wire _w2415_ ;
	wire _w2416_ ;
	wire _w2417_ ;
	wire _w2418_ ;
	wire _w2419_ ;
	wire _w2420_ ;
	wire _w2421_ ;
	wire _w2422_ ;
	wire _w2423_ ;
	wire _w2424_ ;
	wire _w2425_ ;
	wire _w2426_ ;
	wire _w2427_ ;
	wire _w2428_ ;
	wire _w2429_ ;
	wire _w2430_ ;
	wire _w2431_ ;
	wire _w2432_ ;
	wire _w2433_ ;
	wire _w2434_ ;
	wire _w2435_ ;
	wire _w2436_ ;
	wire _w2437_ ;
	wire _w2438_ ;
	wire _w2439_ ;
	wire _w2440_ ;
	wire _w2441_ ;
	wire _w2442_ ;
	wire _w2443_ ;
	wire _w2444_ ;
	wire _w2445_ ;
	wire _w2446_ ;
	wire _w2447_ ;
	wire _w2448_ ;
	wire _w2449_ ;
	wire _w2450_ ;
	wire _w2451_ ;
	wire _w2452_ ;
	wire _w2453_ ;
	wire _w2454_ ;
	wire _w2455_ ;
	wire _w2456_ ;
	wire _w2457_ ;
	wire _w2458_ ;
	wire _w2459_ ;
	wire _w2460_ ;
	wire _w2461_ ;
	wire _w2462_ ;
	wire _w2463_ ;
	wire _w2464_ ;
	wire _w2465_ ;
	wire _w2466_ ;
	wire _w2467_ ;
	wire _w2468_ ;
	wire _w2469_ ;
	wire _w2470_ ;
	wire _w2471_ ;
	wire _w2472_ ;
	wire _w2473_ ;
	wire _w2474_ ;
	wire _w2475_ ;
	wire _w2476_ ;
	wire _w2477_ ;
	wire _w2478_ ;
	wire _w2479_ ;
	wire _w2480_ ;
	wire _w2481_ ;
	wire _w2482_ ;
	wire _w2483_ ;
	wire _w2484_ ;
	wire _w2485_ ;
	wire _w2486_ ;
	wire _w2487_ ;
	wire _w2488_ ;
	wire _w2489_ ;
	wire _w2490_ ;
	wire _w2491_ ;
	wire _w2492_ ;
	wire _w2493_ ;
	wire _w2494_ ;
	wire _w2495_ ;
	wire _w2496_ ;
	wire _w2497_ ;
	wire _w2498_ ;
	wire _w2499_ ;
	wire _w2500_ ;
	wire _w2501_ ;
	wire _w2502_ ;
	wire _w2503_ ;
	wire _w2504_ ;
	wire _w2505_ ;
	wire _w2506_ ;
	wire _w2507_ ;
	wire _w2508_ ;
	wire _w2509_ ;
	wire _w2510_ ;
	wire _w2511_ ;
	wire _w2512_ ;
	wire _w2513_ ;
	wire _w2514_ ;
	wire _w2515_ ;
	wire _w2516_ ;
	wire _w2517_ ;
	wire _w2518_ ;
	wire _w2519_ ;
	wire _w2520_ ;
	wire _w2521_ ;
	wire _w2522_ ;
	wire _w2523_ ;
	wire _w2524_ ;
	wire _w2525_ ;
	wire _w2526_ ;
	wire _w2527_ ;
	wire _w2528_ ;
	wire _w2529_ ;
	wire _w2530_ ;
	wire _w2531_ ;
	wire _w2532_ ;
	wire _w2533_ ;
	wire _w2534_ ;
	wire _w2535_ ;
	wire _w2536_ ;
	wire _w2537_ ;
	wire _w2538_ ;
	wire _w2539_ ;
	wire _w2540_ ;
	wire _w2541_ ;
	wire _w2542_ ;
	wire _w2543_ ;
	wire _w2544_ ;
	wire _w2545_ ;
	wire _w2546_ ;
	wire _w2547_ ;
	wire _w2548_ ;
	wire _w2549_ ;
	wire _w2550_ ;
	wire _w2551_ ;
	wire _w2552_ ;
	wire _w2553_ ;
	wire _w2554_ ;
	wire _w2555_ ;
	wire _w2556_ ;
	wire _w2557_ ;
	wire _w2558_ ;
	wire _w2559_ ;
	wire _w2560_ ;
	wire _w2561_ ;
	wire _w2562_ ;
	wire _w2563_ ;
	wire _w2564_ ;
	wire _w2565_ ;
	wire _w2566_ ;
	wire _w2567_ ;
	wire _w2568_ ;
	wire _w2569_ ;
	wire _w2570_ ;
	wire _w2571_ ;
	wire _w2572_ ;
	wire _w2573_ ;
	wire _w2574_ ;
	wire _w2575_ ;
	wire _w2576_ ;
	wire _w2577_ ;
	wire _w2578_ ;
	wire _w2579_ ;
	wire _w2580_ ;
	wire _w2581_ ;
	wire _w2582_ ;
	wire _w2583_ ;
	wire _w2584_ ;
	wire _w2585_ ;
	wire _w2586_ ;
	wire _w2587_ ;
	wire _w2588_ ;
	wire _w2589_ ;
	wire _w2590_ ;
	wire _w2591_ ;
	wire _w2592_ ;
	wire _w2593_ ;
	wire _w2594_ ;
	wire _w2595_ ;
	wire _w2596_ ;
	wire _w2597_ ;
	wire _w2598_ ;
	wire _w2599_ ;
	wire _w2600_ ;
	wire _w2601_ ;
	wire _w2602_ ;
	wire _w2603_ ;
	wire _w2604_ ;
	wire _w2605_ ;
	wire _w2606_ ;
	wire _w2607_ ;
	wire _w2608_ ;
	wire _w2609_ ;
	wire _w2610_ ;
	wire _w2611_ ;
	wire _w2612_ ;
	wire _w2613_ ;
	wire _w2614_ ;
	wire _w2615_ ;
	wire _w2616_ ;
	wire _w2617_ ;
	wire _w2618_ ;
	wire _w2619_ ;
	wire _w2620_ ;
	wire _w2621_ ;
	wire _w2622_ ;
	wire _w2623_ ;
	wire _w2624_ ;
	wire _w2625_ ;
	wire _w2626_ ;
	wire _w2627_ ;
	wire _w2628_ ;
	wire _w2629_ ;
	wire _w2630_ ;
	wire _w2631_ ;
	wire _w2632_ ;
	wire _w2633_ ;
	wire _w2634_ ;
	wire _w2635_ ;
	wire _w2636_ ;
	wire _w2637_ ;
	wire _w2638_ ;
	wire _w2639_ ;
	wire _w2640_ ;
	wire _w2641_ ;
	wire _w2642_ ;
	wire _w2643_ ;
	wire _w2644_ ;
	wire _w2645_ ;
	wire _w2646_ ;
	wire _w2647_ ;
	wire _w2648_ ;
	wire _w2649_ ;
	wire _w2650_ ;
	wire _w2651_ ;
	wire _w2652_ ;
	wire _w2653_ ;
	wire _w2654_ ;
	wire _w2655_ ;
	wire _w2656_ ;
	wire _w2657_ ;
	wire _w2658_ ;
	wire _w2659_ ;
	wire _w2660_ ;
	wire _w2661_ ;
	wire _w2662_ ;
	wire _w2663_ ;
	wire _w2664_ ;
	wire _w2665_ ;
	wire _w2666_ ;
	wire _w2667_ ;
	wire _w2668_ ;
	wire _w2669_ ;
	wire _w2670_ ;
	wire _w2671_ ;
	wire _w2672_ ;
	wire _w2673_ ;
	wire _w2674_ ;
	wire _w2675_ ;
	wire _w2676_ ;
	wire _w2677_ ;
	wire _w2678_ ;
	wire _w2679_ ;
	wire _w2680_ ;
	wire _w2681_ ;
	wire _w2682_ ;
	wire _w2683_ ;
	wire _w2684_ ;
	wire _w2685_ ;
	wire _w2686_ ;
	wire _w2687_ ;
	wire _w2688_ ;
	wire _w2689_ ;
	wire _w2690_ ;
	wire _w2691_ ;
	wire _w2692_ ;
	wire _w2693_ ;
	wire _w2694_ ;
	wire _w2695_ ;
	wire _w2696_ ;
	wire _w2697_ ;
	wire _w2698_ ;
	wire _w2699_ ;
	wire _w2700_ ;
	wire _w2701_ ;
	wire _w2702_ ;
	wire _w2703_ ;
	wire _w2704_ ;
	wire _w2705_ ;
	wire _w2706_ ;
	wire _w2707_ ;
	wire _w2708_ ;
	wire _w2709_ ;
	wire _w2710_ ;
	wire _w2711_ ;
	wire _w2712_ ;
	wire _w2713_ ;
	wire _w2714_ ;
	wire _w2715_ ;
	wire _w2716_ ;
	wire _w2717_ ;
	wire _w2718_ ;
	wire _w2719_ ;
	wire _w2720_ ;
	wire _w2721_ ;
	wire _w2722_ ;
	wire _w2723_ ;
	wire _w2724_ ;
	wire _w2725_ ;
	wire _w2726_ ;
	wire _w2727_ ;
	wire _w2728_ ;
	wire _w2729_ ;
	wire _w2730_ ;
	wire _w2731_ ;
	wire _w2732_ ;
	wire _w2733_ ;
	wire _w2734_ ;
	wire _w2735_ ;
	wire _w2736_ ;
	wire _w2737_ ;
	wire _w2738_ ;
	wire _w2739_ ;
	wire _w2740_ ;
	wire _w2741_ ;
	wire _w2742_ ;
	wire _w2743_ ;
	wire _w2744_ ;
	wire _w2745_ ;
	wire _w2746_ ;
	wire _w2747_ ;
	wire _w2748_ ;
	wire _w2749_ ;
	wire _w2750_ ;
	wire _w2751_ ;
	wire _w2752_ ;
	wire _w2753_ ;
	wire _w2754_ ;
	wire _w2755_ ;
	wire _w2756_ ;
	wire _w2757_ ;
	wire _w2758_ ;
	wire _w2759_ ;
	wire _w2760_ ;
	wire _w2761_ ;
	wire _w2762_ ;
	wire _w2763_ ;
	wire _w2764_ ;
	wire _w2765_ ;
	wire _w2766_ ;
	wire _w2767_ ;
	wire _w2768_ ;
	wire _w2769_ ;
	wire _w2770_ ;
	wire _w2771_ ;
	wire _w2772_ ;
	wire _w2773_ ;
	wire _w2774_ ;
	wire _w2775_ ;
	wire _w2776_ ;
	wire _w2777_ ;
	wire _w2778_ ;
	wire _w2779_ ;
	wire _w2780_ ;
	wire _w2781_ ;
	wire _w2782_ ;
	wire _w2783_ ;
	wire _w2784_ ;
	wire _w2785_ ;
	wire _w2786_ ;
	wire _w2787_ ;
	wire _w2788_ ;
	wire _w2789_ ;
	wire _w2790_ ;
	wire _w2791_ ;
	wire _w2792_ ;
	wire _w2793_ ;
	wire _w2794_ ;
	wire _w2795_ ;
	wire _w2796_ ;
	wire _w2797_ ;
	wire _w2798_ ;
	wire _w2799_ ;
	wire _w2800_ ;
	wire _w2801_ ;
	wire _w2802_ ;
	wire _w2803_ ;
	wire _w2804_ ;
	wire _w2805_ ;
	wire _w2806_ ;
	wire _w2807_ ;
	wire _w2808_ ;
	wire _w2809_ ;
	wire _w2810_ ;
	wire _w2811_ ;
	wire _w2812_ ;
	wire _w2813_ ;
	wire _w2814_ ;
	wire _w2815_ ;
	wire _w2816_ ;
	wire _w2817_ ;
	wire _w2818_ ;
	wire _w5549_ ;
	wire _w5550_ ;
	wire _w5551_ ;
	wire _w5552_ ;
	wire _w5553_ ;
	wire _w5554_ ;
	wire _w5555_ ;
	wire _w5556_ ;
	wire _w5557_ ;
	wire _w5558_ ;
	wire _w5559_ ;
	wire _w5560_ ;
	wire _w5561_ ;
	wire _w5562_ ;
	wire _w5563_ ;
	wire _w5564_ ;
	wire _w5565_ ;
	wire _w5566_ ;
	wire _w5567_ ;
	wire _w5568_ ;
	wire _w5569_ ;
	wire _w5570_ ;
	wire _w5571_ ;
	wire _w5572_ ;
	wire _w5573_ ;
	wire _w5574_ ;
	wire _w5575_ ;
	wire _w5576_ ;
	wire _w5577_ ;
	wire _w5578_ ;
	wire _w5579_ ;
	wire _w5580_ ;
	wire _w5581_ ;
	wire _w5582_ ;
	wire _w5583_ ;
	wire _w5584_ ;
	wire _w5585_ ;
	wire _w5586_ ;
	wire _w5587_ ;
	wire _w5588_ ;
	wire _w5589_ ;
	wire _w5590_ ;
	wire _w5591_ ;
	wire _w5592_ ;
	wire _w5593_ ;
	wire _w5594_ ;
	wire _w5595_ ;
	wire _w5596_ ;
	wire _w5597_ ;
	wire _w5598_ ;
	wire _w5599_ ;
	wire _w5600_ ;
	wire _w5601_ ;
	wire _w5602_ ;
	wire _w5603_ ;
	wire _w5604_ ;
	wire _w5605_ ;
	wire _w5606_ ;
	wire _w5607_ ;
	wire _w5608_ ;
	wire _w5609_ ;
	wire _w5610_ ;
	wire _w5611_ ;
	wire _w5612_ ;
	wire _w5613_ ;
	wire _w5614_ ;
	wire _w5615_ ;
	wire _w5616_ ;
	wire _w5617_ ;
	wire _w5618_ ;
	wire _w5619_ ;
	wire _w5620_ ;
	wire _w5621_ ;
	wire _w5622_ ;
	wire _w5623_ ;
	wire _w5624_ ;
	wire _w5625_ ;
	wire _w5626_ ;
	wire _w5627_ ;
	wire _w5628_ ;
	wire _w5629_ ;
	wire _w5630_ ;
	wire _w5631_ ;
	wire _w5632_ ;
	wire _w5633_ ;
	wire _w5634_ ;
	wire _w5635_ ;
	wire _w5636_ ;
	wire _w5637_ ;
	wire _w5638_ ;
	wire _w5639_ ;
	wire _w5640_ ;
	wire _w5641_ ;
	wire _w5642_ ;
	wire _w5643_ ;
	wire _w5644_ ;
	wire _w5645_ ;
	wire _w5646_ ;
	wire _w5647_ ;
	wire _w5648_ ;
	wire _w5649_ ;
	wire _w5650_ ;
	wire _w5651_ ;
	wire _w5652_ ;
	wire _w5653_ ;
	wire _w5654_ ;
	wire _w5655_ ;
	wire _w5656_ ;
	wire _w5657_ ;
	wire _w5658_ ;
	wire _w5659_ ;
	wire _w5660_ ;
	wire _w5661_ ;
	wire _w5662_ ;
	wire _w5663_ ;
	wire _w5664_ ;
	wire _w5665_ ;
	wire _w5666_ ;
	wire _w5667_ ;
	wire _w5668_ ;
	wire _w5669_ ;
	wire _w5670_ ;
	wire _w5671_ ;
	wire _w5672_ ;
	wire _w5673_ ;
	wire _w5674_ ;
	wire _w5675_ ;
	wire _w5676_ ;
	wire _w5677_ ;
	wire _w5678_ ;
	wire _w5679_ ;
	wire _w5680_ ;
	wire _w5681_ ;
	wire _w5682_ ;
	wire _w5683_ ;
	wire _w5684_ ;
	wire _w5685_ ;
	wire _w5686_ ;
	wire _w5687_ ;
	wire _w5688_ ;
	wire _w5689_ ;
	wire _w5690_ ;
	wire _w5691_ ;
	wire _w5692_ ;
	wire _w5693_ ;
	wire _w5694_ ;
	wire _w5695_ ;
	wire _w5696_ ;
	wire _w5697_ ;
	wire _w5698_ ;
	wire _w5699_ ;
	wire _w5700_ ;
	wire _w5701_ ;
	wire _w5702_ ;
	wire _w5703_ ;
	wire _w5704_ ;
	wire _w5705_ ;
	wire _w5706_ ;
	wire _w5707_ ;
	wire _w5708_ ;
	wire _w5709_ ;
	wire _w5710_ ;
	wire _w5711_ ;
	wire _w5712_ ;
	wire _w5713_ ;
	wire _w5714_ ;
	wire _w5715_ ;
	wire _w5716_ ;
	wire _w5717_ ;
	wire _w5718_ ;
	wire _w5719_ ;
	wire _w5720_ ;
	wire _w5721_ ;
	wire _w5722_ ;
	wire _w5723_ ;
	wire _w5724_ ;
	wire _w5725_ ;
	wire _w5726_ ;
	wire _w5727_ ;
	wire _w5728_ ;
	wire _w5729_ ;
	wire _w5730_ ;
	wire _w5731_ ;
	wire _w5732_ ;
	wire _w5733_ ;
	wire _w5734_ ;
	wire _w5735_ ;
	wire _w5736_ ;
	wire _w5737_ ;
	wire _w5738_ ;
	wire _w5739_ ;
	wire _w5740_ ;
	wire _w5741_ ;
	wire _w5742_ ;
	wire _w5743_ ;
	wire _w5744_ ;
	wire _w5745_ ;
	wire _w5746_ ;
	wire _w5747_ ;
	wire _w5748_ ;
	wire _w5749_ ;
	wire _w5750_ ;
	wire _w5751_ ;
	wire _w5752_ ;
	wire _w5753_ ;
	wire _w5754_ ;
	wire _w5755_ ;
	wire _w5756_ ;
	wire _w5757_ ;
	wire _w5758_ ;
	wire _w5759_ ;
	wire _w5760_ ;
	wire _w5761_ ;
	wire _w5762_ ;
	wire _w5763_ ;
	wire _w5764_ ;
	wire _w5765_ ;
	wire _w5766_ ;
	wire _w5767_ ;
	wire _w5768_ ;
	wire _w5769_ ;
	wire _w5770_ ;
	wire _w5771_ ;
	wire _w5772_ ;
	wire _w5773_ ;
	wire _w5774_ ;
	wire _w5775_ ;
	wire _w5776_ ;
	wire _w5777_ ;
	wire _w5778_ ;
	wire _w5779_ ;
	wire _w5780_ ;
	wire _w5781_ ;
	wire _w5782_ ;
	wire _w5783_ ;
	wire _w5784_ ;
	wire _w5785_ ;
	wire _w5786_ ;
	wire _w5787_ ;
	wire _w5788_ ;
	wire _w5789_ ;
	wire _w5790_ ;
	wire _w5791_ ;
	wire _w5792_ ;
	wire _w5793_ ;
	wire _w5794_ ;
	wire _w5795_ ;
	wire _w5796_ ;
	wire _w5797_ ;
	wire _w5798_ ;
	wire _w5799_ ;
	wire _w5800_ ;
	wire _w5801_ ;
	wire _w5802_ ;
	wire _w5803_ ;
	wire _w5804_ ;
	wire _w5805_ ;
	wire _w5806_ ;
	wire _w5807_ ;
	wire _w5808_ ;
	wire _w5809_ ;
	wire _w5810_ ;
	wire _w5811_ ;
	wire _w5812_ ;
	wire _w5813_ ;
	wire _w5814_ ;
	wire _w5815_ ;
	wire _w5816_ ;
	wire _w5817_ ;
	wire _w5818_ ;
	wire _w5819_ ;
	wire _w5820_ ;
	wire _w5821_ ;
	wire _w5822_ ;
	wire _w5823_ ;
	wire _w5824_ ;
	wire _w5825_ ;
	wire _w5826_ ;
	wire _w5827_ ;
	wire _w5828_ ;
	wire _w5829_ ;
	wire _w5830_ ;
	wire _w5831_ ;
	wire _w5832_ ;
	wire _w5833_ ;
	wire _w5834_ ;
	wire _w5835_ ;
	wire _w5836_ ;
	wire _w5837_ ;
	wire _w5838_ ;
	wire _w5839_ ;
	wire _w5840_ ;
	wire _w5841_ ;
	wire _w5842_ ;
	wire _w5843_ ;
	wire _w5844_ ;
	wire _w5845_ ;
	wire _w5846_ ;
	wire _w5847_ ;
	wire _w5848_ ;
	wire _w5849_ ;
	wire _w5850_ ;
	wire _w5851_ ;
	wire _w5852_ ;
	wire _w5853_ ;
	wire _w5854_ ;
	wire _w5855_ ;
	wire _w5856_ ;
	wire _w5857_ ;
	wire _w5858_ ;
	wire _w5859_ ;
	wire _w5860_ ;
	wire _w5861_ ;
	wire _w5862_ ;
	wire _w5863_ ;
	wire _w5864_ ;
	wire _w5865_ ;
	wire _w5866_ ;
	wire _w5867_ ;
	wire _w5868_ ;
	wire _w5869_ ;
	wire _w5870_ ;
	wire _w5871_ ;
	wire _w5872_ ;
	wire _w5873_ ;
	wire _w5874_ ;
	wire _w5875_ ;
	wire _w5876_ ;
	wire _w5877_ ;
	wire _w5878_ ;
	wire _w5879_ ;
	wire _w5880_ ;
	wire _w5881_ ;
	wire _w5882_ ;
	wire _w5883_ ;
	wire _w5884_ ;
	wire _w5885_ ;
	wire _w5886_ ;
	wire _w5887_ ;
	wire _w5888_ ;
	wire _w5889_ ;
	wire _w5890_ ;
	wire _w5891_ ;
	wire _w5892_ ;
	wire _w5893_ ;
	wire _w5894_ ;
	wire _w5895_ ;
	wire _w5896_ ;
	wire _w5897_ ;
	wire _w5898_ ;
	wire _w5899_ ;
	wire _w5900_ ;
	wire _w5901_ ;
	wire _w5902_ ;
	wire _w5903_ ;
	wire _w5904_ ;
	wire _w5905_ ;
	wire _w5906_ ;
	wire _w5907_ ;
	wire _w5908_ ;
	wire _w5909_ ;
	wire _w5910_ ;
	wire _w5911_ ;
	wire _w5912_ ;
	wire _w5913_ ;
	wire _w5914_ ;
	wire _w5915_ ;
	wire _w5916_ ;
	wire _w5917_ ;
	wire _w5918_ ;
	wire _w5919_ ;
	wire _w5920_ ;
	wire _w5921_ ;
	wire _w5922_ ;
	wire _w5923_ ;
	wire _w5924_ ;
	wire _w5925_ ;
	wire _w5926_ ;
	wire _w5927_ ;
	wire _w5928_ ;
	wire _w5929_ ;
	wire _w5930_ ;
	wire _w5931_ ;
	wire _w5932_ ;
	wire _w5933_ ;
	wire _w5934_ ;
	wire _w5935_ ;
	wire _w5936_ ;
	wire _w5937_ ;
	wire _w5938_ ;
	wire _w5939_ ;
	wire _w5940_ ;
	wire _w5941_ ;
	wire _w5942_ ;
	wire _w5943_ ;
	wire _w5944_ ;
	wire _w5945_ ;
	wire _w5946_ ;
	wire _w5947_ ;
	wire _w5948_ ;
	wire _w5949_ ;
	wire _w5950_ ;
	wire _w5951_ ;
	wire _w5952_ ;
	wire _w5953_ ;
	wire _w5954_ ;
	wire _w5955_ ;
	wire _w5956_ ;
	wire _w5957_ ;
	wire _w5958_ ;
	wire _w5959_ ;
	wire _w5960_ ;
	wire _w5961_ ;
	wire _w5962_ ;
	wire _w5963_ ;
	wire _w5964_ ;
	wire _w5965_ ;
	wire _w5966_ ;
	wire _w5967_ ;
	wire _w5968_ ;
	wire _w5969_ ;
	wire _w5970_ ;
	wire _w5971_ ;
	wire _w5972_ ;
	wire _w5973_ ;
	wire _w5974_ ;
	wire _w5975_ ;
	wire _w5976_ ;
	wire _w5977_ ;
	wire _w5978_ ;
	wire _w5979_ ;
	wire _w5980_ ;
	wire _w5981_ ;
	wire _w5982_ ;
	wire _w5983_ ;
	wire _w5984_ ;
	wire _w5985_ ;
	wire _w5986_ ;
	wire _w5987_ ;
	wire _w5988_ ;
	wire _w5989_ ;
	wire _w5990_ ;
	wire _w5991_ ;
	wire _w5992_ ;
	wire _w5993_ ;
	wire _w5994_ ;
	wire _w5995_ ;
	wire _w5996_ ;
	wire _w5997_ ;
	wire _w5998_ ;
	wire _w5999_ ;
	wire _w6000_ ;
	wire _w6001_ ;
	wire _w6002_ ;
	wire _w6003_ ;
	wire _w6004_ ;
	wire _w6005_ ;
	wire _w6006_ ;
	wire _w6007_ ;
	wire _w6008_ ;
	wire _w6009_ ;
	wire _w6010_ ;
	wire _w6011_ ;
	wire _w6012_ ;
	wire _w6013_ ;
	wire _w6014_ ;
	wire _w6015_ ;
	wire _w6016_ ;
	wire _w6017_ ;
	wire _w6018_ ;
	wire _w6019_ ;
	wire _w6020_ ;
	wire _w6021_ ;
	wire _w6022_ ;
	wire _w6023_ ;
	wire _w6024_ ;
	wire _w6025_ ;
	wire _w6026_ ;
	wire _w6027_ ;
	wire _w6028_ ;
	wire _w6029_ ;
	wire _w6030_ ;
	wire _w6031_ ;
	wire _w6032_ ;
	wire _w6033_ ;
	wire _w6034_ ;
	wire _w6035_ ;
	wire _w6036_ ;
	wire _w6037_ ;
	wire _w6038_ ;
	wire _w6039_ ;
	wire _w6040_ ;
	wire _w6041_ ;
	wire _w6042_ ;
	wire _w6043_ ;
	wire _w6044_ ;
	wire _w6045_ ;
	wire _w6046_ ;
	wire _w6047_ ;
	wire _w6048_ ;
	wire _w6049_ ;
	wire _w6050_ ;
	wire _w6051_ ;
	wire _w6052_ ;
	wire _w6053_ ;
	wire _w6054_ ;
	wire _w6055_ ;
	wire _w6056_ ;
	wire _w6057_ ;
	wire _w6058_ ;
	wire _w6059_ ;
	wire _w6060_ ;
	wire _w6061_ ;
	wire _w6062_ ;
	wire _w6063_ ;
	wire _w6064_ ;
	wire _w6065_ ;
	wire _w6066_ ;
	wire _w6067_ ;
	wire _w6068_ ;
	wire _w6069_ ;
	wire _w6070_ ;
	wire _w6071_ ;
	wire _w6072_ ;
	wire _w6073_ ;
	wire _w6074_ ;
	wire _w6075_ ;
	wire _w6076_ ;
	wire _w6077_ ;
	wire _w6078_ ;
	wire _w6079_ ;
	wire _w6080_ ;
	wire _w6081_ ;
	wire _w6082_ ;
	wire _w6083_ ;
	wire _w6084_ ;
	wire _w6085_ ;
	wire _w6086_ ;
	wire _w6087_ ;
	wire _w6088_ ;
	wire _w6089_ ;
	wire _w6090_ ;
	wire _w6091_ ;
	wire _w6092_ ;
	wire _w6093_ ;
	wire _w6094_ ;
	wire _w6095_ ;
	wire _w6096_ ;
	wire _w6097_ ;
	wire _w6098_ ;
	wire _w6099_ ;
	wire _w6100_ ;
	wire _w6101_ ;
	wire _w6102_ ;
	wire _w6103_ ;
	wire _w6104_ ;
	wire _w6105_ ;
	wire _w6106_ ;
	wire _w6107_ ;
	wire _w6108_ ;
	wire _w6109_ ;
	wire _w6110_ ;
	wire _w6111_ ;
	wire _w6112_ ;
	wire _w6113_ ;
	wire _w6114_ ;
	wire _w6115_ ;
	wire _w6116_ ;
	wire _w6117_ ;
	wire _w6118_ ;
	wire _w6119_ ;
	wire _w6120_ ;
	wire _w6121_ ;
	wire _w6122_ ;
	wire _w6123_ ;
	wire _w6124_ ;
	wire _w6125_ ;
	wire _w6126_ ;
	wire _w6127_ ;
	wire _w6128_ ;
	wire _w6129_ ;
	wire _w6130_ ;
	wire _w6131_ ;
	wire _w6132_ ;
	wire _w6133_ ;
	wire _w6134_ ;
	wire _w6135_ ;
	wire _w6136_ ;
	wire _w6137_ ;
	wire _w6138_ ;
	wire _w6139_ ;
	wire _w6140_ ;
	wire _w6141_ ;
	wire _w6142_ ;
	wire _w6143_ ;
	wire _w6144_ ;
	wire _w6145_ ;
	wire _w6146_ ;
	wire _w6147_ ;
	wire _w6148_ ;
	wire _w6149_ ;
	wire _w6150_ ;
	wire _w6151_ ;
	wire _w6152_ ;
	wire _w6153_ ;
	wire _w6154_ ;
	wire _w6155_ ;
	wire _w6156_ ;
	wire _w6157_ ;
	wire _w6158_ ;
	wire _w6159_ ;
	wire _w6160_ ;
	wire _w6161_ ;
	wire _w6162_ ;
	wire _w6163_ ;
	wire _w6164_ ;
	wire _w6165_ ;
	wire _w6166_ ;
	wire _w6167_ ;
	wire _w6168_ ;
	wire _w6169_ ;
	wire _w6170_ ;
	wire _w6171_ ;
	wire _w6172_ ;
	wire _w6173_ ;
	wire _w6174_ ;
	wire _w6175_ ;
	wire _w6176_ ;
	wire _w6177_ ;
	wire _w6178_ ;
	wire _w6179_ ;
	wire _w6180_ ;
	wire _w6181_ ;
	wire _w6182_ ;
	wire _w6183_ ;
	wire _w6184_ ;
	wire _w6185_ ;
	wire _w6186_ ;
	wire _w6187_ ;
	wire _w6188_ ;
	wire _w6189_ ;
	wire _w6190_ ;
	wire _w6191_ ;
	wire _w6192_ ;
	wire _w6193_ ;
	wire _w6194_ ;
	wire _w6195_ ;
	wire _w6196_ ;
	wire _w6197_ ;
	wire _w6198_ ;
	wire _w6199_ ;
	wire _w6200_ ;
	wire _w6201_ ;
	wire _w6202_ ;
	wire _w6203_ ;
	wire _w6204_ ;
	wire _w6205_ ;
	wire _w6206_ ;
	wire _w6207_ ;
	wire _w6208_ ;
	wire _w6209_ ;
	wire _w6210_ ;
	wire _w6211_ ;
	wire _w6212_ ;
	wire _w6213_ ;
	wire _w6214_ ;
	wire _w6215_ ;
	wire _w6216_ ;
	wire _w6217_ ;
	wire _w6218_ ;
	wire _w6219_ ;
	wire _w6220_ ;
	wire _w6221_ ;
	wire _w6222_ ;
	wire _w6223_ ;
	wire _w6224_ ;
	wire _w6225_ ;
	wire _w6226_ ;
	wire _w6227_ ;
	wire _w6228_ ;
	wire _w6229_ ;
	wire _w6230_ ;
	wire _w6231_ ;
	wire _w6232_ ;
	wire _w6233_ ;
	wire _w6234_ ;
	wire _w6235_ ;
	wire _w6236_ ;
	wire _w6237_ ;
	wire _w6238_ ;
	wire _w6239_ ;
	wire _w6240_ ;
	wire _w6241_ ;
	wire _w6242_ ;
	wire _w6243_ ;
	wire _w6244_ ;
	wire _w6245_ ;
	wire _w6246_ ;
	wire _w6247_ ;
	wire _w6248_ ;
	wire _w6249_ ;
	wire _w6250_ ;
	wire _w6251_ ;
	wire _w6252_ ;
	wire _w6253_ ;
	wire _w6254_ ;
	wire _w6255_ ;
	wire _w6256_ ;
	wire _w6257_ ;
	wire _w6258_ ;
	wire _w6259_ ;
	wire _w6260_ ;
	wire _w6261_ ;
	wire _w6262_ ;
	wire _w6263_ ;
	wire _w6264_ ;
	wire _w6265_ ;
	wire _w6266_ ;
	wire _w6267_ ;
	wire _w6268_ ;
	wire _w6269_ ;
	wire _w6270_ ;
	wire _w6271_ ;
	wire _w6272_ ;
	wire _w6273_ ;
	wire _w6274_ ;
	wire _w6275_ ;
	wire _w6276_ ;
	wire _w6277_ ;
	wire _w6278_ ;
	wire _w6279_ ;
	wire _w6280_ ;
	wire _w6281_ ;
	wire _w6282_ ;
	wire _w6283_ ;
	wire _w6284_ ;
	wire _w6285_ ;
	wire _w6286_ ;
	wire _w6287_ ;
	wire _w6288_ ;
	wire _w6289_ ;
	wire _w6290_ ;
	wire _w6291_ ;
	wire _w6292_ ;
	wire _w6293_ ;
	wire _w6294_ ;
	wire _w6295_ ;
	wire _w6296_ ;
	wire _w6297_ ;
	wire _w6298_ ;
	wire _w6299_ ;
	wire _w6300_ ;
	wire _w6301_ ;
	wire _w6302_ ;
	wire _w6303_ ;
	wire _w6304_ ;
	wire _w6305_ ;
	wire _w6306_ ;
	wire _w6307_ ;
	wire _w6308_ ;
	wire _w6309_ ;
	wire _w6310_ ;
	wire _w6311_ ;
	wire _w6312_ ;
	wire _w6313_ ;
	wire _w6314_ ;
	wire _w6315_ ;
	wire _w6316_ ;
	wire _w6317_ ;
	wire _w6318_ ;
	wire _w6319_ ;
	wire _w6320_ ;
	wire _w6321_ ;
	wire _w6322_ ;
	wire _w6323_ ;
	wire _w6324_ ;
	wire _w6325_ ;
	wire _w6326_ ;
	wire _w6327_ ;
	wire _w6328_ ;
	wire _w6329_ ;
	wire _w6330_ ;
	wire _w6331_ ;
	wire _w6332_ ;
	wire _w6333_ ;
	wire _w6334_ ;
	wire _w6335_ ;
	wire _w6336_ ;
	wire _w6337_ ;
	wire _w6338_ ;
	wire _w6339_ ;
	wire _w6340_ ;
	wire _w6341_ ;
	wire _w6342_ ;
	wire _w6343_ ;
	wire _w6344_ ;
	wire _w6345_ ;
	wire _w6346_ ;
	wire _w6347_ ;
	wire _w6348_ ;
	wire _w6349_ ;
	wire _w6350_ ;
	wire _w6351_ ;
	wire _w6352_ ;
	wire _w6353_ ;
	wire _w6354_ ;
	wire _w6355_ ;
	wire _w6356_ ;
	wire _w6357_ ;
	wire _w6358_ ;
	wire _w6359_ ;
	wire _w6360_ ;
	wire _w6361_ ;
	wire _w6362_ ;
	wire _w6363_ ;
	wire _w6364_ ;
	wire _w6365_ ;
	wire _w6366_ ;
	wire _w6367_ ;
	wire _w6368_ ;
	wire _w6369_ ;
	wire _w6370_ ;
	wire _w6371_ ;
	wire _w6372_ ;
	wire _w6373_ ;
	wire _w6374_ ;
	wire _w6375_ ;
	wire _w6376_ ;
	wire _w6377_ ;
	wire _w6378_ ;
	wire _w6379_ ;
	wire _w6380_ ;
	wire _w6381_ ;
	wire _w6382_ ;
	wire _w6383_ ;
	wire _w6384_ ;
	wire _w6385_ ;
	wire _w6386_ ;
	wire _w6387_ ;
	wire _w6388_ ;
	wire _w6389_ ;
	wire _w6390_ ;
	wire _w6391_ ;
	wire _w6392_ ;
	wire _w6393_ ;
	wire _w6394_ ;
	wire _w6395_ ;
	wire _w6396_ ;
	wire _w6397_ ;
	wire _w6398_ ;
	wire _w6399_ ;
	wire _w6400_ ;
	wire _w6401_ ;
	wire _w6402_ ;
	wire _w6403_ ;
	wire _w6404_ ;
	wire _w6405_ ;
	wire _w6406_ ;
	wire _w6407_ ;
	wire _w6408_ ;
	wire _w6409_ ;
	wire _w6410_ ;
	wire _w6411_ ;
	wire _w6412_ ;
	wire _w6413_ ;
	wire _w6414_ ;
	wire _w6415_ ;
	wire _w6416_ ;
	wire _w6417_ ;
	wire _w6418_ ;
	wire _w6419_ ;
	wire _w6420_ ;
	wire _w6421_ ;
	wire _w6422_ ;
	wire _w6423_ ;
	wire _w6424_ ;
	wire _w6425_ ;
	wire _w6426_ ;
	wire _w6427_ ;
	wire _w6428_ ;
	wire _w6429_ ;
	wire _w6430_ ;
	wire _w6431_ ;
	wire _w6432_ ;
	wire _w6433_ ;
	wire _w6434_ ;
	wire _w6435_ ;
	wire _w6436_ ;
	wire _w6437_ ;
	wire _w6438_ ;
	wire _w6439_ ;
	wire _w6440_ ;
	wire _w6441_ ;
	wire _w6442_ ;
	wire _w6443_ ;
	wire _w6444_ ;
	wire _w6445_ ;
	wire _w6446_ ;
	wire _w6447_ ;
	wire _w6448_ ;
	wire _w6449_ ;
	wire _w6450_ ;
	wire _w6451_ ;
	wire _w6452_ ;
	wire _w6453_ ;
	wire _w6454_ ;
	wire _w6455_ ;
	wire _w6456_ ;
	wire _w6457_ ;
	wire _w6458_ ;
	wire _w6459_ ;
	wire _w6460_ ;
	wire _w6461_ ;
	wire _w6462_ ;
	wire _w6463_ ;
	wire _w6464_ ;
	wire _w6465_ ;
	wire _w6466_ ;
	wire _w6467_ ;
	wire _w6468_ ;
	wire _w6469_ ;
	wire _w6470_ ;
	wire _w6471_ ;
	wire _w6472_ ;
	wire _w6473_ ;
	wire _w6474_ ;
	wire _w6475_ ;
	wire _w6476_ ;
	wire _w6477_ ;
	wire _w6478_ ;
	wire _w6479_ ;
	wire _w6480_ ;
	wire _w6481_ ;
	wire _w6482_ ;
	wire _w6483_ ;
	wire _w6484_ ;
	wire _w6485_ ;
	wire _w6486_ ;
	wire _w6487_ ;
	wire _w6488_ ;
	wire _w6489_ ;
	wire _w6490_ ;
	wire _w6491_ ;
	wire _w6492_ ;
	wire _w6493_ ;
	wire _w6494_ ;
	wire _w6495_ ;
	wire _w6496_ ;
	wire _w6497_ ;
	wire _w6498_ ;
	wire _w6499_ ;
	wire _w6500_ ;
	wire _w6501_ ;
	wire _w6502_ ;
	wire _w6503_ ;
	wire _w6504_ ;
	wire _w6505_ ;
	wire _w6506_ ;
	wire _w6507_ ;
	wire _w6508_ ;
	wire _w6509_ ;
	wire _w6510_ ;
	wire _w6511_ ;
	wire _w6512_ ;
	wire _w6513_ ;
	wire _w6514_ ;
	wire _w6515_ ;
	wire _w6516_ ;
	wire _w6517_ ;
	wire _w6518_ ;
	wire _w6519_ ;
	wire _w6520_ ;
	wire _w6521_ ;
	wire _w6522_ ;
	wire _w6523_ ;
	wire _w6524_ ;
	wire _w6525_ ;
	wire _w6526_ ;
	wire _w6527_ ;
	wire _w6528_ ;
	wire _w6529_ ;
	wire _w6530_ ;
	wire _w6531_ ;
	wire _w6532_ ;
	wire _w6533_ ;
	wire _w6534_ ;
	wire _w6535_ ;
	wire _w6536_ ;
	wire _w6537_ ;
	wire _w6538_ ;
	wire _w6539_ ;
	wire _w6540_ ;
	wire _w6541_ ;
	wire _w6542_ ;
	wire _w6543_ ;
	wire _w6544_ ;
	wire _w6545_ ;
	wire _w6546_ ;
	wire _w6547_ ;
	wire _w6548_ ;
	wire _w6549_ ;
	wire _w6550_ ;
	wire _w6551_ ;
	wire _w6552_ ;
	wire _w6553_ ;
	wire _w6554_ ;
	wire _w6555_ ;
	wire _w6556_ ;
	wire _w6557_ ;
	wire _w6558_ ;
	wire _w6559_ ;
	wire _w6560_ ;
	wire _w6561_ ;
	wire _w6562_ ;
	wire _w6563_ ;
	wire _w6564_ ;
	wire _w6565_ ;
	wire _w6566_ ;
	wire _w6567_ ;
	wire _w6568_ ;
	wire _w6569_ ;
	wire _w6570_ ;
	wire _w6571_ ;
	wire _w6572_ ;
	wire _w6573_ ;
	wire _w6574_ ;
	wire _w6575_ ;
	wire _w6576_ ;
	wire _w6577_ ;
	wire _w6578_ ;
	wire _w6579_ ;
	wire _w6580_ ;
	wire _w6581_ ;
	wire _w6582_ ;
	wire _w6583_ ;
	wire _w6584_ ;
	wire _w6585_ ;
	wire _w6586_ ;
	wire _w6587_ ;
	wire _w6588_ ;
	wire _w6589_ ;
	wire _w6590_ ;
	wire _w6591_ ;
	wire _w6592_ ;
	wire _w6593_ ;
	wire _w6594_ ;
	wire _w6595_ ;
	wire _w6596_ ;
	wire _w6597_ ;
	wire _w6598_ ;
	wire _w6599_ ;
	wire _w6600_ ;
	wire _w6601_ ;
	wire _w6602_ ;
	wire _w6603_ ;
	wire _w6604_ ;
	wire _w6605_ ;
	wire _w6606_ ;
	wire _w6607_ ;
	wire _w6608_ ;
	wire _w6609_ ;
	wire _w6610_ ;
	wire _w6611_ ;
	wire _w6612_ ;
	wire _w6613_ ;
	wire _w6614_ ;
	wire _w6615_ ;
	wire _w6616_ ;
	wire _w6617_ ;
	wire _w6618_ ;
	wire _w6619_ ;
	wire _w6620_ ;
	wire _w6621_ ;
	wire _w6622_ ;
	wire _w6623_ ;
	wire _w6624_ ;
	wire _w6625_ ;
	wire _w6626_ ;
	wire _w6627_ ;
	wire _w6628_ ;
	wire _w6629_ ;
	wire _w6630_ ;
	wire _w6631_ ;
	wire _w6632_ ;
	wire _w6633_ ;
	wire _w6634_ ;
	wire _w6635_ ;
	wire _w6636_ ;
	wire _w6637_ ;
	wire _w6638_ ;
	wire _w6639_ ;
	wire _w6640_ ;
	wire _w6641_ ;
	wire _w6642_ ;
	wire _w6643_ ;
	wire _w6644_ ;
	wire _w6645_ ;
	wire _w6646_ ;
	wire _w6647_ ;
	wire _w6648_ ;
	wire _w6649_ ;
	wire _w6650_ ;
	wire _w6651_ ;
	wire _w6652_ ;
	wire _w6653_ ;
	wire _w6654_ ;
	wire _w6655_ ;
	wire _w6656_ ;
	wire _w6657_ ;
	wire _w6658_ ;
	wire _w6659_ ;
	wire _w6660_ ;
	wire _w6661_ ;
	wire _w6662_ ;
	wire _w6663_ ;
	wire _w6664_ ;
	wire _w6665_ ;
	wire _w6666_ ;
	wire _w6667_ ;
	wire _w6668_ ;
	wire _w6669_ ;
	wire _w6670_ ;
	wire _w6671_ ;
	wire _w6672_ ;
	wire _w6673_ ;
	wire _w6674_ ;
	wire _w6675_ ;
	wire _w6676_ ;
	wire _w6677_ ;
	wire _w6678_ ;
	wire _w6679_ ;
	wire _w6680_ ;
	wire _w6681_ ;
	wire _w6682_ ;
	wire _w6683_ ;
	wire _w6684_ ;
	wire _w6685_ ;
	wire _w6686_ ;
	wire _w6687_ ;
	wire _w6688_ ;
	wire _w6689_ ;
	wire _w6690_ ;
	wire _w6691_ ;
	wire _w6692_ ;
	wire _w6693_ ;
	wire _w6694_ ;
	wire _w6695_ ;
	wire _w6696_ ;
	wire _w6697_ ;
	wire _w6698_ ;
	wire _w6699_ ;
	wire _w6700_ ;
	wire _w6701_ ;
	wire _w6702_ ;
	wire _w6703_ ;
	wire _w6704_ ;
	wire _w6705_ ;
	wire _w6706_ ;
	wire _w6707_ ;
	wire _w6708_ ;
	wire _w6709_ ;
	wire _w6710_ ;
	wire _w6711_ ;
	wire _w6712_ ;
	wire _w6713_ ;
	wire _w6714_ ;
	wire _w6715_ ;
	wire _w6716_ ;
	wire _w6717_ ;
	wire _w6718_ ;
	wire _w6719_ ;
	wire _w6720_ ;
	wire _w6721_ ;
	wire _w6722_ ;
	wire _w6723_ ;
	wire _w6724_ ;
	wire _w6725_ ;
	wire _w6726_ ;
	wire _w6727_ ;
	wire _w6728_ ;
	wire _w6729_ ;
	wire _w6730_ ;
	wire _w6731_ ;
	wire _w6732_ ;
	wire _w6733_ ;
	wire _w6734_ ;
	wire _w6735_ ;
	wire _w6736_ ;
	wire _w6737_ ;
	wire _w6738_ ;
	wire _w6739_ ;
	wire _w6740_ ;
	wire _w6741_ ;
	wire _w6742_ ;
	wire _w6743_ ;
	wire _w6744_ ;
	wire _w6745_ ;
	wire _w6746_ ;
	wire _w6747_ ;
	wire _w6748_ ;
	wire _w6749_ ;
	wire _w6750_ ;
	wire _w6751_ ;
	wire _w6752_ ;
	wire _w6753_ ;
	wire _w6754_ ;
	wire _w6755_ ;
	wire _w6756_ ;
	wire _w6757_ ;
	wire _w6758_ ;
	wire _w6759_ ;
	wire _w6760_ ;
	wire _w6761_ ;
	wire _w6762_ ;
	wire _w6763_ ;
	wire _w6764_ ;
	wire _w6765_ ;
	wire _w6766_ ;
	wire _w6767_ ;
	wire _w6768_ ;
	wire _w6769_ ;
	wire _w6770_ ;
	wire _w6771_ ;
	wire _w6772_ ;
	wire _w6773_ ;
	wire _w6774_ ;
	wire _w6775_ ;
	wire _w6776_ ;
	wire _w6777_ ;
	wire _w6778_ ;
	wire _w6779_ ;
	wire _w6780_ ;
	wire _w6781_ ;
	wire _w6782_ ;
	wire _w6783_ ;
	wire _w6784_ ;
	wire _w6785_ ;
	wire _w6786_ ;
	wire _w6787_ ;
	wire _w6788_ ;
	wire _w6789_ ;
	wire _w6790_ ;
	wire _w6791_ ;
	wire _w6792_ ;
	wire _w6793_ ;
	wire _w6794_ ;
	wire _w6795_ ;
	wire _w6796_ ;
	wire _w6797_ ;
	wire _w6798_ ;
	wire _w6799_ ;
	wire _w6800_ ;
	wire _w6801_ ;
	wire _w6802_ ;
	wire _w6803_ ;
	wire _w6804_ ;
	wire _w6805_ ;
	wire _w6806_ ;
	wire _w6807_ ;
	wire _w6808_ ;
	wire _w6809_ ;
	wire _w6810_ ;
	wire _w6811_ ;
	wire _w6812_ ;
	wire _w6813_ ;
	wire _w6814_ ;
	wire _w6815_ ;
	wire _w6816_ ;
	wire _w6817_ ;
	wire _w6818_ ;
	wire _w6819_ ;
	wire _w6820_ ;
	wire _w6821_ ;
	wire _w6822_ ;
	wire _w6823_ ;
	wire _w6824_ ;
	wire _w6825_ ;
	wire _w6826_ ;
	wire _w6827_ ;
	wire _w6828_ ;
	wire _w6829_ ;
	wire _w6830_ ;
	wire _w6831_ ;
	wire _w6832_ ;
	wire _w6833_ ;
	wire _w6834_ ;
	wire _w6835_ ;
	wire _w6836_ ;
	wire _w6837_ ;
	wire _w6838_ ;
	wire _w6839_ ;
	wire _w6840_ ;
	wire _w6841_ ;
	wire _w6842_ ;
	wire _w6843_ ;
	wire _w6844_ ;
	wire _w6845_ ;
	wire _w6846_ ;
	wire _w6847_ ;
	wire _w6848_ ;
	wire _w6849_ ;
	wire _w6850_ ;
	wire _w6851_ ;
	wire _w6852_ ;
	wire _w6853_ ;
	wire _w6854_ ;
	wire _w6855_ ;
	wire _w6856_ ;
	wire _w6857_ ;
	wire _w6858_ ;
	wire _w6859_ ;
	wire _w6860_ ;
	wire _w6861_ ;
	wire _w6862_ ;
	wire _w6863_ ;
	wire _w6864_ ;
	wire _w6865_ ;
	wire _w6866_ ;
	wire _w6867_ ;
	wire _w6868_ ;
	wire _w6869_ ;
	wire _w6870_ ;
	wire _w6871_ ;
	wire _w6872_ ;
	wire _w6873_ ;
	wire _w6874_ ;
	wire _w6875_ ;
	wire _w6876_ ;
	wire _w6877_ ;
	wire _w6878_ ;
	wire _w6879_ ;
	wire _w6880_ ;
	wire _w6881_ ;
	wire _w6882_ ;
	wire _w6883_ ;
	wire _w6884_ ;
	wire _w6885_ ;
	wire _w6886_ ;
	wire _w6887_ ;
	wire _w6888_ ;
	wire _w6889_ ;
	wire _w6890_ ;
	wire _w6891_ ;
	wire _w6892_ ;
	wire _w6893_ ;
	wire _w6894_ ;
	wire _w6895_ ;
	wire _w6896_ ;
	wire _w6897_ ;
	wire _w6898_ ;
	wire _w6899_ ;
	wire _w6900_ ;
	wire _w6901_ ;
	wire _w6902_ ;
	wire _w6903_ ;
	wire _w6904_ ;
	wire _w6905_ ;
	wire _w6906_ ;
	wire _w6907_ ;
	wire _w6908_ ;
	wire _w6909_ ;
	wire _w6910_ ;
	wire _w6911_ ;
	wire _w6912_ ;
	wire _w6913_ ;
	wire _w6914_ ;
	wire _w6915_ ;
	wire _w6916_ ;
	wire _w6917_ ;
	wire _w6918_ ;
	wire _w6919_ ;
	wire _w6920_ ;
	wire _w6921_ ;
	wire _w6922_ ;
	wire _w6923_ ;
	wire _w6924_ ;
	wire _w6925_ ;
	wire _w6926_ ;
	wire _w6927_ ;
	wire _w6928_ ;
	wire _w6929_ ;
	wire _w6930_ ;
	wire _w6931_ ;
	wire _w6932_ ;
	wire _w6933_ ;
	wire _w6934_ ;
	wire _w6935_ ;
	wire _w6936_ ;
	wire _w6937_ ;
	wire _w6938_ ;
	wire _w6939_ ;
	wire _w6940_ ;
	wire _w6941_ ;
	wire _w6942_ ;
	wire _w6943_ ;
	wire _w6944_ ;
	wire _w6945_ ;
	wire _w6946_ ;
	wire _w6947_ ;
	wire _w6948_ ;
	wire _w6949_ ;
	wire _w6950_ ;
	wire _w6951_ ;
	wire _w6952_ ;
	wire _w6953_ ;
	wire _w6954_ ;
	wire _w6955_ ;
	wire _w6956_ ;
	wire _w6957_ ;
	wire _w6958_ ;
	wire _w6959_ ;
	wire _w6960_ ;
	wire _w6961_ ;
	wire _w6962_ ;
	wire _w6963_ ;
	wire _w6964_ ;
	wire _w6965_ ;
	wire _w6966_ ;
	wire _w6967_ ;
	wire _w6968_ ;
	wire _w6969_ ;
	wire _w6970_ ;
	wire _w6971_ ;
	wire _w6972_ ;
	wire _w6973_ ;
	wire _w6974_ ;
	wire _w6975_ ;
	wire _w6976_ ;
	wire _w6977_ ;
	wire _w6978_ ;
	wire _w6979_ ;
	wire _w6980_ ;
	wire _w6981_ ;
	wire _w6982_ ;
	wire _w6983_ ;
	wire _w6984_ ;
	wire _w6985_ ;
	wire _w6986_ ;
	wire _w6987_ ;
	wire _w6988_ ;
	wire _w6989_ ;
	wire _w6990_ ;
	wire _w6991_ ;
	wire _w6992_ ;
	wire _w6993_ ;
	wire _w6994_ ;
	wire _w6995_ ;
	wire _w6996_ ;
	wire _w6997_ ;
	wire _w6998_ ;
	wire _w6999_ ;
	wire _w7000_ ;
	wire _w7001_ ;
	wire _w7002_ ;
	wire _w7003_ ;
	wire _w7004_ ;
	wire _w7005_ ;
	wire _w7006_ ;
	wire _w7007_ ;
	wire _w7008_ ;
	wire _w7009_ ;
	wire _w7010_ ;
	wire _w7011_ ;
	wire _w7012_ ;
	wire _w7013_ ;
	wire _w7014_ ;
	wire _w7015_ ;
	wire _w7016_ ;
	wire _w7017_ ;
	wire _w7018_ ;
	wire _w7019_ ;
	wire _w7020_ ;
	wire _w7021_ ;
	wire _w7022_ ;
	wire _w7023_ ;
	wire _w7024_ ;
	wire _w7025_ ;
	wire _w7026_ ;
	wire _w7027_ ;
	wire _w7028_ ;
	wire _w7029_ ;
	wire _w7030_ ;
	wire _w7031_ ;
	wire _w7032_ ;
	wire _w7033_ ;
	wire _w7034_ ;
	wire _w7035_ ;
	wire _w7036_ ;
	wire _w7037_ ;
	wire _w7038_ ;
	wire _w7039_ ;
	wire _w7040_ ;
	wire _w7041_ ;
	wire _w7042_ ;
	wire _w7043_ ;
	wire _w7044_ ;
	wire _w7045_ ;
	wire _w7046_ ;
	wire _w7047_ ;
	wire _w7048_ ;
	wire _w7049_ ;
	wire _w7050_ ;
	wire _w7051_ ;
	wire _w7052_ ;
	wire _w7053_ ;
	wire _w7054_ ;
	wire _w7055_ ;
	wire _w7056_ ;
	wire _w7057_ ;
	wire _w7058_ ;
	wire _w7059_ ;
	wire _w7060_ ;
	wire _w7061_ ;
	wire _w7062_ ;
	wire _w7063_ ;
	wire _w7064_ ;
	wire _w7065_ ;
	wire _w7066_ ;
	wire _w7067_ ;
	wire _w7068_ ;
	wire _w7069_ ;
	wire _w7070_ ;
	wire _w7071_ ;
	wire _w7072_ ;
	wire _w7073_ ;
	wire _w7074_ ;
	wire _w7075_ ;
	wire _w7076_ ;
	wire _w7077_ ;
	wire _w7078_ ;
	wire _w7079_ ;
	wire _w7080_ ;
	wire _w7081_ ;
	wire _w7082_ ;
	wire _w7083_ ;
	wire _w7084_ ;
	wire _w7085_ ;
	wire _w7086_ ;
	wire _w7087_ ;
	wire _w7088_ ;
	wire _w7089_ ;
	wire _w7090_ ;
	wire _w7091_ ;
	wire _w7092_ ;
	wire _w7093_ ;
	wire _w7094_ ;
	wire _w7095_ ;
	wire _w7096_ ;
	wire _w7097_ ;
	wire _w7098_ ;
	wire _w7099_ ;
	wire _w7100_ ;
	wire _w7101_ ;
	wire _w7102_ ;
	wire _w7103_ ;
	wire _w7104_ ;
	wire _w7105_ ;
	wire _w7106_ ;
	wire _w7107_ ;
	wire _w7108_ ;
	wire _w7109_ ;
	wire _w7110_ ;
	wire _w7111_ ;
	wire _w7112_ ;
	wire _w7113_ ;
	wire _w7114_ ;
	wire _w7115_ ;
	wire _w7116_ ;
	wire _w7117_ ;
	wire _w7118_ ;
	wire _w7119_ ;
	wire _w7120_ ;
	wire _w7121_ ;
	wire _w7122_ ;
	wire _w7123_ ;
	wire _w7124_ ;
	wire _w7125_ ;
	wire _w7126_ ;
	wire _w7127_ ;
	wire _w7128_ ;
	wire _w7129_ ;
	wire _w7130_ ;
	wire _w7131_ ;
	wire _w7132_ ;
	wire _w7133_ ;
	wire _w7134_ ;
	wire _w7135_ ;
	wire _w7136_ ;
	wire _w7137_ ;
	wire _w7138_ ;
	wire _w7139_ ;
	wire _w7140_ ;
	wire _w7141_ ;
	wire _w7142_ ;
	wire _w7143_ ;
	wire _w7144_ ;
	wire _w7145_ ;
	wire _w7146_ ;
	wire _w7147_ ;
	wire _w7148_ ;
	wire _w7149_ ;
	wire _w7150_ ;
	wire _w7151_ ;
	wire _w7152_ ;
	wire _w7153_ ;
	wire _w7154_ ;
	wire _w7155_ ;
	wire _w7156_ ;
	wire _w7157_ ;
	wire _w7158_ ;
	wire _w7159_ ;
	wire _w7160_ ;
	wire _w7161_ ;
	wire _w7162_ ;
	wire _w7163_ ;
	wire _w7164_ ;
	wire _w7165_ ;
	wire _w7166_ ;
	wire _w7167_ ;
	wire _w7168_ ;
	wire _w7169_ ;
	wire _w7170_ ;
	wire _w7171_ ;
	wire _w7172_ ;
	wire _w7173_ ;
	wire _w7174_ ;
	wire _w7175_ ;
	wire _w7176_ ;
	wire _w7177_ ;
	wire _w7178_ ;
	wire _w7179_ ;
	wire _w7180_ ;
	wire _w7181_ ;
	wire _w7182_ ;
	wire _w7183_ ;
	wire _w7184_ ;
	wire _w7185_ ;
	wire _w7186_ ;
	wire _w7187_ ;
	wire _w7188_ ;
	wire _w7189_ ;
	wire _w7190_ ;
	wire _w7191_ ;
	wire _w7192_ ;
	wire _w7193_ ;
	wire _w7194_ ;
	wire _w7195_ ;
	wire _w7196_ ;
	wire _w7197_ ;
	wire _w7198_ ;
	wire _w7199_ ;
	wire _w7200_ ;
	wire _w7201_ ;
	wire _w7202_ ;
	wire _w7203_ ;
	wire _w7204_ ;
	wire _w7205_ ;
	wire _w7206_ ;
	wire _w7207_ ;
	wire _w7208_ ;
	wire _w7209_ ;
	wire _w7210_ ;
	wire _w7211_ ;
	wire _w7212_ ;
	wire _w7213_ ;
	wire _w7214_ ;
	wire _w7215_ ;
	wire _w7216_ ;
	wire _w7217_ ;
	wire _w7218_ ;
	wire _w7219_ ;
	wire _w7220_ ;
	wire _w7221_ ;
	wire _w7222_ ;
	wire _w7223_ ;
	wire _w7224_ ;
	wire _w7225_ ;
	wire _w7226_ ;
	wire _w7227_ ;
	wire _w7228_ ;
	wire _w7229_ ;
	wire _w7230_ ;
	wire _w7231_ ;
	wire _w7232_ ;
	wire _w7233_ ;
	wire _w7234_ ;
	wire _w7235_ ;
	wire _w7236_ ;
	wire _w7237_ ;
	wire _w7238_ ;
	wire _w7239_ ;
	wire _w7240_ ;
	wire _w7241_ ;
	wire _w7242_ ;
	wire _w7243_ ;
	wire _w7244_ ;
	wire _w7245_ ;
	wire _w7246_ ;
	wire _w7247_ ;
	wire _w7248_ ;
	wire _w7249_ ;
	wire _w7250_ ;
	wire _w7251_ ;
	wire _w7252_ ;
	wire _w7253_ ;
	wire _w7254_ ;
	wire _w7255_ ;
	wire _w7256_ ;
	wire _w7257_ ;
	wire _w7258_ ;
	wire _w7259_ ;
	wire _w7260_ ;
	wire _w7261_ ;
	wire _w7262_ ;
	wire _w7263_ ;
	wire _w7264_ ;
	wire _w7265_ ;
	wire _w7266_ ;
	wire _w7267_ ;
	wire _w7268_ ;
	wire _w7269_ ;
	wire _w7270_ ;
	wire _w7271_ ;
	wire _w7272_ ;
	wire _w7273_ ;
	wire _w7274_ ;
	wire _w7275_ ;
	wire _w7276_ ;
	wire _w7277_ ;
	wire _w7278_ ;
	wire _w7279_ ;
	wire _w7280_ ;
	wire _w7281_ ;
	wire _w7282_ ;
	wire _w7283_ ;
	wire _w7284_ ;
	wire _w7285_ ;
	wire _w7286_ ;
	wire _w7287_ ;
	wire _w7288_ ;
	wire _w7289_ ;
	wire _w7290_ ;
	wire _w7291_ ;
	wire _w7292_ ;
	wire _w7293_ ;
	wire _w7294_ ;
	wire _w7295_ ;
	wire _w7296_ ;
	wire _w7297_ ;
	wire _w7298_ ;
	wire _w7299_ ;
	wire _w7300_ ;
	wire _w7301_ ;
	wire _w7302_ ;
	wire _w7303_ ;
	wire _w7304_ ;
	wire _w7305_ ;
	wire _w7306_ ;
	wire _w7307_ ;
	wire _w7308_ ;
	wire _w7309_ ;
	wire _w7310_ ;
	wire _w7311_ ;
	wire _w7312_ ;
	wire _w7313_ ;
	wire _w7314_ ;
	wire _w7315_ ;
	wire _w7316_ ;
	wire _w7317_ ;
	wire _w7318_ ;
	wire _w7319_ ;
	wire _w7320_ ;
	wire _w7321_ ;
	wire _w7322_ ;
	wire _w7323_ ;
	wire _w7324_ ;
	wire _w7325_ ;
	wire _w7326_ ;
	wire _w7327_ ;
	wire _w7328_ ;
	wire _w7329_ ;
	wire _w7330_ ;
	wire _w7331_ ;
	wire _w7332_ ;
	wire _w7333_ ;
	wire _w7334_ ;
	wire _w7335_ ;
	wire _w7336_ ;
	wire _w7337_ ;
	wire _w7338_ ;
	wire _w7339_ ;
	wire _w7340_ ;
	wire _w7341_ ;
	wire _w7342_ ;
	wire _w7343_ ;
	wire _w7344_ ;
	wire _w7345_ ;
	wire _w7346_ ;
	wire _w7347_ ;
	wire _w7348_ ;
	wire _w7349_ ;
	wire _w7350_ ;
	wire _w7351_ ;
	wire _w7352_ ;
	wire _w7353_ ;
	wire _w7354_ ;
	wire _w7355_ ;
	wire _w7356_ ;
	wire _w7357_ ;
	wire _w7358_ ;
	wire _w7359_ ;
	wire _w7360_ ;
	wire _w7361_ ;
	wire _w7362_ ;
	wire _w7363_ ;
	wire _w7364_ ;
	wire _w7365_ ;
	wire _w7366_ ;
	wire _w7367_ ;
	wire _w7368_ ;
	wire _w7369_ ;
	wire _w7370_ ;
	wire _w7371_ ;
	wire _w7372_ ;
	wire _w7373_ ;
	wire _w7374_ ;
	wire _w7375_ ;
	wire _w7376_ ;
	wire _w7377_ ;
	wire _w7378_ ;
	wire _w7379_ ;
	wire _w7380_ ;
	wire _w7381_ ;
	wire _w7382_ ;
	wire _w7383_ ;
	wire _w7384_ ;
	wire _w7385_ ;
	wire _w7386_ ;
	wire _w7387_ ;
	wire _w7388_ ;
	wire _w7389_ ;
	wire _w7390_ ;
	wire _w7391_ ;
	wire _w7392_ ;
	wire _w7393_ ;
	wire _w7394_ ;
	wire _w7395_ ;
	wire _w7396_ ;
	wire _w7397_ ;
	wire _w7398_ ;
	wire _w7399_ ;
	wire _w7400_ ;
	wire _w7401_ ;
	wire _w7402_ ;
	wire _w7403_ ;
	wire _w7404_ ;
	wire _w7405_ ;
	wire _w7406_ ;
	wire _w7407_ ;
	wire _w7408_ ;
	wire _w7409_ ;
	wire _w7410_ ;
	wire _w7411_ ;
	wire _w7412_ ;
	wire _w7413_ ;
	wire _w7414_ ;
	wire _w7415_ ;
	wire _w7416_ ;
	wire _w7417_ ;
	wire _w7418_ ;
	wire _w7419_ ;
	wire _w7420_ ;
	wire _w7421_ ;
	wire _w7422_ ;
	wire _w7423_ ;
	wire _w7424_ ;
	wire _w7425_ ;
	wire _w7426_ ;
	wire _w7427_ ;
	wire _w7428_ ;
	wire _w7429_ ;
	wire _w7430_ ;
	wire _w7431_ ;
	wire _w7432_ ;
	wire _w7433_ ;
	wire _w7434_ ;
	wire _w7435_ ;
	wire _w7436_ ;
	wire _w7437_ ;
	wire _w7438_ ;
	wire _w7439_ ;
	wire _w7440_ ;
	wire _w7441_ ;
	wire _w7442_ ;
	wire _w7443_ ;
	wire _w7444_ ;
	wire _w7445_ ;
	wire _w7446_ ;
	wire _w7447_ ;
	wire _w7448_ ;
	wire _w7449_ ;
	wire _w7450_ ;
	wire _w7451_ ;
	wire _w7452_ ;
	wire _w7453_ ;
	wire _w7454_ ;
	wire _w7455_ ;
	wire _w7456_ ;
	wire _w7457_ ;
	wire _w7458_ ;
	wire _w7459_ ;
	wire _w7460_ ;
	wire _w7461_ ;
	wire _w7462_ ;
	wire _w7463_ ;
	wire _w7464_ ;
	wire _w7465_ ;
	wire _w7466_ ;
	wire _w7467_ ;
	wire _w7468_ ;
	wire _w7469_ ;
	wire _w7470_ ;
	wire _w7471_ ;
	wire _w7472_ ;
	wire _w7473_ ;
	wire _w7474_ ;
	wire _w7475_ ;
	wire _w7476_ ;
	wire _w7477_ ;
	wire _w7478_ ;
	wire _w7479_ ;
	wire _w7480_ ;
	wire _w7481_ ;
	wire _w7482_ ;
	wire _w7483_ ;
	wire _w7484_ ;
	wire _w7485_ ;
	wire _w7486_ ;
	wire _w7487_ ;
	wire _w7488_ ;
	wire _w7489_ ;
	wire _w7490_ ;
	wire _w7491_ ;
	wire _w7492_ ;
	wire _w7493_ ;
	wire _w7494_ ;
	wire _w7495_ ;
	wire _w7496_ ;
	wire _w7497_ ;
	wire _w7498_ ;
	wire _w7499_ ;
	wire _w7500_ ;
	wire _w7501_ ;
	wire _w7502_ ;
	wire _w7503_ ;
	wire _w7504_ ;
	wire _w7505_ ;
	wire _w7506_ ;
	wire _w7507_ ;
	wire _w7508_ ;
	wire _w7509_ ;
	wire _w7510_ ;
	wire _w7511_ ;
	wire _w7512_ ;
	wire _w7513_ ;
	wire _w7514_ ;
	wire _w7515_ ;
	wire _w7516_ ;
	wire _w7517_ ;
	wire _w7518_ ;
	wire _w7519_ ;
	wire _w7520_ ;
	wire _w7521_ ;
	wire _w7522_ ;
	wire _w7523_ ;
	wire _w7524_ ;
	wire _w7525_ ;
	wire _w7526_ ;
	wire _w7527_ ;
	wire _w7528_ ;
	wire _w7529_ ;
	wire _w7530_ ;
	wire _w7531_ ;
	wire _w7532_ ;
	wire _w7533_ ;
	wire _w7534_ ;
	wire _w7535_ ;
	wire _w7536_ ;
	wire _w7537_ ;
	wire _w7538_ ;
	wire _w7539_ ;
	wire _w7540_ ;
	wire _w7541_ ;
	wire _w7542_ ;
	wire _w7543_ ;
	wire _w7544_ ;
	wire _w7545_ ;
	wire _w7546_ ;
	wire _w7547_ ;
	wire _w7548_ ;
	wire _w7549_ ;
	wire _w7550_ ;
	wire _w7551_ ;
	wire _w7552_ ;
	wire _w7553_ ;
	wire _w7554_ ;
	wire _w7555_ ;
	wire _w7556_ ;
	wire _w7557_ ;
	wire _w7558_ ;
	wire _w7559_ ;
	wire _w7560_ ;
	wire _w7561_ ;
	wire _w7562_ ;
	wire _w7563_ ;
	wire _w7564_ ;
	wire _w7565_ ;
	wire _w7566_ ;
	wire _w7567_ ;
	wire _w7568_ ;
	wire _w7569_ ;
	wire _w7570_ ;
	wire _w7571_ ;
	wire _w7572_ ;
	wire _w7573_ ;
	wire _w7574_ ;
	wire _w7575_ ;
	wire _w7576_ ;
	wire _w7577_ ;
	wire _w7578_ ;
	wire _w7579_ ;
	wire _w7580_ ;
	wire _w7581_ ;
	wire _w7582_ ;
	wire _w7583_ ;
	wire _w7584_ ;
	wire _w7585_ ;
	wire _w7586_ ;
	wire _w7587_ ;
	wire _w7588_ ;
	wire _w7589_ ;
	wire _w7590_ ;
	wire _w7591_ ;
	wire _w7592_ ;
	wire _w7593_ ;
	wire _w7594_ ;
	wire _w7595_ ;
	wire _w7596_ ;
	wire _w7597_ ;
	wire _w7598_ ;
	wire _w7599_ ;
	wire _w7600_ ;
	wire _w7601_ ;
	wire _w7602_ ;
	wire _w7603_ ;
	wire _w7604_ ;
	wire _w7605_ ;
	wire _w7606_ ;
	wire _w7607_ ;
	wire _w7608_ ;
	wire _w7609_ ;
	wire _w7610_ ;
	wire _w7611_ ;
	wire _w7612_ ;
	wire _w7613_ ;
	wire _w7614_ ;
	wire _w7615_ ;
	wire _w7616_ ;
	wire _w7617_ ;
	wire _w7618_ ;
	wire _w7619_ ;
	wire _w7620_ ;
	wire _w7621_ ;
	wire _w7622_ ;
	wire _w7623_ ;
	wire _w7624_ ;
	wire _w7625_ ;
	wire _w7626_ ;
	wire _w7627_ ;
	wire _w7628_ ;
	wire _w7629_ ;
	wire _w7630_ ;
	wire _w7631_ ;
	wire _w7632_ ;
	wire _w7633_ ;
	wire _w7634_ ;
	wire _w7635_ ;
	wire _w7636_ ;
	wire _w7637_ ;
	wire _w7638_ ;
	wire _w7639_ ;
	wire _w7640_ ;
	wire _w7641_ ;
	wire _w7642_ ;
	wire _w7643_ ;
	wire _w7644_ ;
	wire _w7645_ ;
	wire _w7646_ ;
	wire _w7647_ ;
	wire _w7648_ ;
	wire _w7649_ ;
	wire _w7650_ ;
	wire _w7651_ ;
	wire _w7652_ ;
	wire _w7653_ ;
	wire _w7654_ ;
	wire _w7655_ ;
	wire _w7656_ ;
	wire _w7657_ ;
	wire _w7658_ ;
	wire _w7659_ ;
	wire _w7660_ ;
	wire _w7661_ ;
	wire _w7662_ ;
	wire _w7663_ ;
	wire _w7664_ ;
	wire _w7665_ ;
	wire _w7666_ ;
	wire _w7667_ ;
	wire _w7668_ ;
	wire _w7669_ ;
	wire _w7670_ ;
	wire _w7671_ ;
	wire _w7672_ ;
	wire _w7673_ ;
	wire _w7674_ ;
	wire _w7675_ ;
	wire _w7676_ ;
	wire _w7677_ ;
	wire _w7678_ ;
	wire _w7679_ ;
	wire _w7680_ ;
	wire _w7681_ ;
	wire _w7682_ ;
	wire _w7683_ ;
	wire _w7684_ ;
	wire _w7685_ ;
	wire _w7686_ ;
	wire _w7687_ ;
	wire _w7688_ ;
	wire _w7689_ ;
	wire _w7690_ ;
	wire _w7691_ ;
	wire _w7692_ ;
	wire _w7693_ ;
	wire _w7694_ ;
	wire _w7695_ ;
	wire _w7696_ ;
	wire _w7697_ ;
	wire _w7698_ ;
	wire _w7699_ ;
	wire _w7700_ ;
	wire _w7701_ ;
	wire _w7702_ ;
	wire _w7703_ ;
	wire _w7704_ ;
	wire _w7705_ ;
	wire _w7706_ ;
	wire _w7707_ ;
	wire _w7708_ ;
	wire _w7709_ ;
	wire _w7710_ ;
	wire _w7711_ ;
	wire _w7712_ ;
	wire _w7713_ ;
	wire _w7714_ ;
	wire _w7715_ ;
	wire _w7716_ ;
	wire _w7717_ ;
	wire _w7718_ ;
	wire _w7719_ ;
	wire _w7720_ ;
	wire _w7721_ ;
	wire _w7722_ ;
	wire _w7723_ ;
	wire _w7724_ ;
	wire _w7725_ ;
	wire _w7726_ ;
	wire _w7727_ ;
	wire _w7728_ ;
	wire _w7729_ ;
	wire _w7730_ ;
	wire _w7731_ ;
	wire _w7732_ ;
	wire _w7733_ ;
	wire _w7734_ ;
	wire _w7735_ ;
	wire _w7736_ ;
	wire _w7737_ ;
	wire _w7738_ ;
	wire _w7739_ ;
	wire _w7740_ ;
	wire _w7741_ ;
	wire _w7742_ ;
	wire _w7743_ ;
	wire _w7744_ ;
	wire _w7745_ ;
	wire _w7746_ ;
	wire _w7747_ ;
	wire _w7748_ ;
	wire _w7749_ ;
	wire _w7750_ ;
	wire _w7751_ ;
	wire _w7752_ ;
	wire _w7753_ ;
	wire _w7754_ ;
	wire _w7755_ ;
	wire _w7756_ ;
	wire _w7757_ ;
	wire _w7758_ ;
	wire _w7759_ ;
	wire _w7760_ ;
	wire _w7761_ ;
	wire _w7762_ ;
	wire _w7763_ ;
	wire _w7764_ ;
	wire _w7765_ ;
	wire _w7766_ ;
	wire _w7767_ ;
	wire _w7768_ ;
	wire _w7769_ ;
	wire _w7770_ ;
	wire _w7771_ ;
	wire _w7772_ ;
	wire _w7773_ ;
	wire _w7774_ ;
	wire _w7775_ ;
	wire _w7776_ ;
	wire _w7777_ ;
	wire _w7778_ ;
	wire _w7779_ ;
	wire _w7780_ ;
	wire _w7781_ ;
	wire _w7782_ ;
	wire _w7783_ ;
	wire _w7784_ ;
	wire _w7785_ ;
	wire _w7786_ ;
	wire _w7787_ ;
	wire _w7788_ ;
	wire _w7789_ ;
	wire _w7790_ ;
	wire _w7791_ ;
	wire _w7792_ ;
	wire _w7793_ ;
	wire _w7794_ ;
	wire _w7795_ ;
	wire _w7796_ ;
	wire _w7797_ ;
	wire _w7798_ ;
	wire _w7799_ ;
	wire _w7800_ ;
	wire _w7801_ ;
	wire _w7802_ ;
	wire _w7803_ ;
	wire _w7804_ ;
	wire _w7805_ ;
	wire _w7806_ ;
	wire _w7807_ ;
	wire _w7808_ ;
	wire _w7809_ ;
	wire _w7810_ ;
	wire _w7811_ ;
	wire _w7812_ ;
	wire _w7813_ ;
	wire _w7814_ ;
	wire _w7815_ ;
	wire _w7816_ ;
	wire _w7817_ ;
	wire _w7818_ ;
	wire _w7819_ ;
	wire _w7820_ ;
	wire _w7821_ ;
	wire _w7822_ ;
	wire _w7823_ ;
	wire _w7824_ ;
	wire _w7825_ ;
	wire _w7826_ ;
	wire _w7827_ ;
	wire _w7828_ ;
	wire _w7829_ ;
	wire _w7830_ ;
	wire _w7831_ ;
	wire _w7832_ ;
	wire _w7833_ ;
	wire _w7834_ ;
	wire _w7835_ ;
	wire _w7836_ ;
	wire _w7837_ ;
	wire _w7838_ ;
	wire _w7839_ ;
	wire _w7840_ ;
	wire _w7841_ ;
	wire _w7842_ ;
	wire _w7843_ ;
	wire _w7844_ ;
	wire _w7845_ ;
	wire _w7846_ ;
	wire _w7847_ ;
	wire _w7848_ ;
	wire _w7849_ ;
	wire _w7850_ ;
	wire _w7851_ ;
	wire _w7852_ ;
	wire _w7853_ ;
	wire _w7854_ ;
	wire _w7855_ ;
	wire _w7856_ ;
	wire _w7857_ ;
	wire _w7858_ ;
	wire _w7859_ ;
	wire _w7860_ ;
	wire _w7861_ ;
	wire _w7862_ ;
	wire _w7863_ ;
	wire _w7864_ ;
	wire _w7865_ ;
	wire _w7866_ ;
	wire _w7867_ ;
	wire _w7868_ ;
	wire _w7869_ ;
	wire _w7870_ ;
	wire _w7871_ ;
	wire _w7872_ ;
	wire _w7873_ ;
	wire _w7874_ ;
	wire _w7875_ ;
	wire _w7876_ ;
	wire _w7877_ ;
	wire _w7878_ ;
	wire _w7879_ ;
	wire _w7880_ ;
	wire _w7881_ ;
	wire _w7882_ ;
	wire _w7883_ ;
	wire _w7884_ ;
	wire _w7885_ ;
	wire _w7886_ ;
	wire _w7887_ ;
	wire _w7888_ ;
	wire _w7889_ ;
	wire _w7890_ ;
	wire _w7891_ ;
	wire _w7892_ ;
	wire _w7893_ ;
	wire _w7894_ ;
	wire _w7895_ ;
	wire _w7896_ ;
	wire _w7897_ ;
	wire _w7898_ ;
	wire _w7899_ ;
	wire _w7900_ ;
	wire _w7901_ ;
	wire _w7902_ ;
	wire _w7903_ ;
	wire _w7904_ ;
	wire _w7905_ ;
	wire _w7906_ ;
	wire _w7907_ ;
	wire _w7908_ ;
	wire _w7909_ ;
	wire _w7910_ ;
	wire _w7911_ ;
	wire _w7912_ ;
	wire _w7913_ ;
	wire _w7914_ ;
	wire _w7915_ ;
	wire _w7916_ ;
	wire _w7917_ ;
	wire _w7918_ ;
	wire _w7919_ ;
	wire _w7920_ ;
	wire _w7921_ ;
	wire _w7922_ ;
	wire _w7923_ ;
	wire _w7924_ ;
	wire _w7925_ ;
	wire _w7926_ ;
	wire _w7927_ ;
	wire _w7928_ ;
	wire _w7929_ ;
	wire _w7930_ ;
	wire _w7931_ ;
	wire _w7932_ ;
	wire _w7933_ ;
	wire _w7934_ ;
	wire _w7935_ ;
	wire _w7936_ ;
	wire _w7937_ ;
	wire _w7938_ ;
	wire _w7939_ ;
	wire _w7940_ ;
	wire _w7941_ ;
	wire _w7942_ ;
	wire _w7943_ ;
	wire _w7944_ ;
	wire _w7945_ ;
	wire _w7946_ ;
	wire _w7947_ ;
	wire _w7948_ ;
	wire _w7949_ ;
	wire _w7950_ ;
	wire _w7951_ ;
	wire _w7952_ ;
	wire _w7953_ ;
	wire _w7954_ ;
	wire _w7955_ ;
	wire _w7956_ ;
	wire _w7957_ ;
	wire _w7958_ ;
	wire _w7959_ ;
	wire _w7960_ ;
	wire _w7961_ ;
	wire _w7962_ ;
	wire _w7963_ ;
	wire _w7964_ ;
	wire _w7965_ ;
	wire _w7966_ ;
	wire _w7967_ ;
	wire _w7968_ ;
	wire _w7969_ ;
	wire _w7970_ ;
	wire _w7971_ ;
	wire _w7972_ ;
	wire _w7973_ ;
	wire _w7974_ ;
	wire _w7975_ ;
	wire _w7976_ ;
	wire _w7977_ ;
	wire _w7978_ ;
	wire _w7979_ ;
	wire _w7980_ ;
	wire _w7981_ ;
	wire _w7982_ ;
	wire _w7983_ ;
	wire _w7984_ ;
	wire _w7985_ ;
	wire _w7986_ ;
	wire _w7987_ ;
	wire _w7988_ ;
	wire _w7989_ ;
	wire _w7990_ ;
	wire _w7991_ ;
	wire _w7992_ ;
	wire _w7993_ ;
	wire _w7994_ ;
	wire _w7995_ ;
	wire _w7996_ ;
	wire _w7997_ ;
	wire _w7998_ ;
	wire _w7999_ ;
	wire _w8000_ ;
	wire _w8001_ ;
	wire _w8002_ ;
	wire _w8003_ ;
	wire _w8004_ ;
	wire _w8005_ ;
	wire _w8006_ ;
	wire _w8007_ ;
	wire _w8008_ ;
	wire _w8009_ ;
	wire _w8010_ ;
	wire _w8011_ ;
	wire _w8012_ ;
	wire _w8013_ ;
	wire _w8014_ ;
	wire _w8015_ ;
	wire _w8016_ ;
	wire _w8017_ ;
	wire _w8018_ ;
	wire _w8019_ ;
	wire _w8020_ ;
	wire _w8021_ ;
	wire _w8022_ ;
	wire _w8023_ ;
	wire _w8024_ ;
	wire _w8025_ ;
	wire _w8026_ ;
	wire _w8027_ ;
	wire _w8028_ ;
	wire _w8029_ ;
	wire _w8030_ ;
	wire _w8031_ ;
	wire _w8032_ ;
	wire _w8033_ ;
	wire _w8034_ ;
	wire _w8035_ ;
	wire _w8036_ ;
	wire _w8037_ ;
	wire _w8038_ ;
	wire _w8039_ ;
	wire _w8040_ ;
	wire _w8041_ ;
	wire _w8042_ ;
	wire _w8043_ ;
	wire _w8044_ ;
	wire _w8045_ ;
	wire _w8046_ ;
	wire _w8047_ ;
	wire _w8048_ ;
	wire _w8049_ ;
	wire _w8050_ ;
	wire _w8051_ ;
	wire _w8052_ ;
	wire _w8053_ ;
	wire _w8054_ ;
	wire _w8055_ ;
	wire _w8056_ ;
	wire _w8057_ ;
	wire _w8058_ ;
	wire _w8059_ ;
	wire _w8060_ ;
	wire _w8061_ ;
	wire _w8062_ ;
	wire _w8063_ ;
	wire _w8064_ ;
	wire _w8065_ ;
	wire _w8066_ ;
	wire _w8067_ ;
	wire _w8068_ ;
	wire _w8069_ ;
	wire _w8070_ ;
	wire _w8071_ ;
	wire _w8072_ ;
	wire _w8073_ ;
	wire _w8074_ ;
	wire _w8075_ ;
	wire _w8076_ ;
	wire _w8077_ ;
	wire _w8078_ ;
	wire _w8079_ ;
	wire _w8080_ ;
	wire _w8081_ ;
	wire _w8082_ ;
	wire _w8083_ ;
	wire _w8084_ ;
	wire _w8085_ ;
	wire _w8086_ ;
	wire _w8087_ ;
	wire _w8088_ ;
	wire _w8089_ ;
	wire _w8090_ ;
	wire _w8091_ ;
	wire _w8092_ ;
	wire _w8093_ ;
	wire _w8094_ ;
	wire _w8095_ ;
	wire _w8096_ ;
	wire _w8097_ ;
	wire _w8098_ ;
	wire _w8099_ ;
	wire _w8100_ ;
	wire _w8101_ ;
	wire _w8102_ ;
	wire _w8103_ ;
	wire _w8104_ ;
	wire _w8105_ ;
	wire _w8106_ ;
	wire _w8107_ ;
	wire _w8108_ ;
	wire _w8109_ ;
	wire _w8110_ ;
	wire _w8111_ ;
	wire _w8112_ ;
	wire _w8113_ ;
	wire _w8114_ ;
	wire _w8115_ ;
	wire _w8116_ ;
	wire _w8117_ ;
	wire _w8118_ ;
	wire _w8119_ ;
	wire _w8120_ ;
	wire _w8121_ ;
	wire _w8122_ ;
	wire _w8123_ ;
	wire _w8124_ ;
	wire _w8125_ ;
	wire _w8126_ ;
	wire _w8127_ ;
	wire _w8128_ ;
	wire _w8129_ ;
	wire _w8130_ ;
	wire _w8131_ ;
	wire _w8132_ ;
	wire _w8133_ ;
	wire _w8134_ ;
	wire _w8135_ ;
	wire _w8136_ ;
	wire _w8137_ ;
	wire _w8138_ ;
	wire _w8139_ ;
	wire _w8140_ ;
	wire _w8141_ ;
	wire _w8142_ ;
	wire _w8143_ ;
	wire _w8144_ ;
	wire _w8145_ ;
	wire _w8146_ ;
	wire _w8147_ ;
	wire _w8148_ ;
	wire _w8149_ ;
	wire _w8150_ ;
	wire _w8151_ ;
	wire _w8152_ ;
	wire _w8153_ ;
	wire _w8154_ ;
	wire _w8155_ ;
	wire _w8156_ ;
	wire _w8157_ ;
	wire _w8158_ ;
	wire _w8159_ ;
	wire _w8160_ ;
	wire _w8161_ ;
	wire _w8162_ ;
	wire _w8163_ ;
	wire _w8164_ ;
	wire _w8165_ ;
	wire _w8166_ ;
	wire _w8167_ ;
	wire _w8168_ ;
	wire _w8169_ ;
	wire _w8170_ ;
	wire _w8171_ ;
	wire _w8172_ ;
	wire _w8173_ ;
	wire _w8174_ ;
	wire _w8175_ ;
	wire _w8176_ ;
	wire _w8177_ ;
	wire _w8178_ ;
	wire _w8179_ ;
	wire _w8180_ ;
	wire _w8181_ ;
	wire _w8182_ ;
	wire _w8183_ ;
	wire _w8184_ ;
	wire _w8185_ ;
	wire _w8186_ ;
	wire _w8187_ ;
	wire _w8188_ ;
	wire _w8189_ ;
	wire _w8190_ ;
	wire _w8191_ ;
	wire _w8192_ ;
	wire _w8193_ ;
	wire _w8194_ ;
	wire _w8195_ ;
	wire _w8196_ ;
	wire _w8197_ ;
	wire _w8198_ ;
	wire _w8199_ ;
	wire _w8200_ ;
	wire _w8201_ ;
	wire _w8202_ ;
	wire _w8203_ ;
	wire _w8204_ ;
	wire _w8205_ ;
	wire _w8206_ ;
	wire _w8207_ ;
	wire _w8208_ ;
	wire _w8209_ ;
	wire _w8210_ ;
	wire _w8211_ ;
	wire _w8212_ ;
	wire _w8213_ ;
	wire _w8214_ ;
	wire _w8215_ ;
	wire _w8216_ ;
	wire _w8217_ ;
	wire _w8218_ ;
	wire _w8219_ ;
	wire _w8220_ ;
	wire _w8221_ ;
	wire _w8222_ ;
	wire _w8223_ ;
	wire _w8224_ ;
	wire _w8225_ ;
	wire _w8226_ ;
	wire _w8227_ ;
	wire _w8228_ ;
	wire _w8229_ ;
	wire _w8230_ ;
	wire _w8231_ ;
	wire _w8232_ ;
	wire _w8233_ ;
	wire _w8234_ ;
	wire _w8235_ ;
	wire _w8236_ ;
	wire _w8237_ ;
	wire _w8238_ ;
	wire _w8239_ ;
	wire _w8240_ ;
	wire _w8241_ ;
	wire _w8242_ ;
	wire _w8243_ ;
	wire _w8244_ ;
	wire _w8245_ ;
	wire _w8246_ ;
	wire _w8247_ ;
	wire _w8248_ ;
	wire _w8249_ ;
	wire _w8250_ ;
	wire _w8251_ ;
	wire _w8252_ ;
	wire _w8253_ ;
	wire _w8254_ ;
	wire _w8255_ ;
	wire _w8256_ ;
	wire _w8257_ ;
	wire _w8258_ ;
	wire _w8259_ ;
	wire _w8260_ ;
	wire _w8261_ ;
	wire _w8262_ ;
	wire _w8263_ ;
	wire _w8264_ ;
	wire _w8265_ ;
	wire _w8266_ ;
	wire _w8267_ ;
	wire _w8268_ ;
	wire _w8269_ ;
	wire _w8270_ ;
	wire _w8271_ ;
	wire _w8272_ ;
	wire _w8273_ ;
	wire _w8274_ ;
	wire _w8275_ ;
	wire _w8276_ ;
	wire _w8277_ ;
	wire _w8278_ ;
	wire _w8279_ ;
	wire _w8280_ ;
	wire _w8281_ ;
	wire _w8282_ ;
	wire _w8283_ ;
	wire _w8284_ ;
	wire _w8285_ ;
	wire _w8286_ ;
	wire _w8287_ ;
	wire _w8288_ ;
	wire _w8289_ ;
	wire _w8290_ ;
	wire _w8291_ ;
	wire _w8292_ ;
	wire _w8293_ ;
	wire _w8294_ ;
	wire _w8295_ ;
	wire _w8296_ ;
	wire _w8297_ ;
	wire _w8298_ ;
	wire _w8299_ ;
	wire _w8300_ ;
	wire _w8301_ ;
	wire _w8302_ ;
	wire _w8303_ ;
	wire _w8304_ ;
	wire _w8305_ ;
	wire _w8306_ ;
	wire _w8307_ ;
	wire _w8308_ ;
	wire _w8309_ ;
	wire _w8310_ ;
	wire _w8311_ ;
	wire _w8312_ ;
	wire _w8313_ ;
	wire _w8314_ ;
	wire _w8315_ ;
	wire _w8316_ ;
	wire _w8317_ ;
	wire _w8318_ ;
	wire _w8319_ ;
	wire _w8320_ ;
	wire _w8321_ ;
	wire _w8322_ ;
	wire _w8323_ ;
	wire _w8324_ ;
	wire _w8325_ ;
	wire _w8326_ ;
	wire _w8327_ ;
	wire _w8328_ ;
	wire _w8329_ ;
	wire _w8330_ ;
	wire _w8331_ ;
	wire _w8332_ ;
	wire _w8333_ ;
	wire _w8334_ ;
	wire _w8335_ ;
	wire _w8336_ ;
	wire _w8337_ ;
	wire _w8338_ ;
	wire _w8339_ ;
	wire _w8340_ ;
	wire _w8341_ ;
	wire _w8342_ ;
	wire _w8343_ ;
	wire _w8344_ ;
	wire _w8345_ ;
	wire _w8346_ ;
	wire _w8347_ ;
	wire _w8348_ ;
	wire _w8349_ ;
	wire _w8350_ ;
	wire _w8351_ ;
	wire _w8352_ ;
	wire _w8353_ ;
	wire _w8354_ ;
	wire _w8355_ ;
	wire _w8356_ ;
	wire _w8357_ ;
	wire _w8358_ ;
	wire _w8359_ ;
	wire _w8360_ ;
	wire _w8361_ ;
	wire _w8362_ ;
	wire _w8363_ ;
	wire _w8364_ ;
	wire _w8365_ ;
	wire _w8366_ ;
	wire _w8367_ ;
	wire _w8368_ ;
	wire _w8369_ ;
	wire _w8370_ ;
	wire _w8371_ ;
	wire _w8372_ ;
	wire _w8373_ ;
	wire _w8374_ ;
	wire _w8375_ ;
	wire _w8376_ ;
	wire _w8377_ ;
	wire _w8378_ ;
	wire _w8379_ ;
	wire _w8380_ ;
	wire _w8381_ ;
	wire _w8382_ ;
	wire _w8383_ ;
	wire _w8384_ ;
	wire _w8385_ ;
	wire _w8386_ ;
	wire _w8387_ ;
	wire _w8388_ ;
	wire _w8389_ ;
	wire _w8390_ ;
	wire _w8391_ ;
	wire _w8392_ ;
	wire _w8393_ ;
	wire _w8394_ ;
	wire _w8395_ ;
	wire _w8396_ ;
	wire _w8397_ ;
	wire _w8398_ ;
	wire _w8399_ ;
	wire _w8400_ ;
	wire _w8401_ ;
	wire _w8402_ ;
	wire _w8403_ ;
	wire _w8404_ ;
	wire _w8405_ ;
	wire _w8406_ ;
	wire _w8407_ ;
	wire _w8408_ ;
	wire _w8409_ ;
	wire _w8410_ ;
	wire _w8411_ ;
	wire _w8412_ ;
	wire _w8413_ ;
	wire _w8414_ ;
	wire _w8415_ ;
	wire _w8416_ ;
	wire _w8417_ ;
	wire _w8418_ ;
	wire _w8419_ ;
	wire _w8420_ ;
	wire _w8421_ ;
	wire _w8422_ ;
	wire _w8423_ ;
	wire _w8424_ ;
	wire _w8425_ ;
	wire _w8426_ ;
	wire _w8427_ ;
	wire _w8428_ ;
	wire _w8429_ ;
	wire _w8430_ ;
	wire _w8431_ ;
	wire _w8432_ ;
	wire _w8433_ ;
	wire _w8434_ ;
	wire _w8435_ ;
	wire _w8436_ ;
	wire _w8437_ ;
	wire _w8438_ ;
	wire _w8439_ ;
	wire _w8440_ ;
	wire _w8441_ ;
	wire _w8442_ ;
	wire _w8443_ ;
	wire _w8444_ ;
	wire _w8445_ ;
	wire _w8446_ ;
	wire _w8447_ ;
	wire _w8448_ ;
	wire _w8449_ ;
	wire _w8450_ ;
	wire _w8451_ ;
	wire _w8452_ ;
	wire _w8453_ ;
	wire _w8454_ ;
	wire _w8455_ ;
	wire _w8456_ ;
	wire _w8457_ ;
	wire _w8458_ ;
	wire _w8459_ ;
	wire _w8460_ ;
	wire _w8461_ ;
	wire _w8462_ ;
	wire _w8463_ ;
	wire _w8464_ ;
	wire _w8465_ ;
	wire _w8466_ ;
	wire _w8467_ ;
	wire _w8468_ ;
	wire _w8469_ ;
	wire _w8470_ ;
	wire _w8471_ ;
	wire _w8472_ ;
	wire _w8473_ ;
	wire _w8474_ ;
	wire _w8475_ ;
	wire _w8476_ ;
	wire _w8477_ ;
	wire _w8478_ ;
	wire _w8479_ ;
	wire _w8480_ ;
	wire _w8481_ ;
	wire _w8482_ ;
	wire _w8483_ ;
	wire _w8484_ ;
	wire _w8485_ ;
	wire _w8486_ ;
	wire _w8487_ ;
	wire _w8488_ ;
	wire _w8489_ ;
	wire _w8490_ ;
	wire _w8491_ ;
	wire _w8492_ ;
	wire _w8493_ ;
	wire _w8494_ ;
	wire _w8495_ ;
	wire _w8496_ ;
	wire _w8497_ ;
	wire _w8498_ ;
	wire _w8499_ ;
	wire _w8500_ ;
	wire _w8501_ ;
	wire _w8502_ ;
	wire _w8503_ ;
	wire _w8504_ ;
	wire _w8505_ ;
	wire _w8506_ ;
	wire _w8507_ ;
	wire _w8508_ ;
	wire _w8509_ ;
	wire _w8510_ ;
	wire _w8511_ ;
	wire _w8512_ ;
	wire _w8513_ ;
	wire _w8514_ ;
	wire _w8515_ ;
	wire _w8516_ ;
	wire _w8517_ ;
	wire _w8518_ ;
	wire _w8519_ ;
	wire _w8520_ ;
	wire _w8521_ ;
	wire _w8522_ ;
	wire _w8523_ ;
	wire _w8524_ ;
	wire _w8525_ ;
	wire _w8526_ ;
	wire _w8527_ ;
	wire _w8528_ ;
	wire _w8529_ ;
	wire _w8530_ ;
	wire _w8531_ ;
	wire _w8532_ ;
	wire _w8533_ ;
	wire _w8534_ ;
	wire _w8535_ ;
	wire _w8536_ ;
	wire _w8537_ ;
	wire _w8538_ ;
	wire _w8539_ ;
	wire _w8540_ ;
	wire _w8541_ ;
	wire _w8542_ ;
	wire _w8543_ ;
	wire _w8544_ ;
	wire _w8545_ ;
	wire _w8546_ ;
	wire _w8547_ ;
	wire _w8548_ ;
	wire _w8549_ ;
	wire _w8550_ ;
	wire _w8551_ ;
	wire _w8552_ ;
	wire _w8553_ ;
	wire _w8554_ ;
	wire _w8555_ ;
	wire _w8556_ ;
	wire _w8557_ ;
	wire _w8558_ ;
	wire _w8559_ ;
	wire _w8560_ ;
	wire _w8561_ ;
	wire _w8562_ ;
	wire _w8563_ ;
	wire _w8564_ ;
	wire _w8565_ ;
	wire _w8566_ ;
	wire _w8567_ ;
	wire _w8568_ ;
	wire _w8569_ ;
	wire _w8570_ ;
	wire _w8571_ ;
	wire _w8572_ ;
	wire _w8573_ ;
	wire _w8574_ ;
	wire _w8575_ ;
	wire _w8576_ ;
	wire _w8577_ ;
	wire _w8578_ ;
	wire _w8579_ ;
	wire _w8580_ ;
	wire _w8581_ ;
	wire _w8582_ ;
	wire _w8583_ ;
	wire _w8584_ ;
	wire _w8585_ ;
	wire _w8586_ ;
	wire _w8587_ ;
	wire _w8588_ ;
	wire _w8589_ ;
	wire _w8590_ ;
	wire _w8591_ ;
	wire _w8592_ ;
	wire _w8593_ ;
	wire _w8594_ ;
	wire _w8595_ ;
	wire _w8596_ ;
	wire _w8597_ ;
	wire _w8598_ ;
	wire _w8599_ ;
	wire _w8600_ ;
	wire _w8601_ ;
	wire _w8602_ ;
	wire _w8603_ ;
	wire _w8604_ ;
	wire _w8605_ ;
	wire _w8606_ ;
	wire _w8607_ ;
	wire _w8608_ ;
	wire _w8609_ ;
	wire _w8610_ ;
	wire _w8611_ ;
	wire _w8612_ ;
	wire _w8613_ ;
	wire _w8614_ ;
	wire _w8615_ ;
	wire _w8616_ ;
	wire _w8617_ ;
	wire _w8618_ ;
	wire _w8619_ ;
	wire _w8620_ ;
	wire _w8621_ ;
	wire _w8622_ ;
	wire _w8623_ ;
	wire _w8624_ ;
	wire _w8625_ ;
	wire _w8626_ ;
	wire _w8627_ ;
	wire _w8628_ ;
	wire _w8629_ ;
	wire _w8630_ ;
	wire _w8631_ ;
	wire _w8632_ ;
	wire _w8633_ ;
	wire _w8634_ ;
	wire _w8635_ ;
	wire _w8636_ ;
	wire _w8637_ ;
	wire _w8638_ ;
	wire _w8639_ ;
	wire _w8640_ ;
	wire _w8641_ ;
	wire _w8642_ ;
	wire _w8643_ ;
	wire _w8644_ ;
	wire _w8645_ ;
	wire _w8646_ ;
	wire _w8647_ ;
	wire _w8648_ ;
	wire _w8649_ ;
	wire _w8650_ ;
	wire _w8651_ ;
	wire _w8652_ ;
	wire _w8653_ ;
	wire _w8654_ ;
	wire _w8655_ ;
	wire _w8656_ ;
	wire _w8657_ ;
	wire _w8658_ ;
	wire _w8659_ ;
	wire _w8660_ ;
	wire _w8661_ ;
	wire _w8662_ ;
	wire _w8663_ ;
	wire _w8664_ ;
	wire _w8665_ ;
	wire _w8666_ ;
	wire _w8667_ ;
	wire _w8668_ ;
	wire _w8669_ ;
	wire _w8670_ ;
	wire _w8671_ ;
	wire _w8672_ ;
	wire _w8673_ ;
	wire _w8674_ ;
	wire _w8675_ ;
	wire _w8676_ ;
	wire _w8677_ ;
	wire _w8678_ ;
	wire _w8679_ ;
	wire _w8680_ ;
	wire _w8681_ ;
	wire _w8682_ ;
	wire _w8683_ ;
	wire _w8684_ ;
	wire _w8685_ ;
	wire _w8686_ ;
	wire _w8687_ ;
	wire _w8688_ ;
	wire _w8689_ ;
	wire _w8690_ ;
	wire _w8691_ ;
	wire _w8692_ ;
	wire _w8693_ ;
	wire _w8694_ ;
	wire _w8695_ ;
	wire _w8696_ ;
	wire _w8697_ ;
	wire _w8698_ ;
	wire _w8699_ ;
	wire _w8700_ ;
	wire _w8701_ ;
	wire _w8702_ ;
	wire _w8703_ ;
	wire _w8704_ ;
	wire _w8705_ ;
	wire _w8706_ ;
	wire _w8707_ ;
	wire _w8708_ ;
	wire _w8709_ ;
	wire _w8710_ ;
	wire _w8711_ ;
	wire _w8712_ ;
	wire _w8713_ ;
	wire _w8714_ ;
	wire _w8715_ ;
	wire _w8716_ ;
	wire _w8717_ ;
	wire _w8718_ ;
	wire _w8719_ ;
	wire _w8720_ ;
	wire _w8721_ ;
	wire _w8722_ ;
	wire _w8723_ ;
	wire _w8724_ ;
	wire _w8725_ ;
	wire _w8726_ ;
	wire _w8727_ ;
	wire _w8728_ ;
	wire _w8729_ ;
	wire _w8730_ ;
	wire _w8731_ ;
	wire _w8732_ ;
	wire _w8733_ ;
	wire _w8734_ ;
	wire _w8735_ ;
	wire _w8736_ ;
	wire _w8737_ ;
	wire _w8738_ ;
	wire _w8739_ ;
	wire _w8740_ ;
	wire _w8741_ ;
	wire _w8742_ ;
	wire _w8743_ ;
	wire _w8744_ ;
	wire _w8745_ ;
	wire _w8746_ ;
	wire _w8747_ ;
	wire _w8748_ ;
	wire _w8749_ ;
	wire _w8750_ ;
	wire _w8751_ ;
	wire _w8752_ ;
	wire _w8753_ ;
	wire _w8754_ ;
	wire _w8755_ ;
	wire _w8756_ ;
	wire _w8757_ ;
	wire _w8758_ ;
	wire _w8759_ ;
	wire _w8760_ ;
	wire _w8761_ ;
	wire _w8762_ ;
	wire _w8763_ ;
	wire _w8764_ ;
	wire _w8765_ ;
	wire _w8766_ ;
	wire _w8767_ ;
	wire _w8768_ ;
	wire _w8769_ ;
	wire _w8770_ ;
	wire _w8771_ ;
	wire _w8772_ ;
	wire _w8773_ ;
	wire _w8774_ ;
	wire _w8775_ ;
	wire _w8776_ ;
	wire _w8777_ ;
	wire _w8778_ ;
	wire _w8779_ ;
	wire _w8780_ ;
	wire _w8781_ ;
	wire _w8782_ ;
	wire _w8783_ ;
	wire _w8784_ ;
	wire _w8785_ ;
	wire _w8786_ ;
	wire _w8787_ ;
	wire _w8788_ ;
	wire _w8789_ ;
	wire _w8790_ ;
	wire _w8791_ ;
	wire _w8792_ ;
	wire _w8793_ ;
	wire _w8794_ ;
	wire _w8795_ ;
	wire _w8796_ ;
	wire _w8797_ ;
	wire _w8798_ ;
	wire _w8799_ ;
	wire _w8800_ ;
	wire _w8801_ ;
	wire _w8802_ ;
	wire _w8803_ ;
	wire _w8804_ ;
	wire _w8805_ ;
	wire _w8806_ ;
	wire _w8807_ ;
	wire _w8808_ ;
	wire _w8809_ ;
	wire _w8810_ ;
	wire _w8811_ ;
	wire _w8812_ ;
	wire _w8813_ ;
	wire _w8814_ ;
	wire _w8815_ ;
	wire _w8816_ ;
	wire _w8817_ ;
	wire _w8818_ ;
	wire _w8819_ ;
	wire _w8820_ ;
	wire _w8821_ ;
	wire _w8822_ ;
	wire _w8823_ ;
	wire _w8824_ ;
	wire _w8825_ ;
	wire _w8826_ ;
	wire _w8827_ ;
	wire _w8828_ ;
	wire _w8829_ ;
	wire _w8830_ ;
	wire _w8831_ ;
	wire _w8832_ ;
	wire _w8833_ ;
	wire _w8834_ ;
	wire _w8835_ ;
	wire _w8836_ ;
	wire _w8837_ ;
	wire _w8838_ ;
	wire _w8839_ ;
	wire _w8840_ ;
	wire _w8841_ ;
	wire _w8842_ ;
	wire _w8843_ ;
	wire _w8844_ ;
	wire _w8845_ ;
	wire _w8846_ ;
	wire _w8847_ ;
	wire _w8848_ ;
	wire _w8849_ ;
	wire _w8850_ ;
	wire _w8851_ ;
	wire _w8852_ ;
	wire _w8853_ ;
	wire _w8854_ ;
	wire _w8855_ ;
	wire _w8856_ ;
	wire _w8857_ ;
	wire _w8858_ ;
	wire _w8859_ ;
	wire _w8860_ ;
	wire _w8861_ ;
	wire _w8862_ ;
	wire _w8863_ ;
	wire _w8864_ ;
	wire _w8865_ ;
	wire _w8866_ ;
	wire _w8867_ ;
	wire _w8868_ ;
	wire _w8869_ ;
	wire _w8870_ ;
	wire _w8871_ ;
	wire _w8872_ ;
	wire _w8873_ ;
	wire _w8874_ ;
	wire _w8875_ ;
	wire _w8876_ ;
	wire _w8877_ ;
	wire _w8878_ ;
	wire _w8879_ ;
	wire _w8880_ ;
	wire _w8881_ ;
	wire _w8882_ ;
	wire _w8883_ ;
	wire _w8884_ ;
	wire _w8885_ ;
	wire _w8886_ ;
	wire _w8887_ ;
	wire _w8888_ ;
	wire _w8889_ ;
	wire _w8890_ ;
	wire _w8891_ ;
	wire _w8892_ ;
	wire _w8893_ ;
	wire _w8894_ ;
	wire _w8895_ ;
	wire _w8896_ ;
	wire _w8897_ ;
	wire _w8898_ ;
	wire _w8899_ ;
	wire _w8900_ ;
	wire _w8901_ ;
	wire _w8902_ ;
	wire _w8903_ ;
	wire _w8904_ ;
	wire _w8905_ ;
	wire _w8906_ ;
	wire _w8907_ ;
	wire _w8908_ ;
	wire _w8909_ ;
	wire _w8910_ ;
	wire _w8911_ ;
	wire _w8912_ ;
	wire _w8913_ ;
	wire _w8914_ ;
	wire _w8915_ ;
	wire _w8916_ ;
	wire _w8917_ ;
	wire _w8918_ ;
	wire _w8919_ ;
	wire _w8920_ ;
	wire _w8921_ ;
	wire _w8922_ ;
	wire _w8923_ ;
	wire _w8924_ ;
	wire _w8925_ ;
	wire _w8926_ ;
	wire _w8927_ ;
	wire _w8928_ ;
	wire _w8929_ ;
	wire _w8930_ ;
	wire _w8931_ ;
	wire _w8932_ ;
	wire _w8933_ ;
	wire _w8934_ ;
	wire _w8935_ ;
	wire _w8936_ ;
	wire _w8937_ ;
	wire _w8938_ ;
	wire _w8939_ ;
	wire _w8940_ ;
	wire _w8941_ ;
	wire _w8942_ ;
	wire _w8943_ ;
	wire _w8944_ ;
	wire _w8945_ ;
	wire _w8946_ ;
	wire _w8947_ ;
	wire _w8948_ ;
	wire _w8949_ ;
	wire _w8950_ ;
	wire _w8951_ ;
	wire _w8952_ ;
	wire _w8953_ ;
	wire _w8954_ ;
	wire _w8955_ ;
	wire _w8956_ ;
	wire _w8957_ ;
	wire _w8958_ ;
	wire _w8959_ ;
	wire _w8960_ ;
	wire _w8961_ ;
	wire _w8962_ ;
	wire _w8963_ ;
	wire _w8964_ ;
	wire _w8965_ ;
	wire _w8966_ ;
	wire _w8967_ ;
	wire _w8968_ ;
	wire _w8969_ ;
	wire _w8970_ ;
	wire _w8971_ ;
	wire _w8972_ ;
	wire _w8973_ ;
	wire _w8974_ ;
	wire _w8975_ ;
	wire _w8976_ ;
	wire _w8977_ ;
	wire _w8978_ ;
	wire _w8979_ ;
	wire _w8980_ ;
	wire _w8981_ ;
	wire _w8982_ ;
	wire _w8983_ ;
	wire _w8984_ ;
	wire _w8985_ ;
	wire _w8986_ ;
	wire _w8987_ ;
	wire _w8988_ ;
	wire _w8989_ ;
	wire _w8990_ ;
	wire _w8991_ ;
	wire _w8992_ ;
	wire _w8993_ ;
	wire _w8994_ ;
	wire _w8995_ ;
	wire _w8996_ ;
	wire _w8997_ ;
	wire _w8998_ ;
	wire _w8999_ ;
	wire _w9000_ ;
	wire _w9001_ ;
	wire _w9002_ ;
	wire _w9003_ ;
	wire _w9004_ ;
	wire _w9005_ ;
	wire _w9006_ ;
	wire _w9007_ ;
	wire _w9008_ ;
	wire _w9009_ ;
	wire _w9010_ ;
	wire _w9011_ ;
	wire _w9012_ ;
	wire _w9013_ ;
	wire _w9014_ ;
	wire _w9015_ ;
	wire _w9016_ ;
	wire _w9017_ ;
	wire _w9018_ ;
	wire _w9019_ ;
	wire _w9020_ ;
	wire _w9021_ ;
	wire _w9022_ ;
	wire _w9023_ ;
	wire _w9024_ ;
	wire _w9025_ ;
	wire _w9026_ ;
	wire _w9027_ ;
	wire _w9028_ ;
	wire _w9029_ ;
	wire _w9030_ ;
	wire _w9031_ ;
	wire _w9032_ ;
	wire _w9033_ ;
	wire _w9034_ ;
	wire _w9035_ ;
	wire _w9036_ ;
	wire _w9037_ ;
	wire _w9038_ ;
	wire _w9039_ ;
	wire _w9040_ ;
	wire _w9041_ ;
	wire _w9042_ ;
	wire _w9043_ ;
	wire _w9044_ ;
	wire _w9045_ ;
	wire _w9046_ ;
	wire _w9047_ ;
	wire _w9048_ ;
	wire _w9049_ ;
	wire _w9050_ ;
	wire _w9051_ ;
	wire _w9052_ ;
	wire _w9053_ ;
	wire _w9054_ ;
	wire _w9055_ ;
	wire _w9056_ ;
	wire _w9057_ ;
	wire _w9058_ ;
	wire _w9059_ ;
	wire _w9060_ ;
	wire _w9061_ ;
	wire _w9062_ ;
	wire _w9063_ ;
	wire _w9064_ ;
	wire _w9065_ ;
	wire _w9066_ ;
	wire _w9067_ ;
	wire _w9068_ ;
	wire _w9069_ ;
	wire _w9070_ ;
	wire _w9071_ ;
	wire _w9072_ ;
	wire _w9073_ ;
	wire _w9074_ ;
	wire _w9075_ ;
	wire _w9076_ ;
	wire _w9077_ ;
	wire _w9078_ ;
	wire _w9079_ ;
	wire _w9080_ ;
	wire _w9081_ ;
	wire _w9082_ ;
	wire _w9083_ ;
	wire _w9084_ ;
	wire _w9085_ ;
	wire _w9086_ ;
	wire _w9087_ ;
	wire _w9088_ ;
	wire _w9089_ ;
	wire _w9090_ ;
	wire _w9091_ ;
	wire _w9092_ ;
	wire _w9093_ ;
	wire _w9094_ ;
	wire _w9095_ ;
	wire _w9096_ ;
	wire _w9097_ ;
	wire _w9098_ ;
	wire _w9099_ ;
	wire _w9100_ ;
	wire _w9101_ ;
	wire _w9102_ ;
	wire _w9103_ ;
	wire _w9104_ ;
	wire _w9105_ ;
	wire _w9106_ ;
	wire _w9107_ ;
	wire _w9108_ ;
	wire _w9109_ ;
	wire _w9110_ ;
	wire _w9111_ ;
	wire _w9112_ ;
	wire _w9113_ ;
	wire _w9114_ ;
	wire _w9115_ ;
	wire _w9116_ ;
	wire _w9117_ ;
	wire _w9118_ ;
	wire _w9119_ ;
	wire _w9120_ ;
	wire _w9121_ ;
	wire _w9122_ ;
	wire _w9123_ ;
	wire _w9124_ ;
	wire _w9125_ ;
	wire _w9126_ ;
	wire _w9127_ ;
	wire _w9128_ ;
	wire _w9129_ ;
	wire _w9130_ ;
	wire _w9131_ ;
	wire _w9132_ ;
	wire _w9133_ ;
	wire _w9134_ ;
	wire _w9135_ ;
	wire _w9136_ ;
	wire _w9137_ ;
	wire _w9138_ ;
	wire _w9139_ ;
	wire _w9140_ ;
	wire _w9141_ ;
	wire _w9142_ ;
	wire _w9143_ ;
	wire _w9144_ ;
	wire _w9145_ ;
	wire _w9146_ ;
	wire _w9147_ ;
	wire _w9148_ ;
	wire _w9149_ ;
	wire _w9150_ ;
	wire _w9151_ ;
	wire _w9152_ ;
	wire _w9153_ ;
	wire _w9154_ ;
	wire _w9155_ ;
	wire _w9156_ ;
	wire _w9157_ ;
	wire _w9158_ ;
	wire _w9159_ ;
	wire _w9160_ ;
	wire _w9161_ ;
	wire _w9162_ ;
	wire _w9163_ ;
	wire _w9164_ ;
	wire _w9165_ ;
	wire _w9166_ ;
	wire _w9167_ ;
	wire _w9168_ ;
	wire _w9169_ ;
	wire _w9170_ ;
	wire _w9171_ ;
	wire _w9172_ ;
	wire _w9173_ ;
	wire _w9174_ ;
	wire _w9175_ ;
	wire _w9176_ ;
	wire _w9177_ ;
	wire _w9178_ ;
	wire _w9179_ ;
	wire _w9180_ ;
	wire _w9181_ ;
	wire _w9182_ ;
	wire _w9183_ ;
	wire _w9184_ ;
	wire _w9185_ ;
	wire _w9186_ ;
	wire _w9187_ ;
	wire _w9188_ ;
	wire _w9189_ ;
	wire _w9190_ ;
	wire _w9191_ ;
	wire _w9192_ ;
	wire _w9193_ ;
	wire _w9194_ ;
	wire _w9195_ ;
	wire _w9196_ ;
	wire _w9197_ ;
	wire _w9198_ ;
	wire _w9199_ ;
	wire _w9200_ ;
	wire _w9201_ ;
	wire _w9202_ ;
	wire _w9203_ ;
	wire _w9204_ ;
	wire _w9205_ ;
	wire _w9206_ ;
	wire _w9207_ ;
	wire _w9208_ ;
	wire _w9209_ ;
	wire _w9210_ ;
	wire _w9211_ ;
	wire _w9212_ ;
	wire _w9213_ ;
	wire _w9214_ ;
	wire _w9215_ ;
	wire _w9216_ ;
	wire _w9217_ ;
	wire _w9218_ ;
	wire _w9219_ ;
	wire _w9220_ ;
	wire _w9221_ ;
	wire _w9222_ ;
	wire _w9223_ ;
	wire _w9224_ ;
	wire _w9225_ ;
	wire _w9226_ ;
	wire _w9227_ ;
	wire _w9228_ ;
	wire _w9229_ ;
	wire _w9230_ ;
	wire _w9231_ ;
	wire _w9232_ ;
	wire _w9233_ ;
	wire _w9234_ ;
	wire _w9235_ ;
	wire _w9236_ ;
	wire _w9237_ ;
	wire _w9238_ ;
	wire _w9239_ ;
	wire _w9240_ ;
	wire _w9241_ ;
	wire _w9242_ ;
	wire _w9243_ ;
	wire _w9244_ ;
	wire _w9245_ ;
	wire _w9246_ ;
	wire _w9247_ ;
	wire _w9248_ ;
	wire _w9249_ ;
	wire _w9250_ ;
	wire _w9251_ ;
	wire _w9252_ ;
	wire _w9253_ ;
	wire _w9254_ ;
	wire _w9255_ ;
	wire _w9256_ ;
	wire _w9257_ ;
	wire _w9258_ ;
	wire _w9259_ ;
	wire _w9260_ ;
	wire _w9261_ ;
	wire _w9262_ ;
	wire _w9263_ ;
	wire _w9264_ ;
	wire _w9265_ ;
	wire _w9266_ ;
	wire _w9267_ ;
	wire _w9268_ ;
	wire _w9269_ ;
	wire _w9270_ ;
	wire _w9271_ ;
	wire _w9272_ ;
	wire _w9273_ ;
	wire _w9274_ ;
	wire _w9275_ ;
	wire _w9276_ ;
	wire _w9277_ ;
	wire _w9278_ ;
	wire _w9279_ ;
	wire _w9280_ ;
	wire _w9281_ ;
	wire _w9282_ ;
	wire _w9283_ ;
	wire _w9284_ ;
	wire _w9285_ ;
	wire _w9286_ ;
	wire _w9287_ ;
	wire _w9288_ ;
	wire _w9289_ ;
	wire _w9290_ ;
	wire _w9291_ ;
	wire _w9292_ ;
	wire _w9293_ ;
	wire _w9294_ ;
	wire _w9295_ ;
	wire _w9296_ ;
	wire _w9297_ ;
	wire _w9298_ ;
	wire _w9299_ ;
	wire _w9300_ ;
	wire _w9301_ ;
	wire _w9302_ ;
	wire _w9303_ ;
	wire _w9304_ ;
	wire _w9305_ ;
	wire _w9306_ ;
	wire _w9307_ ;
	wire _w9308_ ;
	wire _w9309_ ;
	wire _w9310_ ;
	wire _w9311_ ;
	wire _w9312_ ;
	wire _w9313_ ;
	wire _w9314_ ;
	wire _w9315_ ;
	wire _w9316_ ;
	wire _w9317_ ;
	wire _w9318_ ;
	wire _w9319_ ;
	wire _w9320_ ;
	wire _w9321_ ;
	wire _w9322_ ;
	wire _w9323_ ;
	wire _w9324_ ;
	wire _w9325_ ;
	wire _w9326_ ;
	wire _w9327_ ;
	wire _w9328_ ;
	wire _w9329_ ;
	wire _w9330_ ;
	wire _w9331_ ;
	wire _w9332_ ;
	wire _w9333_ ;
	wire _w9334_ ;
	wire _w9335_ ;
	wire _w9336_ ;
	wire _w9337_ ;
	wire _w9338_ ;
	wire _w9339_ ;
	wire _w9340_ ;
	wire _w9341_ ;
	wire _w9342_ ;
	wire _w9343_ ;
	wire _w9344_ ;
	wire _w9345_ ;
	wire _w9346_ ;
	wire _w9347_ ;
	wire _w9348_ ;
	wire _w9349_ ;
	wire _w9350_ ;
	wire _w9351_ ;
	wire _w9352_ ;
	wire _w9353_ ;
	wire _w9354_ ;
	wire _w9355_ ;
	wire _w9356_ ;
	wire _w9357_ ;
	wire _w9358_ ;
	wire _w9359_ ;
	wire _w9360_ ;
	wire _w9361_ ;
	wire _w9362_ ;
	wire _w9363_ ;
	wire _w9364_ ;
	wire _w9365_ ;
	wire _w9366_ ;
	wire _w9367_ ;
	wire _w9368_ ;
	wire _w9369_ ;
	wire _w9370_ ;
	wire _w9371_ ;
	wire _w9372_ ;
	wire _w9373_ ;
	wire _w9374_ ;
	wire _w9375_ ;
	wire _w9376_ ;
	wire _w9377_ ;
	wire _w9378_ ;
	wire _w9379_ ;
	wire _w9380_ ;
	wire _w9381_ ;
	wire _w9382_ ;
	wire _w9383_ ;
	wire _w9384_ ;
	wire _w9385_ ;
	wire _w9386_ ;
	wire _w9387_ ;
	wire _w9388_ ;
	wire _w9389_ ;
	wire _w9390_ ;
	wire _w9391_ ;
	wire _w9392_ ;
	wire _w9393_ ;
	wire _w9394_ ;
	wire _w9395_ ;
	wire _w9396_ ;
	wire _w9397_ ;
	wire _w9398_ ;
	wire _w9399_ ;
	wire _w9400_ ;
	wire _w9401_ ;
	wire _w9402_ ;
	wire _w9403_ ;
	wire _w9404_ ;
	wire _w9405_ ;
	wire _w9406_ ;
	wire _w9407_ ;
	wire _w9408_ ;
	wire _w9409_ ;
	wire _w9410_ ;
	wire _w9411_ ;
	wire _w9412_ ;
	wire _w9413_ ;
	wire _w9414_ ;
	wire _w9415_ ;
	wire _w9416_ ;
	wire _w9417_ ;
	wire _w9418_ ;
	wire _w9419_ ;
	wire _w9420_ ;
	wire _w9421_ ;
	wire _w9422_ ;
	wire _w9423_ ;
	wire _w9424_ ;
	wire _w9425_ ;
	wire _w9426_ ;
	wire _w9427_ ;
	wire _w9428_ ;
	wire _w9429_ ;
	wire _w9430_ ;
	wire _w9431_ ;
	wire _w9432_ ;
	wire _w9433_ ;
	wire _w9434_ ;
	wire _w9435_ ;
	wire _w9436_ ;
	wire _w9437_ ;
	wire _w9438_ ;
	wire _w9439_ ;
	wire _w9440_ ;
	wire _w9441_ ;
	wire _w9442_ ;
	wire _w9443_ ;
	wire _w9444_ ;
	wire _w9445_ ;
	wire _w9446_ ;
	wire _w9447_ ;
	wire _w9448_ ;
	wire _w9449_ ;
	wire _w9450_ ;
	wire _w9451_ ;
	wire _w9452_ ;
	wire _w9453_ ;
	wire _w9454_ ;
	wire _w9455_ ;
	wire _w9456_ ;
	wire _w9457_ ;
	wire _w9458_ ;
	wire _w9459_ ;
	wire _w9460_ ;
	wire _w9461_ ;
	wire _w9462_ ;
	wire _w9463_ ;
	wire _w9464_ ;
	wire _w9465_ ;
	wire _w9466_ ;
	wire _w9467_ ;
	wire _w9468_ ;
	wire _w9469_ ;
	wire _w9470_ ;
	wire _w9471_ ;
	wire _w9472_ ;
	wire _w9473_ ;
	wire _w9474_ ;
	wire _w9475_ ;
	wire _w9476_ ;
	wire _w9477_ ;
	wire _w9478_ ;
	wire _w9479_ ;
	wire _w9480_ ;
	wire _w9481_ ;
	wire _w9482_ ;
	wire _w9483_ ;
	wire _w9484_ ;
	wire _w9485_ ;
	wire _w9486_ ;
	wire _w9487_ ;
	wire _w9488_ ;
	wire _w9489_ ;
	wire _w9490_ ;
	wire _w9491_ ;
	wire _w9492_ ;
	wire _w9493_ ;
	wire _w9494_ ;
	wire _w9495_ ;
	wire _w9496_ ;
	wire _w9497_ ;
	wire _w9498_ ;
	wire _w9499_ ;
	wire _w9500_ ;
	wire _w9501_ ;
	wire _w9502_ ;
	wire _w9503_ ;
	wire _w9504_ ;
	wire _w9505_ ;
	wire _w9506_ ;
	wire _w9507_ ;
	wire _w9508_ ;
	wire _w9509_ ;
	wire _w9510_ ;
	wire _w9511_ ;
	wire _w9512_ ;
	wire _w9513_ ;
	wire _w9514_ ;
	wire _w9515_ ;
	wire _w9516_ ;
	wire _w9517_ ;
	wire _w9518_ ;
	wire _w9519_ ;
	wire _w9520_ ;
	wire _w9521_ ;
	wire _w9522_ ;
	wire _w9523_ ;
	wire _w9524_ ;
	wire _w9525_ ;
	wire _w9526_ ;
	wire _w9527_ ;
	wire _w9528_ ;
	wire _w9529_ ;
	wire _w9530_ ;
	wire _w9531_ ;
	wire _w9532_ ;
	wire _w9533_ ;
	wire _w9534_ ;
	wire _w9535_ ;
	wire _w9536_ ;
	wire _w9537_ ;
	wire _w9538_ ;
	wire _w9539_ ;
	wire _w9540_ ;
	wire _w9541_ ;
	wire _w9542_ ;
	wire _w9543_ ;
	wire _w9544_ ;
	wire _w9545_ ;
	wire _w9546_ ;
	wire _w9547_ ;
	wire _w9548_ ;
	wire _w9549_ ;
	wire _w9550_ ;
	wire _w9551_ ;
	wire _w9552_ ;
	wire _w9553_ ;
	wire _w9554_ ;
	wire _w9555_ ;
	wire _w9556_ ;
	wire _w9557_ ;
	wire _w9558_ ;
	wire _w9559_ ;
	wire _w9560_ ;
	wire _w9561_ ;
	wire _w9562_ ;
	wire _w9563_ ;
	wire _w9564_ ;
	wire _w9565_ ;
	wire _w9566_ ;
	wire _w9567_ ;
	wire _w9568_ ;
	wire _w9569_ ;
	wire _w9570_ ;
	wire _w9571_ ;
	wire _w9572_ ;
	wire _w9573_ ;
	wire _w9574_ ;
	wire _w9575_ ;
	wire _w9576_ ;
	wire _w9577_ ;
	wire _w9578_ ;
	wire _w9579_ ;
	wire _w9580_ ;
	wire _w9581_ ;
	wire _w9582_ ;
	wire _w9583_ ;
	wire _w9584_ ;
	wire _w9585_ ;
	wire _w9586_ ;
	wire _w9587_ ;
	wire _w9588_ ;
	wire _w9589_ ;
	wire _w9590_ ;
	wire _w9591_ ;
	wire _w9592_ ;
	wire _w9593_ ;
	wire _w9594_ ;
	wire _w9595_ ;
	wire _w9596_ ;
	wire _w9597_ ;
	wire _w9598_ ;
	wire _w9599_ ;
	wire _w9600_ ;
	wire _w9601_ ;
	wire _w9602_ ;
	wire _w9603_ ;
	wire _w9604_ ;
	wire _w9605_ ;
	wire _w9606_ ;
	wire _w9607_ ;
	wire _w9608_ ;
	wire _w9609_ ;
	wire _w9610_ ;
	wire _w9611_ ;
	wire _w9612_ ;
	wire _w9613_ ;
	wire _w9614_ ;
	wire _w9615_ ;
	wire _w9616_ ;
	wire _w9617_ ;
	wire _w9618_ ;
	wire _w9619_ ;
	wire _w9620_ ;
	wire _w9621_ ;
	wire _w9622_ ;
	wire _w9623_ ;
	wire _w9624_ ;
	wire _w9625_ ;
	wire _w9626_ ;
	wire _w9627_ ;
	wire _w9628_ ;
	wire _w9629_ ;
	wire _w9630_ ;
	wire _w9631_ ;
	wire _w9632_ ;
	wire _w9633_ ;
	wire _w9634_ ;
	wire _w9635_ ;
	wire _w9636_ ;
	wire _w9637_ ;
	wire _w9638_ ;
	wire _w9639_ ;
	wire _w9640_ ;
	wire _w9641_ ;
	wire _w9642_ ;
	wire _w9643_ ;
	wire _w9644_ ;
	wire _w9645_ ;
	wire _w9646_ ;
	wire _w9647_ ;
	wire _w9648_ ;
	wire _w9649_ ;
	wire _w9650_ ;
	wire _w9651_ ;
	wire _w9652_ ;
	wire _w9653_ ;
	wire _w9654_ ;
	wire _w9655_ ;
	wire _w9656_ ;
	wire _w9657_ ;
	wire _w9658_ ;
	wire _w9659_ ;
	wire _w9660_ ;
	wire _w9661_ ;
	wire _w9662_ ;
	wire _w9663_ ;
	wire _w9664_ ;
	wire _w9665_ ;
	wire _w9666_ ;
	wire _w9667_ ;
	wire _w9668_ ;
	wire _w9669_ ;
	wire _w9670_ ;
	wire _w9671_ ;
	wire _w9672_ ;
	wire _w9673_ ;
	wire _w9674_ ;
	wire _w9675_ ;
	wire _w9676_ ;
	wire _w9677_ ;
	wire _w9678_ ;
	wire _w9679_ ;
	wire _w9680_ ;
	wire _w9681_ ;
	wire _w9682_ ;
	wire _w9683_ ;
	wire _w9684_ ;
	wire _w9685_ ;
	wire _w9686_ ;
	wire _w9687_ ;
	wire _w9688_ ;
	wire _w9689_ ;
	wire _w9690_ ;
	wire _w9691_ ;
	wire _w9692_ ;
	wire _w9693_ ;
	wire _w9694_ ;
	wire _w9695_ ;
	wire _w9696_ ;
	wire _w9697_ ;
	wire _w9698_ ;
	wire _w9699_ ;
	wire _w9700_ ;
	wire _w9701_ ;
	wire _w9702_ ;
	wire _w9703_ ;
	wire _w9704_ ;
	wire _w9705_ ;
	wire _w9706_ ;
	wire _w9707_ ;
	wire _w9708_ ;
	wire _w9709_ ;
	wire _w9710_ ;
	wire _w9711_ ;
	wire _w9712_ ;
	wire _w9713_ ;
	wire _w9714_ ;
	wire _w9715_ ;
	wire _w9716_ ;
	wire _w9717_ ;
	wire _w9718_ ;
	wire _w9719_ ;
	wire _w9720_ ;
	wire _w9721_ ;
	wire _w9722_ ;
	wire _w9723_ ;
	wire _w9724_ ;
	wire _w9725_ ;
	wire _w9726_ ;
	wire _w9727_ ;
	wire _w9728_ ;
	wire _w9729_ ;
	wire _w9730_ ;
	wire _w9731_ ;
	wire _w9732_ ;
	wire _w9733_ ;
	wire _w9734_ ;
	wire _w9735_ ;
	wire _w9736_ ;
	wire _w9737_ ;
	wire _w9738_ ;
	wire _w9739_ ;
	wire _w9740_ ;
	wire _w9741_ ;
	wire _w9742_ ;
	wire _w9743_ ;
	wire _w9744_ ;
	wire _w9745_ ;
	wire _w9746_ ;
	wire _w9747_ ;
	wire _w9748_ ;
	wire _w9749_ ;
	wire _w9750_ ;
	wire _w9751_ ;
	wire _w9752_ ;
	wire _w9753_ ;
	wire _w9754_ ;
	wire _w9755_ ;
	wire _w9756_ ;
	wire _w9757_ ;
	wire _w9758_ ;
	wire _w9759_ ;
	wire _w9760_ ;
	wire _w9761_ ;
	wire _w9762_ ;
	wire _w9763_ ;
	wire _w9764_ ;
	wire _w9765_ ;
	wire _w9766_ ;
	wire _w9767_ ;
	wire _w9768_ ;
	wire _w9769_ ;
	wire _w9770_ ;
	wire _w9771_ ;
	wire _w9772_ ;
	wire _w9773_ ;
	wire _w9774_ ;
	wire _w9775_ ;
	wire _w9776_ ;
	wire _w9777_ ;
	wire _w9778_ ;
	wire _w9779_ ;
	wire _w9780_ ;
	wire _w9781_ ;
	wire _w9782_ ;
	wire _w9783_ ;
	wire _w9784_ ;
	wire _w9785_ ;
	wire _w9786_ ;
	wire _w9787_ ;
	wire _w9788_ ;
	wire _w9789_ ;
	wire _w9790_ ;
	wire _w9791_ ;
	wire _w9792_ ;
	wire _w9793_ ;
	wire _w9794_ ;
	wire _w9795_ ;
	wire _w9796_ ;
	wire _w9797_ ;
	wire _w9798_ ;
	wire _w9799_ ;
	wire _w9800_ ;
	wire _w9801_ ;
	wire _w9802_ ;
	wire _w9803_ ;
	wire _w9804_ ;
	wire _w9805_ ;
	wire _w9806_ ;
	wire _w9807_ ;
	wire _w9808_ ;
	wire _w9809_ ;
	wire _w9810_ ;
	wire _w9811_ ;
	wire _w9812_ ;
	wire _w9813_ ;
	wire _w9814_ ;
	wire _w9815_ ;
	wire _w9816_ ;
	wire _w9817_ ;
	wire _w9818_ ;
	wire _w9819_ ;
	wire _w9820_ ;
	wire _w9821_ ;
	wire _w9822_ ;
	wire _w9823_ ;
	wire _w9824_ ;
	wire _w9825_ ;
	wire _w9826_ ;
	wire _w9827_ ;
	wire _w9828_ ;
	wire _w9829_ ;
	wire _w9830_ ;
	wire _w9831_ ;
	wire _w9832_ ;
	wire _w9833_ ;
	wire _w9834_ ;
	wire _w9835_ ;
	wire _w9836_ ;
	wire _w9837_ ;
	wire _w9838_ ;
	wire _w9839_ ;
	wire _w9840_ ;
	wire _w9841_ ;
	wire _w9842_ ;
	wire _w9843_ ;
	wire _w9844_ ;
	wire _w9845_ ;
	wire _w9846_ ;
	wire _w9847_ ;
	wire _w9848_ ;
	wire _w9849_ ;
	wire _w9850_ ;
	wire _w9851_ ;
	wire _w9852_ ;
	wire _w9853_ ;
	wire _w9854_ ;
	wire _w9855_ ;
	wire _w9856_ ;
	wire _w9857_ ;
	wire _w9858_ ;
	wire _w9859_ ;
	wire _w9860_ ;
	wire _w9861_ ;
	wire _w9862_ ;
	wire _w9863_ ;
	wire _w9864_ ;
	wire _w9865_ ;
	wire _w9866_ ;
	wire _w9867_ ;
	wire _w9868_ ;
	wire _w9869_ ;
	wire _w9870_ ;
	wire _w9871_ ;
	wire _w9872_ ;
	wire _w9873_ ;
	wire _w9874_ ;
	wire _w9875_ ;
	wire _w9876_ ;
	wire _w9877_ ;
	wire _w9878_ ;
	wire _w9879_ ;
	wire _w9880_ ;
	wire _w9881_ ;
	wire _w9882_ ;
	wire _w9883_ ;
	wire _w9884_ ;
	wire _w9885_ ;
	wire _w9886_ ;
	wire _w9887_ ;
	wire _w9888_ ;
	wire _w9889_ ;
	wire _w9890_ ;
	wire _w9891_ ;
	wire _w9892_ ;
	wire _w9893_ ;
	wire _w9894_ ;
	wire _w9895_ ;
	wire _w9896_ ;
	wire _w9897_ ;
	wire _w9898_ ;
	wire _w9899_ ;
	wire _w9900_ ;
	wire _w9901_ ;
	wire _w9902_ ;
	wire _w9903_ ;
	wire _w9904_ ;
	wire _w9905_ ;
	wire _w9906_ ;
	wire _w9907_ ;
	wire _w9908_ ;
	wire _w9909_ ;
	wire _w9910_ ;
	wire _w9911_ ;
	wire _w9912_ ;
	wire _w9913_ ;
	wire _w9914_ ;
	wire _w9915_ ;
	wire _w9916_ ;
	wire _w9917_ ;
	wire _w9918_ ;
	wire _w9919_ ;
	wire _w9920_ ;
	wire _w9921_ ;
	wire _w9922_ ;
	wire _w9923_ ;
	wire _w9924_ ;
	wire _w9925_ ;
	wire _w9926_ ;
	wire _w9927_ ;
	wire _w9928_ ;
	wire _w9929_ ;
	wire _w9930_ ;
	wire _w9931_ ;
	wire _w9932_ ;
	wire _w9933_ ;
	wire _w9934_ ;
	wire _w9935_ ;
	wire _w9936_ ;
	wire _w9937_ ;
	wire _w9938_ ;
	wire _w9939_ ;
	wire _w9940_ ;
	wire _w9941_ ;
	wire _w9942_ ;
	wire _w9943_ ;
	wire _w9944_ ;
	wire _w9945_ ;
	wire _w9946_ ;
	wire _w9947_ ;
	wire _w9948_ ;
	wire _w9949_ ;
	wire _w9950_ ;
	wire _w9951_ ;
	wire _w9952_ ;
	wire _w9953_ ;
	wire _w9954_ ;
	wire _w9955_ ;
	wire _w9956_ ;
	wire _w9957_ ;
	wire _w9958_ ;
	wire _w9959_ ;
	wire _w9960_ ;
	wire _w9961_ ;
	wire _w9962_ ;
	wire _w9963_ ;
	wire _w9964_ ;
	wire _w9965_ ;
	wire _w9966_ ;
	wire _w9967_ ;
	wire _w9968_ ;
	wire _w9969_ ;
	wire _w9970_ ;
	wire _w9971_ ;
	wire _w9972_ ;
	wire _w9973_ ;
	wire _w9974_ ;
	wire _w9975_ ;
	wire _w9976_ ;
	wire _w9977_ ;
	wire _w9978_ ;
	wire _w9979_ ;
	wire _w9980_ ;
	wire _w9981_ ;
	wire _w9982_ ;
	wire _w9983_ ;
	wire _w9984_ ;
	wire _w9985_ ;
	wire _w9986_ ;
	wire _w9987_ ;
	wire _w9988_ ;
	wire _w9989_ ;
	wire _w9990_ ;
	wire _w9991_ ;
	wire _w9992_ ;
	wire _w9993_ ;
	wire _w9994_ ;
	wire _w9995_ ;
	wire _w9996_ ;
	wire _w9997_ ;
	wire _w9998_ ;
	wire _w9999_ ;
	wire _w10000_ ;
	wire _w10001_ ;
	wire _w10002_ ;
	wire _w10003_ ;
	wire _w10004_ ;
	wire _w10005_ ;
	wire _w10006_ ;
	wire _w10007_ ;
	wire _w10008_ ;
	wire _w10009_ ;
	wire _w10010_ ;
	wire _w10011_ ;
	wire _w10012_ ;
	wire _w10013_ ;
	wire _w10014_ ;
	wire _w10015_ ;
	wire _w10016_ ;
	wire _w10017_ ;
	wire _w10018_ ;
	wire _w10019_ ;
	wire _w10020_ ;
	wire _w10021_ ;
	wire _w10022_ ;
	wire _w10023_ ;
	wire _w10024_ ;
	wire _w10025_ ;
	wire _w10026_ ;
	wire _w10027_ ;
	wire _w10028_ ;
	wire _w10029_ ;
	wire _w10030_ ;
	wire _w10031_ ;
	wire _w10032_ ;
	wire _w10033_ ;
	wire _w10034_ ;
	wire _w10035_ ;
	wire _w10036_ ;
	wire _w10037_ ;
	wire _w10038_ ;
	wire _w10039_ ;
	wire _w10040_ ;
	wire _w10041_ ;
	wire _w10042_ ;
	wire _w10043_ ;
	wire _w10044_ ;
	wire _w10045_ ;
	wire _w10046_ ;
	wire _w10047_ ;
	wire _w10048_ ;
	wire _w10049_ ;
	wire _w10050_ ;
	wire _w10051_ ;
	wire _w10052_ ;
	wire _w10053_ ;
	wire _w10054_ ;
	wire _w10055_ ;
	wire _w10056_ ;
	wire _w10057_ ;
	wire _w10058_ ;
	wire _w10059_ ;
	wire _w10060_ ;
	wire _w10061_ ;
	wire _w10062_ ;
	wire _w10063_ ;
	wire _w10064_ ;
	wire _w10065_ ;
	wire _w10066_ ;
	wire _w10067_ ;
	wire _w10068_ ;
	wire _w10069_ ;
	wire _w10070_ ;
	wire _w10071_ ;
	wire _w10072_ ;
	wire _w10073_ ;
	wire _w10074_ ;
	wire _w10075_ ;
	wire _w10076_ ;
	wire _w10077_ ;
	wire _w10078_ ;
	wire _w10079_ ;
	wire _w10080_ ;
	wire _w10081_ ;
	wire _w10082_ ;
	wire _w10083_ ;
	wire _w10084_ ;
	wire _w10085_ ;
	wire _w10086_ ;
	wire _w10087_ ;
	wire _w10088_ ;
	wire _w10089_ ;
	wire _w10090_ ;
	wire _w10091_ ;
	wire _w10092_ ;
	wire _w10093_ ;
	wire _w10094_ ;
	wire _w10095_ ;
	wire _w10096_ ;
	wire _w10097_ ;
	wire _w10098_ ;
	wire _w10099_ ;
	wire _w10100_ ;
	wire _w10101_ ;
	wire _w10102_ ;
	wire _w10103_ ;
	wire _w10104_ ;
	wire _w10105_ ;
	wire _w10106_ ;
	wire _w10107_ ;
	wire _w10108_ ;
	wire _w10109_ ;
	wire _w10110_ ;
	wire _w10111_ ;
	wire _w10112_ ;
	wire _w10113_ ;
	wire _w10114_ ;
	wire _w10115_ ;
	wire _w10116_ ;
	wire _w10117_ ;
	wire _w10118_ ;
	wire _w10119_ ;
	wire _w10120_ ;
	wire _w10121_ ;
	wire _w10122_ ;
	wire _w10123_ ;
	wire _w10124_ ;
	wire _w10125_ ;
	wire _w10126_ ;
	wire _w10127_ ;
	wire _w10128_ ;
	wire _w10129_ ;
	wire _w10130_ ;
	wire _w10131_ ;
	wire _w10132_ ;
	wire _w10133_ ;
	wire _w10134_ ;
	wire _w10135_ ;
	wire _w10136_ ;
	wire _w10137_ ;
	wire _w10138_ ;
	wire _w10139_ ;
	wire _w10140_ ;
	wire _w10141_ ;
	wire _w10142_ ;
	wire _w10143_ ;
	wire _w10144_ ;
	wire _w10145_ ;
	wire _w10146_ ;
	wire _w10147_ ;
	wire _w10148_ ;
	wire _w10149_ ;
	wire _w10150_ ;
	wire _w10151_ ;
	wire _w10152_ ;
	wire _w10153_ ;
	wire _w10154_ ;
	wire _w10155_ ;
	wire _w10156_ ;
	wire _w10157_ ;
	wire _w10158_ ;
	wire _w10159_ ;
	wire _w10160_ ;
	wire _w10161_ ;
	wire _w10162_ ;
	wire _w10163_ ;
	wire _w10164_ ;
	wire _w10165_ ;
	wire _w10166_ ;
	wire _w10167_ ;
	wire _w10168_ ;
	wire _w10169_ ;
	wire _w10170_ ;
	wire _w10171_ ;
	wire _w10172_ ;
	wire _w10173_ ;
	wire _w10174_ ;
	wire _w10175_ ;
	wire _w10176_ ;
	wire _w10177_ ;
	wire _w10178_ ;
	wire _w10179_ ;
	wire _w10180_ ;
	wire _w10181_ ;
	wire _w10182_ ;
	wire _w10183_ ;
	wire _w10184_ ;
	wire _w10185_ ;
	wire _w10186_ ;
	wire _w10187_ ;
	wire _w10188_ ;
	wire _w10189_ ;
	wire _w10190_ ;
	wire _w10191_ ;
	wire _w10192_ ;
	wire _w10193_ ;
	wire _w10194_ ;
	wire _w10195_ ;
	wire _w10196_ ;
	wire _w10197_ ;
	wire _w10198_ ;
	wire _w10199_ ;
	wire _w10200_ ;
	wire _w10201_ ;
	wire _w10202_ ;
	wire _w10203_ ;
	wire _w10204_ ;
	wire _w10205_ ;
	wire _w10206_ ;
	wire _w10207_ ;
	wire _w10208_ ;
	wire _w10209_ ;
	wire _w10210_ ;
	wire _w10211_ ;
	wire _w10212_ ;
	wire _w10213_ ;
	wire _w10214_ ;
	wire _w10215_ ;
	wire _w10216_ ;
	wire _w10217_ ;
	wire _w10218_ ;
	wire _w10219_ ;
	wire _w10220_ ;
	wire _w10221_ ;
	wire _w10222_ ;
	wire _w10223_ ;
	wire _w10224_ ;
	wire _w10225_ ;
	wire _w10226_ ;
	wire _w10227_ ;
	wire _w10228_ ;
	wire _w10229_ ;
	wire _w10230_ ;
	wire _w10231_ ;
	wire _w10232_ ;
	wire _w10233_ ;
	wire _w10234_ ;
	wire _w10235_ ;
	wire _w10236_ ;
	wire _w10237_ ;
	wire _w10238_ ;
	wire _w10239_ ;
	wire _w10240_ ;
	wire _w10241_ ;
	wire _w10242_ ;
	wire _w10243_ ;
	wire _w10244_ ;
	wire _w10245_ ;
	wire _w10246_ ;
	wire _w10247_ ;
	wire _w10248_ ;
	wire _w10249_ ;
	wire _w10250_ ;
	wire _w10251_ ;
	wire _w10252_ ;
	wire _w10253_ ;
	wire _w10254_ ;
	wire _w10255_ ;
	wire _w10256_ ;
	wire _w10257_ ;
	wire _w10258_ ;
	wire _w10259_ ;
	wire _w10260_ ;
	wire _w10261_ ;
	wire _w10262_ ;
	wire _w10263_ ;
	wire _w10264_ ;
	wire _w10265_ ;
	wire _w10266_ ;
	wire _w10267_ ;
	wire _w10268_ ;
	wire _w10269_ ;
	wire _w10270_ ;
	wire _w10271_ ;
	wire _w10272_ ;
	wire _w10273_ ;
	wire _w10274_ ;
	wire _w10275_ ;
	wire _w10276_ ;
	wire _w10277_ ;
	wire _w10278_ ;
	wire _w10279_ ;
	wire _w10280_ ;
	wire _w10281_ ;
	wire _w10282_ ;
	wire _w10283_ ;
	wire _w10284_ ;
	wire _w10285_ ;
	wire _w10286_ ;
	wire _w10287_ ;
	wire _w10288_ ;
	wire _w10289_ ;
	wire _w10290_ ;
	wire _w10291_ ;
	wire _w10292_ ;
	wire _w10293_ ;
	wire _w10294_ ;
	wire _w10295_ ;
	wire _w10296_ ;
	wire _w10297_ ;
	wire _w10298_ ;
	wire _w10299_ ;
	wire _w10300_ ;
	wire _w10301_ ;
	wire _w10302_ ;
	wire _w10303_ ;
	wire _w10304_ ;
	wire _w10305_ ;
	wire _w10306_ ;
	wire _w10307_ ;
	wire _w10308_ ;
	wire _w10309_ ;
	wire _w10310_ ;
	wire _w10311_ ;
	wire _w10312_ ;
	wire _w10313_ ;
	wire _w10314_ ;
	wire _w10315_ ;
	wire _w10316_ ;
	wire _w10317_ ;
	wire _w10318_ ;
	wire _w10319_ ;
	wire _w10320_ ;
	wire _w10321_ ;
	wire _w10322_ ;
	wire _w10323_ ;
	wire _w10324_ ;
	wire _w10325_ ;
	wire _w10326_ ;
	wire _w10327_ ;
	wire _w10328_ ;
	wire _w10329_ ;
	wire _w10330_ ;
	wire _w10331_ ;
	wire _w10332_ ;
	wire _w10333_ ;
	wire _w10334_ ;
	wire _w10335_ ;
	wire _w10336_ ;
	wire _w10337_ ;
	wire _w10338_ ;
	wire _w10339_ ;
	wire _w10340_ ;
	wire _w10341_ ;
	wire _w10342_ ;
	wire _w10343_ ;
	wire _w10344_ ;
	wire _w10345_ ;
	wire _w10346_ ;
	wire _w10347_ ;
	wire _w10348_ ;
	wire _w10349_ ;
	wire _w10350_ ;
	wire _w10351_ ;
	wire _w10352_ ;
	wire _w10353_ ;
	wire _w10354_ ;
	wire _w10355_ ;
	wire _w10356_ ;
	wire _w10357_ ;
	wire _w10358_ ;
	wire _w10359_ ;
	wire _w10360_ ;
	wire _w10361_ ;
	wire _w10362_ ;
	wire _w10363_ ;
	wire _w10364_ ;
	wire _w10365_ ;
	wire _w10366_ ;
	wire _w10367_ ;
	wire _w10368_ ;
	wire _w10369_ ;
	wire _w10370_ ;
	wire _w10371_ ;
	wire _w10372_ ;
	wire _w10373_ ;
	wire _w10374_ ;
	wire _w10375_ ;
	wire _w10376_ ;
	wire _w10377_ ;
	wire _w10378_ ;
	wire _w10379_ ;
	wire _w10380_ ;
	wire _w10381_ ;
	wire _w10382_ ;
	wire _w10383_ ;
	wire _w10384_ ;
	wire _w10385_ ;
	wire _w10386_ ;
	wire _w10387_ ;
	wire _w10388_ ;
	wire _w10389_ ;
	wire _w10390_ ;
	wire _w10391_ ;
	wire _w10392_ ;
	wire _w10393_ ;
	wire _w10394_ ;
	wire _w10395_ ;
	wire _w10396_ ;
	wire _w10397_ ;
	wire _w10398_ ;
	wire _w10399_ ;
	wire _w10400_ ;
	wire _w10401_ ;
	wire _w10402_ ;
	wire _w10403_ ;
	wire _w10404_ ;
	wire _w10405_ ;
	wire _w10406_ ;
	wire _w10407_ ;
	wire _w10408_ ;
	wire _w10409_ ;
	wire _w10410_ ;
	wire _w10411_ ;
	wire _w10412_ ;
	wire _w10413_ ;
	wire _w10414_ ;
	wire _w10415_ ;
	wire _w10416_ ;
	wire _w10417_ ;
	wire _w10418_ ;
	wire _w10419_ ;
	wire _w10420_ ;
	wire _w10421_ ;
	wire _w10422_ ;
	wire _w10423_ ;
	wire _w10424_ ;
	wire _w10425_ ;
	wire _w10426_ ;
	wire _w10427_ ;
	wire _w10428_ ;
	wire _w10429_ ;
	wire _w10430_ ;
	wire _w10431_ ;
	wire _w10432_ ;
	wire _w10433_ ;
	wire _w10434_ ;
	wire _w10435_ ;
	wire _w10436_ ;
	wire _w10437_ ;
	wire _w10438_ ;
	wire _w10439_ ;
	wire _w10440_ ;
	wire _w10441_ ;
	wire _w10442_ ;
	wire _w10443_ ;
	wire _w10444_ ;
	wire _w10445_ ;
	wire _w10446_ ;
	wire _w10447_ ;
	wire _w10448_ ;
	wire _w10449_ ;
	wire _w10450_ ;
	wire _w10451_ ;
	wire _w10452_ ;
	wire _w10453_ ;
	wire _w10454_ ;
	wire _w10455_ ;
	wire _w10456_ ;
	wire _w10457_ ;
	wire _w10458_ ;
	wire _w10459_ ;
	wire _w10460_ ;
	wire _w10461_ ;
	wire _w10462_ ;
	wire _w10463_ ;
	wire _w10464_ ;
	wire _w10465_ ;
	wire _w10466_ ;
	wire _w10467_ ;
	wire _w10468_ ;
	wire _w10469_ ;
	wire _w10470_ ;
	wire _w10471_ ;
	wire _w10472_ ;
	wire _w10473_ ;
	wire _w10474_ ;
	wire _w10475_ ;
	wire _w10476_ ;
	wire _w10477_ ;
	wire _w10478_ ;
	wire _w10479_ ;
	wire _w10480_ ;
	wire _w10481_ ;
	wire _w10482_ ;
	wire _w10483_ ;
	wire _w10484_ ;
	wire _w10485_ ;
	wire _w10486_ ;
	wire _w10487_ ;
	wire _w10488_ ;
	wire _w10489_ ;
	wire _w10490_ ;
	wire _w10491_ ;
	wire _w10492_ ;
	wire _w10493_ ;
	wire _w10494_ ;
	wire _w10495_ ;
	wire _w10496_ ;
	wire _w10497_ ;
	wire _w10498_ ;
	wire _w10499_ ;
	wire _w10500_ ;
	wire _w10501_ ;
	wire _w10502_ ;
	wire _w10503_ ;
	wire _w10504_ ;
	wire _w10505_ ;
	wire _w10506_ ;
	wire _w10507_ ;
	wire _w10508_ ;
	wire _w10509_ ;
	wire _w10510_ ;
	wire _w10511_ ;
	wire _w10512_ ;
	wire _w10513_ ;
	wire _w10514_ ;
	wire _w10515_ ;
	wire _w10516_ ;
	wire _w10517_ ;
	wire _w10518_ ;
	wire _w10519_ ;
	wire _w10520_ ;
	wire _w10521_ ;
	wire _w10522_ ;
	wire _w10523_ ;
	wire _w10524_ ;
	wire _w10525_ ;
	wire _w10526_ ;
	wire _w10527_ ;
	wire _w10528_ ;
	wire _w10529_ ;
	wire _w10530_ ;
	wire _w10531_ ;
	wire _w10532_ ;
	wire _w10533_ ;
	wire _w10534_ ;
	wire _w10535_ ;
	wire _w10536_ ;
	wire _w10537_ ;
	wire _w10538_ ;
	wire _w10539_ ;
	wire _w10540_ ;
	wire _w10541_ ;
	wire _w10542_ ;
	wire _w10543_ ;
	wire _w10544_ ;
	wire _w10545_ ;
	wire _w10546_ ;
	wire _w10547_ ;
	wire _w10548_ ;
	wire _w10549_ ;
	wire _w10550_ ;
	wire _w10551_ ;
	wire _w10552_ ;
	wire _w10553_ ;
	wire _w10554_ ;
	wire _w10555_ ;
	wire _w10556_ ;
	wire _w10557_ ;
	wire _w10558_ ;
	wire _w10559_ ;
	wire _w10560_ ;
	wire _w10561_ ;
	wire _w10562_ ;
	wire _w10563_ ;
	wire _w10564_ ;
	wire _w10565_ ;
	wire _w10566_ ;
	wire _w10567_ ;
	wire _w10568_ ;
	wire _w10569_ ;
	wire _w10570_ ;
	wire _w10571_ ;
	wire _w10572_ ;
	wire _w10573_ ;
	wire _w10574_ ;
	wire _w10575_ ;
	wire _w10576_ ;
	wire _w10577_ ;
	wire _w10578_ ;
	wire _w10579_ ;
	wire _w10580_ ;
	wire _w10581_ ;
	wire _w10582_ ;
	wire _w10583_ ;
	wire _w10584_ ;
	wire _w10585_ ;
	wire _w10586_ ;
	wire _w10587_ ;
	wire _w10588_ ;
	wire _w10589_ ;
	wire _w10590_ ;
	wire _w10591_ ;
	wire _w10592_ ;
	wire _w10593_ ;
	wire _w10594_ ;
	wire _w10595_ ;
	wire _w10596_ ;
	wire _w10597_ ;
	wire _w10598_ ;
	wire _w10599_ ;
	wire _w10600_ ;
	wire _w10601_ ;
	wire _w10602_ ;
	wire _w10603_ ;
	wire _w10604_ ;
	wire _w10605_ ;
	wire _w10606_ ;
	wire _w10607_ ;
	wire _w10608_ ;
	wire _w10609_ ;
	wire _w10610_ ;
	wire _w10611_ ;
	wire _w10612_ ;
	wire _w10613_ ;
	wire _w10614_ ;
	wire _w10615_ ;
	wire _w10616_ ;
	wire _w10617_ ;
	wire _w10618_ ;
	wire _w10619_ ;
	wire _w10620_ ;
	wire _w10621_ ;
	wire _w10622_ ;
	wire _w10623_ ;
	wire _w10624_ ;
	wire _w10625_ ;
	wire _w10626_ ;
	wire _w10627_ ;
	wire _w10628_ ;
	wire _w10629_ ;
	wire _w10630_ ;
	wire _w10631_ ;
	wire _w10632_ ;
	wire _w10633_ ;
	wire _w10634_ ;
	wire _w10635_ ;
	wire _w10636_ ;
	wire _w10637_ ;
	wire _w10638_ ;
	wire _w10639_ ;
	wire _w10640_ ;
	wire _w10641_ ;
	wire _w10642_ ;
	wire _w10643_ ;
	wire _w10644_ ;
	wire _w10645_ ;
	wire _w10646_ ;
	wire _w10647_ ;
	wire _w10648_ ;
	wire _w10649_ ;
	wire _w10650_ ;
	wire _w10651_ ;
	wire _w10652_ ;
	wire _w10653_ ;
	wire _w10654_ ;
	wire _w10655_ ;
	wire _w10656_ ;
	wire _w10657_ ;
	wire _w10658_ ;
	wire _w10659_ ;
	wire _w10660_ ;
	wire _w10661_ ;
	wire _w10662_ ;
	wire _w10663_ ;
	wire _w10664_ ;
	wire _w10665_ ;
	wire _w10666_ ;
	wire _w10667_ ;
	wire _w10668_ ;
	wire _w10669_ ;
	wire _w10670_ ;
	wire _w10671_ ;
	wire _w10672_ ;
	wire _w10673_ ;
	wire _w10674_ ;
	wire _w10675_ ;
	wire _w10676_ ;
	wire _w10677_ ;
	wire _w10678_ ;
	wire _w10679_ ;
	wire _w10680_ ;
	wire _w10681_ ;
	wire _w10682_ ;
	wire _w10683_ ;
	wire _w10684_ ;
	wire _w10685_ ;
	wire _w10686_ ;
	wire _w10687_ ;
	wire _w10688_ ;
	wire _w10689_ ;
	wire _w10690_ ;
	wire _w10691_ ;
	wire _w10692_ ;
	wire _w10693_ ;
	wire _w10694_ ;
	wire _w10695_ ;
	wire _w10696_ ;
	wire _w10697_ ;
	wire _w10698_ ;
	wire _w10699_ ;
	wire _w10700_ ;
	wire _w10701_ ;
	wire _w10702_ ;
	wire _w10703_ ;
	wire _w10704_ ;
	wire _w10705_ ;
	wire _w10706_ ;
	wire _w10707_ ;
	wire _w10708_ ;
	wire _w10709_ ;
	wire _w10710_ ;
	wire _w10711_ ;
	wire _w10712_ ;
	wire _w10713_ ;
	wire _w10714_ ;
	wire _w10715_ ;
	wire _w10716_ ;
	wire _w10717_ ;
	wire _w10718_ ;
	wire _w10719_ ;
	wire _w10720_ ;
	wire _w10721_ ;
	wire _w10722_ ;
	wire _w10723_ ;
	wire _w10724_ ;
	wire _w10725_ ;
	wire _w10726_ ;
	wire _w10727_ ;
	wire _w10728_ ;
	wire _w10729_ ;
	wire _w10730_ ;
	wire _w10731_ ;
	wire _w10732_ ;
	wire _w10733_ ;
	wire _w10734_ ;
	LUT2 #(
		.INIT('h1)
	) name0 (
		\P1_IR_reg[6]/NET0131 ,
		\P1_IR_reg[7]/NET0131 ,
		_w462_
	);
	LUT2 #(
		.INIT('h1)
	) name1 (
		\P1_IR_reg[0]/NET0131 ,
		\P1_IR_reg[1]/NET0131 ,
		_w463_
	);
	LUT2 #(
		.INIT('h4)
	) name2 (
		\P1_IR_reg[2]/NET0131 ,
		_w463_,
		_w464_
	);
	LUT2 #(
		.INIT('h1)
	) name3 (
		\P1_IR_reg[3]/NET0131 ,
		\P1_IR_reg[4]/NET0131 ,
		_w465_
	);
	LUT2 #(
		.INIT('h4)
	) name4 (
		\P1_IR_reg[5]/NET0131 ,
		_w465_,
		_w466_
	);
	LUT2 #(
		.INIT('h8)
	) name5 (
		_w464_,
		_w466_,
		_w467_
	);
	LUT2 #(
		.INIT('h8)
	) name6 (
		_w462_,
		_w467_,
		_w468_
	);
	LUT2 #(
		.INIT('h1)
	) name7 (
		\P1_IR_reg[10]/NET0131 ,
		\P1_IR_reg[9]/NET0131 ,
		_w469_
	);
	LUT2 #(
		.INIT('h4)
	) name8 (
		\P1_IR_reg[11]/NET0131 ,
		_w469_,
		_w470_
	);
	LUT2 #(
		.INIT('h4)
	) name9 (
		\P1_IR_reg[12]/NET0131 ,
		_w470_,
		_w471_
	);
	LUT2 #(
		.INIT('h1)
	) name10 (
		\P1_IR_reg[13]/NET0131 ,
		\P1_IR_reg[8]/NET0131 ,
		_w472_
	);
	LUT2 #(
		.INIT('h8)
	) name11 (
		_w471_,
		_w472_,
		_w473_
	);
	LUT2 #(
		.INIT('h8)
	) name12 (
		_w468_,
		_w473_,
		_w474_
	);
	LUT2 #(
		.INIT('h1)
	) name13 (
		\P1_IR_reg[14]/NET0131 ,
		\P1_IR_reg[15]/NET0131 ,
		_w475_
	);
	LUT2 #(
		.INIT('h1)
	) name14 (
		\P1_IR_reg[17]/NET0131 ,
		\P1_IR_reg[18]/NET0131 ,
		_w476_
	);
	LUT2 #(
		.INIT('h4)
	) name15 (
		\P1_IR_reg[19]/NET0131 ,
		_w476_,
		_w477_
	);
	LUT2 #(
		.INIT('h4)
	) name16 (
		\P1_IR_reg[16]/NET0131 ,
		_w477_,
		_w478_
	);
	LUT2 #(
		.INIT('h1)
	) name17 (
		\P1_IR_reg[20]/NET0131 ,
		\P1_IR_reg[21]/NET0131 ,
		_w479_
	);
	LUT2 #(
		.INIT('h8)
	) name18 (
		_w475_,
		_w479_,
		_w480_
	);
	LUT2 #(
		.INIT('h8)
	) name19 (
		_w478_,
		_w480_,
		_w481_
	);
	LUT2 #(
		.INIT('h8)
	) name20 (
		_w474_,
		_w481_,
		_w482_
	);
	LUT2 #(
		.INIT('h2)
	) name21 (
		\P1_IR_reg[31]/NET0131 ,
		_w482_,
		_w483_
	);
	LUT2 #(
		.INIT('h8)
	) name22 (
		\P1_IR_reg[22]/NET0131 ,
		_w483_,
		_w484_
	);
	LUT2 #(
		.INIT('h1)
	) name23 (
		\P1_IR_reg[22]/NET0131 ,
		_w483_,
		_w485_
	);
	LUT2 #(
		.INIT('h1)
	) name24 (
		_w484_,
		_w485_,
		_w486_
	);
	LUT2 #(
		.INIT('h4)
	) name25 (
		\P1_IR_reg[3]/NET0131 ,
		_w464_,
		_w487_
	);
	LUT2 #(
		.INIT('h4)
	) name26 (
		\P1_IR_reg[4]/NET0131 ,
		_w487_,
		_w488_
	);
	LUT2 #(
		.INIT('h4)
	) name27 (
		\P1_IR_reg[8]/NET0131 ,
		_w462_,
		_w489_
	);
	LUT2 #(
		.INIT('h4)
	) name28 (
		\P1_IR_reg[5]/NET0131 ,
		_w489_,
		_w490_
	);
	LUT2 #(
		.INIT('h8)
	) name29 (
		_w488_,
		_w490_,
		_w491_
	);
	LUT2 #(
		.INIT('h1)
	) name30 (
		\P1_IR_reg[13]/NET0131 ,
		\P1_IR_reg[16]/NET0131 ,
		_w492_
	);
	LUT2 #(
		.INIT('h8)
	) name31 (
		_w475_,
		_w492_,
		_w493_
	);
	LUT2 #(
		.INIT('h8)
	) name32 (
		_w471_,
		_w493_,
		_w494_
	);
	LUT2 #(
		.INIT('h8)
	) name33 (
		_w491_,
		_w494_,
		_w495_
	);
	LUT2 #(
		.INIT('h4)
	) name34 (
		\P1_IR_reg[20]/NET0131 ,
		_w477_,
		_w496_
	);
	LUT2 #(
		.INIT('h8)
	) name35 (
		_w495_,
		_w496_,
		_w497_
	);
	LUT2 #(
		.INIT('h2)
	) name36 (
		\P1_IR_reg[31]/NET0131 ,
		_w497_,
		_w498_
	);
	LUT2 #(
		.INIT('h8)
	) name37 (
		\P1_IR_reg[21]/NET0131 ,
		_w498_,
		_w499_
	);
	LUT2 #(
		.INIT('h1)
	) name38 (
		\P1_IR_reg[21]/NET0131 ,
		_w498_,
		_w500_
	);
	LUT2 #(
		.INIT('h1)
	) name39 (
		_w499_,
		_w500_,
		_w501_
	);
	LUT2 #(
		.INIT('h4)
	) name40 (
		\P1_IR_reg[22]/NET0131 ,
		_w479_,
		_w502_
	);
	LUT2 #(
		.INIT('h4)
	) name41 (
		\P1_IR_reg[14]/NET0131 ,
		_w474_,
		_w503_
	);
	LUT2 #(
		.INIT('h1)
	) name42 (
		\P1_IR_reg[15]/NET0131 ,
		\P1_IR_reg[16]/NET0131 ,
		_w504_
	);
	LUT2 #(
		.INIT('h8)
	) name43 (
		_w476_,
		_w504_,
		_w505_
	);
	LUT2 #(
		.INIT('h8)
	) name44 (
		_w503_,
		_w505_,
		_w506_
	);
	LUT2 #(
		.INIT('h4)
	) name45 (
		\P1_IR_reg[19]/NET0131 ,
		_w502_,
		_w507_
	);
	LUT2 #(
		.INIT('h8)
	) name46 (
		_w506_,
		_w507_,
		_w508_
	);
	LUT2 #(
		.INIT('h2)
	) name47 (
		\P1_IR_reg[31]/NET0131 ,
		_w508_,
		_w509_
	);
	LUT2 #(
		.INIT('h4)
	) name48 (
		\P1_IR_reg[23]/NET0131 ,
		_w509_,
		_w510_
	);
	LUT2 #(
		.INIT('h2)
	) name49 (
		\P1_IR_reg[23]/NET0131 ,
		_w509_,
		_w511_
	);
	LUT2 #(
		.INIT('h1)
	) name50 (
		_w510_,
		_w511_,
		_w512_
	);
	LUT2 #(
		.INIT('h2)
	) name51 (
		\P1_B_reg/NET0131 ,
		_w512_,
		_w513_
	);
	LUT2 #(
		.INIT('h8)
	) name52 (
		_w474_,
		_w475_,
		_w514_
	);
	LUT2 #(
		.INIT('h8)
	) name53 (
		_w478_,
		_w514_,
		_w515_
	);
	LUT2 #(
		.INIT('h2)
	) name54 (
		\P1_IR_reg[31]/NET0131 ,
		_w515_,
		_w516_
	);
	LUT2 #(
		.INIT('h8)
	) name55 (
		\P1_IR_reg[20]/NET0131 ,
		_w516_,
		_w517_
	);
	LUT2 #(
		.INIT('h1)
	) name56 (
		\P1_IR_reg[20]/NET0131 ,
		_w516_,
		_w518_
	);
	LUT2 #(
		.INIT('h1)
	) name57 (
		_w517_,
		_w518_,
		_w519_
	);
	LUT2 #(
		.INIT('h1)
	) name58 (
		\P1_IR_reg[23]/NET0131 ,
		\P1_IR_reg[24]/NET0131 ,
		_w520_
	);
	LUT2 #(
		.INIT('h1)
	) name59 (
		\P1_IR_reg[25]/NET0131 ,
		\P1_IR_reg[26]/NET0131 ,
		_w521_
	);
	LUT2 #(
		.INIT('h8)
	) name60 (
		_w520_,
		_w521_,
		_w522_
	);
	LUT2 #(
		.INIT('h8)
	) name61 (
		_w508_,
		_w522_,
		_w523_
	);
	LUT2 #(
		.INIT('h2)
	) name62 (
		\P1_IR_reg[31]/NET0131 ,
		_w523_,
		_w524_
	);
	LUT2 #(
		.INIT('h8)
	) name63 (
		\P1_IR_reg[27]/NET0131 ,
		_w524_,
		_w525_
	);
	LUT2 #(
		.INIT('h1)
	) name64 (
		\P1_IR_reg[27]/NET0131 ,
		_w524_,
		_w526_
	);
	LUT2 #(
		.INIT('h1)
	) name65 (
		_w525_,
		_w526_,
		_w527_
	);
	LUT2 #(
		.INIT('h4)
	) name66 (
		\P1_IR_reg[23]/NET0131 ,
		_w502_,
		_w528_
	);
	LUT2 #(
		.INIT('h8)
	) name67 (
		_w515_,
		_w528_,
		_w529_
	);
	LUT2 #(
		.INIT('h2)
	) name68 (
		\P1_IR_reg[31]/NET0131 ,
		_w529_,
		_w530_
	);
	LUT2 #(
		.INIT('h1)
	) name69 (
		\P1_IR_reg[24]/NET0131 ,
		\P1_IR_reg[27]/NET0131 ,
		_w531_
	);
	LUT2 #(
		.INIT('h8)
	) name70 (
		_w521_,
		_w531_,
		_w532_
	);
	LUT2 #(
		.INIT('h2)
	) name71 (
		\P1_IR_reg[31]/NET0131 ,
		_w532_,
		_w533_
	);
	LUT2 #(
		.INIT('h1)
	) name72 (
		_w530_,
		_w533_,
		_w534_
	);
	LUT2 #(
		.INIT('h2)
	) name73 (
		\P1_IR_reg[28]/NET0131 ,
		_w534_,
		_w535_
	);
	LUT2 #(
		.INIT('h4)
	) name74 (
		\P1_IR_reg[28]/NET0131 ,
		_w534_,
		_w536_
	);
	LUT2 #(
		.INIT('h1)
	) name75 (
		_w535_,
		_w536_,
		_w537_
	);
	LUT2 #(
		.INIT('h1)
	) name76 (
		_w527_,
		_w537_,
		_w538_
	);
	LUT2 #(
		.INIT('h1)
	) name77 (
		\P1_addr_reg[19]/NET0131 ,
		\P2_addr_reg[19]/NET0131 ,
		_w539_
	);
	LUT2 #(
		.INIT('h4)
	) name78 (
		\P1_rd_reg/NET0131 ,
		_w539_,
		_w540_
	);
	LUT2 #(
		.INIT('h8)
	) name79 (
		\P1_addr_reg[19]/NET0131 ,
		\P2_addr_reg[19]/NET0131 ,
		_w541_
	);
	LUT2 #(
		.INIT('h4)
	) name80 (
		\P2_rd_reg/NET0131 ,
		_w541_,
		_w542_
	);
	LUT2 #(
		.INIT('h1)
	) name81 (
		_w540_,
		_w542_,
		_w543_
	);
	LUT2 #(
		.INIT('h1)
	) name82 (
		\P2_datao_reg[22]/NET0131 ,
		\si[22]_pad ,
		_w544_
	);
	LUT2 #(
		.INIT('h8)
	) name83 (
		\P2_datao_reg[22]/NET0131 ,
		\si[22]_pad ,
		_w545_
	);
	LUT2 #(
		.INIT('h8)
	) name84 (
		\P2_datao_reg[21]/NET0131 ,
		\si[21]_pad ,
		_w546_
	);
	LUT2 #(
		.INIT('h1)
	) name85 (
		_w545_,
		_w546_,
		_w547_
	);
	LUT2 #(
		.INIT('h1)
	) name86 (
		_w544_,
		_w547_,
		_w548_
	);
	LUT2 #(
		.INIT('h1)
	) name87 (
		\P2_datao_reg[21]/NET0131 ,
		\si[21]_pad ,
		_w549_
	);
	LUT2 #(
		.INIT('h1)
	) name88 (
		_w544_,
		_w549_,
		_w550_
	);
	LUT2 #(
		.INIT('h1)
	) name89 (
		\P2_datao_reg[20]/NET0131 ,
		\si[20]_pad ,
		_w551_
	);
	LUT2 #(
		.INIT('h8)
	) name90 (
		\P2_datao_reg[20]/NET0131 ,
		\si[20]_pad ,
		_w552_
	);
	LUT2 #(
		.INIT('h8)
	) name91 (
		\P2_datao_reg[19]/NET0131 ,
		\si[19]_pad ,
		_w553_
	);
	LUT2 #(
		.INIT('h1)
	) name92 (
		_w552_,
		_w553_,
		_w554_
	);
	LUT2 #(
		.INIT('h1)
	) name93 (
		_w551_,
		_w554_,
		_w555_
	);
	LUT2 #(
		.INIT('h8)
	) name94 (
		_w550_,
		_w555_,
		_w556_
	);
	LUT2 #(
		.INIT('h1)
	) name95 (
		_w548_,
		_w556_,
		_w557_
	);
	LUT2 #(
		.INIT('h1)
	) name96 (
		\P2_datao_reg[19]/NET0131 ,
		\si[19]_pad ,
		_w558_
	);
	LUT2 #(
		.INIT('h1)
	) name97 (
		_w551_,
		_w558_,
		_w559_
	);
	LUT2 #(
		.INIT('h8)
	) name98 (
		_w550_,
		_w559_,
		_w560_
	);
	LUT2 #(
		.INIT('h1)
	) name99 (
		\P2_datao_reg[18]/NET0131 ,
		\si[18]_pad ,
		_w561_
	);
	LUT2 #(
		.INIT('h8)
	) name100 (
		\P2_datao_reg[18]/NET0131 ,
		\si[18]_pad ,
		_w562_
	);
	LUT2 #(
		.INIT('h8)
	) name101 (
		\P2_datao_reg[17]/NET0131 ,
		\si[17]_pad ,
		_w563_
	);
	LUT2 #(
		.INIT('h1)
	) name102 (
		_w562_,
		_w563_,
		_w564_
	);
	LUT2 #(
		.INIT('h1)
	) name103 (
		_w561_,
		_w564_,
		_w565_
	);
	LUT2 #(
		.INIT('h1)
	) name104 (
		\P2_datao_reg[17]/NET0131 ,
		\si[17]_pad ,
		_w566_
	);
	LUT2 #(
		.INIT('h1)
	) name105 (
		_w561_,
		_w566_,
		_w567_
	);
	LUT2 #(
		.INIT('h1)
	) name106 (
		\P2_datao_reg[16]/NET0131 ,
		\si[16]_pad ,
		_w568_
	);
	LUT2 #(
		.INIT('h8)
	) name107 (
		\P2_datao_reg[15]/NET0131 ,
		\si[15]_pad ,
		_w569_
	);
	LUT2 #(
		.INIT('h8)
	) name108 (
		\P2_datao_reg[16]/NET0131 ,
		\si[16]_pad ,
		_w570_
	);
	LUT2 #(
		.INIT('h1)
	) name109 (
		_w569_,
		_w570_,
		_w571_
	);
	LUT2 #(
		.INIT('h1)
	) name110 (
		_w568_,
		_w571_,
		_w572_
	);
	LUT2 #(
		.INIT('h8)
	) name111 (
		_w567_,
		_w572_,
		_w573_
	);
	LUT2 #(
		.INIT('h1)
	) name112 (
		_w565_,
		_w573_,
		_w574_
	);
	LUT2 #(
		.INIT('h1)
	) name113 (
		\P2_datao_reg[14]/NET0131 ,
		\si[14]_pad ,
		_w575_
	);
	LUT2 #(
		.INIT('h8)
	) name114 (
		\P2_datao_reg[14]/NET0131 ,
		\si[14]_pad ,
		_w576_
	);
	LUT2 #(
		.INIT('h8)
	) name115 (
		\P2_datao_reg[13]/NET0131 ,
		\si[13]_pad ,
		_w577_
	);
	LUT2 #(
		.INIT('h1)
	) name116 (
		_w576_,
		_w577_,
		_w578_
	);
	LUT2 #(
		.INIT('h1)
	) name117 (
		_w575_,
		_w578_,
		_w579_
	);
	LUT2 #(
		.INIT('h1)
	) name118 (
		\P2_datao_reg[13]/NET0131 ,
		\si[13]_pad ,
		_w580_
	);
	LUT2 #(
		.INIT('h1)
	) name119 (
		_w575_,
		_w580_,
		_w581_
	);
	LUT2 #(
		.INIT('h1)
	) name120 (
		\P2_datao_reg[12]/NET0131 ,
		\si[12]_pad ,
		_w582_
	);
	LUT2 #(
		.INIT('h8)
	) name121 (
		\P2_datao_reg[12]/NET0131 ,
		\si[12]_pad ,
		_w583_
	);
	LUT2 #(
		.INIT('h8)
	) name122 (
		\P2_datao_reg[11]/NET0131 ,
		\si[11]_pad ,
		_w584_
	);
	LUT2 #(
		.INIT('h1)
	) name123 (
		_w583_,
		_w584_,
		_w585_
	);
	LUT2 #(
		.INIT('h1)
	) name124 (
		_w582_,
		_w585_,
		_w586_
	);
	LUT2 #(
		.INIT('h8)
	) name125 (
		_w581_,
		_w586_,
		_w587_
	);
	LUT2 #(
		.INIT('h1)
	) name126 (
		_w579_,
		_w587_,
		_w588_
	);
	LUT2 #(
		.INIT('h8)
	) name127 (
		\P2_datao_reg[8]/NET0131 ,
		\si[8]_pad ,
		_w589_
	);
	LUT2 #(
		.INIT('h8)
	) name128 (
		\P2_datao_reg[7]/NET0131 ,
		\si[7]_pad ,
		_w590_
	);
	LUT2 #(
		.INIT('h1)
	) name129 (
		_w589_,
		_w590_,
		_w591_
	);
	LUT2 #(
		.INIT('h1)
	) name130 (
		\P2_datao_reg[9]/NET0131 ,
		\si[9]_pad ,
		_w592_
	);
	LUT2 #(
		.INIT('h1)
	) name131 (
		\P2_datao_reg[10]/NET0131 ,
		\si[10]_pad ,
		_w593_
	);
	LUT2 #(
		.INIT('h1)
	) name132 (
		_w592_,
		_w593_,
		_w594_
	);
	LUT2 #(
		.INIT('h1)
	) name133 (
		\P2_datao_reg[8]/NET0131 ,
		\si[8]_pad ,
		_w595_
	);
	LUT2 #(
		.INIT('h2)
	) name134 (
		_w594_,
		_w595_,
		_w596_
	);
	LUT2 #(
		.INIT('h4)
	) name135 (
		_w591_,
		_w596_,
		_w597_
	);
	LUT2 #(
		.INIT('h8)
	) name136 (
		\P2_datao_reg[9]/NET0131 ,
		\si[9]_pad ,
		_w598_
	);
	LUT2 #(
		.INIT('h8)
	) name137 (
		\P2_datao_reg[10]/NET0131 ,
		\si[10]_pad ,
		_w599_
	);
	LUT2 #(
		.INIT('h1)
	) name138 (
		_w598_,
		_w599_,
		_w600_
	);
	LUT2 #(
		.INIT('h1)
	) name139 (
		_w593_,
		_w600_,
		_w601_
	);
	LUT2 #(
		.INIT('h1)
	) name140 (
		\P2_datao_reg[6]/NET0131 ,
		\si[6]_pad ,
		_w602_
	);
	LUT2 #(
		.INIT('h8)
	) name141 (
		\P2_datao_reg[5]/NET0131 ,
		\si[5]_pad ,
		_w603_
	);
	LUT2 #(
		.INIT('h8)
	) name142 (
		\P2_datao_reg[6]/NET0131 ,
		\si[6]_pad ,
		_w604_
	);
	LUT2 #(
		.INIT('h1)
	) name143 (
		_w603_,
		_w604_,
		_w605_
	);
	LUT2 #(
		.INIT('h1)
	) name144 (
		_w602_,
		_w605_,
		_w606_
	);
	LUT2 #(
		.INIT('h8)
	) name145 (
		\P2_datao_reg[4]/NET0131 ,
		\si[4]_pad ,
		_w607_
	);
	LUT2 #(
		.INIT('h8)
	) name146 (
		\P2_datao_reg[3]/NET0131 ,
		\si[3]_pad ,
		_w608_
	);
	LUT2 #(
		.INIT('h1)
	) name147 (
		\P2_datao_reg[3]/NET0131 ,
		\si[3]_pad ,
		_w609_
	);
	LUT2 #(
		.INIT('h1)
	) name148 (
		\P2_datao_reg[2]/NET0131 ,
		\si[2]_pad ,
		_w610_
	);
	LUT2 #(
		.INIT('h1)
	) name149 (
		_w609_,
		_w610_,
		_w611_
	);
	LUT2 #(
		.INIT('h8)
	) name150 (
		\P2_datao_reg[0]/NET0131 ,
		\si[0]_pad ,
		_w612_
	);
	LUT2 #(
		.INIT('h1)
	) name151 (
		\P2_datao_reg[1]/NET0131 ,
		\si[1]_pad ,
		_w613_
	);
	LUT2 #(
		.INIT('h2)
	) name152 (
		_w612_,
		_w613_,
		_w614_
	);
	LUT2 #(
		.INIT('h8)
	) name153 (
		\P2_datao_reg[1]/NET0131 ,
		\si[1]_pad ,
		_w615_
	);
	LUT2 #(
		.INIT('h8)
	) name154 (
		\P2_datao_reg[2]/NET0131 ,
		\si[2]_pad ,
		_w616_
	);
	LUT2 #(
		.INIT('h1)
	) name155 (
		_w615_,
		_w616_,
		_w617_
	);
	LUT2 #(
		.INIT('h4)
	) name156 (
		_w614_,
		_w617_,
		_w618_
	);
	LUT2 #(
		.INIT('h2)
	) name157 (
		_w611_,
		_w618_,
		_w619_
	);
	LUT2 #(
		.INIT('h1)
	) name158 (
		_w608_,
		_w619_,
		_w620_
	);
	LUT2 #(
		.INIT('h4)
	) name159 (
		_w607_,
		_w620_,
		_w621_
	);
	LUT2 #(
		.INIT('h1)
	) name160 (
		\P2_datao_reg[5]/NET0131 ,
		\si[5]_pad ,
		_w622_
	);
	LUT2 #(
		.INIT('h1)
	) name161 (
		\P2_datao_reg[4]/NET0131 ,
		\si[4]_pad ,
		_w623_
	);
	LUT2 #(
		.INIT('h1)
	) name162 (
		_w622_,
		_w623_,
		_w624_
	);
	LUT2 #(
		.INIT('h4)
	) name163 (
		_w602_,
		_w624_,
		_w625_
	);
	LUT2 #(
		.INIT('h4)
	) name164 (
		_w621_,
		_w625_,
		_w626_
	);
	LUT2 #(
		.INIT('h1)
	) name165 (
		_w606_,
		_w626_,
		_w627_
	);
	LUT2 #(
		.INIT('h1)
	) name166 (
		\P2_datao_reg[7]/NET0131 ,
		\si[7]_pad ,
		_w628_
	);
	LUT2 #(
		.INIT('h1)
	) name167 (
		_w595_,
		_w628_,
		_w629_
	);
	LUT2 #(
		.INIT('h8)
	) name168 (
		_w594_,
		_w629_,
		_w630_
	);
	LUT2 #(
		.INIT('h4)
	) name169 (
		_w627_,
		_w630_,
		_w631_
	);
	LUT2 #(
		.INIT('h1)
	) name170 (
		_w597_,
		_w601_,
		_w632_
	);
	LUT2 #(
		.INIT('h4)
	) name171 (
		_w631_,
		_w632_,
		_w633_
	);
	LUT2 #(
		.INIT('h1)
	) name172 (
		\P2_datao_reg[11]/NET0131 ,
		\si[11]_pad ,
		_w634_
	);
	LUT2 #(
		.INIT('h1)
	) name173 (
		_w582_,
		_w634_,
		_w635_
	);
	LUT2 #(
		.INIT('h8)
	) name174 (
		_w581_,
		_w635_,
		_w636_
	);
	LUT2 #(
		.INIT('h4)
	) name175 (
		_w633_,
		_w636_,
		_w637_
	);
	LUT2 #(
		.INIT('h2)
	) name176 (
		_w588_,
		_w637_,
		_w638_
	);
	LUT2 #(
		.INIT('h1)
	) name177 (
		\P2_datao_reg[15]/NET0131 ,
		\si[15]_pad ,
		_w639_
	);
	LUT2 #(
		.INIT('h1)
	) name178 (
		_w568_,
		_w639_,
		_w640_
	);
	LUT2 #(
		.INIT('h8)
	) name179 (
		_w567_,
		_w640_,
		_w641_
	);
	LUT2 #(
		.INIT('h4)
	) name180 (
		_w638_,
		_w641_,
		_w642_
	);
	LUT2 #(
		.INIT('h2)
	) name181 (
		_w574_,
		_w642_,
		_w643_
	);
	LUT2 #(
		.INIT('h2)
	) name182 (
		_w560_,
		_w643_,
		_w644_
	);
	LUT2 #(
		.INIT('h2)
	) name183 (
		_w557_,
		_w644_,
		_w645_
	);
	LUT2 #(
		.INIT('h1)
	) name184 (
		\P2_datao_reg[30]/NET0131 ,
		\si[30]_pad ,
		_w646_
	);
	LUT2 #(
		.INIT('h1)
	) name185 (
		\P2_datao_reg[29]/NET0131 ,
		\si[29]_pad ,
		_w647_
	);
	LUT2 #(
		.INIT('h1)
	) name186 (
		\P2_datao_reg[27]/NET0131 ,
		\si[27]_pad ,
		_w648_
	);
	LUT2 #(
		.INIT('h1)
	) name187 (
		\P2_datao_reg[28]/NET0131 ,
		\si[28]_pad ,
		_w649_
	);
	LUT2 #(
		.INIT('h1)
	) name188 (
		_w648_,
		_w649_,
		_w650_
	);
	LUT2 #(
		.INIT('h4)
	) name189 (
		_w647_,
		_w650_,
		_w651_
	);
	LUT2 #(
		.INIT('h4)
	) name190 (
		_w646_,
		_w651_,
		_w652_
	);
	LUT2 #(
		.INIT('h1)
	) name191 (
		\P2_datao_reg[26]/NET0131 ,
		\si[26]_pad ,
		_w653_
	);
	LUT2 #(
		.INIT('h1)
	) name192 (
		\P2_datao_reg[25]/NET0131 ,
		\si[25]_pad ,
		_w654_
	);
	LUT2 #(
		.INIT('h1)
	) name193 (
		_w653_,
		_w654_,
		_w655_
	);
	LUT2 #(
		.INIT('h1)
	) name194 (
		\P2_datao_reg[24]/NET0131 ,
		\si[24]_pad ,
		_w656_
	);
	LUT2 #(
		.INIT('h1)
	) name195 (
		\P2_datao_reg[23]/NET0131 ,
		\si[23]_pad ,
		_w657_
	);
	LUT2 #(
		.INIT('h1)
	) name196 (
		_w656_,
		_w657_,
		_w658_
	);
	LUT2 #(
		.INIT('h8)
	) name197 (
		_w655_,
		_w658_,
		_w659_
	);
	LUT2 #(
		.INIT('h8)
	) name198 (
		_w652_,
		_w659_,
		_w660_
	);
	LUT2 #(
		.INIT('h4)
	) name199 (
		_w645_,
		_w660_,
		_w661_
	);
	LUT2 #(
		.INIT('h8)
	) name200 (
		\P2_datao_reg[29]/NET0131 ,
		\si[29]_pad ,
		_w662_
	);
	LUT2 #(
		.INIT('h8)
	) name201 (
		\P2_datao_reg[27]/NET0131 ,
		\si[27]_pad ,
		_w663_
	);
	LUT2 #(
		.INIT('h8)
	) name202 (
		\P2_datao_reg[28]/NET0131 ,
		\si[28]_pad ,
		_w664_
	);
	LUT2 #(
		.INIT('h1)
	) name203 (
		_w663_,
		_w664_,
		_w665_
	);
	LUT2 #(
		.INIT('h1)
	) name204 (
		_w647_,
		_w649_,
		_w666_
	);
	LUT2 #(
		.INIT('h4)
	) name205 (
		_w665_,
		_w666_,
		_w667_
	);
	LUT2 #(
		.INIT('h1)
	) name206 (
		_w662_,
		_w667_,
		_w668_
	);
	LUT2 #(
		.INIT('h1)
	) name207 (
		_w646_,
		_w668_,
		_w669_
	);
	LUT2 #(
		.INIT('h8)
	) name208 (
		\P2_datao_reg[26]/NET0131 ,
		\si[26]_pad ,
		_w670_
	);
	LUT2 #(
		.INIT('h8)
	) name209 (
		\P2_datao_reg[25]/NET0131 ,
		\si[25]_pad ,
		_w671_
	);
	LUT2 #(
		.INIT('h1)
	) name210 (
		_w670_,
		_w671_,
		_w672_
	);
	LUT2 #(
		.INIT('h1)
	) name211 (
		_w653_,
		_w672_,
		_w673_
	);
	LUT2 #(
		.INIT('h8)
	) name212 (
		\P2_datao_reg[24]/NET0131 ,
		\si[24]_pad ,
		_w674_
	);
	LUT2 #(
		.INIT('h8)
	) name213 (
		\P2_datao_reg[23]/NET0131 ,
		\si[23]_pad ,
		_w675_
	);
	LUT2 #(
		.INIT('h1)
	) name214 (
		_w674_,
		_w675_,
		_w676_
	);
	LUT2 #(
		.INIT('h1)
	) name215 (
		_w656_,
		_w676_,
		_w677_
	);
	LUT2 #(
		.INIT('h8)
	) name216 (
		_w655_,
		_w677_,
		_w678_
	);
	LUT2 #(
		.INIT('h1)
	) name217 (
		_w673_,
		_w678_,
		_w679_
	);
	LUT2 #(
		.INIT('h2)
	) name218 (
		_w652_,
		_w679_,
		_w680_
	);
	LUT2 #(
		.INIT('h8)
	) name219 (
		\P2_datao_reg[30]/NET0131 ,
		\si[30]_pad ,
		_w681_
	);
	LUT2 #(
		.INIT('h1)
	) name220 (
		_w669_,
		_w681_,
		_w682_
	);
	LUT2 #(
		.INIT('h4)
	) name221 (
		_w680_,
		_w682_,
		_w683_
	);
	LUT2 #(
		.INIT('h4)
	) name222 (
		_w661_,
		_w683_,
		_w684_
	);
	LUT2 #(
		.INIT('h2)
	) name223 (
		\si[31]_pad ,
		_w684_,
		_w685_
	);
	LUT2 #(
		.INIT('h4)
	) name224 (
		\si[31]_pad ,
		_w684_,
		_w686_
	);
	LUT2 #(
		.INIT('h1)
	) name225 (
		_w543_,
		_w685_,
		_w687_
	);
	LUT2 #(
		.INIT('h4)
	) name226 (
		_w686_,
		_w687_,
		_w688_
	);
	LUT2 #(
		.INIT('h8)
	) name227 (
		\P2_datao_reg[31]/NET0131 ,
		_w688_,
		_w689_
	);
	LUT2 #(
		.INIT('h1)
	) name228 (
		\P2_datao_reg[31]/NET0131 ,
		_w688_,
		_w690_
	);
	LUT2 #(
		.INIT('h1)
	) name229 (
		_w689_,
		_w690_,
		_w691_
	);
	LUT2 #(
		.INIT('h4)
	) name230 (
		_w538_,
		_w691_,
		_w692_
	);
	LUT2 #(
		.INIT('h1)
	) name231 (
		\P1_IR_reg[22]/NET0131 ,
		\P1_IR_reg[25]/NET0131 ,
		_w693_
	);
	LUT2 #(
		.INIT('h8)
	) name232 (
		_w520_,
		_w693_,
		_w694_
	);
	LUT2 #(
		.INIT('h8)
	) name233 (
		_w482_,
		_w694_,
		_w695_
	);
	LUT2 #(
		.INIT('h2)
	) name234 (
		\P1_IR_reg[31]/NET0131 ,
		_w695_,
		_w696_
	);
	LUT2 #(
		.INIT('h1)
	) name235 (
		\P1_IR_reg[27]/NET0131 ,
		\P1_IR_reg[28]/NET0131 ,
		_w697_
	);
	LUT2 #(
		.INIT('h4)
	) name236 (
		\P1_IR_reg[29]/NET0131 ,
		_w697_,
		_w698_
	);
	LUT2 #(
		.INIT('h4)
	) name237 (
		\P1_IR_reg[26]/NET0131 ,
		_w698_,
		_w699_
	);
	LUT2 #(
		.INIT('h2)
	) name238 (
		\P1_IR_reg[31]/NET0131 ,
		_w699_,
		_w700_
	);
	LUT2 #(
		.INIT('h1)
	) name239 (
		_w696_,
		_w700_,
		_w701_
	);
	LUT2 #(
		.INIT('h2)
	) name240 (
		\P1_IR_reg[30]/NET0131 ,
		_w701_,
		_w702_
	);
	LUT2 #(
		.INIT('h4)
	) name241 (
		\P1_IR_reg[30]/NET0131 ,
		_w701_,
		_w703_
	);
	LUT2 #(
		.INIT('h1)
	) name242 (
		_w702_,
		_w703_,
		_w704_
	);
	LUT2 #(
		.INIT('h4)
	) name243 (
		\P1_IR_reg[24]/NET0131 ,
		_w477_,
		_w705_
	);
	LUT2 #(
		.INIT('h8)
	) name244 (
		_w528_,
		_w705_,
		_w706_
	);
	LUT2 #(
		.INIT('h8)
	) name245 (
		_w495_,
		_w706_,
		_w707_
	);
	LUT2 #(
		.INIT('h2)
	) name246 (
		\P1_IR_reg[31]/NET0131 ,
		_w707_,
		_w708_
	);
	LUT2 #(
		.INIT('h8)
	) name247 (
		_w521_,
		_w697_,
		_w709_
	);
	LUT2 #(
		.INIT('h2)
	) name248 (
		\P1_IR_reg[31]/NET0131 ,
		_w709_,
		_w710_
	);
	LUT2 #(
		.INIT('h1)
	) name249 (
		_w708_,
		_w710_,
		_w711_
	);
	LUT2 #(
		.INIT('h2)
	) name250 (
		\P1_IR_reg[29]/NET0131 ,
		_w711_,
		_w712_
	);
	LUT2 #(
		.INIT('h4)
	) name251 (
		\P1_IR_reg[29]/NET0131 ,
		_w711_,
		_w713_
	);
	LUT2 #(
		.INIT('h1)
	) name252 (
		_w712_,
		_w713_,
		_w714_
	);
	LUT2 #(
		.INIT('h8)
	) name253 (
		_w704_,
		_w714_,
		_w715_
	);
	LUT2 #(
		.INIT('h8)
	) name254 (
		\P1_reg3_reg[3]/NET0131 ,
		\P1_reg3_reg[4]/NET0131 ,
		_w716_
	);
	LUT2 #(
		.INIT('h8)
	) name255 (
		\P1_reg3_reg[5]/NET0131 ,
		_w716_,
		_w717_
	);
	LUT2 #(
		.INIT('h8)
	) name256 (
		\P1_reg3_reg[6]/NET0131 ,
		_w717_,
		_w718_
	);
	LUT2 #(
		.INIT('h8)
	) name257 (
		\P1_reg3_reg[7]/NET0131 ,
		_w718_,
		_w719_
	);
	LUT2 #(
		.INIT('h8)
	) name258 (
		\P1_reg3_reg[8]/NET0131 ,
		_w719_,
		_w720_
	);
	LUT2 #(
		.INIT('h8)
	) name259 (
		\P1_reg3_reg[9]/NET0131 ,
		_w720_,
		_w721_
	);
	LUT2 #(
		.INIT('h8)
	) name260 (
		\P1_reg3_reg[10]/NET0131 ,
		_w721_,
		_w722_
	);
	LUT2 #(
		.INIT('h8)
	) name261 (
		\P1_reg3_reg[11]/NET0131 ,
		_w722_,
		_w723_
	);
	LUT2 #(
		.INIT('h8)
	) name262 (
		\P1_reg3_reg[12]/NET0131 ,
		\P1_reg3_reg[13]/NET0131 ,
		_w724_
	);
	LUT2 #(
		.INIT('h8)
	) name263 (
		_w723_,
		_w724_,
		_w725_
	);
	LUT2 #(
		.INIT('h8)
	) name264 (
		\P1_reg3_reg[14]/NET0131 ,
		\P1_reg3_reg[15]/NET0131 ,
		_w726_
	);
	LUT2 #(
		.INIT('h8)
	) name265 (
		\P1_reg3_reg[16]/NET0131 ,
		_w726_,
		_w727_
	);
	LUT2 #(
		.INIT('h8)
	) name266 (
		_w725_,
		_w727_,
		_w728_
	);
	LUT2 #(
		.INIT('h8)
	) name267 (
		\P1_reg3_reg[20]/NET0131 ,
		\P1_reg3_reg[21]/NET0131 ,
		_w729_
	);
	LUT2 #(
		.INIT('h8)
	) name268 (
		\P1_reg3_reg[17]/NET0131 ,
		\P1_reg3_reg[18]/NET0131 ,
		_w730_
	);
	LUT2 #(
		.INIT('h8)
	) name269 (
		\P1_reg3_reg[19]/NET0131 ,
		\P1_reg3_reg[22]/NET0131 ,
		_w731_
	);
	LUT2 #(
		.INIT('h8)
	) name270 (
		\P1_reg3_reg[23]/NET0131 ,
		\P1_reg3_reg[24]/NET0131 ,
		_w732_
	);
	LUT2 #(
		.INIT('h8)
	) name271 (
		_w731_,
		_w732_,
		_w733_
	);
	LUT2 #(
		.INIT('h8)
	) name272 (
		_w729_,
		_w730_,
		_w734_
	);
	LUT2 #(
		.INIT('h8)
	) name273 (
		_w733_,
		_w734_,
		_w735_
	);
	LUT2 #(
		.INIT('h8)
	) name274 (
		_w728_,
		_w735_,
		_w736_
	);
	LUT2 #(
		.INIT('h8)
	) name275 (
		\P1_reg3_reg[25]/NET0131 ,
		\P1_reg3_reg[26]/NET0131 ,
		_w737_
	);
	LUT2 #(
		.INIT('h8)
	) name276 (
		\P1_reg3_reg[27]/NET0131 ,
		\P1_reg3_reg[28]/NET0131 ,
		_w738_
	);
	LUT2 #(
		.INIT('h8)
	) name277 (
		_w737_,
		_w738_,
		_w739_
	);
	LUT2 #(
		.INIT('h8)
	) name278 (
		_w736_,
		_w739_,
		_w740_
	);
	LUT2 #(
		.INIT('h8)
	) name279 (
		_w715_,
		_w740_,
		_w741_
	);
	LUT2 #(
		.INIT('h2)
	) name280 (
		_w704_,
		_w714_,
		_w742_
	);
	LUT2 #(
		.INIT('h8)
	) name281 (
		\P1_reg2_reg[31]/NET0131 ,
		_w742_,
		_w743_
	);
	LUT2 #(
		.INIT('h1)
	) name282 (
		_w704_,
		_w714_,
		_w744_
	);
	LUT2 #(
		.INIT('h8)
	) name283 (
		\P1_reg0_reg[31]/NET0131 ,
		_w744_,
		_w745_
	);
	LUT2 #(
		.INIT('h4)
	) name284 (
		_w704_,
		_w714_,
		_w746_
	);
	LUT2 #(
		.INIT('h8)
	) name285 (
		\P1_reg1_reg[31]/NET0131 ,
		_w746_,
		_w747_
	);
	LUT2 #(
		.INIT('h1)
	) name286 (
		_w741_,
		_w743_,
		_w748_
	);
	LUT2 #(
		.INIT('h1)
	) name287 (
		_w745_,
		_w747_,
		_w749_
	);
	LUT2 #(
		.INIT('h8)
	) name288 (
		_w748_,
		_w749_,
		_w750_
	);
	LUT2 #(
		.INIT('h8)
	) name289 (
		\P2_datao_reg[30]/NET0131 ,
		_w543_,
		_w751_
	);
	LUT2 #(
		.INIT('h1)
	) name290 (
		_w646_,
		_w681_,
		_w752_
	);
	LUT2 #(
		.INIT('h4)
	) name291 (
		_w647_,
		_w664_,
		_w753_
	);
	LUT2 #(
		.INIT('h2)
	) name292 (
		_w651_,
		_w653_,
		_w754_
	);
	LUT2 #(
		.INIT('h1)
	) name293 (
		_w671_,
		_w674_,
		_w755_
	);
	LUT2 #(
		.INIT('h1)
	) name294 (
		_w654_,
		_w755_,
		_w756_
	);
	LUT2 #(
		.INIT('h1)
	) name295 (
		_w654_,
		_w656_,
		_w757_
	);
	LUT2 #(
		.INIT('h1)
	) name296 (
		_w545_,
		_w675_,
		_w758_
	);
	LUT2 #(
		.INIT('h1)
	) name297 (
		_w657_,
		_w758_,
		_w759_
	);
	LUT2 #(
		.INIT('h8)
	) name298 (
		_w757_,
		_w759_,
		_w760_
	);
	LUT2 #(
		.INIT('h1)
	) name299 (
		_w756_,
		_w760_,
		_w761_
	);
	LUT2 #(
		.INIT('h2)
	) name300 (
		_w754_,
		_w761_,
		_w762_
	);
	LUT2 #(
		.INIT('h1)
	) name301 (
		_w663_,
		_w670_,
		_w763_
	);
	LUT2 #(
		.INIT('h2)
	) name302 (
		_w651_,
		_w763_,
		_w764_
	);
	LUT2 #(
		.INIT('h1)
	) name303 (
		_w544_,
		_w657_,
		_w765_
	);
	LUT2 #(
		.INIT('h8)
	) name304 (
		_w757_,
		_w765_,
		_w766_
	);
	LUT2 #(
		.INIT('h1)
	) name305 (
		_w546_,
		_w552_,
		_w767_
	);
	LUT2 #(
		.INIT('h1)
	) name306 (
		_w549_,
		_w767_,
		_w768_
	);
	LUT2 #(
		.INIT('h1)
	) name307 (
		_w549_,
		_w551_,
		_w769_
	);
	LUT2 #(
		.INIT('h1)
	) name308 (
		_w553_,
		_w562_,
		_w770_
	);
	LUT2 #(
		.INIT('h1)
	) name309 (
		_w558_,
		_w770_,
		_w771_
	);
	LUT2 #(
		.INIT('h8)
	) name310 (
		_w769_,
		_w771_,
		_w772_
	);
	LUT2 #(
		.INIT('h1)
	) name311 (
		_w768_,
		_w772_,
		_w773_
	);
	LUT2 #(
		.INIT('h1)
	) name312 (
		_w577_,
		_w583_,
		_w774_
	);
	LUT2 #(
		.INIT('h1)
	) name313 (
		_w584_,
		_w599_,
		_w775_
	);
	LUT2 #(
		.INIT('h2)
	) name314 (
		_w635_,
		_w775_,
		_w776_
	);
	LUT2 #(
		.INIT('h2)
	) name315 (
		_w774_,
		_w776_,
		_w777_
	);
	LUT2 #(
		.INIT('h1)
	) name316 (
		_w580_,
		_w777_,
		_w778_
	);
	LUT2 #(
		.INIT('h1)
	) name317 (
		_w614_,
		_w615_,
		_w779_
	);
	LUT2 #(
		.INIT('h2)
	) name318 (
		_w611_,
		_w779_,
		_w780_
	);
	LUT2 #(
		.INIT('h4)
	) name319 (
		_w609_,
		_w616_,
		_w781_
	);
	LUT2 #(
		.INIT('h1)
	) name320 (
		_w608_,
		_w781_,
		_w782_
	);
	LUT2 #(
		.INIT('h4)
	) name321 (
		_w780_,
		_w782_,
		_w783_
	);
	LUT2 #(
		.INIT('h2)
	) name322 (
		_w624_,
		_w783_,
		_w784_
	);
	LUT2 #(
		.INIT('h1)
	) name323 (
		_w603_,
		_w607_,
		_w785_
	);
	LUT2 #(
		.INIT('h1)
	) name324 (
		_w622_,
		_w785_,
		_w786_
	);
	LUT2 #(
		.INIT('h1)
	) name325 (
		_w784_,
		_w786_,
		_w787_
	);
	LUT2 #(
		.INIT('h4)
	) name326 (
		_w592_,
		_w629_,
		_w788_
	);
	LUT2 #(
		.INIT('h4)
	) name327 (
		_w602_,
		_w788_,
		_w789_
	);
	LUT2 #(
		.INIT('h4)
	) name328 (
		_w787_,
		_w789_,
		_w790_
	);
	LUT2 #(
		.INIT('h1)
	) name329 (
		_w589_,
		_w598_,
		_w791_
	);
	LUT2 #(
		.INIT('h1)
	) name330 (
		_w592_,
		_w791_,
		_w792_
	);
	LUT2 #(
		.INIT('h1)
	) name331 (
		_w590_,
		_w604_,
		_w793_
	);
	LUT2 #(
		.INIT('h2)
	) name332 (
		_w788_,
		_w793_,
		_w794_
	);
	LUT2 #(
		.INIT('h1)
	) name333 (
		_w792_,
		_w794_,
		_w795_
	);
	LUT2 #(
		.INIT('h4)
	) name334 (
		_w790_,
		_w795_,
		_w796_
	);
	LUT2 #(
		.INIT('h1)
	) name335 (
		_w580_,
		_w593_,
		_w797_
	);
	LUT2 #(
		.INIT('h8)
	) name336 (
		_w635_,
		_w797_,
		_w798_
	);
	LUT2 #(
		.INIT('h4)
	) name337 (
		_w796_,
		_w798_,
		_w799_
	);
	LUT2 #(
		.INIT('h1)
	) name338 (
		_w778_,
		_w799_,
		_w800_
	);
	LUT2 #(
		.INIT('h1)
	) name339 (
		_w566_,
		_w575_,
		_w801_
	);
	LUT2 #(
		.INIT('h8)
	) name340 (
		_w640_,
		_w801_,
		_w802_
	);
	LUT2 #(
		.INIT('h4)
	) name341 (
		_w800_,
		_w802_,
		_w803_
	);
	LUT2 #(
		.INIT('h1)
	) name342 (
		_w563_,
		_w570_,
		_w804_
	);
	LUT2 #(
		.INIT('h1)
	) name343 (
		_w569_,
		_w576_,
		_w805_
	);
	LUT2 #(
		.INIT('h2)
	) name344 (
		_w640_,
		_w805_,
		_w806_
	);
	LUT2 #(
		.INIT('h2)
	) name345 (
		_w804_,
		_w806_,
		_w807_
	);
	LUT2 #(
		.INIT('h1)
	) name346 (
		_w566_,
		_w807_,
		_w808_
	);
	LUT2 #(
		.INIT('h1)
	) name347 (
		_w803_,
		_w808_,
		_w809_
	);
	LUT2 #(
		.INIT('h1)
	) name348 (
		_w558_,
		_w561_,
		_w810_
	);
	LUT2 #(
		.INIT('h8)
	) name349 (
		_w769_,
		_w810_,
		_w811_
	);
	LUT2 #(
		.INIT('h4)
	) name350 (
		_w809_,
		_w811_,
		_w812_
	);
	LUT2 #(
		.INIT('h2)
	) name351 (
		_w773_,
		_w812_,
		_w813_
	);
	LUT2 #(
		.INIT('h8)
	) name352 (
		_w754_,
		_w766_,
		_w814_
	);
	LUT2 #(
		.INIT('h4)
	) name353 (
		_w813_,
		_w814_,
		_w815_
	);
	LUT2 #(
		.INIT('h1)
	) name354 (
		_w662_,
		_w753_,
		_w816_
	);
	LUT2 #(
		.INIT('h4)
	) name355 (
		_w764_,
		_w816_,
		_w817_
	);
	LUT2 #(
		.INIT('h4)
	) name356 (
		_w762_,
		_w817_,
		_w818_
	);
	LUT2 #(
		.INIT('h4)
	) name357 (
		_w815_,
		_w818_,
		_w819_
	);
	LUT2 #(
		.INIT('h2)
	) name358 (
		_w752_,
		_w819_,
		_w820_
	);
	LUT2 #(
		.INIT('h4)
	) name359 (
		_w752_,
		_w819_,
		_w821_
	);
	LUT2 #(
		.INIT('h1)
	) name360 (
		_w543_,
		_w820_,
		_w822_
	);
	LUT2 #(
		.INIT('h4)
	) name361 (
		_w821_,
		_w822_,
		_w823_
	);
	LUT2 #(
		.INIT('h1)
	) name362 (
		_w751_,
		_w823_,
		_w824_
	);
	LUT2 #(
		.INIT('h1)
	) name363 (
		_w538_,
		_w824_,
		_w825_
	);
	LUT2 #(
		.INIT('h8)
	) name364 (
		\P1_reg2_reg[30]/NET0131 ,
		_w742_,
		_w826_
	);
	LUT2 #(
		.INIT('h8)
	) name365 (
		\P1_reg0_reg[30]/NET0131 ,
		_w744_,
		_w827_
	);
	LUT2 #(
		.INIT('h8)
	) name366 (
		\P1_reg1_reg[30]/NET0131 ,
		_w746_,
		_w828_
	);
	LUT2 #(
		.INIT('h1)
	) name367 (
		_w741_,
		_w826_,
		_w829_
	);
	LUT2 #(
		.INIT('h1)
	) name368 (
		_w827_,
		_w828_,
		_w830_
	);
	LUT2 #(
		.INIT('h8)
	) name369 (
		_w829_,
		_w830_,
		_w831_
	);
	LUT2 #(
		.INIT('h1)
	) name370 (
		_w825_,
		_w831_,
		_w832_
	);
	LUT2 #(
		.INIT('h1)
	) name371 (
		_w750_,
		_w832_,
		_w833_
	);
	LUT2 #(
		.INIT('h2)
	) name372 (
		_w692_,
		_w833_,
		_w834_
	);
	LUT2 #(
		.INIT('h1)
	) name373 (
		_w692_,
		_w750_,
		_w835_
	);
	LUT2 #(
		.INIT('h1)
	) name374 (
		_w750_,
		_w831_,
		_w836_
	);
	LUT2 #(
		.INIT('h2)
	) name375 (
		_w825_,
		_w836_,
		_w837_
	);
	LUT2 #(
		.INIT('h8)
	) name376 (
		\P2_datao_reg[29]/NET0131 ,
		_w543_,
		_w838_
	);
	LUT2 #(
		.INIT('h1)
	) name377 (
		_w647_,
		_w662_,
		_w839_
	);
	LUT2 #(
		.INIT('h8)
	) name378 (
		_w548_,
		_w658_,
		_w840_
	);
	LUT2 #(
		.INIT('h1)
	) name379 (
		_w677_,
		_w840_,
		_w841_
	);
	LUT2 #(
		.INIT('h2)
	) name380 (
		_w655_,
		_w841_,
		_w842_
	);
	LUT2 #(
		.INIT('h1)
	) name381 (
		_w673_,
		_w842_,
		_w843_
	);
	LUT2 #(
		.INIT('h1)
	) name382 (
		_w648_,
		_w843_,
		_w844_
	);
	LUT2 #(
		.INIT('h2)
	) name383 (
		_w665_,
		_w844_,
		_w845_
	);
	LUT2 #(
		.INIT('h1)
	) name384 (
		_w649_,
		_w845_,
		_w846_
	);
	LUT2 #(
		.INIT('h8)
	) name385 (
		_w559_,
		_w565_,
		_w847_
	);
	LUT2 #(
		.INIT('h1)
	) name386 (
		_w555_,
		_w847_,
		_w848_
	);
	LUT2 #(
		.INIT('h8)
	) name387 (
		_w579_,
		_w640_,
		_w849_
	);
	LUT2 #(
		.INIT('h1)
	) name388 (
		_w572_,
		_w849_,
		_w850_
	);
	LUT2 #(
		.INIT('h1)
	) name389 (
		_w590_,
		_w606_,
		_w851_
	);
	LUT2 #(
		.INIT('h2)
	) name390 (
		_w629_,
		_w851_,
		_w852_
	);
	LUT2 #(
		.INIT('h1)
	) name391 (
		_w620_,
		_w623_,
		_w853_
	);
	LUT2 #(
		.INIT('h1)
	) name392 (
		_w607_,
		_w853_,
		_w854_
	);
	LUT2 #(
		.INIT('h1)
	) name393 (
		_w602_,
		_w628_,
		_w855_
	);
	LUT2 #(
		.INIT('h1)
	) name394 (
		_w595_,
		_w622_,
		_w856_
	);
	LUT2 #(
		.INIT('h8)
	) name395 (
		_w855_,
		_w856_,
		_w857_
	);
	LUT2 #(
		.INIT('h4)
	) name396 (
		_w854_,
		_w857_,
		_w858_
	);
	LUT2 #(
		.INIT('h1)
	) name397 (
		_w589_,
		_w852_,
		_w859_
	);
	LUT2 #(
		.INIT('h4)
	) name398 (
		_w858_,
		_w859_,
		_w860_
	);
	LUT2 #(
		.INIT('h8)
	) name399 (
		_w594_,
		_w635_,
		_w861_
	);
	LUT2 #(
		.INIT('h4)
	) name400 (
		_w860_,
		_w861_,
		_w862_
	);
	LUT2 #(
		.INIT('h8)
	) name401 (
		_w601_,
		_w635_,
		_w863_
	);
	LUT2 #(
		.INIT('h1)
	) name402 (
		_w586_,
		_w863_,
		_w864_
	);
	LUT2 #(
		.INIT('h4)
	) name403 (
		_w862_,
		_w864_,
		_w865_
	);
	LUT2 #(
		.INIT('h8)
	) name404 (
		_w581_,
		_w640_,
		_w866_
	);
	LUT2 #(
		.INIT('h4)
	) name405 (
		_w865_,
		_w866_,
		_w867_
	);
	LUT2 #(
		.INIT('h2)
	) name406 (
		_w850_,
		_w867_,
		_w868_
	);
	LUT2 #(
		.INIT('h8)
	) name407 (
		_w559_,
		_w567_,
		_w869_
	);
	LUT2 #(
		.INIT('h4)
	) name408 (
		_w868_,
		_w869_,
		_w870_
	);
	LUT2 #(
		.INIT('h2)
	) name409 (
		_w848_,
		_w870_,
		_w871_
	);
	LUT2 #(
		.INIT('h8)
	) name410 (
		_w550_,
		_w659_,
		_w872_
	);
	LUT2 #(
		.INIT('h8)
	) name411 (
		_w650_,
		_w872_,
		_w873_
	);
	LUT2 #(
		.INIT('h4)
	) name412 (
		_w871_,
		_w873_,
		_w874_
	);
	LUT2 #(
		.INIT('h1)
	) name413 (
		_w846_,
		_w874_,
		_w875_
	);
	LUT2 #(
		.INIT('h2)
	) name414 (
		_w839_,
		_w875_,
		_w876_
	);
	LUT2 #(
		.INIT('h4)
	) name415 (
		_w839_,
		_w875_,
		_w877_
	);
	LUT2 #(
		.INIT('h1)
	) name416 (
		_w543_,
		_w876_,
		_w878_
	);
	LUT2 #(
		.INIT('h4)
	) name417 (
		_w877_,
		_w878_,
		_w879_
	);
	LUT2 #(
		.INIT('h1)
	) name418 (
		_w838_,
		_w879_,
		_w880_
	);
	LUT2 #(
		.INIT('h1)
	) name419 (
		_w538_,
		_w880_,
		_w881_
	);
	LUT2 #(
		.INIT('h8)
	) name420 (
		\P1_reg1_reg[29]/NET0131 ,
		_w746_,
		_w882_
	);
	LUT2 #(
		.INIT('h8)
	) name421 (
		\P1_reg0_reg[29]/NET0131 ,
		_w744_,
		_w883_
	);
	LUT2 #(
		.INIT('h8)
	) name422 (
		\P1_reg2_reg[29]/NET0131 ,
		_w742_,
		_w884_
	);
	LUT2 #(
		.INIT('h1)
	) name423 (
		_w741_,
		_w882_,
		_w885_
	);
	LUT2 #(
		.INIT('h1)
	) name424 (
		_w883_,
		_w884_,
		_w886_
	);
	LUT2 #(
		.INIT('h8)
	) name425 (
		_w885_,
		_w886_,
		_w887_
	);
	LUT2 #(
		.INIT('h8)
	) name426 (
		_w881_,
		_w887_,
		_w888_
	);
	LUT2 #(
		.INIT('h8)
	) name427 (
		\P2_datao_reg[28]/NET0131 ,
		_w543_,
		_w889_
	);
	LUT2 #(
		.INIT('h1)
	) name428 (
		_w649_,
		_w664_,
		_w890_
	);
	LUT2 #(
		.INIT('h4)
	) name429 (
		_w653_,
		_w756_,
		_w891_
	);
	LUT2 #(
		.INIT('h2)
	) name430 (
		_w763_,
		_w891_,
		_w892_
	);
	LUT2 #(
		.INIT('h1)
	) name431 (
		_w648_,
		_w892_,
		_w893_
	);
	LUT2 #(
		.INIT('h1)
	) name432 (
		_w599_,
		_w792_,
		_w894_
	);
	LUT2 #(
		.INIT('h1)
	) name433 (
		_w593_,
		_w634_,
		_w895_
	);
	LUT2 #(
		.INIT('h4)
	) name434 (
		_w894_,
		_w895_,
		_w896_
	);
	LUT2 #(
		.INIT('h1)
	) name435 (
		_w584_,
		_w896_,
		_w897_
	);
	LUT2 #(
		.INIT('h1)
	) name436 (
		_w582_,
		_w897_,
		_w898_
	);
	LUT2 #(
		.INIT('h2)
	) name437 (
		_w774_,
		_w898_,
		_w899_
	);
	LUT2 #(
		.INIT('h2)
	) name438 (
		_w581_,
		_w899_,
		_w900_
	);
	LUT2 #(
		.INIT('h2)
	) name439 (
		_w805_,
		_w900_,
		_w901_
	);
	LUT2 #(
		.INIT('h1)
	) name440 (
		_w639_,
		_w901_,
		_w902_
	);
	LUT2 #(
		.INIT('h1)
	) name441 (
		_w604_,
		_w786_,
		_w903_
	);
	LUT2 #(
		.INIT('h4)
	) name442 (
		_w784_,
		_w903_,
		_w904_
	);
	LUT2 #(
		.INIT('h2)
	) name443 (
		_w855_,
		_w904_,
		_w905_
	);
	LUT2 #(
		.INIT('h1)
	) name444 (
		_w590_,
		_w905_,
		_w906_
	);
	LUT2 #(
		.INIT('h2)
	) name445 (
		_w596_,
		_w634_,
		_w907_
	);
	LUT2 #(
		.INIT('h4)
	) name446 (
		_w906_,
		_w907_,
		_w908_
	);
	LUT2 #(
		.INIT('h1)
	) name447 (
		_w582_,
		_w639_,
		_w909_
	);
	LUT2 #(
		.INIT('h8)
	) name448 (
		_w581_,
		_w909_,
		_w910_
	);
	LUT2 #(
		.INIT('h8)
	) name449 (
		_w908_,
		_w910_,
		_w911_
	);
	LUT2 #(
		.INIT('h1)
	) name450 (
		_w902_,
		_w911_,
		_w912_
	);
	LUT2 #(
		.INIT('h4)
	) name451 (
		_w558_,
		_w567_,
		_w913_
	);
	LUT2 #(
		.INIT('h4)
	) name452 (
		_w568_,
		_w913_,
		_w914_
	);
	LUT2 #(
		.INIT('h4)
	) name453 (
		_w912_,
		_w914_,
		_w915_
	);
	LUT2 #(
		.INIT('h4)
	) name454 (
		_w804_,
		_w913_,
		_w916_
	);
	LUT2 #(
		.INIT('h1)
	) name455 (
		_w771_,
		_w916_,
		_w917_
	);
	LUT2 #(
		.INIT('h4)
	) name456 (
		_w915_,
		_w917_,
		_w918_
	);
	LUT2 #(
		.INIT('h8)
	) name457 (
		_w765_,
		_w769_,
		_w919_
	);
	LUT2 #(
		.INIT('h4)
	) name458 (
		_w918_,
		_w919_,
		_w920_
	);
	LUT2 #(
		.INIT('h8)
	) name459 (
		_w765_,
		_w768_,
		_w921_
	);
	LUT2 #(
		.INIT('h1)
	) name460 (
		_w759_,
		_w921_,
		_w922_
	);
	LUT2 #(
		.INIT('h4)
	) name461 (
		_w920_,
		_w922_,
		_w923_
	);
	LUT2 #(
		.INIT('h1)
	) name462 (
		_w648_,
		_w656_,
		_w924_
	);
	LUT2 #(
		.INIT('h8)
	) name463 (
		_w655_,
		_w924_,
		_w925_
	);
	LUT2 #(
		.INIT('h4)
	) name464 (
		_w923_,
		_w925_,
		_w926_
	);
	LUT2 #(
		.INIT('h1)
	) name465 (
		_w893_,
		_w926_,
		_w927_
	);
	LUT2 #(
		.INIT('h2)
	) name466 (
		_w890_,
		_w927_,
		_w928_
	);
	LUT2 #(
		.INIT('h4)
	) name467 (
		_w890_,
		_w927_,
		_w929_
	);
	LUT2 #(
		.INIT('h1)
	) name468 (
		_w543_,
		_w928_,
		_w930_
	);
	LUT2 #(
		.INIT('h4)
	) name469 (
		_w929_,
		_w930_,
		_w931_
	);
	LUT2 #(
		.INIT('h1)
	) name470 (
		_w889_,
		_w931_,
		_w932_
	);
	LUT2 #(
		.INIT('h1)
	) name471 (
		_w538_,
		_w932_,
		_w933_
	);
	LUT2 #(
		.INIT('h8)
	) name472 (
		\P1_reg0_reg[28]/NET0131 ,
		_w744_,
		_w934_
	);
	LUT2 #(
		.INIT('h8)
	) name473 (
		\P1_reg1_reg[28]/NET0131 ,
		_w746_,
		_w935_
	);
	LUT2 #(
		.INIT('h8)
	) name474 (
		\P1_reg2_reg[28]/NET0131 ,
		_w742_,
		_w936_
	);
	LUT2 #(
		.INIT('h8)
	) name475 (
		\P1_reg3_reg[25]/NET0131 ,
		_w736_,
		_w937_
	);
	LUT2 #(
		.INIT('h8)
	) name476 (
		\P1_reg3_reg[26]/NET0131 ,
		_w937_,
		_w938_
	);
	LUT2 #(
		.INIT('h8)
	) name477 (
		\P1_reg3_reg[27]/NET0131 ,
		_w938_,
		_w939_
	);
	LUT2 #(
		.INIT('h1)
	) name478 (
		\P1_reg3_reg[28]/NET0131 ,
		_w939_,
		_w940_
	);
	LUT2 #(
		.INIT('h1)
	) name479 (
		_w740_,
		_w940_,
		_w941_
	);
	LUT2 #(
		.INIT('h8)
	) name480 (
		_w715_,
		_w941_,
		_w942_
	);
	LUT2 #(
		.INIT('h1)
	) name481 (
		_w934_,
		_w935_,
		_w943_
	);
	LUT2 #(
		.INIT('h4)
	) name482 (
		_w936_,
		_w943_,
		_w944_
	);
	LUT2 #(
		.INIT('h4)
	) name483 (
		_w942_,
		_w944_,
		_w945_
	);
	LUT2 #(
		.INIT('h1)
	) name484 (
		_w933_,
		_w945_,
		_w946_
	);
	LUT2 #(
		.INIT('h1)
	) name485 (
		_w881_,
		_w887_,
		_w947_
	);
	LUT2 #(
		.INIT('h1)
	) name486 (
		_w946_,
		_w947_,
		_w948_
	);
	LUT2 #(
		.INIT('h1)
	) name487 (
		_w888_,
		_w948_,
		_w949_
	);
	LUT2 #(
		.INIT('h8)
	) name488 (
		_w933_,
		_w945_,
		_w950_
	);
	LUT2 #(
		.INIT('h1)
	) name489 (
		_w888_,
		_w950_,
		_w951_
	);
	LUT2 #(
		.INIT('h8)
	) name490 (
		\P2_datao_reg[27]/NET0131 ,
		_w543_,
		_w952_
	);
	LUT2 #(
		.INIT('h1)
	) name491 (
		_w648_,
		_w663_,
		_w953_
	);
	LUT2 #(
		.INIT('h4)
	) name492 (
		_w588_,
		_w641_,
		_w954_
	);
	LUT2 #(
		.INIT('h2)
	) name493 (
		_w574_,
		_w954_,
		_w955_
	);
	LUT2 #(
		.INIT('h2)
	) name494 (
		_w560_,
		_w955_,
		_w956_
	);
	LUT2 #(
		.INIT('h2)
	) name495 (
		_w557_,
		_w956_,
		_w957_
	);
	LUT2 #(
		.INIT('h2)
	) name496 (
		_w659_,
		_w957_,
		_w958_
	);
	LUT2 #(
		.INIT('h8)
	) name497 (
		_w559_,
		_w641_,
		_w959_
	);
	LUT2 #(
		.INIT('h8)
	) name498 (
		_w872_,
		_w959_,
		_w960_
	);
	LUT2 #(
		.INIT('h8)
	) name499 (
		_w637_,
		_w960_,
		_w961_
	);
	LUT2 #(
		.INIT('h2)
	) name500 (
		_w679_,
		_w958_,
		_w962_
	);
	LUT2 #(
		.INIT('h4)
	) name501 (
		_w961_,
		_w962_,
		_w963_
	);
	LUT2 #(
		.INIT('h2)
	) name502 (
		_w953_,
		_w963_,
		_w964_
	);
	LUT2 #(
		.INIT('h4)
	) name503 (
		_w953_,
		_w963_,
		_w965_
	);
	LUT2 #(
		.INIT('h1)
	) name504 (
		_w543_,
		_w964_,
		_w966_
	);
	LUT2 #(
		.INIT('h4)
	) name505 (
		_w965_,
		_w966_,
		_w967_
	);
	LUT2 #(
		.INIT('h1)
	) name506 (
		_w952_,
		_w967_,
		_w968_
	);
	LUT2 #(
		.INIT('h1)
	) name507 (
		_w538_,
		_w968_,
		_w969_
	);
	LUT2 #(
		.INIT('h8)
	) name508 (
		\P1_reg0_reg[27]/NET0131 ,
		_w744_,
		_w970_
	);
	LUT2 #(
		.INIT('h8)
	) name509 (
		\P1_reg2_reg[27]/NET0131 ,
		_w742_,
		_w971_
	);
	LUT2 #(
		.INIT('h8)
	) name510 (
		\P1_reg1_reg[27]/NET0131 ,
		_w746_,
		_w972_
	);
	LUT2 #(
		.INIT('h1)
	) name511 (
		\P1_reg3_reg[27]/NET0131 ,
		_w938_,
		_w973_
	);
	LUT2 #(
		.INIT('h1)
	) name512 (
		_w939_,
		_w973_,
		_w974_
	);
	LUT2 #(
		.INIT('h8)
	) name513 (
		_w715_,
		_w974_,
		_w975_
	);
	LUT2 #(
		.INIT('h1)
	) name514 (
		_w970_,
		_w971_,
		_w976_
	);
	LUT2 #(
		.INIT('h4)
	) name515 (
		_w972_,
		_w976_,
		_w977_
	);
	LUT2 #(
		.INIT('h4)
	) name516 (
		_w975_,
		_w977_,
		_w978_
	);
	LUT2 #(
		.INIT('h8)
	) name517 (
		_w969_,
		_w978_,
		_w979_
	);
	LUT2 #(
		.INIT('h8)
	) name518 (
		\P2_datao_reg[26]/NET0131 ,
		_w543_,
		_w980_
	);
	LUT2 #(
		.INIT('h1)
	) name519 (
		_w653_,
		_w670_,
		_w981_
	);
	LUT2 #(
		.INIT('h8)
	) name520 (
		_w778_,
		_w802_,
		_w982_
	);
	LUT2 #(
		.INIT('h1)
	) name521 (
		_w808_,
		_w982_,
		_w983_
	);
	LUT2 #(
		.INIT('h2)
	) name522 (
		_w811_,
		_w983_,
		_w984_
	);
	LUT2 #(
		.INIT('h2)
	) name523 (
		_w773_,
		_w984_,
		_w985_
	);
	LUT2 #(
		.INIT('h2)
	) name524 (
		_w766_,
		_w985_,
		_w986_
	);
	LUT2 #(
		.INIT('h8)
	) name525 (
		_w766_,
		_w802_,
		_w987_
	);
	LUT2 #(
		.INIT('h8)
	) name526 (
		_w811_,
		_w987_,
		_w988_
	);
	LUT2 #(
		.INIT('h8)
	) name527 (
		_w799_,
		_w988_,
		_w989_
	);
	LUT2 #(
		.INIT('h2)
	) name528 (
		_w761_,
		_w986_,
		_w990_
	);
	LUT2 #(
		.INIT('h4)
	) name529 (
		_w989_,
		_w990_,
		_w991_
	);
	LUT2 #(
		.INIT('h2)
	) name530 (
		_w981_,
		_w991_,
		_w992_
	);
	LUT2 #(
		.INIT('h4)
	) name531 (
		_w981_,
		_w991_,
		_w993_
	);
	LUT2 #(
		.INIT('h1)
	) name532 (
		_w543_,
		_w992_,
		_w994_
	);
	LUT2 #(
		.INIT('h4)
	) name533 (
		_w993_,
		_w994_,
		_w995_
	);
	LUT2 #(
		.INIT('h1)
	) name534 (
		_w980_,
		_w995_,
		_w996_
	);
	LUT2 #(
		.INIT('h1)
	) name535 (
		_w538_,
		_w996_,
		_w997_
	);
	LUT2 #(
		.INIT('h8)
	) name536 (
		\P1_reg1_reg[26]/NET0131 ,
		_w746_,
		_w998_
	);
	LUT2 #(
		.INIT('h8)
	) name537 (
		\P1_reg2_reg[26]/NET0131 ,
		_w742_,
		_w999_
	);
	LUT2 #(
		.INIT('h8)
	) name538 (
		\P1_reg0_reg[26]/NET0131 ,
		_w744_,
		_w1000_
	);
	LUT2 #(
		.INIT('h1)
	) name539 (
		\P1_reg3_reg[26]/NET0131 ,
		_w937_,
		_w1001_
	);
	LUT2 #(
		.INIT('h1)
	) name540 (
		_w938_,
		_w1001_,
		_w1002_
	);
	LUT2 #(
		.INIT('h8)
	) name541 (
		_w715_,
		_w1002_,
		_w1003_
	);
	LUT2 #(
		.INIT('h1)
	) name542 (
		_w998_,
		_w999_,
		_w1004_
	);
	LUT2 #(
		.INIT('h4)
	) name543 (
		_w1000_,
		_w1004_,
		_w1005_
	);
	LUT2 #(
		.INIT('h4)
	) name544 (
		_w1003_,
		_w1005_,
		_w1006_
	);
	LUT2 #(
		.INIT('h1)
	) name545 (
		_w997_,
		_w1006_,
		_w1007_
	);
	LUT2 #(
		.INIT('h1)
	) name546 (
		_w969_,
		_w978_,
		_w1008_
	);
	LUT2 #(
		.INIT('h1)
	) name547 (
		_w1007_,
		_w1008_,
		_w1009_
	);
	LUT2 #(
		.INIT('h8)
	) name548 (
		_w997_,
		_w1006_,
		_w1010_
	);
	LUT2 #(
		.INIT('h8)
	) name549 (
		\P2_datao_reg[25]/NET0131 ,
		_w543_,
		_w1011_
	);
	LUT2 #(
		.INIT('h1)
	) name550 (
		_w654_,
		_w671_,
		_w1012_
	);
	LUT2 #(
		.INIT('h8)
	) name551 (
		_w550_,
		_w658_,
		_w1013_
	);
	LUT2 #(
		.INIT('h4)
	) name552 (
		_w864_,
		_w866_,
		_w1014_
	);
	LUT2 #(
		.INIT('h2)
	) name553 (
		_w850_,
		_w1014_,
		_w1015_
	);
	LUT2 #(
		.INIT('h2)
	) name554 (
		_w869_,
		_w1015_,
		_w1016_
	);
	LUT2 #(
		.INIT('h2)
	) name555 (
		_w848_,
		_w1016_,
		_w1017_
	);
	LUT2 #(
		.INIT('h2)
	) name556 (
		_w1013_,
		_w1017_,
		_w1018_
	);
	LUT2 #(
		.INIT('h8)
	) name557 (
		_w866_,
		_w869_,
		_w1019_
	);
	LUT2 #(
		.INIT('h8)
	) name558 (
		_w1013_,
		_w1019_,
		_w1020_
	);
	LUT2 #(
		.INIT('h8)
	) name559 (
		_w862_,
		_w1020_,
		_w1021_
	);
	LUT2 #(
		.INIT('h2)
	) name560 (
		_w841_,
		_w1018_,
		_w1022_
	);
	LUT2 #(
		.INIT('h4)
	) name561 (
		_w1021_,
		_w1022_,
		_w1023_
	);
	LUT2 #(
		.INIT('h2)
	) name562 (
		_w1012_,
		_w1023_,
		_w1024_
	);
	LUT2 #(
		.INIT('h4)
	) name563 (
		_w1012_,
		_w1023_,
		_w1025_
	);
	LUT2 #(
		.INIT('h1)
	) name564 (
		_w543_,
		_w1024_,
		_w1026_
	);
	LUT2 #(
		.INIT('h4)
	) name565 (
		_w1025_,
		_w1026_,
		_w1027_
	);
	LUT2 #(
		.INIT('h1)
	) name566 (
		_w1011_,
		_w1027_,
		_w1028_
	);
	LUT2 #(
		.INIT('h1)
	) name567 (
		_w538_,
		_w1028_,
		_w1029_
	);
	LUT2 #(
		.INIT('h8)
	) name568 (
		\P1_reg2_reg[25]/NET0131 ,
		_w742_,
		_w1030_
	);
	LUT2 #(
		.INIT('h8)
	) name569 (
		\P1_reg1_reg[25]/NET0131 ,
		_w746_,
		_w1031_
	);
	LUT2 #(
		.INIT('h8)
	) name570 (
		\P1_reg0_reg[25]/NET0131 ,
		_w744_,
		_w1032_
	);
	LUT2 #(
		.INIT('h1)
	) name571 (
		\P1_reg3_reg[25]/NET0131 ,
		_w736_,
		_w1033_
	);
	LUT2 #(
		.INIT('h1)
	) name572 (
		_w937_,
		_w1033_,
		_w1034_
	);
	LUT2 #(
		.INIT('h8)
	) name573 (
		_w715_,
		_w1034_,
		_w1035_
	);
	LUT2 #(
		.INIT('h1)
	) name574 (
		_w1030_,
		_w1031_,
		_w1036_
	);
	LUT2 #(
		.INIT('h4)
	) name575 (
		_w1032_,
		_w1036_,
		_w1037_
	);
	LUT2 #(
		.INIT('h4)
	) name576 (
		_w1035_,
		_w1037_,
		_w1038_
	);
	LUT2 #(
		.INIT('h8)
	) name577 (
		_w1029_,
		_w1038_,
		_w1039_
	);
	LUT2 #(
		.INIT('h8)
	) name578 (
		\P2_datao_reg[24]/NET0131 ,
		_w543_,
		_w1040_
	);
	LUT2 #(
		.INIT('h1)
	) name579 (
		_w656_,
		_w674_,
		_w1041_
	);
	LUT2 #(
		.INIT('h4)
	) name580 (
		_w923_,
		_w1041_,
		_w1042_
	);
	LUT2 #(
		.INIT('h2)
	) name581 (
		_w923_,
		_w1041_,
		_w1043_
	);
	LUT2 #(
		.INIT('h1)
	) name582 (
		_w543_,
		_w1042_,
		_w1044_
	);
	LUT2 #(
		.INIT('h4)
	) name583 (
		_w1043_,
		_w1044_,
		_w1045_
	);
	LUT2 #(
		.INIT('h1)
	) name584 (
		_w1040_,
		_w1045_,
		_w1046_
	);
	LUT2 #(
		.INIT('h1)
	) name585 (
		_w538_,
		_w1046_,
		_w1047_
	);
	LUT2 #(
		.INIT('h8)
	) name586 (
		\P1_reg2_reg[24]/NET0131 ,
		_w742_,
		_w1048_
	);
	LUT2 #(
		.INIT('h8)
	) name587 (
		\P1_reg0_reg[24]/NET0131 ,
		_w744_,
		_w1049_
	);
	LUT2 #(
		.INIT('h8)
	) name588 (
		\P1_reg1_reg[24]/NET0131 ,
		_w746_,
		_w1050_
	);
	LUT2 #(
		.INIT('h8)
	) name589 (
		\P1_reg3_reg[17]/NET0131 ,
		_w728_,
		_w1051_
	);
	LUT2 #(
		.INIT('h8)
	) name590 (
		\P1_reg3_reg[18]/NET0131 ,
		_w1051_,
		_w1052_
	);
	LUT2 #(
		.INIT('h8)
	) name591 (
		\P1_reg3_reg[19]/NET0131 ,
		_w1052_,
		_w1053_
	);
	LUT2 #(
		.INIT('h8)
	) name592 (
		_w729_,
		_w1053_,
		_w1054_
	);
	LUT2 #(
		.INIT('h8)
	) name593 (
		\P1_reg3_reg[22]/NET0131 ,
		_w1054_,
		_w1055_
	);
	LUT2 #(
		.INIT('h8)
	) name594 (
		\P1_reg3_reg[23]/NET0131 ,
		_w1055_,
		_w1056_
	);
	LUT2 #(
		.INIT('h1)
	) name595 (
		\P1_reg3_reg[24]/NET0131 ,
		_w1056_,
		_w1057_
	);
	LUT2 #(
		.INIT('h1)
	) name596 (
		_w736_,
		_w1057_,
		_w1058_
	);
	LUT2 #(
		.INIT('h8)
	) name597 (
		_w715_,
		_w1058_,
		_w1059_
	);
	LUT2 #(
		.INIT('h1)
	) name598 (
		_w1048_,
		_w1049_,
		_w1060_
	);
	LUT2 #(
		.INIT('h4)
	) name599 (
		_w1050_,
		_w1060_,
		_w1061_
	);
	LUT2 #(
		.INIT('h4)
	) name600 (
		_w1059_,
		_w1061_,
		_w1062_
	);
	LUT2 #(
		.INIT('h1)
	) name601 (
		_w1047_,
		_w1062_,
		_w1063_
	);
	LUT2 #(
		.INIT('h1)
	) name602 (
		_w1029_,
		_w1038_,
		_w1064_
	);
	LUT2 #(
		.INIT('h1)
	) name603 (
		_w1063_,
		_w1064_,
		_w1065_
	);
	LUT2 #(
		.INIT('h1)
	) name604 (
		_w1039_,
		_w1065_,
		_w1066_
	);
	LUT2 #(
		.INIT('h4)
	) name605 (
		_w1010_,
		_w1066_,
		_w1067_
	);
	LUT2 #(
		.INIT('h2)
	) name606 (
		_w1009_,
		_w1067_,
		_w1068_
	);
	LUT2 #(
		.INIT('h1)
	) name607 (
		_w979_,
		_w1068_,
		_w1069_
	);
	LUT2 #(
		.INIT('h2)
	) name608 (
		\P1_IR_reg[31]/NET0131 ,
		_w503_,
		_w1070_
	);
	LUT2 #(
		.INIT('h1)
	) name609 (
		\P1_IR_reg[15]/NET0131 ,
		_w1070_,
		_w1071_
	);
	LUT2 #(
		.INIT('h8)
	) name610 (
		\P1_IR_reg[15]/NET0131 ,
		_w1070_,
		_w1072_
	);
	LUT2 #(
		.INIT('h1)
	) name611 (
		_w1071_,
		_w1072_,
		_w1073_
	);
	LUT2 #(
		.INIT('h2)
	) name612 (
		_w538_,
		_w1073_,
		_w1074_
	);
	LUT2 #(
		.INIT('h8)
	) name613 (
		\P2_datao_reg[15]/NET0131 ,
		_w543_,
		_w1075_
	);
	LUT2 #(
		.INIT('h1)
	) name614 (
		_w569_,
		_w639_,
		_w1076_
	);
	LUT2 #(
		.INIT('h4)
	) name615 (
		_w638_,
		_w1076_,
		_w1077_
	);
	LUT2 #(
		.INIT('h2)
	) name616 (
		_w638_,
		_w1076_,
		_w1078_
	);
	LUT2 #(
		.INIT('h1)
	) name617 (
		_w543_,
		_w1077_,
		_w1079_
	);
	LUT2 #(
		.INIT('h4)
	) name618 (
		_w1078_,
		_w1079_,
		_w1080_
	);
	LUT2 #(
		.INIT('h1)
	) name619 (
		_w1075_,
		_w1080_,
		_w1081_
	);
	LUT2 #(
		.INIT('h4)
	) name620 (
		_w538_,
		_w1081_,
		_w1082_
	);
	LUT2 #(
		.INIT('h1)
	) name621 (
		_w1074_,
		_w1082_,
		_w1083_
	);
	LUT2 #(
		.INIT('h8)
	) name622 (
		\P1_reg1_reg[15]/NET0131 ,
		_w746_,
		_w1084_
	);
	LUT2 #(
		.INIT('h8)
	) name623 (
		\P1_reg3_reg[14]/NET0131 ,
		_w725_,
		_w1085_
	);
	LUT2 #(
		.INIT('h8)
	) name624 (
		\P1_reg3_reg[15]/NET0131 ,
		_w1085_,
		_w1086_
	);
	LUT2 #(
		.INIT('h1)
	) name625 (
		\P1_reg3_reg[15]/NET0131 ,
		_w1085_,
		_w1087_
	);
	LUT2 #(
		.INIT('h1)
	) name626 (
		_w1086_,
		_w1087_,
		_w1088_
	);
	LUT2 #(
		.INIT('h8)
	) name627 (
		_w715_,
		_w1088_,
		_w1089_
	);
	LUT2 #(
		.INIT('h8)
	) name628 (
		\P1_reg0_reg[15]/NET0131 ,
		_w744_,
		_w1090_
	);
	LUT2 #(
		.INIT('h8)
	) name629 (
		\P1_reg2_reg[15]/NET0131 ,
		_w742_,
		_w1091_
	);
	LUT2 #(
		.INIT('h1)
	) name630 (
		_w1084_,
		_w1089_,
		_w1092_
	);
	LUT2 #(
		.INIT('h1)
	) name631 (
		_w1090_,
		_w1091_,
		_w1093_
	);
	LUT2 #(
		.INIT('h8)
	) name632 (
		_w1092_,
		_w1093_,
		_w1094_
	);
	LUT2 #(
		.INIT('h8)
	) name633 (
		_w1083_,
		_w1094_,
		_w1095_
	);
	LUT2 #(
		.INIT('h2)
	) name634 (
		\P1_IR_reg[31]/NET0131 ,
		_w474_,
		_w1096_
	);
	LUT2 #(
		.INIT('h8)
	) name635 (
		\P1_IR_reg[14]/NET0131 ,
		_w1096_,
		_w1097_
	);
	LUT2 #(
		.INIT('h1)
	) name636 (
		\P1_IR_reg[14]/NET0131 ,
		_w1096_,
		_w1098_
	);
	LUT2 #(
		.INIT('h1)
	) name637 (
		_w1097_,
		_w1098_,
		_w1099_
	);
	LUT2 #(
		.INIT('h2)
	) name638 (
		_w538_,
		_w1099_,
		_w1100_
	);
	LUT2 #(
		.INIT('h8)
	) name639 (
		\P2_datao_reg[14]/NET0131 ,
		_w543_,
		_w1101_
	);
	LUT2 #(
		.INIT('h1)
	) name640 (
		_w575_,
		_w576_,
		_w1102_
	);
	LUT2 #(
		.INIT('h4)
	) name641 (
		_w800_,
		_w1102_,
		_w1103_
	);
	LUT2 #(
		.INIT('h2)
	) name642 (
		_w800_,
		_w1102_,
		_w1104_
	);
	LUT2 #(
		.INIT('h1)
	) name643 (
		_w543_,
		_w1103_,
		_w1105_
	);
	LUT2 #(
		.INIT('h4)
	) name644 (
		_w1104_,
		_w1105_,
		_w1106_
	);
	LUT2 #(
		.INIT('h1)
	) name645 (
		_w1101_,
		_w1106_,
		_w1107_
	);
	LUT2 #(
		.INIT('h4)
	) name646 (
		_w538_,
		_w1107_,
		_w1108_
	);
	LUT2 #(
		.INIT('h1)
	) name647 (
		_w1100_,
		_w1108_,
		_w1109_
	);
	LUT2 #(
		.INIT('h8)
	) name648 (
		\P1_reg0_reg[14]/NET0131 ,
		_w744_,
		_w1110_
	);
	LUT2 #(
		.INIT('h8)
	) name649 (
		\P1_reg1_reg[14]/NET0131 ,
		_w746_,
		_w1111_
	);
	LUT2 #(
		.INIT('h1)
	) name650 (
		\P1_reg3_reg[14]/NET0131 ,
		_w725_,
		_w1112_
	);
	LUT2 #(
		.INIT('h1)
	) name651 (
		_w1085_,
		_w1112_,
		_w1113_
	);
	LUT2 #(
		.INIT('h8)
	) name652 (
		_w715_,
		_w1113_,
		_w1114_
	);
	LUT2 #(
		.INIT('h8)
	) name653 (
		\P1_reg2_reg[14]/NET0131 ,
		_w742_,
		_w1115_
	);
	LUT2 #(
		.INIT('h1)
	) name654 (
		_w1110_,
		_w1111_,
		_w1116_
	);
	LUT2 #(
		.INIT('h1)
	) name655 (
		_w1114_,
		_w1115_,
		_w1117_
	);
	LUT2 #(
		.INIT('h8)
	) name656 (
		_w1116_,
		_w1117_,
		_w1118_
	);
	LUT2 #(
		.INIT('h8)
	) name657 (
		_w1109_,
		_w1118_,
		_w1119_
	);
	LUT2 #(
		.INIT('h1)
	) name658 (
		_w1095_,
		_w1119_,
		_w1120_
	);
	LUT2 #(
		.INIT('h2)
	) name659 (
		\P1_IR_reg[31]/NET0131 ,
		_w491_,
		_w1121_
	);
	LUT2 #(
		.INIT('h2)
	) name660 (
		\P1_IR_reg[31]/NET0131 ,
		_w471_,
		_w1122_
	);
	LUT2 #(
		.INIT('h1)
	) name661 (
		_w1121_,
		_w1122_,
		_w1123_
	);
	LUT2 #(
		.INIT('h2)
	) name662 (
		\P1_IR_reg[13]/NET0131 ,
		_w1123_,
		_w1124_
	);
	LUT2 #(
		.INIT('h4)
	) name663 (
		\P1_IR_reg[13]/NET0131 ,
		_w1123_,
		_w1125_
	);
	LUT2 #(
		.INIT('h1)
	) name664 (
		_w1124_,
		_w1125_,
		_w1126_
	);
	LUT2 #(
		.INIT('h2)
	) name665 (
		_w538_,
		_w1126_,
		_w1127_
	);
	LUT2 #(
		.INIT('h8)
	) name666 (
		\P2_datao_reg[13]/NET0131 ,
		_w543_,
		_w1128_
	);
	LUT2 #(
		.INIT('h1)
	) name667 (
		_w577_,
		_w580_,
		_w1129_
	);
	LUT2 #(
		.INIT('h4)
	) name668 (
		_w865_,
		_w1129_,
		_w1130_
	);
	LUT2 #(
		.INIT('h2)
	) name669 (
		_w865_,
		_w1129_,
		_w1131_
	);
	LUT2 #(
		.INIT('h1)
	) name670 (
		_w543_,
		_w1130_,
		_w1132_
	);
	LUT2 #(
		.INIT('h4)
	) name671 (
		_w1131_,
		_w1132_,
		_w1133_
	);
	LUT2 #(
		.INIT('h1)
	) name672 (
		_w1128_,
		_w1133_,
		_w1134_
	);
	LUT2 #(
		.INIT('h4)
	) name673 (
		_w538_,
		_w1134_,
		_w1135_
	);
	LUT2 #(
		.INIT('h1)
	) name674 (
		_w1127_,
		_w1135_,
		_w1136_
	);
	LUT2 #(
		.INIT('h8)
	) name675 (
		\P1_reg2_reg[13]/NET0131 ,
		_w742_,
		_w1137_
	);
	LUT2 #(
		.INIT('h8)
	) name676 (
		\P1_reg3_reg[12]/NET0131 ,
		_w723_,
		_w1138_
	);
	LUT2 #(
		.INIT('h1)
	) name677 (
		\P1_reg3_reg[13]/NET0131 ,
		_w1138_,
		_w1139_
	);
	LUT2 #(
		.INIT('h1)
	) name678 (
		_w725_,
		_w1139_,
		_w1140_
	);
	LUT2 #(
		.INIT('h8)
	) name679 (
		_w715_,
		_w1140_,
		_w1141_
	);
	LUT2 #(
		.INIT('h8)
	) name680 (
		\P1_reg0_reg[13]/NET0131 ,
		_w744_,
		_w1142_
	);
	LUT2 #(
		.INIT('h8)
	) name681 (
		\P1_reg1_reg[13]/NET0131 ,
		_w746_,
		_w1143_
	);
	LUT2 #(
		.INIT('h1)
	) name682 (
		_w1137_,
		_w1141_,
		_w1144_
	);
	LUT2 #(
		.INIT('h1)
	) name683 (
		_w1142_,
		_w1143_,
		_w1145_
	);
	LUT2 #(
		.INIT('h8)
	) name684 (
		_w1144_,
		_w1145_,
		_w1146_
	);
	LUT2 #(
		.INIT('h8)
	) name685 (
		_w1136_,
		_w1146_,
		_w1147_
	);
	LUT2 #(
		.INIT('h1)
	) name686 (
		_w1136_,
		_w1146_,
		_w1148_
	);
	LUT2 #(
		.INIT('h8)
	) name687 (
		_w467_,
		_w489_,
		_w1149_
	);
	LUT2 #(
		.INIT('h8)
	) name688 (
		_w470_,
		_w1149_,
		_w1150_
	);
	LUT2 #(
		.INIT('h2)
	) name689 (
		\P1_IR_reg[31]/NET0131 ,
		_w1150_,
		_w1151_
	);
	LUT2 #(
		.INIT('h8)
	) name690 (
		\P1_IR_reg[12]/NET0131 ,
		_w1151_,
		_w1152_
	);
	LUT2 #(
		.INIT('h1)
	) name691 (
		\P1_IR_reg[12]/NET0131 ,
		_w1151_,
		_w1153_
	);
	LUT2 #(
		.INIT('h1)
	) name692 (
		_w1152_,
		_w1153_,
		_w1154_
	);
	LUT2 #(
		.INIT('h2)
	) name693 (
		_w538_,
		_w1154_,
		_w1155_
	);
	LUT2 #(
		.INIT('h8)
	) name694 (
		\P2_datao_reg[12]/NET0131 ,
		_w543_,
		_w1156_
	);
	LUT2 #(
		.INIT('h1)
	) name695 (
		_w582_,
		_w583_,
		_w1157_
	);
	LUT2 #(
		.INIT('h2)
	) name696 (
		_w897_,
		_w908_,
		_w1158_
	);
	LUT2 #(
		.INIT('h2)
	) name697 (
		_w1157_,
		_w1158_,
		_w1159_
	);
	LUT2 #(
		.INIT('h4)
	) name698 (
		_w1157_,
		_w1158_,
		_w1160_
	);
	LUT2 #(
		.INIT('h1)
	) name699 (
		_w543_,
		_w1159_,
		_w1161_
	);
	LUT2 #(
		.INIT('h4)
	) name700 (
		_w1160_,
		_w1161_,
		_w1162_
	);
	LUT2 #(
		.INIT('h1)
	) name701 (
		_w1156_,
		_w1162_,
		_w1163_
	);
	LUT2 #(
		.INIT('h4)
	) name702 (
		_w538_,
		_w1163_,
		_w1164_
	);
	LUT2 #(
		.INIT('h1)
	) name703 (
		_w1155_,
		_w1164_,
		_w1165_
	);
	LUT2 #(
		.INIT('h8)
	) name704 (
		\P1_reg2_reg[12]/NET0131 ,
		_w742_,
		_w1166_
	);
	LUT2 #(
		.INIT('h8)
	) name705 (
		\P1_reg0_reg[12]/NET0131 ,
		_w744_,
		_w1167_
	);
	LUT2 #(
		.INIT('h8)
	) name706 (
		\P1_reg1_reg[12]/NET0131 ,
		_w746_,
		_w1168_
	);
	LUT2 #(
		.INIT('h1)
	) name707 (
		\P1_reg3_reg[12]/NET0131 ,
		_w723_,
		_w1169_
	);
	LUT2 #(
		.INIT('h1)
	) name708 (
		_w1138_,
		_w1169_,
		_w1170_
	);
	LUT2 #(
		.INIT('h8)
	) name709 (
		_w715_,
		_w1170_,
		_w1171_
	);
	LUT2 #(
		.INIT('h1)
	) name710 (
		_w1166_,
		_w1167_,
		_w1172_
	);
	LUT2 #(
		.INIT('h1)
	) name711 (
		_w1168_,
		_w1171_,
		_w1173_
	);
	LUT2 #(
		.INIT('h8)
	) name712 (
		_w1172_,
		_w1173_,
		_w1174_
	);
	LUT2 #(
		.INIT('h1)
	) name713 (
		_w1165_,
		_w1174_,
		_w1175_
	);
	LUT2 #(
		.INIT('h1)
	) name714 (
		_w1148_,
		_w1175_,
		_w1176_
	);
	LUT2 #(
		.INIT('h1)
	) name715 (
		_w1147_,
		_w1176_,
		_w1177_
	);
	LUT2 #(
		.INIT('h8)
	) name716 (
		_w1120_,
		_w1177_,
		_w1178_
	);
	LUT2 #(
		.INIT('h1)
	) name717 (
		_w1109_,
		_w1118_,
		_w1179_
	);
	LUT2 #(
		.INIT('h1)
	) name718 (
		_w1083_,
		_w1094_,
		_w1180_
	);
	LUT2 #(
		.INIT('h1)
	) name719 (
		_w1179_,
		_w1180_,
		_w1181_
	);
	LUT2 #(
		.INIT('h1)
	) name720 (
		_w1095_,
		_w1181_,
		_w1182_
	);
	LUT2 #(
		.INIT('h1)
	) name721 (
		_w1178_,
		_w1182_,
		_w1183_
	);
	LUT2 #(
		.INIT('h8)
	) name722 (
		_w469_,
		_w1149_,
		_w1184_
	);
	LUT2 #(
		.INIT('h2)
	) name723 (
		\P1_IR_reg[31]/NET0131 ,
		_w1184_,
		_w1185_
	);
	LUT2 #(
		.INIT('h1)
	) name724 (
		\P1_IR_reg[11]/NET0131 ,
		_w1185_,
		_w1186_
	);
	LUT2 #(
		.INIT('h8)
	) name725 (
		\P1_IR_reg[11]/NET0131 ,
		_w1185_,
		_w1187_
	);
	LUT2 #(
		.INIT('h1)
	) name726 (
		_w1186_,
		_w1187_,
		_w1188_
	);
	LUT2 #(
		.INIT('h2)
	) name727 (
		_w538_,
		_w1188_,
		_w1189_
	);
	LUT2 #(
		.INIT('h8)
	) name728 (
		\P2_datao_reg[11]/NET0131 ,
		_w543_,
		_w1190_
	);
	LUT2 #(
		.INIT('h1)
	) name729 (
		_w584_,
		_w634_,
		_w1191_
	);
	LUT2 #(
		.INIT('h4)
	) name730 (
		_w633_,
		_w1191_,
		_w1192_
	);
	LUT2 #(
		.INIT('h2)
	) name731 (
		_w633_,
		_w1191_,
		_w1193_
	);
	LUT2 #(
		.INIT('h1)
	) name732 (
		_w543_,
		_w1192_,
		_w1194_
	);
	LUT2 #(
		.INIT('h4)
	) name733 (
		_w1193_,
		_w1194_,
		_w1195_
	);
	LUT2 #(
		.INIT('h1)
	) name734 (
		_w1190_,
		_w1195_,
		_w1196_
	);
	LUT2 #(
		.INIT('h4)
	) name735 (
		_w538_,
		_w1196_,
		_w1197_
	);
	LUT2 #(
		.INIT('h1)
	) name736 (
		_w1189_,
		_w1197_,
		_w1198_
	);
	LUT2 #(
		.INIT('h8)
	) name737 (
		\P1_reg2_reg[11]/NET0131 ,
		_w742_,
		_w1199_
	);
	LUT2 #(
		.INIT('h8)
	) name738 (
		\P1_reg1_reg[11]/NET0131 ,
		_w746_,
		_w1200_
	);
	LUT2 #(
		.INIT('h8)
	) name739 (
		\P1_reg0_reg[11]/NET0131 ,
		_w744_,
		_w1201_
	);
	LUT2 #(
		.INIT('h1)
	) name740 (
		\P1_reg3_reg[11]/NET0131 ,
		_w722_,
		_w1202_
	);
	LUT2 #(
		.INIT('h1)
	) name741 (
		_w723_,
		_w1202_,
		_w1203_
	);
	LUT2 #(
		.INIT('h8)
	) name742 (
		_w715_,
		_w1203_,
		_w1204_
	);
	LUT2 #(
		.INIT('h1)
	) name743 (
		_w1199_,
		_w1200_,
		_w1205_
	);
	LUT2 #(
		.INIT('h1)
	) name744 (
		_w1201_,
		_w1204_,
		_w1206_
	);
	LUT2 #(
		.INIT('h8)
	) name745 (
		_w1205_,
		_w1206_,
		_w1207_
	);
	LUT2 #(
		.INIT('h1)
	) name746 (
		_w1198_,
		_w1207_,
		_w1208_
	);
	LUT2 #(
		.INIT('h8)
	) name747 (
		_w1198_,
		_w1207_,
		_w1209_
	);
	LUT2 #(
		.INIT('h8)
	) name748 (
		\P1_reg1_reg[10]/NET0131 ,
		_w746_,
		_w1210_
	);
	LUT2 #(
		.INIT('h8)
	) name749 (
		\P1_reg2_reg[10]/NET0131 ,
		_w742_,
		_w1211_
	);
	LUT2 #(
		.INIT('h8)
	) name750 (
		\P1_reg0_reg[10]/NET0131 ,
		_w744_,
		_w1212_
	);
	LUT2 #(
		.INIT('h1)
	) name751 (
		\P1_reg3_reg[10]/NET0131 ,
		_w721_,
		_w1213_
	);
	LUT2 #(
		.INIT('h1)
	) name752 (
		_w722_,
		_w1213_,
		_w1214_
	);
	LUT2 #(
		.INIT('h8)
	) name753 (
		_w715_,
		_w1214_,
		_w1215_
	);
	LUT2 #(
		.INIT('h1)
	) name754 (
		_w1210_,
		_w1211_,
		_w1216_
	);
	LUT2 #(
		.INIT('h1)
	) name755 (
		_w1212_,
		_w1215_,
		_w1217_
	);
	LUT2 #(
		.INIT('h8)
	) name756 (
		_w1216_,
		_w1217_,
		_w1218_
	);
	LUT2 #(
		.INIT('h4)
	) name757 (
		\P1_IR_reg[9]/NET0131 ,
		_w1149_,
		_w1219_
	);
	LUT2 #(
		.INIT('h2)
	) name758 (
		\P1_IR_reg[31]/NET0131 ,
		_w1219_,
		_w1220_
	);
	LUT2 #(
		.INIT('h8)
	) name759 (
		\P1_IR_reg[10]/NET0131 ,
		_w1220_,
		_w1221_
	);
	LUT2 #(
		.INIT('h1)
	) name760 (
		\P1_IR_reg[10]/NET0131 ,
		_w1220_,
		_w1222_
	);
	LUT2 #(
		.INIT('h1)
	) name761 (
		_w1221_,
		_w1222_,
		_w1223_
	);
	LUT2 #(
		.INIT('h2)
	) name762 (
		_w538_,
		_w1223_,
		_w1224_
	);
	LUT2 #(
		.INIT('h8)
	) name763 (
		\P2_datao_reg[10]/NET0131 ,
		_w543_,
		_w1225_
	);
	LUT2 #(
		.INIT('h1)
	) name764 (
		_w593_,
		_w599_,
		_w1226_
	);
	LUT2 #(
		.INIT('h4)
	) name765 (
		_w796_,
		_w1226_,
		_w1227_
	);
	LUT2 #(
		.INIT('h2)
	) name766 (
		_w796_,
		_w1226_,
		_w1228_
	);
	LUT2 #(
		.INIT('h1)
	) name767 (
		_w543_,
		_w1227_,
		_w1229_
	);
	LUT2 #(
		.INIT('h4)
	) name768 (
		_w1228_,
		_w1229_,
		_w1230_
	);
	LUT2 #(
		.INIT('h1)
	) name769 (
		_w1225_,
		_w1230_,
		_w1231_
	);
	LUT2 #(
		.INIT('h4)
	) name770 (
		_w538_,
		_w1231_,
		_w1232_
	);
	LUT2 #(
		.INIT('h1)
	) name771 (
		_w1224_,
		_w1232_,
		_w1233_
	);
	LUT2 #(
		.INIT('h8)
	) name772 (
		_w1218_,
		_w1233_,
		_w1234_
	);
	LUT2 #(
		.INIT('h1)
	) name773 (
		_w1209_,
		_w1234_,
		_w1235_
	);
	LUT2 #(
		.INIT('h8)
	) name774 (
		\P1_reg2_reg[9]/NET0131 ,
		_w742_,
		_w1236_
	);
	LUT2 #(
		.INIT('h8)
	) name775 (
		\P1_reg0_reg[9]/NET0131 ,
		_w744_,
		_w1237_
	);
	LUT2 #(
		.INIT('h1)
	) name776 (
		\P1_reg3_reg[9]/NET0131 ,
		_w720_,
		_w1238_
	);
	LUT2 #(
		.INIT('h1)
	) name777 (
		_w721_,
		_w1238_,
		_w1239_
	);
	LUT2 #(
		.INIT('h8)
	) name778 (
		_w715_,
		_w1239_,
		_w1240_
	);
	LUT2 #(
		.INIT('h8)
	) name779 (
		\P1_reg1_reg[9]/NET0131 ,
		_w746_,
		_w1241_
	);
	LUT2 #(
		.INIT('h1)
	) name780 (
		_w1236_,
		_w1237_,
		_w1242_
	);
	LUT2 #(
		.INIT('h1)
	) name781 (
		_w1240_,
		_w1241_,
		_w1243_
	);
	LUT2 #(
		.INIT('h8)
	) name782 (
		_w1242_,
		_w1243_,
		_w1244_
	);
	LUT2 #(
		.INIT('h1)
	) name783 (
		\P1_IR_reg[9]/NET0131 ,
		_w1121_,
		_w1245_
	);
	LUT2 #(
		.INIT('h8)
	) name784 (
		\P1_IR_reg[9]/NET0131 ,
		_w1121_,
		_w1246_
	);
	LUT2 #(
		.INIT('h1)
	) name785 (
		_w1245_,
		_w1246_,
		_w1247_
	);
	LUT2 #(
		.INIT('h2)
	) name786 (
		_w538_,
		_w1247_,
		_w1248_
	);
	LUT2 #(
		.INIT('h8)
	) name787 (
		\P2_datao_reg[9]/NET0131 ,
		_w543_,
		_w1249_
	);
	LUT2 #(
		.INIT('h1)
	) name788 (
		_w592_,
		_w598_,
		_w1250_
	);
	LUT2 #(
		.INIT('h4)
	) name789 (
		_w860_,
		_w1250_,
		_w1251_
	);
	LUT2 #(
		.INIT('h2)
	) name790 (
		_w860_,
		_w1250_,
		_w1252_
	);
	LUT2 #(
		.INIT('h1)
	) name791 (
		_w543_,
		_w1251_,
		_w1253_
	);
	LUT2 #(
		.INIT('h4)
	) name792 (
		_w1252_,
		_w1253_,
		_w1254_
	);
	LUT2 #(
		.INIT('h1)
	) name793 (
		_w1249_,
		_w1254_,
		_w1255_
	);
	LUT2 #(
		.INIT('h4)
	) name794 (
		_w538_,
		_w1255_,
		_w1256_
	);
	LUT2 #(
		.INIT('h1)
	) name795 (
		_w1248_,
		_w1256_,
		_w1257_
	);
	LUT2 #(
		.INIT('h8)
	) name796 (
		_w1244_,
		_w1257_,
		_w1258_
	);
	LUT2 #(
		.INIT('h8)
	) name797 (
		\P1_reg1_reg[8]/NET0131 ,
		_w746_,
		_w1259_
	);
	LUT2 #(
		.INIT('h8)
	) name798 (
		\P1_reg2_reg[8]/NET0131 ,
		_w742_,
		_w1260_
	);
	LUT2 #(
		.INIT('h1)
	) name799 (
		\P1_reg3_reg[8]/NET0131 ,
		_w719_,
		_w1261_
	);
	LUT2 #(
		.INIT('h1)
	) name800 (
		_w720_,
		_w1261_,
		_w1262_
	);
	LUT2 #(
		.INIT('h8)
	) name801 (
		_w715_,
		_w1262_,
		_w1263_
	);
	LUT2 #(
		.INIT('h8)
	) name802 (
		\P1_reg0_reg[8]/NET0131 ,
		_w744_,
		_w1264_
	);
	LUT2 #(
		.INIT('h1)
	) name803 (
		_w1259_,
		_w1260_,
		_w1265_
	);
	LUT2 #(
		.INIT('h1)
	) name804 (
		_w1263_,
		_w1264_,
		_w1266_
	);
	LUT2 #(
		.INIT('h8)
	) name805 (
		_w1265_,
		_w1266_,
		_w1267_
	);
	LUT2 #(
		.INIT('h2)
	) name806 (
		\P1_IR_reg[31]/NET0131 ,
		_w468_,
		_w1268_
	);
	LUT2 #(
		.INIT('h1)
	) name807 (
		\P1_IR_reg[8]/NET0131 ,
		_w1268_,
		_w1269_
	);
	LUT2 #(
		.INIT('h8)
	) name808 (
		\P1_IR_reg[8]/NET0131 ,
		_w1268_,
		_w1270_
	);
	LUT2 #(
		.INIT('h1)
	) name809 (
		_w1269_,
		_w1270_,
		_w1271_
	);
	LUT2 #(
		.INIT('h2)
	) name810 (
		_w538_,
		_w1271_,
		_w1272_
	);
	LUT2 #(
		.INIT('h8)
	) name811 (
		\P2_datao_reg[8]/NET0131 ,
		_w543_,
		_w1273_
	);
	LUT2 #(
		.INIT('h1)
	) name812 (
		_w589_,
		_w595_,
		_w1274_
	);
	LUT2 #(
		.INIT('h4)
	) name813 (
		_w906_,
		_w1274_,
		_w1275_
	);
	LUT2 #(
		.INIT('h2)
	) name814 (
		_w906_,
		_w1274_,
		_w1276_
	);
	LUT2 #(
		.INIT('h1)
	) name815 (
		_w543_,
		_w1275_,
		_w1277_
	);
	LUT2 #(
		.INIT('h4)
	) name816 (
		_w1276_,
		_w1277_,
		_w1278_
	);
	LUT2 #(
		.INIT('h1)
	) name817 (
		_w1273_,
		_w1278_,
		_w1279_
	);
	LUT2 #(
		.INIT('h4)
	) name818 (
		_w538_,
		_w1279_,
		_w1280_
	);
	LUT2 #(
		.INIT('h1)
	) name819 (
		_w1272_,
		_w1280_,
		_w1281_
	);
	LUT2 #(
		.INIT('h8)
	) name820 (
		_w1267_,
		_w1281_,
		_w1282_
	);
	LUT2 #(
		.INIT('h1)
	) name821 (
		_w1258_,
		_w1282_,
		_w1283_
	);
	LUT2 #(
		.INIT('h1)
	) name822 (
		_w1244_,
		_w1257_,
		_w1284_
	);
	LUT2 #(
		.INIT('h1)
	) name823 (
		_w1218_,
		_w1233_,
		_w1285_
	);
	LUT2 #(
		.INIT('h1)
	) name824 (
		_w1284_,
		_w1285_,
		_w1286_
	);
	LUT2 #(
		.INIT('h4)
	) name825 (
		_w1283_,
		_w1286_,
		_w1287_
	);
	LUT2 #(
		.INIT('h2)
	) name826 (
		_w1235_,
		_w1287_,
		_w1288_
	);
	LUT2 #(
		.INIT('h1)
	) name827 (
		_w1208_,
		_w1288_,
		_w1289_
	);
	LUT2 #(
		.INIT('h8)
	) name828 (
		_w1165_,
		_w1174_,
		_w1290_
	);
	LUT2 #(
		.INIT('h1)
	) name829 (
		_w1147_,
		_w1290_,
		_w1291_
	);
	LUT2 #(
		.INIT('h1)
	) name830 (
		_w1148_,
		_w1179_,
		_w1292_
	);
	LUT2 #(
		.INIT('h4)
	) name831 (
		_w1291_,
		_w1292_,
		_w1293_
	);
	LUT2 #(
		.INIT('h2)
	) name832 (
		_w1120_,
		_w1293_,
		_w1294_
	);
	LUT2 #(
		.INIT('h1)
	) name833 (
		_w1180_,
		_w1294_,
		_w1295_
	);
	LUT2 #(
		.INIT('h1)
	) name834 (
		_w1289_,
		_w1295_,
		_w1296_
	);
	LUT2 #(
		.INIT('h2)
	) name835 (
		_w1183_,
		_w1296_,
		_w1297_
	);
	LUT2 #(
		.INIT('h1)
	) name836 (
		_w979_,
		_w1010_,
		_w1298_
	);
	LUT2 #(
		.INIT('h8)
	) name837 (
		_w1047_,
		_w1062_,
		_w1299_
	);
	LUT2 #(
		.INIT('h1)
	) name838 (
		_w1039_,
		_w1299_,
		_w1300_
	);
	LUT2 #(
		.INIT('h8)
	) name839 (
		_w1298_,
		_w1300_,
		_w1301_
	);
	LUT2 #(
		.INIT('h8)
	) name840 (
		\P2_datao_reg[22]/NET0131 ,
		_w543_,
		_w1302_
	);
	LUT2 #(
		.INIT('h1)
	) name841 (
		_w544_,
		_w545_,
		_w1303_
	);
	LUT2 #(
		.INIT('h4)
	) name842 (
		_w813_,
		_w1303_,
		_w1304_
	);
	LUT2 #(
		.INIT('h2)
	) name843 (
		_w813_,
		_w1303_,
		_w1305_
	);
	LUT2 #(
		.INIT('h1)
	) name844 (
		_w543_,
		_w1304_,
		_w1306_
	);
	LUT2 #(
		.INIT('h4)
	) name845 (
		_w1305_,
		_w1306_,
		_w1307_
	);
	LUT2 #(
		.INIT('h1)
	) name846 (
		_w1302_,
		_w1307_,
		_w1308_
	);
	LUT2 #(
		.INIT('h1)
	) name847 (
		_w538_,
		_w1308_,
		_w1309_
	);
	LUT2 #(
		.INIT('h8)
	) name848 (
		\P1_reg2_reg[22]/NET0131 ,
		_w742_,
		_w1310_
	);
	LUT2 #(
		.INIT('h8)
	) name849 (
		\P1_reg1_reg[22]/NET0131 ,
		_w746_,
		_w1311_
	);
	LUT2 #(
		.INIT('h8)
	) name850 (
		\P1_reg0_reg[22]/NET0131 ,
		_w744_,
		_w1312_
	);
	LUT2 #(
		.INIT('h1)
	) name851 (
		\P1_reg3_reg[22]/NET0131 ,
		_w1054_,
		_w1313_
	);
	LUT2 #(
		.INIT('h1)
	) name852 (
		_w1055_,
		_w1313_,
		_w1314_
	);
	LUT2 #(
		.INIT('h8)
	) name853 (
		_w715_,
		_w1314_,
		_w1315_
	);
	LUT2 #(
		.INIT('h1)
	) name854 (
		_w1310_,
		_w1311_,
		_w1316_
	);
	LUT2 #(
		.INIT('h4)
	) name855 (
		_w1312_,
		_w1316_,
		_w1317_
	);
	LUT2 #(
		.INIT('h4)
	) name856 (
		_w1315_,
		_w1317_,
		_w1318_
	);
	LUT2 #(
		.INIT('h8)
	) name857 (
		_w1309_,
		_w1318_,
		_w1319_
	);
	LUT2 #(
		.INIT('h8)
	) name858 (
		\P2_datao_reg[23]/NET0131 ,
		_w543_,
		_w1320_
	);
	LUT2 #(
		.INIT('h1)
	) name859 (
		_w657_,
		_w675_,
		_w1321_
	);
	LUT2 #(
		.INIT('h4)
	) name860 (
		_w645_,
		_w1321_,
		_w1322_
	);
	LUT2 #(
		.INIT('h2)
	) name861 (
		_w645_,
		_w1321_,
		_w1323_
	);
	LUT2 #(
		.INIT('h1)
	) name862 (
		_w543_,
		_w1322_,
		_w1324_
	);
	LUT2 #(
		.INIT('h4)
	) name863 (
		_w1323_,
		_w1324_,
		_w1325_
	);
	LUT2 #(
		.INIT('h1)
	) name864 (
		_w1320_,
		_w1325_,
		_w1326_
	);
	LUT2 #(
		.INIT('h1)
	) name865 (
		_w538_,
		_w1326_,
		_w1327_
	);
	LUT2 #(
		.INIT('h8)
	) name866 (
		\P1_reg0_reg[23]/NET0131 ,
		_w744_,
		_w1328_
	);
	LUT2 #(
		.INIT('h1)
	) name867 (
		\P1_reg3_reg[23]/NET0131 ,
		_w1055_,
		_w1329_
	);
	LUT2 #(
		.INIT('h1)
	) name868 (
		_w1056_,
		_w1329_,
		_w1330_
	);
	LUT2 #(
		.INIT('h8)
	) name869 (
		_w715_,
		_w1330_,
		_w1331_
	);
	LUT2 #(
		.INIT('h8)
	) name870 (
		\P1_reg1_reg[23]/NET0131 ,
		_w746_,
		_w1332_
	);
	LUT2 #(
		.INIT('h8)
	) name871 (
		\P1_reg2_reg[23]/NET0131 ,
		_w742_,
		_w1333_
	);
	LUT2 #(
		.INIT('h1)
	) name872 (
		_w1328_,
		_w1332_,
		_w1334_
	);
	LUT2 #(
		.INIT('h4)
	) name873 (
		_w1333_,
		_w1334_,
		_w1335_
	);
	LUT2 #(
		.INIT('h4)
	) name874 (
		_w1331_,
		_w1335_,
		_w1336_
	);
	LUT2 #(
		.INIT('h8)
	) name875 (
		_w1327_,
		_w1336_,
		_w1337_
	);
	LUT2 #(
		.INIT('h1)
	) name876 (
		_w1319_,
		_w1337_,
		_w1338_
	);
	LUT2 #(
		.INIT('h8)
	) name877 (
		\P2_datao_reg[21]/NET0131 ,
		_w543_,
		_w1339_
	);
	LUT2 #(
		.INIT('h1)
	) name878 (
		_w546_,
		_w549_,
		_w1340_
	);
	LUT2 #(
		.INIT('h4)
	) name879 (
		_w871_,
		_w1340_,
		_w1341_
	);
	LUT2 #(
		.INIT('h2)
	) name880 (
		_w871_,
		_w1340_,
		_w1342_
	);
	LUT2 #(
		.INIT('h1)
	) name881 (
		_w543_,
		_w1341_,
		_w1343_
	);
	LUT2 #(
		.INIT('h4)
	) name882 (
		_w1342_,
		_w1343_,
		_w1344_
	);
	LUT2 #(
		.INIT('h1)
	) name883 (
		_w1339_,
		_w1344_,
		_w1345_
	);
	LUT2 #(
		.INIT('h1)
	) name884 (
		_w538_,
		_w1345_,
		_w1346_
	);
	LUT2 #(
		.INIT('h8)
	) name885 (
		\P1_reg0_reg[21]/NET0131 ,
		_w744_,
		_w1347_
	);
	LUT2 #(
		.INIT('h8)
	) name886 (
		\P1_reg2_reg[21]/NET0131 ,
		_w742_,
		_w1348_
	);
	LUT2 #(
		.INIT('h8)
	) name887 (
		\P1_reg1_reg[21]/NET0131 ,
		_w746_,
		_w1349_
	);
	LUT2 #(
		.INIT('h8)
	) name888 (
		\P1_reg3_reg[20]/NET0131 ,
		_w1053_,
		_w1350_
	);
	LUT2 #(
		.INIT('h1)
	) name889 (
		\P1_reg3_reg[21]/NET0131 ,
		_w1350_,
		_w1351_
	);
	LUT2 #(
		.INIT('h1)
	) name890 (
		_w1054_,
		_w1351_,
		_w1352_
	);
	LUT2 #(
		.INIT('h8)
	) name891 (
		_w715_,
		_w1352_,
		_w1353_
	);
	LUT2 #(
		.INIT('h1)
	) name892 (
		_w1347_,
		_w1348_,
		_w1354_
	);
	LUT2 #(
		.INIT('h4)
	) name893 (
		_w1349_,
		_w1354_,
		_w1355_
	);
	LUT2 #(
		.INIT('h4)
	) name894 (
		_w1353_,
		_w1355_,
		_w1356_
	);
	LUT2 #(
		.INIT('h8)
	) name895 (
		_w1346_,
		_w1356_,
		_w1357_
	);
	LUT2 #(
		.INIT('h8)
	) name896 (
		\P2_datao_reg[20]/NET0131 ,
		_w543_,
		_w1358_
	);
	LUT2 #(
		.INIT('h1)
	) name897 (
		_w551_,
		_w552_,
		_w1359_
	);
	LUT2 #(
		.INIT('h4)
	) name898 (
		_w918_,
		_w1359_,
		_w1360_
	);
	LUT2 #(
		.INIT('h2)
	) name899 (
		_w918_,
		_w1359_,
		_w1361_
	);
	LUT2 #(
		.INIT('h1)
	) name900 (
		_w543_,
		_w1360_,
		_w1362_
	);
	LUT2 #(
		.INIT('h4)
	) name901 (
		_w1361_,
		_w1362_,
		_w1363_
	);
	LUT2 #(
		.INIT('h1)
	) name902 (
		_w1358_,
		_w1363_,
		_w1364_
	);
	LUT2 #(
		.INIT('h1)
	) name903 (
		_w538_,
		_w1364_,
		_w1365_
	);
	LUT2 #(
		.INIT('h8)
	) name904 (
		\P1_reg0_reg[20]/NET0131 ,
		_w744_,
		_w1366_
	);
	LUT2 #(
		.INIT('h8)
	) name905 (
		\P1_reg2_reg[20]/NET0131 ,
		_w742_,
		_w1367_
	);
	LUT2 #(
		.INIT('h8)
	) name906 (
		\P1_reg1_reg[20]/NET0131 ,
		_w746_,
		_w1368_
	);
	LUT2 #(
		.INIT('h1)
	) name907 (
		\P1_reg3_reg[20]/NET0131 ,
		_w1053_,
		_w1369_
	);
	LUT2 #(
		.INIT('h1)
	) name908 (
		_w1350_,
		_w1369_,
		_w1370_
	);
	LUT2 #(
		.INIT('h8)
	) name909 (
		_w715_,
		_w1370_,
		_w1371_
	);
	LUT2 #(
		.INIT('h1)
	) name910 (
		_w1366_,
		_w1367_,
		_w1372_
	);
	LUT2 #(
		.INIT('h4)
	) name911 (
		_w1368_,
		_w1372_,
		_w1373_
	);
	LUT2 #(
		.INIT('h4)
	) name912 (
		_w1371_,
		_w1373_,
		_w1374_
	);
	LUT2 #(
		.INIT('h8)
	) name913 (
		_w1365_,
		_w1374_,
		_w1375_
	);
	LUT2 #(
		.INIT('h1)
	) name914 (
		_w1357_,
		_w1375_,
		_w1376_
	);
	LUT2 #(
		.INIT('h8)
	) name915 (
		_w1338_,
		_w1376_,
		_w1377_
	);
	LUT2 #(
		.INIT('h2)
	) name916 (
		\P1_IR_reg[31]/NET0131 ,
		_w514_,
		_w1378_
	);
	LUT2 #(
		.INIT('h1)
	) name917 (
		\P1_IR_reg[16]/NET0131 ,
		\P1_IR_reg[17]/NET0131 ,
		_w1379_
	);
	LUT2 #(
		.INIT('h2)
	) name918 (
		\P1_IR_reg[31]/NET0131 ,
		_w1379_,
		_w1380_
	);
	LUT2 #(
		.INIT('h1)
	) name919 (
		_w1378_,
		_w1380_,
		_w1381_
	);
	LUT2 #(
		.INIT('h2)
	) name920 (
		\P1_IR_reg[18]/NET0131 ,
		_w1381_,
		_w1382_
	);
	LUT2 #(
		.INIT('h4)
	) name921 (
		\P1_IR_reg[18]/NET0131 ,
		_w1381_,
		_w1383_
	);
	LUT2 #(
		.INIT('h1)
	) name922 (
		_w1382_,
		_w1383_,
		_w1384_
	);
	LUT2 #(
		.INIT('h2)
	) name923 (
		_w538_,
		_w1384_,
		_w1385_
	);
	LUT2 #(
		.INIT('h8)
	) name924 (
		\P2_datao_reg[18]/NET0131 ,
		_w543_,
		_w1386_
	);
	LUT2 #(
		.INIT('h1)
	) name925 (
		_w561_,
		_w562_,
		_w1387_
	);
	LUT2 #(
		.INIT('h4)
	) name926 (
		_w809_,
		_w1387_,
		_w1388_
	);
	LUT2 #(
		.INIT('h2)
	) name927 (
		_w809_,
		_w1387_,
		_w1389_
	);
	LUT2 #(
		.INIT('h1)
	) name928 (
		_w543_,
		_w1388_,
		_w1390_
	);
	LUT2 #(
		.INIT('h4)
	) name929 (
		_w1389_,
		_w1390_,
		_w1391_
	);
	LUT2 #(
		.INIT('h1)
	) name930 (
		_w1386_,
		_w1391_,
		_w1392_
	);
	LUT2 #(
		.INIT('h4)
	) name931 (
		_w538_,
		_w1392_,
		_w1393_
	);
	LUT2 #(
		.INIT('h1)
	) name932 (
		_w1385_,
		_w1393_,
		_w1394_
	);
	LUT2 #(
		.INIT('h8)
	) name933 (
		\P1_reg1_reg[18]/NET0131 ,
		_w746_,
		_w1395_
	);
	LUT2 #(
		.INIT('h8)
	) name934 (
		\P1_reg0_reg[18]/NET0131 ,
		_w744_,
		_w1396_
	);
	LUT2 #(
		.INIT('h8)
	) name935 (
		\P1_reg2_reg[18]/NET0131 ,
		_w742_,
		_w1397_
	);
	LUT2 #(
		.INIT('h1)
	) name936 (
		\P1_reg3_reg[18]/NET0131 ,
		_w1051_,
		_w1398_
	);
	LUT2 #(
		.INIT('h1)
	) name937 (
		_w1052_,
		_w1398_,
		_w1399_
	);
	LUT2 #(
		.INIT('h8)
	) name938 (
		_w715_,
		_w1399_,
		_w1400_
	);
	LUT2 #(
		.INIT('h1)
	) name939 (
		_w1395_,
		_w1396_,
		_w1401_
	);
	LUT2 #(
		.INIT('h4)
	) name940 (
		_w1397_,
		_w1401_,
		_w1402_
	);
	LUT2 #(
		.INIT('h4)
	) name941 (
		_w1400_,
		_w1402_,
		_w1403_
	);
	LUT2 #(
		.INIT('h8)
	) name942 (
		_w1394_,
		_w1403_,
		_w1404_
	);
	LUT2 #(
		.INIT('h2)
	) name943 (
		\P1_IR_reg[31]/NET0131 ,
		_w506_,
		_w1405_
	);
	LUT2 #(
		.INIT('h1)
	) name944 (
		\P1_IR_reg[19]/NET0131 ,
		_w1405_,
		_w1406_
	);
	LUT2 #(
		.INIT('h8)
	) name945 (
		\P1_IR_reg[19]/NET0131 ,
		_w1405_,
		_w1407_
	);
	LUT2 #(
		.INIT('h1)
	) name946 (
		_w1406_,
		_w1407_,
		_w1408_
	);
	LUT2 #(
		.INIT('h2)
	) name947 (
		_w538_,
		_w1408_,
		_w1409_
	);
	LUT2 #(
		.INIT('h8)
	) name948 (
		\P2_datao_reg[19]/NET0131 ,
		_w543_,
		_w1410_
	);
	LUT2 #(
		.INIT('h1)
	) name949 (
		_w553_,
		_w558_,
		_w1411_
	);
	LUT2 #(
		.INIT('h4)
	) name950 (
		_w643_,
		_w1411_,
		_w1412_
	);
	LUT2 #(
		.INIT('h2)
	) name951 (
		_w643_,
		_w1411_,
		_w1413_
	);
	LUT2 #(
		.INIT('h1)
	) name952 (
		_w543_,
		_w1412_,
		_w1414_
	);
	LUT2 #(
		.INIT('h4)
	) name953 (
		_w1413_,
		_w1414_,
		_w1415_
	);
	LUT2 #(
		.INIT('h1)
	) name954 (
		_w1410_,
		_w1415_,
		_w1416_
	);
	LUT2 #(
		.INIT('h4)
	) name955 (
		_w538_,
		_w1416_,
		_w1417_
	);
	LUT2 #(
		.INIT('h1)
	) name956 (
		_w1409_,
		_w1417_,
		_w1418_
	);
	LUT2 #(
		.INIT('h8)
	) name957 (
		\P1_reg0_reg[19]/NET0131 ,
		_w744_,
		_w1419_
	);
	LUT2 #(
		.INIT('h8)
	) name958 (
		\P1_reg2_reg[19]/NET0131 ,
		_w742_,
		_w1420_
	);
	LUT2 #(
		.INIT('h8)
	) name959 (
		\P1_reg1_reg[19]/NET0131 ,
		_w746_,
		_w1421_
	);
	LUT2 #(
		.INIT('h1)
	) name960 (
		\P1_reg3_reg[19]/NET0131 ,
		_w1052_,
		_w1422_
	);
	LUT2 #(
		.INIT('h1)
	) name961 (
		_w1053_,
		_w1422_,
		_w1423_
	);
	LUT2 #(
		.INIT('h8)
	) name962 (
		_w715_,
		_w1423_,
		_w1424_
	);
	LUT2 #(
		.INIT('h1)
	) name963 (
		_w1419_,
		_w1420_,
		_w1425_
	);
	LUT2 #(
		.INIT('h4)
	) name964 (
		_w1421_,
		_w1425_,
		_w1426_
	);
	LUT2 #(
		.INIT('h4)
	) name965 (
		_w1424_,
		_w1426_,
		_w1427_
	);
	LUT2 #(
		.INIT('h8)
	) name966 (
		_w1418_,
		_w1427_,
		_w1428_
	);
	LUT2 #(
		.INIT('h1)
	) name967 (
		_w1404_,
		_w1428_,
		_w1429_
	);
	LUT2 #(
		.INIT('h2)
	) name968 (
		\P1_IR_reg[31]/NET0131 ,
		_w495_,
		_w1430_
	);
	LUT2 #(
		.INIT('h2)
	) name969 (
		\P1_IR_reg[17]/NET0131 ,
		_w1430_,
		_w1431_
	);
	LUT2 #(
		.INIT('h4)
	) name970 (
		\P1_IR_reg[17]/NET0131 ,
		_w1430_,
		_w1432_
	);
	LUT2 #(
		.INIT('h1)
	) name971 (
		_w1431_,
		_w1432_,
		_w1433_
	);
	LUT2 #(
		.INIT('h8)
	) name972 (
		_w538_,
		_w1433_,
		_w1434_
	);
	LUT2 #(
		.INIT('h8)
	) name973 (
		\P2_datao_reg[17]/NET0131 ,
		_w543_,
		_w1435_
	);
	LUT2 #(
		.INIT('h1)
	) name974 (
		_w563_,
		_w566_,
		_w1436_
	);
	LUT2 #(
		.INIT('h4)
	) name975 (
		_w868_,
		_w1436_,
		_w1437_
	);
	LUT2 #(
		.INIT('h2)
	) name976 (
		_w868_,
		_w1436_,
		_w1438_
	);
	LUT2 #(
		.INIT('h1)
	) name977 (
		_w543_,
		_w1437_,
		_w1439_
	);
	LUT2 #(
		.INIT('h4)
	) name978 (
		_w1438_,
		_w1439_,
		_w1440_
	);
	LUT2 #(
		.INIT('h1)
	) name979 (
		_w1435_,
		_w1440_,
		_w1441_
	);
	LUT2 #(
		.INIT('h4)
	) name980 (
		_w538_,
		_w1441_,
		_w1442_
	);
	LUT2 #(
		.INIT('h1)
	) name981 (
		_w1434_,
		_w1442_,
		_w1443_
	);
	LUT2 #(
		.INIT('h8)
	) name982 (
		\P1_reg0_reg[17]/NET0131 ,
		_w744_,
		_w1444_
	);
	LUT2 #(
		.INIT('h8)
	) name983 (
		\P1_reg1_reg[17]/NET0131 ,
		_w746_,
		_w1445_
	);
	LUT2 #(
		.INIT('h1)
	) name984 (
		\P1_reg3_reg[17]/NET0131 ,
		_w728_,
		_w1446_
	);
	LUT2 #(
		.INIT('h1)
	) name985 (
		_w1051_,
		_w1446_,
		_w1447_
	);
	LUT2 #(
		.INIT('h8)
	) name986 (
		_w715_,
		_w1447_,
		_w1448_
	);
	LUT2 #(
		.INIT('h8)
	) name987 (
		\P1_reg2_reg[17]/NET0131 ,
		_w742_,
		_w1449_
	);
	LUT2 #(
		.INIT('h1)
	) name988 (
		_w1444_,
		_w1445_,
		_w1450_
	);
	LUT2 #(
		.INIT('h1)
	) name989 (
		_w1448_,
		_w1449_,
		_w1451_
	);
	LUT2 #(
		.INIT('h8)
	) name990 (
		_w1450_,
		_w1451_,
		_w1452_
	);
	LUT2 #(
		.INIT('h8)
	) name991 (
		_w1443_,
		_w1452_,
		_w1453_
	);
	LUT2 #(
		.INIT('h1)
	) name992 (
		\P1_IR_reg[16]/NET0131 ,
		_w1378_,
		_w1454_
	);
	LUT2 #(
		.INIT('h8)
	) name993 (
		\P1_IR_reg[16]/NET0131 ,
		_w1378_,
		_w1455_
	);
	LUT2 #(
		.INIT('h1)
	) name994 (
		_w1454_,
		_w1455_,
		_w1456_
	);
	LUT2 #(
		.INIT('h2)
	) name995 (
		_w538_,
		_w1456_,
		_w1457_
	);
	LUT2 #(
		.INIT('h8)
	) name996 (
		\P2_datao_reg[16]/NET0131 ,
		_w543_,
		_w1458_
	);
	LUT2 #(
		.INIT('h1)
	) name997 (
		_w568_,
		_w570_,
		_w1459_
	);
	LUT2 #(
		.INIT('h4)
	) name998 (
		_w912_,
		_w1459_,
		_w1460_
	);
	LUT2 #(
		.INIT('h2)
	) name999 (
		_w912_,
		_w1459_,
		_w1461_
	);
	LUT2 #(
		.INIT('h1)
	) name1000 (
		_w543_,
		_w1460_,
		_w1462_
	);
	LUT2 #(
		.INIT('h4)
	) name1001 (
		_w1461_,
		_w1462_,
		_w1463_
	);
	LUT2 #(
		.INIT('h1)
	) name1002 (
		_w1458_,
		_w1463_,
		_w1464_
	);
	LUT2 #(
		.INIT('h4)
	) name1003 (
		_w538_,
		_w1464_,
		_w1465_
	);
	LUT2 #(
		.INIT('h1)
	) name1004 (
		_w1457_,
		_w1465_,
		_w1466_
	);
	LUT2 #(
		.INIT('h8)
	) name1005 (
		\P1_reg0_reg[16]/NET0131 ,
		_w744_,
		_w1467_
	);
	LUT2 #(
		.INIT('h8)
	) name1006 (
		\P1_reg2_reg[16]/NET0131 ,
		_w742_,
		_w1468_
	);
	LUT2 #(
		.INIT('h8)
	) name1007 (
		\P1_reg1_reg[16]/NET0131 ,
		_w746_,
		_w1469_
	);
	LUT2 #(
		.INIT('h1)
	) name1008 (
		\P1_reg3_reg[16]/NET0131 ,
		_w1086_,
		_w1470_
	);
	LUT2 #(
		.INIT('h1)
	) name1009 (
		_w728_,
		_w1470_,
		_w1471_
	);
	LUT2 #(
		.INIT('h8)
	) name1010 (
		_w715_,
		_w1471_,
		_w1472_
	);
	LUT2 #(
		.INIT('h1)
	) name1011 (
		_w1467_,
		_w1468_,
		_w1473_
	);
	LUT2 #(
		.INIT('h4)
	) name1012 (
		_w1469_,
		_w1473_,
		_w1474_
	);
	LUT2 #(
		.INIT('h4)
	) name1013 (
		_w1472_,
		_w1474_,
		_w1475_
	);
	LUT2 #(
		.INIT('h8)
	) name1014 (
		_w1466_,
		_w1475_,
		_w1476_
	);
	LUT2 #(
		.INIT('h1)
	) name1015 (
		_w1453_,
		_w1476_,
		_w1477_
	);
	LUT2 #(
		.INIT('h8)
	) name1016 (
		_w1429_,
		_w1477_,
		_w1478_
	);
	LUT2 #(
		.INIT('h8)
	) name1017 (
		_w1377_,
		_w1478_,
		_w1479_
	);
	LUT2 #(
		.INIT('h8)
	) name1018 (
		_w1120_,
		_w1291_,
		_w1480_
	);
	LUT2 #(
		.INIT('h1)
	) name1019 (
		_w1267_,
		_w1281_,
		_w1481_
	);
	LUT2 #(
		.INIT('h1)
	) name1020 (
		_w1284_,
		_w1481_,
		_w1482_
	);
	LUT2 #(
		.INIT('h1)
	) name1021 (
		_w1258_,
		_w1482_,
		_w1483_
	);
	LUT2 #(
		.INIT('h8)
	) name1022 (
		_w1235_,
		_w1483_,
		_w1484_
	);
	LUT2 #(
		.INIT('h1)
	) name1023 (
		_w1208_,
		_w1285_,
		_w1485_
	);
	LUT2 #(
		.INIT('h1)
	) name1024 (
		_w1209_,
		_w1485_,
		_w1486_
	);
	LUT2 #(
		.INIT('h1)
	) name1025 (
		_w1484_,
		_w1486_,
		_w1487_
	);
	LUT2 #(
		.INIT('h2)
	) name1026 (
		_w1480_,
		_w1487_,
		_w1488_
	);
	LUT2 #(
		.INIT('h2)
	) name1027 (
		_w1183_,
		_w1488_,
		_w1489_
	);
	LUT2 #(
		.INIT('h1)
	) name1028 (
		\P1_reg3_reg[7]/NET0131 ,
		_w718_,
		_w1490_
	);
	LUT2 #(
		.INIT('h1)
	) name1029 (
		_w719_,
		_w1490_,
		_w1491_
	);
	LUT2 #(
		.INIT('h8)
	) name1030 (
		_w715_,
		_w1491_,
		_w1492_
	);
	LUT2 #(
		.INIT('h8)
	) name1031 (
		\P1_reg2_reg[7]/NET0131 ,
		_w742_,
		_w1493_
	);
	LUT2 #(
		.INIT('h8)
	) name1032 (
		\P1_reg1_reg[7]/NET0131 ,
		_w746_,
		_w1494_
	);
	LUT2 #(
		.INIT('h8)
	) name1033 (
		\P1_reg0_reg[7]/NET0131 ,
		_w744_,
		_w1495_
	);
	LUT2 #(
		.INIT('h1)
	) name1034 (
		_w1492_,
		_w1493_,
		_w1496_
	);
	LUT2 #(
		.INIT('h1)
	) name1035 (
		_w1494_,
		_w1495_,
		_w1497_
	);
	LUT2 #(
		.INIT('h8)
	) name1036 (
		_w1496_,
		_w1497_,
		_w1498_
	);
	LUT2 #(
		.INIT('h8)
	) name1037 (
		\P2_datao_reg[7]/NET0131 ,
		_w543_,
		_w1499_
	);
	LUT2 #(
		.INIT('h1)
	) name1038 (
		_w590_,
		_w628_,
		_w1500_
	);
	LUT2 #(
		.INIT('h4)
	) name1039 (
		_w627_,
		_w1500_,
		_w1501_
	);
	LUT2 #(
		.INIT('h2)
	) name1040 (
		_w627_,
		_w1500_,
		_w1502_
	);
	LUT2 #(
		.INIT('h1)
	) name1041 (
		_w543_,
		_w1501_,
		_w1503_
	);
	LUT2 #(
		.INIT('h4)
	) name1042 (
		_w1502_,
		_w1503_,
		_w1504_
	);
	LUT2 #(
		.INIT('h1)
	) name1043 (
		_w1499_,
		_w1504_,
		_w1505_
	);
	LUT2 #(
		.INIT('h1)
	) name1044 (
		_w538_,
		_w1505_,
		_w1506_
	);
	LUT2 #(
		.INIT('h2)
	) name1045 (
		\P1_IR_reg[31]/NET0131 ,
		_w467_,
		_w1507_
	);
	LUT2 #(
		.INIT('h8)
	) name1046 (
		\P1_IR_reg[31]/NET0131 ,
		\P1_IR_reg[6]/NET0131 ,
		_w1508_
	);
	LUT2 #(
		.INIT('h1)
	) name1047 (
		_w1507_,
		_w1508_,
		_w1509_
	);
	LUT2 #(
		.INIT('h2)
	) name1048 (
		\P1_IR_reg[7]/NET0131 ,
		_w1509_,
		_w1510_
	);
	LUT2 #(
		.INIT('h4)
	) name1049 (
		\P1_IR_reg[7]/NET0131 ,
		_w1509_,
		_w1511_
	);
	LUT2 #(
		.INIT('h1)
	) name1050 (
		_w1510_,
		_w1511_,
		_w1512_
	);
	LUT2 #(
		.INIT('h8)
	) name1051 (
		_w538_,
		_w1512_,
		_w1513_
	);
	LUT2 #(
		.INIT('h1)
	) name1052 (
		_w1506_,
		_w1513_,
		_w1514_
	);
	LUT2 #(
		.INIT('h2)
	) name1053 (
		_w1498_,
		_w1514_,
		_w1515_
	);
	LUT2 #(
		.INIT('h8)
	) name1054 (
		\P1_reg0_reg[6]/NET0131 ,
		_w744_,
		_w1516_
	);
	LUT2 #(
		.INIT('h1)
	) name1055 (
		\P1_reg3_reg[6]/NET0131 ,
		_w717_,
		_w1517_
	);
	LUT2 #(
		.INIT('h1)
	) name1056 (
		_w718_,
		_w1517_,
		_w1518_
	);
	LUT2 #(
		.INIT('h8)
	) name1057 (
		_w715_,
		_w1518_,
		_w1519_
	);
	LUT2 #(
		.INIT('h8)
	) name1058 (
		\P1_reg1_reg[6]/NET0131 ,
		_w746_,
		_w1520_
	);
	LUT2 #(
		.INIT('h8)
	) name1059 (
		\P1_reg2_reg[6]/NET0131 ,
		_w742_,
		_w1521_
	);
	LUT2 #(
		.INIT('h1)
	) name1060 (
		_w1516_,
		_w1519_,
		_w1522_
	);
	LUT2 #(
		.INIT('h1)
	) name1061 (
		_w1520_,
		_w1521_,
		_w1523_
	);
	LUT2 #(
		.INIT('h8)
	) name1062 (
		_w1522_,
		_w1523_,
		_w1524_
	);
	LUT2 #(
		.INIT('h8)
	) name1063 (
		\P2_datao_reg[6]/NET0131 ,
		_w543_,
		_w1525_
	);
	LUT2 #(
		.INIT('h1)
	) name1064 (
		_w602_,
		_w604_,
		_w1526_
	);
	LUT2 #(
		.INIT('h4)
	) name1065 (
		_w787_,
		_w1526_,
		_w1527_
	);
	LUT2 #(
		.INIT('h2)
	) name1066 (
		_w787_,
		_w1526_,
		_w1528_
	);
	LUT2 #(
		.INIT('h1)
	) name1067 (
		_w543_,
		_w1527_,
		_w1529_
	);
	LUT2 #(
		.INIT('h4)
	) name1068 (
		_w1528_,
		_w1529_,
		_w1530_
	);
	LUT2 #(
		.INIT('h1)
	) name1069 (
		_w1525_,
		_w1530_,
		_w1531_
	);
	LUT2 #(
		.INIT('h1)
	) name1070 (
		_w538_,
		_w1531_,
		_w1532_
	);
	LUT2 #(
		.INIT('h2)
	) name1071 (
		\P1_IR_reg[6]/NET0131 ,
		_w1507_,
		_w1533_
	);
	LUT2 #(
		.INIT('h4)
	) name1072 (
		\P1_IR_reg[6]/NET0131 ,
		_w1507_,
		_w1534_
	);
	LUT2 #(
		.INIT('h1)
	) name1073 (
		_w1533_,
		_w1534_,
		_w1535_
	);
	LUT2 #(
		.INIT('h2)
	) name1074 (
		_w538_,
		_w1535_,
		_w1536_
	);
	LUT2 #(
		.INIT('h1)
	) name1075 (
		_w1532_,
		_w1536_,
		_w1537_
	);
	LUT2 #(
		.INIT('h2)
	) name1076 (
		_w1524_,
		_w1537_,
		_w1538_
	);
	LUT2 #(
		.INIT('h1)
	) name1077 (
		_w1515_,
		_w1538_,
		_w1539_
	);
	LUT2 #(
		.INIT('h8)
	) name1078 (
		\P1_reg0_reg[5]/NET0131 ,
		_w744_,
		_w1540_
	);
	LUT2 #(
		.INIT('h8)
	) name1079 (
		\P1_reg1_reg[5]/NET0131 ,
		_w746_,
		_w1541_
	);
	LUT2 #(
		.INIT('h1)
	) name1080 (
		\P1_reg3_reg[5]/NET0131 ,
		_w716_,
		_w1542_
	);
	LUT2 #(
		.INIT('h1)
	) name1081 (
		_w717_,
		_w1542_,
		_w1543_
	);
	LUT2 #(
		.INIT('h8)
	) name1082 (
		_w715_,
		_w1543_,
		_w1544_
	);
	LUT2 #(
		.INIT('h8)
	) name1083 (
		\P1_reg2_reg[5]/NET0131 ,
		_w742_,
		_w1545_
	);
	LUT2 #(
		.INIT('h1)
	) name1084 (
		_w1540_,
		_w1541_,
		_w1546_
	);
	LUT2 #(
		.INIT('h1)
	) name1085 (
		_w1544_,
		_w1545_,
		_w1547_
	);
	LUT2 #(
		.INIT('h8)
	) name1086 (
		_w1546_,
		_w1547_,
		_w1548_
	);
	LUT2 #(
		.INIT('h8)
	) name1087 (
		\P2_datao_reg[5]/NET0131 ,
		_w543_,
		_w1549_
	);
	LUT2 #(
		.INIT('h1)
	) name1088 (
		_w603_,
		_w622_,
		_w1550_
	);
	LUT2 #(
		.INIT('h4)
	) name1089 (
		_w854_,
		_w1550_,
		_w1551_
	);
	LUT2 #(
		.INIT('h2)
	) name1090 (
		_w854_,
		_w1550_,
		_w1552_
	);
	LUT2 #(
		.INIT('h1)
	) name1091 (
		_w543_,
		_w1551_,
		_w1553_
	);
	LUT2 #(
		.INIT('h4)
	) name1092 (
		_w1552_,
		_w1553_,
		_w1554_
	);
	LUT2 #(
		.INIT('h1)
	) name1093 (
		_w1549_,
		_w1554_,
		_w1555_
	);
	LUT2 #(
		.INIT('h1)
	) name1094 (
		_w538_,
		_w1555_,
		_w1556_
	);
	LUT2 #(
		.INIT('h2)
	) name1095 (
		\P1_IR_reg[31]/NET0131 ,
		_w488_,
		_w1557_
	);
	LUT2 #(
		.INIT('h4)
	) name1096 (
		\P1_IR_reg[5]/NET0131 ,
		_w1557_,
		_w1558_
	);
	LUT2 #(
		.INIT('h2)
	) name1097 (
		\P1_IR_reg[5]/NET0131 ,
		_w1557_,
		_w1559_
	);
	LUT2 #(
		.INIT('h1)
	) name1098 (
		_w1558_,
		_w1559_,
		_w1560_
	);
	LUT2 #(
		.INIT('h2)
	) name1099 (
		_w538_,
		_w1560_,
		_w1561_
	);
	LUT2 #(
		.INIT('h1)
	) name1100 (
		_w1556_,
		_w1561_,
		_w1562_
	);
	LUT2 #(
		.INIT('h2)
	) name1101 (
		_w1548_,
		_w1562_,
		_w1563_
	);
	LUT2 #(
		.INIT('h8)
	) name1102 (
		\P1_reg1_reg[4]/NET0131 ,
		_w746_,
		_w1564_
	);
	LUT2 #(
		.INIT('h8)
	) name1103 (
		\P1_reg2_reg[4]/NET0131 ,
		_w742_,
		_w1565_
	);
	LUT2 #(
		.INIT('h8)
	) name1104 (
		\P1_reg0_reg[4]/NET0131 ,
		_w744_,
		_w1566_
	);
	LUT2 #(
		.INIT('h1)
	) name1105 (
		\P1_reg3_reg[3]/NET0131 ,
		\P1_reg3_reg[4]/NET0131 ,
		_w1567_
	);
	LUT2 #(
		.INIT('h1)
	) name1106 (
		_w716_,
		_w1567_,
		_w1568_
	);
	LUT2 #(
		.INIT('h8)
	) name1107 (
		_w715_,
		_w1568_,
		_w1569_
	);
	LUT2 #(
		.INIT('h1)
	) name1108 (
		_w1564_,
		_w1565_,
		_w1570_
	);
	LUT2 #(
		.INIT('h1)
	) name1109 (
		_w1566_,
		_w1569_,
		_w1571_
	);
	LUT2 #(
		.INIT('h8)
	) name1110 (
		_w1570_,
		_w1571_,
		_w1572_
	);
	LUT2 #(
		.INIT('h8)
	) name1111 (
		\P2_datao_reg[4]/NET0131 ,
		_w543_,
		_w1573_
	);
	LUT2 #(
		.INIT('h1)
	) name1112 (
		_w607_,
		_w623_,
		_w1574_
	);
	LUT2 #(
		.INIT('h4)
	) name1113 (
		_w783_,
		_w1574_,
		_w1575_
	);
	LUT2 #(
		.INIT('h2)
	) name1114 (
		_w783_,
		_w1574_,
		_w1576_
	);
	LUT2 #(
		.INIT('h1)
	) name1115 (
		_w543_,
		_w1575_,
		_w1577_
	);
	LUT2 #(
		.INIT('h4)
	) name1116 (
		_w1576_,
		_w1577_,
		_w1578_
	);
	LUT2 #(
		.INIT('h1)
	) name1117 (
		_w1573_,
		_w1578_,
		_w1579_
	);
	LUT2 #(
		.INIT('h1)
	) name1118 (
		_w538_,
		_w1579_,
		_w1580_
	);
	LUT2 #(
		.INIT('h2)
	) name1119 (
		\P1_IR_reg[31]/NET0131 ,
		_w487_,
		_w1581_
	);
	LUT2 #(
		.INIT('h2)
	) name1120 (
		\P1_IR_reg[4]/NET0131 ,
		_w1581_,
		_w1582_
	);
	LUT2 #(
		.INIT('h4)
	) name1121 (
		\P1_IR_reg[4]/NET0131 ,
		_w1581_,
		_w1583_
	);
	LUT2 #(
		.INIT('h1)
	) name1122 (
		_w1582_,
		_w1583_,
		_w1584_
	);
	LUT2 #(
		.INIT('h2)
	) name1123 (
		_w538_,
		_w1584_,
		_w1585_
	);
	LUT2 #(
		.INIT('h1)
	) name1124 (
		_w1580_,
		_w1585_,
		_w1586_
	);
	LUT2 #(
		.INIT('h2)
	) name1125 (
		_w1572_,
		_w1586_,
		_w1587_
	);
	LUT2 #(
		.INIT('h1)
	) name1126 (
		_w1563_,
		_w1587_,
		_w1588_
	);
	LUT2 #(
		.INIT('h8)
	) name1127 (
		\P1_reg0_reg[2]/NET0131 ,
		_w744_,
		_w1589_
	);
	LUT2 #(
		.INIT('h8)
	) name1128 (
		\P1_reg1_reg[2]/NET0131 ,
		_w746_,
		_w1590_
	);
	LUT2 #(
		.INIT('h8)
	) name1129 (
		\P1_reg2_reg[2]/NET0131 ,
		_w742_,
		_w1591_
	);
	LUT2 #(
		.INIT('h8)
	) name1130 (
		\P1_reg3_reg[2]/NET0131 ,
		_w715_,
		_w1592_
	);
	LUT2 #(
		.INIT('h1)
	) name1131 (
		_w1589_,
		_w1590_,
		_w1593_
	);
	LUT2 #(
		.INIT('h1)
	) name1132 (
		_w1591_,
		_w1592_,
		_w1594_
	);
	LUT2 #(
		.INIT('h8)
	) name1133 (
		_w1593_,
		_w1594_,
		_w1595_
	);
	LUT2 #(
		.INIT('h8)
	) name1134 (
		\P2_datao_reg[2]/NET0131 ,
		_w543_,
		_w1596_
	);
	LUT2 #(
		.INIT('h1)
	) name1135 (
		_w610_,
		_w616_,
		_w1597_
	);
	LUT2 #(
		.INIT('h4)
	) name1136 (
		_w779_,
		_w1597_,
		_w1598_
	);
	LUT2 #(
		.INIT('h2)
	) name1137 (
		_w779_,
		_w1597_,
		_w1599_
	);
	LUT2 #(
		.INIT('h1)
	) name1138 (
		_w543_,
		_w1598_,
		_w1600_
	);
	LUT2 #(
		.INIT('h4)
	) name1139 (
		_w1599_,
		_w1600_,
		_w1601_
	);
	LUT2 #(
		.INIT('h1)
	) name1140 (
		_w1596_,
		_w1601_,
		_w1602_
	);
	LUT2 #(
		.INIT('h1)
	) name1141 (
		_w538_,
		_w1602_,
		_w1603_
	);
	LUT2 #(
		.INIT('h2)
	) name1142 (
		\P1_IR_reg[31]/NET0131 ,
		_w463_,
		_w1604_
	);
	LUT2 #(
		.INIT('h8)
	) name1143 (
		\P1_IR_reg[2]/NET0131 ,
		_w1604_,
		_w1605_
	);
	LUT2 #(
		.INIT('h1)
	) name1144 (
		\P1_IR_reg[2]/NET0131 ,
		_w1604_,
		_w1606_
	);
	LUT2 #(
		.INIT('h1)
	) name1145 (
		_w1605_,
		_w1606_,
		_w1607_
	);
	LUT2 #(
		.INIT('h8)
	) name1146 (
		_w538_,
		_w1607_,
		_w1608_
	);
	LUT2 #(
		.INIT('h1)
	) name1147 (
		_w1603_,
		_w1608_,
		_w1609_
	);
	LUT2 #(
		.INIT('h2)
	) name1148 (
		_w1595_,
		_w1609_,
		_w1610_
	);
	LUT2 #(
		.INIT('h8)
	) name1149 (
		\P1_reg1_reg[3]/NET0131 ,
		_w746_,
		_w1611_
	);
	LUT2 #(
		.INIT('h8)
	) name1150 (
		\P1_reg2_reg[3]/NET0131 ,
		_w742_,
		_w1612_
	);
	LUT2 #(
		.INIT('h8)
	) name1151 (
		\P1_reg0_reg[3]/NET0131 ,
		_w744_,
		_w1613_
	);
	LUT2 #(
		.INIT('h4)
	) name1152 (
		\P1_reg3_reg[3]/NET0131 ,
		_w715_,
		_w1614_
	);
	LUT2 #(
		.INIT('h1)
	) name1153 (
		_w1611_,
		_w1612_,
		_w1615_
	);
	LUT2 #(
		.INIT('h1)
	) name1154 (
		_w1613_,
		_w1614_,
		_w1616_
	);
	LUT2 #(
		.INIT('h8)
	) name1155 (
		_w1615_,
		_w1616_,
		_w1617_
	);
	LUT2 #(
		.INIT('h2)
	) name1156 (
		\P1_IR_reg[31]/NET0131 ,
		_w464_,
		_w1618_
	);
	LUT2 #(
		.INIT('h2)
	) name1157 (
		\P1_IR_reg[3]/NET0131 ,
		_w1618_,
		_w1619_
	);
	LUT2 #(
		.INIT('h4)
	) name1158 (
		\P1_IR_reg[3]/NET0131 ,
		_w1618_,
		_w1620_
	);
	LUT2 #(
		.INIT('h1)
	) name1159 (
		_w1619_,
		_w1620_,
		_w1621_
	);
	LUT2 #(
		.INIT('h2)
	) name1160 (
		_w538_,
		_w1621_,
		_w1622_
	);
	LUT2 #(
		.INIT('h4)
	) name1161 (
		\P2_datao_reg[3]/NET0131 ,
		_w543_,
		_w1623_
	);
	LUT2 #(
		.INIT('h1)
	) name1162 (
		_w610_,
		_w618_,
		_w1624_
	);
	LUT2 #(
		.INIT('h1)
	) name1163 (
		_w608_,
		_w609_,
		_w1625_
	);
	LUT2 #(
		.INIT('h2)
	) name1164 (
		_w1624_,
		_w1625_,
		_w1626_
	);
	LUT2 #(
		.INIT('h4)
	) name1165 (
		_w1624_,
		_w1625_,
		_w1627_
	);
	LUT2 #(
		.INIT('h1)
	) name1166 (
		_w543_,
		_w1626_,
		_w1628_
	);
	LUT2 #(
		.INIT('h4)
	) name1167 (
		_w1627_,
		_w1628_,
		_w1629_
	);
	LUT2 #(
		.INIT('h1)
	) name1168 (
		_w1623_,
		_w1629_,
		_w1630_
	);
	LUT2 #(
		.INIT('h4)
	) name1169 (
		_w538_,
		_w1630_,
		_w1631_
	);
	LUT2 #(
		.INIT('h1)
	) name1170 (
		_w1622_,
		_w1631_,
		_w1632_
	);
	LUT2 #(
		.INIT('h2)
	) name1171 (
		_w1617_,
		_w1632_,
		_w1633_
	);
	LUT2 #(
		.INIT('h1)
	) name1172 (
		_w1610_,
		_w1633_,
		_w1634_
	);
	LUT2 #(
		.INIT('h8)
	) name1173 (
		\P1_reg1_reg[1]/NET0131 ,
		_w746_,
		_w1635_
	);
	LUT2 #(
		.INIT('h8)
	) name1174 (
		\P1_reg0_reg[1]/NET0131 ,
		_w744_,
		_w1636_
	);
	LUT2 #(
		.INIT('h8)
	) name1175 (
		\P1_reg3_reg[1]/NET0131 ,
		_w715_,
		_w1637_
	);
	LUT2 #(
		.INIT('h8)
	) name1176 (
		\P1_reg2_reg[1]/NET0131 ,
		_w742_,
		_w1638_
	);
	LUT2 #(
		.INIT('h1)
	) name1177 (
		_w1635_,
		_w1636_,
		_w1639_
	);
	LUT2 #(
		.INIT('h1)
	) name1178 (
		_w1637_,
		_w1638_,
		_w1640_
	);
	LUT2 #(
		.INIT('h8)
	) name1179 (
		_w1639_,
		_w1640_,
		_w1641_
	);
	LUT2 #(
		.INIT('h8)
	) name1180 (
		\P1_IR_reg[0]/NET0131 ,
		\P1_IR_reg[31]/NET0131 ,
		_w1642_
	);
	LUT2 #(
		.INIT('h1)
	) name1181 (
		\P1_IR_reg[1]/NET0131 ,
		_w1642_,
		_w1643_
	);
	LUT2 #(
		.INIT('h8)
	) name1182 (
		\P1_IR_reg[1]/NET0131 ,
		_w1642_,
		_w1644_
	);
	LUT2 #(
		.INIT('h1)
	) name1183 (
		_w1643_,
		_w1644_,
		_w1645_
	);
	LUT2 #(
		.INIT('h8)
	) name1184 (
		_w538_,
		_w1645_,
		_w1646_
	);
	LUT2 #(
		.INIT('h4)
	) name1185 (
		\P2_datao_reg[1]/NET0131 ,
		_w543_,
		_w1647_
	);
	LUT2 #(
		.INIT('h1)
	) name1186 (
		_w613_,
		_w615_,
		_w1648_
	);
	LUT2 #(
		.INIT('h4)
	) name1187 (
		_w612_,
		_w1648_,
		_w1649_
	);
	LUT2 #(
		.INIT('h2)
	) name1188 (
		_w612_,
		_w1648_,
		_w1650_
	);
	LUT2 #(
		.INIT('h1)
	) name1189 (
		_w543_,
		_w1649_,
		_w1651_
	);
	LUT2 #(
		.INIT('h4)
	) name1190 (
		_w1650_,
		_w1651_,
		_w1652_
	);
	LUT2 #(
		.INIT('h1)
	) name1191 (
		_w1647_,
		_w1652_,
		_w1653_
	);
	LUT2 #(
		.INIT('h4)
	) name1192 (
		_w538_,
		_w1653_,
		_w1654_
	);
	LUT2 #(
		.INIT('h1)
	) name1193 (
		_w1646_,
		_w1654_,
		_w1655_
	);
	LUT2 #(
		.INIT('h4)
	) name1194 (
		_w1641_,
		_w1655_,
		_w1656_
	);
	LUT2 #(
		.INIT('h2)
	) name1195 (
		_w1641_,
		_w1655_,
		_w1657_
	);
	LUT2 #(
		.INIT('h8)
	) name1196 (
		\P1_reg3_reg[0]/NET0131 ,
		_w715_,
		_w1658_
	);
	LUT2 #(
		.INIT('h8)
	) name1197 (
		\P1_reg2_reg[0]/NET0131 ,
		_w742_,
		_w1659_
	);
	LUT2 #(
		.INIT('h8)
	) name1198 (
		\P1_reg0_reg[0]/NET0131 ,
		_w744_,
		_w1660_
	);
	LUT2 #(
		.INIT('h8)
	) name1199 (
		\P1_reg1_reg[0]/NET0131 ,
		_w746_,
		_w1661_
	);
	LUT2 #(
		.INIT('h1)
	) name1200 (
		_w1658_,
		_w1659_,
		_w1662_
	);
	LUT2 #(
		.INIT('h1)
	) name1201 (
		_w1660_,
		_w1661_,
		_w1663_
	);
	LUT2 #(
		.INIT('h8)
	) name1202 (
		_w1662_,
		_w1663_,
		_w1664_
	);
	LUT2 #(
		.INIT('h2)
	) name1203 (
		\si[0]_pad ,
		_w543_,
		_w1665_
	);
	LUT2 #(
		.INIT('h1)
	) name1204 (
		\P2_datao_reg[0]/NET0131 ,
		_w1665_,
		_w1666_
	);
	LUT2 #(
		.INIT('h4)
	) name1205 (
		_w543_,
		_w612_,
		_w1667_
	);
	LUT2 #(
		.INIT('h1)
	) name1206 (
		_w1666_,
		_w1667_,
		_w1668_
	);
	LUT2 #(
		.INIT('h4)
	) name1207 (
		_w538_,
		_w1668_,
		_w1669_
	);
	LUT2 #(
		.INIT('h8)
	) name1208 (
		\P1_IR_reg[0]/NET0131 ,
		_w538_,
		_w1670_
	);
	LUT2 #(
		.INIT('h1)
	) name1209 (
		_w1669_,
		_w1670_,
		_w1671_
	);
	LUT2 #(
		.INIT('h2)
	) name1210 (
		_w1664_,
		_w1671_,
		_w1672_
	);
	LUT2 #(
		.INIT('h1)
	) name1211 (
		_w1657_,
		_w1672_,
		_w1673_
	);
	LUT2 #(
		.INIT('h1)
	) name1212 (
		_w1656_,
		_w1673_,
		_w1674_
	);
	LUT2 #(
		.INIT('h2)
	) name1213 (
		_w1634_,
		_w1674_,
		_w1675_
	);
	LUT2 #(
		.INIT('h4)
	) name1214 (
		_w1617_,
		_w1632_,
		_w1676_
	);
	LUT2 #(
		.INIT('h4)
	) name1215 (
		_w1595_,
		_w1609_,
		_w1677_
	);
	LUT2 #(
		.INIT('h1)
	) name1216 (
		_w1676_,
		_w1677_,
		_w1678_
	);
	LUT2 #(
		.INIT('h1)
	) name1217 (
		_w1633_,
		_w1678_,
		_w1679_
	);
	LUT2 #(
		.INIT('h1)
	) name1218 (
		_w1675_,
		_w1679_,
		_w1680_
	);
	LUT2 #(
		.INIT('h2)
	) name1219 (
		_w1588_,
		_w1680_,
		_w1681_
	);
	LUT2 #(
		.INIT('h4)
	) name1220 (
		_w1548_,
		_w1562_,
		_w1682_
	);
	LUT2 #(
		.INIT('h4)
	) name1221 (
		_w1572_,
		_w1586_,
		_w1683_
	);
	LUT2 #(
		.INIT('h4)
	) name1222 (
		_w1563_,
		_w1683_,
		_w1684_
	);
	LUT2 #(
		.INIT('h1)
	) name1223 (
		_w1682_,
		_w1684_,
		_w1685_
	);
	LUT2 #(
		.INIT('h4)
	) name1224 (
		_w1681_,
		_w1685_,
		_w1686_
	);
	LUT2 #(
		.INIT('h2)
	) name1225 (
		_w1539_,
		_w1686_,
		_w1687_
	);
	LUT2 #(
		.INIT('h4)
	) name1226 (
		_w1498_,
		_w1514_,
		_w1688_
	);
	LUT2 #(
		.INIT('h4)
	) name1227 (
		_w1524_,
		_w1537_,
		_w1689_
	);
	LUT2 #(
		.INIT('h4)
	) name1228 (
		_w1515_,
		_w1689_,
		_w1690_
	);
	LUT2 #(
		.INIT('h1)
	) name1229 (
		_w1688_,
		_w1690_,
		_w1691_
	);
	LUT2 #(
		.INIT('h8)
	) name1230 (
		_w1489_,
		_w1691_,
		_w1692_
	);
	LUT2 #(
		.INIT('h4)
	) name1231 (
		_w1687_,
		_w1692_,
		_w1693_
	);
	LUT2 #(
		.INIT('h4)
	) name1232 (
		_w1297_,
		_w1301_,
		_w1694_
	);
	LUT2 #(
		.INIT('h8)
	) name1233 (
		_w1479_,
		_w1694_,
		_w1695_
	);
	LUT2 #(
		.INIT('h4)
	) name1234 (
		_w1693_,
		_w1695_,
		_w1696_
	);
	LUT2 #(
		.INIT('h1)
	) name1235 (
		_w1327_,
		_w1336_,
		_w1697_
	);
	LUT2 #(
		.INIT('h1)
	) name1236 (
		_w1346_,
		_w1356_,
		_w1698_
	);
	LUT2 #(
		.INIT('h1)
	) name1237 (
		_w1309_,
		_w1318_,
		_w1699_
	);
	LUT2 #(
		.INIT('h1)
	) name1238 (
		_w1698_,
		_w1699_,
		_w1700_
	);
	LUT2 #(
		.INIT('h4)
	) name1239 (
		_w1376_,
		_w1700_,
		_w1701_
	);
	LUT2 #(
		.INIT('h2)
	) name1240 (
		_w1338_,
		_w1701_,
		_w1702_
	);
	LUT2 #(
		.INIT('h1)
	) name1241 (
		_w1697_,
		_w1702_,
		_w1703_
	);
	LUT2 #(
		.INIT('h1)
	) name1242 (
		_w1365_,
		_w1374_,
		_w1704_
	);
	LUT2 #(
		.INIT('h1)
	) name1243 (
		_w1698_,
		_w1704_,
		_w1705_
	);
	LUT2 #(
		.INIT('h1)
	) name1244 (
		_w1357_,
		_w1705_,
		_w1706_
	);
	LUT2 #(
		.INIT('h8)
	) name1245 (
		_w1338_,
		_w1706_,
		_w1707_
	);
	LUT2 #(
		.INIT('h1)
	) name1246 (
		_w1697_,
		_w1699_,
		_w1708_
	);
	LUT2 #(
		.INIT('h1)
	) name1247 (
		_w1337_,
		_w1708_,
		_w1709_
	);
	LUT2 #(
		.INIT('h1)
	) name1248 (
		_w1707_,
		_w1709_,
		_w1710_
	);
	LUT2 #(
		.INIT('h1)
	) name1249 (
		_w1443_,
		_w1452_,
		_w1711_
	);
	LUT2 #(
		.INIT('h1)
	) name1250 (
		_w1466_,
		_w1475_,
		_w1712_
	);
	LUT2 #(
		.INIT('h1)
	) name1251 (
		_w1711_,
		_w1712_,
		_w1713_
	);
	LUT2 #(
		.INIT('h1)
	) name1252 (
		_w1453_,
		_w1713_,
		_w1714_
	);
	LUT2 #(
		.INIT('h8)
	) name1253 (
		_w1429_,
		_w1714_,
		_w1715_
	);
	LUT2 #(
		.INIT('h1)
	) name1254 (
		_w1418_,
		_w1427_,
		_w1716_
	);
	LUT2 #(
		.INIT('h1)
	) name1255 (
		_w1394_,
		_w1403_,
		_w1717_
	);
	LUT2 #(
		.INIT('h1)
	) name1256 (
		_w1716_,
		_w1717_,
		_w1718_
	);
	LUT2 #(
		.INIT('h1)
	) name1257 (
		_w1428_,
		_w1718_,
		_w1719_
	);
	LUT2 #(
		.INIT('h1)
	) name1258 (
		_w1715_,
		_w1719_,
		_w1720_
	);
	LUT2 #(
		.INIT('h8)
	) name1259 (
		_w1710_,
		_w1720_,
		_w1721_
	);
	LUT2 #(
		.INIT('h2)
	) name1260 (
		_w1301_,
		_w1703_,
		_w1722_
	);
	LUT2 #(
		.INIT('h4)
	) name1261 (
		_w1721_,
		_w1722_,
		_w1723_
	);
	LUT2 #(
		.INIT('h1)
	) name1262 (
		_w1069_,
		_w1696_,
		_w1724_
	);
	LUT2 #(
		.INIT('h4)
	) name1263 (
		_w1723_,
		_w1724_,
		_w1725_
	);
	LUT2 #(
		.INIT('h2)
	) name1264 (
		_w951_,
		_w1725_,
		_w1726_
	);
	LUT2 #(
		.INIT('h1)
	) name1265 (
		_w949_,
		_w1726_,
		_w1727_
	);
	LUT2 #(
		.INIT('h1)
	) name1266 (
		_w835_,
		_w837_,
		_w1728_
	);
	LUT2 #(
		.INIT('h4)
	) name1267 (
		_w1727_,
		_w1728_,
		_w1729_
	);
	LUT2 #(
		.INIT('h1)
	) name1268 (
		_w834_,
		_w1729_,
		_w1730_
	);
	LUT2 #(
		.INIT('h4)
	) name1269 (
		_w519_,
		_w1730_,
		_w1731_
	);
	LUT2 #(
		.INIT('h2)
	) name1270 (
		_w519_,
		_w1730_,
		_w1732_
	);
	LUT2 #(
		.INIT('h1)
	) name1271 (
		_w513_,
		_w1731_,
		_w1733_
	);
	LUT2 #(
		.INIT('h4)
	) name1272 (
		_w1732_,
		_w1733_,
		_w1734_
	);
	LUT2 #(
		.INIT('h8)
	) name1273 (
		_w486_,
		_w501_,
		_w1735_
	);
	LUT2 #(
		.INIT('h4)
	) name1274 (
		_w1734_,
		_w1735_,
		_w1736_
	);
	LUT2 #(
		.INIT('h8)
	) name1275 (
		_w692_,
		_w750_,
		_w1737_
	);
	LUT2 #(
		.INIT('h1)
	) name1276 (
		_w832_,
		_w1737_,
		_w1738_
	);
	LUT2 #(
		.INIT('h8)
	) name1277 (
		_w825_,
		_w831_,
		_w1739_
	);
	LUT2 #(
		.INIT('h2)
	) name1278 (
		_w949_,
		_w1739_,
		_w1740_
	);
	LUT2 #(
		.INIT('h2)
	) name1279 (
		_w1738_,
		_w1740_,
		_w1741_
	);
	LUT2 #(
		.INIT('h1)
	) name1280 (
		_w835_,
		_w1741_,
		_w1742_
	);
	LUT2 #(
		.INIT('h8)
	) name1281 (
		_w1539_,
		_w1681_,
		_w1743_
	);
	LUT2 #(
		.INIT('h2)
	) name1282 (
		_w1539_,
		_w1685_,
		_w1744_
	);
	LUT2 #(
		.INIT('h2)
	) name1283 (
		_w1691_,
		_w1744_,
		_w1745_
	);
	LUT2 #(
		.INIT('h4)
	) name1284 (
		_w1743_,
		_w1745_,
		_w1746_
	);
	LUT2 #(
		.INIT('h8)
	) name1285 (
		_w1235_,
		_w1283_,
		_w1747_
	);
	LUT2 #(
		.INIT('h4)
	) name1286 (
		_w1746_,
		_w1747_,
		_w1748_
	);
	LUT2 #(
		.INIT('h8)
	) name1287 (
		_w1480_,
		_w1748_,
		_w1749_
	);
	LUT2 #(
		.INIT('h2)
	) name1288 (
		_w1489_,
		_w1749_,
		_w1750_
	);
	LUT2 #(
		.INIT('h2)
	) name1289 (
		_w1479_,
		_w1750_,
		_w1751_
	);
	LUT2 #(
		.INIT('h2)
	) name1290 (
		_w1377_,
		_w1720_,
		_w1752_
	);
	LUT2 #(
		.INIT('h2)
	) name1291 (
		_w1710_,
		_w1752_,
		_w1753_
	);
	LUT2 #(
		.INIT('h4)
	) name1292 (
		_w1751_,
		_w1753_,
		_w1754_
	);
	LUT2 #(
		.INIT('h2)
	) name1293 (
		_w1301_,
		_w1754_,
		_w1755_
	);
	LUT2 #(
		.INIT('h1)
	) name1294 (
		_w1069_,
		_w1755_,
		_w1756_
	);
	LUT2 #(
		.INIT('h1)
	) name1295 (
		_w835_,
		_w1739_,
		_w1757_
	);
	LUT2 #(
		.INIT('h8)
	) name1296 (
		_w951_,
		_w1757_,
		_w1758_
	);
	LUT2 #(
		.INIT('h4)
	) name1297 (
		_w1756_,
		_w1758_,
		_w1759_
	);
	LUT2 #(
		.INIT('h1)
	) name1298 (
		_w1742_,
		_w1759_,
		_w1760_
	);
	LUT2 #(
		.INIT('h4)
	) name1299 (
		_w501_,
		_w519_,
		_w1761_
	);
	LUT2 #(
		.INIT('h4)
	) name1300 (
		_w486_,
		_w512_,
		_w1762_
	);
	LUT2 #(
		.INIT('h8)
	) name1301 (
		_w1761_,
		_w1762_,
		_w1763_
	);
	LUT2 #(
		.INIT('h4)
	) name1302 (
		_w1760_,
		_w1763_,
		_w1764_
	);
	LUT2 #(
		.INIT('h1)
	) name1303 (
		_w486_,
		_w512_,
		_w1765_
	);
	LUT2 #(
		.INIT('h4)
	) name1304 (
		_w519_,
		_w1765_,
		_w1766_
	);
	LUT2 #(
		.INIT('h4)
	) name1305 (
		_w969_,
		_w978_,
		_w1767_
	);
	LUT2 #(
		.INIT('h2)
	) name1306 (
		_w969_,
		_w978_,
		_w1768_
	);
	LUT2 #(
		.INIT('h1)
	) name1307 (
		_w1767_,
		_w1768_,
		_w1769_
	);
	LUT2 #(
		.INIT('h4)
	) name1308 (
		_w1198_,
		_w1207_,
		_w1770_
	);
	LUT2 #(
		.INIT('h2)
	) name1309 (
		_w1198_,
		_w1207_,
		_w1771_
	);
	LUT2 #(
		.INIT('h1)
	) name1310 (
		_w1770_,
		_w1771_,
		_w1772_
	);
	LUT2 #(
		.INIT('h1)
	) name1311 (
		_w1633_,
		_w1676_,
		_w1773_
	);
	LUT2 #(
		.INIT('h8)
	) name1312 (
		_w1498_,
		_w1514_,
		_w1774_
	);
	LUT2 #(
		.INIT('h1)
	) name1313 (
		_w1498_,
		_w1514_,
		_w1775_
	);
	LUT2 #(
		.INIT('h1)
	) name1314 (
		_w1774_,
		_w1775_,
		_w1776_
	);
	LUT2 #(
		.INIT('h1)
	) name1315 (
		_w1595_,
		_w1609_,
		_w1777_
	);
	LUT2 #(
		.INIT('h8)
	) name1316 (
		_w1595_,
		_w1609_,
		_w1778_
	);
	LUT2 #(
		.INIT('h1)
	) name1317 (
		_w1777_,
		_w1778_,
		_w1779_
	);
	LUT2 #(
		.INIT('h4)
	) name1318 (
		_w1244_,
		_w1257_,
		_w1780_
	);
	LUT2 #(
		.INIT('h2)
	) name1319 (
		_w1244_,
		_w1257_,
		_w1781_
	);
	LUT2 #(
		.INIT('h1)
	) name1320 (
		_w1780_,
		_w1781_,
		_w1782_
	);
	LUT2 #(
		.INIT('h4)
	) name1321 (
		_w1466_,
		_w1475_,
		_w1783_
	);
	LUT2 #(
		.INIT('h2)
	) name1322 (
		_w1466_,
		_w1475_,
		_w1784_
	);
	LUT2 #(
		.INIT('h1)
	) name1323 (
		_w1783_,
		_w1784_,
		_w1785_
	);
	LUT2 #(
		.INIT('h4)
	) name1324 (
		_w1083_,
		_w1094_,
		_w1786_
	);
	LUT2 #(
		.INIT('h2)
	) name1325 (
		_w1083_,
		_w1094_,
		_w1787_
	);
	LUT2 #(
		.INIT('h1)
	) name1326 (
		_w1786_,
		_w1787_,
		_w1788_
	);
	LUT2 #(
		.INIT('h4)
	) name1327 (
		_w1218_,
		_w1233_,
		_w1789_
	);
	LUT2 #(
		.INIT('h2)
	) name1328 (
		_w1218_,
		_w1233_,
		_w1790_
	);
	LUT2 #(
		.INIT('h1)
	) name1329 (
		_w1789_,
		_w1790_,
		_w1791_
	);
	LUT2 #(
		.INIT('h1)
	) name1330 (
		_w1656_,
		_w1657_,
		_w1792_
	);
	LUT2 #(
		.INIT('h1)
	) name1331 (
		_w1538_,
		_w1689_,
		_w1793_
	);
	LUT2 #(
		.INIT('h4)
	) name1332 (
		_w1165_,
		_w1174_,
		_w1794_
	);
	LUT2 #(
		.INIT('h2)
	) name1333 (
		_w1165_,
		_w1174_,
		_w1795_
	);
	LUT2 #(
		.INIT('h1)
	) name1334 (
		_w1794_,
		_w1795_,
		_w1796_
	);
	LUT2 #(
		.INIT('h4)
	) name1335 (
		_w1136_,
		_w1146_,
		_w1797_
	);
	LUT2 #(
		.INIT('h2)
	) name1336 (
		_w1136_,
		_w1146_,
		_w1798_
	);
	LUT2 #(
		.INIT('h1)
	) name1337 (
		_w1797_,
		_w1798_,
		_w1799_
	);
	LUT2 #(
		.INIT('h2)
	) name1338 (
		_w1267_,
		_w1281_,
		_w1800_
	);
	LUT2 #(
		.INIT('h4)
	) name1339 (
		_w1267_,
		_w1281_,
		_w1801_
	);
	LUT2 #(
		.INIT('h1)
	) name1340 (
		_w1800_,
		_w1801_,
		_w1802_
	);
	LUT2 #(
		.INIT('h4)
	) name1341 (
		_w1664_,
		_w1671_,
		_w1803_
	);
	LUT2 #(
		.INIT('h1)
	) name1342 (
		_w1672_,
		_w1803_,
		_w1804_
	);
	LUT2 #(
		.INIT('h1)
	) name1343 (
		_w1563_,
		_w1682_,
		_w1805_
	);
	LUT2 #(
		.INIT('h1)
	) name1344 (
		_w1587_,
		_w1683_,
		_w1806_
	);
	LUT2 #(
		.INIT('h2)
	) name1345 (
		_w997_,
		_w1006_,
		_w1807_
	);
	LUT2 #(
		.INIT('h4)
	) name1346 (
		_w997_,
		_w1006_,
		_w1808_
	);
	LUT2 #(
		.INIT('h1)
	) name1347 (
		_w1807_,
		_w1808_,
		_w1809_
	);
	LUT2 #(
		.INIT('h4)
	) name1348 (
		_w1029_,
		_w1038_,
		_w1810_
	);
	LUT2 #(
		.INIT('h2)
	) name1349 (
		_w1029_,
		_w1038_,
		_w1811_
	);
	LUT2 #(
		.INIT('h1)
	) name1350 (
		_w1810_,
		_w1811_,
		_w1812_
	);
	LUT2 #(
		.INIT('h4)
	) name1351 (
		_w1109_,
		_w1118_,
		_w1813_
	);
	LUT2 #(
		.INIT('h2)
	) name1352 (
		_w1109_,
		_w1118_,
		_w1814_
	);
	LUT2 #(
		.INIT('h1)
	) name1353 (
		_w1813_,
		_w1814_,
		_w1815_
	);
	LUT2 #(
		.INIT('h4)
	) name1354 (
		_w1047_,
		_w1062_,
		_w1816_
	);
	LUT2 #(
		.INIT('h2)
	) name1355 (
		_w1047_,
		_w1062_,
		_w1817_
	);
	LUT2 #(
		.INIT('h1)
	) name1356 (
		_w1816_,
		_w1817_,
		_w1818_
	);
	LUT2 #(
		.INIT('h2)
	) name1357 (
		_w1327_,
		_w1336_,
		_w1819_
	);
	LUT2 #(
		.INIT('h4)
	) name1358 (
		_w1327_,
		_w1336_,
		_w1820_
	);
	LUT2 #(
		.INIT('h1)
	) name1359 (
		_w1819_,
		_w1820_,
		_w1821_
	);
	LUT2 #(
		.INIT('h4)
	) name1360 (
		_w1394_,
		_w1403_,
		_w1822_
	);
	LUT2 #(
		.INIT('h2)
	) name1361 (
		_w1394_,
		_w1403_,
		_w1823_
	);
	LUT2 #(
		.INIT('h1)
	) name1362 (
		_w1822_,
		_w1823_,
		_w1824_
	);
	LUT2 #(
		.INIT('h1)
	) name1363 (
		_w1453_,
		_w1711_,
		_w1825_
	);
	LUT2 #(
		.INIT('h4)
	) name1364 (
		_w1365_,
		_w1374_,
		_w1826_
	);
	LUT2 #(
		.INIT('h2)
	) name1365 (
		_w1365_,
		_w1374_,
		_w1827_
	);
	LUT2 #(
		.INIT('h1)
	) name1366 (
		_w1826_,
		_w1827_,
		_w1828_
	);
	LUT2 #(
		.INIT('h4)
	) name1367 (
		_w933_,
		_w945_,
		_w1829_
	);
	LUT2 #(
		.INIT('h2)
	) name1368 (
		_w933_,
		_w945_,
		_w1830_
	);
	LUT2 #(
		.INIT('h1)
	) name1369 (
		_w1829_,
		_w1830_,
		_w1831_
	);
	LUT2 #(
		.INIT('h1)
	) name1370 (
		_w888_,
		_w947_,
		_w1832_
	);
	LUT2 #(
		.INIT('h4)
	) name1371 (
		_w1418_,
		_w1427_,
		_w1833_
	);
	LUT2 #(
		.INIT('h2)
	) name1372 (
		_w1418_,
		_w1427_,
		_w1834_
	);
	LUT2 #(
		.INIT('h1)
	) name1373 (
		_w1833_,
		_w1834_,
		_w1835_
	);
	LUT2 #(
		.INIT('h4)
	) name1374 (
		_w1309_,
		_w1318_,
		_w1836_
	);
	LUT2 #(
		.INIT('h2)
	) name1375 (
		_w1309_,
		_w1318_,
		_w1837_
	);
	LUT2 #(
		.INIT('h1)
	) name1376 (
		_w1836_,
		_w1837_,
		_w1838_
	);
	LUT2 #(
		.INIT('h4)
	) name1377 (
		_w1346_,
		_w1356_,
		_w1839_
	);
	LUT2 #(
		.INIT('h2)
	) name1378 (
		_w1346_,
		_w1356_,
		_w1840_
	);
	LUT2 #(
		.INIT('h1)
	) name1379 (
		_w1839_,
		_w1840_,
		_w1841_
	);
	LUT2 #(
		.INIT('h2)
	) name1380 (
		_w1773_,
		_w1776_,
		_w1842_
	);
	LUT2 #(
		.INIT('h1)
	) name1381 (
		_w1779_,
		_w1782_,
		_w1843_
	);
	LUT2 #(
		.INIT('h4)
	) name1382 (
		_w1791_,
		_w1792_,
		_w1844_
	);
	LUT2 #(
		.INIT('h2)
	) name1383 (
		_w1793_,
		_w1802_,
		_w1845_
	);
	LUT2 #(
		.INIT('h8)
	) name1384 (
		_w1804_,
		_w1805_,
		_w1846_
	);
	LUT2 #(
		.INIT('h8)
	) name1385 (
		_w1806_,
		_w1846_,
		_w1847_
	);
	LUT2 #(
		.INIT('h8)
	) name1386 (
		_w1844_,
		_w1845_,
		_w1848_
	);
	LUT2 #(
		.INIT('h8)
	) name1387 (
		_w1842_,
		_w1843_,
		_w1849_
	);
	LUT2 #(
		.INIT('h4)
	) name1388 (
		_w1772_,
		_w1849_,
		_w1850_
	);
	LUT2 #(
		.INIT('h8)
	) name1389 (
		_w1847_,
		_w1848_,
		_w1851_
	);
	LUT2 #(
		.INIT('h1)
	) name1390 (
		_w1796_,
		_w1799_,
		_w1852_
	);
	LUT2 #(
		.INIT('h1)
	) name1391 (
		_w1809_,
		_w1812_,
		_w1853_
	);
	LUT2 #(
		.INIT('h4)
	) name1392 (
		_w1815_,
		_w1853_,
		_w1854_
	);
	LUT2 #(
		.INIT('h8)
	) name1393 (
		_w1851_,
		_w1852_,
		_w1855_
	);
	LUT2 #(
		.INIT('h4)
	) name1394 (
		_w1769_,
		_w1850_,
		_w1856_
	);
	LUT2 #(
		.INIT('h1)
	) name1395 (
		_w1785_,
		_w1788_,
		_w1857_
	);
	LUT2 #(
		.INIT('h8)
	) name1396 (
		_w1856_,
		_w1857_,
		_w1858_
	);
	LUT2 #(
		.INIT('h8)
	) name1397 (
		_w1854_,
		_w1855_,
		_w1859_
	);
	LUT2 #(
		.INIT('h4)
	) name1398 (
		_w1824_,
		_w1825_,
		_w1860_
	);
	LUT2 #(
		.INIT('h4)
	) name1399 (
		_w1828_,
		_w1860_,
		_w1861_
	);
	LUT2 #(
		.INIT('h8)
	) name1400 (
		_w1858_,
		_w1859_,
		_w1862_
	);
	LUT2 #(
		.INIT('h1)
	) name1401 (
		_w1835_,
		_w1838_,
		_w1863_
	);
	LUT2 #(
		.INIT('h4)
	) name1402 (
		_w1841_,
		_w1863_,
		_w1864_
	);
	LUT2 #(
		.INIT('h8)
	) name1403 (
		_w1861_,
		_w1862_,
		_w1865_
	);
	LUT2 #(
		.INIT('h1)
	) name1404 (
		_w1818_,
		_w1821_,
		_w1866_
	);
	LUT2 #(
		.INIT('h8)
	) name1405 (
		_w1865_,
		_w1866_,
		_w1867_
	);
	LUT2 #(
		.INIT('h8)
	) name1406 (
		_w1832_,
		_w1864_,
		_w1868_
	);
	LUT2 #(
		.INIT('h8)
	) name1407 (
		_w1867_,
		_w1868_,
		_w1869_
	);
	LUT2 #(
		.INIT('h4)
	) name1408 (
		_w1831_,
		_w1869_,
		_w1870_
	);
	LUT2 #(
		.INIT('h8)
	) name1409 (
		_w1738_,
		_w1757_,
		_w1871_
	);
	LUT2 #(
		.INIT('h8)
	) name1410 (
		_w1870_,
		_w1871_,
		_w1872_
	);
	LUT2 #(
		.INIT('h8)
	) name1411 (
		_w501_,
		_w1872_,
		_w1873_
	);
	LUT2 #(
		.INIT('h1)
	) name1412 (
		\P1_B_reg/NET0131 ,
		_w1873_,
		_w1874_
	);
	LUT2 #(
		.INIT('h2)
	) name1413 (
		_w1766_,
		_w1874_,
		_w1875_
	);
	LUT2 #(
		.INIT('h4)
	) name1414 (
		\P1_B_reg/NET0131 ,
		_w1872_,
		_w1876_
	);
	LUT2 #(
		.INIT('h8)
	) name1415 (
		_w519_,
		_w1765_,
		_w1877_
	);
	LUT2 #(
		.INIT('h8)
	) name1416 (
		_w501_,
		_w1877_,
		_w1878_
	);
	LUT2 #(
		.INIT('h4)
	) name1417 (
		_w1876_,
		_w1878_,
		_w1879_
	);
	LUT2 #(
		.INIT('h8)
	) name1418 (
		_w501_,
		_w1762_,
		_w1880_
	);
	LUT2 #(
		.INIT('h1)
	) name1419 (
		_w519_,
		_w1872_,
		_w1881_
	);
	LUT2 #(
		.INIT('h8)
	) name1420 (
		_w519_,
		_w1872_,
		_w1882_
	);
	LUT2 #(
		.INIT('h2)
	) name1421 (
		_w1880_,
		_w1881_,
		_w1883_
	);
	LUT2 #(
		.INIT('h4)
	) name1422 (
		_w1882_,
		_w1883_,
		_w1884_
	);
	LUT2 #(
		.INIT('h1)
	) name1423 (
		_w501_,
		_w519_,
		_w1885_
	);
	LUT2 #(
		.INIT('h4)
	) name1424 (
		_w486_,
		_w1885_,
		_w1886_
	);
	LUT2 #(
		.INIT('h8)
	) name1425 (
		_w1760_,
		_w1886_,
		_w1887_
	);
	LUT2 #(
		.INIT('h8)
	) name1426 (
		_w486_,
		_w512_,
		_w1888_
	);
	LUT2 #(
		.INIT('h1)
	) name1427 (
		_w1007_,
		_w1064_,
		_w1889_
	);
	LUT2 #(
		.INIT('h4)
	) name1428 (
		_w1300_,
		_w1889_,
		_w1890_
	);
	LUT2 #(
		.INIT('h2)
	) name1429 (
		_w1298_,
		_w1890_,
		_w1891_
	);
	LUT2 #(
		.INIT('h1)
	) name1430 (
		_w946_,
		_w1008_,
		_w1892_
	);
	LUT2 #(
		.INIT('h4)
	) name1431 (
		_w1891_,
		_w1892_,
		_w1893_
	);
	LUT2 #(
		.INIT('h2)
	) name1432 (
		_w951_,
		_w1893_,
		_w1894_
	);
	LUT2 #(
		.INIT('h1)
	) name1433 (
		_w947_,
		_w1894_,
		_w1895_
	);
	LUT2 #(
		.INIT('h1)
	) name1434 (
		_w1682_,
		_w1689_,
		_w1896_
	);
	LUT2 #(
		.INIT('h1)
	) name1435 (
		_w1676_,
		_w1683_,
		_w1897_
	);
	LUT2 #(
		.INIT('h4)
	) name1436 (
		_w1657_,
		_w1803_,
		_w1898_
	);
	LUT2 #(
		.INIT('h1)
	) name1437 (
		_w1656_,
		_w1677_,
		_w1899_
	);
	LUT2 #(
		.INIT('h4)
	) name1438 (
		_w1898_,
		_w1899_,
		_w1900_
	);
	LUT2 #(
		.INIT('h2)
	) name1439 (
		_w1634_,
		_w1900_,
		_w1901_
	);
	LUT2 #(
		.INIT('h2)
	) name1440 (
		_w1897_,
		_w1901_,
		_w1902_
	);
	LUT2 #(
		.INIT('h2)
	) name1441 (
		_w1588_,
		_w1902_,
		_w1903_
	);
	LUT2 #(
		.INIT('h2)
	) name1442 (
		_w1896_,
		_w1903_,
		_w1904_
	);
	LUT2 #(
		.INIT('h2)
	) name1443 (
		_w1539_,
		_w1904_,
		_w1905_
	);
	LUT2 #(
		.INIT('h2)
	) name1444 (
		_w1482_,
		_w1688_,
		_w1906_
	);
	LUT2 #(
		.INIT('h8)
	) name1445 (
		_w1485_,
		_w1906_,
		_w1907_
	);
	LUT2 #(
		.INIT('h8)
	) name1446 (
		_w1176_,
		_w1907_,
		_w1908_
	);
	LUT2 #(
		.INIT('h8)
	) name1447 (
		_w1181_,
		_w1908_,
		_w1909_
	);
	LUT2 #(
		.INIT('h4)
	) name1448 (
		_w1905_,
		_w1909_,
		_w1910_
	);
	LUT2 #(
		.INIT('h1)
	) name1449 (
		_w1297_,
		_w1910_,
		_w1911_
	);
	LUT2 #(
		.INIT('h8)
	) name1450 (
		_w1705_,
		_w1708_,
		_w1912_
	);
	LUT2 #(
		.INIT('h8)
	) name1451 (
		_w1713_,
		_w1718_,
		_w1913_
	);
	LUT2 #(
		.INIT('h8)
	) name1452 (
		_w1912_,
		_w1913_,
		_w1914_
	);
	LUT2 #(
		.INIT('h4)
	) name1453 (
		_w1911_,
		_w1914_,
		_w1915_
	);
	LUT2 #(
		.INIT('h1)
	) name1454 (
		_w1711_,
		_w1717_,
		_w1916_
	);
	LUT2 #(
		.INIT('h4)
	) name1455 (
		_w1477_,
		_w1916_,
		_w1917_
	);
	LUT2 #(
		.INIT('h2)
	) name1456 (
		_w1429_,
		_w1917_,
		_w1918_
	);
	LUT2 #(
		.INIT('h1)
	) name1457 (
		_w1716_,
		_w1918_,
		_w1919_
	);
	LUT2 #(
		.INIT('h8)
	) name1458 (
		_w1912_,
		_w1919_,
		_w1920_
	);
	LUT2 #(
		.INIT('h1)
	) name1459 (
		_w1703_,
		_w1920_,
		_w1921_
	);
	LUT2 #(
		.INIT('h4)
	) name1460 (
		_w1915_,
		_w1921_,
		_w1922_
	);
	LUT2 #(
		.INIT('h8)
	) name1461 (
		_w1009_,
		_w1065_,
		_w1923_
	);
	LUT2 #(
		.INIT('h8)
	) name1462 (
		_w948_,
		_w1923_,
		_w1924_
	);
	LUT2 #(
		.INIT('h4)
	) name1463 (
		_w1922_,
		_w1924_,
		_w1925_
	);
	LUT2 #(
		.INIT('h1)
	) name1464 (
		_w1895_,
		_w1925_,
		_w1926_
	);
	LUT2 #(
		.INIT('h1)
	) name1465 (
		_w832_,
		_w1926_,
		_w1927_
	);
	LUT2 #(
		.INIT('h2)
	) name1466 (
		_w1757_,
		_w1927_,
		_w1928_
	);
	LUT2 #(
		.INIT('h1)
	) name1467 (
		_w1737_,
		_w1928_,
		_w1929_
	);
	LUT2 #(
		.INIT('h1)
	) name1468 (
		_w1761_,
		_w1929_,
		_w1930_
	);
	LUT2 #(
		.INIT('h4)
	) name1469 (
		_w1885_,
		_w1929_,
		_w1931_
	);
	LUT2 #(
		.INIT('h2)
	) name1470 (
		_w1888_,
		_w1930_,
		_w1932_
	);
	LUT2 #(
		.INIT('h4)
	) name1471 (
		_w1931_,
		_w1932_,
		_w1933_
	);
	LUT2 #(
		.INIT('h1)
	) name1472 (
		\P1_B_reg/NET0131 ,
		_w1929_,
		_w1934_
	);
	LUT2 #(
		.INIT('h2)
	) name1473 (
		_w486_,
		_w512_,
		_w1935_
	);
	LUT2 #(
		.INIT('h8)
	) name1474 (
		_w1885_,
		_w1935_,
		_w1936_
	);
	LUT2 #(
		.INIT('h4)
	) name1475 (
		_w1934_,
		_w1936_,
		_w1937_
	);
	LUT2 #(
		.INIT('h4)
	) name1476 (
		\P1_B_reg/NET0131 ,
		_w1929_,
		_w1938_
	);
	LUT2 #(
		.INIT('h8)
	) name1477 (
		_w1761_,
		_w1935_,
		_w1939_
	);
	LUT2 #(
		.INIT('h4)
	) name1478 (
		_w1938_,
		_w1939_,
		_w1940_
	);
	LUT2 #(
		.INIT('h4)
	) name1479 (
		\P1_B_reg/NET0131 ,
		_w1760_,
		_w1941_
	);
	LUT2 #(
		.INIT('h8)
	) name1480 (
		_w1761_,
		_w1765_,
		_w1942_
	);
	LUT2 #(
		.INIT('h4)
	) name1481 (
		_w1941_,
		_w1942_,
		_w1943_
	);
	LUT2 #(
		.INIT('h1)
	) name1482 (
		_w1875_,
		_w1879_,
		_w1944_
	);
	LUT2 #(
		.INIT('h4)
	) name1483 (
		_w1884_,
		_w1944_,
		_w1945_
	);
	LUT2 #(
		.INIT('h4)
	) name1484 (
		_w1764_,
		_w1945_,
		_w1946_
	);
	LUT2 #(
		.INIT('h4)
	) name1485 (
		_w1887_,
		_w1946_,
		_w1947_
	);
	LUT2 #(
		.INIT('h1)
	) name1486 (
		_w1937_,
		_w1940_,
		_w1948_
	);
	LUT2 #(
		.INIT('h4)
	) name1487 (
		_w1943_,
		_w1948_,
		_w1949_
	);
	LUT2 #(
		.INIT('h4)
	) name1488 (
		_w1933_,
		_w1947_,
		_w1950_
	);
	LUT2 #(
		.INIT('h8)
	) name1489 (
		_w1949_,
		_w1950_,
		_w1951_
	);
	LUT2 #(
		.INIT('h4)
	) name1490 (
		_w1736_,
		_w1951_,
		_w1952_
	);
	LUT2 #(
		.INIT('h2)
	) name1491 (
		\P1_state_reg[0]/NET0131 ,
		_w512_,
		_w1953_
	);
	LUT2 #(
		.INIT('h4)
	) name1492 (
		_w1952_,
		_w1953_,
		_w1954_
	);
	LUT2 #(
		.INIT('h2)
	) name1493 (
		\P1_B_reg/NET0131 ,
		_w1953_,
		_w1955_
	);
	LUT2 #(
		.INIT('h1)
	) name1494 (
		_w1954_,
		_w1955_,
		_w1956_
	);
	LUT2 #(
		.INIT('h1)
	) name1495 (
		\P2_IR_reg[20]/NET0131 ,
		\P2_IR_reg[21]/NET0131 ,
		_w1957_
	);
	LUT2 #(
		.INIT('h4)
	) name1496 (
		\P2_IR_reg[22]/NET0131 ,
		_w1957_,
		_w1958_
	);
	LUT2 #(
		.INIT('h1)
	) name1497 (
		\P2_IR_reg[10]/NET0131 ,
		\P2_IR_reg[11]/NET0131 ,
		_w1959_
	);
	LUT2 #(
		.INIT('h4)
	) name1498 (
		\P2_IR_reg[12]/NET0131 ,
		_w1959_,
		_w1960_
	);
	LUT2 #(
		.INIT('h1)
	) name1499 (
		\P2_IR_reg[0]/NET0131 ,
		\P2_IR_reg[1]/NET0131 ,
		_w1961_
	);
	LUT2 #(
		.INIT('h4)
	) name1500 (
		\P2_IR_reg[2]/NET0131 ,
		_w1961_,
		_w1962_
	);
	LUT2 #(
		.INIT('h1)
	) name1501 (
		\P2_IR_reg[3]/NET0131 ,
		\P2_IR_reg[4]/NET0131 ,
		_w1963_
	);
	LUT2 #(
		.INIT('h8)
	) name1502 (
		_w1962_,
		_w1963_,
		_w1964_
	);
	LUT2 #(
		.INIT('h1)
	) name1503 (
		\P2_IR_reg[5]/NET0131 ,
		\P2_IR_reg[6]/NET0131 ,
		_w1965_
	);
	LUT2 #(
		.INIT('h4)
	) name1504 (
		\P2_IR_reg[7]/NET0131 ,
		_w1965_,
		_w1966_
	);
	LUT2 #(
		.INIT('h1)
	) name1505 (
		\P2_IR_reg[8]/NET0131 ,
		\P2_IR_reg[9]/NET0131 ,
		_w1967_
	);
	LUT2 #(
		.INIT('h8)
	) name1506 (
		_w1966_,
		_w1967_,
		_w1968_
	);
	LUT2 #(
		.INIT('h8)
	) name1507 (
		_w1964_,
		_w1968_,
		_w1969_
	);
	LUT2 #(
		.INIT('h4)
	) name1508 (
		\P2_IR_reg[13]/NET0131 ,
		_w1960_,
		_w1970_
	);
	LUT2 #(
		.INIT('h8)
	) name1509 (
		_w1969_,
		_w1970_,
		_w1971_
	);
	LUT2 #(
		.INIT('h4)
	) name1510 (
		\P2_IR_reg[14]/NET0131 ,
		_w1971_,
		_w1972_
	);
	LUT2 #(
		.INIT('h4)
	) name1511 (
		\P2_IR_reg[15]/NET0131 ,
		_w1972_,
		_w1973_
	);
	LUT2 #(
		.INIT('h1)
	) name1512 (
		\P2_IR_reg[16]/NET0131 ,
		\P2_IR_reg[17]/NET0131 ,
		_w1974_
	);
	LUT2 #(
		.INIT('h4)
	) name1513 (
		\P2_IR_reg[18]/NET0131 ,
		_w1974_,
		_w1975_
	);
	LUT2 #(
		.INIT('h8)
	) name1514 (
		_w1973_,
		_w1975_,
		_w1976_
	);
	LUT2 #(
		.INIT('h4)
	) name1515 (
		\P2_IR_reg[19]/NET0131 ,
		_w1958_,
		_w1977_
	);
	LUT2 #(
		.INIT('h8)
	) name1516 (
		_w1976_,
		_w1977_,
		_w1978_
	);
	LUT2 #(
		.INIT('h2)
	) name1517 (
		\P2_IR_reg[31]/NET0131 ,
		_w1978_,
		_w1979_
	);
	LUT2 #(
		.INIT('h1)
	) name1518 (
		\P2_IR_reg[23]/NET0131 ,
		_w1979_,
		_w1980_
	);
	LUT2 #(
		.INIT('h8)
	) name1519 (
		\P2_IR_reg[23]/NET0131 ,
		_w1979_,
		_w1981_
	);
	LUT2 #(
		.INIT('h1)
	) name1520 (
		_w1980_,
		_w1981_,
		_w1982_
	);
	LUT2 #(
		.INIT('h2)
	) name1521 (
		\P1_state_reg[0]/NET0131 ,
		_w1982_,
		_w1983_
	);
	LUT2 #(
		.INIT('h2)
	) name1522 (
		\P2_reg0_reg[29]/NET0131 ,
		_w1983_,
		_w1984_
	);
	LUT2 #(
		.INIT('h1)
	) name1523 (
		\P2_IR_reg[23]/NET0131 ,
		\P2_IR_reg[24]/NET0131 ,
		_w1985_
	);
	LUT2 #(
		.INIT('h4)
	) name1524 (
		\P2_IR_reg[22]/NET0131 ,
		_w1985_,
		_w1986_
	);
	LUT2 #(
		.INIT('h1)
	) name1525 (
		\P2_IR_reg[13]/NET0131 ,
		\P2_IR_reg[14]/NET0131 ,
		_w1987_
	);
	LUT2 #(
		.INIT('h1)
	) name1526 (
		\P2_IR_reg[15]/NET0131 ,
		\P2_IR_reg[16]/NET0131 ,
		_w1988_
	);
	LUT2 #(
		.INIT('h8)
	) name1527 (
		_w1987_,
		_w1988_,
		_w1989_
	);
	LUT2 #(
		.INIT('h4)
	) name1528 (
		\P2_IR_reg[17]/NET0131 ,
		_w1989_,
		_w1990_
	);
	LUT2 #(
		.INIT('h8)
	) name1529 (
		_w1960_,
		_w1990_,
		_w1991_
	);
	LUT2 #(
		.INIT('h8)
	) name1530 (
		_w1969_,
		_w1991_,
		_w1992_
	);
	LUT2 #(
		.INIT('h1)
	) name1531 (
		\P2_IR_reg[18]/NET0131 ,
		\P2_IR_reg[19]/NET0131 ,
		_w1993_
	);
	LUT2 #(
		.INIT('h8)
	) name1532 (
		_w1957_,
		_w1993_,
		_w1994_
	);
	LUT2 #(
		.INIT('h8)
	) name1533 (
		_w1992_,
		_w1994_,
		_w1995_
	);
	LUT2 #(
		.INIT('h4)
	) name1534 (
		\P2_IR_reg[25]/NET0131 ,
		_w1986_,
		_w1996_
	);
	LUT2 #(
		.INIT('h8)
	) name1535 (
		_w1995_,
		_w1996_,
		_w1997_
	);
	LUT2 #(
		.INIT('h2)
	) name1536 (
		\P2_IR_reg[31]/NET0131 ,
		_w1997_,
		_w1998_
	);
	LUT2 #(
		.INIT('h8)
	) name1537 (
		\P2_IR_reg[26]/NET0131 ,
		_w1998_,
		_w1999_
	);
	LUT2 #(
		.INIT('h1)
	) name1538 (
		\P2_IR_reg[26]/NET0131 ,
		_w1998_,
		_w2000_
	);
	LUT2 #(
		.INIT('h1)
	) name1539 (
		_w1999_,
		_w2000_,
		_w2001_
	);
	LUT2 #(
		.INIT('h8)
	) name1540 (
		_w1992_,
		_w1993_,
		_w2002_
	);
	LUT2 #(
		.INIT('h4)
	) name1541 (
		\P2_IR_reg[23]/NET0131 ,
		_w1958_,
		_w2003_
	);
	LUT2 #(
		.INIT('h8)
	) name1542 (
		_w2002_,
		_w2003_,
		_w2004_
	);
	LUT2 #(
		.INIT('h2)
	) name1543 (
		\P2_IR_reg[31]/NET0131 ,
		_w2004_,
		_w2005_
	);
	LUT2 #(
		.INIT('h1)
	) name1544 (
		\P2_IR_reg[24]/NET0131 ,
		_w2005_,
		_w2006_
	);
	LUT2 #(
		.INIT('h8)
	) name1545 (
		\P2_IR_reg[24]/NET0131 ,
		_w2005_,
		_w2007_
	);
	LUT2 #(
		.INIT('h1)
	) name1546 (
		_w2006_,
		_w2007_,
		_w2008_
	);
	LUT2 #(
		.INIT('h8)
	) name1547 (
		_w2001_,
		_w2008_,
		_w2009_
	);
	LUT2 #(
		.INIT('h4)
	) name1548 (
		\P2_IR_reg[8]/NET0131 ,
		_w1966_,
		_w2010_
	);
	LUT2 #(
		.INIT('h8)
	) name1549 (
		_w1964_,
		_w2010_,
		_w2011_
	);
	LUT2 #(
		.INIT('h4)
	) name1550 (
		\P2_IR_reg[9]/NET0131 ,
		_w1960_,
		_w2012_
	);
	LUT2 #(
		.INIT('h8)
	) name1551 (
		_w2011_,
		_w2012_,
		_w2013_
	);
	LUT2 #(
		.INIT('h4)
	) name1552 (
		\P2_IR_reg[20]/NET0131 ,
		_w1993_,
		_w2014_
	);
	LUT2 #(
		.INIT('h8)
	) name1553 (
		_w1990_,
		_w2014_,
		_w2015_
	);
	LUT2 #(
		.INIT('h8)
	) name1554 (
		_w2013_,
		_w2015_,
		_w2016_
	);
	LUT2 #(
		.INIT('h4)
	) name1555 (
		\P2_IR_reg[21]/NET0131 ,
		_w1986_,
		_w2017_
	);
	LUT2 #(
		.INIT('h8)
	) name1556 (
		_w2016_,
		_w2017_,
		_w2018_
	);
	LUT2 #(
		.INIT('h2)
	) name1557 (
		\P2_IR_reg[31]/NET0131 ,
		_w2018_,
		_w2019_
	);
	LUT2 #(
		.INIT('h8)
	) name1558 (
		\P2_IR_reg[25]/NET0131 ,
		_w2019_,
		_w2020_
	);
	LUT2 #(
		.INIT('h1)
	) name1559 (
		\P2_IR_reg[25]/NET0131 ,
		_w2019_,
		_w2021_
	);
	LUT2 #(
		.INIT('h1)
	) name1560 (
		_w2020_,
		_w2021_,
		_w2022_
	);
	LUT2 #(
		.INIT('h8)
	) name1561 (
		_w2009_,
		_w2022_,
		_w2023_
	);
	LUT2 #(
		.INIT('h4)
	) name1562 (
		_w1982_,
		_w2023_,
		_w2024_
	);
	LUT2 #(
		.INIT('h8)
	) name1563 (
		\P2_reg0_reg[29]/NET0131 ,
		_w2024_,
		_w2025_
	);
	LUT2 #(
		.INIT('h1)
	) name1564 (
		_w1982_,
		_w2023_,
		_w2026_
	);
	LUT2 #(
		.INIT('h2)
	) name1565 (
		\P2_B_reg/NET0131 ,
		_w2008_,
		_w2027_
	);
	LUT2 #(
		.INIT('h4)
	) name1566 (
		_w2022_,
		_w2027_,
		_w2028_
	);
	LUT2 #(
		.INIT('h1)
	) name1567 (
		\P2_d_reg[1]/NET0131 ,
		_w2028_,
		_w2029_
	);
	LUT2 #(
		.INIT('h2)
	) name1568 (
		_w2001_,
		_w2029_,
		_w2030_
	);
	LUT2 #(
		.INIT('h1)
	) name1569 (
		\P2_B_reg/NET0131 ,
		_w2022_,
		_w2031_
	);
	LUT2 #(
		.INIT('h2)
	) name1570 (
		_w2001_,
		_w2031_,
		_w2032_
	);
	LUT2 #(
		.INIT('h1)
	) name1571 (
		_w2009_,
		_w2022_,
		_w2033_
	);
	LUT2 #(
		.INIT('h1)
	) name1572 (
		_w2032_,
		_w2033_,
		_w2034_
	);
	LUT2 #(
		.INIT('h1)
	) name1573 (
		_w2030_,
		_w2034_,
		_w2035_
	);
	LUT2 #(
		.INIT('h1)
	) name1574 (
		\P2_d_reg[0]/NET0131 ,
		_w2028_,
		_w2036_
	);
	LUT2 #(
		.INIT('h2)
	) name1575 (
		_w2001_,
		_w2036_,
		_w2037_
	);
	LUT2 #(
		.INIT('h2)
	) name1576 (
		_w2008_,
		_w2032_,
		_w2038_
	);
	LUT2 #(
		.INIT('h1)
	) name1577 (
		_w2037_,
		_w2038_,
		_w2039_
	);
	LUT2 #(
		.INIT('h8)
	) name1578 (
		_w2035_,
		_w2039_,
		_w2040_
	);
	LUT2 #(
		.INIT('h2)
	) name1579 (
		\P2_reg0_reg[29]/NET0131 ,
		_w2040_,
		_w2041_
	);
	LUT2 #(
		.INIT('h2)
	) name1580 (
		\P2_IR_reg[31]/NET0131 ,
		_w2002_,
		_w2042_
	);
	LUT2 #(
		.INIT('h1)
	) name1581 (
		\P2_IR_reg[25]/NET0131 ,
		\P2_IR_reg[26]/NET0131 ,
		_w2043_
	);
	LUT2 #(
		.INIT('h8)
	) name1582 (
		_w1985_,
		_w2043_,
		_w2044_
	);
	LUT2 #(
		.INIT('h4)
	) name1583 (
		\P2_IR_reg[22]/NET0131 ,
		_w2044_,
		_w2045_
	);
	LUT2 #(
		.INIT('h8)
	) name1584 (
		_w1957_,
		_w2045_,
		_w2046_
	);
	LUT2 #(
		.INIT('h2)
	) name1585 (
		\P2_IR_reg[31]/NET0131 ,
		_w2046_,
		_w2047_
	);
	LUT2 #(
		.INIT('h1)
	) name1586 (
		_w2042_,
		_w2047_,
		_w2048_
	);
	LUT2 #(
		.INIT('h2)
	) name1587 (
		\P2_IR_reg[27]/NET0131 ,
		_w2048_,
		_w2049_
	);
	LUT2 #(
		.INIT('h4)
	) name1588 (
		\P2_IR_reg[27]/NET0131 ,
		_w2048_,
		_w2050_
	);
	LUT2 #(
		.INIT('h1)
	) name1589 (
		_w2049_,
		_w2050_,
		_w2051_
	);
	LUT2 #(
		.INIT('h1)
	) name1590 (
		\P2_IR_reg[24]/NET0131 ,
		\P2_IR_reg[27]/NET0131 ,
		_w2052_
	);
	LUT2 #(
		.INIT('h8)
	) name1591 (
		_w2043_,
		_w2052_,
		_w2053_
	);
	LUT2 #(
		.INIT('h2)
	) name1592 (
		\P2_IR_reg[31]/NET0131 ,
		_w2053_,
		_w2054_
	);
	LUT2 #(
		.INIT('h1)
	) name1593 (
		_w2005_,
		_w2054_,
		_w2055_
	);
	LUT2 #(
		.INIT('h2)
	) name1594 (
		\P2_IR_reg[28]/NET0131 ,
		_w2055_,
		_w2056_
	);
	LUT2 #(
		.INIT('h4)
	) name1595 (
		\P2_IR_reg[28]/NET0131 ,
		_w2055_,
		_w2057_
	);
	LUT2 #(
		.INIT('h1)
	) name1596 (
		_w2056_,
		_w2057_,
		_w2058_
	);
	LUT2 #(
		.INIT('h1)
	) name1597 (
		_w2051_,
		_w2058_,
		_w2059_
	);
	LUT2 #(
		.INIT('h2)
	) name1598 (
		\P1_datao_reg[29]/NET0131 ,
		_w543_,
		_w2060_
	);
	LUT2 #(
		.INIT('h8)
	) name1599 (
		\P1_datao_reg[29]/NET0131 ,
		\si[29]_pad ,
		_w2061_
	);
	LUT2 #(
		.INIT('h1)
	) name1600 (
		\P1_datao_reg[29]/NET0131 ,
		\si[29]_pad ,
		_w2062_
	);
	LUT2 #(
		.INIT('h1)
	) name1601 (
		_w2061_,
		_w2062_,
		_w2063_
	);
	LUT2 #(
		.INIT('h1)
	) name1602 (
		\P1_datao_reg[28]/NET0131 ,
		\si[28]_pad ,
		_w2064_
	);
	LUT2 #(
		.INIT('h1)
	) name1603 (
		\P1_datao_reg[23]/NET0131 ,
		\si[23]_pad ,
		_w2065_
	);
	LUT2 #(
		.INIT('h1)
	) name1604 (
		\P1_datao_reg[24]/NET0131 ,
		\si[24]_pad ,
		_w2066_
	);
	LUT2 #(
		.INIT('h1)
	) name1605 (
		_w2065_,
		_w2066_,
		_w2067_
	);
	LUT2 #(
		.INIT('h1)
	) name1606 (
		\P1_datao_reg[22]/NET0131 ,
		\si[22]_pad ,
		_w2068_
	);
	LUT2 #(
		.INIT('h1)
	) name1607 (
		\P1_datao_reg[21]/NET0131 ,
		\si[21]_pad ,
		_w2069_
	);
	LUT2 #(
		.INIT('h1)
	) name1608 (
		_w2068_,
		_w2069_,
		_w2070_
	);
	LUT2 #(
		.INIT('h8)
	) name1609 (
		_w2067_,
		_w2070_,
		_w2071_
	);
	LUT2 #(
		.INIT('h1)
	) name1610 (
		\P1_datao_reg[27]/NET0131 ,
		\si[27]_pad ,
		_w2072_
	);
	LUT2 #(
		.INIT('h1)
	) name1611 (
		\P1_datao_reg[26]/NET0131 ,
		\si[26]_pad ,
		_w2073_
	);
	LUT2 #(
		.INIT('h1)
	) name1612 (
		\P1_datao_reg[25]/NET0131 ,
		\si[25]_pad ,
		_w2074_
	);
	LUT2 #(
		.INIT('h1)
	) name1613 (
		_w2073_,
		_w2074_,
		_w2075_
	);
	LUT2 #(
		.INIT('h4)
	) name1614 (
		_w2072_,
		_w2075_,
		_w2076_
	);
	LUT2 #(
		.INIT('h1)
	) name1615 (
		\P1_datao_reg[17]/NET0131 ,
		\si[17]_pad ,
		_w2077_
	);
	LUT2 #(
		.INIT('h1)
	) name1616 (
		\P1_datao_reg[20]/NET0131 ,
		\si[20]_pad ,
		_w2078_
	);
	LUT2 #(
		.INIT('h1)
	) name1617 (
		\P1_datao_reg[18]/NET0131 ,
		\si[18]_pad ,
		_w2079_
	);
	LUT2 #(
		.INIT('h1)
	) name1618 (
		\P1_datao_reg[19]/NET0131 ,
		\si[19]_pad ,
		_w2080_
	);
	LUT2 #(
		.INIT('h1)
	) name1619 (
		_w2079_,
		_w2080_,
		_w2081_
	);
	LUT2 #(
		.INIT('h4)
	) name1620 (
		_w2078_,
		_w2081_,
		_w2082_
	);
	LUT2 #(
		.INIT('h4)
	) name1621 (
		_w2077_,
		_w2082_,
		_w2083_
	);
	LUT2 #(
		.INIT('h1)
	) name1622 (
		\P1_datao_reg[16]/NET0131 ,
		\si[16]_pad ,
		_w2084_
	);
	LUT2 #(
		.INIT('h8)
	) name1623 (
		\P1_datao_reg[15]/NET0131 ,
		\si[15]_pad ,
		_w2085_
	);
	LUT2 #(
		.INIT('h8)
	) name1624 (
		\P1_datao_reg[16]/NET0131 ,
		\si[16]_pad ,
		_w2086_
	);
	LUT2 #(
		.INIT('h1)
	) name1625 (
		_w2085_,
		_w2086_,
		_w2087_
	);
	LUT2 #(
		.INIT('h1)
	) name1626 (
		\P1_datao_reg[14]/NET0131 ,
		\si[14]_pad ,
		_w2088_
	);
	LUT2 #(
		.INIT('h1)
	) name1627 (
		\P1_datao_reg[15]/NET0131 ,
		\si[15]_pad ,
		_w2089_
	);
	LUT2 #(
		.INIT('h1)
	) name1628 (
		_w2088_,
		_w2089_,
		_w2090_
	);
	LUT2 #(
		.INIT('h8)
	) name1629 (
		\P1_datao_reg[13]/NET0131 ,
		\si[13]_pad ,
		_w2091_
	);
	LUT2 #(
		.INIT('h8)
	) name1630 (
		\P1_datao_reg[14]/NET0131 ,
		\si[14]_pad ,
		_w2092_
	);
	LUT2 #(
		.INIT('h1)
	) name1631 (
		_w2091_,
		_w2092_,
		_w2093_
	);
	LUT2 #(
		.INIT('h2)
	) name1632 (
		_w2090_,
		_w2093_,
		_w2094_
	);
	LUT2 #(
		.INIT('h2)
	) name1633 (
		_w2087_,
		_w2094_,
		_w2095_
	);
	LUT2 #(
		.INIT('h1)
	) name1634 (
		_w2084_,
		_w2095_,
		_w2096_
	);
	LUT2 #(
		.INIT('h8)
	) name1635 (
		_w2083_,
		_w2096_,
		_w2097_
	);
	LUT2 #(
		.INIT('h8)
	) name1636 (
		\P1_datao_reg[19]/NET0131 ,
		\si[19]_pad ,
		_w2098_
	);
	LUT2 #(
		.INIT('h8)
	) name1637 (
		\P1_datao_reg[20]/NET0131 ,
		\si[20]_pad ,
		_w2099_
	);
	LUT2 #(
		.INIT('h1)
	) name1638 (
		_w2098_,
		_w2099_,
		_w2100_
	);
	LUT2 #(
		.INIT('h1)
	) name1639 (
		_w2078_,
		_w2100_,
		_w2101_
	);
	LUT2 #(
		.INIT('h8)
	) name1640 (
		\P1_datao_reg[17]/NET0131 ,
		\si[17]_pad ,
		_w2102_
	);
	LUT2 #(
		.INIT('h8)
	) name1641 (
		\P1_datao_reg[18]/NET0131 ,
		\si[18]_pad ,
		_w2103_
	);
	LUT2 #(
		.INIT('h1)
	) name1642 (
		_w2102_,
		_w2103_,
		_w2104_
	);
	LUT2 #(
		.INIT('h2)
	) name1643 (
		_w2082_,
		_w2104_,
		_w2105_
	);
	LUT2 #(
		.INIT('h1)
	) name1644 (
		_w2101_,
		_w2105_,
		_w2106_
	);
	LUT2 #(
		.INIT('h8)
	) name1645 (
		\P1_datao_reg[8]/NET0131 ,
		\si[8]_pad ,
		_w2107_
	);
	LUT2 #(
		.INIT('h1)
	) name1646 (
		\P1_datao_reg[7]/NET0131 ,
		\si[7]_pad ,
		_w2108_
	);
	LUT2 #(
		.INIT('h1)
	) name1647 (
		\P1_datao_reg[8]/NET0131 ,
		\si[8]_pad ,
		_w2109_
	);
	LUT2 #(
		.INIT('h1)
	) name1648 (
		_w2108_,
		_w2109_,
		_w2110_
	);
	LUT2 #(
		.INIT('h8)
	) name1649 (
		\P1_datao_reg[7]/NET0131 ,
		\si[7]_pad ,
		_w2111_
	);
	LUT2 #(
		.INIT('h1)
	) name1650 (
		\P1_datao_reg[6]/NET0131 ,
		\si[6]_pad ,
		_w2112_
	);
	LUT2 #(
		.INIT('h8)
	) name1651 (
		\P1_datao_reg[5]/NET0131 ,
		\si[5]_pad ,
		_w2113_
	);
	LUT2 #(
		.INIT('h8)
	) name1652 (
		\P1_datao_reg[6]/NET0131 ,
		\si[6]_pad ,
		_w2114_
	);
	LUT2 #(
		.INIT('h1)
	) name1653 (
		_w2113_,
		_w2114_,
		_w2115_
	);
	LUT2 #(
		.INIT('h1)
	) name1654 (
		_w2112_,
		_w2115_,
		_w2116_
	);
	LUT2 #(
		.INIT('h1)
	) name1655 (
		_w2111_,
		_w2116_,
		_w2117_
	);
	LUT2 #(
		.INIT('h2)
	) name1656 (
		_w2110_,
		_w2117_,
		_w2118_
	);
	LUT2 #(
		.INIT('h1)
	) name1657 (
		\P1_datao_reg[4]/NET0131 ,
		\si[4]_pad ,
		_w2119_
	);
	LUT2 #(
		.INIT('h1)
	) name1658 (
		\P1_datao_reg[3]/NET0131 ,
		\si[3]_pad ,
		_w2120_
	);
	LUT2 #(
		.INIT('h8)
	) name1659 (
		\P1_datao_reg[2]/NET0131 ,
		\si[2]_pad ,
		_w2121_
	);
	LUT2 #(
		.INIT('h1)
	) name1660 (
		\P1_datao_reg[2]/NET0131 ,
		\si[2]_pad ,
		_w2122_
	);
	LUT2 #(
		.INIT('h1)
	) name1661 (
		\P1_datao_reg[1]/NET0131 ,
		\si[1]_pad ,
		_w2123_
	);
	LUT2 #(
		.INIT('h8)
	) name1662 (
		\P1_datao_reg[1]/NET0131 ,
		\si[1]_pad ,
		_w2124_
	);
	LUT2 #(
		.INIT('h8)
	) name1663 (
		\P1_datao_reg[0]/NET0131 ,
		\si[0]_pad ,
		_w2125_
	);
	LUT2 #(
		.INIT('h1)
	) name1664 (
		_w2124_,
		_w2125_,
		_w2126_
	);
	LUT2 #(
		.INIT('h1)
	) name1665 (
		_w2123_,
		_w2126_,
		_w2127_
	);
	LUT2 #(
		.INIT('h4)
	) name1666 (
		_w2122_,
		_w2127_,
		_w2128_
	);
	LUT2 #(
		.INIT('h1)
	) name1667 (
		_w2121_,
		_w2128_,
		_w2129_
	);
	LUT2 #(
		.INIT('h1)
	) name1668 (
		_w2120_,
		_w2129_,
		_w2130_
	);
	LUT2 #(
		.INIT('h8)
	) name1669 (
		\P1_datao_reg[4]/NET0131 ,
		\si[4]_pad ,
		_w2131_
	);
	LUT2 #(
		.INIT('h8)
	) name1670 (
		\P1_datao_reg[3]/NET0131 ,
		\si[3]_pad ,
		_w2132_
	);
	LUT2 #(
		.INIT('h1)
	) name1671 (
		_w2131_,
		_w2132_,
		_w2133_
	);
	LUT2 #(
		.INIT('h4)
	) name1672 (
		_w2130_,
		_w2133_,
		_w2134_
	);
	LUT2 #(
		.INIT('h1)
	) name1673 (
		_w2119_,
		_w2134_,
		_w2135_
	);
	LUT2 #(
		.INIT('h1)
	) name1674 (
		\P1_datao_reg[5]/NET0131 ,
		\si[5]_pad ,
		_w2136_
	);
	LUT2 #(
		.INIT('h1)
	) name1675 (
		_w2112_,
		_w2136_,
		_w2137_
	);
	LUT2 #(
		.INIT('h8)
	) name1676 (
		_w2110_,
		_w2137_,
		_w2138_
	);
	LUT2 #(
		.INIT('h8)
	) name1677 (
		_w2135_,
		_w2138_,
		_w2139_
	);
	LUT2 #(
		.INIT('h1)
	) name1678 (
		_w2107_,
		_w2118_,
		_w2140_
	);
	LUT2 #(
		.INIT('h4)
	) name1679 (
		_w2139_,
		_w2140_,
		_w2141_
	);
	LUT2 #(
		.INIT('h1)
	) name1680 (
		\P1_datao_reg[12]/NET0131 ,
		\si[12]_pad ,
		_w2142_
	);
	LUT2 #(
		.INIT('h1)
	) name1681 (
		\P1_datao_reg[11]/NET0131 ,
		\si[11]_pad ,
		_w2143_
	);
	LUT2 #(
		.INIT('h1)
	) name1682 (
		\P1_datao_reg[10]/NET0131 ,
		\si[10]_pad ,
		_w2144_
	);
	LUT2 #(
		.INIT('h1)
	) name1683 (
		_w2143_,
		_w2144_,
		_w2145_
	);
	LUT2 #(
		.INIT('h1)
	) name1684 (
		\P1_datao_reg[9]/NET0131 ,
		\si[9]_pad ,
		_w2146_
	);
	LUT2 #(
		.INIT('h1)
	) name1685 (
		_w2142_,
		_w2146_,
		_w2147_
	);
	LUT2 #(
		.INIT('h8)
	) name1686 (
		_w2145_,
		_w2147_,
		_w2148_
	);
	LUT2 #(
		.INIT('h4)
	) name1687 (
		_w2141_,
		_w2148_,
		_w2149_
	);
	LUT2 #(
		.INIT('h8)
	) name1688 (
		\P1_datao_reg[12]/NET0131 ,
		\si[12]_pad ,
		_w2150_
	);
	LUT2 #(
		.INIT('h8)
	) name1689 (
		\P1_datao_reg[11]/NET0131 ,
		\si[11]_pad ,
		_w2151_
	);
	LUT2 #(
		.INIT('h8)
	) name1690 (
		\P1_datao_reg[10]/NET0131 ,
		\si[10]_pad ,
		_w2152_
	);
	LUT2 #(
		.INIT('h8)
	) name1691 (
		\P1_datao_reg[9]/NET0131 ,
		\si[9]_pad ,
		_w2153_
	);
	LUT2 #(
		.INIT('h1)
	) name1692 (
		_w2152_,
		_w2153_,
		_w2154_
	);
	LUT2 #(
		.INIT('h1)
	) name1693 (
		_w2144_,
		_w2154_,
		_w2155_
	);
	LUT2 #(
		.INIT('h1)
	) name1694 (
		_w2151_,
		_w2155_,
		_w2156_
	);
	LUT2 #(
		.INIT('h1)
	) name1695 (
		_w2142_,
		_w2143_,
		_w2157_
	);
	LUT2 #(
		.INIT('h4)
	) name1696 (
		_w2156_,
		_w2157_,
		_w2158_
	);
	LUT2 #(
		.INIT('h1)
	) name1697 (
		_w2150_,
		_w2158_,
		_w2159_
	);
	LUT2 #(
		.INIT('h4)
	) name1698 (
		_w2149_,
		_w2159_,
		_w2160_
	);
	LUT2 #(
		.INIT('h1)
	) name1699 (
		\P1_datao_reg[13]/NET0131 ,
		\si[13]_pad ,
		_w2161_
	);
	LUT2 #(
		.INIT('h1)
	) name1700 (
		_w2084_,
		_w2161_,
		_w2162_
	);
	LUT2 #(
		.INIT('h8)
	) name1701 (
		_w2090_,
		_w2162_,
		_w2163_
	);
	LUT2 #(
		.INIT('h8)
	) name1702 (
		_w2083_,
		_w2163_,
		_w2164_
	);
	LUT2 #(
		.INIT('h4)
	) name1703 (
		_w2160_,
		_w2164_,
		_w2165_
	);
	LUT2 #(
		.INIT('h4)
	) name1704 (
		_w2097_,
		_w2106_,
		_w2166_
	);
	LUT2 #(
		.INIT('h4)
	) name1705 (
		_w2165_,
		_w2166_,
		_w2167_
	);
	LUT2 #(
		.INIT('h8)
	) name1706 (
		_w2071_,
		_w2076_,
		_w2168_
	);
	LUT2 #(
		.INIT('h4)
	) name1707 (
		_w2167_,
		_w2168_,
		_w2169_
	);
	LUT2 #(
		.INIT('h8)
	) name1708 (
		\P1_datao_reg[27]/NET0131 ,
		\si[27]_pad ,
		_w2170_
	);
	LUT2 #(
		.INIT('h8)
	) name1709 (
		\P1_datao_reg[28]/NET0131 ,
		\si[28]_pad ,
		_w2171_
	);
	LUT2 #(
		.INIT('h1)
	) name1710 (
		_w2170_,
		_w2171_,
		_w2172_
	);
	LUT2 #(
		.INIT('h8)
	) name1711 (
		\P1_datao_reg[26]/NET0131 ,
		\si[26]_pad ,
		_w2173_
	);
	LUT2 #(
		.INIT('h8)
	) name1712 (
		\P1_datao_reg[25]/NET0131 ,
		\si[25]_pad ,
		_w2174_
	);
	LUT2 #(
		.INIT('h1)
	) name1713 (
		_w2173_,
		_w2174_,
		_w2175_
	);
	LUT2 #(
		.INIT('h1)
	) name1714 (
		_w2073_,
		_w2175_,
		_w2176_
	);
	LUT2 #(
		.INIT('h8)
	) name1715 (
		\P1_datao_reg[22]/NET0131 ,
		\si[22]_pad ,
		_w2177_
	);
	LUT2 #(
		.INIT('h8)
	) name1716 (
		\P1_datao_reg[21]/NET0131 ,
		\si[21]_pad ,
		_w2178_
	);
	LUT2 #(
		.INIT('h1)
	) name1717 (
		_w2177_,
		_w2178_,
		_w2179_
	);
	LUT2 #(
		.INIT('h1)
	) name1718 (
		_w2068_,
		_w2179_,
		_w2180_
	);
	LUT2 #(
		.INIT('h8)
	) name1719 (
		_w2067_,
		_w2180_,
		_w2181_
	);
	LUT2 #(
		.INIT('h8)
	) name1720 (
		\P1_datao_reg[23]/NET0131 ,
		\si[23]_pad ,
		_w2182_
	);
	LUT2 #(
		.INIT('h8)
	) name1721 (
		\P1_datao_reg[24]/NET0131 ,
		\si[24]_pad ,
		_w2183_
	);
	LUT2 #(
		.INIT('h1)
	) name1722 (
		_w2182_,
		_w2183_,
		_w2184_
	);
	LUT2 #(
		.INIT('h1)
	) name1723 (
		_w2066_,
		_w2184_,
		_w2185_
	);
	LUT2 #(
		.INIT('h1)
	) name1724 (
		_w2181_,
		_w2185_,
		_w2186_
	);
	LUT2 #(
		.INIT('h2)
	) name1725 (
		_w2075_,
		_w2186_,
		_w2187_
	);
	LUT2 #(
		.INIT('h1)
	) name1726 (
		_w2176_,
		_w2187_,
		_w2188_
	);
	LUT2 #(
		.INIT('h1)
	) name1727 (
		_w2072_,
		_w2188_,
		_w2189_
	);
	LUT2 #(
		.INIT('h2)
	) name1728 (
		_w2172_,
		_w2189_,
		_w2190_
	);
	LUT2 #(
		.INIT('h4)
	) name1729 (
		_w2169_,
		_w2190_,
		_w2191_
	);
	LUT2 #(
		.INIT('h1)
	) name1730 (
		_w2064_,
		_w2191_,
		_w2192_
	);
	LUT2 #(
		.INIT('h1)
	) name1731 (
		_w2063_,
		_w2192_,
		_w2193_
	);
	LUT2 #(
		.INIT('h8)
	) name1732 (
		_w2063_,
		_w2192_,
		_w2194_
	);
	LUT2 #(
		.INIT('h2)
	) name1733 (
		_w543_,
		_w2193_,
		_w2195_
	);
	LUT2 #(
		.INIT('h4)
	) name1734 (
		_w2194_,
		_w2195_,
		_w2196_
	);
	LUT2 #(
		.INIT('h1)
	) name1735 (
		_w2060_,
		_w2196_,
		_w2197_
	);
	LUT2 #(
		.INIT('h1)
	) name1736 (
		_w2059_,
		_w2197_,
		_w2198_
	);
	LUT2 #(
		.INIT('h2)
	) name1737 (
		\P2_IR_reg[31]/NET0131 ,
		_w1995_,
		_w2199_
	);
	LUT2 #(
		.INIT('h1)
	) name1738 (
		\P2_IR_reg[27]/NET0131 ,
		\P2_IR_reg[28]/NET0131 ,
		_w2200_
	);
	LUT2 #(
		.INIT('h4)
	) name1739 (
		\P2_IR_reg[29]/NET0131 ,
		_w2200_,
		_w2201_
	);
	LUT2 #(
		.INIT('h8)
	) name1740 (
		_w2045_,
		_w2201_,
		_w2202_
	);
	LUT2 #(
		.INIT('h2)
	) name1741 (
		\P2_IR_reg[31]/NET0131 ,
		_w2202_,
		_w2203_
	);
	LUT2 #(
		.INIT('h1)
	) name1742 (
		_w2199_,
		_w2203_,
		_w2204_
	);
	LUT2 #(
		.INIT('h2)
	) name1743 (
		\P2_IR_reg[30]/NET0131 ,
		_w2204_,
		_w2205_
	);
	LUT2 #(
		.INIT('h4)
	) name1744 (
		\P2_IR_reg[30]/NET0131 ,
		_w2204_,
		_w2206_
	);
	LUT2 #(
		.INIT('h1)
	) name1745 (
		_w2205_,
		_w2206_,
		_w2207_
	);
	LUT2 #(
		.INIT('h2)
	) name1746 (
		\P2_IR_reg[31]/NET0131 ,
		_w2016_,
		_w2208_
	);
	LUT2 #(
		.INIT('h4)
	) name1747 (
		\P2_IR_reg[21]/NET0131 ,
		_w2200_,
		_w2209_
	);
	LUT2 #(
		.INIT('h8)
	) name1748 (
		_w2045_,
		_w2209_,
		_w2210_
	);
	LUT2 #(
		.INIT('h2)
	) name1749 (
		\P2_IR_reg[31]/NET0131 ,
		_w2210_,
		_w2211_
	);
	LUT2 #(
		.INIT('h1)
	) name1750 (
		_w2208_,
		_w2211_,
		_w2212_
	);
	LUT2 #(
		.INIT('h2)
	) name1751 (
		\P2_IR_reg[29]/NET0131 ,
		_w2212_,
		_w2213_
	);
	LUT2 #(
		.INIT('h4)
	) name1752 (
		\P2_IR_reg[29]/NET0131 ,
		_w2212_,
		_w2214_
	);
	LUT2 #(
		.INIT('h1)
	) name1753 (
		_w2213_,
		_w2214_,
		_w2215_
	);
	LUT2 #(
		.INIT('h8)
	) name1754 (
		_w2207_,
		_w2215_,
		_w2216_
	);
	LUT2 #(
		.INIT('h8)
	) name1755 (
		\P2_reg3_reg[3]/NET0131 ,
		\P2_reg3_reg[4]/NET0131 ,
		_w2217_
	);
	LUT2 #(
		.INIT('h8)
	) name1756 (
		\P2_reg3_reg[5]/NET0131 ,
		_w2217_,
		_w2218_
	);
	LUT2 #(
		.INIT('h8)
	) name1757 (
		\P2_reg3_reg[6]/NET0131 ,
		_w2218_,
		_w2219_
	);
	LUT2 #(
		.INIT('h8)
	) name1758 (
		\P2_reg3_reg[7]/NET0131 ,
		_w2219_,
		_w2220_
	);
	LUT2 #(
		.INIT('h8)
	) name1759 (
		\P2_reg3_reg[8]/NET0131 ,
		_w2220_,
		_w2221_
	);
	LUT2 #(
		.INIT('h8)
	) name1760 (
		\P2_reg3_reg[9]/NET0131 ,
		_w2221_,
		_w2222_
	);
	LUT2 #(
		.INIT('h8)
	) name1761 (
		\P2_reg3_reg[10]/NET0131 ,
		_w2222_,
		_w2223_
	);
	LUT2 #(
		.INIT('h8)
	) name1762 (
		\P2_reg3_reg[11]/NET0131 ,
		\P2_reg3_reg[12]/NET0131 ,
		_w2224_
	);
	LUT2 #(
		.INIT('h8)
	) name1763 (
		\P2_reg3_reg[13]/NET0131 ,
		\P2_reg3_reg[14]/NET0131 ,
		_w2225_
	);
	LUT2 #(
		.INIT('h8)
	) name1764 (
		_w2224_,
		_w2225_,
		_w2226_
	);
	LUT2 #(
		.INIT('h8)
	) name1765 (
		_w2223_,
		_w2226_,
		_w2227_
	);
	LUT2 #(
		.INIT('h8)
	) name1766 (
		\P2_reg3_reg[15]/NET0131 ,
		\P2_reg3_reg[16]/NET0131 ,
		_w2228_
	);
	LUT2 #(
		.INIT('h8)
	) name1767 (
		_w2227_,
		_w2228_,
		_w2229_
	);
	LUT2 #(
		.INIT('h8)
	) name1768 (
		\P2_reg3_reg[20]/NET0131 ,
		\P2_reg3_reg[21]/NET0131 ,
		_w2230_
	);
	LUT2 #(
		.INIT('h8)
	) name1769 (
		\P2_reg3_reg[22]/NET0131 ,
		_w2230_,
		_w2231_
	);
	LUT2 #(
		.INIT('h8)
	) name1770 (
		\P2_reg3_reg[17]/NET0131 ,
		\P2_reg3_reg[18]/NET0131 ,
		_w2232_
	);
	LUT2 #(
		.INIT('h8)
	) name1771 (
		\P2_reg3_reg[19]/NET0131 ,
		\P2_reg3_reg[23]/NET0131 ,
		_w2233_
	);
	LUT2 #(
		.INIT('h8)
	) name1772 (
		\P2_reg3_reg[24]/NET0131 ,
		_w2233_,
		_w2234_
	);
	LUT2 #(
		.INIT('h8)
	) name1773 (
		_w2232_,
		_w2234_,
		_w2235_
	);
	LUT2 #(
		.INIT('h8)
	) name1774 (
		_w2231_,
		_w2235_,
		_w2236_
	);
	LUT2 #(
		.INIT('h8)
	) name1775 (
		_w2229_,
		_w2236_,
		_w2237_
	);
	LUT2 #(
		.INIT('h8)
	) name1776 (
		\P2_reg3_reg[25]/NET0131 ,
		\P2_reg3_reg[26]/NET0131 ,
		_w2238_
	);
	LUT2 #(
		.INIT('h8)
	) name1777 (
		\P2_reg3_reg[27]/NET0131 ,
		\P2_reg3_reg[28]/NET0131 ,
		_w2239_
	);
	LUT2 #(
		.INIT('h8)
	) name1778 (
		_w2238_,
		_w2239_,
		_w2240_
	);
	LUT2 #(
		.INIT('h8)
	) name1779 (
		_w2237_,
		_w2240_,
		_w2241_
	);
	LUT2 #(
		.INIT('h8)
	) name1780 (
		_w2216_,
		_w2241_,
		_w2242_
	);
	LUT2 #(
		.INIT('h2)
	) name1781 (
		_w2207_,
		_w2215_,
		_w2243_
	);
	LUT2 #(
		.INIT('h8)
	) name1782 (
		\P2_reg2_reg[29]/NET0131 ,
		_w2243_,
		_w2244_
	);
	LUT2 #(
		.INIT('h1)
	) name1783 (
		_w2207_,
		_w2215_,
		_w2245_
	);
	LUT2 #(
		.INIT('h8)
	) name1784 (
		\P2_reg0_reg[29]/NET0131 ,
		_w2245_,
		_w2246_
	);
	LUT2 #(
		.INIT('h4)
	) name1785 (
		_w2207_,
		_w2215_,
		_w2247_
	);
	LUT2 #(
		.INIT('h8)
	) name1786 (
		\P2_reg1_reg[29]/NET0131 ,
		_w2247_,
		_w2248_
	);
	LUT2 #(
		.INIT('h1)
	) name1787 (
		_w2242_,
		_w2244_,
		_w2249_
	);
	LUT2 #(
		.INIT('h1)
	) name1788 (
		_w2246_,
		_w2248_,
		_w2250_
	);
	LUT2 #(
		.INIT('h8)
	) name1789 (
		_w2249_,
		_w2250_,
		_w2251_
	);
	LUT2 #(
		.INIT('h8)
	) name1790 (
		_w2198_,
		_w2251_,
		_w2252_
	);
	LUT2 #(
		.INIT('h1)
	) name1791 (
		_w2198_,
		_w2251_,
		_w2253_
	);
	LUT2 #(
		.INIT('h1)
	) name1792 (
		_w2252_,
		_w2253_,
		_w2254_
	);
	LUT2 #(
		.INIT('h2)
	) name1793 (
		\P2_IR_reg[31]/NET0131 ,
		_w1976_,
		_w2255_
	);
	LUT2 #(
		.INIT('h1)
	) name1794 (
		\P2_IR_reg[19]/NET0131 ,
		_w2255_,
		_w2256_
	);
	LUT2 #(
		.INIT('h8)
	) name1795 (
		\P2_IR_reg[19]/NET0131 ,
		_w2255_,
		_w2257_
	);
	LUT2 #(
		.INIT('h1)
	) name1796 (
		_w2256_,
		_w2257_,
		_w2258_
	);
	LUT2 #(
		.INIT('h2)
	) name1797 (
		_w2059_,
		_w2258_,
		_w2259_
	);
	LUT2 #(
		.INIT('h2)
	) name1798 (
		\P1_datao_reg[19]/NET0131 ,
		_w543_,
		_w2260_
	);
	LUT2 #(
		.INIT('h1)
	) name1799 (
		_w2077_,
		_w2084_,
		_w2261_
	);
	LUT2 #(
		.INIT('h4)
	) name1800 (
		_w2079_,
		_w2261_,
		_w2262_
	);
	LUT2 #(
		.INIT('h4)
	) name1801 (
		_w2089_,
		_w2262_,
		_w2263_
	);
	LUT2 #(
		.INIT('h1)
	) name1802 (
		_w2119_,
		_w2136_,
		_w2264_
	);
	LUT2 #(
		.INIT('h4)
	) name1803 (
		_w2112_,
		_w2264_,
		_w2265_
	);
	LUT2 #(
		.INIT('h4)
	) name1804 (
		_w2134_,
		_w2265_,
		_w2266_
	);
	LUT2 #(
		.INIT('h1)
	) name1805 (
		_w2116_,
		_w2266_,
		_w2267_
	);
	LUT2 #(
		.INIT('h1)
	) name1806 (
		_w2109_,
		_w2146_,
		_w2268_
	);
	LUT2 #(
		.INIT('h4)
	) name1807 (
		_w2108_,
		_w2268_,
		_w2269_
	);
	LUT2 #(
		.INIT('h4)
	) name1808 (
		_w2144_,
		_w2269_,
		_w2270_
	);
	LUT2 #(
		.INIT('h4)
	) name1809 (
		_w2267_,
		_w2270_,
		_w2271_
	);
	LUT2 #(
		.INIT('h1)
	) name1810 (
		_w2107_,
		_w2111_,
		_w2272_
	);
	LUT2 #(
		.INIT('h4)
	) name1811 (
		_w2144_,
		_w2268_,
		_w2273_
	);
	LUT2 #(
		.INIT('h4)
	) name1812 (
		_w2272_,
		_w2273_,
		_w2274_
	);
	LUT2 #(
		.INIT('h1)
	) name1813 (
		_w2155_,
		_w2274_,
		_w2275_
	);
	LUT2 #(
		.INIT('h4)
	) name1814 (
		_w2271_,
		_w2275_,
		_w2276_
	);
	LUT2 #(
		.INIT('h2)
	) name1815 (
		_w2157_,
		_w2161_,
		_w2277_
	);
	LUT2 #(
		.INIT('h4)
	) name1816 (
		_w2088_,
		_w2277_,
		_w2278_
	);
	LUT2 #(
		.INIT('h4)
	) name1817 (
		_w2276_,
		_w2278_,
		_w2279_
	);
	LUT2 #(
		.INIT('h8)
	) name1818 (
		_w2263_,
		_w2279_,
		_w2280_
	);
	LUT2 #(
		.INIT('h1)
	) name1819 (
		_w2142_,
		_w2161_,
		_w2281_
	);
	LUT2 #(
		.INIT('h1)
	) name1820 (
		_w2150_,
		_w2151_,
		_w2282_
	);
	LUT2 #(
		.INIT('h2)
	) name1821 (
		_w2281_,
		_w2282_,
		_w2283_
	);
	LUT2 #(
		.INIT('h2)
	) name1822 (
		_w2093_,
		_w2283_,
		_w2284_
	);
	LUT2 #(
		.INIT('h1)
	) name1823 (
		_w2088_,
		_w2284_,
		_w2285_
	);
	LUT2 #(
		.INIT('h8)
	) name1824 (
		_w2263_,
		_w2285_,
		_w2286_
	);
	LUT2 #(
		.INIT('h4)
	) name1825 (
		_w2087_,
		_w2261_,
		_w2287_
	);
	LUT2 #(
		.INIT('h2)
	) name1826 (
		_w2104_,
		_w2287_,
		_w2288_
	);
	LUT2 #(
		.INIT('h1)
	) name1827 (
		_w2079_,
		_w2288_,
		_w2289_
	);
	LUT2 #(
		.INIT('h1)
	) name1828 (
		_w2286_,
		_w2289_,
		_w2290_
	);
	LUT2 #(
		.INIT('h4)
	) name1829 (
		_w2280_,
		_w2290_,
		_w2291_
	);
	LUT2 #(
		.INIT('h1)
	) name1830 (
		_w2080_,
		_w2098_,
		_w2292_
	);
	LUT2 #(
		.INIT('h2)
	) name1831 (
		_w2291_,
		_w2292_,
		_w2293_
	);
	LUT2 #(
		.INIT('h4)
	) name1832 (
		_w2291_,
		_w2292_,
		_w2294_
	);
	LUT2 #(
		.INIT('h2)
	) name1833 (
		_w543_,
		_w2293_,
		_w2295_
	);
	LUT2 #(
		.INIT('h4)
	) name1834 (
		_w2294_,
		_w2295_,
		_w2296_
	);
	LUT2 #(
		.INIT('h1)
	) name1835 (
		_w2260_,
		_w2296_,
		_w2297_
	);
	LUT2 #(
		.INIT('h4)
	) name1836 (
		_w2059_,
		_w2297_,
		_w2298_
	);
	LUT2 #(
		.INIT('h1)
	) name1837 (
		_w2259_,
		_w2298_,
		_w2299_
	);
	LUT2 #(
		.INIT('h8)
	) name1838 (
		\P2_reg0_reg[19]/NET0131 ,
		_w2245_,
		_w2300_
	);
	LUT2 #(
		.INIT('h8)
	) name1839 (
		\P2_reg2_reg[19]/NET0131 ,
		_w2243_,
		_w2301_
	);
	LUT2 #(
		.INIT('h8)
	) name1840 (
		\P2_reg1_reg[19]/NET0131 ,
		_w2247_,
		_w2302_
	);
	LUT2 #(
		.INIT('h8)
	) name1841 (
		\P2_reg3_reg[17]/NET0131 ,
		_w2229_,
		_w2303_
	);
	LUT2 #(
		.INIT('h8)
	) name1842 (
		\P2_reg3_reg[18]/NET0131 ,
		_w2303_,
		_w2304_
	);
	LUT2 #(
		.INIT('h1)
	) name1843 (
		\P2_reg3_reg[19]/NET0131 ,
		_w2304_,
		_w2305_
	);
	LUT2 #(
		.INIT('h8)
	) name1844 (
		\P2_reg3_reg[19]/NET0131 ,
		_w2304_,
		_w2306_
	);
	LUT2 #(
		.INIT('h1)
	) name1845 (
		_w2305_,
		_w2306_,
		_w2307_
	);
	LUT2 #(
		.INIT('h8)
	) name1846 (
		_w2216_,
		_w2307_,
		_w2308_
	);
	LUT2 #(
		.INIT('h1)
	) name1847 (
		_w2300_,
		_w2301_,
		_w2309_
	);
	LUT2 #(
		.INIT('h4)
	) name1848 (
		_w2302_,
		_w2309_,
		_w2310_
	);
	LUT2 #(
		.INIT('h4)
	) name1849 (
		_w2308_,
		_w2310_,
		_w2311_
	);
	LUT2 #(
		.INIT('h4)
	) name1850 (
		_w2299_,
		_w2311_,
		_w2312_
	);
	LUT2 #(
		.INIT('h2)
	) name1851 (
		\P1_datao_reg[20]/NET0131 ,
		_w543_,
		_w2313_
	);
	LUT2 #(
		.INIT('h1)
	) name1852 (
		_w2098_,
		_w2103_,
		_w2314_
	);
	LUT2 #(
		.INIT('h1)
	) name1853 (
		_w2080_,
		_w2314_,
		_w2315_
	);
	LUT2 #(
		.INIT('h1)
	) name1854 (
		_w2086_,
		_w2102_,
		_w2316_
	);
	LUT2 #(
		.INIT('h1)
	) name1855 (
		_w2077_,
		_w2316_,
		_w2317_
	);
	LUT2 #(
		.INIT('h8)
	) name1856 (
		_w2081_,
		_w2317_,
		_w2318_
	);
	LUT2 #(
		.INIT('h8)
	) name1857 (
		_w2090_,
		_w2281_,
		_w2319_
	);
	LUT2 #(
		.INIT('h1)
	) name1858 (
		_w2121_,
		_w2132_,
		_w2320_
	);
	LUT2 #(
		.INIT('h4)
	) name1859 (
		_w2128_,
		_w2320_,
		_w2321_
	);
	LUT2 #(
		.INIT('h1)
	) name1860 (
		_w2120_,
		_w2321_,
		_w2322_
	);
	LUT2 #(
		.INIT('h8)
	) name1861 (
		_w2265_,
		_w2322_,
		_w2323_
	);
	LUT2 #(
		.INIT('h1)
	) name1862 (
		_w2111_,
		_w2114_,
		_w2324_
	);
	LUT2 #(
		.INIT('h1)
	) name1863 (
		_w2113_,
		_w2131_,
		_w2325_
	);
	LUT2 #(
		.INIT('h1)
	) name1864 (
		_w2136_,
		_w2325_,
		_w2326_
	);
	LUT2 #(
		.INIT('h4)
	) name1865 (
		_w2112_,
		_w2326_,
		_w2327_
	);
	LUT2 #(
		.INIT('h2)
	) name1866 (
		_w2324_,
		_w2327_,
		_w2328_
	);
	LUT2 #(
		.INIT('h4)
	) name1867 (
		_w2323_,
		_w2328_,
		_w2329_
	);
	LUT2 #(
		.INIT('h1)
	) name1868 (
		_w2108_,
		_w2329_,
		_w2330_
	);
	LUT2 #(
		.INIT('h8)
	) name1869 (
		_w2145_,
		_w2268_,
		_w2331_
	);
	LUT2 #(
		.INIT('h8)
	) name1870 (
		_w2330_,
		_w2331_,
		_w2332_
	);
	LUT2 #(
		.INIT('h8)
	) name1871 (
		_w2319_,
		_w2332_,
		_w2333_
	);
	LUT2 #(
		.INIT('h1)
	) name1872 (
		_w2091_,
		_w2150_,
		_w2334_
	);
	LUT2 #(
		.INIT('h1)
	) name1873 (
		_w2161_,
		_w2334_,
		_w2335_
	);
	LUT2 #(
		.INIT('h8)
	) name1874 (
		_w2090_,
		_w2335_,
		_w2336_
	);
	LUT2 #(
		.INIT('h1)
	) name1875 (
		_w2107_,
		_w2153_,
		_w2337_
	);
	LUT2 #(
		.INIT('h1)
	) name1876 (
		_w2146_,
		_w2337_,
		_w2338_
	);
	LUT2 #(
		.INIT('h1)
	) name1877 (
		_w2152_,
		_w2338_,
		_w2339_
	);
	LUT2 #(
		.INIT('h2)
	) name1878 (
		_w2145_,
		_w2339_,
		_w2340_
	);
	LUT2 #(
		.INIT('h1)
	) name1879 (
		_w2151_,
		_w2340_,
		_w2341_
	);
	LUT2 #(
		.INIT('h2)
	) name1880 (
		_w2319_,
		_w2341_,
		_w2342_
	);
	LUT2 #(
		.INIT('h1)
	) name1881 (
		_w2085_,
		_w2092_,
		_w2343_
	);
	LUT2 #(
		.INIT('h1)
	) name1882 (
		_w2089_,
		_w2343_,
		_w2344_
	);
	LUT2 #(
		.INIT('h1)
	) name1883 (
		_w2336_,
		_w2344_,
		_w2345_
	);
	LUT2 #(
		.INIT('h4)
	) name1884 (
		_w2342_,
		_w2345_,
		_w2346_
	);
	LUT2 #(
		.INIT('h4)
	) name1885 (
		_w2333_,
		_w2346_,
		_w2347_
	);
	LUT2 #(
		.INIT('h4)
	) name1886 (
		_w2080_,
		_w2262_,
		_w2348_
	);
	LUT2 #(
		.INIT('h4)
	) name1887 (
		_w2347_,
		_w2348_,
		_w2349_
	);
	LUT2 #(
		.INIT('h1)
	) name1888 (
		_w2315_,
		_w2318_,
		_w2350_
	);
	LUT2 #(
		.INIT('h4)
	) name1889 (
		_w2349_,
		_w2350_,
		_w2351_
	);
	LUT2 #(
		.INIT('h1)
	) name1890 (
		_w2078_,
		_w2099_,
		_w2352_
	);
	LUT2 #(
		.INIT('h2)
	) name1891 (
		_w2351_,
		_w2352_,
		_w2353_
	);
	LUT2 #(
		.INIT('h4)
	) name1892 (
		_w2351_,
		_w2352_,
		_w2354_
	);
	LUT2 #(
		.INIT('h2)
	) name1893 (
		_w543_,
		_w2353_,
		_w2355_
	);
	LUT2 #(
		.INIT('h4)
	) name1894 (
		_w2354_,
		_w2355_,
		_w2356_
	);
	LUT2 #(
		.INIT('h1)
	) name1895 (
		_w2313_,
		_w2356_,
		_w2357_
	);
	LUT2 #(
		.INIT('h1)
	) name1896 (
		_w2059_,
		_w2357_,
		_w2358_
	);
	LUT2 #(
		.INIT('h8)
	) name1897 (
		\P2_reg1_reg[20]/NET0131 ,
		_w2247_,
		_w2359_
	);
	LUT2 #(
		.INIT('h8)
	) name1898 (
		\P2_reg0_reg[20]/NET0131 ,
		_w2245_,
		_w2360_
	);
	LUT2 #(
		.INIT('h8)
	) name1899 (
		\P2_reg2_reg[20]/NET0131 ,
		_w2243_,
		_w2361_
	);
	LUT2 #(
		.INIT('h8)
	) name1900 (
		\P2_reg3_reg[20]/NET0131 ,
		_w2306_,
		_w2362_
	);
	LUT2 #(
		.INIT('h1)
	) name1901 (
		\P2_reg3_reg[20]/NET0131 ,
		_w2306_,
		_w2363_
	);
	LUT2 #(
		.INIT('h1)
	) name1902 (
		_w2362_,
		_w2363_,
		_w2364_
	);
	LUT2 #(
		.INIT('h8)
	) name1903 (
		_w2216_,
		_w2364_,
		_w2365_
	);
	LUT2 #(
		.INIT('h1)
	) name1904 (
		_w2359_,
		_w2360_,
		_w2366_
	);
	LUT2 #(
		.INIT('h4)
	) name1905 (
		_w2361_,
		_w2366_,
		_w2367_
	);
	LUT2 #(
		.INIT('h4)
	) name1906 (
		_w2365_,
		_w2367_,
		_w2368_
	);
	LUT2 #(
		.INIT('h4)
	) name1907 (
		_w2358_,
		_w2368_,
		_w2369_
	);
	LUT2 #(
		.INIT('h1)
	) name1908 (
		_w2312_,
		_w2369_,
		_w2370_
	);
	LUT2 #(
		.INIT('h8)
	) name1909 (
		\P2_reg1_reg[17]/NET0131 ,
		_w2247_,
		_w2371_
	);
	LUT2 #(
		.INIT('h1)
	) name1910 (
		\P2_reg3_reg[17]/NET0131 ,
		_w2229_,
		_w2372_
	);
	LUT2 #(
		.INIT('h1)
	) name1911 (
		_w2303_,
		_w2372_,
		_w2373_
	);
	LUT2 #(
		.INIT('h8)
	) name1912 (
		_w2216_,
		_w2373_,
		_w2374_
	);
	LUT2 #(
		.INIT('h8)
	) name1913 (
		\P2_reg2_reg[17]/NET0131 ,
		_w2243_,
		_w2375_
	);
	LUT2 #(
		.INIT('h8)
	) name1914 (
		\P2_reg0_reg[17]/NET0131 ,
		_w2245_,
		_w2376_
	);
	LUT2 #(
		.INIT('h1)
	) name1915 (
		_w2371_,
		_w2374_,
		_w2377_
	);
	LUT2 #(
		.INIT('h1)
	) name1916 (
		_w2375_,
		_w2376_,
		_w2378_
	);
	LUT2 #(
		.INIT('h8)
	) name1917 (
		_w2377_,
		_w2378_,
		_w2379_
	);
	LUT2 #(
		.INIT('h2)
	) name1918 (
		\P2_IR_reg[31]/NET0131 ,
		_w2013_,
		_w2380_
	);
	LUT2 #(
		.INIT('h2)
	) name1919 (
		\P2_IR_reg[31]/NET0131 ,
		_w1989_,
		_w2381_
	);
	LUT2 #(
		.INIT('h1)
	) name1920 (
		_w2380_,
		_w2381_,
		_w2382_
	);
	LUT2 #(
		.INIT('h2)
	) name1921 (
		\P2_IR_reg[17]/NET0131 ,
		_w2382_,
		_w2383_
	);
	LUT2 #(
		.INIT('h4)
	) name1922 (
		\P2_IR_reg[17]/NET0131 ,
		_w2382_,
		_w2384_
	);
	LUT2 #(
		.INIT('h1)
	) name1923 (
		_w2383_,
		_w2384_,
		_w2385_
	);
	LUT2 #(
		.INIT('h2)
	) name1924 (
		_w2059_,
		_w2385_,
		_w2386_
	);
	LUT2 #(
		.INIT('h2)
	) name1925 (
		\P1_datao_reg[17]/NET0131 ,
		_w543_,
		_w2387_
	);
	LUT2 #(
		.INIT('h8)
	) name1926 (
		_w2149_,
		_w2163_,
		_w2388_
	);
	LUT2 #(
		.INIT('h4)
	) name1927 (
		_w2159_,
		_w2163_,
		_w2389_
	);
	LUT2 #(
		.INIT('h1)
	) name1928 (
		_w2096_,
		_w2389_,
		_w2390_
	);
	LUT2 #(
		.INIT('h4)
	) name1929 (
		_w2388_,
		_w2390_,
		_w2391_
	);
	LUT2 #(
		.INIT('h1)
	) name1930 (
		_w2077_,
		_w2102_,
		_w2392_
	);
	LUT2 #(
		.INIT('h2)
	) name1931 (
		_w2391_,
		_w2392_,
		_w2393_
	);
	LUT2 #(
		.INIT('h4)
	) name1932 (
		_w2391_,
		_w2392_,
		_w2394_
	);
	LUT2 #(
		.INIT('h2)
	) name1933 (
		_w543_,
		_w2393_,
		_w2395_
	);
	LUT2 #(
		.INIT('h4)
	) name1934 (
		_w2394_,
		_w2395_,
		_w2396_
	);
	LUT2 #(
		.INIT('h1)
	) name1935 (
		_w2387_,
		_w2396_,
		_w2397_
	);
	LUT2 #(
		.INIT('h4)
	) name1936 (
		_w2059_,
		_w2397_,
		_w2398_
	);
	LUT2 #(
		.INIT('h1)
	) name1937 (
		_w2386_,
		_w2398_,
		_w2399_
	);
	LUT2 #(
		.INIT('h2)
	) name1938 (
		_w2379_,
		_w2399_,
		_w2400_
	);
	LUT2 #(
		.INIT('h2)
	) name1939 (
		\P2_IR_reg[31]/NET0131 ,
		_w1992_,
		_w2401_
	);
	LUT2 #(
		.INIT('h1)
	) name1940 (
		\P2_IR_reg[18]/NET0131 ,
		_w2401_,
		_w2402_
	);
	LUT2 #(
		.INIT('h8)
	) name1941 (
		\P2_IR_reg[18]/NET0131 ,
		_w2401_,
		_w2403_
	);
	LUT2 #(
		.INIT('h1)
	) name1942 (
		_w2402_,
		_w2403_,
		_w2404_
	);
	LUT2 #(
		.INIT('h2)
	) name1943 (
		_w2059_,
		_w2404_,
		_w2405_
	);
	LUT2 #(
		.INIT('h2)
	) name1944 (
		\P1_datao_reg[18]/NET0131 ,
		_w543_,
		_w2406_
	);
	LUT2 #(
		.INIT('h1)
	) name1945 (
		_w2079_,
		_w2103_,
		_w2407_
	);
	LUT2 #(
		.INIT('h8)
	) name1946 (
		_w2264_,
		_w2322_,
		_w2408_
	);
	LUT2 #(
		.INIT('h1)
	) name1947 (
		_w2326_,
		_w2408_,
		_w2409_
	);
	LUT2 #(
		.INIT('h4)
	) name1948 (
		_w2112_,
		_w2269_,
		_w2410_
	);
	LUT2 #(
		.INIT('h4)
	) name1949 (
		_w2409_,
		_w2410_,
		_w2411_
	);
	LUT2 #(
		.INIT('h2)
	) name1950 (
		_w2269_,
		_w2324_,
		_w2412_
	);
	LUT2 #(
		.INIT('h1)
	) name1951 (
		_w2338_,
		_w2412_,
		_w2413_
	);
	LUT2 #(
		.INIT('h4)
	) name1952 (
		_w2411_,
		_w2413_,
		_w2414_
	);
	LUT2 #(
		.INIT('h4)
	) name1953 (
		_w2144_,
		_w2277_,
		_w2415_
	);
	LUT2 #(
		.INIT('h4)
	) name1954 (
		_w2414_,
		_w2415_,
		_w2416_
	);
	LUT2 #(
		.INIT('h8)
	) name1955 (
		_w2090_,
		_w2261_,
		_w2417_
	);
	LUT2 #(
		.INIT('h8)
	) name1956 (
		_w2416_,
		_w2417_,
		_w2418_
	);
	LUT2 #(
		.INIT('h8)
	) name1957 (
		_w2261_,
		_w2344_,
		_w2419_
	);
	LUT2 #(
		.INIT('h1)
	) name1958 (
		_w2317_,
		_w2419_,
		_w2420_
	);
	LUT2 #(
		.INIT('h1)
	) name1959 (
		_w2151_,
		_w2152_,
		_w2421_
	);
	LUT2 #(
		.INIT('h2)
	) name1960 (
		_w2277_,
		_w2421_,
		_w2422_
	);
	LUT2 #(
		.INIT('h1)
	) name1961 (
		_w2335_,
		_w2422_,
		_w2423_
	);
	LUT2 #(
		.INIT('h2)
	) name1962 (
		_w2417_,
		_w2423_,
		_w2424_
	);
	LUT2 #(
		.INIT('h2)
	) name1963 (
		_w2420_,
		_w2424_,
		_w2425_
	);
	LUT2 #(
		.INIT('h4)
	) name1964 (
		_w2418_,
		_w2425_,
		_w2426_
	);
	LUT2 #(
		.INIT('h2)
	) name1965 (
		_w2407_,
		_w2426_,
		_w2427_
	);
	LUT2 #(
		.INIT('h4)
	) name1966 (
		_w2407_,
		_w2426_,
		_w2428_
	);
	LUT2 #(
		.INIT('h2)
	) name1967 (
		_w543_,
		_w2427_,
		_w2429_
	);
	LUT2 #(
		.INIT('h4)
	) name1968 (
		_w2428_,
		_w2429_,
		_w2430_
	);
	LUT2 #(
		.INIT('h1)
	) name1969 (
		_w2406_,
		_w2430_,
		_w2431_
	);
	LUT2 #(
		.INIT('h4)
	) name1970 (
		_w2059_,
		_w2431_,
		_w2432_
	);
	LUT2 #(
		.INIT('h1)
	) name1971 (
		_w2405_,
		_w2432_,
		_w2433_
	);
	LUT2 #(
		.INIT('h8)
	) name1972 (
		\P2_reg2_reg[18]/NET0131 ,
		_w2243_,
		_w2434_
	);
	LUT2 #(
		.INIT('h8)
	) name1973 (
		\P2_reg0_reg[18]/NET0131 ,
		_w2245_,
		_w2435_
	);
	LUT2 #(
		.INIT('h8)
	) name1974 (
		\P2_reg1_reg[18]/NET0131 ,
		_w2247_,
		_w2436_
	);
	LUT2 #(
		.INIT('h1)
	) name1975 (
		\P2_reg3_reg[18]/NET0131 ,
		_w2303_,
		_w2437_
	);
	LUT2 #(
		.INIT('h1)
	) name1976 (
		_w2304_,
		_w2437_,
		_w2438_
	);
	LUT2 #(
		.INIT('h8)
	) name1977 (
		_w2216_,
		_w2438_,
		_w2439_
	);
	LUT2 #(
		.INIT('h1)
	) name1978 (
		_w2434_,
		_w2435_,
		_w2440_
	);
	LUT2 #(
		.INIT('h4)
	) name1979 (
		_w2436_,
		_w2440_,
		_w2441_
	);
	LUT2 #(
		.INIT('h4)
	) name1980 (
		_w2439_,
		_w2441_,
		_w2442_
	);
	LUT2 #(
		.INIT('h4)
	) name1981 (
		_w2433_,
		_w2442_,
		_w2443_
	);
	LUT2 #(
		.INIT('h1)
	) name1982 (
		_w2400_,
		_w2443_,
		_w2444_
	);
	LUT2 #(
		.INIT('h8)
	) name1983 (
		_w2370_,
		_w2444_,
		_w2445_
	);
	LUT2 #(
		.INIT('h1)
	) name1984 (
		\P2_reg3_reg[8]/NET0131 ,
		_w2220_,
		_w2446_
	);
	LUT2 #(
		.INIT('h1)
	) name1985 (
		_w2221_,
		_w2446_,
		_w2447_
	);
	LUT2 #(
		.INIT('h8)
	) name1986 (
		_w2216_,
		_w2447_,
		_w2448_
	);
	LUT2 #(
		.INIT('h8)
	) name1987 (
		\P2_reg1_reg[8]/NET0131 ,
		_w2247_,
		_w2449_
	);
	LUT2 #(
		.INIT('h8)
	) name1988 (
		\P2_reg0_reg[8]/NET0131 ,
		_w2245_,
		_w2450_
	);
	LUT2 #(
		.INIT('h8)
	) name1989 (
		\P2_reg2_reg[8]/NET0131 ,
		_w2243_,
		_w2451_
	);
	LUT2 #(
		.INIT('h1)
	) name1990 (
		_w2448_,
		_w2449_,
		_w2452_
	);
	LUT2 #(
		.INIT('h1)
	) name1991 (
		_w2450_,
		_w2451_,
		_w2453_
	);
	LUT2 #(
		.INIT('h8)
	) name1992 (
		_w2452_,
		_w2453_,
		_w2454_
	);
	LUT2 #(
		.INIT('h2)
	) name1993 (
		\P2_IR_reg[31]/NET0131 ,
		_w1964_,
		_w2455_
	);
	LUT2 #(
		.INIT('h2)
	) name1994 (
		\P2_IR_reg[31]/NET0131 ,
		_w1966_,
		_w2456_
	);
	LUT2 #(
		.INIT('h1)
	) name1995 (
		_w2455_,
		_w2456_,
		_w2457_
	);
	LUT2 #(
		.INIT('h2)
	) name1996 (
		\P2_IR_reg[8]/NET0131 ,
		_w2457_,
		_w2458_
	);
	LUT2 #(
		.INIT('h4)
	) name1997 (
		\P2_IR_reg[8]/NET0131 ,
		_w2457_,
		_w2459_
	);
	LUT2 #(
		.INIT('h1)
	) name1998 (
		_w2458_,
		_w2459_,
		_w2460_
	);
	LUT2 #(
		.INIT('h2)
	) name1999 (
		_w2059_,
		_w2460_,
		_w2461_
	);
	LUT2 #(
		.INIT('h2)
	) name2000 (
		\P1_datao_reg[8]/NET0131 ,
		_w543_,
		_w2462_
	);
	LUT2 #(
		.INIT('h1)
	) name2001 (
		_w2107_,
		_w2109_,
		_w2463_
	);
	LUT2 #(
		.INIT('h1)
	) name2002 (
		_w2330_,
		_w2463_,
		_w2464_
	);
	LUT2 #(
		.INIT('h8)
	) name2003 (
		_w2330_,
		_w2463_,
		_w2465_
	);
	LUT2 #(
		.INIT('h2)
	) name2004 (
		_w543_,
		_w2464_,
		_w2466_
	);
	LUT2 #(
		.INIT('h4)
	) name2005 (
		_w2465_,
		_w2466_,
		_w2467_
	);
	LUT2 #(
		.INIT('h1)
	) name2006 (
		_w2462_,
		_w2467_,
		_w2468_
	);
	LUT2 #(
		.INIT('h4)
	) name2007 (
		_w2059_,
		_w2468_,
		_w2469_
	);
	LUT2 #(
		.INIT('h1)
	) name2008 (
		_w2461_,
		_w2469_,
		_w2470_
	);
	LUT2 #(
		.INIT('h2)
	) name2009 (
		_w2454_,
		_w2470_,
		_w2471_
	);
	LUT2 #(
		.INIT('h8)
	) name2010 (
		\P2_reg2_reg[7]/NET0131 ,
		_w2243_,
		_w2472_
	);
	LUT2 #(
		.INIT('h8)
	) name2011 (
		\P2_reg1_reg[7]/NET0131 ,
		_w2247_,
		_w2473_
	);
	LUT2 #(
		.INIT('h8)
	) name2012 (
		\P2_reg0_reg[7]/NET0131 ,
		_w2245_,
		_w2474_
	);
	LUT2 #(
		.INIT('h1)
	) name2013 (
		\P2_reg3_reg[7]/NET0131 ,
		_w2219_,
		_w2475_
	);
	LUT2 #(
		.INIT('h1)
	) name2014 (
		_w2220_,
		_w2475_,
		_w2476_
	);
	LUT2 #(
		.INIT('h8)
	) name2015 (
		_w2216_,
		_w2476_,
		_w2477_
	);
	LUT2 #(
		.INIT('h1)
	) name2016 (
		_w2472_,
		_w2473_,
		_w2478_
	);
	LUT2 #(
		.INIT('h1)
	) name2017 (
		_w2474_,
		_w2477_,
		_w2479_
	);
	LUT2 #(
		.INIT('h8)
	) name2018 (
		_w2478_,
		_w2479_,
		_w2480_
	);
	LUT2 #(
		.INIT('h2)
	) name2019 (
		\P2_IR_reg[31]/NET0131 ,
		_w1965_,
		_w2481_
	);
	LUT2 #(
		.INIT('h1)
	) name2020 (
		_w2455_,
		_w2481_,
		_w2482_
	);
	LUT2 #(
		.INIT('h2)
	) name2021 (
		\P2_IR_reg[7]/NET0131 ,
		_w2482_,
		_w2483_
	);
	LUT2 #(
		.INIT('h4)
	) name2022 (
		\P2_IR_reg[7]/NET0131 ,
		_w2482_,
		_w2484_
	);
	LUT2 #(
		.INIT('h1)
	) name2023 (
		_w2483_,
		_w2484_,
		_w2485_
	);
	LUT2 #(
		.INIT('h2)
	) name2024 (
		_w2059_,
		_w2485_,
		_w2486_
	);
	LUT2 #(
		.INIT('h2)
	) name2025 (
		\P1_datao_reg[7]/NET0131 ,
		_w543_,
		_w2487_
	);
	LUT2 #(
		.INIT('h1)
	) name2026 (
		_w2108_,
		_w2111_,
		_w2488_
	);
	LUT2 #(
		.INIT('h4)
	) name2027 (
		_w2267_,
		_w2488_,
		_w2489_
	);
	LUT2 #(
		.INIT('h2)
	) name2028 (
		_w2267_,
		_w2488_,
		_w2490_
	);
	LUT2 #(
		.INIT('h2)
	) name2029 (
		_w543_,
		_w2489_,
		_w2491_
	);
	LUT2 #(
		.INIT('h4)
	) name2030 (
		_w2490_,
		_w2491_,
		_w2492_
	);
	LUT2 #(
		.INIT('h1)
	) name2031 (
		_w2487_,
		_w2492_,
		_w2493_
	);
	LUT2 #(
		.INIT('h4)
	) name2032 (
		_w2059_,
		_w2493_,
		_w2494_
	);
	LUT2 #(
		.INIT('h1)
	) name2033 (
		_w2486_,
		_w2494_,
		_w2495_
	);
	LUT2 #(
		.INIT('h2)
	) name2034 (
		_w2480_,
		_w2495_,
		_w2496_
	);
	LUT2 #(
		.INIT('h1)
	) name2035 (
		_w2471_,
		_w2496_,
		_w2497_
	);
	LUT2 #(
		.INIT('h1)
	) name2036 (
		\P2_reg3_reg[6]/NET0131 ,
		_w2218_,
		_w2498_
	);
	LUT2 #(
		.INIT('h1)
	) name2037 (
		_w2219_,
		_w2498_,
		_w2499_
	);
	LUT2 #(
		.INIT('h8)
	) name2038 (
		_w2216_,
		_w2499_,
		_w2500_
	);
	LUT2 #(
		.INIT('h8)
	) name2039 (
		\P2_reg0_reg[6]/NET0131 ,
		_w2245_,
		_w2501_
	);
	LUT2 #(
		.INIT('h8)
	) name2040 (
		\P2_reg1_reg[6]/NET0131 ,
		_w2247_,
		_w2502_
	);
	LUT2 #(
		.INIT('h8)
	) name2041 (
		\P2_reg2_reg[6]/NET0131 ,
		_w2243_,
		_w2503_
	);
	LUT2 #(
		.INIT('h1)
	) name2042 (
		_w2500_,
		_w2501_,
		_w2504_
	);
	LUT2 #(
		.INIT('h1)
	) name2043 (
		_w2502_,
		_w2503_,
		_w2505_
	);
	LUT2 #(
		.INIT('h8)
	) name2044 (
		_w2504_,
		_w2505_,
		_w2506_
	);
	LUT2 #(
		.INIT('h2)
	) name2045 (
		\P1_datao_reg[6]/NET0131 ,
		_w543_,
		_w2507_
	);
	LUT2 #(
		.INIT('h1)
	) name2046 (
		_w2112_,
		_w2114_,
		_w2508_
	);
	LUT2 #(
		.INIT('h4)
	) name2047 (
		_w2409_,
		_w2508_,
		_w2509_
	);
	LUT2 #(
		.INIT('h2)
	) name2048 (
		_w2409_,
		_w2508_,
		_w2510_
	);
	LUT2 #(
		.INIT('h2)
	) name2049 (
		_w543_,
		_w2509_,
		_w2511_
	);
	LUT2 #(
		.INIT('h4)
	) name2050 (
		_w2510_,
		_w2511_,
		_w2512_
	);
	LUT2 #(
		.INIT('h1)
	) name2051 (
		_w2507_,
		_w2512_,
		_w2513_
	);
	LUT2 #(
		.INIT('h1)
	) name2052 (
		_w2059_,
		_w2513_,
		_w2514_
	);
	LUT2 #(
		.INIT('h8)
	) name2053 (
		\P2_IR_reg[31]/NET0131 ,
		\P2_IR_reg[5]/NET0131 ,
		_w2515_
	);
	LUT2 #(
		.INIT('h1)
	) name2054 (
		_w2455_,
		_w2515_,
		_w2516_
	);
	LUT2 #(
		.INIT('h2)
	) name2055 (
		\P2_IR_reg[6]/NET0131 ,
		_w2516_,
		_w2517_
	);
	LUT2 #(
		.INIT('h4)
	) name2056 (
		\P2_IR_reg[6]/NET0131 ,
		_w2516_,
		_w2518_
	);
	LUT2 #(
		.INIT('h1)
	) name2057 (
		_w2517_,
		_w2518_,
		_w2519_
	);
	LUT2 #(
		.INIT('h8)
	) name2058 (
		_w2059_,
		_w2519_,
		_w2520_
	);
	LUT2 #(
		.INIT('h1)
	) name2059 (
		_w2514_,
		_w2520_,
		_w2521_
	);
	LUT2 #(
		.INIT('h8)
	) name2060 (
		_w2506_,
		_w2521_,
		_w2522_
	);
	LUT2 #(
		.INIT('h8)
	) name2061 (
		\P2_reg0_reg[5]/NET0131 ,
		_w2245_,
		_w2523_
	);
	LUT2 #(
		.INIT('h8)
	) name2062 (
		\P2_reg2_reg[5]/NET0131 ,
		_w2243_,
		_w2524_
	);
	LUT2 #(
		.INIT('h1)
	) name2063 (
		\P2_reg3_reg[5]/NET0131 ,
		_w2217_,
		_w2525_
	);
	LUT2 #(
		.INIT('h1)
	) name2064 (
		_w2218_,
		_w2525_,
		_w2526_
	);
	LUT2 #(
		.INIT('h8)
	) name2065 (
		_w2216_,
		_w2526_,
		_w2527_
	);
	LUT2 #(
		.INIT('h8)
	) name2066 (
		\P2_reg1_reg[5]/NET0131 ,
		_w2247_,
		_w2528_
	);
	LUT2 #(
		.INIT('h1)
	) name2067 (
		_w2523_,
		_w2524_,
		_w2529_
	);
	LUT2 #(
		.INIT('h1)
	) name2068 (
		_w2527_,
		_w2528_,
		_w2530_
	);
	LUT2 #(
		.INIT('h8)
	) name2069 (
		_w2529_,
		_w2530_,
		_w2531_
	);
	LUT2 #(
		.INIT('h2)
	) name2070 (
		\P1_datao_reg[5]/NET0131 ,
		_w543_,
		_w2532_
	);
	LUT2 #(
		.INIT('h1)
	) name2071 (
		_w2113_,
		_w2136_,
		_w2533_
	);
	LUT2 #(
		.INIT('h1)
	) name2072 (
		_w2135_,
		_w2533_,
		_w2534_
	);
	LUT2 #(
		.INIT('h8)
	) name2073 (
		_w2135_,
		_w2533_,
		_w2535_
	);
	LUT2 #(
		.INIT('h2)
	) name2074 (
		_w543_,
		_w2534_,
		_w2536_
	);
	LUT2 #(
		.INIT('h4)
	) name2075 (
		_w2535_,
		_w2536_,
		_w2537_
	);
	LUT2 #(
		.INIT('h1)
	) name2076 (
		_w2532_,
		_w2537_,
		_w2538_
	);
	LUT2 #(
		.INIT('h1)
	) name2077 (
		_w2059_,
		_w2538_,
		_w2539_
	);
	LUT2 #(
		.INIT('h2)
	) name2078 (
		\P2_IR_reg[5]/NET0131 ,
		_w2455_,
		_w2540_
	);
	LUT2 #(
		.INIT('h4)
	) name2079 (
		\P2_IR_reg[5]/NET0131 ,
		_w2455_,
		_w2541_
	);
	LUT2 #(
		.INIT('h1)
	) name2080 (
		_w2540_,
		_w2541_,
		_w2542_
	);
	LUT2 #(
		.INIT('h2)
	) name2081 (
		_w2059_,
		_w2542_,
		_w2543_
	);
	LUT2 #(
		.INIT('h1)
	) name2082 (
		_w2539_,
		_w2543_,
		_w2544_
	);
	LUT2 #(
		.INIT('h8)
	) name2083 (
		_w2531_,
		_w2544_,
		_w2545_
	);
	LUT2 #(
		.INIT('h8)
	) name2084 (
		\P2_reg0_reg[2]/NET0131 ,
		_w2245_,
		_w2546_
	);
	LUT2 #(
		.INIT('h8)
	) name2085 (
		\P2_reg1_reg[2]/NET0131 ,
		_w2247_,
		_w2547_
	);
	LUT2 #(
		.INIT('h8)
	) name2086 (
		\P2_reg2_reg[2]/NET0131 ,
		_w2243_,
		_w2548_
	);
	LUT2 #(
		.INIT('h8)
	) name2087 (
		\P2_reg3_reg[2]/NET0131 ,
		_w2216_,
		_w2549_
	);
	LUT2 #(
		.INIT('h1)
	) name2088 (
		_w2546_,
		_w2547_,
		_w2550_
	);
	LUT2 #(
		.INIT('h1)
	) name2089 (
		_w2548_,
		_w2549_,
		_w2551_
	);
	LUT2 #(
		.INIT('h8)
	) name2090 (
		_w2550_,
		_w2551_,
		_w2552_
	);
	LUT2 #(
		.INIT('h2)
	) name2091 (
		\P1_datao_reg[2]/NET0131 ,
		_w543_,
		_w2553_
	);
	LUT2 #(
		.INIT('h1)
	) name2092 (
		_w2121_,
		_w2122_,
		_w2554_
	);
	LUT2 #(
		.INIT('h1)
	) name2093 (
		_w2127_,
		_w2554_,
		_w2555_
	);
	LUT2 #(
		.INIT('h8)
	) name2094 (
		_w2127_,
		_w2554_,
		_w2556_
	);
	LUT2 #(
		.INIT('h2)
	) name2095 (
		_w543_,
		_w2555_,
		_w2557_
	);
	LUT2 #(
		.INIT('h4)
	) name2096 (
		_w2556_,
		_w2557_,
		_w2558_
	);
	LUT2 #(
		.INIT('h1)
	) name2097 (
		_w2553_,
		_w2558_,
		_w2559_
	);
	LUT2 #(
		.INIT('h1)
	) name2098 (
		_w2059_,
		_w2559_,
		_w2560_
	);
	LUT2 #(
		.INIT('h2)
	) name2099 (
		\P2_IR_reg[31]/NET0131 ,
		_w1961_,
		_w2561_
	);
	LUT2 #(
		.INIT('h8)
	) name2100 (
		\P2_IR_reg[2]/NET0131 ,
		_w2561_,
		_w2562_
	);
	LUT2 #(
		.INIT('h1)
	) name2101 (
		\P2_IR_reg[2]/NET0131 ,
		_w2561_,
		_w2563_
	);
	LUT2 #(
		.INIT('h1)
	) name2102 (
		_w2562_,
		_w2563_,
		_w2564_
	);
	LUT2 #(
		.INIT('h8)
	) name2103 (
		_w2059_,
		_w2564_,
		_w2565_
	);
	LUT2 #(
		.INIT('h1)
	) name2104 (
		_w2560_,
		_w2565_,
		_w2566_
	);
	LUT2 #(
		.INIT('h1)
	) name2105 (
		_w2552_,
		_w2566_,
		_w2567_
	);
	LUT2 #(
		.INIT('h8)
	) name2106 (
		\P2_reg3_reg[1]/NET0131 ,
		_w2216_,
		_w2568_
	);
	LUT2 #(
		.INIT('h8)
	) name2107 (
		\P2_reg0_reg[1]/NET0131 ,
		_w2245_,
		_w2569_
	);
	LUT2 #(
		.INIT('h8)
	) name2108 (
		\P2_reg2_reg[1]/NET0131 ,
		_w2243_,
		_w2570_
	);
	LUT2 #(
		.INIT('h8)
	) name2109 (
		\P2_reg1_reg[1]/NET0131 ,
		_w2247_,
		_w2571_
	);
	LUT2 #(
		.INIT('h1)
	) name2110 (
		_w2568_,
		_w2569_,
		_w2572_
	);
	LUT2 #(
		.INIT('h1)
	) name2111 (
		_w2570_,
		_w2571_,
		_w2573_
	);
	LUT2 #(
		.INIT('h8)
	) name2112 (
		_w2572_,
		_w2573_,
		_w2574_
	);
	LUT2 #(
		.INIT('h8)
	) name2113 (
		\P2_IR_reg[0]/NET0131 ,
		\P2_IR_reg[31]/NET0131 ,
		_w2575_
	);
	LUT2 #(
		.INIT('h1)
	) name2114 (
		\P2_IR_reg[1]/NET0131 ,
		_w2575_,
		_w2576_
	);
	LUT2 #(
		.INIT('h8)
	) name2115 (
		\P2_IR_reg[1]/NET0131 ,
		_w2575_,
		_w2577_
	);
	LUT2 #(
		.INIT('h1)
	) name2116 (
		_w2576_,
		_w2577_,
		_w2578_
	);
	LUT2 #(
		.INIT('h8)
	) name2117 (
		_w2059_,
		_w2578_,
		_w2579_
	);
	LUT2 #(
		.INIT('h1)
	) name2118 (
		\P1_datao_reg[1]/NET0131 ,
		_w543_,
		_w2580_
	);
	LUT2 #(
		.INIT('h1)
	) name2119 (
		_w2123_,
		_w2124_,
		_w2581_
	);
	LUT2 #(
		.INIT('h4)
	) name2120 (
		_w2125_,
		_w2581_,
		_w2582_
	);
	LUT2 #(
		.INIT('h2)
	) name2121 (
		_w2125_,
		_w2581_,
		_w2583_
	);
	LUT2 #(
		.INIT('h2)
	) name2122 (
		_w543_,
		_w2582_,
		_w2584_
	);
	LUT2 #(
		.INIT('h4)
	) name2123 (
		_w2583_,
		_w2584_,
		_w2585_
	);
	LUT2 #(
		.INIT('h1)
	) name2124 (
		_w2580_,
		_w2585_,
		_w2586_
	);
	LUT2 #(
		.INIT('h4)
	) name2125 (
		_w2059_,
		_w2586_,
		_w2587_
	);
	LUT2 #(
		.INIT('h1)
	) name2126 (
		_w2579_,
		_w2587_,
		_w2588_
	);
	LUT2 #(
		.INIT('h8)
	) name2127 (
		_w2574_,
		_w2588_,
		_w2589_
	);
	LUT2 #(
		.INIT('h1)
	) name2128 (
		_w2574_,
		_w2588_,
		_w2590_
	);
	LUT2 #(
		.INIT('h8)
	) name2129 (
		\P2_reg2_reg[0]/NET0131 ,
		_w2243_,
		_w2591_
	);
	LUT2 #(
		.INIT('h8)
	) name2130 (
		\P2_reg0_reg[0]/NET0131 ,
		_w2245_,
		_w2592_
	);
	LUT2 #(
		.INIT('h8)
	) name2131 (
		\P2_reg1_reg[0]/NET0131 ,
		_w2247_,
		_w2593_
	);
	LUT2 #(
		.INIT('h8)
	) name2132 (
		\P2_reg3_reg[0]/NET0131 ,
		_w2216_,
		_w2594_
	);
	LUT2 #(
		.INIT('h1)
	) name2133 (
		_w2591_,
		_w2592_,
		_w2595_
	);
	LUT2 #(
		.INIT('h1)
	) name2134 (
		_w2593_,
		_w2594_,
		_w2596_
	);
	LUT2 #(
		.INIT('h8)
	) name2135 (
		_w2595_,
		_w2596_,
		_w2597_
	);
	LUT2 #(
		.INIT('h8)
	) name2136 (
		\si[0]_pad ,
		_w543_,
		_w2598_
	);
	LUT2 #(
		.INIT('h1)
	) name2137 (
		\P1_datao_reg[0]/NET0131 ,
		_w2598_,
		_w2599_
	);
	LUT2 #(
		.INIT('h8)
	) name2138 (
		\P1_datao_reg[0]/NET0131 ,
		_w2598_,
		_w2600_
	);
	LUT2 #(
		.INIT('h1)
	) name2139 (
		_w2599_,
		_w2600_,
		_w2601_
	);
	LUT2 #(
		.INIT('h4)
	) name2140 (
		_w2059_,
		_w2601_,
		_w2602_
	);
	LUT2 #(
		.INIT('h8)
	) name2141 (
		\P2_IR_reg[0]/NET0131 ,
		_w2059_,
		_w2603_
	);
	LUT2 #(
		.INIT('h1)
	) name2142 (
		_w2602_,
		_w2603_,
		_w2604_
	);
	LUT2 #(
		.INIT('h1)
	) name2143 (
		_w2597_,
		_w2604_,
		_w2605_
	);
	LUT2 #(
		.INIT('h1)
	) name2144 (
		_w2590_,
		_w2605_,
		_w2606_
	);
	LUT2 #(
		.INIT('h1)
	) name2145 (
		_w2589_,
		_w2606_,
		_w2607_
	);
	LUT2 #(
		.INIT('h1)
	) name2146 (
		_w2567_,
		_w2607_,
		_w2608_
	);
	LUT2 #(
		.INIT('h8)
	) name2147 (
		_w2552_,
		_w2566_,
		_w2609_
	);
	LUT2 #(
		.INIT('h8)
	) name2148 (
		\P2_reg1_reg[3]/NET0131 ,
		_w2247_,
		_w2610_
	);
	LUT2 #(
		.INIT('h8)
	) name2149 (
		\P2_reg2_reg[3]/NET0131 ,
		_w2243_,
		_w2611_
	);
	LUT2 #(
		.INIT('h8)
	) name2150 (
		\P2_reg0_reg[3]/NET0131 ,
		_w2245_,
		_w2612_
	);
	LUT2 #(
		.INIT('h4)
	) name2151 (
		\P2_reg3_reg[3]/NET0131 ,
		_w2216_,
		_w2613_
	);
	LUT2 #(
		.INIT('h1)
	) name2152 (
		_w2610_,
		_w2611_,
		_w2614_
	);
	LUT2 #(
		.INIT('h1)
	) name2153 (
		_w2612_,
		_w2613_,
		_w2615_
	);
	LUT2 #(
		.INIT('h8)
	) name2154 (
		_w2614_,
		_w2615_,
		_w2616_
	);
	LUT2 #(
		.INIT('h2)
	) name2155 (
		\P1_datao_reg[3]/NET0131 ,
		_w543_,
		_w2617_
	);
	LUT2 #(
		.INIT('h1)
	) name2156 (
		_w2120_,
		_w2132_,
		_w2618_
	);
	LUT2 #(
		.INIT('h2)
	) name2157 (
		_w2129_,
		_w2618_,
		_w2619_
	);
	LUT2 #(
		.INIT('h4)
	) name2158 (
		_w2129_,
		_w2618_,
		_w2620_
	);
	LUT2 #(
		.INIT('h2)
	) name2159 (
		_w543_,
		_w2619_,
		_w2621_
	);
	LUT2 #(
		.INIT('h4)
	) name2160 (
		_w2620_,
		_w2621_,
		_w2622_
	);
	LUT2 #(
		.INIT('h1)
	) name2161 (
		_w2617_,
		_w2622_,
		_w2623_
	);
	LUT2 #(
		.INIT('h1)
	) name2162 (
		_w2059_,
		_w2623_,
		_w2624_
	);
	LUT2 #(
		.INIT('h2)
	) name2163 (
		\P2_IR_reg[31]/NET0131 ,
		_w1962_,
		_w2625_
	);
	LUT2 #(
		.INIT('h1)
	) name2164 (
		\P2_IR_reg[3]/NET0131 ,
		_w2625_,
		_w2626_
	);
	LUT2 #(
		.INIT('h8)
	) name2165 (
		\P2_IR_reg[31]/NET0131 ,
		\P2_IR_reg[3]/NET0131 ,
		_w2627_
	);
	LUT2 #(
		.INIT('h4)
	) name2166 (
		_w1962_,
		_w2627_,
		_w2628_
	);
	LUT2 #(
		.INIT('h1)
	) name2167 (
		_w2626_,
		_w2628_,
		_w2629_
	);
	LUT2 #(
		.INIT('h8)
	) name2168 (
		_w2059_,
		_w2629_,
		_w2630_
	);
	LUT2 #(
		.INIT('h1)
	) name2169 (
		_w2624_,
		_w2630_,
		_w2631_
	);
	LUT2 #(
		.INIT('h8)
	) name2170 (
		_w2616_,
		_w2631_,
		_w2632_
	);
	LUT2 #(
		.INIT('h1)
	) name2171 (
		_w2609_,
		_w2632_,
		_w2633_
	);
	LUT2 #(
		.INIT('h1)
	) name2172 (
		\P2_reg3_reg[3]/NET0131 ,
		\P2_reg3_reg[4]/NET0131 ,
		_w2634_
	);
	LUT2 #(
		.INIT('h1)
	) name2173 (
		_w2217_,
		_w2634_,
		_w2635_
	);
	LUT2 #(
		.INIT('h8)
	) name2174 (
		_w2216_,
		_w2635_,
		_w2636_
	);
	LUT2 #(
		.INIT('h8)
	) name2175 (
		\P2_reg2_reg[4]/NET0131 ,
		_w2243_,
		_w2637_
	);
	LUT2 #(
		.INIT('h8)
	) name2176 (
		\P2_reg1_reg[4]/NET0131 ,
		_w2247_,
		_w2638_
	);
	LUT2 #(
		.INIT('h8)
	) name2177 (
		\P2_reg0_reg[4]/NET0131 ,
		_w2245_,
		_w2639_
	);
	LUT2 #(
		.INIT('h1)
	) name2178 (
		_w2636_,
		_w2637_,
		_w2640_
	);
	LUT2 #(
		.INIT('h1)
	) name2179 (
		_w2638_,
		_w2639_,
		_w2641_
	);
	LUT2 #(
		.INIT('h8)
	) name2180 (
		_w2640_,
		_w2641_,
		_w2642_
	);
	LUT2 #(
		.INIT('h1)
	) name2181 (
		_w2625_,
		_w2627_,
		_w2643_
	);
	LUT2 #(
		.INIT('h2)
	) name2182 (
		\P2_IR_reg[4]/NET0131 ,
		_w2643_,
		_w2644_
	);
	LUT2 #(
		.INIT('h4)
	) name2183 (
		\P2_IR_reg[4]/NET0131 ,
		_w2643_,
		_w2645_
	);
	LUT2 #(
		.INIT('h1)
	) name2184 (
		_w2644_,
		_w2645_,
		_w2646_
	);
	LUT2 #(
		.INIT('h8)
	) name2185 (
		_w2059_,
		_w2646_,
		_w2647_
	);
	LUT2 #(
		.INIT('h1)
	) name2186 (
		\P1_datao_reg[4]/NET0131 ,
		_w543_,
		_w2648_
	);
	LUT2 #(
		.INIT('h1)
	) name2187 (
		_w2119_,
		_w2131_,
		_w2649_
	);
	LUT2 #(
		.INIT('h4)
	) name2188 (
		_w2322_,
		_w2649_,
		_w2650_
	);
	LUT2 #(
		.INIT('h2)
	) name2189 (
		_w2322_,
		_w2649_,
		_w2651_
	);
	LUT2 #(
		.INIT('h2)
	) name2190 (
		_w543_,
		_w2650_,
		_w2652_
	);
	LUT2 #(
		.INIT('h4)
	) name2191 (
		_w2651_,
		_w2652_,
		_w2653_
	);
	LUT2 #(
		.INIT('h1)
	) name2192 (
		_w2648_,
		_w2653_,
		_w2654_
	);
	LUT2 #(
		.INIT('h4)
	) name2193 (
		_w2059_,
		_w2654_,
		_w2655_
	);
	LUT2 #(
		.INIT('h1)
	) name2194 (
		_w2647_,
		_w2655_,
		_w2656_
	);
	LUT2 #(
		.INIT('h8)
	) name2195 (
		_w2642_,
		_w2656_,
		_w2657_
	);
	LUT2 #(
		.INIT('h2)
	) name2196 (
		_w2633_,
		_w2657_,
		_w2658_
	);
	LUT2 #(
		.INIT('h4)
	) name2197 (
		_w2608_,
		_w2658_,
		_w2659_
	);
	LUT2 #(
		.INIT('h1)
	) name2198 (
		_w2642_,
		_w2656_,
		_w2660_
	);
	LUT2 #(
		.INIT('h1)
	) name2199 (
		_w2616_,
		_w2631_,
		_w2661_
	);
	LUT2 #(
		.INIT('h1)
	) name2200 (
		_w2660_,
		_w2661_,
		_w2662_
	);
	LUT2 #(
		.INIT('h1)
	) name2201 (
		_w2657_,
		_w2662_,
		_w2663_
	);
	LUT2 #(
		.INIT('h1)
	) name2202 (
		_w2659_,
		_w2663_,
		_w2664_
	);
	LUT2 #(
		.INIT('h1)
	) name2203 (
		_w2522_,
		_w2545_,
		_w2665_
	);
	LUT2 #(
		.INIT('h4)
	) name2204 (
		_w2664_,
		_w2665_,
		_w2666_
	);
	LUT2 #(
		.INIT('h8)
	) name2205 (
		_w2497_,
		_w2666_,
		_w2667_
	);
	LUT2 #(
		.INIT('h1)
	) name2206 (
		_w2506_,
		_w2521_,
		_w2668_
	);
	LUT2 #(
		.INIT('h1)
	) name2207 (
		_w2531_,
		_w2544_,
		_w2669_
	);
	LUT2 #(
		.INIT('h4)
	) name2208 (
		_w2522_,
		_w2669_,
		_w2670_
	);
	LUT2 #(
		.INIT('h1)
	) name2209 (
		_w2668_,
		_w2670_,
		_w2671_
	);
	LUT2 #(
		.INIT('h2)
	) name2210 (
		_w2497_,
		_w2671_,
		_w2672_
	);
	LUT2 #(
		.INIT('h4)
	) name2211 (
		_w2454_,
		_w2470_,
		_w2673_
	);
	LUT2 #(
		.INIT('h4)
	) name2212 (
		_w2480_,
		_w2495_,
		_w2674_
	);
	LUT2 #(
		.INIT('h1)
	) name2213 (
		_w2673_,
		_w2674_,
		_w2675_
	);
	LUT2 #(
		.INIT('h1)
	) name2214 (
		_w2471_,
		_w2675_,
		_w2676_
	);
	LUT2 #(
		.INIT('h1)
	) name2215 (
		_w2672_,
		_w2676_,
		_w2677_
	);
	LUT2 #(
		.INIT('h4)
	) name2216 (
		_w2667_,
		_w2677_,
		_w2678_
	);
	LUT2 #(
		.INIT('h8)
	) name2217 (
		\P2_reg3_reg[11]/NET0131 ,
		_w2223_,
		_w2679_
	);
	LUT2 #(
		.INIT('h1)
	) name2218 (
		\P2_reg3_reg[11]/NET0131 ,
		_w2223_,
		_w2680_
	);
	LUT2 #(
		.INIT('h1)
	) name2219 (
		_w2679_,
		_w2680_,
		_w2681_
	);
	LUT2 #(
		.INIT('h8)
	) name2220 (
		_w2216_,
		_w2681_,
		_w2682_
	);
	LUT2 #(
		.INIT('h8)
	) name2221 (
		\P2_reg0_reg[11]/NET0131 ,
		_w2245_,
		_w2683_
	);
	LUT2 #(
		.INIT('h8)
	) name2222 (
		\P2_reg1_reg[11]/NET0131 ,
		_w2247_,
		_w2684_
	);
	LUT2 #(
		.INIT('h8)
	) name2223 (
		\P2_reg2_reg[11]/NET0131 ,
		_w2243_,
		_w2685_
	);
	LUT2 #(
		.INIT('h1)
	) name2224 (
		_w2682_,
		_w2683_,
		_w2686_
	);
	LUT2 #(
		.INIT('h1)
	) name2225 (
		_w2684_,
		_w2685_,
		_w2687_
	);
	LUT2 #(
		.INIT('h8)
	) name2226 (
		_w2686_,
		_w2687_,
		_w2688_
	);
	LUT2 #(
		.INIT('h2)
	) name2227 (
		\P2_IR_reg[31]/NET0131 ,
		_w1969_,
		_w2689_
	);
	LUT2 #(
		.INIT('h8)
	) name2228 (
		\P2_IR_reg[10]/NET0131 ,
		\P2_IR_reg[31]/NET0131 ,
		_w2690_
	);
	LUT2 #(
		.INIT('h1)
	) name2229 (
		_w2689_,
		_w2690_,
		_w2691_
	);
	LUT2 #(
		.INIT('h2)
	) name2230 (
		\P2_IR_reg[11]/NET0131 ,
		_w2691_,
		_w2692_
	);
	LUT2 #(
		.INIT('h4)
	) name2231 (
		\P2_IR_reg[11]/NET0131 ,
		_w2691_,
		_w2693_
	);
	LUT2 #(
		.INIT('h1)
	) name2232 (
		_w2692_,
		_w2693_,
		_w2694_
	);
	LUT2 #(
		.INIT('h2)
	) name2233 (
		_w2059_,
		_w2694_,
		_w2695_
	);
	LUT2 #(
		.INIT('h2)
	) name2234 (
		\P1_datao_reg[11]/NET0131 ,
		_w543_,
		_w2696_
	);
	LUT2 #(
		.INIT('h1)
	) name2235 (
		_w2143_,
		_w2151_,
		_w2697_
	);
	LUT2 #(
		.INIT('h4)
	) name2236 (
		_w2276_,
		_w2697_,
		_w2698_
	);
	LUT2 #(
		.INIT('h2)
	) name2237 (
		_w2276_,
		_w2697_,
		_w2699_
	);
	LUT2 #(
		.INIT('h2)
	) name2238 (
		_w543_,
		_w2698_,
		_w2700_
	);
	LUT2 #(
		.INIT('h4)
	) name2239 (
		_w2699_,
		_w2700_,
		_w2701_
	);
	LUT2 #(
		.INIT('h1)
	) name2240 (
		_w2696_,
		_w2701_,
		_w2702_
	);
	LUT2 #(
		.INIT('h4)
	) name2241 (
		_w2059_,
		_w2702_,
		_w2703_
	);
	LUT2 #(
		.INIT('h1)
	) name2242 (
		_w2695_,
		_w2703_,
		_w2704_
	);
	LUT2 #(
		.INIT('h2)
	) name2243 (
		_w2688_,
		_w2704_,
		_w2705_
	);
	LUT2 #(
		.INIT('h8)
	) name2244 (
		\P2_reg1_reg[12]/NET0131 ,
		_w2247_,
		_w2706_
	);
	LUT2 #(
		.INIT('h8)
	) name2245 (
		\P2_reg3_reg[12]/NET0131 ,
		_w2679_,
		_w2707_
	);
	LUT2 #(
		.INIT('h1)
	) name2246 (
		\P2_reg3_reg[12]/NET0131 ,
		_w2679_,
		_w2708_
	);
	LUT2 #(
		.INIT('h1)
	) name2247 (
		_w2707_,
		_w2708_,
		_w2709_
	);
	LUT2 #(
		.INIT('h8)
	) name2248 (
		_w2216_,
		_w2709_,
		_w2710_
	);
	LUT2 #(
		.INIT('h8)
	) name2249 (
		\P2_reg2_reg[12]/NET0131 ,
		_w2243_,
		_w2711_
	);
	LUT2 #(
		.INIT('h8)
	) name2250 (
		\P2_reg0_reg[12]/NET0131 ,
		_w2245_,
		_w2712_
	);
	LUT2 #(
		.INIT('h1)
	) name2251 (
		_w2706_,
		_w2710_,
		_w2713_
	);
	LUT2 #(
		.INIT('h1)
	) name2252 (
		_w2711_,
		_w2712_,
		_w2714_
	);
	LUT2 #(
		.INIT('h8)
	) name2253 (
		_w2713_,
		_w2714_,
		_w2715_
	);
	LUT2 #(
		.INIT('h2)
	) name2254 (
		\P2_IR_reg[31]/NET0131 ,
		_w1959_,
		_w2716_
	);
	LUT2 #(
		.INIT('h1)
	) name2255 (
		_w2689_,
		_w2716_,
		_w2717_
	);
	LUT2 #(
		.INIT('h2)
	) name2256 (
		\P2_IR_reg[12]/NET0131 ,
		_w2717_,
		_w2718_
	);
	LUT2 #(
		.INIT('h4)
	) name2257 (
		\P2_IR_reg[12]/NET0131 ,
		_w2717_,
		_w2719_
	);
	LUT2 #(
		.INIT('h1)
	) name2258 (
		_w2718_,
		_w2719_,
		_w2720_
	);
	LUT2 #(
		.INIT('h2)
	) name2259 (
		_w2059_,
		_w2720_,
		_w2721_
	);
	LUT2 #(
		.INIT('h2)
	) name2260 (
		\P1_datao_reg[12]/NET0131 ,
		_w543_,
		_w2722_
	);
	LUT2 #(
		.INIT('h1)
	) name2261 (
		_w2142_,
		_w2150_,
		_w2723_
	);
	LUT2 #(
		.INIT('h4)
	) name2262 (
		_w2332_,
		_w2341_,
		_w2724_
	);
	LUT2 #(
		.INIT('h2)
	) name2263 (
		_w2723_,
		_w2724_,
		_w2725_
	);
	LUT2 #(
		.INIT('h4)
	) name2264 (
		_w2723_,
		_w2724_,
		_w2726_
	);
	LUT2 #(
		.INIT('h2)
	) name2265 (
		_w543_,
		_w2725_,
		_w2727_
	);
	LUT2 #(
		.INIT('h4)
	) name2266 (
		_w2726_,
		_w2727_,
		_w2728_
	);
	LUT2 #(
		.INIT('h1)
	) name2267 (
		_w2722_,
		_w2728_,
		_w2729_
	);
	LUT2 #(
		.INIT('h4)
	) name2268 (
		_w2059_,
		_w2729_,
		_w2730_
	);
	LUT2 #(
		.INIT('h1)
	) name2269 (
		_w2721_,
		_w2730_,
		_w2731_
	);
	LUT2 #(
		.INIT('h2)
	) name2270 (
		_w2715_,
		_w2731_,
		_w2732_
	);
	LUT2 #(
		.INIT('h1)
	) name2271 (
		_w2705_,
		_w2732_,
		_w2733_
	);
	LUT2 #(
		.INIT('h1)
	) name2272 (
		\P2_reg3_reg[10]/NET0131 ,
		_w2222_,
		_w2734_
	);
	LUT2 #(
		.INIT('h1)
	) name2273 (
		_w2223_,
		_w2734_,
		_w2735_
	);
	LUT2 #(
		.INIT('h8)
	) name2274 (
		_w2216_,
		_w2735_,
		_w2736_
	);
	LUT2 #(
		.INIT('h8)
	) name2275 (
		\P2_reg1_reg[10]/NET0131 ,
		_w2247_,
		_w2737_
	);
	LUT2 #(
		.INIT('h8)
	) name2276 (
		\P2_reg0_reg[10]/NET0131 ,
		_w2245_,
		_w2738_
	);
	LUT2 #(
		.INIT('h8)
	) name2277 (
		\P2_reg2_reg[10]/NET0131 ,
		_w2243_,
		_w2739_
	);
	LUT2 #(
		.INIT('h1)
	) name2278 (
		_w2736_,
		_w2737_,
		_w2740_
	);
	LUT2 #(
		.INIT('h1)
	) name2279 (
		_w2738_,
		_w2739_,
		_w2741_
	);
	LUT2 #(
		.INIT('h8)
	) name2280 (
		_w2740_,
		_w2741_,
		_w2742_
	);
	LUT2 #(
		.INIT('h4)
	) name2281 (
		\P2_IR_reg[10]/NET0131 ,
		_w2689_,
		_w2743_
	);
	LUT2 #(
		.INIT('h2)
	) name2282 (
		\P2_IR_reg[10]/NET0131 ,
		_w2689_,
		_w2744_
	);
	LUT2 #(
		.INIT('h1)
	) name2283 (
		_w2743_,
		_w2744_,
		_w2745_
	);
	LUT2 #(
		.INIT('h8)
	) name2284 (
		_w2059_,
		_w2745_,
		_w2746_
	);
	LUT2 #(
		.INIT('h2)
	) name2285 (
		\P1_datao_reg[10]/NET0131 ,
		_w543_,
		_w2747_
	);
	LUT2 #(
		.INIT('h1)
	) name2286 (
		_w2144_,
		_w2152_,
		_w2748_
	);
	LUT2 #(
		.INIT('h4)
	) name2287 (
		_w2414_,
		_w2748_,
		_w2749_
	);
	LUT2 #(
		.INIT('h2)
	) name2288 (
		_w2414_,
		_w2748_,
		_w2750_
	);
	LUT2 #(
		.INIT('h2)
	) name2289 (
		_w543_,
		_w2749_,
		_w2751_
	);
	LUT2 #(
		.INIT('h4)
	) name2290 (
		_w2750_,
		_w2751_,
		_w2752_
	);
	LUT2 #(
		.INIT('h1)
	) name2291 (
		_w2747_,
		_w2752_,
		_w2753_
	);
	LUT2 #(
		.INIT('h4)
	) name2292 (
		_w2059_,
		_w2753_,
		_w2754_
	);
	LUT2 #(
		.INIT('h1)
	) name2293 (
		_w2746_,
		_w2754_,
		_w2755_
	);
	LUT2 #(
		.INIT('h2)
	) name2294 (
		_w2742_,
		_w2755_,
		_w2756_
	);
	LUT2 #(
		.INIT('h8)
	) name2295 (
		\P2_reg2_reg[9]/NET0131 ,
		_w2243_,
		_w2757_
	);
	LUT2 #(
		.INIT('h8)
	) name2296 (
		\P2_reg1_reg[9]/NET0131 ,
		_w2247_,
		_w2758_
	);
	LUT2 #(
		.INIT('h1)
	) name2297 (
		\P2_reg3_reg[9]/NET0131 ,
		_w2221_,
		_w2759_
	);
	LUT2 #(
		.INIT('h1)
	) name2298 (
		_w2222_,
		_w2759_,
		_w2760_
	);
	LUT2 #(
		.INIT('h8)
	) name2299 (
		_w2216_,
		_w2760_,
		_w2761_
	);
	LUT2 #(
		.INIT('h8)
	) name2300 (
		\P2_reg0_reg[9]/NET0131 ,
		_w2245_,
		_w2762_
	);
	LUT2 #(
		.INIT('h1)
	) name2301 (
		_w2757_,
		_w2758_,
		_w2763_
	);
	LUT2 #(
		.INIT('h1)
	) name2302 (
		_w2761_,
		_w2762_,
		_w2764_
	);
	LUT2 #(
		.INIT('h8)
	) name2303 (
		_w2763_,
		_w2764_,
		_w2765_
	);
	LUT2 #(
		.INIT('h2)
	) name2304 (
		\P2_IR_reg[31]/NET0131 ,
		_w2011_,
		_w2766_
	);
	LUT2 #(
		.INIT('h4)
	) name2305 (
		\P2_IR_reg[9]/NET0131 ,
		_w2766_,
		_w2767_
	);
	LUT2 #(
		.INIT('h2)
	) name2306 (
		\P2_IR_reg[9]/NET0131 ,
		_w2766_,
		_w2768_
	);
	LUT2 #(
		.INIT('h1)
	) name2307 (
		_w2767_,
		_w2768_,
		_w2769_
	);
	LUT2 #(
		.INIT('h8)
	) name2308 (
		_w2059_,
		_w2769_,
		_w2770_
	);
	LUT2 #(
		.INIT('h2)
	) name2309 (
		\P1_datao_reg[9]/NET0131 ,
		_w543_,
		_w2771_
	);
	LUT2 #(
		.INIT('h1)
	) name2310 (
		_w2146_,
		_w2153_,
		_w2772_
	);
	LUT2 #(
		.INIT('h4)
	) name2311 (
		_w2141_,
		_w2772_,
		_w2773_
	);
	LUT2 #(
		.INIT('h2)
	) name2312 (
		_w2141_,
		_w2772_,
		_w2774_
	);
	LUT2 #(
		.INIT('h2)
	) name2313 (
		_w543_,
		_w2773_,
		_w2775_
	);
	LUT2 #(
		.INIT('h4)
	) name2314 (
		_w2774_,
		_w2775_,
		_w2776_
	);
	LUT2 #(
		.INIT('h1)
	) name2315 (
		_w2771_,
		_w2776_,
		_w2777_
	);
	LUT2 #(
		.INIT('h4)
	) name2316 (
		_w2059_,
		_w2777_,
		_w2778_
	);
	LUT2 #(
		.INIT('h1)
	) name2317 (
		_w2770_,
		_w2778_,
		_w2779_
	);
	LUT2 #(
		.INIT('h2)
	) name2318 (
		_w2765_,
		_w2779_,
		_w2780_
	);
	LUT2 #(
		.INIT('h1)
	) name2319 (
		_w2756_,
		_w2780_,
		_w2781_
	);
	LUT2 #(
		.INIT('h8)
	) name2320 (
		_w2733_,
		_w2781_,
		_w2782_
	);
	LUT2 #(
		.INIT('h4)
	) name2321 (
		_w2678_,
		_w2782_,
		_w2783_
	);
	LUT2 #(
		.INIT('h4)
	) name2322 (
		_w2742_,
		_w2755_,
		_w2784_
	);
	LUT2 #(
		.INIT('h4)
	) name2323 (
		_w2765_,
		_w2779_,
		_w2785_
	);
	LUT2 #(
		.INIT('h4)
	) name2324 (
		_w2756_,
		_w2785_,
		_w2786_
	);
	LUT2 #(
		.INIT('h1)
	) name2325 (
		_w2784_,
		_w2786_,
		_w2787_
	);
	LUT2 #(
		.INIT('h2)
	) name2326 (
		_w2733_,
		_w2787_,
		_w2788_
	);
	LUT2 #(
		.INIT('h4)
	) name2327 (
		_w2715_,
		_w2731_,
		_w2789_
	);
	LUT2 #(
		.INIT('h4)
	) name2328 (
		_w2688_,
		_w2704_,
		_w2790_
	);
	LUT2 #(
		.INIT('h1)
	) name2329 (
		_w2789_,
		_w2790_,
		_w2791_
	);
	LUT2 #(
		.INIT('h1)
	) name2330 (
		_w2732_,
		_w2791_,
		_w2792_
	);
	LUT2 #(
		.INIT('h1)
	) name2331 (
		_w2788_,
		_w2792_,
		_w2793_
	);
	LUT2 #(
		.INIT('h4)
	) name2332 (
		_w2783_,
		_w2793_,
		_w2794_
	);
	LUT2 #(
		.INIT('h8)
	) name2333 (
		\P2_reg3_reg[15]/NET0131 ,
		_w2227_,
		_w2795_
	);
	LUT2 #(
		.INIT('h1)
	) name2334 (
		\P2_reg3_reg[16]/NET0131 ,
		_w2795_,
		_w2796_
	);
	LUT2 #(
		.INIT('h1)
	) name2335 (
		_w2229_,
		_w2796_,
		_w2797_
	);
	LUT2 #(
		.INIT('h8)
	) name2336 (
		_w2216_,
		_w2797_,
		_w2798_
	);
	LUT2 #(
		.INIT('h8)
	) name2337 (
		\P2_reg0_reg[16]/NET0131 ,
		_w2245_,
		_w2799_
	);
	LUT2 #(
		.INIT('h8)
	) name2338 (
		\P2_reg2_reg[16]/NET0131 ,
		_w2243_,
		_w2800_
	);
	LUT2 #(
		.INIT('h8)
	) name2339 (
		\P2_reg1_reg[16]/NET0131 ,
		_w2247_,
		_w2801_
	);
	LUT2 #(
		.INIT('h1)
	) name2340 (
		_w2798_,
		_w2799_,
		_w2802_
	);
	LUT2 #(
		.INIT('h1)
	) name2341 (
		_w2800_,
		_w2801_,
		_w2803_
	);
	LUT2 #(
		.INIT('h8)
	) name2342 (
		_w2802_,
		_w2803_,
		_w2804_
	);
	LUT2 #(
		.INIT('h2)
	) name2343 (
		\P2_IR_reg[31]/NET0131 ,
		_w1973_,
		_w2805_
	);
	LUT2 #(
		.INIT('h8)
	) name2344 (
		\P2_IR_reg[16]/NET0131 ,
		_w2805_,
		_w2806_
	);
	LUT2 #(
		.INIT('h1)
	) name2345 (
		\P2_IR_reg[16]/NET0131 ,
		_w2805_,
		_w2807_
	);
	LUT2 #(
		.INIT('h1)
	) name2346 (
		_w2806_,
		_w2807_,
		_w2808_
	);
	LUT2 #(
		.INIT('h2)
	) name2347 (
		_w2059_,
		_w2808_,
		_w2809_
	);
	LUT2 #(
		.INIT('h2)
	) name2348 (
		\P1_datao_reg[16]/NET0131 ,
		_w543_,
		_w2810_
	);
	LUT2 #(
		.INIT('h1)
	) name2349 (
		_w2084_,
		_w2086_,
		_w2811_
	);
	LUT2 #(
		.INIT('h4)
	) name2350 (
		_w2347_,
		_w2811_,
		_w2812_
	);
	LUT2 #(
		.INIT('h2)
	) name2351 (
		_w2347_,
		_w2811_,
		_w2813_
	);
	LUT2 #(
		.INIT('h2)
	) name2352 (
		_w543_,
		_w2812_,
		_w2814_
	);
	LUT2 #(
		.INIT('h4)
	) name2353 (
		_w2813_,
		_w2814_,
		_w2815_
	);
	LUT2 #(
		.INIT('h1)
	) name2354 (
		_w2810_,
		_w2815_,
		_w2816_
	);
	LUT2 #(
		.INIT('h4)
	) name2355 (
		_w2059_,
		_w2816_,
		_w2817_
	);
	LUT2 #(
		.INIT('h1)
	) name2356 (
		_w2809_,
		_w2817_,
		_w2818_
	);
	LUT2 #(
		.INIT('h2)
	) name2357 (
		_w2804_,
		_w2818_,
		_w2819_
	);
	LUT2 #(
		.INIT('h8)
	) name2358 (
		\P2_reg2_reg[15]/NET0131 ,
		_w2243_,
		_w2820_
	);
	LUT2 #(
		.INIT('h1)
	) name2359 (
		\P2_reg3_reg[15]/NET0131 ,
		_w2227_,
		_w2821_
	);
	LUT2 #(
		.INIT('h1)
	) name2360 (
		_w2795_,
		_w2821_,
		_w2822_
	);
	LUT2 #(
		.INIT('h8)
	) name2361 (
		_w2216_,
		_w2822_,
		_w2823_
	);
	LUT2 #(
		.INIT('h8)
	) name2362 (
		\P2_reg1_reg[15]/NET0131 ,
		_w2247_,
		_w2824_
	);
	LUT2 #(
		.INIT('h8)
	) name2363 (
		\P2_reg0_reg[15]/NET0131 ,
		_w2245_,
		_w2825_
	);
	LUT2 #(
		.INIT('h1)
	) name2364 (
		_w2820_,
		_w2823_,
		_w2826_
	);
	LUT2 #(
		.INIT('h1)
	) name2365 (
		_w2824_,
		_w2825_,
		_w2827_
	);
	LUT2 #(
		.INIT('h8)
	) name2366 (
		_w2826_,
		_w2827_,
		_w2828_
	);
	LUT2 #(
		.INIT('h2)
	) name2367 (
		\P2_IR_reg[31]/NET0131 ,
		_w1972_,
		_w2829_
	);
	LUT2 #(
		.INIT('h8)
	) name2368 (
		\P2_IR_reg[15]/NET0131 ,
		_w2829_,
		_w2830_
	);
	LUT2 #(
		.INIT('h1)
	) name2369 (
		\P2_IR_reg[15]/NET0131 ,
		_w2829_,
		_w2831_
	);
	LUT2 #(
		.INIT('h1)
	) name2370 (
		_w2830_,
		_w2831_,
		_w2832_
	);
	LUT2 #(
		.INIT('h2)
	) name2371 (
		_w2059_,
		_w2832_,
		_w2833_
	);
	LUT2 #(
		.INIT('h2)
	) name2372 (
		\P1_datao_reg[15]/NET0131 ,
		_w543_,
		_w2834_
	);
	LUT2 #(
		.INIT('h1)
	) name2373 (
		_w2279_,
		_w2285_,
		_w2835_
	);
	LUT2 #(
		.INIT('h1)
	) name2374 (
		_w2085_,
		_w2089_,
		_w2836_
	);
	LUT2 #(
		.INIT('h2)
	) name2375 (
		_w2835_,
		_w2836_,
		_w2837_
	);
	LUT2 #(
		.INIT('h4)
	) name2376 (
		_w2835_,
		_w2836_,
		_w2838_
	);
	LUT2 #(
		.INIT('h2)
	) name2377 (
		_w543_,
		_w2837_,
		_w2839_
	);
	LUT2 #(
		.INIT('h4)
	) name2378 (
		_w2838_,
		_w2839_,
		_w2840_
	);
	LUT2 #(
		.INIT('h1)
	) name2379 (
		_w2834_,
		_w2840_,
		_w2841_
	);
	LUT2 #(
		.INIT('h4)
	) name2380 (
		_w2059_,
		_w2841_,
		_w2842_
	);
	LUT2 #(
		.INIT('h1)
	) name2381 (
		_w2833_,
		_w2842_,
		_w2843_
	);
	LUT2 #(
		.INIT('h2)
	) name2382 (
		_w2828_,
		_w2843_,
		_w2844_
	);
	LUT2 #(
		.INIT('h1)
	) name2383 (
		_w2819_,
		_w2844_,
		_w2845_
	);
	LUT2 #(
		.INIT('h2)
	) name2384 (
		\P2_IR_reg[31]/NET0131 ,
		_w1971_,
		_w2846_
	);
	LUT2 #(
		.INIT('h8)
	) name2385 (
		\P2_IR_reg[14]/NET0131 ,
		_w2846_,
		_w2847_
	);
	LUT2 #(
		.INIT('h1)
	) name2386 (
		\P2_IR_reg[14]/NET0131 ,
		_w2846_,
		_w2848_
	);
	LUT2 #(
		.INIT('h1)
	) name2387 (
		_w2847_,
		_w2848_,
		_w2849_
	);
	LUT2 #(
		.INIT('h2)
	) name2388 (
		_w2059_,
		_w2849_,
		_w2850_
	);
	LUT2 #(
		.INIT('h2)
	) name2389 (
		\P1_datao_reg[14]/NET0131 ,
		_w543_,
		_w2851_
	);
	LUT2 #(
		.INIT('h4)
	) name2390 (
		_w2416_,
		_w2423_,
		_w2852_
	);
	LUT2 #(
		.INIT('h1)
	) name2391 (
		_w2088_,
		_w2092_,
		_w2853_
	);
	LUT2 #(
		.INIT('h2)
	) name2392 (
		_w2852_,
		_w2853_,
		_w2854_
	);
	LUT2 #(
		.INIT('h4)
	) name2393 (
		_w2852_,
		_w2853_,
		_w2855_
	);
	LUT2 #(
		.INIT('h2)
	) name2394 (
		_w543_,
		_w2854_,
		_w2856_
	);
	LUT2 #(
		.INIT('h4)
	) name2395 (
		_w2855_,
		_w2856_,
		_w2857_
	);
	LUT2 #(
		.INIT('h1)
	) name2396 (
		_w2851_,
		_w2857_,
		_w2858_
	);
	LUT2 #(
		.INIT('h4)
	) name2397 (
		_w2059_,
		_w2858_,
		_w2859_
	);
	LUT2 #(
		.INIT('h1)
	) name2398 (
		_w2850_,
		_w2859_,
		_w2860_
	);
	LUT2 #(
		.INIT('h8)
	) name2399 (
		\P2_reg2_reg[14]/NET0131 ,
		_w2243_,
		_w2861_
	);
	LUT2 #(
		.INIT('h8)
	) name2400 (
		\P2_reg1_reg[14]/NET0131 ,
		_w2247_,
		_w2862_
	);
	LUT2 #(
		.INIT('h8)
	) name2401 (
		\P2_reg0_reg[14]/NET0131 ,
		_w2245_,
		_w2863_
	);
	LUT2 #(
		.INIT('h8)
	) name2402 (
		\P2_reg3_reg[13]/NET0131 ,
		_w2707_,
		_w2864_
	);
	LUT2 #(
		.INIT('h1)
	) name2403 (
		\P2_reg3_reg[14]/NET0131 ,
		_w2864_,
		_w2865_
	);
	LUT2 #(
		.INIT('h1)
	) name2404 (
		_w2227_,
		_w2865_,
		_w2866_
	);
	LUT2 #(
		.INIT('h8)
	) name2405 (
		_w2216_,
		_w2866_,
		_w2867_
	);
	LUT2 #(
		.INIT('h1)
	) name2406 (
		_w2861_,
		_w2862_,
		_w2868_
	);
	LUT2 #(
		.INIT('h4)
	) name2407 (
		_w2863_,
		_w2868_,
		_w2869_
	);
	LUT2 #(
		.INIT('h4)
	) name2408 (
		_w2867_,
		_w2869_,
		_w2870_
	);
	LUT2 #(
		.INIT('h4)
	) name2409 (
		_w2860_,
		_w2870_,
		_w2871_
	);
	LUT2 #(
		.INIT('h8)
	) name2410 (
		\P2_reg2_reg[13]/NET0131 ,
		_w2243_,
		_w2872_
	);
	LUT2 #(
		.INIT('h1)
	) name2411 (
		\P2_reg3_reg[13]/NET0131 ,
		_w2707_,
		_w2873_
	);
	LUT2 #(
		.INIT('h1)
	) name2412 (
		_w2864_,
		_w2873_,
		_w2874_
	);
	LUT2 #(
		.INIT('h8)
	) name2413 (
		_w2216_,
		_w2874_,
		_w2875_
	);
	LUT2 #(
		.INIT('h8)
	) name2414 (
		\P2_reg1_reg[13]/NET0131 ,
		_w2247_,
		_w2876_
	);
	LUT2 #(
		.INIT('h8)
	) name2415 (
		\P2_reg0_reg[13]/NET0131 ,
		_w2245_,
		_w2877_
	);
	LUT2 #(
		.INIT('h1)
	) name2416 (
		_w2872_,
		_w2875_,
		_w2878_
	);
	LUT2 #(
		.INIT('h1)
	) name2417 (
		_w2876_,
		_w2877_,
		_w2879_
	);
	LUT2 #(
		.INIT('h8)
	) name2418 (
		_w2878_,
		_w2879_,
		_w2880_
	);
	LUT2 #(
		.INIT('h2)
	) name2419 (
		\P2_IR_reg[13]/NET0131 ,
		_w2380_,
		_w2881_
	);
	LUT2 #(
		.INIT('h4)
	) name2420 (
		\P2_IR_reg[13]/NET0131 ,
		_w2380_,
		_w2882_
	);
	LUT2 #(
		.INIT('h1)
	) name2421 (
		_w2881_,
		_w2882_,
		_w2883_
	);
	LUT2 #(
		.INIT('h8)
	) name2422 (
		_w2059_,
		_w2883_,
		_w2884_
	);
	LUT2 #(
		.INIT('h2)
	) name2423 (
		\P1_datao_reg[13]/NET0131 ,
		_w543_,
		_w2885_
	);
	LUT2 #(
		.INIT('h1)
	) name2424 (
		_w2091_,
		_w2161_,
		_w2886_
	);
	LUT2 #(
		.INIT('h4)
	) name2425 (
		_w2160_,
		_w2886_,
		_w2887_
	);
	LUT2 #(
		.INIT('h2)
	) name2426 (
		_w2160_,
		_w2886_,
		_w2888_
	);
	LUT2 #(
		.INIT('h2)
	) name2427 (
		_w543_,
		_w2887_,
		_w2889_
	);
	LUT2 #(
		.INIT('h4)
	) name2428 (
		_w2888_,
		_w2889_,
		_w2890_
	);
	LUT2 #(
		.INIT('h1)
	) name2429 (
		_w2885_,
		_w2890_,
		_w2891_
	);
	LUT2 #(
		.INIT('h4)
	) name2430 (
		_w2059_,
		_w2891_,
		_w2892_
	);
	LUT2 #(
		.INIT('h1)
	) name2431 (
		_w2884_,
		_w2892_,
		_w2893_
	);
	LUT2 #(
		.INIT('h2)
	) name2432 (
		_w2880_,
		_w2893_,
		_w2894_
	);
	LUT2 #(
		.INIT('h1)
	) name2433 (
		_w2871_,
		_w2894_,
		_w2895_
	);
	LUT2 #(
		.INIT('h8)
	) name2434 (
		_w2845_,
		_w2895_,
		_w2896_
	);
	LUT2 #(
		.INIT('h4)
	) name2435 (
		_w2794_,
		_w2896_,
		_w2897_
	);
	LUT2 #(
		.INIT('h8)
	) name2436 (
		_w2445_,
		_w2897_,
		_w2898_
	);
	LUT2 #(
		.INIT('h2)
	) name2437 (
		_w2860_,
		_w2870_,
		_w2899_
	);
	LUT2 #(
		.INIT('h4)
	) name2438 (
		_w2880_,
		_w2893_,
		_w2900_
	);
	LUT2 #(
		.INIT('h4)
	) name2439 (
		_w2871_,
		_w2900_,
		_w2901_
	);
	LUT2 #(
		.INIT('h1)
	) name2440 (
		_w2899_,
		_w2901_,
		_w2902_
	);
	LUT2 #(
		.INIT('h2)
	) name2441 (
		_w2845_,
		_w2902_,
		_w2903_
	);
	LUT2 #(
		.INIT('h4)
	) name2442 (
		_w2804_,
		_w2818_,
		_w2904_
	);
	LUT2 #(
		.INIT('h4)
	) name2443 (
		_w2828_,
		_w2843_,
		_w2905_
	);
	LUT2 #(
		.INIT('h4)
	) name2444 (
		_w2819_,
		_w2905_,
		_w2906_
	);
	LUT2 #(
		.INIT('h1)
	) name2445 (
		_w2904_,
		_w2906_,
		_w2907_
	);
	LUT2 #(
		.INIT('h4)
	) name2446 (
		_w2903_,
		_w2907_,
		_w2908_
	);
	LUT2 #(
		.INIT('h2)
	) name2447 (
		_w2445_,
		_w2908_,
		_w2909_
	);
	LUT2 #(
		.INIT('h2)
	) name2448 (
		_w2433_,
		_w2442_,
		_w2910_
	);
	LUT2 #(
		.INIT('h4)
	) name2449 (
		_w2379_,
		_w2399_,
		_w2911_
	);
	LUT2 #(
		.INIT('h1)
	) name2450 (
		_w2910_,
		_w2911_,
		_w2912_
	);
	LUT2 #(
		.INIT('h1)
	) name2451 (
		_w2443_,
		_w2912_,
		_w2913_
	);
	LUT2 #(
		.INIT('h8)
	) name2452 (
		_w2370_,
		_w2913_,
		_w2914_
	);
	LUT2 #(
		.INIT('h2)
	) name2453 (
		_w2358_,
		_w2368_,
		_w2915_
	);
	LUT2 #(
		.INIT('h2)
	) name2454 (
		_w2299_,
		_w2311_,
		_w2916_
	);
	LUT2 #(
		.INIT('h4)
	) name2455 (
		_w2369_,
		_w2916_,
		_w2917_
	);
	LUT2 #(
		.INIT('h1)
	) name2456 (
		_w2915_,
		_w2917_,
		_w2918_
	);
	LUT2 #(
		.INIT('h4)
	) name2457 (
		_w2914_,
		_w2918_,
		_w2919_
	);
	LUT2 #(
		.INIT('h4)
	) name2458 (
		_w2909_,
		_w2919_,
		_w2920_
	);
	LUT2 #(
		.INIT('h4)
	) name2459 (
		_w2898_,
		_w2920_,
		_w2921_
	);
	LUT2 #(
		.INIT('h2)
	) name2460 (
		\P1_datao_reg[28]/NET0131 ,
		_w543_,
		_w2922_
	);
	LUT2 #(
		.INIT('h1)
	) name2461 (
		_w2064_,
		_w2171_,
		_w2923_
	);
	LUT2 #(
		.INIT('h1)
	) name2462 (
		_w2170_,
		_w2173_,
		_w2924_
	);
	LUT2 #(
		.INIT('h1)
	) name2463 (
		_w2174_,
		_w2183_,
		_w2925_
	);
	LUT2 #(
		.INIT('h1)
	) name2464 (
		_w2074_,
		_w2925_,
		_w2926_
	);
	LUT2 #(
		.INIT('h4)
	) name2465 (
		_w2073_,
		_w2926_,
		_w2927_
	);
	LUT2 #(
		.INIT('h2)
	) name2466 (
		_w2924_,
		_w2927_,
		_w2928_
	);
	LUT2 #(
		.INIT('h1)
	) name2467 (
		_w2072_,
		_w2928_,
		_w2929_
	);
	LUT2 #(
		.INIT('h1)
	) name2468 (
		_w2065_,
		_w2068_,
		_w2930_
	);
	LUT2 #(
		.INIT('h1)
	) name2469 (
		_w2069_,
		_w2078_,
		_w2931_
	);
	LUT2 #(
		.INIT('h8)
	) name2470 (
		_w2930_,
		_w2931_,
		_w2932_
	);
	LUT2 #(
		.INIT('h4)
	) name2471 (
		_w2351_,
		_w2932_,
		_w2933_
	);
	LUT2 #(
		.INIT('h1)
	) name2472 (
		_w2177_,
		_w2182_,
		_w2934_
	);
	LUT2 #(
		.INIT('h1)
	) name2473 (
		_w2065_,
		_w2934_,
		_w2935_
	);
	LUT2 #(
		.INIT('h1)
	) name2474 (
		_w2099_,
		_w2178_,
		_w2936_
	);
	LUT2 #(
		.INIT('h1)
	) name2475 (
		_w2069_,
		_w2936_,
		_w2937_
	);
	LUT2 #(
		.INIT('h8)
	) name2476 (
		_w2930_,
		_w2937_,
		_w2938_
	);
	LUT2 #(
		.INIT('h1)
	) name2477 (
		_w2935_,
		_w2938_,
		_w2939_
	);
	LUT2 #(
		.INIT('h4)
	) name2478 (
		_w2933_,
		_w2939_,
		_w2940_
	);
	LUT2 #(
		.INIT('h4)
	) name2479 (
		_w2066_,
		_w2076_,
		_w2941_
	);
	LUT2 #(
		.INIT('h4)
	) name2480 (
		_w2940_,
		_w2941_,
		_w2942_
	);
	LUT2 #(
		.INIT('h1)
	) name2481 (
		_w2929_,
		_w2942_,
		_w2943_
	);
	LUT2 #(
		.INIT('h2)
	) name2482 (
		_w2923_,
		_w2943_,
		_w2944_
	);
	LUT2 #(
		.INIT('h4)
	) name2483 (
		_w2923_,
		_w2943_,
		_w2945_
	);
	LUT2 #(
		.INIT('h2)
	) name2484 (
		_w543_,
		_w2944_,
		_w2946_
	);
	LUT2 #(
		.INIT('h4)
	) name2485 (
		_w2945_,
		_w2946_,
		_w2947_
	);
	LUT2 #(
		.INIT('h1)
	) name2486 (
		_w2922_,
		_w2947_,
		_w2948_
	);
	LUT2 #(
		.INIT('h1)
	) name2487 (
		_w2059_,
		_w2948_,
		_w2949_
	);
	LUT2 #(
		.INIT('h8)
	) name2488 (
		\P2_reg0_reg[28]/NET0131 ,
		_w2245_,
		_w2950_
	);
	LUT2 #(
		.INIT('h8)
	) name2489 (
		\P2_reg2_reg[28]/NET0131 ,
		_w2243_,
		_w2951_
	);
	LUT2 #(
		.INIT('h8)
	) name2490 (
		\P2_reg1_reg[28]/NET0131 ,
		_w2247_,
		_w2952_
	);
	LUT2 #(
		.INIT('h8)
	) name2491 (
		\P2_reg3_reg[25]/NET0131 ,
		_w2237_,
		_w2953_
	);
	LUT2 #(
		.INIT('h8)
	) name2492 (
		\P2_reg3_reg[26]/NET0131 ,
		_w2953_,
		_w2954_
	);
	LUT2 #(
		.INIT('h8)
	) name2493 (
		\P2_reg3_reg[27]/NET0131 ,
		_w2954_,
		_w2955_
	);
	LUT2 #(
		.INIT('h2)
	) name2494 (
		\P2_reg3_reg[28]/NET0131 ,
		_w2955_,
		_w2956_
	);
	LUT2 #(
		.INIT('h4)
	) name2495 (
		\P2_reg3_reg[28]/NET0131 ,
		_w2955_,
		_w2957_
	);
	LUT2 #(
		.INIT('h1)
	) name2496 (
		_w2956_,
		_w2957_,
		_w2958_
	);
	LUT2 #(
		.INIT('h2)
	) name2497 (
		_w2216_,
		_w2958_,
		_w2959_
	);
	LUT2 #(
		.INIT('h1)
	) name2498 (
		_w2950_,
		_w2951_,
		_w2960_
	);
	LUT2 #(
		.INIT('h4)
	) name2499 (
		_w2952_,
		_w2960_,
		_w2961_
	);
	LUT2 #(
		.INIT('h4)
	) name2500 (
		_w2959_,
		_w2961_,
		_w2962_
	);
	LUT2 #(
		.INIT('h4)
	) name2501 (
		_w2949_,
		_w2962_,
		_w2963_
	);
	LUT2 #(
		.INIT('h2)
	) name2502 (
		\P1_datao_reg[27]/NET0131 ,
		_w543_,
		_w2964_
	);
	LUT2 #(
		.INIT('h1)
	) name2503 (
		_w2072_,
		_w2170_,
		_w2965_
	);
	LUT2 #(
		.INIT('h8)
	) name2504 (
		_w2075_,
		_w2185_,
		_w2966_
	);
	LUT2 #(
		.INIT('h1)
	) name2505 (
		_w2176_,
		_w2966_,
		_w2967_
	);
	LUT2 #(
		.INIT('h8)
	) name2506 (
		_w2067_,
		_w2075_,
		_w2968_
	);
	LUT2 #(
		.INIT('h8)
	) name2507 (
		_w2070_,
		_w2101_,
		_w2969_
	);
	LUT2 #(
		.INIT('h1)
	) name2508 (
		_w2180_,
		_w2969_,
		_w2970_
	);
	LUT2 #(
		.INIT('h1)
	) name2509 (
		_w2068_,
		_w2080_,
		_w2971_
	);
	LUT2 #(
		.INIT('h8)
	) name2510 (
		_w2931_,
		_w2971_,
		_w2972_
	);
	LUT2 #(
		.INIT('h4)
	) name2511 (
		_w2291_,
		_w2972_,
		_w2973_
	);
	LUT2 #(
		.INIT('h2)
	) name2512 (
		_w2970_,
		_w2973_,
		_w2974_
	);
	LUT2 #(
		.INIT('h2)
	) name2513 (
		_w2968_,
		_w2974_,
		_w2975_
	);
	LUT2 #(
		.INIT('h2)
	) name2514 (
		_w2967_,
		_w2975_,
		_w2976_
	);
	LUT2 #(
		.INIT('h2)
	) name2515 (
		_w2965_,
		_w2976_,
		_w2977_
	);
	LUT2 #(
		.INIT('h4)
	) name2516 (
		_w2965_,
		_w2976_,
		_w2978_
	);
	LUT2 #(
		.INIT('h2)
	) name2517 (
		_w543_,
		_w2977_,
		_w2979_
	);
	LUT2 #(
		.INIT('h4)
	) name2518 (
		_w2978_,
		_w2979_,
		_w2980_
	);
	LUT2 #(
		.INIT('h1)
	) name2519 (
		_w2964_,
		_w2980_,
		_w2981_
	);
	LUT2 #(
		.INIT('h1)
	) name2520 (
		_w2059_,
		_w2981_,
		_w2982_
	);
	LUT2 #(
		.INIT('h8)
	) name2521 (
		\P2_reg0_reg[27]/NET0131 ,
		_w2245_,
		_w2983_
	);
	LUT2 #(
		.INIT('h8)
	) name2522 (
		\P2_reg1_reg[27]/NET0131 ,
		_w2247_,
		_w2984_
	);
	LUT2 #(
		.INIT('h8)
	) name2523 (
		\P2_reg2_reg[27]/NET0131 ,
		_w2243_,
		_w2985_
	);
	LUT2 #(
		.INIT('h1)
	) name2524 (
		\P2_reg3_reg[27]/NET0131 ,
		_w2954_,
		_w2986_
	);
	LUT2 #(
		.INIT('h1)
	) name2525 (
		_w2955_,
		_w2986_,
		_w2987_
	);
	LUT2 #(
		.INIT('h8)
	) name2526 (
		_w2216_,
		_w2987_,
		_w2988_
	);
	LUT2 #(
		.INIT('h1)
	) name2527 (
		_w2983_,
		_w2984_,
		_w2989_
	);
	LUT2 #(
		.INIT('h4)
	) name2528 (
		_w2985_,
		_w2989_,
		_w2990_
	);
	LUT2 #(
		.INIT('h4)
	) name2529 (
		_w2988_,
		_w2990_,
		_w2991_
	);
	LUT2 #(
		.INIT('h4)
	) name2530 (
		_w2982_,
		_w2991_,
		_w2992_
	);
	LUT2 #(
		.INIT('h1)
	) name2531 (
		_w2963_,
		_w2992_,
		_w2993_
	);
	LUT2 #(
		.INIT('h2)
	) name2532 (
		\P1_datao_reg[26]/NET0131 ,
		_w543_,
		_w2994_
	);
	LUT2 #(
		.INIT('h1)
	) name2533 (
		_w2073_,
		_w2173_,
		_w2995_
	);
	LUT2 #(
		.INIT('h1)
	) name2534 (
		_w2066_,
		_w2074_,
		_w2996_
	);
	LUT2 #(
		.INIT('h8)
	) name2535 (
		_w2935_,
		_w2996_,
		_w2997_
	);
	LUT2 #(
		.INIT('h1)
	) name2536 (
		_w2926_,
		_w2997_,
		_w2998_
	);
	LUT2 #(
		.INIT('h8)
	) name2537 (
		_w2930_,
		_w2996_,
		_w2999_
	);
	LUT2 #(
		.INIT('h4)
	) name2538 (
		_w2069_,
		_w2082_,
		_w3000_
	);
	LUT2 #(
		.INIT('h4)
	) name2539 (
		_w2426_,
		_w3000_,
		_w3001_
	);
	LUT2 #(
		.INIT('h8)
	) name2540 (
		_w2315_,
		_w2931_,
		_w3002_
	);
	LUT2 #(
		.INIT('h1)
	) name2541 (
		_w2937_,
		_w3002_,
		_w3003_
	);
	LUT2 #(
		.INIT('h4)
	) name2542 (
		_w3001_,
		_w3003_,
		_w3004_
	);
	LUT2 #(
		.INIT('h2)
	) name2543 (
		_w2999_,
		_w3004_,
		_w3005_
	);
	LUT2 #(
		.INIT('h2)
	) name2544 (
		_w2998_,
		_w3005_,
		_w3006_
	);
	LUT2 #(
		.INIT('h2)
	) name2545 (
		_w2995_,
		_w3006_,
		_w3007_
	);
	LUT2 #(
		.INIT('h4)
	) name2546 (
		_w2995_,
		_w3006_,
		_w3008_
	);
	LUT2 #(
		.INIT('h2)
	) name2547 (
		_w543_,
		_w3007_,
		_w3009_
	);
	LUT2 #(
		.INIT('h4)
	) name2548 (
		_w3008_,
		_w3009_,
		_w3010_
	);
	LUT2 #(
		.INIT('h1)
	) name2549 (
		_w2994_,
		_w3010_,
		_w3011_
	);
	LUT2 #(
		.INIT('h1)
	) name2550 (
		_w2059_,
		_w3011_,
		_w3012_
	);
	LUT2 #(
		.INIT('h8)
	) name2551 (
		\P2_reg0_reg[26]/NET0131 ,
		_w2245_,
		_w3013_
	);
	LUT2 #(
		.INIT('h8)
	) name2552 (
		\P2_reg1_reg[26]/NET0131 ,
		_w2247_,
		_w3014_
	);
	LUT2 #(
		.INIT('h8)
	) name2553 (
		\P2_reg2_reg[26]/NET0131 ,
		_w2243_,
		_w3015_
	);
	LUT2 #(
		.INIT('h1)
	) name2554 (
		\P2_reg3_reg[26]/NET0131 ,
		_w2953_,
		_w3016_
	);
	LUT2 #(
		.INIT('h1)
	) name2555 (
		_w2954_,
		_w3016_,
		_w3017_
	);
	LUT2 #(
		.INIT('h8)
	) name2556 (
		_w2216_,
		_w3017_,
		_w3018_
	);
	LUT2 #(
		.INIT('h1)
	) name2557 (
		_w3013_,
		_w3014_,
		_w3019_
	);
	LUT2 #(
		.INIT('h4)
	) name2558 (
		_w3015_,
		_w3019_,
		_w3020_
	);
	LUT2 #(
		.INIT('h4)
	) name2559 (
		_w3018_,
		_w3020_,
		_w3021_
	);
	LUT2 #(
		.INIT('h4)
	) name2560 (
		_w3012_,
		_w3021_,
		_w3022_
	);
	LUT2 #(
		.INIT('h2)
	) name2561 (
		\P1_datao_reg[25]/NET0131 ,
		_w543_,
		_w3023_
	);
	LUT2 #(
		.INIT('h1)
	) name2562 (
		_w2074_,
		_w2174_,
		_w3024_
	);
	LUT2 #(
		.INIT('h2)
	) name2563 (
		_w2083_,
		_w2391_,
		_w3025_
	);
	LUT2 #(
		.INIT('h2)
	) name2564 (
		_w2106_,
		_w3025_,
		_w3026_
	);
	LUT2 #(
		.INIT('h2)
	) name2565 (
		_w2071_,
		_w3026_,
		_w3027_
	);
	LUT2 #(
		.INIT('h2)
	) name2566 (
		_w2186_,
		_w3027_,
		_w3028_
	);
	LUT2 #(
		.INIT('h2)
	) name2567 (
		_w3024_,
		_w3028_,
		_w3029_
	);
	LUT2 #(
		.INIT('h4)
	) name2568 (
		_w3024_,
		_w3028_,
		_w3030_
	);
	LUT2 #(
		.INIT('h2)
	) name2569 (
		_w543_,
		_w3029_,
		_w3031_
	);
	LUT2 #(
		.INIT('h4)
	) name2570 (
		_w3030_,
		_w3031_,
		_w3032_
	);
	LUT2 #(
		.INIT('h1)
	) name2571 (
		_w3023_,
		_w3032_,
		_w3033_
	);
	LUT2 #(
		.INIT('h1)
	) name2572 (
		_w2059_,
		_w3033_,
		_w3034_
	);
	LUT2 #(
		.INIT('h8)
	) name2573 (
		\P2_reg0_reg[25]/NET0131 ,
		_w2245_,
		_w3035_
	);
	LUT2 #(
		.INIT('h8)
	) name2574 (
		\P2_reg1_reg[25]/NET0131 ,
		_w2247_,
		_w3036_
	);
	LUT2 #(
		.INIT('h8)
	) name2575 (
		\P2_reg2_reg[25]/NET0131 ,
		_w2243_,
		_w3037_
	);
	LUT2 #(
		.INIT('h1)
	) name2576 (
		\P2_reg3_reg[25]/NET0131 ,
		_w2237_,
		_w3038_
	);
	LUT2 #(
		.INIT('h1)
	) name2577 (
		_w2953_,
		_w3038_,
		_w3039_
	);
	LUT2 #(
		.INIT('h8)
	) name2578 (
		_w2216_,
		_w3039_,
		_w3040_
	);
	LUT2 #(
		.INIT('h1)
	) name2579 (
		_w3035_,
		_w3036_,
		_w3041_
	);
	LUT2 #(
		.INIT('h4)
	) name2580 (
		_w3037_,
		_w3041_,
		_w3042_
	);
	LUT2 #(
		.INIT('h4)
	) name2581 (
		_w3040_,
		_w3042_,
		_w3043_
	);
	LUT2 #(
		.INIT('h4)
	) name2582 (
		_w3034_,
		_w3043_,
		_w3044_
	);
	LUT2 #(
		.INIT('h1)
	) name2583 (
		_w3022_,
		_w3044_,
		_w3045_
	);
	LUT2 #(
		.INIT('h8)
	) name2584 (
		_w2993_,
		_w3045_,
		_w3046_
	);
	LUT2 #(
		.INIT('h2)
	) name2585 (
		\P1_datao_reg[24]/NET0131 ,
		_w543_,
		_w3047_
	);
	LUT2 #(
		.INIT('h1)
	) name2586 (
		_w2066_,
		_w2183_,
		_w3048_
	);
	LUT2 #(
		.INIT('h4)
	) name2587 (
		_w2940_,
		_w3048_,
		_w3049_
	);
	LUT2 #(
		.INIT('h2)
	) name2588 (
		_w2940_,
		_w3048_,
		_w3050_
	);
	LUT2 #(
		.INIT('h2)
	) name2589 (
		_w543_,
		_w3049_,
		_w3051_
	);
	LUT2 #(
		.INIT('h4)
	) name2590 (
		_w3050_,
		_w3051_,
		_w3052_
	);
	LUT2 #(
		.INIT('h1)
	) name2591 (
		_w3047_,
		_w3052_,
		_w3053_
	);
	LUT2 #(
		.INIT('h1)
	) name2592 (
		_w2059_,
		_w3053_,
		_w3054_
	);
	LUT2 #(
		.INIT('h8)
	) name2593 (
		_w2231_,
		_w2306_,
		_w3055_
	);
	LUT2 #(
		.INIT('h8)
	) name2594 (
		\P2_reg3_reg[23]/NET0131 ,
		_w3055_,
		_w3056_
	);
	LUT2 #(
		.INIT('h1)
	) name2595 (
		\P2_reg3_reg[24]/NET0131 ,
		_w3056_,
		_w3057_
	);
	LUT2 #(
		.INIT('h1)
	) name2596 (
		_w2237_,
		_w3057_,
		_w3058_
	);
	LUT2 #(
		.INIT('h8)
	) name2597 (
		_w2216_,
		_w3058_,
		_w3059_
	);
	LUT2 #(
		.INIT('h8)
	) name2598 (
		\P2_reg1_reg[24]/NET0131 ,
		_w2247_,
		_w3060_
	);
	LUT2 #(
		.INIT('h8)
	) name2599 (
		\P2_reg2_reg[24]/NET0131 ,
		_w2243_,
		_w3061_
	);
	LUT2 #(
		.INIT('h8)
	) name2600 (
		\P2_reg0_reg[24]/NET0131 ,
		_w2245_,
		_w3062_
	);
	LUT2 #(
		.INIT('h1)
	) name2601 (
		_w3060_,
		_w3061_,
		_w3063_
	);
	LUT2 #(
		.INIT('h4)
	) name2602 (
		_w3062_,
		_w3063_,
		_w3064_
	);
	LUT2 #(
		.INIT('h4)
	) name2603 (
		_w3059_,
		_w3064_,
		_w3065_
	);
	LUT2 #(
		.INIT('h4)
	) name2604 (
		_w3054_,
		_w3065_,
		_w3066_
	);
	LUT2 #(
		.INIT('h2)
	) name2605 (
		\P1_datao_reg[23]/NET0131 ,
		_w543_,
		_w3067_
	);
	LUT2 #(
		.INIT('h1)
	) name2606 (
		_w2065_,
		_w2182_,
		_w3068_
	);
	LUT2 #(
		.INIT('h8)
	) name2607 (
		_w2289_,
		_w2972_,
		_w3069_
	);
	LUT2 #(
		.INIT('h8)
	) name2608 (
		_w2263_,
		_w2972_,
		_w3070_
	);
	LUT2 #(
		.INIT('h4)
	) name2609 (
		_w2835_,
		_w3070_,
		_w3071_
	);
	LUT2 #(
		.INIT('h2)
	) name2610 (
		_w2970_,
		_w3069_,
		_w3072_
	);
	LUT2 #(
		.INIT('h4)
	) name2611 (
		_w3071_,
		_w3072_,
		_w3073_
	);
	LUT2 #(
		.INIT('h2)
	) name2612 (
		_w3068_,
		_w3073_,
		_w3074_
	);
	LUT2 #(
		.INIT('h4)
	) name2613 (
		_w3068_,
		_w3073_,
		_w3075_
	);
	LUT2 #(
		.INIT('h2)
	) name2614 (
		_w543_,
		_w3074_,
		_w3076_
	);
	LUT2 #(
		.INIT('h4)
	) name2615 (
		_w3075_,
		_w3076_,
		_w3077_
	);
	LUT2 #(
		.INIT('h1)
	) name2616 (
		_w3067_,
		_w3077_,
		_w3078_
	);
	LUT2 #(
		.INIT('h1)
	) name2617 (
		_w2059_,
		_w3078_,
		_w3079_
	);
	LUT2 #(
		.INIT('h8)
	) name2618 (
		\P2_reg0_reg[23]/NET0131 ,
		_w2245_,
		_w3080_
	);
	LUT2 #(
		.INIT('h8)
	) name2619 (
		\P2_reg2_reg[23]/NET0131 ,
		_w2243_,
		_w3081_
	);
	LUT2 #(
		.INIT('h8)
	) name2620 (
		\P2_reg1_reg[23]/NET0131 ,
		_w2247_,
		_w3082_
	);
	LUT2 #(
		.INIT('h1)
	) name2621 (
		\P2_reg3_reg[23]/NET0131 ,
		_w3055_,
		_w3083_
	);
	LUT2 #(
		.INIT('h1)
	) name2622 (
		_w3056_,
		_w3083_,
		_w3084_
	);
	LUT2 #(
		.INIT('h8)
	) name2623 (
		_w2216_,
		_w3084_,
		_w3085_
	);
	LUT2 #(
		.INIT('h1)
	) name2624 (
		_w3080_,
		_w3081_,
		_w3086_
	);
	LUT2 #(
		.INIT('h4)
	) name2625 (
		_w3082_,
		_w3086_,
		_w3087_
	);
	LUT2 #(
		.INIT('h4)
	) name2626 (
		_w3085_,
		_w3087_,
		_w3088_
	);
	LUT2 #(
		.INIT('h4)
	) name2627 (
		_w3079_,
		_w3088_,
		_w3089_
	);
	LUT2 #(
		.INIT('h1)
	) name2628 (
		_w3066_,
		_w3089_,
		_w3090_
	);
	LUT2 #(
		.INIT('h2)
	) name2629 (
		\P1_datao_reg[22]/NET0131 ,
		_w543_,
		_w3091_
	);
	LUT2 #(
		.INIT('h1)
	) name2630 (
		_w2068_,
		_w2177_,
		_w3092_
	);
	LUT2 #(
		.INIT('h2)
	) name2631 (
		_w2417_,
		_w2852_,
		_w3093_
	);
	LUT2 #(
		.INIT('h2)
	) name2632 (
		_w2420_,
		_w3093_,
		_w3094_
	);
	LUT2 #(
		.INIT('h2)
	) name2633 (
		_w3000_,
		_w3094_,
		_w3095_
	);
	LUT2 #(
		.INIT('h2)
	) name2634 (
		_w3003_,
		_w3095_,
		_w3096_
	);
	LUT2 #(
		.INIT('h2)
	) name2635 (
		_w3092_,
		_w3096_,
		_w3097_
	);
	LUT2 #(
		.INIT('h4)
	) name2636 (
		_w3092_,
		_w3096_,
		_w3098_
	);
	LUT2 #(
		.INIT('h2)
	) name2637 (
		_w543_,
		_w3097_,
		_w3099_
	);
	LUT2 #(
		.INIT('h4)
	) name2638 (
		_w3098_,
		_w3099_,
		_w3100_
	);
	LUT2 #(
		.INIT('h1)
	) name2639 (
		_w3091_,
		_w3100_,
		_w3101_
	);
	LUT2 #(
		.INIT('h1)
	) name2640 (
		_w2059_,
		_w3101_,
		_w3102_
	);
	LUT2 #(
		.INIT('h8)
	) name2641 (
		\P2_reg0_reg[22]/NET0131 ,
		_w2245_,
		_w3103_
	);
	LUT2 #(
		.INIT('h8)
	) name2642 (
		\P2_reg1_reg[22]/NET0131 ,
		_w2247_,
		_w3104_
	);
	LUT2 #(
		.INIT('h8)
	) name2643 (
		\P2_reg2_reg[22]/NET0131 ,
		_w2243_,
		_w3105_
	);
	LUT2 #(
		.INIT('h8)
	) name2644 (
		_w2230_,
		_w2306_,
		_w3106_
	);
	LUT2 #(
		.INIT('h1)
	) name2645 (
		\P2_reg3_reg[22]/NET0131 ,
		_w3106_,
		_w3107_
	);
	LUT2 #(
		.INIT('h1)
	) name2646 (
		_w3055_,
		_w3107_,
		_w3108_
	);
	LUT2 #(
		.INIT('h8)
	) name2647 (
		_w2216_,
		_w3108_,
		_w3109_
	);
	LUT2 #(
		.INIT('h1)
	) name2648 (
		_w3103_,
		_w3104_,
		_w3110_
	);
	LUT2 #(
		.INIT('h4)
	) name2649 (
		_w3105_,
		_w3110_,
		_w3111_
	);
	LUT2 #(
		.INIT('h4)
	) name2650 (
		_w3109_,
		_w3111_,
		_w3112_
	);
	LUT2 #(
		.INIT('h4)
	) name2651 (
		_w3102_,
		_w3112_,
		_w3113_
	);
	LUT2 #(
		.INIT('h2)
	) name2652 (
		\P1_datao_reg[21]/NET0131 ,
		_w543_,
		_w3114_
	);
	LUT2 #(
		.INIT('h1)
	) name2653 (
		_w2069_,
		_w2178_,
		_w3115_
	);
	LUT2 #(
		.INIT('h4)
	) name2654 (
		_w2167_,
		_w3115_,
		_w3116_
	);
	LUT2 #(
		.INIT('h2)
	) name2655 (
		_w2167_,
		_w3115_,
		_w3117_
	);
	LUT2 #(
		.INIT('h2)
	) name2656 (
		_w543_,
		_w3116_,
		_w3118_
	);
	LUT2 #(
		.INIT('h4)
	) name2657 (
		_w3117_,
		_w3118_,
		_w3119_
	);
	LUT2 #(
		.INIT('h1)
	) name2658 (
		_w3114_,
		_w3119_,
		_w3120_
	);
	LUT2 #(
		.INIT('h1)
	) name2659 (
		_w2059_,
		_w3120_,
		_w3121_
	);
	LUT2 #(
		.INIT('h8)
	) name2660 (
		\P2_reg2_reg[21]/NET0131 ,
		_w2243_,
		_w3122_
	);
	LUT2 #(
		.INIT('h8)
	) name2661 (
		\P2_reg0_reg[21]/NET0131 ,
		_w2245_,
		_w3123_
	);
	LUT2 #(
		.INIT('h8)
	) name2662 (
		\P2_reg1_reg[21]/NET0131 ,
		_w2247_,
		_w3124_
	);
	LUT2 #(
		.INIT('h1)
	) name2663 (
		\P2_reg3_reg[21]/NET0131 ,
		_w2362_,
		_w3125_
	);
	LUT2 #(
		.INIT('h1)
	) name2664 (
		_w3106_,
		_w3125_,
		_w3126_
	);
	LUT2 #(
		.INIT('h8)
	) name2665 (
		_w2216_,
		_w3126_,
		_w3127_
	);
	LUT2 #(
		.INIT('h1)
	) name2666 (
		_w3122_,
		_w3123_,
		_w3128_
	);
	LUT2 #(
		.INIT('h4)
	) name2667 (
		_w3124_,
		_w3128_,
		_w3129_
	);
	LUT2 #(
		.INIT('h4)
	) name2668 (
		_w3127_,
		_w3129_,
		_w3130_
	);
	LUT2 #(
		.INIT('h4)
	) name2669 (
		_w3121_,
		_w3130_,
		_w3131_
	);
	LUT2 #(
		.INIT('h1)
	) name2670 (
		_w3113_,
		_w3131_,
		_w3132_
	);
	LUT2 #(
		.INIT('h8)
	) name2671 (
		_w3090_,
		_w3132_,
		_w3133_
	);
	LUT2 #(
		.INIT('h8)
	) name2672 (
		_w3046_,
		_w3133_,
		_w3134_
	);
	LUT2 #(
		.INIT('h4)
	) name2673 (
		_w2921_,
		_w3134_,
		_w3135_
	);
	LUT2 #(
		.INIT('h2)
	) name2674 (
		_w2982_,
		_w2991_,
		_w3136_
	);
	LUT2 #(
		.INIT('h4)
	) name2675 (
		_w2963_,
		_w3136_,
		_w3137_
	);
	LUT2 #(
		.INIT('h2)
	) name2676 (
		_w3102_,
		_w3112_,
		_w3138_
	);
	LUT2 #(
		.INIT('h2)
	) name2677 (
		_w3121_,
		_w3130_,
		_w3139_
	);
	LUT2 #(
		.INIT('h4)
	) name2678 (
		_w3113_,
		_w3139_,
		_w3140_
	);
	LUT2 #(
		.INIT('h1)
	) name2679 (
		_w3138_,
		_w3140_,
		_w3141_
	);
	LUT2 #(
		.INIT('h2)
	) name2680 (
		_w3090_,
		_w3141_,
		_w3142_
	);
	LUT2 #(
		.INIT('h2)
	) name2681 (
		_w3054_,
		_w3065_,
		_w3143_
	);
	LUT2 #(
		.INIT('h2)
	) name2682 (
		_w3079_,
		_w3088_,
		_w3144_
	);
	LUT2 #(
		.INIT('h4)
	) name2683 (
		_w3066_,
		_w3144_,
		_w3145_
	);
	LUT2 #(
		.INIT('h1)
	) name2684 (
		_w3143_,
		_w3145_,
		_w3146_
	);
	LUT2 #(
		.INIT('h4)
	) name2685 (
		_w3142_,
		_w3146_,
		_w3147_
	);
	LUT2 #(
		.INIT('h2)
	) name2686 (
		_w3046_,
		_w3147_,
		_w3148_
	);
	LUT2 #(
		.INIT('h2)
	) name2687 (
		_w3012_,
		_w3021_,
		_w3149_
	);
	LUT2 #(
		.INIT('h2)
	) name2688 (
		_w3034_,
		_w3043_,
		_w3150_
	);
	LUT2 #(
		.INIT('h4)
	) name2689 (
		_w3022_,
		_w3150_,
		_w3151_
	);
	LUT2 #(
		.INIT('h1)
	) name2690 (
		_w3149_,
		_w3151_,
		_w3152_
	);
	LUT2 #(
		.INIT('h2)
	) name2691 (
		_w2993_,
		_w3152_,
		_w3153_
	);
	LUT2 #(
		.INIT('h2)
	) name2692 (
		_w2949_,
		_w2962_,
		_w3154_
	);
	LUT2 #(
		.INIT('h1)
	) name2693 (
		_w3137_,
		_w3154_,
		_w3155_
	);
	LUT2 #(
		.INIT('h4)
	) name2694 (
		_w3153_,
		_w3155_,
		_w3156_
	);
	LUT2 #(
		.INIT('h4)
	) name2695 (
		_w3148_,
		_w3156_,
		_w3157_
	);
	LUT2 #(
		.INIT('h4)
	) name2696 (
		_w3135_,
		_w3157_,
		_w3158_
	);
	LUT2 #(
		.INIT('h2)
	) name2697 (
		_w2254_,
		_w3158_,
		_w3159_
	);
	LUT2 #(
		.INIT('h4)
	) name2698 (
		_w2254_,
		_w3158_,
		_w3160_
	);
	LUT2 #(
		.INIT('h1)
	) name2699 (
		_w3159_,
		_w3160_,
		_w3161_
	);
	LUT2 #(
		.INIT('h2)
	) name2700 (
		_w2040_,
		_w3161_,
		_w3162_
	);
	LUT2 #(
		.INIT('h1)
	) name2701 (
		_w2041_,
		_w3162_,
		_w3163_
	);
	LUT2 #(
		.INIT('h1)
	) name2702 (
		\P2_IR_reg[22]/NET0131 ,
		_w2199_,
		_w3164_
	);
	LUT2 #(
		.INIT('h8)
	) name2703 (
		\P2_IR_reg[22]/NET0131 ,
		_w2199_,
		_w3165_
	);
	LUT2 #(
		.INIT('h1)
	) name2704 (
		_w3164_,
		_w3165_,
		_w3166_
	);
	LUT2 #(
		.INIT('h4)
	) name2705 (
		_w1982_,
		_w3166_,
		_w3167_
	);
	LUT2 #(
		.INIT('h2)
	) name2706 (
		\P2_IR_reg[21]/NET0131 ,
		_w2208_,
		_w3168_
	);
	LUT2 #(
		.INIT('h4)
	) name2707 (
		\P2_IR_reg[21]/NET0131 ,
		_w2208_,
		_w3169_
	);
	LUT2 #(
		.INIT('h1)
	) name2708 (
		_w3168_,
		_w3169_,
		_w3170_
	);
	LUT2 #(
		.INIT('h8)
	) name2709 (
		_w3167_,
		_w3170_,
		_w3171_
	);
	LUT2 #(
		.INIT('h2)
	) name2710 (
		_w1982_,
		_w3166_,
		_w3172_
	);
	LUT2 #(
		.INIT('h2)
	) name2711 (
		\P2_IR_reg[20]/NET0131 ,
		_w2042_,
		_w3173_
	);
	LUT2 #(
		.INIT('h4)
	) name2712 (
		\P2_IR_reg[20]/NET0131 ,
		_w2042_,
		_w3174_
	);
	LUT2 #(
		.INIT('h1)
	) name2713 (
		_w3173_,
		_w3174_,
		_w3175_
	);
	LUT2 #(
		.INIT('h8)
	) name2714 (
		_w3172_,
		_w3175_,
		_w3176_
	);
	LUT2 #(
		.INIT('h1)
	) name2715 (
		_w3171_,
		_w3176_,
		_w3177_
	);
	LUT2 #(
		.INIT('h1)
	) name2716 (
		_w3163_,
		_w3177_,
		_w3178_
	);
	LUT2 #(
		.INIT('h8)
	) name2717 (
		_w2949_,
		_w2962_,
		_w3179_
	);
	LUT2 #(
		.INIT('h8)
	) name2718 (
		_w2982_,
		_w2991_,
		_w3180_
	);
	LUT2 #(
		.INIT('h1)
	) name2719 (
		_w3179_,
		_w3180_,
		_w3181_
	);
	LUT2 #(
		.INIT('h8)
	) name2720 (
		_w3012_,
		_w3021_,
		_w3182_
	);
	LUT2 #(
		.INIT('h8)
	) name2721 (
		_w3034_,
		_w3043_,
		_w3183_
	);
	LUT2 #(
		.INIT('h1)
	) name2722 (
		_w3182_,
		_w3183_,
		_w3184_
	);
	LUT2 #(
		.INIT('h8)
	) name2723 (
		_w3181_,
		_w3184_,
		_w3185_
	);
	LUT2 #(
		.INIT('h8)
	) name2724 (
		_w3079_,
		_w3088_,
		_w3186_
	);
	LUT2 #(
		.INIT('h8)
	) name2725 (
		_w3054_,
		_w3065_,
		_w3187_
	);
	LUT2 #(
		.INIT('h1)
	) name2726 (
		_w3186_,
		_w3187_,
		_w3188_
	);
	LUT2 #(
		.INIT('h8)
	) name2727 (
		_w3102_,
		_w3112_,
		_w3189_
	);
	LUT2 #(
		.INIT('h1)
	) name2728 (
		_w3102_,
		_w3112_,
		_w3190_
	);
	LUT2 #(
		.INIT('h1)
	) name2729 (
		_w3121_,
		_w3130_,
		_w3191_
	);
	LUT2 #(
		.INIT('h1)
	) name2730 (
		_w3190_,
		_w3191_,
		_w3192_
	);
	LUT2 #(
		.INIT('h1)
	) name2731 (
		_w3189_,
		_w3192_,
		_w3193_
	);
	LUT2 #(
		.INIT('h8)
	) name2732 (
		_w3188_,
		_w3193_,
		_w3194_
	);
	LUT2 #(
		.INIT('h1)
	) name2733 (
		_w3054_,
		_w3065_,
		_w3195_
	);
	LUT2 #(
		.INIT('h1)
	) name2734 (
		_w3079_,
		_w3088_,
		_w3196_
	);
	LUT2 #(
		.INIT('h4)
	) name2735 (
		_w3187_,
		_w3196_,
		_w3197_
	);
	LUT2 #(
		.INIT('h1)
	) name2736 (
		_w3195_,
		_w3197_,
		_w3198_
	);
	LUT2 #(
		.INIT('h4)
	) name2737 (
		_w3194_,
		_w3198_,
		_w3199_
	);
	LUT2 #(
		.INIT('h2)
	) name2738 (
		_w3185_,
		_w3199_,
		_w3200_
	);
	LUT2 #(
		.INIT('h1)
	) name2739 (
		_w3012_,
		_w3021_,
		_w3201_
	);
	LUT2 #(
		.INIT('h1)
	) name2740 (
		_w3034_,
		_w3043_,
		_w3202_
	);
	LUT2 #(
		.INIT('h1)
	) name2741 (
		_w3201_,
		_w3202_,
		_w3203_
	);
	LUT2 #(
		.INIT('h1)
	) name2742 (
		_w3182_,
		_w3203_,
		_w3204_
	);
	LUT2 #(
		.INIT('h8)
	) name2743 (
		_w3181_,
		_w3204_,
		_w3205_
	);
	LUT2 #(
		.INIT('h1)
	) name2744 (
		_w2949_,
		_w2962_,
		_w3206_
	);
	LUT2 #(
		.INIT('h1)
	) name2745 (
		_w2982_,
		_w2991_,
		_w3207_
	);
	LUT2 #(
		.INIT('h1)
	) name2746 (
		_w3206_,
		_w3207_,
		_w3208_
	);
	LUT2 #(
		.INIT('h1)
	) name2747 (
		_w3179_,
		_w3208_,
		_w3209_
	);
	LUT2 #(
		.INIT('h8)
	) name2748 (
		_w2299_,
		_w2311_,
		_w3210_
	);
	LUT2 #(
		.INIT('h8)
	) name2749 (
		_w2358_,
		_w2368_,
		_w3211_
	);
	LUT2 #(
		.INIT('h1)
	) name2750 (
		_w3210_,
		_w3211_,
		_w3212_
	);
	LUT2 #(
		.INIT('h8)
	) name2751 (
		_w2379_,
		_w2399_,
		_w3213_
	);
	LUT2 #(
		.INIT('h8)
	) name2752 (
		_w2433_,
		_w2442_,
		_w3214_
	);
	LUT2 #(
		.INIT('h1)
	) name2753 (
		_w3213_,
		_w3214_,
		_w3215_
	);
	LUT2 #(
		.INIT('h8)
	) name2754 (
		_w3212_,
		_w3215_,
		_w3216_
	);
	LUT2 #(
		.INIT('h8)
	) name2755 (
		_w2804_,
		_w2818_,
		_w3217_
	);
	LUT2 #(
		.INIT('h8)
	) name2756 (
		_w2828_,
		_w2843_,
		_w3218_
	);
	LUT2 #(
		.INIT('h1)
	) name2757 (
		_w3217_,
		_w3218_,
		_w3219_
	);
	LUT2 #(
		.INIT('h8)
	) name2758 (
		_w2860_,
		_w2870_,
		_w3220_
	);
	LUT2 #(
		.INIT('h8)
	) name2759 (
		_w2880_,
		_w2893_,
		_w3221_
	);
	LUT2 #(
		.INIT('h1)
	) name2760 (
		_w3220_,
		_w3221_,
		_w3222_
	);
	LUT2 #(
		.INIT('h8)
	) name2761 (
		_w3219_,
		_w3222_,
		_w3223_
	);
	LUT2 #(
		.INIT('h8)
	) name2762 (
		_w3216_,
		_w3223_,
		_w3224_
	);
	LUT2 #(
		.INIT('h8)
	) name2763 (
		_w2688_,
		_w2704_,
		_w3225_
	);
	LUT2 #(
		.INIT('h8)
	) name2764 (
		_w2715_,
		_w2731_,
		_w3226_
	);
	LUT2 #(
		.INIT('h1)
	) name2765 (
		_w3225_,
		_w3226_,
		_w3227_
	);
	LUT2 #(
		.INIT('h1)
	) name2766 (
		_w2742_,
		_w2755_,
		_w3228_
	);
	LUT2 #(
		.INIT('h8)
	) name2767 (
		_w2742_,
		_w2755_,
		_w3229_
	);
	LUT2 #(
		.INIT('h1)
	) name2768 (
		_w2765_,
		_w2779_,
		_w3230_
	);
	LUT2 #(
		.INIT('h4)
	) name2769 (
		_w3229_,
		_w3230_,
		_w3231_
	);
	LUT2 #(
		.INIT('h1)
	) name2770 (
		_w3228_,
		_w3231_,
		_w3232_
	);
	LUT2 #(
		.INIT('h2)
	) name2771 (
		_w3227_,
		_w3232_,
		_w3233_
	);
	LUT2 #(
		.INIT('h1)
	) name2772 (
		_w2715_,
		_w2731_,
		_w3234_
	);
	LUT2 #(
		.INIT('h1)
	) name2773 (
		_w2688_,
		_w2704_,
		_w3235_
	);
	LUT2 #(
		.INIT('h4)
	) name2774 (
		_w3226_,
		_w3235_,
		_w3236_
	);
	LUT2 #(
		.INIT('h1)
	) name2775 (
		_w3234_,
		_w3236_,
		_w3237_
	);
	LUT2 #(
		.INIT('h4)
	) name2776 (
		_w3233_,
		_w3237_,
		_w3238_
	);
	LUT2 #(
		.INIT('h8)
	) name2777 (
		_w2765_,
		_w2779_,
		_w3239_
	);
	LUT2 #(
		.INIT('h1)
	) name2778 (
		_w3229_,
		_w3239_,
		_w3240_
	);
	LUT2 #(
		.INIT('h8)
	) name2779 (
		_w2480_,
		_w2495_,
		_w3241_
	);
	LUT2 #(
		.INIT('h8)
	) name2780 (
		_w2454_,
		_w2470_,
		_w3242_
	);
	LUT2 #(
		.INIT('h1)
	) name2781 (
		_w3241_,
		_w3242_,
		_w3243_
	);
	LUT2 #(
		.INIT('h2)
	) name2782 (
		_w2506_,
		_w2521_,
		_w3244_
	);
	LUT2 #(
		.INIT('h4)
	) name2783 (
		_w2506_,
		_w2521_,
		_w3245_
	);
	LUT2 #(
		.INIT('h4)
	) name2784 (
		_w2531_,
		_w2544_,
		_w3246_
	);
	LUT2 #(
		.INIT('h1)
	) name2785 (
		_w3245_,
		_w3246_,
		_w3247_
	);
	LUT2 #(
		.INIT('h1)
	) name2786 (
		_w3244_,
		_w3247_,
		_w3248_
	);
	LUT2 #(
		.INIT('h8)
	) name2787 (
		_w3243_,
		_w3248_,
		_w3249_
	);
	LUT2 #(
		.INIT('h1)
	) name2788 (
		_w2454_,
		_w2470_,
		_w3250_
	);
	LUT2 #(
		.INIT('h1)
	) name2789 (
		_w2480_,
		_w2495_,
		_w3251_
	);
	LUT2 #(
		.INIT('h4)
	) name2790 (
		_w3242_,
		_w3251_,
		_w3252_
	);
	LUT2 #(
		.INIT('h1)
	) name2791 (
		_w3250_,
		_w3252_,
		_w3253_
	);
	LUT2 #(
		.INIT('h4)
	) name2792 (
		_w2552_,
		_w2566_,
		_w3254_
	);
	LUT2 #(
		.INIT('h4)
	) name2793 (
		_w2574_,
		_w2588_,
		_w3255_
	);
	LUT2 #(
		.INIT('h1)
	) name2794 (
		_w3254_,
		_w3255_,
		_w3256_
	);
	LUT2 #(
		.INIT('h2)
	) name2795 (
		_w2574_,
		_w2588_,
		_w3257_
	);
	LUT2 #(
		.INIT('h2)
	) name2796 (
		_w2597_,
		_w2604_,
		_w3258_
	);
	LUT2 #(
		.INIT('h1)
	) name2797 (
		_w3257_,
		_w3258_,
		_w3259_
	);
	LUT2 #(
		.INIT('h2)
	) name2798 (
		_w3256_,
		_w3259_,
		_w3260_
	);
	LUT2 #(
		.INIT('h2)
	) name2799 (
		_w2552_,
		_w2566_,
		_w3261_
	);
	LUT2 #(
		.INIT('h2)
	) name2800 (
		_w2616_,
		_w2631_,
		_w3262_
	);
	LUT2 #(
		.INIT('h1)
	) name2801 (
		_w3261_,
		_w3262_,
		_w3263_
	);
	LUT2 #(
		.INIT('h2)
	) name2802 (
		_w2642_,
		_w2656_,
		_w3264_
	);
	LUT2 #(
		.INIT('h2)
	) name2803 (
		_w3263_,
		_w3264_,
		_w3265_
	);
	LUT2 #(
		.INIT('h4)
	) name2804 (
		_w3260_,
		_w3265_,
		_w3266_
	);
	LUT2 #(
		.INIT('h4)
	) name2805 (
		_w2642_,
		_w2656_,
		_w3267_
	);
	LUT2 #(
		.INIT('h4)
	) name2806 (
		_w2616_,
		_w2631_,
		_w3268_
	);
	LUT2 #(
		.INIT('h1)
	) name2807 (
		_w3267_,
		_w3268_,
		_w3269_
	);
	LUT2 #(
		.INIT('h1)
	) name2808 (
		_w3264_,
		_w3269_,
		_w3270_
	);
	LUT2 #(
		.INIT('h1)
	) name2809 (
		_w3266_,
		_w3270_,
		_w3271_
	);
	LUT2 #(
		.INIT('h2)
	) name2810 (
		_w2531_,
		_w2544_,
		_w3272_
	);
	LUT2 #(
		.INIT('h1)
	) name2811 (
		_w3244_,
		_w3272_,
		_w3273_
	);
	LUT2 #(
		.INIT('h8)
	) name2812 (
		_w3243_,
		_w3273_,
		_w3274_
	);
	LUT2 #(
		.INIT('h4)
	) name2813 (
		_w3271_,
		_w3274_,
		_w3275_
	);
	LUT2 #(
		.INIT('h4)
	) name2814 (
		_w3249_,
		_w3253_,
		_w3276_
	);
	LUT2 #(
		.INIT('h4)
	) name2815 (
		_w3275_,
		_w3276_,
		_w3277_
	);
	LUT2 #(
		.INIT('h8)
	) name2816 (
		_w3227_,
		_w3240_,
		_w3278_
	);
	LUT2 #(
		.INIT('h4)
	) name2817 (
		_w3277_,
		_w3278_,
		_w3279_
	);
	LUT2 #(
		.INIT('h2)
	) name2818 (
		_w3238_,
		_w3279_,
		_w3280_
	);
	LUT2 #(
		.INIT('h2)
	) name2819 (
		_w3224_,
		_w3280_,
		_w3281_
	);
	LUT2 #(
		.INIT('h1)
	) name2820 (
		_w2860_,
		_w2870_,
		_w3282_
	);
	LUT2 #(
		.INIT('h1)
	) name2821 (
		_w2880_,
		_w2893_,
		_w3283_
	);
	LUT2 #(
		.INIT('h1)
	) name2822 (
		_w3282_,
		_w3283_,
		_w3284_
	);
	LUT2 #(
		.INIT('h1)
	) name2823 (
		_w3220_,
		_w3284_,
		_w3285_
	);
	LUT2 #(
		.INIT('h8)
	) name2824 (
		_w3219_,
		_w3285_,
		_w3286_
	);
	LUT2 #(
		.INIT('h1)
	) name2825 (
		_w2804_,
		_w2818_,
		_w3287_
	);
	LUT2 #(
		.INIT('h1)
	) name2826 (
		_w2828_,
		_w2843_,
		_w3288_
	);
	LUT2 #(
		.INIT('h1)
	) name2827 (
		_w3287_,
		_w3288_,
		_w3289_
	);
	LUT2 #(
		.INIT('h1)
	) name2828 (
		_w3217_,
		_w3289_,
		_w3290_
	);
	LUT2 #(
		.INIT('h1)
	) name2829 (
		_w3286_,
		_w3290_,
		_w3291_
	);
	LUT2 #(
		.INIT('h2)
	) name2830 (
		_w3216_,
		_w3291_,
		_w3292_
	);
	LUT2 #(
		.INIT('h1)
	) name2831 (
		_w2433_,
		_w2442_,
		_w3293_
	);
	LUT2 #(
		.INIT('h1)
	) name2832 (
		_w2379_,
		_w2399_,
		_w3294_
	);
	LUT2 #(
		.INIT('h1)
	) name2833 (
		_w3293_,
		_w3294_,
		_w3295_
	);
	LUT2 #(
		.INIT('h1)
	) name2834 (
		_w3214_,
		_w3295_,
		_w3296_
	);
	LUT2 #(
		.INIT('h8)
	) name2835 (
		_w3212_,
		_w3296_,
		_w3297_
	);
	LUT2 #(
		.INIT('h1)
	) name2836 (
		_w2358_,
		_w2368_,
		_w3298_
	);
	LUT2 #(
		.INIT('h1)
	) name2837 (
		_w2299_,
		_w2311_,
		_w3299_
	);
	LUT2 #(
		.INIT('h1)
	) name2838 (
		_w3298_,
		_w3299_,
		_w3300_
	);
	LUT2 #(
		.INIT('h1)
	) name2839 (
		_w3211_,
		_w3300_,
		_w3301_
	);
	LUT2 #(
		.INIT('h1)
	) name2840 (
		_w3297_,
		_w3301_,
		_w3302_
	);
	LUT2 #(
		.INIT('h4)
	) name2841 (
		_w3292_,
		_w3302_,
		_w3303_
	);
	LUT2 #(
		.INIT('h4)
	) name2842 (
		_w3281_,
		_w3303_,
		_w3304_
	);
	LUT2 #(
		.INIT('h8)
	) name2843 (
		_w3121_,
		_w3130_,
		_w3305_
	);
	LUT2 #(
		.INIT('h1)
	) name2844 (
		_w3189_,
		_w3305_,
		_w3306_
	);
	LUT2 #(
		.INIT('h8)
	) name2845 (
		_w3188_,
		_w3306_,
		_w3307_
	);
	LUT2 #(
		.INIT('h8)
	) name2846 (
		_w3185_,
		_w3307_,
		_w3308_
	);
	LUT2 #(
		.INIT('h4)
	) name2847 (
		_w3304_,
		_w3308_,
		_w3309_
	);
	LUT2 #(
		.INIT('h1)
	) name2848 (
		_w3205_,
		_w3209_,
		_w3310_
	);
	LUT2 #(
		.INIT('h4)
	) name2849 (
		_w3200_,
		_w3310_,
		_w3311_
	);
	LUT2 #(
		.INIT('h4)
	) name2850 (
		_w3309_,
		_w3311_,
		_w3312_
	);
	LUT2 #(
		.INIT('h2)
	) name2851 (
		_w2254_,
		_w3312_,
		_w3313_
	);
	LUT2 #(
		.INIT('h4)
	) name2852 (
		_w2254_,
		_w3312_,
		_w3314_
	);
	LUT2 #(
		.INIT('h1)
	) name2853 (
		_w3313_,
		_w3314_,
		_w3315_
	);
	LUT2 #(
		.INIT('h8)
	) name2854 (
		_w2040_,
		_w3315_,
		_w3316_
	);
	LUT2 #(
		.INIT('h1)
	) name2855 (
		_w2041_,
		_w3316_,
		_w3317_
	);
	LUT2 #(
		.INIT('h2)
	) name2856 (
		_w3172_,
		_w3175_,
		_w3318_
	);
	LUT2 #(
		.INIT('h2)
	) name2857 (
		_w3167_,
		_w3170_,
		_w3319_
	);
	LUT2 #(
		.INIT('h1)
	) name2858 (
		_w3318_,
		_w3319_,
		_w3320_
	);
	LUT2 #(
		.INIT('h1)
	) name2859 (
		_w3317_,
		_w3320_,
		_w3321_
	);
	LUT2 #(
		.INIT('h1)
	) name2860 (
		_w2299_,
		_w2358_,
		_w3322_
	);
	LUT2 #(
		.INIT('h1)
	) name2861 (
		_w3079_,
		_w3121_,
		_w3323_
	);
	LUT2 #(
		.INIT('h4)
	) name2862 (
		_w3102_,
		_w3323_,
		_w3324_
	);
	LUT2 #(
		.INIT('h8)
	) name2863 (
		_w3322_,
		_w3324_,
		_w3325_
	);
	LUT2 #(
		.INIT('h8)
	) name2864 (
		_w2588_,
		_w2604_,
		_w3326_
	);
	LUT2 #(
		.INIT('h8)
	) name2865 (
		_w2566_,
		_w3326_,
		_w3327_
	);
	LUT2 #(
		.INIT('h8)
	) name2866 (
		_w2631_,
		_w3327_,
		_w3328_
	);
	LUT2 #(
		.INIT('h8)
	) name2867 (
		_w2656_,
		_w3328_,
		_w3329_
	);
	LUT2 #(
		.INIT('h8)
	) name2868 (
		_w2544_,
		_w3329_,
		_w3330_
	);
	LUT2 #(
		.INIT('h8)
	) name2869 (
		_w2521_,
		_w3330_,
		_w3331_
	);
	LUT2 #(
		.INIT('h4)
	) name2870 (
		_w2495_,
		_w3331_,
		_w3332_
	);
	LUT2 #(
		.INIT('h1)
	) name2871 (
		_w2470_,
		_w2779_,
		_w3333_
	);
	LUT2 #(
		.INIT('h8)
	) name2872 (
		_w3332_,
		_w3333_,
		_w3334_
	);
	LUT2 #(
		.INIT('h1)
	) name2873 (
		_w2704_,
		_w2755_,
		_w3335_
	);
	LUT2 #(
		.INIT('h8)
	) name2874 (
		_w3334_,
		_w3335_,
		_w3336_
	);
	LUT2 #(
		.INIT('h4)
	) name2875 (
		_w2731_,
		_w3336_,
		_w3337_
	);
	LUT2 #(
		.INIT('h1)
	) name2876 (
		_w2860_,
		_w2893_,
		_w3338_
	);
	LUT2 #(
		.INIT('h8)
	) name2877 (
		_w3337_,
		_w3338_,
		_w3339_
	);
	LUT2 #(
		.INIT('h1)
	) name2878 (
		_w2399_,
		_w2818_,
		_w3340_
	);
	LUT2 #(
		.INIT('h1)
	) name2879 (
		_w2433_,
		_w2843_,
		_w3341_
	);
	LUT2 #(
		.INIT('h8)
	) name2880 (
		_w3340_,
		_w3341_,
		_w3342_
	);
	LUT2 #(
		.INIT('h8)
	) name2881 (
		_w3339_,
		_w3342_,
		_w3343_
	);
	LUT2 #(
		.INIT('h1)
	) name2882 (
		_w3034_,
		_w3054_,
		_w3344_
	);
	LUT2 #(
		.INIT('h8)
	) name2883 (
		_w3325_,
		_w3344_,
		_w3345_
	);
	LUT2 #(
		.INIT('h8)
	) name2884 (
		_w3343_,
		_w3345_,
		_w3346_
	);
	LUT2 #(
		.INIT('h1)
	) name2885 (
		_w2982_,
		_w3012_,
		_w3347_
	);
	LUT2 #(
		.INIT('h4)
	) name2886 (
		_w2949_,
		_w3347_,
		_w3348_
	);
	LUT2 #(
		.INIT('h8)
	) name2887 (
		_w3346_,
		_w3348_,
		_w3349_
	);
	LUT2 #(
		.INIT('h4)
	) name2888 (
		_w2198_,
		_w3349_,
		_w3350_
	);
	LUT2 #(
		.INIT('h2)
	) name2889 (
		_w2198_,
		_w3349_,
		_w3351_
	);
	LUT2 #(
		.INIT('h1)
	) name2890 (
		_w3350_,
		_w3351_,
		_w3352_
	);
	LUT2 #(
		.INIT('h8)
	) name2891 (
		_w3170_,
		_w3175_,
		_w3353_
	);
	LUT2 #(
		.INIT('h4)
	) name2892 (
		_w3166_,
		_w3353_,
		_w3354_
	);
	LUT2 #(
		.INIT('h4)
	) name2893 (
		_w1982_,
		_w3354_,
		_w3355_
	);
	LUT2 #(
		.INIT('h8)
	) name2894 (
		_w3352_,
		_w3355_,
		_w3356_
	);
	LUT2 #(
		.INIT('h1)
	) name2895 (
		_w1982_,
		_w3166_,
		_w3357_
	);
	LUT2 #(
		.INIT('h4)
	) name2896 (
		_w3170_,
		_w3357_,
		_w3358_
	);
	LUT2 #(
		.INIT('h8)
	) name2897 (
		_w2198_,
		_w3358_,
		_w3359_
	);
	LUT2 #(
		.INIT('h2)
	) name2898 (
		_w2058_,
		_w2962_,
		_w3360_
	);
	LUT2 #(
		.INIT('h1)
	) name2899 (
		_w3021_,
		_w3043_,
		_w3361_
	);
	LUT2 #(
		.INIT('h1)
	) name2900 (
		_w3088_,
		_w3112_,
		_w3362_
	);
	LUT2 #(
		.INIT('h4)
	) name2901 (
		_w3065_,
		_w3362_,
		_w3363_
	);
	LUT2 #(
		.INIT('h4)
	) name2902 (
		_w2991_,
		_w3361_,
		_w3364_
	);
	LUT2 #(
		.INIT('h8)
	) name2903 (
		_w3363_,
		_w3364_,
		_w3365_
	);
	LUT2 #(
		.INIT('h4)
	) name2904 (
		_w2962_,
		_w3365_,
		_w3366_
	);
	LUT2 #(
		.INIT('h8)
	) name2905 (
		\P2_reg2_reg[31]/NET0131 ,
		_w2243_,
		_w3367_
	);
	LUT2 #(
		.INIT('h8)
	) name2906 (
		\P2_reg0_reg[31]/NET0131 ,
		_w2245_,
		_w3368_
	);
	LUT2 #(
		.INIT('h8)
	) name2907 (
		\P2_reg1_reg[31]/NET0131 ,
		_w2247_,
		_w3369_
	);
	LUT2 #(
		.INIT('h1)
	) name2908 (
		_w2242_,
		_w3367_,
		_w3370_
	);
	LUT2 #(
		.INIT('h1)
	) name2909 (
		_w3368_,
		_w3369_,
		_w3371_
	);
	LUT2 #(
		.INIT('h8)
	) name2910 (
		_w3370_,
		_w3371_,
		_w3372_
	);
	LUT2 #(
		.INIT('h1)
	) name2911 (
		_w2597_,
		_w3372_,
		_w3373_
	);
	LUT2 #(
		.INIT('h4)
	) name2912 (
		_w2574_,
		_w3373_,
		_w3374_
	);
	LUT2 #(
		.INIT('h4)
	) name2913 (
		_w2552_,
		_w3374_,
		_w3375_
	);
	LUT2 #(
		.INIT('h4)
	) name2914 (
		_w2616_,
		_w3375_,
		_w3376_
	);
	LUT2 #(
		.INIT('h1)
	) name2915 (
		_w2531_,
		_w2642_,
		_w3377_
	);
	LUT2 #(
		.INIT('h8)
	) name2916 (
		_w3376_,
		_w3377_,
		_w3378_
	);
	LUT2 #(
		.INIT('h4)
	) name2917 (
		_w2506_,
		_w3378_,
		_w3379_
	);
	LUT2 #(
		.INIT('h4)
	) name2918 (
		_w2480_,
		_w3379_,
		_w3380_
	);
	LUT2 #(
		.INIT('h1)
	) name2919 (
		_w2454_,
		_w2742_,
		_w3381_
	);
	LUT2 #(
		.INIT('h4)
	) name2920 (
		_w2765_,
		_w3381_,
		_w3382_
	);
	LUT2 #(
		.INIT('h8)
	) name2921 (
		_w3380_,
		_w3382_,
		_w3383_
	);
	LUT2 #(
		.INIT('h1)
	) name2922 (
		_w2688_,
		_w2715_,
		_w3384_
	);
	LUT2 #(
		.INIT('h4)
	) name2923 (
		_w2880_,
		_w3384_,
		_w3385_
	);
	LUT2 #(
		.INIT('h4)
	) name2924 (
		_w2870_,
		_w3385_,
		_w3386_
	);
	LUT2 #(
		.INIT('h8)
	) name2925 (
		_w3383_,
		_w3386_,
		_w3387_
	);
	LUT2 #(
		.INIT('h1)
	) name2926 (
		_w2379_,
		_w2804_,
		_w3388_
	);
	LUT2 #(
		.INIT('h4)
	) name2927 (
		_w2828_,
		_w3388_,
		_w3389_
	);
	LUT2 #(
		.INIT('h4)
	) name2928 (
		_w2442_,
		_w3389_,
		_w3390_
	);
	LUT2 #(
		.INIT('h1)
	) name2929 (
		_w2311_,
		_w2368_,
		_w3391_
	);
	LUT2 #(
		.INIT('h4)
	) name2930 (
		_w3130_,
		_w3391_,
		_w3392_
	);
	LUT2 #(
		.INIT('h8)
	) name2931 (
		_w3390_,
		_w3392_,
		_w3393_
	);
	LUT2 #(
		.INIT('h8)
	) name2932 (
		_w3387_,
		_w3393_,
		_w3394_
	);
	LUT2 #(
		.INIT('h4)
	) name2933 (
		_w2251_,
		_w3366_,
		_w3395_
	);
	LUT2 #(
		.INIT('h8)
	) name2934 (
		_w3394_,
		_w3395_,
		_w3396_
	);
	LUT2 #(
		.INIT('h8)
	) name2935 (
		\P2_reg2_reg[30]/NET0131 ,
		_w2243_,
		_w3397_
	);
	LUT2 #(
		.INIT('h8)
	) name2936 (
		\P2_reg0_reg[30]/NET0131 ,
		_w2245_,
		_w3398_
	);
	LUT2 #(
		.INIT('h8)
	) name2937 (
		\P2_reg1_reg[30]/NET0131 ,
		_w2247_,
		_w3399_
	);
	LUT2 #(
		.INIT('h1)
	) name2938 (
		_w2242_,
		_w3397_,
		_w3400_
	);
	LUT2 #(
		.INIT('h1)
	) name2939 (
		_w3398_,
		_w3399_,
		_w3401_
	);
	LUT2 #(
		.INIT('h8)
	) name2940 (
		_w3400_,
		_w3401_,
		_w3402_
	);
	LUT2 #(
		.INIT('h4)
	) name2941 (
		_w3396_,
		_w3402_,
		_w3403_
	);
	LUT2 #(
		.INIT('h2)
	) name2942 (
		_w3396_,
		_w3402_,
		_w3404_
	);
	LUT2 #(
		.INIT('h8)
	) name2943 (
		\P2_B_reg/NET0131 ,
		_w2051_,
		_w3405_
	);
	LUT2 #(
		.INIT('h1)
	) name2944 (
		_w2058_,
		_w3405_,
		_w3406_
	);
	LUT2 #(
		.INIT('h4)
	) name2945 (
		_w3404_,
		_w3406_,
		_w3407_
	);
	LUT2 #(
		.INIT('h4)
	) name2946 (
		_w3403_,
		_w3407_,
		_w3408_
	);
	LUT2 #(
		.INIT('h1)
	) name2947 (
		_w3360_,
		_w3408_,
		_w3409_
	);
	LUT2 #(
		.INIT('h8)
	) name2948 (
		_w1982_,
		_w3166_,
		_w3410_
	);
	LUT2 #(
		.INIT('h8)
	) name2949 (
		_w3353_,
		_w3410_,
		_w3411_
	);
	LUT2 #(
		.INIT('h4)
	) name2950 (
		_w3409_,
		_w3411_,
		_w3412_
	);
	LUT2 #(
		.INIT('h1)
	) name2951 (
		_w3359_,
		_w3412_,
		_w3413_
	);
	LUT2 #(
		.INIT('h4)
	) name2952 (
		_w3356_,
		_w3413_,
		_w3414_
	);
	LUT2 #(
		.INIT('h2)
	) name2953 (
		_w2040_,
		_w3414_,
		_w3415_
	);
	LUT2 #(
		.INIT('h4)
	) name2954 (
		_w2040_,
		_w3411_,
		_w3416_
	);
	LUT2 #(
		.INIT('h4)
	) name2955 (
		_w3353_,
		_w3410_,
		_w3417_
	);
	LUT2 #(
		.INIT('h2)
	) name2956 (
		_w3170_,
		_w3175_,
		_w3418_
	);
	LUT2 #(
		.INIT('h4)
	) name2957 (
		_w3166_,
		_w3418_,
		_w3419_
	);
	LUT2 #(
		.INIT('h4)
	) name2958 (
		_w1982_,
		_w3419_,
		_w3420_
	);
	LUT2 #(
		.INIT('h1)
	) name2959 (
		_w3417_,
		_w3420_,
		_w3421_
	);
	LUT2 #(
		.INIT('h4)
	) name2960 (
		_w2040_,
		_w3358_,
		_w3422_
	);
	LUT2 #(
		.INIT('h2)
	) name2961 (
		_w3421_,
		_w3422_,
		_w3423_
	);
	LUT2 #(
		.INIT('h4)
	) name2962 (
		_w2040_,
		_w3355_,
		_w3424_
	);
	LUT2 #(
		.INIT('h2)
	) name2963 (
		_w3423_,
		_w3424_,
		_w3425_
	);
	LUT2 #(
		.INIT('h4)
	) name2964 (
		_w3416_,
		_w3425_,
		_w3426_
	);
	LUT2 #(
		.INIT('h2)
	) name2965 (
		\P2_reg0_reg[29]/NET0131 ,
		_w3426_,
		_w3427_
	);
	LUT2 #(
		.INIT('h1)
	) name2966 (
		_w3415_,
		_w3427_,
		_w3428_
	);
	LUT2 #(
		.INIT('h4)
	) name2967 (
		_w3321_,
		_w3428_,
		_w3429_
	);
	LUT2 #(
		.INIT('h4)
	) name2968 (
		_w3178_,
		_w3429_,
		_w3430_
	);
	LUT2 #(
		.INIT('h2)
	) name2969 (
		_w2026_,
		_w3430_,
		_w3431_
	);
	LUT2 #(
		.INIT('h1)
	) name2970 (
		_w2025_,
		_w3431_,
		_w3432_
	);
	LUT2 #(
		.INIT('h2)
	) name2971 (
		\P1_state_reg[0]/NET0131 ,
		_w3432_,
		_w3433_
	);
	LUT2 #(
		.INIT('h1)
	) name2972 (
		_w1984_,
		_w3433_,
		_w3434_
	);
	LUT2 #(
		.INIT('h8)
	) name2973 (
		\P1_state_reg[0]/NET0131 ,
		_w512_,
		_w3435_
	);
	LUT2 #(
		.INIT('h2)
	) name2974 (
		\P1_reg2_reg[29]/NET0131 ,
		_w3435_,
		_w3436_
	);
	LUT2 #(
		.INIT('h2)
	) name2975 (
		\P1_IR_reg[25]/NET0131 ,
		_w708_,
		_w3437_
	);
	LUT2 #(
		.INIT('h4)
	) name2976 (
		\P1_IR_reg[25]/NET0131 ,
		_w708_,
		_w3438_
	);
	LUT2 #(
		.INIT('h1)
	) name2977 (
		_w3437_,
		_w3438_,
		_w3439_
	);
	LUT2 #(
		.INIT('h2)
	) name2978 (
		\P1_IR_reg[26]/NET0131 ,
		_w696_,
		_w3440_
	);
	LUT2 #(
		.INIT('h4)
	) name2979 (
		\P1_IR_reg[26]/NET0131 ,
		_w696_,
		_w3441_
	);
	LUT2 #(
		.INIT('h1)
	) name2980 (
		_w3440_,
		_w3441_,
		_w3442_
	);
	LUT2 #(
		.INIT('h1)
	) name2981 (
		\P1_IR_reg[24]/NET0131 ,
		_w530_,
		_w3443_
	);
	LUT2 #(
		.INIT('h8)
	) name2982 (
		\P1_IR_reg[24]/NET0131 ,
		_w530_,
		_w3444_
	);
	LUT2 #(
		.INIT('h1)
	) name2983 (
		_w3443_,
		_w3444_,
		_w3445_
	);
	LUT2 #(
		.INIT('h1)
	) name2984 (
		_w3439_,
		_w3442_,
		_w3446_
	);
	LUT2 #(
		.INIT('h8)
	) name2985 (
		_w3445_,
		_w3446_,
		_w3447_
	);
	LUT2 #(
		.INIT('h8)
	) name2986 (
		_w512_,
		_w3447_,
		_w3448_
	);
	LUT2 #(
		.INIT('h8)
	) name2987 (
		\P1_reg2_reg[29]/NET0131 ,
		_w3448_,
		_w3449_
	);
	LUT2 #(
		.INIT('h2)
	) name2988 (
		_w512_,
		_w3447_,
		_w3450_
	);
	LUT2 #(
		.INIT('h2)
	) name2989 (
		_w3439_,
		_w3442_,
		_w3451_
	);
	LUT2 #(
		.INIT('h4)
	) name2990 (
		\P1_B_reg/NET0131 ,
		_w3445_,
		_w3452_
	);
	LUT2 #(
		.INIT('h8)
	) name2991 (
		_w3451_,
		_w3452_,
		_w3453_
	);
	LUT2 #(
		.INIT('h1)
	) name2992 (
		\P1_d_reg[0]/NET0131 ,
		_w3453_,
		_w3454_
	);
	LUT2 #(
		.INIT('h1)
	) name2993 (
		_w3442_,
		_w3454_,
		_w3455_
	);
	LUT2 #(
		.INIT('h2)
	) name2994 (
		\P1_B_reg/NET0131 ,
		_w3445_,
		_w3456_
	);
	LUT2 #(
		.INIT('h8)
	) name2995 (
		_w3451_,
		_w3456_,
		_w3457_
	);
	LUT2 #(
		.INIT('h8)
	) name2996 (
		_w3442_,
		_w3445_,
		_w3458_
	);
	LUT2 #(
		.INIT('h1)
	) name2997 (
		_w3457_,
		_w3458_,
		_w3459_
	);
	LUT2 #(
		.INIT('h4)
	) name2998 (
		_w3455_,
		_w3459_,
		_w3460_
	);
	LUT2 #(
		.INIT('h2)
	) name2999 (
		\P1_d_reg[1]/NET0131 ,
		_w3442_,
		_w3461_
	);
	LUT2 #(
		.INIT('h4)
	) name3000 (
		_w3439_,
		_w3442_,
		_w3462_
	);
	LUT2 #(
		.INIT('h1)
	) name3001 (
		_w3461_,
		_w3462_,
		_w3463_
	);
	LUT2 #(
		.INIT('h4)
	) name3002 (
		_w3453_,
		_w3463_,
		_w3464_
	);
	LUT2 #(
		.INIT('h4)
	) name3003 (
		_w3457_,
		_w3464_,
		_w3465_
	);
	LUT2 #(
		.INIT('h2)
	) name3004 (
		_w3460_,
		_w3465_,
		_w3466_
	);
	LUT2 #(
		.INIT('h2)
	) name3005 (
		\P1_reg2_reg[29]/NET0131 ,
		_w3466_,
		_w3467_
	);
	LUT2 #(
		.INIT('h1)
	) name3006 (
		_w1816_,
		_w1820_,
		_w3468_
	);
	LUT2 #(
		.INIT('h4)
	) name3007 (
		_w1836_,
		_w1840_,
		_w3469_
	);
	LUT2 #(
		.INIT('h1)
	) name3008 (
		_w1837_,
		_w3469_,
		_w3470_
	);
	LUT2 #(
		.INIT('h2)
	) name3009 (
		_w3468_,
		_w3470_,
		_w3471_
	);
	LUT2 #(
		.INIT('h4)
	) name3010 (
		_w1816_,
		_w1819_,
		_w3472_
	);
	LUT2 #(
		.INIT('h1)
	) name3011 (
		_w1817_,
		_w3472_,
		_w3473_
	);
	LUT2 #(
		.INIT('h4)
	) name3012 (
		_w3471_,
		_w3473_,
		_w3474_
	);
	LUT2 #(
		.INIT('h1)
	) name3013 (
		_w1767_,
		_w1808_,
		_w3475_
	);
	LUT2 #(
		.INIT('h4)
	) name3014 (
		_w1810_,
		_w3475_,
		_w3476_
	);
	LUT2 #(
		.INIT('h4)
	) name3015 (
		_w3474_,
		_w3476_,
		_w3477_
	);
	LUT2 #(
		.INIT('h1)
	) name3016 (
		_w1807_,
		_w1811_,
		_w3478_
	);
	LUT2 #(
		.INIT('h2)
	) name3017 (
		_w3475_,
		_w3478_,
		_w3479_
	);
	LUT2 #(
		.INIT('h1)
	) name3018 (
		_w1768_,
		_w3479_,
		_w3480_
	);
	LUT2 #(
		.INIT('h4)
	) name3019 (
		_w1830_,
		_w3480_,
		_w3481_
	);
	LUT2 #(
		.INIT('h4)
	) name3020 (
		_w3477_,
		_w3481_,
		_w3482_
	);
	LUT2 #(
		.INIT('h1)
	) name3021 (
		_w1829_,
		_w3482_,
		_w3483_
	);
	LUT2 #(
		.INIT('h1)
	) name3022 (
		_w1826_,
		_w1833_,
		_w3484_
	);
	LUT2 #(
		.INIT('h4)
	) name3023 (
		_w1443_,
		_w1452_,
		_w3485_
	);
	LUT2 #(
		.INIT('h1)
	) name3024 (
		_w1822_,
		_w3485_,
		_w3486_
	);
	LUT2 #(
		.INIT('h8)
	) name3025 (
		_w3484_,
		_w3486_,
		_w3487_
	);
	LUT2 #(
		.INIT('h1)
	) name3026 (
		_w1797_,
		_w1813_,
		_w3488_
	);
	LUT2 #(
		.INIT('h1)
	) name3027 (
		_w1783_,
		_w1786_,
		_w3489_
	);
	LUT2 #(
		.INIT('h8)
	) name3028 (
		_w3488_,
		_w3489_,
		_w3490_
	);
	LUT2 #(
		.INIT('h8)
	) name3029 (
		_w3487_,
		_w3490_,
		_w3491_
	);
	LUT2 #(
		.INIT('h1)
	) name3030 (
		_w1770_,
		_w1794_,
		_w3492_
	);
	LUT2 #(
		.INIT('h2)
	) name3031 (
		_w1780_,
		_w1790_,
		_w3493_
	);
	LUT2 #(
		.INIT('h1)
	) name3032 (
		_w1789_,
		_w3493_,
		_w3494_
	);
	LUT2 #(
		.INIT('h2)
	) name3033 (
		_w3492_,
		_w3494_,
		_w3495_
	);
	LUT2 #(
		.INIT('h2)
	) name3034 (
		_w1771_,
		_w1794_,
		_w3496_
	);
	LUT2 #(
		.INIT('h1)
	) name3035 (
		_w1795_,
		_w3496_,
		_w3497_
	);
	LUT2 #(
		.INIT('h4)
	) name3036 (
		_w3495_,
		_w3497_,
		_w3498_
	);
	LUT2 #(
		.INIT('h8)
	) name3037 (
		_w1524_,
		_w1537_,
		_w3499_
	);
	LUT2 #(
		.INIT('h8)
	) name3038 (
		_w1548_,
		_w1562_,
		_w3500_
	);
	LUT2 #(
		.INIT('h1)
	) name3039 (
		_w3499_,
		_w3500_,
		_w3501_
	);
	LUT2 #(
		.INIT('h1)
	) name3040 (
		_w1774_,
		_w1800_,
		_w3502_
	);
	LUT2 #(
		.INIT('h8)
	) name3041 (
		_w1641_,
		_w1655_,
		_w3503_
	);
	LUT2 #(
		.INIT('h1)
	) name3042 (
		_w1641_,
		_w1655_,
		_w3504_
	);
	LUT2 #(
		.INIT('h1)
	) name3043 (
		_w1664_,
		_w1671_,
		_w3505_
	);
	LUT2 #(
		.INIT('h1)
	) name3044 (
		_w3504_,
		_w3505_,
		_w3506_
	);
	LUT2 #(
		.INIT('h1)
	) name3045 (
		_w3503_,
		_w3506_,
		_w3507_
	);
	LUT2 #(
		.INIT('h1)
	) name3046 (
		_w1777_,
		_w3507_,
		_w3508_
	);
	LUT2 #(
		.INIT('h8)
	) name3047 (
		_w1617_,
		_w1632_,
		_w3509_
	);
	LUT2 #(
		.INIT('h1)
	) name3048 (
		_w1778_,
		_w3509_,
		_w3510_
	);
	LUT2 #(
		.INIT('h8)
	) name3049 (
		_w1572_,
		_w1586_,
		_w3511_
	);
	LUT2 #(
		.INIT('h2)
	) name3050 (
		_w3510_,
		_w3511_,
		_w3512_
	);
	LUT2 #(
		.INIT('h4)
	) name3051 (
		_w3508_,
		_w3512_,
		_w3513_
	);
	LUT2 #(
		.INIT('h1)
	) name3052 (
		_w1572_,
		_w1586_,
		_w3514_
	);
	LUT2 #(
		.INIT('h1)
	) name3053 (
		_w1617_,
		_w1632_,
		_w3515_
	);
	LUT2 #(
		.INIT('h4)
	) name3054 (
		_w3511_,
		_w3515_,
		_w3516_
	);
	LUT2 #(
		.INIT('h1)
	) name3055 (
		_w3514_,
		_w3516_,
		_w3517_
	);
	LUT2 #(
		.INIT('h4)
	) name3056 (
		_w3513_,
		_w3517_,
		_w3518_
	);
	LUT2 #(
		.INIT('h8)
	) name3057 (
		_w3501_,
		_w3502_,
		_w3519_
	);
	LUT2 #(
		.INIT('h4)
	) name3058 (
		_w3518_,
		_w3519_,
		_w3520_
	);
	LUT2 #(
		.INIT('h1)
	) name3059 (
		_w1524_,
		_w1537_,
		_w3521_
	);
	LUT2 #(
		.INIT('h1)
	) name3060 (
		_w1548_,
		_w1562_,
		_w3522_
	);
	LUT2 #(
		.INIT('h4)
	) name3061 (
		_w3499_,
		_w3522_,
		_w3523_
	);
	LUT2 #(
		.INIT('h1)
	) name3062 (
		_w3521_,
		_w3523_,
		_w3524_
	);
	LUT2 #(
		.INIT('h2)
	) name3063 (
		_w3502_,
		_w3524_,
		_w3525_
	);
	LUT2 #(
		.INIT('h2)
	) name3064 (
		_w1775_,
		_w1800_,
		_w3526_
	);
	LUT2 #(
		.INIT('h1)
	) name3065 (
		_w1801_,
		_w3526_,
		_w3527_
	);
	LUT2 #(
		.INIT('h4)
	) name3066 (
		_w3525_,
		_w3527_,
		_w3528_
	);
	LUT2 #(
		.INIT('h4)
	) name3067 (
		_w3520_,
		_w3528_,
		_w3529_
	);
	LUT2 #(
		.INIT('h1)
	) name3068 (
		_w1781_,
		_w1790_,
		_w3530_
	);
	LUT2 #(
		.INIT('h8)
	) name3069 (
		_w3492_,
		_w3530_,
		_w3531_
	);
	LUT2 #(
		.INIT('h4)
	) name3070 (
		_w3529_,
		_w3531_,
		_w3532_
	);
	LUT2 #(
		.INIT('h2)
	) name3071 (
		_w3498_,
		_w3532_,
		_w3533_
	);
	LUT2 #(
		.INIT('h2)
	) name3072 (
		_w3491_,
		_w3533_,
		_w3534_
	);
	LUT2 #(
		.INIT('h2)
	) name3073 (
		_w1798_,
		_w1813_,
		_w3535_
	);
	LUT2 #(
		.INIT('h1)
	) name3074 (
		_w1814_,
		_w3535_,
		_w3536_
	);
	LUT2 #(
		.INIT('h2)
	) name3075 (
		_w3489_,
		_w3536_,
		_w3537_
	);
	LUT2 #(
		.INIT('h1)
	) name3076 (
		_w1784_,
		_w1787_,
		_w3538_
	);
	LUT2 #(
		.INIT('h1)
	) name3077 (
		_w1783_,
		_w3538_,
		_w3539_
	);
	LUT2 #(
		.INIT('h1)
	) name3078 (
		_w3537_,
		_w3539_,
		_w3540_
	);
	LUT2 #(
		.INIT('h2)
	) name3079 (
		_w3487_,
		_w3540_,
		_w3541_
	);
	LUT2 #(
		.INIT('h2)
	) name3080 (
		_w1443_,
		_w1452_,
		_w3542_
	);
	LUT2 #(
		.INIT('h4)
	) name3081 (
		_w1822_,
		_w3542_,
		_w3543_
	);
	LUT2 #(
		.INIT('h1)
	) name3082 (
		_w1823_,
		_w3543_,
		_w3544_
	);
	LUT2 #(
		.INIT('h2)
	) name3083 (
		_w3484_,
		_w3544_,
		_w3545_
	);
	LUT2 #(
		.INIT('h4)
	) name3084 (
		_w1826_,
		_w1834_,
		_w3546_
	);
	LUT2 #(
		.INIT('h1)
	) name3085 (
		_w1827_,
		_w3546_,
		_w3547_
	);
	LUT2 #(
		.INIT('h4)
	) name3086 (
		_w3545_,
		_w3547_,
		_w3548_
	);
	LUT2 #(
		.INIT('h4)
	) name3087 (
		_w3541_,
		_w3548_,
		_w3549_
	);
	LUT2 #(
		.INIT('h4)
	) name3088 (
		_w3534_,
		_w3549_,
		_w3550_
	);
	LUT2 #(
		.INIT('h1)
	) name3089 (
		_w1836_,
		_w1839_,
		_w3551_
	);
	LUT2 #(
		.INIT('h8)
	) name3090 (
		_w3468_,
		_w3551_,
		_w3552_
	);
	LUT2 #(
		.INIT('h4)
	) name3091 (
		_w1829_,
		_w3476_,
		_w3553_
	);
	LUT2 #(
		.INIT('h8)
	) name3092 (
		_w3552_,
		_w3553_,
		_w3554_
	);
	LUT2 #(
		.INIT('h4)
	) name3093 (
		_w3550_,
		_w3554_,
		_w3555_
	);
	LUT2 #(
		.INIT('h1)
	) name3094 (
		_w3483_,
		_w3555_,
		_w3556_
	);
	LUT2 #(
		.INIT('h2)
	) name3095 (
		_w1832_,
		_w3556_,
		_w3557_
	);
	LUT2 #(
		.INIT('h4)
	) name3096 (
		_w1832_,
		_w3556_,
		_w3558_
	);
	LUT2 #(
		.INIT('h1)
	) name3097 (
		_w3557_,
		_w3558_,
		_w3559_
	);
	LUT2 #(
		.INIT('h2)
	) name3098 (
		_w3466_,
		_w3559_,
		_w3560_
	);
	LUT2 #(
		.INIT('h1)
	) name3099 (
		_w3467_,
		_w3560_,
		_w3561_
	);
	LUT2 #(
		.INIT('h4)
	) name3100 (
		_w501_,
		_w1888_,
		_w3562_
	);
	LUT2 #(
		.INIT('h1)
	) name3101 (
		_w1766_,
		_w3562_,
		_w3563_
	);
	LUT2 #(
		.INIT('h1)
	) name3102 (
		_w3561_,
		_w3563_,
		_w3564_
	);
	LUT2 #(
		.INIT('h2)
	) name3103 (
		_w537_,
		_w945_,
		_w3565_
	);
	LUT2 #(
		.INIT('h1)
	) name3104 (
		\P1_B_reg/NET0131 ,
		_w537_,
		_w3566_
	);
	LUT2 #(
		.INIT('h1)
	) name3105 (
		_w538_,
		_w3566_,
		_w3567_
	);
	LUT2 #(
		.INIT('h1)
	) name3106 (
		_w1452_,
		_w1475_,
		_w3568_
	);
	LUT2 #(
		.INIT('h1)
	) name3107 (
		_w1094_,
		_w1118_,
		_w3569_
	);
	LUT2 #(
		.INIT('h1)
	) name3108 (
		_w750_,
		_w1664_,
		_w3570_
	);
	LUT2 #(
		.INIT('h4)
	) name3109 (
		_w1641_,
		_w3570_,
		_w3571_
	);
	LUT2 #(
		.INIT('h4)
	) name3110 (
		_w1595_,
		_w3571_,
		_w3572_
	);
	LUT2 #(
		.INIT('h4)
	) name3111 (
		_w1617_,
		_w3572_,
		_w3573_
	);
	LUT2 #(
		.INIT('h1)
	) name3112 (
		_w1548_,
		_w1572_,
		_w3574_
	);
	LUT2 #(
		.INIT('h8)
	) name3113 (
		_w3573_,
		_w3574_,
		_w3575_
	);
	LUT2 #(
		.INIT('h1)
	) name3114 (
		_w1498_,
		_w1524_,
		_w3576_
	);
	LUT2 #(
		.INIT('h8)
	) name3115 (
		_w3575_,
		_w3576_,
		_w3577_
	);
	LUT2 #(
		.INIT('h1)
	) name3116 (
		_w1218_,
		_w1244_,
		_w3578_
	);
	LUT2 #(
		.INIT('h4)
	) name3117 (
		_w1267_,
		_w3578_,
		_w3579_
	);
	LUT2 #(
		.INIT('h8)
	) name3118 (
		_w3577_,
		_w3579_,
		_w3580_
	);
	LUT2 #(
		.INIT('h1)
	) name3119 (
		_w1146_,
		_w1174_,
		_w3581_
	);
	LUT2 #(
		.INIT('h4)
	) name3120 (
		_w1207_,
		_w3581_,
		_w3582_
	);
	LUT2 #(
		.INIT('h8)
	) name3121 (
		_w3580_,
		_w3582_,
		_w3583_
	);
	LUT2 #(
		.INIT('h8)
	) name3122 (
		_w3568_,
		_w3569_,
		_w3584_
	);
	LUT2 #(
		.INIT('h8)
	) name3123 (
		_w3583_,
		_w3584_,
		_w3585_
	);
	LUT2 #(
		.INIT('h1)
	) name3124 (
		_w1318_,
		_w1336_,
		_w3586_
	);
	LUT2 #(
		.INIT('h1)
	) name3125 (
		_w1374_,
		_w1427_,
		_w3587_
	);
	LUT2 #(
		.INIT('h1)
	) name3126 (
		_w1356_,
		_w1403_,
		_w3588_
	);
	LUT2 #(
		.INIT('h8)
	) name3127 (
		_w3587_,
		_w3588_,
		_w3589_
	);
	LUT2 #(
		.INIT('h8)
	) name3128 (
		_w3586_,
		_w3589_,
		_w3590_
	);
	LUT2 #(
		.INIT('h4)
	) name3129 (
		_w1062_,
		_w3590_,
		_w3591_
	);
	LUT2 #(
		.INIT('h4)
	) name3130 (
		_w1038_,
		_w3591_,
		_w3592_
	);
	LUT2 #(
		.INIT('h8)
	) name3131 (
		_w3585_,
		_w3592_,
		_w3593_
	);
	LUT2 #(
		.INIT('h4)
	) name3132 (
		_w1006_,
		_w3593_,
		_w3594_
	);
	LUT2 #(
		.INIT('h1)
	) name3133 (
		_w945_,
		_w978_,
		_w3595_
	);
	LUT2 #(
		.INIT('h4)
	) name3134 (
		_w887_,
		_w3595_,
		_w3596_
	);
	LUT2 #(
		.INIT('h8)
	) name3135 (
		_w3594_,
		_w3596_,
		_w3597_
	);
	LUT2 #(
		.INIT('h2)
	) name3136 (
		_w831_,
		_w3597_,
		_w3598_
	);
	LUT2 #(
		.INIT('h4)
	) name3137 (
		_w831_,
		_w3597_,
		_w3599_
	);
	LUT2 #(
		.INIT('h1)
	) name3138 (
		_w3567_,
		_w3598_,
		_w3600_
	);
	LUT2 #(
		.INIT('h4)
	) name3139 (
		_w3599_,
		_w3600_,
		_w3601_
	);
	LUT2 #(
		.INIT('h1)
	) name3140 (
		_w3565_,
		_w3601_,
		_w3602_
	);
	LUT2 #(
		.INIT('h2)
	) name3141 (
		_w3466_,
		_w3602_,
		_w3603_
	);
	LUT2 #(
		.INIT('h1)
	) name3142 (
		_w3467_,
		_w3603_,
		_w3604_
	);
	LUT2 #(
		.INIT('h2)
	) name3143 (
		_w1936_,
		_w3604_,
		_w3605_
	);
	LUT2 #(
		.INIT('h1)
	) name3144 (
		_w1299_,
		_w1337_,
		_w3606_
	);
	LUT2 #(
		.INIT('h1)
	) name3145 (
		_w1319_,
		_w1700_,
		_w3607_
	);
	LUT2 #(
		.INIT('h8)
	) name3146 (
		_w3606_,
		_w3607_,
		_w3608_
	);
	LUT2 #(
		.INIT('h1)
	) name3147 (
		_w1063_,
		_w1697_,
		_w3609_
	);
	LUT2 #(
		.INIT('h1)
	) name3148 (
		_w1299_,
		_w3609_,
		_w3610_
	);
	LUT2 #(
		.INIT('h1)
	) name3149 (
		_w3608_,
		_w3610_,
		_w3611_
	);
	LUT2 #(
		.INIT('h1)
	) name3150 (
		_w1010_,
		_w1039_,
		_w3612_
	);
	LUT2 #(
		.INIT('h4)
	) name3151 (
		_w979_,
		_w3612_,
		_w3613_
	);
	LUT2 #(
		.INIT('h4)
	) name3152 (
		_w3611_,
		_w3613_,
		_w3614_
	);
	LUT2 #(
		.INIT('h1)
	) name3153 (
		_w1010_,
		_w1889_,
		_w3615_
	);
	LUT2 #(
		.INIT('h4)
	) name3154 (
		_w979_,
		_w3615_,
		_w3616_
	);
	LUT2 #(
		.INIT('h2)
	) name3155 (
		_w1892_,
		_w3616_,
		_w3617_
	);
	LUT2 #(
		.INIT('h4)
	) name3156 (
		_w3614_,
		_w3617_,
		_w3618_
	);
	LUT2 #(
		.INIT('h1)
	) name3157 (
		_w950_,
		_w3618_,
		_w3619_
	);
	LUT2 #(
		.INIT('h1)
	) name3158 (
		_w1375_,
		_w1428_,
		_w3620_
	);
	LUT2 #(
		.INIT('h1)
	) name3159 (
		_w1404_,
		_w1453_,
		_w3621_
	);
	LUT2 #(
		.INIT('h8)
	) name3160 (
		_w3620_,
		_w3621_,
		_w3622_
	);
	LUT2 #(
		.INIT('h1)
	) name3161 (
		_w1095_,
		_w1476_,
		_w3623_
	);
	LUT2 #(
		.INIT('h1)
	) name3162 (
		_w1119_,
		_w1147_,
		_w3624_
	);
	LUT2 #(
		.INIT('h8)
	) name3163 (
		_w3623_,
		_w3624_,
		_w3625_
	);
	LUT2 #(
		.INIT('h8)
	) name3164 (
		_w3622_,
		_w3625_,
		_w3626_
	);
	LUT2 #(
		.INIT('h1)
	) name3165 (
		_w1209_,
		_w1290_,
		_w3627_
	);
	LUT2 #(
		.INIT('h1)
	) name3166 (
		_w1234_,
		_w1286_,
		_w3628_
	);
	LUT2 #(
		.INIT('h8)
	) name3167 (
		_w3627_,
		_w3628_,
		_w3629_
	);
	LUT2 #(
		.INIT('h1)
	) name3168 (
		_w1175_,
		_w1208_,
		_w3630_
	);
	LUT2 #(
		.INIT('h1)
	) name3169 (
		_w1290_,
		_w3630_,
		_w3631_
	);
	LUT2 #(
		.INIT('h1)
	) name3170 (
		_w3629_,
		_w3631_,
		_w3632_
	);
	LUT2 #(
		.INIT('h4)
	) name3171 (
		_w1673_,
		_w1899_,
		_w3633_
	);
	LUT2 #(
		.INIT('h2)
	) name3172 (
		_w1634_,
		_w3633_,
		_w3634_
	);
	LUT2 #(
		.INIT('h2)
	) name3173 (
		_w1897_,
		_w3634_,
		_w3635_
	);
	LUT2 #(
		.INIT('h1)
	) name3174 (
		_w1587_,
		_w3635_,
		_w3636_
	);
	LUT2 #(
		.INIT('h1)
	) name3175 (
		_w1538_,
		_w1563_,
		_w3637_
	);
	LUT2 #(
		.INIT('h1)
	) name3176 (
		_w1282_,
		_w1515_,
		_w3638_
	);
	LUT2 #(
		.INIT('h8)
	) name3177 (
		_w3637_,
		_w3638_,
		_w3639_
	);
	LUT2 #(
		.INIT('h8)
	) name3178 (
		_w3636_,
		_w3639_,
		_w3640_
	);
	LUT2 #(
		.INIT('h1)
	) name3179 (
		_w1538_,
		_w1896_,
		_w3641_
	);
	LUT2 #(
		.INIT('h8)
	) name3180 (
		_w3638_,
		_w3641_,
		_w3642_
	);
	LUT2 #(
		.INIT('h1)
	) name3181 (
		_w1481_,
		_w1688_,
		_w3643_
	);
	LUT2 #(
		.INIT('h1)
	) name3182 (
		_w1282_,
		_w3643_,
		_w3644_
	);
	LUT2 #(
		.INIT('h1)
	) name3183 (
		_w3642_,
		_w3644_,
		_w3645_
	);
	LUT2 #(
		.INIT('h4)
	) name3184 (
		_w3640_,
		_w3645_,
		_w3646_
	);
	LUT2 #(
		.INIT('h1)
	) name3185 (
		_w1234_,
		_w1258_,
		_w3647_
	);
	LUT2 #(
		.INIT('h8)
	) name3186 (
		_w3627_,
		_w3647_,
		_w3648_
	);
	LUT2 #(
		.INIT('h4)
	) name3187 (
		_w3646_,
		_w3648_,
		_w3649_
	);
	LUT2 #(
		.INIT('h2)
	) name3188 (
		_w3632_,
		_w3649_,
		_w3650_
	);
	LUT2 #(
		.INIT('h2)
	) name3189 (
		_w3626_,
		_w3650_,
		_w3651_
	);
	LUT2 #(
		.INIT('h1)
	) name3190 (
		_w1119_,
		_w1292_,
		_w3652_
	);
	LUT2 #(
		.INIT('h8)
	) name3191 (
		_w3623_,
		_w3652_,
		_w3653_
	);
	LUT2 #(
		.INIT('h1)
	) name3192 (
		_w1180_,
		_w1712_,
		_w3654_
	);
	LUT2 #(
		.INIT('h1)
	) name3193 (
		_w1476_,
		_w3654_,
		_w3655_
	);
	LUT2 #(
		.INIT('h1)
	) name3194 (
		_w3653_,
		_w3655_,
		_w3656_
	);
	LUT2 #(
		.INIT('h2)
	) name3195 (
		_w3622_,
		_w3656_,
		_w3657_
	);
	LUT2 #(
		.INIT('h1)
	) name3196 (
		_w1404_,
		_w1916_,
		_w3658_
	);
	LUT2 #(
		.INIT('h8)
	) name3197 (
		_w3620_,
		_w3658_,
		_w3659_
	);
	LUT2 #(
		.INIT('h4)
	) name3198 (
		_w1375_,
		_w1716_,
		_w3660_
	);
	LUT2 #(
		.INIT('h1)
	) name3199 (
		_w1704_,
		_w3660_,
		_w3661_
	);
	LUT2 #(
		.INIT('h4)
	) name3200 (
		_w3659_,
		_w3661_,
		_w3662_
	);
	LUT2 #(
		.INIT('h4)
	) name3201 (
		_w3657_,
		_w3662_,
		_w3663_
	);
	LUT2 #(
		.INIT('h4)
	) name3202 (
		_w3651_,
		_w3663_,
		_w3664_
	);
	LUT2 #(
		.INIT('h1)
	) name3203 (
		_w1319_,
		_w1357_,
		_w3665_
	);
	LUT2 #(
		.INIT('h8)
	) name3204 (
		_w3606_,
		_w3665_,
		_w3666_
	);
	LUT2 #(
		.INIT('h4)
	) name3205 (
		_w950_,
		_w3613_,
		_w3667_
	);
	LUT2 #(
		.INIT('h8)
	) name3206 (
		_w3666_,
		_w3667_,
		_w3668_
	);
	LUT2 #(
		.INIT('h4)
	) name3207 (
		_w3664_,
		_w3668_,
		_w3669_
	);
	LUT2 #(
		.INIT('h1)
	) name3208 (
		_w3619_,
		_w3669_,
		_w3670_
	);
	LUT2 #(
		.INIT('h4)
	) name3209 (
		_w1832_,
		_w3670_,
		_w3671_
	);
	LUT2 #(
		.INIT('h2)
	) name3210 (
		_w1832_,
		_w3670_,
		_w3672_
	);
	LUT2 #(
		.INIT('h1)
	) name3211 (
		_w3671_,
		_w3672_,
		_w3673_
	);
	LUT2 #(
		.INIT('h8)
	) name3212 (
		_w3466_,
		_w3673_,
		_w3674_
	);
	LUT2 #(
		.INIT('h1)
	) name3213 (
		_w3467_,
		_w3674_,
		_w3675_
	);
	LUT2 #(
		.INIT('h8)
	) name3214 (
		_w501_,
		_w1888_,
		_w3676_
	);
	LUT2 #(
		.INIT('h1)
	) name3215 (
		_w1877_,
		_w3676_,
		_w3677_
	);
	LUT2 #(
		.INIT('h1)
	) name3216 (
		_w3675_,
		_w3677_,
		_w3678_
	);
	LUT2 #(
		.INIT('h8)
	) name3217 (
		_w1655_,
		_w1671_,
		_w3679_
	);
	LUT2 #(
		.INIT('h8)
	) name3218 (
		_w1609_,
		_w3679_,
		_w3680_
	);
	LUT2 #(
		.INIT('h8)
	) name3219 (
		_w1632_,
		_w3680_,
		_w3681_
	);
	LUT2 #(
		.INIT('h8)
	) name3220 (
		_w1586_,
		_w3681_,
		_w3682_
	);
	LUT2 #(
		.INIT('h8)
	) name3221 (
		_w1562_,
		_w3682_,
		_w3683_
	);
	LUT2 #(
		.INIT('h8)
	) name3222 (
		_w1537_,
		_w3683_,
		_w3684_
	);
	LUT2 #(
		.INIT('h4)
	) name3223 (
		_w1281_,
		_w1514_,
		_w3685_
	);
	LUT2 #(
		.INIT('h4)
	) name3224 (
		_w1257_,
		_w3685_,
		_w3686_
	);
	LUT2 #(
		.INIT('h8)
	) name3225 (
		_w3684_,
		_w3686_,
		_w3687_
	);
	LUT2 #(
		.INIT('h1)
	) name3226 (
		_w1198_,
		_w1233_,
		_w3688_
	);
	LUT2 #(
		.INIT('h4)
	) name3227 (
		_w1165_,
		_w3688_,
		_w3689_
	);
	LUT2 #(
		.INIT('h8)
	) name3228 (
		_w3687_,
		_w3689_,
		_w3690_
	);
	LUT2 #(
		.INIT('h1)
	) name3229 (
		_w1083_,
		_w1109_,
		_w3691_
	);
	LUT2 #(
		.INIT('h1)
	) name3230 (
		_w1136_,
		_w1466_,
		_w3692_
	);
	LUT2 #(
		.INIT('h4)
	) name3231 (
		_w1394_,
		_w3692_,
		_w3693_
	);
	LUT2 #(
		.INIT('h4)
	) name3232 (
		_w1443_,
		_w3691_,
		_w3694_
	);
	LUT2 #(
		.INIT('h8)
	) name3233 (
		_w3693_,
		_w3694_,
		_w3695_
	);
	LUT2 #(
		.INIT('h8)
	) name3234 (
		_w3690_,
		_w3695_,
		_w3696_
	);
	LUT2 #(
		.INIT('h1)
	) name3235 (
		_w1365_,
		_w1418_,
		_w3697_
	);
	LUT2 #(
		.INIT('h8)
	) name3236 (
		_w3696_,
		_w3697_,
		_w3698_
	);
	LUT2 #(
		.INIT('h1)
	) name3237 (
		_w1309_,
		_w1346_,
		_w3699_
	);
	LUT2 #(
		.INIT('h8)
	) name3238 (
		_w3698_,
		_w3699_,
		_w3700_
	);
	LUT2 #(
		.INIT('h1)
	) name3239 (
		_w1047_,
		_w1327_,
		_w3701_
	);
	LUT2 #(
		.INIT('h1)
	) name3240 (
		_w997_,
		_w1029_,
		_w3702_
	);
	LUT2 #(
		.INIT('h8)
	) name3241 (
		_w3701_,
		_w3702_,
		_w3703_
	);
	LUT2 #(
		.INIT('h8)
	) name3242 (
		_w3700_,
		_w3703_,
		_w3704_
	);
	LUT2 #(
		.INIT('h1)
	) name3243 (
		_w933_,
		_w969_,
		_w3705_
	);
	LUT2 #(
		.INIT('h8)
	) name3244 (
		_w3704_,
		_w3705_,
		_w3706_
	);
	LUT2 #(
		.INIT('h2)
	) name3245 (
		_w881_,
		_w3706_,
		_w3707_
	);
	LUT2 #(
		.INIT('h4)
	) name3246 (
		_w881_,
		_w3706_,
		_w3708_
	);
	LUT2 #(
		.INIT('h1)
	) name3247 (
		_w3707_,
		_w3708_,
		_w3709_
	);
	LUT2 #(
		.INIT('h8)
	) name3248 (
		_w3466_,
		_w3709_,
		_w3710_
	);
	LUT2 #(
		.INIT('h1)
	) name3249 (
		_w3467_,
		_w3710_,
		_w3711_
	);
	LUT2 #(
		.INIT('h8)
	) name3250 (
		_w512_,
		_w1886_,
		_w3712_
	);
	LUT2 #(
		.INIT('h4)
	) name3251 (
		_w3711_,
		_w3712_,
		_w3713_
	);
	LUT2 #(
		.INIT('h8)
	) name3252 (
		_w881_,
		_w1880_,
		_w3714_
	);
	LUT2 #(
		.INIT('h8)
	) name3253 (
		_w3466_,
		_w3714_,
		_w3715_
	);
	LUT2 #(
		.INIT('h4)
	) name3254 (
		_w1885_,
		_w1935_,
		_w3716_
	);
	LUT2 #(
		.INIT('h2)
	) name3255 (
		_w1880_,
		_w3466_,
		_w3717_
	);
	LUT2 #(
		.INIT('h1)
	) name3256 (
		_w3716_,
		_w3717_,
		_w3718_
	);
	LUT2 #(
		.INIT('h2)
	) name3257 (
		\P1_reg2_reg[29]/NET0131 ,
		_w3718_,
		_w3719_
	);
	LUT2 #(
		.INIT('h8)
	) name3258 (
		_w740_,
		_w1763_,
		_w3720_
	);
	LUT2 #(
		.INIT('h1)
	) name3259 (
		_w3719_,
		_w3720_,
		_w3721_
	);
	LUT2 #(
		.INIT('h4)
	) name3260 (
		_w3715_,
		_w3721_,
		_w3722_
	);
	LUT2 #(
		.INIT('h4)
	) name3261 (
		_w3713_,
		_w3722_,
		_w3723_
	);
	LUT2 #(
		.INIT('h4)
	) name3262 (
		_w3564_,
		_w3723_,
		_w3724_
	);
	LUT2 #(
		.INIT('h1)
	) name3263 (
		_w3605_,
		_w3678_,
		_w3725_
	);
	LUT2 #(
		.INIT('h8)
	) name3264 (
		_w3724_,
		_w3725_,
		_w3726_
	);
	LUT2 #(
		.INIT('h2)
	) name3265 (
		_w3450_,
		_w3726_,
		_w3727_
	);
	LUT2 #(
		.INIT('h1)
	) name3266 (
		_w3449_,
		_w3727_,
		_w3728_
	);
	LUT2 #(
		.INIT('h2)
	) name3267 (
		\P1_state_reg[0]/NET0131 ,
		_w3728_,
		_w3729_
	);
	LUT2 #(
		.INIT('h1)
	) name3268 (
		_w3436_,
		_w3729_,
		_w3730_
	);
	LUT2 #(
		.INIT('h2)
	) name3269 (
		\P2_reg1_reg[29]/NET0131 ,
		_w1983_,
		_w3731_
	);
	LUT2 #(
		.INIT('h8)
	) name3270 (
		\P2_reg1_reg[29]/NET0131 ,
		_w2024_,
		_w3732_
	);
	LUT2 #(
		.INIT('h2)
	) name3271 (
		_w2035_,
		_w2039_,
		_w3733_
	);
	LUT2 #(
		.INIT('h2)
	) name3272 (
		\P2_reg1_reg[29]/NET0131 ,
		_w3733_,
		_w3734_
	);
	LUT2 #(
		.INIT('h4)
	) name3273 (
		_w3161_,
		_w3733_,
		_w3735_
	);
	LUT2 #(
		.INIT('h1)
	) name3274 (
		_w3734_,
		_w3735_,
		_w3736_
	);
	LUT2 #(
		.INIT('h1)
	) name3275 (
		_w3177_,
		_w3736_,
		_w3737_
	);
	LUT2 #(
		.INIT('h8)
	) name3276 (
		_w3315_,
		_w3733_,
		_w3738_
	);
	LUT2 #(
		.INIT('h1)
	) name3277 (
		_w3734_,
		_w3738_,
		_w3739_
	);
	LUT2 #(
		.INIT('h1)
	) name3278 (
		_w3320_,
		_w3739_,
		_w3740_
	);
	LUT2 #(
		.INIT('h4)
	) name3279 (
		_w3414_,
		_w3733_,
		_w3741_
	);
	LUT2 #(
		.INIT('h2)
	) name3280 (
		_w3358_,
		_w3733_,
		_w3742_
	);
	LUT2 #(
		.INIT('h2)
	) name3281 (
		_w3421_,
		_w3742_,
		_w3743_
	);
	LUT2 #(
		.INIT('h1)
	) name3282 (
		_w3167_,
		_w3172_,
		_w3744_
	);
	LUT2 #(
		.INIT('h8)
	) name3283 (
		_w3353_,
		_w3744_,
		_w3745_
	);
	LUT2 #(
		.INIT('h4)
	) name3284 (
		_w3733_,
		_w3745_,
		_w3746_
	);
	LUT2 #(
		.INIT('h2)
	) name3285 (
		_w3743_,
		_w3746_,
		_w3747_
	);
	LUT2 #(
		.INIT('h2)
	) name3286 (
		\P2_reg1_reg[29]/NET0131 ,
		_w3747_,
		_w3748_
	);
	LUT2 #(
		.INIT('h1)
	) name3287 (
		_w3741_,
		_w3748_,
		_w3749_
	);
	LUT2 #(
		.INIT('h4)
	) name3288 (
		_w3740_,
		_w3749_,
		_w3750_
	);
	LUT2 #(
		.INIT('h4)
	) name3289 (
		_w3737_,
		_w3750_,
		_w3751_
	);
	LUT2 #(
		.INIT('h2)
	) name3290 (
		_w2026_,
		_w3751_,
		_w3752_
	);
	LUT2 #(
		.INIT('h1)
	) name3291 (
		_w3732_,
		_w3752_,
		_w3753_
	);
	LUT2 #(
		.INIT('h2)
	) name3292 (
		\P1_state_reg[0]/NET0131 ,
		_w3753_,
		_w3754_
	);
	LUT2 #(
		.INIT('h1)
	) name3293 (
		_w3731_,
		_w3754_,
		_w3755_
	);
	LUT2 #(
		.INIT('h2)
	) name3294 (
		\P2_reg2_reg[29]/NET0131 ,
		_w1983_,
		_w3756_
	);
	LUT2 #(
		.INIT('h8)
	) name3295 (
		\P2_reg2_reg[29]/NET0131 ,
		_w2024_,
		_w3757_
	);
	LUT2 #(
		.INIT('h4)
	) name3296 (
		_w2035_,
		_w2039_,
		_w3758_
	);
	LUT2 #(
		.INIT('h2)
	) name3297 (
		\P2_reg2_reg[29]/NET0131 ,
		_w3758_,
		_w3759_
	);
	LUT2 #(
		.INIT('h4)
	) name3298 (
		_w3161_,
		_w3758_,
		_w3760_
	);
	LUT2 #(
		.INIT('h1)
	) name3299 (
		_w3759_,
		_w3760_,
		_w3761_
	);
	LUT2 #(
		.INIT('h1)
	) name3300 (
		_w3177_,
		_w3761_,
		_w3762_
	);
	LUT2 #(
		.INIT('h8)
	) name3301 (
		_w3315_,
		_w3758_,
		_w3763_
	);
	LUT2 #(
		.INIT('h1)
	) name3302 (
		_w3759_,
		_w3763_,
		_w3764_
	);
	LUT2 #(
		.INIT('h1)
	) name3303 (
		_w3320_,
		_w3764_,
		_w3765_
	);
	LUT2 #(
		.INIT('h8)
	) name3304 (
		_w3352_,
		_w3758_,
		_w3766_
	);
	LUT2 #(
		.INIT('h1)
	) name3305 (
		_w3759_,
		_w3766_,
		_w3767_
	);
	LUT2 #(
		.INIT('h2)
	) name3306 (
		_w3355_,
		_w3767_,
		_w3768_
	);
	LUT2 #(
		.INIT('h4)
	) name3307 (
		_w3409_,
		_w3758_,
		_w3769_
	);
	LUT2 #(
		.INIT('h1)
	) name3308 (
		_w3759_,
		_w3769_,
		_w3770_
	);
	LUT2 #(
		.INIT('h2)
	) name3309 (
		_w3411_,
		_w3770_,
		_w3771_
	);
	LUT2 #(
		.INIT('h8)
	) name3310 (
		_w3359_,
		_w3758_,
		_w3772_
	);
	LUT2 #(
		.INIT('h2)
	) name3311 (
		_w3358_,
		_w3758_,
		_w3773_
	);
	LUT2 #(
		.INIT('h1)
	) name3312 (
		_w3417_,
		_w3773_,
		_w3774_
	);
	LUT2 #(
		.INIT('h2)
	) name3313 (
		\P2_reg2_reg[29]/NET0131 ,
		_w3774_,
		_w3775_
	);
	LUT2 #(
		.INIT('h8)
	) name3314 (
		_w2241_,
		_w3420_,
		_w3776_
	);
	LUT2 #(
		.INIT('h1)
	) name3315 (
		_w3775_,
		_w3776_,
		_w3777_
	);
	LUT2 #(
		.INIT('h4)
	) name3316 (
		_w3772_,
		_w3777_,
		_w3778_
	);
	LUT2 #(
		.INIT('h4)
	) name3317 (
		_w3771_,
		_w3778_,
		_w3779_
	);
	LUT2 #(
		.INIT('h4)
	) name3318 (
		_w3768_,
		_w3779_,
		_w3780_
	);
	LUT2 #(
		.INIT('h4)
	) name3319 (
		_w3765_,
		_w3780_,
		_w3781_
	);
	LUT2 #(
		.INIT('h4)
	) name3320 (
		_w3762_,
		_w3781_,
		_w3782_
	);
	LUT2 #(
		.INIT('h2)
	) name3321 (
		_w2026_,
		_w3782_,
		_w3783_
	);
	LUT2 #(
		.INIT('h1)
	) name3322 (
		_w3757_,
		_w3783_,
		_w3784_
	);
	LUT2 #(
		.INIT('h2)
	) name3323 (
		\P1_state_reg[0]/NET0131 ,
		_w3784_,
		_w3785_
	);
	LUT2 #(
		.INIT('h1)
	) name3324 (
		_w3756_,
		_w3785_,
		_w3786_
	);
	LUT2 #(
		.INIT('h2)
	) name3325 (
		_w2024_,
		_w2958_,
		_w3787_
	);
	LUT2 #(
		.INIT('h1)
	) name3326 (
		_w2035_,
		_w2039_,
		_w3788_
	);
	LUT2 #(
		.INIT('h1)
	) name3327 (
		_w2958_,
		_w3788_,
		_w3789_
	);
	LUT2 #(
		.INIT('h1)
	) name3328 (
		_w3183_,
		_w3187_,
		_w3790_
	);
	LUT2 #(
		.INIT('h1)
	) name3329 (
		_w3180_,
		_w3182_,
		_w3791_
	);
	LUT2 #(
		.INIT('h8)
	) name3330 (
		_w3790_,
		_w3791_,
		_w3792_
	);
	LUT2 #(
		.INIT('h1)
	) name3331 (
		_w3186_,
		_w3189_,
		_w3793_
	);
	LUT2 #(
		.INIT('h1)
	) name3332 (
		_w3211_,
		_w3305_,
		_w3794_
	);
	LUT2 #(
		.INIT('h8)
	) name3333 (
		_w3793_,
		_w3794_,
		_w3795_
	);
	LUT2 #(
		.INIT('h8)
	) name3334 (
		_w3792_,
		_w3795_,
		_w3796_
	);
	LUT2 #(
		.INIT('h1)
	) name3335 (
		_w3210_,
		_w3214_,
		_w3797_
	);
	LUT2 #(
		.INIT('h1)
	) name3336 (
		_w3213_,
		_w3217_,
		_w3798_
	);
	LUT2 #(
		.INIT('h8)
	) name3337 (
		_w3797_,
		_w3798_,
		_w3799_
	);
	LUT2 #(
		.INIT('h1)
	) name3338 (
		_w3218_,
		_w3220_,
		_w3800_
	);
	LUT2 #(
		.INIT('h1)
	) name3339 (
		_w3234_,
		_w3283_,
		_w3801_
	);
	LUT2 #(
		.INIT('h1)
	) name3340 (
		_w3221_,
		_w3801_,
		_w3802_
	);
	LUT2 #(
		.INIT('h8)
	) name3341 (
		_w3800_,
		_w3802_,
		_w3803_
	);
	LUT2 #(
		.INIT('h1)
	) name3342 (
		_w3282_,
		_w3288_,
		_w3804_
	);
	LUT2 #(
		.INIT('h1)
	) name3343 (
		_w3218_,
		_w3804_,
		_w3805_
	);
	LUT2 #(
		.INIT('h1)
	) name3344 (
		_w3803_,
		_w3805_,
		_w3806_
	);
	LUT2 #(
		.INIT('h2)
	) name3345 (
		_w3799_,
		_w3806_,
		_w3807_
	);
	LUT2 #(
		.INIT('h4)
	) name3346 (
		_w3213_,
		_w3287_,
		_w3808_
	);
	LUT2 #(
		.INIT('h1)
	) name3347 (
		_w3294_,
		_w3808_,
		_w3809_
	);
	LUT2 #(
		.INIT('h2)
	) name3348 (
		_w3797_,
		_w3809_,
		_w3810_
	);
	LUT2 #(
		.INIT('h4)
	) name3349 (
		_w3210_,
		_w3293_,
		_w3811_
	);
	LUT2 #(
		.INIT('h1)
	) name3350 (
		_w3299_,
		_w3811_,
		_w3812_
	);
	LUT2 #(
		.INIT('h4)
	) name3351 (
		_w3810_,
		_w3812_,
		_w3813_
	);
	LUT2 #(
		.INIT('h1)
	) name3352 (
		_w3239_,
		_w3242_,
		_w3814_
	);
	LUT2 #(
		.INIT('h1)
	) name3353 (
		_w3225_,
		_w3229_,
		_w3815_
	);
	LUT2 #(
		.INIT('h8)
	) name3354 (
		_w3814_,
		_w3815_,
		_w3816_
	);
	LUT2 #(
		.INIT('h1)
	) name3355 (
		_w3241_,
		_w3244_,
		_w3817_
	);
	LUT2 #(
		.INIT('h1)
	) name3356 (
		_w3264_,
		_w3272_,
		_w3818_
	);
	LUT2 #(
		.INIT('h1)
	) name3357 (
		_w3255_,
		_w3259_,
		_w3819_
	);
	LUT2 #(
		.INIT('h2)
	) name3358 (
		_w3263_,
		_w3819_,
		_w3820_
	);
	LUT2 #(
		.INIT('h1)
	) name3359 (
		_w3254_,
		_w3268_,
		_w3821_
	);
	LUT2 #(
		.INIT('h1)
	) name3360 (
		_w3262_,
		_w3821_,
		_w3822_
	);
	LUT2 #(
		.INIT('h1)
	) name3361 (
		_w3820_,
		_w3822_,
		_w3823_
	);
	LUT2 #(
		.INIT('h2)
	) name3362 (
		_w3818_,
		_w3823_,
		_w3824_
	);
	LUT2 #(
		.INIT('h2)
	) name3363 (
		_w3267_,
		_w3272_,
		_w3825_
	);
	LUT2 #(
		.INIT('h1)
	) name3364 (
		_w3246_,
		_w3825_,
		_w3826_
	);
	LUT2 #(
		.INIT('h4)
	) name3365 (
		_w3824_,
		_w3826_,
		_w3827_
	);
	LUT2 #(
		.INIT('h2)
	) name3366 (
		_w3817_,
		_w3827_,
		_w3828_
	);
	LUT2 #(
		.INIT('h1)
	) name3367 (
		_w3245_,
		_w3251_,
		_w3829_
	);
	LUT2 #(
		.INIT('h1)
	) name3368 (
		_w3241_,
		_w3829_,
		_w3830_
	);
	LUT2 #(
		.INIT('h1)
	) name3369 (
		_w3828_,
		_w3830_,
		_w3831_
	);
	LUT2 #(
		.INIT('h2)
	) name3370 (
		_w3816_,
		_w3831_,
		_w3832_
	);
	LUT2 #(
		.INIT('h1)
	) name3371 (
		_w3230_,
		_w3250_,
		_w3833_
	);
	LUT2 #(
		.INIT('h1)
	) name3372 (
		_w3239_,
		_w3833_,
		_w3834_
	);
	LUT2 #(
		.INIT('h8)
	) name3373 (
		_w3815_,
		_w3834_,
		_w3835_
	);
	LUT2 #(
		.INIT('h1)
	) name3374 (
		_w3228_,
		_w3235_,
		_w3836_
	);
	LUT2 #(
		.INIT('h1)
	) name3375 (
		_w3225_,
		_w3836_,
		_w3837_
	);
	LUT2 #(
		.INIT('h1)
	) name3376 (
		_w3835_,
		_w3837_,
		_w3838_
	);
	LUT2 #(
		.INIT('h4)
	) name3377 (
		_w3832_,
		_w3838_,
		_w3839_
	);
	LUT2 #(
		.INIT('h1)
	) name3378 (
		_w3221_,
		_w3226_,
		_w3840_
	);
	LUT2 #(
		.INIT('h8)
	) name3379 (
		_w3800_,
		_w3840_,
		_w3841_
	);
	LUT2 #(
		.INIT('h8)
	) name3380 (
		_w3799_,
		_w3841_,
		_w3842_
	);
	LUT2 #(
		.INIT('h4)
	) name3381 (
		_w3839_,
		_w3842_,
		_w3843_
	);
	LUT2 #(
		.INIT('h4)
	) name3382 (
		_w3807_,
		_w3813_,
		_w3844_
	);
	LUT2 #(
		.INIT('h4)
	) name3383 (
		_w3843_,
		_w3844_,
		_w3845_
	);
	LUT2 #(
		.INIT('h2)
	) name3384 (
		_w3796_,
		_w3845_,
		_w3846_
	);
	LUT2 #(
		.INIT('h2)
	) name3385 (
		_w3298_,
		_w3305_,
		_w3847_
	);
	LUT2 #(
		.INIT('h1)
	) name3386 (
		_w3191_,
		_w3847_,
		_w3848_
	);
	LUT2 #(
		.INIT('h2)
	) name3387 (
		_w3793_,
		_w3848_,
		_w3849_
	);
	LUT2 #(
		.INIT('h1)
	) name3388 (
		_w3190_,
		_w3196_,
		_w3850_
	);
	LUT2 #(
		.INIT('h1)
	) name3389 (
		_w3186_,
		_w3850_,
		_w3851_
	);
	LUT2 #(
		.INIT('h1)
	) name3390 (
		_w3849_,
		_w3851_,
		_w3852_
	);
	LUT2 #(
		.INIT('h2)
	) name3391 (
		_w3792_,
		_w3852_,
		_w3853_
	);
	LUT2 #(
		.INIT('h1)
	) name3392 (
		_w3201_,
		_w3207_,
		_w3854_
	);
	LUT2 #(
		.INIT('h1)
	) name3393 (
		_w3195_,
		_w3202_,
		_w3855_
	);
	LUT2 #(
		.INIT('h1)
	) name3394 (
		_w3183_,
		_w3855_,
		_w3856_
	);
	LUT2 #(
		.INIT('h4)
	) name3395 (
		_w3182_,
		_w3856_,
		_w3857_
	);
	LUT2 #(
		.INIT('h2)
	) name3396 (
		_w3854_,
		_w3857_,
		_w3858_
	);
	LUT2 #(
		.INIT('h1)
	) name3397 (
		_w3180_,
		_w3858_,
		_w3859_
	);
	LUT2 #(
		.INIT('h1)
	) name3398 (
		_w3846_,
		_w3853_,
		_w3860_
	);
	LUT2 #(
		.INIT('h4)
	) name3399 (
		_w3859_,
		_w3860_,
		_w3861_
	);
	LUT2 #(
		.INIT('h1)
	) name3400 (
		_w2963_,
		_w3154_,
		_w3862_
	);
	LUT2 #(
		.INIT('h4)
	) name3401 (
		_w3861_,
		_w3862_,
		_w3863_
	);
	LUT2 #(
		.INIT('h2)
	) name3402 (
		_w3861_,
		_w3862_,
		_w3864_
	);
	LUT2 #(
		.INIT('h1)
	) name3403 (
		_w3863_,
		_w3864_,
		_w3865_
	);
	LUT2 #(
		.INIT('h2)
	) name3404 (
		_w3788_,
		_w3865_,
		_w3866_
	);
	LUT2 #(
		.INIT('h1)
	) name3405 (
		_w3789_,
		_w3866_,
		_w3867_
	);
	LUT2 #(
		.INIT('h1)
	) name3406 (
		_w3320_,
		_w3867_,
		_w3868_
	);
	LUT2 #(
		.INIT('h1)
	) name3407 (
		_w2705_,
		_w2756_,
		_w3869_
	);
	LUT2 #(
		.INIT('h2)
	) name3408 (
		_w2673_,
		_w2780_,
		_w3870_
	);
	LUT2 #(
		.INIT('h1)
	) name3409 (
		_w2785_,
		_w3870_,
		_w3871_
	);
	LUT2 #(
		.INIT('h2)
	) name3410 (
		_w3869_,
		_w3871_,
		_w3872_
	);
	LUT2 #(
		.INIT('h4)
	) name3411 (
		_w2705_,
		_w2784_,
		_w3873_
	);
	LUT2 #(
		.INIT('h1)
	) name3412 (
		_w2790_,
		_w3873_,
		_w3874_
	);
	LUT2 #(
		.INIT('h4)
	) name3413 (
		_w3872_,
		_w3874_,
		_w3875_
	);
	LUT2 #(
		.INIT('h1)
	) name3414 (
		_w2496_,
		_w2522_,
		_w3876_
	);
	LUT2 #(
		.INIT('h8)
	) name3415 (
		_w2607_,
		_w2633_,
		_w3877_
	);
	LUT2 #(
		.INIT('h1)
	) name3416 (
		_w2567_,
		_w2661_,
		_w3878_
	);
	LUT2 #(
		.INIT('h1)
	) name3417 (
		_w2632_,
		_w3878_,
		_w3879_
	);
	LUT2 #(
		.INIT('h1)
	) name3418 (
		_w3877_,
		_w3879_,
		_w3880_
	);
	LUT2 #(
		.INIT('h1)
	) name3419 (
		_w2545_,
		_w2657_,
		_w3881_
	);
	LUT2 #(
		.INIT('h4)
	) name3420 (
		_w3880_,
		_w3881_,
		_w3882_
	);
	LUT2 #(
		.INIT('h1)
	) name3421 (
		_w2660_,
		_w2669_,
		_w3883_
	);
	LUT2 #(
		.INIT('h1)
	) name3422 (
		_w2545_,
		_w3883_,
		_w3884_
	);
	LUT2 #(
		.INIT('h1)
	) name3423 (
		_w3882_,
		_w3884_,
		_w3885_
	);
	LUT2 #(
		.INIT('h2)
	) name3424 (
		_w3876_,
		_w3885_,
		_w3886_
	);
	LUT2 #(
		.INIT('h1)
	) name3425 (
		_w2668_,
		_w2674_,
		_w3887_
	);
	LUT2 #(
		.INIT('h1)
	) name3426 (
		_w2496_,
		_w3887_,
		_w3888_
	);
	LUT2 #(
		.INIT('h1)
	) name3427 (
		_w3886_,
		_w3888_,
		_w3889_
	);
	LUT2 #(
		.INIT('h1)
	) name3428 (
		_w2471_,
		_w2780_,
		_w3890_
	);
	LUT2 #(
		.INIT('h8)
	) name3429 (
		_w3869_,
		_w3890_,
		_w3891_
	);
	LUT2 #(
		.INIT('h4)
	) name3430 (
		_w3889_,
		_w3891_,
		_w3892_
	);
	LUT2 #(
		.INIT('h2)
	) name3431 (
		_w3875_,
		_w3892_,
		_w3893_
	);
	LUT2 #(
		.INIT('h1)
	) name3432 (
		_w2844_,
		_w2871_,
		_w3894_
	);
	LUT2 #(
		.INIT('h1)
	) name3433 (
		_w2732_,
		_w2894_,
		_w3895_
	);
	LUT2 #(
		.INIT('h8)
	) name3434 (
		_w3894_,
		_w3895_,
		_w3896_
	);
	LUT2 #(
		.INIT('h1)
	) name3435 (
		_w2400_,
		_w2819_,
		_w3897_
	);
	LUT2 #(
		.INIT('h1)
	) name3436 (
		_w2312_,
		_w2443_,
		_w3898_
	);
	LUT2 #(
		.INIT('h8)
	) name3437 (
		_w3897_,
		_w3898_,
		_w3899_
	);
	LUT2 #(
		.INIT('h8)
	) name3438 (
		_w3896_,
		_w3899_,
		_w3900_
	);
	LUT2 #(
		.INIT('h4)
	) name3439 (
		_w3893_,
		_w3900_,
		_w3901_
	);
	LUT2 #(
		.INIT('h1)
	) name3440 (
		_w2789_,
		_w2900_,
		_w3902_
	);
	LUT2 #(
		.INIT('h1)
	) name3441 (
		_w2894_,
		_w3902_,
		_w3903_
	);
	LUT2 #(
		.INIT('h8)
	) name3442 (
		_w3894_,
		_w3903_,
		_w3904_
	);
	LUT2 #(
		.INIT('h1)
	) name3443 (
		_w2899_,
		_w2905_,
		_w3905_
	);
	LUT2 #(
		.INIT('h1)
	) name3444 (
		_w2844_,
		_w3905_,
		_w3906_
	);
	LUT2 #(
		.INIT('h1)
	) name3445 (
		_w3904_,
		_w3906_,
		_w3907_
	);
	LUT2 #(
		.INIT('h2)
	) name3446 (
		_w3899_,
		_w3907_,
		_w3908_
	);
	LUT2 #(
		.INIT('h1)
	) name3447 (
		_w2904_,
		_w2911_,
		_w3909_
	);
	LUT2 #(
		.INIT('h1)
	) name3448 (
		_w2400_,
		_w3909_,
		_w3910_
	);
	LUT2 #(
		.INIT('h8)
	) name3449 (
		_w3898_,
		_w3910_,
		_w3911_
	);
	LUT2 #(
		.INIT('h4)
	) name3450 (
		_w2312_,
		_w2910_,
		_w3912_
	);
	LUT2 #(
		.INIT('h1)
	) name3451 (
		_w2916_,
		_w3912_,
		_w3913_
	);
	LUT2 #(
		.INIT('h4)
	) name3452 (
		_w3911_,
		_w3913_,
		_w3914_
	);
	LUT2 #(
		.INIT('h4)
	) name3453 (
		_w3908_,
		_w3914_,
		_w3915_
	);
	LUT2 #(
		.INIT('h4)
	) name3454 (
		_w3901_,
		_w3915_,
		_w3916_
	);
	LUT2 #(
		.INIT('h1)
	) name3455 (
		_w3044_,
		_w3066_,
		_w3917_
	);
	LUT2 #(
		.INIT('h1)
	) name3456 (
		_w2992_,
		_w3022_,
		_w3918_
	);
	LUT2 #(
		.INIT('h8)
	) name3457 (
		_w3917_,
		_w3918_,
		_w3919_
	);
	LUT2 #(
		.INIT('h1)
	) name3458 (
		_w3089_,
		_w3113_,
		_w3920_
	);
	LUT2 #(
		.INIT('h1)
	) name3459 (
		_w2369_,
		_w3131_,
		_w3921_
	);
	LUT2 #(
		.INIT('h8)
	) name3460 (
		_w3920_,
		_w3921_,
		_w3922_
	);
	LUT2 #(
		.INIT('h8)
	) name3461 (
		_w3919_,
		_w3922_,
		_w3923_
	);
	LUT2 #(
		.INIT('h4)
	) name3462 (
		_w3916_,
		_w3923_,
		_w3924_
	);
	LUT2 #(
		.INIT('h2)
	) name3463 (
		_w2915_,
		_w3131_,
		_w3925_
	);
	LUT2 #(
		.INIT('h1)
	) name3464 (
		_w3139_,
		_w3925_,
		_w3926_
	);
	LUT2 #(
		.INIT('h2)
	) name3465 (
		_w3920_,
		_w3926_,
		_w3927_
	);
	LUT2 #(
		.INIT('h4)
	) name3466 (
		_w3089_,
		_w3138_,
		_w3928_
	);
	LUT2 #(
		.INIT('h1)
	) name3467 (
		_w3144_,
		_w3928_,
		_w3929_
	);
	LUT2 #(
		.INIT('h4)
	) name3468 (
		_w3927_,
		_w3929_,
		_w3930_
	);
	LUT2 #(
		.INIT('h2)
	) name3469 (
		_w3919_,
		_w3930_,
		_w3931_
	);
	LUT2 #(
		.INIT('h4)
	) name3470 (
		_w3044_,
		_w3143_,
		_w3932_
	);
	LUT2 #(
		.INIT('h1)
	) name3471 (
		_w3150_,
		_w3932_,
		_w3933_
	);
	LUT2 #(
		.INIT('h2)
	) name3472 (
		_w3918_,
		_w3933_,
		_w3934_
	);
	LUT2 #(
		.INIT('h4)
	) name3473 (
		_w2992_,
		_w3149_,
		_w3935_
	);
	LUT2 #(
		.INIT('h1)
	) name3474 (
		_w3136_,
		_w3935_,
		_w3936_
	);
	LUT2 #(
		.INIT('h4)
	) name3475 (
		_w3934_,
		_w3936_,
		_w3937_
	);
	LUT2 #(
		.INIT('h4)
	) name3476 (
		_w3931_,
		_w3937_,
		_w3938_
	);
	LUT2 #(
		.INIT('h4)
	) name3477 (
		_w3924_,
		_w3938_,
		_w3939_
	);
	LUT2 #(
		.INIT('h8)
	) name3478 (
		_w3862_,
		_w3939_,
		_w3940_
	);
	LUT2 #(
		.INIT('h1)
	) name3479 (
		_w3862_,
		_w3939_,
		_w3941_
	);
	LUT2 #(
		.INIT('h1)
	) name3480 (
		_w3940_,
		_w3941_,
		_w3942_
	);
	LUT2 #(
		.INIT('h2)
	) name3481 (
		_w3788_,
		_w3942_,
		_w3943_
	);
	LUT2 #(
		.INIT('h1)
	) name3482 (
		_w3789_,
		_w3943_,
		_w3944_
	);
	LUT2 #(
		.INIT('h1)
	) name3483 (
		_w3177_,
		_w3944_,
		_w3945_
	);
	LUT2 #(
		.INIT('h8)
	) name3484 (
		_w3346_,
		_w3347_,
		_w3946_
	);
	LUT2 #(
		.INIT('h2)
	) name3485 (
		_w2949_,
		_w3946_,
		_w3947_
	);
	LUT2 #(
		.INIT('h1)
	) name3486 (
		_w3349_,
		_w3947_,
		_w3948_
	);
	LUT2 #(
		.INIT('h8)
	) name3487 (
		_w3788_,
		_w3948_,
		_w3949_
	);
	LUT2 #(
		.INIT('h1)
	) name3488 (
		_w3789_,
		_w3949_,
		_w3950_
	);
	LUT2 #(
		.INIT('h2)
	) name3489 (
		_w3355_,
		_w3950_,
		_w3951_
	);
	LUT2 #(
		.INIT('h8)
	) name3490 (
		_w3366_,
		_w3394_,
		_w3952_
	);
	LUT2 #(
		.INIT('h2)
	) name3491 (
		_w2251_,
		_w3952_,
		_w3953_
	);
	LUT2 #(
		.INIT('h1)
	) name3492 (
		_w3396_,
		_w3953_,
		_w3954_
	);
	LUT2 #(
		.INIT('h1)
	) name3493 (
		_w2058_,
		_w3954_,
		_w3955_
	);
	LUT2 #(
		.INIT('h8)
	) name3494 (
		_w2058_,
		_w2991_,
		_w3956_
	);
	LUT2 #(
		.INIT('h1)
	) name3495 (
		_w3955_,
		_w3956_,
		_w3957_
	);
	LUT2 #(
		.INIT('h8)
	) name3496 (
		_w3788_,
		_w3957_,
		_w3958_
	);
	LUT2 #(
		.INIT('h1)
	) name3497 (
		_w3789_,
		_w3958_,
		_w3959_
	);
	LUT2 #(
		.INIT('h2)
	) name3498 (
		_w3411_,
		_w3959_,
		_w3960_
	);
	LUT2 #(
		.INIT('h2)
	) name3499 (
		_w3358_,
		_w3788_,
		_w3961_
	);
	LUT2 #(
		.INIT('h1)
	) name3500 (
		_w3417_,
		_w3961_,
		_w3962_
	);
	LUT2 #(
		.INIT('h1)
	) name3501 (
		_w2958_,
		_w3962_,
		_w3963_
	);
	LUT2 #(
		.INIT('h8)
	) name3502 (
		_w3358_,
		_w3788_,
		_w3964_
	);
	LUT2 #(
		.INIT('h1)
	) name3503 (
		_w3420_,
		_w3964_,
		_w3965_
	);
	LUT2 #(
		.INIT('h2)
	) name3504 (
		_w2949_,
		_w3965_,
		_w3966_
	);
	LUT2 #(
		.INIT('h1)
	) name3505 (
		_w3963_,
		_w3966_,
		_w3967_
	);
	LUT2 #(
		.INIT('h4)
	) name3506 (
		_w3960_,
		_w3967_,
		_w3968_
	);
	LUT2 #(
		.INIT('h4)
	) name3507 (
		_w3951_,
		_w3968_,
		_w3969_
	);
	LUT2 #(
		.INIT('h4)
	) name3508 (
		_w3945_,
		_w3969_,
		_w3970_
	);
	LUT2 #(
		.INIT('h4)
	) name3509 (
		_w3868_,
		_w3970_,
		_w3971_
	);
	LUT2 #(
		.INIT('h2)
	) name3510 (
		_w2026_,
		_w3971_,
		_w3972_
	);
	LUT2 #(
		.INIT('h1)
	) name3511 (
		_w3787_,
		_w3972_,
		_w3973_
	);
	LUT2 #(
		.INIT('h2)
	) name3512 (
		\P1_state_reg[0]/NET0131 ,
		_w3973_,
		_w3974_
	);
	LUT2 #(
		.INIT('h4)
	) name3513 (
		\P1_state_reg[0]/NET0131 ,
		\P2_reg3_reg[28]/NET0131 ,
		_w3975_
	);
	LUT2 #(
		.INIT('h8)
	) name3514 (
		\P1_state_reg[0]/NET0131 ,
		_w1982_,
		_w3976_
	);
	LUT2 #(
		.INIT('h4)
	) name3515 (
		_w2958_,
		_w3976_,
		_w3977_
	);
	LUT2 #(
		.INIT('h1)
	) name3516 (
		_w3975_,
		_w3977_,
		_w3978_
	);
	LUT2 #(
		.INIT('h4)
	) name3517 (
		_w3974_,
		_w3978_,
		_w3979_
	);
	LUT2 #(
		.INIT('h1)
	) name3518 (
		_w3460_,
		_w3465_,
		_w3980_
	);
	LUT2 #(
		.INIT('h2)
	) name3519 (
		_w941_,
		_w3980_,
		_w3981_
	);
	LUT2 #(
		.INIT('h1)
	) name3520 (
		_w1774_,
		_w3499_,
		_w3982_
	);
	LUT2 #(
		.INIT('h8)
	) name3521 (
		_w3507_,
		_w3510_,
		_w3983_
	);
	LUT2 #(
		.INIT('h1)
	) name3522 (
		_w1777_,
		_w3515_,
		_w3984_
	);
	LUT2 #(
		.INIT('h1)
	) name3523 (
		_w3509_,
		_w3984_,
		_w3985_
	);
	LUT2 #(
		.INIT('h1)
	) name3524 (
		_w3983_,
		_w3985_,
		_w3986_
	);
	LUT2 #(
		.INIT('h1)
	) name3525 (
		_w3500_,
		_w3511_,
		_w3987_
	);
	LUT2 #(
		.INIT('h4)
	) name3526 (
		_w3986_,
		_w3987_,
		_w3988_
	);
	LUT2 #(
		.INIT('h8)
	) name3527 (
		_w3982_,
		_w3988_,
		_w3989_
	);
	LUT2 #(
		.INIT('h4)
	) name3528 (
		_w3500_,
		_w3514_,
		_w3990_
	);
	LUT2 #(
		.INIT('h1)
	) name3529 (
		_w3522_,
		_w3990_,
		_w3991_
	);
	LUT2 #(
		.INIT('h2)
	) name3530 (
		_w3982_,
		_w3991_,
		_w3992_
	);
	LUT2 #(
		.INIT('h4)
	) name3531 (
		_w1774_,
		_w3521_,
		_w3993_
	);
	LUT2 #(
		.INIT('h1)
	) name3532 (
		_w1775_,
		_w3993_,
		_w3994_
	);
	LUT2 #(
		.INIT('h4)
	) name3533 (
		_w3992_,
		_w3994_,
		_w3995_
	);
	LUT2 #(
		.INIT('h4)
	) name3534 (
		_w3989_,
		_w3995_,
		_w3996_
	);
	LUT2 #(
		.INIT('h1)
	) name3535 (
		_w1781_,
		_w1800_,
		_w3997_
	);
	LUT2 #(
		.INIT('h1)
	) name3536 (
		_w1770_,
		_w1790_,
		_w3998_
	);
	LUT2 #(
		.INIT('h8)
	) name3537 (
		_w3997_,
		_w3998_,
		_w3999_
	);
	LUT2 #(
		.INIT('h4)
	) name3538 (
		_w3996_,
		_w3999_,
		_w4000_
	);
	LUT2 #(
		.INIT('h4)
	) name3539 (
		_w1781_,
		_w1801_,
		_w4001_
	);
	LUT2 #(
		.INIT('h1)
	) name3540 (
		_w1780_,
		_w4001_,
		_w4002_
	);
	LUT2 #(
		.INIT('h2)
	) name3541 (
		_w3998_,
		_w4002_,
		_w4003_
	);
	LUT2 #(
		.INIT('h1)
	) name3542 (
		_w1771_,
		_w1789_,
		_w4004_
	);
	LUT2 #(
		.INIT('h1)
	) name3543 (
		_w1770_,
		_w4004_,
		_w4005_
	);
	LUT2 #(
		.INIT('h1)
	) name3544 (
		_w4003_,
		_w4005_,
		_w4006_
	);
	LUT2 #(
		.INIT('h4)
	) name3545 (
		_w4000_,
		_w4006_,
		_w4007_
	);
	LUT2 #(
		.INIT('h1)
	) name3546 (
		_w1794_,
		_w1797_,
		_w4008_
	);
	LUT2 #(
		.INIT('h1)
	) name3547 (
		_w1786_,
		_w1813_,
		_w4009_
	);
	LUT2 #(
		.INIT('h8)
	) name3548 (
		_w4008_,
		_w4009_,
		_w4010_
	);
	LUT2 #(
		.INIT('h1)
	) name3549 (
		_w1783_,
		_w3485_,
		_w4011_
	);
	LUT2 #(
		.INIT('h1)
	) name3550 (
		_w1822_,
		_w1833_,
		_w4012_
	);
	LUT2 #(
		.INIT('h8)
	) name3551 (
		_w4011_,
		_w4012_,
		_w4013_
	);
	LUT2 #(
		.INIT('h8)
	) name3552 (
		_w4010_,
		_w4013_,
		_w4014_
	);
	LUT2 #(
		.INIT('h4)
	) name3553 (
		_w4007_,
		_w4014_,
		_w4015_
	);
	LUT2 #(
		.INIT('h2)
	) name3554 (
		_w1795_,
		_w1797_,
		_w4016_
	);
	LUT2 #(
		.INIT('h1)
	) name3555 (
		_w1798_,
		_w4016_,
		_w4017_
	);
	LUT2 #(
		.INIT('h2)
	) name3556 (
		_w4009_,
		_w4017_,
		_w4018_
	);
	LUT2 #(
		.INIT('h4)
	) name3557 (
		_w1786_,
		_w1814_,
		_w4019_
	);
	LUT2 #(
		.INIT('h1)
	) name3558 (
		_w1787_,
		_w4019_,
		_w4020_
	);
	LUT2 #(
		.INIT('h4)
	) name3559 (
		_w4018_,
		_w4020_,
		_w4021_
	);
	LUT2 #(
		.INIT('h2)
	) name3560 (
		_w4013_,
		_w4021_,
		_w4022_
	);
	LUT2 #(
		.INIT('h1)
	) name3561 (
		_w1784_,
		_w3542_,
		_w4023_
	);
	LUT2 #(
		.INIT('h1)
	) name3562 (
		_w3485_,
		_w4023_,
		_w4024_
	);
	LUT2 #(
		.INIT('h8)
	) name3563 (
		_w4012_,
		_w4024_,
		_w4025_
	);
	LUT2 #(
		.INIT('h1)
	) name3564 (
		_w1823_,
		_w1834_,
		_w4026_
	);
	LUT2 #(
		.INIT('h1)
	) name3565 (
		_w1833_,
		_w4026_,
		_w4027_
	);
	LUT2 #(
		.INIT('h1)
	) name3566 (
		_w4025_,
		_w4027_,
		_w4028_
	);
	LUT2 #(
		.INIT('h4)
	) name3567 (
		_w4022_,
		_w4028_,
		_w4029_
	);
	LUT2 #(
		.INIT('h4)
	) name3568 (
		_w4015_,
		_w4029_,
		_w4030_
	);
	LUT2 #(
		.INIT('h1)
	) name3569 (
		_w1820_,
		_w1836_,
		_w4031_
	);
	LUT2 #(
		.INIT('h1)
	) name3570 (
		_w1826_,
		_w1839_,
		_w4032_
	);
	LUT2 #(
		.INIT('h8)
	) name3571 (
		_w4031_,
		_w4032_,
		_w4033_
	);
	LUT2 #(
		.INIT('h4)
	) name3572 (
		_w1816_,
		_w3476_,
		_w4034_
	);
	LUT2 #(
		.INIT('h8)
	) name3573 (
		_w4033_,
		_w4034_,
		_w4035_
	);
	LUT2 #(
		.INIT('h4)
	) name3574 (
		_w4030_,
		_w4035_,
		_w4036_
	);
	LUT2 #(
		.INIT('h4)
	) name3575 (
		_w1767_,
		_w1807_,
		_w4037_
	);
	LUT2 #(
		.INIT('h2)
	) name3576 (
		_w1827_,
		_w1839_,
		_w4038_
	);
	LUT2 #(
		.INIT('h1)
	) name3577 (
		_w1840_,
		_w4038_,
		_w4039_
	);
	LUT2 #(
		.INIT('h2)
	) name3578 (
		_w4031_,
		_w4039_,
		_w4040_
	);
	LUT2 #(
		.INIT('h4)
	) name3579 (
		_w1820_,
		_w1837_,
		_w4041_
	);
	LUT2 #(
		.INIT('h1)
	) name3580 (
		_w1819_,
		_w4041_,
		_w4042_
	);
	LUT2 #(
		.INIT('h4)
	) name3581 (
		_w4040_,
		_w4042_,
		_w4043_
	);
	LUT2 #(
		.INIT('h2)
	) name3582 (
		_w4034_,
		_w4043_,
		_w4044_
	);
	LUT2 #(
		.INIT('h1)
	) name3583 (
		_w1811_,
		_w1817_,
		_w4045_
	);
	LUT2 #(
		.INIT('h2)
	) name3584 (
		_w3476_,
		_w4045_,
		_w4046_
	);
	LUT2 #(
		.INIT('h1)
	) name3585 (
		_w1768_,
		_w4037_,
		_w4047_
	);
	LUT2 #(
		.INIT('h4)
	) name3586 (
		_w4046_,
		_w4047_,
		_w4048_
	);
	LUT2 #(
		.INIT('h4)
	) name3587 (
		_w4044_,
		_w4048_,
		_w4049_
	);
	LUT2 #(
		.INIT('h4)
	) name3588 (
		_w4036_,
		_w4049_,
		_w4050_
	);
	LUT2 #(
		.INIT('h8)
	) name3589 (
		_w1831_,
		_w4050_,
		_w4051_
	);
	LUT2 #(
		.INIT('h1)
	) name3590 (
		_w1831_,
		_w4050_,
		_w4052_
	);
	LUT2 #(
		.INIT('h1)
	) name3591 (
		_w4051_,
		_w4052_,
		_w4053_
	);
	LUT2 #(
		.INIT('h2)
	) name3592 (
		_w3980_,
		_w4053_,
		_w4054_
	);
	LUT2 #(
		.INIT('h1)
	) name3593 (
		_w3981_,
		_w4054_,
		_w4055_
	);
	LUT2 #(
		.INIT('h1)
	) name3594 (
		_w3563_,
		_w4055_,
		_w4056_
	);
	LUT2 #(
		.INIT('h4)
	) name3595 (
		_w969_,
		_w3704_,
		_w4057_
	);
	LUT2 #(
		.INIT('h2)
	) name3596 (
		_w933_,
		_w4057_,
		_w4058_
	);
	LUT2 #(
		.INIT('h1)
	) name3597 (
		_w3706_,
		_w4058_,
		_w4059_
	);
	LUT2 #(
		.INIT('h8)
	) name3598 (
		_w3980_,
		_w4059_,
		_w4060_
	);
	LUT2 #(
		.INIT('h1)
	) name3599 (
		_w3981_,
		_w4060_,
		_w4061_
	);
	LUT2 #(
		.INIT('h2)
	) name3600 (
		_w3712_,
		_w4061_,
		_w4062_
	);
	LUT2 #(
		.INIT('h2)
	) name3601 (
		_w1880_,
		_w3980_,
		_w4063_
	);
	LUT2 #(
		.INIT('h1)
	) name3602 (
		_w3716_,
		_w4063_,
		_w4064_
	);
	LUT2 #(
		.INIT('h2)
	) name3603 (
		_w941_,
		_w4064_,
		_w4065_
	);
	LUT2 #(
		.INIT('h8)
	) name3604 (
		_w1880_,
		_w3980_,
		_w4066_
	);
	LUT2 #(
		.INIT('h1)
	) name3605 (
		_w1763_,
		_w4066_,
		_w4067_
	);
	LUT2 #(
		.INIT('h2)
	) name3606 (
		_w933_,
		_w4067_,
		_w4068_
	);
	LUT2 #(
		.INIT('h4)
	) name3607 (
		_w1207_,
		_w3580_,
		_w4069_
	);
	LUT2 #(
		.INIT('h4)
	) name3608 (
		_w1174_,
		_w4069_,
		_w4070_
	);
	LUT2 #(
		.INIT('h4)
	) name3609 (
		_w1146_,
		_w3569_,
		_w4071_
	);
	LUT2 #(
		.INIT('h4)
	) name3610 (
		_w1475_,
		_w4071_,
		_w4072_
	);
	LUT2 #(
		.INIT('h8)
	) name3611 (
		_w4070_,
		_w4072_,
		_w4073_
	);
	LUT2 #(
		.INIT('h4)
	) name3612 (
		_w1452_,
		_w3591_,
		_w4074_
	);
	LUT2 #(
		.INIT('h8)
	) name3613 (
		_w4073_,
		_w4074_,
		_w4075_
	);
	LUT2 #(
		.INIT('h1)
	) name3614 (
		_w1006_,
		_w1038_,
		_w4076_
	);
	LUT2 #(
		.INIT('h8)
	) name3615 (
		_w3595_,
		_w4076_,
		_w4077_
	);
	LUT2 #(
		.INIT('h8)
	) name3616 (
		_w4075_,
		_w4077_,
		_w4078_
	);
	LUT2 #(
		.INIT('h1)
	) name3617 (
		_w887_,
		_w4078_,
		_w4079_
	);
	LUT2 #(
		.INIT('h8)
	) name3618 (
		_w887_,
		_w4078_,
		_w4080_
	);
	LUT2 #(
		.INIT('h1)
	) name3619 (
		_w4079_,
		_w4080_,
		_w4081_
	);
	LUT2 #(
		.INIT('h1)
	) name3620 (
		_w537_,
		_w4081_,
		_w4082_
	);
	LUT2 #(
		.INIT('h2)
	) name3621 (
		_w537_,
		_w978_,
		_w4083_
	);
	LUT2 #(
		.INIT('h1)
	) name3622 (
		_w4082_,
		_w4083_,
		_w4084_
	);
	LUT2 #(
		.INIT('h2)
	) name3623 (
		_w3980_,
		_w4084_,
		_w4085_
	);
	LUT2 #(
		.INIT('h1)
	) name3624 (
		_w3981_,
		_w4085_,
		_w4086_
	);
	LUT2 #(
		.INIT('h2)
	) name3625 (
		_w1936_,
		_w4086_,
		_w4087_
	);
	LUT2 #(
		.INIT('h2)
	) name3626 (
		_w1487_,
		_w1748_,
		_w4088_
	);
	LUT2 #(
		.INIT('h8)
	) name3627 (
		_w1478_,
		_w1480_,
		_w4089_
	);
	LUT2 #(
		.INIT('h4)
	) name3628 (
		_w4088_,
		_w4089_,
		_w4090_
	);
	LUT2 #(
		.INIT('h4)
	) name3629 (
		_w1183_,
		_w1478_,
		_w4091_
	);
	LUT2 #(
		.INIT('h2)
	) name3630 (
		_w1720_,
		_w4091_,
		_w4092_
	);
	LUT2 #(
		.INIT('h4)
	) name3631 (
		_w4090_,
		_w4092_,
		_w4093_
	);
	LUT2 #(
		.INIT('h8)
	) name3632 (
		_w1301_,
		_w1377_,
		_w4094_
	);
	LUT2 #(
		.INIT('h4)
	) name3633 (
		_w4093_,
		_w4094_,
		_w4095_
	);
	LUT2 #(
		.INIT('h2)
	) name3634 (
		_w1301_,
		_w1710_,
		_w4096_
	);
	LUT2 #(
		.INIT('h1)
	) name3635 (
		_w1069_,
		_w4096_,
		_w4097_
	);
	LUT2 #(
		.INIT('h4)
	) name3636 (
		_w4095_,
		_w4097_,
		_w4098_
	);
	LUT2 #(
		.INIT('h2)
	) name3637 (
		_w1831_,
		_w4098_,
		_w4099_
	);
	LUT2 #(
		.INIT('h4)
	) name3638 (
		_w1831_,
		_w4098_,
		_w4100_
	);
	LUT2 #(
		.INIT('h1)
	) name3639 (
		_w4099_,
		_w4100_,
		_w4101_
	);
	LUT2 #(
		.INIT('h2)
	) name3640 (
		_w3980_,
		_w4101_,
		_w4102_
	);
	LUT2 #(
		.INIT('h1)
	) name3641 (
		_w3981_,
		_w4102_,
		_w4103_
	);
	LUT2 #(
		.INIT('h1)
	) name3642 (
		_w3677_,
		_w4103_,
		_w4104_
	);
	LUT2 #(
		.INIT('h1)
	) name3643 (
		_w4065_,
		_w4068_,
		_w4105_
	);
	LUT2 #(
		.INIT('h4)
	) name3644 (
		_w4062_,
		_w4105_,
		_w4106_
	);
	LUT2 #(
		.INIT('h4)
	) name3645 (
		_w4056_,
		_w4106_,
		_w4107_
	);
	LUT2 #(
		.INIT('h1)
	) name3646 (
		_w4087_,
		_w4104_,
		_w4108_
	);
	LUT2 #(
		.INIT('h8)
	) name3647 (
		_w4107_,
		_w4108_,
		_w4109_
	);
	LUT2 #(
		.INIT('h2)
	) name3648 (
		_w3450_,
		_w4109_,
		_w4110_
	);
	LUT2 #(
		.INIT('h8)
	) name3649 (
		_w941_,
		_w3448_,
		_w4111_
	);
	LUT2 #(
		.INIT('h1)
	) name3650 (
		_w4110_,
		_w4111_,
		_w4112_
	);
	LUT2 #(
		.INIT('h2)
	) name3651 (
		\P1_state_reg[0]/NET0131 ,
		_w4112_,
		_w4113_
	);
	LUT2 #(
		.INIT('h2)
	) name3652 (
		\P1_reg3_reg[28]/NET0131 ,
		\P1_state_reg[0]/NET0131 ,
		_w4114_
	);
	LUT2 #(
		.INIT('h8)
	) name3653 (
		_w941_,
		_w1953_,
		_w4115_
	);
	LUT2 #(
		.INIT('h1)
	) name3654 (
		_w4114_,
		_w4115_,
		_w4116_
	);
	LUT2 #(
		.INIT('h4)
	) name3655 (
		_w4113_,
		_w4116_,
		_w4117_
	);
	LUT2 #(
		.INIT('h4)
	) name3656 (
		_w3419_,
		_w3976_,
		_w4118_
	);
	LUT2 #(
		.INIT('h2)
	) name3657 (
		\P2_B_reg/NET0131 ,
		_w4118_,
		_w4119_
	);
	LUT2 #(
		.INIT('h1)
	) name3658 (
		\P1_datao_reg[30]/NET0131 ,
		\si[30]_pad ,
		_w4120_
	);
	LUT2 #(
		.INIT('h1)
	) name3659 (
		_w2062_,
		_w2064_,
		_w4121_
	);
	LUT2 #(
		.INIT('h4)
	) name3660 (
		_w2072_,
		_w4121_,
		_w4122_
	);
	LUT2 #(
		.INIT('h4)
	) name3661 (
		_w4120_,
		_w4122_,
		_w4123_
	);
	LUT2 #(
		.INIT('h8)
	) name3662 (
		_w2968_,
		_w4123_,
		_w4124_
	);
	LUT2 #(
		.INIT('h4)
	) name3663 (
		_w3073_,
		_w4124_,
		_w4125_
	);
	LUT2 #(
		.INIT('h4)
	) name3664 (
		_w2172_,
		_w4121_,
		_w4126_
	);
	LUT2 #(
		.INIT('h1)
	) name3665 (
		_w2061_,
		_w4126_,
		_w4127_
	);
	LUT2 #(
		.INIT('h1)
	) name3666 (
		_w4120_,
		_w4127_,
		_w4128_
	);
	LUT2 #(
		.INIT('h4)
	) name3667 (
		_w2967_,
		_w4123_,
		_w4129_
	);
	LUT2 #(
		.INIT('h8)
	) name3668 (
		\P1_datao_reg[30]/NET0131 ,
		\si[30]_pad ,
		_w4130_
	);
	LUT2 #(
		.INIT('h1)
	) name3669 (
		_w4128_,
		_w4130_,
		_w4131_
	);
	LUT2 #(
		.INIT('h4)
	) name3670 (
		_w4129_,
		_w4131_,
		_w4132_
	);
	LUT2 #(
		.INIT('h4)
	) name3671 (
		_w4125_,
		_w4132_,
		_w4133_
	);
	LUT2 #(
		.INIT('h2)
	) name3672 (
		\si[31]_pad ,
		_w4133_,
		_w4134_
	);
	LUT2 #(
		.INIT('h4)
	) name3673 (
		\si[31]_pad ,
		_w4133_,
		_w4135_
	);
	LUT2 #(
		.INIT('h2)
	) name3674 (
		_w543_,
		_w4134_,
		_w4136_
	);
	LUT2 #(
		.INIT('h4)
	) name3675 (
		_w4135_,
		_w4136_,
		_w4137_
	);
	LUT2 #(
		.INIT('h8)
	) name3676 (
		\P1_datao_reg[31]/NET0131 ,
		_w4137_,
		_w4138_
	);
	LUT2 #(
		.INIT('h1)
	) name3677 (
		\P1_datao_reg[31]/NET0131 ,
		_w4137_,
		_w4139_
	);
	LUT2 #(
		.INIT('h1)
	) name3678 (
		_w4138_,
		_w4139_,
		_w4140_
	);
	LUT2 #(
		.INIT('h4)
	) name3679 (
		_w2059_,
		_w4140_,
		_w4141_
	);
	LUT2 #(
		.INIT('h2)
	) name3680 (
		\P1_datao_reg[30]/NET0131 ,
		_w543_,
		_w4142_
	);
	LUT2 #(
		.INIT('h1)
	) name3681 (
		_w4120_,
		_w4130_,
		_w4143_
	);
	LUT2 #(
		.INIT('h4)
	) name3682 (
		_w2062_,
		_w2171_,
		_w4144_
	);
	LUT2 #(
		.INIT('h4)
	) name3683 (
		_w2073_,
		_w4122_,
		_w4145_
	);
	LUT2 #(
		.INIT('h4)
	) name3684 (
		_w2998_,
		_w4145_,
		_w4146_
	);
	LUT2 #(
		.INIT('h4)
	) name3685 (
		_w2924_,
		_w4122_,
		_w4147_
	);
	LUT2 #(
		.INIT('h8)
	) name3686 (
		_w2999_,
		_w4145_,
		_w4148_
	);
	LUT2 #(
		.INIT('h4)
	) name3687 (
		_w3096_,
		_w4148_,
		_w4149_
	);
	LUT2 #(
		.INIT('h1)
	) name3688 (
		_w2061_,
		_w4144_,
		_w4150_
	);
	LUT2 #(
		.INIT('h4)
	) name3689 (
		_w4147_,
		_w4150_,
		_w4151_
	);
	LUT2 #(
		.INIT('h4)
	) name3690 (
		_w4146_,
		_w4151_,
		_w4152_
	);
	LUT2 #(
		.INIT('h4)
	) name3691 (
		_w4149_,
		_w4152_,
		_w4153_
	);
	LUT2 #(
		.INIT('h2)
	) name3692 (
		_w4143_,
		_w4153_,
		_w4154_
	);
	LUT2 #(
		.INIT('h4)
	) name3693 (
		_w4143_,
		_w4153_,
		_w4155_
	);
	LUT2 #(
		.INIT('h2)
	) name3694 (
		_w543_,
		_w4154_,
		_w4156_
	);
	LUT2 #(
		.INIT('h4)
	) name3695 (
		_w4155_,
		_w4156_,
		_w4157_
	);
	LUT2 #(
		.INIT('h1)
	) name3696 (
		_w4142_,
		_w4157_,
		_w4158_
	);
	LUT2 #(
		.INIT('h1)
	) name3697 (
		_w2059_,
		_w4158_,
		_w4159_
	);
	LUT2 #(
		.INIT('h1)
	) name3698 (
		_w3402_,
		_w4159_,
		_w4160_
	);
	LUT2 #(
		.INIT('h1)
	) name3699 (
		_w3372_,
		_w4160_,
		_w4161_
	);
	LUT2 #(
		.INIT('h2)
	) name3700 (
		_w4141_,
		_w4161_,
		_w4162_
	);
	LUT2 #(
		.INIT('h1)
	) name3701 (
		_w2253_,
		_w3206_,
		_w4163_
	);
	LUT2 #(
		.INIT('h1)
	) name3702 (
		_w2252_,
		_w4163_,
		_w4164_
	);
	LUT2 #(
		.INIT('h1)
	) name3703 (
		_w2252_,
		_w3179_,
		_w4165_
	);
	LUT2 #(
		.INIT('h4)
	) name3704 (
		_w3838_,
		_w3841_,
		_w4166_
	);
	LUT2 #(
		.INIT('h2)
	) name3705 (
		_w3806_,
		_w4166_,
		_w4167_
	);
	LUT2 #(
		.INIT('h8)
	) name3706 (
		_w3832_,
		_w3841_,
		_w4168_
	);
	LUT2 #(
		.INIT('h2)
	) name3707 (
		_w4167_,
		_w4168_,
		_w4169_
	);
	LUT2 #(
		.INIT('h2)
	) name3708 (
		_w3799_,
		_w4169_,
		_w4170_
	);
	LUT2 #(
		.INIT('h8)
	) name3709 (
		_w3796_,
		_w4170_,
		_w4171_
	);
	LUT2 #(
		.INIT('h2)
	) name3710 (
		_w3795_,
		_w3813_,
		_w4172_
	);
	LUT2 #(
		.INIT('h2)
	) name3711 (
		_w3852_,
		_w4172_,
		_w4173_
	);
	LUT2 #(
		.INIT('h2)
	) name3712 (
		_w3792_,
		_w4173_,
		_w4174_
	);
	LUT2 #(
		.INIT('h1)
	) name3713 (
		_w3859_,
		_w4174_,
		_w4175_
	);
	LUT2 #(
		.INIT('h4)
	) name3714 (
		_w4171_,
		_w4175_,
		_w4176_
	);
	LUT2 #(
		.INIT('h2)
	) name3715 (
		_w4165_,
		_w4176_,
		_w4177_
	);
	LUT2 #(
		.INIT('h1)
	) name3716 (
		_w4164_,
		_w4177_,
		_w4178_
	);
	LUT2 #(
		.INIT('h1)
	) name3717 (
		_w3372_,
		_w4141_,
		_w4179_
	);
	LUT2 #(
		.INIT('h1)
	) name3718 (
		_w3372_,
		_w3402_,
		_w4180_
	);
	LUT2 #(
		.INIT('h2)
	) name3719 (
		_w4159_,
		_w4180_,
		_w4181_
	);
	LUT2 #(
		.INIT('h1)
	) name3720 (
		_w4179_,
		_w4181_,
		_w4182_
	);
	LUT2 #(
		.INIT('h4)
	) name3721 (
		_w4178_,
		_w4182_,
		_w4183_
	);
	LUT2 #(
		.INIT('h1)
	) name3722 (
		_w4162_,
		_w4183_,
		_w4184_
	);
	LUT2 #(
		.INIT('h4)
	) name3723 (
		_w3175_,
		_w4184_,
		_w4185_
	);
	LUT2 #(
		.INIT('h2)
	) name3724 (
		_w3175_,
		_w4184_,
		_w4186_
	);
	LUT2 #(
		.INIT('h2)
	) name3725 (
		_w3166_,
		_w3170_,
		_w4187_
	);
	LUT2 #(
		.INIT('h4)
	) name3726 (
		_w4185_,
		_w4187_,
		_w4188_
	);
	LUT2 #(
		.INIT('h4)
	) name3727 (
		_w4186_,
		_w4188_,
		_w4189_
	);
	LUT2 #(
		.INIT('h8)
	) name3728 (
		\P2_B_reg/NET0131 ,
		_w1982_,
		_w4190_
	);
	LUT2 #(
		.INIT('h1)
	) name3729 (
		_w2400_,
		_w2911_,
		_w4191_
	);
	LUT2 #(
		.INIT('h1)
	) name3730 (
		_w2894_,
		_w2900_,
		_w4192_
	);
	LUT2 #(
		.INIT('h1)
	) name3731 (
		_w3262_,
		_w3268_,
		_w4193_
	);
	LUT2 #(
		.INIT('h1)
	) name3732 (
		_w3246_,
		_w3272_,
		_w4194_
	);
	LUT2 #(
		.INIT('h1)
	) name3733 (
		_w3228_,
		_w3229_,
		_w4195_
	);
	LUT2 #(
		.INIT('h1)
	) name3734 (
		_w3089_,
		_w3144_,
		_w4196_
	);
	LUT2 #(
		.INIT('h1)
	) name3735 (
		_w2312_,
		_w2916_,
		_w4197_
	);
	LUT2 #(
		.INIT('h1)
	) name3736 (
		_w3230_,
		_w3239_,
		_w4198_
	);
	LUT2 #(
		.INIT('h1)
	) name3737 (
		_w3255_,
		_w3257_,
		_w4199_
	);
	LUT2 #(
		.INIT('h1)
	) name3738 (
		_w3066_,
		_w3143_,
		_w4200_
	);
	LUT2 #(
		.INIT('h1)
	) name3739 (
		_w2705_,
		_w2790_,
		_w4201_
	);
	LUT2 #(
		.INIT('h1)
	) name3740 (
		_w2567_,
		_w2609_,
		_w4202_
	);
	LUT2 #(
		.INIT('h4)
	) name3741 (
		_w2597_,
		_w2604_,
		_w4203_
	);
	LUT2 #(
		.INIT('h1)
	) name3742 (
		_w3258_,
		_w4203_,
		_w4204_
	);
	LUT2 #(
		.INIT('h1)
	) name3743 (
		_w2522_,
		_w2668_,
		_w4205_
	);
	LUT2 #(
		.INIT('h1)
	) name3744 (
		_w2657_,
		_w2660_,
		_w4206_
	);
	LUT2 #(
		.INIT('h1)
	) name3745 (
		_w2496_,
		_w2674_,
		_w4207_
	);
	LUT2 #(
		.INIT('h1)
	) name3746 (
		_w2471_,
		_w2673_,
		_w4208_
	);
	LUT2 #(
		.INIT('h1)
	) name3747 (
		_w3113_,
		_w3138_,
		_w4209_
	);
	LUT2 #(
		.INIT('h1)
	) name3748 (
		_w2871_,
		_w2899_,
		_w4210_
	);
	LUT2 #(
		.INIT('h1)
	) name3749 (
		_w2819_,
		_w2904_,
		_w4211_
	);
	LUT2 #(
		.INIT('h1)
	) name3750 (
		_w2732_,
		_w2789_,
		_w4212_
	);
	LUT2 #(
		.INIT('h1)
	) name3751 (
		_w3044_,
		_w3150_,
		_w4213_
	);
	LUT2 #(
		.INIT('h1)
	) name3752 (
		_w3022_,
		_w3149_,
		_w4214_
	);
	LUT2 #(
		.INIT('h1)
	) name3753 (
		_w2844_,
		_w2905_,
		_w4215_
	);
	LUT2 #(
		.INIT('h1)
	) name3754 (
		_w3131_,
		_w3139_,
		_w4216_
	);
	LUT2 #(
		.INIT('h1)
	) name3755 (
		_w2369_,
		_w2915_,
		_w4217_
	);
	LUT2 #(
		.INIT('h1)
	) name3756 (
		_w2443_,
		_w2910_,
		_w4218_
	);
	LUT2 #(
		.INIT('h1)
	) name3757 (
		_w2992_,
		_w3136_,
		_w4219_
	);
	LUT2 #(
		.INIT('h8)
	) name3758 (
		_w3402_,
		_w4159_,
		_w4220_
	);
	LUT2 #(
		.INIT('h1)
	) name3759 (
		_w4179_,
		_w4220_,
		_w4221_
	);
	LUT2 #(
		.INIT('h8)
	) name3760 (
		_w3372_,
		_w4141_,
		_w4222_
	);
	LUT2 #(
		.INIT('h1)
	) name3761 (
		_w4160_,
		_w4222_,
		_w4223_
	);
	LUT2 #(
		.INIT('h8)
	) name3762 (
		_w4193_,
		_w4194_,
		_w4224_
	);
	LUT2 #(
		.INIT('h2)
	) name3763 (
		_w4199_,
		_w4202_,
		_w4225_
	);
	LUT2 #(
		.INIT('h2)
	) name3764 (
		_w4204_,
		_w4205_,
		_w4226_
	);
	LUT2 #(
		.INIT('h4)
	) name3765 (
		_w4206_,
		_w4226_,
		_w4227_
	);
	LUT2 #(
		.INIT('h8)
	) name3766 (
		_w4224_,
		_w4225_,
		_w4228_
	);
	LUT2 #(
		.INIT('h1)
	) name3767 (
		_w4207_,
		_w4208_,
		_w4229_
	);
	LUT2 #(
		.INIT('h8)
	) name3768 (
		_w4228_,
		_w4229_,
		_w4230_
	);
	LUT2 #(
		.INIT('h8)
	) name3769 (
		_w4195_,
		_w4227_,
		_w4231_
	);
	LUT2 #(
		.INIT('h8)
	) name3770 (
		_w4198_,
		_w4231_,
		_w4232_
	);
	LUT2 #(
		.INIT('h4)
	) name3771 (
		_w4201_,
		_w4230_,
		_w4233_
	);
	LUT2 #(
		.INIT('h4)
	) name3772 (
		_w4212_,
		_w4233_,
		_w4234_
	);
	LUT2 #(
		.INIT('h4)
	) name3773 (
		_w4192_,
		_w4232_,
		_w4235_
	);
	LUT2 #(
		.INIT('h1)
	) name3774 (
		_w4210_,
		_w4211_,
		_w4236_
	);
	LUT2 #(
		.INIT('h8)
	) name3775 (
		_w4235_,
		_w4236_,
		_w4237_
	);
	LUT2 #(
		.INIT('h4)
	) name3776 (
		_w4191_,
		_w4234_,
		_w4238_
	);
	LUT2 #(
		.INIT('h1)
	) name3777 (
		_w4215_,
		_w4216_,
		_w4239_
	);
	LUT2 #(
		.INIT('h1)
	) name3778 (
		_w4217_,
		_w4218_,
		_w4240_
	);
	LUT2 #(
		.INIT('h8)
	) name3779 (
		_w4239_,
		_w4240_,
		_w4241_
	);
	LUT2 #(
		.INIT('h8)
	) name3780 (
		_w4237_,
		_w4238_,
		_w4242_
	);
	LUT2 #(
		.INIT('h1)
	) name3781 (
		_w4196_,
		_w4197_,
		_w4243_
	);
	LUT2 #(
		.INIT('h8)
	) name3782 (
		_w4242_,
		_w4243_,
		_w4244_
	);
	LUT2 #(
		.INIT('h4)
	) name3783 (
		_w4200_,
		_w4241_,
		_w4245_
	);
	LUT2 #(
		.INIT('h4)
	) name3784 (
		_w4209_,
		_w4245_,
		_w4246_
	);
	LUT2 #(
		.INIT('h8)
	) name3785 (
		_w2254_,
		_w4244_,
		_w4247_
	);
	LUT2 #(
		.INIT('h1)
	) name3786 (
		_w4213_,
		_w4214_,
		_w4248_
	);
	LUT2 #(
		.INIT('h8)
	) name3787 (
		_w4247_,
		_w4248_,
		_w4249_
	);
	LUT2 #(
		.INIT('h4)
	) name3788 (
		_w3862_,
		_w4246_,
		_w4250_
	);
	LUT2 #(
		.INIT('h4)
	) name3789 (
		_w4219_,
		_w4221_,
		_w4251_
	);
	LUT2 #(
		.INIT('h8)
	) name3790 (
		_w4223_,
		_w4251_,
		_w4252_
	);
	LUT2 #(
		.INIT('h8)
	) name3791 (
		_w4249_,
		_w4250_,
		_w4253_
	);
	LUT2 #(
		.INIT('h8)
	) name3792 (
		_w4252_,
		_w4253_,
		_w4254_
	);
	LUT2 #(
		.INIT('h4)
	) name3793 (
		_w3175_,
		_w4254_,
		_w4255_
	);
	LUT2 #(
		.INIT('h2)
	) name3794 (
		_w3175_,
		_w4254_,
		_w4256_
	);
	LUT2 #(
		.INIT('h1)
	) name3795 (
		_w3166_,
		_w4255_,
		_w4257_
	);
	LUT2 #(
		.INIT('h4)
	) name3796 (
		_w4256_,
		_w4257_,
		_w4258_
	);
	LUT2 #(
		.INIT('h1)
	) name3797 (
		_w4190_,
		_w4258_,
		_w4259_
	);
	LUT2 #(
		.INIT('h1)
	) name3798 (
		_w3170_,
		_w4259_,
		_w4260_
	);
	LUT2 #(
		.INIT('h1)
	) name3799 (
		_w2253_,
		_w4160_,
		_w4261_
	);
	LUT2 #(
		.INIT('h4)
	) name3800 (
		_w4165_,
		_w4261_,
		_w4262_
	);
	LUT2 #(
		.INIT('h2)
	) name3801 (
		_w4221_,
		_w4262_,
		_w4263_
	);
	LUT2 #(
		.INIT('h1)
	) name3802 (
		_w4222_,
		_w4263_,
		_w4264_
	);
	LUT2 #(
		.INIT('h8)
	) name3803 (
		_w4163_,
		_w4223_,
		_w4265_
	);
	LUT2 #(
		.INIT('h8)
	) name3804 (
		_w3854_,
		_w3855_,
		_w4266_
	);
	LUT2 #(
		.INIT('h8)
	) name3805 (
		_w4265_,
		_w4266_,
		_w4267_
	);
	LUT2 #(
		.INIT('h8)
	) name3806 (
		_w3816_,
		_w3841_,
		_w4268_
	);
	LUT2 #(
		.INIT('h2)
	) name3807 (
		_w4167_,
		_w4268_,
		_w4269_
	);
	LUT2 #(
		.INIT('h4)
	) name3808 (
		_w3257_,
		_w4203_,
		_w4270_
	);
	LUT2 #(
		.INIT('h2)
	) name3809 (
		_w3256_,
		_w4270_,
		_w4271_
	);
	LUT2 #(
		.INIT('h2)
	) name3810 (
		_w3263_,
		_w4271_,
		_w4272_
	);
	LUT2 #(
		.INIT('h2)
	) name3811 (
		_w3269_,
		_w4272_,
		_w4273_
	);
	LUT2 #(
		.INIT('h2)
	) name3812 (
		_w3818_,
		_w4273_,
		_w4274_
	);
	LUT2 #(
		.INIT('h2)
	) name3813 (
		_w3247_,
		_w4274_,
		_w4275_
	);
	LUT2 #(
		.INIT('h2)
	) name3814 (
		_w3817_,
		_w4275_,
		_w4276_
	);
	LUT2 #(
		.INIT('h4)
	) name3815 (
		_w3251_,
		_w3833_,
		_w4277_
	);
	LUT2 #(
		.INIT('h8)
	) name3816 (
		_w3836_,
		_w4277_,
		_w4278_
	);
	LUT2 #(
		.INIT('h8)
	) name3817 (
		_w3801_,
		_w4278_,
		_w4279_
	);
	LUT2 #(
		.INIT('h8)
	) name3818 (
		_w3804_,
		_w4279_,
		_w4280_
	);
	LUT2 #(
		.INIT('h4)
	) name3819 (
		_w4276_,
		_w4280_,
		_w4281_
	);
	LUT2 #(
		.INIT('h1)
	) name3820 (
		_w4269_,
		_w4281_,
		_w4282_
	);
	LUT2 #(
		.INIT('h4)
	) name3821 (
		_w3191_,
		_w3300_,
		_w4283_
	);
	LUT2 #(
		.INIT('h8)
	) name3822 (
		_w3850_,
		_w4283_,
		_w4284_
	);
	LUT2 #(
		.INIT('h4)
	) name3823 (
		_w3287_,
		_w3295_,
		_w4285_
	);
	LUT2 #(
		.INIT('h8)
	) name3824 (
		_w4284_,
		_w4285_,
		_w4286_
	);
	LUT2 #(
		.INIT('h4)
	) name3825 (
		_w4282_,
		_w4286_,
		_w4287_
	);
	LUT2 #(
		.INIT('h8)
	) name3826 (
		_w4267_,
		_w4287_,
		_w4288_
	);
	LUT2 #(
		.INIT('h2)
	) name3827 (
		_w3192_,
		_w3794_,
		_w4289_
	);
	LUT2 #(
		.INIT('h2)
	) name3828 (
		_w3793_,
		_w4289_,
		_w4290_
	);
	LUT2 #(
		.INIT('h1)
	) name3829 (
		_w3196_,
		_w4290_,
		_w4291_
	);
	LUT2 #(
		.INIT('h2)
	) name3830 (
		_w3295_,
		_w3798_,
		_w4292_
	);
	LUT2 #(
		.INIT('h2)
	) name3831 (
		_w3797_,
		_w4292_,
		_w4293_
	);
	LUT2 #(
		.INIT('h2)
	) name3832 (
		_w4284_,
		_w4293_,
		_w4294_
	);
	LUT2 #(
		.INIT('h1)
	) name3833 (
		_w4291_,
		_w4294_,
		_w4295_
	);
	LUT2 #(
		.INIT('h2)
	) name3834 (
		_w4267_,
		_w4295_,
		_w4296_
	);
	LUT2 #(
		.INIT('h2)
	) name3835 (
		_w3203_,
		_w3790_,
		_w4297_
	);
	LUT2 #(
		.INIT('h2)
	) name3836 (
		_w3791_,
		_w4297_,
		_w4298_
	);
	LUT2 #(
		.INIT('h4)
	) name3837 (
		_w3207_,
		_w4265_,
		_w4299_
	);
	LUT2 #(
		.INIT('h4)
	) name3838 (
		_w4298_,
		_w4299_,
		_w4300_
	);
	LUT2 #(
		.INIT('h1)
	) name3839 (
		_w4264_,
		_w4288_,
		_w4301_
	);
	LUT2 #(
		.INIT('h1)
	) name3840 (
		_w4296_,
		_w4300_,
		_w4302_
	);
	LUT2 #(
		.INIT('h8)
	) name3841 (
		_w4301_,
		_w4302_,
		_w4303_
	);
	LUT2 #(
		.INIT('h1)
	) name3842 (
		\P2_B_reg/NET0131 ,
		_w4303_,
		_w4304_
	);
	LUT2 #(
		.INIT('h8)
	) name3843 (
		_w3410_,
		_w3418_,
		_w4305_
	);
	LUT2 #(
		.INIT('h4)
	) name3844 (
		_w4304_,
		_w4305_,
		_w4306_
	);
	LUT2 #(
		.INIT('h2)
	) name3845 (
		_w3411_,
		_w4303_,
		_w4307_
	);
	LUT2 #(
		.INIT('h1)
	) name3846 (
		_w3176_,
		_w3411_,
		_w4308_
	);
	LUT2 #(
		.INIT('h2)
	) name3847 (
		\P2_B_reg/NET0131 ,
		_w4308_,
		_w4309_
	);
	LUT2 #(
		.INIT('h1)
	) name3848 (
		_w3175_,
		_w4303_,
		_w4310_
	);
	LUT2 #(
		.INIT('h8)
	) name3849 (
		_w3175_,
		_w4303_,
		_w4311_
	);
	LUT2 #(
		.INIT('h2)
	) name3850 (
		_w3171_,
		_w4310_,
		_w4312_
	);
	LUT2 #(
		.INIT('h4)
	) name3851 (
		_w4311_,
		_w4312_,
		_w4313_
	);
	LUT2 #(
		.INIT('h1)
	) name3852 (
		_w4264_,
		_w4265_,
		_w4314_
	);
	LUT2 #(
		.INIT('h8)
	) name3853 (
		_w4177_,
		_w4221_,
		_w4315_
	);
	LUT2 #(
		.INIT('h1)
	) name3854 (
		_w4314_,
		_w4315_,
		_w4316_
	);
	LUT2 #(
		.INIT('h8)
	) name3855 (
		_w3354_,
		_w4316_,
		_w4317_
	);
	LUT2 #(
		.INIT('h2)
	) name3856 (
		_w3419_,
		_w4316_,
		_w4318_
	);
	LUT2 #(
		.INIT('h1)
	) name3857 (
		_w4307_,
		_w4309_,
		_w4319_
	);
	LUT2 #(
		.INIT('h4)
	) name3858 (
		_w4306_,
		_w4319_,
		_w4320_
	);
	LUT2 #(
		.INIT('h4)
	) name3859 (
		_w4260_,
		_w4320_,
		_w4321_
	);
	LUT2 #(
		.INIT('h4)
	) name3860 (
		_w4313_,
		_w4321_,
		_w4322_
	);
	LUT2 #(
		.INIT('h1)
	) name3861 (
		_w4317_,
		_w4318_,
		_w4323_
	);
	LUT2 #(
		.INIT('h8)
	) name3862 (
		_w4322_,
		_w4323_,
		_w4324_
	);
	LUT2 #(
		.INIT('h4)
	) name3863 (
		_w4189_,
		_w4324_,
		_w4325_
	);
	LUT2 #(
		.INIT('h2)
	) name3864 (
		_w3976_,
		_w4325_,
		_w4326_
	);
	LUT2 #(
		.INIT('h1)
	) name3865 (
		_w4119_,
		_w4326_,
		_w4327_
	);
	LUT2 #(
		.INIT('h2)
	) name3866 (
		\P2_reg0_reg[28]/NET0131 ,
		_w1983_,
		_w4328_
	);
	LUT2 #(
		.INIT('h8)
	) name3867 (
		\P2_reg0_reg[28]/NET0131 ,
		_w2024_,
		_w4329_
	);
	LUT2 #(
		.INIT('h2)
	) name3868 (
		\P2_reg0_reg[28]/NET0131 ,
		_w2040_,
		_w4330_
	);
	LUT2 #(
		.INIT('h2)
	) name3869 (
		_w2040_,
		_w3865_,
		_w4331_
	);
	LUT2 #(
		.INIT('h1)
	) name3870 (
		_w4330_,
		_w4331_,
		_w4332_
	);
	LUT2 #(
		.INIT('h1)
	) name3871 (
		_w3320_,
		_w4332_,
		_w4333_
	);
	LUT2 #(
		.INIT('h2)
	) name3872 (
		_w2040_,
		_w3942_,
		_w4334_
	);
	LUT2 #(
		.INIT('h1)
	) name3873 (
		_w4330_,
		_w4334_,
		_w4335_
	);
	LUT2 #(
		.INIT('h1)
	) name3874 (
		_w3177_,
		_w4335_,
		_w4336_
	);
	LUT2 #(
		.INIT('h8)
	) name3875 (
		_w3355_,
		_w3948_,
		_w4337_
	);
	LUT2 #(
		.INIT('h8)
	) name3876 (
		_w2949_,
		_w3358_,
		_w4338_
	);
	LUT2 #(
		.INIT('h8)
	) name3877 (
		_w3411_,
		_w3957_,
		_w4339_
	);
	LUT2 #(
		.INIT('h1)
	) name3878 (
		_w4338_,
		_w4339_,
		_w4340_
	);
	LUT2 #(
		.INIT('h4)
	) name3879 (
		_w4337_,
		_w4340_,
		_w4341_
	);
	LUT2 #(
		.INIT('h2)
	) name3880 (
		_w2040_,
		_w4341_,
		_w4342_
	);
	LUT2 #(
		.INIT('h2)
	) name3881 (
		\P2_reg0_reg[28]/NET0131 ,
		_w3426_,
		_w4343_
	);
	LUT2 #(
		.INIT('h1)
	) name3882 (
		_w4342_,
		_w4343_,
		_w4344_
	);
	LUT2 #(
		.INIT('h4)
	) name3883 (
		_w4336_,
		_w4344_,
		_w4345_
	);
	LUT2 #(
		.INIT('h4)
	) name3884 (
		_w4333_,
		_w4345_,
		_w4346_
	);
	LUT2 #(
		.INIT('h2)
	) name3885 (
		_w2026_,
		_w4346_,
		_w4347_
	);
	LUT2 #(
		.INIT('h1)
	) name3886 (
		_w4329_,
		_w4347_,
		_w4348_
	);
	LUT2 #(
		.INIT('h2)
	) name3887 (
		\P1_state_reg[0]/NET0131 ,
		_w4348_,
		_w4349_
	);
	LUT2 #(
		.INIT('h1)
	) name3888 (
		_w4328_,
		_w4349_,
		_w4350_
	);
	LUT2 #(
		.INIT('h2)
	) name3889 (
		\P2_reg1_reg[28]/NET0131 ,
		_w1983_,
		_w4351_
	);
	LUT2 #(
		.INIT('h8)
	) name3890 (
		\P2_reg1_reg[28]/NET0131 ,
		_w2024_,
		_w4352_
	);
	LUT2 #(
		.INIT('h2)
	) name3891 (
		\P2_reg1_reg[28]/NET0131 ,
		_w3733_,
		_w4353_
	);
	LUT2 #(
		.INIT('h2)
	) name3892 (
		_w3733_,
		_w3865_,
		_w4354_
	);
	LUT2 #(
		.INIT('h1)
	) name3893 (
		_w4353_,
		_w4354_,
		_w4355_
	);
	LUT2 #(
		.INIT('h1)
	) name3894 (
		_w3320_,
		_w4355_,
		_w4356_
	);
	LUT2 #(
		.INIT('h2)
	) name3895 (
		_w3733_,
		_w3942_,
		_w4357_
	);
	LUT2 #(
		.INIT('h1)
	) name3896 (
		_w4353_,
		_w4357_,
		_w4358_
	);
	LUT2 #(
		.INIT('h1)
	) name3897 (
		_w3177_,
		_w4358_,
		_w4359_
	);
	LUT2 #(
		.INIT('h2)
	) name3898 (
		_w3733_,
		_w4341_,
		_w4360_
	);
	LUT2 #(
		.INIT('h2)
	) name3899 (
		\P2_reg1_reg[28]/NET0131 ,
		_w3747_,
		_w4361_
	);
	LUT2 #(
		.INIT('h1)
	) name3900 (
		_w4360_,
		_w4361_,
		_w4362_
	);
	LUT2 #(
		.INIT('h4)
	) name3901 (
		_w4359_,
		_w4362_,
		_w4363_
	);
	LUT2 #(
		.INIT('h4)
	) name3902 (
		_w4356_,
		_w4363_,
		_w4364_
	);
	LUT2 #(
		.INIT('h2)
	) name3903 (
		_w2026_,
		_w4364_,
		_w4365_
	);
	LUT2 #(
		.INIT('h1)
	) name3904 (
		_w4352_,
		_w4365_,
		_w4366_
	);
	LUT2 #(
		.INIT('h2)
	) name3905 (
		\P1_state_reg[0]/NET0131 ,
		_w4366_,
		_w4367_
	);
	LUT2 #(
		.INIT('h1)
	) name3906 (
		_w4351_,
		_w4367_,
		_w4368_
	);
	LUT2 #(
		.INIT('h2)
	) name3907 (
		\P2_reg2_reg[28]/NET0131 ,
		_w1983_,
		_w4369_
	);
	LUT2 #(
		.INIT('h8)
	) name3908 (
		\P2_reg2_reg[28]/NET0131 ,
		_w2024_,
		_w4370_
	);
	LUT2 #(
		.INIT('h2)
	) name3909 (
		\P2_reg2_reg[28]/NET0131 ,
		_w3758_,
		_w4371_
	);
	LUT2 #(
		.INIT('h2)
	) name3910 (
		_w3758_,
		_w3865_,
		_w4372_
	);
	LUT2 #(
		.INIT('h1)
	) name3911 (
		_w4371_,
		_w4372_,
		_w4373_
	);
	LUT2 #(
		.INIT('h1)
	) name3912 (
		_w3320_,
		_w4373_,
		_w4374_
	);
	LUT2 #(
		.INIT('h2)
	) name3913 (
		_w3758_,
		_w3942_,
		_w4375_
	);
	LUT2 #(
		.INIT('h1)
	) name3914 (
		_w4371_,
		_w4375_,
		_w4376_
	);
	LUT2 #(
		.INIT('h1)
	) name3915 (
		_w3177_,
		_w4376_,
		_w4377_
	);
	LUT2 #(
		.INIT('h2)
	) name3916 (
		_w3758_,
		_w4341_,
		_w4378_
	);
	LUT2 #(
		.INIT('h4)
	) name3917 (
		_w2958_,
		_w3420_,
		_w4379_
	);
	LUT2 #(
		.INIT('h2)
	) name3918 (
		_w3411_,
		_w3758_,
		_w4380_
	);
	LUT2 #(
		.INIT('h2)
	) name3919 (
		_w3354_,
		_w3758_,
		_w4381_
	);
	LUT2 #(
		.INIT('h4)
	) name3920 (
		_w1982_,
		_w4381_,
		_w4382_
	);
	LUT2 #(
		.INIT('h2)
	) name3921 (
		_w3774_,
		_w4382_,
		_w4383_
	);
	LUT2 #(
		.INIT('h4)
	) name3922 (
		_w4380_,
		_w4383_,
		_w4384_
	);
	LUT2 #(
		.INIT('h2)
	) name3923 (
		\P2_reg2_reg[28]/NET0131 ,
		_w4384_,
		_w4385_
	);
	LUT2 #(
		.INIT('h1)
	) name3924 (
		_w4379_,
		_w4385_,
		_w4386_
	);
	LUT2 #(
		.INIT('h4)
	) name3925 (
		_w4378_,
		_w4386_,
		_w4387_
	);
	LUT2 #(
		.INIT('h4)
	) name3926 (
		_w4377_,
		_w4387_,
		_w4388_
	);
	LUT2 #(
		.INIT('h4)
	) name3927 (
		_w4374_,
		_w4388_,
		_w4389_
	);
	LUT2 #(
		.INIT('h2)
	) name3928 (
		_w2026_,
		_w4389_,
		_w4390_
	);
	LUT2 #(
		.INIT('h1)
	) name3929 (
		_w4370_,
		_w4390_,
		_w4391_
	);
	LUT2 #(
		.INIT('h2)
	) name3930 (
		\P1_state_reg[0]/NET0131 ,
		_w4391_,
		_w4392_
	);
	LUT2 #(
		.INIT('h1)
	) name3931 (
		_w4369_,
		_w4392_,
		_w4393_
	);
	LUT2 #(
		.INIT('h2)
	) name3932 (
		\P1_reg0_reg[27]/NET0131 ,
		_w3435_,
		_w4394_
	);
	LUT2 #(
		.INIT('h8)
	) name3933 (
		\P1_reg0_reg[27]/NET0131 ,
		_w3448_,
		_w4395_
	);
	LUT2 #(
		.INIT('h8)
	) name3934 (
		_w3460_,
		_w3465_,
		_w4396_
	);
	LUT2 #(
		.INIT('h2)
	) name3935 (
		\P1_reg0_reg[27]/NET0131 ,
		_w4396_,
		_w4397_
	);
	LUT2 #(
		.INIT('h8)
	) name3936 (
		_w3636_,
		_w3637_,
		_w4398_
	);
	LUT2 #(
		.INIT('h1)
	) name3937 (
		_w3641_,
		_w4398_,
		_w4399_
	);
	LUT2 #(
		.INIT('h8)
	) name3938 (
		_w3638_,
		_w3647_,
		_w4400_
	);
	LUT2 #(
		.INIT('h4)
	) name3939 (
		_w4399_,
		_w4400_,
		_w4401_
	);
	LUT2 #(
		.INIT('h8)
	) name3940 (
		_w3644_,
		_w3647_,
		_w4402_
	);
	LUT2 #(
		.INIT('h1)
	) name3941 (
		_w3628_,
		_w4402_,
		_w4403_
	);
	LUT2 #(
		.INIT('h4)
	) name3942 (
		_w4401_,
		_w4403_,
		_w4404_
	);
	LUT2 #(
		.INIT('h8)
	) name3943 (
		_w3621_,
		_w3623_,
		_w4405_
	);
	LUT2 #(
		.INIT('h8)
	) name3944 (
		_w3624_,
		_w3627_,
		_w4406_
	);
	LUT2 #(
		.INIT('h8)
	) name3945 (
		_w4405_,
		_w4406_,
		_w4407_
	);
	LUT2 #(
		.INIT('h4)
	) name3946 (
		_w4404_,
		_w4407_,
		_w4408_
	);
	LUT2 #(
		.INIT('h8)
	) name3947 (
		_w3624_,
		_w3631_,
		_w4409_
	);
	LUT2 #(
		.INIT('h1)
	) name3948 (
		_w3652_,
		_w4409_,
		_w4410_
	);
	LUT2 #(
		.INIT('h2)
	) name3949 (
		_w4405_,
		_w4410_,
		_w4411_
	);
	LUT2 #(
		.INIT('h8)
	) name3950 (
		_w3621_,
		_w3655_,
		_w4412_
	);
	LUT2 #(
		.INIT('h1)
	) name3951 (
		_w3658_,
		_w4412_,
		_w4413_
	);
	LUT2 #(
		.INIT('h4)
	) name3952 (
		_w4411_,
		_w4413_,
		_w4414_
	);
	LUT2 #(
		.INIT('h4)
	) name3953 (
		_w4408_,
		_w4414_,
		_w4415_
	);
	LUT2 #(
		.INIT('h8)
	) name3954 (
		_w3606_,
		_w3612_,
		_w4416_
	);
	LUT2 #(
		.INIT('h8)
	) name3955 (
		_w3620_,
		_w3665_,
		_w4417_
	);
	LUT2 #(
		.INIT('h8)
	) name3956 (
		_w4416_,
		_w4417_,
		_w4418_
	);
	LUT2 #(
		.INIT('h4)
	) name3957 (
		_w4415_,
		_w4418_,
		_w4419_
	);
	LUT2 #(
		.INIT('h8)
	) name3958 (
		_w3610_,
		_w3612_,
		_w4420_
	);
	LUT2 #(
		.INIT('h4)
	) name3959 (
		_w3661_,
		_w3665_,
		_w4421_
	);
	LUT2 #(
		.INIT('h1)
	) name3960 (
		_w3607_,
		_w4421_,
		_w4422_
	);
	LUT2 #(
		.INIT('h2)
	) name3961 (
		_w4416_,
		_w4422_,
		_w4423_
	);
	LUT2 #(
		.INIT('h1)
	) name3962 (
		_w3615_,
		_w4420_,
		_w4424_
	);
	LUT2 #(
		.INIT('h4)
	) name3963 (
		_w4423_,
		_w4424_,
		_w4425_
	);
	LUT2 #(
		.INIT('h4)
	) name3964 (
		_w4419_,
		_w4425_,
		_w4426_
	);
	LUT2 #(
		.INIT('h2)
	) name3965 (
		_w1769_,
		_w4426_,
		_w4427_
	);
	LUT2 #(
		.INIT('h4)
	) name3966 (
		_w1769_,
		_w4426_,
		_w4428_
	);
	LUT2 #(
		.INIT('h1)
	) name3967 (
		_w4427_,
		_w4428_,
		_w4429_
	);
	LUT2 #(
		.INIT('h2)
	) name3968 (
		_w4396_,
		_w4429_,
		_w4430_
	);
	LUT2 #(
		.INIT('h1)
	) name3969 (
		_w4397_,
		_w4430_,
		_w4431_
	);
	LUT2 #(
		.INIT('h1)
	) name3970 (
		_w3677_,
		_w4431_,
		_w4432_
	);
	LUT2 #(
		.INIT('h4)
	) name3971 (
		_w1810_,
		_w3468_,
		_w4433_
	);
	LUT2 #(
		.INIT('h4)
	) name3972 (
		_w3547_,
		_w3551_,
		_w4434_
	);
	LUT2 #(
		.INIT('h2)
	) name3973 (
		_w3470_,
		_w4434_,
		_w4435_
	);
	LUT2 #(
		.INIT('h2)
	) name3974 (
		_w4433_,
		_w4435_,
		_w4436_
	);
	LUT2 #(
		.INIT('h1)
	) name3975 (
		_w1810_,
		_w3473_,
		_w4437_
	);
	LUT2 #(
		.INIT('h2)
	) name3976 (
		_w3478_,
		_w4437_,
		_w4438_
	);
	LUT2 #(
		.INIT('h4)
	) name3977 (
		_w4436_,
		_w4438_,
		_w4439_
	);
	LUT2 #(
		.INIT('h1)
	) name3978 (
		_w1808_,
		_w4439_,
		_w4440_
	);
	LUT2 #(
		.INIT('h2)
	) name3979 (
		_w3501_,
		_w3518_,
		_w4441_
	);
	LUT2 #(
		.INIT('h2)
	) name3980 (
		_w3524_,
		_w4441_,
		_w4442_
	);
	LUT2 #(
		.INIT('h8)
	) name3981 (
		_w3502_,
		_w3530_,
		_w4443_
	);
	LUT2 #(
		.INIT('h4)
	) name3982 (
		_w4442_,
		_w4443_,
		_w4444_
	);
	LUT2 #(
		.INIT('h4)
	) name3983 (
		_w3527_,
		_w3530_,
		_w4445_
	);
	LUT2 #(
		.INIT('h2)
	) name3984 (
		_w3494_,
		_w4445_,
		_w4446_
	);
	LUT2 #(
		.INIT('h4)
	) name3985 (
		_w4444_,
		_w4446_,
		_w4447_
	);
	LUT2 #(
		.INIT('h8)
	) name3986 (
		_w3488_,
		_w3492_,
		_w4448_
	);
	LUT2 #(
		.INIT('h8)
	) name3987 (
		_w3486_,
		_w3489_,
		_w4449_
	);
	LUT2 #(
		.INIT('h8)
	) name3988 (
		_w4448_,
		_w4449_,
		_w4450_
	);
	LUT2 #(
		.INIT('h4)
	) name3989 (
		_w4447_,
		_w4450_,
		_w4451_
	);
	LUT2 #(
		.INIT('h2)
	) name3990 (
		_w3488_,
		_w3497_,
		_w4452_
	);
	LUT2 #(
		.INIT('h2)
	) name3991 (
		_w3536_,
		_w4452_,
		_w4453_
	);
	LUT2 #(
		.INIT('h2)
	) name3992 (
		_w4449_,
		_w4453_,
		_w4454_
	);
	LUT2 #(
		.INIT('h8)
	) name3993 (
		_w3486_,
		_w3539_,
		_w4455_
	);
	LUT2 #(
		.INIT('h2)
	) name3994 (
		_w3544_,
		_w4455_,
		_w4456_
	);
	LUT2 #(
		.INIT('h4)
	) name3995 (
		_w4454_,
		_w4456_,
		_w4457_
	);
	LUT2 #(
		.INIT('h4)
	) name3996 (
		_w4451_,
		_w4457_,
		_w4458_
	);
	LUT2 #(
		.INIT('h8)
	) name3997 (
		_w3484_,
		_w3551_,
		_w4459_
	);
	LUT2 #(
		.INIT('h4)
	) name3998 (
		_w1808_,
		_w4459_,
		_w4460_
	);
	LUT2 #(
		.INIT('h8)
	) name3999 (
		_w4433_,
		_w4460_,
		_w4461_
	);
	LUT2 #(
		.INIT('h4)
	) name4000 (
		_w4458_,
		_w4461_,
		_w4462_
	);
	LUT2 #(
		.INIT('h1)
	) name4001 (
		_w4440_,
		_w4462_,
		_w4463_
	);
	LUT2 #(
		.INIT('h8)
	) name4002 (
		_w1769_,
		_w4463_,
		_w4464_
	);
	LUT2 #(
		.INIT('h1)
	) name4003 (
		_w1769_,
		_w4463_,
		_w4465_
	);
	LUT2 #(
		.INIT('h1)
	) name4004 (
		_w4464_,
		_w4465_,
		_w4466_
	);
	LUT2 #(
		.INIT('h2)
	) name4005 (
		_w4396_,
		_w4466_,
		_w4467_
	);
	LUT2 #(
		.INIT('h1)
	) name4006 (
		_w4397_,
		_w4467_,
		_w4468_
	);
	LUT2 #(
		.INIT('h1)
	) name4007 (
		_w3563_,
		_w4468_,
		_w4469_
	);
	LUT2 #(
		.INIT('h8)
	) name4008 (
		_w4070_,
		_w4071_,
		_w4470_
	);
	LUT2 #(
		.INIT('h8)
	) name4009 (
		_w3568_,
		_w3590_,
		_w4471_
	);
	LUT2 #(
		.INIT('h8)
	) name4010 (
		_w4470_,
		_w4471_,
		_w4472_
	);
	LUT2 #(
		.INIT('h4)
	) name4011 (
		_w1062_,
		_w4076_,
		_w4473_
	);
	LUT2 #(
		.INIT('h4)
	) name4012 (
		_w978_,
		_w4473_,
		_w4474_
	);
	LUT2 #(
		.INIT('h8)
	) name4013 (
		_w4472_,
		_w4474_,
		_w4475_
	);
	LUT2 #(
		.INIT('h2)
	) name4014 (
		_w945_,
		_w4475_,
		_w4476_
	);
	LUT2 #(
		.INIT('h1)
	) name4015 (
		_w4078_,
		_w4476_,
		_w4477_
	);
	LUT2 #(
		.INIT('h1)
	) name4016 (
		_w537_,
		_w4477_,
		_w4478_
	);
	LUT2 #(
		.INIT('h8)
	) name4017 (
		_w537_,
		_w1006_,
		_w4479_
	);
	LUT2 #(
		.INIT('h1)
	) name4018 (
		_w4478_,
		_w4479_,
		_w4480_
	);
	LUT2 #(
		.INIT('h8)
	) name4019 (
		_w4396_,
		_w4480_,
		_w4481_
	);
	LUT2 #(
		.INIT('h1)
	) name4020 (
		_w4397_,
		_w4481_,
		_w4482_
	);
	LUT2 #(
		.INIT('h2)
	) name4021 (
		_w1936_,
		_w4482_,
		_w4483_
	);
	LUT2 #(
		.INIT('h2)
	) name4022 (
		_w969_,
		_w3704_,
		_w4484_
	);
	LUT2 #(
		.INIT('h1)
	) name4023 (
		_w4057_,
		_w4484_,
		_w4485_
	);
	LUT2 #(
		.INIT('h8)
	) name4024 (
		_w3712_,
		_w4485_,
		_w4486_
	);
	LUT2 #(
		.INIT('h8)
	) name4025 (
		_w969_,
		_w1880_,
		_w4487_
	);
	LUT2 #(
		.INIT('h1)
	) name4026 (
		_w4486_,
		_w4487_,
		_w4488_
	);
	LUT2 #(
		.INIT('h2)
	) name4027 (
		_w4396_,
		_w4488_,
		_w4489_
	);
	LUT2 #(
		.INIT('h2)
	) name4028 (
		_w3712_,
		_w4396_,
		_w4490_
	);
	LUT2 #(
		.INIT('h1)
	) name4029 (
		_w1763_,
		_w3716_,
		_w4491_
	);
	LUT2 #(
		.INIT('h2)
	) name4030 (
		_w1880_,
		_w4396_,
		_w4492_
	);
	LUT2 #(
		.INIT('h2)
	) name4031 (
		_w4491_,
		_w4492_,
		_w4493_
	);
	LUT2 #(
		.INIT('h4)
	) name4032 (
		_w4490_,
		_w4493_,
		_w4494_
	);
	LUT2 #(
		.INIT('h2)
	) name4033 (
		\P1_reg0_reg[27]/NET0131 ,
		_w4494_,
		_w4495_
	);
	LUT2 #(
		.INIT('h1)
	) name4034 (
		_w4489_,
		_w4495_,
		_w4496_
	);
	LUT2 #(
		.INIT('h4)
	) name4035 (
		_w4432_,
		_w4496_,
		_w4497_
	);
	LUT2 #(
		.INIT('h1)
	) name4036 (
		_w4469_,
		_w4483_,
		_w4498_
	);
	LUT2 #(
		.INIT('h8)
	) name4037 (
		_w4497_,
		_w4498_,
		_w4499_
	);
	LUT2 #(
		.INIT('h2)
	) name4038 (
		_w3450_,
		_w4499_,
		_w4500_
	);
	LUT2 #(
		.INIT('h1)
	) name4039 (
		_w4395_,
		_w4500_,
		_w4501_
	);
	LUT2 #(
		.INIT('h2)
	) name4040 (
		\P1_state_reg[0]/NET0131 ,
		_w4501_,
		_w4502_
	);
	LUT2 #(
		.INIT('h1)
	) name4041 (
		_w4394_,
		_w4502_,
		_w4503_
	);
	LUT2 #(
		.INIT('h2)
	) name4042 (
		\P1_reg0_reg[29]/NET0131 ,
		_w3435_,
		_w4504_
	);
	LUT2 #(
		.INIT('h8)
	) name4043 (
		\P1_reg0_reg[29]/NET0131 ,
		_w3448_,
		_w4505_
	);
	LUT2 #(
		.INIT('h2)
	) name4044 (
		\P1_reg0_reg[29]/NET0131 ,
		_w4396_,
		_w4506_
	);
	LUT2 #(
		.INIT('h4)
	) name4045 (
		_w3559_,
		_w4396_,
		_w4507_
	);
	LUT2 #(
		.INIT('h1)
	) name4046 (
		_w4506_,
		_w4507_,
		_w4508_
	);
	LUT2 #(
		.INIT('h1)
	) name4047 (
		_w3563_,
		_w4508_,
		_w4509_
	);
	LUT2 #(
		.INIT('h8)
	) name4048 (
		_w3709_,
		_w4396_,
		_w4510_
	);
	LUT2 #(
		.INIT('h1)
	) name4049 (
		_w4506_,
		_w4510_,
		_w4511_
	);
	LUT2 #(
		.INIT('h2)
	) name4050 (
		_w3712_,
		_w4511_,
		_w4512_
	);
	LUT2 #(
		.INIT('h2)
	) name4051 (
		\P1_reg0_reg[29]/NET0131 ,
		_w4493_,
		_w4513_
	);
	LUT2 #(
		.INIT('h8)
	) name4052 (
		_w3714_,
		_w4396_,
		_w4514_
	);
	LUT2 #(
		.INIT('h4)
	) name4053 (
		_w3602_,
		_w4396_,
		_w4515_
	);
	LUT2 #(
		.INIT('h1)
	) name4054 (
		_w4506_,
		_w4515_,
		_w4516_
	);
	LUT2 #(
		.INIT('h2)
	) name4055 (
		_w1936_,
		_w4516_,
		_w4517_
	);
	LUT2 #(
		.INIT('h8)
	) name4056 (
		_w3673_,
		_w4396_,
		_w4518_
	);
	LUT2 #(
		.INIT('h1)
	) name4057 (
		_w4506_,
		_w4518_,
		_w4519_
	);
	LUT2 #(
		.INIT('h1)
	) name4058 (
		_w3677_,
		_w4519_,
		_w4520_
	);
	LUT2 #(
		.INIT('h1)
	) name4059 (
		_w4513_,
		_w4514_,
		_w4521_
	);
	LUT2 #(
		.INIT('h4)
	) name4060 (
		_w4512_,
		_w4521_,
		_w4522_
	);
	LUT2 #(
		.INIT('h4)
	) name4061 (
		_w4509_,
		_w4522_,
		_w4523_
	);
	LUT2 #(
		.INIT('h1)
	) name4062 (
		_w4517_,
		_w4520_,
		_w4524_
	);
	LUT2 #(
		.INIT('h8)
	) name4063 (
		_w4523_,
		_w4524_,
		_w4525_
	);
	LUT2 #(
		.INIT('h2)
	) name4064 (
		_w3450_,
		_w4525_,
		_w4526_
	);
	LUT2 #(
		.INIT('h1)
	) name4065 (
		_w4505_,
		_w4526_,
		_w4527_
	);
	LUT2 #(
		.INIT('h2)
	) name4066 (
		\P1_state_reg[0]/NET0131 ,
		_w4527_,
		_w4528_
	);
	LUT2 #(
		.INIT('h1)
	) name4067 (
		_w4504_,
		_w4528_,
		_w4529_
	);
	LUT2 #(
		.INIT('h2)
	) name4068 (
		\P1_reg1_reg[29]/NET0131 ,
		_w3435_,
		_w4530_
	);
	LUT2 #(
		.INIT('h8)
	) name4069 (
		\P1_reg1_reg[29]/NET0131 ,
		_w3448_,
		_w4531_
	);
	LUT2 #(
		.INIT('h4)
	) name4070 (
		_w3460_,
		_w3465_,
		_w4532_
	);
	LUT2 #(
		.INIT('h2)
	) name4071 (
		\P1_reg1_reg[29]/NET0131 ,
		_w4532_,
		_w4533_
	);
	LUT2 #(
		.INIT('h4)
	) name4072 (
		_w3559_,
		_w4532_,
		_w4534_
	);
	LUT2 #(
		.INIT('h1)
	) name4073 (
		_w4533_,
		_w4534_,
		_w4535_
	);
	LUT2 #(
		.INIT('h1)
	) name4074 (
		_w3563_,
		_w4535_,
		_w4536_
	);
	LUT2 #(
		.INIT('h8)
	) name4075 (
		_w3709_,
		_w4532_,
		_w4537_
	);
	LUT2 #(
		.INIT('h1)
	) name4076 (
		_w4533_,
		_w4537_,
		_w4538_
	);
	LUT2 #(
		.INIT('h2)
	) name4077 (
		_w3712_,
		_w4538_,
		_w4539_
	);
	LUT2 #(
		.INIT('h2)
	) name4078 (
		_w1880_,
		_w4532_,
		_w4540_
	);
	LUT2 #(
		.INIT('h2)
	) name4079 (
		_w4491_,
		_w4540_,
		_w4541_
	);
	LUT2 #(
		.INIT('h2)
	) name4080 (
		\P1_reg1_reg[29]/NET0131 ,
		_w4541_,
		_w4542_
	);
	LUT2 #(
		.INIT('h8)
	) name4081 (
		_w3714_,
		_w4532_,
		_w4543_
	);
	LUT2 #(
		.INIT('h4)
	) name4082 (
		_w3602_,
		_w4532_,
		_w4544_
	);
	LUT2 #(
		.INIT('h1)
	) name4083 (
		_w4533_,
		_w4544_,
		_w4545_
	);
	LUT2 #(
		.INIT('h2)
	) name4084 (
		_w1936_,
		_w4545_,
		_w4546_
	);
	LUT2 #(
		.INIT('h8)
	) name4085 (
		_w3673_,
		_w4532_,
		_w4547_
	);
	LUT2 #(
		.INIT('h1)
	) name4086 (
		_w4533_,
		_w4547_,
		_w4548_
	);
	LUT2 #(
		.INIT('h1)
	) name4087 (
		_w3677_,
		_w4548_,
		_w4549_
	);
	LUT2 #(
		.INIT('h1)
	) name4088 (
		_w4542_,
		_w4543_,
		_w4550_
	);
	LUT2 #(
		.INIT('h4)
	) name4089 (
		_w4539_,
		_w4550_,
		_w4551_
	);
	LUT2 #(
		.INIT('h4)
	) name4090 (
		_w4536_,
		_w4551_,
		_w4552_
	);
	LUT2 #(
		.INIT('h1)
	) name4091 (
		_w4546_,
		_w4549_,
		_w4553_
	);
	LUT2 #(
		.INIT('h8)
	) name4092 (
		_w4552_,
		_w4553_,
		_w4554_
	);
	LUT2 #(
		.INIT('h2)
	) name4093 (
		_w3450_,
		_w4554_,
		_w4555_
	);
	LUT2 #(
		.INIT('h1)
	) name4094 (
		_w4531_,
		_w4555_,
		_w4556_
	);
	LUT2 #(
		.INIT('h2)
	) name4095 (
		\P1_state_reg[0]/NET0131 ,
		_w4556_,
		_w4557_
	);
	LUT2 #(
		.INIT('h1)
	) name4096 (
		_w4530_,
		_w4557_,
		_w4558_
	);
	LUT2 #(
		.INIT('h2)
	) name4097 (
		\P1_reg1_reg[27]/NET0131 ,
		_w3435_,
		_w4559_
	);
	LUT2 #(
		.INIT('h8)
	) name4098 (
		\P1_reg1_reg[27]/NET0131 ,
		_w3448_,
		_w4560_
	);
	LUT2 #(
		.INIT('h2)
	) name4099 (
		\P1_reg1_reg[27]/NET0131 ,
		_w4532_,
		_w4561_
	);
	LUT2 #(
		.INIT('h4)
	) name4100 (
		_w4429_,
		_w4532_,
		_w4562_
	);
	LUT2 #(
		.INIT('h1)
	) name4101 (
		_w4561_,
		_w4562_,
		_w4563_
	);
	LUT2 #(
		.INIT('h1)
	) name4102 (
		_w3677_,
		_w4563_,
		_w4564_
	);
	LUT2 #(
		.INIT('h4)
	) name4103 (
		_w4466_,
		_w4532_,
		_w4565_
	);
	LUT2 #(
		.INIT('h1)
	) name4104 (
		_w4561_,
		_w4565_,
		_w4566_
	);
	LUT2 #(
		.INIT('h1)
	) name4105 (
		_w3563_,
		_w4566_,
		_w4567_
	);
	LUT2 #(
		.INIT('h8)
	) name4106 (
		_w4480_,
		_w4532_,
		_w4568_
	);
	LUT2 #(
		.INIT('h1)
	) name4107 (
		_w4561_,
		_w4568_,
		_w4569_
	);
	LUT2 #(
		.INIT('h2)
	) name4108 (
		_w1936_,
		_w4569_,
		_w4570_
	);
	LUT2 #(
		.INIT('h4)
	) name4109 (
		_w4488_,
		_w4532_,
		_w4571_
	);
	LUT2 #(
		.INIT('h2)
	) name4110 (
		_w3712_,
		_w4532_,
		_w4572_
	);
	LUT2 #(
		.INIT('h2)
	) name4111 (
		_w4541_,
		_w4572_,
		_w4573_
	);
	LUT2 #(
		.INIT('h2)
	) name4112 (
		\P1_reg1_reg[27]/NET0131 ,
		_w4573_,
		_w4574_
	);
	LUT2 #(
		.INIT('h1)
	) name4113 (
		_w4571_,
		_w4574_,
		_w4575_
	);
	LUT2 #(
		.INIT('h4)
	) name4114 (
		_w4564_,
		_w4575_,
		_w4576_
	);
	LUT2 #(
		.INIT('h1)
	) name4115 (
		_w4567_,
		_w4570_,
		_w4577_
	);
	LUT2 #(
		.INIT('h8)
	) name4116 (
		_w4576_,
		_w4577_,
		_w4578_
	);
	LUT2 #(
		.INIT('h2)
	) name4117 (
		_w3450_,
		_w4578_,
		_w4579_
	);
	LUT2 #(
		.INIT('h1)
	) name4118 (
		_w4560_,
		_w4579_,
		_w4580_
	);
	LUT2 #(
		.INIT('h2)
	) name4119 (
		\P1_state_reg[0]/NET0131 ,
		_w4580_,
		_w4581_
	);
	LUT2 #(
		.INIT('h1)
	) name4120 (
		_w4559_,
		_w4581_,
		_w4582_
	);
	LUT2 #(
		.INIT('h4)
	) name4121 (
		\P1_state_reg[0]/NET0131 ,
		\P2_reg3_reg[25]/NET0131 ,
		_w4583_
	);
	LUT2 #(
		.INIT('h8)
	) name4122 (
		_w3039_,
		_w3976_,
		_w4584_
	);
	LUT2 #(
		.INIT('h8)
	) name4123 (
		_w2024_,
		_w3039_,
		_w4585_
	);
	LUT2 #(
		.INIT('h2)
	) name4124 (
		_w3039_,
		_w3788_,
		_w4586_
	);
	LUT2 #(
		.INIT('h4)
	) name4125 (
		_w2897_,
		_w2908_,
		_w4587_
	);
	LUT2 #(
		.INIT('h8)
	) name4126 (
		_w2445_,
		_w3133_,
		_w4588_
	);
	LUT2 #(
		.INIT('h4)
	) name4127 (
		_w4587_,
		_w4588_,
		_w4589_
	);
	LUT2 #(
		.INIT('h4)
	) name4128 (
		_w2919_,
		_w3133_,
		_w4590_
	);
	LUT2 #(
		.INIT('h2)
	) name4129 (
		_w3147_,
		_w4590_,
		_w4591_
	);
	LUT2 #(
		.INIT('h4)
	) name4130 (
		_w4589_,
		_w4591_,
		_w4592_
	);
	LUT2 #(
		.INIT('h8)
	) name4131 (
		_w4213_,
		_w4592_,
		_w4593_
	);
	LUT2 #(
		.INIT('h1)
	) name4132 (
		_w4213_,
		_w4592_,
		_w4594_
	);
	LUT2 #(
		.INIT('h1)
	) name4133 (
		_w4593_,
		_w4594_,
		_w4595_
	);
	LUT2 #(
		.INIT('h2)
	) name4134 (
		_w3788_,
		_w4595_,
		_w4596_
	);
	LUT2 #(
		.INIT('h1)
	) name4135 (
		_w4586_,
		_w4596_,
		_w4597_
	);
	LUT2 #(
		.INIT('h1)
	) name4136 (
		_w3177_,
		_w4597_,
		_w4598_
	);
	LUT2 #(
		.INIT('h2)
	) name4137 (
		_w3223_,
		_w3238_,
		_w4599_
	);
	LUT2 #(
		.INIT('h2)
	) name4138 (
		_w3291_,
		_w4599_,
		_w4600_
	);
	LUT2 #(
		.INIT('h2)
	) name4139 (
		_w3216_,
		_w4600_,
		_w4601_
	);
	LUT2 #(
		.INIT('h8)
	) name4140 (
		_w3224_,
		_w3279_,
		_w4602_
	);
	LUT2 #(
		.INIT('h2)
	) name4141 (
		_w3302_,
		_w4601_,
		_w4603_
	);
	LUT2 #(
		.INIT('h4)
	) name4142 (
		_w4602_,
		_w4603_,
		_w4604_
	);
	LUT2 #(
		.INIT('h2)
	) name4143 (
		_w3307_,
		_w4604_,
		_w4605_
	);
	LUT2 #(
		.INIT('h2)
	) name4144 (
		_w3199_,
		_w4605_,
		_w4606_
	);
	LUT2 #(
		.INIT('h2)
	) name4145 (
		_w4213_,
		_w4606_,
		_w4607_
	);
	LUT2 #(
		.INIT('h4)
	) name4146 (
		_w4213_,
		_w4606_,
		_w4608_
	);
	LUT2 #(
		.INIT('h1)
	) name4147 (
		_w4607_,
		_w4608_,
		_w4609_
	);
	LUT2 #(
		.INIT('h2)
	) name4148 (
		_w3788_,
		_w4609_,
		_w4610_
	);
	LUT2 #(
		.INIT('h1)
	) name4149 (
		_w4586_,
		_w4610_,
		_w4611_
	);
	LUT2 #(
		.INIT('h1)
	) name4150 (
		_w3320_,
		_w4611_,
		_w4612_
	);
	LUT2 #(
		.INIT('h2)
	) name4151 (
		_w3034_,
		_w3965_,
		_w4613_
	);
	LUT2 #(
		.INIT('h8)
	) name4152 (
		_w3325_,
		_w3343_,
		_w4614_
	);
	LUT2 #(
		.INIT('h4)
	) name4153 (
		_w3054_,
		_w4614_,
		_w4615_
	);
	LUT2 #(
		.INIT('h2)
	) name4154 (
		_w3034_,
		_w4615_,
		_w4616_
	);
	LUT2 #(
		.INIT('h1)
	) name4155 (
		_w3346_,
		_w4616_,
		_w4617_
	);
	LUT2 #(
		.INIT('h8)
	) name4156 (
		_w3788_,
		_w4617_,
		_w4618_
	);
	LUT2 #(
		.INIT('h1)
	) name4157 (
		_w4586_,
		_w4618_,
		_w4619_
	);
	LUT2 #(
		.INIT('h2)
	) name4158 (
		_w3355_,
		_w4619_,
		_w4620_
	);
	LUT2 #(
		.INIT('h8)
	) name4159 (
		_w2058_,
		_w3065_,
		_w4621_
	);
	LUT2 #(
		.INIT('h8)
	) name4160 (
		_w3363_,
		_w3394_,
		_w4622_
	);
	LUT2 #(
		.INIT('h4)
	) name4161 (
		_w3043_,
		_w4622_,
		_w4623_
	);
	LUT2 #(
		.INIT('h2)
	) name4162 (
		_w3021_,
		_w4623_,
		_w4624_
	);
	LUT2 #(
		.INIT('h8)
	) name4163 (
		_w3361_,
		_w4622_,
		_w4625_
	);
	LUT2 #(
		.INIT('h1)
	) name4164 (
		_w4624_,
		_w4625_,
		_w4626_
	);
	LUT2 #(
		.INIT('h1)
	) name4165 (
		_w2058_,
		_w4626_,
		_w4627_
	);
	LUT2 #(
		.INIT('h2)
	) name4166 (
		_w3411_,
		_w4621_,
		_w4628_
	);
	LUT2 #(
		.INIT('h4)
	) name4167 (
		_w4627_,
		_w4628_,
		_w4629_
	);
	LUT2 #(
		.INIT('h8)
	) name4168 (
		_w3788_,
		_w4629_,
		_w4630_
	);
	LUT2 #(
		.INIT('h2)
	) name4169 (
		_w3411_,
		_w3788_,
		_w4631_
	);
	LUT2 #(
		.INIT('h2)
	) name4170 (
		_w3962_,
		_w4631_,
		_w4632_
	);
	LUT2 #(
		.INIT('h2)
	) name4171 (
		_w3039_,
		_w4632_,
		_w4633_
	);
	LUT2 #(
		.INIT('h1)
	) name4172 (
		_w4613_,
		_w4633_,
		_w4634_
	);
	LUT2 #(
		.INIT('h4)
	) name4173 (
		_w4630_,
		_w4634_,
		_w4635_
	);
	LUT2 #(
		.INIT('h4)
	) name4174 (
		_w4620_,
		_w4635_,
		_w4636_
	);
	LUT2 #(
		.INIT('h4)
	) name4175 (
		_w4598_,
		_w4636_,
		_w4637_
	);
	LUT2 #(
		.INIT('h4)
	) name4176 (
		_w4612_,
		_w4637_,
		_w4638_
	);
	LUT2 #(
		.INIT('h2)
	) name4177 (
		_w2026_,
		_w4638_,
		_w4639_
	);
	LUT2 #(
		.INIT('h1)
	) name4178 (
		_w4585_,
		_w4639_,
		_w4640_
	);
	LUT2 #(
		.INIT('h2)
	) name4179 (
		\P1_state_reg[0]/NET0131 ,
		_w4640_,
		_w4641_
	);
	LUT2 #(
		.INIT('h1)
	) name4180 (
		_w4583_,
		_w4584_,
		_w4642_
	);
	LUT2 #(
		.INIT('h4)
	) name4181 (
		_w4641_,
		_w4642_,
		_w4643_
	);
	LUT2 #(
		.INIT('h2)
	) name4182 (
		\P1_reg3_reg[25]/NET0131 ,
		\P1_state_reg[0]/NET0131 ,
		_w4644_
	);
	LUT2 #(
		.INIT('h8)
	) name4183 (
		_w1034_,
		_w1953_,
		_w4645_
	);
	LUT2 #(
		.INIT('h8)
	) name4184 (
		_w1034_,
		_w3448_,
		_w4646_
	);
	LUT2 #(
		.INIT('h2)
	) name4185 (
		_w1034_,
		_w3980_,
		_w4647_
	);
	LUT2 #(
		.INIT('h8)
	) name4186 (
		_w3626_,
		_w3649_,
		_w4648_
	);
	LUT2 #(
		.INIT('h2)
	) name4187 (
		_w3625_,
		_w3632_,
		_w4649_
	);
	LUT2 #(
		.INIT('h2)
	) name4188 (
		_w3656_,
		_w4649_,
		_w4650_
	);
	LUT2 #(
		.INIT('h2)
	) name4189 (
		_w3622_,
		_w4650_,
		_w4651_
	);
	LUT2 #(
		.INIT('h2)
	) name4190 (
		_w3662_,
		_w4651_,
		_w4652_
	);
	LUT2 #(
		.INIT('h4)
	) name4191 (
		_w4648_,
		_w4652_,
		_w4653_
	);
	LUT2 #(
		.INIT('h2)
	) name4192 (
		_w3666_,
		_w4653_,
		_w4654_
	);
	LUT2 #(
		.INIT('h2)
	) name4193 (
		_w3611_,
		_w4654_,
		_w4655_
	);
	LUT2 #(
		.INIT('h2)
	) name4194 (
		_w1812_,
		_w4655_,
		_w4656_
	);
	LUT2 #(
		.INIT('h4)
	) name4195 (
		_w1812_,
		_w4655_,
		_w4657_
	);
	LUT2 #(
		.INIT('h1)
	) name4196 (
		_w4656_,
		_w4657_,
		_w4658_
	);
	LUT2 #(
		.INIT('h2)
	) name4197 (
		_w3980_,
		_w4658_,
		_w4659_
	);
	LUT2 #(
		.INIT('h1)
	) name4198 (
		_w4647_,
		_w4659_,
		_w4660_
	);
	LUT2 #(
		.INIT('h1)
	) name4199 (
		_w3677_,
		_w4660_,
		_w4661_
	);
	LUT2 #(
		.INIT('h8)
	) name4200 (
		_w3491_,
		_w3532_,
		_w4662_
	);
	LUT2 #(
		.INIT('h2)
	) name4201 (
		_w3490_,
		_w3498_,
		_w4663_
	);
	LUT2 #(
		.INIT('h2)
	) name4202 (
		_w3540_,
		_w4663_,
		_w4664_
	);
	LUT2 #(
		.INIT('h2)
	) name4203 (
		_w3487_,
		_w4664_,
		_w4665_
	);
	LUT2 #(
		.INIT('h2)
	) name4204 (
		_w3548_,
		_w4665_,
		_w4666_
	);
	LUT2 #(
		.INIT('h4)
	) name4205 (
		_w4662_,
		_w4666_,
		_w4667_
	);
	LUT2 #(
		.INIT('h2)
	) name4206 (
		_w3552_,
		_w4667_,
		_w4668_
	);
	LUT2 #(
		.INIT('h2)
	) name4207 (
		_w3474_,
		_w4668_,
		_w4669_
	);
	LUT2 #(
		.INIT('h8)
	) name4208 (
		_w1812_,
		_w4669_,
		_w4670_
	);
	LUT2 #(
		.INIT('h1)
	) name4209 (
		_w1812_,
		_w4669_,
		_w4671_
	);
	LUT2 #(
		.INIT('h1)
	) name4210 (
		_w4670_,
		_w4671_,
		_w4672_
	);
	LUT2 #(
		.INIT('h2)
	) name4211 (
		_w3980_,
		_w4672_,
		_w4673_
	);
	LUT2 #(
		.INIT('h1)
	) name4212 (
		_w4647_,
		_w4673_,
		_w4674_
	);
	LUT2 #(
		.INIT('h1)
	) name4213 (
		_w3563_,
		_w4674_,
		_w4675_
	);
	LUT2 #(
		.INIT('h2)
	) name4214 (
		_w1029_,
		_w4067_,
		_w4676_
	);
	LUT2 #(
		.INIT('h2)
	) name4215 (
		_w1034_,
		_w4064_,
		_w4677_
	);
	LUT2 #(
		.INIT('h2)
	) name4216 (
		_w1006_,
		_w3593_,
		_w4678_
	);
	LUT2 #(
		.INIT('h1)
	) name4217 (
		_w3594_,
		_w4678_,
		_w4679_
	);
	LUT2 #(
		.INIT('h1)
	) name4218 (
		_w537_,
		_w4679_,
		_w4680_
	);
	LUT2 #(
		.INIT('h8)
	) name4219 (
		_w537_,
		_w1062_,
		_w4681_
	);
	LUT2 #(
		.INIT('h1)
	) name4220 (
		_w4680_,
		_w4681_,
		_w4682_
	);
	LUT2 #(
		.INIT('h8)
	) name4221 (
		_w3980_,
		_w4682_,
		_w4683_
	);
	LUT2 #(
		.INIT('h1)
	) name4222 (
		_w4647_,
		_w4683_,
		_w4684_
	);
	LUT2 #(
		.INIT('h2)
	) name4223 (
		_w1936_,
		_w4684_,
		_w4685_
	);
	LUT2 #(
		.INIT('h8)
	) name4224 (
		_w3700_,
		_w3701_,
		_w4686_
	);
	LUT2 #(
		.INIT('h2)
	) name4225 (
		_w1029_,
		_w4686_,
		_w4687_
	);
	LUT2 #(
		.INIT('h4)
	) name4226 (
		_w1029_,
		_w4686_,
		_w4688_
	);
	LUT2 #(
		.INIT('h1)
	) name4227 (
		_w4687_,
		_w4688_,
		_w4689_
	);
	LUT2 #(
		.INIT('h8)
	) name4228 (
		_w3980_,
		_w4689_,
		_w4690_
	);
	LUT2 #(
		.INIT('h1)
	) name4229 (
		_w4647_,
		_w4690_,
		_w4691_
	);
	LUT2 #(
		.INIT('h2)
	) name4230 (
		_w3712_,
		_w4691_,
		_w4692_
	);
	LUT2 #(
		.INIT('h1)
	) name4231 (
		_w4676_,
		_w4677_,
		_w4693_
	);
	LUT2 #(
		.INIT('h4)
	) name4232 (
		_w4685_,
		_w4693_,
		_w4694_
	);
	LUT2 #(
		.INIT('h4)
	) name4233 (
		_w4692_,
		_w4694_,
		_w4695_
	);
	LUT2 #(
		.INIT('h1)
	) name4234 (
		_w4661_,
		_w4675_,
		_w4696_
	);
	LUT2 #(
		.INIT('h8)
	) name4235 (
		_w4695_,
		_w4696_,
		_w4697_
	);
	LUT2 #(
		.INIT('h2)
	) name4236 (
		_w3450_,
		_w4697_,
		_w4698_
	);
	LUT2 #(
		.INIT('h1)
	) name4237 (
		_w4646_,
		_w4698_,
		_w4699_
	);
	LUT2 #(
		.INIT('h2)
	) name4238 (
		\P1_state_reg[0]/NET0131 ,
		_w4699_,
		_w4700_
	);
	LUT2 #(
		.INIT('h1)
	) name4239 (
		_w4644_,
		_w4645_,
		_w4701_
	);
	LUT2 #(
		.INIT('h4)
	) name4240 (
		_w4700_,
		_w4701_,
		_w4702_
	);
	LUT2 #(
		.INIT('h2)
	) name4241 (
		_w3017_,
		_w3788_,
		_w4703_
	);
	LUT2 #(
		.INIT('h8)
	) name4242 (
		_w3790_,
		_w3793_,
		_w4704_
	);
	LUT2 #(
		.INIT('h8)
	) name4243 (
		_w3814_,
		_w3817_,
		_w4705_
	);
	LUT2 #(
		.INIT('h4)
	) name4244 (
		_w3827_,
		_w4705_,
		_w4706_
	);
	LUT2 #(
		.INIT('h8)
	) name4245 (
		_w3814_,
		_w3830_,
		_w4707_
	);
	LUT2 #(
		.INIT('h1)
	) name4246 (
		_w3834_,
		_w4707_,
		_w4708_
	);
	LUT2 #(
		.INIT('h4)
	) name4247 (
		_w4706_,
		_w4708_,
		_w4709_
	);
	LUT2 #(
		.INIT('h8)
	) name4248 (
		_w3815_,
		_w3840_,
		_w4710_
	);
	LUT2 #(
		.INIT('h4)
	) name4249 (
		_w4709_,
		_w4710_,
		_w4711_
	);
	LUT2 #(
		.INIT('h8)
	) name4250 (
		_w3837_,
		_w3840_,
		_w4712_
	);
	LUT2 #(
		.INIT('h1)
	) name4251 (
		_w3802_,
		_w4712_,
		_w4713_
	);
	LUT2 #(
		.INIT('h4)
	) name4252 (
		_w4711_,
		_w4713_,
		_w4714_
	);
	LUT2 #(
		.INIT('h8)
	) name4253 (
		_w3798_,
		_w3800_,
		_w4715_
	);
	LUT2 #(
		.INIT('h4)
	) name4254 (
		_w4714_,
		_w4715_,
		_w4716_
	);
	LUT2 #(
		.INIT('h8)
	) name4255 (
		_w3798_,
		_w3805_,
		_w4717_
	);
	LUT2 #(
		.INIT('h2)
	) name4256 (
		_w3809_,
		_w4717_,
		_w4718_
	);
	LUT2 #(
		.INIT('h4)
	) name4257 (
		_w4716_,
		_w4718_,
		_w4719_
	);
	LUT2 #(
		.INIT('h8)
	) name4258 (
		_w3794_,
		_w3797_,
		_w4720_
	);
	LUT2 #(
		.INIT('h4)
	) name4259 (
		_w4719_,
		_w4720_,
		_w4721_
	);
	LUT2 #(
		.INIT('h8)
	) name4260 (
		_w4704_,
		_w4721_,
		_w4722_
	);
	LUT2 #(
		.INIT('h8)
	) name4261 (
		_w3790_,
		_w3851_,
		_w4723_
	);
	LUT2 #(
		.INIT('h2)
	) name4262 (
		_w3794_,
		_w3812_,
		_w4724_
	);
	LUT2 #(
		.INIT('h2)
	) name4263 (
		_w3848_,
		_w4724_,
		_w4725_
	);
	LUT2 #(
		.INIT('h2)
	) name4264 (
		_w4704_,
		_w4725_,
		_w4726_
	);
	LUT2 #(
		.INIT('h1)
	) name4265 (
		_w3856_,
		_w4723_,
		_w4727_
	);
	LUT2 #(
		.INIT('h4)
	) name4266 (
		_w4726_,
		_w4727_,
		_w4728_
	);
	LUT2 #(
		.INIT('h4)
	) name4267 (
		_w4722_,
		_w4728_,
		_w4729_
	);
	LUT2 #(
		.INIT('h2)
	) name4268 (
		_w4214_,
		_w4729_,
		_w4730_
	);
	LUT2 #(
		.INIT('h4)
	) name4269 (
		_w4214_,
		_w4729_,
		_w4731_
	);
	LUT2 #(
		.INIT('h1)
	) name4270 (
		_w4730_,
		_w4731_,
		_w4732_
	);
	LUT2 #(
		.INIT('h2)
	) name4271 (
		_w3788_,
		_w4732_,
		_w4733_
	);
	LUT2 #(
		.INIT('h1)
	) name4272 (
		_w4703_,
		_w4733_,
		_w4734_
	);
	LUT2 #(
		.INIT('h1)
	) name4273 (
		_w3320_,
		_w4734_,
		_w4735_
	);
	LUT2 #(
		.INIT('h8)
	) name4274 (
		_w3876_,
		_w3890_,
		_w4736_
	);
	LUT2 #(
		.INIT('h4)
	) name4275 (
		_w3885_,
		_w4736_,
		_w4737_
	);
	LUT2 #(
		.INIT('h8)
	) name4276 (
		_w3888_,
		_w3890_,
		_w4738_
	);
	LUT2 #(
		.INIT('h2)
	) name4277 (
		_w3871_,
		_w4738_,
		_w4739_
	);
	LUT2 #(
		.INIT('h4)
	) name4278 (
		_w4737_,
		_w4739_,
		_w4740_
	);
	LUT2 #(
		.INIT('h8)
	) name4279 (
		_w3869_,
		_w3895_,
		_w4741_
	);
	LUT2 #(
		.INIT('h4)
	) name4280 (
		_w4740_,
		_w4741_,
		_w4742_
	);
	LUT2 #(
		.INIT('h4)
	) name4281 (
		_w3874_,
		_w3895_,
		_w4743_
	);
	LUT2 #(
		.INIT('h1)
	) name4282 (
		_w3903_,
		_w4743_,
		_w4744_
	);
	LUT2 #(
		.INIT('h4)
	) name4283 (
		_w4742_,
		_w4744_,
		_w4745_
	);
	LUT2 #(
		.INIT('h8)
	) name4284 (
		_w3894_,
		_w3897_,
		_w4746_
	);
	LUT2 #(
		.INIT('h4)
	) name4285 (
		_w4745_,
		_w4746_,
		_w4747_
	);
	LUT2 #(
		.INIT('h8)
	) name4286 (
		_w3897_,
		_w3906_,
		_w4748_
	);
	LUT2 #(
		.INIT('h1)
	) name4287 (
		_w3910_,
		_w4748_,
		_w4749_
	);
	LUT2 #(
		.INIT('h4)
	) name4288 (
		_w4747_,
		_w4749_,
		_w4750_
	);
	LUT2 #(
		.INIT('h8)
	) name4289 (
		_w3917_,
		_w3920_,
		_w4751_
	);
	LUT2 #(
		.INIT('h8)
	) name4290 (
		_w3898_,
		_w3921_,
		_w4752_
	);
	LUT2 #(
		.INIT('h8)
	) name4291 (
		_w4751_,
		_w4752_,
		_w4753_
	);
	LUT2 #(
		.INIT('h4)
	) name4292 (
		_w4750_,
		_w4753_,
		_w4754_
	);
	LUT2 #(
		.INIT('h2)
	) name4293 (
		_w3917_,
		_w3929_,
		_w4755_
	);
	LUT2 #(
		.INIT('h4)
	) name4294 (
		_w3913_,
		_w3921_,
		_w4756_
	);
	LUT2 #(
		.INIT('h2)
	) name4295 (
		_w3926_,
		_w4756_,
		_w4757_
	);
	LUT2 #(
		.INIT('h2)
	) name4296 (
		_w4751_,
		_w4757_,
		_w4758_
	);
	LUT2 #(
		.INIT('h2)
	) name4297 (
		_w3933_,
		_w4755_,
		_w4759_
	);
	LUT2 #(
		.INIT('h4)
	) name4298 (
		_w4758_,
		_w4759_,
		_w4760_
	);
	LUT2 #(
		.INIT('h4)
	) name4299 (
		_w4754_,
		_w4760_,
		_w4761_
	);
	LUT2 #(
		.INIT('h8)
	) name4300 (
		_w4214_,
		_w4761_,
		_w4762_
	);
	LUT2 #(
		.INIT('h1)
	) name4301 (
		_w4214_,
		_w4761_,
		_w4763_
	);
	LUT2 #(
		.INIT('h1)
	) name4302 (
		_w4762_,
		_w4763_,
		_w4764_
	);
	LUT2 #(
		.INIT('h2)
	) name4303 (
		_w3788_,
		_w4764_,
		_w4765_
	);
	LUT2 #(
		.INIT('h1)
	) name4304 (
		_w4703_,
		_w4765_,
		_w4766_
	);
	LUT2 #(
		.INIT('h1)
	) name4305 (
		_w3177_,
		_w4766_,
		_w4767_
	);
	LUT2 #(
		.INIT('h2)
	) name4306 (
		_w2991_,
		_w4625_,
		_w4768_
	);
	LUT2 #(
		.INIT('h8)
	) name4307 (
		_w3365_,
		_w3394_,
		_w4769_
	);
	LUT2 #(
		.INIT('h1)
	) name4308 (
		_w4768_,
		_w4769_,
		_w4770_
	);
	LUT2 #(
		.INIT('h1)
	) name4309 (
		_w2058_,
		_w4770_,
		_w4771_
	);
	LUT2 #(
		.INIT('h8)
	) name4310 (
		_w2058_,
		_w3043_,
		_w4772_
	);
	LUT2 #(
		.INIT('h1)
	) name4311 (
		_w4771_,
		_w4772_,
		_w4773_
	);
	LUT2 #(
		.INIT('h8)
	) name4312 (
		_w3788_,
		_w4773_,
		_w4774_
	);
	LUT2 #(
		.INIT('h1)
	) name4313 (
		_w4703_,
		_w4774_,
		_w4775_
	);
	LUT2 #(
		.INIT('h2)
	) name4314 (
		_w3411_,
		_w4775_,
		_w4776_
	);
	LUT2 #(
		.INIT('h2)
	) name4315 (
		_w3012_,
		_w3346_,
		_w4777_
	);
	LUT2 #(
		.INIT('h4)
	) name4316 (
		_w3012_,
		_w3346_,
		_w4778_
	);
	LUT2 #(
		.INIT('h1)
	) name4317 (
		_w4777_,
		_w4778_,
		_w4779_
	);
	LUT2 #(
		.INIT('h8)
	) name4318 (
		_w3788_,
		_w4779_,
		_w4780_
	);
	LUT2 #(
		.INIT('h1)
	) name4319 (
		_w4703_,
		_w4780_,
		_w4781_
	);
	LUT2 #(
		.INIT('h2)
	) name4320 (
		_w3355_,
		_w4781_,
		_w4782_
	);
	LUT2 #(
		.INIT('h2)
	) name4321 (
		_w3017_,
		_w3962_,
		_w4783_
	);
	LUT2 #(
		.INIT('h2)
	) name4322 (
		_w3012_,
		_w3965_,
		_w4784_
	);
	LUT2 #(
		.INIT('h1)
	) name4323 (
		_w4783_,
		_w4784_,
		_w4785_
	);
	LUT2 #(
		.INIT('h4)
	) name4324 (
		_w4782_,
		_w4785_,
		_w4786_
	);
	LUT2 #(
		.INIT('h4)
	) name4325 (
		_w4776_,
		_w4786_,
		_w4787_
	);
	LUT2 #(
		.INIT('h4)
	) name4326 (
		_w4767_,
		_w4787_,
		_w4788_
	);
	LUT2 #(
		.INIT('h4)
	) name4327 (
		_w4735_,
		_w4788_,
		_w4789_
	);
	LUT2 #(
		.INIT('h2)
	) name4328 (
		_w2026_,
		_w4789_,
		_w4790_
	);
	LUT2 #(
		.INIT('h8)
	) name4329 (
		_w2024_,
		_w3017_,
		_w4791_
	);
	LUT2 #(
		.INIT('h1)
	) name4330 (
		_w4790_,
		_w4791_,
		_w4792_
	);
	LUT2 #(
		.INIT('h2)
	) name4331 (
		\P1_state_reg[0]/NET0131 ,
		_w4792_,
		_w4793_
	);
	LUT2 #(
		.INIT('h8)
	) name4332 (
		_w3017_,
		_w3976_,
		_w4794_
	);
	LUT2 #(
		.INIT('h4)
	) name4333 (
		\P1_state_reg[0]/NET0131 ,
		\P2_reg3_reg[26]/NET0131 ,
		_w4795_
	);
	LUT2 #(
		.INIT('h1)
	) name4334 (
		_w4794_,
		_w4795_,
		_w4796_
	);
	LUT2 #(
		.INIT('h4)
	) name4335 (
		_w4793_,
		_w4796_,
		_w4797_
	);
	LUT2 #(
		.INIT('h2)
	) name4336 (
		_w2987_,
		_w3788_,
		_w4798_
	);
	LUT2 #(
		.INIT('h4)
	) name4337 (
		_w2666_,
		_w2671_,
		_w4799_
	);
	LUT2 #(
		.INIT('h8)
	) name4338 (
		_w2497_,
		_w2781_,
		_w4800_
	);
	LUT2 #(
		.INIT('h4)
	) name4339 (
		_w4799_,
		_w4800_,
		_w4801_
	);
	LUT2 #(
		.INIT('h8)
	) name4340 (
		_w2676_,
		_w2781_,
		_w4802_
	);
	LUT2 #(
		.INIT('h2)
	) name4341 (
		_w2787_,
		_w4802_,
		_w4803_
	);
	LUT2 #(
		.INIT('h4)
	) name4342 (
		_w4801_,
		_w4803_,
		_w4804_
	);
	LUT2 #(
		.INIT('h8)
	) name4343 (
		_w2733_,
		_w2895_,
		_w4805_
	);
	LUT2 #(
		.INIT('h4)
	) name4344 (
		_w4804_,
		_w4805_,
		_w4806_
	);
	LUT2 #(
		.INIT('h8)
	) name4345 (
		_w2792_,
		_w2895_,
		_w4807_
	);
	LUT2 #(
		.INIT('h2)
	) name4346 (
		_w2902_,
		_w4807_,
		_w4808_
	);
	LUT2 #(
		.INIT('h4)
	) name4347 (
		_w4806_,
		_w4808_,
		_w4809_
	);
	LUT2 #(
		.INIT('h8)
	) name4348 (
		_w2444_,
		_w2845_,
		_w4810_
	);
	LUT2 #(
		.INIT('h4)
	) name4349 (
		_w4809_,
		_w4810_,
		_w4811_
	);
	LUT2 #(
		.INIT('h2)
	) name4350 (
		_w2444_,
		_w2907_,
		_w4812_
	);
	LUT2 #(
		.INIT('h1)
	) name4351 (
		_w2913_,
		_w4812_,
		_w4813_
	);
	LUT2 #(
		.INIT('h4)
	) name4352 (
		_w4811_,
		_w4813_,
		_w4814_
	);
	LUT2 #(
		.INIT('h8)
	) name4353 (
		_w3045_,
		_w3090_,
		_w4815_
	);
	LUT2 #(
		.INIT('h8)
	) name4354 (
		_w2370_,
		_w3132_,
		_w4816_
	);
	LUT2 #(
		.INIT('h8)
	) name4355 (
		_w4815_,
		_w4816_,
		_w4817_
	);
	LUT2 #(
		.INIT('h4)
	) name4356 (
		_w4814_,
		_w4817_,
		_w4818_
	);
	LUT2 #(
		.INIT('h2)
	) name4357 (
		_w3045_,
		_w3146_,
		_w4819_
	);
	LUT2 #(
		.INIT('h4)
	) name4358 (
		_w2918_,
		_w3132_,
		_w4820_
	);
	LUT2 #(
		.INIT('h2)
	) name4359 (
		_w3141_,
		_w4820_,
		_w4821_
	);
	LUT2 #(
		.INIT('h2)
	) name4360 (
		_w4815_,
		_w4821_,
		_w4822_
	);
	LUT2 #(
		.INIT('h2)
	) name4361 (
		_w3152_,
		_w4819_,
		_w4823_
	);
	LUT2 #(
		.INIT('h4)
	) name4362 (
		_w4822_,
		_w4823_,
		_w4824_
	);
	LUT2 #(
		.INIT('h4)
	) name4363 (
		_w4818_,
		_w4824_,
		_w4825_
	);
	LUT2 #(
		.INIT('h2)
	) name4364 (
		_w4219_,
		_w4825_,
		_w4826_
	);
	LUT2 #(
		.INIT('h4)
	) name4365 (
		_w4219_,
		_w4825_,
		_w4827_
	);
	LUT2 #(
		.INIT('h1)
	) name4366 (
		_w4826_,
		_w4827_,
		_w4828_
	);
	LUT2 #(
		.INIT('h8)
	) name4367 (
		_w3788_,
		_w4828_,
		_w4829_
	);
	LUT2 #(
		.INIT('h1)
	) name4368 (
		_w4798_,
		_w4829_,
		_w4830_
	);
	LUT2 #(
		.INIT('h1)
	) name4369 (
		_w3177_,
		_w4830_,
		_w4831_
	);
	LUT2 #(
		.INIT('h8)
	) name4370 (
		_w3266_,
		_w3273_,
		_w4832_
	);
	LUT2 #(
		.INIT('h8)
	) name4371 (
		_w3270_,
		_w3273_,
		_w4833_
	);
	LUT2 #(
		.INIT('h1)
	) name4372 (
		_w3248_,
		_w4833_,
		_w4834_
	);
	LUT2 #(
		.INIT('h4)
	) name4373 (
		_w4832_,
		_w4834_,
		_w4835_
	);
	LUT2 #(
		.INIT('h8)
	) name4374 (
		_w3240_,
		_w3243_,
		_w4836_
	);
	LUT2 #(
		.INIT('h4)
	) name4375 (
		_w4835_,
		_w4836_,
		_w4837_
	);
	LUT2 #(
		.INIT('h2)
	) name4376 (
		_w3240_,
		_w3253_,
		_w4838_
	);
	LUT2 #(
		.INIT('h2)
	) name4377 (
		_w3232_,
		_w4838_,
		_w4839_
	);
	LUT2 #(
		.INIT('h4)
	) name4378 (
		_w4837_,
		_w4839_,
		_w4840_
	);
	LUT2 #(
		.INIT('h8)
	) name4379 (
		_w3222_,
		_w3227_,
		_w4841_
	);
	LUT2 #(
		.INIT('h4)
	) name4380 (
		_w4840_,
		_w4841_,
		_w4842_
	);
	LUT2 #(
		.INIT('h2)
	) name4381 (
		_w3222_,
		_w3237_,
		_w4843_
	);
	LUT2 #(
		.INIT('h1)
	) name4382 (
		_w3285_,
		_w4843_,
		_w4844_
	);
	LUT2 #(
		.INIT('h4)
	) name4383 (
		_w4842_,
		_w4844_,
		_w4845_
	);
	LUT2 #(
		.INIT('h8)
	) name4384 (
		_w3215_,
		_w3219_,
		_w4846_
	);
	LUT2 #(
		.INIT('h4)
	) name4385 (
		_w4845_,
		_w4846_,
		_w4847_
	);
	LUT2 #(
		.INIT('h8)
	) name4386 (
		_w3215_,
		_w3290_,
		_w4848_
	);
	LUT2 #(
		.INIT('h1)
	) name4387 (
		_w3296_,
		_w4848_,
		_w4849_
	);
	LUT2 #(
		.INIT('h4)
	) name4388 (
		_w4847_,
		_w4849_,
		_w4850_
	);
	LUT2 #(
		.INIT('h8)
	) name4389 (
		_w3212_,
		_w3306_,
		_w4851_
	);
	LUT2 #(
		.INIT('h8)
	) name4390 (
		_w3184_,
		_w3188_,
		_w4852_
	);
	LUT2 #(
		.INIT('h8)
	) name4391 (
		_w4851_,
		_w4852_,
		_w4853_
	);
	LUT2 #(
		.INIT('h4)
	) name4392 (
		_w4850_,
		_w4853_,
		_w4854_
	);
	LUT2 #(
		.INIT('h8)
	) name4393 (
		_w3301_,
		_w3306_,
		_w4855_
	);
	LUT2 #(
		.INIT('h1)
	) name4394 (
		_w3193_,
		_w4855_,
		_w4856_
	);
	LUT2 #(
		.INIT('h2)
	) name4395 (
		_w4852_,
		_w4856_,
		_w4857_
	);
	LUT2 #(
		.INIT('h2)
	) name4396 (
		_w3184_,
		_w3198_,
		_w4858_
	);
	LUT2 #(
		.INIT('h1)
	) name4397 (
		_w3204_,
		_w4858_,
		_w4859_
	);
	LUT2 #(
		.INIT('h4)
	) name4398 (
		_w4857_,
		_w4859_,
		_w4860_
	);
	LUT2 #(
		.INIT('h4)
	) name4399 (
		_w4854_,
		_w4860_,
		_w4861_
	);
	LUT2 #(
		.INIT('h2)
	) name4400 (
		_w4219_,
		_w4861_,
		_w4862_
	);
	LUT2 #(
		.INIT('h4)
	) name4401 (
		_w4219_,
		_w4861_,
		_w4863_
	);
	LUT2 #(
		.INIT('h1)
	) name4402 (
		_w4862_,
		_w4863_,
		_w4864_
	);
	LUT2 #(
		.INIT('h2)
	) name4403 (
		_w3788_,
		_w4864_,
		_w4865_
	);
	LUT2 #(
		.INIT('h1)
	) name4404 (
		_w4798_,
		_w4865_,
		_w4866_
	);
	LUT2 #(
		.INIT('h1)
	) name4405 (
		_w3320_,
		_w4866_,
		_w4867_
	);
	LUT2 #(
		.INIT('h2)
	) name4406 (
		_w2982_,
		_w4778_,
		_w4868_
	);
	LUT2 #(
		.INIT('h1)
	) name4407 (
		_w3946_,
		_w4868_,
		_w4869_
	);
	LUT2 #(
		.INIT('h8)
	) name4408 (
		_w3788_,
		_w4869_,
		_w4870_
	);
	LUT2 #(
		.INIT('h1)
	) name4409 (
		_w4798_,
		_w4870_,
		_w4871_
	);
	LUT2 #(
		.INIT('h2)
	) name4410 (
		_w3355_,
		_w4871_,
		_w4872_
	);
	LUT2 #(
		.INIT('h2)
	) name4411 (
		_w2962_,
		_w4769_,
		_w4873_
	);
	LUT2 #(
		.INIT('h1)
	) name4412 (
		_w3952_,
		_w4873_,
		_w4874_
	);
	LUT2 #(
		.INIT('h1)
	) name4413 (
		_w2058_,
		_w4874_,
		_w4875_
	);
	LUT2 #(
		.INIT('h8)
	) name4414 (
		_w2058_,
		_w3021_,
		_w4876_
	);
	LUT2 #(
		.INIT('h1)
	) name4415 (
		_w4875_,
		_w4876_,
		_w4877_
	);
	LUT2 #(
		.INIT('h8)
	) name4416 (
		_w3788_,
		_w4877_,
		_w4878_
	);
	LUT2 #(
		.INIT('h1)
	) name4417 (
		_w4798_,
		_w4878_,
		_w4879_
	);
	LUT2 #(
		.INIT('h2)
	) name4418 (
		_w3411_,
		_w4879_,
		_w4880_
	);
	LUT2 #(
		.INIT('h2)
	) name4419 (
		_w2982_,
		_w3965_,
		_w4881_
	);
	LUT2 #(
		.INIT('h2)
	) name4420 (
		_w2987_,
		_w3962_,
		_w4882_
	);
	LUT2 #(
		.INIT('h1)
	) name4421 (
		_w4881_,
		_w4882_,
		_w4883_
	);
	LUT2 #(
		.INIT('h4)
	) name4422 (
		_w4880_,
		_w4883_,
		_w4884_
	);
	LUT2 #(
		.INIT('h4)
	) name4423 (
		_w4867_,
		_w4884_,
		_w4885_
	);
	LUT2 #(
		.INIT('h4)
	) name4424 (
		_w4872_,
		_w4885_,
		_w4886_
	);
	LUT2 #(
		.INIT('h4)
	) name4425 (
		_w4831_,
		_w4886_,
		_w4887_
	);
	LUT2 #(
		.INIT('h2)
	) name4426 (
		_w2026_,
		_w4887_,
		_w4888_
	);
	LUT2 #(
		.INIT('h8)
	) name4427 (
		_w2024_,
		_w2987_,
		_w4889_
	);
	LUT2 #(
		.INIT('h1)
	) name4428 (
		_w4888_,
		_w4889_,
		_w4890_
	);
	LUT2 #(
		.INIT('h2)
	) name4429 (
		\P1_state_reg[0]/NET0131 ,
		_w4890_,
		_w4891_
	);
	LUT2 #(
		.INIT('h4)
	) name4430 (
		\P1_state_reg[0]/NET0131 ,
		\P2_reg3_reg[27]/NET0131 ,
		_w4892_
	);
	LUT2 #(
		.INIT('h8)
	) name4431 (
		_w2987_,
		_w3976_,
		_w4893_
	);
	LUT2 #(
		.INIT('h1)
	) name4432 (
		_w4892_,
		_w4893_,
		_w4894_
	);
	LUT2 #(
		.INIT('h4)
	) name4433 (
		_w4891_,
		_w4894_,
		_w4895_
	);
	LUT2 #(
		.INIT('h2)
	) name4434 (
		\P1_reg3_reg[27]/NET0131 ,
		\P1_state_reg[0]/NET0131 ,
		_w4896_
	);
	LUT2 #(
		.INIT('h8)
	) name4435 (
		_w974_,
		_w1953_,
		_w4897_
	);
	LUT2 #(
		.INIT('h8)
	) name4436 (
		_w974_,
		_w3448_,
		_w4898_
	);
	LUT2 #(
		.INIT('h2)
	) name4437 (
		_w974_,
		_w3980_,
		_w4899_
	);
	LUT2 #(
		.INIT('h2)
	) name4438 (
		_w3980_,
		_w4429_,
		_w4900_
	);
	LUT2 #(
		.INIT('h1)
	) name4439 (
		_w4899_,
		_w4900_,
		_w4901_
	);
	LUT2 #(
		.INIT('h1)
	) name4440 (
		_w3677_,
		_w4901_,
		_w4902_
	);
	LUT2 #(
		.INIT('h8)
	) name4441 (
		_w3980_,
		_w4480_,
		_w4903_
	);
	LUT2 #(
		.INIT('h1)
	) name4442 (
		_w4899_,
		_w4903_,
		_w4904_
	);
	LUT2 #(
		.INIT('h2)
	) name4443 (
		_w1936_,
		_w4904_,
		_w4905_
	);
	LUT2 #(
		.INIT('h2)
	) name4444 (
		_w3980_,
		_w4466_,
		_w4906_
	);
	LUT2 #(
		.INIT('h1)
	) name4445 (
		_w4899_,
		_w4906_,
		_w4907_
	);
	LUT2 #(
		.INIT('h1)
	) name4446 (
		_w3563_,
		_w4907_,
		_w4908_
	);
	LUT2 #(
		.INIT('h2)
	) name4447 (
		_w3712_,
		_w3980_,
		_w4909_
	);
	LUT2 #(
		.INIT('h2)
	) name4448 (
		_w4064_,
		_w4909_,
		_w4910_
	);
	LUT2 #(
		.INIT('h2)
	) name4449 (
		_w974_,
		_w4910_,
		_w4911_
	);
	LUT2 #(
		.INIT('h8)
	) name4450 (
		_w3980_,
		_w4486_,
		_w4912_
	);
	LUT2 #(
		.INIT('h2)
	) name4451 (
		_w969_,
		_w4067_,
		_w4913_
	);
	LUT2 #(
		.INIT('h1)
	) name4452 (
		_w4911_,
		_w4913_,
		_w4914_
	);
	LUT2 #(
		.INIT('h4)
	) name4453 (
		_w4912_,
		_w4914_,
		_w4915_
	);
	LUT2 #(
		.INIT('h4)
	) name4454 (
		_w4902_,
		_w4915_,
		_w4916_
	);
	LUT2 #(
		.INIT('h1)
	) name4455 (
		_w4905_,
		_w4908_,
		_w4917_
	);
	LUT2 #(
		.INIT('h8)
	) name4456 (
		_w4916_,
		_w4917_,
		_w4918_
	);
	LUT2 #(
		.INIT('h2)
	) name4457 (
		_w3450_,
		_w4918_,
		_w4919_
	);
	LUT2 #(
		.INIT('h1)
	) name4458 (
		_w4898_,
		_w4919_,
		_w4920_
	);
	LUT2 #(
		.INIT('h2)
	) name4459 (
		\P1_state_reg[0]/NET0131 ,
		_w4920_,
		_w4921_
	);
	LUT2 #(
		.INIT('h1)
	) name4460 (
		_w4896_,
		_w4897_,
		_w4922_
	);
	LUT2 #(
		.INIT('h4)
	) name4461 (
		_w4921_,
		_w4922_,
		_w4923_
	);
	LUT2 #(
		.INIT('h2)
	) name4462 (
		\P2_reg2_reg[25]/NET0131 ,
		_w1983_,
		_w4924_
	);
	LUT2 #(
		.INIT('h8)
	) name4463 (
		\P2_reg2_reg[25]/NET0131 ,
		_w2024_,
		_w4925_
	);
	LUT2 #(
		.INIT('h8)
	) name4464 (
		_w3355_,
		_w4617_,
		_w4926_
	);
	LUT2 #(
		.INIT('h8)
	) name4465 (
		_w3034_,
		_w3358_,
		_w4927_
	);
	LUT2 #(
		.INIT('h1)
	) name4466 (
		_w4629_,
		_w4927_,
		_w4928_
	);
	LUT2 #(
		.INIT('h4)
	) name4467 (
		_w4926_,
		_w4928_,
		_w4929_
	);
	LUT2 #(
		.INIT('h2)
	) name4468 (
		_w3758_,
		_w4929_,
		_w4930_
	);
	LUT2 #(
		.INIT('h8)
	) name4469 (
		_w3039_,
		_w3420_,
		_w4931_
	);
	LUT2 #(
		.INIT('h2)
	) name4470 (
		_w3745_,
		_w3758_,
		_w4932_
	);
	LUT2 #(
		.INIT('h2)
	) name4471 (
		_w3774_,
		_w4932_,
		_w4933_
	);
	LUT2 #(
		.INIT('h2)
	) name4472 (
		\P2_reg2_reg[25]/NET0131 ,
		_w4933_,
		_w4934_
	);
	LUT2 #(
		.INIT('h2)
	) name4473 (
		\P2_reg2_reg[25]/NET0131 ,
		_w3758_,
		_w4935_
	);
	LUT2 #(
		.INIT('h2)
	) name4474 (
		_w3758_,
		_w4595_,
		_w4936_
	);
	LUT2 #(
		.INIT('h1)
	) name4475 (
		_w4935_,
		_w4936_,
		_w4937_
	);
	LUT2 #(
		.INIT('h1)
	) name4476 (
		_w3177_,
		_w4937_,
		_w4938_
	);
	LUT2 #(
		.INIT('h2)
	) name4477 (
		_w3758_,
		_w4609_,
		_w4939_
	);
	LUT2 #(
		.INIT('h1)
	) name4478 (
		_w4935_,
		_w4939_,
		_w4940_
	);
	LUT2 #(
		.INIT('h1)
	) name4479 (
		_w3320_,
		_w4940_,
		_w4941_
	);
	LUT2 #(
		.INIT('h1)
	) name4480 (
		_w4931_,
		_w4934_,
		_w4942_
	);
	LUT2 #(
		.INIT('h4)
	) name4481 (
		_w4930_,
		_w4942_,
		_w4943_
	);
	LUT2 #(
		.INIT('h4)
	) name4482 (
		_w4938_,
		_w4943_,
		_w4944_
	);
	LUT2 #(
		.INIT('h4)
	) name4483 (
		_w4941_,
		_w4944_,
		_w4945_
	);
	LUT2 #(
		.INIT('h2)
	) name4484 (
		_w2026_,
		_w4945_,
		_w4946_
	);
	LUT2 #(
		.INIT('h1)
	) name4485 (
		_w4925_,
		_w4946_,
		_w4947_
	);
	LUT2 #(
		.INIT('h2)
	) name4486 (
		\P1_state_reg[0]/NET0131 ,
		_w4947_,
		_w4948_
	);
	LUT2 #(
		.INIT('h1)
	) name4487 (
		_w4924_,
		_w4948_,
		_w4949_
	);
	LUT2 #(
		.INIT('h8)
	) name4488 (
		\P2_reg2_reg[26]/NET0131 ,
		_w2024_,
		_w4950_
	);
	LUT2 #(
		.INIT('h2)
	) name4489 (
		\P2_reg2_reg[26]/NET0131 ,
		_w3758_,
		_w4951_
	);
	LUT2 #(
		.INIT('h2)
	) name4490 (
		_w3758_,
		_w4732_,
		_w4952_
	);
	LUT2 #(
		.INIT('h1)
	) name4491 (
		_w4951_,
		_w4952_,
		_w4953_
	);
	LUT2 #(
		.INIT('h1)
	) name4492 (
		_w3320_,
		_w4953_,
		_w4954_
	);
	LUT2 #(
		.INIT('h2)
	) name4493 (
		_w3758_,
		_w4764_,
		_w4955_
	);
	LUT2 #(
		.INIT('h1)
	) name4494 (
		_w4951_,
		_w4955_,
		_w4956_
	);
	LUT2 #(
		.INIT('h1)
	) name4495 (
		_w3177_,
		_w4956_,
		_w4957_
	);
	LUT2 #(
		.INIT('h8)
	) name4496 (
		_w3411_,
		_w4773_,
		_w4958_
	);
	LUT2 #(
		.INIT('h8)
	) name4497 (
		_w3012_,
		_w3358_,
		_w4959_
	);
	LUT2 #(
		.INIT('h8)
	) name4498 (
		_w3355_,
		_w4779_,
		_w4960_
	);
	LUT2 #(
		.INIT('h1)
	) name4499 (
		_w4959_,
		_w4960_,
		_w4961_
	);
	LUT2 #(
		.INIT('h4)
	) name4500 (
		_w4958_,
		_w4961_,
		_w4962_
	);
	LUT2 #(
		.INIT('h2)
	) name4501 (
		_w3758_,
		_w4962_,
		_w4963_
	);
	LUT2 #(
		.INIT('h8)
	) name4502 (
		_w3017_,
		_w3420_,
		_w4964_
	);
	LUT2 #(
		.INIT('h2)
	) name4503 (
		\P2_reg2_reg[26]/NET0131 ,
		_w4384_,
		_w4965_
	);
	LUT2 #(
		.INIT('h1)
	) name4504 (
		_w4964_,
		_w4965_,
		_w4966_
	);
	LUT2 #(
		.INIT('h4)
	) name4505 (
		_w4963_,
		_w4966_,
		_w4967_
	);
	LUT2 #(
		.INIT('h4)
	) name4506 (
		_w4957_,
		_w4967_,
		_w4968_
	);
	LUT2 #(
		.INIT('h4)
	) name4507 (
		_w4954_,
		_w4968_,
		_w4969_
	);
	LUT2 #(
		.INIT('h2)
	) name4508 (
		_w2026_,
		_w4969_,
		_w4970_
	);
	LUT2 #(
		.INIT('h1)
	) name4509 (
		_w4950_,
		_w4970_,
		_w4971_
	);
	LUT2 #(
		.INIT('h2)
	) name4510 (
		\P1_state_reg[0]/NET0131 ,
		_w4971_,
		_w4972_
	);
	LUT2 #(
		.INIT('h2)
	) name4511 (
		\P2_reg2_reg[26]/NET0131 ,
		_w1983_,
		_w4973_
	);
	LUT2 #(
		.INIT('h1)
	) name4512 (
		_w4972_,
		_w4973_,
		_w4974_
	);
	LUT2 #(
		.INIT('h2)
	) name4513 (
		\P2_reg0_reg[24]/NET0131 ,
		_w1983_,
		_w4975_
	);
	LUT2 #(
		.INIT('h8)
	) name4514 (
		\P2_reg0_reg[24]/NET0131 ,
		_w2024_,
		_w4976_
	);
	LUT2 #(
		.INIT('h2)
	) name4515 (
		\P2_reg0_reg[24]/NET0131 ,
		_w2040_,
		_w4977_
	);
	LUT2 #(
		.INIT('h2)
	) name4516 (
		_w3813_,
		_w4170_,
		_w4978_
	);
	LUT2 #(
		.INIT('h2)
	) name4517 (
		_w3795_,
		_w4978_,
		_w4979_
	);
	LUT2 #(
		.INIT('h2)
	) name4518 (
		_w3852_,
		_w4979_,
		_w4980_
	);
	LUT2 #(
		.INIT('h2)
	) name4519 (
		_w4200_,
		_w4980_,
		_w4981_
	);
	LUT2 #(
		.INIT('h4)
	) name4520 (
		_w4200_,
		_w4980_,
		_w4982_
	);
	LUT2 #(
		.INIT('h1)
	) name4521 (
		_w4981_,
		_w4982_,
		_w4983_
	);
	LUT2 #(
		.INIT('h2)
	) name4522 (
		_w2040_,
		_w4983_,
		_w4984_
	);
	LUT2 #(
		.INIT('h1)
	) name4523 (
		_w4977_,
		_w4984_,
		_w4985_
	);
	LUT2 #(
		.INIT('h1)
	) name4524 (
		_w3320_,
		_w4985_,
		_w4986_
	);
	LUT2 #(
		.INIT('h4)
	) name4525 (
		_w3875_,
		_w3896_,
		_w4987_
	);
	LUT2 #(
		.INIT('h2)
	) name4526 (
		_w3907_,
		_w4987_,
		_w4988_
	);
	LUT2 #(
		.INIT('h2)
	) name4527 (
		_w3899_,
		_w4988_,
		_w4989_
	);
	LUT2 #(
		.INIT('h8)
	) name4528 (
		_w3892_,
		_w3900_,
		_w4990_
	);
	LUT2 #(
		.INIT('h2)
	) name4529 (
		_w3914_,
		_w4989_,
		_w4991_
	);
	LUT2 #(
		.INIT('h4)
	) name4530 (
		_w4990_,
		_w4991_,
		_w4992_
	);
	LUT2 #(
		.INIT('h2)
	) name4531 (
		_w3922_,
		_w4992_,
		_w4993_
	);
	LUT2 #(
		.INIT('h2)
	) name4532 (
		_w3930_,
		_w4993_,
		_w4994_
	);
	LUT2 #(
		.INIT('h8)
	) name4533 (
		_w4200_,
		_w4994_,
		_w4995_
	);
	LUT2 #(
		.INIT('h1)
	) name4534 (
		_w4200_,
		_w4994_,
		_w4996_
	);
	LUT2 #(
		.INIT('h1)
	) name4535 (
		_w4995_,
		_w4996_,
		_w4997_
	);
	LUT2 #(
		.INIT('h2)
	) name4536 (
		_w2040_,
		_w4997_,
		_w4998_
	);
	LUT2 #(
		.INIT('h1)
	) name4537 (
		_w4977_,
		_w4998_,
		_w4999_
	);
	LUT2 #(
		.INIT('h1)
	) name4538 (
		_w3177_,
		_w4999_,
		_w5000_
	);
	LUT2 #(
		.INIT('h2)
	) name4539 (
		_w3054_,
		_w4614_,
		_w5001_
	);
	LUT2 #(
		.INIT('h1)
	) name4540 (
		_w4615_,
		_w5001_,
		_w5002_
	);
	LUT2 #(
		.INIT('h8)
	) name4541 (
		_w3355_,
		_w5002_,
		_w5003_
	);
	LUT2 #(
		.INIT('h2)
	) name4542 (
		_w3043_,
		_w4622_,
		_w5004_
	);
	LUT2 #(
		.INIT('h1)
	) name4543 (
		_w4623_,
		_w5004_,
		_w5005_
	);
	LUT2 #(
		.INIT('h1)
	) name4544 (
		_w2058_,
		_w5005_,
		_w5006_
	);
	LUT2 #(
		.INIT('h8)
	) name4545 (
		_w2058_,
		_w3088_,
		_w5007_
	);
	LUT2 #(
		.INIT('h1)
	) name4546 (
		_w5006_,
		_w5007_,
		_w5008_
	);
	LUT2 #(
		.INIT('h8)
	) name4547 (
		_w3411_,
		_w5008_,
		_w5009_
	);
	LUT2 #(
		.INIT('h8)
	) name4548 (
		_w3054_,
		_w3358_,
		_w5010_
	);
	LUT2 #(
		.INIT('h1)
	) name4549 (
		_w5003_,
		_w5010_,
		_w5011_
	);
	LUT2 #(
		.INIT('h4)
	) name4550 (
		_w5009_,
		_w5011_,
		_w5012_
	);
	LUT2 #(
		.INIT('h2)
	) name4551 (
		_w2040_,
		_w5012_,
		_w5013_
	);
	LUT2 #(
		.INIT('h2)
	) name4552 (
		\P2_reg0_reg[24]/NET0131 ,
		_w3426_,
		_w5014_
	);
	LUT2 #(
		.INIT('h1)
	) name4553 (
		_w5013_,
		_w5014_,
		_w5015_
	);
	LUT2 #(
		.INIT('h4)
	) name4554 (
		_w5000_,
		_w5015_,
		_w5016_
	);
	LUT2 #(
		.INIT('h4)
	) name4555 (
		_w4986_,
		_w5016_,
		_w5017_
	);
	LUT2 #(
		.INIT('h2)
	) name4556 (
		_w2026_,
		_w5017_,
		_w5018_
	);
	LUT2 #(
		.INIT('h1)
	) name4557 (
		_w4976_,
		_w5018_,
		_w5019_
	);
	LUT2 #(
		.INIT('h2)
	) name4558 (
		\P1_state_reg[0]/NET0131 ,
		_w5019_,
		_w5020_
	);
	LUT2 #(
		.INIT('h1)
	) name4559 (
		_w4975_,
		_w5020_,
		_w5021_
	);
	LUT2 #(
		.INIT('h8)
	) name4560 (
		\P2_reg0_reg[27]/NET0131 ,
		_w2024_,
		_w5022_
	);
	LUT2 #(
		.INIT('h2)
	) name4561 (
		\P2_reg0_reg[27]/NET0131 ,
		_w2040_,
		_w5023_
	);
	LUT2 #(
		.INIT('h8)
	) name4562 (
		_w2040_,
		_w4828_,
		_w5024_
	);
	LUT2 #(
		.INIT('h1)
	) name4563 (
		_w5023_,
		_w5024_,
		_w5025_
	);
	LUT2 #(
		.INIT('h1)
	) name4564 (
		_w3177_,
		_w5025_,
		_w5026_
	);
	LUT2 #(
		.INIT('h8)
	) name4565 (
		_w2040_,
		_w4869_,
		_w5027_
	);
	LUT2 #(
		.INIT('h1)
	) name4566 (
		_w5023_,
		_w5027_,
		_w5028_
	);
	LUT2 #(
		.INIT('h2)
	) name4567 (
		_w3355_,
		_w5028_,
		_w5029_
	);
	LUT2 #(
		.INIT('h2)
	) name4568 (
		_w2040_,
		_w4864_,
		_w5030_
	);
	LUT2 #(
		.INIT('h1)
	) name4569 (
		_w5023_,
		_w5030_,
		_w5031_
	);
	LUT2 #(
		.INIT('h1)
	) name4570 (
		_w3320_,
		_w5031_,
		_w5032_
	);
	LUT2 #(
		.INIT('h8)
	) name4571 (
		_w2040_,
		_w4877_,
		_w5033_
	);
	LUT2 #(
		.INIT('h1)
	) name4572 (
		_w5023_,
		_w5033_,
		_w5034_
	);
	LUT2 #(
		.INIT('h2)
	) name4573 (
		_w3411_,
		_w5034_,
		_w5035_
	);
	LUT2 #(
		.INIT('h8)
	) name4574 (
		_w2982_,
		_w3358_,
		_w5036_
	);
	LUT2 #(
		.INIT('h8)
	) name4575 (
		_w2040_,
		_w5036_,
		_w5037_
	);
	LUT2 #(
		.INIT('h2)
	) name4576 (
		\P2_reg0_reg[27]/NET0131 ,
		_w3423_,
		_w5038_
	);
	LUT2 #(
		.INIT('h1)
	) name4577 (
		_w5037_,
		_w5038_,
		_w5039_
	);
	LUT2 #(
		.INIT('h4)
	) name4578 (
		_w5035_,
		_w5039_,
		_w5040_
	);
	LUT2 #(
		.INIT('h4)
	) name4579 (
		_w5029_,
		_w5040_,
		_w5041_
	);
	LUT2 #(
		.INIT('h4)
	) name4580 (
		_w5032_,
		_w5041_,
		_w5042_
	);
	LUT2 #(
		.INIT('h4)
	) name4581 (
		_w5026_,
		_w5042_,
		_w5043_
	);
	LUT2 #(
		.INIT('h2)
	) name4582 (
		_w2026_,
		_w5043_,
		_w5044_
	);
	LUT2 #(
		.INIT('h1)
	) name4583 (
		_w5022_,
		_w5044_,
		_w5045_
	);
	LUT2 #(
		.INIT('h2)
	) name4584 (
		\P1_state_reg[0]/NET0131 ,
		_w5045_,
		_w5046_
	);
	LUT2 #(
		.INIT('h2)
	) name4585 (
		\P2_reg0_reg[27]/NET0131 ,
		_w1983_,
		_w5047_
	);
	LUT2 #(
		.INIT('h1)
	) name4586 (
		_w5046_,
		_w5047_,
		_w5048_
	);
	LUT2 #(
		.INIT('h2)
	) name4587 (
		\P1_reg2_reg[27]/NET0131 ,
		_w3435_,
		_w5049_
	);
	LUT2 #(
		.INIT('h8)
	) name4588 (
		\P1_reg2_reg[27]/NET0131 ,
		_w3448_,
		_w5050_
	);
	LUT2 #(
		.INIT('h2)
	) name4589 (
		\P1_reg2_reg[27]/NET0131 ,
		_w3466_,
		_w5051_
	);
	LUT2 #(
		.INIT('h2)
	) name4590 (
		_w3466_,
		_w4429_,
		_w5052_
	);
	LUT2 #(
		.INIT('h1)
	) name4591 (
		_w5051_,
		_w5052_,
		_w5053_
	);
	LUT2 #(
		.INIT('h1)
	) name4592 (
		_w3677_,
		_w5053_,
		_w5054_
	);
	LUT2 #(
		.INIT('h8)
	) name4593 (
		_w3466_,
		_w4480_,
		_w5055_
	);
	LUT2 #(
		.INIT('h1)
	) name4594 (
		_w5051_,
		_w5055_,
		_w5056_
	);
	LUT2 #(
		.INIT('h2)
	) name4595 (
		_w1936_,
		_w5056_,
		_w5057_
	);
	LUT2 #(
		.INIT('h2)
	) name4596 (
		_w3466_,
		_w4466_,
		_w5058_
	);
	LUT2 #(
		.INIT('h1)
	) name4597 (
		_w5051_,
		_w5058_,
		_w5059_
	);
	LUT2 #(
		.INIT('h1)
	) name4598 (
		_w3563_,
		_w5059_,
		_w5060_
	);
	LUT2 #(
		.INIT('h8)
	) name4599 (
		_w974_,
		_w1763_,
		_w5061_
	);
	LUT2 #(
		.INIT('h8)
	) name4600 (
		_w3466_,
		_w4485_,
		_w5062_
	);
	LUT2 #(
		.INIT('h1)
	) name4601 (
		_w5051_,
		_w5062_,
		_w5063_
	);
	LUT2 #(
		.INIT('h2)
	) name4602 (
		_w3712_,
		_w5063_,
		_w5064_
	);
	LUT2 #(
		.INIT('h8)
	) name4603 (
		_w969_,
		_w3466_,
		_w5065_
	);
	LUT2 #(
		.INIT('h1)
	) name4604 (
		_w5051_,
		_w5065_,
		_w5066_
	);
	LUT2 #(
		.INIT('h2)
	) name4605 (
		_w1880_,
		_w5066_,
		_w5067_
	);
	LUT2 #(
		.INIT('h8)
	) name4606 (
		\P1_reg2_reg[27]/NET0131 ,
		_w3716_,
		_w5068_
	);
	LUT2 #(
		.INIT('h1)
	) name4607 (
		_w5061_,
		_w5068_,
		_w5069_
	);
	LUT2 #(
		.INIT('h4)
	) name4608 (
		_w5067_,
		_w5069_,
		_w5070_
	);
	LUT2 #(
		.INIT('h4)
	) name4609 (
		_w5064_,
		_w5070_,
		_w5071_
	);
	LUT2 #(
		.INIT('h4)
	) name4610 (
		_w5054_,
		_w5071_,
		_w5072_
	);
	LUT2 #(
		.INIT('h1)
	) name4611 (
		_w5057_,
		_w5060_,
		_w5073_
	);
	LUT2 #(
		.INIT('h8)
	) name4612 (
		_w5072_,
		_w5073_,
		_w5074_
	);
	LUT2 #(
		.INIT('h2)
	) name4613 (
		_w3450_,
		_w5074_,
		_w5075_
	);
	LUT2 #(
		.INIT('h1)
	) name4614 (
		_w5050_,
		_w5075_,
		_w5076_
	);
	LUT2 #(
		.INIT('h2)
	) name4615 (
		\P1_state_reg[0]/NET0131 ,
		_w5076_,
		_w5077_
	);
	LUT2 #(
		.INIT('h1)
	) name4616 (
		_w5049_,
		_w5077_,
		_w5078_
	);
	LUT2 #(
		.INIT('h2)
	) name4617 (
		\P2_reg1_reg[24]/NET0131 ,
		_w1983_,
		_w5079_
	);
	LUT2 #(
		.INIT('h8)
	) name4618 (
		\P2_reg1_reg[24]/NET0131 ,
		_w2024_,
		_w5080_
	);
	LUT2 #(
		.INIT('h2)
	) name4619 (
		\P2_reg1_reg[24]/NET0131 ,
		_w3733_,
		_w5081_
	);
	LUT2 #(
		.INIT('h2)
	) name4620 (
		_w3733_,
		_w4983_,
		_w5082_
	);
	LUT2 #(
		.INIT('h1)
	) name4621 (
		_w5081_,
		_w5082_,
		_w5083_
	);
	LUT2 #(
		.INIT('h1)
	) name4622 (
		_w3320_,
		_w5083_,
		_w5084_
	);
	LUT2 #(
		.INIT('h2)
	) name4623 (
		_w3733_,
		_w4997_,
		_w5085_
	);
	LUT2 #(
		.INIT('h1)
	) name4624 (
		_w5081_,
		_w5085_,
		_w5086_
	);
	LUT2 #(
		.INIT('h1)
	) name4625 (
		_w3177_,
		_w5086_,
		_w5087_
	);
	LUT2 #(
		.INIT('h2)
	) name4626 (
		_w3733_,
		_w5012_,
		_w5088_
	);
	LUT2 #(
		.INIT('h2)
	) name4627 (
		\P2_reg1_reg[24]/NET0131 ,
		_w3747_,
		_w5089_
	);
	LUT2 #(
		.INIT('h1)
	) name4628 (
		_w5088_,
		_w5089_,
		_w5090_
	);
	LUT2 #(
		.INIT('h4)
	) name4629 (
		_w5087_,
		_w5090_,
		_w5091_
	);
	LUT2 #(
		.INIT('h4)
	) name4630 (
		_w5084_,
		_w5091_,
		_w5092_
	);
	LUT2 #(
		.INIT('h2)
	) name4631 (
		_w2026_,
		_w5092_,
		_w5093_
	);
	LUT2 #(
		.INIT('h1)
	) name4632 (
		_w5080_,
		_w5093_,
		_w5094_
	);
	LUT2 #(
		.INIT('h2)
	) name4633 (
		\P1_state_reg[0]/NET0131 ,
		_w5094_,
		_w5095_
	);
	LUT2 #(
		.INIT('h1)
	) name4634 (
		_w5079_,
		_w5095_,
		_w5096_
	);
	LUT2 #(
		.INIT('h2)
	) name4635 (
		\P2_reg1_reg[25]/NET0131 ,
		_w1983_,
		_w5097_
	);
	LUT2 #(
		.INIT('h8)
	) name4636 (
		\P2_reg1_reg[25]/NET0131 ,
		_w2024_,
		_w5098_
	);
	LUT2 #(
		.INIT('h2)
	) name4637 (
		\P2_reg1_reg[25]/NET0131 ,
		_w3747_,
		_w5099_
	);
	LUT2 #(
		.INIT('h2)
	) name4638 (
		_w3733_,
		_w4929_,
		_w5100_
	);
	LUT2 #(
		.INIT('h2)
	) name4639 (
		\P2_reg1_reg[25]/NET0131 ,
		_w3733_,
		_w5101_
	);
	LUT2 #(
		.INIT('h2)
	) name4640 (
		_w3733_,
		_w4595_,
		_w5102_
	);
	LUT2 #(
		.INIT('h1)
	) name4641 (
		_w5101_,
		_w5102_,
		_w5103_
	);
	LUT2 #(
		.INIT('h1)
	) name4642 (
		_w3177_,
		_w5103_,
		_w5104_
	);
	LUT2 #(
		.INIT('h2)
	) name4643 (
		_w3733_,
		_w4609_,
		_w5105_
	);
	LUT2 #(
		.INIT('h1)
	) name4644 (
		_w5101_,
		_w5105_,
		_w5106_
	);
	LUT2 #(
		.INIT('h1)
	) name4645 (
		_w3320_,
		_w5106_,
		_w5107_
	);
	LUT2 #(
		.INIT('h1)
	) name4646 (
		_w5099_,
		_w5100_,
		_w5108_
	);
	LUT2 #(
		.INIT('h4)
	) name4647 (
		_w5104_,
		_w5108_,
		_w5109_
	);
	LUT2 #(
		.INIT('h4)
	) name4648 (
		_w5107_,
		_w5109_,
		_w5110_
	);
	LUT2 #(
		.INIT('h2)
	) name4649 (
		_w2026_,
		_w5110_,
		_w5111_
	);
	LUT2 #(
		.INIT('h1)
	) name4650 (
		_w5098_,
		_w5111_,
		_w5112_
	);
	LUT2 #(
		.INIT('h2)
	) name4651 (
		\P1_state_reg[0]/NET0131 ,
		_w5112_,
		_w5113_
	);
	LUT2 #(
		.INIT('h1)
	) name4652 (
		_w5097_,
		_w5113_,
		_w5114_
	);
	LUT2 #(
		.INIT('h2)
	) name4653 (
		\P2_reg1_reg[26]/NET0131 ,
		_w1983_,
		_w5115_
	);
	LUT2 #(
		.INIT('h2)
	) name4654 (
		\P2_reg1_reg[26]/NET0131 ,
		_w3733_,
		_w5116_
	);
	LUT2 #(
		.INIT('h2)
	) name4655 (
		_w3733_,
		_w4732_,
		_w5117_
	);
	LUT2 #(
		.INIT('h1)
	) name4656 (
		_w5116_,
		_w5117_,
		_w5118_
	);
	LUT2 #(
		.INIT('h1)
	) name4657 (
		_w3320_,
		_w5118_,
		_w5119_
	);
	LUT2 #(
		.INIT('h2)
	) name4658 (
		_w3733_,
		_w4764_,
		_w5120_
	);
	LUT2 #(
		.INIT('h1)
	) name4659 (
		_w5116_,
		_w5120_,
		_w5121_
	);
	LUT2 #(
		.INIT('h1)
	) name4660 (
		_w3177_,
		_w5121_,
		_w5122_
	);
	LUT2 #(
		.INIT('h2)
	) name4661 (
		_w3733_,
		_w4962_,
		_w5123_
	);
	LUT2 #(
		.INIT('h2)
	) name4662 (
		\P2_reg1_reg[26]/NET0131 ,
		_w3747_,
		_w5124_
	);
	LUT2 #(
		.INIT('h1)
	) name4663 (
		_w5123_,
		_w5124_,
		_w5125_
	);
	LUT2 #(
		.INIT('h4)
	) name4664 (
		_w5122_,
		_w5125_,
		_w5126_
	);
	LUT2 #(
		.INIT('h4)
	) name4665 (
		_w5119_,
		_w5126_,
		_w5127_
	);
	LUT2 #(
		.INIT('h2)
	) name4666 (
		_w2026_,
		_w5127_,
		_w5128_
	);
	LUT2 #(
		.INIT('h8)
	) name4667 (
		\P2_reg1_reg[26]/NET0131 ,
		_w2024_,
		_w5129_
	);
	LUT2 #(
		.INIT('h1)
	) name4668 (
		_w5128_,
		_w5129_,
		_w5130_
	);
	LUT2 #(
		.INIT('h2)
	) name4669 (
		\P1_state_reg[0]/NET0131 ,
		_w5130_,
		_w5131_
	);
	LUT2 #(
		.INIT('h1)
	) name4670 (
		_w5115_,
		_w5131_,
		_w5132_
	);
	LUT2 #(
		.INIT('h2)
	) name4671 (
		\P2_reg1_reg[27]/NET0131 ,
		_w3733_,
		_w5133_
	);
	LUT2 #(
		.INIT('h8)
	) name4672 (
		_w3733_,
		_w4828_,
		_w5134_
	);
	LUT2 #(
		.INIT('h1)
	) name4673 (
		_w5133_,
		_w5134_,
		_w5135_
	);
	LUT2 #(
		.INIT('h1)
	) name4674 (
		_w3177_,
		_w5135_,
		_w5136_
	);
	LUT2 #(
		.INIT('h2)
	) name4675 (
		_w3733_,
		_w4864_,
		_w5137_
	);
	LUT2 #(
		.INIT('h1)
	) name4676 (
		_w5133_,
		_w5137_,
		_w5138_
	);
	LUT2 #(
		.INIT('h1)
	) name4677 (
		_w3320_,
		_w5138_,
		_w5139_
	);
	LUT2 #(
		.INIT('h8)
	) name4678 (
		_w3733_,
		_w4869_,
		_w5140_
	);
	LUT2 #(
		.INIT('h1)
	) name4679 (
		_w5133_,
		_w5140_,
		_w5141_
	);
	LUT2 #(
		.INIT('h2)
	) name4680 (
		_w3355_,
		_w5141_,
		_w5142_
	);
	LUT2 #(
		.INIT('h8)
	) name4681 (
		_w3733_,
		_w4877_,
		_w5143_
	);
	LUT2 #(
		.INIT('h1)
	) name4682 (
		_w5133_,
		_w5143_,
		_w5144_
	);
	LUT2 #(
		.INIT('h2)
	) name4683 (
		_w3411_,
		_w5144_,
		_w5145_
	);
	LUT2 #(
		.INIT('h8)
	) name4684 (
		_w3733_,
		_w5036_,
		_w5146_
	);
	LUT2 #(
		.INIT('h2)
	) name4685 (
		\P2_reg1_reg[27]/NET0131 ,
		_w3743_,
		_w5147_
	);
	LUT2 #(
		.INIT('h1)
	) name4686 (
		_w5146_,
		_w5147_,
		_w5148_
	);
	LUT2 #(
		.INIT('h4)
	) name4687 (
		_w5145_,
		_w5148_,
		_w5149_
	);
	LUT2 #(
		.INIT('h4)
	) name4688 (
		_w5139_,
		_w5149_,
		_w5150_
	);
	LUT2 #(
		.INIT('h4)
	) name4689 (
		_w5142_,
		_w5150_,
		_w5151_
	);
	LUT2 #(
		.INIT('h4)
	) name4690 (
		_w5136_,
		_w5151_,
		_w5152_
	);
	LUT2 #(
		.INIT('h2)
	) name4691 (
		_w2026_,
		_w5152_,
		_w5153_
	);
	LUT2 #(
		.INIT('h8)
	) name4692 (
		\P2_reg1_reg[27]/NET0131 ,
		_w2024_,
		_w5154_
	);
	LUT2 #(
		.INIT('h1)
	) name4693 (
		_w5153_,
		_w5154_,
		_w5155_
	);
	LUT2 #(
		.INIT('h2)
	) name4694 (
		\P1_state_reg[0]/NET0131 ,
		_w5155_,
		_w5156_
	);
	LUT2 #(
		.INIT('h2)
	) name4695 (
		\P2_reg1_reg[27]/NET0131 ,
		_w1983_,
		_w5157_
	);
	LUT2 #(
		.INIT('h1)
	) name4696 (
		_w5156_,
		_w5157_,
		_w5158_
	);
	LUT2 #(
		.INIT('h2)
	) name4697 (
		\P1_reg2_reg[24]/NET0131 ,
		_w3435_,
		_w5159_
	);
	LUT2 #(
		.INIT('h8)
	) name4698 (
		\P1_reg2_reg[24]/NET0131 ,
		_w3448_,
		_w5160_
	);
	LUT2 #(
		.INIT('h2)
	) name4699 (
		\P1_reg2_reg[24]/NET0131 ,
		_w3466_,
		_w5161_
	);
	LUT2 #(
		.INIT('h8)
	) name4700 (
		_w4000_,
		_w4014_,
		_w5162_
	);
	LUT2 #(
		.INIT('h4)
	) name4701 (
		_w4006_,
		_w4010_,
		_w5163_
	);
	LUT2 #(
		.INIT('h2)
	) name4702 (
		_w4021_,
		_w5163_,
		_w5164_
	);
	LUT2 #(
		.INIT('h2)
	) name4703 (
		_w4013_,
		_w5164_,
		_w5165_
	);
	LUT2 #(
		.INIT('h2)
	) name4704 (
		_w4028_,
		_w5165_,
		_w5166_
	);
	LUT2 #(
		.INIT('h4)
	) name4705 (
		_w5162_,
		_w5166_,
		_w5167_
	);
	LUT2 #(
		.INIT('h2)
	) name4706 (
		_w4033_,
		_w5167_,
		_w5168_
	);
	LUT2 #(
		.INIT('h2)
	) name4707 (
		_w4043_,
		_w5168_,
		_w5169_
	);
	LUT2 #(
		.INIT('h8)
	) name4708 (
		_w1818_,
		_w5169_,
		_w5170_
	);
	LUT2 #(
		.INIT('h1)
	) name4709 (
		_w1818_,
		_w5169_,
		_w5171_
	);
	LUT2 #(
		.INIT('h1)
	) name4710 (
		_w5170_,
		_w5171_,
		_w5172_
	);
	LUT2 #(
		.INIT('h2)
	) name4711 (
		_w3466_,
		_w5172_,
		_w5173_
	);
	LUT2 #(
		.INIT('h1)
	) name4712 (
		_w5161_,
		_w5173_,
		_w5174_
	);
	LUT2 #(
		.INIT('h1)
	) name4713 (
		_w3563_,
		_w5174_,
		_w5175_
	);
	LUT2 #(
		.INIT('h8)
	) name4714 (
		_w1479_,
		_w1749_,
		_w5176_
	);
	LUT2 #(
		.INIT('h2)
	) name4715 (
		_w1478_,
		_w1489_,
		_w5177_
	);
	LUT2 #(
		.INIT('h2)
	) name4716 (
		_w1720_,
		_w5177_,
		_w5178_
	);
	LUT2 #(
		.INIT('h2)
	) name4717 (
		_w1377_,
		_w5178_,
		_w5179_
	);
	LUT2 #(
		.INIT('h2)
	) name4718 (
		_w1710_,
		_w5176_,
		_w5180_
	);
	LUT2 #(
		.INIT('h4)
	) name4719 (
		_w5179_,
		_w5180_,
		_w5181_
	);
	LUT2 #(
		.INIT('h2)
	) name4720 (
		_w1818_,
		_w5181_,
		_w5182_
	);
	LUT2 #(
		.INIT('h4)
	) name4721 (
		_w1818_,
		_w5181_,
		_w5183_
	);
	LUT2 #(
		.INIT('h1)
	) name4722 (
		_w5182_,
		_w5183_,
		_w5184_
	);
	LUT2 #(
		.INIT('h2)
	) name4723 (
		_w3466_,
		_w5184_,
		_w5185_
	);
	LUT2 #(
		.INIT('h1)
	) name4724 (
		_w5161_,
		_w5185_,
		_w5186_
	);
	LUT2 #(
		.INIT('h1)
	) name4725 (
		_w3677_,
		_w5186_,
		_w5187_
	);
	LUT2 #(
		.INIT('h4)
	) name4726 (
		_w1327_,
		_w3700_,
		_w5188_
	);
	LUT2 #(
		.INIT('h2)
	) name4727 (
		_w1047_,
		_w5188_,
		_w5189_
	);
	LUT2 #(
		.INIT('h1)
	) name4728 (
		_w4686_,
		_w5189_,
		_w5190_
	);
	LUT2 #(
		.INIT('h8)
	) name4729 (
		_w3466_,
		_w5190_,
		_w5191_
	);
	LUT2 #(
		.INIT('h1)
	) name4730 (
		_w5161_,
		_w5191_,
		_w5192_
	);
	LUT2 #(
		.INIT('h2)
	) name4731 (
		_w3712_,
		_w5192_,
		_w5193_
	);
	LUT2 #(
		.INIT('h2)
	) name4732 (
		_w1038_,
		_w4075_,
		_w5194_
	);
	LUT2 #(
		.INIT('h8)
	) name4733 (
		_w3568_,
		_w4470_,
		_w5195_
	);
	LUT2 #(
		.INIT('h8)
	) name4734 (
		_w3592_,
		_w5195_,
		_w5196_
	);
	LUT2 #(
		.INIT('h1)
	) name4735 (
		_w5194_,
		_w5196_,
		_w5197_
	);
	LUT2 #(
		.INIT('h1)
	) name4736 (
		_w537_,
		_w5197_,
		_w5198_
	);
	LUT2 #(
		.INIT('h8)
	) name4737 (
		_w537_,
		_w1336_,
		_w5199_
	);
	LUT2 #(
		.INIT('h1)
	) name4738 (
		_w5198_,
		_w5199_,
		_w5200_
	);
	LUT2 #(
		.INIT('h8)
	) name4739 (
		_w3466_,
		_w5200_,
		_w5201_
	);
	LUT2 #(
		.INIT('h1)
	) name4740 (
		_w5161_,
		_w5201_,
		_w5202_
	);
	LUT2 #(
		.INIT('h2)
	) name4741 (
		_w1936_,
		_w5202_,
		_w5203_
	);
	LUT2 #(
		.INIT('h2)
	) name4742 (
		\P1_reg2_reg[24]/NET0131 ,
		_w3718_,
		_w5204_
	);
	LUT2 #(
		.INIT('h8)
	) name4743 (
		_w1058_,
		_w1763_,
		_w5205_
	);
	LUT2 #(
		.INIT('h8)
	) name4744 (
		_w1047_,
		_w1880_,
		_w5206_
	);
	LUT2 #(
		.INIT('h8)
	) name4745 (
		_w3466_,
		_w5206_,
		_w5207_
	);
	LUT2 #(
		.INIT('h1)
	) name4746 (
		_w5204_,
		_w5205_,
		_w5208_
	);
	LUT2 #(
		.INIT('h4)
	) name4747 (
		_w5207_,
		_w5208_,
		_w5209_
	);
	LUT2 #(
		.INIT('h4)
	) name4748 (
		_w5193_,
		_w5209_,
		_w5210_
	);
	LUT2 #(
		.INIT('h4)
	) name4749 (
		_w5175_,
		_w5210_,
		_w5211_
	);
	LUT2 #(
		.INIT('h1)
	) name4750 (
		_w5187_,
		_w5203_,
		_w5212_
	);
	LUT2 #(
		.INIT('h8)
	) name4751 (
		_w5211_,
		_w5212_,
		_w5213_
	);
	LUT2 #(
		.INIT('h2)
	) name4752 (
		_w3450_,
		_w5213_,
		_w5214_
	);
	LUT2 #(
		.INIT('h1)
	) name4753 (
		_w5160_,
		_w5214_,
		_w5215_
	);
	LUT2 #(
		.INIT('h2)
	) name4754 (
		\P1_state_reg[0]/NET0131 ,
		_w5215_,
		_w5216_
	);
	LUT2 #(
		.INIT('h1)
	) name4755 (
		_w5159_,
		_w5216_,
		_w5217_
	);
	LUT2 #(
		.INIT('h2)
	) name4756 (
		\P1_reg2_reg[28]/NET0131 ,
		_w3435_,
		_w5218_
	);
	LUT2 #(
		.INIT('h8)
	) name4757 (
		\P1_reg2_reg[28]/NET0131 ,
		_w3448_,
		_w5219_
	);
	LUT2 #(
		.INIT('h2)
	) name4758 (
		\P1_reg2_reg[28]/NET0131 ,
		_w3466_,
		_w5220_
	);
	LUT2 #(
		.INIT('h2)
	) name4759 (
		_w3466_,
		_w4101_,
		_w5221_
	);
	LUT2 #(
		.INIT('h1)
	) name4760 (
		_w5220_,
		_w5221_,
		_w5222_
	);
	LUT2 #(
		.INIT('h1)
	) name4761 (
		_w3677_,
		_w5222_,
		_w5223_
	);
	LUT2 #(
		.INIT('h8)
	) name4762 (
		_w3466_,
		_w4059_,
		_w5224_
	);
	LUT2 #(
		.INIT('h1)
	) name4763 (
		_w5220_,
		_w5224_,
		_w5225_
	);
	LUT2 #(
		.INIT('h2)
	) name4764 (
		_w3712_,
		_w5225_,
		_w5226_
	);
	LUT2 #(
		.INIT('h2)
	) name4765 (
		\P1_reg2_reg[28]/NET0131 ,
		_w3718_,
		_w5227_
	);
	LUT2 #(
		.INIT('h8)
	) name4766 (
		_w941_,
		_w1763_,
		_w5228_
	);
	LUT2 #(
		.INIT('h8)
	) name4767 (
		_w933_,
		_w1880_,
		_w5229_
	);
	LUT2 #(
		.INIT('h8)
	) name4768 (
		_w3466_,
		_w5229_,
		_w5230_
	);
	LUT2 #(
		.INIT('h2)
	) name4769 (
		_w3466_,
		_w4084_,
		_w5231_
	);
	LUT2 #(
		.INIT('h1)
	) name4770 (
		_w5220_,
		_w5231_,
		_w5232_
	);
	LUT2 #(
		.INIT('h2)
	) name4771 (
		_w1936_,
		_w5232_,
		_w5233_
	);
	LUT2 #(
		.INIT('h2)
	) name4772 (
		_w3466_,
		_w4053_,
		_w5234_
	);
	LUT2 #(
		.INIT('h1)
	) name4773 (
		_w5220_,
		_w5234_,
		_w5235_
	);
	LUT2 #(
		.INIT('h1)
	) name4774 (
		_w3563_,
		_w5235_,
		_w5236_
	);
	LUT2 #(
		.INIT('h1)
	) name4775 (
		_w5227_,
		_w5228_,
		_w5237_
	);
	LUT2 #(
		.INIT('h4)
	) name4776 (
		_w5230_,
		_w5237_,
		_w5238_
	);
	LUT2 #(
		.INIT('h4)
	) name4777 (
		_w5226_,
		_w5238_,
		_w5239_
	);
	LUT2 #(
		.INIT('h4)
	) name4778 (
		_w5223_,
		_w5239_,
		_w5240_
	);
	LUT2 #(
		.INIT('h1)
	) name4779 (
		_w5233_,
		_w5236_,
		_w5241_
	);
	LUT2 #(
		.INIT('h8)
	) name4780 (
		_w5240_,
		_w5241_,
		_w5242_
	);
	LUT2 #(
		.INIT('h2)
	) name4781 (
		_w3450_,
		_w5242_,
		_w5243_
	);
	LUT2 #(
		.INIT('h1)
	) name4782 (
		_w5219_,
		_w5243_,
		_w5244_
	);
	LUT2 #(
		.INIT('h2)
	) name4783 (
		\P1_state_reg[0]/NET0131 ,
		_w5244_,
		_w5245_
	);
	LUT2 #(
		.INIT('h1)
	) name4784 (
		_w5218_,
		_w5245_,
		_w5246_
	);
	LUT2 #(
		.INIT('h2)
	) name4785 (
		\P2_reg2_reg[27]/NET0131 ,
		_w3758_,
		_w5247_
	);
	LUT2 #(
		.INIT('h8)
	) name4786 (
		_w3758_,
		_w4828_,
		_w5248_
	);
	LUT2 #(
		.INIT('h1)
	) name4787 (
		_w5247_,
		_w5248_,
		_w5249_
	);
	LUT2 #(
		.INIT('h1)
	) name4788 (
		_w3177_,
		_w5249_,
		_w5250_
	);
	LUT2 #(
		.INIT('h8)
	) name4789 (
		_w3758_,
		_w4869_,
		_w5251_
	);
	LUT2 #(
		.INIT('h1)
	) name4790 (
		_w5247_,
		_w5251_,
		_w5252_
	);
	LUT2 #(
		.INIT('h2)
	) name4791 (
		_w3355_,
		_w5252_,
		_w5253_
	);
	LUT2 #(
		.INIT('h2)
	) name4792 (
		_w3758_,
		_w4864_,
		_w5254_
	);
	LUT2 #(
		.INIT('h1)
	) name4793 (
		_w5247_,
		_w5254_,
		_w5255_
	);
	LUT2 #(
		.INIT('h1)
	) name4794 (
		_w3320_,
		_w5255_,
		_w5256_
	);
	LUT2 #(
		.INIT('h8)
	) name4795 (
		_w3758_,
		_w4877_,
		_w5257_
	);
	LUT2 #(
		.INIT('h1)
	) name4796 (
		_w5247_,
		_w5257_,
		_w5258_
	);
	LUT2 #(
		.INIT('h2)
	) name4797 (
		_w3411_,
		_w5258_,
		_w5259_
	);
	LUT2 #(
		.INIT('h8)
	) name4798 (
		_w3758_,
		_w5036_,
		_w5260_
	);
	LUT2 #(
		.INIT('h8)
	) name4799 (
		_w2987_,
		_w3420_,
		_w5261_
	);
	LUT2 #(
		.INIT('h2)
	) name4800 (
		\P2_reg2_reg[27]/NET0131 ,
		_w3774_,
		_w5262_
	);
	LUT2 #(
		.INIT('h1)
	) name4801 (
		_w5261_,
		_w5262_,
		_w5263_
	);
	LUT2 #(
		.INIT('h4)
	) name4802 (
		_w5260_,
		_w5263_,
		_w5264_
	);
	LUT2 #(
		.INIT('h4)
	) name4803 (
		_w5259_,
		_w5264_,
		_w5265_
	);
	LUT2 #(
		.INIT('h4)
	) name4804 (
		_w5253_,
		_w5265_,
		_w5266_
	);
	LUT2 #(
		.INIT('h4)
	) name4805 (
		_w5256_,
		_w5266_,
		_w5267_
	);
	LUT2 #(
		.INIT('h4)
	) name4806 (
		_w5250_,
		_w5267_,
		_w5268_
	);
	LUT2 #(
		.INIT('h2)
	) name4807 (
		_w2026_,
		_w5268_,
		_w5269_
	);
	LUT2 #(
		.INIT('h8)
	) name4808 (
		\P2_reg2_reg[27]/NET0131 ,
		_w2024_,
		_w5270_
	);
	LUT2 #(
		.INIT('h1)
	) name4809 (
		_w5269_,
		_w5270_,
		_w5271_
	);
	LUT2 #(
		.INIT('h2)
	) name4810 (
		\P1_state_reg[0]/NET0131 ,
		_w5271_,
		_w5272_
	);
	LUT2 #(
		.INIT('h2)
	) name4811 (
		\P2_reg2_reg[27]/NET0131 ,
		_w1983_,
		_w5273_
	);
	LUT2 #(
		.INIT('h1)
	) name4812 (
		_w5272_,
		_w5273_,
		_w5274_
	);
	LUT2 #(
		.INIT('h8)
	) name4813 (
		_w3358_,
		_w4141_,
		_w5275_
	);
	LUT2 #(
		.INIT('h4)
	) name4814 (
		_w3372_,
		_w3411_,
		_w5276_
	);
	LUT2 #(
		.INIT('h8)
	) name4815 (
		_w3407_,
		_w5276_,
		_w5277_
	);
	LUT2 #(
		.INIT('h1)
	) name4816 (
		_w5275_,
		_w5277_,
		_w5278_
	);
	LUT2 #(
		.INIT('h2)
	) name4817 (
		_w3350_,
		_w4159_,
		_w5279_
	);
	LUT2 #(
		.INIT('h2)
	) name4818 (
		_w4141_,
		_w5279_,
		_w5280_
	);
	LUT2 #(
		.INIT('h4)
	) name4819 (
		_w4141_,
		_w5279_,
		_w5281_
	);
	LUT2 #(
		.INIT('h1)
	) name4820 (
		_w5280_,
		_w5281_,
		_w5282_
	);
	LUT2 #(
		.INIT('h8)
	) name4821 (
		_w3354_,
		_w5282_,
		_w5283_
	);
	LUT2 #(
		.INIT('h2)
	) name4822 (
		_w5278_,
		_w5283_,
		_w5284_
	);
	LUT2 #(
		.INIT('h2)
	) name4823 (
		_w3758_,
		_w5284_,
		_w5285_
	);
	LUT2 #(
		.INIT('h1)
	) name4824 (
		_w3776_,
		_w5285_,
		_w5286_
	);
	LUT2 #(
		.INIT('h2)
	) name4825 (
		_w1983_,
		_w2023_,
		_w5287_
	);
	LUT2 #(
		.INIT('h4)
	) name4826 (
		_w5286_,
		_w5287_,
		_w5288_
	);
	LUT2 #(
		.INIT('h1)
	) name4827 (
		_w3357_,
		_w3758_,
		_w5289_
	);
	LUT2 #(
		.INIT('h2)
	) name4828 (
		_w3774_,
		_w5289_,
		_w5290_
	);
	LUT2 #(
		.INIT('h4)
	) name4829 (
		_w4381_,
		_w5287_,
		_w5291_
	);
	LUT2 #(
		.INIT('h8)
	) name4830 (
		_w5290_,
		_w5291_,
		_w5292_
	);
	LUT2 #(
		.INIT('h2)
	) name4831 (
		\P2_reg2_reg[31]/NET0131 ,
		_w5292_,
		_w5293_
	);
	LUT2 #(
		.INIT('h1)
	) name4832 (
		_w5288_,
		_w5293_,
		_w5294_
	);
	LUT2 #(
		.INIT('h2)
	) name4833 (
		\P1_reg0_reg[25]/NET0131 ,
		_w3435_,
		_w5295_
	);
	LUT2 #(
		.INIT('h8)
	) name4834 (
		\P1_reg0_reg[25]/NET0131 ,
		_w3448_,
		_w5296_
	);
	LUT2 #(
		.INIT('h2)
	) name4835 (
		\P1_reg0_reg[25]/NET0131 ,
		_w4396_,
		_w5297_
	);
	LUT2 #(
		.INIT('h2)
	) name4836 (
		_w4396_,
		_w4658_,
		_w5298_
	);
	LUT2 #(
		.INIT('h1)
	) name4837 (
		_w5297_,
		_w5298_,
		_w5299_
	);
	LUT2 #(
		.INIT('h1)
	) name4838 (
		_w3677_,
		_w5299_,
		_w5300_
	);
	LUT2 #(
		.INIT('h2)
	) name4839 (
		_w4396_,
		_w4672_,
		_w5301_
	);
	LUT2 #(
		.INIT('h1)
	) name4840 (
		_w5297_,
		_w5301_,
		_w5302_
	);
	LUT2 #(
		.INIT('h1)
	) name4841 (
		_w3563_,
		_w5302_,
		_w5303_
	);
	LUT2 #(
		.INIT('h8)
	) name4842 (
		_w1029_,
		_w1880_,
		_w5304_
	);
	LUT2 #(
		.INIT('h8)
	) name4843 (
		_w4396_,
		_w5304_,
		_w5305_
	);
	LUT2 #(
		.INIT('h2)
	) name4844 (
		\P1_reg0_reg[25]/NET0131 ,
		_w4493_,
		_w5306_
	);
	LUT2 #(
		.INIT('h8)
	) name4845 (
		_w4396_,
		_w4682_,
		_w5307_
	);
	LUT2 #(
		.INIT('h1)
	) name4846 (
		_w5297_,
		_w5307_,
		_w5308_
	);
	LUT2 #(
		.INIT('h2)
	) name4847 (
		_w1936_,
		_w5308_,
		_w5309_
	);
	LUT2 #(
		.INIT('h8)
	) name4848 (
		_w4396_,
		_w4689_,
		_w5310_
	);
	LUT2 #(
		.INIT('h1)
	) name4849 (
		_w5297_,
		_w5310_,
		_w5311_
	);
	LUT2 #(
		.INIT('h2)
	) name4850 (
		_w3712_,
		_w5311_,
		_w5312_
	);
	LUT2 #(
		.INIT('h1)
	) name4851 (
		_w5305_,
		_w5306_,
		_w5313_
	);
	LUT2 #(
		.INIT('h4)
	) name4852 (
		_w5309_,
		_w5313_,
		_w5314_
	);
	LUT2 #(
		.INIT('h4)
	) name4853 (
		_w5312_,
		_w5314_,
		_w5315_
	);
	LUT2 #(
		.INIT('h1)
	) name4854 (
		_w5300_,
		_w5303_,
		_w5316_
	);
	LUT2 #(
		.INIT('h8)
	) name4855 (
		_w5315_,
		_w5316_,
		_w5317_
	);
	LUT2 #(
		.INIT('h2)
	) name4856 (
		_w3450_,
		_w5317_,
		_w5318_
	);
	LUT2 #(
		.INIT('h1)
	) name4857 (
		_w5296_,
		_w5318_,
		_w5319_
	);
	LUT2 #(
		.INIT('h2)
	) name4858 (
		\P1_state_reg[0]/NET0131 ,
		_w5319_,
		_w5320_
	);
	LUT2 #(
		.INIT('h1)
	) name4859 (
		_w5295_,
		_w5320_,
		_w5321_
	);
	LUT2 #(
		.INIT('h8)
	) name4860 (
		\P1_reg0_reg[28]/NET0131 ,
		_w3448_,
		_w5322_
	);
	LUT2 #(
		.INIT('h2)
	) name4861 (
		\P1_reg0_reg[28]/NET0131 ,
		_w4396_,
		_w5323_
	);
	LUT2 #(
		.INIT('h4)
	) name4862 (
		_w4101_,
		_w4396_,
		_w5324_
	);
	LUT2 #(
		.INIT('h1)
	) name4863 (
		_w5323_,
		_w5324_,
		_w5325_
	);
	LUT2 #(
		.INIT('h1)
	) name4864 (
		_w3677_,
		_w5325_,
		_w5326_
	);
	LUT2 #(
		.INIT('h8)
	) name4865 (
		_w4059_,
		_w4396_,
		_w5327_
	);
	LUT2 #(
		.INIT('h1)
	) name4866 (
		_w5323_,
		_w5327_,
		_w5328_
	);
	LUT2 #(
		.INIT('h2)
	) name4867 (
		_w3712_,
		_w5328_,
		_w5329_
	);
	LUT2 #(
		.INIT('h2)
	) name4868 (
		\P1_reg0_reg[28]/NET0131 ,
		_w4493_,
		_w5330_
	);
	LUT2 #(
		.INIT('h8)
	) name4869 (
		_w4396_,
		_w5229_,
		_w5331_
	);
	LUT2 #(
		.INIT('h4)
	) name4870 (
		_w4084_,
		_w4396_,
		_w5332_
	);
	LUT2 #(
		.INIT('h1)
	) name4871 (
		_w5323_,
		_w5332_,
		_w5333_
	);
	LUT2 #(
		.INIT('h2)
	) name4872 (
		_w1936_,
		_w5333_,
		_w5334_
	);
	LUT2 #(
		.INIT('h4)
	) name4873 (
		_w4053_,
		_w4396_,
		_w5335_
	);
	LUT2 #(
		.INIT('h1)
	) name4874 (
		_w5323_,
		_w5335_,
		_w5336_
	);
	LUT2 #(
		.INIT('h1)
	) name4875 (
		_w3563_,
		_w5336_,
		_w5337_
	);
	LUT2 #(
		.INIT('h1)
	) name4876 (
		_w5330_,
		_w5331_,
		_w5338_
	);
	LUT2 #(
		.INIT('h4)
	) name4877 (
		_w5329_,
		_w5338_,
		_w5339_
	);
	LUT2 #(
		.INIT('h4)
	) name4878 (
		_w5326_,
		_w5339_,
		_w5340_
	);
	LUT2 #(
		.INIT('h1)
	) name4879 (
		_w5334_,
		_w5337_,
		_w5341_
	);
	LUT2 #(
		.INIT('h8)
	) name4880 (
		_w5340_,
		_w5341_,
		_w5342_
	);
	LUT2 #(
		.INIT('h2)
	) name4881 (
		_w3450_,
		_w5342_,
		_w5343_
	);
	LUT2 #(
		.INIT('h1)
	) name4882 (
		_w5322_,
		_w5343_,
		_w5344_
	);
	LUT2 #(
		.INIT('h2)
	) name4883 (
		\P1_state_reg[0]/NET0131 ,
		_w5344_,
		_w5345_
	);
	LUT2 #(
		.INIT('h2)
	) name4884 (
		\P1_reg0_reg[28]/NET0131 ,
		_w3435_,
		_w5346_
	);
	LUT2 #(
		.INIT('h1)
	) name4885 (
		_w5345_,
		_w5346_,
		_w5347_
	);
	LUT2 #(
		.INIT('h2)
	) name4886 (
		\P1_reg1_reg[24]/NET0131 ,
		_w3435_,
		_w5348_
	);
	LUT2 #(
		.INIT('h8)
	) name4887 (
		\P1_reg1_reg[24]/NET0131 ,
		_w3448_,
		_w5349_
	);
	LUT2 #(
		.INIT('h2)
	) name4888 (
		\P1_reg1_reg[24]/NET0131 ,
		_w4532_,
		_w5350_
	);
	LUT2 #(
		.INIT('h2)
	) name4889 (
		_w4532_,
		_w5172_,
		_w5351_
	);
	LUT2 #(
		.INIT('h1)
	) name4890 (
		_w5350_,
		_w5351_,
		_w5352_
	);
	LUT2 #(
		.INIT('h1)
	) name4891 (
		_w3563_,
		_w5352_,
		_w5353_
	);
	LUT2 #(
		.INIT('h8)
	) name4892 (
		_w4532_,
		_w5200_,
		_w5354_
	);
	LUT2 #(
		.INIT('h1)
	) name4893 (
		_w5350_,
		_w5354_,
		_w5355_
	);
	LUT2 #(
		.INIT('h2)
	) name4894 (
		_w1936_,
		_w5355_,
		_w5356_
	);
	LUT2 #(
		.INIT('h2)
	) name4895 (
		\P1_reg1_reg[24]/NET0131 ,
		_w4541_,
		_w5357_
	);
	LUT2 #(
		.INIT('h8)
	) name4896 (
		_w4532_,
		_w5206_,
		_w5358_
	);
	LUT2 #(
		.INIT('h8)
	) name4897 (
		_w4532_,
		_w5190_,
		_w5359_
	);
	LUT2 #(
		.INIT('h1)
	) name4898 (
		_w5350_,
		_w5359_,
		_w5360_
	);
	LUT2 #(
		.INIT('h2)
	) name4899 (
		_w3712_,
		_w5360_,
		_w5361_
	);
	LUT2 #(
		.INIT('h2)
	) name4900 (
		_w4532_,
		_w5184_,
		_w5362_
	);
	LUT2 #(
		.INIT('h1)
	) name4901 (
		_w5350_,
		_w5362_,
		_w5363_
	);
	LUT2 #(
		.INIT('h1)
	) name4902 (
		_w3677_,
		_w5363_,
		_w5364_
	);
	LUT2 #(
		.INIT('h1)
	) name4903 (
		_w5357_,
		_w5358_,
		_w5365_
	);
	LUT2 #(
		.INIT('h4)
	) name4904 (
		_w5361_,
		_w5365_,
		_w5366_
	);
	LUT2 #(
		.INIT('h4)
	) name4905 (
		_w5353_,
		_w5366_,
		_w5367_
	);
	LUT2 #(
		.INIT('h1)
	) name4906 (
		_w5356_,
		_w5364_,
		_w5368_
	);
	LUT2 #(
		.INIT('h8)
	) name4907 (
		_w5367_,
		_w5368_,
		_w5369_
	);
	LUT2 #(
		.INIT('h2)
	) name4908 (
		_w3450_,
		_w5369_,
		_w5370_
	);
	LUT2 #(
		.INIT('h1)
	) name4909 (
		_w5349_,
		_w5370_,
		_w5371_
	);
	LUT2 #(
		.INIT('h2)
	) name4910 (
		\P1_state_reg[0]/NET0131 ,
		_w5371_,
		_w5372_
	);
	LUT2 #(
		.INIT('h1)
	) name4911 (
		_w5348_,
		_w5372_,
		_w5373_
	);
	LUT2 #(
		.INIT('h2)
	) name4912 (
		\P1_reg1_reg[25]/NET0131 ,
		_w3435_,
		_w5374_
	);
	LUT2 #(
		.INIT('h8)
	) name4913 (
		\P1_reg1_reg[25]/NET0131 ,
		_w3448_,
		_w5375_
	);
	LUT2 #(
		.INIT('h2)
	) name4914 (
		\P1_reg1_reg[25]/NET0131 ,
		_w4532_,
		_w5376_
	);
	LUT2 #(
		.INIT('h2)
	) name4915 (
		_w4532_,
		_w4658_,
		_w5377_
	);
	LUT2 #(
		.INIT('h1)
	) name4916 (
		_w5376_,
		_w5377_,
		_w5378_
	);
	LUT2 #(
		.INIT('h1)
	) name4917 (
		_w3677_,
		_w5378_,
		_w5379_
	);
	LUT2 #(
		.INIT('h2)
	) name4918 (
		_w4532_,
		_w4672_,
		_w5380_
	);
	LUT2 #(
		.INIT('h1)
	) name4919 (
		_w5376_,
		_w5380_,
		_w5381_
	);
	LUT2 #(
		.INIT('h1)
	) name4920 (
		_w3563_,
		_w5381_,
		_w5382_
	);
	LUT2 #(
		.INIT('h8)
	) name4921 (
		_w4532_,
		_w5304_,
		_w5383_
	);
	LUT2 #(
		.INIT('h2)
	) name4922 (
		\P1_reg1_reg[25]/NET0131 ,
		_w4541_,
		_w5384_
	);
	LUT2 #(
		.INIT('h8)
	) name4923 (
		_w4532_,
		_w4682_,
		_w5385_
	);
	LUT2 #(
		.INIT('h1)
	) name4924 (
		_w5376_,
		_w5385_,
		_w5386_
	);
	LUT2 #(
		.INIT('h2)
	) name4925 (
		_w1936_,
		_w5386_,
		_w5387_
	);
	LUT2 #(
		.INIT('h8)
	) name4926 (
		_w4532_,
		_w4689_,
		_w5388_
	);
	LUT2 #(
		.INIT('h1)
	) name4927 (
		_w5376_,
		_w5388_,
		_w5389_
	);
	LUT2 #(
		.INIT('h2)
	) name4928 (
		_w3712_,
		_w5389_,
		_w5390_
	);
	LUT2 #(
		.INIT('h1)
	) name4929 (
		_w5383_,
		_w5384_,
		_w5391_
	);
	LUT2 #(
		.INIT('h4)
	) name4930 (
		_w5387_,
		_w5391_,
		_w5392_
	);
	LUT2 #(
		.INIT('h4)
	) name4931 (
		_w5390_,
		_w5392_,
		_w5393_
	);
	LUT2 #(
		.INIT('h1)
	) name4932 (
		_w5379_,
		_w5382_,
		_w5394_
	);
	LUT2 #(
		.INIT('h8)
	) name4933 (
		_w5393_,
		_w5394_,
		_w5395_
	);
	LUT2 #(
		.INIT('h2)
	) name4934 (
		_w3450_,
		_w5395_,
		_w5396_
	);
	LUT2 #(
		.INIT('h1)
	) name4935 (
		_w5375_,
		_w5396_,
		_w5397_
	);
	LUT2 #(
		.INIT('h2)
	) name4936 (
		\P1_state_reg[0]/NET0131 ,
		_w5397_,
		_w5398_
	);
	LUT2 #(
		.INIT('h1)
	) name4937 (
		_w5374_,
		_w5398_,
		_w5399_
	);
	LUT2 #(
		.INIT('h8)
	) name4938 (
		\P1_reg1_reg[28]/NET0131 ,
		_w3448_,
		_w5400_
	);
	LUT2 #(
		.INIT('h2)
	) name4939 (
		\P1_reg1_reg[28]/NET0131 ,
		_w4532_,
		_w5401_
	);
	LUT2 #(
		.INIT('h4)
	) name4940 (
		_w4101_,
		_w4532_,
		_w5402_
	);
	LUT2 #(
		.INIT('h1)
	) name4941 (
		_w5401_,
		_w5402_,
		_w5403_
	);
	LUT2 #(
		.INIT('h1)
	) name4942 (
		_w3677_,
		_w5403_,
		_w5404_
	);
	LUT2 #(
		.INIT('h8)
	) name4943 (
		_w4059_,
		_w4532_,
		_w5405_
	);
	LUT2 #(
		.INIT('h1)
	) name4944 (
		_w5401_,
		_w5405_,
		_w5406_
	);
	LUT2 #(
		.INIT('h2)
	) name4945 (
		_w3712_,
		_w5406_,
		_w5407_
	);
	LUT2 #(
		.INIT('h2)
	) name4946 (
		\P1_reg1_reg[28]/NET0131 ,
		_w4541_,
		_w5408_
	);
	LUT2 #(
		.INIT('h8)
	) name4947 (
		_w4532_,
		_w5229_,
		_w5409_
	);
	LUT2 #(
		.INIT('h4)
	) name4948 (
		_w4084_,
		_w4532_,
		_w5410_
	);
	LUT2 #(
		.INIT('h1)
	) name4949 (
		_w5401_,
		_w5410_,
		_w5411_
	);
	LUT2 #(
		.INIT('h2)
	) name4950 (
		_w1936_,
		_w5411_,
		_w5412_
	);
	LUT2 #(
		.INIT('h4)
	) name4951 (
		_w4053_,
		_w4532_,
		_w5413_
	);
	LUT2 #(
		.INIT('h1)
	) name4952 (
		_w5401_,
		_w5413_,
		_w5414_
	);
	LUT2 #(
		.INIT('h1)
	) name4953 (
		_w3563_,
		_w5414_,
		_w5415_
	);
	LUT2 #(
		.INIT('h1)
	) name4954 (
		_w5408_,
		_w5409_,
		_w5416_
	);
	LUT2 #(
		.INIT('h4)
	) name4955 (
		_w5407_,
		_w5416_,
		_w5417_
	);
	LUT2 #(
		.INIT('h4)
	) name4956 (
		_w5404_,
		_w5417_,
		_w5418_
	);
	LUT2 #(
		.INIT('h1)
	) name4957 (
		_w5412_,
		_w5415_,
		_w5419_
	);
	LUT2 #(
		.INIT('h8)
	) name4958 (
		_w5418_,
		_w5419_,
		_w5420_
	);
	LUT2 #(
		.INIT('h2)
	) name4959 (
		_w3450_,
		_w5420_,
		_w5421_
	);
	LUT2 #(
		.INIT('h1)
	) name4960 (
		_w5400_,
		_w5421_,
		_w5422_
	);
	LUT2 #(
		.INIT('h2)
	) name4961 (
		\P1_state_reg[0]/NET0131 ,
		_w5422_,
		_w5423_
	);
	LUT2 #(
		.INIT('h2)
	) name4962 (
		\P1_reg1_reg[28]/NET0131 ,
		_w3435_,
		_w5424_
	);
	LUT2 #(
		.INIT('h1)
	) name4963 (
		_w5423_,
		_w5424_,
		_w5425_
	);
	LUT2 #(
		.INIT('h2)
	) name4964 (
		\P1_reg3_reg[17]/NET0131 ,
		\P1_state_reg[0]/NET0131 ,
		_w5426_
	);
	LUT2 #(
		.INIT('h8)
	) name4965 (
		_w1447_,
		_w1953_,
		_w5427_
	);
	LUT2 #(
		.INIT('h8)
	) name4966 (
		_w1447_,
		_w3448_,
		_w5428_
	);
	LUT2 #(
		.INIT('h2)
	) name4967 (
		_w1447_,
		_w4064_,
		_w5429_
	);
	LUT2 #(
		.INIT('h2)
	) name4968 (
		_w1443_,
		_w4067_,
		_w5430_
	);
	LUT2 #(
		.INIT('h2)
	) name4969 (
		_w1447_,
		_w3980_,
		_w5431_
	);
	LUT2 #(
		.INIT('h2)
	) name4970 (
		_w3625_,
		_w3650_,
		_w5432_
	);
	LUT2 #(
		.INIT('h2)
	) name4971 (
		_w3656_,
		_w5432_,
		_w5433_
	);
	LUT2 #(
		.INIT('h2)
	) name4972 (
		_w1825_,
		_w5433_,
		_w5434_
	);
	LUT2 #(
		.INIT('h4)
	) name4973 (
		_w1825_,
		_w5433_,
		_w5435_
	);
	LUT2 #(
		.INIT('h1)
	) name4974 (
		_w5434_,
		_w5435_,
		_w5436_
	);
	LUT2 #(
		.INIT('h8)
	) name4975 (
		_w3980_,
		_w5436_,
		_w5437_
	);
	LUT2 #(
		.INIT('h1)
	) name4976 (
		_w5431_,
		_w5437_,
		_w5438_
	);
	LUT2 #(
		.INIT('h1)
	) name4977 (
		_w3677_,
		_w5438_,
		_w5439_
	);
	LUT2 #(
		.INIT('h4)
	) name4978 (
		_w1136_,
		_w3690_,
		_w5440_
	);
	LUT2 #(
		.INIT('h8)
	) name4979 (
		_w3691_,
		_w5440_,
		_w5441_
	);
	LUT2 #(
		.INIT('h4)
	) name4980 (
		_w1466_,
		_w5441_,
		_w5442_
	);
	LUT2 #(
		.INIT('h2)
	) name4981 (
		_w1443_,
		_w5442_,
		_w5443_
	);
	LUT2 #(
		.INIT('h4)
	) name4982 (
		_w1443_,
		_w5442_,
		_w5444_
	);
	LUT2 #(
		.INIT('h1)
	) name4983 (
		_w5443_,
		_w5444_,
		_w5445_
	);
	LUT2 #(
		.INIT('h8)
	) name4984 (
		_w3980_,
		_w5445_,
		_w5446_
	);
	LUT2 #(
		.INIT('h1)
	) name4985 (
		_w5431_,
		_w5446_,
		_w5447_
	);
	LUT2 #(
		.INIT('h2)
	) name4986 (
		_w3712_,
		_w5447_,
		_w5448_
	);
	LUT2 #(
		.INIT('h2)
	) name4987 (
		_w3490_,
		_w3533_,
		_w5449_
	);
	LUT2 #(
		.INIT('h2)
	) name4988 (
		_w3540_,
		_w5449_,
		_w5450_
	);
	LUT2 #(
		.INIT('h2)
	) name4989 (
		_w1825_,
		_w5450_,
		_w5451_
	);
	LUT2 #(
		.INIT('h4)
	) name4990 (
		_w1825_,
		_w5450_,
		_w5452_
	);
	LUT2 #(
		.INIT('h1)
	) name4991 (
		_w5451_,
		_w5452_,
		_w5453_
	);
	LUT2 #(
		.INIT('h2)
	) name4992 (
		_w3980_,
		_w5453_,
		_w5454_
	);
	LUT2 #(
		.INIT('h1)
	) name4993 (
		_w5431_,
		_w5454_,
		_w5455_
	);
	LUT2 #(
		.INIT('h1)
	) name4994 (
		_w3563_,
		_w5455_,
		_w5456_
	);
	LUT2 #(
		.INIT('h2)
	) name4995 (
		_w1403_,
		_w3585_,
		_w5457_
	);
	LUT2 #(
		.INIT('h4)
	) name4996 (
		_w1403_,
		_w3585_,
		_w5458_
	);
	LUT2 #(
		.INIT('h1)
	) name4997 (
		_w5457_,
		_w5458_,
		_w5459_
	);
	LUT2 #(
		.INIT('h1)
	) name4998 (
		_w537_,
		_w5459_,
		_w5460_
	);
	LUT2 #(
		.INIT('h8)
	) name4999 (
		_w537_,
		_w1475_,
		_w5461_
	);
	LUT2 #(
		.INIT('h1)
	) name5000 (
		_w5460_,
		_w5461_,
		_w5462_
	);
	LUT2 #(
		.INIT('h8)
	) name5001 (
		_w3980_,
		_w5462_,
		_w5463_
	);
	LUT2 #(
		.INIT('h1)
	) name5002 (
		_w5431_,
		_w5463_,
		_w5464_
	);
	LUT2 #(
		.INIT('h2)
	) name5003 (
		_w1936_,
		_w5464_,
		_w5465_
	);
	LUT2 #(
		.INIT('h1)
	) name5004 (
		_w5429_,
		_w5430_,
		_w5466_
	);
	LUT2 #(
		.INIT('h4)
	) name5005 (
		_w5448_,
		_w5466_,
		_w5467_
	);
	LUT2 #(
		.INIT('h4)
	) name5006 (
		_w5465_,
		_w5467_,
		_w5468_
	);
	LUT2 #(
		.INIT('h1)
	) name5007 (
		_w5439_,
		_w5456_,
		_w5469_
	);
	LUT2 #(
		.INIT('h8)
	) name5008 (
		_w5468_,
		_w5469_,
		_w5470_
	);
	LUT2 #(
		.INIT('h2)
	) name5009 (
		_w3450_,
		_w5470_,
		_w5471_
	);
	LUT2 #(
		.INIT('h1)
	) name5010 (
		_w5428_,
		_w5471_,
		_w5472_
	);
	LUT2 #(
		.INIT('h2)
	) name5011 (
		\P1_state_reg[0]/NET0131 ,
		_w5472_,
		_w5473_
	);
	LUT2 #(
		.INIT('h1)
	) name5012 (
		_w5426_,
		_w5427_,
		_w5474_
	);
	LUT2 #(
		.INIT('h4)
	) name5013 (
		_w5473_,
		_w5474_,
		_w5475_
	);
	LUT2 #(
		.INIT('h8)
	) name5014 (
		_w1399_,
		_w1953_,
		_w5476_
	);
	LUT2 #(
		.INIT('h2)
	) name5015 (
		\P1_reg3_reg[18]/NET0131 ,
		\P1_state_reg[0]/NET0131 ,
		_w5477_
	);
	LUT2 #(
		.INIT('h8)
	) name5016 (
		_w1399_,
		_w3448_,
		_w5478_
	);
	LUT2 #(
		.INIT('h2)
	) name5017 (
		_w1399_,
		_w4064_,
		_w5479_
	);
	LUT2 #(
		.INIT('h2)
	) name5018 (
		_w1399_,
		_w3980_,
		_w5480_
	);
	LUT2 #(
		.INIT('h2)
	) name5019 (
		_w1394_,
		_w5444_,
		_w5481_
	);
	LUT2 #(
		.INIT('h1)
	) name5020 (
		_w3696_,
		_w5481_,
		_w5482_
	);
	LUT2 #(
		.INIT('h8)
	) name5021 (
		_w3980_,
		_w5482_,
		_w5483_
	);
	LUT2 #(
		.INIT('h1)
	) name5022 (
		_w5480_,
		_w5483_,
		_w5484_
	);
	LUT2 #(
		.INIT('h2)
	) name5023 (
		_w3712_,
		_w5484_,
		_w5485_
	);
	LUT2 #(
		.INIT('h8)
	) name5024 (
		_w1120_,
		_w1477_,
		_w5486_
	);
	LUT2 #(
		.INIT('h8)
	) name5025 (
		_w1283_,
		_w1539_,
		_w5487_
	);
	LUT2 #(
		.INIT('h4)
	) name5026 (
		_w1686_,
		_w5487_,
		_w5488_
	);
	LUT2 #(
		.INIT('h2)
	) name5027 (
		_w1283_,
		_w1691_,
		_w5489_
	);
	LUT2 #(
		.INIT('h1)
	) name5028 (
		_w1483_,
		_w5489_,
		_w5490_
	);
	LUT2 #(
		.INIT('h4)
	) name5029 (
		_w5488_,
		_w5490_,
		_w5491_
	);
	LUT2 #(
		.INIT('h8)
	) name5030 (
		_w1235_,
		_w1291_,
		_w5492_
	);
	LUT2 #(
		.INIT('h4)
	) name5031 (
		_w5491_,
		_w5492_,
		_w5493_
	);
	LUT2 #(
		.INIT('h8)
	) name5032 (
		_w5486_,
		_w5493_,
		_w5494_
	);
	LUT2 #(
		.INIT('h8)
	) name5033 (
		_w1291_,
		_w1486_,
		_w5495_
	);
	LUT2 #(
		.INIT('h1)
	) name5034 (
		_w1177_,
		_w5495_,
		_w5496_
	);
	LUT2 #(
		.INIT('h2)
	) name5035 (
		_w5486_,
		_w5496_,
		_w5497_
	);
	LUT2 #(
		.INIT('h8)
	) name5036 (
		_w1182_,
		_w1477_,
		_w5498_
	);
	LUT2 #(
		.INIT('h1)
	) name5037 (
		_w1714_,
		_w5498_,
		_w5499_
	);
	LUT2 #(
		.INIT('h4)
	) name5038 (
		_w5497_,
		_w5499_,
		_w5500_
	);
	LUT2 #(
		.INIT('h4)
	) name5039 (
		_w5494_,
		_w5500_,
		_w5501_
	);
	LUT2 #(
		.INIT('h2)
	) name5040 (
		_w1824_,
		_w5501_,
		_w5502_
	);
	LUT2 #(
		.INIT('h4)
	) name5041 (
		_w1824_,
		_w5501_,
		_w5503_
	);
	LUT2 #(
		.INIT('h1)
	) name5042 (
		_w5502_,
		_w5503_,
		_w5504_
	);
	LUT2 #(
		.INIT('h2)
	) name5043 (
		_w3980_,
		_w5504_,
		_w5505_
	);
	LUT2 #(
		.INIT('h1)
	) name5044 (
		_w5480_,
		_w5505_,
		_w5506_
	);
	LUT2 #(
		.INIT('h1)
	) name5045 (
		_w3677_,
		_w5506_,
		_w5507_
	);
	LUT2 #(
		.INIT('h8)
	) name5046 (
		_w4009_,
		_w4011_,
		_w5508_
	);
	LUT2 #(
		.INIT('h4)
	) name5047 (
		_w3988_,
		_w3991_,
		_w5509_
	);
	LUT2 #(
		.INIT('h8)
	) name5048 (
		_w3982_,
		_w3997_,
		_w5510_
	);
	LUT2 #(
		.INIT('h4)
	) name5049 (
		_w5509_,
		_w5510_,
		_w5511_
	);
	LUT2 #(
		.INIT('h4)
	) name5050 (
		_w3994_,
		_w3997_,
		_w5512_
	);
	LUT2 #(
		.INIT('h2)
	) name5051 (
		_w4002_,
		_w5512_,
		_w5513_
	);
	LUT2 #(
		.INIT('h4)
	) name5052 (
		_w5511_,
		_w5513_,
		_w5514_
	);
	LUT2 #(
		.INIT('h8)
	) name5053 (
		_w3998_,
		_w4008_,
		_w5515_
	);
	LUT2 #(
		.INIT('h4)
	) name5054 (
		_w5514_,
		_w5515_,
		_w5516_
	);
	LUT2 #(
		.INIT('h8)
	) name5055 (
		_w5508_,
		_w5516_,
		_w5517_
	);
	LUT2 #(
		.INIT('h8)
	) name5056 (
		_w4005_,
		_w4008_,
		_w5518_
	);
	LUT2 #(
		.INIT('h2)
	) name5057 (
		_w4017_,
		_w5518_,
		_w5519_
	);
	LUT2 #(
		.INIT('h2)
	) name5058 (
		_w5508_,
		_w5519_,
		_w5520_
	);
	LUT2 #(
		.INIT('h2)
	) name5059 (
		_w4011_,
		_w4020_,
		_w5521_
	);
	LUT2 #(
		.INIT('h1)
	) name5060 (
		_w4024_,
		_w5521_,
		_w5522_
	);
	LUT2 #(
		.INIT('h4)
	) name5061 (
		_w5520_,
		_w5522_,
		_w5523_
	);
	LUT2 #(
		.INIT('h4)
	) name5062 (
		_w5517_,
		_w5523_,
		_w5524_
	);
	LUT2 #(
		.INIT('h2)
	) name5063 (
		_w1824_,
		_w5524_,
		_w5525_
	);
	LUT2 #(
		.INIT('h4)
	) name5064 (
		_w1824_,
		_w5524_,
		_w5526_
	);
	LUT2 #(
		.INIT('h1)
	) name5065 (
		_w5525_,
		_w5526_,
		_w5527_
	);
	LUT2 #(
		.INIT('h8)
	) name5066 (
		_w3980_,
		_w5527_,
		_w5528_
	);
	LUT2 #(
		.INIT('h1)
	) name5067 (
		_w5480_,
		_w5528_,
		_w5529_
	);
	LUT2 #(
		.INIT('h1)
	) name5068 (
		_w3563_,
		_w5529_,
		_w5530_
	);
	LUT2 #(
		.INIT('h1)
	) name5069 (
		_w1427_,
		_w5458_,
		_w5531_
	);
	LUT2 #(
		.INIT('h8)
	) name5070 (
		_w1427_,
		_w5458_,
		_w5532_
	);
	LUT2 #(
		.INIT('h1)
	) name5071 (
		_w5531_,
		_w5532_,
		_w5533_
	);
	LUT2 #(
		.INIT('h1)
	) name5072 (
		_w537_,
		_w5533_,
		_w5534_
	);
	LUT2 #(
		.INIT('h2)
	) name5073 (
		_w537_,
		_w1452_,
		_w5535_
	);
	LUT2 #(
		.INIT('h1)
	) name5074 (
		_w5534_,
		_w5535_,
		_w5536_
	);
	LUT2 #(
		.INIT('h2)
	) name5075 (
		_w3980_,
		_w5536_,
		_w5537_
	);
	LUT2 #(
		.INIT('h1)
	) name5076 (
		_w5480_,
		_w5537_,
		_w5538_
	);
	LUT2 #(
		.INIT('h2)
	) name5077 (
		_w1936_,
		_w5538_,
		_w5539_
	);
	LUT2 #(
		.INIT('h2)
	) name5078 (
		_w1394_,
		_w4067_,
		_w5540_
	);
	LUT2 #(
		.INIT('h1)
	) name5079 (
		_w5479_,
		_w5540_,
		_w5541_
	);
	LUT2 #(
		.INIT('h4)
	) name5080 (
		_w5485_,
		_w5541_,
		_w5542_
	);
	LUT2 #(
		.INIT('h1)
	) name5081 (
		_w5507_,
		_w5530_,
		_w5543_
	);
	LUT2 #(
		.INIT('h4)
	) name5082 (
		_w5539_,
		_w5543_,
		_w5544_
	);
	LUT2 #(
		.INIT('h8)
	) name5083 (
		_w5542_,
		_w5544_,
		_w5545_
	);
	LUT2 #(
		.INIT('h2)
	) name5084 (
		_w3450_,
		_w5545_,
		_w5546_
	);
	LUT2 #(
		.INIT('h1)
	) name5085 (
		_w5478_,
		_w5546_,
		_w5547_
	);
	LUT2 #(
		.INIT('h2)
	) name5086 (
		\P1_state_reg[0]/NET0131 ,
		_w5547_,
		_w5548_
	);
	LUT2 #(
		.INIT('h1)
	) name5087 (
		_w5476_,
		_w5477_,
		_w5549_
	);
	LUT2 #(
		.INIT('h4)
	) name5088 (
		_w5548_,
		_w5549_,
		_w5550_
	);
	LUT2 #(
		.INIT('h4)
	) name5089 (
		\P1_state_reg[0]/NET0131 ,
		\P2_reg3_reg[17]/NET0131 ,
		_w5551_
	);
	LUT2 #(
		.INIT('h8)
	) name5090 (
		_w2373_,
		_w3976_,
		_w5552_
	);
	LUT2 #(
		.INIT('h8)
	) name5091 (
		_w2024_,
		_w2373_,
		_w5553_
	);
	LUT2 #(
		.INIT('h2)
	) name5092 (
		_w2399_,
		_w3965_,
		_w5554_
	);
	LUT2 #(
		.INIT('h2)
	) name5093 (
		_w2373_,
		_w3788_,
		_w5555_
	);
	LUT2 #(
		.INIT('h2)
	) name5094 (
		_w4191_,
		_w4587_,
		_w5556_
	);
	LUT2 #(
		.INIT('h4)
	) name5095 (
		_w4191_,
		_w4587_,
		_w5557_
	);
	LUT2 #(
		.INIT('h1)
	) name5096 (
		_w5556_,
		_w5557_,
		_w5558_
	);
	LUT2 #(
		.INIT('h8)
	) name5097 (
		_w3788_,
		_w5558_,
		_w5559_
	);
	LUT2 #(
		.INIT('h1)
	) name5098 (
		_w5555_,
		_w5559_,
		_w5560_
	);
	LUT2 #(
		.INIT('h1)
	) name5099 (
		_w3177_,
		_w5560_,
		_w5561_
	);
	LUT2 #(
		.INIT('h2)
	) name5100 (
		_w2058_,
		_w2804_,
		_w5562_
	);
	LUT2 #(
		.INIT('h8)
	) name5101 (
		_w3387_,
		_w3390_,
		_w5563_
	);
	LUT2 #(
		.INIT('h4)
	) name5102 (
		_w2828_,
		_w3387_,
		_w5564_
	);
	LUT2 #(
		.INIT('h4)
	) name5103 (
		_w2804_,
		_w5564_,
		_w5565_
	);
	LUT2 #(
		.INIT('h4)
	) name5104 (
		_w2379_,
		_w5565_,
		_w5566_
	);
	LUT2 #(
		.INIT('h2)
	) name5105 (
		_w2442_,
		_w5566_,
		_w5567_
	);
	LUT2 #(
		.INIT('h1)
	) name5106 (
		_w2058_,
		_w5563_,
		_w5568_
	);
	LUT2 #(
		.INIT('h4)
	) name5107 (
		_w5567_,
		_w5568_,
		_w5569_
	);
	LUT2 #(
		.INIT('h1)
	) name5108 (
		_w5562_,
		_w5569_,
		_w5570_
	);
	LUT2 #(
		.INIT('h2)
	) name5109 (
		_w3788_,
		_w5570_,
		_w5571_
	);
	LUT2 #(
		.INIT('h1)
	) name5110 (
		_w5555_,
		_w5571_,
		_w5572_
	);
	LUT2 #(
		.INIT('h2)
	) name5111 (
		_w3411_,
		_w5572_,
		_w5573_
	);
	LUT2 #(
		.INIT('h4)
	) name5112 (
		_w2843_,
		_w3339_,
		_w5574_
	);
	LUT2 #(
		.INIT('h4)
	) name5113 (
		_w2818_,
		_w5574_,
		_w5575_
	);
	LUT2 #(
		.INIT('h2)
	) name5114 (
		_w2399_,
		_w5575_,
		_w5576_
	);
	LUT2 #(
		.INIT('h4)
	) name5115 (
		_w2399_,
		_w5575_,
		_w5577_
	);
	LUT2 #(
		.INIT('h1)
	) name5116 (
		_w5576_,
		_w5577_,
		_w5578_
	);
	LUT2 #(
		.INIT('h8)
	) name5117 (
		_w3788_,
		_w5578_,
		_w5579_
	);
	LUT2 #(
		.INIT('h1)
	) name5118 (
		_w5555_,
		_w5579_,
		_w5580_
	);
	LUT2 #(
		.INIT('h2)
	) name5119 (
		_w3355_,
		_w5580_,
		_w5581_
	);
	LUT2 #(
		.INIT('h2)
	) name5120 (
		_w3223_,
		_w3280_,
		_w5582_
	);
	LUT2 #(
		.INIT('h2)
	) name5121 (
		_w3291_,
		_w5582_,
		_w5583_
	);
	LUT2 #(
		.INIT('h8)
	) name5122 (
		_w4191_,
		_w5583_,
		_w5584_
	);
	LUT2 #(
		.INIT('h1)
	) name5123 (
		_w4191_,
		_w5583_,
		_w5585_
	);
	LUT2 #(
		.INIT('h1)
	) name5124 (
		_w5584_,
		_w5585_,
		_w5586_
	);
	LUT2 #(
		.INIT('h8)
	) name5125 (
		_w3788_,
		_w5586_,
		_w5587_
	);
	LUT2 #(
		.INIT('h1)
	) name5126 (
		_w5555_,
		_w5587_,
		_w5588_
	);
	LUT2 #(
		.INIT('h1)
	) name5127 (
		_w3320_,
		_w5588_,
		_w5589_
	);
	LUT2 #(
		.INIT('h2)
	) name5128 (
		_w2373_,
		_w3962_,
		_w5590_
	);
	LUT2 #(
		.INIT('h1)
	) name5129 (
		_w5554_,
		_w5590_,
		_w5591_
	);
	LUT2 #(
		.INIT('h4)
	) name5130 (
		_w5589_,
		_w5591_,
		_w5592_
	);
	LUT2 #(
		.INIT('h4)
	) name5131 (
		_w5561_,
		_w5592_,
		_w5593_
	);
	LUT2 #(
		.INIT('h1)
	) name5132 (
		_w5573_,
		_w5581_,
		_w5594_
	);
	LUT2 #(
		.INIT('h8)
	) name5133 (
		_w5593_,
		_w5594_,
		_w5595_
	);
	LUT2 #(
		.INIT('h2)
	) name5134 (
		_w2026_,
		_w5595_,
		_w5596_
	);
	LUT2 #(
		.INIT('h1)
	) name5135 (
		_w5553_,
		_w5596_,
		_w5597_
	);
	LUT2 #(
		.INIT('h2)
	) name5136 (
		\P1_state_reg[0]/NET0131 ,
		_w5597_,
		_w5598_
	);
	LUT2 #(
		.INIT('h1)
	) name5137 (
		_w5551_,
		_w5552_,
		_w5599_
	);
	LUT2 #(
		.INIT('h4)
	) name5138 (
		_w5598_,
		_w5599_,
		_w5600_
	);
	LUT2 #(
		.INIT('h8)
	) name5139 (
		_w2307_,
		_w3976_,
		_w5601_
	);
	LUT2 #(
		.INIT('h4)
	) name5140 (
		\P1_state_reg[0]/NET0131 ,
		\P2_reg3_reg[19]/NET0131 ,
		_w5602_
	);
	LUT2 #(
		.INIT('h8)
	) name5141 (
		_w2024_,
		_w2307_,
		_w5603_
	);
	LUT2 #(
		.INIT('h2)
	) name5142 (
		_w2307_,
		_w3962_,
		_w5604_
	);
	LUT2 #(
		.INIT('h2)
	) name5143 (
		_w2307_,
		_w3788_,
		_w5605_
	);
	LUT2 #(
		.INIT('h2)
	) name5144 (
		_w4197_,
		_w4814_,
		_w5606_
	);
	LUT2 #(
		.INIT('h4)
	) name5145 (
		_w4197_,
		_w4814_,
		_w5607_
	);
	LUT2 #(
		.INIT('h1)
	) name5146 (
		_w5606_,
		_w5607_,
		_w5608_
	);
	LUT2 #(
		.INIT('h8)
	) name5147 (
		_w3788_,
		_w5608_,
		_w5609_
	);
	LUT2 #(
		.INIT('h1)
	) name5148 (
		_w5605_,
		_w5609_,
		_w5610_
	);
	LUT2 #(
		.INIT('h1)
	) name5149 (
		_w3177_,
		_w5610_,
		_w5611_
	);
	LUT2 #(
		.INIT('h2)
	) name5150 (
		_w4197_,
		_w4850_,
		_w5612_
	);
	LUT2 #(
		.INIT('h4)
	) name5151 (
		_w4197_,
		_w4850_,
		_w5613_
	);
	LUT2 #(
		.INIT('h1)
	) name5152 (
		_w5612_,
		_w5613_,
		_w5614_
	);
	LUT2 #(
		.INIT('h2)
	) name5153 (
		_w3788_,
		_w5614_,
		_w5615_
	);
	LUT2 #(
		.INIT('h1)
	) name5154 (
		_w5605_,
		_w5615_,
		_w5616_
	);
	LUT2 #(
		.INIT('h1)
	) name5155 (
		_w3320_,
		_w5616_,
		_w5617_
	);
	LUT2 #(
		.INIT('h4)
	) name5156 (
		_w2311_,
		_w5563_,
		_w5618_
	);
	LUT2 #(
		.INIT('h2)
	) name5157 (
		_w2368_,
		_w5618_,
		_w5619_
	);
	LUT2 #(
		.INIT('h4)
	) name5158 (
		_w2368_,
		_w5618_,
		_w5620_
	);
	LUT2 #(
		.INIT('h1)
	) name5159 (
		_w5619_,
		_w5620_,
		_w5621_
	);
	LUT2 #(
		.INIT('h1)
	) name5160 (
		_w2058_,
		_w5621_,
		_w5622_
	);
	LUT2 #(
		.INIT('h8)
	) name5161 (
		_w2058_,
		_w2442_,
		_w5623_
	);
	LUT2 #(
		.INIT('h1)
	) name5162 (
		_w5622_,
		_w5623_,
		_w5624_
	);
	LUT2 #(
		.INIT('h8)
	) name5163 (
		_w3788_,
		_w5624_,
		_w5625_
	);
	LUT2 #(
		.INIT('h1)
	) name5164 (
		_w5605_,
		_w5625_,
		_w5626_
	);
	LUT2 #(
		.INIT('h2)
	) name5165 (
		_w3411_,
		_w5626_,
		_w5627_
	);
	LUT2 #(
		.INIT('h2)
	) name5166 (
		_w2299_,
		_w3343_,
		_w5628_
	);
	LUT2 #(
		.INIT('h4)
	) name5167 (
		_w2299_,
		_w3343_,
		_w5629_
	);
	LUT2 #(
		.INIT('h1)
	) name5168 (
		_w5628_,
		_w5629_,
		_w5630_
	);
	LUT2 #(
		.INIT('h8)
	) name5169 (
		_w3788_,
		_w5630_,
		_w5631_
	);
	LUT2 #(
		.INIT('h1)
	) name5170 (
		_w5605_,
		_w5631_,
		_w5632_
	);
	LUT2 #(
		.INIT('h2)
	) name5171 (
		_w3355_,
		_w5632_,
		_w5633_
	);
	LUT2 #(
		.INIT('h2)
	) name5172 (
		_w2299_,
		_w3965_,
		_w5634_
	);
	LUT2 #(
		.INIT('h1)
	) name5173 (
		_w5604_,
		_w5634_,
		_w5635_
	);
	LUT2 #(
		.INIT('h4)
	) name5174 (
		_w5617_,
		_w5635_,
		_w5636_
	);
	LUT2 #(
		.INIT('h4)
	) name5175 (
		_w5633_,
		_w5636_,
		_w5637_
	);
	LUT2 #(
		.INIT('h4)
	) name5176 (
		_w5627_,
		_w5637_,
		_w5638_
	);
	LUT2 #(
		.INIT('h4)
	) name5177 (
		_w5611_,
		_w5638_,
		_w5639_
	);
	LUT2 #(
		.INIT('h2)
	) name5178 (
		_w2026_,
		_w5639_,
		_w5640_
	);
	LUT2 #(
		.INIT('h1)
	) name5179 (
		_w5603_,
		_w5640_,
		_w5641_
	);
	LUT2 #(
		.INIT('h2)
	) name5180 (
		\P1_state_reg[0]/NET0131 ,
		_w5641_,
		_w5642_
	);
	LUT2 #(
		.INIT('h1)
	) name5181 (
		_w5601_,
		_w5602_,
		_w5643_
	);
	LUT2 #(
		.INIT('h4)
	) name5182 (
		_w5642_,
		_w5643_,
		_w5644_
	);
	LUT2 #(
		.INIT('h8)
	) name5183 (
		_w1423_,
		_w3448_,
		_w5645_
	);
	LUT2 #(
		.INIT('h2)
	) name5184 (
		_w1423_,
		_w3980_,
		_w5646_
	);
	LUT2 #(
		.INIT('h2)
	) name5185 (
		_w537_,
		_w1403_,
		_w5647_
	);
	LUT2 #(
		.INIT('h4)
	) name5186 (
		_w1403_,
		_w5195_,
		_w5648_
	);
	LUT2 #(
		.INIT('h8)
	) name5187 (
		_w3587_,
		_w5648_,
		_w5649_
	);
	LUT2 #(
		.INIT('h4)
	) name5188 (
		_w1427_,
		_w5648_,
		_w5650_
	);
	LUT2 #(
		.INIT('h2)
	) name5189 (
		_w1374_,
		_w5650_,
		_w5651_
	);
	LUT2 #(
		.INIT('h1)
	) name5190 (
		_w537_,
		_w5649_,
		_w5652_
	);
	LUT2 #(
		.INIT('h4)
	) name5191 (
		_w5651_,
		_w5652_,
		_w5653_
	);
	LUT2 #(
		.INIT('h1)
	) name5192 (
		_w5647_,
		_w5653_,
		_w5654_
	);
	LUT2 #(
		.INIT('h2)
	) name5193 (
		_w3980_,
		_w5654_,
		_w5655_
	);
	LUT2 #(
		.INIT('h1)
	) name5194 (
		_w5646_,
		_w5655_,
		_w5656_
	);
	LUT2 #(
		.INIT('h2)
	) name5195 (
		_w1936_,
		_w5656_,
		_w5657_
	);
	LUT2 #(
		.INIT('h2)
	) name5196 (
		_w1423_,
		_w4910_,
		_w5658_
	);
	LUT2 #(
		.INIT('h2)
	) name5197 (
		_w1835_,
		_w4458_,
		_w5659_
	);
	LUT2 #(
		.INIT('h4)
	) name5198 (
		_w1835_,
		_w4458_,
		_w5660_
	);
	LUT2 #(
		.INIT('h1)
	) name5199 (
		_w5659_,
		_w5660_,
		_w5661_
	);
	LUT2 #(
		.INIT('h8)
	) name5200 (
		_w3980_,
		_w5661_,
		_w5662_
	);
	LUT2 #(
		.INIT('h1)
	) name5201 (
		_w5646_,
		_w5662_,
		_w5663_
	);
	LUT2 #(
		.INIT('h1)
	) name5202 (
		_w3563_,
		_w5663_,
		_w5664_
	);
	LUT2 #(
		.INIT('h2)
	) name5203 (
		_w1835_,
		_w4415_,
		_w5665_
	);
	LUT2 #(
		.INIT('h4)
	) name5204 (
		_w1835_,
		_w4415_,
		_w5666_
	);
	LUT2 #(
		.INIT('h1)
	) name5205 (
		_w5665_,
		_w5666_,
		_w5667_
	);
	LUT2 #(
		.INIT('h2)
	) name5206 (
		_w3980_,
		_w5667_,
		_w5668_
	);
	LUT2 #(
		.INIT('h1)
	) name5207 (
		_w5646_,
		_w5668_,
		_w5669_
	);
	LUT2 #(
		.INIT('h1)
	) name5208 (
		_w3677_,
		_w5669_,
		_w5670_
	);
	LUT2 #(
		.INIT('h4)
	) name5209 (
		_w1418_,
		_w3696_,
		_w5671_
	);
	LUT2 #(
		.INIT('h2)
	) name5210 (
		_w1418_,
		_w3696_,
		_w5672_
	);
	LUT2 #(
		.INIT('h1)
	) name5211 (
		_w5671_,
		_w5672_,
		_w5673_
	);
	LUT2 #(
		.INIT('h8)
	) name5212 (
		_w3712_,
		_w5673_,
		_w5674_
	);
	LUT2 #(
		.INIT('h8)
	) name5213 (
		_w3980_,
		_w5674_,
		_w5675_
	);
	LUT2 #(
		.INIT('h2)
	) name5214 (
		_w1418_,
		_w4067_,
		_w5676_
	);
	LUT2 #(
		.INIT('h1)
	) name5215 (
		_w5658_,
		_w5676_,
		_w5677_
	);
	LUT2 #(
		.INIT('h4)
	) name5216 (
		_w5675_,
		_w5677_,
		_w5678_
	);
	LUT2 #(
		.INIT('h4)
	) name5217 (
		_w5664_,
		_w5678_,
		_w5679_
	);
	LUT2 #(
		.INIT('h4)
	) name5218 (
		_w5670_,
		_w5679_,
		_w5680_
	);
	LUT2 #(
		.INIT('h4)
	) name5219 (
		_w5657_,
		_w5680_,
		_w5681_
	);
	LUT2 #(
		.INIT('h2)
	) name5220 (
		_w3450_,
		_w5681_,
		_w5682_
	);
	LUT2 #(
		.INIT('h1)
	) name5221 (
		_w5645_,
		_w5682_,
		_w5683_
	);
	LUT2 #(
		.INIT('h2)
	) name5222 (
		\P1_state_reg[0]/NET0131 ,
		_w5683_,
		_w5684_
	);
	LUT2 #(
		.INIT('h2)
	) name5223 (
		\P1_reg3_reg[19]/NET0131 ,
		\P1_state_reg[0]/NET0131 ,
		_w5685_
	);
	LUT2 #(
		.INIT('h8)
	) name5224 (
		_w1423_,
		_w1953_,
		_w5686_
	);
	LUT2 #(
		.INIT('h1)
	) name5225 (
		_w5685_,
		_w5686_,
		_w5687_
	);
	LUT2 #(
		.INIT('h4)
	) name5226 (
		_w5684_,
		_w5687_,
		_w5688_
	);
	LUT2 #(
		.INIT('h8)
	) name5227 (
		_w2024_,
		_w3058_,
		_w5689_
	);
	LUT2 #(
		.INIT('h2)
	) name5228 (
		_w3058_,
		_w3788_,
		_w5690_
	);
	LUT2 #(
		.INIT('h2)
	) name5229 (
		_w3788_,
		_w4983_,
		_w5691_
	);
	LUT2 #(
		.INIT('h1)
	) name5230 (
		_w5690_,
		_w5691_,
		_w5692_
	);
	LUT2 #(
		.INIT('h1)
	) name5231 (
		_w3320_,
		_w5692_,
		_w5693_
	);
	LUT2 #(
		.INIT('h2)
	) name5232 (
		_w3788_,
		_w4997_,
		_w5694_
	);
	LUT2 #(
		.INIT('h1)
	) name5233 (
		_w5690_,
		_w5694_,
		_w5695_
	);
	LUT2 #(
		.INIT('h1)
	) name5234 (
		_w3177_,
		_w5695_,
		_w5696_
	);
	LUT2 #(
		.INIT('h2)
	) name5235 (
		_w3355_,
		_w3788_,
		_w5697_
	);
	LUT2 #(
		.INIT('h2)
	) name5236 (
		_w3962_,
		_w5697_,
		_w5698_
	);
	LUT2 #(
		.INIT('h2)
	) name5237 (
		_w3058_,
		_w5698_,
		_w5699_
	);
	LUT2 #(
		.INIT('h8)
	) name5238 (
		_w3788_,
		_w5008_,
		_w5700_
	);
	LUT2 #(
		.INIT('h1)
	) name5239 (
		_w5690_,
		_w5700_,
		_w5701_
	);
	LUT2 #(
		.INIT('h2)
	) name5240 (
		_w3411_,
		_w5701_,
		_w5702_
	);
	LUT2 #(
		.INIT('h8)
	) name5241 (
		_w3788_,
		_w5003_,
		_w5703_
	);
	LUT2 #(
		.INIT('h2)
	) name5242 (
		_w3054_,
		_w3965_,
		_w5704_
	);
	LUT2 #(
		.INIT('h1)
	) name5243 (
		_w5699_,
		_w5704_,
		_w5705_
	);
	LUT2 #(
		.INIT('h4)
	) name5244 (
		_w5703_,
		_w5705_,
		_w5706_
	);
	LUT2 #(
		.INIT('h4)
	) name5245 (
		_w5702_,
		_w5706_,
		_w5707_
	);
	LUT2 #(
		.INIT('h4)
	) name5246 (
		_w5696_,
		_w5707_,
		_w5708_
	);
	LUT2 #(
		.INIT('h4)
	) name5247 (
		_w5693_,
		_w5708_,
		_w5709_
	);
	LUT2 #(
		.INIT('h2)
	) name5248 (
		_w2026_,
		_w5709_,
		_w5710_
	);
	LUT2 #(
		.INIT('h1)
	) name5249 (
		_w5689_,
		_w5710_,
		_w5711_
	);
	LUT2 #(
		.INIT('h2)
	) name5250 (
		\P1_state_reg[0]/NET0131 ,
		_w5711_,
		_w5712_
	);
	LUT2 #(
		.INIT('h4)
	) name5251 (
		\P1_state_reg[0]/NET0131 ,
		\P2_reg3_reg[24]/NET0131 ,
		_w5713_
	);
	LUT2 #(
		.INIT('h8)
	) name5252 (
		_w3058_,
		_w3976_,
		_w5714_
	);
	LUT2 #(
		.INIT('h1)
	) name5253 (
		_w5713_,
		_w5714_,
		_w5715_
	);
	LUT2 #(
		.INIT('h4)
	) name5254 (
		_w5712_,
		_w5715_,
		_w5716_
	);
	LUT2 #(
		.INIT('h2)
	) name5255 (
		\P1_reg3_reg[24]/NET0131 ,
		\P1_state_reg[0]/NET0131 ,
		_w5717_
	);
	LUT2 #(
		.INIT('h8)
	) name5256 (
		_w1058_,
		_w1953_,
		_w5718_
	);
	LUT2 #(
		.INIT('h8)
	) name5257 (
		_w1058_,
		_w3448_,
		_w5719_
	);
	LUT2 #(
		.INIT('h2)
	) name5258 (
		_w1058_,
		_w3980_,
		_w5720_
	);
	LUT2 #(
		.INIT('h2)
	) name5259 (
		_w3980_,
		_w5172_,
		_w5721_
	);
	LUT2 #(
		.INIT('h1)
	) name5260 (
		_w5720_,
		_w5721_,
		_w5722_
	);
	LUT2 #(
		.INIT('h1)
	) name5261 (
		_w3563_,
		_w5722_,
		_w5723_
	);
	LUT2 #(
		.INIT('h2)
	) name5262 (
		_w3980_,
		_w5184_,
		_w5724_
	);
	LUT2 #(
		.INIT('h1)
	) name5263 (
		_w5720_,
		_w5724_,
		_w5725_
	);
	LUT2 #(
		.INIT('h1)
	) name5264 (
		_w3677_,
		_w5725_,
		_w5726_
	);
	LUT2 #(
		.INIT('h2)
	) name5265 (
		_w1058_,
		_w4064_,
		_w5727_
	);
	LUT2 #(
		.INIT('h2)
	) name5266 (
		_w1047_,
		_w4067_,
		_w5728_
	);
	LUT2 #(
		.INIT('h8)
	) name5267 (
		_w3980_,
		_w5190_,
		_w5729_
	);
	LUT2 #(
		.INIT('h1)
	) name5268 (
		_w5720_,
		_w5729_,
		_w5730_
	);
	LUT2 #(
		.INIT('h2)
	) name5269 (
		_w3712_,
		_w5730_,
		_w5731_
	);
	LUT2 #(
		.INIT('h8)
	) name5270 (
		_w3980_,
		_w5200_,
		_w5732_
	);
	LUT2 #(
		.INIT('h1)
	) name5271 (
		_w5720_,
		_w5732_,
		_w5733_
	);
	LUT2 #(
		.INIT('h2)
	) name5272 (
		_w1936_,
		_w5733_,
		_w5734_
	);
	LUT2 #(
		.INIT('h1)
	) name5273 (
		_w5727_,
		_w5728_,
		_w5735_
	);
	LUT2 #(
		.INIT('h4)
	) name5274 (
		_w5731_,
		_w5735_,
		_w5736_
	);
	LUT2 #(
		.INIT('h4)
	) name5275 (
		_w5723_,
		_w5736_,
		_w5737_
	);
	LUT2 #(
		.INIT('h1)
	) name5276 (
		_w5726_,
		_w5734_,
		_w5738_
	);
	LUT2 #(
		.INIT('h8)
	) name5277 (
		_w5737_,
		_w5738_,
		_w5739_
	);
	LUT2 #(
		.INIT('h2)
	) name5278 (
		_w3450_,
		_w5739_,
		_w5740_
	);
	LUT2 #(
		.INIT('h1)
	) name5279 (
		_w5719_,
		_w5740_,
		_w5741_
	);
	LUT2 #(
		.INIT('h2)
	) name5280 (
		\P1_state_reg[0]/NET0131 ,
		_w5741_,
		_w5742_
	);
	LUT2 #(
		.INIT('h1)
	) name5281 (
		_w5717_,
		_w5718_,
		_w5743_
	);
	LUT2 #(
		.INIT('h4)
	) name5282 (
		_w5742_,
		_w5743_,
		_w5744_
	);
	LUT2 #(
		.INIT('h4)
	) name5283 (
		\P1_state_reg[0]/NET0131 ,
		\P2_reg3_reg[22]/NET0131 ,
		_w5745_
	);
	LUT2 #(
		.INIT('h8)
	) name5284 (
		_w3108_,
		_w3976_,
		_w5746_
	);
	LUT2 #(
		.INIT('h8)
	) name5285 (
		_w2024_,
		_w3108_,
		_w5747_
	);
	LUT2 #(
		.INIT('h2)
	) name5286 (
		_w3108_,
		_w3788_,
		_w5748_
	);
	LUT2 #(
		.INIT('h4)
	) name5287 (
		_w4750_,
		_w4752_,
		_w5749_
	);
	LUT2 #(
		.INIT('h2)
	) name5288 (
		_w4757_,
		_w5749_,
		_w5750_
	);
	LUT2 #(
		.INIT('h8)
	) name5289 (
		_w4209_,
		_w5750_,
		_w5751_
	);
	LUT2 #(
		.INIT('h1)
	) name5290 (
		_w4209_,
		_w5750_,
		_w5752_
	);
	LUT2 #(
		.INIT('h1)
	) name5291 (
		_w5751_,
		_w5752_,
		_w5753_
	);
	LUT2 #(
		.INIT('h2)
	) name5292 (
		_w3788_,
		_w5753_,
		_w5754_
	);
	LUT2 #(
		.INIT('h1)
	) name5293 (
		_w5748_,
		_w5754_,
		_w5755_
	);
	LUT2 #(
		.INIT('h1)
	) name5294 (
		_w3177_,
		_w5755_,
		_w5756_
	);
	LUT2 #(
		.INIT('h4)
	) name5295 (
		_w4721_,
		_w4725_,
		_w5757_
	);
	LUT2 #(
		.INIT('h8)
	) name5296 (
		_w4209_,
		_w5757_,
		_w5758_
	);
	LUT2 #(
		.INIT('h1)
	) name5297 (
		_w4209_,
		_w5757_,
		_w5759_
	);
	LUT2 #(
		.INIT('h1)
	) name5298 (
		_w5758_,
		_w5759_,
		_w5760_
	);
	LUT2 #(
		.INIT('h8)
	) name5299 (
		_w3788_,
		_w5760_,
		_w5761_
	);
	LUT2 #(
		.INIT('h1)
	) name5300 (
		_w5748_,
		_w5761_,
		_w5762_
	);
	LUT2 #(
		.INIT('h1)
	) name5301 (
		_w3320_,
		_w5762_,
		_w5763_
	);
	LUT2 #(
		.INIT('h2)
	) name5302 (
		_w3108_,
		_w3962_,
		_w5764_
	);
	LUT2 #(
		.INIT('h8)
	) name5303 (
		_w3322_,
		_w3343_,
		_w5765_
	);
	LUT2 #(
		.INIT('h4)
	) name5304 (
		_w3121_,
		_w5765_,
		_w5766_
	);
	LUT2 #(
		.INIT('h2)
	) name5305 (
		_w3102_,
		_w5766_,
		_w5767_
	);
	LUT2 #(
		.INIT('h4)
	) name5306 (
		_w3102_,
		_w5766_,
		_w5768_
	);
	LUT2 #(
		.INIT('h1)
	) name5307 (
		_w5767_,
		_w5768_,
		_w5769_
	);
	LUT2 #(
		.INIT('h8)
	) name5308 (
		_w3788_,
		_w5769_,
		_w5770_
	);
	LUT2 #(
		.INIT('h1)
	) name5309 (
		_w5748_,
		_w5770_,
		_w5771_
	);
	LUT2 #(
		.INIT('h2)
	) name5310 (
		_w3355_,
		_w5771_,
		_w5772_
	);
	LUT2 #(
		.INIT('h4)
	) name5311 (
		_w3112_,
		_w3394_,
		_w5773_
	);
	LUT2 #(
		.INIT('h2)
	) name5312 (
		_w3088_,
		_w5773_,
		_w5774_
	);
	LUT2 #(
		.INIT('h4)
	) name5313 (
		_w3088_,
		_w5773_,
		_w5775_
	);
	LUT2 #(
		.INIT('h1)
	) name5314 (
		_w5774_,
		_w5775_,
		_w5776_
	);
	LUT2 #(
		.INIT('h1)
	) name5315 (
		_w2058_,
		_w5776_,
		_w5777_
	);
	LUT2 #(
		.INIT('h8)
	) name5316 (
		_w2058_,
		_w3130_,
		_w5778_
	);
	LUT2 #(
		.INIT('h1)
	) name5317 (
		_w5777_,
		_w5778_,
		_w5779_
	);
	LUT2 #(
		.INIT('h8)
	) name5318 (
		_w3788_,
		_w5779_,
		_w5780_
	);
	LUT2 #(
		.INIT('h1)
	) name5319 (
		_w5748_,
		_w5780_,
		_w5781_
	);
	LUT2 #(
		.INIT('h2)
	) name5320 (
		_w3411_,
		_w5781_,
		_w5782_
	);
	LUT2 #(
		.INIT('h2)
	) name5321 (
		_w3102_,
		_w3965_,
		_w5783_
	);
	LUT2 #(
		.INIT('h1)
	) name5322 (
		_w5764_,
		_w5783_,
		_w5784_
	);
	LUT2 #(
		.INIT('h4)
	) name5323 (
		_w5782_,
		_w5784_,
		_w5785_
	);
	LUT2 #(
		.INIT('h4)
	) name5324 (
		_w5772_,
		_w5785_,
		_w5786_
	);
	LUT2 #(
		.INIT('h4)
	) name5325 (
		_w5756_,
		_w5786_,
		_w5787_
	);
	LUT2 #(
		.INIT('h4)
	) name5326 (
		_w5763_,
		_w5787_,
		_w5788_
	);
	LUT2 #(
		.INIT('h2)
	) name5327 (
		_w2026_,
		_w5788_,
		_w5789_
	);
	LUT2 #(
		.INIT('h1)
	) name5328 (
		_w5747_,
		_w5789_,
		_w5790_
	);
	LUT2 #(
		.INIT('h2)
	) name5329 (
		\P1_state_reg[0]/NET0131 ,
		_w5790_,
		_w5791_
	);
	LUT2 #(
		.INIT('h1)
	) name5330 (
		_w5745_,
		_w5746_,
		_w5792_
	);
	LUT2 #(
		.INIT('h4)
	) name5331 (
		_w5791_,
		_w5792_,
		_w5793_
	);
	LUT2 #(
		.INIT('h8)
	) name5332 (
		_w692_,
		_w1880_,
		_w5794_
	);
	LUT2 #(
		.INIT('h8)
	) name5333 (
		_w3585_,
		_w3589_,
		_w5795_
	);
	LUT2 #(
		.INIT('h8)
	) name5334 (
		_w3586_,
		_w5795_,
		_w5796_
	);
	LUT2 #(
		.INIT('h8)
	) name5335 (
		_w4473_,
		_w5796_,
		_w5797_
	);
	LUT2 #(
		.INIT('h4)
	) name5336 (
		_w831_,
		_w3596_,
		_w5798_
	);
	LUT2 #(
		.INIT('h8)
	) name5337 (
		_w5797_,
		_w5798_,
		_w5799_
	);
	LUT2 #(
		.INIT('h2)
	) name5338 (
		_w1936_,
		_w3567_,
		_w5800_
	);
	LUT2 #(
		.INIT('h4)
	) name5339 (
		_w750_,
		_w5800_,
		_w5801_
	);
	LUT2 #(
		.INIT('h4)
	) name5340 (
		_w5799_,
		_w5801_,
		_w5802_
	);
	LUT2 #(
		.INIT('h4)
	) name5341 (
		_w825_,
		_w3708_,
		_w5803_
	);
	LUT2 #(
		.INIT('h2)
	) name5342 (
		_w692_,
		_w5803_,
		_w5804_
	);
	LUT2 #(
		.INIT('h4)
	) name5343 (
		_w692_,
		_w5803_,
		_w5805_
	);
	LUT2 #(
		.INIT('h2)
	) name5344 (
		_w3712_,
		_w5804_,
		_w5806_
	);
	LUT2 #(
		.INIT('h4)
	) name5345 (
		_w5805_,
		_w5806_,
		_w5807_
	);
	LUT2 #(
		.INIT('h1)
	) name5346 (
		_w5794_,
		_w5802_,
		_w5808_
	);
	LUT2 #(
		.INIT('h4)
	) name5347 (
		_w5807_,
		_w5808_,
		_w5809_
	);
	LUT2 #(
		.INIT('h2)
	) name5348 (
		_w3466_,
		_w5809_,
		_w5810_
	);
	LUT2 #(
		.INIT('h1)
	) name5349 (
		_w3720_,
		_w5810_,
		_w5811_
	);
	LUT2 #(
		.INIT('h2)
	) name5350 (
		_w3435_,
		_w3447_,
		_w5812_
	);
	LUT2 #(
		.INIT('h4)
	) name5351 (
		_w5811_,
		_w5812_,
		_w5813_
	);
	LUT2 #(
		.INIT('h1)
	) name5352 (
		_w1763_,
		_w3466_,
		_w5814_
	);
	LUT2 #(
		.INIT('h4)
	) name5353 (
		_w3716_,
		_w5812_,
		_w5815_
	);
	LUT2 #(
		.INIT('h4)
	) name5354 (
		_w5814_,
		_w5815_,
		_w5816_
	);
	LUT2 #(
		.INIT('h2)
	) name5355 (
		\P1_reg2_reg[31]/NET0131 ,
		_w5816_,
		_w5817_
	);
	LUT2 #(
		.INIT('h1)
	) name5356 (
		_w5813_,
		_w5817_,
		_w5818_
	);
	LUT2 #(
		.INIT('h2)
	) name5357 (
		\P2_reg0_reg[25]/NET0131 ,
		_w1983_,
		_w5819_
	);
	LUT2 #(
		.INIT('h8)
	) name5358 (
		\P2_reg0_reg[25]/NET0131 ,
		_w2024_,
		_w5820_
	);
	LUT2 #(
		.INIT('h2)
	) name5359 (
		\P2_reg0_reg[25]/NET0131 ,
		_w2040_,
		_w5821_
	);
	LUT2 #(
		.INIT('h2)
	) name5360 (
		_w2040_,
		_w4595_,
		_w5822_
	);
	LUT2 #(
		.INIT('h1)
	) name5361 (
		_w5821_,
		_w5822_,
		_w5823_
	);
	LUT2 #(
		.INIT('h1)
	) name5362 (
		_w3177_,
		_w5823_,
		_w5824_
	);
	LUT2 #(
		.INIT('h2)
	) name5363 (
		_w2040_,
		_w4609_,
		_w5825_
	);
	LUT2 #(
		.INIT('h1)
	) name5364 (
		_w5821_,
		_w5825_,
		_w5826_
	);
	LUT2 #(
		.INIT('h1)
	) name5365 (
		_w3320_,
		_w5826_,
		_w5827_
	);
	LUT2 #(
		.INIT('h2)
	) name5366 (
		_w2040_,
		_w4928_,
		_w5828_
	);
	LUT2 #(
		.INIT('h8)
	) name5367 (
		_w2040_,
		_w4617_,
		_w5829_
	);
	LUT2 #(
		.INIT('h1)
	) name5368 (
		_w5821_,
		_w5829_,
		_w5830_
	);
	LUT2 #(
		.INIT('h2)
	) name5369 (
		_w3355_,
		_w5830_,
		_w5831_
	);
	LUT2 #(
		.INIT('h4)
	) name5370 (
		_w3416_,
		_w3423_,
		_w5832_
	);
	LUT2 #(
		.INIT('h2)
	) name5371 (
		\P2_reg0_reg[25]/NET0131 ,
		_w5832_,
		_w5833_
	);
	LUT2 #(
		.INIT('h1)
	) name5372 (
		_w5828_,
		_w5833_,
		_w5834_
	);
	LUT2 #(
		.INIT('h4)
	) name5373 (
		_w5831_,
		_w5834_,
		_w5835_
	);
	LUT2 #(
		.INIT('h4)
	) name5374 (
		_w5824_,
		_w5835_,
		_w5836_
	);
	LUT2 #(
		.INIT('h4)
	) name5375 (
		_w5827_,
		_w5836_,
		_w5837_
	);
	LUT2 #(
		.INIT('h2)
	) name5376 (
		_w2026_,
		_w5837_,
		_w5838_
	);
	LUT2 #(
		.INIT('h1)
	) name5377 (
		_w5820_,
		_w5838_,
		_w5839_
	);
	LUT2 #(
		.INIT('h2)
	) name5378 (
		\P1_state_reg[0]/NET0131 ,
		_w5839_,
		_w5840_
	);
	LUT2 #(
		.INIT('h1)
	) name5379 (
		_w5819_,
		_w5840_,
		_w5841_
	);
	LUT2 #(
		.INIT('h2)
	) name5380 (
		\P2_reg0_reg[26]/NET0131 ,
		_w1983_,
		_w5842_
	);
	LUT2 #(
		.INIT('h2)
	) name5381 (
		\P2_reg0_reg[26]/NET0131 ,
		_w2040_,
		_w5843_
	);
	LUT2 #(
		.INIT('h2)
	) name5382 (
		_w2040_,
		_w4732_,
		_w5844_
	);
	LUT2 #(
		.INIT('h1)
	) name5383 (
		_w5843_,
		_w5844_,
		_w5845_
	);
	LUT2 #(
		.INIT('h1)
	) name5384 (
		_w3320_,
		_w5845_,
		_w5846_
	);
	LUT2 #(
		.INIT('h2)
	) name5385 (
		_w2040_,
		_w4764_,
		_w5847_
	);
	LUT2 #(
		.INIT('h1)
	) name5386 (
		_w5843_,
		_w5847_,
		_w5848_
	);
	LUT2 #(
		.INIT('h1)
	) name5387 (
		_w3177_,
		_w5848_,
		_w5849_
	);
	LUT2 #(
		.INIT('h2)
	) name5388 (
		_w2040_,
		_w4962_,
		_w5850_
	);
	LUT2 #(
		.INIT('h2)
	) name5389 (
		\P2_reg0_reg[26]/NET0131 ,
		_w3426_,
		_w5851_
	);
	LUT2 #(
		.INIT('h1)
	) name5390 (
		_w5850_,
		_w5851_,
		_w5852_
	);
	LUT2 #(
		.INIT('h4)
	) name5391 (
		_w5849_,
		_w5852_,
		_w5853_
	);
	LUT2 #(
		.INIT('h4)
	) name5392 (
		_w5846_,
		_w5853_,
		_w5854_
	);
	LUT2 #(
		.INIT('h2)
	) name5393 (
		_w2026_,
		_w5854_,
		_w5855_
	);
	LUT2 #(
		.INIT('h8)
	) name5394 (
		\P2_reg0_reg[26]/NET0131 ,
		_w2024_,
		_w5856_
	);
	LUT2 #(
		.INIT('h1)
	) name5395 (
		_w5855_,
		_w5856_,
		_w5857_
	);
	LUT2 #(
		.INIT('h2)
	) name5396 (
		\P1_state_reg[0]/NET0131 ,
		_w5857_,
		_w5858_
	);
	LUT2 #(
		.INIT('h1)
	) name5397 (
		_w5842_,
		_w5858_,
		_w5859_
	);
	LUT2 #(
		.INIT('h8)
	) name5398 (
		_w2040_,
		_w5287_,
		_w5860_
	);
	LUT2 #(
		.INIT('h8)
	) name5399 (
		_w3421_,
		_w5860_,
		_w5861_
	);
	LUT2 #(
		.INIT('h2)
	) name5400 (
		\P2_reg0_reg[31]/NET0131 ,
		_w5861_,
		_w5862_
	);
	LUT2 #(
		.INIT('h8)
	) name5401 (
		_w3355_,
		_w5282_,
		_w5863_
	);
	LUT2 #(
		.INIT('h2)
	) name5402 (
		_w5278_,
		_w5863_,
		_w5864_
	);
	LUT2 #(
		.INIT('h2)
	) name5403 (
		_w5860_,
		_w5864_,
		_w5865_
	);
	LUT2 #(
		.INIT('h1)
	) name5404 (
		_w5862_,
		_w5865_,
		_w5866_
	);
	LUT2 #(
		.INIT('h2)
	) name5405 (
		\P1_reg2_reg[25]/NET0131 ,
		_w3435_,
		_w5867_
	);
	LUT2 #(
		.INIT('h8)
	) name5406 (
		\P1_reg2_reg[25]/NET0131 ,
		_w3448_,
		_w5868_
	);
	LUT2 #(
		.INIT('h2)
	) name5407 (
		\P1_reg2_reg[25]/NET0131 ,
		_w3466_,
		_w5869_
	);
	LUT2 #(
		.INIT('h2)
	) name5408 (
		_w3466_,
		_w4658_,
		_w5870_
	);
	LUT2 #(
		.INIT('h1)
	) name5409 (
		_w5869_,
		_w5870_,
		_w5871_
	);
	LUT2 #(
		.INIT('h1)
	) name5410 (
		_w3677_,
		_w5871_,
		_w5872_
	);
	LUT2 #(
		.INIT('h2)
	) name5411 (
		_w3466_,
		_w4672_,
		_w5873_
	);
	LUT2 #(
		.INIT('h1)
	) name5412 (
		_w5869_,
		_w5873_,
		_w5874_
	);
	LUT2 #(
		.INIT('h1)
	) name5413 (
		_w3563_,
		_w5874_,
		_w5875_
	);
	LUT2 #(
		.INIT('h8)
	) name5414 (
		_w3466_,
		_w5304_,
		_w5876_
	);
	LUT2 #(
		.INIT('h8)
	) name5415 (
		_w3466_,
		_w4682_,
		_w5877_
	);
	LUT2 #(
		.INIT('h1)
	) name5416 (
		_w5869_,
		_w5877_,
		_w5878_
	);
	LUT2 #(
		.INIT('h2)
	) name5417 (
		_w1936_,
		_w5878_,
		_w5879_
	);
	LUT2 #(
		.INIT('h8)
	) name5418 (
		_w3466_,
		_w4689_,
		_w5880_
	);
	LUT2 #(
		.INIT('h1)
	) name5419 (
		_w5869_,
		_w5880_,
		_w5881_
	);
	LUT2 #(
		.INIT('h2)
	) name5420 (
		_w3712_,
		_w5881_,
		_w5882_
	);
	LUT2 #(
		.INIT('h8)
	) name5421 (
		_w1034_,
		_w1763_,
		_w5883_
	);
	LUT2 #(
		.INIT('h2)
	) name5422 (
		\P1_reg2_reg[25]/NET0131 ,
		_w3718_,
		_w5884_
	);
	LUT2 #(
		.INIT('h1)
	) name5423 (
		_w5876_,
		_w5883_,
		_w5885_
	);
	LUT2 #(
		.INIT('h4)
	) name5424 (
		_w5884_,
		_w5885_,
		_w5886_
	);
	LUT2 #(
		.INIT('h4)
	) name5425 (
		_w5879_,
		_w5886_,
		_w5887_
	);
	LUT2 #(
		.INIT('h4)
	) name5426 (
		_w5882_,
		_w5887_,
		_w5888_
	);
	LUT2 #(
		.INIT('h1)
	) name5427 (
		_w5872_,
		_w5875_,
		_w5889_
	);
	LUT2 #(
		.INIT('h8)
	) name5428 (
		_w5888_,
		_w5889_,
		_w5890_
	);
	LUT2 #(
		.INIT('h2)
	) name5429 (
		_w3450_,
		_w5890_,
		_w5891_
	);
	LUT2 #(
		.INIT('h1)
	) name5430 (
		_w5868_,
		_w5891_,
		_w5892_
	);
	LUT2 #(
		.INIT('h2)
	) name5431 (
		\P1_state_reg[0]/NET0131 ,
		_w5892_,
		_w5893_
	);
	LUT2 #(
		.INIT('h1)
	) name5432 (
		_w5867_,
		_w5893_,
		_w5894_
	);
	LUT2 #(
		.INIT('h2)
	) name5433 (
		\P1_reg2_reg[26]/NET0131 ,
		_w3435_,
		_w5895_
	);
	LUT2 #(
		.INIT('h8)
	) name5434 (
		\P1_reg2_reg[26]/NET0131 ,
		_w3448_,
		_w5896_
	);
	LUT2 #(
		.INIT('h2)
	) name5435 (
		\P1_reg2_reg[26]/NET0131 ,
		_w3466_,
		_w5897_
	);
	LUT2 #(
		.INIT('h1)
	) name5436 (
		_w978_,
		_w5797_,
		_w5898_
	);
	LUT2 #(
		.INIT('h8)
	) name5437 (
		_w978_,
		_w5797_,
		_w5899_
	);
	LUT2 #(
		.INIT('h1)
	) name5438 (
		_w5898_,
		_w5899_,
		_w5900_
	);
	LUT2 #(
		.INIT('h1)
	) name5439 (
		_w537_,
		_w5900_,
		_w5901_
	);
	LUT2 #(
		.INIT('h2)
	) name5440 (
		_w537_,
		_w1038_,
		_w5902_
	);
	LUT2 #(
		.INIT('h1)
	) name5441 (
		_w5901_,
		_w5902_,
		_w5903_
	);
	LUT2 #(
		.INIT('h2)
	) name5442 (
		_w3466_,
		_w5903_,
		_w5904_
	);
	LUT2 #(
		.INIT('h1)
	) name5443 (
		_w5897_,
		_w5904_,
		_w5905_
	);
	LUT2 #(
		.INIT('h2)
	) name5444 (
		_w1936_,
		_w5905_,
		_w5906_
	);
	LUT2 #(
		.INIT('h2)
	) name5445 (
		_w997_,
		_w4688_,
		_w5907_
	);
	LUT2 #(
		.INIT('h1)
	) name5446 (
		_w3704_,
		_w5907_,
		_w5908_
	);
	LUT2 #(
		.INIT('h8)
	) name5447 (
		_w3712_,
		_w5908_,
		_w5909_
	);
	LUT2 #(
		.INIT('h8)
	) name5448 (
		_w997_,
		_w1880_,
		_w5910_
	);
	LUT2 #(
		.INIT('h1)
	) name5449 (
		_w5909_,
		_w5910_,
		_w5911_
	);
	LUT2 #(
		.INIT('h2)
	) name5450 (
		_w3466_,
		_w5911_,
		_w5912_
	);
	LUT2 #(
		.INIT('h4)
	) name5451 (
		_w3466_,
		_w3712_,
		_w5913_
	);
	LUT2 #(
		.INIT('h2)
	) name5452 (
		_w3718_,
		_w5913_,
		_w5914_
	);
	LUT2 #(
		.INIT('h2)
	) name5453 (
		\P1_reg2_reg[26]/NET0131 ,
		_w5914_,
		_w5915_
	);
	LUT2 #(
		.INIT('h8)
	) name5454 (
		_w1002_,
		_w1763_,
		_w5916_
	);
	LUT2 #(
		.INIT('h8)
	) name5455 (
		_w1300_,
		_w1338_,
		_w5917_
	);
	LUT2 #(
		.INIT('h8)
	) name5456 (
		_w1376_,
		_w1429_,
		_w5918_
	);
	LUT2 #(
		.INIT('h8)
	) name5457 (
		_w5917_,
		_w5918_,
		_w5919_
	);
	LUT2 #(
		.INIT('h4)
	) name5458 (
		_w5501_,
		_w5919_,
		_w5920_
	);
	LUT2 #(
		.INIT('h8)
	) name5459 (
		_w1300_,
		_w1709_,
		_w5921_
	);
	LUT2 #(
		.INIT('h8)
	) name5460 (
		_w1376_,
		_w1719_,
		_w5922_
	);
	LUT2 #(
		.INIT('h1)
	) name5461 (
		_w1706_,
		_w5922_,
		_w5923_
	);
	LUT2 #(
		.INIT('h2)
	) name5462 (
		_w5917_,
		_w5923_,
		_w5924_
	);
	LUT2 #(
		.INIT('h1)
	) name5463 (
		_w1066_,
		_w5921_,
		_w5925_
	);
	LUT2 #(
		.INIT('h4)
	) name5464 (
		_w5924_,
		_w5925_,
		_w5926_
	);
	LUT2 #(
		.INIT('h4)
	) name5465 (
		_w5920_,
		_w5926_,
		_w5927_
	);
	LUT2 #(
		.INIT('h2)
	) name5466 (
		_w1809_,
		_w5927_,
		_w5928_
	);
	LUT2 #(
		.INIT('h4)
	) name5467 (
		_w1809_,
		_w5927_,
		_w5929_
	);
	LUT2 #(
		.INIT('h1)
	) name5468 (
		_w5928_,
		_w5929_,
		_w5930_
	);
	LUT2 #(
		.INIT('h2)
	) name5469 (
		_w3466_,
		_w5930_,
		_w5931_
	);
	LUT2 #(
		.INIT('h1)
	) name5470 (
		_w5897_,
		_w5931_,
		_w5932_
	);
	LUT2 #(
		.INIT('h1)
	) name5471 (
		_w3677_,
		_w5932_,
		_w5933_
	);
	LUT2 #(
		.INIT('h8)
	) name5472 (
		_w4012_,
		_w4032_,
		_w5934_
	);
	LUT2 #(
		.INIT('h4)
	) name5473 (
		_w1836_,
		_w4433_,
		_w5935_
	);
	LUT2 #(
		.INIT('h8)
	) name5474 (
		_w5934_,
		_w5935_,
		_w5936_
	);
	LUT2 #(
		.INIT('h4)
	) name5475 (
		_w5524_,
		_w5936_,
		_w5937_
	);
	LUT2 #(
		.INIT('h8)
	) name5476 (
		_w4027_,
		_w4032_,
		_w5938_
	);
	LUT2 #(
		.INIT('h2)
	) name5477 (
		_w4039_,
		_w5938_,
		_w5939_
	);
	LUT2 #(
		.INIT('h2)
	) name5478 (
		_w5935_,
		_w5939_,
		_w5940_
	);
	LUT2 #(
		.INIT('h1)
	) name5479 (
		_w1816_,
		_w4042_,
		_w5941_
	);
	LUT2 #(
		.INIT('h2)
	) name5480 (
		_w4045_,
		_w5941_,
		_w5942_
	);
	LUT2 #(
		.INIT('h1)
	) name5481 (
		_w1810_,
		_w5942_,
		_w5943_
	);
	LUT2 #(
		.INIT('h1)
	) name5482 (
		_w5940_,
		_w5943_,
		_w5944_
	);
	LUT2 #(
		.INIT('h4)
	) name5483 (
		_w5937_,
		_w5944_,
		_w5945_
	);
	LUT2 #(
		.INIT('h8)
	) name5484 (
		_w1809_,
		_w5945_,
		_w5946_
	);
	LUT2 #(
		.INIT('h1)
	) name5485 (
		_w1809_,
		_w5945_,
		_w5947_
	);
	LUT2 #(
		.INIT('h1)
	) name5486 (
		_w5946_,
		_w5947_,
		_w5948_
	);
	LUT2 #(
		.INIT('h2)
	) name5487 (
		_w3466_,
		_w5948_,
		_w5949_
	);
	LUT2 #(
		.INIT('h1)
	) name5488 (
		_w5897_,
		_w5949_,
		_w5950_
	);
	LUT2 #(
		.INIT('h1)
	) name5489 (
		_w3563_,
		_w5950_,
		_w5951_
	);
	LUT2 #(
		.INIT('h1)
	) name5490 (
		_w5915_,
		_w5916_,
		_w5952_
	);
	LUT2 #(
		.INIT('h4)
	) name5491 (
		_w5912_,
		_w5952_,
		_w5953_
	);
	LUT2 #(
		.INIT('h4)
	) name5492 (
		_w5906_,
		_w5953_,
		_w5954_
	);
	LUT2 #(
		.INIT('h1)
	) name5493 (
		_w5933_,
		_w5951_,
		_w5955_
	);
	LUT2 #(
		.INIT('h8)
	) name5494 (
		_w5954_,
		_w5955_,
		_w5956_
	);
	LUT2 #(
		.INIT('h2)
	) name5495 (
		_w3450_,
		_w5956_,
		_w5957_
	);
	LUT2 #(
		.INIT('h1)
	) name5496 (
		_w5896_,
		_w5957_,
		_w5958_
	);
	LUT2 #(
		.INIT('h2)
	) name5497 (
		\P1_state_reg[0]/NET0131 ,
		_w5958_,
		_w5959_
	);
	LUT2 #(
		.INIT('h1)
	) name5498 (
		_w5895_,
		_w5959_,
		_w5960_
	);
	LUT2 #(
		.INIT('h8)
	) name5499 (
		_w3421_,
		_w5287_,
		_w5961_
	);
	LUT2 #(
		.INIT('h8)
	) name5500 (
		_w3733_,
		_w5961_,
		_w5962_
	);
	LUT2 #(
		.INIT('h2)
	) name5501 (
		\P2_reg1_reg[31]/NET0131 ,
		_w5962_,
		_w5963_
	);
	LUT2 #(
		.INIT('h8)
	) name5502 (
		_w3733_,
		_w5287_,
		_w5964_
	);
	LUT2 #(
		.INIT('h4)
	) name5503 (
		_w5864_,
		_w5964_,
		_w5965_
	);
	LUT2 #(
		.INIT('h1)
	) name5504 (
		_w5963_,
		_w5965_,
		_w5966_
	);
	LUT2 #(
		.INIT('h2)
	) name5505 (
		\P1_reg0_reg[24]/NET0131 ,
		_w3435_,
		_w5967_
	);
	LUT2 #(
		.INIT('h8)
	) name5506 (
		\P1_reg0_reg[24]/NET0131 ,
		_w3448_,
		_w5968_
	);
	LUT2 #(
		.INIT('h2)
	) name5507 (
		\P1_reg0_reg[24]/NET0131 ,
		_w4396_,
		_w5969_
	);
	LUT2 #(
		.INIT('h2)
	) name5508 (
		_w4396_,
		_w5172_,
		_w5970_
	);
	LUT2 #(
		.INIT('h1)
	) name5509 (
		_w5969_,
		_w5970_,
		_w5971_
	);
	LUT2 #(
		.INIT('h1)
	) name5510 (
		_w3563_,
		_w5971_,
		_w5972_
	);
	LUT2 #(
		.INIT('h8)
	) name5511 (
		_w4396_,
		_w5200_,
		_w5973_
	);
	LUT2 #(
		.INIT('h1)
	) name5512 (
		_w5969_,
		_w5973_,
		_w5974_
	);
	LUT2 #(
		.INIT('h2)
	) name5513 (
		_w1936_,
		_w5974_,
		_w5975_
	);
	LUT2 #(
		.INIT('h2)
	) name5514 (
		\P1_reg0_reg[24]/NET0131 ,
		_w4493_,
		_w5976_
	);
	LUT2 #(
		.INIT('h8)
	) name5515 (
		_w4396_,
		_w5206_,
		_w5977_
	);
	LUT2 #(
		.INIT('h8)
	) name5516 (
		_w4396_,
		_w5190_,
		_w5978_
	);
	LUT2 #(
		.INIT('h1)
	) name5517 (
		_w5969_,
		_w5978_,
		_w5979_
	);
	LUT2 #(
		.INIT('h2)
	) name5518 (
		_w3712_,
		_w5979_,
		_w5980_
	);
	LUT2 #(
		.INIT('h2)
	) name5519 (
		_w4396_,
		_w5184_,
		_w5981_
	);
	LUT2 #(
		.INIT('h1)
	) name5520 (
		_w5969_,
		_w5981_,
		_w5982_
	);
	LUT2 #(
		.INIT('h1)
	) name5521 (
		_w3677_,
		_w5982_,
		_w5983_
	);
	LUT2 #(
		.INIT('h1)
	) name5522 (
		_w5976_,
		_w5977_,
		_w5984_
	);
	LUT2 #(
		.INIT('h4)
	) name5523 (
		_w5980_,
		_w5984_,
		_w5985_
	);
	LUT2 #(
		.INIT('h4)
	) name5524 (
		_w5972_,
		_w5985_,
		_w5986_
	);
	LUT2 #(
		.INIT('h1)
	) name5525 (
		_w5975_,
		_w5983_,
		_w5987_
	);
	LUT2 #(
		.INIT('h8)
	) name5526 (
		_w5986_,
		_w5987_,
		_w5988_
	);
	LUT2 #(
		.INIT('h2)
	) name5527 (
		_w3450_,
		_w5988_,
		_w5989_
	);
	LUT2 #(
		.INIT('h1)
	) name5528 (
		_w5968_,
		_w5989_,
		_w5990_
	);
	LUT2 #(
		.INIT('h2)
	) name5529 (
		\P1_state_reg[0]/NET0131 ,
		_w5990_,
		_w5991_
	);
	LUT2 #(
		.INIT('h1)
	) name5530 (
		_w5967_,
		_w5991_,
		_w5992_
	);
	LUT2 #(
		.INIT('h2)
	) name5531 (
		\P1_reg0_reg[26]/NET0131 ,
		_w3435_,
		_w5993_
	);
	LUT2 #(
		.INIT('h8)
	) name5532 (
		\P1_reg0_reg[26]/NET0131 ,
		_w3448_,
		_w5994_
	);
	LUT2 #(
		.INIT('h2)
	) name5533 (
		\P1_reg0_reg[26]/NET0131 ,
		_w4396_,
		_w5995_
	);
	LUT2 #(
		.INIT('h2)
	) name5534 (
		_w4396_,
		_w5903_,
		_w5996_
	);
	LUT2 #(
		.INIT('h1)
	) name5535 (
		_w5995_,
		_w5996_,
		_w5997_
	);
	LUT2 #(
		.INIT('h2)
	) name5536 (
		_w1936_,
		_w5997_,
		_w5998_
	);
	LUT2 #(
		.INIT('h2)
	) name5537 (
		\P1_reg0_reg[26]/NET0131 ,
		_w4494_,
		_w5999_
	);
	LUT2 #(
		.INIT('h2)
	) name5538 (
		_w4396_,
		_w5911_,
		_w6000_
	);
	LUT2 #(
		.INIT('h2)
	) name5539 (
		_w4396_,
		_w5948_,
		_w6001_
	);
	LUT2 #(
		.INIT('h1)
	) name5540 (
		_w5995_,
		_w6001_,
		_w6002_
	);
	LUT2 #(
		.INIT('h1)
	) name5541 (
		_w3563_,
		_w6002_,
		_w6003_
	);
	LUT2 #(
		.INIT('h2)
	) name5542 (
		_w4396_,
		_w5930_,
		_w6004_
	);
	LUT2 #(
		.INIT('h1)
	) name5543 (
		_w5995_,
		_w6004_,
		_w6005_
	);
	LUT2 #(
		.INIT('h1)
	) name5544 (
		_w3677_,
		_w6005_,
		_w6006_
	);
	LUT2 #(
		.INIT('h1)
	) name5545 (
		_w5999_,
		_w6000_,
		_w6007_
	);
	LUT2 #(
		.INIT('h4)
	) name5546 (
		_w5998_,
		_w6007_,
		_w6008_
	);
	LUT2 #(
		.INIT('h1)
	) name5547 (
		_w6003_,
		_w6006_,
		_w6009_
	);
	LUT2 #(
		.INIT('h8)
	) name5548 (
		_w6008_,
		_w6009_,
		_w6010_
	);
	LUT2 #(
		.INIT('h2)
	) name5549 (
		_w3450_,
		_w6010_,
		_w6011_
	);
	LUT2 #(
		.INIT('h1)
	) name5550 (
		_w5994_,
		_w6011_,
		_w6012_
	);
	LUT2 #(
		.INIT('h2)
	) name5551 (
		\P1_state_reg[0]/NET0131 ,
		_w6012_,
		_w6013_
	);
	LUT2 #(
		.INIT('h1)
	) name5552 (
		_w5993_,
		_w6013_,
		_w6014_
	);
	LUT2 #(
		.INIT('h2)
	) name5553 (
		\P1_reg1_reg[22]/NET0131 ,
		_w3435_,
		_w6015_
	);
	LUT2 #(
		.INIT('h8)
	) name5554 (
		\P1_reg1_reg[22]/NET0131 ,
		_w3448_,
		_w6016_
	);
	LUT2 #(
		.INIT('h2)
	) name5555 (
		\P1_reg1_reg[22]/NET0131 ,
		_w4532_,
		_w6017_
	);
	LUT2 #(
		.INIT('h4)
	) name5556 (
		_w5499_,
		_w5918_,
		_w6018_
	);
	LUT2 #(
		.INIT('h4)
	) name5557 (
		_w5493_,
		_w5496_,
		_w6019_
	);
	LUT2 #(
		.INIT('h8)
	) name5558 (
		_w5486_,
		_w5918_,
		_w6020_
	);
	LUT2 #(
		.INIT('h4)
	) name5559 (
		_w6019_,
		_w6020_,
		_w6021_
	);
	LUT2 #(
		.INIT('h2)
	) name5560 (
		_w5923_,
		_w6018_,
		_w6022_
	);
	LUT2 #(
		.INIT('h4)
	) name5561 (
		_w6021_,
		_w6022_,
		_w6023_
	);
	LUT2 #(
		.INIT('h8)
	) name5562 (
		_w1838_,
		_w6023_,
		_w6024_
	);
	LUT2 #(
		.INIT('h1)
	) name5563 (
		_w1838_,
		_w6023_,
		_w6025_
	);
	LUT2 #(
		.INIT('h1)
	) name5564 (
		_w6024_,
		_w6025_,
		_w6026_
	);
	LUT2 #(
		.INIT('h8)
	) name5565 (
		_w4532_,
		_w6026_,
		_w6027_
	);
	LUT2 #(
		.INIT('h1)
	) name5566 (
		_w6017_,
		_w6027_,
		_w6028_
	);
	LUT2 #(
		.INIT('h1)
	) name5567 (
		_w3677_,
		_w6028_,
		_w6029_
	);
	LUT2 #(
		.INIT('h4)
	) name5568 (
		_w5522_,
		_w5934_,
		_w6030_
	);
	LUT2 #(
		.INIT('h4)
	) name5569 (
		_w5516_,
		_w5519_,
		_w6031_
	);
	LUT2 #(
		.INIT('h8)
	) name5570 (
		_w5508_,
		_w5934_,
		_w6032_
	);
	LUT2 #(
		.INIT('h4)
	) name5571 (
		_w6031_,
		_w6032_,
		_w6033_
	);
	LUT2 #(
		.INIT('h2)
	) name5572 (
		_w5939_,
		_w6030_,
		_w6034_
	);
	LUT2 #(
		.INIT('h4)
	) name5573 (
		_w6033_,
		_w6034_,
		_w6035_
	);
	LUT2 #(
		.INIT('h8)
	) name5574 (
		_w1838_,
		_w6035_,
		_w6036_
	);
	LUT2 #(
		.INIT('h1)
	) name5575 (
		_w1838_,
		_w6035_,
		_w6037_
	);
	LUT2 #(
		.INIT('h1)
	) name5576 (
		_w6036_,
		_w6037_,
		_w6038_
	);
	LUT2 #(
		.INIT('h2)
	) name5577 (
		_w4532_,
		_w6038_,
		_w6039_
	);
	LUT2 #(
		.INIT('h1)
	) name5578 (
		_w6017_,
		_w6039_,
		_w6040_
	);
	LUT2 #(
		.INIT('h1)
	) name5579 (
		_w3563_,
		_w6040_,
		_w6041_
	);
	LUT2 #(
		.INIT('h2)
	) name5580 (
		\P1_reg1_reg[22]/NET0131 ,
		_w4573_,
		_w6042_
	);
	LUT2 #(
		.INIT('h2)
	) name5581 (
		_w537_,
		_w1356_,
		_w6043_
	);
	LUT2 #(
		.INIT('h4)
	) name5582 (
		_w1318_,
		_w5795_,
		_w6044_
	);
	LUT2 #(
		.INIT('h2)
	) name5583 (
		_w1336_,
		_w6044_,
		_w6045_
	);
	LUT2 #(
		.INIT('h1)
	) name5584 (
		_w537_,
		_w5796_,
		_w6046_
	);
	LUT2 #(
		.INIT('h4)
	) name5585 (
		_w6045_,
		_w6046_,
		_w6047_
	);
	LUT2 #(
		.INIT('h1)
	) name5586 (
		_w6043_,
		_w6047_,
		_w6048_
	);
	LUT2 #(
		.INIT('h2)
	) name5587 (
		_w4532_,
		_w6048_,
		_w6049_
	);
	LUT2 #(
		.INIT('h1)
	) name5588 (
		_w6017_,
		_w6049_,
		_w6050_
	);
	LUT2 #(
		.INIT('h2)
	) name5589 (
		_w1936_,
		_w6050_,
		_w6051_
	);
	LUT2 #(
		.INIT('h4)
	) name5590 (
		_w1346_,
		_w3698_,
		_w6052_
	);
	LUT2 #(
		.INIT('h2)
	) name5591 (
		_w1309_,
		_w6052_,
		_w6053_
	);
	LUT2 #(
		.INIT('h1)
	) name5592 (
		_w3700_,
		_w6053_,
		_w6054_
	);
	LUT2 #(
		.INIT('h8)
	) name5593 (
		_w3712_,
		_w6054_,
		_w6055_
	);
	LUT2 #(
		.INIT('h8)
	) name5594 (
		_w1309_,
		_w1880_,
		_w6056_
	);
	LUT2 #(
		.INIT('h1)
	) name5595 (
		_w6055_,
		_w6056_,
		_w6057_
	);
	LUT2 #(
		.INIT('h2)
	) name5596 (
		_w4532_,
		_w6057_,
		_w6058_
	);
	LUT2 #(
		.INIT('h1)
	) name5597 (
		_w6042_,
		_w6058_,
		_w6059_
	);
	LUT2 #(
		.INIT('h4)
	) name5598 (
		_w6051_,
		_w6059_,
		_w6060_
	);
	LUT2 #(
		.INIT('h4)
	) name5599 (
		_w6029_,
		_w6060_,
		_w6061_
	);
	LUT2 #(
		.INIT('h4)
	) name5600 (
		_w6041_,
		_w6061_,
		_w6062_
	);
	LUT2 #(
		.INIT('h2)
	) name5601 (
		_w3450_,
		_w6062_,
		_w6063_
	);
	LUT2 #(
		.INIT('h1)
	) name5602 (
		_w6016_,
		_w6063_,
		_w6064_
	);
	LUT2 #(
		.INIT('h2)
	) name5603 (
		\P1_state_reg[0]/NET0131 ,
		_w6064_,
		_w6065_
	);
	LUT2 #(
		.INIT('h1)
	) name5604 (
		_w6015_,
		_w6065_,
		_w6066_
	);
	LUT2 #(
		.INIT('h2)
	) name5605 (
		\P1_reg1_reg[26]/NET0131 ,
		_w3435_,
		_w6067_
	);
	LUT2 #(
		.INIT('h8)
	) name5606 (
		\P1_reg1_reg[26]/NET0131 ,
		_w3448_,
		_w6068_
	);
	LUT2 #(
		.INIT('h2)
	) name5607 (
		\P1_reg1_reg[26]/NET0131 ,
		_w4532_,
		_w6069_
	);
	LUT2 #(
		.INIT('h2)
	) name5608 (
		_w4532_,
		_w5903_,
		_w6070_
	);
	LUT2 #(
		.INIT('h1)
	) name5609 (
		_w6069_,
		_w6070_,
		_w6071_
	);
	LUT2 #(
		.INIT('h2)
	) name5610 (
		_w1936_,
		_w6071_,
		_w6072_
	);
	LUT2 #(
		.INIT('h2)
	) name5611 (
		\P1_reg1_reg[26]/NET0131 ,
		_w4573_,
		_w6073_
	);
	LUT2 #(
		.INIT('h2)
	) name5612 (
		_w4532_,
		_w5911_,
		_w6074_
	);
	LUT2 #(
		.INIT('h2)
	) name5613 (
		_w4532_,
		_w5948_,
		_w6075_
	);
	LUT2 #(
		.INIT('h1)
	) name5614 (
		_w6069_,
		_w6075_,
		_w6076_
	);
	LUT2 #(
		.INIT('h1)
	) name5615 (
		_w3563_,
		_w6076_,
		_w6077_
	);
	LUT2 #(
		.INIT('h2)
	) name5616 (
		_w4532_,
		_w5930_,
		_w6078_
	);
	LUT2 #(
		.INIT('h1)
	) name5617 (
		_w6069_,
		_w6078_,
		_w6079_
	);
	LUT2 #(
		.INIT('h1)
	) name5618 (
		_w3677_,
		_w6079_,
		_w6080_
	);
	LUT2 #(
		.INIT('h1)
	) name5619 (
		_w6073_,
		_w6074_,
		_w6081_
	);
	LUT2 #(
		.INIT('h4)
	) name5620 (
		_w6072_,
		_w6081_,
		_w6082_
	);
	LUT2 #(
		.INIT('h1)
	) name5621 (
		_w6077_,
		_w6080_,
		_w6083_
	);
	LUT2 #(
		.INIT('h8)
	) name5622 (
		_w6082_,
		_w6083_,
		_w6084_
	);
	LUT2 #(
		.INIT('h2)
	) name5623 (
		_w3450_,
		_w6084_,
		_w6085_
	);
	LUT2 #(
		.INIT('h1)
	) name5624 (
		_w6068_,
		_w6085_,
		_w6086_
	);
	LUT2 #(
		.INIT('h2)
	) name5625 (
		\P1_state_reg[0]/NET0131 ,
		_w6086_,
		_w6087_
	);
	LUT2 #(
		.INIT('h1)
	) name5626 (
		_w6067_,
		_w6087_,
		_w6088_
	);
	LUT2 #(
		.INIT('h2)
	) name5627 (
		\P1_reg3_reg[12]/NET0131 ,
		\P1_state_reg[0]/NET0131 ,
		_w6089_
	);
	LUT2 #(
		.INIT('h8)
	) name5628 (
		_w1170_,
		_w1953_,
		_w6090_
	);
	LUT2 #(
		.INIT('h8)
	) name5629 (
		_w1170_,
		_w3448_,
		_w6091_
	);
	LUT2 #(
		.INIT('h2)
	) name5630 (
		_w1165_,
		_w4067_,
		_w6092_
	);
	LUT2 #(
		.INIT('h2)
	) name5631 (
		_w1170_,
		_w3980_,
		_w6093_
	);
	LUT2 #(
		.INIT('h2)
	) name5632 (
		_w1146_,
		_w4070_,
		_w6094_
	);
	LUT2 #(
		.INIT('h1)
	) name5633 (
		_w3583_,
		_w6094_,
		_w6095_
	);
	LUT2 #(
		.INIT('h1)
	) name5634 (
		_w537_,
		_w6095_,
		_w6096_
	);
	LUT2 #(
		.INIT('h8)
	) name5635 (
		_w537_,
		_w1207_,
		_w6097_
	);
	LUT2 #(
		.INIT('h1)
	) name5636 (
		_w6096_,
		_w6097_,
		_w6098_
	);
	LUT2 #(
		.INIT('h8)
	) name5637 (
		_w3980_,
		_w6098_,
		_w6099_
	);
	LUT2 #(
		.INIT('h1)
	) name5638 (
		_w6093_,
		_w6099_,
		_w6100_
	);
	LUT2 #(
		.INIT('h2)
	) name5639 (
		_w1936_,
		_w6100_,
		_w6101_
	);
	LUT2 #(
		.INIT('h2)
	) name5640 (
		_w1796_,
		_w4007_,
		_w6102_
	);
	LUT2 #(
		.INIT('h4)
	) name5641 (
		_w1796_,
		_w4007_,
		_w6103_
	);
	LUT2 #(
		.INIT('h1)
	) name5642 (
		_w6102_,
		_w6103_,
		_w6104_
	);
	LUT2 #(
		.INIT('h8)
	) name5643 (
		_w3980_,
		_w6104_,
		_w6105_
	);
	LUT2 #(
		.INIT('h1)
	) name5644 (
		_w6093_,
		_w6105_,
		_w6106_
	);
	LUT2 #(
		.INIT('h1)
	) name5645 (
		_w3563_,
		_w6106_,
		_w6107_
	);
	LUT2 #(
		.INIT('h2)
	) name5646 (
		_w1796_,
		_w4088_,
		_w6108_
	);
	LUT2 #(
		.INIT('h4)
	) name5647 (
		_w1796_,
		_w4088_,
		_w6109_
	);
	LUT2 #(
		.INIT('h1)
	) name5648 (
		_w6108_,
		_w6109_,
		_w6110_
	);
	LUT2 #(
		.INIT('h2)
	) name5649 (
		_w3980_,
		_w6110_,
		_w6111_
	);
	LUT2 #(
		.INIT('h1)
	) name5650 (
		_w6093_,
		_w6111_,
		_w6112_
	);
	LUT2 #(
		.INIT('h1)
	) name5651 (
		_w3677_,
		_w6112_,
		_w6113_
	);
	LUT2 #(
		.INIT('h4)
	) name5652 (
		_w1233_,
		_w3687_,
		_w6114_
	);
	LUT2 #(
		.INIT('h4)
	) name5653 (
		_w1198_,
		_w6114_,
		_w6115_
	);
	LUT2 #(
		.INIT('h2)
	) name5654 (
		_w1165_,
		_w6115_,
		_w6116_
	);
	LUT2 #(
		.INIT('h1)
	) name5655 (
		_w3690_,
		_w6116_,
		_w6117_
	);
	LUT2 #(
		.INIT('h8)
	) name5656 (
		_w3980_,
		_w6117_,
		_w6118_
	);
	LUT2 #(
		.INIT('h1)
	) name5657 (
		_w6093_,
		_w6118_,
		_w6119_
	);
	LUT2 #(
		.INIT('h2)
	) name5658 (
		_w3712_,
		_w6119_,
		_w6120_
	);
	LUT2 #(
		.INIT('h2)
	) name5659 (
		_w1170_,
		_w4064_,
		_w6121_
	);
	LUT2 #(
		.INIT('h1)
	) name5660 (
		_w6092_,
		_w6121_,
		_w6122_
	);
	LUT2 #(
		.INIT('h4)
	) name5661 (
		_w6120_,
		_w6122_,
		_w6123_
	);
	LUT2 #(
		.INIT('h4)
	) name5662 (
		_w6107_,
		_w6123_,
		_w6124_
	);
	LUT2 #(
		.INIT('h4)
	) name5663 (
		_w6113_,
		_w6124_,
		_w6125_
	);
	LUT2 #(
		.INIT('h4)
	) name5664 (
		_w6101_,
		_w6125_,
		_w6126_
	);
	LUT2 #(
		.INIT('h2)
	) name5665 (
		_w3450_,
		_w6126_,
		_w6127_
	);
	LUT2 #(
		.INIT('h1)
	) name5666 (
		_w6091_,
		_w6127_,
		_w6128_
	);
	LUT2 #(
		.INIT('h2)
	) name5667 (
		\P1_state_reg[0]/NET0131 ,
		_w6128_,
		_w6129_
	);
	LUT2 #(
		.INIT('h1)
	) name5668 (
		_w6089_,
		_w6090_,
		_w6130_
	);
	LUT2 #(
		.INIT('h4)
	) name5669 (
		_w6129_,
		_w6130_,
		_w6131_
	);
	LUT2 #(
		.INIT('h2)
	) name5670 (
		\P1_reg3_reg[16]/NET0131 ,
		\P1_state_reg[0]/NET0131 ,
		_w6132_
	);
	LUT2 #(
		.INIT('h8)
	) name5671 (
		_w1471_,
		_w1953_,
		_w6133_
	);
	LUT2 #(
		.INIT('h8)
	) name5672 (
		_w1471_,
		_w3448_,
		_w6134_
	);
	LUT2 #(
		.INIT('h2)
	) name5673 (
		_w1471_,
		_w4910_,
		_w6135_
	);
	LUT2 #(
		.INIT('h2)
	) name5674 (
		_w1471_,
		_w3980_,
		_w6136_
	);
	LUT2 #(
		.INIT('h4)
	) name5675 (
		_w4007_,
		_w4010_,
		_w6137_
	);
	LUT2 #(
		.INIT('h2)
	) name5676 (
		_w4021_,
		_w6137_,
		_w6138_
	);
	LUT2 #(
		.INIT('h8)
	) name5677 (
		_w1785_,
		_w6138_,
		_w6139_
	);
	LUT2 #(
		.INIT('h1)
	) name5678 (
		_w1785_,
		_w6138_,
		_w6140_
	);
	LUT2 #(
		.INIT('h1)
	) name5679 (
		_w6139_,
		_w6140_,
		_w6141_
	);
	LUT2 #(
		.INIT('h2)
	) name5680 (
		_w3980_,
		_w6141_,
		_w6142_
	);
	LUT2 #(
		.INIT('h1)
	) name5681 (
		_w6136_,
		_w6142_,
		_w6143_
	);
	LUT2 #(
		.INIT('h1)
	) name5682 (
		_w3563_,
		_w6143_,
		_w6144_
	);
	LUT2 #(
		.INIT('h2)
	) name5683 (
		_w1452_,
		_w4073_,
		_w6145_
	);
	LUT2 #(
		.INIT('h1)
	) name5684 (
		_w5195_,
		_w6145_,
		_w6146_
	);
	LUT2 #(
		.INIT('h1)
	) name5685 (
		_w537_,
		_w6146_,
		_w6147_
	);
	LUT2 #(
		.INIT('h8)
	) name5686 (
		_w537_,
		_w1094_,
		_w6148_
	);
	LUT2 #(
		.INIT('h1)
	) name5687 (
		_w6147_,
		_w6148_,
		_w6149_
	);
	LUT2 #(
		.INIT('h8)
	) name5688 (
		_w3980_,
		_w6149_,
		_w6150_
	);
	LUT2 #(
		.INIT('h1)
	) name5689 (
		_w6136_,
		_w6150_,
		_w6151_
	);
	LUT2 #(
		.INIT('h2)
	) name5690 (
		_w1936_,
		_w6151_,
		_w6152_
	);
	LUT2 #(
		.INIT('h4)
	) name5691 (
		_w1750_,
		_w1785_,
		_w6153_
	);
	LUT2 #(
		.INIT('h2)
	) name5692 (
		_w1750_,
		_w1785_,
		_w6154_
	);
	LUT2 #(
		.INIT('h1)
	) name5693 (
		_w6153_,
		_w6154_,
		_w6155_
	);
	LUT2 #(
		.INIT('h2)
	) name5694 (
		_w3980_,
		_w6155_,
		_w6156_
	);
	LUT2 #(
		.INIT('h1)
	) name5695 (
		_w6136_,
		_w6156_,
		_w6157_
	);
	LUT2 #(
		.INIT('h1)
	) name5696 (
		_w3677_,
		_w6157_,
		_w6158_
	);
	LUT2 #(
		.INIT('h2)
	) name5697 (
		_w1466_,
		_w5441_,
		_w6159_
	);
	LUT2 #(
		.INIT('h1)
	) name5698 (
		_w5442_,
		_w6159_,
		_w6160_
	);
	LUT2 #(
		.INIT('h8)
	) name5699 (
		_w3712_,
		_w6160_,
		_w6161_
	);
	LUT2 #(
		.INIT('h8)
	) name5700 (
		_w3980_,
		_w6161_,
		_w6162_
	);
	LUT2 #(
		.INIT('h2)
	) name5701 (
		_w1466_,
		_w4067_,
		_w6163_
	);
	LUT2 #(
		.INIT('h1)
	) name5702 (
		_w6135_,
		_w6163_,
		_w6164_
	);
	LUT2 #(
		.INIT('h4)
	) name5703 (
		_w6162_,
		_w6164_,
		_w6165_
	);
	LUT2 #(
		.INIT('h4)
	) name5704 (
		_w6158_,
		_w6165_,
		_w6166_
	);
	LUT2 #(
		.INIT('h4)
	) name5705 (
		_w6144_,
		_w6166_,
		_w6167_
	);
	LUT2 #(
		.INIT('h4)
	) name5706 (
		_w6152_,
		_w6167_,
		_w6168_
	);
	LUT2 #(
		.INIT('h2)
	) name5707 (
		_w3450_,
		_w6168_,
		_w6169_
	);
	LUT2 #(
		.INIT('h1)
	) name5708 (
		_w6134_,
		_w6169_,
		_w6170_
	);
	LUT2 #(
		.INIT('h2)
	) name5709 (
		\P1_state_reg[0]/NET0131 ,
		_w6170_,
		_w6171_
	);
	LUT2 #(
		.INIT('h1)
	) name5710 (
		_w6132_,
		_w6133_,
		_w6172_
	);
	LUT2 #(
		.INIT('h4)
	) name5711 (
		_w6171_,
		_w6172_,
		_w6173_
	);
	LUT2 #(
		.INIT('h4)
	) name5712 (
		\P1_state_reg[0]/NET0131 ,
		\P2_reg3_reg[12]/NET0131 ,
		_w6174_
	);
	LUT2 #(
		.INIT('h8)
	) name5713 (
		_w2709_,
		_w3976_,
		_w6175_
	);
	LUT2 #(
		.INIT('h8)
	) name5714 (
		_w2024_,
		_w2709_,
		_w6176_
	);
	LUT2 #(
		.INIT('h2)
	) name5715 (
		_w2709_,
		_w5698_,
		_w6177_
	);
	LUT2 #(
		.INIT('h2)
	) name5716 (
		_w2709_,
		_w3788_,
		_w6178_
	);
	LUT2 #(
		.INIT('h4)
	) name5717 (
		_w2688_,
		_w3383_,
		_w6179_
	);
	LUT2 #(
		.INIT('h4)
	) name5718 (
		_w2715_,
		_w6179_,
		_w6180_
	);
	LUT2 #(
		.INIT('h2)
	) name5719 (
		_w2880_,
		_w6180_,
		_w6181_
	);
	LUT2 #(
		.INIT('h4)
	) name5720 (
		_w2880_,
		_w6180_,
		_w6182_
	);
	LUT2 #(
		.INIT('h1)
	) name5721 (
		_w6181_,
		_w6182_,
		_w6183_
	);
	LUT2 #(
		.INIT('h1)
	) name5722 (
		_w2058_,
		_w6183_,
		_w6184_
	);
	LUT2 #(
		.INIT('h8)
	) name5723 (
		_w2058_,
		_w2688_,
		_w6185_
	);
	LUT2 #(
		.INIT('h1)
	) name5724 (
		_w6184_,
		_w6185_,
		_w6186_
	);
	LUT2 #(
		.INIT('h8)
	) name5725 (
		_w3788_,
		_w6186_,
		_w6187_
	);
	LUT2 #(
		.INIT('h1)
	) name5726 (
		_w6178_,
		_w6187_,
		_w6188_
	);
	LUT2 #(
		.INIT('h2)
	) name5727 (
		_w3411_,
		_w6188_,
		_w6189_
	);
	LUT2 #(
		.INIT('h4)
	) name5728 (
		_w3893_,
		_w4212_,
		_w6190_
	);
	LUT2 #(
		.INIT('h2)
	) name5729 (
		_w3893_,
		_w4212_,
		_w6191_
	);
	LUT2 #(
		.INIT('h1)
	) name5730 (
		_w6190_,
		_w6191_,
		_w6192_
	);
	LUT2 #(
		.INIT('h8)
	) name5731 (
		_w3788_,
		_w6192_,
		_w6193_
	);
	LUT2 #(
		.INIT('h1)
	) name5732 (
		_w6178_,
		_w6193_,
		_w6194_
	);
	LUT2 #(
		.INIT('h1)
	) name5733 (
		_w3177_,
		_w6194_,
		_w6195_
	);
	LUT2 #(
		.INIT('h4)
	) name5734 (
		_w3839_,
		_w4212_,
		_w6196_
	);
	LUT2 #(
		.INIT('h2)
	) name5735 (
		_w3839_,
		_w4212_,
		_w6197_
	);
	LUT2 #(
		.INIT('h1)
	) name5736 (
		_w6196_,
		_w6197_,
		_w6198_
	);
	LUT2 #(
		.INIT('h2)
	) name5737 (
		_w3788_,
		_w6198_,
		_w6199_
	);
	LUT2 #(
		.INIT('h1)
	) name5738 (
		_w6178_,
		_w6199_,
		_w6200_
	);
	LUT2 #(
		.INIT('h1)
	) name5739 (
		_w3320_,
		_w6200_,
		_w6201_
	);
	LUT2 #(
		.INIT('h2)
	) name5740 (
		_w2731_,
		_w3336_,
		_w6202_
	);
	LUT2 #(
		.INIT('h1)
	) name5741 (
		_w3337_,
		_w6202_,
		_w6203_
	);
	LUT2 #(
		.INIT('h8)
	) name5742 (
		_w3355_,
		_w6203_,
		_w6204_
	);
	LUT2 #(
		.INIT('h8)
	) name5743 (
		_w3788_,
		_w6204_,
		_w6205_
	);
	LUT2 #(
		.INIT('h2)
	) name5744 (
		_w2731_,
		_w3965_,
		_w6206_
	);
	LUT2 #(
		.INIT('h1)
	) name5745 (
		_w6177_,
		_w6206_,
		_w6207_
	);
	LUT2 #(
		.INIT('h4)
	) name5746 (
		_w6205_,
		_w6207_,
		_w6208_
	);
	LUT2 #(
		.INIT('h4)
	) name5747 (
		_w6195_,
		_w6208_,
		_w6209_
	);
	LUT2 #(
		.INIT('h4)
	) name5748 (
		_w6201_,
		_w6209_,
		_w6210_
	);
	LUT2 #(
		.INIT('h4)
	) name5749 (
		_w6189_,
		_w6210_,
		_w6211_
	);
	LUT2 #(
		.INIT('h2)
	) name5750 (
		_w2026_,
		_w6211_,
		_w6212_
	);
	LUT2 #(
		.INIT('h1)
	) name5751 (
		_w6176_,
		_w6212_,
		_w6213_
	);
	LUT2 #(
		.INIT('h2)
	) name5752 (
		\P1_state_reg[0]/NET0131 ,
		_w6213_,
		_w6214_
	);
	LUT2 #(
		.INIT('h1)
	) name5753 (
		_w6174_,
		_w6175_,
		_w6215_
	);
	LUT2 #(
		.INIT('h4)
	) name5754 (
		_w6214_,
		_w6215_,
		_w6216_
	);
	LUT2 #(
		.INIT('h8)
	) name5755 (
		_w2797_,
		_w3976_,
		_w6217_
	);
	LUT2 #(
		.INIT('h4)
	) name5756 (
		\P1_state_reg[0]/NET0131 ,
		\P2_reg3_reg[16]/NET0131 ,
		_w6218_
	);
	LUT2 #(
		.INIT('h8)
	) name5757 (
		_w2024_,
		_w2797_,
		_w6219_
	);
	LUT2 #(
		.INIT('h2)
	) name5758 (
		_w2797_,
		_w3962_,
		_w6220_
	);
	LUT2 #(
		.INIT('h2)
	) name5759 (
		_w2797_,
		_w3788_,
		_w6221_
	);
	LUT2 #(
		.INIT('h4)
	) name5760 (
		_w3893_,
		_w3896_,
		_w6222_
	);
	LUT2 #(
		.INIT('h2)
	) name5761 (
		_w3907_,
		_w6222_,
		_w6223_
	);
	LUT2 #(
		.INIT('h8)
	) name5762 (
		_w4211_,
		_w6223_,
		_w6224_
	);
	LUT2 #(
		.INIT('h1)
	) name5763 (
		_w4211_,
		_w6223_,
		_w6225_
	);
	LUT2 #(
		.INIT('h1)
	) name5764 (
		_w6224_,
		_w6225_,
		_w6226_
	);
	LUT2 #(
		.INIT('h2)
	) name5765 (
		_w3788_,
		_w6226_,
		_w6227_
	);
	LUT2 #(
		.INIT('h1)
	) name5766 (
		_w6221_,
		_w6227_,
		_w6228_
	);
	LUT2 #(
		.INIT('h1)
	) name5767 (
		_w3177_,
		_w6228_,
		_w6229_
	);
	LUT2 #(
		.INIT('h2)
	) name5768 (
		_w2379_,
		_w5565_,
		_w6230_
	);
	LUT2 #(
		.INIT('h1)
	) name5769 (
		_w5566_,
		_w6230_,
		_w6231_
	);
	LUT2 #(
		.INIT('h1)
	) name5770 (
		_w2058_,
		_w6231_,
		_w6232_
	);
	LUT2 #(
		.INIT('h8)
	) name5771 (
		_w2058_,
		_w2828_,
		_w6233_
	);
	LUT2 #(
		.INIT('h1)
	) name5772 (
		_w6232_,
		_w6233_,
		_w6234_
	);
	LUT2 #(
		.INIT('h8)
	) name5773 (
		_w3788_,
		_w6234_,
		_w6235_
	);
	LUT2 #(
		.INIT('h1)
	) name5774 (
		_w6221_,
		_w6235_,
		_w6236_
	);
	LUT2 #(
		.INIT('h2)
	) name5775 (
		_w3411_,
		_w6236_,
		_w6237_
	);
	LUT2 #(
		.INIT('h2)
	) name5776 (
		_w2818_,
		_w3965_,
		_w6238_
	);
	LUT2 #(
		.INIT('h2)
	) name5777 (
		_w2818_,
		_w5574_,
		_w6239_
	);
	LUT2 #(
		.INIT('h1)
	) name5778 (
		_w5575_,
		_w6239_,
		_w6240_
	);
	LUT2 #(
		.INIT('h8)
	) name5779 (
		_w3788_,
		_w6240_,
		_w6241_
	);
	LUT2 #(
		.INIT('h1)
	) name5780 (
		_w6221_,
		_w6241_,
		_w6242_
	);
	LUT2 #(
		.INIT('h2)
	) name5781 (
		_w3355_,
		_w6242_,
		_w6243_
	);
	LUT2 #(
		.INIT('h4)
	) name5782 (
		_w4169_,
		_w4211_,
		_w6244_
	);
	LUT2 #(
		.INIT('h2)
	) name5783 (
		_w4169_,
		_w4211_,
		_w6245_
	);
	LUT2 #(
		.INIT('h1)
	) name5784 (
		_w6244_,
		_w6245_,
		_w6246_
	);
	LUT2 #(
		.INIT('h2)
	) name5785 (
		_w3788_,
		_w6246_,
		_w6247_
	);
	LUT2 #(
		.INIT('h1)
	) name5786 (
		_w6221_,
		_w6247_,
		_w6248_
	);
	LUT2 #(
		.INIT('h1)
	) name5787 (
		_w3320_,
		_w6248_,
		_w6249_
	);
	LUT2 #(
		.INIT('h1)
	) name5788 (
		_w6220_,
		_w6238_,
		_w6250_
	);
	LUT2 #(
		.INIT('h4)
	) name5789 (
		_w6243_,
		_w6250_,
		_w6251_
	);
	LUT2 #(
		.INIT('h4)
	) name5790 (
		_w6249_,
		_w6251_,
		_w6252_
	);
	LUT2 #(
		.INIT('h1)
	) name5791 (
		_w6229_,
		_w6237_,
		_w6253_
	);
	LUT2 #(
		.INIT('h8)
	) name5792 (
		_w6252_,
		_w6253_,
		_w6254_
	);
	LUT2 #(
		.INIT('h2)
	) name5793 (
		_w2026_,
		_w6254_,
		_w6255_
	);
	LUT2 #(
		.INIT('h1)
	) name5794 (
		_w6219_,
		_w6255_,
		_w6256_
	);
	LUT2 #(
		.INIT('h2)
	) name5795 (
		\P1_state_reg[0]/NET0131 ,
		_w6256_,
		_w6257_
	);
	LUT2 #(
		.INIT('h1)
	) name5796 (
		_w6217_,
		_w6218_,
		_w6258_
	);
	LUT2 #(
		.INIT('h4)
	) name5797 (
		_w6257_,
		_w6258_,
		_w6259_
	);
	LUT2 #(
		.INIT('h2)
	) name5798 (
		\P1_reg3_reg[22]/NET0131 ,
		\P1_state_reg[0]/NET0131 ,
		_w6260_
	);
	LUT2 #(
		.INIT('h8)
	) name5799 (
		_w1314_,
		_w1953_,
		_w6261_
	);
	LUT2 #(
		.INIT('h8)
	) name5800 (
		_w1314_,
		_w3448_,
		_w6262_
	);
	LUT2 #(
		.INIT('h2)
	) name5801 (
		_w1314_,
		_w3980_,
		_w6263_
	);
	LUT2 #(
		.INIT('h2)
	) name5802 (
		_w3980_,
		_w6038_,
		_w6264_
	);
	LUT2 #(
		.INIT('h1)
	) name5803 (
		_w6263_,
		_w6264_,
		_w6265_
	);
	LUT2 #(
		.INIT('h1)
	) name5804 (
		_w3563_,
		_w6265_,
		_w6266_
	);
	LUT2 #(
		.INIT('h8)
	) name5805 (
		_w3980_,
		_w6026_,
		_w6267_
	);
	LUT2 #(
		.INIT('h1)
	) name5806 (
		_w6263_,
		_w6267_,
		_w6268_
	);
	LUT2 #(
		.INIT('h1)
	) name5807 (
		_w3677_,
		_w6268_,
		_w6269_
	);
	LUT2 #(
		.INIT('h2)
	) name5808 (
		_w1314_,
		_w4910_,
		_w6270_
	);
	LUT2 #(
		.INIT('h2)
	) name5809 (
		_w3980_,
		_w6048_,
		_w6271_
	);
	LUT2 #(
		.INIT('h1)
	) name5810 (
		_w6263_,
		_w6271_,
		_w6272_
	);
	LUT2 #(
		.INIT('h2)
	) name5811 (
		_w1936_,
		_w6272_,
		_w6273_
	);
	LUT2 #(
		.INIT('h8)
	) name5812 (
		_w3980_,
		_w6055_,
		_w6274_
	);
	LUT2 #(
		.INIT('h2)
	) name5813 (
		_w1309_,
		_w4067_,
		_w6275_
	);
	LUT2 #(
		.INIT('h1)
	) name5814 (
		_w6270_,
		_w6275_,
		_w6276_
	);
	LUT2 #(
		.INIT('h4)
	) name5815 (
		_w6274_,
		_w6276_,
		_w6277_
	);
	LUT2 #(
		.INIT('h4)
	) name5816 (
		_w6273_,
		_w6277_,
		_w6278_
	);
	LUT2 #(
		.INIT('h4)
	) name5817 (
		_w6266_,
		_w6278_,
		_w6279_
	);
	LUT2 #(
		.INIT('h4)
	) name5818 (
		_w6269_,
		_w6279_,
		_w6280_
	);
	LUT2 #(
		.INIT('h2)
	) name5819 (
		_w3450_,
		_w6280_,
		_w6281_
	);
	LUT2 #(
		.INIT('h1)
	) name5820 (
		_w6262_,
		_w6281_,
		_w6282_
	);
	LUT2 #(
		.INIT('h2)
	) name5821 (
		\P1_state_reg[0]/NET0131 ,
		_w6282_,
		_w6283_
	);
	LUT2 #(
		.INIT('h1)
	) name5822 (
		_w6260_,
		_w6261_,
		_w6284_
	);
	LUT2 #(
		.INIT('h4)
	) name5823 (
		_w6283_,
		_w6284_,
		_w6285_
	);
	LUT2 #(
		.INIT('h8)
	) name5824 (
		_w2024_,
		_w3126_,
		_w6286_
	);
	LUT2 #(
		.INIT('h2)
	) name5825 (
		_w3121_,
		_w3965_,
		_w6287_
	);
	LUT2 #(
		.INIT('h8)
	) name5826 (
		_w2921_,
		_w4216_,
		_w6288_
	);
	LUT2 #(
		.INIT('h1)
	) name5827 (
		_w2921_,
		_w4216_,
		_w6289_
	);
	LUT2 #(
		.INIT('h1)
	) name5828 (
		_w6288_,
		_w6289_,
		_w6290_
	);
	LUT2 #(
		.INIT('h8)
	) name5829 (
		_w3788_,
		_w6290_,
		_w6291_
	);
	LUT2 #(
		.INIT('h1)
	) name5830 (
		_w3126_,
		_w3788_,
		_w6292_
	);
	LUT2 #(
		.INIT('h1)
	) name5831 (
		_w3177_,
		_w6292_,
		_w6293_
	);
	LUT2 #(
		.INIT('h4)
	) name5832 (
		_w6291_,
		_w6293_,
		_w6294_
	);
	LUT2 #(
		.INIT('h8)
	) name5833 (
		_w2058_,
		_w2368_,
		_w6295_
	);
	LUT2 #(
		.INIT('h2)
	) name5834 (
		_w3112_,
		_w3394_,
		_w6296_
	);
	LUT2 #(
		.INIT('h1)
	) name5835 (
		_w5773_,
		_w6296_,
		_w6297_
	);
	LUT2 #(
		.INIT('h1)
	) name5836 (
		_w2058_,
		_w6297_,
		_w6298_
	);
	LUT2 #(
		.INIT('h2)
	) name5837 (
		_w3411_,
		_w6295_,
		_w6299_
	);
	LUT2 #(
		.INIT('h4)
	) name5838 (
		_w6298_,
		_w6299_,
		_w6300_
	);
	LUT2 #(
		.INIT('h2)
	) name5839 (
		_w3121_,
		_w5765_,
		_w6301_
	);
	LUT2 #(
		.INIT('h2)
	) name5840 (
		_w3355_,
		_w5766_,
		_w6302_
	);
	LUT2 #(
		.INIT('h4)
	) name5841 (
		_w6301_,
		_w6302_,
		_w6303_
	);
	LUT2 #(
		.INIT('h1)
	) name5842 (
		_w3304_,
		_w4216_,
		_w6304_
	);
	LUT2 #(
		.INIT('h8)
	) name5843 (
		_w3304_,
		_w4216_,
		_w6305_
	);
	LUT2 #(
		.INIT('h1)
	) name5844 (
		_w3320_,
		_w6304_,
		_w6306_
	);
	LUT2 #(
		.INIT('h4)
	) name5845 (
		_w6305_,
		_w6306_,
		_w6307_
	);
	LUT2 #(
		.INIT('h1)
	) name5846 (
		_w6300_,
		_w6307_,
		_w6308_
	);
	LUT2 #(
		.INIT('h4)
	) name5847 (
		_w6303_,
		_w6308_,
		_w6309_
	);
	LUT2 #(
		.INIT('h2)
	) name5848 (
		_w3788_,
		_w6309_,
		_w6310_
	);
	LUT2 #(
		.INIT('h1)
	) name5849 (
		_w3320_,
		_w3788_,
		_w6311_
	);
	LUT2 #(
		.INIT('h2)
	) name5850 (
		_w3962_,
		_w6311_,
		_w6312_
	);
	LUT2 #(
		.INIT('h2)
	) name5851 (
		_w3745_,
		_w3788_,
		_w6313_
	);
	LUT2 #(
		.INIT('h2)
	) name5852 (
		_w6312_,
		_w6313_,
		_w6314_
	);
	LUT2 #(
		.INIT('h2)
	) name5853 (
		_w3126_,
		_w6314_,
		_w6315_
	);
	LUT2 #(
		.INIT('h1)
	) name5854 (
		_w6287_,
		_w6315_,
		_w6316_
	);
	LUT2 #(
		.INIT('h4)
	) name5855 (
		_w6294_,
		_w6316_,
		_w6317_
	);
	LUT2 #(
		.INIT('h4)
	) name5856 (
		_w6310_,
		_w6317_,
		_w6318_
	);
	LUT2 #(
		.INIT('h2)
	) name5857 (
		_w2026_,
		_w6318_,
		_w6319_
	);
	LUT2 #(
		.INIT('h1)
	) name5858 (
		_w6286_,
		_w6319_,
		_w6320_
	);
	LUT2 #(
		.INIT('h2)
	) name5859 (
		\P1_state_reg[0]/NET0131 ,
		_w6320_,
		_w6321_
	);
	LUT2 #(
		.INIT('h8)
	) name5860 (
		_w3126_,
		_w3976_,
		_w6322_
	);
	LUT2 #(
		.INIT('h4)
	) name5861 (
		\P1_state_reg[0]/NET0131 ,
		\P2_reg3_reg[21]/NET0131 ,
		_w6323_
	);
	LUT2 #(
		.INIT('h1)
	) name5862 (
		_w6322_,
		_w6323_,
		_w6324_
	);
	LUT2 #(
		.INIT('h4)
	) name5863 (
		_w6321_,
		_w6324_,
		_w6325_
	);
	LUT2 #(
		.INIT('h2)
	) name5864 (
		\P2_reg2_reg[18]/NET0131 ,
		_w1983_,
		_w6326_
	);
	LUT2 #(
		.INIT('h8)
	) name5865 (
		\P2_reg2_reg[18]/NET0131 ,
		_w2024_,
		_w6327_
	);
	LUT2 #(
		.INIT('h2)
	) name5866 (
		\P2_reg2_reg[18]/NET0131 ,
		_w3774_,
		_w6328_
	);
	LUT2 #(
		.INIT('h2)
	) name5867 (
		\P2_reg2_reg[18]/NET0131 ,
		_w3758_,
		_w6329_
	);
	LUT2 #(
		.INIT('h2)
	) name5868 (
		_w2433_,
		_w5577_,
		_w6330_
	);
	LUT2 #(
		.INIT('h1)
	) name5869 (
		_w3343_,
		_w6330_,
		_w6331_
	);
	LUT2 #(
		.INIT('h8)
	) name5870 (
		_w3758_,
		_w6331_,
		_w6332_
	);
	LUT2 #(
		.INIT('h1)
	) name5871 (
		_w6329_,
		_w6332_,
		_w6333_
	);
	LUT2 #(
		.INIT('h2)
	) name5872 (
		_w3355_,
		_w6333_,
		_w6334_
	);
	LUT2 #(
		.INIT('h2)
	) name5873 (
		_w4218_,
		_w4750_,
		_w6335_
	);
	LUT2 #(
		.INIT('h4)
	) name5874 (
		_w4218_,
		_w4750_,
		_w6336_
	);
	LUT2 #(
		.INIT('h1)
	) name5875 (
		_w6335_,
		_w6336_,
		_w6337_
	);
	LUT2 #(
		.INIT('h8)
	) name5876 (
		_w3758_,
		_w6337_,
		_w6338_
	);
	LUT2 #(
		.INIT('h1)
	) name5877 (
		_w6329_,
		_w6338_,
		_w6339_
	);
	LUT2 #(
		.INIT('h1)
	) name5878 (
		_w3177_,
		_w6339_,
		_w6340_
	);
	LUT2 #(
		.INIT('h2)
	) name5879 (
		_w4218_,
		_w4719_,
		_w6341_
	);
	LUT2 #(
		.INIT('h4)
	) name5880 (
		_w4218_,
		_w4719_,
		_w6342_
	);
	LUT2 #(
		.INIT('h1)
	) name5881 (
		_w6341_,
		_w6342_,
		_w6343_
	);
	LUT2 #(
		.INIT('h2)
	) name5882 (
		_w3758_,
		_w6343_,
		_w6344_
	);
	LUT2 #(
		.INIT('h1)
	) name5883 (
		_w6329_,
		_w6344_,
		_w6345_
	);
	LUT2 #(
		.INIT('h1)
	) name5884 (
		_w3320_,
		_w6345_,
		_w6346_
	);
	LUT2 #(
		.INIT('h2)
	) name5885 (
		_w2311_,
		_w5563_,
		_w6347_
	);
	LUT2 #(
		.INIT('h1)
	) name5886 (
		_w5618_,
		_w6347_,
		_w6348_
	);
	LUT2 #(
		.INIT('h1)
	) name5887 (
		_w2058_,
		_w6348_,
		_w6349_
	);
	LUT2 #(
		.INIT('h8)
	) name5888 (
		_w2058_,
		_w2379_,
		_w6350_
	);
	LUT2 #(
		.INIT('h1)
	) name5889 (
		_w6349_,
		_w6350_,
		_w6351_
	);
	LUT2 #(
		.INIT('h8)
	) name5890 (
		_w3758_,
		_w6351_,
		_w6352_
	);
	LUT2 #(
		.INIT('h1)
	) name5891 (
		_w6329_,
		_w6352_,
		_w6353_
	);
	LUT2 #(
		.INIT('h2)
	) name5892 (
		_w3411_,
		_w6353_,
		_w6354_
	);
	LUT2 #(
		.INIT('h8)
	) name5893 (
		_w2438_,
		_w3420_,
		_w6355_
	);
	LUT2 #(
		.INIT('h8)
	) name5894 (
		_w2433_,
		_w3358_,
		_w6356_
	);
	LUT2 #(
		.INIT('h8)
	) name5895 (
		_w3758_,
		_w6356_,
		_w6357_
	);
	LUT2 #(
		.INIT('h1)
	) name5896 (
		_w6328_,
		_w6355_,
		_w6358_
	);
	LUT2 #(
		.INIT('h4)
	) name5897 (
		_w6357_,
		_w6358_,
		_w6359_
	);
	LUT2 #(
		.INIT('h4)
	) name5898 (
		_w6354_,
		_w6359_,
		_w6360_
	);
	LUT2 #(
		.INIT('h4)
	) name5899 (
		_w6340_,
		_w6360_,
		_w6361_
	);
	LUT2 #(
		.INIT('h4)
	) name5900 (
		_w6346_,
		_w6361_,
		_w6362_
	);
	LUT2 #(
		.INIT('h4)
	) name5901 (
		_w6334_,
		_w6362_,
		_w6363_
	);
	LUT2 #(
		.INIT('h2)
	) name5902 (
		_w2026_,
		_w6363_,
		_w6364_
	);
	LUT2 #(
		.INIT('h1)
	) name5903 (
		_w6327_,
		_w6364_,
		_w6365_
	);
	LUT2 #(
		.INIT('h2)
	) name5904 (
		\P1_state_reg[0]/NET0131 ,
		_w6365_,
		_w6366_
	);
	LUT2 #(
		.INIT('h1)
	) name5905 (
		_w6326_,
		_w6366_,
		_w6367_
	);
	LUT2 #(
		.INIT('h8)
	) name5906 (
		_w4532_,
		_w5812_,
		_w6368_
	);
	LUT2 #(
		.INIT('h4)
	) name5907 (
		_w5809_,
		_w6368_,
		_w6369_
	);
	LUT2 #(
		.INIT('h8)
	) name5908 (
		_w4491_,
		_w6368_,
		_w6370_
	);
	LUT2 #(
		.INIT('h2)
	) name5909 (
		\P1_reg1_reg[31]/NET0131 ,
		_w6370_,
		_w6371_
	);
	LUT2 #(
		.INIT('h1)
	) name5910 (
		_w6369_,
		_w6371_,
		_w6372_
	);
	LUT2 #(
		.INIT('h2)
	) name5911 (
		\P2_reg0_reg[22]/NET0131 ,
		_w1983_,
		_w6373_
	);
	LUT2 #(
		.INIT('h8)
	) name5912 (
		\P2_reg0_reg[22]/NET0131 ,
		_w2024_,
		_w6374_
	);
	LUT2 #(
		.INIT('h8)
	) name5913 (
		_w3411_,
		_w5779_,
		_w6375_
	);
	LUT2 #(
		.INIT('h8)
	) name5914 (
		_w3355_,
		_w5769_,
		_w6376_
	);
	LUT2 #(
		.INIT('h8)
	) name5915 (
		_w3102_,
		_w3358_,
		_w6377_
	);
	LUT2 #(
		.INIT('h1)
	) name5916 (
		_w6375_,
		_w6377_,
		_w6378_
	);
	LUT2 #(
		.INIT('h4)
	) name5917 (
		_w6376_,
		_w6378_,
		_w6379_
	);
	LUT2 #(
		.INIT('h2)
	) name5918 (
		_w2040_,
		_w6379_,
		_w6380_
	);
	LUT2 #(
		.INIT('h2)
	) name5919 (
		\P2_reg0_reg[22]/NET0131 ,
		_w3426_,
		_w6381_
	);
	LUT2 #(
		.INIT('h2)
	) name5920 (
		\P2_reg0_reg[22]/NET0131 ,
		_w2040_,
		_w6382_
	);
	LUT2 #(
		.INIT('h2)
	) name5921 (
		_w2040_,
		_w5753_,
		_w6383_
	);
	LUT2 #(
		.INIT('h1)
	) name5922 (
		_w6382_,
		_w6383_,
		_w6384_
	);
	LUT2 #(
		.INIT('h1)
	) name5923 (
		_w3177_,
		_w6384_,
		_w6385_
	);
	LUT2 #(
		.INIT('h8)
	) name5924 (
		_w2040_,
		_w5760_,
		_w6386_
	);
	LUT2 #(
		.INIT('h1)
	) name5925 (
		_w6382_,
		_w6386_,
		_w6387_
	);
	LUT2 #(
		.INIT('h1)
	) name5926 (
		_w3320_,
		_w6387_,
		_w6388_
	);
	LUT2 #(
		.INIT('h1)
	) name5927 (
		_w6380_,
		_w6381_,
		_w6389_
	);
	LUT2 #(
		.INIT('h4)
	) name5928 (
		_w6385_,
		_w6389_,
		_w6390_
	);
	LUT2 #(
		.INIT('h4)
	) name5929 (
		_w6388_,
		_w6390_,
		_w6391_
	);
	LUT2 #(
		.INIT('h2)
	) name5930 (
		_w2026_,
		_w6391_,
		_w6392_
	);
	LUT2 #(
		.INIT('h1)
	) name5931 (
		_w6374_,
		_w6392_,
		_w6393_
	);
	LUT2 #(
		.INIT('h2)
	) name5932 (
		\P1_state_reg[0]/NET0131 ,
		_w6393_,
		_w6394_
	);
	LUT2 #(
		.INIT('h1)
	) name5933 (
		_w6373_,
		_w6394_,
		_w6395_
	);
	LUT2 #(
		.INIT('h2)
	) name5934 (
		\P1_reg2_reg[18]/NET0131 ,
		_w3435_,
		_w6396_
	);
	LUT2 #(
		.INIT('h8)
	) name5935 (
		\P1_reg2_reg[18]/NET0131 ,
		_w3448_,
		_w6397_
	);
	LUT2 #(
		.INIT('h2)
	) name5936 (
		\P1_reg2_reg[18]/NET0131 ,
		_w3718_,
		_w6398_
	);
	LUT2 #(
		.INIT('h2)
	) name5937 (
		\P1_reg2_reg[18]/NET0131 ,
		_w3466_,
		_w6399_
	);
	LUT2 #(
		.INIT('h8)
	) name5938 (
		_w3466_,
		_w5482_,
		_w6400_
	);
	LUT2 #(
		.INIT('h1)
	) name5939 (
		_w6399_,
		_w6400_,
		_w6401_
	);
	LUT2 #(
		.INIT('h2)
	) name5940 (
		_w3712_,
		_w6401_,
		_w6402_
	);
	LUT2 #(
		.INIT('h2)
	) name5941 (
		_w3466_,
		_w5504_,
		_w6403_
	);
	LUT2 #(
		.INIT('h1)
	) name5942 (
		_w6399_,
		_w6403_,
		_w6404_
	);
	LUT2 #(
		.INIT('h1)
	) name5943 (
		_w3677_,
		_w6404_,
		_w6405_
	);
	LUT2 #(
		.INIT('h8)
	) name5944 (
		_w3466_,
		_w5527_,
		_w6406_
	);
	LUT2 #(
		.INIT('h1)
	) name5945 (
		_w6399_,
		_w6406_,
		_w6407_
	);
	LUT2 #(
		.INIT('h1)
	) name5946 (
		_w3563_,
		_w6407_,
		_w6408_
	);
	LUT2 #(
		.INIT('h2)
	) name5947 (
		_w3466_,
		_w5536_,
		_w6409_
	);
	LUT2 #(
		.INIT('h1)
	) name5948 (
		_w6399_,
		_w6409_,
		_w6410_
	);
	LUT2 #(
		.INIT('h2)
	) name5949 (
		_w1936_,
		_w6410_,
		_w6411_
	);
	LUT2 #(
		.INIT('h8)
	) name5950 (
		_w1399_,
		_w1763_,
		_w6412_
	);
	LUT2 #(
		.INIT('h8)
	) name5951 (
		_w1394_,
		_w1880_,
		_w6413_
	);
	LUT2 #(
		.INIT('h8)
	) name5952 (
		_w3466_,
		_w6413_,
		_w6414_
	);
	LUT2 #(
		.INIT('h1)
	) name5953 (
		_w6398_,
		_w6412_,
		_w6415_
	);
	LUT2 #(
		.INIT('h4)
	) name5954 (
		_w6414_,
		_w6415_,
		_w6416_
	);
	LUT2 #(
		.INIT('h4)
	) name5955 (
		_w6402_,
		_w6416_,
		_w6417_
	);
	LUT2 #(
		.INIT('h1)
	) name5956 (
		_w6405_,
		_w6408_,
		_w6418_
	);
	LUT2 #(
		.INIT('h4)
	) name5957 (
		_w6411_,
		_w6418_,
		_w6419_
	);
	LUT2 #(
		.INIT('h8)
	) name5958 (
		_w6417_,
		_w6419_,
		_w6420_
	);
	LUT2 #(
		.INIT('h2)
	) name5959 (
		_w3450_,
		_w6420_,
		_w6421_
	);
	LUT2 #(
		.INIT('h1)
	) name5960 (
		_w6397_,
		_w6421_,
		_w6422_
	);
	LUT2 #(
		.INIT('h2)
	) name5961 (
		\P1_state_reg[0]/NET0131 ,
		_w6422_,
		_w6423_
	);
	LUT2 #(
		.INIT('h1)
	) name5962 (
		_w6396_,
		_w6423_,
		_w6424_
	);
	LUT2 #(
		.INIT('h2)
	) name5963 (
		\P1_reg2_reg[17]/NET0131 ,
		_w3435_,
		_w6425_
	);
	LUT2 #(
		.INIT('h8)
	) name5964 (
		\P1_reg2_reg[17]/NET0131 ,
		_w3448_,
		_w6426_
	);
	LUT2 #(
		.INIT('h2)
	) name5965 (
		\P1_reg2_reg[17]/NET0131 ,
		_w3466_,
		_w6427_
	);
	LUT2 #(
		.INIT('h2)
	) name5966 (
		_w3466_,
		_w5453_,
		_w6428_
	);
	LUT2 #(
		.INIT('h1)
	) name5967 (
		_w6427_,
		_w6428_,
		_w6429_
	);
	LUT2 #(
		.INIT('h1)
	) name5968 (
		_w3563_,
		_w6429_,
		_w6430_
	);
	LUT2 #(
		.INIT('h8)
	) name5969 (
		_w3466_,
		_w5445_,
		_w6431_
	);
	LUT2 #(
		.INIT('h1)
	) name5970 (
		_w6427_,
		_w6431_,
		_w6432_
	);
	LUT2 #(
		.INIT('h2)
	) name5971 (
		_w3712_,
		_w6432_,
		_w6433_
	);
	LUT2 #(
		.INIT('h8)
	) name5972 (
		_w3466_,
		_w5436_,
		_w6434_
	);
	LUT2 #(
		.INIT('h1)
	) name5973 (
		_w6427_,
		_w6434_,
		_w6435_
	);
	LUT2 #(
		.INIT('h1)
	) name5974 (
		_w3677_,
		_w6435_,
		_w6436_
	);
	LUT2 #(
		.INIT('h8)
	) name5975 (
		_w3466_,
		_w5462_,
		_w6437_
	);
	LUT2 #(
		.INIT('h1)
	) name5976 (
		_w6427_,
		_w6437_,
		_w6438_
	);
	LUT2 #(
		.INIT('h2)
	) name5977 (
		_w1936_,
		_w6438_,
		_w6439_
	);
	LUT2 #(
		.INIT('h2)
	) name5978 (
		\P1_reg2_reg[17]/NET0131 ,
		_w3718_,
		_w6440_
	);
	LUT2 #(
		.INIT('h8)
	) name5979 (
		_w1447_,
		_w1763_,
		_w6441_
	);
	LUT2 #(
		.INIT('h8)
	) name5980 (
		_w1443_,
		_w1880_,
		_w6442_
	);
	LUT2 #(
		.INIT('h8)
	) name5981 (
		_w3466_,
		_w6442_,
		_w6443_
	);
	LUT2 #(
		.INIT('h1)
	) name5982 (
		_w6440_,
		_w6441_,
		_w6444_
	);
	LUT2 #(
		.INIT('h4)
	) name5983 (
		_w6443_,
		_w6444_,
		_w6445_
	);
	LUT2 #(
		.INIT('h4)
	) name5984 (
		_w6433_,
		_w6445_,
		_w6446_
	);
	LUT2 #(
		.INIT('h4)
	) name5985 (
		_w6439_,
		_w6446_,
		_w6447_
	);
	LUT2 #(
		.INIT('h1)
	) name5986 (
		_w6430_,
		_w6436_,
		_w6448_
	);
	LUT2 #(
		.INIT('h8)
	) name5987 (
		_w6447_,
		_w6448_,
		_w6449_
	);
	LUT2 #(
		.INIT('h2)
	) name5988 (
		_w3450_,
		_w6449_,
		_w6450_
	);
	LUT2 #(
		.INIT('h1)
	) name5989 (
		_w6426_,
		_w6450_,
		_w6451_
	);
	LUT2 #(
		.INIT('h2)
	) name5990 (
		\P1_state_reg[0]/NET0131 ,
		_w6451_,
		_w6452_
	);
	LUT2 #(
		.INIT('h1)
	) name5991 (
		_w6425_,
		_w6452_,
		_w6453_
	);
	LUT2 #(
		.INIT('h8)
	) name5992 (
		\P1_reg2_reg[19]/NET0131 ,
		_w3448_,
		_w6454_
	);
	LUT2 #(
		.INIT('h2)
	) name5993 (
		\P1_reg2_reg[19]/NET0131 ,
		_w3466_,
		_w6455_
	);
	LUT2 #(
		.INIT('h2)
	) name5994 (
		_w3466_,
		_w5654_,
		_w6456_
	);
	LUT2 #(
		.INIT('h1)
	) name5995 (
		_w6455_,
		_w6456_,
		_w6457_
	);
	LUT2 #(
		.INIT('h2)
	) name5996 (
		_w1936_,
		_w6457_,
		_w6458_
	);
	LUT2 #(
		.INIT('h8)
	) name5997 (
		_w1423_,
		_w1763_,
		_w6459_
	);
	LUT2 #(
		.INIT('h8)
	) name5998 (
		_w3466_,
		_w5661_,
		_w6460_
	);
	LUT2 #(
		.INIT('h1)
	) name5999 (
		_w6455_,
		_w6460_,
		_w6461_
	);
	LUT2 #(
		.INIT('h1)
	) name6000 (
		_w3563_,
		_w6461_,
		_w6462_
	);
	LUT2 #(
		.INIT('h2)
	) name6001 (
		_w3466_,
		_w5667_,
		_w6463_
	);
	LUT2 #(
		.INIT('h1)
	) name6002 (
		_w6455_,
		_w6463_,
		_w6464_
	);
	LUT2 #(
		.INIT('h1)
	) name6003 (
		_w3677_,
		_w6464_,
		_w6465_
	);
	LUT2 #(
		.INIT('h8)
	) name6004 (
		_w3466_,
		_w5673_,
		_w6466_
	);
	LUT2 #(
		.INIT('h1)
	) name6005 (
		_w6455_,
		_w6466_,
		_w6467_
	);
	LUT2 #(
		.INIT('h2)
	) name6006 (
		_w3712_,
		_w6467_,
		_w6468_
	);
	LUT2 #(
		.INIT('h8)
	) name6007 (
		_w1418_,
		_w3466_,
		_w6469_
	);
	LUT2 #(
		.INIT('h1)
	) name6008 (
		_w6455_,
		_w6469_,
		_w6470_
	);
	LUT2 #(
		.INIT('h2)
	) name6009 (
		_w1880_,
		_w6470_,
		_w6471_
	);
	LUT2 #(
		.INIT('h8)
	) name6010 (
		\P1_reg2_reg[19]/NET0131 ,
		_w3716_,
		_w6472_
	);
	LUT2 #(
		.INIT('h1)
	) name6011 (
		_w6459_,
		_w6472_,
		_w6473_
	);
	LUT2 #(
		.INIT('h4)
	) name6012 (
		_w6471_,
		_w6473_,
		_w6474_
	);
	LUT2 #(
		.INIT('h4)
	) name6013 (
		_w6468_,
		_w6474_,
		_w6475_
	);
	LUT2 #(
		.INIT('h4)
	) name6014 (
		_w6462_,
		_w6475_,
		_w6476_
	);
	LUT2 #(
		.INIT('h4)
	) name6015 (
		_w6465_,
		_w6476_,
		_w6477_
	);
	LUT2 #(
		.INIT('h4)
	) name6016 (
		_w6458_,
		_w6477_,
		_w6478_
	);
	LUT2 #(
		.INIT('h2)
	) name6017 (
		_w3450_,
		_w6478_,
		_w6479_
	);
	LUT2 #(
		.INIT('h1)
	) name6018 (
		_w6454_,
		_w6479_,
		_w6480_
	);
	LUT2 #(
		.INIT('h2)
	) name6019 (
		\P1_state_reg[0]/NET0131 ,
		_w6480_,
		_w6481_
	);
	LUT2 #(
		.INIT('h2)
	) name6020 (
		\P1_reg2_reg[19]/NET0131 ,
		_w3435_,
		_w6482_
	);
	LUT2 #(
		.INIT('h1)
	) name6021 (
		_w6481_,
		_w6482_,
		_w6483_
	);
	LUT2 #(
		.INIT('h2)
	) name6022 (
		\P1_reg2_reg[20]/NET0131 ,
		_w3435_,
		_w6484_
	);
	LUT2 #(
		.INIT('h8)
	) name6023 (
		\P1_reg2_reg[20]/NET0131 ,
		_w3448_,
		_w6485_
	);
	LUT2 #(
		.INIT('h2)
	) name6024 (
		\P1_reg2_reg[20]/NET0131 ,
		_w3466_,
		_w6486_
	);
	LUT2 #(
		.INIT('h2)
	) name6025 (
		_w1356_,
		_w5649_,
		_w6487_
	);
	LUT2 #(
		.INIT('h8)
	) name6026 (
		_w3589_,
		_w5195_,
		_w6488_
	);
	LUT2 #(
		.INIT('h1)
	) name6027 (
		_w6487_,
		_w6488_,
		_w6489_
	);
	LUT2 #(
		.INIT('h1)
	) name6028 (
		_w537_,
		_w6489_,
		_w6490_
	);
	LUT2 #(
		.INIT('h8)
	) name6029 (
		_w537_,
		_w1427_,
		_w6491_
	);
	LUT2 #(
		.INIT('h1)
	) name6030 (
		_w6490_,
		_w6491_,
		_w6492_
	);
	LUT2 #(
		.INIT('h8)
	) name6031 (
		_w3466_,
		_w6492_,
		_w6493_
	);
	LUT2 #(
		.INIT('h1)
	) name6032 (
		_w6486_,
		_w6493_,
		_w6494_
	);
	LUT2 #(
		.INIT('h2)
	) name6033 (
		_w1936_,
		_w6494_,
		_w6495_
	);
	LUT2 #(
		.INIT('h2)
	) name6034 (
		\P1_reg2_reg[20]/NET0131 ,
		_w3718_,
		_w6496_
	);
	LUT2 #(
		.INIT('h2)
	) name6035 (
		_w1828_,
		_w4093_,
		_w6497_
	);
	LUT2 #(
		.INIT('h4)
	) name6036 (
		_w1828_,
		_w4093_,
		_w6498_
	);
	LUT2 #(
		.INIT('h1)
	) name6037 (
		_w6497_,
		_w6498_,
		_w6499_
	);
	LUT2 #(
		.INIT('h2)
	) name6038 (
		_w3466_,
		_w6499_,
		_w6500_
	);
	LUT2 #(
		.INIT('h1)
	) name6039 (
		_w6486_,
		_w6500_,
		_w6501_
	);
	LUT2 #(
		.INIT('h1)
	) name6040 (
		_w3677_,
		_w6501_,
		_w6502_
	);
	LUT2 #(
		.INIT('h8)
	) name6041 (
		_w1828_,
		_w4030_,
		_w6503_
	);
	LUT2 #(
		.INIT('h1)
	) name6042 (
		_w1828_,
		_w4030_,
		_w6504_
	);
	LUT2 #(
		.INIT('h1)
	) name6043 (
		_w6503_,
		_w6504_,
		_w6505_
	);
	LUT2 #(
		.INIT('h2)
	) name6044 (
		_w3466_,
		_w6505_,
		_w6506_
	);
	LUT2 #(
		.INIT('h1)
	) name6045 (
		_w6486_,
		_w6506_,
		_w6507_
	);
	LUT2 #(
		.INIT('h1)
	) name6046 (
		_w3563_,
		_w6507_,
		_w6508_
	);
	LUT2 #(
		.INIT('h2)
	) name6047 (
		_w1365_,
		_w5671_,
		_w6509_
	);
	LUT2 #(
		.INIT('h1)
	) name6048 (
		_w3698_,
		_w6509_,
		_w6510_
	);
	LUT2 #(
		.INIT('h8)
	) name6049 (
		_w3466_,
		_w6510_,
		_w6511_
	);
	LUT2 #(
		.INIT('h1)
	) name6050 (
		_w6486_,
		_w6511_,
		_w6512_
	);
	LUT2 #(
		.INIT('h2)
	) name6051 (
		_w3712_,
		_w6512_,
		_w6513_
	);
	LUT2 #(
		.INIT('h8)
	) name6052 (
		_w1370_,
		_w1763_,
		_w6514_
	);
	LUT2 #(
		.INIT('h8)
	) name6053 (
		_w1365_,
		_w1880_,
		_w6515_
	);
	LUT2 #(
		.INIT('h8)
	) name6054 (
		_w3466_,
		_w6515_,
		_w6516_
	);
	LUT2 #(
		.INIT('h1)
	) name6055 (
		_w6496_,
		_w6514_,
		_w6517_
	);
	LUT2 #(
		.INIT('h4)
	) name6056 (
		_w6516_,
		_w6517_,
		_w6518_
	);
	LUT2 #(
		.INIT('h4)
	) name6057 (
		_w6513_,
		_w6518_,
		_w6519_
	);
	LUT2 #(
		.INIT('h4)
	) name6058 (
		_w6502_,
		_w6519_,
		_w6520_
	);
	LUT2 #(
		.INIT('h4)
	) name6059 (
		_w6508_,
		_w6520_,
		_w6521_
	);
	LUT2 #(
		.INIT('h4)
	) name6060 (
		_w6495_,
		_w6521_,
		_w6522_
	);
	LUT2 #(
		.INIT('h2)
	) name6061 (
		_w3450_,
		_w6522_,
		_w6523_
	);
	LUT2 #(
		.INIT('h1)
	) name6062 (
		_w6485_,
		_w6523_,
		_w6524_
	);
	LUT2 #(
		.INIT('h2)
	) name6063 (
		\P1_state_reg[0]/NET0131 ,
		_w6524_,
		_w6525_
	);
	LUT2 #(
		.INIT('h1)
	) name6064 (
		_w6484_,
		_w6525_,
		_w6526_
	);
	LUT2 #(
		.INIT('h2)
	) name6065 (
		\P2_reg1_reg[17]/NET0131 ,
		_w1983_,
		_w6527_
	);
	LUT2 #(
		.INIT('h8)
	) name6066 (
		\P2_reg1_reg[17]/NET0131 ,
		_w2024_,
		_w6528_
	);
	LUT2 #(
		.INIT('h8)
	) name6067 (
		_w2399_,
		_w3358_,
		_w6529_
	);
	LUT2 #(
		.INIT('h8)
	) name6068 (
		_w3733_,
		_w6529_,
		_w6530_
	);
	LUT2 #(
		.INIT('h2)
	) name6069 (
		\P2_reg1_reg[17]/NET0131 ,
		_w3733_,
		_w6531_
	);
	LUT2 #(
		.INIT('h8)
	) name6070 (
		_w3733_,
		_w5558_,
		_w6532_
	);
	LUT2 #(
		.INIT('h1)
	) name6071 (
		_w6531_,
		_w6532_,
		_w6533_
	);
	LUT2 #(
		.INIT('h1)
	) name6072 (
		_w3177_,
		_w6533_,
		_w6534_
	);
	LUT2 #(
		.INIT('h2)
	) name6073 (
		_w3733_,
		_w5570_,
		_w6535_
	);
	LUT2 #(
		.INIT('h1)
	) name6074 (
		_w6531_,
		_w6535_,
		_w6536_
	);
	LUT2 #(
		.INIT('h2)
	) name6075 (
		_w3411_,
		_w6536_,
		_w6537_
	);
	LUT2 #(
		.INIT('h8)
	) name6076 (
		_w3733_,
		_w5578_,
		_w6538_
	);
	LUT2 #(
		.INIT('h1)
	) name6077 (
		_w6531_,
		_w6538_,
		_w6539_
	);
	LUT2 #(
		.INIT('h2)
	) name6078 (
		_w3355_,
		_w6539_,
		_w6540_
	);
	LUT2 #(
		.INIT('h8)
	) name6079 (
		_w3733_,
		_w5586_,
		_w6541_
	);
	LUT2 #(
		.INIT('h1)
	) name6080 (
		_w6531_,
		_w6541_,
		_w6542_
	);
	LUT2 #(
		.INIT('h1)
	) name6081 (
		_w3320_,
		_w6542_,
		_w6543_
	);
	LUT2 #(
		.INIT('h2)
	) name6082 (
		\P2_reg1_reg[17]/NET0131 ,
		_w3743_,
		_w6544_
	);
	LUT2 #(
		.INIT('h1)
	) name6083 (
		_w6530_,
		_w6544_,
		_w6545_
	);
	LUT2 #(
		.INIT('h4)
	) name6084 (
		_w6543_,
		_w6545_,
		_w6546_
	);
	LUT2 #(
		.INIT('h4)
	) name6085 (
		_w6534_,
		_w6546_,
		_w6547_
	);
	LUT2 #(
		.INIT('h1)
	) name6086 (
		_w6537_,
		_w6540_,
		_w6548_
	);
	LUT2 #(
		.INIT('h8)
	) name6087 (
		_w6547_,
		_w6548_,
		_w6549_
	);
	LUT2 #(
		.INIT('h2)
	) name6088 (
		_w2026_,
		_w6549_,
		_w6550_
	);
	LUT2 #(
		.INIT('h1)
	) name6089 (
		_w6528_,
		_w6550_,
		_w6551_
	);
	LUT2 #(
		.INIT('h2)
	) name6090 (
		\P1_state_reg[0]/NET0131 ,
		_w6551_,
		_w6552_
	);
	LUT2 #(
		.INIT('h1)
	) name6091 (
		_w6527_,
		_w6552_,
		_w6553_
	);
	LUT2 #(
		.INIT('h2)
	) name6092 (
		\P1_reg2_reg[22]/NET0131 ,
		_w3435_,
		_w6554_
	);
	LUT2 #(
		.INIT('h8)
	) name6093 (
		\P1_reg2_reg[22]/NET0131 ,
		_w3448_,
		_w6555_
	);
	LUT2 #(
		.INIT('h2)
	) name6094 (
		\P1_reg2_reg[22]/NET0131 ,
		_w3466_,
		_w6556_
	);
	LUT2 #(
		.INIT('h8)
	) name6095 (
		_w3466_,
		_w6026_,
		_w6557_
	);
	LUT2 #(
		.INIT('h1)
	) name6096 (
		_w6556_,
		_w6557_,
		_w6558_
	);
	LUT2 #(
		.INIT('h1)
	) name6097 (
		_w3677_,
		_w6558_,
		_w6559_
	);
	LUT2 #(
		.INIT('h2)
	) name6098 (
		_w3466_,
		_w6038_,
		_w6560_
	);
	LUT2 #(
		.INIT('h1)
	) name6099 (
		_w6556_,
		_w6560_,
		_w6561_
	);
	LUT2 #(
		.INIT('h1)
	) name6100 (
		_w3563_,
		_w6561_,
		_w6562_
	);
	LUT2 #(
		.INIT('h8)
	) name6101 (
		\P1_reg2_reg[22]/NET0131 ,
		_w3716_,
		_w6563_
	);
	LUT2 #(
		.INIT('h2)
	) name6102 (
		_w3466_,
		_w6048_,
		_w6564_
	);
	LUT2 #(
		.INIT('h1)
	) name6103 (
		_w6556_,
		_w6564_,
		_w6565_
	);
	LUT2 #(
		.INIT('h2)
	) name6104 (
		_w1936_,
		_w6565_,
		_w6566_
	);
	LUT2 #(
		.INIT('h8)
	) name6105 (
		_w3466_,
		_w6054_,
		_w6567_
	);
	LUT2 #(
		.INIT('h1)
	) name6106 (
		_w6556_,
		_w6567_,
		_w6568_
	);
	LUT2 #(
		.INIT('h2)
	) name6107 (
		_w3712_,
		_w6568_,
		_w6569_
	);
	LUT2 #(
		.INIT('h8)
	) name6108 (
		_w1309_,
		_w3466_,
		_w6570_
	);
	LUT2 #(
		.INIT('h1)
	) name6109 (
		_w6556_,
		_w6570_,
		_w6571_
	);
	LUT2 #(
		.INIT('h2)
	) name6110 (
		_w1880_,
		_w6571_,
		_w6572_
	);
	LUT2 #(
		.INIT('h8)
	) name6111 (
		_w1314_,
		_w1763_,
		_w6573_
	);
	LUT2 #(
		.INIT('h1)
	) name6112 (
		_w6563_,
		_w6573_,
		_w6574_
	);
	LUT2 #(
		.INIT('h4)
	) name6113 (
		_w6572_,
		_w6574_,
		_w6575_
	);
	LUT2 #(
		.INIT('h4)
	) name6114 (
		_w6569_,
		_w6575_,
		_w6576_
	);
	LUT2 #(
		.INIT('h4)
	) name6115 (
		_w6566_,
		_w6576_,
		_w6577_
	);
	LUT2 #(
		.INIT('h4)
	) name6116 (
		_w6559_,
		_w6577_,
		_w6578_
	);
	LUT2 #(
		.INIT('h4)
	) name6117 (
		_w6562_,
		_w6578_,
		_w6579_
	);
	LUT2 #(
		.INIT('h2)
	) name6118 (
		_w3450_,
		_w6579_,
		_w6580_
	);
	LUT2 #(
		.INIT('h1)
	) name6119 (
		_w6555_,
		_w6580_,
		_w6581_
	);
	LUT2 #(
		.INIT('h2)
	) name6120 (
		\P1_state_reg[0]/NET0131 ,
		_w6581_,
		_w6582_
	);
	LUT2 #(
		.INIT('h1)
	) name6121 (
		_w6554_,
		_w6582_,
		_w6583_
	);
	LUT2 #(
		.INIT('h2)
	) name6122 (
		\P2_reg1_reg[18]/NET0131 ,
		_w1983_,
		_w6584_
	);
	LUT2 #(
		.INIT('h8)
	) name6123 (
		\P2_reg1_reg[18]/NET0131 ,
		_w2024_,
		_w6585_
	);
	LUT2 #(
		.INIT('h2)
	) name6124 (
		\P2_reg1_reg[18]/NET0131 ,
		_w3743_,
		_w6586_
	);
	LUT2 #(
		.INIT('h2)
	) name6125 (
		\P2_reg1_reg[18]/NET0131 ,
		_w3733_,
		_w6587_
	);
	LUT2 #(
		.INIT('h8)
	) name6126 (
		_w3733_,
		_w6331_,
		_w6588_
	);
	LUT2 #(
		.INIT('h1)
	) name6127 (
		_w6587_,
		_w6588_,
		_w6589_
	);
	LUT2 #(
		.INIT('h2)
	) name6128 (
		_w3355_,
		_w6589_,
		_w6590_
	);
	LUT2 #(
		.INIT('h8)
	) name6129 (
		_w3733_,
		_w6337_,
		_w6591_
	);
	LUT2 #(
		.INIT('h1)
	) name6130 (
		_w6587_,
		_w6591_,
		_w6592_
	);
	LUT2 #(
		.INIT('h1)
	) name6131 (
		_w3177_,
		_w6592_,
		_w6593_
	);
	LUT2 #(
		.INIT('h2)
	) name6132 (
		_w3733_,
		_w6343_,
		_w6594_
	);
	LUT2 #(
		.INIT('h1)
	) name6133 (
		_w6587_,
		_w6594_,
		_w6595_
	);
	LUT2 #(
		.INIT('h1)
	) name6134 (
		_w3320_,
		_w6595_,
		_w6596_
	);
	LUT2 #(
		.INIT('h8)
	) name6135 (
		_w3733_,
		_w6351_,
		_w6597_
	);
	LUT2 #(
		.INIT('h1)
	) name6136 (
		_w6587_,
		_w6597_,
		_w6598_
	);
	LUT2 #(
		.INIT('h2)
	) name6137 (
		_w3411_,
		_w6598_,
		_w6599_
	);
	LUT2 #(
		.INIT('h8)
	) name6138 (
		_w3733_,
		_w6356_,
		_w6600_
	);
	LUT2 #(
		.INIT('h1)
	) name6139 (
		_w6586_,
		_w6600_,
		_w6601_
	);
	LUT2 #(
		.INIT('h4)
	) name6140 (
		_w6599_,
		_w6601_,
		_w6602_
	);
	LUT2 #(
		.INIT('h4)
	) name6141 (
		_w6593_,
		_w6602_,
		_w6603_
	);
	LUT2 #(
		.INIT('h4)
	) name6142 (
		_w6596_,
		_w6603_,
		_w6604_
	);
	LUT2 #(
		.INIT('h4)
	) name6143 (
		_w6590_,
		_w6604_,
		_w6605_
	);
	LUT2 #(
		.INIT('h2)
	) name6144 (
		_w2026_,
		_w6605_,
		_w6606_
	);
	LUT2 #(
		.INIT('h1)
	) name6145 (
		_w6585_,
		_w6606_,
		_w6607_
	);
	LUT2 #(
		.INIT('h2)
	) name6146 (
		\P1_state_reg[0]/NET0131 ,
		_w6607_,
		_w6608_
	);
	LUT2 #(
		.INIT('h1)
	) name6147 (
		_w6584_,
		_w6608_,
		_w6609_
	);
	LUT2 #(
		.INIT('h2)
	) name6148 (
		\P2_reg1_reg[19]/NET0131 ,
		_w1983_,
		_w6610_
	);
	LUT2 #(
		.INIT('h8)
	) name6149 (
		\P2_reg1_reg[19]/NET0131 ,
		_w2024_,
		_w6611_
	);
	LUT2 #(
		.INIT('h2)
	) name6150 (
		\P2_reg1_reg[19]/NET0131 ,
		_w3743_,
		_w6612_
	);
	LUT2 #(
		.INIT('h2)
	) name6151 (
		\P2_reg1_reg[19]/NET0131 ,
		_w3733_,
		_w6613_
	);
	LUT2 #(
		.INIT('h8)
	) name6152 (
		_w3733_,
		_w5608_,
		_w6614_
	);
	LUT2 #(
		.INIT('h1)
	) name6153 (
		_w6613_,
		_w6614_,
		_w6615_
	);
	LUT2 #(
		.INIT('h1)
	) name6154 (
		_w3177_,
		_w6615_,
		_w6616_
	);
	LUT2 #(
		.INIT('h2)
	) name6155 (
		_w3733_,
		_w5614_,
		_w6617_
	);
	LUT2 #(
		.INIT('h1)
	) name6156 (
		_w6613_,
		_w6617_,
		_w6618_
	);
	LUT2 #(
		.INIT('h1)
	) name6157 (
		_w3320_,
		_w6618_,
		_w6619_
	);
	LUT2 #(
		.INIT('h8)
	) name6158 (
		_w3733_,
		_w5624_,
		_w6620_
	);
	LUT2 #(
		.INIT('h1)
	) name6159 (
		_w6613_,
		_w6620_,
		_w6621_
	);
	LUT2 #(
		.INIT('h2)
	) name6160 (
		_w3411_,
		_w6621_,
		_w6622_
	);
	LUT2 #(
		.INIT('h8)
	) name6161 (
		_w3733_,
		_w5630_,
		_w6623_
	);
	LUT2 #(
		.INIT('h1)
	) name6162 (
		_w6613_,
		_w6623_,
		_w6624_
	);
	LUT2 #(
		.INIT('h2)
	) name6163 (
		_w3355_,
		_w6624_,
		_w6625_
	);
	LUT2 #(
		.INIT('h8)
	) name6164 (
		_w2299_,
		_w3358_,
		_w6626_
	);
	LUT2 #(
		.INIT('h8)
	) name6165 (
		_w3733_,
		_w6626_,
		_w6627_
	);
	LUT2 #(
		.INIT('h1)
	) name6166 (
		_w6612_,
		_w6627_,
		_w6628_
	);
	LUT2 #(
		.INIT('h4)
	) name6167 (
		_w6619_,
		_w6628_,
		_w6629_
	);
	LUT2 #(
		.INIT('h4)
	) name6168 (
		_w6625_,
		_w6629_,
		_w6630_
	);
	LUT2 #(
		.INIT('h4)
	) name6169 (
		_w6622_,
		_w6630_,
		_w6631_
	);
	LUT2 #(
		.INIT('h4)
	) name6170 (
		_w6616_,
		_w6631_,
		_w6632_
	);
	LUT2 #(
		.INIT('h2)
	) name6171 (
		_w2026_,
		_w6632_,
		_w6633_
	);
	LUT2 #(
		.INIT('h1)
	) name6172 (
		_w6611_,
		_w6633_,
		_w6634_
	);
	LUT2 #(
		.INIT('h2)
	) name6173 (
		\P1_state_reg[0]/NET0131 ,
		_w6634_,
		_w6635_
	);
	LUT2 #(
		.INIT('h1)
	) name6174 (
		_w6610_,
		_w6635_,
		_w6636_
	);
	LUT2 #(
		.INIT('h2)
	) name6175 (
		\P2_reg1_reg[21]/NET0131 ,
		_w1983_,
		_w6637_
	);
	LUT2 #(
		.INIT('h8)
	) name6176 (
		\P2_reg1_reg[21]/NET0131 ,
		_w2024_,
		_w6638_
	);
	LUT2 #(
		.INIT('h2)
	) name6177 (
		_w3320_,
		_w3358_,
		_w6639_
	);
	LUT2 #(
		.INIT('h2)
	) name6178 (
		_w3177_,
		_w3745_,
		_w6640_
	);
	LUT2 #(
		.INIT('h8)
	) name6179 (
		_w6639_,
		_w6640_,
		_w6641_
	);
	LUT2 #(
		.INIT('h1)
	) name6180 (
		_w3733_,
		_w6641_,
		_w6642_
	);
	LUT2 #(
		.INIT('h2)
	) name6181 (
		_w3421_,
		_w6642_,
		_w6643_
	);
	LUT2 #(
		.INIT('h2)
	) name6182 (
		\P2_reg1_reg[21]/NET0131 ,
		_w6643_,
		_w6644_
	);
	LUT2 #(
		.INIT('h8)
	) name6183 (
		_w3121_,
		_w3358_,
		_w6645_
	);
	LUT2 #(
		.INIT('h1)
	) name6184 (
		_w3177_,
		_w6290_,
		_w6646_
	);
	LUT2 #(
		.INIT('h2)
	) name6185 (
		_w6309_,
		_w6645_,
		_w6647_
	);
	LUT2 #(
		.INIT('h4)
	) name6186 (
		_w6646_,
		_w6647_,
		_w6648_
	);
	LUT2 #(
		.INIT('h2)
	) name6187 (
		_w3733_,
		_w6648_,
		_w6649_
	);
	LUT2 #(
		.INIT('h1)
	) name6188 (
		_w6644_,
		_w6649_,
		_w6650_
	);
	LUT2 #(
		.INIT('h2)
	) name6189 (
		_w2026_,
		_w6650_,
		_w6651_
	);
	LUT2 #(
		.INIT('h1)
	) name6190 (
		_w6638_,
		_w6651_,
		_w6652_
	);
	LUT2 #(
		.INIT('h2)
	) name6191 (
		\P1_state_reg[0]/NET0131 ,
		_w6652_,
		_w6653_
	);
	LUT2 #(
		.INIT('h1)
	) name6192 (
		_w6637_,
		_w6653_,
		_w6654_
	);
	LUT2 #(
		.INIT('h2)
	) name6193 (
		\P2_reg1_reg[22]/NET0131 ,
		_w1983_,
		_w6655_
	);
	LUT2 #(
		.INIT('h8)
	) name6194 (
		\P2_reg1_reg[22]/NET0131 ,
		_w2024_,
		_w6656_
	);
	LUT2 #(
		.INIT('h2)
	) name6195 (
		_w3733_,
		_w6379_,
		_w6657_
	);
	LUT2 #(
		.INIT('h2)
	) name6196 (
		\P2_reg1_reg[22]/NET0131 ,
		_w3747_,
		_w6658_
	);
	LUT2 #(
		.INIT('h2)
	) name6197 (
		\P2_reg1_reg[22]/NET0131 ,
		_w3733_,
		_w6659_
	);
	LUT2 #(
		.INIT('h2)
	) name6198 (
		_w3733_,
		_w5753_,
		_w6660_
	);
	LUT2 #(
		.INIT('h1)
	) name6199 (
		_w6659_,
		_w6660_,
		_w6661_
	);
	LUT2 #(
		.INIT('h1)
	) name6200 (
		_w3177_,
		_w6661_,
		_w6662_
	);
	LUT2 #(
		.INIT('h8)
	) name6201 (
		_w3733_,
		_w5760_,
		_w6663_
	);
	LUT2 #(
		.INIT('h1)
	) name6202 (
		_w6659_,
		_w6663_,
		_w6664_
	);
	LUT2 #(
		.INIT('h1)
	) name6203 (
		_w3320_,
		_w6664_,
		_w6665_
	);
	LUT2 #(
		.INIT('h1)
	) name6204 (
		_w6657_,
		_w6658_,
		_w6666_
	);
	LUT2 #(
		.INIT('h4)
	) name6205 (
		_w6662_,
		_w6666_,
		_w6667_
	);
	LUT2 #(
		.INIT('h4)
	) name6206 (
		_w6665_,
		_w6667_,
		_w6668_
	);
	LUT2 #(
		.INIT('h2)
	) name6207 (
		_w2026_,
		_w6668_,
		_w6669_
	);
	LUT2 #(
		.INIT('h1)
	) name6208 (
		_w6656_,
		_w6669_,
		_w6670_
	);
	LUT2 #(
		.INIT('h2)
	) name6209 (
		\P1_state_reg[0]/NET0131 ,
		_w6670_,
		_w6671_
	);
	LUT2 #(
		.INIT('h1)
	) name6210 (
		_w6655_,
		_w6671_,
		_w6672_
	);
	LUT2 #(
		.INIT('h2)
	) name6211 (
		\P2_reg2_reg[17]/NET0131 ,
		_w1983_,
		_w6673_
	);
	LUT2 #(
		.INIT('h8)
	) name6212 (
		\P2_reg2_reg[17]/NET0131 ,
		_w2024_,
		_w6674_
	);
	LUT2 #(
		.INIT('h2)
	) name6213 (
		\P2_reg2_reg[17]/NET0131 ,
		_w3774_,
		_w6675_
	);
	LUT2 #(
		.INIT('h2)
	) name6214 (
		\P2_reg2_reg[17]/NET0131 ,
		_w3758_,
		_w6676_
	);
	LUT2 #(
		.INIT('h8)
	) name6215 (
		_w3758_,
		_w5558_,
		_w6677_
	);
	LUT2 #(
		.INIT('h1)
	) name6216 (
		_w6676_,
		_w6677_,
		_w6678_
	);
	LUT2 #(
		.INIT('h1)
	) name6217 (
		_w3177_,
		_w6678_,
		_w6679_
	);
	LUT2 #(
		.INIT('h2)
	) name6218 (
		_w3758_,
		_w5570_,
		_w6680_
	);
	LUT2 #(
		.INIT('h1)
	) name6219 (
		_w6676_,
		_w6680_,
		_w6681_
	);
	LUT2 #(
		.INIT('h2)
	) name6220 (
		_w3411_,
		_w6681_,
		_w6682_
	);
	LUT2 #(
		.INIT('h8)
	) name6221 (
		_w3758_,
		_w5578_,
		_w6683_
	);
	LUT2 #(
		.INIT('h1)
	) name6222 (
		_w6676_,
		_w6683_,
		_w6684_
	);
	LUT2 #(
		.INIT('h2)
	) name6223 (
		_w3355_,
		_w6684_,
		_w6685_
	);
	LUT2 #(
		.INIT('h8)
	) name6224 (
		_w3758_,
		_w5586_,
		_w6686_
	);
	LUT2 #(
		.INIT('h1)
	) name6225 (
		_w6676_,
		_w6686_,
		_w6687_
	);
	LUT2 #(
		.INIT('h1)
	) name6226 (
		_w3320_,
		_w6687_,
		_w6688_
	);
	LUT2 #(
		.INIT('h8)
	) name6227 (
		_w2373_,
		_w3420_,
		_w6689_
	);
	LUT2 #(
		.INIT('h8)
	) name6228 (
		_w3758_,
		_w6529_,
		_w6690_
	);
	LUT2 #(
		.INIT('h1)
	) name6229 (
		_w6675_,
		_w6689_,
		_w6691_
	);
	LUT2 #(
		.INIT('h4)
	) name6230 (
		_w6690_,
		_w6691_,
		_w6692_
	);
	LUT2 #(
		.INIT('h4)
	) name6231 (
		_w6688_,
		_w6692_,
		_w6693_
	);
	LUT2 #(
		.INIT('h4)
	) name6232 (
		_w6679_,
		_w6693_,
		_w6694_
	);
	LUT2 #(
		.INIT('h1)
	) name6233 (
		_w6682_,
		_w6685_,
		_w6695_
	);
	LUT2 #(
		.INIT('h8)
	) name6234 (
		_w6694_,
		_w6695_,
		_w6696_
	);
	LUT2 #(
		.INIT('h2)
	) name6235 (
		_w2026_,
		_w6696_,
		_w6697_
	);
	LUT2 #(
		.INIT('h1)
	) name6236 (
		_w6674_,
		_w6697_,
		_w6698_
	);
	LUT2 #(
		.INIT('h2)
	) name6237 (
		\P1_state_reg[0]/NET0131 ,
		_w6698_,
		_w6699_
	);
	LUT2 #(
		.INIT('h1)
	) name6238 (
		_w6673_,
		_w6699_,
		_w6700_
	);
	LUT2 #(
		.INIT('h2)
	) name6239 (
		\P2_reg2_reg[19]/NET0131 ,
		_w1983_,
		_w6701_
	);
	LUT2 #(
		.INIT('h8)
	) name6240 (
		\P2_reg2_reg[19]/NET0131 ,
		_w2024_,
		_w6702_
	);
	LUT2 #(
		.INIT('h8)
	) name6241 (
		_w3758_,
		_w6626_,
		_w6703_
	);
	LUT2 #(
		.INIT('h2)
	) name6242 (
		\P2_reg2_reg[19]/NET0131 ,
		_w3758_,
		_w6704_
	);
	LUT2 #(
		.INIT('h8)
	) name6243 (
		_w3758_,
		_w5608_,
		_w6705_
	);
	LUT2 #(
		.INIT('h1)
	) name6244 (
		_w6704_,
		_w6705_,
		_w6706_
	);
	LUT2 #(
		.INIT('h1)
	) name6245 (
		_w3177_,
		_w6706_,
		_w6707_
	);
	LUT2 #(
		.INIT('h2)
	) name6246 (
		_w3758_,
		_w5614_,
		_w6708_
	);
	LUT2 #(
		.INIT('h1)
	) name6247 (
		_w6704_,
		_w6708_,
		_w6709_
	);
	LUT2 #(
		.INIT('h1)
	) name6248 (
		_w3320_,
		_w6709_,
		_w6710_
	);
	LUT2 #(
		.INIT('h8)
	) name6249 (
		_w3758_,
		_w5624_,
		_w6711_
	);
	LUT2 #(
		.INIT('h1)
	) name6250 (
		_w6704_,
		_w6711_,
		_w6712_
	);
	LUT2 #(
		.INIT('h2)
	) name6251 (
		_w3411_,
		_w6712_,
		_w6713_
	);
	LUT2 #(
		.INIT('h8)
	) name6252 (
		_w3758_,
		_w5630_,
		_w6714_
	);
	LUT2 #(
		.INIT('h1)
	) name6253 (
		_w6704_,
		_w6714_,
		_w6715_
	);
	LUT2 #(
		.INIT('h2)
	) name6254 (
		_w3355_,
		_w6715_,
		_w6716_
	);
	LUT2 #(
		.INIT('h8)
	) name6255 (
		_w2307_,
		_w3420_,
		_w6717_
	);
	LUT2 #(
		.INIT('h2)
	) name6256 (
		\P2_reg2_reg[19]/NET0131 ,
		_w3774_,
		_w6718_
	);
	LUT2 #(
		.INIT('h1)
	) name6257 (
		_w6717_,
		_w6718_,
		_w6719_
	);
	LUT2 #(
		.INIT('h4)
	) name6258 (
		_w6703_,
		_w6719_,
		_w6720_
	);
	LUT2 #(
		.INIT('h4)
	) name6259 (
		_w6710_,
		_w6720_,
		_w6721_
	);
	LUT2 #(
		.INIT('h4)
	) name6260 (
		_w6716_,
		_w6721_,
		_w6722_
	);
	LUT2 #(
		.INIT('h4)
	) name6261 (
		_w6713_,
		_w6722_,
		_w6723_
	);
	LUT2 #(
		.INIT('h4)
	) name6262 (
		_w6707_,
		_w6723_,
		_w6724_
	);
	LUT2 #(
		.INIT('h2)
	) name6263 (
		_w2026_,
		_w6724_,
		_w6725_
	);
	LUT2 #(
		.INIT('h1)
	) name6264 (
		_w6702_,
		_w6725_,
		_w6726_
	);
	LUT2 #(
		.INIT('h2)
	) name6265 (
		\P1_state_reg[0]/NET0131 ,
		_w6726_,
		_w6727_
	);
	LUT2 #(
		.INIT('h1)
	) name6266 (
		_w6701_,
		_w6727_,
		_w6728_
	);
	LUT2 #(
		.INIT('h2)
	) name6267 (
		\P2_reg2_reg[20]/NET0131 ,
		_w1983_,
		_w6729_
	);
	LUT2 #(
		.INIT('h8)
	) name6268 (
		\P2_reg2_reg[20]/NET0131 ,
		_w2024_,
		_w6730_
	);
	LUT2 #(
		.INIT('h2)
	) name6269 (
		\P2_reg2_reg[20]/NET0131 ,
		_w3774_,
		_w6731_
	);
	LUT2 #(
		.INIT('h2)
	) name6270 (
		\P2_reg2_reg[20]/NET0131 ,
		_w3758_,
		_w6732_
	);
	LUT2 #(
		.INIT('h2)
	) name6271 (
		_w3130_,
		_w5620_,
		_w6733_
	);
	LUT2 #(
		.INIT('h1)
	) name6272 (
		_w3394_,
		_w6733_,
		_w6734_
	);
	LUT2 #(
		.INIT('h1)
	) name6273 (
		_w2058_,
		_w6734_,
		_w6735_
	);
	LUT2 #(
		.INIT('h8)
	) name6274 (
		_w2058_,
		_w2311_,
		_w6736_
	);
	LUT2 #(
		.INIT('h1)
	) name6275 (
		_w6735_,
		_w6736_,
		_w6737_
	);
	LUT2 #(
		.INIT('h8)
	) name6276 (
		_w3758_,
		_w6737_,
		_w6738_
	);
	LUT2 #(
		.INIT('h1)
	) name6277 (
		_w6732_,
		_w6738_,
		_w6739_
	);
	LUT2 #(
		.INIT('h2)
	) name6278 (
		_w3411_,
		_w6739_,
		_w6740_
	);
	LUT2 #(
		.INIT('h8)
	) name6279 (
		_w3916_,
		_w4217_,
		_w6741_
	);
	LUT2 #(
		.INIT('h1)
	) name6280 (
		_w3916_,
		_w4217_,
		_w6742_
	);
	LUT2 #(
		.INIT('h1)
	) name6281 (
		_w6741_,
		_w6742_,
		_w6743_
	);
	LUT2 #(
		.INIT('h2)
	) name6282 (
		_w3758_,
		_w6743_,
		_w6744_
	);
	LUT2 #(
		.INIT('h1)
	) name6283 (
		_w6732_,
		_w6744_,
		_w6745_
	);
	LUT2 #(
		.INIT('h1)
	) name6284 (
		_w3177_,
		_w6745_,
		_w6746_
	);
	LUT2 #(
		.INIT('h4)
	) name6285 (
		_w3845_,
		_w4217_,
		_w6747_
	);
	LUT2 #(
		.INIT('h2)
	) name6286 (
		_w3845_,
		_w4217_,
		_w6748_
	);
	LUT2 #(
		.INIT('h1)
	) name6287 (
		_w6747_,
		_w6748_,
		_w6749_
	);
	LUT2 #(
		.INIT('h2)
	) name6288 (
		_w3758_,
		_w6749_,
		_w6750_
	);
	LUT2 #(
		.INIT('h1)
	) name6289 (
		_w6732_,
		_w6750_,
		_w6751_
	);
	LUT2 #(
		.INIT('h1)
	) name6290 (
		_w3320_,
		_w6751_,
		_w6752_
	);
	LUT2 #(
		.INIT('h2)
	) name6291 (
		_w2358_,
		_w5629_,
		_w6753_
	);
	LUT2 #(
		.INIT('h1)
	) name6292 (
		_w5765_,
		_w6753_,
		_w6754_
	);
	LUT2 #(
		.INIT('h8)
	) name6293 (
		_w3758_,
		_w6754_,
		_w6755_
	);
	LUT2 #(
		.INIT('h1)
	) name6294 (
		_w6732_,
		_w6755_,
		_w6756_
	);
	LUT2 #(
		.INIT('h2)
	) name6295 (
		_w3355_,
		_w6756_,
		_w6757_
	);
	LUT2 #(
		.INIT('h8)
	) name6296 (
		_w2364_,
		_w3420_,
		_w6758_
	);
	LUT2 #(
		.INIT('h8)
	) name6297 (
		_w2358_,
		_w3358_,
		_w6759_
	);
	LUT2 #(
		.INIT('h8)
	) name6298 (
		_w3758_,
		_w6759_,
		_w6760_
	);
	LUT2 #(
		.INIT('h1)
	) name6299 (
		_w6731_,
		_w6758_,
		_w6761_
	);
	LUT2 #(
		.INIT('h4)
	) name6300 (
		_w6760_,
		_w6761_,
		_w6762_
	);
	LUT2 #(
		.INIT('h4)
	) name6301 (
		_w6746_,
		_w6762_,
		_w6763_
	);
	LUT2 #(
		.INIT('h1)
	) name6302 (
		_w6752_,
		_w6757_,
		_w6764_
	);
	LUT2 #(
		.INIT('h8)
	) name6303 (
		_w6763_,
		_w6764_,
		_w6765_
	);
	LUT2 #(
		.INIT('h4)
	) name6304 (
		_w6740_,
		_w6765_,
		_w6766_
	);
	LUT2 #(
		.INIT('h2)
	) name6305 (
		_w2026_,
		_w6766_,
		_w6767_
	);
	LUT2 #(
		.INIT('h1)
	) name6306 (
		_w6730_,
		_w6767_,
		_w6768_
	);
	LUT2 #(
		.INIT('h2)
	) name6307 (
		\P1_state_reg[0]/NET0131 ,
		_w6768_,
		_w6769_
	);
	LUT2 #(
		.INIT('h1)
	) name6308 (
		_w6729_,
		_w6769_,
		_w6770_
	);
	LUT2 #(
		.INIT('h2)
	) name6309 (
		\P2_reg2_reg[22]/NET0131 ,
		_w1983_,
		_w6771_
	);
	LUT2 #(
		.INIT('h8)
	) name6310 (
		\P2_reg2_reg[22]/NET0131 ,
		_w2024_,
		_w6772_
	);
	LUT2 #(
		.INIT('h2)
	) name6311 (
		_w3758_,
		_w6379_,
		_w6773_
	);
	LUT2 #(
		.INIT('h2)
	) name6312 (
		\P2_reg2_reg[22]/NET0131 ,
		_w4933_,
		_w6774_
	);
	LUT2 #(
		.INIT('h8)
	) name6313 (
		_w3108_,
		_w3420_,
		_w6775_
	);
	LUT2 #(
		.INIT('h2)
	) name6314 (
		\P2_reg2_reg[22]/NET0131 ,
		_w3758_,
		_w6776_
	);
	LUT2 #(
		.INIT('h2)
	) name6315 (
		_w3758_,
		_w5753_,
		_w6777_
	);
	LUT2 #(
		.INIT('h1)
	) name6316 (
		_w6776_,
		_w6777_,
		_w6778_
	);
	LUT2 #(
		.INIT('h1)
	) name6317 (
		_w3177_,
		_w6778_,
		_w6779_
	);
	LUT2 #(
		.INIT('h8)
	) name6318 (
		_w3758_,
		_w5760_,
		_w6780_
	);
	LUT2 #(
		.INIT('h1)
	) name6319 (
		_w6776_,
		_w6780_,
		_w6781_
	);
	LUT2 #(
		.INIT('h1)
	) name6320 (
		_w3320_,
		_w6781_,
		_w6782_
	);
	LUT2 #(
		.INIT('h1)
	) name6321 (
		_w6774_,
		_w6775_,
		_w6783_
	);
	LUT2 #(
		.INIT('h4)
	) name6322 (
		_w6773_,
		_w6783_,
		_w6784_
	);
	LUT2 #(
		.INIT('h4)
	) name6323 (
		_w6779_,
		_w6784_,
		_w6785_
	);
	LUT2 #(
		.INIT('h4)
	) name6324 (
		_w6782_,
		_w6785_,
		_w6786_
	);
	LUT2 #(
		.INIT('h2)
	) name6325 (
		_w2026_,
		_w6786_,
		_w6787_
	);
	LUT2 #(
		.INIT('h1)
	) name6326 (
		_w6772_,
		_w6787_,
		_w6788_
	);
	LUT2 #(
		.INIT('h2)
	) name6327 (
		\P1_state_reg[0]/NET0131 ,
		_w6788_,
		_w6789_
	);
	LUT2 #(
		.INIT('h1)
	) name6328 (
		_w6771_,
		_w6789_,
		_w6790_
	);
	LUT2 #(
		.INIT('h2)
	) name6329 (
		\P1_reg0_reg[17]/NET0131 ,
		_w3435_,
		_w6791_
	);
	LUT2 #(
		.INIT('h8)
	) name6330 (
		\P1_reg0_reg[17]/NET0131 ,
		_w3448_,
		_w6792_
	);
	LUT2 #(
		.INIT('h2)
	) name6331 (
		\P1_reg0_reg[17]/NET0131 ,
		_w4493_,
		_w6793_
	);
	LUT2 #(
		.INIT('h8)
	) name6332 (
		_w4396_,
		_w6442_,
		_w6794_
	);
	LUT2 #(
		.INIT('h2)
	) name6333 (
		\P1_reg0_reg[17]/NET0131 ,
		_w4396_,
		_w6795_
	);
	LUT2 #(
		.INIT('h8)
	) name6334 (
		_w4396_,
		_w5436_,
		_w6796_
	);
	LUT2 #(
		.INIT('h1)
	) name6335 (
		_w6795_,
		_w6796_,
		_w6797_
	);
	LUT2 #(
		.INIT('h1)
	) name6336 (
		_w3677_,
		_w6797_,
		_w6798_
	);
	LUT2 #(
		.INIT('h8)
	) name6337 (
		_w4396_,
		_w5445_,
		_w6799_
	);
	LUT2 #(
		.INIT('h1)
	) name6338 (
		_w6795_,
		_w6799_,
		_w6800_
	);
	LUT2 #(
		.INIT('h2)
	) name6339 (
		_w3712_,
		_w6800_,
		_w6801_
	);
	LUT2 #(
		.INIT('h2)
	) name6340 (
		_w4396_,
		_w5453_,
		_w6802_
	);
	LUT2 #(
		.INIT('h1)
	) name6341 (
		_w6795_,
		_w6802_,
		_w6803_
	);
	LUT2 #(
		.INIT('h1)
	) name6342 (
		_w3563_,
		_w6803_,
		_w6804_
	);
	LUT2 #(
		.INIT('h8)
	) name6343 (
		_w4396_,
		_w5462_,
		_w6805_
	);
	LUT2 #(
		.INIT('h1)
	) name6344 (
		_w6795_,
		_w6805_,
		_w6806_
	);
	LUT2 #(
		.INIT('h2)
	) name6345 (
		_w1936_,
		_w6806_,
		_w6807_
	);
	LUT2 #(
		.INIT('h1)
	) name6346 (
		_w6793_,
		_w6794_,
		_w6808_
	);
	LUT2 #(
		.INIT('h4)
	) name6347 (
		_w6801_,
		_w6808_,
		_w6809_
	);
	LUT2 #(
		.INIT('h4)
	) name6348 (
		_w6807_,
		_w6809_,
		_w6810_
	);
	LUT2 #(
		.INIT('h1)
	) name6349 (
		_w6798_,
		_w6804_,
		_w6811_
	);
	LUT2 #(
		.INIT('h8)
	) name6350 (
		_w6810_,
		_w6811_,
		_w6812_
	);
	LUT2 #(
		.INIT('h2)
	) name6351 (
		_w3450_,
		_w6812_,
		_w6813_
	);
	LUT2 #(
		.INIT('h1)
	) name6352 (
		_w6792_,
		_w6813_,
		_w6814_
	);
	LUT2 #(
		.INIT('h2)
	) name6353 (
		\P1_state_reg[0]/NET0131 ,
		_w6814_,
		_w6815_
	);
	LUT2 #(
		.INIT('h1)
	) name6354 (
		_w6791_,
		_w6815_,
		_w6816_
	);
	LUT2 #(
		.INIT('h2)
	) name6355 (
		\P1_reg0_reg[18]/NET0131 ,
		_w3435_,
		_w6817_
	);
	LUT2 #(
		.INIT('h8)
	) name6356 (
		\P1_reg0_reg[18]/NET0131 ,
		_w3448_,
		_w6818_
	);
	LUT2 #(
		.INIT('h8)
	) name6357 (
		_w4396_,
		_w6413_,
		_w6819_
	);
	LUT2 #(
		.INIT('h2)
	) name6358 (
		\P1_reg0_reg[18]/NET0131 ,
		_w4396_,
		_w6820_
	);
	LUT2 #(
		.INIT('h8)
	) name6359 (
		_w4396_,
		_w5482_,
		_w6821_
	);
	LUT2 #(
		.INIT('h1)
	) name6360 (
		_w6820_,
		_w6821_,
		_w6822_
	);
	LUT2 #(
		.INIT('h2)
	) name6361 (
		_w3712_,
		_w6822_,
		_w6823_
	);
	LUT2 #(
		.INIT('h2)
	) name6362 (
		_w4396_,
		_w5504_,
		_w6824_
	);
	LUT2 #(
		.INIT('h1)
	) name6363 (
		_w6820_,
		_w6824_,
		_w6825_
	);
	LUT2 #(
		.INIT('h1)
	) name6364 (
		_w3677_,
		_w6825_,
		_w6826_
	);
	LUT2 #(
		.INIT('h8)
	) name6365 (
		_w4396_,
		_w5527_,
		_w6827_
	);
	LUT2 #(
		.INIT('h1)
	) name6366 (
		_w6820_,
		_w6827_,
		_w6828_
	);
	LUT2 #(
		.INIT('h1)
	) name6367 (
		_w3563_,
		_w6828_,
		_w6829_
	);
	LUT2 #(
		.INIT('h2)
	) name6368 (
		_w4396_,
		_w5536_,
		_w6830_
	);
	LUT2 #(
		.INIT('h1)
	) name6369 (
		_w6820_,
		_w6830_,
		_w6831_
	);
	LUT2 #(
		.INIT('h2)
	) name6370 (
		_w1936_,
		_w6831_,
		_w6832_
	);
	LUT2 #(
		.INIT('h2)
	) name6371 (
		\P1_reg0_reg[18]/NET0131 ,
		_w4493_,
		_w6833_
	);
	LUT2 #(
		.INIT('h1)
	) name6372 (
		_w6819_,
		_w6833_,
		_w6834_
	);
	LUT2 #(
		.INIT('h4)
	) name6373 (
		_w6823_,
		_w6834_,
		_w6835_
	);
	LUT2 #(
		.INIT('h1)
	) name6374 (
		_w6826_,
		_w6829_,
		_w6836_
	);
	LUT2 #(
		.INIT('h4)
	) name6375 (
		_w6832_,
		_w6836_,
		_w6837_
	);
	LUT2 #(
		.INIT('h8)
	) name6376 (
		_w6835_,
		_w6837_,
		_w6838_
	);
	LUT2 #(
		.INIT('h2)
	) name6377 (
		_w3450_,
		_w6838_,
		_w6839_
	);
	LUT2 #(
		.INIT('h1)
	) name6378 (
		_w6818_,
		_w6839_,
		_w6840_
	);
	LUT2 #(
		.INIT('h2)
	) name6379 (
		\P1_state_reg[0]/NET0131 ,
		_w6840_,
		_w6841_
	);
	LUT2 #(
		.INIT('h1)
	) name6380 (
		_w6817_,
		_w6841_,
		_w6842_
	);
	LUT2 #(
		.INIT('h2)
	) name6381 (
		\P1_reg0_reg[19]/NET0131 ,
		_w3435_,
		_w6843_
	);
	LUT2 #(
		.INIT('h8)
	) name6382 (
		\P1_reg0_reg[19]/NET0131 ,
		_w3448_,
		_w6844_
	);
	LUT2 #(
		.INIT('h4)
	) name6383 (
		_w1936_,
		_w3563_,
		_w6845_
	);
	LUT2 #(
		.INIT('h8)
	) name6384 (
		_w3677_,
		_w6845_,
		_w6846_
	);
	LUT2 #(
		.INIT('h1)
	) name6385 (
		_w4396_,
		_w6846_,
		_w6847_
	);
	LUT2 #(
		.INIT('h2)
	) name6386 (
		_w4494_,
		_w6847_,
		_w6848_
	);
	LUT2 #(
		.INIT('h2)
	) name6387 (
		\P1_reg0_reg[19]/NET0131 ,
		_w6848_,
		_w6849_
	);
	LUT2 #(
		.INIT('h2)
	) name6388 (
		_w1936_,
		_w5654_,
		_w6850_
	);
	LUT2 #(
		.INIT('h8)
	) name6389 (
		_w1418_,
		_w1880_,
		_w6851_
	);
	LUT2 #(
		.INIT('h4)
	) name6390 (
		_w3563_,
		_w5661_,
		_w6852_
	);
	LUT2 #(
		.INIT('h1)
	) name6391 (
		_w3677_,
		_w5667_,
		_w6853_
	);
	LUT2 #(
		.INIT('h1)
	) name6392 (
		_w5674_,
		_w6851_,
		_w6854_
	);
	LUT2 #(
		.INIT('h4)
	) name6393 (
		_w6852_,
		_w6854_,
		_w6855_
	);
	LUT2 #(
		.INIT('h4)
	) name6394 (
		_w6853_,
		_w6855_,
		_w6856_
	);
	LUT2 #(
		.INIT('h4)
	) name6395 (
		_w6850_,
		_w6856_,
		_w6857_
	);
	LUT2 #(
		.INIT('h2)
	) name6396 (
		_w4396_,
		_w6857_,
		_w6858_
	);
	LUT2 #(
		.INIT('h1)
	) name6397 (
		_w6849_,
		_w6858_,
		_w6859_
	);
	LUT2 #(
		.INIT('h2)
	) name6398 (
		_w3450_,
		_w6859_,
		_w6860_
	);
	LUT2 #(
		.INIT('h1)
	) name6399 (
		_w6844_,
		_w6860_,
		_w6861_
	);
	LUT2 #(
		.INIT('h2)
	) name6400 (
		\P1_state_reg[0]/NET0131 ,
		_w6861_,
		_w6862_
	);
	LUT2 #(
		.INIT('h1)
	) name6401 (
		_w6843_,
		_w6862_,
		_w6863_
	);
	LUT2 #(
		.INIT('h2)
	) name6402 (
		\P1_reg0_reg[22]/NET0131 ,
		_w3435_,
		_w6864_
	);
	LUT2 #(
		.INIT('h8)
	) name6403 (
		\P1_reg0_reg[22]/NET0131 ,
		_w3448_,
		_w6865_
	);
	LUT2 #(
		.INIT('h2)
	) name6404 (
		\P1_reg0_reg[22]/NET0131 ,
		_w4396_,
		_w6866_
	);
	LUT2 #(
		.INIT('h2)
	) name6405 (
		_w4396_,
		_w6038_,
		_w6867_
	);
	LUT2 #(
		.INIT('h1)
	) name6406 (
		_w6866_,
		_w6867_,
		_w6868_
	);
	LUT2 #(
		.INIT('h1)
	) name6407 (
		_w3563_,
		_w6868_,
		_w6869_
	);
	LUT2 #(
		.INIT('h8)
	) name6408 (
		_w4396_,
		_w6026_,
		_w6870_
	);
	LUT2 #(
		.INIT('h1)
	) name6409 (
		_w6866_,
		_w6870_,
		_w6871_
	);
	LUT2 #(
		.INIT('h1)
	) name6410 (
		_w3677_,
		_w6871_,
		_w6872_
	);
	LUT2 #(
		.INIT('h2)
	) name6411 (
		\P1_reg0_reg[22]/NET0131 ,
		_w4494_,
		_w6873_
	);
	LUT2 #(
		.INIT('h2)
	) name6412 (
		_w4396_,
		_w6048_,
		_w6874_
	);
	LUT2 #(
		.INIT('h1)
	) name6413 (
		_w6866_,
		_w6874_,
		_w6875_
	);
	LUT2 #(
		.INIT('h2)
	) name6414 (
		_w1936_,
		_w6875_,
		_w6876_
	);
	LUT2 #(
		.INIT('h2)
	) name6415 (
		_w4396_,
		_w6057_,
		_w6877_
	);
	LUT2 #(
		.INIT('h1)
	) name6416 (
		_w6873_,
		_w6877_,
		_w6878_
	);
	LUT2 #(
		.INIT('h4)
	) name6417 (
		_w6876_,
		_w6878_,
		_w6879_
	);
	LUT2 #(
		.INIT('h4)
	) name6418 (
		_w6869_,
		_w6879_,
		_w6880_
	);
	LUT2 #(
		.INIT('h4)
	) name6419 (
		_w6872_,
		_w6880_,
		_w6881_
	);
	LUT2 #(
		.INIT('h2)
	) name6420 (
		_w3450_,
		_w6881_,
		_w6882_
	);
	LUT2 #(
		.INIT('h1)
	) name6421 (
		_w6865_,
		_w6882_,
		_w6883_
	);
	LUT2 #(
		.INIT('h2)
	) name6422 (
		\P1_state_reg[0]/NET0131 ,
		_w6883_,
		_w6884_
	);
	LUT2 #(
		.INIT('h1)
	) name6423 (
		_w6864_,
		_w6884_,
		_w6885_
	);
	LUT2 #(
		.INIT('h8)
	) name6424 (
		_w4396_,
		_w5812_,
		_w6886_
	);
	LUT2 #(
		.INIT('h8)
	) name6425 (
		_w4491_,
		_w6886_,
		_w6887_
	);
	LUT2 #(
		.INIT('h2)
	) name6426 (
		\P1_reg0_reg[31]/NET0131 ,
		_w6887_,
		_w6888_
	);
	LUT2 #(
		.INIT('h4)
	) name6427 (
		_w5809_,
		_w6886_,
		_w6889_
	);
	LUT2 #(
		.INIT('h1)
	) name6428 (
		_w6888_,
		_w6889_,
		_w6890_
	);
	LUT2 #(
		.INIT('h2)
	) name6429 (
		\P1_reg1_reg[17]/NET0131 ,
		_w3435_,
		_w6891_
	);
	LUT2 #(
		.INIT('h8)
	) name6430 (
		\P1_reg1_reg[17]/NET0131 ,
		_w3448_,
		_w6892_
	);
	LUT2 #(
		.INIT('h2)
	) name6431 (
		\P1_reg1_reg[17]/NET0131 ,
		_w4541_,
		_w6893_
	);
	LUT2 #(
		.INIT('h8)
	) name6432 (
		_w4532_,
		_w6442_,
		_w6894_
	);
	LUT2 #(
		.INIT('h2)
	) name6433 (
		\P1_reg1_reg[17]/NET0131 ,
		_w4532_,
		_w6895_
	);
	LUT2 #(
		.INIT('h8)
	) name6434 (
		_w4532_,
		_w5436_,
		_w6896_
	);
	LUT2 #(
		.INIT('h1)
	) name6435 (
		_w6895_,
		_w6896_,
		_w6897_
	);
	LUT2 #(
		.INIT('h1)
	) name6436 (
		_w3677_,
		_w6897_,
		_w6898_
	);
	LUT2 #(
		.INIT('h8)
	) name6437 (
		_w4532_,
		_w5445_,
		_w6899_
	);
	LUT2 #(
		.INIT('h1)
	) name6438 (
		_w6895_,
		_w6899_,
		_w6900_
	);
	LUT2 #(
		.INIT('h2)
	) name6439 (
		_w3712_,
		_w6900_,
		_w6901_
	);
	LUT2 #(
		.INIT('h2)
	) name6440 (
		_w4532_,
		_w5453_,
		_w6902_
	);
	LUT2 #(
		.INIT('h1)
	) name6441 (
		_w6895_,
		_w6902_,
		_w6903_
	);
	LUT2 #(
		.INIT('h1)
	) name6442 (
		_w3563_,
		_w6903_,
		_w6904_
	);
	LUT2 #(
		.INIT('h8)
	) name6443 (
		_w4532_,
		_w5462_,
		_w6905_
	);
	LUT2 #(
		.INIT('h1)
	) name6444 (
		_w6895_,
		_w6905_,
		_w6906_
	);
	LUT2 #(
		.INIT('h2)
	) name6445 (
		_w1936_,
		_w6906_,
		_w6907_
	);
	LUT2 #(
		.INIT('h1)
	) name6446 (
		_w6893_,
		_w6894_,
		_w6908_
	);
	LUT2 #(
		.INIT('h4)
	) name6447 (
		_w6901_,
		_w6908_,
		_w6909_
	);
	LUT2 #(
		.INIT('h4)
	) name6448 (
		_w6907_,
		_w6909_,
		_w6910_
	);
	LUT2 #(
		.INIT('h1)
	) name6449 (
		_w6898_,
		_w6904_,
		_w6911_
	);
	LUT2 #(
		.INIT('h8)
	) name6450 (
		_w6910_,
		_w6911_,
		_w6912_
	);
	LUT2 #(
		.INIT('h2)
	) name6451 (
		_w3450_,
		_w6912_,
		_w6913_
	);
	LUT2 #(
		.INIT('h1)
	) name6452 (
		_w6892_,
		_w6913_,
		_w6914_
	);
	LUT2 #(
		.INIT('h2)
	) name6453 (
		\P1_state_reg[0]/NET0131 ,
		_w6914_,
		_w6915_
	);
	LUT2 #(
		.INIT('h1)
	) name6454 (
		_w6891_,
		_w6915_,
		_w6916_
	);
	LUT2 #(
		.INIT('h2)
	) name6455 (
		\P1_reg1_reg[18]/NET0131 ,
		_w3435_,
		_w6917_
	);
	LUT2 #(
		.INIT('h8)
	) name6456 (
		\P1_reg1_reg[18]/NET0131 ,
		_w3448_,
		_w6918_
	);
	LUT2 #(
		.INIT('h8)
	) name6457 (
		_w4532_,
		_w6413_,
		_w6919_
	);
	LUT2 #(
		.INIT('h2)
	) name6458 (
		\P1_reg1_reg[18]/NET0131 ,
		_w4532_,
		_w6920_
	);
	LUT2 #(
		.INIT('h8)
	) name6459 (
		_w4532_,
		_w5482_,
		_w6921_
	);
	LUT2 #(
		.INIT('h1)
	) name6460 (
		_w6920_,
		_w6921_,
		_w6922_
	);
	LUT2 #(
		.INIT('h2)
	) name6461 (
		_w3712_,
		_w6922_,
		_w6923_
	);
	LUT2 #(
		.INIT('h2)
	) name6462 (
		_w4532_,
		_w5504_,
		_w6924_
	);
	LUT2 #(
		.INIT('h1)
	) name6463 (
		_w6920_,
		_w6924_,
		_w6925_
	);
	LUT2 #(
		.INIT('h1)
	) name6464 (
		_w3677_,
		_w6925_,
		_w6926_
	);
	LUT2 #(
		.INIT('h8)
	) name6465 (
		_w4532_,
		_w5527_,
		_w6927_
	);
	LUT2 #(
		.INIT('h1)
	) name6466 (
		_w6920_,
		_w6927_,
		_w6928_
	);
	LUT2 #(
		.INIT('h1)
	) name6467 (
		_w3563_,
		_w6928_,
		_w6929_
	);
	LUT2 #(
		.INIT('h2)
	) name6468 (
		_w4532_,
		_w5536_,
		_w6930_
	);
	LUT2 #(
		.INIT('h1)
	) name6469 (
		_w6920_,
		_w6930_,
		_w6931_
	);
	LUT2 #(
		.INIT('h2)
	) name6470 (
		_w1936_,
		_w6931_,
		_w6932_
	);
	LUT2 #(
		.INIT('h2)
	) name6471 (
		\P1_reg1_reg[18]/NET0131 ,
		_w4541_,
		_w6933_
	);
	LUT2 #(
		.INIT('h1)
	) name6472 (
		_w6919_,
		_w6933_,
		_w6934_
	);
	LUT2 #(
		.INIT('h4)
	) name6473 (
		_w6923_,
		_w6934_,
		_w6935_
	);
	LUT2 #(
		.INIT('h1)
	) name6474 (
		_w6926_,
		_w6929_,
		_w6936_
	);
	LUT2 #(
		.INIT('h4)
	) name6475 (
		_w6932_,
		_w6936_,
		_w6937_
	);
	LUT2 #(
		.INIT('h8)
	) name6476 (
		_w6935_,
		_w6937_,
		_w6938_
	);
	LUT2 #(
		.INIT('h2)
	) name6477 (
		_w3450_,
		_w6938_,
		_w6939_
	);
	LUT2 #(
		.INIT('h1)
	) name6478 (
		_w6918_,
		_w6939_,
		_w6940_
	);
	LUT2 #(
		.INIT('h2)
	) name6479 (
		\P1_state_reg[0]/NET0131 ,
		_w6940_,
		_w6941_
	);
	LUT2 #(
		.INIT('h1)
	) name6480 (
		_w6917_,
		_w6941_,
		_w6942_
	);
	LUT2 #(
		.INIT('h2)
	) name6481 (
		\P1_reg1_reg[19]/NET0131 ,
		_w3435_,
		_w6943_
	);
	LUT2 #(
		.INIT('h8)
	) name6482 (
		\P1_reg1_reg[19]/NET0131 ,
		_w3448_,
		_w6944_
	);
	LUT2 #(
		.INIT('h8)
	) name6483 (
		_w4491_,
		_w4532_,
		_w6945_
	);
	LUT2 #(
		.INIT('h2)
	) name6484 (
		\P1_reg1_reg[19]/NET0131 ,
		_w6945_,
		_w6946_
	);
	LUT2 #(
		.INIT('h2)
	) name6485 (
		_w4532_,
		_w6857_,
		_w6947_
	);
	LUT2 #(
		.INIT('h1)
	) name6486 (
		_w6946_,
		_w6947_,
		_w6948_
	);
	LUT2 #(
		.INIT('h2)
	) name6487 (
		_w3450_,
		_w6948_,
		_w6949_
	);
	LUT2 #(
		.INIT('h1)
	) name6488 (
		_w6944_,
		_w6949_,
		_w6950_
	);
	LUT2 #(
		.INIT('h2)
	) name6489 (
		\P1_state_reg[0]/NET0131 ,
		_w6950_,
		_w6951_
	);
	LUT2 #(
		.INIT('h1)
	) name6490 (
		_w6943_,
		_w6951_,
		_w6952_
	);
	LUT2 #(
		.INIT('h2)
	) name6491 (
		\P1_reg1_reg[21]/NET0131 ,
		_w3435_,
		_w6953_
	);
	LUT2 #(
		.INIT('h8)
	) name6492 (
		\P1_reg1_reg[21]/NET0131 ,
		_w3448_,
		_w6954_
	);
	LUT2 #(
		.INIT('h8)
	) name6493 (
		_w1346_,
		_w1880_,
		_w6955_
	);
	LUT2 #(
		.INIT('h8)
	) name6494 (
		_w4532_,
		_w6955_,
		_w6956_
	);
	LUT2 #(
		.INIT('h2)
	) name6495 (
		\P1_reg1_reg[21]/NET0131 ,
		_w4532_,
		_w6957_
	);
	LUT2 #(
		.INIT('h2)
	) name6496 (
		_w1318_,
		_w5795_,
		_w6958_
	);
	LUT2 #(
		.INIT('h1)
	) name6497 (
		_w6044_,
		_w6958_,
		_w6959_
	);
	LUT2 #(
		.INIT('h1)
	) name6498 (
		_w537_,
		_w6959_,
		_w6960_
	);
	LUT2 #(
		.INIT('h8)
	) name6499 (
		_w537_,
		_w1374_,
		_w6961_
	);
	LUT2 #(
		.INIT('h1)
	) name6500 (
		_w6960_,
		_w6961_,
		_w6962_
	);
	LUT2 #(
		.INIT('h8)
	) name6501 (
		_w4532_,
		_w6962_,
		_w6963_
	);
	LUT2 #(
		.INIT('h1)
	) name6502 (
		_w6957_,
		_w6963_,
		_w6964_
	);
	LUT2 #(
		.INIT('h2)
	) name6503 (
		_w1936_,
		_w6964_,
		_w6965_
	);
	LUT2 #(
		.INIT('h8)
	) name6504 (
		_w1841_,
		_w3550_,
		_w6966_
	);
	LUT2 #(
		.INIT('h1)
	) name6505 (
		_w1841_,
		_w3550_,
		_w6967_
	);
	LUT2 #(
		.INIT('h1)
	) name6506 (
		_w6966_,
		_w6967_,
		_w6968_
	);
	LUT2 #(
		.INIT('h2)
	) name6507 (
		_w4532_,
		_w6968_,
		_w6969_
	);
	LUT2 #(
		.INIT('h1)
	) name6508 (
		_w6957_,
		_w6969_,
		_w6970_
	);
	LUT2 #(
		.INIT('h1)
	) name6509 (
		_w3563_,
		_w6970_,
		_w6971_
	);
	LUT2 #(
		.INIT('h8)
	) name6510 (
		_w1841_,
		_w3664_,
		_w6972_
	);
	LUT2 #(
		.INIT('h1)
	) name6511 (
		_w1841_,
		_w3664_,
		_w6973_
	);
	LUT2 #(
		.INIT('h1)
	) name6512 (
		_w6972_,
		_w6973_,
		_w6974_
	);
	LUT2 #(
		.INIT('h8)
	) name6513 (
		_w4532_,
		_w6974_,
		_w6975_
	);
	LUT2 #(
		.INIT('h1)
	) name6514 (
		_w6957_,
		_w6975_,
		_w6976_
	);
	LUT2 #(
		.INIT('h1)
	) name6515 (
		_w3677_,
		_w6976_,
		_w6977_
	);
	LUT2 #(
		.INIT('h2)
	) name6516 (
		_w1346_,
		_w3698_,
		_w6978_
	);
	LUT2 #(
		.INIT('h1)
	) name6517 (
		_w6052_,
		_w6978_,
		_w6979_
	);
	LUT2 #(
		.INIT('h8)
	) name6518 (
		_w4532_,
		_w6979_,
		_w6980_
	);
	LUT2 #(
		.INIT('h1)
	) name6519 (
		_w6957_,
		_w6980_,
		_w6981_
	);
	LUT2 #(
		.INIT('h2)
	) name6520 (
		_w3712_,
		_w6981_,
		_w6982_
	);
	LUT2 #(
		.INIT('h2)
	) name6521 (
		\P1_reg1_reg[21]/NET0131 ,
		_w4541_,
		_w6983_
	);
	LUT2 #(
		.INIT('h1)
	) name6522 (
		_w6956_,
		_w6983_,
		_w6984_
	);
	LUT2 #(
		.INIT('h4)
	) name6523 (
		_w6982_,
		_w6984_,
		_w6985_
	);
	LUT2 #(
		.INIT('h4)
	) name6524 (
		_w6965_,
		_w6985_,
		_w6986_
	);
	LUT2 #(
		.INIT('h1)
	) name6525 (
		_w6971_,
		_w6977_,
		_w6987_
	);
	LUT2 #(
		.INIT('h8)
	) name6526 (
		_w6986_,
		_w6987_,
		_w6988_
	);
	LUT2 #(
		.INIT('h2)
	) name6527 (
		_w3450_,
		_w6988_,
		_w6989_
	);
	LUT2 #(
		.INIT('h1)
	) name6528 (
		_w6954_,
		_w6989_,
		_w6990_
	);
	LUT2 #(
		.INIT('h2)
	) name6529 (
		\P1_state_reg[0]/NET0131 ,
		_w6990_,
		_w6991_
	);
	LUT2 #(
		.INIT('h1)
	) name6530 (
		_w6953_,
		_w6991_,
		_w6992_
	);
	LUT2 #(
		.INIT('h2)
	) name6531 (
		\P2_reg0_reg[17]/NET0131 ,
		_w1983_,
		_w6993_
	);
	LUT2 #(
		.INIT('h8)
	) name6532 (
		\P2_reg0_reg[17]/NET0131 ,
		_w2024_,
		_w6994_
	);
	LUT2 #(
		.INIT('h2)
	) name6533 (
		\P2_reg0_reg[17]/NET0131 ,
		_w3423_,
		_w6995_
	);
	LUT2 #(
		.INIT('h2)
	) name6534 (
		\P2_reg0_reg[17]/NET0131 ,
		_w2040_,
		_w6996_
	);
	LUT2 #(
		.INIT('h8)
	) name6535 (
		_w2040_,
		_w5558_,
		_w6997_
	);
	LUT2 #(
		.INIT('h1)
	) name6536 (
		_w6996_,
		_w6997_,
		_w6998_
	);
	LUT2 #(
		.INIT('h1)
	) name6537 (
		_w3177_,
		_w6998_,
		_w6999_
	);
	LUT2 #(
		.INIT('h2)
	) name6538 (
		_w2040_,
		_w5570_,
		_w7000_
	);
	LUT2 #(
		.INIT('h1)
	) name6539 (
		_w6996_,
		_w7000_,
		_w7001_
	);
	LUT2 #(
		.INIT('h2)
	) name6540 (
		_w3411_,
		_w7001_,
		_w7002_
	);
	LUT2 #(
		.INIT('h8)
	) name6541 (
		_w2040_,
		_w5578_,
		_w7003_
	);
	LUT2 #(
		.INIT('h1)
	) name6542 (
		_w6996_,
		_w7003_,
		_w7004_
	);
	LUT2 #(
		.INIT('h2)
	) name6543 (
		_w3355_,
		_w7004_,
		_w7005_
	);
	LUT2 #(
		.INIT('h8)
	) name6544 (
		_w2040_,
		_w5586_,
		_w7006_
	);
	LUT2 #(
		.INIT('h1)
	) name6545 (
		_w6996_,
		_w7006_,
		_w7007_
	);
	LUT2 #(
		.INIT('h1)
	) name6546 (
		_w3320_,
		_w7007_,
		_w7008_
	);
	LUT2 #(
		.INIT('h8)
	) name6547 (
		_w2040_,
		_w6529_,
		_w7009_
	);
	LUT2 #(
		.INIT('h1)
	) name6548 (
		_w6995_,
		_w7009_,
		_w7010_
	);
	LUT2 #(
		.INIT('h4)
	) name6549 (
		_w7008_,
		_w7010_,
		_w7011_
	);
	LUT2 #(
		.INIT('h4)
	) name6550 (
		_w6999_,
		_w7011_,
		_w7012_
	);
	LUT2 #(
		.INIT('h1)
	) name6551 (
		_w7002_,
		_w7005_,
		_w7013_
	);
	LUT2 #(
		.INIT('h8)
	) name6552 (
		_w7012_,
		_w7013_,
		_w7014_
	);
	LUT2 #(
		.INIT('h2)
	) name6553 (
		_w2026_,
		_w7014_,
		_w7015_
	);
	LUT2 #(
		.INIT('h1)
	) name6554 (
		_w6994_,
		_w7015_,
		_w7016_
	);
	LUT2 #(
		.INIT('h2)
	) name6555 (
		\P1_state_reg[0]/NET0131 ,
		_w7016_,
		_w7017_
	);
	LUT2 #(
		.INIT('h1)
	) name6556 (
		_w6993_,
		_w7017_,
		_w7018_
	);
	LUT2 #(
		.INIT('h2)
	) name6557 (
		\P2_reg0_reg[18]/NET0131 ,
		_w1983_,
		_w7019_
	);
	LUT2 #(
		.INIT('h8)
	) name6558 (
		\P2_reg0_reg[18]/NET0131 ,
		_w2024_,
		_w7020_
	);
	LUT2 #(
		.INIT('h8)
	) name6559 (
		_w2040_,
		_w6356_,
		_w7021_
	);
	LUT2 #(
		.INIT('h2)
	) name6560 (
		\P2_reg0_reg[18]/NET0131 ,
		_w2040_,
		_w7022_
	);
	LUT2 #(
		.INIT('h8)
	) name6561 (
		_w2040_,
		_w6331_,
		_w7023_
	);
	LUT2 #(
		.INIT('h1)
	) name6562 (
		_w7022_,
		_w7023_,
		_w7024_
	);
	LUT2 #(
		.INIT('h2)
	) name6563 (
		_w3355_,
		_w7024_,
		_w7025_
	);
	LUT2 #(
		.INIT('h8)
	) name6564 (
		_w2040_,
		_w6337_,
		_w7026_
	);
	LUT2 #(
		.INIT('h1)
	) name6565 (
		_w7022_,
		_w7026_,
		_w7027_
	);
	LUT2 #(
		.INIT('h1)
	) name6566 (
		_w3177_,
		_w7027_,
		_w7028_
	);
	LUT2 #(
		.INIT('h2)
	) name6567 (
		_w2040_,
		_w6343_,
		_w7029_
	);
	LUT2 #(
		.INIT('h1)
	) name6568 (
		_w7022_,
		_w7029_,
		_w7030_
	);
	LUT2 #(
		.INIT('h1)
	) name6569 (
		_w3320_,
		_w7030_,
		_w7031_
	);
	LUT2 #(
		.INIT('h8)
	) name6570 (
		_w2040_,
		_w6351_,
		_w7032_
	);
	LUT2 #(
		.INIT('h1)
	) name6571 (
		_w7022_,
		_w7032_,
		_w7033_
	);
	LUT2 #(
		.INIT('h2)
	) name6572 (
		_w3411_,
		_w7033_,
		_w7034_
	);
	LUT2 #(
		.INIT('h2)
	) name6573 (
		\P2_reg0_reg[18]/NET0131 ,
		_w3423_,
		_w7035_
	);
	LUT2 #(
		.INIT('h1)
	) name6574 (
		_w7021_,
		_w7035_,
		_w7036_
	);
	LUT2 #(
		.INIT('h4)
	) name6575 (
		_w7034_,
		_w7036_,
		_w7037_
	);
	LUT2 #(
		.INIT('h4)
	) name6576 (
		_w7028_,
		_w7037_,
		_w7038_
	);
	LUT2 #(
		.INIT('h4)
	) name6577 (
		_w7031_,
		_w7038_,
		_w7039_
	);
	LUT2 #(
		.INIT('h4)
	) name6578 (
		_w7025_,
		_w7039_,
		_w7040_
	);
	LUT2 #(
		.INIT('h2)
	) name6579 (
		_w2026_,
		_w7040_,
		_w7041_
	);
	LUT2 #(
		.INIT('h1)
	) name6580 (
		_w7020_,
		_w7041_,
		_w7042_
	);
	LUT2 #(
		.INIT('h2)
	) name6581 (
		\P1_state_reg[0]/NET0131 ,
		_w7042_,
		_w7043_
	);
	LUT2 #(
		.INIT('h1)
	) name6582 (
		_w7019_,
		_w7043_,
		_w7044_
	);
	LUT2 #(
		.INIT('h2)
	) name6583 (
		\P2_reg0_reg[19]/NET0131 ,
		_w1983_,
		_w7045_
	);
	LUT2 #(
		.INIT('h8)
	) name6584 (
		\P2_reg0_reg[19]/NET0131 ,
		_w2024_,
		_w7046_
	);
	LUT2 #(
		.INIT('h8)
	) name6585 (
		_w2040_,
		_w6626_,
		_w7047_
	);
	LUT2 #(
		.INIT('h2)
	) name6586 (
		\P2_reg0_reg[19]/NET0131 ,
		_w2040_,
		_w7048_
	);
	LUT2 #(
		.INIT('h8)
	) name6587 (
		_w2040_,
		_w5608_,
		_w7049_
	);
	LUT2 #(
		.INIT('h1)
	) name6588 (
		_w7048_,
		_w7049_,
		_w7050_
	);
	LUT2 #(
		.INIT('h1)
	) name6589 (
		_w3177_,
		_w7050_,
		_w7051_
	);
	LUT2 #(
		.INIT('h2)
	) name6590 (
		_w2040_,
		_w5614_,
		_w7052_
	);
	LUT2 #(
		.INIT('h1)
	) name6591 (
		_w7048_,
		_w7052_,
		_w7053_
	);
	LUT2 #(
		.INIT('h1)
	) name6592 (
		_w3320_,
		_w7053_,
		_w7054_
	);
	LUT2 #(
		.INIT('h8)
	) name6593 (
		_w2040_,
		_w5624_,
		_w7055_
	);
	LUT2 #(
		.INIT('h1)
	) name6594 (
		_w7048_,
		_w7055_,
		_w7056_
	);
	LUT2 #(
		.INIT('h2)
	) name6595 (
		_w3411_,
		_w7056_,
		_w7057_
	);
	LUT2 #(
		.INIT('h8)
	) name6596 (
		_w2040_,
		_w5630_,
		_w7058_
	);
	LUT2 #(
		.INIT('h1)
	) name6597 (
		_w7048_,
		_w7058_,
		_w7059_
	);
	LUT2 #(
		.INIT('h2)
	) name6598 (
		_w3355_,
		_w7059_,
		_w7060_
	);
	LUT2 #(
		.INIT('h2)
	) name6599 (
		\P2_reg0_reg[19]/NET0131 ,
		_w3423_,
		_w7061_
	);
	LUT2 #(
		.INIT('h1)
	) name6600 (
		_w7047_,
		_w7061_,
		_w7062_
	);
	LUT2 #(
		.INIT('h4)
	) name6601 (
		_w7054_,
		_w7062_,
		_w7063_
	);
	LUT2 #(
		.INIT('h4)
	) name6602 (
		_w7060_,
		_w7063_,
		_w7064_
	);
	LUT2 #(
		.INIT('h4)
	) name6603 (
		_w7057_,
		_w7064_,
		_w7065_
	);
	LUT2 #(
		.INIT('h4)
	) name6604 (
		_w7051_,
		_w7065_,
		_w7066_
	);
	LUT2 #(
		.INIT('h2)
	) name6605 (
		_w2026_,
		_w7066_,
		_w7067_
	);
	LUT2 #(
		.INIT('h1)
	) name6606 (
		_w7046_,
		_w7067_,
		_w7068_
	);
	LUT2 #(
		.INIT('h2)
	) name6607 (
		\P1_state_reg[0]/NET0131 ,
		_w7068_,
		_w7069_
	);
	LUT2 #(
		.INIT('h1)
	) name6608 (
		_w7045_,
		_w7069_,
		_w7070_
	);
	LUT2 #(
		.INIT('h2)
	) name6609 (
		\P1_reg3_reg[10]/NET0131 ,
		\P1_state_reg[0]/NET0131 ,
		_w7071_
	);
	LUT2 #(
		.INIT('h8)
	) name6610 (
		_w1214_,
		_w1953_,
		_w7072_
	);
	LUT2 #(
		.INIT('h8)
	) name6611 (
		_w1214_,
		_w3448_,
		_w7073_
	);
	LUT2 #(
		.INIT('h2)
	) name6612 (
		_w1233_,
		_w4067_,
		_w7074_
	);
	LUT2 #(
		.INIT('h2)
	) name6613 (
		_w1214_,
		_w3980_,
		_w7075_
	);
	LUT2 #(
		.INIT('h2)
	) name6614 (
		_w1791_,
		_w5491_,
		_w7076_
	);
	LUT2 #(
		.INIT('h4)
	) name6615 (
		_w1791_,
		_w5491_,
		_w7077_
	);
	LUT2 #(
		.INIT('h1)
	) name6616 (
		_w7076_,
		_w7077_,
		_w7078_
	);
	LUT2 #(
		.INIT('h2)
	) name6617 (
		_w3980_,
		_w7078_,
		_w7079_
	);
	LUT2 #(
		.INIT('h1)
	) name6618 (
		_w7075_,
		_w7079_,
		_w7080_
	);
	LUT2 #(
		.INIT('h1)
	) name6619 (
		_w3677_,
		_w7080_,
		_w7081_
	);
	LUT2 #(
		.INIT('h2)
	) name6620 (
		_w1207_,
		_w3580_,
		_w7082_
	);
	LUT2 #(
		.INIT('h1)
	) name6621 (
		_w4069_,
		_w7082_,
		_w7083_
	);
	LUT2 #(
		.INIT('h1)
	) name6622 (
		_w537_,
		_w7083_,
		_w7084_
	);
	LUT2 #(
		.INIT('h8)
	) name6623 (
		_w537_,
		_w1244_,
		_w7085_
	);
	LUT2 #(
		.INIT('h1)
	) name6624 (
		_w7084_,
		_w7085_,
		_w7086_
	);
	LUT2 #(
		.INIT('h8)
	) name6625 (
		_w3980_,
		_w7086_,
		_w7087_
	);
	LUT2 #(
		.INIT('h1)
	) name6626 (
		_w7075_,
		_w7087_,
		_w7088_
	);
	LUT2 #(
		.INIT('h2)
	) name6627 (
		_w1936_,
		_w7088_,
		_w7089_
	);
	LUT2 #(
		.INIT('h2)
	) name6628 (
		_w1791_,
		_w5514_,
		_w7090_
	);
	LUT2 #(
		.INIT('h4)
	) name6629 (
		_w1791_,
		_w5514_,
		_w7091_
	);
	LUT2 #(
		.INIT('h1)
	) name6630 (
		_w7090_,
		_w7091_,
		_w7092_
	);
	LUT2 #(
		.INIT('h8)
	) name6631 (
		_w3980_,
		_w7092_,
		_w7093_
	);
	LUT2 #(
		.INIT('h1)
	) name6632 (
		_w7075_,
		_w7093_,
		_w7094_
	);
	LUT2 #(
		.INIT('h1)
	) name6633 (
		_w3563_,
		_w7094_,
		_w7095_
	);
	LUT2 #(
		.INIT('h2)
	) name6634 (
		_w1233_,
		_w3687_,
		_w7096_
	);
	LUT2 #(
		.INIT('h1)
	) name6635 (
		_w6114_,
		_w7096_,
		_w7097_
	);
	LUT2 #(
		.INIT('h8)
	) name6636 (
		_w3980_,
		_w7097_,
		_w7098_
	);
	LUT2 #(
		.INIT('h1)
	) name6637 (
		_w7075_,
		_w7098_,
		_w7099_
	);
	LUT2 #(
		.INIT('h2)
	) name6638 (
		_w3712_,
		_w7099_,
		_w7100_
	);
	LUT2 #(
		.INIT('h2)
	) name6639 (
		_w1214_,
		_w4064_,
		_w7101_
	);
	LUT2 #(
		.INIT('h1)
	) name6640 (
		_w7074_,
		_w7101_,
		_w7102_
	);
	LUT2 #(
		.INIT('h4)
	) name6641 (
		_w7100_,
		_w7102_,
		_w7103_
	);
	LUT2 #(
		.INIT('h4)
	) name6642 (
		_w7081_,
		_w7103_,
		_w7104_
	);
	LUT2 #(
		.INIT('h1)
	) name6643 (
		_w7089_,
		_w7095_,
		_w7105_
	);
	LUT2 #(
		.INIT('h8)
	) name6644 (
		_w7104_,
		_w7105_,
		_w7106_
	);
	LUT2 #(
		.INIT('h2)
	) name6645 (
		_w3450_,
		_w7106_,
		_w7107_
	);
	LUT2 #(
		.INIT('h1)
	) name6646 (
		_w7073_,
		_w7107_,
		_w7108_
	);
	LUT2 #(
		.INIT('h2)
	) name6647 (
		\P1_state_reg[0]/NET0131 ,
		_w7108_,
		_w7109_
	);
	LUT2 #(
		.INIT('h1)
	) name6648 (
		_w7071_,
		_w7072_,
		_w7110_
	);
	LUT2 #(
		.INIT('h4)
	) name6649 (
		_w7109_,
		_w7110_,
		_w7111_
	);
	LUT2 #(
		.INIT('h8)
	) name6650 (
		_w1140_,
		_w1953_,
		_w7112_
	);
	LUT2 #(
		.INIT('h2)
	) name6651 (
		\P1_reg3_reg[13]/NET0131 ,
		\P1_state_reg[0]/NET0131 ,
		_w7113_
	);
	LUT2 #(
		.INIT('h8)
	) name6652 (
		_w1140_,
		_w3448_,
		_w7114_
	);
	LUT2 #(
		.INIT('h2)
	) name6653 (
		_w1136_,
		_w4067_,
		_w7115_
	);
	LUT2 #(
		.INIT('h2)
	) name6654 (
		_w1140_,
		_w3980_,
		_w7116_
	);
	LUT2 #(
		.INIT('h2)
	) name6655 (
		_w1799_,
		_w3650_,
		_w7117_
	);
	LUT2 #(
		.INIT('h4)
	) name6656 (
		_w1799_,
		_w3650_,
		_w7118_
	);
	LUT2 #(
		.INIT('h1)
	) name6657 (
		_w7117_,
		_w7118_,
		_w7119_
	);
	LUT2 #(
		.INIT('h2)
	) name6658 (
		_w3980_,
		_w7119_,
		_w7120_
	);
	LUT2 #(
		.INIT('h1)
	) name6659 (
		_w7116_,
		_w7120_,
		_w7121_
	);
	LUT2 #(
		.INIT('h1)
	) name6660 (
		_w3677_,
		_w7121_,
		_w7122_
	);
	LUT2 #(
		.INIT('h2)
	) name6661 (
		_w1799_,
		_w3533_,
		_w7123_
	);
	LUT2 #(
		.INIT('h4)
	) name6662 (
		_w1799_,
		_w3533_,
		_w7124_
	);
	LUT2 #(
		.INIT('h1)
	) name6663 (
		_w7123_,
		_w7124_,
		_w7125_
	);
	LUT2 #(
		.INIT('h8)
	) name6664 (
		_w3980_,
		_w7125_,
		_w7126_
	);
	LUT2 #(
		.INIT('h1)
	) name6665 (
		_w7116_,
		_w7126_,
		_w7127_
	);
	LUT2 #(
		.INIT('h1)
	) name6666 (
		_w3563_,
		_w7127_,
		_w7128_
	);
	LUT2 #(
		.INIT('h2)
	) name6667 (
		_w1118_,
		_w3583_,
		_w7129_
	);
	LUT2 #(
		.INIT('h4)
	) name6668 (
		_w1118_,
		_w3583_,
		_w7130_
	);
	LUT2 #(
		.INIT('h1)
	) name6669 (
		_w7129_,
		_w7130_,
		_w7131_
	);
	LUT2 #(
		.INIT('h1)
	) name6670 (
		_w537_,
		_w7131_,
		_w7132_
	);
	LUT2 #(
		.INIT('h8)
	) name6671 (
		_w537_,
		_w1174_,
		_w7133_
	);
	LUT2 #(
		.INIT('h1)
	) name6672 (
		_w7132_,
		_w7133_,
		_w7134_
	);
	LUT2 #(
		.INIT('h8)
	) name6673 (
		_w3980_,
		_w7134_,
		_w7135_
	);
	LUT2 #(
		.INIT('h1)
	) name6674 (
		_w7116_,
		_w7135_,
		_w7136_
	);
	LUT2 #(
		.INIT('h2)
	) name6675 (
		_w1936_,
		_w7136_,
		_w7137_
	);
	LUT2 #(
		.INIT('h2)
	) name6676 (
		_w1136_,
		_w3690_,
		_w7138_
	);
	LUT2 #(
		.INIT('h1)
	) name6677 (
		_w5440_,
		_w7138_,
		_w7139_
	);
	LUT2 #(
		.INIT('h8)
	) name6678 (
		_w3980_,
		_w7139_,
		_w7140_
	);
	LUT2 #(
		.INIT('h1)
	) name6679 (
		_w7116_,
		_w7140_,
		_w7141_
	);
	LUT2 #(
		.INIT('h2)
	) name6680 (
		_w3712_,
		_w7141_,
		_w7142_
	);
	LUT2 #(
		.INIT('h2)
	) name6681 (
		_w1140_,
		_w4064_,
		_w7143_
	);
	LUT2 #(
		.INIT('h1)
	) name6682 (
		_w7115_,
		_w7143_,
		_w7144_
	);
	LUT2 #(
		.INIT('h4)
	) name6683 (
		_w7142_,
		_w7144_,
		_w7145_
	);
	LUT2 #(
		.INIT('h4)
	) name6684 (
		_w7122_,
		_w7145_,
		_w7146_
	);
	LUT2 #(
		.INIT('h1)
	) name6685 (
		_w7128_,
		_w7137_,
		_w7147_
	);
	LUT2 #(
		.INIT('h8)
	) name6686 (
		_w7146_,
		_w7147_,
		_w7148_
	);
	LUT2 #(
		.INIT('h2)
	) name6687 (
		_w3450_,
		_w7148_,
		_w7149_
	);
	LUT2 #(
		.INIT('h1)
	) name6688 (
		_w7114_,
		_w7149_,
		_w7150_
	);
	LUT2 #(
		.INIT('h2)
	) name6689 (
		\P1_state_reg[0]/NET0131 ,
		_w7150_,
		_w7151_
	);
	LUT2 #(
		.INIT('h1)
	) name6690 (
		_w7112_,
		_w7113_,
		_w7152_
	);
	LUT2 #(
		.INIT('h4)
	) name6691 (
		_w7151_,
		_w7152_,
		_w7153_
	);
	LUT2 #(
		.INIT('h4)
	) name6692 (
		\P1_state_reg[0]/NET0131 ,
		\P2_reg3_reg[10]/NET0131 ,
		_w7154_
	);
	LUT2 #(
		.INIT('h8)
	) name6693 (
		_w2735_,
		_w3976_,
		_w7155_
	);
	LUT2 #(
		.INIT('h8)
	) name6694 (
		_w2024_,
		_w2735_,
		_w7156_
	);
	LUT2 #(
		.INIT('h2)
	) name6695 (
		_w2755_,
		_w3965_,
		_w7157_
	);
	LUT2 #(
		.INIT('h2)
	) name6696 (
		_w2735_,
		_w3788_,
		_w7158_
	);
	LUT2 #(
		.INIT('h2)
	) name6697 (
		_w2688_,
		_w3383_,
		_w7159_
	);
	LUT2 #(
		.INIT('h1)
	) name6698 (
		_w6179_,
		_w7159_,
		_w7160_
	);
	LUT2 #(
		.INIT('h1)
	) name6699 (
		_w2058_,
		_w7160_,
		_w7161_
	);
	LUT2 #(
		.INIT('h8)
	) name6700 (
		_w2058_,
		_w2765_,
		_w7162_
	);
	LUT2 #(
		.INIT('h1)
	) name6701 (
		_w7161_,
		_w7162_,
		_w7163_
	);
	LUT2 #(
		.INIT('h8)
	) name6702 (
		_w3788_,
		_w7163_,
		_w7164_
	);
	LUT2 #(
		.INIT('h1)
	) name6703 (
		_w7158_,
		_w7164_,
		_w7165_
	);
	LUT2 #(
		.INIT('h2)
	) name6704 (
		_w3411_,
		_w7165_,
		_w7166_
	);
	LUT2 #(
		.INIT('h2)
	) name6705 (
		_w4195_,
		_w4740_,
		_w7167_
	);
	LUT2 #(
		.INIT('h4)
	) name6706 (
		_w4195_,
		_w4740_,
		_w7168_
	);
	LUT2 #(
		.INIT('h1)
	) name6707 (
		_w7167_,
		_w7168_,
		_w7169_
	);
	LUT2 #(
		.INIT('h2)
	) name6708 (
		_w3788_,
		_w7169_,
		_w7170_
	);
	LUT2 #(
		.INIT('h1)
	) name6709 (
		_w7158_,
		_w7170_,
		_w7171_
	);
	LUT2 #(
		.INIT('h1)
	) name6710 (
		_w3177_,
		_w7171_,
		_w7172_
	);
	LUT2 #(
		.INIT('h2)
	) name6711 (
		_w4195_,
		_w4709_,
		_w7173_
	);
	LUT2 #(
		.INIT('h4)
	) name6712 (
		_w4195_,
		_w4709_,
		_w7174_
	);
	LUT2 #(
		.INIT('h1)
	) name6713 (
		_w7173_,
		_w7174_,
		_w7175_
	);
	LUT2 #(
		.INIT('h8)
	) name6714 (
		_w3788_,
		_w7175_,
		_w7176_
	);
	LUT2 #(
		.INIT('h1)
	) name6715 (
		_w7158_,
		_w7176_,
		_w7177_
	);
	LUT2 #(
		.INIT('h1)
	) name6716 (
		_w3320_,
		_w7177_,
		_w7178_
	);
	LUT2 #(
		.INIT('h4)
	) name6717 (
		_w2755_,
		_w3334_,
		_w7179_
	);
	LUT2 #(
		.INIT('h2)
	) name6718 (
		_w2755_,
		_w3334_,
		_w7180_
	);
	LUT2 #(
		.INIT('h1)
	) name6719 (
		_w7179_,
		_w7180_,
		_w7181_
	);
	LUT2 #(
		.INIT('h8)
	) name6720 (
		_w3788_,
		_w7181_,
		_w7182_
	);
	LUT2 #(
		.INIT('h1)
	) name6721 (
		_w7158_,
		_w7182_,
		_w7183_
	);
	LUT2 #(
		.INIT('h2)
	) name6722 (
		_w3355_,
		_w7183_,
		_w7184_
	);
	LUT2 #(
		.INIT('h2)
	) name6723 (
		_w2735_,
		_w3962_,
		_w7185_
	);
	LUT2 #(
		.INIT('h1)
	) name6724 (
		_w7157_,
		_w7185_,
		_w7186_
	);
	LUT2 #(
		.INIT('h4)
	) name6725 (
		_w7184_,
		_w7186_,
		_w7187_
	);
	LUT2 #(
		.INIT('h4)
	) name6726 (
		_w7172_,
		_w7187_,
		_w7188_
	);
	LUT2 #(
		.INIT('h4)
	) name6727 (
		_w7178_,
		_w7188_,
		_w7189_
	);
	LUT2 #(
		.INIT('h4)
	) name6728 (
		_w7166_,
		_w7189_,
		_w7190_
	);
	LUT2 #(
		.INIT('h2)
	) name6729 (
		_w2026_,
		_w7190_,
		_w7191_
	);
	LUT2 #(
		.INIT('h1)
	) name6730 (
		_w7156_,
		_w7191_,
		_w7192_
	);
	LUT2 #(
		.INIT('h2)
	) name6731 (
		\P1_state_reg[0]/NET0131 ,
		_w7192_,
		_w7193_
	);
	LUT2 #(
		.INIT('h1)
	) name6732 (
		_w7154_,
		_w7155_,
		_w7194_
	);
	LUT2 #(
		.INIT('h4)
	) name6733 (
		_w7193_,
		_w7194_,
		_w7195_
	);
	LUT2 #(
		.INIT('h8)
	) name6734 (
		_w2874_,
		_w3976_,
		_w7196_
	);
	LUT2 #(
		.INIT('h4)
	) name6735 (
		\P1_state_reg[0]/NET0131 ,
		\P2_reg3_reg[13]/NET0131 ,
		_w7197_
	);
	LUT2 #(
		.INIT('h8)
	) name6736 (
		_w2024_,
		_w2874_,
		_w7198_
	);
	LUT2 #(
		.INIT('h2)
	) name6737 (
		_w2893_,
		_w3965_,
		_w7199_
	);
	LUT2 #(
		.INIT('h2)
	) name6738 (
		_w2874_,
		_w3788_,
		_w7200_
	);
	LUT2 #(
		.INIT('h2)
	) name6739 (
		_w2058_,
		_w2715_,
		_w7201_
	);
	LUT2 #(
		.INIT('h2)
	) name6740 (
		_w2870_,
		_w6182_,
		_w7202_
	);
	LUT2 #(
		.INIT('h1)
	) name6741 (
		_w2058_,
		_w3387_,
		_w7203_
	);
	LUT2 #(
		.INIT('h4)
	) name6742 (
		_w7202_,
		_w7203_,
		_w7204_
	);
	LUT2 #(
		.INIT('h1)
	) name6743 (
		_w7201_,
		_w7204_,
		_w7205_
	);
	LUT2 #(
		.INIT('h2)
	) name6744 (
		_w3788_,
		_w7205_,
		_w7206_
	);
	LUT2 #(
		.INIT('h1)
	) name6745 (
		_w7200_,
		_w7206_,
		_w7207_
	);
	LUT2 #(
		.INIT('h2)
	) name6746 (
		_w3411_,
		_w7207_,
		_w7208_
	);
	LUT2 #(
		.INIT('h4)
	) name6747 (
		_w2794_,
		_w4192_,
		_w7209_
	);
	LUT2 #(
		.INIT('h2)
	) name6748 (
		_w2794_,
		_w4192_,
		_w7210_
	);
	LUT2 #(
		.INIT('h1)
	) name6749 (
		_w7209_,
		_w7210_,
		_w7211_
	);
	LUT2 #(
		.INIT('h8)
	) name6750 (
		_w3788_,
		_w7211_,
		_w7212_
	);
	LUT2 #(
		.INIT('h1)
	) name6751 (
		_w7200_,
		_w7212_,
		_w7213_
	);
	LUT2 #(
		.INIT('h1)
	) name6752 (
		_w3177_,
		_w7213_,
		_w7214_
	);
	LUT2 #(
		.INIT('h4)
	) name6753 (
		_w2893_,
		_w3337_,
		_w7215_
	);
	LUT2 #(
		.INIT('h2)
	) name6754 (
		_w2893_,
		_w3337_,
		_w7216_
	);
	LUT2 #(
		.INIT('h1)
	) name6755 (
		_w7215_,
		_w7216_,
		_w7217_
	);
	LUT2 #(
		.INIT('h8)
	) name6756 (
		_w3788_,
		_w7217_,
		_w7218_
	);
	LUT2 #(
		.INIT('h1)
	) name6757 (
		_w7200_,
		_w7218_,
		_w7219_
	);
	LUT2 #(
		.INIT('h2)
	) name6758 (
		_w3355_,
		_w7219_,
		_w7220_
	);
	LUT2 #(
		.INIT('h4)
	) name6759 (
		_w3280_,
		_w4192_,
		_w7221_
	);
	LUT2 #(
		.INIT('h2)
	) name6760 (
		_w3280_,
		_w4192_,
		_w7222_
	);
	LUT2 #(
		.INIT('h1)
	) name6761 (
		_w7221_,
		_w7222_,
		_w7223_
	);
	LUT2 #(
		.INIT('h2)
	) name6762 (
		_w3788_,
		_w7223_,
		_w7224_
	);
	LUT2 #(
		.INIT('h1)
	) name6763 (
		_w7200_,
		_w7224_,
		_w7225_
	);
	LUT2 #(
		.INIT('h1)
	) name6764 (
		_w3320_,
		_w7225_,
		_w7226_
	);
	LUT2 #(
		.INIT('h2)
	) name6765 (
		_w2874_,
		_w3962_,
		_w7227_
	);
	LUT2 #(
		.INIT('h1)
	) name6766 (
		_w7199_,
		_w7227_,
		_w7228_
	);
	LUT2 #(
		.INIT('h4)
	) name6767 (
		_w7226_,
		_w7228_,
		_w7229_
	);
	LUT2 #(
		.INIT('h4)
	) name6768 (
		_w7220_,
		_w7229_,
		_w7230_
	);
	LUT2 #(
		.INIT('h4)
	) name6769 (
		_w7214_,
		_w7230_,
		_w7231_
	);
	LUT2 #(
		.INIT('h4)
	) name6770 (
		_w7208_,
		_w7231_,
		_w7232_
	);
	LUT2 #(
		.INIT('h2)
	) name6771 (
		_w2026_,
		_w7232_,
		_w7233_
	);
	LUT2 #(
		.INIT('h1)
	) name6772 (
		_w7198_,
		_w7233_,
		_w7234_
	);
	LUT2 #(
		.INIT('h2)
	) name6773 (
		\P1_state_reg[0]/NET0131 ,
		_w7234_,
		_w7235_
	);
	LUT2 #(
		.INIT('h1)
	) name6774 (
		_w7196_,
		_w7197_,
		_w7236_
	);
	LUT2 #(
		.INIT('h4)
	) name6775 (
		_w7235_,
		_w7236_,
		_w7237_
	);
	LUT2 #(
		.INIT('h4)
	) name6776 (
		\P1_state_reg[0]/NET0131 ,
		\P2_reg3_reg[9]/NET0131 ,
		_w7238_
	);
	LUT2 #(
		.INIT('h8)
	) name6777 (
		_w2024_,
		_w2760_,
		_w7239_
	);
	LUT2 #(
		.INIT('h2)
	) name6778 (
		_w2760_,
		_w6312_,
		_w7240_
	);
	LUT2 #(
		.INIT('h2)
	) name6779 (
		_w2760_,
		_w3788_,
		_w7241_
	);
	LUT2 #(
		.INIT('h4)
	) name6780 (
		_w2454_,
		_w3380_,
		_w7242_
	);
	LUT2 #(
		.INIT('h4)
	) name6781 (
		_w2765_,
		_w7242_,
		_w7243_
	);
	LUT2 #(
		.INIT('h2)
	) name6782 (
		_w2742_,
		_w7243_,
		_w7244_
	);
	LUT2 #(
		.INIT('h1)
	) name6783 (
		_w3383_,
		_w7244_,
		_w7245_
	);
	LUT2 #(
		.INIT('h1)
	) name6784 (
		_w2058_,
		_w7245_,
		_w7246_
	);
	LUT2 #(
		.INIT('h8)
	) name6785 (
		_w2058_,
		_w2454_,
		_w7247_
	);
	LUT2 #(
		.INIT('h1)
	) name6786 (
		_w7246_,
		_w7247_,
		_w7248_
	);
	LUT2 #(
		.INIT('h8)
	) name6787 (
		_w3788_,
		_w7248_,
		_w7249_
	);
	LUT2 #(
		.INIT('h1)
	) name6788 (
		_w7241_,
		_w7249_,
		_w7250_
	);
	LUT2 #(
		.INIT('h2)
	) name6789 (
		_w3411_,
		_w7250_,
		_w7251_
	);
	LUT2 #(
		.INIT('h2)
	) name6790 (
		_w2678_,
		_w4198_,
		_w7252_
	);
	LUT2 #(
		.INIT('h4)
	) name6791 (
		_w2678_,
		_w4198_,
		_w7253_
	);
	LUT2 #(
		.INIT('h1)
	) name6792 (
		_w7252_,
		_w7253_,
		_w7254_
	);
	LUT2 #(
		.INIT('h2)
	) name6793 (
		_w3788_,
		_w7254_,
		_w7255_
	);
	LUT2 #(
		.INIT('h1)
	) name6794 (
		_w7241_,
		_w7255_,
		_w7256_
	);
	LUT2 #(
		.INIT('h1)
	) name6795 (
		_w3177_,
		_w7256_,
		_w7257_
	);
	LUT2 #(
		.INIT('h4)
	) name6796 (
		_w2470_,
		_w3332_,
		_w7258_
	);
	LUT2 #(
		.INIT('h2)
	) name6797 (
		_w2779_,
		_w7258_,
		_w7259_
	);
	LUT2 #(
		.INIT('h1)
	) name6798 (
		_w3334_,
		_w7259_,
		_w7260_
	);
	LUT2 #(
		.INIT('h8)
	) name6799 (
		_w3788_,
		_w7260_,
		_w7261_
	);
	LUT2 #(
		.INIT('h1)
	) name6800 (
		_w7241_,
		_w7261_,
		_w7262_
	);
	LUT2 #(
		.INIT('h2)
	) name6801 (
		_w3355_,
		_w7262_,
		_w7263_
	);
	LUT2 #(
		.INIT('h2)
	) name6802 (
		_w3277_,
		_w4198_,
		_w7264_
	);
	LUT2 #(
		.INIT('h4)
	) name6803 (
		_w3277_,
		_w4198_,
		_w7265_
	);
	LUT2 #(
		.INIT('h1)
	) name6804 (
		_w7264_,
		_w7265_,
		_w7266_
	);
	LUT2 #(
		.INIT('h4)
	) name6805 (
		_w3320_,
		_w7266_,
		_w7267_
	);
	LUT2 #(
		.INIT('h8)
	) name6806 (
		_w3788_,
		_w7267_,
		_w7268_
	);
	LUT2 #(
		.INIT('h2)
	) name6807 (
		_w2779_,
		_w3965_,
		_w7269_
	);
	LUT2 #(
		.INIT('h1)
	) name6808 (
		_w7240_,
		_w7269_,
		_w7270_
	);
	LUT2 #(
		.INIT('h4)
	) name6809 (
		_w7268_,
		_w7270_,
		_w7271_
	);
	LUT2 #(
		.INIT('h4)
	) name6810 (
		_w7263_,
		_w7271_,
		_w7272_
	);
	LUT2 #(
		.INIT('h4)
	) name6811 (
		_w7257_,
		_w7272_,
		_w7273_
	);
	LUT2 #(
		.INIT('h4)
	) name6812 (
		_w7251_,
		_w7273_,
		_w7274_
	);
	LUT2 #(
		.INIT('h2)
	) name6813 (
		_w2026_,
		_w7274_,
		_w7275_
	);
	LUT2 #(
		.INIT('h1)
	) name6814 (
		_w7239_,
		_w7275_,
		_w7276_
	);
	LUT2 #(
		.INIT('h2)
	) name6815 (
		\P1_state_reg[0]/NET0131 ,
		_w7276_,
		_w7277_
	);
	LUT2 #(
		.INIT('h8)
	) name6816 (
		_w2760_,
		_w3976_,
		_w7278_
	);
	LUT2 #(
		.INIT('h1)
	) name6817 (
		_w7238_,
		_w7278_,
		_w7279_
	);
	LUT2 #(
		.INIT('h4)
	) name6818 (
		_w7277_,
		_w7279_,
		_w7280_
	);
	LUT2 #(
		.INIT('h2)
	) name6819 (
		\P1_reg3_reg[9]/NET0131 ,
		\P1_state_reg[0]/NET0131 ,
		_w7281_
	);
	LUT2 #(
		.INIT('h8)
	) name6820 (
		_w1239_,
		_w1953_,
		_w7282_
	);
	LUT2 #(
		.INIT('h8)
	) name6821 (
		_w1239_,
		_w3448_,
		_w7283_
	);
	LUT2 #(
		.INIT('h2)
	) name6822 (
		_w1257_,
		_w4067_,
		_w7284_
	);
	LUT2 #(
		.INIT('h2)
	) name6823 (
		_w1239_,
		_w3980_,
		_w7285_
	);
	LUT2 #(
		.INIT('h2)
	) name6824 (
		_w1782_,
		_w3646_,
		_w7286_
	);
	LUT2 #(
		.INIT('h4)
	) name6825 (
		_w1782_,
		_w3646_,
		_w7287_
	);
	LUT2 #(
		.INIT('h1)
	) name6826 (
		_w7286_,
		_w7287_,
		_w7288_
	);
	LUT2 #(
		.INIT('h2)
	) name6827 (
		_w3980_,
		_w7288_,
		_w7289_
	);
	LUT2 #(
		.INIT('h1)
	) name6828 (
		_w7285_,
		_w7289_,
		_w7290_
	);
	LUT2 #(
		.INIT('h1)
	) name6829 (
		_w3677_,
		_w7290_,
		_w7291_
	);
	LUT2 #(
		.INIT('h2)
	) name6830 (
		_w1782_,
		_w3529_,
		_w7292_
	);
	LUT2 #(
		.INIT('h4)
	) name6831 (
		_w1782_,
		_w3529_,
		_w7293_
	);
	LUT2 #(
		.INIT('h1)
	) name6832 (
		_w7292_,
		_w7293_,
		_w7294_
	);
	LUT2 #(
		.INIT('h8)
	) name6833 (
		_w3980_,
		_w7294_,
		_w7295_
	);
	LUT2 #(
		.INIT('h1)
	) name6834 (
		_w7285_,
		_w7295_,
		_w7296_
	);
	LUT2 #(
		.INIT('h1)
	) name6835 (
		_w3563_,
		_w7296_,
		_w7297_
	);
	LUT2 #(
		.INIT('h8)
	) name6836 (
		_w3684_,
		_w3685_,
		_w7298_
	);
	LUT2 #(
		.INIT('h2)
	) name6837 (
		_w1257_,
		_w7298_,
		_w7299_
	);
	LUT2 #(
		.INIT('h1)
	) name6838 (
		_w3687_,
		_w7299_,
		_w7300_
	);
	LUT2 #(
		.INIT('h8)
	) name6839 (
		_w3980_,
		_w7300_,
		_w7301_
	);
	LUT2 #(
		.INIT('h1)
	) name6840 (
		_w7285_,
		_w7301_,
		_w7302_
	);
	LUT2 #(
		.INIT('h2)
	) name6841 (
		_w3712_,
		_w7302_,
		_w7303_
	);
	LUT2 #(
		.INIT('h2)
	) name6842 (
		_w537_,
		_w1267_,
		_w7304_
	);
	LUT2 #(
		.INIT('h4)
	) name6843 (
		_w1267_,
		_w3577_,
		_w7305_
	);
	LUT2 #(
		.INIT('h4)
	) name6844 (
		_w1244_,
		_w7305_,
		_w7306_
	);
	LUT2 #(
		.INIT('h2)
	) name6845 (
		_w1218_,
		_w7306_,
		_w7307_
	);
	LUT2 #(
		.INIT('h1)
	) name6846 (
		_w537_,
		_w3580_,
		_w7308_
	);
	LUT2 #(
		.INIT('h4)
	) name6847 (
		_w7307_,
		_w7308_,
		_w7309_
	);
	LUT2 #(
		.INIT('h1)
	) name6848 (
		_w7304_,
		_w7309_,
		_w7310_
	);
	LUT2 #(
		.INIT('h2)
	) name6849 (
		_w3980_,
		_w7310_,
		_w7311_
	);
	LUT2 #(
		.INIT('h1)
	) name6850 (
		_w7285_,
		_w7311_,
		_w7312_
	);
	LUT2 #(
		.INIT('h2)
	) name6851 (
		_w1936_,
		_w7312_,
		_w7313_
	);
	LUT2 #(
		.INIT('h2)
	) name6852 (
		_w1239_,
		_w4064_,
		_w7314_
	);
	LUT2 #(
		.INIT('h1)
	) name6853 (
		_w7284_,
		_w7314_,
		_w7315_
	);
	LUT2 #(
		.INIT('h4)
	) name6854 (
		_w7303_,
		_w7315_,
		_w7316_
	);
	LUT2 #(
		.INIT('h4)
	) name6855 (
		_w7291_,
		_w7316_,
		_w7317_
	);
	LUT2 #(
		.INIT('h4)
	) name6856 (
		_w7297_,
		_w7317_,
		_w7318_
	);
	LUT2 #(
		.INIT('h4)
	) name6857 (
		_w7313_,
		_w7318_,
		_w7319_
	);
	LUT2 #(
		.INIT('h2)
	) name6858 (
		_w3450_,
		_w7319_,
		_w7320_
	);
	LUT2 #(
		.INIT('h1)
	) name6859 (
		_w7283_,
		_w7320_,
		_w7321_
	);
	LUT2 #(
		.INIT('h2)
	) name6860 (
		\P1_state_reg[0]/NET0131 ,
		_w7321_,
		_w7322_
	);
	LUT2 #(
		.INIT('h1)
	) name6861 (
		_w7281_,
		_w7282_,
		_w7323_
	);
	LUT2 #(
		.INIT('h4)
	) name6862 (
		_w7322_,
		_w7323_,
		_w7324_
	);
	LUT2 #(
		.INIT('h8)
	) name6863 (
		_w2364_,
		_w3976_,
		_w7325_
	);
	LUT2 #(
		.INIT('h4)
	) name6864 (
		\P1_state_reg[0]/NET0131 ,
		\P2_reg3_reg[20]/NET0131 ,
		_w7326_
	);
	LUT2 #(
		.INIT('h8)
	) name6865 (
		_w2024_,
		_w2364_,
		_w7327_
	);
	LUT2 #(
		.INIT('h2)
	) name6866 (
		_w2364_,
		_w3962_,
		_w7328_
	);
	LUT2 #(
		.INIT('h2)
	) name6867 (
		_w2364_,
		_w3788_,
		_w7329_
	);
	LUT2 #(
		.INIT('h8)
	) name6868 (
		_w3788_,
		_w6737_,
		_w7330_
	);
	LUT2 #(
		.INIT('h1)
	) name6869 (
		_w7329_,
		_w7330_,
		_w7331_
	);
	LUT2 #(
		.INIT('h2)
	) name6870 (
		_w3411_,
		_w7331_,
		_w7332_
	);
	LUT2 #(
		.INIT('h2)
	) name6871 (
		_w3788_,
		_w6743_,
		_w7333_
	);
	LUT2 #(
		.INIT('h1)
	) name6872 (
		_w7329_,
		_w7333_,
		_w7334_
	);
	LUT2 #(
		.INIT('h1)
	) name6873 (
		_w3177_,
		_w7334_,
		_w7335_
	);
	LUT2 #(
		.INIT('h2)
	) name6874 (
		_w3788_,
		_w6749_,
		_w7336_
	);
	LUT2 #(
		.INIT('h1)
	) name6875 (
		_w7329_,
		_w7336_,
		_w7337_
	);
	LUT2 #(
		.INIT('h1)
	) name6876 (
		_w3320_,
		_w7337_,
		_w7338_
	);
	LUT2 #(
		.INIT('h8)
	) name6877 (
		_w3788_,
		_w6754_,
		_w7339_
	);
	LUT2 #(
		.INIT('h1)
	) name6878 (
		_w7329_,
		_w7339_,
		_w7340_
	);
	LUT2 #(
		.INIT('h2)
	) name6879 (
		_w3355_,
		_w7340_,
		_w7341_
	);
	LUT2 #(
		.INIT('h2)
	) name6880 (
		_w2358_,
		_w3965_,
		_w7342_
	);
	LUT2 #(
		.INIT('h1)
	) name6881 (
		_w7328_,
		_w7342_,
		_w7343_
	);
	LUT2 #(
		.INIT('h4)
	) name6882 (
		_w7335_,
		_w7343_,
		_w7344_
	);
	LUT2 #(
		.INIT('h1)
	) name6883 (
		_w7338_,
		_w7341_,
		_w7345_
	);
	LUT2 #(
		.INIT('h8)
	) name6884 (
		_w7344_,
		_w7345_,
		_w7346_
	);
	LUT2 #(
		.INIT('h4)
	) name6885 (
		_w7332_,
		_w7346_,
		_w7347_
	);
	LUT2 #(
		.INIT('h2)
	) name6886 (
		_w2026_,
		_w7347_,
		_w7348_
	);
	LUT2 #(
		.INIT('h1)
	) name6887 (
		_w7327_,
		_w7348_,
		_w7349_
	);
	LUT2 #(
		.INIT('h2)
	) name6888 (
		\P1_state_reg[0]/NET0131 ,
		_w7349_,
		_w7350_
	);
	LUT2 #(
		.INIT('h1)
	) name6889 (
		_w7325_,
		_w7326_,
		_w7351_
	);
	LUT2 #(
		.INIT('h4)
	) name6890 (
		_w7350_,
		_w7351_,
		_w7352_
	);
	LUT2 #(
		.INIT('h2)
	) name6891 (
		\P1_reg3_reg[20]/NET0131 ,
		\P1_state_reg[0]/NET0131 ,
		_w7353_
	);
	LUT2 #(
		.INIT('h8)
	) name6892 (
		_w1370_,
		_w1953_,
		_w7354_
	);
	LUT2 #(
		.INIT('h8)
	) name6893 (
		_w1370_,
		_w3448_,
		_w7355_
	);
	LUT2 #(
		.INIT('h2)
	) name6894 (
		_w1370_,
		_w3980_,
		_w7356_
	);
	LUT2 #(
		.INIT('h8)
	) name6895 (
		_w3980_,
		_w6492_,
		_w7357_
	);
	LUT2 #(
		.INIT('h1)
	) name6896 (
		_w7356_,
		_w7357_,
		_w7358_
	);
	LUT2 #(
		.INIT('h2)
	) name6897 (
		_w1936_,
		_w7358_,
		_w7359_
	);
	LUT2 #(
		.INIT('h2)
	) name6898 (
		_w1365_,
		_w4067_,
		_w7360_
	);
	LUT2 #(
		.INIT('h2)
	) name6899 (
		_w3980_,
		_w6505_,
		_w7361_
	);
	LUT2 #(
		.INIT('h1)
	) name6900 (
		_w7356_,
		_w7361_,
		_w7362_
	);
	LUT2 #(
		.INIT('h1)
	) name6901 (
		_w3563_,
		_w7362_,
		_w7363_
	);
	LUT2 #(
		.INIT('h2)
	) name6902 (
		_w3980_,
		_w6499_,
		_w7364_
	);
	LUT2 #(
		.INIT('h1)
	) name6903 (
		_w7356_,
		_w7364_,
		_w7365_
	);
	LUT2 #(
		.INIT('h1)
	) name6904 (
		_w3677_,
		_w7365_,
		_w7366_
	);
	LUT2 #(
		.INIT('h8)
	) name6905 (
		_w3980_,
		_w6510_,
		_w7367_
	);
	LUT2 #(
		.INIT('h1)
	) name6906 (
		_w7356_,
		_w7367_,
		_w7368_
	);
	LUT2 #(
		.INIT('h2)
	) name6907 (
		_w3712_,
		_w7368_,
		_w7369_
	);
	LUT2 #(
		.INIT('h2)
	) name6908 (
		_w1370_,
		_w4064_,
		_w7370_
	);
	LUT2 #(
		.INIT('h1)
	) name6909 (
		_w7360_,
		_w7370_,
		_w7371_
	);
	LUT2 #(
		.INIT('h4)
	) name6910 (
		_w7369_,
		_w7371_,
		_w7372_
	);
	LUT2 #(
		.INIT('h4)
	) name6911 (
		_w7363_,
		_w7372_,
		_w7373_
	);
	LUT2 #(
		.INIT('h4)
	) name6912 (
		_w7366_,
		_w7373_,
		_w7374_
	);
	LUT2 #(
		.INIT('h4)
	) name6913 (
		_w7359_,
		_w7374_,
		_w7375_
	);
	LUT2 #(
		.INIT('h2)
	) name6914 (
		_w3450_,
		_w7375_,
		_w7376_
	);
	LUT2 #(
		.INIT('h1)
	) name6915 (
		_w7355_,
		_w7376_,
		_w7377_
	);
	LUT2 #(
		.INIT('h2)
	) name6916 (
		\P1_state_reg[0]/NET0131 ,
		_w7377_,
		_w7378_
	);
	LUT2 #(
		.INIT('h1)
	) name6917 (
		_w7353_,
		_w7354_,
		_w7379_
	);
	LUT2 #(
		.INIT('h4)
	) name6918 (
		_w7378_,
		_w7379_,
		_w7380_
	);
	LUT2 #(
		.INIT('h8)
	) name6919 (
		_w1352_,
		_w1953_,
		_w7381_
	);
	LUT2 #(
		.INIT('h2)
	) name6920 (
		\P1_reg3_reg[21]/NET0131 ,
		\P1_state_reg[0]/NET0131 ,
		_w7382_
	);
	LUT2 #(
		.INIT('h8)
	) name6921 (
		_w1352_,
		_w3448_,
		_w7383_
	);
	LUT2 #(
		.INIT('h2)
	) name6922 (
		_w1346_,
		_w4067_,
		_w7384_
	);
	LUT2 #(
		.INIT('h2)
	) name6923 (
		_w1352_,
		_w3980_,
		_w7385_
	);
	LUT2 #(
		.INIT('h8)
	) name6924 (
		_w3980_,
		_w6962_,
		_w7386_
	);
	LUT2 #(
		.INIT('h1)
	) name6925 (
		_w7385_,
		_w7386_,
		_w7387_
	);
	LUT2 #(
		.INIT('h2)
	) name6926 (
		_w1936_,
		_w7387_,
		_w7388_
	);
	LUT2 #(
		.INIT('h2)
	) name6927 (
		_w3980_,
		_w6968_,
		_w7389_
	);
	LUT2 #(
		.INIT('h1)
	) name6928 (
		_w7385_,
		_w7389_,
		_w7390_
	);
	LUT2 #(
		.INIT('h1)
	) name6929 (
		_w3563_,
		_w7390_,
		_w7391_
	);
	LUT2 #(
		.INIT('h8)
	) name6930 (
		_w3980_,
		_w6974_,
		_w7392_
	);
	LUT2 #(
		.INIT('h1)
	) name6931 (
		_w7385_,
		_w7392_,
		_w7393_
	);
	LUT2 #(
		.INIT('h1)
	) name6932 (
		_w3677_,
		_w7393_,
		_w7394_
	);
	LUT2 #(
		.INIT('h8)
	) name6933 (
		_w3980_,
		_w6979_,
		_w7395_
	);
	LUT2 #(
		.INIT('h1)
	) name6934 (
		_w7385_,
		_w7395_,
		_w7396_
	);
	LUT2 #(
		.INIT('h2)
	) name6935 (
		_w3712_,
		_w7396_,
		_w7397_
	);
	LUT2 #(
		.INIT('h2)
	) name6936 (
		_w1352_,
		_w4064_,
		_w7398_
	);
	LUT2 #(
		.INIT('h1)
	) name6937 (
		_w7384_,
		_w7398_,
		_w7399_
	);
	LUT2 #(
		.INIT('h4)
	) name6938 (
		_w7397_,
		_w7399_,
		_w7400_
	);
	LUT2 #(
		.INIT('h4)
	) name6939 (
		_w7388_,
		_w7400_,
		_w7401_
	);
	LUT2 #(
		.INIT('h1)
	) name6940 (
		_w7391_,
		_w7394_,
		_w7402_
	);
	LUT2 #(
		.INIT('h8)
	) name6941 (
		_w7401_,
		_w7402_,
		_w7403_
	);
	LUT2 #(
		.INIT('h2)
	) name6942 (
		_w3450_,
		_w7403_,
		_w7404_
	);
	LUT2 #(
		.INIT('h1)
	) name6943 (
		_w7383_,
		_w7404_,
		_w7405_
	);
	LUT2 #(
		.INIT('h2)
	) name6944 (
		\P1_state_reg[0]/NET0131 ,
		_w7405_,
		_w7406_
	);
	LUT2 #(
		.INIT('h1)
	) name6945 (
		_w7381_,
		_w7382_,
		_w7407_
	);
	LUT2 #(
		.INIT('h4)
	) name6946 (
		_w7406_,
		_w7407_,
		_w7408_
	);
	LUT2 #(
		.INIT('h2)
	) name6947 (
		\P1_reg3_reg[23]/NET0131 ,
		\P1_state_reg[0]/NET0131 ,
		_w7409_
	);
	LUT2 #(
		.INIT('h8)
	) name6948 (
		_w1330_,
		_w1953_,
		_w7410_
	);
	LUT2 #(
		.INIT('h8)
	) name6949 (
		_w1330_,
		_w3448_,
		_w7411_
	);
	LUT2 #(
		.INIT('h2)
	) name6950 (
		_w1330_,
		_w3980_,
		_w7412_
	);
	LUT2 #(
		.INIT('h4)
	) name6951 (
		_w4404_,
		_w4406_,
		_w7413_
	);
	LUT2 #(
		.INIT('h2)
	) name6952 (
		_w4410_,
		_w7413_,
		_w7414_
	);
	LUT2 #(
		.INIT('h8)
	) name6953 (
		_w4405_,
		_w4417_,
		_w7415_
	);
	LUT2 #(
		.INIT('h4)
	) name6954 (
		_w7414_,
		_w7415_,
		_w7416_
	);
	LUT2 #(
		.INIT('h4)
	) name6955 (
		_w4413_,
		_w4417_,
		_w7417_
	);
	LUT2 #(
		.INIT('h2)
	) name6956 (
		_w4422_,
		_w7417_,
		_w7418_
	);
	LUT2 #(
		.INIT('h4)
	) name6957 (
		_w7416_,
		_w7418_,
		_w7419_
	);
	LUT2 #(
		.INIT('h2)
	) name6958 (
		_w1821_,
		_w7419_,
		_w7420_
	);
	LUT2 #(
		.INIT('h4)
	) name6959 (
		_w1821_,
		_w7419_,
		_w7421_
	);
	LUT2 #(
		.INIT('h1)
	) name6960 (
		_w7420_,
		_w7421_,
		_w7422_
	);
	LUT2 #(
		.INIT('h2)
	) name6961 (
		_w3980_,
		_w7422_,
		_w7423_
	);
	LUT2 #(
		.INIT('h1)
	) name6962 (
		_w7412_,
		_w7423_,
		_w7424_
	);
	LUT2 #(
		.INIT('h1)
	) name6963 (
		_w3677_,
		_w7424_,
		_w7425_
	);
	LUT2 #(
		.INIT('h4)
	) name6964 (
		_w4447_,
		_w4448_,
		_w7426_
	);
	LUT2 #(
		.INIT('h2)
	) name6965 (
		_w4453_,
		_w7426_,
		_w7427_
	);
	LUT2 #(
		.INIT('h8)
	) name6966 (
		_w4449_,
		_w4459_,
		_w7428_
	);
	LUT2 #(
		.INIT('h4)
	) name6967 (
		_w7427_,
		_w7428_,
		_w7429_
	);
	LUT2 #(
		.INIT('h4)
	) name6968 (
		_w4456_,
		_w4459_,
		_w7430_
	);
	LUT2 #(
		.INIT('h2)
	) name6969 (
		_w4435_,
		_w7430_,
		_w7431_
	);
	LUT2 #(
		.INIT('h4)
	) name6970 (
		_w7429_,
		_w7431_,
		_w7432_
	);
	LUT2 #(
		.INIT('h8)
	) name6971 (
		_w1821_,
		_w7432_,
		_w7433_
	);
	LUT2 #(
		.INIT('h1)
	) name6972 (
		_w1821_,
		_w7432_,
		_w7434_
	);
	LUT2 #(
		.INIT('h1)
	) name6973 (
		_w7433_,
		_w7434_,
		_w7435_
	);
	LUT2 #(
		.INIT('h2)
	) name6974 (
		_w3980_,
		_w7435_,
		_w7436_
	);
	LUT2 #(
		.INIT('h1)
	) name6975 (
		_w7412_,
		_w7436_,
		_w7437_
	);
	LUT2 #(
		.INIT('h1)
	) name6976 (
		_w3563_,
		_w7437_,
		_w7438_
	);
	LUT2 #(
		.INIT('h2)
	) name6977 (
		_w1330_,
		_w4910_,
		_w7439_
	);
	LUT2 #(
		.INIT('h2)
	) name6978 (
		_w1062_,
		_w4472_,
		_w7440_
	);
	LUT2 #(
		.INIT('h1)
	) name6979 (
		_w4075_,
		_w7440_,
		_w7441_
	);
	LUT2 #(
		.INIT('h1)
	) name6980 (
		_w537_,
		_w7441_,
		_w7442_
	);
	LUT2 #(
		.INIT('h8)
	) name6981 (
		_w537_,
		_w1318_,
		_w7443_
	);
	LUT2 #(
		.INIT('h1)
	) name6982 (
		_w7442_,
		_w7443_,
		_w7444_
	);
	LUT2 #(
		.INIT('h8)
	) name6983 (
		_w3980_,
		_w7444_,
		_w7445_
	);
	LUT2 #(
		.INIT('h1)
	) name6984 (
		_w7412_,
		_w7445_,
		_w7446_
	);
	LUT2 #(
		.INIT('h2)
	) name6985 (
		_w1936_,
		_w7446_,
		_w7447_
	);
	LUT2 #(
		.INIT('h2)
	) name6986 (
		_w1327_,
		_w3700_,
		_w7448_
	);
	LUT2 #(
		.INIT('h1)
	) name6987 (
		_w5188_,
		_w7448_,
		_w7449_
	);
	LUT2 #(
		.INIT('h8)
	) name6988 (
		_w3712_,
		_w7449_,
		_w7450_
	);
	LUT2 #(
		.INIT('h8)
	) name6989 (
		_w3980_,
		_w7450_,
		_w7451_
	);
	LUT2 #(
		.INIT('h2)
	) name6990 (
		_w1327_,
		_w4067_,
		_w7452_
	);
	LUT2 #(
		.INIT('h1)
	) name6991 (
		_w7439_,
		_w7452_,
		_w7453_
	);
	LUT2 #(
		.INIT('h4)
	) name6992 (
		_w7451_,
		_w7453_,
		_w7454_
	);
	LUT2 #(
		.INIT('h4)
	) name6993 (
		_w7447_,
		_w7454_,
		_w7455_
	);
	LUT2 #(
		.INIT('h4)
	) name6994 (
		_w7425_,
		_w7455_,
		_w7456_
	);
	LUT2 #(
		.INIT('h4)
	) name6995 (
		_w7438_,
		_w7456_,
		_w7457_
	);
	LUT2 #(
		.INIT('h2)
	) name6996 (
		_w3450_,
		_w7457_,
		_w7458_
	);
	LUT2 #(
		.INIT('h1)
	) name6997 (
		_w7411_,
		_w7458_,
		_w7459_
	);
	LUT2 #(
		.INIT('h2)
	) name6998 (
		\P1_state_reg[0]/NET0131 ,
		_w7459_,
		_w7460_
	);
	LUT2 #(
		.INIT('h1)
	) name6999 (
		_w7409_,
		_w7410_,
		_w7461_
	);
	LUT2 #(
		.INIT('h4)
	) name7000 (
		_w7460_,
		_w7461_,
		_w7462_
	);
	LUT2 #(
		.INIT('h2)
	) name7001 (
		\P2_reg0_reg[20]/NET0131 ,
		_w1983_,
		_w7463_
	);
	LUT2 #(
		.INIT('h8)
	) name7002 (
		\P2_reg0_reg[20]/NET0131 ,
		_w2024_,
		_w7464_
	);
	LUT2 #(
		.INIT('h2)
	) name7003 (
		\P2_reg0_reg[20]/NET0131 ,
		_w3423_,
		_w7465_
	);
	LUT2 #(
		.INIT('h2)
	) name7004 (
		\P2_reg0_reg[20]/NET0131 ,
		_w2040_,
		_w7466_
	);
	LUT2 #(
		.INIT('h8)
	) name7005 (
		_w2040_,
		_w6737_,
		_w7467_
	);
	LUT2 #(
		.INIT('h1)
	) name7006 (
		_w7466_,
		_w7467_,
		_w7468_
	);
	LUT2 #(
		.INIT('h2)
	) name7007 (
		_w3411_,
		_w7468_,
		_w7469_
	);
	LUT2 #(
		.INIT('h2)
	) name7008 (
		_w2040_,
		_w6743_,
		_w7470_
	);
	LUT2 #(
		.INIT('h1)
	) name7009 (
		_w7466_,
		_w7470_,
		_w7471_
	);
	LUT2 #(
		.INIT('h1)
	) name7010 (
		_w3177_,
		_w7471_,
		_w7472_
	);
	LUT2 #(
		.INIT('h2)
	) name7011 (
		_w2040_,
		_w6749_,
		_w7473_
	);
	LUT2 #(
		.INIT('h1)
	) name7012 (
		_w7466_,
		_w7473_,
		_w7474_
	);
	LUT2 #(
		.INIT('h1)
	) name7013 (
		_w3320_,
		_w7474_,
		_w7475_
	);
	LUT2 #(
		.INIT('h8)
	) name7014 (
		_w2040_,
		_w6754_,
		_w7476_
	);
	LUT2 #(
		.INIT('h1)
	) name7015 (
		_w7466_,
		_w7476_,
		_w7477_
	);
	LUT2 #(
		.INIT('h2)
	) name7016 (
		_w3355_,
		_w7477_,
		_w7478_
	);
	LUT2 #(
		.INIT('h8)
	) name7017 (
		_w2040_,
		_w6759_,
		_w7479_
	);
	LUT2 #(
		.INIT('h1)
	) name7018 (
		_w7465_,
		_w7479_,
		_w7480_
	);
	LUT2 #(
		.INIT('h4)
	) name7019 (
		_w7472_,
		_w7480_,
		_w7481_
	);
	LUT2 #(
		.INIT('h1)
	) name7020 (
		_w7475_,
		_w7478_,
		_w7482_
	);
	LUT2 #(
		.INIT('h8)
	) name7021 (
		_w7481_,
		_w7482_,
		_w7483_
	);
	LUT2 #(
		.INIT('h4)
	) name7022 (
		_w7469_,
		_w7483_,
		_w7484_
	);
	LUT2 #(
		.INIT('h2)
	) name7023 (
		_w2026_,
		_w7484_,
		_w7485_
	);
	LUT2 #(
		.INIT('h1)
	) name7024 (
		_w7464_,
		_w7485_,
		_w7486_
	);
	LUT2 #(
		.INIT('h2)
	) name7025 (
		\P1_state_reg[0]/NET0131 ,
		_w7486_,
		_w7487_
	);
	LUT2 #(
		.INIT('h1)
	) name7026 (
		_w7463_,
		_w7487_,
		_w7488_
	);
	LUT2 #(
		.INIT('h8)
	) name7027 (
		_w825_,
		_w1880_,
		_w7489_
	);
	LUT2 #(
		.INIT('h1)
	) name7028 (
		_w5802_,
		_w7489_,
		_w7490_
	);
	LUT2 #(
		.INIT('h2)
	) name7029 (
		_w825_,
		_w3708_,
		_w7491_
	);
	LUT2 #(
		.INIT('h1)
	) name7030 (
		_w5803_,
		_w7491_,
		_w7492_
	);
	LUT2 #(
		.INIT('h8)
	) name7031 (
		_w3712_,
		_w7492_,
		_w7493_
	);
	LUT2 #(
		.INIT('h2)
	) name7032 (
		_w7490_,
		_w7493_,
		_w7494_
	);
	LUT2 #(
		.INIT('h2)
	) name7033 (
		_w4532_,
		_w7494_,
		_w7495_
	);
	LUT2 #(
		.INIT('h2)
	) name7034 (
		\P1_reg1_reg[30]/NET0131 ,
		_w6945_,
		_w7496_
	);
	LUT2 #(
		.INIT('h1)
	) name7035 (
		_w7495_,
		_w7496_,
		_w7497_
	);
	LUT2 #(
		.INIT('h2)
	) name7036 (
		_w3450_,
		_w7497_,
		_w7498_
	);
	LUT2 #(
		.INIT('h8)
	) name7037 (
		\P1_reg1_reg[30]/NET0131 ,
		_w3448_,
		_w7499_
	);
	LUT2 #(
		.INIT('h1)
	) name7038 (
		_w7498_,
		_w7499_,
		_w7500_
	);
	LUT2 #(
		.INIT('h2)
	) name7039 (
		\P1_state_reg[0]/NET0131 ,
		_w7500_,
		_w7501_
	);
	LUT2 #(
		.INIT('h2)
	) name7040 (
		\P1_reg1_reg[30]/NET0131 ,
		_w3435_,
		_w7502_
	);
	LUT2 #(
		.INIT('h1)
	) name7041 (
		_w7501_,
		_w7502_,
		_w7503_
	);
	LUT2 #(
		.INIT('h2)
	) name7042 (
		_w5860_,
		_w6648_,
		_w7504_
	);
	LUT2 #(
		.INIT('h1)
	) name7043 (
		_w2040_,
		_w6639_,
		_w7505_
	);
	LUT2 #(
		.INIT('h2)
	) name7044 (
		_w3421_,
		_w7505_,
		_w7506_
	);
	LUT2 #(
		.INIT('h4)
	) name7045 (
		_w2040_,
		_w3354_,
		_w7507_
	);
	LUT2 #(
		.INIT('h4)
	) name7046 (
		_w3171_,
		_w4308_,
		_w7508_
	);
	LUT2 #(
		.INIT('h1)
	) name7047 (
		_w2040_,
		_w7508_,
		_w7509_
	);
	LUT2 #(
		.INIT('h2)
	) name7048 (
		_w5287_,
		_w7509_,
		_w7510_
	);
	LUT2 #(
		.INIT('h2)
	) name7049 (
		_w7506_,
		_w7507_,
		_w7511_
	);
	LUT2 #(
		.INIT('h8)
	) name7050 (
		_w7510_,
		_w7511_,
		_w7512_
	);
	LUT2 #(
		.INIT('h2)
	) name7051 (
		\P2_reg0_reg[21]/NET0131 ,
		_w7512_,
		_w7513_
	);
	LUT2 #(
		.INIT('h1)
	) name7052 (
		_w7504_,
		_w7513_,
		_w7514_
	);
	LUT2 #(
		.INIT('h2)
	) name7053 (
		\P1_reg2_reg[12]/NET0131 ,
		_w3435_,
		_w7515_
	);
	LUT2 #(
		.INIT('h8)
	) name7054 (
		\P1_reg2_reg[12]/NET0131 ,
		_w3448_,
		_w7516_
	);
	LUT2 #(
		.INIT('h2)
	) name7055 (
		\P1_reg2_reg[12]/NET0131 ,
		_w3718_,
		_w7517_
	);
	LUT2 #(
		.INIT('h2)
	) name7056 (
		\P1_reg2_reg[12]/NET0131 ,
		_w3466_,
		_w7518_
	);
	LUT2 #(
		.INIT('h8)
	) name7057 (
		_w3466_,
		_w6098_,
		_w7519_
	);
	LUT2 #(
		.INIT('h1)
	) name7058 (
		_w7518_,
		_w7519_,
		_w7520_
	);
	LUT2 #(
		.INIT('h2)
	) name7059 (
		_w1936_,
		_w7520_,
		_w7521_
	);
	LUT2 #(
		.INIT('h8)
	) name7060 (
		_w3466_,
		_w6104_,
		_w7522_
	);
	LUT2 #(
		.INIT('h1)
	) name7061 (
		_w7518_,
		_w7522_,
		_w7523_
	);
	LUT2 #(
		.INIT('h1)
	) name7062 (
		_w3563_,
		_w7523_,
		_w7524_
	);
	LUT2 #(
		.INIT('h2)
	) name7063 (
		_w3466_,
		_w6110_,
		_w7525_
	);
	LUT2 #(
		.INIT('h1)
	) name7064 (
		_w7518_,
		_w7525_,
		_w7526_
	);
	LUT2 #(
		.INIT('h1)
	) name7065 (
		_w3677_,
		_w7526_,
		_w7527_
	);
	LUT2 #(
		.INIT('h8)
	) name7066 (
		_w3466_,
		_w6117_,
		_w7528_
	);
	LUT2 #(
		.INIT('h1)
	) name7067 (
		_w7518_,
		_w7528_,
		_w7529_
	);
	LUT2 #(
		.INIT('h2)
	) name7068 (
		_w3712_,
		_w7529_,
		_w7530_
	);
	LUT2 #(
		.INIT('h8)
	) name7069 (
		_w1170_,
		_w1763_,
		_w7531_
	);
	LUT2 #(
		.INIT('h8)
	) name7070 (
		_w1165_,
		_w1880_,
		_w7532_
	);
	LUT2 #(
		.INIT('h8)
	) name7071 (
		_w3466_,
		_w7532_,
		_w7533_
	);
	LUT2 #(
		.INIT('h1)
	) name7072 (
		_w7531_,
		_w7533_,
		_w7534_
	);
	LUT2 #(
		.INIT('h4)
	) name7073 (
		_w7517_,
		_w7534_,
		_w7535_
	);
	LUT2 #(
		.INIT('h4)
	) name7074 (
		_w7530_,
		_w7535_,
		_w7536_
	);
	LUT2 #(
		.INIT('h4)
	) name7075 (
		_w7524_,
		_w7536_,
		_w7537_
	);
	LUT2 #(
		.INIT('h4)
	) name7076 (
		_w7527_,
		_w7537_,
		_w7538_
	);
	LUT2 #(
		.INIT('h4)
	) name7077 (
		_w7521_,
		_w7538_,
		_w7539_
	);
	LUT2 #(
		.INIT('h2)
	) name7078 (
		_w3450_,
		_w7539_,
		_w7540_
	);
	LUT2 #(
		.INIT('h1)
	) name7079 (
		_w7516_,
		_w7540_,
		_w7541_
	);
	LUT2 #(
		.INIT('h2)
	) name7080 (
		\P1_state_reg[0]/NET0131 ,
		_w7541_,
		_w7542_
	);
	LUT2 #(
		.INIT('h1)
	) name7081 (
		_w7515_,
		_w7542_,
		_w7543_
	);
	LUT2 #(
		.INIT('h2)
	) name7082 (
		\P2_reg0_reg[30]/NET0131 ,
		_w5861_,
		_w7544_
	);
	LUT2 #(
		.INIT('h8)
	) name7083 (
		_w3358_,
		_w4159_,
		_w7545_
	);
	LUT2 #(
		.INIT('h1)
	) name7084 (
		_w5277_,
		_w7545_,
		_w7546_
	);
	LUT2 #(
		.INIT('h4)
	) name7085 (
		_w3350_,
		_w4159_,
		_w7547_
	);
	LUT2 #(
		.INIT('h1)
	) name7086 (
		_w5279_,
		_w7547_,
		_w7548_
	);
	LUT2 #(
		.INIT('h8)
	) name7087 (
		_w3355_,
		_w7548_,
		_w7549_
	);
	LUT2 #(
		.INIT('h2)
	) name7088 (
		_w7546_,
		_w7549_,
		_w7550_
	);
	LUT2 #(
		.INIT('h2)
	) name7089 (
		_w5860_,
		_w7550_,
		_w7551_
	);
	LUT2 #(
		.INIT('h1)
	) name7090 (
		_w7544_,
		_w7551_,
		_w7552_
	);
	LUT2 #(
		.INIT('h2)
	) name7091 (
		\P1_reg2_reg[16]/NET0131 ,
		_w3435_,
		_w7553_
	);
	LUT2 #(
		.INIT('h8)
	) name7092 (
		\P1_reg2_reg[16]/NET0131 ,
		_w3448_,
		_w7554_
	);
	LUT2 #(
		.INIT('h2)
	) name7093 (
		\P1_reg2_reg[16]/NET0131 ,
		_w3718_,
		_w7555_
	);
	LUT2 #(
		.INIT('h2)
	) name7094 (
		\P1_reg2_reg[16]/NET0131 ,
		_w3466_,
		_w7556_
	);
	LUT2 #(
		.INIT('h2)
	) name7095 (
		_w3466_,
		_w6141_,
		_w7557_
	);
	LUT2 #(
		.INIT('h1)
	) name7096 (
		_w7556_,
		_w7557_,
		_w7558_
	);
	LUT2 #(
		.INIT('h1)
	) name7097 (
		_w3563_,
		_w7558_,
		_w7559_
	);
	LUT2 #(
		.INIT('h8)
	) name7098 (
		_w3466_,
		_w6149_,
		_w7560_
	);
	LUT2 #(
		.INIT('h1)
	) name7099 (
		_w7556_,
		_w7560_,
		_w7561_
	);
	LUT2 #(
		.INIT('h2)
	) name7100 (
		_w1936_,
		_w7561_,
		_w7562_
	);
	LUT2 #(
		.INIT('h8)
	) name7101 (
		_w3466_,
		_w6160_,
		_w7563_
	);
	LUT2 #(
		.INIT('h1)
	) name7102 (
		_w7556_,
		_w7563_,
		_w7564_
	);
	LUT2 #(
		.INIT('h2)
	) name7103 (
		_w3712_,
		_w7564_,
		_w7565_
	);
	LUT2 #(
		.INIT('h2)
	) name7104 (
		_w3466_,
		_w6155_,
		_w7566_
	);
	LUT2 #(
		.INIT('h1)
	) name7105 (
		_w7556_,
		_w7566_,
		_w7567_
	);
	LUT2 #(
		.INIT('h1)
	) name7106 (
		_w3677_,
		_w7567_,
		_w7568_
	);
	LUT2 #(
		.INIT('h8)
	) name7107 (
		_w1471_,
		_w1763_,
		_w7569_
	);
	LUT2 #(
		.INIT('h8)
	) name7108 (
		_w1466_,
		_w1880_,
		_w7570_
	);
	LUT2 #(
		.INIT('h8)
	) name7109 (
		_w3466_,
		_w7570_,
		_w7571_
	);
	LUT2 #(
		.INIT('h1)
	) name7110 (
		_w7555_,
		_w7569_,
		_w7572_
	);
	LUT2 #(
		.INIT('h4)
	) name7111 (
		_w7571_,
		_w7572_,
		_w7573_
	);
	LUT2 #(
		.INIT('h4)
	) name7112 (
		_w7565_,
		_w7573_,
		_w7574_
	);
	LUT2 #(
		.INIT('h4)
	) name7113 (
		_w7568_,
		_w7574_,
		_w7575_
	);
	LUT2 #(
		.INIT('h4)
	) name7114 (
		_w7559_,
		_w7575_,
		_w7576_
	);
	LUT2 #(
		.INIT('h4)
	) name7115 (
		_w7562_,
		_w7576_,
		_w7577_
	);
	LUT2 #(
		.INIT('h2)
	) name7116 (
		_w3450_,
		_w7577_,
		_w7578_
	);
	LUT2 #(
		.INIT('h1)
	) name7117 (
		_w7554_,
		_w7578_,
		_w7579_
	);
	LUT2 #(
		.INIT('h2)
	) name7118 (
		\P1_state_reg[0]/NET0131 ,
		_w7579_,
		_w7580_
	);
	LUT2 #(
		.INIT('h1)
	) name7119 (
		_w7553_,
		_w7580_,
		_w7581_
	);
	LUT2 #(
		.INIT('h2)
	) name7120 (
		\P2_reg1_reg[12]/NET0131 ,
		_w1983_,
		_w7582_
	);
	LUT2 #(
		.INIT('h8)
	) name7121 (
		\P2_reg1_reg[12]/NET0131 ,
		_w2024_,
		_w7583_
	);
	LUT2 #(
		.INIT('h8)
	) name7122 (
		_w2731_,
		_w3358_,
		_w7584_
	);
	LUT2 #(
		.INIT('h1)
	) name7123 (
		_w6204_,
		_w7584_,
		_w7585_
	);
	LUT2 #(
		.INIT('h2)
	) name7124 (
		_w3733_,
		_w7585_,
		_w7586_
	);
	LUT2 #(
		.INIT('h2)
	) name7125 (
		\P2_reg1_reg[12]/NET0131 ,
		_w3733_,
		_w7587_
	);
	LUT2 #(
		.INIT('h8)
	) name7126 (
		_w3733_,
		_w6186_,
		_w7588_
	);
	LUT2 #(
		.INIT('h1)
	) name7127 (
		_w7587_,
		_w7588_,
		_w7589_
	);
	LUT2 #(
		.INIT('h2)
	) name7128 (
		_w3411_,
		_w7589_,
		_w7590_
	);
	LUT2 #(
		.INIT('h8)
	) name7129 (
		_w3733_,
		_w6192_,
		_w7591_
	);
	LUT2 #(
		.INIT('h1)
	) name7130 (
		_w7587_,
		_w7591_,
		_w7592_
	);
	LUT2 #(
		.INIT('h1)
	) name7131 (
		_w3177_,
		_w7592_,
		_w7593_
	);
	LUT2 #(
		.INIT('h2)
	) name7132 (
		_w3733_,
		_w6198_,
		_w7594_
	);
	LUT2 #(
		.INIT('h1)
	) name7133 (
		_w7587_,
		_w7594_,
		_w7595_
	);
	LUT2 #(
		.INIT('h1)
	) name7134 (
		_w3320_,
		_w7595_,
		_w7596_
	);
	LUT2 #(
		.INIT('h2)
	) name7135 (
		_w3355_,
		_w3733_,
		_w7597_
	);
	LUT2 #(
		.INIT('h2)
	) name7136 (
		_w3743_,
		_w7597_,
		_w7598_
	);
	LUT2 #(
		.INIT('h2)
	) name7137 (
		\P2_reg1_reg[12]/NET0131 ,
		_w7598_,
		_w7599_
	);
	LUT2 #(
		.INIT('h1)
	) name7138 (
		_w7586_,
		_w7599_,
		_w7600_
	);
	LUT2 #(
		.INIT('h4)
	) name7139 (
		_w7593_,
		_w7600_,
		_w7601_
	);
	LUT2 #(
		.INIT('h4)
	) name7140 (
		_w7596_,
		_w7601_,
		_w7602_
	);
	LUT2 #(
		.INIT('h4)
	) name7141 (
		_w7590_,
		_w7602_,
		_w7603_
	);
	LUT2 #(
		.INIT('h2)
	) name7142 (
		_w2026_,
		_w7603_,
		_w7604_
	);
	LUT2 #(
		.INIT('h1)
	) name7143 (
		_w7583_,
		_w7604_,
		_w7605_
	);
	LUT2 #(
		.INIT('h2)
	) name7144 (
		\P1_state_reg[0]/NET0131 ,
		_w7605_,
		_w7606_
	);
	LUT2 #(
		.INIT('h1)
	) name7145 (
		_w7582_,
		_w7606_,
		_w7607_
	);
	LUT2 #(
		.INIT('h2)
	) name7146 (
		\P1_reg2_reg[21]/NET0131 ,
		_w3435_,
		_w7608_
	);
	LUT2 #(
		.INIT('h8)
	) name7147 (
		\P1_reg2_reg[21]/NET0131 ,
		_w3448_,
		_w7609_
	);
	LUT2 #(
		.INIT('h2)
	) name7148 (
		\P1_reg2_reg[21]/NET0131 ,
		_w3718_,
		_w7610_
	);
	LUT2 #(
		.INIT('h2)
	) name7149 (
		\P1_reg2_reg[21]/NET0131 ,
		_w3466_,
		_w7611_
	);
	LUT2 #(
		.INIT('h8)
	) name7150 (
		_w3466_,
		_w6962_,
		_w7612_
	);
	LUT2 #(
		.INIT('h1)
	) name7151 (
		_w7611_,
		_w7612_,
		_w7613_
	);
	LUT2 #(
		.INIT('h2)
	) name7152 (
		_w1936_,
		_w7613_,
		_w7614_
	);
	LUT2 #(
		.INIT('h2)
	) name7153 (
		_w3466_,
		_w6968_,
		_w7615_
	);
	LUT2 #(
		.INIT('h1)
	) name7154 (
		_w7611_,
		_w7615_,
		_w7616_
	);
	LUT2 #(
		.INIT('h1)
	) name7155 (
		_w3563_,
		_w7616_,
		_w7617_
	);
	LUT2 #(
		.INIT('h8)
	) name7156 (
		_w3466_,
		_w6974_,
		_w7618_
	);
	LUT2 #(
		.INIT('h1)
	) name7157 (
		_w7611_,
		_w7618_,
		_w7619_
	);
	LUT2 #(
		.INIT('h1)
	) name7158 (
		_w3677_,
		_w7619_,
		_w7620_
	);
	LUT2 #(
		.INIT('h8)
	) name7159 (
		_w3466_,
		_w6979_,
		_w7621_
	);
	LUT2 #(
		.INIT('h1)
	) name7160 (
		_w7611_,
		_w7621_,
		_w7622_
	);
	LUT2 #(
		.INIT('h2)
	) name7161 (
		_w3712_,
		_w7622_,
		_w7623_
	);
	LUT2 #(
		.INIT('h8)
	) name7162 (
		_w1352_,
		_w1763_,
		_w7624_
	);
	LUT2 #(
		.INIT('h8)
	) name7163 (
		_w3466_,
		_w6955_,
		_w7625_
	);
	LUT2 #(
		.INIT('h1)
	) name7164 (
		_w7610_,
		_w7624_,
		_w7626_
	);
	LUT2 #(
		.INIT('h4)
	) name7165 (
		_w7625_,
		_w7626_,
		_w7627_
	);
	LUT2 #(
		.INIT('h4)
	) name7166 (
		_w7623_,
		_w7627_,
		_w7628_
	);
	LUT2 #(
		.INIT('h4)
	) name7167 (
		_w7614_,
		_w7628_,
		_w7629_
	);
	LUT2 #(
		.INIT('h1)
	) name7168 (
		_w7617_,
		_w7620_,
		_w7630_
	);
	LUT2 #(
		.INIT('h8)
	) name7169 (
		_w7629_,
		_w7630_,
		_w7631_
	);
	LUT2 #(
		.INIT('h2)
	) name7170 (
		_w3450_,
		_w7631_,
		_w7632_
	);
	LUT2 #(
		.INIT('h1)
	) name7171 (
		_w7609_,
		_w7632_,
		_w7633_
	);
	LUT2 #(
		.INIT('h2)
	) name7172 (
		\P1_state_reg[0]/NET0131 ,
		_w7633_,
		_w7634_
	);
	LUT2 #(
		.INIT('h1)
	) name7173 (
		_w7608_,
		_w7634_,
		_w7635_
	);
	LUT2 #(
		.INIT('h2)
	) name7174 (
		\P1_reg2_reg[23]/NET0131 ,
		_w3435_,
		_w7636_
	);
	LUT2 #(
		.INIT('h8)
	) name7175 (
		\P1_reg2_reg[23]/NET0131 ,
		_w3448_,
		_w7637_
	);
	LUT2 #(
		.INIT('h2)
	) name7176 (
		\P1_reg2_reg[23]/NET0131 ,
		_w3466_,
		_w7638_
	);
	LUT2 #(
		.INIT('h2)
	) name7177 (
		_w3466_,
		_w7422_,
		_w7639_
	);
	LUT2 #(
		.INIT('h1)
	) name7178 (
		_w7638_,
		_w7639_,
		_w7640_
	);
	LUT2 #(
		.INIT('h1)
	) name7179 (
		_w3677_,
		_w7640_,
		_w7641_
	);
	LUT2 #(
		.INIT('h2)
	) name7180 (
		_w3466_,
		_w7435_,
		_w7642_
	);
	LUT2 #(
		.INIT('h1)
	) name7181 (
		_w7638_,
		_w7642_,
		_w7643_
	);
	LUT2 #(
		.INIT('h1)
	) name7182 (
		_w3563_,
		_w7643_,
		_w7644_
	);
	LUT2 #(
		.INIT('h2)
	) name7183 (
		\P1_reg2_reg[23]/NET0131 ,
		_w3718_,
		_w7645_
	);
	LUT2 #(
		.INIT('h8)
	) name7184 (
		_w3466_,
		_w7444_,
		_w7646_
	);
	LUT2 #(
		.INIT('h1)
	) name7185 (
		_w7638_,
		_w7646_,
		_w7647_
	);
	LUT2 #(
		.INIT('h2)
	) name7186 (
		_w1936_,
		_w7647_,
		_w7648_
	);
	LUT2 #(
		.INIT('h8)
	) name7187 (
		_w3466_,
		_w7449_,
		_w7649_
	);
	LUT2 #(
		.INIT('h1)
	) name7188 (
		_w7638_,
		_w7649_,
		_w7650_
	);
	LUT2 #(
		.INIT('h2)
	) name7189 (
		_w3712_,
		_w7650_,
		_w7651_
	);
	LUT2 #(
		.INIT('h8)
	) name7190 (
		_w1330_,
		_w1763_,
		_w7652_
	);
	LUT2 #(
		.INIT('h8)
	) name7191 (
		_w1327_,
		_w1880_,
		_w7653_
	);
	LUT2 #(
		.INIT('h8)
	) name7192 (
		_w3466_,
		_w7653_,
		_w7654_
	);
	LUT2 #(
		.INIT('h1)
	) name7193 (
		_w7645_,
		_w7652_,
		_w7655_
	);
	LUT2 #(
		.INIT('h4)
	) name7194 (
		_w7654_,
		_w7655_,
		_w7656_
	);
	LUT2 #(
		.INIT('h4)
	) name7195 (
		_w7651_,
		_w7656_,
		_w7657_
	);
	LUT2 #(
		.INIT('h4)
	) name7196 (
		_w7648_,
		_w7657_,
		_w7658_
	);
	LUT2 #(
		.INIT('h4)
	) name7197 (
		_w7641_,
		_w7658_,
		_w7659_
	);
	LUT2 #(
		.INIT('h4)
	) name7198 (
		_w7644_,
		_w7659_,
		_w7660_
	);
	LUT2 #(
		.INIT('h2)
	) name7199 (
		_w3450_,
		_w7660_,
		_w7661_
	);
	LUT2 #(
		.INIT('h1)
	) name7200 (
		_w7637_,
		_w7661_,
		_w7662_
	);
	LUT2 #(
		.INIT('h2)
	) name7201 (
		\P1_state_reg[0]/NET0131 ,
		_w7662_,
		_w7663_
	);
	LUT2 #(
		.INIT('h1)
	) name7202 (
		_w7636_,
		_w7663_,
		_w7664_
	);
	LUT2 #(
		.INIT('h2)
	) name7203 (
		\P2_reg1_reg[20]/NET0131 ,
		_w1983_,
		_w7665_
	);
	LUT2 #(
		.INIT('h8)
	) name7204 (
		\P2_reg1_reg[20]/NET0131 ,
		_w2024_,
		_w7666_
	);
	LUT2 #(
		.INIT('h2)
	) name7205 (
		\P2_reg1_reg[20]/NET0131 ,
		_w3743_,
		_w7667_
	);
	LUT2 #(
		.INIT('h2)
	) name7206 (
		\P2_reg1_reg[20]/NET0131 ,
		_w3733_,
		_w7668_
	);
	LUT2 #(
		.INIT('h8)
	) name7207 (
		_w3733_,
		_w6737_,
		_w7669_
	);
	LUT2 #(
		.INIT('h1)
	) name7208 (
		_w7668_,
		_w7669_,
		_w7670_
	);
	LUT2 #(
		.INIT('h2)
	) name7209 (
		_w3411_,
		_w7670_,
		_w7671_
	);
	LUT2 #(
		.INIT('h2)
	) name7210 (
		_w3733_,
		_w6743_,
		_w7672_
	);
	LUT2 #(
		.INIT('h1)
	) name7211 (
		_w7668_,
		_w7672_,
		_w7673_
	);
	LUT2 #(
		.INIT('h1)
	) name7212 (
		_w3177_,
		_w7673_,
		_w7674_
	);
	LUT2 #(
		.INIT('h2)
	) name7213 (
		_w3733_,
		_w6749_,
		_w7675_
	);
	LUT2 #(
		.INIT('h1)
	) name7214 (
		_w7668_,
		_w7675_,
		_w7676_
	);
	LUT2 #(
		.INIT('h1)
	) name7215 (
		_w3320_,
		_w7676_,
		_w7677_
	);
	LUT2 #(
		.INIT('h8)
	) name7216 (
		_w3733_,
		_w6754_,
		_w7678_
	);
	LUT2 #(
		.INIT('h1)
	) name7217 (
		_w7668_,
		_w7678_,
		_w7679_
	);
	LUT2 #(
		.INIT('h2)
	) name7218 (
		_w3355_,
		_w7679_,
		_w7680_
	);
	LUT2 #(
		.INIT('h8)
	) name7219 (
		_w3733_,
		_w6759_,
		_w7681_
	);
	LUT2 #(
		.INIT('h1)
	) name7220 (
		_w7667_,
		_w7681_,
		_w7682_
	);
	LUT2 #(
		.INIT('h4)
	) name7221 (
		_w7674_,
		_w7682_,
		_w7683_
	);
	LUT2 #(
		.INIT('h1)
	) name7222 (
		_w7677_,
		_w7680_,
		_w7684_
	);
	LUT2 #(
		.INIT('h8)
	) name7223 (
		_w7683_,
		_w7684_,
		_w7685_
	);
	LUT2 #(
		.INIT('h4)
	) name7224 (
		_w7671_,
		_w7685_,
		_w7686_
	);
	LUT2 #(
		.INIT('h2)
	) name7225 (
		_w2026_,
		_w7686_,
		_w7687_
	);
	LUT2 #(
		.INIT('h1)
	) name7226 (
		_w7666_,
		_w7687_,
		_w7688_
	);
	LUT2 #(
		.INIT('h2)
	) name7227 (
		\P1_state_reg[0]/NET0131 ,
		_w7688_,
		_w7689_
	);
	LUT2 #(
		.INIT('h1)
	) name7228 (
		_w7665_,
		_w7689_,
		_w7690_
	);
	LUT2 #(
		.INIT('h2)
	) name7229 (
		\P2_reg1_reg[30]/NET0131 ,
		_w5962_,
		_w7691_
	);
	LUT2 #(
		.INIT('h2)
	) name7230 (
		_w5964_,
		_w7550_,
		_w7692_
	);
	LUT2 #(
		.INIT('h1)
	) name7231 (
		_w7691_,
		_w7692_,
		_w7693_
	);
	LUT2 #(
		.INIT('h2)
	) name7232 (
		\P1_reg2_reg[30]/NET0131 ,
		_w3466_,
		_w7694_
	);
	LUT2 #(
		.INIT('h8)
	) name7233 (
		_w3466_,
		_w5812_,
		_w7695_
	);
	LUT2 #(
		.INIT('h8)
	) name7234 (
		_w7492_,
		_w7695_,
		_w7696_
	);
	LUT2 #(
		.INIT('h1)
	) name7235 (
		_w7694_,
		_w7696_,
		_w7697_
	);
	LUT2 #(
		.INIT('h2)
	) name7236 (
		_w3712_,
		_w7697_,
		_w7698_
	);
	LUT2 #(
		.INIT('h2)
	) name7237 (
		_w3466_,
		_w7490_,
		_w7699_
	);
	LUT2 #(
		.INIT('h1)
	) name7238 (
		_w3720_,
		_w7699_,
		_w7700_
	);
	LUT2 #(
		.INIT('h2)
	) name7239 (
		_w5812_,
		_w7700_,
		_w7701_
	);
	LUT2 #(
		.INIT('h4)
	) name7240 (
		_w501_,
		_w1762_,
		_w7702_
	);
	LUT2 #(
		.INIT('h1)
	) name7241 (
		_w3466_,
		_w7702_,
		_w7703_
	);
	LUT2 #(
		.INIT('h2)
	) name7242 (
		_w5815_,
		_w7703_,
		_w7704_
	);
	LUT2 #(
		.INIT('h2)
	) name7243 (
		\P1_reg2_reg[30]/NET0131 ,
		_w7704_,
		_w7705_
	);
	LUT2 #(
		.INIT('h1)
	) name7244 (
		_w7701_,
		_w7705_,
		_w7706_
	);
	LUT2 #(
		.INIT('h4)
	) name7245 (
		_w7698_,
		_w7706_,
		_w7707_
	);
	LUT2 #(
		.INIT('h2)
	) name7246 (
		\P2_reg2_reg[12]/NET0131 ,
		_w1983_,
		_w7708_
	);
	LUT2 #(
		.INIT('h8)
	) name7247 (
		\P2_reg2_reg[12]/NET0131 ,
		_w2024_,
		_w7709_
	);
	LUT2 #(
		.INIT('h2)
	) name7248 (
		\P2_reg2_reg[12]/NET0131 ,
		_w3774_,
		_w7710_
	);
	LUT2 #(
		.INIT('h2)
	) name7249 (
		\P2_reg2_reg[12]/NET0131 ,
		_w3758_,
		_w7711_
	);
	LUT2 #(
		.INIT('h8)
	) name7250 (
		_w3758_,
		_w6186_,
		_w7712_
	);
	LUT2 #(
		.INIT('h1)
	) name7251 (
		_w7711_,
		_w7712_,
		_w7713_
	);
	LUT2 #(
		.INIT('h2)
	) name7252 (
		_w3411_,
		_w7713_,
		_w7714_
	);
	LUT2 #(
		.INIT('h8)
	) name7253 (
		_w3758_,
		_w6192_,
		_w7715_
	);
	LUT2 #(
		.INIT('h1)
	) name7254 (
		_w7711_,
		_w7715_,
		_w7716_
	);
	LUT2 #(
		.INIT('h1)
	) name7255 (
		_w3177_,
		_w7716_,
		_w7717_
	);
	LUT2 #(
		.INIT('h2)
	) name7256 (
		_w3758_,
		_w6198_,
		_w7718_
	);
	LUT2 #(
		.INIT('h1)
	) name7257 (
		_w7711_,
		_w7718_,
		_w7719_
	);
	LUT2 #(
		.INIT('h1)
	) name7258 (
		_w3320_,
		_w7719_,
		_w7720_
	);
	LUT2 #(
		.INIT('h8)
	) name7259 (
		_w3758_,
		_w6203_,
		_w7721_
	);
	LUT2 #(
		.INIT('h1)
	) name7260 (
		_w7711_,
		_w7721_,
		_w7722_
	);
	LUT2 #(
		.INIT('h2)
	) name7261 (
		_w3355_,
		_w7722_,
		_w7723_
	);
	LUT2 #(
		.INIT('h8)
	) name7262 (
		_w2709_,
		_w3420_,
		_w7724_
	);
	LUT2 #(
		.INIT('h8)
	) name7263 (
		_w3758_,
		_w7584_,
		_w7725_
	);
	LUT2 #(
		.INIT('h1)
	) name7264 (
		_w7710_,
		_w7724_,
		_w7726_
	);
	LUT2 #(
		.INIT('h4)
	) name7265 (
		_w7725_,
		_w7726_,
		_w7727_
	);
	LUT2 #(
		.INIT('h4)
	) name7266 (
		_w7723_,
		_w7727_,
		_w7728_
	);
	LUT2 #(
		.INIT('h4)
	) name7267 (
		_w7717_,
		_w7728_,
		_w7729_
	);
	LUT2 #(
		.INIT('h4)
	) name7268 (
		_w7720_,
		_w7729_,
		_w7730_
	);
	LUT2 #(
		.INIT('h4)
	) name7269 (
		_w7714_,
		_w7730_,
		_w7731_
	);
	LUT2 #(
		.INIT('h2)
	) name7270 (
		_w2026_,
		_w7731_,
		_w7732_
	);
	LUT2 #(
		.INIT('h1)
	) name7271 (
		_w7709_,
		_w7732_,
		_w7733_
	);
	LUT2 #(
		.INIT('h2)
	) name7272 (
		\P1_state_reg[0]/NET0131 ,
		_w7733_,
		_w7734_
	);
	LUT2 #(
		.INIT('h1)
	) name7273 (
		_w7708_,
		_w7734_,
		_w7735_
	);
	LUT2 #(
		.INIT('h2)
	) name7274 (
		\P2_reg2_reg[16]/NET0131 ,
		_w1983_,
		_w7736_
	);
	LUT2 #(
		.INIT('h8)
	) name7275 (
		\P2_reg2_reg[16]/NET0131 ,
		_w2024_,
		_w7737_
	);
	LUT2 #(
		.INIT('h2)
	) name7276 (
		\P2_reg2_reg[16]/NET0131 ,
		_w3774_,
		_w7738_
	);
	LUT2 #(
		.INIT('h2)
	) name7277 (
		\P2_reg2_reg[16]/NET0131 ,
		_w3758_,
		_w7739_
	);
	LUT2 #(
		.INIT('h2)
	) name7278 (
		_w3758_,
		_w6226_,
		_w7740_
	);
	LUT2 #(
		.INIT('h1)
	) name7279 (
		_w7739_,
		_w7740_,
		_w7741_
	);
	LUT2 #(
		.INIT('h1)
	) name7280 (
		_w3177_,
		_w7741_,
		_w7742_
	);
	LUT2 #(
		.INIT('h8)
	) name7281 (
		_w3758_,
		_w6234_,
		_w7743_
	);
	LUT2 #(
		.INIT('h1)
	) name7282 (
		_w7739_,
		_w7743_,
		_w7744_
	);
	LUT2 #(
		.INIT('h2)
	) name7283 (
		_w3411_,
		_w7744_,
		_w7745_
	);
	LUT2 #(
		.INIT('h8)
	) name7284 (
		_w3758_,
		_w6240_,
		_w7746_
	);
	LUT2 #(
		.INIT('h1)
	) name7285 (
		_w7739_,
		_w7746_,
		_w7747_
	);
	LUT2 #(
		.INIT('h2)
	) name7286 (
		_w3355_,
		_w7747_,
		_w7748_
	);
	LUT2 #(
		.INIT('h2)
	) name7287 (
		_w3758_,
		_w6246_,
		_w7749_
	);
	LUT2 #(
		.INIT('h1)
	) name7288 (
		_w7739_,
		_w7749_,
		_w7750_
	);
	LUT2 #(
		.INIT('h1)
	) name7289 (
		_w3320_,
		_w7750_,
		_w7751_
	);
	LUT2 #(
		.INIT('h8)
	) name7290 (
		_w2818_,
		_w3358_,
		_w7752_
	);
	LUT2 #(
		.INIT('h8)
	) name7291 (
		_w3758_,
		_w7752_,
		_w7753_
	);
	LUT2 #(
		.INIT('h8)
	) name7292 (
		_w2797_,
		_w3420_,
		_w7754_
	);
	LUT2 #(
		.INIT('h1)
	) name7293 (
		_w7738_,
		_w7754_,
		_w7755_
	);
	LUT2 #(
		.INIT('h4)
	) name7294 (
		_w7753_,
		_w7755_,
		_w7756_
	);
	LUT2 #(
		.INIT('h4)
	) name7295 (
		_w7748_,
		_w7756_,
		_w7757_
	);
	LUT2 #(
		.INIT('h4)
	) name7296 (
		_w7751_,
		_w7757_,
		_w7758_
	);
	LUT2 #(
		.INIT('h1)
	) name7297 (
		_w7742_,
		_w7745_,
		_w7759_
	);
	LUT2 #(
		.INIT('h8)
	) name7298 (
		_w7758_,
		_w7759_,
		_w7760_
	);
	LUT2 #(
		.INIT('h2)
	) name7299 (
		_w2026_,
		_w7760_,
		_w7761_
	);
	LUT2 #(
		.INIT('h1)
	) name7300 (
		_w7737_,
		_w7761_,
		_w7762_
	);
	LUT2 #(
		.INIT('h2)
	) name7301 (
		\P1_state_reg[0]/NET0131 ,
		_w7762_,
		_w7763_
	);
	LUT2 #(
		.INIT('h1)
	) name7302 (
		_w7736_,
		_w7763_,
		_w7764_
	);
	LUT2 #(
		.INIT('h2)
	) name7303 (
		_w3758_,
		_w6648_,
		_w7765_
	);
	LUT2 #(
		.INIT('h8)
	) name7304 (
		_w3126_,
		_w3419_,
		_w7766_
	);
	LUT2 #(
		.INIT('h1)
	) name7305 (
		_w7765_,
		_w7766_,
		_w7767_
	);
	LUT2 #(
		.INIT('h2)
	) name7306 (
		_w5287_,
		_w7767_,
		_w7768_
	);
	LUT2 #(
		.INIT('h1)
	) name7307 (
		_w3320_,
		_w3758_,
		_w7769_
	);
	LUT2 #(
		.INIT('h2)
	) name7308 (
		_w3774_,
		_w7769_,
		_w7770_
	);
	LUT2 #(
		.INIT('h1)
	) name7309 (
		_w3758_,
		_w6640_,
		_w7771_
	);
	LUT2 #(
		.INIT('h2)
	) name7310 (
		_w5287_,
		_w7771_,
		_w7772_
	);
	LUT2 #(
		.INIT('h8)
	) name7311 (
		_w7770_,
		_w7772_,
		_w7773_
	);
	LUT2 #(
		.INIT('h2)
	) name7312 (
		\P2_reg2_reg[21]/NET0131 ,
		_w7773_,
		_w7774_
	);
	LUT2 #(
		.INIT('h1)
	) name7313 (
		_w7768_,
		_w7774_,
		_w7775_
	);
	LUT2 #(
		.INIT('h2)
	) name7314 (
		\P2_reg2_reg[30]/NET0131 ,
		_w1983_,
		_w7776_
	);
	LUT2 #(
		.INIT('h8)
	) name7315 (
		\P2_reg2_reg[30]/NET0131 ,
		_w2024_,
		_w7777_
	);
	LUT2 #(
		.INIT('h2)
	) name7316 (
		\P2_reg2_reg[30]/NET0131 ,
		_w5290_,
		_w7778_
	);
	LUT2 #(
		.INIT('h2)
	) name7317 (
		_w3758_,
		_w7548_,
		_w7779_
	);
	LUT2 #(
		.INIT('h1)
	) name7318 (
		\P2_reg2_reg[30]/NET0131 ,
		_w3758_,
		_w7780_
	);
	LUT2 #(
		.INIT('h2)
	) name7319 (
		_w3355_,
		_w7780_,
		_w7781_
	);
	LUT2 #(
		.INIT('h4)
	) name7320 (
		_w7779_,
		_w7781_,
		_w7782_
	);
	LUT2 #(
		.INIT('h2)
	) name7321 (
		_w3758_,
		_w7546_,
		_w7783_
	);
	LUT2 #(
		.INIT('h1)
	) name7322 (
		_w3776_,
		_w7778_,
		_w7784_
	);
	LUT2 #(
		.INIT('h4)
	) name7323 (
		_w7783_,
		_w7784_,
		_w7785_
	);
	LUT2 #(
		.INIT('h4)
	) name7324 (
		_w7782_,
		_w7785_,
		_w7786_
	);
	LUT2 #(
		.INIT('h2)
	) name7325 (
		_w2026_,
		_w7786_,
		_w7787_
	);
	LUT2 #(
		.INIT('h1)
	) name7326 (
		_w7777_,
		_w7787_,
		_w7788_
	);
	LUT2 #(
		.INIT('h2)
	) name7327 (
		\P1_state_reg[0]/NET0131 ,
		_w7788_,
		_w7789_
	);
	LUT2 #(
		.INIT('h1)
	) name7328 (
		_w7776_,
		_w7789_,
		_w7790_
	);
	LUT2 #(
		.INIT('h2)
	) name7329 (
		\P1_reg0_reg[12]/NET0131 ,
		_w3435_,
		_w7791_
	);
	LUT2 #(
		.INIT('h8)
	) name7330 (
		\P1_reg0_reg[12]/NET0131 ,
		_w3448_,
		_w7792_
	);
	LUT2 #(
		.INIT('h8)
	) name7331 (
		_w4396_,
		_w7532_,
		_w7793_
	);
	LUT2 #(
		.INIT('h2)
	) name7332 (
		\P1_reg0_reg[12]/NET0131 ,
		_w4396_,
		_w7794_
	);
	LUT2 #(
		.INIT('h8)
	) name7333 (
		_w4396_,
		_w6098_,
		_w7795_
	);
	LUT2 #(
		.INIT('h1)
	) name7334 (
		_w7794_,
		_w7795_,
		_w7796_
	);
	LUT2 #(
		.INIT('h2)
	) name7335 (
		_w1936_,
		_w7796_,
		_w7797_
	);
	LUT2 #(
		.INIT('h8)
	) name7336 (
		_w4396_,
		_w6104_,
		_w7798_
	);
	LUT2 #(
		.INIT('h1)
	) name7337 (
		_w7794_,
		_w7798_,
		_w7799_
	);
	LUT2 #(
		.INIT('h1)
	) name7338 (
		_w3563_,
		_w7799_,
		_w7800_
	);
	LUT2 #(
		.INIT('h2)
	) name7339 (
		_w4396_,
		_w6110_,
		_w7801_
	);
	LUT2 #(
		.INIT('h1)
	) name7340 (
		_w7794_,
		_w7801_,
		_w7802_
	);
	LUT2 #(
		.INIT('h1)
	) name7341 (
		_w3677_,
		_w7802_,
		_w7803_
	);
	LUT2 #(
		.INIT('h8)
	) name7342 (
		_w4396_,
		_w6117_,
		_w7804_
	);
	LUT2 #(
		.INIT('h1)
	) name7343 (
		_w7794_,
		_w7804_,
		_w7805_
	);
	LUT2 #(
		.INIT('h2)
	) name7344 (
		_w3712_,
		_w7805_,
		_w7806_
	);
	LUT2 #(
		.INIT('h2)
	) name7345 (
		\P1_reg0_reg[12]/NET0131 ,
		_w4493_,
		_w7807_
	);
	LUT2 #(
		.INIT('h1)
	) name7346 (
		_w7793_,
		_w7807_,
		_w7808_
	);
	LUT2 #(
		.INIT('h4)
	) name7347 (
		_w7806_,
		_w7808_,
		_w7809_
	);
	LUT2 #(
		.INIT('h4)
	) name7348 (
		_w7800_,
		_w7809_,
		_w7810_
	);
	LUT2 #(
		.INIT('h4)
	) name7349 (
		_w7803_,
		_w7810_,
		_w7811_
	);
	LUT2 #(
		.INIT('h4)
	) name7350 (
		_w7797_,
		_w7811_,
		_w7812_
	);
	LUT2 #(
		.INIT('h2)
	) name7351 (
		_w3450_,
		_w7812_,
		_w7813_
	);
	LUT2 #(
		.INIT('h1)
	) name7352 (
		_w7792_,
		_w7813_,
		_w7814_
	);
	LUT2 #(
		.INIT('h2)
	) name7353 (
		\P1_state_reg[0]/NET0131 ,
		_w7814_,
		_w7815_
	);
	LUT2 #(
		.INIT('h1)
	) name7354 (
		_w7791_,
		_w7815_,
		_w7816_
	);
	LUT2 #(
		.INIT('h2)
	) name7355 (
		\P1_reg0_reg[16]/NET0131 ,
		_w3435_,
		_w7817_
	);
	LUT2 #(
		.INIT('h8)
	) name7356 (
		\P1_reg0_reg[16]/NET0131 ,
		_w3448_,
		_w7818_
	);
	LUT2 #(
		.INIT('h2)
	) name7357 (
		\P1_reg0_reg[16]/NET0131 ,
		_w6848_,
		_w7819_
	);
	LUT2 #(
		.INIT('h8)
	) name7358 (
		_w1936_,
		_w6149_,
		_w7820_
	);
	LUT2 #(
		.INIT('h1)
	) name7359 (
		_w3677_,
		_w6155_,
		_w7821_
	);
	LUT2 #(
		.INIT('h1)
	) name7360 (
		_w3563_,
		_w6141_,
		_w7822_
	);
	LUT2 #(
		.INIT('h1)
	) name7361 (
		_w6161_,
		_w7570_,
		_w7823_
	);
	LUT2 #(
		.INIT('h4)
	) name7362 (
		_w7821_,
		_w7823_,
		_w7824_
	);
	LUT2 #(
		.INIT('h4)
	) name7363 (
		_w7820_,
		_w7824_,
		_w7825_
	);
	LUT2 #(
		.INIT('h4)
	) name7364 (
		_w7822_,
		_w7825_,
		_w7826_
	);
	LUT2 #(
		.INIT('h2)
	) name7365 (
		_w4396_,
		_w7826_,
		_w7827_
	);
	LUT2 #(
		.INIT('h1)
	) name7366 (
		_w7819_,
		_w7827_,
		_w7828_
	);
	LUT2 #(
		.INIT('h2)
	) name7367 (
		_w3450_,
		_w7828_,
		_w7829_
	);
	LUT2 #(
		.INIT('h1)
	) name7368 (
		_w7818_,
		_w7829_,
		_w7830_
	);
	LUT2 #(
		.INIT('h2)
	) name7369 (
		\P1_state_reg[0]/NET0131 ,
		_w7830_,
		_w7831_
	);
	LUT2 #(
		.INIT('h1)
	) name7370 (
		_w7817_,
		_w7831_,
		_w7832_
	);
	LUT2 #(
		.INIT('h2)
	) name7371 (
		\P1_reg0_reg[20]/NET0131 ,
		_w3435_,
		_w7833_
	);
	LUT2 #(
		.INIT('h8)
	) name7372 (
		\P1_reg0_reg[20]/NET0131 ,
		_w3448_,
		_w7834_
	);
	LUT2 #(
		.INIT('h2)
	) name7373 (
		\P1_reg0_reg[20]/NET0131 ,
		_w4396_,
		_w7835_
	);
	LUT2 #(
		.INIT('h8)
	) name7374 (
		_w4396_,
		_w6492_,
		_w7836_
	);
	LUT2 #(
		.INIT('h1)
	) name7375 (
		_w7835_,
		_w7836_,
		_w7837_
	);
	LUT2 #(
		.INIT('h2)
	) name7376 (
		_w1936_,
		_w7837_,
		_w7838_
	);
	LUT2 #(
		.INIT('h8)
	) name7377 (
		_w4396_,
		_w6515_,
		_w7839_
	);
	LUT2 #(
		.INIT('h2)
	) name7378 (
		_w4396_,
		_w6499_,
		_w7840_
	);
	LUT2 #(
		.INIT('h1)
	) name7379 (
		_w7835_,
		_w7840_,
		_w7841_
	);
	LUT2 #(
		.INIT('h1)
	) name7380 (
		_w3677_,
		_w7841_,
		_w7842_
	);
	LUT2 #(
		.INIT('h2)
	) name7381 (
		_w4396_,
		_w6505_,
		_w7843_
	);
	LUT2 #(
		.INIT('h1)
	) name7382 (
		_w7835_,
		_w7843_,
		_w7844_
	);
	LUT2 #(
		.INIT('h1)
	) name7383 (
		_w3563_,
		_w7844_,
		_w7845_
	);
	LUT2 #(
		.INIT('h8)
	) name7384 (
		_w4396_,
		_w6510_,
		_w7846_
	);
	LUT2 #(
		.INIT('h1)
	) name7385 (
		_w7835_,
		_w7846_,
		_w7847_
	);
	LUT2 #(
		.INIT('h2)
	) name7386 (
		_w3712_,
		_w7847_,
		_w7848_
	);
	LUT2 #(
		.INIT('h2)
	) name7387 (
		\P1_reg0_reg[20]/NET0131 ,
		_w4493_,
		_w7849_
	);
	LUT2 #(
		.INIT('h1)
	) name7388 (
		_w7839_,
		_w7849_,
		_w7850_
	);
	LUT2 #(
		.INIT('h4)
	) name7389 (
		_w7848_,
		_w7850_,
		_w7851_
	);
	LUT2 #(
		.INIT('h4)
	) name7390 (
		_w7842_,
		_w7851_,
		_w7852_
	);
	LUT2 #(
		.INIT('h4)
	) name7391 (
		_w7845_,
		_w7852_,
		_w7853_
	);
	LUT2 #(
		.INIT('h4)
	) name7392 (
		_w7838_,
		_w7853_,
		_w7854_
	);
	LUT2 #(
		.INIT('h2)
	) name7393 (
		_w3450_,
		_w7854_,
		_w7855_
	);
	LUT2 #(
		.INIT('h1)
	) name7394 (
		_w7834_,
		_w7855_,
		_w7856_
	);
	LUT2 #(
		.INIT('h2)
	) name7395 (
		\P1_state_reg[0]/NET0131 ,
		_w7856_,
		_w7857_
	);
	LUT2 #(
		.INIT('h1)
	) name7396 (
		_w7833_,
		_w7857_,
		_w7858_
	);
	LUT2 #(
		.INIT('h2)
	) name7397 (
		\P1_reg0_reg[21]/NET0131 ,
		_w3435_,
		_w7859_
	);
	LUT2 #(
		.INIT('h8)
	) name7398 (
		\P1_reg0_reg[21]/NET0131 ,
		_w3448_,
		_w7860_
	);
	LUT2 #(
		.INIT('h8)
	) name7399 (
		_w4396_,
		_w6955_,
		_w7861_
	);
	LUT2 #(
		.INIT('h2)
	) name7400 (
		\P1_reg0_reg[21]/NET0131 ,
		_w4396_,
		_w7862_
	);
	LUT2 #(
		.INIT('h8)
	) name7401 (
		_w4396_,
		_w6962_,
		_w7863_
	);
	LUT2 #(
		.INIT('h1)
	) name7402 (
		_w7862_,
		_w7863_,
		_w7864_
	);
	LUT2 #(
		.INIT('h2)
	) name7403 (
		_w1936_,
		_w7864_,
		_w7865_
	);
	LUT2 #(
		.INIT('h2)
	) name7404 (
		_w4396_,
		_w6968_,
		_w7866_
	);
	LUT2 #(
		.INIT('h1)
	) name7405 (
		_w7862_,
		_w7866_,
		_w7867_
	);
	LUT2 #(
		.INIT('h1)
	) name7406 (
		_w3563_,
		_w7867_,
		_w7868_
	);
	LUT2 #(
		.INIT('h8)
	) name7407 (
		_w4396_,
		_w6974_,
		_w7869_
	);
	LUT2 #(
		.INIT('h1)
	) name7408 (
		_w7862_,
		_w7869_,
		_w7870_
	);
	LUT2 #(
		.INIT('h1)
	) name7409 (
		_w3677_,
		_w7870_,
		_w7871_
	);
	LUT2 #(
		.INIT('h8)
	) name7410 (
		_w4396_,
		_w6979_,
		_w7872_
	);
	LUT2 #(
		.INIT('h1)
	) name7411 (
		_w7862_,
		_w7872_,
		_w7873_
	);
	LUT2 #(
		.INIT('h2)
	) name7412 (
		_w3712_,
		_w7873_,
		_w7874_
	);
	LUT2 #(
		.INIT('h2)
	) name7413 (
		\P1_reg0_reg[21]/NET0131 ,
		_w4493_,
		_w7875_
	);
	LUT2 #(
		.INIT('h1)
	) name7414 (
		_w7861_,
		_w7875_,
		_w7876_
	);
	LUT2 #(
		.INIT('h4)
	) name7415 (
		_w7874_,
		_w7876_,
		_w7877_
	);
	LUT2 #(
		.INIT('h4)
	) name7416 (
		_w7865_,
		_w7877_,
		_w7878_
	);
	LUT2 #(
		.INIT('h1)
	) name7417 (
		_w7868_,
		_w7871_,
		_w7879_
	);
	LUT2 #(
		.INIT('h8)
	) name7418 (
		_w7878_,
		_w7879_,
		_w7880_
	);
	LUT2 #(
		.INIT('h2)
	) name7419 (
		_w3450_,
		_w7880_,
		_w7881_
	);
	LUT2 #(
		.INIT('h1)
	) name7420 (
		_w7860_,
		_w7881_,
		_w7882_
	);
	LUT2 #(
		.INIT('h2)
	) name7421 (
		\P1_state_reg[0]/NET0131 ,
		_w7882_,
		_w7883_
	);
	LUT2 #(
		.INIT('h1)
	) name7422 (
		_w7859_,
		_w7883_,
		_w7884_
	);
	LUT2 #(
		.INIT('h2)
	) name7423 (
		\P1_reg0_reg[30]/NET0131 ,
		_w6887_,
		_w7885_
	);
	LUT2 #(
		.INIT('h2)
	) name7424 (
		_w6886_,
		_w7494_,
		_w7886_
	);
	LUT2 #(
		.INIT('h1)
	) name7425 (
		_w7885_,
		_w7886_,
		_w7887_
	);
	LUT2 #(
		.INIT('h2)
	) name7426 (
		\P1_reg1_reg[12]/NET0131 ,
		_w3435_,
		_w7888_
	);
	LUT2 #(
		.INIT('h8)
	) name7427 (
		\P1_reg1_reg[12]/NET0131 ,
		_w3448_,
		_w7889_
	);
	LUT2 #(
		.INIT('h8)
	) name7428 (
		_w4532_,
		_w7532_,
		_w7890_
	);
	LUT2 #(
		.INIT('h2)
	) name7429 (
		\P1_reg1_reg[12]/NET0131 ,
		_w4532_,
		_w7891_
	);
	LUT2 #(
		.INIT('h8)
	) name7430 (
		_w4532_,
		_w6098_,
		_w7892_
	);
	LUT2 #(
		.INIT('h1)
	) name7431 (
		_w7891_,
		_w7892_,
		_w7893_
	);
	LUT2 #(
		.INIT('h2)
	) name7432 (
		_w1936_,
		_w7893_,
		_w7894_
	);
	LUT2 #(
		.INIT('h8)
	) name7433 (
		_w4532_,
		_w6104_,
		_w7895_
	);
	LUT2 #(
		.INIT('h1)
	) name7434 (
		_w7891_,
		_w7895_,
		_w7896_
	);
	LUT2 #(
		.INIT('h1)
	) name7435 (
		_w3563_,
		_w7896_,
		_w7897_
	);
	LUT2 #(
		.INIT('h2)
	) name7436 (
		_w4532_,
		_w6110_,
		_w7898_
	);
	LUT2 #(
		.INIT('h1)
	) name7437 (
		_w7891_,
		_w7898_,
		_w7899_
	);
	LUT2 #(
		.INIT('h1)
	) name7438 (
		_w3677_,
		_w7899_,
		_w7900_
	);
	LUT2 #(
		.INIT('h8)
	) name7439 (
		_w4532_,
		_w6117_,
		_w7901_
	);
	LUT2 #(
		.INIT('h1)
	) name7440 (
		_w7891_,
		_w7901_,
		_w7902_
	);
	LUT2 #(
		.INIT('h2)
	) name7441 (
		_w3712_,
		_w7902_,
		_w7903_
	);
	LUT2 #(
		.INIT('h2)
	) name7442 (
		\P1_reg1_reg[12]/NET0131 ,
		_w4541_,
		_w7904_
	);
	LUT2 #(
		.INIT('h1)
	) name7443 (
		_w7890_,
		_w7904_,
		_w7905_
	);
	LUT2 #(
		.INIT('h4)
	) name7444 (
		_w7903_,
		_w7905_,
		_w7906_
	);
	LUT2 #(
		.INIT('h4)
	) name7445 (
		_w7897_,
		_w7906_,
		_w7907_
	);
	LUT2 #(
		.INIT('h4)
	) name7446 (
		_w7900_,
		_w7907_,
		_w7908_
	);
	LUT2 #(
		.INIT('h4)
	) name7447 (
		_w7894_,
		_w7908_,
		_w7909_
	);
	LUT2 #(
		.INIT('h2)
	) name7448 (
		_w3450_,
		_w7909_,
		_w7910_
	);
	LUT2 #(
		.INIT('h1)
	) name7449 (
		_w7889_,
		_w7910_,
		_w7911_
	);
	LUT2 #(
		.INIT('h2)
	) name7450 (
		\P1_state_reg[0]/NET0131 ,
		_w7911_,
		_w7912_
	);
	LUT2 #(
		.INIT('h1)
	) name7451 (
		_w7888_,
		_w7912_,
		_w7913_
	);
	LUT2 #(
		.INIT('h2)
	) name7452 (
		\P1_reg1_reg[16]/NET0131 ,
		_w3435_,
		_w7914_
	);
	LUT2 #(
		.INIT('h8)
	) name7453 (
		\P1_reg1_reg[16]/NET0131 ,
		_w3448_,
		_w7915_
	);
	LUT2 #(
		.INIT('h2)
	) name7454 (
		_w4532_,
		_w7826_,
		_w7916_
	);
	LUT2 #(
		.INIT('h1)
	) name7455 (
		_w4532_,
		_w6846_,
		_w7917_
	);
	LUT2 #(
		.INIT('h2)
	) name7456 (
		_w4573_,
		_w7917_,
		_w7918_
	);
	LUT2 #(
		.INIT('h2)
	) name7457 (
		\P1_reg1_reg[16]/NET0131 ,
		_w7918_,
		_w7919_
	);
	LUT2 #(
		.INIT('h1)
	) name7458 (
		_w7916_,
		_w7919_,
		_w7920_
	);
	LUT2 #(
		.INIT('h2)
	) name7459 (
		_w3450_,
		_w7920_,
		_w7921_
	);
	LUT2 #(
		.INIT('h1)
	) name7460 (
		_w7915_,
		_w7921_,
		_w7922_
	);
	LUT2 #(
		.INIT('h2)
	) name7461 (
		\P1_state_reg[0]/NET0131 ,
		_w7922_,
		_w7923_
	);
	LUT2 #(
		.INIT('h1)
	) name7462 (
		_w7914_,
		_w7923_,
		_w7924_
	);
	LUT2 #(
		.INIT('h2)
	) name7463 (
		\P1_reg1_reg[20]/NET0131 ,
		_w3435_,
		_w7925_
	);
	LUT2 #(
		.INIT('h8)
	) name7464 (
		\P1_reg1_reg[20]/NET0131 ,
		_w3448_,
		_w7926_
	);
	LUT2 #(
		.INIT('h2)
	) name7465 (
		\P1_reg1_reg[20]/NET0131 ,
		_w4532_,
		_w7927_
	);
	LUT2 #(
		.INIT('h8)
	) name7466 (
		_w4532_,
		_w6492_,
		_w7928_
	);
	LUT2 #(
		.INIT('h1)
	) name7467 (
		_w7927_,
		_w7928_,
		_w7929_
	);
	LUT2 #(
		.INIT('h2)
	) name7468 (
		_w1936_,
		_w7929_,
		_w7930_
	);
	LUT2 #(
		.INIT('h8)
	) name7469 (
		_w4532_,
		_w6515_,
		_w7931_
	);
	LUT2 #(
		.INIT('h2)
	) name7470 (
		_w4532_,
		_w6499_,
		_w7932_
	);
	LUT2 #(
		.INIT('h1)
	) name7471 (
		_w7927_,
		_w7932_,
		_w7933_
	);
	LUT2 #(
		.INIT('h1)
	) name7472 (
		_w3677_,
		_w7933_,
		_w7934_
	);
	LUT2 #(
		.INIT('h2)
	) name7473 (
		_w4532_,
		_w6505_,
		_w7935_
	);
	LUT2 #(
		.INIT('h1)
	) name7474 (
		_w7927_,
		_w7935_,
		_w7936_
	);
	LUT2 #(
		.INIT('h1)
	) name7475 (
		_w3563_,
		_w7936_,
		_w7937_
	);
	LUT2 #(
		.INIT('h8)
	) name7476 (
		_w4532_,
		_w6510_,
		_w7938_
	);
	LUT2 #(
		.INIT('h1)
	) name7477 (
		_w7927_,
		_w7938_,
		_w7939_
	);
	LUT2 #(
		.INIT('h2)
	) name7478 (
		_w3712_,
		_w7939_,
		_w7940_
	);
	LUT2 #(
		.INIT('h2)
	) name7479 (
		\P1_reg1_reg[20]/NET0131 ,
		_w4541_,
		_w7941_
	);
	LUT2 #(
		.INIT('h1)
	) name7480 (
		_w7931_,
		_w7941_,
		_w7942_
	);
	LUT2 #(
		.INIT('h4)
	) name7481 (
		_w7940_,
		_w7942_,
		_w7943_
	);
	LUT2 #(
		.INIT('h4)
	) name7482 (
		_w7934_,
		_w7943_,
		_w7944_
	);
	LUT2 #(
		.INIT('h4)
	) name7483 (
		_w7937_,
		_w7944_,
		_w7945_
	);
	LUT2 #(
		.INIT('h4)
	) name7484 (
		_w7930_,
		_w7945_,
		_w7946_
	);
	LUT2 #(
		.INIT('h2)
	) name7485 (
		_w3450_,
		_w7946_,
		_w7947_
	);
	LUT2 #(
		.INIT('h1)
	) name7486 (
		_w7926_,
		_w7947_,
		_w7948_
	);
	LUT2 #(
		.INIT('h2)
	) name7487 (
		\P1_state_reg[0]/NET0131 ,
		_w7948_,
		_w7949_
	);
	LUT2 #(
		.INIT('h1)
	) name7488 (
		_w7925_,
		_w7949_,
		_w7950_
	);
	LUT2 #(
		.INIT('h2)
	) name7489 (
		\P2_reg0_reg[12]/NET0131 ,
		_w1983_,
		_w7951_
	);
	LUT2 #(
		.INIT('h8)
	) name7490 (
		\P2_reg0_reg[12]/NET0131 ,
		_w2024_,
		_w7952_
	);
	LUT2 #(
		.INIT('h2)
	) name7491 (
		_w2040_,
		_w7585_,
		_w7953_
	);
	LUT2 #(
		.INIT('h2)
	) name7492 (
		\P2_reg0_reg[12]/NET0131 ,
		_w2040_,
		_w7954_
	);
	LUT2 #(
		.INIT('h8)
	) name7493 (
		_w2040_,
		_w6186_,
		_w7955_
	);
	LUT2 #(
		.INIT('h1)
	) name7494 (
		_w7954_,
		_w7955_,
		_w7956_
	);
	LUT2 #(
		.INIT('h2)
	) name7495 (
		_w3411_,
		_w7956_,
		_w7957_
	);
	LUT2 #(
		.INIT('h8)
	) name7496 (
		_w2040_,
		_w6192_,
		_w7958_
	);
	LUT2 #(
		.INIT('h1)
	) name7497 (
		_w7954_,
		_w7958_,
		_w7959_
	);
	LUT2 #(
		.INIT('h1)
	) name7498 (
		_w3177_,
		_w7959_,
		_w7960_
	);
	LUT2 #(
		.INIT('h2)
	) name7499 (
		_w2040_,
		_w6198_,
		_w7961_
	);
	LUT2 #(
		.INIT('h1)
	) name7500 (
		_w7954_,
		_w7961_,
		_w7962_
	);
	LUT2 #(
		.INIT('h1)
	) name7501 (
		_w3320_,
		_w7962_,
		_w7963_
	);
	LUT2 #(
		.INIT('h2)
	) name7502 (
		\P2_reg0_reg[12]/NET0131 ,
		_w3425_,
		_w7964_
	);
	LUT2 #(
		.INIT('h1)
	) name7503 (
		_w7953_,
		_w7964_,
		_w7965_
	);
	LUT2 #(
		.INIT('h4)
	) name7504 (
		_w7960_,
		_w7965_,
		_w7966_
	);
	LUT2 #(
		.INIT('h4)
	) name7505 (
		_w7963_,
		_w7966_,
		_w7967_
	);
	LUT2 #(
		.INIT('h4)
	) name7506 (
		_w7957_,
		_w7967_,
		_w7968_
	);
	LUT2 #(
		.INIT('h2)
	) name7507 (
		_w2026_,
		_w7968_,
		_w7969_
	);
	LUT2 #(
		.INIT('h1)
	) name7508 (
		_w7952_,
		_w7969_,
		_w7970_
	);
	LUT2 #(
		.INIT('h2)
	) name7509 (
		\P1_state_reg[0]/NET0131 ,
		_w7970_,
		_w7971_
	);
	LUT2 #(
		.INIT('h1)
	) name7510 (
		_w7951_,
		_w7971_,
		_w7972_
	);
	LUT2 #(
		.INIT('h2)
	) name7511 (
		\P2_reg0_reg[16]/NET0131 ,
		_w1983_,
		_w7973_
	);
	LUT2 #(
		.INIT('h8)
	) name7512 (
		\P2_reg0_reg[16]/NET0131 ,
		_w2024_,
		_w7974_
	);
	LUT2 #(
		.INIT('h2)
	) name7513 (
		\P2_reg0_reg[16]/NET0131 ,
		_w2040_,
		_w7975_
	);
	LUT2 #(
		.INIT('h2)
	) name7514 (
		_w2040_,
		_w6226_,
		_w7976_
	);
	LUT2 #(
		.INIT('h1)
	) name7515 (
		_w7975_,
		_w7976_,
		_w7977_
	);
	LUT2 #(
		.INIT('h1)
	) name7516 (
		_w3177_,
		_w7977_,
		_w7978_
	);
	LUT2 #(
		.INIT('h8)
	) name7517 (
		_w2040_,
		_w6240_,
		_w7979_
	);
	LUT2 #(
		.INIT('h1)
	) name7518 (
		_w7975_,
		_w7979_,
		_w7980_
	);
	LUT2 #(
		.INIT('h2)
	) name7519 (
		_w3355_,
		_w7980_,
		_w7981_
	);
	LUT2 #(
		.INIT('h1)
	) name7520 (
		_w3320_,
		_w6246_,
		_w7982_
	);
	LUT2 #(
		.INIT('h1)
	) name7521 (
		_w7752_,
		_w7982_,
		_w7983_
	);
	LUT2 #(
		.INIT('h2)
	) name7522 (
		_w2040_,
		_w7983_,
		_w7984_
	);
	LUT2 #(
		.INIT('h2)
	) name7523 (
		\P2_reg0_reg[16]/NET0131 ,
		_w7506_,
		_w7985_
	);
	LUT2 #(
		.INIT('h8)
	) name7524 (
		_w2040_,
		_w6234_,
		_w7986_
	);
	LUT2 #(
		.INIT('h1)
	) name7525 (
		_w7975_,
		_w7986_,
		_w7987_
	);
	LUT2 #(
		.INIT('h2)
	) name7526 (
		_w3411_,
		_w7987_,
		_w7988_
	);
	LUT2 #(
		.INIT('h1)
	) name7527 (
		_w7981_,
		_w7985_,
		_w7989_
	);
	LUT2 #(
		.INIT('h4)
	) name7528 (
		_w7984_,
		_w7989_,
		_w7990_
	);
	LUT2 #(
		.INIT('h1)
	) name7529 (
		_w7978_,
		_w7988_,
		_w7991_
	);
	LUT2 #(
		.INIT('h8)
	) name7530 (
		_w7990_,
		_w7991_,
		_w7992_
	);
	LUT2 #(
		.INIT('h2)
	) name7531 (
		_w2026_,
		_w7992_,
		_w7993_
	);
	LUT2 #(
		.INIT('h1)
	) name7532 (
		_w7974_,
		_w7993_,
		_w7994_
	);
	LUT2 #(
		.INIT('h2)
	) name7533 (
		\P1_state_reg[0]/NET0131 ,
		_w7994_,
		_w7995_
	);
	LUT2 #(
		.INIT('h1)
	) name7534 (
		_w7973_,
		_w7995_,
		_w7996_
	);
	LUT2 #(
		.INIT('h2)
	) name7535 (
		\P1_reg3_reg[11]/NET0131 ,
		\P1_state_reg[0]/NET0131 ,
		_w7997_
	);
	LUT2 #(
		.INIT('h8)
	) name7536 (
		_w1203_,
		_w1953_,
		_w7998_
	);
	LUT2 #(
		.INIT('h8)
	) name7537 (
		_w1203_,
		_w3448_,
		_w7999_
	);
	LUT2 #(
		.INIT('h2)
	) name7538 (
		_w1203_,
		_w4910_,
		_w8000_
	);
	LUT2 #(
		.INIT('h2)
	) name7539 (
		_w1203_,
		_w3980_,
		_w8001_
	);
	LUT2 #(
		.INIT('h2)
	) name7540 (
		_w1772_,
		_w4404_,
		_w8002_
	);
	LUT2 #(
		.INIT('h4)
	) name7541 (
		_w1772_,
		_w4404_,
		_w8003_
	);
	LUT2 #(
		.INIT('h1)
	) name7542 (
		_w8002_,
		_w8003_,
		_w8004_
	);
	LUT2 #(
		.INIT('h2)
	) name7543 (
		_w3980_,
		_w8004_,
		_w8005_
	);
	LUT2 #(
		.INIT('h1)
	) name7544 (
		_w8001_,
		_w8005_,
		_w8006_
	);
	LUT2 #(
		.INIT('h1)
	) name7545 (
		_w3677_,
		_w8006_,
		_w8007_
	);
	LUT2 #(
		.INIT('h2)
	) name7546 (
		_w1772_,
		_w4447_,
		_w8008_
	);
	LUT2 #(
		.INIT('h4)
	) name7547 (
		_w1772_,
		_w4447_,
		_w8009_
	);
	LUT2 #(
		.INIT('h1)
	) name7548 (
		_w8008_,
		_w8009_,
		_w8010_
	);
	LUT2 #(
		.INIT('h8)
	) name7549 (
		_w3980_,
		_w8010_,
		_w8011_
	);
	LUT2 #(
		.INIT('h1)
	) name7550 (
		_w8001_,
		_w8011_,
		_w8012_
	);
	LUT2 #(
		.INIT('h1)
	) name7551 (
		_w3563_,
		_w8012_,
		_w8013_
	);
	LUT2 #(
		.INIT('h2)
	) name7552 (
		_w1174_,
		_w4069_,
		_w8014_
	);
	LUT2 #(
		.INIT('h1)
	) name7553 (
		_w4070_,
		_w8014_,
		_w8015_
	);
	LUT2 #(
		.INIT('h1)
	) name7554 (
		_w537_,
		_w8015_,
		_w8016_
	);
	LUT2 #(
		.INIT('h8)
	) name7555 (
		_w537_,
		_w1218_,
		_w8017_
	);
	LUT2 #(
		.INIT('h1)
	) name7556 (
		_w8016_,
		_w8017_,
		_w8018_
	);
	LUT2 #(
		.INIT('h8)
	) name7557 (
		_w3980_,
		_w8018_,
		_w8019_
	);
	LUT2 #(
		.INIT('h1)
	) name7558 (
		_w8001_,
		_w8019_,
		_w8020_
	);
	LUT2 #(
		.INIT('h2)
	) name7559 (
		_w1936_,
		_w8020_,
		_w8021_
	);
	LUT2 #(
		.INIT('h2)
	) name7560 (
		_w1198_,
		_w6114_,
		_w8022_
	);
	LUT2 #(
		.INIT('h1)
	) name7561 (
		_w6115_,
		_w8022_,
		_w8023_
	);
	LUT2 #(
		.INIT('h8)
	) name7562 (
		_w3712_,
		_w8023_,
		_w8024_
	);
	LUT2 #(
		.INIT('h8)
	) name7563 (
		_w3980_,
		_w8024_,
		_w8025_
	);
	LUT2 #(
		.INIT('h2)
	) name7564 (
		_w1198_,
		_w4067_,
		_w8026_
	);
	LUT2 #(
		.INIT('h1)
	) name7565 (
		_w8000_,
		_w8026_,
		_w8027_
	);
	LUT2 #(
		.INIT('h4)
	) name7566 (
		_w8025_,
		_w8027_,
		_w8028_
	);
	LUT2 #(
		.INIT('h4)
	) name7567 (
		_w8007_,
		_w8028_,
		_w8029_
	);
	LUT2 #(
		.INIT('h1)
	) name7568 (
		_w8013_,
		_w8021_,
		_w8030_
	);
	LUT2 #(
		.INIT('h8)
	) name7569 (
		_w8029_,
		_w8030_,
		_w8031_
	);
	LUT2 #(
		.INIT('h2)
	) name7570 (
		_w3450_,
		_w8031_,
		_w8032_
	);
	LUT2 #(
		.INIT('h1)
	) name7571 (
		_w7999_,
		_w8032_,
		_w8033_
	);
	LUT2 #(
		.INIT('h2)
	) name7572 (
		\P1_state_reg[0]/NET0131 ,
		_w8033_,
		_w8034_
	);
	LUT2 #(
		.INIT('h1)
	) name7573 (
		_w7997_,
		_w7998_,
		_w8035_
	);
	LUT2 #(
		.INIT('h4)
	) name7574 (
		_w8034_,
		_w8035_,
		_w8036_
	);
	LUT2 #(
		.INIT('h8)
	) name7575 (
		_w1113_,
		_w1953_,
		_w8037_
	);
	LUT2 #(
		.INIT('h2)
	) name7576 (
		\P1_reg3_reg[14]/NET0131 ,
		\P1_state_reg[0]/NET0131 ,
		_w8038_
	);
	LUT2 #(
		.INIT('h8)
	) name7577 (
		_w1113_,
		_w3448_,
		_w8039_
	);
	LUT2 #(
		.INIT('h2)
	) name7578 (
		_w1113_,
		_w4064_,
		_w8040_
	);
	LUT2 #(
		.INIT('h2)
	) name7579 (
		_w1113_,
		_w3980_,
		_w8041_
	);
	LUT2 #(
		.INIT('h1)
	) name7580 (
		_w1094_,
		_w7130_,
		_w8042_
	);
	LUT2 #(
		.INIT('h8)
	) name7581 (
		_w1094_,
		_w7130_,
		_w8043_
	);
	LUT2 #(
		.INIT('h1)
	) name7582 (
		_w8042_,
		_w8043_,
		_w8044_
	);
	LUT2 #(
		.INIT('h1)
	) name7583 (
		_w537_,
		_w8044_,
		_w8045_
	);
	LUT2 #(
		.INIT('h2)
	) name7584 (
		_w537_,
		_w1146_,
		_w8046_
	);
	LUT2 #(
		.INIT('h1)
	) name7585 (
		_w8045_,
		_w8046_,
		_w8047_
	);
	LUT2 #(
		.INIT('h2)
	) name7586 (
		_w3980_,
		_w8047_,
		_w8048_
	);
	LUT2 #(
		.INIT('h1)
	) name7587 (
		_w8041_,
		_w8048_,
		_w8049_
	);
	LUT2 #(
		.INIT('h2)
	) name7588 (
		_w1936_,
		_w8049_,
		_w8050_
	);
	LUT2 #(
		.INIT('h1)
	) name7589 (
		_w1815_,
		_w6031_,
		_w8051_
	);
	LUT2 #(
		.INIT('h8)
	) name7590 (
		_w1815_,
		_w6031_,
		_w8052_
	);
	LUT2 #(
		.INIT('h1)
	) name7591 (
		_w8051_,
		_w8052_,
		_w8053_
	);
	LUT2 #(
		.INIT('h1)
	) name7592 (
		_w3563_,
		_w8053_,
		_w8054_
	);
	LUT2 #(
		.INIT('h2)
	) name7593 (
		_w1815_,
		_w6019_,
		_w8055_
	);
	LUT2 #(
		.INIT('h4)
	) name7594 (
		_w1815_,
		_w6019_,
		_w8056_
	);
	LUT2 #(
		.INIT('h1)
	) name7595 (
		_w8055_,
		_w8056_,
		_w8057_
	);
	LUT2 #(
		.INIT('h4)
	) name7596 (
		_w8054_,
		_w8057_,
		_w8058_
	);
	LUT2 #(
		.INIT('h2)
	) name7597 (
		_w3980_,
		_w8058_,
		_w8059_
	);
	LUT2 #(
		.INIT('h1)
	) name7598 (
		_w8041_,
		_w8059_,
		_w8060_
	);
	LUT2 #(
		.INIT('h1)
	) name7599 (
		_w3563_,
		_w3980_,
		_w8061_
	);
	LUT2 #(
		.INIT('h2)
	) name7600 (
		_w3677_,
		_w8054_,
		_w8062_
	);
	LUT2 #(
		.INIT('h4)
	) name7601 (
		_w8061_,
		_w8062_,
		_w8063_
	);
	LUT2 #(
		.INIT('h1)
	) name7602 (
		_w8060_,
		_w8063_,
		_w8064_
	);
	LUT2 #(
		.INIT('h4)
	) name7603 (
		_w1109_,
		_w5440_,
		_w8065_
	);
	LUT2 #(
		.INIT('h2)
	) name7604 (
		_w1109_,
		_w5440_,
		_w8066_
	);
	LUT2 #(
		.INIT('h1)
	) name7605 (
		_w8065_,
		_w8066_,
		_w8067_
	);
	LUT2 #(
		.INIT('h8)
	) name7606 (
		_w3980_,
		_w8067_,
		_w8068_
	);
	LUT2 #(
		.INIT('h1)
	) name7607 (
		_w8041_,
		_w8068_,
		_w8069_
	);
	LUT2 #(
		.INIT('h2)
	) name7608 (
		_w3712_,
		_w8069_,
		_w8070_
	);
	LUT2 #(
		.INIT('h2)
	) name7609 (
		_w1109_,
		_w4067_,
		_w8071_
	);
	LUT2 #(
		.INIT('h1)
	) name7610 (
		_w8040_,
		_w8071_,
		_w8072_
	);
	LUT2 #(
		.INIT('h4)
	) name7611 (
		_w8070_,
		_w8072_,
		_w8073_
	);
	LUT2 #(
		.INIT('h4)
	) name7612 (
		_w8050_,
		_w8073_,
		_w8074_
	);
	LUT2 #(
		.INIT('h4)
	) name7613 (
		_w8064_,
		_w8074_,
		_w8075_
	);
	LUT2 #(
		.INIT('h2)
	) name7614 (
		_w3450_,
		_w8075_,
		_w8076_
	);
	LUT2 #(
		.INIT('h1)
	) name7615 (
		_w8039_,
		_w8076_,
		_w8077_
	);
	LUT2 #(
		.INIT('h2)
	) name7616 (
		\P1_state_reg[0]/NET0131 ,
		_w8077_,
		_w8078_
	);
	LUT2 #(
		.INIT('h1)
	) name7617 (
		_w8037_,
		_w8038_,
		_w8079_
	);
	LUT2 #(
		.INIT('h4)
	) name7618 (
		_w8078_,
		_w8079_,
		_w8080_
	);
	LUT2 #(
		.INIT('h8)
	) name7619 (
		_w1088_,
		_w1953_,
		_w8081_
	);
	LUT2 #(
		.INIT('h2)
	) name7620 (
		\P1_reg3_reg[15]/NET0131 ,
		\P1_state_reg[0]/NET0131 ,
		_w8082_
	);
	LUT2 #(
		.INIT('h8)
	) name7621 (
		_w1088_,
		_w3448_,
		_w8083_
	);
	LUT2 #(
		.INIT('h2)
	) name7622 (
		_w1088_,
		_w4910_,
		_w8084_
	);
	LUT2 #(
		.INIT('h2)
	) name7623 (
		_w1088_,
		_w3980_,
		_w8085_
	);
	LUT2 #(
		.INIT('h2)
	) name7624 (
		_w1788_,
		_w7414_,
		_w8086_
	);
	LUT2 #(
		.INIT('h4)
	) name7625 (
		_w1788_,
		_w7414_,
		_w8087_
	);
	LUT2 #(
		.INIT('h1)
	) name7626 (
		_w8086_,
		_w8087_,
		_w8088_
	);
	LUT2 #(
		.INIT('h2)
	) name7627 (
		_w3980_,
		_w8088_,
		_w8089_
	);
	LUT2 #(
		.INIT('h1)
	) name7628 (
		_w8085_,
		_w8089_,
		_w8090_
	);
	LUT2 #(
		.INIT('h1)
	) name7629 (
		_w3677_,
		_w8090_,
		_w8091_
	);
	LUT2 #(
		.INIT('h2)
	) name7630 (
		_w1788_,
		_w7427_,
		_w8092_
	);
	LUT2 #(
		.INIT('h4)
	) name7631 (
		_w1788_,
		_w7427_,
		_w8093_
	);
	LUT2 #(
		.INIT('h1)
	) name7632 (
		_w8092_,
		_w8093_,
		_w8094_
	);
	LUT2 #(
		.INIT('h8)
	) name7633 (
		_w3980_,
		_w8094_,
		_w8095_
	);
	LUT2 #(
		.INIT('h1)
	) name7634 (
		_w8085_,
		_w8095_,
		_w8096_
	);
	LUT2 #(
		.INIT('h1)
	) name7635 (
		_w3563_,
		_w8096_,
		_w8097_
	);
	LUT2 #(
		.INIT('h2)
	) name7636 (
		_w1475_,
		_w4470_,
		_w8098_
	);
	LUT2 #(
		.INIT('h1)
	) name7637 (
		_w4073_,
		_w8098_,
		_w8099_
	);
	LUT2 #(
		.INIT('h1)
	) name7638 (
		_w537_,
		_w8099_,
		_w8100_
	);
	LUT2 #(
		.INIT('h8)
	) name7639 (
		_w537_,
		_w1118_,
		_w8101_
	);
	LUT2 #(
		.INIT('h1)
	) name7640 (
		_w8100_,
		_w8101_,
		_w8102_
	);
	LUT2 #(
		.INIT('h8)
	) name7641 (
		_w3980_,
		_w8102_,
		_w8103_
	);
	LUT2 #(
		.INIT('h1)
	) name7642 (
		_w8085_,
		_w8103_,
		_w8104_
	);
	LUT2 #(
		.INIT('h2)
	) name7643 (
		_w1936_,
		_w8104_,
		_w8105_
	);
	LUT2 #(
		.INIT('h2)
	) name7644 (
		_w1083_,
		_w8065_,
		_w8106_
	);
	LUT2 #(
		.INIT('h1)
	) name7645 (
		_w5441_,
		_w8106_,
		_w8107_
	);
	LUT2 #(
		.INIT('h8)
	) name7646 (
		_w3712_,
		_w8107_,
		_w8108_
	);
	LUT2 #(
		.INIT('h8)
	) name7647 (
		_w3980_,
		_w8108_,
		_w8109_
	);
	LUT2 #(
		.INIT('h2)
	) name7648 (
		_w1083_,
		_w4067_,
		_w8110_
	);
	LUT2 #(
		.INIT('h1)
	) name7649 (
		_w8084_,
		_w8110_,
		_w8111_
	);
	LUT2 #(
		.INIT('h4)
	) name7650 (
		_w8109_,
		_w8111_,
		_w8112_
	);
	LUT2 #(
		.INIT('h4)
	) name7651 (
		_w8091_,
		_w8112_,
		_w8113_
	);
	LUT2 #(
		.INIT('h1)
	) name7652 (
		_w8097_,
		_w8105_,
		_w8114_
	);
	LUT2 #(
		.INIT('h8)
	) name7653 (
		_w8113_,
		_w8114_,
		_w8115_
	);
	LUT2 #(
		.INIT('h2)
	) name7654 (
		_w3450_,
		_w8115_,
		_w8116_
	);
	LUT2 #(
		.INIT('h1)
	) name7655 (
		_w8083_,
		_w8116_,
		_w8117_
	);
	LUT2 #(
		.INIT('h2)
	) name7656 (
		\P1_state_reg[0]/NET0131 ,
		_w8117_,
		_w8118_
	);
	LUT2 #(
		.INIT('h1)
	) name7657 (
		_w8081_,
		_w8082_,
		_w8119_
	);
	LUT2 #(
		.INIT('h4)
	) name7658 (
		_w8118_,
		_w8119_,
		_w8120_
	);
	LUT2 #(
		.INIT('h4)
	) name7659 (
		\P1_state_reg[0]/NET0131 ,
		\P2_reg3_reg[11]/NET0131 ,
		_w8121_
	);
	LUT2 #(
		.INIT('h8)
	) name7660 (
		_w2024_,
		_w2681_,
		_w8122_
	);
	LUT2 #(
		.INIT('h2)
	) name7661 (
		_w2681_,
		_w6312_,
		_w8123_
	);
	LUT2 #(
		.INIT('h2)
	) name7662 (
		_w2681_,
		_w3788_,
		_w8124_
	);
	LUT2 #(
		.INIT('h2)
	) name7663 (
		_w2715_,
		_w6179_,
		_w8125_
	);
	LUT2 #(
		.INIT('h1)
	) name7664 (
		_w6180_,
		_w8125_,
		_w8126_
	);
	LUT2 #(
		.INIT('h1)
	) name7665 (
		_w2058_,
		_w8126_,
		_w8127_
	);
	LUT2 #(
		.INIT('h8)
	) name7666 (
		_w2058_,
		_w2742_,
		_w8128_
	);
	LUT2 #(
		.INIT('h1)
	) name7667 (
		_w8127_,
		_w8128_,
		_w8129_
	);
	LUT2 #(
		.INIT('h8)
	) name7668 (
		_w3788_,
		_w8129_,
		_w8130_
	);
	LUT2 #(
		.INIT('h1)
	) name7669 (
		_w8124_,
		_w8130_,
		_w8131_
	);
	LUT2 #(
		.INIT('h2)
	) name7670 (
		_w3411_,
		_w8131_,
		_w8132_
	);
	LUT2 #(
		.INIT('h2)
	) name7671 (
		_w4201_,
		_w4804_,
		_w8133_
	);
	LUT2 #(
		.INIT('h4)
	) name7672 (
		_w4201_,
		_w4804_,
		_w8134_
	);
	LUT2 #(
		.INIT('h1)
	) name7673 (
		_w8133_,
		_w8134_,
		_w8135_
	);
	LUT2 #(
		.INIT('h8)
	) name7674 (
		_w3788_,
		_w8135_,
		_w8136_
	);
	LUT2 #(
		.INIT('h1)
	) name7675 (
		_w8124_,
		_w8136_,
		_w8137_
	);
	LUT2 #(
		.INIT('h1)
	) name7676 (
		_w3177_,
		_w8137_,
		_w8138_
	);
	LUT2 #(
		.INIT('h2)
	) name7677 (
		_w2704_,
		_w7179_,
		_w8139_
	);
	LUT2 #(
		.INIT('h1)
	) name7678 (
		_w3336_,
		_w8139_,
		_w8140_
	);
	LUT2 #(
		.INIT('h8)
	) name7679 (
		_w3788_,
		_w8140_,
		_w8141_
	);
	LUT2 #(
		.INIT('h1)
	) name7680 (
		_w8124_,
		_w8141_,
		_w8142_
	);
	LUT2 #(
		.INIT('h2)
	) name7681 (
		_w3355_,
		_w8142_,
		_w8143_
	);
	LUT2 #(
		.INIT('h2)
	) name7682 (
		_w4201_,
		_w4840_,
		_w8144_
	);
	LUT2 #(
		.INIT('h4)
	) name7683 (
		_w4201_,
		_w4840_,
		_w8145_
	);
	LUT2 #(
		.INIT('h1)
	) name7684 (
		_w8144_,
		_w8145_,
		_w8146_
	);
	LUT2 #(
		.INIT('h1)
	) name7685 (
		_w3320_,
		_w8146_,
		_w8147_
	);
	LUT2 #(
		.INIT('h8)
	) name7686 (
		_w3788_,
		_w8147_,
		_w8148_
	);
	LUT2 #(
		.INIT('h2)
	) name7687 (
		_w2704_,
		_w3965_,
		_w8149_
	);
	LUT2 #(
		.INIT('h1)
	) name7688 (
		_w8123_,
		_w8149_,
		_w8150_
	);
	LUT2 #(
		.INIT('h4)
	) name7689 (
		_w8148_,
		_w8150_,
		_w8151_
	);
	LUT2 #(
		.INIT('h4)
	) name7690 (
		_w8143_,
		_w8151_,
		_w8152_
	);
	LUT2 #(
		.INIT('h4)
	) name7691 (
		_w8138_,
		_w8152_,
		_w8153_
	);
	LUT2 #(
		.INIT('h4)
	) name7692 (
		_w8132_,
		_w8153_,
		_w8154_
	);
	LUT2 #(
		.INIT('h2)
	) name7693 (
		_w2026_,
		_w8154_,
		_w8155_
	);
	LUT2 #(
		.INIT('h1)
	) name7694 (
		_w8122_,
		_w8155_,
		_w8156_
	);
	LUT2 #(
		.INIT('h2)
	) name7695 (
		\P1_state_reg[0]/NET0131 ,
		_w8156_,
		_w8157_
	);
	LUT2 #(
		.INIT('h8)
	) name7696 (
		_w2681_,
		_w3976_,
		_w8158_
	);
	LUT2 #(
		.INIT('h1)
	) name7697 (
		_w8121_,
		_w8158_,
		_w8159_
	);
	LUT2 #(
		.INIT('h4)
	) name7698 (
		_w8157_,
		_w8159_,
		_w8160_
	);
	LUT2 #(
		.INIT('h8)
	) name7699 (
		_w2866_,
		_w3976_,
		_w8161_
	);
	LUT2 #(
		.INIT('h4)
	) name7700 (
		\P1_state_reg[0]/NET0131 ,
		\P2_reg3_reg[14]/NET0131 ,
		_w8162_
	);
	LUT2 #(
		.INIT('h8)
	) name7701 (
		_w2024_,
		_w2866_,
		_w8163_
	);
	LUT2 #(
		.INIT('h2)
	) name7702 (
		_w2860_,
		_w3965_,
		_w8164_
	);
	LUT2 #(
		.INIT('h2)
	) name7703 (
		_w2866_,
		_w3962_,
		_w8165_
	);
	LUT2 #(
		.INIT('h2)
	) name7704 (
		_w2866_,
		_w3788_,
		_w8166_
	);
	LUT2 #(
		.INIT('h2)
	) name7705 (
		_w2828_,
		_w3387_,
		_w8167_
	);
	LUT2 #(
		.INIT('h1)
	) name7706 (
		_w5564_,
		_w8167_,
		_w8168_
	);
	LUT2 #(
		.INIT('h1)
	) name7707 (
		_w2058_,
		_w8168_,
		_w8169_
	);
	LUT2 #(
		.INIT('h8)
	) name7708 (
		_w2058_,
		_w2880_,
		_w8170_
	);
	LUT2 #(
		.INIT('h1)
	) name7709 (
		_w8169_,
		_w8170_,
		_w8171_
	);
	LUT2 #(
		.INIT('h8)
	) name7710 (
		_w3788_,
		_w8171_,
		_w8172_
	);
	LUT2 #(
		.INIT('h1)
	) name7711 (
		_w8166_,
		_w8172_,
		_w8173_
	);
	LUT2 #(
		.INIT('h2)
	) name7712 (
		_w3411_,
		_w8173_,
		_w8174_
	);
	LUT2 #(
		.INIT('h2)
	) name7713 (
		_w2860_,
		_w7215_,
		_w8175_
	);
	LUT2 #(
		.INIT('h1)
	) name7714 (
		_w3339_,
		_w8175_,
		_w8176_
	);
	LUT2 #(
		.INIT('h8)
	) name7715 (
		_w3788_,
		_w8176_,
		_w8177_
	);
	LUT2 #(
		.INIT('h1)
	) name7716 (
		_w8166_,
		_w8177_,
		_w8178_
	);
	LUT2 #(
		.INIT('h2)
	) name7717 (
		_w3355_,
		_w8178_,
		_w8179_
	);
	LUT2 #(
		.INIT('h2)
	) name7718 (
		_w4210_,
		_w4745_,
		_w8180_
	);
	LUT2 #(
		.INIT('h4)
	) name7719 (
		_w4210_,
		_w4745_,
		_w8181_
	);
	LUT2 #(
		.INIT('h1)
	) name7720 (
		_w8180_,
		_w8181_,
		_w8182_
	);
	LUT2 #(
		.INIT('h8)
	) name7721 (
		_w3788_,
		_w8182_,
		_w8183_
	);
	LUT2 #(
		.INIT('h1)
	) name7722 (
		_w8166_,
		_w8183_,
		_w8184_
	);
	LUT2 #(
		.INIT('h1)
	) name7723 (
		_w3177_,
		_w8184_,
		_w8185_
	);
	LUT2 #(
		.INIT('h2)
	) name7724 (
		_w4210_,
		_w4714_,
		_w8186_
	);
	LUT2 #(
		.INIT('h4)
	) name7725 (
		_w4210_,
		_w4714_,
		_w8187_
	);
	LUT2 #(
		.INIT('h1)
	) name7726 (
		_w8186_,
		_w8187_,
		_w8188_
	);
	LUT2 #(
		.INIT('h2)
	) name7727 (
		_w3788_,
		_w8188_,
		_w8189_
	);
	LUT2 #(
		.INIT('h1)
	) name7728 (
		_w8166_,
		_w8189_,
		_w8190_
	);
	LUT2 #(
		.INIT('h1)
	) name7729 (
		_w3320_,
		_w8190_,
		_w8191_
	);
	LUT2 #(
		.INIT('h1)
	) name7730 (
		_w8164_,
		_w8165_,
		_w8192_
	);
	LUT2 #(
		.INIT('h4)
	) name7731 (
		_w8174_,
		_w8192_,
		_w8193_
	);
	LUT2 #(
		.INIT('h1)
	) name7732 (
		_w8179_,
		_w8185_,
		_w8194_
	);
	LUT2 #(
		.INIT('h4)
	) name7733 (
		_w8191_,
		_w8194_,
		_w8195_
	);
	LUT2 #(
		.INIT('h8)
	) name7734 (
		_w8193_,
		_w8195_,
		_w8196_
	);
	LUT2 #(
		.INIT('h2)
	) name7735 (
		_w2026_,
		_w8196_,
		_w8197_
	);
	LUT2 #(
		.INIT('h1)
	) name7736 (
		_w8163_,
		_w8197_,
		_w8198_
	);
	LUT2 #(
		.INIT('h2)
	) name7737 (
		\P1_state_reg[0]/NET0131 ,
		_w8198_,
		_w8199_
	);
	LUT2 #(
		.INIT('h1)
	) name7738 (
		_w8161_,
		_w8162_,
		_w8200_
	);
	LUT2 #(
		.INIT('h4)
	) name7739 (
		_w8199_,
		_w8200_,
		_w8201_
	);
	LUT2 #(
		.INIT('h8)
	) name7740 (
		_w2822_,
		_w3976_,
		_w8202_
	);
	LUT2 #(
		.INIT('h4)
	) name7741 (
		\P1_state_reg[0]/NET0131 ,
		\P2_reg3_reg[15]/NET0131 ,
		_w8203_
	);
	LUT2 #(
		.INIT('h8)
	) name7742 (
		_w2024_,
		_w2822_,
		_w8204_
	);
	LUT2 #(
		.INIT('h2)
	) name7743 (
		_w2843_,
		_w3965_,
		_w8205_
	);
	LUT2 #(
		.INIT('h2)
	) name7744 (
		_w2822_,
		_w3788_,
		_w8206_
	);
	LUT2 #(
		.INIT('h2)
	) name7745 (
		_w2804_,
		_w5564_,
		_w8207_
	);
	LUT2 #(
		.INIT('h1)
	) name7746 (
		_w5565_,
		_w8207_,
		_w8208_
	);
	LUT2 #(
		.INIT('h1)
	) name7747 (
		_w2058_,
		_w8208_,
		_w8209_
	);
	LUT2 #(
		.INIT('h8)
	) name7748 (
		_w2058_,
		_w2870_,
		_w8210_
	);
	LUT2 #(
		.INIT('h1)
	) name7749 (
		_w8209_,
		_w8210_,
		_w8211_
	);
	LUT2 #(
		.INIT('h8)
	) name7750 (
		_w3788_,
		_w8211_,
		_w8212_
	);
	LUT2 #(
		.INIT('h1)
	) name7751 (
		_w8206_,
		_w8212_,
		_w8213_
	);
	LUT2 #(
		.INIT('h2)
	) name7752 (
		_w3411_,
		_w8213_,
		_w8214_
	);
	LUT2 #(
		.INIT('h2)
	) name7753 (
		_w4215_,
		_w4809_,
		_w8215_
	);
	LUT2 #(
		.INIT('h4)
	) name7754 (
		_w4215_,
		_w4809_,
		_w8216_
	);
	LUT2 #(
		.INIT('h1)
	) name7755 (
		_w8215_,
		_w8216_,
		_w8217_
	);
	LUT2 #(
		.INIT('h8)
	) name7756 (
		_w3788_,
		_w8217_,
		_w8218_
	);
	LUT2 #(
		.INIT('h1)
	) name7757 (
		_w8206_,
		_w8218_,
		_w8219_
	);
	LUT2 #(
		.INIT('h1)
	) name7758 (
		_w3177_,
		_w8219_,
		_w8220_
	);
	LUT2 #(
		.INIT('h2)
	) name7759 (
		_w2843_,
		_w3339_,
		_w8221_
	);
	LUT2 #(
		.INIT('h1)
	) name7760 (
		_w5574_,
		_w8221_,
		_w8222_
	);
	LUT2 #(
		.INIT('h8)
	) name7761 (
		_w3788_,
		_w8222_,
		_w8223_
	);
	LUT2 #(
		.INIT('h1)
	) name7762 (
		_w8206_,
		_w8223_,
		_w8224_
	);
	LUT2 #(
		.INIT('h2)
	) name7763 (
		_w3355_,
		_w8224_,
		_w8225_
	);
	LUT2 #(
		.INIT('h2)
	) name7764 (
		_w4215_,
		_w4845_,
		_w8226_
	);
	LUT2 #(
		.INIT('h4)
	) name7765 (
		_w4215_,
		_w4845_,
		_w8227_
	);
	LUT2 #(
		.INIT('h1)
	) name7766 (
		_w8226_,
		_w8227_,
		_w8228_
	);
	LUT2 #(
		.INIT('h2)
	) name7767 (
		_w3788_,
		_w8228_,
		_w8229_
	);
	LUT2 #(
		.INIT('h1)
	) name7768 (
		_w8206_,
		_w8229_,
		_w8230_
	);
	LUT2 #(
		.INIT('h1)
	) name7769 (
		_w3320_,
		_w8230_,
		_w8231_
	);
	LUT2 #(
		.INIT('h2)
	) name7770 (
		_w2822_,
		_w3962_,
		_w8232_
	);
	LUT2 #(
		.INIT('h1)
	) name7771 (
		_w8205_,
		_w8232_,
		_w8233_
	);
	LUT2 #(
		.INIT('h4)
	) name7772 (
		_w8231_,
		_w8233_,
		_w8234_
	);
	LUT2 #(
		.INIT('h4)
	) name7773 (
		_w8225_,
		_w8234_,
		_w8235_
	);
	LUT2 #(
		.INIT('h4)
	) name7774 (
		_w8214_,
		_w8235_,
		_w8236_
	);
	LUT2 #(
		.INIT('h4)
	) name7775 (
		_w8220_,
		_w8236_,
		_w8237_
	);
	LUT2 #(
		.INIT('h2)
	) name7776 (
		_w2026_,
		_w8237_,
		_w8238_
	);
	LUT2 #(
		.INIT('h1)
	) name7777 (
		_w8204_,
		_w8238_,
		_w8239_
	);
	LUT2 #(
		.INIT('h2)
	) name7778 (
		\P1_state_reg[0]/NET0131 ,
		_w8239_,
		_w8240_
	);
	LUT2 #(
		.INIT('h1)
	) name7779 (
		_w8202_,
		_w8203_,
		_w8241_
	);
	LUT2 #(
		.INIT('h4)
	) name7780 (
		_w8240_,
		_w8241_,
		_w8242_
	);
	LUT2 #(
		.INIT('h4)
	) name7781 (
		\P1_state_reg[0]/NET0131 ,
		\P2_reg3_reg[8]/NET0131 ,
		_w8243_
	);
	LUT2 #(
		.INIT('h8)
	) name7782 (
		_w2447_,
		_w3976_,
		_w8244_
	);
	LUT2 #(
		.INIT('h8)
	) name7783 (
		_w2024_,
		_w2447_,
		_w8245_
	);
	LUT2 #(
		.INIT('h2)
	) name7784 (
		_w2447_,
		_w5698_,
		_w8246_
	);
	LUT2 #(
		.INIT('h2)
	) name7785 (
		_w2447_,
		_w3788_,
		_w8247_
	);
	LUT2 #(
		.INIT('h2)
	) name7786 (
		_w2765_,
		_w7242_,
		_w8248_
	);
	LUT2 #(
		.INIT('h1)
	) name7787 (
		_w7243_,
		_w8248_,
		_w8249_
	);
	LUT2 #(
		.INIT('h1)
	) name7788 (
		_w2058_,
		_w8249_,
		_w8250_
	);
	LUT2 #(
		.INIT('h8)
	) name7789 (
		_w2058_,
		_w2480_,
		_w8251_
	);
	LUT2 #(
		.INIT('h1)
	) name7790 (
		_w8250_,
		_w8251_,
		_w8252_
	);
	LUT2 #(
		.INIT('h8)
	) name7791 (
		_w3788_,
		_w8252_,
		_w8253_
	);
	LUT2 #(
		.INIT('h1)
	) name7792 (
		_w8247_,
		_w8253_,
		_w8254_
	);
	LUT2 #(
		.INIT('h2)
	) name7793 (
		_w3411_,
		_w8254_,
		_w8255_
	);
	LUT2 #(
		.INIT('h4)
	) name7794 (
		_w3889_,
		_w4208_,
		_w8256_
	);
	LUT2 #(
		.INIT('h2)
	) name7795 (
		_w3889_,
		_w4208_,
		_w8257_
	);
	LUT2 #(
		.INIT('h1)
	) name7796 (
		_w8256_,
		_w8257_,
		_w8258_
	);
	LUT2 #(
		.INIT('h8)
	) name7797 (
		_w3788_,
		_w8258_,
		_w8259_
	);
	LUT2 #(
		.INIT('h1)
	) name7798 (
		_w8247_,
		_w8259_,
		_w8260_
	);
	LUT2 #(
		.INIT('h1)
	) name7799 (
		_w3177_,
		_w8260_,
		_w8261_
	);
	LUT2 #(
		.INIT('h4)
	) name7800 (
		_w3831_,
		_w4208_,
		_w8262_
	);
	LUT2 #(
		.INIT('h2)
	) name7801 (
		_w3831_,
		_w4208_,
		_w8263_
	);
	LUT2 #(
		.INIT('h1)
	) name7802 (
		_w8262_,
		_w8263_,
		_w8264_
	);
	LUT2 #(
		.INIT('h2)
	) name7803 (
		_w3788_,
		_w8264_,
		_w8265_
	);
	LUT2 #(
		.INIT('h1)
	) name7804 (
		_w8247_,
		_w8265_,
		_w8266_
	);
	LUT2 #(
		.INIT('h1)
	) name7805 (
		_w3320_,
		_w8266_,
		_w8267_
	);
	LUT2 #(
		.INIT('h2)
	) name7806 (
		_w2470_,
		_w3332_,
		_w8268_
	);
	LUT2 #(
		.INIT('h1)
	) name7807 (
		_w7258_,
		_w8268_,
		_w8269_
	);
	LUT2 #(
		.INIT('h8)
	) name7808 (
		_w3355_,
		_w8269_,
		_w8270_
	);
	LUT2 #(
		.INIT('h8)
	) name7809 (
		_w3788_,
		_w8270_,
		_w8271_
	);
	LUT2 #(
		.INIT('h2)
	) name7810 (
		_w2470_,
		_w3965_,
		_w8272_
	);
	LUT2 #(
		.INIT('h1)
	) name7811 (
		_w8246_,
		_w8272_,
		_w8273_
	);
	LUT2 #(
		.INIT('h4)
	) name7812 (
		_w8271_,
		_w8273_,
		_w8274_
	);
	LUT2 #(
		.INIT('h4)
	) name7813 (
		_w8261_,
		_w8274_,
		_w8275_
	);
	LUT2 #(
		.INIT('h4)
	) name7814 (
		_w8267_,
		_w8275_,
		_w8276_
	);
	LUT2 #(
		.INIT('h4)
	) name7815 (
		_w8255_,
		_w8276_,
		_w8277_
	);
	LUT2 #(
		.INIT('h2)
	) name7816 (
		_w2026_,
		_w8277_,
		_w8278_
	);
	LUT2 #(
		.INIT('h1)
	) name7817 (
		_w8245_,
		_w8278_,
		_w8279_
	);
	LUT2 #(
		.INIT('h2)
	) name7818 (
		\P1_state_reg[0]/NET0131 ,
		_w8279_,
		_w8280_
	);
	LUT2 #(
		.INIT('h1)
	) name7819 (
		_w8243_,
		_w8244_,
		_w8281_
	);
	LUT2 #(
		.INIT('h4)
	) name7820 (
		_w8280_,
		_w8281_,
		_w8282_
	);
	LUT2 #(
		.INIT('h2)
	) name7821 (
		\P1_reg3_reg[8]/NET0131 ,
		\P1_state_reg[0]/NET0131 ,
		_w8283_
	);
	LUT2 #(
		.INIT('h8)
	) name7822 (
		_w1262_,
		_w1953_,
		_w8284_
	);
	LUT2 #(
		.INIT('h8)
	) name7823 (
		_w1262_,
		_w3448_,
		_w8285_
	);
	LUT2 #(
		.INIT('h2)
	) name7824 (
		_w1281_,
		_w4067_,
		_w8286_
	);
	LUT2 #(
		.INIT('h2)
	) name7825 (
		_w1262_,
		_w3980_,
		_w8287_
	);
	LUT2 #(
		.INIT('h2)
	) name7826 (
		_w1244_,
		_w7305_,
		_w8288_
	);
	LUT2 #(
		.INIT('h1)
	) name7827 (
		_w7306_,
		_w8288_,
		_w8289_
	);
	LUT2 #(
		.INIT('h1)
	) name7828 (
		_w537_,
		_w8289_,
		_w8290_
	);
	LUT2 #(
		.INIT('h8)
	) name7829 (
		_w537_,
		_w1498_,
		_w8291_
	);
	LUT2 #(
		.INIT('h1)
	) name7830 (
		_w8290_,
		_w8291_,
		_w8292_
	);
	LUT2 #(
		.INIT('h8)
	) name7831 (
		_w3980_,
		_w8292_,
		_w8293_
	);
	LUT2 #(
		.INIT('h1)
	) name7832 (
		_w8287_,
		_w8293_,
		_w8294_
	);
	LUT2 #(
		.INIT('h2)
	) name7833 (
		_w1936_,
		_w8294_,
		_w8295_
	);
	LUT2 #(
		.INIT('h2)
	) name7834 (
		_w1802_,
		_w3996_,
		_w8296_
	);
	LUT2 #(
		.INIT('h4)
	) name7835 (
		_w1802_,
		_w3996_,
		_w8297_
	);
	LUT2 #(
		.INIT('h1)
	) name7836 (
		_w8296_,
		_w8297_,
		_w8298_
	);
	LUT2 #(
		.INIT('h8)
	) name7837 (
		_w3980_,
		_w8298_,
		_w8299_
	);
	LUT2 #(
		.INIT('h1)
	) name7838 (
		_w8287_,
		_w8299_,
		_w8300_
	);
	LUT2 #(
		.INIT('h1)
	) name7839 (
		_w3563_,
		_w8300_,
		_w8301_
	);
	LUT2 #(
		.INIT('h4)
	) name7840 (
		_w1746_,
		_w1802_,
		_w8302_
	);
	LUT2 #(
		.INIT('h2)
	) name7841 (
		_w1746_,
		_w1802_,
		_w8303_
	);
	LUT2 #(
		.INIT('h1)
	) name7842 (
		_w8302_,
		_w8303_,
		_w8304_
	);
	LUT2 #(
		.INIT('h2)
	) name7843 (
		_w3980_,
		_w8304_,
		_w8305_
	);
	LUT2 #(
		.INIT('h1)
	) name7844 (
		_w8287_,
		_w8305_,
		_w8306_
	);
	LUT2 #(
		.INIT('h1)
	) name7845 (
		_w3677_,
		_w8306_,
		_w8307_
	);
	LUT2 #(
		.INIT('h8)
	) name7846 (
		_w1514_,
		_w3684_,
		_w8308_
	);
	LUT2 #(
		.INIT('h2)
	) name7847 (
		_w1281_,
		_w8308_,
		_w8309_
	);
	LUT2 #(
		.INIT('h1)
	) name7848 (
		_w7298_,
		_w8309_,
		_w8310_
	);
	LUT2 #(
		.INIT('h8)
	) name7849 (
		_w3980_,
		_w8310_,
		_w8311_
	);
	LUT2 #(
		.INIT('h1)
	) name7850 (
		_w8287_,
		_w8311_,
		_w8312_
	);
	LUT2 #(
		.INIT('h2)
	) name7851 (
		_w3712_,
		_w8312_,
		_w8313_
	);
	LUT2 #(
		.INIT('h2)
	) name7852 (
		_w1262_,
		_w4064_,
		_w8314_
	);
	LUT2 #(
		.INIT('h1)
	) name7853 (
		_w8286_,
		_w8314_,
		_w8315_
	);
	LUT2 #(
		.INIT('h4)
	) name7854 (
		_w8313_,
		_w8315_,
		_w8316_
	);
	LUT2 #(
		.INIT('h4)
	) name7855 (
		_w8301_,
		_w8316_,
		_w8317_
	);
	LUT2 #(
		.INIT('h4)
	) name7856 (
		_w8307_,
		_w8317_,
		_w8318_
	);
	LUT2 #(
		.INIT('h4)
	) name7857 (
		_w8295_,
		_w8318_,
		_w8319_
	);
	LUT2 #(
		.INIT('h2)
	) name7858 (
		_w3450_,
		_w8319_,
		_w8320_
	);
	LUT2 #(
		.INIT('h1)
	) name7859 (
		_w8285_,
		_w8320_,
		_w8321_
	);
	LUT2 #(
		.INIT('h2)
	) name7860 (
		\P1_state_reg[0]/NET0131 ,
		_w8321_,
		_w8322_
	);
	LUT2 #(
		.INIT('h1)
	) name7861 (
		_w8283_,
		_w8284_,
		_w8323_
	);
	LUT2 #(
		.INIT('h4)
	) name7862 (
		_w8322_,
		_w8323_,
		_w8324_
	);
	LUT2 #(
		.INIT('h8)
	) name7863 (
		_w2024_,
		_w3084_,
		_w8325_
	);
	LUT2 #(
		.INIT('h2)
	) name7864 (
		_w3084_,
		_w3788_,
		_w8326_
	);
	LUT2 #(
		.INIT('h4)
	) name7865 (
		_w4814_,
		_w4816_,
		_w8327_
	);
	LUT2 #(
		.INIT('h2)
	) name7866 (
		_w4821_,
		_w8327_,
		_w8328_
	);
	LUT2 #(
		.INIT('h2)
	) name7867 (
		_w4196_,
		_w8328_,
		_w8329_
	);
	LUT2 #(
		.INIT('h4)
	) name7868 (
		_w4196_,
		_w8328_,
		_w8330_
	);
	LUT2 #(
		.INIT('h1)
	) name7869 (
		_w8329_,
		_w8330_,
		_w8331_
	);
	LUT2 #(
		.INIT('h8)
	) name7870 (
		_w3788_,
		_w8331_,
		_w8332_
	);
	LUT2 #(
		.INIT('h1)
	) name7871 (
		_w8326_,
		_w8332_,
		_w8333_
	);
	LUT2 #(
		.INIT('h1)
	) name7872 (
		_w3177_,
		_w8333_,
		_w8334_
	);
	LUT2 #(
		.INIT('h2)
	) name7873 (
		_w3079_,
		_w5768_,
		_w8335_
	);
	LUT2 #(
		.INIT('h1)
	) name7874 (
		_w4614_,
		_w8335_,
		_w8336_
	);
	LUT2 #(
		.INIT('h8)
	) name7875 (
		_w3788_,
		_w8336_,
		_w8337_
	);
	LUT2 #(
		.INIT('h1)
	) name7876 (
		_w8326_,
		_w8337_,
		_w8338_
	);
	LUT2 #(
		.INIT('h2)
	) name7877 (
		_w3355_,
		_w8338_,
		_w8339_
	);
	LUT2 #(
		.INIT('h4)
	) name7878 (
		_w4850_,
		_w4851_,
		_w8340_
	);
	LUT2 #(
		.INIT('h2)
	) name7879 (
		_w4856_,
		_w8340_,
		_w8341_
	);
	LUT2 #(
		.INIT('h2)
	) name7880 (
		_w4196_,
		_w8341_,
		_w8342_
	);
	LUT2 #(
		.INIT('h4)
	) name7881 (
		_w4196_,
		_w8341_,
		_w8343_
	);
	LUT2 #(
		.INIT('h1)
	) name7882 (
		_w8342_,
		_w8343_,
		_w8344_
	);
	LUT2 #(
		.INIT('h2)
	) name7883 (
		_w3788_,
		_w8344_,
		_w8345_
	);
	LUT2 #(
		.INIT('h1)
	) name7884 (
		_w8326_,
		_w8345_,
		_w8346_
	);
	LUT2 #(
		.INIT('h1)
	) name7885 (
		_w3320_,
		_w8346_,
		_w8347_
	);
	LUT2 #(
		.INIT('h2)
	) name7886 (
		_w2058_,
		_w3112_,
		_w8348_
	);
	LUT2 #(
		.INIT('h2)
	) name7887 (
		_w3065_,
		_w5775_,
		_w8349_
	);
	LUT2 #(
		.INIT('h1)
	) name7888 (
		_w2058_,
		_w4622_,
		_w8350_
	);
	LUT2 #(
		.INIT('h4)
	) name7889 (
		_w8349_,
		_w8350_,
		_w8351_
	);
	LUT2 #(
		.INIT('h1)
	) name7890 (
		_w8348_,
		_w8351_,
		_w8352_
	);
	LUT2 #(
		.INIT('h2)
	) name7891 (
		_w3788_,
		_w8352_,
		_w8353_
	);
	LUT2 #(
		.INIT('h1)
	) name7892 (
		_w8326_,
		_w8353_,
		_w8354_
	);
	LUT2 #(
		.INIT('h2)
	) name7893 (
		_w3411_,
		_w8354_,
		_w8355_
	);
	LUT2 #(
		.INIT('h2)
	) name7894 (
		_w3084_,
		_w3962_,
		_w8356_
	);
	LUT2 #(
		.INIT('h2)
	) name7895 (
		_w3079_,
		_w3965_,
		_w8357_
	);
	LUT2 #(
		.INIT('h1)
	) name7896 (
		_w8356_,
		_w8357_,
		_w8358_
	);
	LUT2 #(
		.INIT('h4)
	) name7897 (
		_w8355_,
		_w8358_,
		_w8359_
	);
	LUT2 #(
		.INIT('h4)
	) name7898 (
		_w8347_,
		_w8359_,
		_w8360_
	);
	LUT2 #(
		.INIT('h4)
	) name7899 (
		_w8339_,
		_w8360_,
		_w8361_
	);
	LUT2 #(
		.INIT('h4)
	) name7900 (
		_w8334_,
		_w8361_,
		_w8362_
	);
	LUT2 #(
		.INIT('h2)
	) name7901 (
		_w2026_,
		_w8362_,
		_w8363_
	);
	LUT2 #(
		.INIT('h1)
	) name7902 (
		_w8325_,
		_w8363_,
		_w8364_
	);
	LUT2 #(
		.INIT('h2)
	) name7903 (
		\P1_state_reg[0]/NET0131 ,
		_w8364_,
		_w8365_
	);
	LUT2 #(
		.INIT('h4)
	) name7904 (
		\P1_state_reg[0]/NET0131 ,
		\P2_reg3_reg[23]/NET0131 ,
		_w8366_
	);
	LUT2 #(
		.INIT('h8)
	) name7905 (
		_w3084_,
		_w3976_,
		_w8367_
	);
	LUT2 #(
		.INIT('h1)
	) name7906 (
		_w8366_,
		_w8367_,
		_w8368_
	);
	LUT2 #(
		.INIT('h4)
	) name7907 (
		_w8365_,
		_w8368_,
		_w8369_
	);
	LUT2 #(
		.INIT('h2)
	) name7908 (
		\P2_reg0_reg[23]/NET0131 ,
		_w1983_,
		_w8370_
	);
	LUT2 #(
		.INIT('h8)
	) name7909 (
		\P2_reg0_reg[23]/NET0131 ,
		_w2024_,
		_w8371_
	);
	LUT2 #(
		.INIT('h2)
	) name7910 (
		\P2_reg0_reg[23]/NET0131 ,
		_w2040_,
		_w8372_
	);
	LUT2 #(
		.INIT('h8)
	) name7911 (
		_w2040_,
		_w8331_,
		_w8373_
	);
	LUT2 #(
		.INIT('h1)
	) name7912 (
		_w8372_,
		_w8373_,
		_w8374_
	);
	LUT2 #(
		.INIT('h1)
	) name7913 (
		_w3177_,
		_w8374_,
		_w8375_
	);
	LUT2 #(
		.INIT('h8)
	) name7914 (
		_w3355_,
		_w8336_,
		_w8376_
	);
	LUT2 #(
		.INIT('h8)
	) name7915 (
		_w3079_,
		_w3358_,
		_w8377_
	);
	LUT2 #(
		.INIT('h1)
	) name7916 (
		_w3320_,
		_w8344_,
		_w8378_
	);
	LUT2 #(
		.INIT('h1)
	) name7917 (
		_w8377_,
		_w8378_,
		_w8379_
	);
	LUT2 #(
		.INIT('h4)
	) name7918 (
		_w8376_,
		_w8379_,
		_w8380_
	);
	LUT2 #(
		.INIT('h2)
	) name7919 (
		_w2040_,
		_w8380_,
		_w8381_
	);
	LUT2 #(
		.INIT('h2)
	) name7920 (
		_w2040_,
		_w8352_,
		_w8382_
	);
	LUT2 #(
		.INIT('h1)
	) name7921 (
		_w8372_,
		_w8382_,
		_w8383_
	);
	LUT2 #(
		.INIT('h2)
	) name7922 (
		_w3411_,
		_w8383_,
		_w8384_
	);
	LUT2 #(
		.INIT('h4)
	) name7923 (
		_w3424_,
		_w7506_,
		_w8385_
	);
	LUT2 #(
		.INIT('h2)
	) name7924 (
		\P2_reg0_reg[23]/NET0131 ,
		_w8385_,
		_w8386_
	);
	LUT2 #(
		.INIT('h1)
	) name7925 (
		_w8384_,
		_w8386_,
		_w8387_
	);
	LUT2 #(
		.INIT('h4)
	) name7926 (
		_w8381_,
		_w8387_,
		_w8388_
	);
	LUT2 #(
		.INIT('h4)
	) name7927 (
		_w8375_,
		_w8388_,
		_w8389_
	);
	LUT2 #(
		.INIT('h2)
	) name7928 (
		_w2026_,
		_w8389_,
		_w8390_
	);
	LUT2 #(
		.INIT('h1)
	) name7929 (
		_w8371_,
		_w8390_,
		_w8391_
	);
	LUT2 #(
		.INIT('h2)
	) name7930 (
		\P1_state_reg[0]/NET0131 ,
		_w8391_,
		_w8392_
	);
	LUT2 #(
		.INIT('h1)
	) name7931 (
		_w8370_,
		_w8392_,
		_w8393_
	);
	LUT2 #(
		.INIT('h2)
	) name7932 (
		\P1_reg1_reg[9]/NET0131 ,
		_w3435_,
		_w8394_
	);
	LUT2 #(
		.INIT('h8)
	) name7933 (
		\P1_reg1_reg[9]/NET0131 ,
		_w3448_,
		_w8395_
	);
	LUT2 #(
		.INIT('h8)
	) name7934 (
		_w1257_,
		_w1880_,
		_w8396_
	);
	LUT2 #(
		.INIT('h8)
	) name7935 (
		_w4532_,
		_w8396_,
		_w8397_
	);
	LUT2 #(
		.INIT('h2)
	) name7936 (
		\P1_reg1_reg[9]/NET0131 ,
		_w4532_,
		_w8398_
	);
	LUT2 #(
		.INIT('h8)
	) name7937 (
		_w4532_,
		_w7294_,
		_w8399_
	);
	LUT2 #(
		.INIT('h1)
	) name7938 (
		_w8398_,
		_w8399_,
		_w8400_
	);
	LUT2 #(
		.INIT('h1)
	) name7939 (
		_w3563_,
		_w8400_,
		_w8401_
	);
	LUT2 #(
		.INIT('h2)
	) name7940 (
		_w4532_,
		_w7288_,
		_w8402_
	);
	LUT2 #(
		.INIT('h1)
	) name7941 (
		_w8398_,
		_w8402_,
		_w8403_
	);
	LUT2 #(
		.INIT('h1)
	) name7942 (
		_w3677_,
		_w8403_,
		_w8404_
	);
	LUT2 #(
		.INIT('h8)
	) name7943 (
		_w4532_,
		_w7300_,
		_w8405_
	);
	LUT2 #(
		.INIT('h1)
	) name7944 (
		_w8398_,
		_w8405_,
		_w8406_
	);
	LUT2 #(
		.INIT('h2)
	) name7945 (
		_w3712_,
		_w8406_,
		_w8407_
	);
	LUT2 #(
		.INIT('h2)
	) name7946 (
		_w4532_,
		_w7310_,
		_w8408_
	);
	LUT2 #(
		.INIT('h1)
	) name7947 (
		_w8398_,
		_w8408_,
		_w8409_
	);
	LUT2 #(
		.INIT('h2)
	) name7948 (
		_w1936_,
		_w8409_,
		_w8410_
	);
	LUT2 #(
		.INIT('h2)
	) name7949 (
		\P1_reg1_reg[9]/NET0131 ,
		_w4541_,
		_w8411_
	);
	LUT2 #(
		.INIT('h1)
	) name7950 (
		_w8397_,
		_w8411_,
		_w8412_
	);
	LUT2 #(
		.INIT('h4)
	) name7951 (
		_w8407_,
		_w8412_,
		_w8413_
	);
	LUT2 #(
		.INIT('h4)
	) name7952 (
		_w8401_,
		_w8413_,
		_w8414_
	);
	LUT2 #(
		.INIT('h4)
	) name7953 (
		_w8404_,
		_w8414_,
		_w8415_
	);
	LUT2 #(
		.INIT('h4)
	) name7954 (
		_w8410_,
		_w8415_,
		_w8416_
	);
	LUT2 #(
		.INIT('h2)
	) name7955 (
		_w3450_,
		_w8416_,
		_w8417_
	);
	LUT2 #(
		.INIT('h1)
	) name7956 (
		_w8395_,
		_w8417_,
		_w8418_
	);
	LUT2 #(
		.INIT('h2)
	) name7957 (
		\P1_state_reg[0]/NET0131 ,
		_w8418_,
		_w8419_
	);
	LUT2 #(
		.INIT('h1)
	) name7958 (
		_w8394_,
		_w8419_,
		_w8420_
	);
	LUT2 #(
		.INIT('h2)
	) name7959 (
		\P1_reg2_reg[10]/NET0131 ,
		_w3435_,
		_w8421_
	);
	LUT2 #(
		.INIT('h8)
	) name7960 (
		\P1_reg2_reg[10]/NET0131 ,
		_w3448_,
		_w8422_
	);
	LUT2 #(
		.INIT('h8)
	) name7961 (
		_w1233_,
		_w1880_,
		_w8423_
	);
	LUT2 #(
		.INIT('h8)
	) name7962 (
		_w3466_,
		_w8423_,
		_w8424_
	);
	LUT2 #(
		.INIT('h2)
	) name7963 (
		\P1_reg2_reg[10]/NET0131 ,
		_w3466_,
		_w8425_
	);
	LUT2 #(
		.INIT('h8)
	) name7964 (
		_w3466_,
		_w7086_,
		_w8426_
	);
	LUT2 #(
		.INIT('h1)
	) name7965 (
		_w8425_,
		_w8426_,
		_w8427_
	);
	LUT2 #(
		.INIT('h2)
	) name7966 (
		_w1936_,
		_w8427_,
		_w8428_
	);
	LUT2 #(
		.INIT('h8)
	) name7967 (
		_w3466_,
		_w7092_,
		_w8429_
	);
	LUT2 #(
		.INIT('h1)
	) name7968 (
		_w8425_,
		_w8429_,
		_w8430_
	);
	LUT2 #(
		.INIT('h1)
	) name7969 (
		_w3563_,
		_w8430_,
		_w8431_
	);
	LUT2 #(
		.INIT('h2)
	) name7970 (
		_w3466_,
		_w7078_,
		_w8432_
	);
	LUT2 #(
		.INIT('h1)
	) name7971 (
		_w8425_,
		_w8432_,
		_w8433_
	);
	LUT2 #(
		.INIT('h1)
	) name7972 (
		_w3677_,
		_w8433_,
		_w8434_
	);
	LUT2 #(
		.INIT('h8)
	) name7973 (
		_w3466_,
		_w7097_,
		_w8435_
	);
	LUT2 #(
		.INIT('h1)
	) name7974 (
		_w8425_,
		_w8435_,
		_w8436_
	);
	LUT2 #(
		.INIT('h2)
	) name7975 (
		_w3712_,
		_w8436_,
		_w8437_
	);
	LUT2 #(
		.INIT('h8)
	) name7976 (
		_w1214_,
		_w1763_,
		_w8438_
	);
	LUT2 #(
		.INIT('h2)
	) name7977 (
		\P1_reg2_reg[10]/NET0131 ,
		_w3718_,
		_w8439_
	);
	LUT2 #(
		.INIT('h1)
	) name7978 (
		_w8424_,
		_w8438_,
		_w8440_
	);
	LUT2 #(
		.INIT('h4)
	) name7979 (
		_w8439_,
		_w8440_,
		_w8441_
	);
	LUT2 #(
		.INIT('h4)
	) name7980 (
		_w8437_,
		_w8441_,
		_w8442_
	);
	LUT2 #(
		.INIT('h4)
	) name7981 (
		_w8428_,
		_w8442_,
		_w8443_
	);
	LUT2 #(
		.INIT('h1)
	) name7982 (
		_w8431_,
		_w8434_,
		_w8444_
	);
	LUT2 #(
		.INIT('h8)
	) name7983 (
		_w8443_,
		_w8444_,
		_w8445_
	);
	LUT2 #(
		.INIT('h2)
	) name7984 (
		_w3450_,
		_w8445_,
		_w8446_
	);
	LUT2 #(
		.INIT('h1)
	) name7985 (
		_w8422_,
		_w8446_,
		_w8447_
	);
	LUT2 #(
		.INIT('h2)
	) name7986 (
		\P1_state_reg[0]/NET0131 ,
		_w8447_,
		_w8448_
	);
	LUT2 #(
		.INIT('h1)
	) name7987 (
		_w8421_,
		_w8448_,
		_w8449_
	);
	LUT2 #(
		.INIT('h2)
	) name7988 (
		\P1_reg2_reg[13]/NET0131 ,
		_w3435_,
		_w8450_
	);
	LUT2 #(
		.INIT('h8)
	) name7989 (
		\P1_reg2_reg[13]/NET0131 ,
		_w3448_,
		_w8451_
	);
	LUT2 #(
		.INIT('h2)
	) name7990 (
		\P1_reg2_reg[13]/NET0131 ,
		_w3718_,
		_w8452_
	);
	LUT2 #(
		.INIT('h2)
	) name7991 (
		\P1_reg2_reg[13]/NET0131 ,
		_w3466_,
		_w8453_
	);
	LUT2 #(
		.INIT('h8)
	) name7992 (
		_w3466_,
		_w7125_,
		_w8454_
	);
	LUT2 #(
		.INIT('h1)
	) name7993 (
		_w8453_,
		_w8454_,
		_w8455_
	);
	LUT2 #(
		.INIT('h1)
	) name7994 (
		_w3563_,
		_w8455_,
		_w8456_
	);
	LUT2 #(
		.INIT('h8)
	) name7995 (
		_w3466_,
		_w7134_,
		_w8457_
	);
	LUT2 #(
		.INIT('h1)
	) name7996 (
		_w8453_,
		_w8457_,
		_w8458_
	);
	LUT2 #(
		.INIT('h2)
	) name7997 (
		_w1936_,
		_w8458_,
		_w8459_
	);
	LUT2 #(
		.INIT('h2)
	) name7998 (
		_w3466_,
		_w7119_,
		_w8460_
	);
	LUT2 #(
		.INIT('h1)
	) name7999 (
		_w8453_,
		_w8460_,
		_w8461_
	);
	LUT2 #(
		.INIT('h1)
	) name8000 (
		_w3677_,
		_w8461_,
		_w8462_
	);
	LUT2 #(
		.INIT('h8)
	) name8001 (
		_w3466_,
		_w7139_,
		_w8463_
	);
	LUT2 #(
		.INIT('h1)
	) name8002 (
		_w8453_,
		_w8463_,
		_w8464_
	);
	LUT2 #(
		.INIT('h2)
	) name8003 (
		_w3712_,
		_w8464_,
		_w8465_
	);
	LUT2 #(
		.INIT('h8)
	) name8004 (
		_w1140_,
		_w1763_,
		_w8466_
	);
	LUT2 #(
		.INIT('h8)
	) name8005 (
		_w1136_,
		_w1880_,
		_w8467_
	);
	LUT2 #(
		.INIT('h8)
	) name8006 (
		_w3466_,
		_w8467_,
		_w8468_
	);
	LUT2 #(
		.INIT('h1)
	) name8007 (
		_w8466_,
		_w8468_,
		_w8469_
	);
	LUT2 #(
		.INIT('h4)
	) name8008 (
		_w8452_,
		_w8469_,
		_w8470_
	);
	LUT2 #(
		.INIT('h4)
	) name8009 (
		_w8465_,
		_w8470_,
		_w8471_
	);
	LUT2 #(
		.INIT('h4)
	) name8010 (
		_w8456_,
		_w8471_,
		_w8472_
	);
	LUT2 #(
		.INIT('h1)
	) name8011 (
		_w8459_,
		_w8462_,
		_w8473_
	);
	LUT2 #(
		.INIT('h8)
	) name8012 (
		_w8472_,
		_w8473_,
		_w8474_
	);
	LUT2 #(
		.INIT('h2)
	) name8013 (
		_w3450_,
		_w8474_,
		_w8475_
	);
	LUT2 #(
		.INIT('h1)
	) name8014 (
		_w8451_,
		_w8475_,
		_w8476_
	);
	LUT2 #(
		.INIT('h2)
	) name8015 (
		\P1_state_reg[0]/NET0131 ,
		_w8476_,
		_w8477_
	);
	LUT2 #(
		.INIT('h1)
	) name8016 (
		_w8450_,
		_w8477_,
		_w8478_
	);
	LUT2 #(
		.INIT('h2)
	) name8017 (
		\P2_reg0_reg[9]/NET0131 ,
		_w1983_,
		_w8479_
	);
	LUT2 #(
		.INIT('h8)
	) name8018 (
		\P2_reg0_reg[9]/NET0131 ,
		_w2024_,
		_w8480_
	);
	LUT2 #(
		.INIT('h2)
	) name8019 (
		\P2_reg0_reg[9]/NET0131 ,
		_w8385_,
		_w8481_
	);
	LUT2 #(
		.INIT('h2)
	) name8020 (
		\P2_reg0_reg[9]/NET0131 ,
		_w2040_,
		_w8482_
	);
	LUT2 #(
		.INIT('h8)
	) name8021 (
		_w2040_,
		_w7248_,
		_w8483_
	);
	LUT2 #(
		.INIT('h1)
	) name8022 (
		_w8482_,
		_w8483_,
		_w8484_
	);
	LUT2 #(
		.INIT('h2)
	) name8023 (
		_w3411_,
		_w8484_,
		_w8485_
	);
	LUT2 #(
		.INIT('h2)
	) name8024 (
		_w2040_,
		_w7254_,
		_w8486_
	);
	LUT2 #(
		.INIT('h1)
	) name8025 (
		_w8482_,
		_w8486_,
		_w8487_
	);
	LUT2 #(
		.INIT('h1)
	) name8026 (
		_w3177_,
		_w8487_,
		_w8488_
	);
	LUT2 #(
		.INIT('h8)
	) name8027 (
		_w2779_,
		_w3358_,
		_w8489_
	);
	LUT2 #(
		.INIT('h8)
	) name8028 (
		_w3355_,
		_w7260_,
		_w8490_
	);
	LUT2 #(
		.INIT('h1)
	) name8029 (
		_w7267_,
		_w8489_,
		_w8491_
	);
	LUT2 #(
		.INIT('h4)
	) name8030 (
		_w8490_,
		_w8491_,
		_w8492_
	);
	LUT2 #(
		.INIT('h2)
	) name8031 (
		_w2040_,
		_w8492_,
		_w8493_
	);
	LUT2 #(
		.INIT('h1)
	) name8032 (
		_w8481_,
		_w8493_,
		_w8494_
	);
	LUT2 #(
		.INIT('h4)
	) name8033 (
		_w8488_,
		_w8494_,
		_w8495_
	);
	LUT2 #(
		.INIT('h4)
	) name8034 (
		_w8485_,
		_w8495_,
		_w8496_
	);
	LUT2 #(
		.INIT('h2)
	) name8035 (
		_w2026_,
		_w8496_,
		_w8497_
	);
	LUT2 #(
		.INIT('h1)
	) name8036 (
		_w8480_,
		_w8497_,
		_w8498_
	);
	LUT2 #(
		.INIT('h2)
	) name8037 (
		\P1_state_reg[0]/NET0131 ,
		_w8498_,
		_w8499_
	);
	LUT2 #(
		.INIT('h1)
	) name8038 (
		_w8479_,
		_w8499_,
		_w8500_
	);
	LUT2 #(
		.INIT('h2)
	) name8039 (
		\P2_reg1_reg[10]/NET0131 ,
		_w1983_,
		_w8501_
	);
	LUT2 #(
		.INIT('h8)
	) name8040 (
		\P2_reg1_reg[10]/NET0131 ,
		_w2024_,
		_w8502_
	);
	LUT2 #(
		.INIT('h8)
	) name8041 (
		_w2755_,
		_w3358_,
		_w8503_
	);
	LUT2 #(
		.INIT('h8)
	) name8042 (
		_w3733_,
		_w8503_,
		_w8504_
	);
	LUT2 #(
		.INIT('h2)
	) name8043 (
		\P2_reg1_reg[10]/NET0131 ,
		_w3733_,
		_w8505_
	);
	LUT2 #(
		.INIT('h8)
	) name8044 (
		_w3733_,
		_w7163_,
		_w8506_
	);
	LUT2 #(
		.INIT('h1)
	) name8045 (
		_w8505_,
		_w8506_,
		_w8507_
	);
	LUT2 #(
		.INIT('h2)
	) name8046 (
		_w3411_,
		_w8507_,
		_w8508_
	);
	LUT2 #(
		.INIT('h2)
	) name8047 (
		_w3733_,
		_w7169_,
		_w8509_
	);
	LUT2 #(
		.INIT('h1)
	) name8048 (
		_w8505_,
		_w8509_,
		_w8510_
	);
	LUT2 #(
		.INIT('h1)
	) name8049 (
		_w3177_,
		_w8510_,
		_w8511_
	);
	LUT2 #(
		.INIT('h8)
	) name8050 (
		_w3733_,
		_w7175_,
		_w8512_
	);
	LUT2 #(
		.INIT('h1)
	) name8051 (
		_w8505_,
		_w8512_,
		_w8513_
	);
	LUT2 #(
		.INIT('h1)
	) name8052 (
		_w3320_,
		_w8513_,
		_w8514_
	);
	LUT2 #(
		.INIT('h8)
	) name8053 (
		_w3733_,
		_w7181_,
		_w8515_
	);
	LUT2 #(
		.INIT('h1)
	) name8054 (
		_w8505_,
		_w8515_,
		_w8516_
	);
	LUT2 #(
		.INIT('h2)
	) name8055 (
		_w3355_,
		_w8516_,
		_w8517_
	);
	LUT2 #(
		.INIT('h2)
	) name8056 (
		\P2_reg1_reg[10]/NET0131 ,
		_w3743_,
		_w8518_
	);
	LUT2 #(
		.INIT('h1)
	) name8057 (
		_w8504_,
		_w8518_,
		_w8519_
	);
	LUT2 #(
		.INIT('h4)
	) name8058 (
		_w8517_,
		_w8519_,
		_w8520_
	);
	LUT2 #(
		.INIT('h4)
	) name8059 (
		_w8511_,
		_w8520_,
		_w8521_
	);
	LUT2 #(
		.INIT('h4)
	) name8060 (
		_w8514_,
		_w8521_,
		_w8522_
	);
	LUT2 #(
		.INIT('h4)
	) name8061 (
		_w8508_,
		_w8522_,
		_w8523_
	);
	LUT2 #(
		.INIT('h2)
	) name8062 (
		_w2026_,
		_w8523_,
		_w8524_
	);
	LUT2 #(
		.INIT('h1)
	) name8063 (
		_w8502_,
		_w8524_,
		_w8525_
	);
	LUT2 #(
		.INIT('h2)
	) name8064 (
		\P1_state_reg[0]/NET0131 ,
		_w8525_,
		_w8526_
	);
	LUT2 #(
		.INIT('h1)
	) name8065 (
		_w8501_,
		_w8526_,
		_w8527_
	);
	LUT2 #(
		.INIT('h2)
	) name8066 (
		\P2_reg1_reg[13]/NET0131 ,
		_w1983_,
		_w8528_
	);
	LUT2 #(
		.INIT('h8)
	) name8067 (
		\P2_reg1_reg[13]/NET0131 ,
		_w2024_,
		_w8529_
	);
	LUT2 #(
		.INIT('h1)
	) name8068 (
		_w3733_,
		_w6639_,
		_w8530_
	);
	LUT2 #(
		.INIT('h2)
	) name8069 (
		_w3421_,
		_w8530_,
		_w8531_
	);
	LUT2 #(
		.INIT('h4)
	) name8070 (
		_w7597_,
		_w8531_,
		_w8532_
	);
	LUT2 #(
		.INIT('h1)
	) name8071 (
		_w3733_,
		_w7508_,
		_w8533_
	);
	LUT2 #(
		.INIT('h2)
	) name8072 (
		_w8532_,
		_w8533_,
		_w8534_
	);
	LUT2 #(
		.INIT('h2)
	) name8073 (
		\P2_reg1_reg[13]/NET0131 ,
		_w8534_,
		_w8535_
	);
	LUT2 #(
		.INIT('h8)
	) name8074 (
		_w2893_,
		_w3358_,
		_w8536_
	);
	LUT2 #(
		.INIT('h1)
	) name8075 (
		_w3320_,
		_w7223_,
		_w8537_
	);
	LUT2 #(
		.INIT('h1)
	) name8076 (
		_w8536_,
		_w8537_,
		_w8538_
	);
	LUT2 #(
		.INIT('h8)
	) name8077 (
		_w3355_,
		_w7217_,
		_w8539_
	);
	LUT2 #(
		.INIT('h2)
	) name8078 (
		_w8538_,
		_w8539_,
		_w8540_
	);
	LUT2 #(
		.INIT('h2)
	) name8079 (
		_w3411_,
		_w7205_,
		_w8541_
	);
	LUT2 #(
		.INIT('h4)
	) name8080 (
		_w3177_,
		_w7211_,
		_w8542_
	);
	LUT2 #(
		.INIT('h2)
	) name8081 (
		_w8540_,
		_w8542_,
		_w8543_
	);
	LUT2 #(
		.INIT('h4)
	) name8082 (
		_w8541_,
		_w8543_,
		_w8544_
	);
	LUT2 #(
		.INIT('h2)
	) name8083 (
		_w3733_,
		_w8544_,
		_w8545_
	);
	LUT2 #(
		.INIT('h1)
	) name8084 (
		_w8535_,
		_w8545_,
		_w8546_
	);
	LUT2 #(
		.INIT('h2)
	) name8085 (
		_w2026_,
		_w8546_,
		_w8547_
	);
	LUT2 #(
		.INIT('h1)
	) name8086 (
		_w8529_,
		_w8547_,
		_w8548_
	);
	LUT2 #(
		.INIT('h2)
	) name8087 (
		\P1_state_reg[0]/NET0131 ,
		_w8548_,
		_w8549_
	);
	LUT2 #(
		.INIT('h1)
	) name8088 (
		_w8528_,
		_w8549_,
		_w8550_
	);
	LUT2 #(
		.INIT('h2)
	) name8089 (
		\P2_reg1_reg[23]/NET0131 ,
		_w1983_,
		_w8551_
	);
	LUT2 #(
		.INIT('h8)
	) name8090 (
		\P2_reg1_reg[23]/NET0131 ,
		_w2024_,
		_w8552_
	);
	LUT2 #(
		.INIT('h2)
	) name8091 (
		\P2_reg1_reg[23]/NET0131 ,
		_w3733_,
		_w8553_
	);
	LUT2 #(
		.INIT('h8)
	) name8092 (
		_w3733_,
		_w8331_,
		_w8554_
	);
	LUT2 #(
		.INIT('h1)
	) name8093 (
		_w8553_,
		_w8554_,
		_w8555_
	);
	LUT2 #(
		.INIT('h1)
	) name8094 (
		_w3177_,
		_w8555_,
		_w8556_
	);
	LUT2 #(
		.INIT('h2)
	) name8095 (
		_w3733_,
		_w8380_,
		_w8557_
	);
	LUT2 #(
		.INIT('h2)
	) name8096 (
		_w3733_,
		_w8352_,
		_w8558_
	);
	LUT2 #(
		.INIT('h1)
	) name8097 (
		_w8553_,
		_w8558_,
		_w8559_
	);
	LUT2 #(
		.INIT('h2)
	) name8098 (
		_w3411_,
		_w8559_,
		_w8560_
	);
	LUT2 #(
		.INIT('h2)
	) name8099 (
		\P2_reg1_reg[23]/NET0131 ,
		_w8532_,
		_w8561_
	);
	LUT2 #(
		.INIT('h1)
	) name8100 (
		_w8560_,
		_w8561_,
		_w8562_
	);
	LUT2 #(
		.INIT('h4)
	) name8101 (
		_w8557_,
		_w8562_,
		_w8563_
	);
	LUT2 #(
		.INIT('h4)
	) name8102 (
		_w8556_,
		_w8563_,
		_w8564_
	);
	LUT2 #(
		.INIT('h2)
	) name8103 (
		_w2026_,
		_w8564_,
		_w8565_
	);
	LUT2 #(
		.INIT('h1)
	) name8104 (
		_w8552_,
		_w8565_,
		_w8566_
	);
	LUT2 #(
		.INIT('h2)
	) name8105 (
		\P1_state_reg[0]/NET0131 ,
		_w8566_,
		_w8567_
	);
	LUT2 #(
		.INIT('h1)
	) name8106 (
		_w8551_,
		_w8567_,
		_w8568_
	);
	LUT2 #(
		.INIT('h2)
	) name8107 (
		\P1_reg0_reg[10]/NET0131 ,
		_w3435_,
		_w8569_
	);
	LUT2 #(
		.INIT('h8)
	) name8108 (
		\P1_reg0_reg[10]/NET0131 ,
		_w3448_,
		_w8570_
	);
	LUT2 #(
		.INIT('h8)
	) name8109 (
		_w4396_,
		_w8423_,
		_w8571_
	);
	LUT2 #(
		.INIT('h2)
	) name8110 (
		\P1_reg0_reg[10]/NET0131 ,
		_w4396_,
		_w8572_
	);
	LUT2 #(
		.INIT('h8)
	) name8111 (
		_w4396_,
		_w7092_,
		_w8573_
	);
	LUT2 #(
		.INIT('h1)
	) name8112 (
		_w8572_,
		_w8573_,
		_w8574_
	);
	LUT2 #(
		.INIT('h1)
	) name8113 (
		_w3563_,
		_w8574_,
		_w8575_
	);
	LUT2 #(
		.INIT('h8)
	) name8114 (
		_w4396_,
		_w7086_,
		_w8576_
	);
	LUT2 #(
		.INIT('h1)
	) name8115 (
		_w8572_,
		_w8576_,
		_w8577_
	);
	LUT2 #(
		.INIT('h2)
	) name8116 (
		_w1936_,
		_w8577_,
		_w8578_
	);
	LUT2 #(
		.INIT('h2)
	) name8117 (
		_w4396_,
		_w7078_,
		_w8579_
	);
	LUT2 #(
		.INIT('h1)
	) name8118 (
		_w8572_,
		_w8579_,
		_w8580_
	);
	LUT2 #(
		.INIT('h1)
	) name8119 (
		_w3677_,
		_w8580_,
		_w8581_
	);
	LUT2 #(
		.INIT('h8)
	) name8120 (
		_w4396_,
		_w7097_,
		_w8582_
	);
	LUT2 #(
		.INIT('h1)
	) name8121 (
		_w8572_,
		_w8582_,
		_w8583_
	);
	LUT2 #(
		.INIT('h2)
	) name8122 (
		_w3712_,
		_w8583_,
		_w8584_
	);
	LUT2 #(
		.INIT('h2)
	) name8123 (
		\P1_reg0_reg[10]/NET0131 ,
		_w4493_,
		_w8585_
	);
	LUT2 #(
		.INIT('h1)
	) name8124 (
		_w8571_,
		_w8585_,
		_w8586_
	);
	LUT2 #(
		.INIT('h4)
	) name8125 (
		_w8584_,
		_w8586_,
		_w8587_
	);
	LUT2 #(
		.INIT('h4)
	) name8126 (
		_w8575_,
		_w8587_,
		_w8588_
	);
	LUT2 #(
		.INIT('h1)
	) name8127 (
		_w8578_,
		_w8581_,
		_w8589_
	);
	LUT2 #(
		.INIT('h8)
	) name8128 (
		_w8588_,
		_w8589_,
		_w8590_
	);
	LUT2 #(
		.INIT('h2)
	) name8129 (
		_w3450_,
		_w8590_,
		_w8591_
	);
	LUT2 #(
		.INIT('h1)
	) name8130 (
		_w8570_,
		_w8591_,
		_w8592_
	);
	LUT2 #(
		.INIT('h2)
	) name8131 (
		\P1_state_reg[0]/NET0131 ,
		_w8592_,
		_w8593_
	);
	LUT2 #(
		.INIT('h1)
	) name8132 (
		_w8569_,
		_w8593_,
		_w8594_
	);
	LUT2 #(
		.INIT('h2)
	) name8133 (
		\P2_reg1_reg[9]/NET0131 ,
		_w1983_,
		_w8595_
	);
	LUT2 #(
		.INIT('h8)
	) name8134 (
		\P2_reg1_reg[9]/NET0131 ,
		_w2024_,
		_w8596_
	);
	LUT2 #(
		.INIT('h2)
	) name8135 (
		\P2_reg1_reg[9]/NET0131 ,
		_w8532_,
		_w8597_
	);
	LUT2 #(
		.INIT('h2)
	) name8136 (
		\P2_reg1_reg[9]/NET0131 ,
		_w3733_,
		_w8598_
	);
	LUT2 #(
		.INIT('h8)
	) name8137 (
		_w3733_,
		_w7248_,
		_w8599_
	);
	LUT2 #(
		.INIT('h1)
	) name8138 (
		_w8598_,
		_w8599_,
		_w8600_
	);
	LUT2 #(
		.INIT('h2)
	) name8139 (
		_w3411_,
		_w8600_,
		_w8601_
	);
	LUT2 #(
		.INIT('h2)
	) name8140 (
		_w3733_,
		_w7254_,
		_w8602_
	);
	LUT2 #(
		.INIT('h1)
	) name8141 (
		_w8598_,
		_w8602_,
		_w8603_
	);
	LUT2 #(
		.INIT('h1)
	) name8142 (
		_w3177_,
		_w8603_,
		_w8604_
	);
	LUT2 #(
		.INIT('h2)
	) name8143 (
		_w3733_,
		_w8492_,
		_w8605_
	);
	LUT2 #(
		.INIT('h1)
	) name8144 (
		_w8597_,
		_w8605_,
		_w8606_
	);
	LUT2 #(
		.INIT('h4)
	) name8145 (
		_w8604_,
		_w8606_,
		_w8607_
	);
	LUT2 #(
		.INIT('h4)
	) name8146 (
		_w8601_,
		_w8607_,
		_w8608_
	);
	LUT2 #(
		.INIT('h2)
	) name8147 (
		_w2026_,
		_w8608_,
		_w8609_
	);
	LUT2 #(
		.INIT('h1)
	) name8148 (
		_w8596_,
		_w8609_,
		_w8610_
	);
	LUT2 #(
		.INIT('h2)
	) name8149 (
		\P1_state_reg[0]/NET0131 ,
		_w8610_,
		_w8611_
	);
	LUT2 #(
		.INIT('h1)
	) name8150 (
		_w8595_,
		_w8611_,
		_w8612_
	);
	LUT2 #(
		.INIT('h2)
	) name8151 (
		\P2_reg2_reg[10]/NET0131 ,
		_w1983_,
		_w8613_
	);
	LUT2 #(
		.INIT('h8)
	) name8152 (
		\P2_reg2_reg[10]/NET0131 ,
		_w2024_,
		_w8614_
	);
	LUT2 #(
		.INIT('h8)
	) name8153 (
		_w3758_,
		_w8503_,
		_w8615_
	);
	LUT2 #(
		.INIT('h2)
	) name8154 (
		\P2_reg2_reg[10]/NET0131 ,
		_w3758_,
		_w8616_
	);
	LUT2 #(
		.INIT('h8)
	) name8155 (
		_w3758_,
		_w7163_,
		_w8617_
	);
	LUT2 #(
		.INIT('h1)
	) name8156 (
		_w8616_,
		_w8617_,
		_w8618_
	);
	LUT2 #(
		.INIT('h2)
	) name8157 (
		_w3411_,
		_w8618_,
		_w8619_
	);
	LUT2 #(
		.INIT('h2)
	) name8158 (
		_w3758_,
		_w7169_,
		_w8620_
	);
	LUT2 #(
		.INIT('h1)
	) name8159 (
		_w8616_,
		_w8620_,
		_w8621_
	);
	LUT2 #(
		.INIT('h1)
	) name8160 (
		_w3177_,
		_w8621_,
		_w8622_
	);
	LUT2 #(
		.INIT('h8)
	) name8161 (
		_w3758_,
		_w7175_,
		_w8623_
	);
	LUT2 #(
		.INIT('h1)
	) name8162 (
		_w8616_,
		_w8623_,
		_w8624_
	);
	LUT2 #(
		.INIT('h1)
	) name8163 (
		_w3320_,
		_w8624_,
		_w8625_
	);
	LUT2 #(
		.INIT('h8)
	) name8164 (
		_w3758_,
		_w7181_,
		_w8626_
	);
	LUT2 #(
		.INIT('h1)
	) name8165 (
		_w8616_,
		_w8626_,
		_w8627_
	);
	LUT2 #(
		.INIT('h2)
	) name8166 (
		_w3355_,
		_w8627_,
		_w8628_
	);
	LUT2 #(
		.INIT('h8)
	) name8167 (
		_w2735_,
		_w3420_,
		_w8629_
	);
	LUT2 #(
		.INIT('h2)
	) name8168 (
		\P2_reg2_reg[10]/NET0131 ,
		_w3774_,
		_w8630_
	);
	LUT2 #(
		.INIT('h1)
	) name8169 (
		_w8615_,
		_w8629_,
		_w8631_
	);
	LUT2 #(
		.INIT('h4)
	) name8170 (
		_w8630_,
		_w8631_,
		_w8632_
	);
	LUT2 #(
		.INIT('h4)
	) name8171 (
		_w8628_,
		_w8632_,
		_w8633_
	);
	LUT2 #(
		.INIT('h4)
	) name8172 (
		_w8622_,
		_w8633_,
		_w8634_
	);
	LUT2 #(
		.INIT('h4)
	) name8173 (
		_w8625_,
		_w8634_,
		_w8635_
	);
	LUT2 #(
		.INIT('h4)
	) name8174 (
		_w8619_,
		_w8635_,
		_w8636_
	);
	LUT2 #(
		.INIT('h2)
	) name8175 (
		_w2026_,
		_w8636_,
		_w8637_
	);
	LUT2 #(
		.INIT('h1)
	) name8176 (
		_w8614_,
		_w8637_,
		_w8638_
	);
	LUT2 #(
		.INIT('h2)
	) name8177 (
		\P1_state_reg[0]/NET0131 ,
		_w8638_,
		_w8639_
	);
	LUT2 #(
		.INIT('h1)
	) name8178 (
		_w8613_,
		_w8639_,
		_w8640_
	);
	LUT2 #(
		.INIT('h2)
	) name8179 (
		\P2_reg2_reg[13]/NET0131 ,
		_w1983_,
		_w8641_
	);
	LUT2 #(
		.INIT('h8)
	) name8180 (
		\P2_reg2_reg[13]/NET0131 ,
		_w2024_,
		_w8642_
	);
	LUT2 #(
		.INIT('h2)
	) name8181 (
		\P2_reg2_reg[13]/NET0131 ,
		_w7770_,
		_w8643_
	);
	LUT2 #(
		.INIT('h2)
	) name8182 (
		\P2_reg2_reg[13]/NET0131 ,
		_w3758_,
		_w8644_
	);
	LUT2 #(
		.INIT('h2)
	) name8183 (
		_w3758_,
		_w7205_,
		_w8645_
	);
	LUT2 #(
		.INIT('h1)
	) name8184 (
		_w8644_,
		_w8645_,
		_w8646_
	);
	LUT2 #(
		.INIT('h2)
	) name8185 (
		_w3411_,
		_w8646_,
		_w8647_
	);
	LUT2 #(
		.INIT('h8)
	) name8186 (
		_w3758_,
		_w7211_,
		_w8648_
	);
	LUT2 #(
		.INIT('h1)
	) name8187 (
		_w8644_,
		_w8648_,
		_w8649_
	);
	LUT2 #(
		.INIT('h1)
	) name8188 (
		_w3177_,
		_w8649_,
		_w8650_
	);
	LUT2 #(
		.INIT('h8)
	) name8189 (
		_w3758_,
		_w7217_,
		_w8651_
	);
	LUT2 #(
		.INIT('h1)
	) name8190 (
		_w8644_,
		_w8651_,
		_w8652_
	);
	LUT2 #(
		.INIT('h2)
	) name8191 (
		_w3355_,
		_w8652_,
		_w8653_
	);
	LUT2 #(
		.INIT('h2)
	) name8192 (
		_w3758_,
		_w8538_,
		_w8654_
	);
	LUT2 #(
		.INIT('h8)
	) name8193 (
		_w2874_,
		_w3420_,
		_w8655_
	);
	LUT2 #(
		.INIT('h1)
	) name8194 (
		_w8643_,
		_w8655_,
		_w8656_
	);
	LUT2 #(
		.INIT('h4)
	) name8195 (
		_w8654_,
		_w8656_,
		_w8657_
	);
	LUT2 #(
		.INIT('h4)
	) name8196 (
		_w8653_,
		_w8657_,
		_w8658_
	);
	LUT2 #(
		.INIT('h4)
	) name8197 (
		_w8650_,
		_w8658_,
		_w8659_
	);
	LUT2 #(
		.INIT('h4)
	) name8198 (
		_w8647_,
		_w8659_,
		_w8660_
	);
	LUT2 #(
		.INIT('h2)
	) name8199 (
		_w2026_,
		_w8660_,
		_w8661_
	);
	LUT2 #(
		.INIT('h1)
	) name8200 (
		_w8642_,
		_w8661_,
		_w8662_
	);
	LUT2 #(
		.INIT('h2)
	) name8201 (
		\P1_state_reg[0]/NET0131 ,
		_w8662_,
		_w8663_
	);
	LUT2 #(
		.INIT('h1)
	) name8202 (
		_w8641_,
		_w8663_,
		_w8664_
	);
	LUT2 #(
		.INIT('h2)
	) name8203 (
		\P1_reg2_reg[9]/NET0131 ,
		_w3435_,
		_w8665_
	);
	LUT2 #(
		.INIT('h8)
	) name8204 (
		\P1_reg2_reg[9]/NET0131 ,
		_w3448_,
		_w8666_
	);
	LUT2 #(
		.INIT('h8)
	) name8205 (
		_w3466_,
		_w8396_,
		_w8667_
	);
	LUT2 #(
		.INIT('h2)
	) name8206 (
		\P1_reg2_reg[9]/NET0131 ,
		_w3466_,
		_w8668_
	);
	LUT2 #(
		.INIT('h8)
	) name8207 (
		_w3466_,
		_w7294_,
		_w8669_
	);
	LUT2 #(
		.INIT('h1)
	) name8208 (
		_w8668_,
		_w8669_,
		_w8670_
	);
	LUT2 #(
		.INIT('h1)
	) name8209 (
		_w3563_,
		_w8670_,
		_w8671_
	);
	LUT2 #(
		.INIT('h2)
	) name8210 (
		_w3466_,
		_w7288_,
		_w8672_
	);
	LUT2 #(
		.INIT('h1)
	) name8211 (
		_w8668_,
		_w8672_,
		_w8673_
	);
	LUT2 #(
		.INIT('h1)
	) name8212 (
		_w3677_,
		_w8673_,
		_w8674_
	);
	LUT2 #(
		.INIT('h8)
	) name8213 (
		_w3466_,
		_w7300_,
		_w8675_
	);
	LUT2 #(
		.INIT('h1)
	) name8214 (
		_w8668_,
		_w8675_,
		_w8676_
	);
	LUT2 #(
		.INIT('h2)
	) name8215 (
		_w3712_,
		_w8676_,
		_w8677_
	);
	LUT2 #(
		.INIT('h2)
	) name8216 (
		_w3466_,
		_w7310_,
		_w8678_
	);
	LUT2 #(
		.INIT('h1)
	) name8217 (
		_w8668_,
		_w8678_,
		_w8679_
	);
	LUT2 #(
		.INIT('h2)
	) name8218 (
		_w1936_,
		_w8679_,
		_w8680_
	);
	LUT2 #(
		.INIT('h8)
	) name8219 (
		_w1239_,
		_w1763_,
		_w8681_
	);
	LUT2 #(
		.INIT('h2)
	) name8220 (
		\P1_reg2_reg[9]/NET0131 ,
		_w3718_,
		_w8682_
	);
	LUT2 #(
		.INIT('h1)
	) name8221 (
		_w8667_,
		_w8681_,
		_w8683_
	);
	LUT2 #(
		.INIT('h4)
	) name8222 (
		_w8682_,
		_w8683_,
		_w8684_
	);
	LUT2 #(
		.INIT('h4)
	) name8223 (
		_w8677_,
		_w8684_,
		_w8685_
	);
	LUT2 #(
		.INIT('h4)
	) name8224 (
		_w8671_,
		_w8685_,
		_w8686_
	);
	LUT2 #(
		.INIT('h4)
	) name8225 (
		_w8674_,
		_w8686_,
		_w8687_
	);
	LUT2 #(
		.INIT('h4)
	) name8226 (
		_w8680_,
		_w8687_,
		_w8688_
	);
	LUT2 #(
		.INIT('h2)
	) name8227 (
		_w3450_,
		_w8688_,
		_w8689_
	);
	LUT2 #(
		.INIT('h1)
	) name8228 (
		_w8666_,
		_w8689_,
		_w8690_
	);
	LUT2 #(
		.INIT('h2)
	) name8229 (
		\P1_state_reg[0]/NET0131 ,
		_w8690_,
		_w8691_
	);
	LUT2 #(
		.INIT('h1)
	) name8230 (
		_w8665_,
		_w8691_,
		_w8692_
	);
	LUT2 #(
		.INIT('h2)
	) name8231 (
		\P2_reg2_reg[23]/NET0131 ,
		_w1983_,
		_w8693_
	);
	LUT2 #(
		.INIT('h8)
	) name8232 (
		\P2_reg2_reg[23]/NET0131 ,
		_w2024_,
		_w8694_
	);
	LUT2 #(
		.INIT('h2)
	) name8233 (
		\P2_reg2_reg[23]/NET0131 ,
		_w3758_,
		_w8695_
	);
	LUT2 #(
		.INIT('h8)
	) name8234 (
		_w3758_,
		_w8331_,
		_w8696_
	);
	LUT2 #(
		.INIT('h1)
	) name8235 (
		_w8695_,
		_w8696_,
		_w8697_
	);
	LUT2 #(
		.INIT('h1)
	) name8236 (
		_w3177_,
		_w8697_,
		_w8698_
	);
	LUT2 #(
		.INIT('h2)
	) name8237 (
		_w3758_,
		_w8380_,
		_w8699_
	);
	LUT2 #(
		.INIT('h8)
	) name8238 (
		_w3084_,
		_w3420_,
		_w8700_
	);
	LUT2 #(
		.INIT('h2)
	) name8239 (
		_w3758_,
		_w8352_,
		_w8701_
	);
	LUT2 #(
		.INIT('h1)
	) name8240 (
		_w8695_,
		_w8701_,
		_w8702_
	);
	LUT2 #(
		.INIT('h2)
	) name8241 (
		_w3411_,
		_w8702_,
		_w8703_
	);
	LUT2 #(
		.INIT('h4)
	) name8242 (
		_w4382_,
		_w7770_,
		_w8704_
	);
	LUT2 #(
		.INIT('h2)
	) name8243 (
		\P2_reg2_reg[23]/NET0131 ,
		_w8704_,
		_w8705_
	);
	LUT2 #(
		.INIT('h1)
	) name8244 (
		_w8700_,
		_w8705_,
		_w8706_
	);
	LUT2 #(
		.INIT('h4)
	) name8245 (
		_w8703_,
		_w8706_,
		_w8707_
	);
	LUT2 #(
		.INIT('h4)
	) name8246 (
		_w8699_,
		_w8707_,
		_w8708_
	);
	LUT2 #(
		.INIT('h4)
	) name8247 (
		_w8698_,
		_w8708_,
		_w8709_
	);
	LUT2 #(
		.INIT('h2)
	) name8248 (
		_w2026_,
		_w8709_,
		_w8710_
	);
	LUT2 #(
		.INIT('h1)
	) name8249 (
		_w8694_,
		_w8710_,
		_w8711_
	);
	LUT2 #(
		.INIT('h2)
	) name8250 (
		\P1_state_reg[0]/NET0131 ,
		_w8711_,
		_w8712_
	);
	LUT2 #(
		.INIT('h1)
	) name8251 (
		_w8693_,
		_w8712_,
		_w8713_
	);
	LUT2 #(
		.INIT('h2)
	) name8252 (
		\P2_reg2_reg[9]/NET0131 ,
		_w1983_,
		_w8714_
	);
	LUT2 #(
		.INIT('h8)
	) name8253 (
		\P2_reg2_reg[9]/NET0131 ,
		_w2024_,
		_w8715_
	);
	LUT2 #(
		.INIT('h8)
	) name8254 (
		_w3758_,
		_w8489_,
		_w8716_
	);
	LUT2 #(
		.INIT('h2)
	) name8255 (
		\P2_reg2_reg[9]/NET0131 ,
		_w3758_,
		_w8717_
	);
	LUT2 #(
		.INIT('h8)
	) name8256 (
		_w3758_,
		_w7248_,
		_w8718_
	);
	LUT2 #(
		.INIT('h1)
	) name8257 (
		_w8717_,
		_w8718_,
		_w8719_
	);
	LUT2 #(
		.INIT('h2)
	) name8258 (
		_w3411_,
		_w8719_,
		_w8720_
	);
	LUT2 #(
		.INIT('h2)
	) name8259 (
		_w3758_,
		_w7254_,
		_w8721_
	);
	LUT2 #(
		.INIT('h1)
	) name8260 (
		_w8717_,
		_w8721_,
		_w8722_
	);
	LUT2 #(
		.INIT('h1)
	) name8261 (
		_w3177_,
		_w8722_,
		_w8723_
	);
	LUT2 #(
		.INIT('h8)
	) name8262 (
		_w3758_,
		_w7260_,
		_w8724_
	);
	LUT2 #(
		.INIT('h1)
	) name8263 (
		_w8717_,
		_w8724_,
		_w8725_
	);
	LUT2 #(
		.INIT('h2)
	) name8264 (
		_w3355_,
		_w8725_,
		_w8726_
	);
	LUT2 #(
		.INIT('h8)
	) name8265 (
		_w3758_,
		_w7266_,
		_w8727_
	);
	LUT2 #(
		.INIT('h1)
	) name8266 (
		_w8717_,
		_w8727_,
		_w8728_
	);
	LUT2 #(
		.INIT('h1)
	) name8267 (
		_w3320_,
		_w8728_,
		_w8729_
	);
	LUT2 #(
		.INIT('h8)
	) name8268 (
		_w2760_,
		_w3420_,
		_w8730_
	);
	LUT2 #(
		.INIT('h2)
	) name8269 (
		\P2_reg2_reg[9]/NET0131 ,
		_w3774_,
		_w8731_
	);
	LUT2 #(
		.INIT('h1)
	) name8270 (
		_w8716_,
		_w8730_,
		_w8732_
	);
	LUT2 #(
		.INIT('h4)
	) name8271 (
		_w8731_,
		_w8732_,
		_w8733_
	);
	LUT2 #(
		.INIT('h4)
	) name8272 (
		_w8729_,
		_w8733_,
		_w8734_
	);
	LUT2 #(
		.INIT('h4)
	) name8273 (
		_w8726_,
		_w8734_,
		_w8735_
	);
	LUT2 #(
		.INIT('h4)
	) name8274 (
		_w8723_,
		_w8735_,
		_w8736_
	);
	LUT2 #(
		.INIT('h4)
	) name8275 (
		_w8720_,
		_w8736_,
		_w8737_
	);
	LUT2 #(
		.INIT('h2)
	) name8276 (
		_w2026_,
		_w8737_,
		_w8738_
	);
	LUT2 #(
		.INIT('h1)
	) name8277 (
		_w8715_,
		_w8738_,
		_w8739_
	);
	LUT2 #(
		.INIT('h2)
	) name8278 (
		\P1_state_reg[0]/NET0131 ,
		_w8739_,
		_w8740_
	);
	LUT2 #(
		.INIT('h1)
	) name8279 (
		_w8714_,
		_w8740_,
		_w8741_
	);
	LUT2 #(
		.INIT('h2)
	) name8280 (
		\P1_reg0_reg[13]/NET0131 ,
		_w3435_,
		_w8742_
	);
	LUT2 #(
		.INIT('h8)
	) name8281 (
		\P1_reg0_reg[13]/NET0131 ,
		_w3448_,
		_w8743_
	);
	LUT2 #(
		.INIT('h8)
	) name8282 (
		_w4396_,
		_w8467_,
		_w8744_
	);
	LUT2 #(
		.INIT('h2)
	) name8283 (
		\P1_reg0_reg[13]/NET0131 ,
		_w4396_,
		_w8745_
	);
	LUT2 #(
		.INIT('h2)
	) name8284 (
		_w4396_,
		_w7119_,
		_w8746_
	);
	LUT2 #(
		.INIT('h1)
	) name8285 (
		_w8745_,
		_w8746_,
		_w8747_
	);
	LUT2 #(
		.INIT('h1)
	) name8286 (
		_w3677_,
		_w8747_,
		_w8748_
	);
	LUT2 #(
		.INIT('h8)
	) name8287 (
		_w4396_,
		_w7125_,
		_w8749_
	);
	LUT2 #(
		.INIT('h1)
	) name8288 (
		_w8745_,
		_w8749_,
		_w8750_
	);
	LUT2 #(
		.INIT('h1)
	) name8289 (
		_w3563_,
		_w8750_,
		_w8751_
	);
	LUT2 #(
		.INIT('h8)
	) name8290 (
		_w4396_,
		_w7134_,
		_w8752_
	);
	LUT2 #(
		.INIT('h1)
	) name8291 (
		_w8745_,
		_w8752_,
		_w8753_
	);
	LUT2 #(
		.INIT('h2)
	) name8292 (
		_w1936_,
		_w8753_,
		_w8754_
	);
	LUT2 #(
		.INIT('h8)
	) name8293 (
		_w4396_,
		_w7139_,
		_w8755_
	);
	LUT2 #(
		.INIT('h1)
	) name8294 (
		_w8745_,
		_w8755_,
		_w8756_
	);
	LUT2 #(
		.INIT('h2)
	) name8295 (
		_w3712_,
		_w8756_,
		_w8757_
	);
	LUT2 #(
		.INIT('h2)
	) name8296 (
		\P1_reg0_reg[13]/NET0131 ,
		_w4493_,
		_w8758_
	);
	LUT2 #(
		.INIT('h1)
	) name8297 (
		_w8744_,
		_w8758_,
		_w8759_
	);
	LUT2 #(
		.INIT('h4)
	) name8298 (
		_w8757_,
		_w8759_,
		_w8760_
	);
	LUT2 #(
		.INIT('h4)
	) name8299 (
		_w8748_,
		_w8760_,
		_w8761_
	);
	LUT2 #(
		.INIT('h1)
	) name8300 (
		_w8751_,
		_w8754_,
		_w8762_
	);
	LUT2 #(
		.INIT('h8)
	) name8301 (
		_w8761_,
		_w8762_,
		_w8763_
	);
	LUT2 #(
		.INIT('h2)
	) name8302 (
		_w3450_,
		_w8763_,
		_w8764_
	);
	LUT2 #(
		.INIT('h1)
	) name8303 (
		_w8743_,
		_w8764_,
		_w8765_
	);
	LUT2 #(
		.INIT('h2)
	) name8304 (
		\P1_state_reg[0]/NET0131 ,
		_w8765_,
		_w8766_
	);
	LUT2 #(
		.INIT('h1)
	) name8305 (
		_w8742_,
		_w8766_,
		_w8767_
	);
	LUT2 #(
		.INIT('h2)
	) name8306 (
		\P1_reg0_reg[23]/NET0131 ,
		_w3435_,
		_w8768_
	);
	LUT2 #(
		.INIT('h8)
	) name8307 (
		\P1_reg0_reg[23]/NET0131 ,
		_w3448_,
		_w8769_
	);
	LUT2 #(
		.INIT('h2)
	) name8308 (
		\P1_reg0_reg[23]/NET0131 ,
		_w4396_,
		_w8770_
	);
	LUT2 #(
		.INIT('h2)
	) name8309 (
		_w4396_,
		_w7422_,
		_w8771_
	);
	LUT2 #(
		.INIT('h1)
	) name8310 (
		_w8770_,
		_w8771_,
		_w8772_
	);
	LUT2 #(
		.INIT('h1)
	) name8311 (
		_w3677_,
		_w8772_,
		_w8773_
	);
	LUT2 #(
		.INIT('h2)
	) name8312 (
		_w4396_,
		_w7435_,
		_w8774_
	);
	LUT2 #(
		.INIT('h1)
	) name8313 (
		_w8770_,
		_w8774_,
		_w8775_
	);
	LUT2 #(
		.INIT('h1)
	) name8314 (
		_w3563_,
		_w8775_,
		_w8776_
	);
	LUT2 #(
		.INIT('h1)
	) name8315 (
		_w7450_,
		_w7653_,
		_w8777_
	);
	LUT2 #(
		.INIT('h2)
	) name8316 (
		_w4396_,
		_w8777_,
		_w8778_
	);
	LUT2 #(
		.INIT('h8)
	) name8317 (
		_w4396_,
		_w7444_,
		_w8779_
	);
	LUT2 #(
		.INIT('h1)
	) name8318 (
		_w8770_,
		_w8779_,
		_w8780_
	);
	LUT2 #(
		.INIT('h2)
	) name8319 (
		_w1936_,
		_w8780_,
		_w8781_
	);
	LUT2 #(
		.INIT('h2)
	) name8320 (
		\P1_reg0_reg[23]/NET0131 ,
		_w4494_,
		_w8782_
	);
	LUT2 #(
		.INIT('h1)
	) name8321 (
		_w8778_,
		_w8782_,
		_w8783_
	);
	LUT2 #(
		.INIT('h4)
	) name8322 (
		_w8781_,
		_w8783_,
		_w8784_
	);
	LUT2 #(
		.INIT('h4)
	) name8323 (
		_w8773_,
		_w8784_,
		_w8785_
	);
	LUT2 #(
		.INIT('h4)
	) name8324 (
		_w8776_,
		_w8785_,
		_w8786_
	);
	LUT2 #(
		.INIT('h2)
	) name8325 (
		_w3450_,
		_w8786_,
		_w8787_
	);
	LUT2 #(
		.INIT('h1)
	) name8326 (
		_w8769_,
		_w8787_,
		_w8788_
	);
	LUT2 #(
		.INIT('h2)
	) name8327 (
		\P1_state_reg[0]/NET0131 ,
		_w8788_,
		_w8789_
	);
	LUT2 #(
		.INIT('h1)
	) name8328 (
		_w8768_,
		_w8789_,
		_w8790_
	);
	LUT2 #(
		.INIT('h2)
	) name8329 (
		\P1_reg0_reg[9]/NET0131 ,
		_w3435_,
		_w8791_
	);
	LUT2 #(
		.INIT('h8)
	) name8330 (
		\P1_reg0_reg[9]/NET0131 ,
		_w3448_,
		_w8792_
	);
	LUT2 #(
		.INIT('h8)
	) name8331 (
		_w4396_,
		_w8396_,
		_w8793_
	);
	LUT2 #(
		.INIT('h2)
	) name8332 (
		\P1_reg0_reg[9]/NET0131 ,
		_w4396_,
		_w8794_
	);
	LUT2 #(
		.INIT('h8)
	) name8333 (
		_w4396_,
		_w7294_,
		_w8795_
	);
	LUT2 #(
		.INIT('h1)
	) name8334 (
		_w8794_,
		_w8795_,
		_w8796_
	);
	LUT2 #(
		.INIT('h1)
	) name8335 (
		_w3563_,
		_w8796_,
		_w8797_
	);
	LUT2 #(
		.INIT('h2)
	) name8336 (
		_w4396_,
		_w7288_,
		_w8798_
	);
	LUT2 #(
		.INIT('h1)
	) name8337 (
		_w8794_,
		_w8798_,
		_w8799_
	);
	LUT2 #(
		.INIT('h1)
	) name8338 (
		_w3677_,
		_w8799_,
		_w8800_
	);
	LUT2 #(
		.INIT('h8)
	) name8339 (
		_w4396_,
		_w7300_,
		_w8801_
	);
	LUT2 #(
		.INIT('h1)
	) name8340 (
		_w8794_,
		_w8801_,
		_w8802_
	);
	LUT2 #(
		.INIT('h2)
	) name8341 (
		_w3712_,
		_w8802_,
		_w8803_
	);
	LUT2 #(
		.INIT('h2)
	) name8342 (
		_w4396_,
		_w7310_,
		_w8804_
	);
	LUT2 #(
		.INIT('h1)
	) name8343 (
		_w8794_,
		_w8804_,
		_w8805_
	);
	LUT2 #(
		.INIT('h2)
	) name8344 (
		_w1936_,
		_w8805_,
		_w8806_
	);
	LUT2 #(
		.INIT('h2)
	) name8345 (
		\P1_reg0_reg[9]/NET0131 ,
		_w4493_,
		_w8807_
	);
	LUT2 #(
		.INIT('h1)
	) name8346 (
		_w8793_,
		_w8807_,
		_w8808_
	);
	LUT2 #(
		.INIT('h4)
	) name8347 (
		_w8803_,
		_w8808_,
		_w8809_
	);
	LUT2 #(
		.INIT('h4)
	) name8348 (
		_w8797_,
		_w8809_,
		_w8810_
	);
	LUT2 #(
		.INIT('h4)
	) name8349 (
		_w8800_,
		_w8810_,
		_w8811_
	);
	LUT2 #(
		.INIT('h4)
	) name8350 (
		_w8806_,
		_w8811_,
		_w8812_
	);
	LUT2 #(
		.INIT('h2)
	) name8351 (
		_w3450_,
		_w8812_,
		_w8813_
	);
	LUT2 #(
		.INIT('h1)
	) name8352 (
		_w8792_,
		_w8813_,
		_w8814_
	);
	LUT2 #(
		.INIT('h2)
	) name8353 (
		\P1_state_reg[0]/NET0131 ,
		_w8814_,
		_w8815_
	);
	LUT2 #(
		.INIT('h1)
	) name8354 (
		_w8791_,
		_w8815_,
		_w8816_
	);
	LUT2 #(
		.INIT('h2)
	) name8355 (
		\P1_reg1_reg[10]/NET0131 ,
		_w3435_,
		_w8817_
	);
	LUT2 #(
		.INIT('h8)
	) name8356 (
		\P1_reg1_reg[10]/NET0131 ,
		_w3448_,
		_w8818_
	);
	LUT2 #(
		.INIT('h8)
	) name8357 (
		_w4532_,
		_w8423_,
		_w8819_
	);
	LUT2 #(
		.INIT('h2)
	) name8358 (
		\P1_reg1_reg[10]/NET0131 ,
		_w4532_,
		_w8820_
	);
	LUT2 #(
		.INIT('h8)
	) name8359 (
		_w4532_,
		_w7092_,
		_w8821_
	);
	LUT2 #(
		.INIT('h1)
	) name8360 (
		_w8820_,
		_w8821_,
		_w8822_
	);
	LUT2 #(
		.INIT('h1)
	) name8361 (
		_w3563_,
		_w8822_,
		_w8823_
	);
	LUT2 #(
		.INIT('h8)
	) name8362 (
		_w4532_,
		_w7086_,
		_w8824_
	);
	LUT2 #(
		.INIT('h1)
	) name8363 (
		_w8820_,
		_w8824_,
		_w8825_
	);
	LUT2 #(
		.INIT('h2)
	) name8364 (
		_w1936_,
		_w8825_,
		_w8826_
	);
	LUT2 #(
		.INIT('h2)
	) name8365 (
		_w4532_,
		_w7078_,
		_w8827_
	);
	LUT2 #(
		.INIT('h1)
	) name8366 (
		_w8820_,
		_w8827_,
		_w8828_
	);
	LUT2 #(
		.INIT('h1)
	) name8367 (
		_w3677_,
		_w8828_,
		_w8829_
	);
	LUT2 #(
		.INIT('h8)
	) name8368 (
		_w4532_,
		_w7097_,
		_w8830_
	);
	LUT2 #(
		.INIT('h1)
	) name8369 (
		_w8820_,
		_w8830_,
		_w8831_
	);
	LUT2 #(
		.INIT('h2)
	) name8370 (
		_w3712_,
		_w8831_,
		_w8832_
	);
	LUT2 #(
		.INIT('h2)
	) name8371 (
		\P1_reg1_reg[10]/NET0131 ,
		_w4541_,
		_w8833_
	);
	LUT2 #(
		.INIT('h1)
	) name8372 (
		_w8819_,
		_w8833_,
		_w8834_
	);
	LUT2 #(
		.INIT('h4)
	) name8373 (
		_w8832_,
		_w8834_,
		_w8835_
	);
	LUT2 #(
		.INIT('h4)
	) name8374 (
		_w8823_,
		_w8835_,
		_w8836_
	);
	LUT2 #(
		.INIT('h1)
	) name8375 (
		_w8826_,
		_w8829_,
		_w8837_
	);
	LUT2 #(
		.INIT('h8)
	) name8376 (
		_w8836_,
		_w8837_,
		_w8838_
	);
	LUT2 #(
		.INIT('h2)
	) name8377 (
		_w3450_,
		_w8838_,
		_w8839_
	);
	LUT2 #(
		.INIT('h1)
	) name8378 (
		_w8818_,
		_w8839_,
		_w8840_
	);
	LUT2 #(
		.INIT('h2)
	) name8379 (
		\P1_state_reg[0]/NET0131 ,
		_w8840_,
		_w8841_
	);
	LUT2 #(
		.INIT('h1)
	) name8380 (
		_w8817_,
		_w8841_,
		_w8842_
	);
	LUT2 #(
		.INIT('h2)
	) name8381 (
		\P1_reg1_reg[13]/NET0131 ,
		_w3435_,
		_w8843_
	);
	LUT2 #(
		.INIT('h8)
	) name8382 (
		\P1_reg1_reg[13]/NET0131 ,
		_w3448_,
		_w8844_
	);
	LUT2 #(
		.INIT('h8)
	) name8383 (
		_w4532_,
		_w8467_,
		_w8845_
	);
	LUT2 #(
		.INIT('h2)
	) name8384 (
		\P1_reg1_reg[13]/NET0131 ,
		_w4532_,
		_w8846_
	);
	LUT2 #(
		.INIT('h2)
	) name8385 (
		_w4532_,
		_w7119_,
		_w8847_
	);
	LUT2 #(
		.INIT('h1)
	) name8386 (
		_w8846_,
		_w8847_,
		_w8848_
	);
	LUT2 #(
		.INIT('h1)
	) name8387 (
		_w3677_,
		_w8848_,
		_w8849_
	);
	LUT2 #(
		.INIT('h8)
	) name8388 (
		_w4532_,
		_w7125_,
		_w8850_
	);
	LUT2 #(
		.INIT('h1)
	) name8389 (
		_w8846_,
		_w8850_,
		_w8851_
	);
	LUT2 #(
		.INIT('h1)
	) name8390 (
		_w3563_,
		_w8851_,
		_w8852_
	);
	LUT2 #(
		.INIT('h8)
	) name8391 (
		_w4532_,
		_w7134_,
		_w8853_
	);
	LUT2 #(
		.INIT('h1)
	) name8392 (
		_w8846_,
		_w8853_,
		_w8854_
	);
	LUT2 #(
		.INIT('h2)
	) name8393 (
		_w1936_,
		_w8854_,
		_w8855_
	);
	LUT2 #(
		.INIT('h8)
	) name8394 (
		_w4532_,
		_w7139_,
		_w8856_
	);
	LUT2 #(
		.INIT('h1)
	) name8395 (
		_w8846_,
		_w8856_,
		_w8857_
	);
	LUT2 #(
		.INIT('h2)
	) name8396 (
		_w3712_,
		_w8857_,
		_w8858_
	);
	LUT2 #(
		.INIT('h2)
	) name8397 (
		\P1_reg1_reg[13]/NET0131 ,
		_w4541_,
		_w8859_
	);
	LUT2 #(
		.INIT('h1)
	) name8398 (
		_w8845_,
		_w8859_,
		_w8860_
	);
	LUT2 #(
		.INIT('h4)
	) name8399 (
		_w8858_,
		_w8860_,
		_w8861_
	);
	LUT2 #(
		.INIT('h4)
	) name8400 (
		_w8849_,
		_w8861_,
		_w8862_
	);
	LUT2 #(
		.INIT('h1)
	) name8401 (
		_w8852_,
		_w8855_,
		_w8863_
	);
	LUT2 #(
		.INIT('h8)
	) name8402 (
		_w8862_,
		_w8863_,
		_w8864_
	);
	LUT2 #(
		.INIT('h2)
	) name8403 (
		_w3450_,
		_w8864_,
		_w8865_
	);
	LUT2 #(
		.INIT('h1)
	) name8404 (
		_w8844_,
		_w8865_,
		_w8866_
	);
	LUT2 #(
		.INIT('h2)
	) name8405 (
		\P1_state_reg[0]/NET0131 ,
		_w8866_,
		_w8867_
	);
	LUT2 #(
		.INIT('h1)
	) name8406 (
		_w8843_,
		_w8867_,
		_w8868_
	);
	LUT2 #(
		.INIT('h2)
	) name8407 (
		\P2_reg0_reg[10]/NET0131 ,
		_w1983_,
		_w8869_
	);
	LUT2 #(
		.INIT('h8)
	) name8408 (
		\P2_reg0_reg[10]/NET0131 ,
		_w2024_,
		_w8870_
	);
	LUT2 #(
		.INIT('h2)
	) name8409 (
		\P2_reg0_reg[10]/NET0131 ,
		_w3423_,
		_w8871_
	);
	LUT2 #(
		.INIT('h2)
	) name8410 (
		\P2_reg0_reg[10]/NET0131 ,
		_w2040_,
		_w8872_
	);
	LUT2 #(
		.INIT('h8)
	) name8411 (
		_w2040_,
		_w7163_,
		_w8873_
	);
	LUT2 #(
		.INIT('h1)
	) name8412 (
		_w8872_,
		_w8873_,
		_w8874_
	);
	LUT2 #(
		.INIT('h2)
	) name8413 (
		_w3411_,
		_w8874_,
		_w8875_
	);
	LUT2 #(
		.INIT('h2)
	) name8414 (
		_w2040_,
		_w7169_,
		_w8876_
	);
	LUT2 #(
		.INIT('h1)
	) name8415 (
		_w8872_,
		_w8876_,
		_w8877_
	);
	LUT2 #(
		.INIT('h1)
	) name8416 (
		_w3177_,
		_w8877_,
		_w8878_
	);
	LUT2 #(
		.INIT('h8)
	) name8417 (
		_w2040_,
		_w7175_,
		_w8879_
	);
	LUT2 #(
		.INIT('h1)
	) name8418 (
		_w8872_,
		_w8879_,
		_w8880_
	);
	LUT2 #(
		.INIT('h1)
	) name8419 (
		_w3320_,
		_w8880_,
		_w8881_
	);
	LUT2 #(
		.INIT('h8)
	) name8420 (
		_w2040_,
		_w7181_,
		_w8882_
	);
	LUT2 #(
		.INIT('h1)
	) name8421 (
		_w8872_,
		_w8882_,
		_w8883_
	);
	LUT2 #(
		.INIT('h2)
	) name8422 (
		_w3355_,
		_w8883_,
		_w8884_
	);
	LUT2 #(
		.INIT('h8)
	) name8423 (
		_w2040_,
		_w8503_,
		_w8885_
	);
	LUT2 #(
		.INIT('h1)
	) name8424 (
		_w8871_,
		_w8885_,
		_w8886_
	);
	LUT2 #(
		.INIT('h4)
	) name8425 (
		_w8884_,
		_w8886_,
		_w8887_
	);
	LUT2 #(
		.INIT('h4)
	) name8426 (
		_w8878_,
		_w8887_,
		_w8888_
	);
	LUT2 #(
		.INIT('h4)
	) name8427 (
		_w8881_,
		_w8888_,
		_w8889_
	);
	LUT2 #(
		.INIT('h4)
	) name8428 (
		_w8875_,
		_w8889_,
		_w8890_
	);
	LUT2 #(
		.INIT('h2)
	) name8429 (
		_w2026_,
		_w8890_,
		_w8891_
	);
	LUT2 #(
		.INIT('h1)
	) name8430 (
		_w8870_,
		_w8891_,
		_w8892_
	);
	LUT2 #(
		.INIT('h2)
	) name8431 (
		\P1_state_reg[0]/NET0131 ,
		_w8892_,
		_w8893_
	);
	LUT2 #(
		.INIT('h1)
	) name8432 (
		_w8869_,
		_w8893_,
		_w8894_
	);
	LUT2 #(
		.INIT('h2)
	) name8433 (
		\P2_reg0_reg[13]/NET0131 ,
		_w1983_,
		_w8895_
	);
	LUT2 #(
		.INIT('h8)
	) name8434 (
		\P2_reg0_reg[13]/NET0131 ,
		_w2024_,
		_w8896_
	);
	LUT2 #(
		.INIT('h2)
	) name8435 (
		_w2040_,
		_w8540_,
		_w8897_
	);
	LUT2 #(
		.INIT('h2)
	) name8436 (
		\P2_reg0_reg[13]/NET0131 ,
		_w2040_,
		_w8898_
	);
	LUT2 #(
		.INIT('h2)
	) name8437 (
		_w2040_,
		_w7205_,
		_w8899_
	);
	LUT2 #(
		.INIT('h1)
	) name8438 (
		_w8898_,
		_w8899_,
		_w8900_
	);
	LUT2 #(
		.INIT('h2)
	) name8439 (
		_w3411_,
		_w8900_,
		_w8901_
	);
	LUT2 #(
		.INIT('h2)
	) name8440 (
		\P2_reg0_reg[13]/NET0131 ,
		_w8385_,
		_w8902_
	);
	LUT2 #(
		.INIT('h8)
	) name8441 (
		_w2040_,
		_w7211_,
		_w8903_
	);
	LUT2 #(
		.INIT('h1)
	) name8442 (
		_w8898_,
		_w8903_,
		_w8904_
	);
	LUT2 #(
		.INIT('h1)
	) name8443 (
		_w3177_,
		_w8904_,
		_w8905_
	);
	LUT2 #(
		.INIT('h1)
	) name8444 (
		_w8897_,
		_w8902_,
		_w8906_
	);
	LUT2 #(
		.INIT('h4)
	) name8445 (
		_w8905_,
		_w8906_,
		_w8907_
	);
	LUT2 #(
		.INIT('h4)
	) name8446 (
		_w8901_,
		_w8907_,
		_w8908_
	);
	LUT2 #(
		.INIT('h2)
	) name8447 (
		_w2026_,
		_w8908_,
		_w8909_
	);
	LUT2 #(
		.INIT('h1)
	) name8448 (
		_w8896_,
		_w8909_,
		_w8910_
	);
	LUT2 #(
		.INIT('h2)
	) name8449 (
		\P1_state_reg[0]/NET0131 ,
		_w8910_,
		_w8911_
	);
	LUT2 #(
		.INIT('h1)
	) name8450 (
		_w8895_,
		_w8911_,
		_w8912_
	);
	LUT2 #(
		.INIT('h2)
	) name8451 (
		\P1_reg1_reg[23]/NET0131 ,
		_w3435_,
		_w8913_
	);
	LUT2 #(
		.INIT('h8)
	) name8452 (
		\P1_reg1_reg[23]/NET0131 ,
		_w3448_,
		_w8914_
	);
	LUT2 #(
		.INIT('h2)
	) name8453 (
		\P1_reg1_reg[23]/NET0131 ,
		_w4532_,
		_w8915_
	);
	LUT2 #(
		.INIT('h2)
	) name8454 (
		_w4532_,
		_w7422_,
		_w8916_
	);
	LUT2 #(
		.INIT('h1)
	) name8455 (
		_w8915_,
		_w8916_,
		_w8917_
	);
	LUT2 #(
		.INIT('h1)
	) name8456 (
		_w3677_,
		_w8917_,
		_w8918_
	);
	LUT2 #(
		.INIT('h2)
	) name8457 (
		_w4532_,
		_w7435_,
		_w8919_
	);
	LUT2 #(
		.INIT('h1)
	) name8458 (
		_w8915_,
		_w8919_,
		_w8920_
	);
	LUT2 #(
		.INIT('h1)
	) name8459 (
		_w3563_,
		_w8920_,
		_w8921_
	);
	LUT2 #(
		.INIT('h2)
	) name8460 (
		_w4532_,
		_w8777_,
		_w8922_
	);
	LUT2 #(
		.INIT('h8)
	) name8461 (
		_w4532_,
		_w7444_,
		_w8923_
	);
	LUT2 #(
		.INIT('h1)
	) name8462 (
		_w8915_,
		_w8923_,
		_w8924_
	);
	LUT2 #(
		.INIT('h2)
	) name8463 (
		_w1936_,
		_w8924_,
		_w8925_
	);
	LUT2 #(
		.INIT('h2)
	) name8464 (
		\P1_reg1_reg[23]/NET0131 ,
		_w4573_,
		_w8926_
	);
	LUT2 #(
		.INIT('h1)
	) name8465 (
		_w8922_,
		_w8926_,
		_w8927_
	);
	LUT2 #(
		.INIT('h4)
	) name8466 (
		_w8925_,
		_w8927_,
		_w8928_
	);
	LUT2 #(
		.INIT('h4)
	) name8467 (
		_w8918_,
		_w8928_,
		_w8929_
	);
	LUT2 #(
		.INIT('h4)
	) name8468 (
		_w8921_,
		_w8929_,
		_w8930_
	);
	LUT2 #(
		.INIT('h2)
	) name8469 (
		_w3450_,
		_w8930_,
		_w8931_
	);
	LUT2 #(
		.INIT('h1)
	) name8470 (
		_w8914_,
		_w8931_,
		_w8932_
	);
	LUT2 #(
		.INIT('h2)
	) name8471 (
		\P1_state_reg[0]/NET0131 ,
		_w8932_,
		_w8933_
	);
	LUT2 #(
		.INIT('h1)
	) name8472 (
		_w8913_,
		_w8933_,
		_w8934_
	);
	LUT2 #(
		.INIT('h4)
	) name8473 (
		\P1_state_reg[0]/NET0131 ,
		\P2_reg3_reg[4]/NET0131 ,
		_w8935_
	);
	LUT2 #(
		.INIT('h8)
	) name8474 (
		_w2635_,
		_w3976_,
		_w8936_
	);
	LUT2 #(
		.INIT('h8)
	) name8475 (
		_w2024_,
		_w2635_,
		_w8937_
	);
	LUT2 #(
		.INIT('h1)
	) name8476 (
		_w2656_,
		_w3965_,
		_w8938_
	);
	LUT2 #(
		.INIT('h2)
	) name8477 (
		_w2635_,
		_w3788_,
		_w8939_
	);
	LUT2 #(
		.INIT('h2)
	) name8478 (
		_w2058_,
		_w2616_,
		_w8940_
	);
	LUT2 #(
		.INIT('h4)
	) name8479 (
		_w2642_,
		_w3376_,
		_w8941_
	);
	LUT2 #(
		.INIT('h2)
	) name8480 (
		_w2531_,
		_w8941_,
		_w8942_
	);
	LUT2 #(
		.INIT('h1)
	) name8481 (
		_w2058_,
		_w3378_,
		_w8943_
	);
	LUT2 #(
		.INIT('h4)
	) name8482 (
		_w8942_,
		_w8943_,
		_w8944_
	);
	LUT2 #(
		.INIT('h1)
	) name8483 (
		_w8940_,
		_w8944_,
		_w8945_
	);
	LUT2 #(
		.INIT('h2)
	) name8484 (
		_w3788_,
		_w8945_,
		_w8946_
	);
	LUT2 #(
		.INIT('h1)
	) name8485 (
		_w8939_,
		_w8946_,
		_w8947_
	);
	LUT2 #(
		.INIT('h2)
	) name8486 (
		_w3411_,
		_w8947_,
		_w8948_
	);
	LUT2 #(
		.INIT('h2)
	) name8487 (
		_w3880_,
		_w4206_,
		_w8949_
	);
	LUT2 #(
		.INIT('h4)
	) name8488 (
		_w3880_,
		_w4206_,
		_w8950_
	);
	LUT2 #(
		.INIT('h1)
	) name8489 (
		_w8949_,
		_w8950_,
		_w8951_
	);
	LUT2 #(
		.INIT('h8)
	) name8490 (
		_w3788_,
		_w8951_,
		_w8952_
	);
	LUT2 #(
		.INIT('h1)
	) name8491 (
		_w8939_,
		_w8952_,
		_w8953_
	);
	LUT2 #(
		.INIT('h1)
	) name8492 (
		_w3177_,
		_w8953_,
		_w8954_
	);
	LUT2 #(
		.INIT('h2)
	) name8493 (
		_w3823_,
		_w4206_,
		_w8955_
	);
	LUT2 #(
		.INIT('h4)
	) name8494 (
		_w3823_,
		_w4206_,
		_w8956_
	);
	LUT2 #(
		.INIT('h1)
	) name8495 (
		_w8955_,
		_w8956_,
		_w8957_
	);
	LUT2 #(
		.INIT('h2)
	) name8496 (
		_w3788_,
		_w8957_,
		_w8958_
	);
	LUT2 #(
		.INIT('h1)
	) name8497 (
		_w8939_,
		_w8958_,
		_w8959_
	);
	LUT2 #(
		.INIT('h1)
	) name8498 (
		_w3320_,
		_w8959_,
		_w8960_
	);
	LUT2 #(
		.INIT('h1)
	) name8499 (
		_w2656_,
		_w3328_,
		_w8961_
	);
	LUT2 #(
		.INIT('h1)
	) name8500 (
		_w3329_,
		_w8961_,
		_w8962_
	);
	LUT2 #(
		.INIT('h8)
	) name8501 (
		_w3788_,
		_w8962_,
		_w8963_
	);
	LUT2 #(
		.INIT('h1)
	) name8502 (
		_w8939_,
		_w8963_,
		_w8964_
	);
	LUT2 #(
		.INIT('h2)
	) name8503 (
		_w3355_,
		_w8964_,
		_w8965_
	);
	LUT2 #(
		.INIT('h2)
	) name8504 (
		_w2635_,
		_w3962_,
		_w8966_
	);
	LUT2 #(
		.INIT('h1)
	) name8505 (
		_w8938_,
		_w8966_,
		_w8967_
	);
	LUT2 #(
		.INIT('h4)
	) name8506 (
		_w8965_,
		_w8967_,
		_w8968_
	);
	LUT2 #(
		.INIT('h4)
	) name8507 (
		_w8954_,
		_w8968_,
		_w8969_
	);
	LUT2 #(
		.INIT('h4)
	) name8508 (
		_w8960_,
		_w8969_,
		_w8970_
	);
	LUT2 #(
		.INIT('h4)
	) name8509 (
		_w8948_,
		_w8970_,
		_w8971_
	);
	LUT2 #(
		.INIT('h2)
	) name8510 (
		_w2026_,
		_w8971_,
		_w8972_
	);
	LUT2 #(
		.INIT('h1)
	) name8511 (
		_w8937_,
		_w8972_,
		_w8973_
	);
	LUT2 #(
		.INIT('h2)
	) name8512 (
		\P1_state_reg[0]/NET0131 ,
		_w8973_,
		_w8974_
	);
	LUT2 #(
		.INIT('h1)
	) name8513 (
		_w8935_,
		_w8936_,
		_w8975_
	);
	LUT2 #(
		.INIT('h4)
	) name8514 (
		_w8974_,
		_w8975_,
		_w8976_
	);
	LUT2 #(
		.INIT('h4)
	) name8515 (
		\P1_state_reg[0]/NET0131 ,
		\P2_reg3_reg[5]/NET0131 ,
		_w8977_
	);
	LUT2 #(
		.INIT('h8)
	) name8516 (
		_w2024_,
		_w2526_,
		_w8978_
	);
	LUT2 #(
		.INIT('h1)
	) name8517 (
		_w2544_,
		_w3965_,
		_w8979_
	);
	LUT2 #(
		.INIT('h2)
	) name8518 (
		_w2526_,
		_w3788_,
		_w8980_
	);
	LUT2 #(
		.INIT('h2)
	) name8519 (
		_w2506_,
		_w3378_,
		_w8981_
	);
	LUT2 #(
		.INIT('h1)
	) name8520 (
		_w3379_,
		_w8981_,
		_w8982_
	);
	LUT2 #(
		.INIT('h1)
	) name8521 (
		_w2058_,
		_w8982_,
		_w8983_
	);
	LUT2 #(
		.INIT('h8)
	) name8522 (
		_w2058_,
		_w2642_,
		_w8984_
	);
	LUT2 #(
		.INIT('h1)
	) name8523 (
		_w8983_,
		_w8984_,
		_w8985_
	);
	LUT2 #(
		.INIT('h8)
	) name8524 (
		_w3788_,
		_w8985_,
		_w8986_
	);
	LUT2 #(
		.INIT('h1)
	) name8525 (
		_w8980_,
		_w8986_,
		_w8987_
	);
	LUT2 #(
		.INIT('h2)
	) name8526 (
		_w3411_,
		_w8987_,
		_w8988_
	);
	LUT2 #(
		.INIT('h4)
	) name8527 (
		_w2664_,
		_w4194_,
		_w8989_
	);
	LUT2 #(
		.INIT('h2)
	) name8528 (
		_w2664_,
		_w4194_,
		_w8990_
	);
	LUT2 #(
		.INIT('h1)
	) name8529 (
		_w8989_,
		_w8990_,
		_w8991_
	);
	LUT2 #(
		.INIT('h2)
	) name8530 (
		_w3788_,
		_w8991_,
		_w8992_
	);
	LUT2 #(
		.INIT('h1)
	) name8531 (
		_w8980_,
		_w8992_,
		_w8993_
	);
	LUT2 #(
		.INIT('h1)
	) name8532 (
		_w3177_,
		_w8993_,
		_w8994_
	);
	LUT2 #(
		.INIT('h1)
	) name8533 (
		_w2544_,
		_w3329_,
		_w8995_
	);
	LUT2 #(
		.INIT('h4)
	) name8534 (
		_w3330_,
		_w3355_,
		_w8996_
	);
	LUT2 #(
		.INIT('h4)
	) name8535 (
		_w8995_,
		_w8996_,
		_w8997_
	);
	LUT2 #(
		.INIT('h2)
	) name8536 (
		_w3271_,
		_w4194_,
		_w8998_
	);
	LUT2 #(
		.INIT('h4)
	) name8537 (
		_w3271_,
		_w4194_,
		_w8999_
	);
	LUT2 #(
		.INIT('h1)
	) name8538 (
		_w3320_,
		_w8998_,
		_w9000_
	);
	LUT2 #(
		.INIT('h4)
	) name8539 (
		_w8999_,
		_w9000_,
		_w9001_
	);
	LUT2 #(
		.INIT('h1)
	) name8540 (
		_w8997_,
		_w9001_,
		_w9002_
	);
	LUT2 #(
		.INIT('h2)
	) name8541 (
		_w3788_,
		_w9002_,
		_w9003_
	);
	LUT2 #(
		.INIT('h2)
	) name8542 (
		_w5698_,
		_w6311_,
		_w9004_
	);
	LUT2 #(
		.INIT('h2)
	) name8543 (
		_w2526_,
		_w9004_,
		_w9005_
	);
	LUT2 #(
		.INIT('h1)
	) name8544 (
		_w8979_,
		_w9005_,
		_w9006_
	);
	LUT2 #(
		.INIT('h4)
	) name8545 (
		_w9003_,
		_w9006_,
		_w9007_
	);
	LUT2 #(
		.INIT('h4)
	) name8546 (
		_w8994_,
		_w9007_,
		_w9008_
	);
	LUT2 #(
		.INIT('h4)
	) name8547 (
		_w8988_,
		_w9008_,
		_w9009_
	);
	LUT2 #(
		.INIT('h2)
	) name8548 (
		_w2026_,
		_w9009_,
		_w9010_
	);
	LUT2 #(
		.INIT('h1)
	) name8549 (
		_w8978_,
		_w9010_,
		_w9011_
	);
	LUT2 #(
		.INIT('h2)
	) name8550 (
		\P1_state_reg[0]/NET0131 ,
		_w9011_,
		_w9012_
	);
	LUT2 #(
		.INIT('h8)
	) name8551 (
		_w2526_,
		_w3976_,
		_w9013_
	);
	LUT2 #(
		.INIT('h1)
	) name8552 (
		_w8977_,
		_w9013_,
		_w9014_
	);
	LUT2 #(
		.INIT('h4)
	) name8553 (
		_w9012_,
		_w9014_,
		_w9015_
	);
	LUT2 #(
		.INIT('h2)
	) name8554 (
		\P1_reg3_reg[4]/NET0131 ,
		\P1_state_reg[0]/NET0131 ,
		_w9016_
	);
	LUT2 #(
		.INIT('h8)
	) name8555 (
		_w1568_,
		_w1953_,
		_w9017_
	);
	LUT2 #(
		.INIT('h8)
	) name8556 (
		_w1568_,
		_w3448_,
		_w9018_
	);
	LUT2 #(
		.INIT('h1)
	) name8557 (
		_w1586_,
		_w4067_,
		_w9019_
	);
	LUT2 #(
		.INIT('h2)
	) name8558 (
		_w1568_,
		_w3980_,
		_w9020_
	);
	LUT2 #(
		.INIT('h2)
	) name8559 (
		_w537_,
		_w1617_,
		_w9021_
	);
	LUT2 #(
		.INIT('h4)
	) name8560 (
		_w1572_,
		_w3573_,
		_w9022_
	);
	LUT2 #(
		.INIT('h2)
	) name8561 (
		_w1548_,
		_w9022_,
		_w9023_
	);
	LUT2 #(
		.INIT('h1)
	) name8562 (
		_w537_,
		_w3575_,
		_w9024_
	);
	LUT2 #(
		.INIT('h4)
	) name8563 (
		_w9023_,
		_w9024_,
		_w9025_
	);
	LUT2 #(
		.INIT('h1)
	) name8564 (
		_w9021_,
		_w9025_,
		_w9026_
	);
	LUT2 #(
		.INIT('h2)
	) name8565 (
		_w3980_,
		_w9026_,
		_w9027_
	);
	LUT2 #(
		.INIT('h1)
	) name8566 (
		_w9020_,
		_w9027_,
		_w9028_
	);
	LUT2 #(
		.INIT('h2)
	) name8567 (
		_w1936_,
		_w9028_,
		_w9029_
	);
	LUT2 #(
		.INIT('h2)
	) name8568 (
		_w1806_,
		_w3986_,
		_w9030_
	);
	LUT2 #(
		.INIT('h4)
	) name8569 (
		_w1806_,
		_w3986_,
		_w9031_
	);
	LUT2 #(
		.INIT('h1)
	) name8570 (
		_w9030_,
		_w9031_,
		_w9032_
	);
	LUT2 #(
		.INIT('h2)
	) name8571 (
		_w3980_,
		_w9032_,
		_w9033_
	);
	LUT2 #(
		.INIT('h1)
	) name8572 (
		_w9020_,
		_w9033_,
		_w9034_
	);
	LUT2 #(
		.INIT('h1)
	) name8573 (
		_w3563_,
		_w9034_,
		_w9035_
	);
	LUT2 #(
		.INIT('h4)
	) name8574 (
		_w1680_,
		_w1806_,
		_w9036_
	);
	LUT2 #(
		.INIT('h2)
	) name8575 (
		_w1680_,
		_w1806_,
		_w9037_
	);
	LUT2 #(
		.INIT('h1)
	) name8576 (
		_w9036_,
		_w9037_,
		_w9038_
	);
	LUT2 #(
		.INIT('h8)
	) name8577 (
		_w3980_,
		_w9038_,
		_w9039_
	);
	LUT2 #(
		.INIT('h1)
	) name8578 (
		_w9020_,
		_w9039_,
		_w9040_
	);
	LUT2 #(
		.INIT('h1)
	) name8579 (
		_w3677_,
		_w9040_,
		_w9041_
	);
	LUT2 #(
		.INIT('h1)
	) name8580 (
		_w1586_,
		_w3681_,
		_w9042_
	);
	LUT2 #(
		.INIT('h1)
	) name8581 (
		_w3682_,
		_w9042_,
		_w9043_
	);
	LUT2 #(
		.INIT('h8)
	) name8582 (
		_w3980_,
		_w9043_,
		_w9044_
	);
	LUT2 #(
		.INIT('h1)
	) name8583 (
		_w9020_,
		_w9044_,
		_w9045_
	);
	LUT2 #(
		.INIT('h2)
	) name8584 (
		_w3712_,
		_w9045_,
		_w9046_
	);
	LUT2 #(
		.INIT('h2)
	) name8585 (
		_w1568_,
		_w4064_,
		_w9047_
	);
	LUT2 #(
		.INIT('h1)
	) name8586 (
		_w9019_,
		_w9047_,
		_w9048_
	);
	LUT2 #(
		.INIT('h4)
	) name8587 (
		_w9046_,
		_w9048_,
		_w9049_
	);
	LUT2 #(
		.INIT('h4)
	) name8588 (
		_w9035_,
		_w9049_,
		_w9050_
	);
	LUT2 #(
		.INIT('h4)
	) name8589 (
		_w9041_,
		_w9050_,
		_w9051_
	);
	LUT2 #(
		.INIT('h4)
	) name8590 (
		_w9029_,
		_w9051_,
		_w9052_
	);
	LUT2 #(
		.INIT('h2)
	) name8591 (
		_w3450_,
		_w9052_,
		_w9053_
	);
	LUT2 #(
		.INIT('h1)
	) name8592 (
		_w9018_,
		_w9053_,
		_w9054_
	);
	LUT2 #(
		.INIT('h2)
	) name8593 (
		\P1_state_reg[0]/NET0131 ,
		_w9054_,
		_w9055_
	);
	LUT2 #(
		.INIT('h1)
	) name8594 (
		_w9016_,
		_w9017_,
		_w9056_
	);
	LUT2 #(
		.INIT('h4)
	) name8595 (
		_w9055_,
		_w9056_,
		_w9057_
	);
	LUT2 #(
		.INIT('h2)
	) name8596 (
		\P1_reg3_reg[5]/NET0131 ,
		\P1_state_reg[0]/NET0131 ,
		_w9058_
	);
	LUT2 #(
		.INIT('h8)
	) name8597 (
		_w1543_,
		_w1953_,
		_w9059_
	);
	LUT2 #(
		.INIT('h8)
	) name8598 (
		_w1543_,
		_w3448_,
		_w9060_
	);
	LUT2 #(
		.INIT('h4)
	) name8599 (
		_w1562_,
		_w1880_,
		_w9061_
	);
	LUT2 #(
		.INIT('h1)
	) name8600 (
		_w1562_,
		_w3682_,
		_w9062_
	);
	LUT2 #(
		.INIT('h1)
	) name8601 (
		_w3683_,
		_w9062_,
		_w9063_
	);
	LUT2 #(
		.INIT('h8)
	) name8602 (
		_w3712_,
		_w9063_,
		_w9064_
	);
	LUT2 #(
		.INIT('h1)
	) name8603 (
		_w9061_,
		_w9064_,
		_w9065_
	);
	LUT2 #(
		.INIT('h2)
	) name8604 (
		_w3980_,
		_w9065_,
		_w9066_
	);
	LUT2 #(
		.INIT('h2)
	) name8605 (
		_w1543_,
		_w3980_,
		_w9067_
	);
	LUT2 #(
		.INIT('h2)
	) name8606 (
		_w1524_,
		_w3575_,
		_w9068_
	);
	LUT2 #(
		.INIT('h4)
	) name8607 (
		_w1524_,
		_w3575_,
		_w9069_
	);
	LUT2 #(
		.INIT('h1)
	) name8608 (
		_w9068_,
		_w9069_,
		_w9070_
	);
	LUT2 #(
		.INIT('h1)
	) name8609 (
		_w537_,
		_w9070_,
		_w9071_
	);
	LUT2 #(
		.INIT('h8)
	) name8610 (
		_w537_,
		_w1572_,
		_w9072_
	);
	LUT2 #(
		.INIT('h1)
	) name8611 (
		_w9071_,
		_w9072_,
		_w9073_
	);
	LUT2 #(
		.INIT('h8)
	) name8612 (
		_w3980_,
		_w9073_,
		_w9074_
	);
	LUT2 #(
		.INIT('h1)
	) name8613 (
		_w9067_,
		_w9074_,
		_w9075_
	);
	LUT2 #(
		.INIT('h2)
	) name8614 (
		_w1936_,
		_w9075_,
		_w9076_
	);
	LUT2 #(
		.INIT('h2)
	) name8615 (
		_w1805_,
		_w3518_,
		_w9077_
	);
	LUT2 #(
		.INIT('h4)
	) name8616 (
		_w1805_,
		_w3518_,
		_w9078_
	);
	LUT2 #(
		.INIT('h1)
	) name8617 (
		_w9077_,
		_w9078_,
		_w9079_
	);
	LUT2 #(
		.INIT('h2)
	) name8618 (
		_w3980_,
		_w9079_,
		_w9080_
	);
	LUT2 #(
		.INIT('h1)
	) name8619 (
		_w9067_,
		_w9080_,
		_w9081_
	);
	LUT2 #(
		.INIT('h1)
	) name8620 (
		_w3563_,
		_w9081_,
		_w9082_
	);
	LUT2 #(
		.INIT('h2)
	) name8621 (
		_w1805_,
		_w3636_,
		_w9083_
	);
	LUT2 #(
		.INIT('h4)
	) name8622 (
		_w1805_,
		_w3636_,
		_w9084_
	);
	LUT2 #(
		.INIT('h1)
	) name8623 (
		_w9083_,
		_w9084_,
		_w9085_
	);
	LUT2 #(
		.INIT('h2)
	) name8624 (
		_w3980_,
		_w9085_,
		_w9086_
	);
	LUT2 #(
		.INIT('h1)
	) name8625 (
		_w9067_,
		_w9086_,
		_w9087_
	);
	LUT2 #(
		.INIT('h1)
	) name8626 (
		_w3677_,
		_w9087_,
		_w9088_
	);
	LUT2 #(
		.INIT('h4)
	) name8627 (
		_w1562_,
		_w1763_,
		_w9089_
	);
	LUT2 #(
		.INIT('h4)
	) name8628 (
		_w1761_,
		_w1762_,
		_w9090_
	);
	LUT2 #(
		.INIT('h4)
	) name8629 (
		_w3980_,
		_w9090_,
		_w9091_
	);
	LUT2 #(
		.INIT('h1)
	) name8630 (
		_w3716_,
		_w9091_,
		_w9092_
	);
	LUT2 #(
		.INIT('h2)
	) name8631 (
		_w1543_,
		_w9092_,
		_w9093_
	);
	LUT2 #(
		.INIT('h1)
	) name8632 (
		_w9089_,
		_w9093_,
		_w9094_
	);
	LUT2 #(
		.INIT('h4)
	) name8633 (
		_w9066_,
		_w9094_,
		_w9095_
	);
	LUT2 #(
		.INIT('h4)
	) name8634 (
		_w9082_,
		_w9095_,
		_w9096_
	);
	LUT2 #(
		.INIT('h4)
	) name8635 (
		_w9088_,
		_w9096_,
		_w9097_
	);
	LUT2 #(
		.INIT('h4)
	) name8636 (
		_w9076_,
		_w9097_,
		_w9098_
	);
	LUT2 #(
		.INIT('h2)
	) name8637 (
		_w3450_,
		_w9098_,
		_w9099_
	);
	LUT2 #(
		.INIT('h1)
	) name8638 (
		_w9060_,
		_w9099_,
		_w9100_
	);
	LUT2 #(
		.INIT('h2)
	) name8639 (
		\P1_state_reg[0]/NET0131 ,
		_w9100_,
		_w9101_
	);
	LUT2 #(
		.INIT('h1)
	) name8640 (
		_w9058_,
		_w9059_,
		_w9102_
	);
	LUT2 #(
		.INIT('h4)
	) name8641 (
		_w9101_,
		_w9102_,
		_w9103_
	);
	LUT2 #(
		.INIT('h2)
	) name8642 (
		\P1_reg1_reg[4]/NET0131 ,
		_w3435_,
		_w9104_
	);
	LUT2 #(
		.INIT('h8)
	) name8643 (
		\P1_reg1_reg[4]/NET0131 ,
		_w3448_,
		_w9105_
	);
	LUT2 #(
		.INIT('h4)
	) name8644 (
		_w1586_,
		_w1880_,
		_w9106_
	);
	LUT2 #(
		.INIT('h8)
	) name8645 (
		_w4532_,
		_w9106_,
		_w9107_
	);
	LUT2 #(
		.INIT('h2)
	) name8646 (
		\P1_reg1_reg[4]/NET0131 ,
		_w4532_,
		_w9108_
	);
	LUT2 #(
		.INIT('h2)
	) name8647 (
		_w4532_,
		_w9026_,
		_w9109_
	);
	LUT2 #(
		.INIT('h1)
	) name8648 (
		_w9108_,
		_w9109_,
		_w9110_
	);
	LUT2 #(
		.INIT('h2)
	) name8649 (
		_w1936_,
		_w9110_,
		_w9111_
	);
	LUT2 #(
		.INIT('h2)
	) name8650 (
		_w4532_,
		_w9032_,
		_w9112_
	);
	LUT2 #(
		.INIT('h1)
	) name8651 (
		_w9108_,
		_w9112_,
		_w9113_
	);
	LUT2 #(
		.INIT('h1)
	) name8652 (
		_w3563_,
		_w9113_,
		_w9114_
	);
	LUT2 #(
		.INIT('h8)
	) name8653 (
		_w4532_,
		_w9038_,
		_w9115_
	);
	LUT2 #(
		.INIT('h1)
	) name8654 (
		_w9108_,
		_w9115_,
		_w9116_
	);
	LUT2 #(
		.INIT('h1)
	) name8655 (
		_w3677_,
		_w9116_,
		_w9117_
	);
	LUT2 #(
		.INIT('h8)
	) name8656 (
		_w4532_,
		_w9043_,
		_w9118_
	);
	LUT2 #(
		.INIT('h1)
	) name8657 (
		_w9108_,
		_w9118_,
		_w9119_
	);
	LUT2 #(
		.INIT('h2)
	) name8658 (
		_w3712_,
		_w9119_,
		_w9120_
	);
	LUT2 #(
		.INIT('h2)
	) name8659 (
		\P1_reg1_reg[4]/NET0131 ,
		_w4541_,
		_w9121_
	);
	LUT2 #(
		.INIT('h1)
	) name8660 (
		_w9107_,
		_w9121_,
		_w9122_
	);
	LUT2 #(
		.INIT('h4)
	) name8661 (
		_w9120_,
		_w9122_,
		_w9123_
	);
	LUT2 #(
		.INIT('h4)
	) name8662 (
		_w9114_,
		_w9123_,
		_w9124_
	);
	LUT2 #(
		.INIT('h4)
	) name8663 (
		_w9117_,
		_w9124_,
		_w9125_
	);
	LUT2 #(
		.INIT('h4)
	) name8664 (
		_w9111_,
		_w9125_,
		_w9126_
	);
	LUT2 #(
		.INIT('h2)
	) name8665 (
		_w3450_,
		_w9126_,
		_w9127_
	);
	LUT2 #(
		.INIT('h1)
	) name8666 (
		_w9105_,
		_w9127_,
		_w9128_
	);
	LUT2 #(
		.INIT('h2)
	) name8667 (
		\P1_state_reg[0]/NET0131 ,
		_w9128_,
		_w9129_
	);
	LUT2 #(
		.INIT('h1)
	) name8668 (
		_w9104_,
		_w9129_,
		_w9130_
	);
	LUT2 #(
		.INIT('h2)
	) name8669 (
		\P1_reg0_reg[4]/NET0131 ,
		_w3435_,
		_w9131_
	);
	LUT2 #(
		.INIT('h8)
	) name8670 (
		\P1_reg0_reg[4]/NET0131 ,
		_w3448_,
		_w9132_
	);
	LUT2 #(
		.INIT('h8)
	) name8671 (
		_w4396_,
		_w9106_,
		_w9133_
	);
	LUT2 #(
		.INIT('h2)
	) name8672 (
		\P1_reg0_reg[4]/NET0131 ,
		_w4396_,
		_w9134_
	);
	LUT2 #(
		.INIT('h2)
	) name8673 (
		_w4396_,
		_w9026_,
		_w9135_
	);
	LUT2 #(
		.INIT('h1)
	) name8674 (
		_w9134_,
		_w9135_,
		_w9136_
	);
	LUT2 #(
		.INIT('h2)
	) name8675 (
		_w1936_,
		_w9136_,
		_w9137_
	);
	LUT2 #(
		.INIT('h2)
	) name8676 (
		_w4396_,
		_w9032_,
		_w9138_
	);
	LUT2 #(
		.INIT('h1)
	) name8677 (
		_w9134_,
		_w9138_,
		_w9139_
	);
	LUT2 #(
		.INIT('h1)
	) name8678 (
		_w3563_,
		_w9139_,
		_w9140_
	);
	LUT2 #(
		.INIT('h8)
	) name8679 (
		_w4396_,
		_w9038_,
		_w9141_
	);
	LUT2 #(
		.INIT('h1)
	) name8680 (
		_w9134_,
		_w9141_,
		_w9142_
	);
	LUT2 #(
		.INIT('h1)
	) name8681 (
		_w3677_,
		_w9142_,
		_w9143_
	);
	LUT2 #(
		.INIT('h8)
	) name8682 (
		_w4396_,
		_w9043_,
		_w9144_
	);
	LUT2 #(
		.INIT('h1)
	) name8683 (
		_w9134_,
		_w9144_,
		_w9145_
	);
	LUT2 #(
		.INIT('h2)
	) name8684 (
		_w3712_,
		_w9145_,
		_w9146_
	);
	LUT2 #(
		.INIT('h2)
	) name8685 (
		\P1_reg0_reg[4]/NET0131 ,
		_w4493_,
		_w9147_
	);
	LUT2 #(
		.INIT('h1)
	) name8686 (
		_w9133_,
		_w9147_,
		_w9148_
	);
	LUT2 #(
		.INIT('h4)
	) name8687 (
		_w9146_,
		_w9148_,
		_w9149_
	);
	LUT2 #(
		.INIT('h4)
	) name8688 (
		_w9140_,
		_w9149_,
		_w9150_
	);
	LUT2 #(
		.INIT('h4)
	) name8689 (
		_w9143_,
		_w9150_,
		_w9151_
	);
	LUT2 #(
		.INIT('h4)
	) name8690 (
		_w9137_,
		_w9151_,
		_w9152_
	);
	LUT2 #(
		.INIT('h2)
	) name8691 (
		_w3450_,
		_w9152_,
		_w9153_
	);
	LUT2 #(
		.INIT('h1)
	) name8692 (
		_w9132_,
		_w9153_,
		_w9154_
	);
	LUT2 #(
		.INIT('h2)
	) name8693 (
		\P1_state_reg[0]/NET0131 ,
		_w9154_,
		_w9155_
	);
	LUT2 #(
		.INIT('h1)
	) name8694 (
		_w9131_,
		_w9155_,
		_w9156_
	);
	LUT2 #(
		.INIT('h2)
	) name8695 (
		\P2_reg0_reg[4]/NET0131 ,
		_w1983_,
		_w9157_
	);
	LUT2 #(
		.INIT('h8)
	) name8696 (
		\P2_reg0_reg[4]/NET0131 ,
		_w2024_,
		_w9158_
	);
	LUT2 #(
		.INIT('h4)
	) name8697 (
		_w2656_,
		_w3358_,
		_w9159_
	);
	LUT2 #(
		.INIT('h8)
	) name8698 (
		_w2040_,
		_w9159_,
		_w9160_
	);
	LUT2 #(
		.INIT('h2)
	) name8699 (
		\P2_reg0_reg[4]/NET0131 ,
		_w2040_,
		_w9161_
	);
	LUT2 #(
		.INIT('h2)
	) name8700 (
		_w2040_,
		_w8945_,
		_w9162_
	);
	LUT2 #(
		.INIT('h1)
	) name8701 (
		_w9161_,
		_w9162_,
		_w9163_
	);
	LUT2 #(
		.INIT('h2)
	) name8702 (
		_w3411_,
		_w9163_,
		_w9164_
	);
	LUT2 #(
		.INIT('h2)
	) name8703 (
		_w2040_,
		_w8957_,
		_w9165_
	);
	LUT2 #(
		.INIT('h1)
	) name8704 (
		_w9161_,
		_w9165_,
		_w9166_
	);
	LUT2 #(
		.INIT('h1)
	) name8705 (
		_w3320_,
		_w9166_,
		_w9167_
	);
	LUT2 #(
		.INIT('h8)
	) name8706 (
		_w2040_,
		_w8951_,
		_w9168_
	);
	LUT2 #(
		.INIT('h1)
	) name8707 (
		_w9161_,
		_w9168_,
		_w9169_
	);
	LUT2 #(
		.INIT('h1)
	) name8708 (
		_w3177_,
		_w9169_,
		_w9170_
	);
	LUT2 #(
		.INIT('h8)
	) name8709 (
		_w2040_,
		_w8962_,
		_w9171_
	);
	LUT2 #(
		.INIT('h1)
	) name8710 (
		_w9161_,
		_w9171_,
		_w9172_
	);
	LUT2 #(
		.INIT('h2)
	) name8711 (
		_w3355_,
		_w9172_,
		_w9173_
	);
	LUT2 #(
		.INIT('h2)
	) name8712 (
		\P2_reg0_reg[4]/NET0131 ,
		_w3423_,
		_w9174_
	);
	LUT2 #(
		.INIT('h1)
	) name8713 (
		_w9160_,
		_w9174_,
		_w9175_
	);
	LUT2 #(
		.INIT('h4)
	) name8714 (
		_w9173_,
		_w9175_,
		_w9176_
	);
	LUT2 #(
		.INIT('h4)
	) name8715 (
		_w9167_,
		_w9176_,
		_w9177_
	);
	LUT2 #(
		.INIT('h4)
	) name8716 (
		_w9170_,
		_w9177_,
		_w9178_
	);
	LUT2 #(
		.INIT('h4)
	) name8717 (
		_w9164_,
		_w9178_,
		_w9179_
	);
	LUT2 #(
		.INIT('h2)
	) name8718 (
		_w2026_,
		_w9179_,
		_w9180_
	);
	LUT2 #(
		.INIT('h1)
	) name8719 (
		_w9158_,
		_w9180_,
		_w9181_
	);
	LUT2 #(
		.INIT('h2)
	) name8720 (
		\P1_state_reg[0]/NET0131 ,
		_w9181_,
		_w9182_
	);
	LUT2 #(
		.INIT('h1)
	) name8721 (
		_w9157_,
		_w9182_,
		_w9183_
	);
	LUT2 #(
		.INIT('h2)
	) name8722 (
		\P2_reg1_reg[4]/NET0131 ,
		_w1983_,
		_w9184_
	);
	LUT2 #(
		.INIT('h8)
	) name8723 (
		\P2_reg1_reg[4]/NET0131 ,
		_w2024_,
		_w9185_
	);
	LUT2 #(
		.INIT('h8)
	) name8724 (
		_w3733_,
		_w9159_,
		_w9186_
	);
	LUT2 #(
		.INIT('h2)
	) name8725 (
		\P2_reg1_reg[4]/NET0131 ,
		_w3733_,
		_w9187_
	);
	LUT2 #(
		.INIT('h2)
	) name8726 (
		_w3733_,
		_w8945_,
		_w9188_
	);
	LUT2 #(
		.INIT('h1)
	) name8727 (
		_w9187_,
		_w9188_,
		_w9189_
	);
	LUT2 #(
		.INIT('h2)
	) name8728 (
		_w3411_,
		_w9189_,
		_w9190_
	);
	LUT2 #(
		.INIT('h8)
	) name8729 (
		_w3733_,
		_w8951_,
		_w9191_
	);
	LUT2 #(
		.INIT('h1)
	) name8730 (
		_w9187_,
		_w9191_,
		_w9192_
	);
	LUT2 #(
		.INIT('h1)
	) name8731 (
		_w3177_,
		_w9192_,
		_w9193_
	);
	LUT2 #(
		.INIT('h2)
	) name8732 (
		_w3733_,
		_w8957_,
		_w9194_
	);
	LUT2 #(
		.INIT('h1)
	) name8733 (
		_w9187_,
		_w9194_,
		_w9195_
	);
	LUT2 #(
		.INIT('h1)
	) name8734 (
		_w3320_,
		_w9195_,
		_w9196_
	);
	LUT2 #(
		.INIT('h8)
	) name8735 (
		_w3733_,
		_w8962_,
		_w9197_
	);
	LUT2 #(
		.INIT('h1)
	) name8736 (
		_w9187_,
		_w9197_,
		_w9198_
	);
	LUT2 #(
		.INIT('h2)
	) name8737 (
		_w3355_,
		_w9198_,
		_w9199_
	);
	LUT2 #(
		.INIT('h2)
	) name8738 (
		\P2_reg1_reg[4]/NET0131 ,
		_w3743_,
		_w9200_
	);
	LUT2 #(
		.INIT('h1)
	) name8739 (
		_w9186_,
		_w9200_,
		_w9201_
	);
	LUT2 #(
		.INIT('h4)
	) name8740 (
		_w9199_,
		_w9201_,
		_w9202_
	);
	LUT2 #(
		.INIT('h4)
	) name8741 (
		_w9193_,
		_w9202_,
		_w9203_
	);
	LUT2 #(
		.INIT('h4)
	) name8742 (
		_w9196_,
		_w9203_,
		_w9204_
	);
	LUT2 #(
		.INIT('h4)
	) name8743 (
		_w9190_,
		_w9204_,
		_w9205_
	);
	LUT2 #(
		.INIT('h2)
	) name8744 (
		_w2026_,
		_w9205_,
		_w9206_
	);
	LUT2 #(
		.INIT('h1)
	) name8745 (
		_w9185_,
		_w9206_,
		_w9207_
	);
	LUT2 #(
		.INIT('h2)
	) name8746 (
		\P1_state_reg[0]/NET0131 ,
		_w9207_,
		_w9208_
	);
	LUT2 #(
		.INIT('h1)
	) name8747 (
		_w9184_,
		_w9208_,
		_w9209_
	);
	LUT2 #(
		.INIT('h2)
	) name8748 (
		\P1_reg2_reg[8]/NET0131 ,
		_w3435_,
		_w9210_
	);
	LUT2 #(
		.INIT('h8)
	) name8749 (
		\P1_reg2_reg[8]/NET0131 ,
		_w3448_,
		_w9211_
	);
	LUT2 #(
		.INIT('h8)
	) name8750 (
		_w1281_,
		_w1880_,
		_w9212_
	);
	LUT2 #(
		.INIT('h8)
	) name8751 (
		_w3466_,
		_w9212_,
		_w9213_
	);
	LUT2 #(
		.INIT('h2)
	) name8752 (
		\P1_reg2_reg[8]/NET0131 ,
		_w3466_,
		_w9214_
	);
	LUT2 #(
		.INIT('h8)
	) name8753 (
		_w3466_,
		_w8292_,
		_w9215_
	);
	LUT2 #(
		.INIT('h1)
	) name8754 (
		_w9214_,
		_w9215_,
		_w9216_
	);
	LUT2 #(
		.INIT('h2)
	) name8755 (
		_w1936_,
		_w9216_,
		_w9217_
	);
	LUT2 #(
		.INIT('h8)
	) name8756 (
		_w3466_,
		_w8298_,
		_w9218_
	);
	LUT2 #(
		.INIT('h1)
	) name8757 (
		_w9214_,
		_w9218_,
		_w9219_
	);
	LUT2 #(
		.INIT('h1)
	) name8758 (
		_w3563_,
		_w9219_,
		_w9220_
	);
	LUT2 #(
		.INIT('h2)
	) name8759 (
		_w3466_,
		_w8304_,
		_w9221_
	);
	LUT2 #(
		.INIT('h1)
	) name8760 (
		_w9214_,
		_w9221_,
		_w9222_
	);
	LUT2 #(
		.INIT('h1)
	) name8761 (
		_w3677_,
		_w9222_,
		_w9223_
	);
	LUT2 #(
		.INIT('h8)
	) name8762 (
		_w3466_,
		_w8310_,
		_w9224_
	);
	LUT2 #(
		.INIT('h1)
	) name8763 (
		_w9214_,
		_w9224_,
		_w9225_
	);
	LUT2 #(
		.INIT('h2)
	) name8764 (
		_w3712_,
		_w9225_,
		_w9226_
	);
	LUT2 #(
		.INIT('h8)
	) name8765 (
		_w1262_,
		_w1763_,
		_w9227_
	);
	LUT2 #(
		.INIT('h2)
	) name8766 (
		\P1_reg2_reg[8]/NET0131 ,
		_w3718_,
		_w9228_
	);
	LUT2 #(
		.INIT('h1)
	) name8767 (
		_w9213_,
		_w9227_,
		_w9229_
	);
	LUT2 #(
		.INIT('h4)
	) name8768 (
		_w9228_,
		_w9229_,
		_w9230_
	);
	LUT2 #(
		.INIT('h4)
	) name8769 (
		_w9226_,
		_w9230_,
		_w9231_
	);
	LUT2 #(
		.INIT('h4)
	) name8770 (
		_w9220_,
		_w9231_,
		_w9232_
	);
	LUT2 #(
		.INIT('h4)
	) name8771 (
		_w9223_,
		_w9232_,
		_w9233_
	);
	LUT2 #(
		.INIT('h4)
	) name8772 (
		_w9217_,
		_w9233_,
		_w9234_
	);
	LUT2 #(
		.INIT('h2)
	) name8773 (
		_w3450_,
		_w9234_,
		_w9235_
	);
	LUT2 #(
		.INIT('h1)
	) name8774 (
		_w9211_,
		_w9235_,
		_w9236_
	);
	LUT2 #(
		.INIT('h2)
	) name8775 (
		\P1_state_reg[0]/NET0131 ,
		_w9236_,
		_w9237_
	);
	LUT2 #(
		.INIT('h1)
	) name8776 (
		_w9210_,
		_w9237_,
		_w9238_
	);
	LUT2 #(
		.INIT('h2)
	) name8777 (
		\P1_reg1_reg[8]/NET0131 ,
		_w3435_,
		_w9239_
	);
	LUT2 #(
		.INIT('h8)
	) name8778 (
		\P1_reg1_reg[8]/NET0131 ,
		_w3448_,
		_w9240_
	);
	LUT2 #(
		.INIT('h8)
	) name8779 (
		_w4532_,
		_w9212_,
		_w9241_
	);
	LUT2 #(
		.INIT('h2)
	) name8780 (
		\P1_reg1_reg[8]/NET0131 ,
		_w4532_,
		_w9242_
	);
	LUT2 #(
		.INIT('h8)
	) name8781 (
		_w4532_,
		_w8292_,
		_w9243_
	);
	LUT2 #(
		.INIT('h1)
	) name8782 (
		_w9242_,
		_w9243_,
		_w9244_
	);
	LUT2 #(
		.INIT('h2)
	) name8783 (
		_w1936_,
		_w9244_,
		_w9245_
	);
	LUT2 #(
		.INIT('h2)
	) name8784 (
		_w4532_,
		_w8304_,
		_w9246_
	);
	LUT2 #(
		.INIT('h1)
	) name8785 (
		_w9242_,
		_w9246_,
		_w9247_
	);
	LUT2 #(
		.INIT('h1)
	) name8786 (
		_w3677_,
		_w9247_,
		_w9248_
	);
	LUT2 #(
		.INIT('h8)
	) name8787 (
		_w4532_,
		_w8298_,
		_w9249_
	);
	LUT2 #(
		.INIT('h1)
	) name8788 (
		_w9242_,
		_w9249_,
		_w9250_
	);
	LUT2 #(
		.INIT('h1)
	) name8789 (
		_w3563_,
		_w9250_,
		_w9251_
	);
	LUT2 #(
		.INIT('h8)
	) name8790 (
		_w4532_,
		_w8310_,
		_w9252_
	);
	LUT2 #(
		.INIT('h1)
	) name8791 (
		_w9242_,
		_w9252_,
		_w9253_
	);
	LUT2 #(
		.INIT('h2)
	) name8792 (
		_w3712_,
		_w9253_,
		_w9254_
	);
	LUT2 #(
		.INIT('h2)
	) name8793 (
		\P1_reg1_reg[8]/NET0131 ,
		_w4541_,
		_w9255_
	);
	LUT2 #(
		.INIT('h1)
	) name8794 (
		_w9241_,
		_w9255_,
		_w9256_
	);
	LUT2 #(
		.INIT('h4)
	) name8795 (
		_w9254_,
		_w9256_,
		_w9257_
	);
	LUT2 #(
		.INIT('h4)
	) name8796 (
		_w9248_,
		_w9257_,
		_w9258_
	);
	LUT2 #(
		.INIT('h4)
	) name8797 (
		_w9251_,
		_w9258_,
		_w9259_
	);
	LUT2 #(
		.INIT('h4)
	) name8798 (
		_w9245_,
		_w9259_,
		_w9260_
	);
	LUT2 #(
		.INIT('h2)
	) name8799 (
		_w3450_,
		_w9260_,
		_w9261_
	);
	LUT2 #(
		.INIT('h1)
	) name8800 (
		_w9240_,
		_w9261_,
		_w9262_
	);
	LUT2 #(
		.INIT('h2)
	) name8801 (
		\P1_state_reg[0]/NET0131 ,
		_w9262_,
		_w9263_
	);
	LUT2 #(
		.INIT('h1)
	) name8802 (
		_w9239_,
		_w9263_,
		_w9264_
	);
	LUT2 #(
		.INIT('h2)
	) name8803 (
		\P1_reg2_reg[11]/NET0131 ,
		_w3435_,
		_w9265_
	);
	LUT2 #(
		.INIT('h8)
	) name8804 (
		\P1_reg2_reg[11]/NET0131 ,
		_w3448_,
		_w9266_
	);
	LUT2 #(
		.INIT('h2)
	) name8805 (
		\P1_reg2_reg[11]/NET0131 ,
		_w5914_,
		_w9267_
	);
	LUT2 #(
		.INIT('h2)
	) name8806 (
		\P1_reg2_reg[11]/NET0131 ,
		_w3466_,
		_w9268_
	);
	LUT2 #(
		.INIT('h8)
	) name8807 (
		_w3466_,
		_w8010_,
		_w9269_
	);
	LUT2 #(
		.INIT('h1)
	) name8808 (
		_w9268_,
		_w9269_,
		_w9270_
	);
	LUT2 #(
		.INIT('h1)
	) name8809 (
		_w3563_,
		_w9270_,
		_w9271_
	);
	LUT2 #(
		.INIT('h8)
	) name8810 (
		_w3466_,
		_w8018_,
		_w9272_
	);
	LUT2 #(
		.INIT('h1)
	) name8811 (
		_w9268_,
		_w9272_,
		_w9273_
	);
	LUT2 #(
		.INIT('h2)
	) name8812 (
		_w1936_,
		_w9273_,
		_w9274_
	);
	LUT2 #(
		.INIT('h2)
	) name8813 (
		_w3466_,
		_w8004_,
		_w9275_
	);
	LUT2 #(
		.INIT('h1)
	) name8814 (
		_w9268_,
		_w9275_,
		_w9276_
	);
	LUT2 #(
		.INIT('h1)
	) name8815 (
		_w3677_,
		_w9276_,
		_w9277_
	);
	LUT2 #(
		.INIT('h8)
	) name8816 (
		_w1198_,
		_w1880_,
		_w9278_
	);
	LUT2 #(
		.INIT('h1)
	) name8817 (
		_w8024_,
		_w9278_,
		_w9279_
	);
	LUT2 #(
		.INIT('h2)
	) name8818 (
		_w3466_,
		_w9279_,
		_w9280_
	);
	LUT2 #(
		.INIT('h8)
	) name8819 (
		_w1203_,
		_w1763_,
		_w9281_
	);
	LUT2 #(
		.INIT('h1)
	) name8820 (
		_w9267_,
		_w9281_,
		_w9282_
	);
	LUT2 #(
		.INIT('h4)
	) name8821 (
		_w9280_,
		_w9282_,
		_w9283_
	);
	LUT2 #(
		.INIT('h4)
	) name8822 (
		_w9271_,
		_w9283_,
		_w9284_
	);
	LUT2 #(
		.INIT('h1)
	) name8823 (
		_w9274_,
		_w9277_,
		_w9285_
	);
	LUT2 #(
		.INIT('h8)
	) name8824 (
		_w9284_,
		_w9285_,
		_w9286_
	);
	LUT2 #(
		.INIT('h2)
	) name8825 (
		_w3450_,
		_w9286_,
		_w9287_
	);
	LUT2 #(
		.INIT('h1)
	) name8826 (
		_w9266_,
		_w9287_,
		_w9288_
	);
	LUT2 #(
		.INIT('h2)
	) name8827 (
		\P1_state_reg[0]/NET0131 ,
		_w9288_,
		_w9289_
	);
	LUT2 #(
		.INIT('h1)
	) name8828 (
		_w9265_,
		_w9289_,
		_w9290_
	);
	LUT2 #(
		.INIT('h2)
	) name8829 (
		\P1_reg2_reg[14]/NET0131 ,
		_w3435_,
		_w9291_
	);
	LUT2 #(
		.INIT('h8)
	) name8830 (
		\P1_reg2_reg[14]/NET0131 ,
		_w3448_,
		_w9292_
	);
	LUT2 #(
		.INIT('h2)
	) name8831 (
		\P1_reg2_reg[14]/NET0131 ,
		_w3718_,
		_w9293_
	);
	LUT2 #(
		.INIT('h2)
	) name8832 (
		\P1_reg2_reg[14]/NET0131 ,
		_w3466_,
		_w9294_
	);
	LUT2 #(
		.INIT('h2)
	) name8833 (
		_w3466_,
		_w8047_,
		_w9295_
	);
	LUT2 #(
		.INIT('h1)
	) name8834 (
		_w9294_,
		_w9295_,
		_w9296_
	);
	LUT2 #(
		.INIT('h2)
	) name8835 (
		_w1936_,
		_w9296_,
		_w9297_
	);
	LUT2 #(
		.INIT('h2)
	) name8836 (
		_w3466_,
		_w8058_,
		_w9298_
	);
	LUT2 #(
		.INIT('h1)
	) name8837 (
		_w9294_,
		_w9298_,
		_w9299_
	);
	LUT2 #(
		.INIT('h1)
	) name8838 (
		_w3466_,
		_w3563_,
		_w9300_
	);
	LUT2 #(
		.INIT('h2)
	) name8839 (
		_w8062_,
		_w9300_,
		_w9301_
	);
	LUT2 #(
		.INIT('h1)
	) name8840 (
		_w9299_,
		_w9301_,
		_w9302_
	);
	LUT2 #(
		.INIT('h8)
	) name8841 (
		_w3466_,
		_w8067_,
		_w9303_
	);
	LUT2 #(
		.INIT('h1)
	) name8842 (
		_w9294_,
		_w9303_,
		_w9304_
	);
	LUT2 #(
		.INIT('h2)
	) name8843 (
		_w3712_,
		_w9304_,
		_w9305_
	);
	LUT2 #(
		.INIT('h8)
	) name8844 (
		_w1113_,
		_w1763_,
		_w9306_
	);
	LUT2 #(
		.INIT('h8)
	) name8845 (
		_w1109_,
		_w1880_,
		_w9307_
	);
	LUT2 #(
		.INIT('h8)
	) name8846 (
		_w3466_,
		_w9307_,
		_w9308_
	);
	LUT2 #(
		.INIT('h1)
	) name8847 (
		_w9306_,
		_w9308_,
		_w9309_
	);
	LUT2 #(
		.INIT('h4)
	) name8848 (
		_w9293_,
		_w9309_,
		_w9310_
	);
	LUT2 #(
		.INIT('h4)
	) name8849 (
		_w9305_,
		_w9310_,
		_w9311_
	);
	LUT2 #(
		.INIT('h4)
	) name8850 (
		_w9297_,
		_w9311_,
		_w9312_
	);
	LUT2 #(
		.INIT('h4)
	) name8851 (
		_w9302_,
		_w9312_,
		_w9313_
	);
	LUT2 #(
		.INIT('h2)
	) name8852 (
		_w3450_,
		_w9313_,
		_w9314_
	);
	LUT2 #(
		.INIT('h1)
	) name8853 (
		_w9292_,
		_w9314_,
		_w9315_
	);
	LUT2 #(
		.INIT('h2)
	) name8854 (
		\P1_state_reg[0]/NET0131 ,
		_w9315_,
		_w9316_
	);
	LUT2 #(
		.INIT('h1)
	) name8855 (
		_w9291_,
		_w9316_,
		_w9317_
	);
	LUT2 #(
		.INIT('h2)
	) name8856 (
		\P1_reg2_reg[15]/NET0131 ,
		_w3435_,
		_w9318_
	);
	LUT2 #(
		.INIT('h8)
	) name8857 (
		\P1_reg2_reg[15]/NET0131 ,
		_w3448_,
		_w9319_
	);
	LUT2 #(
		.INIT('h2)
	) name8858 (
		\P1_reg2_reg[15]/NET0131 ,
		_w5914_,
		_w9320_
	);
	LUT2 #(
		.INIT('h2)
	) name8859 (
		\P1_reg2_reg[15]/NET0131 ,
		_w3466_,
		_w9321_
	);
	LUT2 #(
		.INIT('h8)
	) name8860 (
		_w3466_,
		_w8094_,
		_w9322_
	);
	LUT2 #(
		.INIT('h1)
	) name8861 (
		_w9321_,
		_w9322_,
		_w9323_
	);
	LUT2 #(
		.INIT('h1)
	) name8862 (
		_w3563_,
		_w9323_,
		_w9324_
	);
	LUT2 #(
		.INIT('h8)
	) name8863 (
		_w3466_,
		_w8102_,
		_w9325_
	);
	LUT2 #(
		.INIT('h1)
	) name8864 (
		_w9321_,
		_w9325_,
		_w9326_
	);
	LUT2 #(
		.INIT('h2)
	) name8865 (
		_w1936_,
		_w9326_,
		_w9327_
	);
	LUT2 #(
		.INIT('h2)
	) name8866 (
		_w3466_,
		_w8088_,
		_w9328_
	);
	LUT2 #(
		.INIT('h1)
	) name8867 (
		_w9321_,
		_w9328_,
		_w9329_
	);
	LUT2 #(
		.INIT('h1)
	) name8868 (
		_w3677_,
		_w9329_,
		_w9330_
	);
	LUT2 #(
		.INIT('h8)
	) name8869 (
		_w1083_,
		_w1880_,
		_w9331_
	);
	LUT2 #(
		.INIT('h1)
	) name8870 (
		_w8108_,
		_w9331_,
		_w9332_
	);
	LUT2 #(
		.INIT('h2)
	) name8871 (
		_w3466_,
		_w9332_,
		_w9333_
	);
	LUT2 #(
		.INIT('h8)
	) name8872 (
		_w1088_,
		_w1763_,
		_w9334_
	);
	LUT2 #(
		.INIT('h1)
	) name8873 (
		_w9320_,
		_w9334_,
		_w9335_
	);
	LUT2 #(
		.INIT('h4)
	) name8874 (
		_w9333_,
		_w9335_,
		_w9336_
	);
	LUT2 #(
		.INIT('h4)
	) name8875 (
		_w9324_,
		_w9336_,
		_w9337_
	);
	LUT2 #(
		.INIT('h1)
	) name8876 (
		_w9327_,
		_w9330_,
		_w9338_
	);
	LUT2 #(
		.INIT('h8)
	) name8877 (
		_w9337_,
		_w9338_,
		_w9339_
	);
	LUT2 #(
		.INIT('h2)
	) name8878 (
		_w3450_,
		_w9339_,
		_w9340_
	);
	LUT2 #(
		.INIT('h1)
	) name8879 (
		_w9319_,
		_w9340_,
		_w9341_
	);
	LUT2 #(
		.INIT('h2)
	) name8880 (
		\P1_state_reg[0]/NET0131 ,
		_w9341_,
		_w9342_
	);
	LUT2 #(
		.INIT('h1)
	) name8881 (
		_w9318_,
		_w9342_,
		_w9343_
	);
	LUT2 #(
		.INIT('h8)
	) name8882 (
		_w3411_,
		_w8252_,
		_w9344_
	);
	LUT2 #(
		.INIT('h8)
	) name8883 (
		_w2470_,
		_w3358_,
		_w9345_
	);
	LUT2 #(
		.INIT('h1)
	) name8884 (
		_w3320_,
		_w8264_,
		_w9346_
	);
	LUT2 #(
		.INIT('h4)
	) name8885 (
		_w3177_,
		_w8258_,
		_w9347_
	);
	LUT2 #(
		.INIT('h1)
	) name8886 (
		_w8270_,
		_w9345_,
		_w9348_
	);
	LUT2 #(
		.INIT('h4)
	) name8887 (
		_w9346_,
		_w9348_,
		_w9349_
	);
	LUT2 #(
		.INIT('h4)
	) name8888 (
		_w9347_,
		_w9349_,
		_w9350_
	);
	LUT2 #(
		.INIT('h4)
	) name8889 (
		_w9344_,
		_w9350_,
		_w9351_
	);
	LUT2 #(
		.INIT('h2)
	) name8890 (
		_w5860_,
		_w9351_,
		_w9352_
	);
	LUT2 #(
		.INIT('h8)
	) name8891 (
		_w7510_,
		_w8385_,
		_w9353_
	);
	LUT2 #(
		.INIT('h4)
	) name8892 (
		_w9344_,
		_w9353_,
		_w9354_
	);
	LUT2 #(
		.INIT('h2)
	) name8893 (
		\P2_reg0_reg[8]/NET0131 ,
		_w9354_,
		_w9355_
	);
	LUT2 #(
		.INIT('h1)
	) name8894 (
		_w9352_,
		_w9355_,
		_w9356_
	);
	LUT2 #(
		.INIT('h2)
	) name8895 (
		\P2_reg1_reg[15]/NET0131 ,
		_w1983_,
		_w9357_
	);
	LUT2 #(
		.INIT('h8)
	) name8896 (
		\P2_reg1_reg[15]/NET0131 ,
		_w2024_,
		_w9358_
	);
	LUT2 #(
		.INIT('h8)
	) name8897 (
		_w2843_,
		_w3358_,
		_w9359_
	);
	LUT2 #(
		.INIT('h1)
	) name8898 (
		_w3320_,
		_w8228_,
		_w9360_
	);
	LUT2 #(
		.INIT('h1)
	) name8899 (
		_w9359_,
		_w9360_,
		_w9361_
	);
	LUT2 #(
		.INIT('h2)
	) name8900 (
		_w3733_,
		_w9361_,
		_w9362_
	);
	LUT2 #(
		.INIT('h2)
	) name8901 (
		\P2_reg1_reg[15]/NET0131 ,
		_w3733_,
		_w9363_
	);
	LUT2 #(
		.INIT('h8)
	) name8902 (
		_w3733_,
		_w8211_,
		_w9364_
	);
	LUT2 #(
		.INIT('h1)
	) name8903 (
		_w9363_,
		_w9364_,
		_w9365_
	);
	LUT2 #(
		.INIT('h2)
	) name8904 (
		_w3411_,
		_w9365_,
		_w9366_
	);
	LUT2 #(
		.INIT('h8)
	) name8905 (
		_w3733_,
		_w8217_,
		_w9367_
	);
	LUT2 #(
		.INIT('h1)
	) name8906 (
		_w9363_,
		_w9367_,
		_w9368_
	);
	LUT2 #(
		.INIT('h1)
	) name8907 (
		_w3177_,
		_w9368_,
		_w9369_
	);
	LUT2 #(
		.INIT('h8)
	) name8908 (
		_w3733_,
		_w8222_,
		_w9370_
	);
	LUT2 #(
		.INIT('h1)
	) name8909 (
		_w9363_,
		_w9370_,
		_w9371_
	);
	LUT2 #(
		.INIT('h2)
	) name8910 (
		_w3355_,
		_w9371_,
		_w9372_
	);
	LUT2 #(
		.INIT('h2)
	) name8911 (
		\P2_reg1_reg[15]/NET0131 ,
		_w8531_,
		_w9373_
	);
	LUT2 #(
		.INIT('h1)
	) name8912 (
		_w9362_,
		_w9373_,
		_w9374_
	);
	LUT2 #(
		.INIT('h4)
	) name8913 (
		_w9372_,
		_w9374_,
		_w9375_
	);
	LUT2 #(
		.INIT('h4)
	) name8914 (
		_w9366_,
		_w9375_,
		_w9376_
	);
	LUT2 #(
		.INIT('h4)
	) name8915 (
		_w9369_,
		_w9376_,
		_w9377_
	);
	LUT2 #(
		.INIT('h2)
	) name8916 (
		_w2026_,
		_w9377_,
		_w9378_
	);
	LUT2 #(
		.INIT('h1)
	) name8917 (
		_w9358_,
		_w9378_,
		_w9379_
	);
	LUT2 #(
		.INIT('h2)
	) name8918 (
		\P1_state_reg[0]/NET0131 ,
		_w9379_,
		_w9380_
	);
	LUT2 #(
		.INIT('h1)
	) name8919 (
		_w9357_,
		_w9380_,
		_w9381_
	);
	LUT2 #(
		.INIT('h2)
	) name8920 (
		\P2_reg1_reg[8]/NET0131 ,
		_w1983_,
		_w9382_
	);
	LUT2 #(
		.INIT('h8)
	) name8921 (
		\P2_reg1_reg[8]/NET0131 ,
		_w2024_,
		_w9383_
	);
	LUT2 #(
		.INIT('h2)
	) name8922 (
		\P2_reg1_reg[8]/NET0131 ,
		_w8534_,
		_w9384_
	);
	LUT2 #(
		.INIT('h2)
	) name8923 (
		_w3733_,
		_w9351_,
		_w9385_
	);
	LUT2 #(
		.INIT('h1)
	) name8924 (
		_w9384_,
		_w9385_,
		_w9386_
	);
	LUT2 #(
		.INIT('h2)
	) name8925 (
		_w2026_,
		_w9386_,
		_w9387_
	);
	LUT2 #(
		.INIT('h1)
	) name8926 (
		_w9383_,
		_w9387_,
		_w9388_
	);
	LUT2 #(
		.INIT('h2)
	) name8927 (
		\P1_state_reg[0]/NET0131 ,
		_w9388_,
		_w9389_
	);
	LUT2 #(
		.INIT('h1)
	) name8928 (
		_w9382_,
		_w9389_,
		_w9390_
	);
	LUT2 #(
		.INIT('h2)
	) name8929 (
		\P2_reg2_reg[11]/NET0131 ,
		_w1983_,
		_w9391_
	);
	LUT2 #(
		.INIT('h8)
	) name8930 (
		\P2_reg2_reg[11]/NET0131 ,
		_w2024_,
		_w9392_
	);
	LUT2 #(
		.INIT('h2)
	) name8931 (
		\P2_reg2_reg[11]/NET0131 ,
		_w3774_,
		_w9393_
	);
	LUT2 #(
		.INIT('h2)
	) name8932 (
		\P2_reg2_reg[11]/NET0131 ,
		_w3758_,
		_w9394_
	);
	LUT2 #(
		.INIT('h8)
	) name8933 (
		_w3758_,
		_w8129_,
		_w9395_
	);
	LUT2 #(
		.INIT('h1)
	) name8934 (
		_w9394_,
		_w9395_,
		_w9396_
	);
	LUT2 #(
		.INIT('h2)
	) name8935 (
		_w3411_,
		_w9396_,
		_w9397_
	);
	LUT2 #(
		.INIT('h8)
	) name8936 (
		_w3758_,
		_w8135_,
		_w9398_
	);
	LUT2 #(
		.INIT('h1)
	) name8937 (
		_w9394_,
		_w9398_,
		_w9399_
	);
	LUT2 #(
		.INIT('h1)
	) name8938 (
		_w3177_,
		_w9399_,
		_w9400_
	);
	LUT2 #(
		.INIT('h8)
	) name8939 (
		_w3758_,
		_w8140_,
		_w9401_
	);
	LUT2 #(
		.INIT('h1)
	) name8940 (
		_w9394_,
		_w9401_,
		_w9402_
	);
	LUT2 #(
		.INIT('h2)
	) name8941 (
		_w3355_,
		_w9402_,
		_w9403_
	);
	LUT2 #(
		.INIT('h2)
	) name8942 (
		_w3758_,
		_w8146_,
		_w9404_
	);
	LUT2 #(
		.INIT('h1)
	) name8943 (
		_w9394_,
		_w9404_,
		_w9405_
	);
	LUT2 #(
		.INIT('h1)
	) name8944 (
		_w3320_,
		_w9405_,
		_w9406_
	);
	LUT2 #(
		.INIT('h8)
	) name8945 (
		_w2681_,
		_w3420_,
		_w9407_
	);
	LUT2 #(
		.INIT('h8)
	) name8946 (
		_w2704_,
		_w3358_,
		_w9408_
	);
	LUT2 #(
		.INIT('h8)
	) name8947 (
		_w3758_,
		_w9408_,
		_w9409_
	);
	LUT2 #(
		.INIT('h1)
	) name8948 (
		_w9393_,
		_w9407_,
		_w9410_
	);
	LUT2 #(
		.INIT('h4)
	) name8949 (
		_w9409_,
		_w9410_,
		_w9411_
	);
	LUT2 #(
		.INIT('h4)
	) name8950 (
		_w9406_,
		_w9411_,
		_w9412_
	);
	LUT2 #(
		.INIT('h4)
	) name8951 (
		_w9403_,
		_w9412_,
		_w9413_
	);
	LUT2 #(
		.INIT('h4)
	) name8952 (
		_w9400_,
		_w9413_,
		_w9414_
	);
	LUT2 #(
		.INIT('h4)
	) name8953 (
		_w9397_,
		_w9414_,
		_w9415_
	);
	LUT2 #(
		.INIT('h2)
	) name8954 (
		_w2026_,
		_w9415_,
		_w9416_
	);
	LUT2 #(
		.INIT('h1)
	) name8955 (
		_w9392_,
		_w9416_,
		_w9417_
	);
	LUT2 #(
		.INIT('h2)
	) name8956 (
		\P1_state_reg[0]/NET0131 ,
		_w9417_,
		_w9418_
	);
	LUT2 #(
		.INIT('h1)
	) name8957 (
		_w9391_,
		_w9418_,
		_w9419_
	);
	LUT2 #(
		.INIT('h2)
	) name8958 (
		\P2_reg2_reg[14]/NET0131 ,
		_w1983_,
		_w9420_
	);
	LUT2 #(
		.INIT('h8)
	) name8959 (
		\P2_reg2_reg[14]/NET0131 ,
		_w2024_,
		_w9421_
	);
	LUT2 #(
		.INIT('h2)
	) name8960 (
		\P2_reg2_reg[14]/NET0131 ,
		_w3774_,
		_w9422_
	);
	LUT2 #(
		.INIT('h2)
	) name8961 (
		\P2_reg2_reg[14]/NET0131 ,
		_w3758_,
		_w9423_
	);
	LUT2 #(
		.INIT('h8)
	) name8962 (
		_w3758_,
		_w8171_,
		_w9424_
	);
	LUT2 #(
		.INIT('h1)
	) name8963 (
		_w9423_,
		_w9424_,
		_w9425_
	);
	LUT2 #(
		.INIT('h2)
	) name8964 (
		_w3411_,
		_w9425_,
		_w9426_
	);
	LUT2 #(
		.INIT('h8)
	) name8965 (
		_w3758_,
		_w8176_,
		_w9427_
	);
	LUT2 #(
		.INIT('h1)
	) name8966 (
		_w9423_,
		_w9427_,
		_w9428_
	);
	LUT2 #(
		.INIT('h2)
	) name8967 (
		_w3355_,
		_w9428_,
		_w9429_
	);
	LUT2 #(
		.INIT('h8)
	) name8968 (
		_w3758_,
		_w8182_,
		_w9430_
	);
	LUT2 #(
		.INIT('h1)
	) name8969 (
		_w9423_,
		_w9430_,
		_w9431_
	);
	LUT2 #(
		.INIT('h1)
	) name8970 (
		_w3177_,
		_w9431_,
		_w9432_
	);
	LUT2 #(
		.INIT('h2)
	) name8971 (
		_w3758_,
		_w8188_,
		_w9433_
	);
	LUT2 #(
		.INIT('h1)
	) name8972 (
		_w9423_,
		_w9433_,
		_w9434_
	);
	LUT2 #(
		.INIT('h1)
	) name8973 (
		_w3320_,
		_w9434_,
		_w9435_
	);
	LUT2 #(
		.INIT('h8)
	) name8974 (
		_w2866_,
		_w3420_,
		_w9436_
	);
	LUT2 #(
		.INIT('h8)
	) name8975 (
		_w2860_,
		_w3358_,
		_w9437_
	);
	LUT2 #(
		.INIT('h8)
	) name8976 (
		_w3758_,
		_w9437_,
		_w9438_
	);
	LUT2 #(
		.INIT('h1)
	) name8977 (
		_w9422_,
		_w9436_,
		_w9439_
	);
	LUT2 #(
		.INIT('h4)
	) name8978 (
		_w9438_,
		_w9439_,
		_w9440_
	);
	LUT2 #(
		.INIT('h4)
	) name8979 (
		_w9426_,
		_w9440_,
		_w9441_
	);
	LUT2 #(
		.INIT('h1)
	) name8980 (
		_w9429_,
		_w9432_,
		_w9442_
	);
	LUT2 #(
		.INIT('h4)
	) name8981 (
		_w9435_,
		_w9442_,
		_w9443_
	);
	LUT2 #(
		.INIT('h8)
	) name8982 (
		_w9441_,
		_w9443_,
		_w9444_
	);
	LUT2 #(
		.INIT('h2)
	) name8983 (
		_w2026_,
		_w9444_,
		_w9445_
	);
	LUT2 #(
		.INIT('h1)
	) name8984 (
		_w9421_,
		_w9445_,
		_w9446_
	);
	LUT2 #(
		.INIT('h2)
	) name8985 (
		\P1_state_reg[0]/NET0131 ,
		_w9446_,
		_w9447_
	);
	LUT2 #(
		.INIT('h1)
	) name8986 (
		_w9420_,
		_w9447_,
		_w9448_
	);
	LUT2 #(
		.INIT('h2)
	) name8987 (
		\P2_reg2_reg[8]/NET0131 ,
		_w1983_,
		_w9449_
	);
	LUT2 #(
		.INIT('h8)
	) name8988 (
		\P2_reg2_reg[8]/NET0131 ,
		_w2024_,
		_w9450_
	);
	LUT2 #(
		.INIT('h8)
	) name8989 (
		_w3758_,
		_w9345_,
		_w9451_
	);
	LUT2 #(
		.INIT('h2)
	) name8990 (
		\P2_reg2_reg[8]/NET0131 ,
		_w3758_,
		_w9452_
	);
	LUT2 #(
		.INIT('h8)
	) name8991 (
		_w3758_,
		_w8252_,
		_w9453_
	);
	LUT2 #(
		.INIT('h1)
	) name8992 (
		_w9452_,
		_w9453_,
		_w9454_
	);
	LUT2 #(
		.INIT('h2)
	) name8993 (
		_w3411_,
		_w9454_,
		_w9455_
	);
	LUT2 #(
		.INIT('h8)
	) name8994 (
		_w3758_,
		_w8258_,
		_w9456_
	);
	LUT2 #(
		.INIT('h1)
	) name8995 (
		_w9452_,
		_w9456_,
		_w9457_
	);
	LUT2 #(
		.INIT('h1)
	) name8996 (
		_w3177_,
		_w9457_,
		_w9458_
	);
	LUT2 #(
		.INIT('h2)
	) name8997 (
		_w3758_,
		_w8264_,
		_w9459_
	);
	LUT2 #(
		.INIT('h1)
	) name8998 (
		_w9452_,
		_w9459_,
		_w9460_
	);
	LUT2 #(
		.INIT('h1)
	) name8999 (
		_w3320_,
		_w9460_,
		_w9461_
	);
	LUT2 #(
		.INIT('h8)
	) name9000 (
		_w3758_,
		_w8269_,
		_w9462_
	);
	LUT2 #(
		.INIT('h1)
	) name9001 (
		_w9452_,
		_w9462_,
		_w9463_
	);
	LUT2 #(
		.INIT('h2)
	) name9002 (
		_w3355_,
		_w9463_,
		_w9464_
	);
	LUT2 #(
		.INIT('h8)
	) name9003 (
		_w2447_,
		_w3420_,
		_w9465_
	);
	LUT2 #(
		.INIT('h2)
	) name9004 (
		\P2_reg2_reg[8]/NET0131 ,
		_w3774_,
		_w9466_
	);
	LUT2 #(
		.INIT('h1)
	) name9005 (
		_w9451_,
		_w9465_,
		_w9467_
	);
	LUT2 #(
		.INIT('h4)
	) name9006 (
		_w9466_,
		_w9467_,
		_w9468_
	);
	LUT2 #(
		.INIT('h4)
	) name9007 (
		_w9464_,
		_w9468_,
		_w9469_
	);
	LUT2 #(
		.INIT('h4)
	) name9008 (
		_w9458_,
		_w9469_,
		_w9470_
	);
	LUT2 #(
		.INIT('h4)
	) name9009 (
		_w9461_,
		_w9470_,
		_w9471_
	);
	LUT2 #(
		.INIT('h4)
	) name9010 (
		_w9455_,
		_w9471_,
		_w9472_
	);
	LUT2 #(
		.INIT('h2)
	) name9011 (
		_w2026_,
		_w9472_,
		_w9473_
	);
	LUT2 #(
		.INIT('h1)
	) name9012 (
		_w9450_,
		_w9473_,
		_w9474_
	);
	LUT2 #(
		.INIT('h2)
	) name9013 (
		\P1_state_reg[0]/NET0131 ,
		_w9474_,
		_w9475_
	);
	LUT2 #(
		.INIT('h1)
	) name9014 (
		_w9449_,
		_w9475_,
		_w9476_
	);
	LUT2 #(
		.INIT('h2)
	) name9015 (
		\P1_reg0_reg[15]/NET0131 ,
		_w3435_,
		_w9477_
	);
	LUT2 #(
		.INIT('h8)
	) name9016 (
		\P1_reg0_reg[15]/NET0131 ,
		_w3448_,
		_w9478_
	);
	LUT2 #(
		.INIT('h2)
	) name9017 (
		\P1_reg0_reg[15]/NET0131 ,
		_w4494_,
		_w9479_
	);
	LUT2 #(
		.INIT('h2)
	) name9018 (
		\P1_reg0_reg[15]/NET0131 ,
		_w4396_,
		_w9480_
	);
	LUT2 #(
		.INIT('h8)
	) name9019 (
		_w4396_,
		_w8094_,
		_w9481_
	);
	LUT2 #(
		.INIT('h1)
	) name9020 (
		_w9480_,
		_w9481_,
		_w9482_
	);
	LUT2 #(
		.INIT('h1)
	) name9021 (
		_w3563_,
		_w9482_,
		_w9483_
	);
	LUT2 #(
		.INIT('h8)
	) name9022 (
		_w4396_,
		_w8102_,
		_w9484_
	);
	LUT2 #(
		.INIT('h1)
	) name9023 (
		_w9480_,
		_w9484_,
		_w9485_
	);
	LUT2 #(
		.INIT('h2)
	) name9024 (
		_w1936_,
		_w9485_,
		_w9486_
	);
	LUT2 #(
		.INIT('h2)
	) name9025 (
		_w4396_,
		_w8088_,
		_w9487_
	);
	LUT2 #(
		.INIT('h1)
	) name9026 (
		_w9480_,
		_w9487_,
		_w9488_
	);
	LUT2 #(
		.INIT('h1)
	) name9027 (
		_w3677_,
		_w9488_,
		_w9489_
	);
	LUT2 #(
		.INIT('h2)
	) name9028 (
		_w4396_,
		_w9332_,
		_w9490_
	);
	LUT2 #(
		.INIT('h1)
	) name9029 (
		_w9479_,
		_w9490_,
		_w9491_
	);
	LUT2 #(
		.INIT('h4)
	) name9030 (
		_w9483_,
		_w9491_,
		_w9492_
	);
	LUT2 #(
		.INIT('h1)
	) name9031 (
		_w9486_,
		_w9489_,
		_w9493_
	);
	LUT2 #(
		.INIT('h8)
	) name9032 (
		_w9492_,
		_w9493_,
		_w9494_
	);
	LUT2 #(
		.INIT('h2)
	) name9033 (
		_w3450_,
		_w9494_,
		_w9495_
	);
	LUT2 #(
		.INIT('h1)
	) name9034 (
		_w9478_,
		_w9495_,
		_w9496_
	);
	LUT2 #(
		.INIT('h2)
	) name9035 (
		\P1_state_reg[0]/NET0131 ,
		_w9496_,
		_w9497_
	);
	LUT2 #(
		.INIT('h1)
	) name9036 (
		_w9477_,
		_w9497_,
		_w9498_
	);
	LUT2 #(
		.INIT('h2)
	) name9037 (
		\P1_reg0_reg[8]/NET0131 ,
		_w3435_,
		_w9499_
	);
	LUT2 #(
		.INIT('h8)
	) name9038 (
		\P1_reg0_reg[8]/NET0131 ,
		_w3448_,
		_w9500_
	);
	LUT2 #(
		.INIT('h8)
	) name9039 (
		_w4396_,
		_w9212_,
		_w9501_
	);
	LUT2 #(
		.INIT('h2)
	) name9040 (
		\P1_reg0_reg[8]/NET0131 ,
		_w4396_,
		_w9502_
	);
	LUT2 #(
		.INIT('h8)
	) name9041 (
		_w4396_,
		_w8292_,
		_w9503_
	);
	LUT2 #(
		.INIT('h1)
	) name9042 (
		_w9502_,
		_w9503_,
		_w9504_
	);
	LUT2 #(
		.INIT('h2)
	) name9043 (
		_w1936_,
		_w9504_,
		_w9505_
	);
	LUT2 #(
		.INIT('h8)
	) name9044 (
		_w4396_,
		_w8298_,
		_w9506_
	);
	LUT2 #(
		.INIT('h1)
	) name9045 (
		_w9502_,
		_w9506_,
		_w9507_
	);
	LUT2 #(
		.INIT('h1)
	) name9046 (
		_w3563_,
		_w9507_,
		_w9508_
	);
	LUT2 #(
		.INIT('h2)
	) name9047 (
		_w4396_,
		_w8304_,
		_w9509_
	);
	LUT2 #(
		.INIT('h1)
	) name9048 (
		_w9502_,
		_w9509_,
		_w9510_
	);
	LUT2 #(
		.INIT('h1)
	) name9049 (
		_w3677_,
		_w9510_,
		_w9511_
	);
	LUT2 #(
		.INIT('h8)
	) name9050 (
		_w4396_,
		_w8310_,
		_w9512_
	);
	LUT2 #(
		.INIT('h1)
	) name9051 (
		_w9502_,
		_w9512_,
		_w9513_
	);
	LUT2 #(
		.INIT('h2)
	) name9052 (
		_w3712_,
		_w9513_,
		_w9514_
	);
	LUT2 #(
		.INIT('h2)
	) name9053 (
		\P1_reg0_reg[8]/NET0131 ,
		_w4493_,
		_w9515_
	);
	LUT2 #(
		.INIT('h1)
	) name9054 (
		_w9501_,
		_w9515_,
		_w9516_
	);
	LUT2 #(
		.INIT('h4)
	) name9055 (
		_w9514_,
		_w9516_,
		_w9517_
	);
	LUT2 #(
		.INIT('h4)
	) name9056 (
		_w9508_,
		_w9517_,
		_w9518_
	);
	LUT2 #(
		.INIT('h4)
	) name9057 (
		_w9511_,
		_w9518_,
		_w9519_
	);
	LUT2 #(
		.INIT('h4)
	) name9058 (
		_w9505_,
		_w9519_,
		_w9520_
	);
	LUT2 #(
		.INIT('h2)
	) name9059 (
		_w3450_,
		_w9520_,
		_w9521_
	);
	LUT2 #(
		.INIT('h1)
	) name9060 (
		_w9500_,
		_w9521_,
		_w9522_
	);
	LUT2 #(
		.INIT('h2)
	) name9061 (
		\P1_state_reg[0]/NET0131 ,
		_w9522_,
		_w9523_
	);
	LUT2 #(
		.INIT('h1)
	) name9062 (
		_w9499_,
		_w9523_,
		_w9524_
	);
	LUT2 #(
		.INIT('h2)
	) name9063 (
		\P1_reg1_reg[15]/NET0131 ,
		_w3435_,
		_w9525_
	);
	LUT2 #(
		.INIT('h8)
	) name9064 (
		\P1_reg1_reg[15]/NET0131 ,
		_w3448_,
		_w9526_
	);
	LUT2 #(
		.INIT('h2)
	) name9065 (
		\P1_reg1_reg[15]/NET0131 ,
		_w4491_,
		_w9527_
	);
	LUT2 #(
		.INIT('h2)
	) name9066 (
		\P1_reg1_reg[15]/NET0131 ,
		_w4532_,
		_w9528_
	);
	LUT2 #(
		.INIT('h8)
	) name9067 (
		_w4532_,
		_w8094_,
		_w9529_
	);
	LUT2 #(
		.INIT('h1)
	) name9068 (
		_w9528_,
		_w9529_,
		_w9530_
	);
	LUT2 #(
		.INIT('h1)
	) name9069 (
		_w3563_,
		_w9530_,
		_w9531_
	);
	LUT2 #(
		.INIT('h8)
	) name9070 (
		_w4532_,
		_w8102_,
		_w9532_
	);
	LUT2 #(
		.INIT('h1)
	) name9071 (
		_w9528_,
		_w9532_,
		_w9533_
	);
	LUT2 #(
		.INIT('h2)
	) name9072 (
		_w1936_,
		_w9533_,
		_w9534_
	);
	LUT2 #(
		.INIT('h2)
	) name9073 (
		_w4532_,
		_w8088_,
		_w9535_
	);
	LUT2 #(
		.INIT('h1)
	) name9074 (
		_w9528_,
		_w9535_,
		_w9536_
	);
	LUT2 #(
		.INIT('h1)
	) name9075 (
		_w3677_,
		_w9536_,
		_w9537_
	);
	LUT2 #(
		.INIT('h8)
	) name9076 (
		_w4532_,
		_w8107_,
		_w9538_
	);
	LUT2 #(
		.INIT('h1)
	) name9077 (
		_w9528_,
		_w9538_,
		_w9539_
	);
	LUT2 #(
		.INIT('h2)
	) name9078 (
		_w3712_,
		_w9539_,
		_w9540_
	);
	LUT2 #(
		.INIT('h8)
	) name9079 (
		_w1083_,
		_w4532_,
		_w9541_
	);
	LUT2 #(
		.INIT('h1)
	) name9080 (
		_w9528_,
		_w9541_,
		_w9542_
	);
	LUT2 #(
		.INIT('h2)
	) name9081 (
		_w1880_,
		_w9542_,
		_w9543_
	);
	LUT2 #(
		.INIT('h1)
	) name9082 (
		_w9527_,
		_w9543_,
		_w9544_
	);
	LUT2 #(
		.INIT('h4)
	) name9083 (
		_w9540_,
		_w9544_,
		_w9545_
	);
	LUT2 #(
		.INIT('h4)
	) name9084 (
		_w9531_,
		_w9545_,
		_w9546_
	);
	LUT2 #(
		.INIT('h1)
	) name9085 (
		_w9534_,
		_w9537_,
		_w9547_
	);
	LUT2 #(
		.INIT('h8)
	) name9086 (
		_w9546_,
		_w9547_,
		_w9548_
	);
	LUT2 #(
		.INIT('h2)
	) name9087 (
		_w3450_,
		_w9548_,
		_w9549_
	);
	LUT2 #(
		.INIT('h1)
	) name9088 (
		_w9526_,
		_w9549_,
		_w9550_
	);
	LUT2 #(
		.INIT('h2)
	) name9089 (
		\P1_state_reg[0]/NET0131 ,
		_w9550_,
		_w9551_
	);
	LUT2 #(
		.INIT('h1)
	) name9090 (
		_w9525_,
		_w9551_,
		_w9552_
	);
	LUT2 #(
		.INIT('h2)
	) name9091 (
		\P2_reg0_reg[15]/NET0131 ,
		_w1983_,
		_w9553_
	);
	LUT2 #(
		.INIT('h8)
	) name9092 (
		\P2_reg0_reg[15]/NET0131 ,
		_w2024_,
		_w9554_
	);
	LUT2 #(
		.INIT('h2)
	) name9093 (
		_w2040_,
		_w9361_,
		_w9555_
	);
	LUT2 #(
		.INIT('h2)
	) name9094 (
		\P2_reg0_reg[15]/NET0131 ,
		_w2040_,
		_w9556_
	);
	LUT2 #(
		.INIT('h8)
	) name9095 (
		_w2040_,
		_w8211_,
		_w9557_
	);
	LUT2 #(
		.INIT('h1)
	) name9096 (
		_w9556_,
		_w9557_,
		_w9558_
	);
	LUT2 #(
		.INIT('h2)
	) name9097 (
		_w3411_,
		_w9558_,
		_w9559_
	);
	LUT2 #(
		.INIT('h8)
	) name9098 (
		_w2040_,
		_w8217_,
		_w9560_
	);
	LUT2 #(
		.INIT('h1)
	) name9099 (
		_w9556_,
		_w9560_,
		_w9561_
	);
	LUT2 #(
		.INIT('h1)
	) name9100 (
		_w3177_,
		_w9561_,
		_w9562_
	);
	LUT2 #(
		.INIT('h8)
	) name9101 (
		_w2040_,
		_w8222_,
		_w9563_
	);
	LUT2 #(
		.INIT('h1)
	) name9102 (
		_w9556_,
		_w9563_,
		_w9564_
	);
	LUT2 #(
		.INIT('h2)
	) name9103 (
		_w3355_,
		_w9564_,
		_w9565_
	);
	LUT2 #(
		.INIT('h2)
	) name9104 (
		\P2_reg0_reg[15]/NET0131 ,
		_w7506_,
		_w9566_
	);
	LUT2 #(
		.INIT('h1)
	) name9105 (
		_w9555_,
		_w9566_,
		_w9567_
	);
	LUT2 #(
		.INIT('h4)
	) name9106 (
		_w9565_,
		_w9567_,
		_w9568_
	);
	LUT2 #(
		.INIT('h4)
	) name9107 (
		_w9559_,
		_w9568_,
		_w9569_
	);
	LUT2 #(
		.INIT('h4)
	) name9108 (
		_w9562_,
		_w9569_,
		_w9570_
	);
	LUT2 #(
		.INIT('h2)
	) name9109 (
		_w2026_,
		_w9570_,
		_w9571_
	);
	LUT2 #(
		.INIT('h1)
	) name9110 (
		_w9554_,
		_w9571_,
		_w9572_
	);
	LUT2 #(
		.INIT('h2)
	) name9111 (
		\P1_state_reg[0]/NET0131 ,
		_w9572_,
		_w9573_
	);
	LUT2 #(
		.INIT('h1)
	) name9112 (
		_w9553_,
		_w9573_,
		_w9574_
	);
	LUT2 #(
		.INIT('h4)
	) name9113 (
		\P1_state_reg[0]/NET0131 ,
		\P2_reg3_reg[3]/NET0131 ,
		_w9575_
	);
	LUT2 #(
		.INIT('h4)
	) name9114 (
		\P2_reg3_reg[3]/NET0131 ,
		_w2024_,
		_w9576_
	);
	LUT2 #(
		.INIT('h4)
	) name9115 (
		_w2631_,
		_w3358_,
		_w9577_
	);
	LUT2 #(
		.INIT('h1)
	) name9116 (
		_w3260_,
		_w3261_,
		_w9578_
	);
	LUT2 #(
		.INIT('h4)
	) name9117 (
		_w4193_,
		_w9578_,
		_w9579_
	);
	LUT2 #(
		.INIT('h2)
	) name9118 (
		_w4193_,
		_w9578_,
		_w9580_
	);
	LUT2 #(
		.INIT('h1)
	) name9119 (
		_w9579_,
		_w9580_,
		_w9581_
	);
	LUT2 #(
		.INIT('h1)
	) name9120 (
		_w3320_,
		_w9581_,
		_w9582_
	);
	LUT2 #(
		.INIT('h1)
	) name9121 (
		_w2631_,
		_w3327_,
		_w9583_
	);
	LUT2 #(
		.INIT('h4)
	) name9122 (
		_w3328_,
		_w3355_,
		_w9584_
	);
	LUT2 #(
		.INIT('h4)
	) name9123 (
		_w9583_,
		_w9584_,
		_w9585_
	);
	LUT2 #(
		.INIT('h1)
	) name9124 (
		_w9577_,
		_w9585_,
		_w9586_
	);
	LUT2 #(
		.INIT('h4)
	) name9125 (
		_w9582_,
		_w9586_,
		_w9587_
	);
	LUT2 #(
		.INIT('h1)
	) name9126 (
		_w2608_,
		_w2609_,
		_w9588_
	);
	LUT2 #(
		.INIT('h8)
	) name9127 (
		_w4193_,
		_w9588_,
		_w9589_
	);
	LUT2 #(
		.INIT('h1)
	) name9128 (
		_w4193_,
		_w9588_,
		_w9590_
	);
	LUT2 #(
		.INIT('h1)
	) name9129 (
		_w9589_,
		_w9590_,
		_w9591_
	);
	LUT2 #(
		.INIT('h1)
	) name9130 (
		_w3177_,
		_w9591_,
		_w9592_
	);
	LUT2 #(
		.INIT('h2)
	) name9131 (
		_w2642_,
		_w3376_,
		_w9593_
	);
	LUT2 #(
		.INIT('h1)
	) name9132 (
		_w8941_,
		_w9593_,
		_w9594_
	);
	LUT2 #(
		.INIT('h1)
	) name9133 (
		_w2058_,
		_w9594_,
		_w9595_
	);
	LUT2 #(
		.INIT('h8)
	) name9134 (
		_w2058_,
		_w2552_,
		_w9596_
	);
	LUT2 #(
		.INIT('h1)
	) name9135 (
		_w9595_,
		_w9596_,
		_w9597_
	);
	LUT2 #(
		.INIT('h8)
	) name9136 (
		_w3411_,
		_w9597_,
		_w9598_
	);
	LUT2 #(
		.INIT('h2)
	) name9137 (
		_w9587_,
		_w9592_,
		_w9599_
	);
	LUT2 #(
		.INIT('h4)
	) name9138 (
		_w9598_,
		_w9599_,
		_w9600_
	);
	LUT2 #(
		.INIT('h2)
	) name9139 (
		_w3788_,
		_w9600_,
		_w9601_
	);
	LUT2 #(
		.INIT('h4)
	) name9140 (
		\P2_reg3_reg[3]/NET0131 ,
		_w3417_,
		_w9602_
	);
	LUT2 #(
		.INIT('h4)
	) name9141 (
		_w2631_,
		_w3420_,
		_w9603_
	);
	LUT2 #(
		.INIT('h1)
	) name9142 (
		\P2_reg3_reg[3]/NET0131 ,
		_w3788_,
		_w9604_
	);
	LUT2 #(
		.INIT('h4)
	) name9143 (
		_w6641_,
		_w9604_,
		_w9605_
	);
	LUT2 #(
		.INIT('h1)
	) name9144 (
		_w9602_,
		_w9603_,
		_w9606_
	);
	LUT2 #(
		.INIT('h4)
	) name9145 (
		_w9605_,
		_w9606_,
		_w9607_
	);
	LUT2 #(
		.INIT('h4)
	) name9146 (
		_w9601_,
		_w9607_,
		_w9608_
	);
	LUT2 #(
		.INIT('h2)
	) name9147 (
		_w2026_,
		_w9608_,
		_w9609_
	);
	LUT2 #(
		.INIT('h1)
	) name9148 (
		_w9576_,
		_w9609_,
		_w9610_
	);
	LUT2 #(
		.INIT('h2)
	) name9149 (
		\P1_state_reg[0]/NET0131 ,
		_w9610_,
		_w9611_
	);
	LUT2 #(
		.INIT('h4)
	) name9150 (
		\P2_reg3_reg[3]/NET0131 ,
		_w3976_,
		_w9612_
	);
	LUT2 #(
		.INIT('h1)
	) name9151 (
		_w9575_,
		_w9612_,
		_w9613_
	);
	LUT2 #(
		.INIT('h4)
	) name9152 (
		_w9611_,
		_w9613_,
		_w9614_
	);
	LUT2 #(
		.INIT('h4)
	) name9153 (
		\P1_state_reg[0]/NET0131 ,
		\P2_reg3_reg[6]/NET0131 ,
		_w9615_
	);
	LUT2 #(
		.INIT('h8)
	) name9154 (
		_w2499_,
		_w3976_,
		_w9616_
	);
	LUT2 #(
		.INIT('h8)
	) name9155 (
		_w2024_,
		_w2499_,
		_w9617_
	);
	LUT2 #(
		.INIT('h1)
	) name9156 (
		_w2521_,
		_w3965_,
		_w9618_
	);
	LUT2 #(
		.INIT('h2)
	) name9157 (
		_w2499_,
		_w3788_,
		_w9619_
	);
	LUT2 #(
		.INIT('h2)
	) name9158 (
		_w2480_,
		_w3379_,
		_w9620_
	);
	LUT2 #(
		.INIT('h1)
	) name9159 (
		_w3380_,
		_w9620_,
		_w9621_
	);
	LUT2 #(
		.INIT('h1)
	) name9160 (
		_w2058_,
		_w9621_,
		_w9622_
	);
	LUT2 #(
		.INIT('h8)
	) name9161 (
		_w2058_,
		_w2531_,
		_w9623_
	);
	LUT2 #(
		.INIT('h1)
	) name9162 (
		_w9622_,
		_w9623_,
		_w9624_
	);
	LUT2 #(
		.INIT('h8)
	) name9163 (
		_w3788_,
		_w9624_,
		_w9625_
	);
	LUT2 #(
		.INIT('h1)
	) name9164 (
		_w9619_,
		_w9625_,
		_w9626_
	);
	LUT2 #(
		.INIT('h2)
	) name9165 (
		_w3411_,
		_w9626_,
		_w9627_
	);
	LUT2 #(
		.INIT('h2)
	) name9166 (
		_w3827_,
		_w4205_,
		_w9628_
	);
	LUT2 #(
		.INIT('h4)
	) name9167 (
		_w3827_,
		_w4205_,
		_w9629_
	);
	LUT2 #(
		.INIT('h1)
	) name9168 (
		_w9628_,
		_w9629_,
		_w9630_
	);
	LUT2 #(
		.INIT('h2)
	) name9169 (
		_w3788_,
		_w9630_,
		_w9631_
	);
	LUT2 #(
		.INIT('h1)
	) name9170 (
		_w9619_,
		_w9631_,
		_w9632_
	);
	LUT2 #(
		.INIT('h1)
	) name9171 (
		_w3320_,
		_w9632_,
		_w9633_
	);
	LUT2 #(
		.INIT('h2)
	) name9172 (
		_w3885_,
		_w4205_,
		_w9634_
	);
	LUT2 #(
		.INIT('h4)
	) name9173 (
		_w3885_,
		_w4205_,
		_w9635_
	);
	LUT2 #(
		.INIT('h1)
	) name9174 (
		_w9634_,
		_w9635_,
		_w9636_
	);
	LUT2 #(
		.INIT('h8)
	) name9175 (
		_w3788_,
		_w9636_,
		_w9637_
	);
	LUT2 #(
		.INIT('h1)
	) name9176 (
		_w9619_,
		_w9637_,
		_w9638_
	);
	LUT2 #(
		.INIT('h1)
	) name9177 (
		_w3177_,
		_w9638_,
		_w9639_
	);
	LUT2 #(
		.INIT('h1)
	) name9178 (
		_w2521_,
		_w3330_,
		_w9640_
	);
	LUT2 #(
		.INIT('h1)
	) name9179 (
		_w3331_,
		_w9640_,
		_w9641_
	);
	LUT2 #(
		.INIT('h8)
	) name9180 (
		_w3788_,
		_w9641_,
		_w9642_
	);
	LUT2 #(
		.INIT('h1)
	) name9181 (
		_w9619_,
		_w9642_,
		_w9643_
	);
	LUT2 #(
		.INIT('h2)
	) name9182 (
		_w3355_,
		_w9643_,
		_w9644_
	);
	LUT2 #(
		.INIT('h2)
	) name9183 (
		_w2499_,
		_w3962_,
		_w9645_
	);
	LUT2 #(
		.INIT('h1)
	) name9184 (
		_w9618_,
		_w9645_,
		_w9646_
	);
	LUT2 #(
		.INIT('h4)
	) name9185 (
		_w9644_,
		_w9646_,
		_w9647_
	);
	LUT2 #(
		.INIT('h4)
	) name9186 (
		_w9633_,
		_w9647_,
		_w9648_
	);
	LUT2 #(
		.INIT('h4)
	) name9187 (
		_w9639_,
		_w9648_,
		_w9649_
	);
	LUT2 #(
		.INIT('h4)
	) name9188 (
		_w9627_,
		_w9649_,
		_w9650_
	);
	LUT2 #(
		.INIT('h2)
	) name9189 (
		_w2026_,
		_w9650_,
		_w9651_
	);
	LUT2 #(
		.INIT('h1)
	) name9190 (
		_w9617_,
		_w9651_,
		_w9652_
	);
	LUT2 #(
		.INIT('h2)
	) name9191 (
		\P1_state_reg[0]/NET0131 ,
		_w9652_,
		_w9653_
	);
	LUT2 #(
		.INIT('h1)
	) name9192 (
		_w9615_,
		_w9616_,
		_w9654_
	);
	LUT2 #(
		.INIT('h4)
	) name9193 (
		_w9653_,
		_w9654_,
		_w9655_
	);
	LUT2 #(
		.INIT('h4)
	) name9194 (
		\P1_state_reg[0]/NET0131 ,
		\P2_reg3_reg[7]/NET0131 ,
		_w9656_
	);
	LUT2 #(
		.INIT('h8)
	) name9195 (
		_w2024_,
		_w2476_,
		_w9657_
	);
	LUT2 #(
		.INIT('h2)
	) name9196 (
		_w2476_,
		_w5698_,
		_w9658_
	);
	LUT2 #(
		.INIT('h2)
	) name9197 (
		_w2476_,
		_w3788_,
		_w9659_
	);
	LUT2 #(
		.INIT('h2)
	) name9198 (
		_w2454_,
		_w3380_,
		_w9660_
	);
	LUT2 #(
		.INIT('h1)
	) name9199 (
		_w7242_,
		_w9660_,
		_w9661_
	);
	LUT2 #(
		.INIT('h1)
	) name9200 (
		_w2058_,
		_w9661_,
		_w9662_
	);
	LUT2 #(
		.INIT('h8)
	) name9201 (
		_w2058_,
		_w2506_,
		_w9663_
	);
	LUT2 #(
		.INIT('h1)
	) name9202 (
		_w9662_,
		_w9663_,
		_w9664_
	);
	LUT2 #(
		.INIT('h8)
	) name9203 (
		_w3788_,
		_w9664_,
		_w9665_
	);
	LUT2 #(
		.INIT('h1)
	) name9204 (
		_w9659_,
		_w9665_,
		_w9666_
	);
	LUT2 #(
		.INIT('h2)
	) name9205 (
		_w3411_,
		_w9666_,
		_w9667_
	);
	LUT2 #(
		.INIT('h2)
	) name9206 (
		_w4207_,
		_w4799_,
		_w9668_
	);
	LUT2 #(
		.INIT('h4)
	) name9207 (
		_w4207_,
		_w4799_,
		_w9669_
	);
	LUT2 #(
		.INIT('h1)
	) name9208 (
		_w9668_,
		_w9669_,
		_w9670_
	);
	LUT2 #(
		.INIT('h8)
	) name9209 (
		_w3788_,
		_w9670_,
		_w9671_
	);
	LUT2 #(
		.INIT('h1)
	) name9210 (
		_w9659_,
		_w9671_,
		_w9672_
	);
	LUT2 #(
		.INIT('h1)
	) name9211 (
		_w3177_,
		_w9672_,
		_w9673_
	);
	LUT2 #(
		.INIT('h2)
	) name9212 (
		_w4207_,
		_w4835_,
		_w9674_
	);
	LUT2 #(
		.INIT('h4)
	) name9213 (
		_w4207_,
		_w4835_,
		_w9675_
	);
	LUT2 #(
		.INIT('h1)
	) name9214 (
		_w9674_,
		_w9675_,
		_w9676_
	);
	LUT2 #(
		.INIT('h2)
	) name9215 (
		_w3788_,
		_w9676_,
		_w9677_
	);
	LUT2 #(
		.INIT('h1)
	) name9216 (
		_w9659_,
		_w9677_,
		_w9678_
	);
	LUT2 #(
		.INIT('h1)
	) name9217 (
		_w3320_,
		_w9678_,
		_w9679_
	);
	LUT2 #(
		.INIT('h2)
	) name9218 (
		_w2495_,
		_w3331_,
		_w9680_
	);
	LUT2 #(
		.INIT('h1)
	) name9219 (
		_w3332_,
		_w9680_,
		_w9681_
	);
	LUT2 #(
		.INIT('h8)
	) name9220 (
		_w3355_,
		_w9681_,
		_w9682_
	);
	LUT2 #(
		.INIT('h8)
	) name9221 (
		_w3788_,
		_w9682_,
		_w9683_
	);
	LUT2 #(
		.INIT('h2)
	) name9222 (
		_w2495_,
		_w3965_,
		_w9684_
	);
	LUT2 #(
		.INIT('h1)
	) name9223 (
		_w9658_,
		_w9684_,
		_w9685_
	);
	LUT2 #(
		.INIT('h4)
	) name9224 (
		_w9683_,
		_w9685_,
		_w9686_
	);
	LUT2 #(
		.INIT('h4)
	) name9225 (
		_w9679_,
		_w9686_,
		_w9687_
	);
	LUT2 #(
		.INIT('h4)
	) name9226 (
		_w9673_,
		_w9687_,
		_w9688_
	);
	LUT2 #(
		.INIT('h4)
	) name9227 (
		_w9667_,
		_w9688_,
		_w9689_
	);
	LUT2 #(
		.INIT('h2)
	) name9228 (
		_w2026_,
		_w9689_,
		_w9690_
	);
	LUT2 #(
		.INIT('h1)
	) name9229 (
		_w9657_,
		_w9690_,
		_w9691_
	);
	LUT2 #(
		.INIT('h2)
	) name9230 (
		\P1_state_reg[0]/NET0131 ,
		_w9691_,
		_w9692_
	);
	LUT2 #(
		.INIT('h8)
	) name9231 (
		_w2476_,
		_w3976_,
		_w9693_
	);
	LUT2 #(
		.INIT('h1)
	) name9232 (
		_w9656_,
		_w9693_,
		_w9694_
	);
	LUT2 #(
		.INIT('h4)
	) name9233 (
		_w9692_,
		_w9694_,
		_w9695_
	);
	LUT2 #(
		.INIT('h2)
	) name9234 (
		\P1_reg3_reg[3]/NET0131 ,
		\P1_state_reg[0]/NET0131 ,
		_w9696_
	);
	LUT2 #(
		.INIT('h4)
	) name9235 (
		\P1_reg3_reg[3]/NET0131 ,
		_w3448_,
		_w9697_
	);
	LUT2 #(
		.INIT('h4)
	) name9236 (
		_w1632_,
		_w1880_,
		_w9698_
	);
	LUT2 #(
		.INIT('h1)
	) name9237 (
		_w1632_,
		_w3680_,
		_w9699_
	);
	LUT2 #(
		.INIT('h4)
	) name9238 (
		_w3681_,
		_w3712_,
		_w9700_
	);
	LUT2 #(
		.INIT('h4)
	) name9239 (
		_w9699_,
		_w9700_,
		_w9701_
	);
	LUT2 #(
		.INIT('h1)
	) name9240 (
		_w9698_,
		_w9701_,
		_w9702_
	);
	LUT2 #(
		.INIT('h2)
	) name9241 (
		_w3980_,
		_w9702_,
		_w9703_
	);
	LUT2 #(
		.INIT('h1)
	) name9242 (
		\P1_reg3_reg[3]/NET0131 ,
		_w3980_,
		_w9704_
	);
	LUT2 #(
		.INIT('h2)
	) name9243 (
		_w1572_,
		_w3573_,
		_w9705_
	);
	LUT2 #(
		.INIT('h1)
	) name9244 (
		_w9022_,
		_w9705_,
		_w9706_
	);
	LUT2 #(
		.INIT('h1)
	) name9245 (
		_w537_,
		_w9706_,
		_w9707_
	);
	LUT2 #(
		.INIT('h8)
	) name9246 (
		_w537_,
		_w1595_,
		_w9708_
	);
	LUT2 #(
		.INIT('h1)
	) name9247 (
		_w9707_,
		_w9708_,
		_w9709_
	);
	LUT2 #(
		.INIT('h8)
	) name9248 (
		_w3980_,
		_w9709_,
		_w9710_
	);
	LUT2 #(
		.INIT('h1)
	) name9249 (
		_w9704_,
		_w9710_,
		_w9711_
	);
	LUT2 #(
		.INIT('h2)
	) name9250 (
		_w1936_,
		_w9711_,
		_w9712_
	);
	LUT2 #(
		.INIT('h1)
	) name9251 (
		_w1778_,
		_w3508_,
		_w9713_
	);
	LUT2 #(
		.INIT('h8)
	) name9252 (
		_w1773_,
		_w9713_,
		_w9714_
	);
	LUT2 #(
		.INIT('h1)
	) name9253 (
		_w1773_,
		_w9713_,
		_w9715_
	);
	LUT2 #(
		.INIT('h1)
	) name9254 (
		_w9714_,
		_w9715_,
		_w9716_
	);
	LUT2 #(
		.INIT('h2)
	) name9255 (
		_w3980_,
		_w9716_,
		_w9717_
	);
	LUT2 #(
		.INIT('h1)
	) name9256 (
		_w9704_,
		_w9717_,
		_w9718_
	);
	LUT2 #(
		.INIT('h1)
	) name9257 (
		_w3563_,
		_w9718_,
		_w9719_
	);
	LUT2 #(
		.INIT('h1)
	) name9258 (
		_w1610_,
		_w3633_,
		_w9720_
	);
	LUT2 #(
		.INIT('h8)
	) name9259 (
		_w1773_,
		_w9720_,
		_w9721_
	);
	LUT2 #(
		.INIT('h1)
	) name9260 (
		_w1773_,
		_w9720_,
		_w9722_
	);
	LUT2 #(
		.INIT('h1)
	) name9261 (
		_w9721_,
		_w9722_,
		_w9723_
	);
	LUT2 #(
		.INIT('h8)
	) name9262 (
		_w3980_,
		_w9723_,
		_w9724_
	);
	LUT2 #(
		.INIT('h1)
	) name9263 (
		_w9704_,
		_w9724_,
		_w9725_
	);
	LUT2 #(
		.INIT('h1)
	) name9264 (
		_w3677_,
		_w9725_,
		_w9726_
	);
	LUT2 #(
		.INIT('h4)
	) name9265 (
		_w1632_,
		_w1763_,
		_w9727_
	);
	LUT2 #(
		.INIT('h1)
	) name9266 (
		\P1_reg3_reg[3]/NET0131 ,
		_w9092_,
		_w9728_
	);
	LUT2 #(
		.INIT('h1)
	) name9267 (
		_w9727_,
		_w9728_,
		_w9729_
	);
	LUT2 #(
		.INIT('h4)
	) name9268 (
		_w9703_,
		_w9729_,
		_w9730_
	);
	LUT2 #(
		.INIT('h4)
	) name9269 (
		_w9726_,
		_w9730_,
		_w9731_
	);
	LUT2 #(
		.INIT('h4)
	) name9270 (
		_w9719_,
		_w9731_,
		_w9732_
	);
	LUT2 #(
		.INIT('h4)
	) name9271 (
		_w9712_,
		_w9732_,
		_w9733_
	);
	LUT2 #(
		.INIT('h2)
	) name9272 (
		_w3450_,
		_w9733_,
		_w9734_
	);
	LUT2 #(
		.INIT('h1)
	) name9273 (
		_w9697_,
		_w9734_,
		_w9735_
	);
	LUT2 #(
		.INIT('h2)
	) name9274 (
		\P1_state_reg[0]/NET0131 ,
		_w9735_,
		_w9736_
	);
	LUT2 #(
		.INIT('h4)
	) name9275 (
		\P1_reg3_reg[3]/NET0131 ,
		_w1953_,
		_w9737_
	);
	LUT2 #(
		.INIT('h1)
	) name9276 (
		_w9696_,
		_w9737_,
		_w9738_
	);
	LUT2 #(
		.INIT('h4)
	) name9277 (
		_w9736_,
		_w9738_,
		_w9739_
	);
	LUT2 #(
		.INIT('h2)
	) name9278 (
		\P1_reg3_reg[6]/NET0131 ,
		\P1_state_reg[0]/NET0131 ,
		_w9740_
	);
	LUT2 #(
		.INIT('h8)
	) name9279 (
		_w1518_,
		_w1953_,
		_w9741_
	);
	LUT2 #(
		.INIT('h8)
	) name9280 (
		_w1518_,
		_w3448_,
		_w9742_
	);
	LUT2 #(
		.INIT('h1)
	) name9281 (
		_w1537_,
		_w4067_,
		_w9743_
	);
	LUT2 #(
		.INIT('h2)
	) name9282 (
		_w1518_,
		_w3980_,
		_w9744_
	);
	LUT2 #(
		.INIT('h2)
	) name9283 (
		_w537_,
		_w1548_,
		_w9745_
	);
	LUT2 #(
		.INIT('h2)
	) name9284 (
		_w1498_,
		_w9069_,
		_w9746_
	);
	LUT2 #(
		.INIT('h1)
	) name9285 (
		_w537_,
		_w3577_,
		_w9747_
	);
	LUT2 #(
		.INIT('h4)
	) name9286 (
		_w9746_,
		_w9747_,
		_w9748_
	);
	LUT2 #(
		.INIT('h1)
	) name9287 (
		_w9745_,
		_w9748_,
		_w9749_
	);
	LUT2 #(
		.INIT('h2)
	) name9288 (
		_w3980_,
		_w9749_,
		_w9750_
	);
	LUT2 #(
		.INIT('h1)
	) name9289 (
		_w9744_,
		_w9750_,
		_w9751_
	);
	LUT2 #(
		.INIT('h2)
	) name9290 (
		_w1936_,
		_w9751_,
		_w9752_
	);
	LUT2 #(
		.INIT('h4)
	) name9291 (
		_w1686_,
		_w1793_,
		_w9753_
	);
	LUT2 #(
		.INIT('h2)
	) name9292 (
		_w1686_,
		_w1793_,
		_w9754_
	);
	LUT2 #(
		.INIT('h1)
	) name9293 (
		_w9753_,
		_w9754_,
		_w9755_
	);
	LUT2 #(
		.INIT('h8)
	) name9294 (
		_w3980_,
		_w9755_,
		_w9756_
	);
	LUT2 #(
		.INIT('h1)
	) name9295 (
		_w9744_,
		_w9756_,
		_w9757_
	);
	LUT2 #(
		.INIT('h1)
	) name9296 (
		_w3677_,
		_w9757_,
		_w9758_
	);
	LUT2 #(
		.INIT('h2)
	) name9297 (
		_w1793_,
		_w5509_,
		_w9759_
	);
	LUT2 #(
		.INIT('h4)
	) name9298 (
		_w1793_,
		_w5509_,
		_w9760_
	);
	LUT2 #(
		.INIT('h1)
	) name9299 (
		_w9759_,
		_w9760_,
		_w9761_
	);
	LUT2 #(
		.INIT('h2)
	) name9300 (
		_w3980_,
		_w9761_,
		_w9762_
	);
	LUT2 #(
		.INIT('h1)
	) name9301 (
		_w9744_,
		_w9762_,
		_w9763_
	);
	LUT2 #(
		.INIT('h1)
	) name9302 (
		_w3563_,
		_w9763_,
		_w9764_
	);
	LUT2 #(
		.INIT('h1)
	) name9303 (
		_w1537_,
		_w3683_,
		_w9765_
	);
	LUT2 #(
		.INIT('h1)
	) name9304 (
		_w3684_,
		_w9765_,
		_w9766_
	);
	LUT2 #(
		.INIT('h8)
	) name9305 (
		_w3980_,
		_w9766_,
		_w9767_
	);
	LUT2 #(
		.INIT('h1)
	) name9306 (
		_w9744_,
		_w9767_,
		_w9768_
	);
	LUT2 #(
		.INIT('h2)
	) name9307 (
		_w3712_,
		_w9768_,
		_w9769_
	);
	LUT2 #(
		.INIT('h2)
	) name9308 (
		_w1518_,
		_w4064_,
		_w9770_
	);
	LUT2 #(
		.INIT('h1)
	) name9309 (
		_w9743_,
		_w9770_,
		_w9771_
	);
	LUT2 #(
		.INIT('h4)
	) name9310 (
		_w9769_,
		_w9771_,
		_w9772_
	);
	LUT2 #(
		.INIT('h4)
	) name9311 (
		_w9752_,
		_w9772_,
		_w9773_
	);
	LUT2 #(
		.INIT('h1)
	) name9312 (
		_w9758_,
		_w9764_,
		_w9774_
	);
	LUT2 #(
		.INIT('h8)
	) name9313 (
		_w9773_,
		_w9774_,
		_w9775_
	);
	LUT2 #(
		.INIT('h2)
	) name9314 (
		_w3450_,
		_w9775_,
		_w9776_
	);
	LUT2 #(
		.INIT('h1)
	) name9315 (
		_w9742_,
		_w9776_,
		_w9777_
	);
	LUT2 #(
		.INIT('h2)
	) name9316 (
		\P1_state_reg[0]/NET0131 ,
		_w9777_,
		_w9778_
	);
	LUT2 #(
		.INIT('h1)
	) name9317 (
		_w9740_,
		_w9741_,
		_w9779_
	);
	LUT2 #(
		.INIT('h4)
	) name9318 (
		_w9778_,
		_w9779_,
		_w9780_
	);
	LUT2 #(
		.INIT('h2)
	) name9319 (
		\P1_reg3_reg[7]/NET0131 ,
		\P1_state_reg[0]/NET0131 ,
		_w9781_
	);
	LUT2 #(
		.INIT('h8)
	) name9320 (
		_w1491_,
		_w1953_,
		_w9782_
	);
	LUT2 #(
		.INIT('h8)
	) name9321 (
		_w1491_,
		_w3448_,
		_w9783_
	);
	LUT2 #(
		.INIT('h2)
	) name9322 (
		_w1491_,
		_w4910_,
		_w9784_
	);
	LUT2 #(
		.INIT('h2)
	) name9323 (
		_w1491_,
		_w3980_,
		_w9785_
	);
	LUT2 #(
		.INIT('h2)
	) name9324 (
		_w1776_,
		_w4399_,
		_w9786_
	);
	LUT2 #(
		.INIT('h4)
	) name9325 (
		_w1776_,
		_w4399_,
		_w9787_
	);
	LUT2 #(
		.INIT('h1)
	) name9326 (
		_w9786_,
		_w9787_,
		_w9788_
	);
	LUT2 #(
		.INIT('h2)
	) name9327 (
		_w3980_,
		_w9788_,
		_w9789_
	);
	LUT2 #(
		.INIT('h1)
	) name9328 (
		_w9785_,
		_w9789_,
		_w9790_
	);
	LUT2 #(
		.INIT('h1)
	) name9329 (
		_w3677_,
		_w9790_,
		_w9791_
	);
	LUT2 #(
		.INIT('h2)
	) name9330 (
		_w1776_,
		_w4442_,
		_w9792_
	);
	LUT2 #(
		.INIT('h4)
	) name9331 (
		_w1776_,
		_w4442_,
		_w9793_
	);
	LUT2 #(
		.INIT('h1)
	) name9332 (
		_w9792_,
		_w9793_,
		_w9794_
	);
	LUT2 #(
		.INIT('h8)
	) name9333 (
		_w3980_,
		_w9794_,
		_w9795_
	);
	LUT2 #(
		.INIT('h1)
	) name9334 (
		_w9785_,
		_w9795_,
		_w9796_
	);
	LUT2 #(
		.INIT('h1)
	) name9335 (
		_w3563_,
		_w9796_,
		_w9797_
	);
	LUT2 #(
		.INIT('h2)
	) name9336 (
		_w1267_,
		_w3577_,
		_w9798_
	);
	LUT2 #(
		.INIT('h1)
	) name9337 (
		_w7305_,
		_w9798_,
		_w9799_
	);
	LUT2 #(
		.INIT('h1)
	) name9338 (
		_w537_,
		_w9799_,
		_w9800_
	);
	LUT2 #(
		.INIT('h8)
	) name9339 (
		_w537_,
		_w1524_,
		_w9801_
	);
	LUT2 #(
		.INIT('h1)
	) name9340 (
		_w9800_,
		_w9801_,
		_w9802_
	);
	LUT2 #(
		.INIT('h8)
	) name9341 (
		_w3980_,
		_w9802_,
		_w9803_
	);
	LUT2 #(
		.INIT('h1)
	) name9342 (
		_w9785_,
		_w9803_,
		_w9804_
	);
	LUT2 #(
		.INIT('h2)
	) name9343 (
		_w1936_,
		_w9804_,
		_w9805_
	);
	LUT2 #(
		.INIT('h1)
	) name9344 (
		_w1514_,
		_w3684_,
		_w9806_
	);
	LUT2 #(
		.INIT('h1)
	) name9345 (
		_w8308_,
		_w9806_,
		_w9807_
	);
	LUT2 #(
		.INIT('h8)
	) name9346 (
		_w3712_,
		_w9807_,
		_w9808_
	);
	LUT2 #(
		.INIT('h8)
	) name9347 (
		_w3980_,
		_w9808_,
		_w9809_
	);
	LUT2 #(
		.INIT('h1)
	) name9348 (
		_w1514_,
		_w4067_,
		_w9810_
	);
	LUT2 #(
		.INIT('h1)
	) name9349 (
		_w9784_,
		_w9810_,
		_w9811_
	);
	LUT2 #(
		.INIT('h4)
	) name9350 (
		_w9809_,
		_w9811_,
		_w9812_
	);
	LUT2 #(
		.INIT('h4)
	) name9351 (
		_w9791_,
		_w9812_,
		_w9813_
	);
	LUT2 #(
		.INIT('h1)
	) name9352 (
		_w9797_,
		_w9805_,
		_w9814_
	);
	LUT2 #(
		.INIT('h8)
	) name9353 (
		_w9813_,
		_w9814_,
		_w9815_
	);
	LUT2 #(
		.INIT('h2)
	) name9354 (
		_w3450_,
		_w9815_,
		_w9816_
	);
	LUT2 #(
		.INIT('h1)
	) name9355 (
		_w9783_,
		_w9816_,
		_w9817_
	);
	LUT2 #(
		.INIT('h2)
	) name9356 (
		\P1_state_reg[0]/NET0131 ,
		_w9817_,
		_w9818_
	);
	LUT2 #(
		.INIT('h1)
	) name9357 (
		_w9781_,
		_w9782_,
		_w9819_
	);
	LUT2 #(
		.INIT('h4)
	) name9358 (
		_w9818_,
		_w9819_,
		_w9820_
	);
	LUT2 #(
		.INIT('h2)
	) name9359 (
		\P1_reg1_reg[5]/NET0131 ,
		_w3435_,
		_w9821_
	);
	LUT2 #(
		.INIT('h8)
	) name9360 (
		\P1_reg1_reg[5]/NET0131 ,
		_w3448_,
		_w9822_
	);
	LUT2 #(
		.INIT('h2)
	) name9361 (
		_w4532_,
		_w9065_,
		_w9823_
	);
	LUT2 #(
		.INIT('h2)
	) name9362 (
		\P1_reg1_reg[5]/NET0131 ,
		_w4532_,
		_w9824_
	);
	LUT2 #(
		.INIT('h8)
	) name9363 (
		_w4532_,
		_w9073_,
		_w9825_
	);
	LUT2 #(
		.INIT('h1)
	) name9364 (
		_w9824_,
		_w9825_,
		_w9826_
	);
	LUT2 #(
		.INIT('h2)
	) name9365 (
		_w1936_,
		_w9826_,
		_w9827_
	);
	LUT2 #(
		.INIT('h2)
	) name9366 (
		_w4532_,
		_w9079_,
		_w9828_
	);
	LUT2 #(
		.INIT('h1)
	) name9367 (
		_w9824_,
		_w9828_,
		_w9829_
	);
	LUT2 #(
		.INIT('h1)
	) name9368 (
		_w3563_,
		_w9829_,
		_w9830_
	);
	LUT2 #(
		.INIT('h2)
	) name9369 (
		_w4532_,
		_w9085_,
		_w9831_
	);
	LUT2 #(
		.INIT('h1)
	) name9370 (
		_w9824_,
		_w9831_,
		_w9832_
	);
	LUT2 #(
		.INIT('h1)
	) name9371 (
		_w3677_,
		_w9832_,
		_w9833_
	);
	LUT2 #(
		.INIT('h4)
	) name9372 (
		_w4532_,
		_w9090_,
		_w9834_
	);
	LUT2 #(
		.INIT('h2)
	) name9373 (
		_w4491_,
		_w9834_,
		_w9835_
	);
	LUT2 #(
		.INIT('h2)
	) name9374 (
		\P1_reg1_reg[5]/NET0131 ,
		_w9835_,
		_w9836_
	);
	LUT2 #(
		.INIT('h1)
	) name9375 (
		_w9823_,
		_w9836_,
		_w9837_
	);
	LUT2 #(
		.INIT('h4)
	) name9376 (
		_w9830_,
		_w9837_,
		_w9838_
	);
	LUT2 #(
		.INIT('h4)
	) name9377 (
		_w9833_,
		_w9838_,
		_w9839_
	);
	LUT2 #(
		.INIT('h4)
	) name9378 (
		_w9827_,
		_w9839_,
		_w9840_
	);
	LUT2 #(
		.INIT('h2)
	) name9379 (
		_w3450_,
		_w9840_,
		_w9841_
	);
	LUT2 #(
		.INIT('h1)
	) name9380 (
		_w9822_,
		_w9841_,
		_w9842_
	);
	LUT2 #(
		.INIT('h2)
	) name9381 (
		\P1_state_reg[0]/NET0131 ,
		_w9842_,
		_w9843_
	);
	LUT2 #(
		.INIT('h1)
	) name9382 (
		_w9821_,
		_w9843_,
		_w9844_
	);
	LUT2 #(
		.INIT('h8)
	) name9383 (
		_w3411_,
		_w8985_,
		_w9845_
	);
	LUT2 #(
		.INIT('h2)
	) name9384 (
		_w9353_,
		_w9845_,
		_w9846_
	);
	LUT2 #(
		.INIT('h2)
	) name9385 (
		\P2_reg0_reg[5]/NET0131 ,
		_w9846_,
		_w9847_
	);
	LUT2 #(
		.INIT('h4)
	) name9386 (
		_w2544_,
		_w3358_,
		_w9848_
	);
	LUT2 #(
		.INIT('h1)
	) name9387 (
		_w3177_,
		_w8991_,
		_w9849_
	);
	LUT2 #(
		.INIT('h2)
	) name9388 (
		_w9002_,
		_w9848_,
		_w9850_
	);
	LUT2 #(
		.INIT('h4)
	) name9389 (
		_w9849_,
		_w9850_,
		_w9851_
	);
	LUT2 #(
		.INIT('h4)
	) name9390 (
		_w9845_,
		_w9851_,
		_w9852_
	);
	LUT2 #(
		.INIT('h2)
	) name9391 (
		_w5860_,
		_w9852_,
		_w9853_
	);
	LUT2 #(
		.INIT('h1)
	) name9392 (
		_w9847_,
		_w9853_,
		_w9854_
	);
	LUT2 #(
		.INIT('h2)
	) name9393 (
		\P2_reg1_reg[11]/NET0131 ,
		_w1983_,
		_w9855_
	);
	LUT2 #(
		.INIT('h8)
	) name9394 (
		\P2_reg1_reg[11]/NET0131 ,
		_w2024_,
		_w9856_
	);
	LUT2 #(
		.INIT('h2)
	) name9395 (
		\P2_reg1_reg[11]/NET0131 ,
		_w8532_,
		_w9857_
	);
	LUT2 #(
		.INIT('h2)
	) name9396 (
		\P2_reg1_reg[11]/NET0131 ,
		_w3733_,
		_w9858_
	);
	LUT2 #(
		.INIT('h8)
	) name9397 (
		_w3733_,
		_w8129_,
		_w9859_
	);
	LUT2 #(
		.INIT('h1)
	) name9398 (
		_w9858_,
		_w9859_,
		_w9860_
	);
	LUT2 #(
		.INIT('h2)
	) name9399 (
		_w3411_,
		_w9860_,
		_w9861_
	);
	LUT2 #(
		.INIT('h8)
	) name9400 (
		_w3733_,
		_w8135_,
		_w9862_
	);
	LUT2 #(
		.INIT('h1)
	) name9401 (
		_w9858_,
		_w9862_,
		_w9863_
	);
	LUT2 #(
		.INIT('h1)
	) name9402 (
		_w3177_,
		_w9863_,
		_w9864_
	);
	LUT2 #(
		.INIT('h8)
	) name9403 (
		_w3355_,
		_w8140_,
		_w9865_
	);
	LUT2 #(
		.INIT('h1)
	) name9404 (
		_w8147_,
		_w9408_,
		_w9866_
	);
	LUT2 #(
		.INIT('h4)
	) name9405 (
		_w9865_,
		_w9866_,
		_w9867_
	);
	LUT2 #(
		.INIT('h2)
	) name9406 (
		_w3733_,
		_w9867_,
		_w9868_
	);
	LUT2 #(
		.INIT('h1)
	) name9407 (
		_w9857_,
		_w9868_,
		_w9869_
	);
	LUT2 #(
		.INIT('h4)
	) name9408 (
		_w9864_,
		_w9869_,
		_w9870_
	);
	LUT2 #(
		.INIT('h4)
	) name9409 (
		_w9861_,
		_w9870_,
		_w9871_
	);
	LUT2 #(
		.INIT('h2)
	) name9410 (
		_w2026_,
		_w9871_,
		_w9872_
	);
	LUT2 #(
		.INIT('h1)
	) name9411 (
		_w9856_,
		_w9872_,
		_w9873_
	);
	LUT2 #(
		.INIT('h2)
	) name9412 (
		\P1_state_reg[0]/NET0131 ,
		_w9873_,
		_w9874_
	);
	LUT2 #(
		.INIT('h1)
	) name9413 (
		_w9855_,
		_w9874_,
		_w9875_
	);
	LUT2 #(
		.INIT('h2)
	) name9414 (
		\P2_reg1_reg[14]/NET0131 ,
		_w1983_,
		_w9876_
	);
	LUT2 #(
		.INIT('h8)
	) name9415 (
		\P2_reg1_reg[14]/NET0131 ,
		_w2024_,
		_w9877_
	);
	LUT2 #(
		.INIT('h8)
	) name9416 (
		_w3733_,
		_w9437_,
		_w9878_
	);
	LUT2 #(
		.INIT('h2)
	) name9417 (
		\P2_reg1_reg[14]/NET0131 ,
		_w3743_,
		_w9879_
	);
	LUT2 #(
		.INIT('h2)
	) name9418 (
		\P2_reg1_reg[14]/NET0131 ,
		_w3733_,
		_w9880_
	);
	LUT2 #(
		.INIT('h8)
	) name9419 (
		_w3733_,
		_w8176_,
		_w9881_
	);
	LUT2 #(
		.INIT('h1)
	) name9420 (
		_w9880_,
		_w9881_,
		_w9882_
	);
	LUT2 #(
		.INIT('h2)
	) name9421 (
		_w3355_,
		_w9882_,
		_w9883_
	);
	LUT2 #(
		.INIT('h8)
	) name9422 (
		_w3733_,
		_w8182_,
		_w9884_
	);
	LUT2 #(
		.INIT('h1)
	) name9423 (
		_w9880_,
		_w9884_,
		_w9885_
	);
	LUT2 #(
		.INIT('h1)
	) name9424 (
		_w3177_,
		_w9885_,
		_w9886_
	);
	LUT2 #(
		.INIT('h2)
	) name9425 (
		_w3733_,
		_w8188_,
		_w9887_
	);
	LUT2 #(
		.INIT('h1)
	) name9426 (
		_w9880_,
		_w9887_,
		_w9888_
	);
	LUT2 #(
		.INIT('h1)
	) name9427 (
		_w3320_,
		_w9888_,
		_w9889_
	);
	LUT2 #(
		.INIT('h8)
	) name9428 (
		_w3733_,
		_w8171_,
		_w9890_
	);
	LUT2 #(
		.INIT('h1)
	) name9429 (
		_w9880_,
		_w9890_,
		_w9891_
	);
	LUT2 #(
		.INIT('h2)
	) name9430 (
		_w3411_,
		_w9891_,
		_w9892_
	);
	LUT2 #(
		.INIT('h1)
	) name9431 (
		_w9878_,
		_w9879_,
		_w9893_
	);
	LUT2 #(
		.INIT('h4)
	) name9432 (
		_w9883_,
		_w9893_,
		_w9894_
	);
	LUT2 #(
		.INIT('h1)
	) name9433 (
		_w9886_,
		_w9889_,
		_w9895_
	);
	LUT2 #(
		.INIT('h4)
	) name9434 (
		_w9892_,
		_w9895_,
		_w9896_
	);
	LUT2 #(
		.INIT('h8)
	) name9435 (
		_w9894_,
		_w9896_,
		_w9897_
	);
	LUT2 #(
		.INIT('h2)
	) name9436 (
		_w2026_,
		_w9897_,
		_w9898_
	);
	LUT2 #(
		.INIT('h1)
	) name9437 (
		_w9877_,
		_w9898_,
		_w9899_
	);
	LUT2 #(
		.INIT('h2)
	) name9438 (
		\P1_state_reg[0]/NET0131 ,
		_w9899_,
		_w9900_
	);
	LUT2 #(
		.INIT('h1)
	) name9439 (
		_w9876_,
		_w9900_,
		_w9901_
	);
	LUT2 #(
		.INIT('h2)
	) name9440 (
		_w5964_,
		_w9852_,
		_w9902_
	);
	LUT2 #(
		.INIT('h2)
	) name9441 (
		_w3357_,
		_w3418_,
		_w9903_
	);
	LUT2 #(
		.INIT('h2)
	) name9442 (
		_w3320_,
		_w9903_,
		_w9904_
	);
	LUT2 #(
		.INIT('h1)
	) name9443 (
		_w3733_,
		_w9904_,
		_w9905_
	);
	LUT2 #(
		.INIT('h2)
	) name9444 (
		_w3421_,
		_w9905_,
		_w9906_
	);
	LUT2 #(
		.INIT('h2)
	) name9445 (
		_w5287_,
		_w8533_,
		_w9907_
	);
	LUT2 #(
		.INIT('h8)
	) name9446 (
		_w9906_,
		_w9907_,
		_w9908_
	);
	LUT2 #(
		.INIT('h2)
	) name9447 (
		\P2_reg1_reg[5]/NET0131 ,
		_w9908_,
		_w9909_
	);
	LUT2 #(
		.INIT('h1)
	) name9448 (
		_w9902_,
		_w9909_,
		_w9910_
	);
	LUT2 #(
		.INIT('h2)
	) name9449 (
		\P1_reg2_reg[4]/NET0131 ,
		_w3435_,
		_w9911_
	);
	LUT2 #(
		.INIT('h8)
	) name9450 (
		\P1_reg2_reg[4]/NET0131 ,
		_w3448_,
		_w9912_
	);
	LUT2 #(
		.INIT('h8)
	) name9451 (
		_w3466_,
		_w9106_,
		_w9913_
	);
	LUT2 #(
		.INIT('h2)
	) name9452 (
		\P1_reg2_reg[4]/NET0131 ,
		_w3466_,
		_w9914_
	);
	LUT2 #(
		.INIT('h2)
	) name9453 (
		_w3466_,
		_w9026_,
		_w9915_
	);
	LUT2 #(
		.INIT('h1)
	) name9454 (
		_w9914_,
		_w9915_,
		_w9916_
	);
	LUT2 #(
		.INIT('h2)
	) name9455 (
		_w1936_,
		_w9916_,
		_w9917_
	);
	LUT2 #(
		.INIT('h2)
	) name9456 (
		_w3466_,
		_w9032_,
		_w9918_
	);
	LUT2 #(
		.INIT('h1)
	) name9457 (
		_w9914_,
		_w9918_,
		_w9919_
	);
	LUT2 #(
		.INIT('h1)
	) name9458 (
		_w3563_,
		_w9919_,
		_w9920_
	);
	LUT2 #(
		.INIT('h8)
	) name9459 (
		_w3466_,
		_w9038_,
		_w9921_
	);
	LUT2 #(
		.INIT('h1)
	) name9460 (
		_w9914_,
		_w9921_,
		_w9922_
	);
	LUT2 #(
		.INIT('h1)
	) name9461 (
		_w3677_,
		_w9922_,
		_w9923_
	);
	LUT2 #(
		.INIT('h8)
	) name9462 (
		_w3466_,
		_w9043_,
		_w9924_
	);
	LUT2 #(
		.INIT('h1)
	) name9463 (
		_w9914_,
		_w9924_,
		_w9925_
	);
	LUT2 #(
		.INIT('h2)
	) name9464 (
		_w3712_,
		_w9925_,
		_w9926_
	);
	LUT2 #(
		.INIT('h8)
	) name9465 (
		_w1568_,
		_w1763_,
		_w9927_
	);
	LUT2 #(
		.INIT('h2)
	) name9466 (
		\P1_reg2_reg[4]/NET0131 ,
		_w3718_,
		_w9928_
	);
	LUT2 #(
		.INIT('h1)
	) name9467 (
		_w9913_,
		_w9927_,
		_w9929_
	);
	LUT2 #(
		.INIT('h4)
	) name9468 (
		_w9928_,
		_w9929_,
		_w9930_
	);
	LUT2 #(
		.INIT('h4)
	) name9469 (
		_w9926_,
		_w9930_,
		_w9931_
	);
	LUT2 #(
		.INIT('h4)
	) name9470 (
		_w9920_,
		_w9931_,
		_w9932_
	);
	LUT2 #(
		.INIT('h4)
	) name9471 (
		_w9923_,
		_w9932_,
		_w9933_
	);
	LUT2 #(
		.INIT('h4)
	) name9472 (
		_w9917_,
		_w9933_,
		_w9934_
	);
	LUT2 #(
		.INIT('h2)
	) name9473 (
		_w3450_,
		_w9934_,
		_w9935_
	);
	LUT2 #(
		.INIT('h1)
	) name9474 (
		_w9912_,
		_w9935_,
		_w9936_
	);
	LUT2 #(
		.INIT('h2)
	) name9475 (
		\P1_state_reg[0]/NET0131 ,
		_w9936_,
		_w9937_
	);
	LUT2 #(
		.INIT('h1)
	) name9476 (
		_w9911_,
		_w9937_,
		_w9938_
	);
	LUT2 #(
		.INIT('h2)
	) name9477 (
		\P1_reg2_reg[5]/NET0131 ,
		_w3435_,
		_w9939_
	);
	LUT2 #(
		.INIT('h8)
	) name9478 (
		\P1_reg2_reg[5]/NET0131 ,
		_w3448_,
		_w9940_
	);
	LUT2 #(
		.INIT('h2)
	) name9479 (
		_w3466_,
		_w9065_,
		_w9941_
	);
	LUT2 #(
		.INIT('h2)
	) name9480 (
		\P1_reg2_reg[5]/NET0131 ,
		_w3466_,
		_w9942_
	);
	LUT2 #(
		.INIT('h8)
	) name9481 (
		_w3466_,
		_w9073_,
		_w9943_
	);
	LUT2 #(
		.INIT('h1)
	) name9482 (
		_w9942_,
		_w9943_,
		_w9944_
	);
	LUT2 #(
		.INIT('h2)
	) name9483 (
		_w1936_,
		_w9944_,
		_w9945_
	);
	LUT2 #(
		.INIT('h2)
	) name9484 (
		_w3466_,
		_w9079_,
		_w9946_
	);
	LUT2 #(
		.INIT('h1)
	) name9485 (
		_w9942_,
		_w9946_,
		_w9947_
	);
	LUT2 #(
		.INIT('h1)
	) name9486 (
		_w3563_,
		_w9947_,
		_w9948_
	);
	LUT2 #(
		.INIT('h2)
	) name9487 (
		_w3466_,
		_w9085_,
		_w9949_
	);
	LUT2 #(
		.INIT('h1)
	) name9488 (
		_w9942_,
		_w9949_,
		_w9950_
	);
	LUT2 #(
		.INIT('h1)
	) name9489 (
		_w3677_,
		_w9950_,
		_w9951_
	);
	LUT2 #(
		.INIT('h8)
	) name9490 (
		_w1543_,
		_w1763_,
		_w9952_
	);
	LUT2 #(
		.INIT('h4)
	) name9491 (
		_w3466_,
		_w9090_,
		_w9953_
	);
	LUT2 #(
		.INIT('h1)
	) name9492 (
		_w3716_,
		_w9953_,
		_w9954_
	);
	LUT2 #(
		.INIT('h2)
	) name9493 (
		\P1_reg2_reg[5]/NET0131 ,
		_w9954_,
		_w9955_
	);
	LUT2 #(
		.INIT('h1)
	) name9494 (
		_w9952_,
		_w9955_,
		_w9956_
	);
	LUT2 #(
		.INIT('h4)
	) name9495 (
		_w9941_,
		_w9956_,
		_w9957_
	);
	LUT2 #(
		.INIT('h4)
	) name9496 (
		_w9948_,
		_w9957_,
		_w9958_
	);
	LUT2 #(
		.INIT('h4)
	) name9497 (
		_w9951_,
		_w9958_,
		_w9959_
	);
	LUT2 #(
		.INIT('h4)
	) name9498 (
		_w9945_,
		_w9959_,
		_w9960_
	);
	LUT2 #(
		.INIT('h2)
	) name9499 (
		_w3450_,
		_w9960_,
		_w9961_
	);
	LUT2 #(
		.INIT('h1)
	) name9500 (
		_w9940_,
		_w9961_,
		_w9962_
	);
	LUT2 #(
		.INIT('h2)
	) name9501 (
		\P1_state_reg[0]/NET0131 ,
		_w9962_,
		_w9963_
	);
	LUT2 #(
		.INIT('h1)
	) name9502 (
		_w9939_,
		_w9963_,
		_w9964_
	);
	LUT2 #(
		.INIT('h2)
	) name9503 (
		\P1_reg0_reg[11]/NET0131 ,
		_w3435_,
		_w9965_
	);
	LUT2 #(
		.INIT('h8)
	) name9504 (
		\P1_reg0_reg[11]/NET0131 ,
		_w3448_,
		_w9966_
	);
	LUT2 #(
		.INIT('h2)
	) name9505 (
		\P1_reg0_reg[11]/NET0131 ,
		_w4494_,
		_w9967_
	);
	LUT2 #(
		.INIT('h2)
	) name9506 (
		\P1_reg0_reg[11]/NET0131 ,
		_w4396_,
		_w9968_
	);
	LUT2 #(
		.INIT('h8)
	) name9507 (
		_w4396_,
		_w8010_,
		_w9969_
	);
	LUT2 #(
		.INIT('h1)
	) name9508 (
		_w9968_,
		_w9969_,
		_w9970_
	);
	LUT2 #(
		.INIT('h1)
	) name9509 (
		_w3563_,
		_w9970_,
		_w9971_
	);
	LUT2 #(
		.INIT('h8)
	) name9510 (
		_w4396_,
		_w8018_,
		_w9972_
	);
	LUT2 #(
		.INIT('h1)
	) name9511 (
		_w9968_,
		_w9972_,
		_w9973_
	);
	LUT2 #(
		.INIT('h2)
	) name9512 (
		_w1936_,
		_w9973_,
		_w9974_
	);
	LUT2 #(
		.INIT('h2)
	) name9513 (
		_w4396_,
		_w8004_,
		_w9975_
	);
	LUT2 #(
		.INIT('h1)
	) name9514 (
		_w9968_,
		_w9975_,
		_w9976_
	);
	LUT2 #(
		.INIT('h1)
	) name9515 (
		_w3677_,
		_w9976_,
		_w9977_
	);
	LUT2 #(
		.INIT('h2)
	) name9516 (
		_w4396_,
		_w9279_,
		_w9978_
	);
	LUT2 #(
		.INIT('h1)
	) name9517 (
		_w9967_,
		_w9978_,
		_w9979_
	);
	LUT2 #(
		.INIT('h4)
	) name9518 (
		_w9971_,
		_w9979_,
		_w9980_
	);
	LUT2 #(
		.INIT('h1)
	) name9519 (
		_w9974_,
		_w9977_,
		_w9981_
	);
	LUT2 #(
		.INIT('h8)
	) name9520 (
		_w9980_,
		_w9981_,
		_w9982_
	);
	LUT2 #(
		.INIT('h2)
	) name9521 (
		_w3450_,
		_w9982_,
		_w9983_
	);
	LUT2 #(
		.INIT('h1)
	) name9522 (
		_w9966_,
		_w9983_,
		_w9984_
	);
	LUT2 #(
		.INIT('h2)
	) name9523 (
		\P1_state_reg[0]/NET0131 ,
		_w9984_,
		_w9985_
	);
	LUT2 #(
		.INIT('h1)
	) name9524 (
		_w9965_,
		_w9985_,
		_w9986_
	);
	LUT2 #(
		.INIT('h2)
	) name9525 (
		\P2_reg2_reg[4]/NET0131 ,
		_w1983_,
		_w9987_
	);
	LUT2 #(
		.INIT('h8)
	) name9526 (
		\P2_reg2_reg[4]/NET0131 ,
		_w2024_,
		_w9988_
	);
	LUT2 #(
		.INIT('h8)
	) name9527 (
		_w3758_,
		_w9159_,
		_w9989_
	);
	LUT2 #(
		.INIT('h2)
	) name9528 (
		\P2_reg2_reg[4]/NET0131 ,
		_w3758_,
		_w9990_
	);
	LUT2 #(
		.INIT('h2)
	) name9529 (
		_w3758_,
		_w8945_,
		_w9991_
	);
	LUT2 #(
		.INIT('h1)
	) name9530 (
		_w9990_,
		_w9991_,
		_w9992_
	);
	LUT2 #(
		.INIT('h2)
	) name9531 (
		_w3411_,
		_w9992_,
		_w9993_
	);
	LUT2 #(
		.INIT('h8)
	) name9532 (
		_w3758_,
		_w8951_,
		_w9994_
	);
	LUT2 #(
		.INIT('h1)
	) name9533 (
		_w9990_,
		_w9994_,
		_w9995_
	);
	LUT2 #(
		.INIT('h1)
	) name9534 (
		_w3177_,
		_w9995_,
		_w9996_
	);
	LUT2 #(
		.INIT('h2)
	) name9535 (
		_w3758_,
		_w8957_,
		_w9997_
	);
	LUT2 #(
		.INIT('h1)
	) name9536 (
		_w9990_,
		_w9997_,
		_w9998_
	);
	LUT2 #(
		.INIT('h1)
	) name9537 (
		_w3320_,
		_w9998_,
		_w9999_
	);
	LUT2 #(
		.INIT('h8)
	) name9538 (
		_w3758_,
		_w8962_,
		_w10000_
	);
	LUT2 #(
		.INIT('h1)
	) name9539 (
		_w9990_,
		_w10000_,
		_w10001_
	);
	LUT2 #(
		.INIT('h2)
	) name9540 (
		_w3355_,
		_w10001_,
		_w10002_
	);
	LUT2 #(
		.INIT('h8)
	) name9541 (
		_w2635_,
		_w3420_,
		_w10003_
	);
	LUT2 #(
		.INIT('h2)
	) name9542 (
		\P2_reg2_reg[4]/NET0131 ,
		_w3774_,
		_w10004_
	);
	LUT2 #(
		.INIT('h1)
	) name9543 (
		_w9989_,
		_w10003_,
		_w10005_
	);
	LUT2 #(
		.INIT('h4)
	) name9544 (
		_w10004_,
		_w10005_,
		_w10006_
	);
	LUT2 #(
		.INIT('h4)
	) name9545 (
		_w10002_,
		_w10006_,
		_w10007_
	);
	LUT2 #(
		.INIT('h4)
	) name9546 (
		_w9996_,
		_w10007_,
		_w10008_
	);
	LUT2 #(
		.INIT('h4)
	) name9547 (
		_w9999_,
		_w10008_,
		_w10009_
	);
	LUT2 #(
		.INIT('h4)
	) name9548 (
		_w9993_,
		_w10009_,
		_w10010_
	);
	LUT2 #(
		.INIT('h2)
	) name9549 (
		_w2026_,
		_w10010_,
		_w10011_
	);
	LUT2 #(
		.INIT('h1)
	) name9550 (
		_w9988_,
		_w10011_,
		_w10012_
	);
	LUT2 #(
		.INIT('h2)
	) name9551 (
		\P1_state_reg[0]/NET0131 ,
		_w10012_,
		_w10013_
	);
	LUT2 #(
		.INIT('h1)
	) name9552 (
		_w9987_,
		_w10013_,
		_w10014_
	);
	LUT2 #(
		.INIT('h4)
	) name9553 (
		_w3758_,
		_w9903_,
		_w10015_
	);
	LUT2 #(
		.INIT('h1)
	) name9554 (
		_w3417_,
		_w10015_,
		_w10016_
	);
	LUT2 #(
		.INIT('h2)
	) name9555 (
		_w5287_,
		_w5289_,
		_w10017_
	);
	LUT2 #(
		.INIT('h8)
	) name9556 (
		_w10016_,
		_w10017_,
		_w10018_
	);
	LUT2 #(
		.INIT('h2)
	) name9557 (
		\P2_reg2_reg[5]/NET0131 ,
		_w10018_,
		_w10019_
	);
	LUT2 #(
		.INIT('h8)
	) name9558 (
		_w2526_,
		_w3420_,
		_w10020_
	);
	LUT2 #(
		.INIT('h2)
	) name9559 (
		_w3758_,
		_w9852_,
		_w10021_
	);
	LUT2 #(
		.INIT('h1)
	) name9560 (
		_w10020_,
		_w10021_,
		_w10022_
	);
	LUT2 #(
		.INIT('h2)
	) name9561 (
		_w5287_,
		_w10022_,
		_w10023_
	);
	LUT2 #(
		.INIT('h1)
	) name9562 (
		_w10019_,
		_w10023_,
		_w10024_
	);
	LUT2 #(
		.INIT('h2)
	) name9563 (
		\P1_reg0_reg[14]/NET0131 ,
		_w3435_,
		_w10025_
	);
	LUT2 #(
		.INIT('h8)
	) name9564 (
		\P1_reg0_reg[14]/NET0131 ,
		_w3448_,
		_w10026_
	);
	LUT2 #(
		.INIT('h8)
	) name9565 (
		_w4396_,
		_w9307_,
		_w10027_
	);
	LUT2 #(
		.INIT('h2)
	) name9566 (
		\P1_reg0_reg[14]/NET0131 ,
		_w4396_,
		_w10028_
	);
	LUT2 #(
		.INIT('h2)
	) name9567 (
		_w4396_,
		_w8047_,
		_w10029_
	);
	LUT2 #(
		.INIT('h1)
	) name9568 (
		_w10028_,
		_w10029_,
		_w10030_
	);
	LUT2 #(
		.INIT('h2)
	) name9569 (
		_w1936_,
		_w10030_,
		_w10031_
	);
	LUT2 #(
		.INIT('h2)
	) name9570 (
		_w4396_,
		_w8058_,
		_w10032_
	);
	LUT2 #(
		.INIT('h1)
	) name9571 (
		_w10028_,
		_w10032_,
		_w10033_
	);
	LUT2 #(
		.INIT('h1)
	) name9572 (
		_w3563_,
		_w4396_,
		_w10034_
	);
	LUT2 #(
		.INIT('h2)
	) name9573 (
		_w8062_,
		_w10034_,
		_w10035_
	);
	LUT2 #(
		.INIT('h1)
	) name9574 (
		_w10033_,
		_w10035_,
		_w10036_
	);
	LUT2 #(
		.INIT('h8)
	) name9575 (
		_w4396_,
		_w8067_,
		_w10037_
	);
	LUT2 #(
		.INIT('h1)
	) name9576 (
		_w10028_,
		_w10037_,
		_w10038_
	);
	LUT2 #(
		.INIT('h2)
	) name9577 (
		_w3712_,
		_w10038_,
		_w10039_
	);
	LUT2 #(
		.INIT('h2)
	) name9578 (
		\P1_reg0_reg[14]/NET0131 ,
		_w4493_,
		_w10040_
	);
	LUT2 #(
		.INIT('h1)
	) name9579 (
		_w10027_,
		_w10040_,
		_w10041_
	);
	LUT2 #(
		.INIT('h4)
	) name9580 (
		_w10039_,
		_w10041_,
		_w10042_
	);
	LUT2 #(
		.INIT('h4)
	) name9581 (
		_w10031_,
		_w10042_,
		_w10043_
	);
	LUT2 #(
		.INIT('h4)
	) name9582 (
		_w10036_,
		_w10043_,
		_w10044_
	);
	LUT2 #(
		.INIT('h2)
	) name9583 (
		_w3450_,
		_w10044_,
		_w10045_
	);
	LUT2 #(
		.INIT('h1)
	) name9584 (
		_w10026_,
		_w10045_,
		_w10046_
	);
	LUT2 #(
		.INIT('h2)
	) name9585 (
		\P1_state_reg[0]/NET0131 ,
		_w10046_,
		_w10047_
	);
	LUT2 #(
		.INIT('h1)
	) name9586 (
		_w10025_,
		_w10047_,
		_w10048_
	);
	LUT2 #(
		.INIT('h2)
	) name9587 (
		\P1_reg0_reg[5]/NET0131 ,
		_w3435_,
		_w10049_
	);
	LUT2 #(
		.INIT('h8)
	) name9588 (
		\P1_reg0_reg[5]/NET0131 ,
		_w3448_,
		_w10050_
	);
	LUT2 #(
		.INIT('h2)
	) name9589 (
		\P1_reg0_reg[5]/NET0131 ,
		_w4491_,
		_w10051_
	);
	LUT2 #(
		.INIT('h2)
	) name9590 (
		\P1_reg0_reg[5]/NET0131 ,
		_w4396_,
		_w10052_
	);
	LUT2 #(
		.INIT('h8)
	) name9591 (
		_w4396_,
		_w9073_,
		_w10053_
	);
	LUT2 #(
		.INIT('h1)
	) name9592 (
		_w10052_,
		_w10053_,
		_w10054_
	);
	LUT2 #(
		.INIT('h2)
	) name9593 (
		_w1936_,
		_w10054_,
		_w10055_
	);
	LUT2 #(
		.INIT('h2)
	) name9594 (
		_w4396_,
		_w9079_,
		_w10056_
	);
	LUT2 #(
		.INIT('h1)
	) name9595 (
		_w10052_,
		_w10056_,
		_w10057_
	);
	LUT2 #(
		.INIT('h1)
	) name9596 (
		_w3563_,
		_w10057_,
		_w10058_
	);
	LUT2 #(
		.INIT('h2)
	) name9597 (
		_w4396_,
		_w9085_,
		_w10059_
	);
	LUT2 #(
		.INIT('h1)
	) name9598 (
		_w10052_,
		_w10059_,
		_w10060_
	);
	LUT2 #(
		.INIT('h1)
	) name9599 (
		_w3677_,
		_w10060_,
		_w10061_
	);
	LUT2 #(
		.INIT('h8)
	) name9600 (
		_w4396_,
		_w9063_,
		_w10062_
	);
	LUT2 #(
		.INIT('h1)
	) name9601 (
		_w10052_,
		_w10062_,
		_w10063_
	);
	LUT2 #(
		.INIT('h2)
	) name9602 (
		_w3712_,
		_w10063_,
		_w10064_
	);
	LUT2 #(
		.INIT('h4)
	) name9603 (
		_w1562_,
		_w4396_,
		_w10065_
	);
	LUT2 #(
		.INIT('h1)
	) name9604 (
		_w10052_,
		_w10065_,
		_w10066_
	);
	LUT2 #(
		.INIT('h2)
	) name9605 (
		_w1880_,
		_w10066_,
		_w10067_
	);
	LUT2 #(
		.INIT('h1)
	) name9606 (
		_w10051_,
		_w10067_,
		_w10068_
	);
	LUT2 #(
		.INIT('h4)
	) name9607 (
		_w10064_,
		_w10068_,
		_w10069_
	);
	LUT2 #(
		.INIT('h4)
	) name9608 (
		_w10058_,
		_w10069_,
		_w10070_
	);
	LUT2 #(
		.INIT('h4)
	) name9609 (
		_w10061_,
		_w10070_,
		_w10071_
	);
	LUT2 #(
		.INIT('h4)
	) name9610 (
		_w10055_,
		_w10071_,
		_w10072_
	);
	LUT2 #(
		.INIT('h2)
	) name9611 (
		_w3450_,
		_w10072_,
		_w10073_
	);
	LUT2 #(
		.INIT('h1)
	) name9612 (
		_w10050_,
		_w10073_,
		_w10074_
	);
	LUT2 #(
		.INIT('h2)
	) name9613 (
		\P1_state_reg[0]/NET0131 ,
		_w10074_,
		_w10075_
	);
	LUT2 #(
		.INIT('h1)
	) name9614 (
		_w10049_,
		_w10075_,
		_w10076_
	);
	LUT2 #(
		.INIT('h2)
	) name9615 (
		\P1_reg1_reg[11]/NET0131 ,
		_w3435_,
		_w10077_
	);
	LUT2 #(
		.INIT('h8)
	) name9616 (
		\P1_reg1_reg[11]/NET0131 ,
		_w3448_,
		_w10078_
	);
	LUT2 #(
		.INIT('h2)
	) name9617 (
		\P1_reg1_reg[11]/NET0131 ,
		_w4491_,
		_w10079_
	);
	LUT2 #(
		.INIT('h2)
	) name9618 (
		\P1_reg1_reg[11]/NET0131 ,
		_w4532_,
		_w10080_
	);
	LUT2 #(
		.INIT('h8)
	) name9619 (
		_w4532_,
		_w8010_,
		_w10081_
	);
	LUT2 #(
		.INIT('h1)
	) name9620 (
		_w10080_,
		_w10081_,
		_w10082_
	);
	LUT2 #(
		.INIT('h1)
	) name9621 (
		_w3563_,
		_w10082_,
		_w10083_
	);
	LUT2 #(
		.INIT('h8)
	) name9622 (
		_w4532_,
		_w8018_,
		_w10084_
	);
	LUT2 #(
		.INIT('h1)
	) name9623 (
		_w10080_,
		_w10084_,
		_w10085_
	);
	LUT2 #(
		.INIT('h2)
	) name9624 (
		_w1936_,
		_w10085_,
		_w10086_
	);
	LUT2 #(
		.INIT('h2)
	) name9625 (
		_w4532_,
		_w8004_,
		_w10087_
	);
	LUT2 #(
		.INIT('h1)
	) name9626 (
		_w10080_,
		_w10087_,
		_w10088_
	);
	LUT2 #(
		.INIT('h1)
	) name9627 (
		_w3677_,
		_w10088_,
		_w10089_
	);
	LUT2 #(
		.INIT('h8)
	) name9628 (
		_w4532_,
		_w8023_,
		_w10090_
	);
	LUT2 #(
		.INIT('h1)
	) name9629 (
		_w10080_,
		_w10090_,
		_w10091_
	);
	LUT2 #(
		.INIT('h2)
	) name9630 (
		_w3712_,
		_w10091_,
		_w10092_
	);
	LUT2 #(
		.INIT('h8)
	) name9631 (
		_w1198_,
		_w4532_,
		_w10093_
	);
	LUT2 #(
		.INIT('h1)
	) name9632 (
		_w10080_,
		_w10093_,
		_w10094_
	);
	LUT2 #(
		.INIT('h2)
	) name9633 (
		_w1880_,
		_w10094_,
		_w10095_
	);
	LUT2 #(
		.INIT('h1)
	) name9634 (
		_w10079_,
		_w10095_,
		_w10096_
	);
	LUT2 #(
		.INIT('h4)
	) name9635 (
		_w10092_,
		_w10096_,
		_w10097_
	);
	LUT2 #(
		.INIT('h4)
	) name9636 (
		_w10083_,
		_w10097_,
		_w10098_
	);
	LUT2 #(
		.INIT('h1)
	) name9637 (
		_w10086_,
		_w10089_,
		_w10099_
	);
	LUT2 #(
		.INIT('h8)
	) name9638 (
		_w10098_,
		_w10099_,
		_w10100_
	);
	LUT2 #(
		.INIT('h2)
	) name9639 (
		_w3450_,
		_w10100_,
		_w10101_
	);
	LUT2 #(
		.INIT('h1)
	) name9640 (
		_w10078_,
		_w10101_,
		_w10102_
	);
	LUT2 #(
		.INIT('h2)
	) name9641 (
		\P1_state_reg[0]/NET0131 ,
		_w10102_,
		_w10103_
	);
	LUT2 #(
		.INIT('h1)
	) name9642 (
		_w10077_,
		_w10103_,
		_w10104_
	);
	LUT2 #(
		.INIT('h2)
	) name9643 (
		\P1_reg1_reg[14]/NET0131 ,
		_w3435_,
		_w10105_
	);
	LUT2 #(
		.INIT('h8)
	) name9644 (
		\P1_reg1_reg[14]/NET0131 ,
		_w3448_,
		_w10106_
	);
	LUT2 #(
		.INIT('h8)
	) name9645 (
		_w4532_,
		_w9307_,
		_w10107_
	);
	LUT2 #(
		.INIT('h2)
	) name9646 (
		\P1_reg1_reg[14]/NET0131 ,
		_w4532_,
		_w10108_
	);
	LUT2 #(
		.INIT('h2)
	) name9647 (
		_w4532_,
		_w8047_,
		_w10109_
	);
	LUT2 #(
		.INIT('h1)
	) name9648 (
		_w10108_,
		_w10109_,
		_w10110_
	);
	LUT2 #(
		.INIT('h2)
	) name9649 (
		_w1936_,
		_w10110_,
		_w10111_
	);
	LUT2 #(
		.INIT('h2)
	) name9650 (
		_w4532_,
		_w8058_,
		_w10112_
	);
	LUT2 #(
		.INIT('h1)
	) name9651 (
		_w10108_,
		_w10112_,
		_w10113_
	);
	LUT2 #(
		.INIT('h1)
	) name9652 (
		_w3563_,
		_w4532_,
		_w10114_
	);
	LUT2 #(
		.INIT('h2)
	) name9653 (
		_w8062_,
		_w10114_,
		_w10115_
	);
	LUT2 #(
		.INIT('h1)
	) name9654 (
		_w10113_,
		_w10115_,
		_w10116_
	);
	LUT2 #(
		.INIT('h8)
	) name9655 (
		_w4532_,
		_w8067_,
		_w10117_
	);
	LUT2 #(
		.INIT('h1)
	) name9656 (
		_w10108_,
		_w10117_,
		_w10118_
	);
	LUT2 #(
		.INIT('h2)
	) name9657 (
		_w3712_,
		_w10118_,
		_w10119_
	);
	LUT2 #(
		.INIT('h2)
	) name9658 (
		\P1_reg1_reg[14]/NET0131 ,
		_w4541_,
		_w10120_
	);
	LUT2 #(
		.INIT('h1)
	) name9659 (
		_w10107_,
		_w10120_,
		_w10121_
	);
	LUT2 #(
		.INIT('h4)
	) name9660 (
		_w10119_,
		_w10121_,
		_w10122_
	);
	LUT2 #(
		.INIT('h4)
	) name9661 (
		_w10111_,
		_w10122_,
		_w10123_
	);
	LUT2 #(
		.INIT('h4)
	) name9662 (
		_w10116_,
		_w10123_,
		_w10124_
	);
	LUT2 #(
		.INIT('h2)
	) name9663 (
		_w3450_,
		_w10124_,
		_w10125_
	);
	LUT2 #(
		.INIT('h1)
	) name9664 (
		_w10106_,
		_w10125_,
		_w10126_
	);
	LUT2 #(
		.INIT('h2)
	) name9665 (
		\P1_state_reg[0]/NET0131 ,
		_w10126_,
		_w10127_
	);
	LUT2 #(
		.INIT('h1)
	) name9666 (
		_w10105_,
		_w10127_,
		_w10128_
	);
	LUT2 #(
		.INIT('h2)
	) name9667 (
		\P2_reg0_reg[11]/NET0131 ,
		_w1983_,
		_w10129_
	);
	LUT2 #(
		.INIT('h8)
	) name9668 (
		\P2_reg0_reg[11]/NET0131 ,
		_w2024_,
		_w10130_
	);
	LUT2 #(
		.INIT('h2)
	) name9669 (
		\P2_reg0_reg[11]/NET0131 ,
		_w8385_,
		_w10131_
	);
	LUT2 #(
		.INIT('h2)
	) name9670 (
		\P2_reg0_reg[11]/NET0131 ,
		_w2040_,
		_w10132_
	);
	LUT2 #(
		.INIT('h8)
	) name9671 (
		_w2040_,
		_w8129_,
		_w10133_
	);
	LUT2 #(
		.INIT('h1)
	) name9672 (
		_w10132_,
		_w10133_,
		_w10134_
	);
	LUT2 #(
		.INIT('h2)
	) name9673 (
		_w3411_,
		_w10134_,
		_w10135_
	);
	LUT2 #(
		.INIT('h8)
	) name9674 (
		_w2040_,
		_w8135_,
		_w10136_
	);
	LUT2 #(
		.INIT('h1)
	) name9675 (
		_w10132_,
		_w10136_,
		_w10137_
	);
	LUT2 #(
		.INIT('h1)
	) name9676 (
		_w3177_,
		_w10137_,
		_w10138_
	);
	LUT2 #(
		.INIT('h2)
	) name9677 (
		_w2040_,
		_w9867_,
		_w10139_
	);
	LUT2 #(
		.INIT('h1)
	) name9678 (
		_w10131_,
		_w10139_,
		_w10140_
	);
	LUT2 #(
		.INIT('h4)
	) name9679 (
		_w10138_,
		_w10140_,
		_w10141_
	);
	LUT2 #(
		.INIT('h4)
	) name9680 (
		_w10135_,
		_w10141_,
		_w10142_
	);
	LUT2 #(
		.INIT('h2)
	) name9681 (
		_w2026_,
		_w10142_,
		_w10143_
	);
	LUT2 #(
		.INIT('h1)
	) name9682 (
		_w10130_,
		_w10143_,
		_w10144_
	);
	LUT2 #(
		.INIT('h2)
	) name9683 (
		\P1_state_reg[0]/NET0131 ,
		_w10144_,
		_w10145_
	);
	LUT2 #(
		.INIT('h1)
	) name9684 (
		_w10129_,
		_w10145_,
		_w10146_
	);
	LUT2 #(
		.INIT('h2)
	) name9685 (
		\P2_reg0_reg[14]/NET0131 ,
		_w1983_,
		_w10147_
	);
	LUT2 #(
		.INIT('h8)
	) name9686 (
		\P2_reg0_reg[14]/NET0131 ,
		_w2024_,
		_w10148_
	);
	LUT2 #(
		.INIT('h2)
	) name9687 (
		\P2_reg0_reg[14]/NET0131 ,
		_w3423_,
		_w10149_
	);
	LUT2 #(
		.INIT('h8)
	) name9688 (
		_w2040_,
		_w9437_,
		_w10150_
	);
	LUT2 #(
		.INIT('h2)
	) name9689 (
		\P2_reg0_reg[14]/NET0131 ,
		_w2040_,
		_w10151_
	);
	LUT2 #(
		.INIT('h8)
	) name9690 (
		_w2040_,
		_w8176_,
		_w10152_
	);
	LUT2 #(
		.INIT('h1)
	) name9691 (
		_w10151_,
		_w10152_,
		_w10153_
	);
	LUT2 #(
		.INIT('h2)
	) name9692 (
		_w3355_,
		_w10153_,
		_w10154_
	);
	LUT2 #(
		.INIT('h8)
	) name9693 (
		_w2040_,
		_w8182_,
		_w10155_
	);
	LUT2 #(
		.INIT('h1)
	) name9694 (
		_w10151_,
		_w10155_,
		_w10156_
	);
	LUT2 #(
		.INIT('h1)
	) name9695 (
		_w3177_,
		_w10156_,
		_w10157_
	);
	LUT2 #(
		.INIT('h2)
	) name9696 (
		_w2040_,
		_w8188_,
		_w10158_
	);
	LUT2 #(
		.INIT('h1)
	) name9697 (
		_w10151_,
		_w10158_,
		_w10159_
	);
	LUT2 #(
		.INIT('h1)
	) name9698 (
		_w3320_,
		_w10159_,
		_w10160_
	);
	LUT2 #(
		.INIT('h8)
	) name9699 (
		_w2040_,
		_w8171_,
		_w10161_
	);
	LUT2 #(
		.INIT('h1)
	) name9700 (
		_w10151_,
		_w10161_,
		_w10162_
	);
	LUT2 #(
		.INIT('h2)
	) name9701 (
		_w3411_,
		_w10162_,
		_w10163_
	);
	LUT2 #(
		.INIT('h1)
	) name9702 (
		_w10149_,
		_w10150_,
		_w10164_
	);
	LUT2 #(
		.INIT('h4)
	) name9703 (
		_w10154_,
		_w10164_,
		_w10165_
	);
	LUT2 #(
		.INIT('h1)
	) name9704 (
		_w10157_,
		_w10160_,
		_w10166_
	);
	LUT2 #(
		.INIT('h4)
	) name9705 (
		_w10163_,
		_w10166_,
		_w10167_
	);
	LUT2 #(
		.INIT('h8)
	) name9706 (
		_w10165_,
		_w10167_,
		_w10168_
	);
	LUT2 #(
		.INIT('h2)
	) name9707 (
		_w2026_,
		_w10168_,
		_w10169_
	);
	LUT2 #(
		.INIT('h1)
	) name9708 (
		_w10148_,
		_w10169_,
		_w10170_
	);
	LUT2 #(
		.INIT('h2)
	) name9709 (
		\P1_state_reg[0]/NET0131 ,
		_w10170_,
		_w10171_
	);
	LUT2 #(
		.INIT('h1)
	) name9710 (
		_w10147_,
		_w10171_,
		_w10172_
	);
	LUT2 #(
		.INIT('h2)
	) name9711 (
		\P1_reg1_reg[3]/NET0131 ,
		_w3435_,
		_w10173_
	);
	LUT2 #(
		.INIT('h8)
	) name9712 (
		\P1_reg1_reg[3]/NET0131 ,
		_w3448_,
		_w10174_
	);
	LUT2 #(
		.INIT('h4)
	) name9713 (
		_w3677_,
		_w9723_,
		_w10175_
	);
	LUT2 #(
		.INIT('h2)
	) name9714 (
		_w9702_,
		_w10175_,
		_w10176_
	);
	LUT2 #(
		.INIT('h2)
	) name9715 (
		_w4532_,
		_w10176_,
		_w10177_
	);
	LUT2 #(
		.INIT('h2)
	) name9716 (
		\P1_reg1_reg[3]/NET0131 ,
		_w4532_,
		_w10178_
	);
	LUT2 #(
		.INIT('h8)
	) name9717 (
		_w4532_,
		_w9709_,
		_w10179_
	);
	LUT2 #(
		.INIT('h1)
	) name9718 (
		_w10178_,
		_w10179_,
		_w10180_
	);
	LUT2 #(
		.INIT('h2)
	) name9719 (
		_w1936_,
		_w10180_,
		_w10181_
	);
	LUT2 #(
		.INIT('h2)
	) name9720 (
		_w4532_,
		_w9716_,
		_w10182_
	);
	LUT2 #(
		.INIT('h1)
	) name9721 (
		_w10178_,
		_w10182_,
		_w10183_
	);
	LUT2 #(
		.INIT('h1)
	) name9722 (
		_w3563_,
		_w10183_,
		_w10184_
	);
	LUT2 #(
		.INIT('h1)
	) name9723 (
		_w3677_,
		_w4532_,
		_w10185_
	);
	LUT2 #(
		.INIT('h2)
	) name9724 (
		_w9835_,
		_w10185_,
		_w10186_
	);
	LUT2 #(
		.INIT('h2)
	) name9725 (
		\P1_reg1_reg[3]/NET0131 ,
		_w10186_,
		_w10187_
	);
	LUT2 #(
		.INIT('h1)
	) name9726 (
		_w10177_,
		_w10187_,
		_w10188_
	);
	LUT2 #(
		.INIT('h4)
	) name9727 (
		_w10184_,
		_w10188_,
		_w10189_
	);
	LUT2 #(
		.INIT('h4)
	) name9728 (
		_w10181_,
		_w10189_,
		_w10190_
	);
	LUT2 #(
		.INIT('h2)
	) name9729 (
		_w3450_,
		_w10190_,
		_w10191_
	);
	LUT2 #(
		.INIT('h1)
	) name9730 (
		_w10174_,
		_w10191_,
		_w10192_
	);
	LUT2 #(
		.INIT('h2)
	) name9731 (
		\P1_state_reg[0]/NET0131 ,
		_w10192_,
		_w10193_
	);
	LUT2 #(
		.INIT('h1)
	) name9732 (
		_w10173_,
		_w10193_,
		_w10194_
	);
	LUT2 #(
		.INIT('h2)
	) name9733 (
		\P1_reg1_reg[7]/NET0131 ,
		_w3435_,
		_w10195_
	);
	LUT2 #(
		.INIT('h8)
	) name9734 (
		\P1_reg1_reg[7]/NET0131 ,
		_w3448_,
		_w10196_
	);
	LUT2 #(
		.INIT('h2)
	) name9735 (
		\P1_reg1_reg[7]/NET0131 ,
		_w4573_,
		_w10197_
	);
	LUT2 #(
		.INIT('h2)
	) name9736 (
		\P1_reg1_reg[7]/NET0131 ,
		_w4532_,
		_w10198_
	);
	LUT2 #(
		.INIT('h8)
	) name9737 (
		_w4532_,
		_w9794_,
		_w10199_
	);
	LUT2 #(
		.INIT('h1)
	) name9738 (
		_w10198_,
		_w10199_,
		_w10200_
	);
	LUT2 #(
		.INIT('h1)
	) name9739 (
		_w3563_,
		_w10200_,
		_w10201_
	);
	LUT2 #(
		.INIT('h8)
	) name9740 (
		_w4532_,
		_w9802_,
		_w10202_
	);
	LUT2 #(
		.INIT('h1)
	) name9741 (
		_w10198_,
		_w10202_,
		_w10203_
	);
	LUT2 #(
		.INIT('h2)
	) name9742 (
		_w1936_,
		_w10203_,
		_w10204_
	);
	LUT2 #(
		.INIT('h2)
	) name9743 (
		_w4532_,
		_w9788_,
		_w10205_
	);
	LUT2 #(
		.INIT('h1)
	) name9744 (
		_w10198_,
		_w10205_,
		_w10206_
	);
	LUT2 #(
		.INIT('h1)
	) name9745 (
		_w3677_,
		_w10206_,
		_w10207_
	);
	LUT2 #(
		.INIT('h4)
	) name9746 (
		_w1514_,
		_w1880_,
		_w10208_
	);
	LUT2 #(
		.INIT('h1)
	) name9747 (
		_w9808_,
		_w10208_,
		_w10209_
	);
	LUT2 #(
		.INIT('h2)
	) name9748 (
		_w4532_,
		_w10209_,
		_w10210_
	);
	LUT2 #(
		.INIT('h1)
	) name9749 (
		_w10197_,
		_w10210_,
		_w10211_
	);
	LUT2 #(
		.INIT('h4)
	) name9750 (
		_w10201_,
		_w10211_,
		_w10212_
	);
	LUT2 #(
		.INIT('h1)
	) name9751 (
		_w10204_,
		_w10207_,
		_w10213_
	);
	LUT2 #(
		.INIT('h8)
	) name9752 (
		_w10212_,
		_w10213_,
		_w10214_
	);
	LUT2 #(
		.INIT('h2)
	) name9753 (
		_w3450_,
		_w10214_,
		_w10215_
	);
	LUT2 #(
		.INIT('h1)
	) name9754 (
		_w10196_,
		_w10215_,
		_w10216_
	);
	LUT2 #(
		.INIT('h2)
	) name9755 (
		\P1_state_reg[0]/NET0131 ,
		_w10216_,
		_w10217_
	);
	LUT2 #(
		.INIT('h1)
	) name9756 (
		_w10195_,
		_w10217_,
		_w10218_
	);
	LUT2 #(
		.INIT('h2)
	) name9757 (
		\P2_reg0_reg[3]/NET0131 ,
		_w1983_,
		_w10219_
	);
	LUT2 #(
		.INIT('h8)
	) name9758 (
		\P2_reg0_reg[3]/NET0131 ,
		_w2024_,
		_w10220_
	);
	LUT2 #(
		.INIT('h2)
	) name9759 (
		_w2040_,
		_w9587_,
		_w10221_
	);
	LUT2 #(
		.INIT('h2)
	) name9760 (
		\P2_reg0_reg[3]/NET0131 ,
		_w2040_,
		_w10222_
	);
	LUT2 #(
		.INIT('h8)
	) name9761 (
		_w2040_,
		_w9597_,
		_w10223_
	);
	LUT2 #(
		.INIT('h1)
	) name9762 (
		_w10222_,
		_w10223_,
		_w10224_
	);
	LUT2 #(
		.INIT('h2)
	) name9763 (
		_w3411_,
		_w10224_,
		_w10225_
	);
	LUT2 #(
		.INIT('h2)
	) name9764 (
		_w2040_,
		_w9591_,
		_w10226_
	);
	LUT2 #(
		.INIT('h1)
	) name9765 (
		_w10222_,
		_w10226_,
		_w10227_
	);
	LUT2 #(
		.INIT('h1)
	) name9766 (
		_w3177_,
		_w10227_,
		_w10228_
	);
	LUT2 #(
		.INIT('h1)
	) name9767 (
		_w2040_,
		_w9904_,
		_w10229_
	);
	LUT2 #(
		.INIT('h2)
	) name9768 (
		_w3421_,
		_w10229_,
		_w10230_
	);
	LUT2 #(
		.INIT('h2)
	) name9769 (
		\P2_reg0_reg[3]/NET0131 ,
		_w10230_,
		_w10231_
	);
	LUT2 #(
		.INIT('h1)
	) name9770 (
		_w10221_,
		_w10231_,
		_w10232_
	);
	LUT2 #(
		.INIT('h4)
	) name9771 (
		_w10228_,
		_w10232_,
		_w10233_
	);
	LUT2 #(
		.INIT('h4)
	) name9772 (
		_w10225_,
		_w10233_,
		_w10234_
	);
	LUT2 #(
		.INIT('h2)
	) name9773 (
		_w2026_,
		_w10234_,
		_w10235_
	);
	LUT2 #(
		.INIT('h1)
	) name9774 (
		_w10220_,
		_w10235_,
		_w10236_
	);
	LUT2 #(
		.INIT('h2)
	) name9775 (
		\P1_state_reg[0]/NET0131 ,
		_w10236_,
		_w10237_
	);
	LUT2 #(
		.INIT('h1)
	) name9776 (
		_w10219_,
		_w10237_,
		_w10238_
	);
	LUT2 #(
		.INIT('h2)
	) name9777 (
		\P2_reg0_reg[7]/NET0131 ,
		_w1983_,
		_w10239_
	);
	LUT2 #(
		.INIT('h8)
	) name9778 (
		\P2_reg0_reg[7]/NET0131 ,
		_w2024_,
		_w10240_
	);
	LUT2 #(
		.INIT('h2)
	) name9779 (
		\P2_reg0_reg[7]/NET0131 ,
		_w8385_,
		_w10241_
	);
	LUT2 #(
		.INIT('h2)
	) name9780 (
		\P2_reg0_reg[7]/NET0131 ,
		_w2040_,
		_w10242_
	);
	LUT2 #(
		.INIT('h8)
	) name9781 (
		_w2040_,
		_w9664_,
		_w10243_
	);
	LUT2 #(
		.INIT('h1)
	) name9782 (
		_w10242_,
		_w10243_,
		_w10244_
	);
	LUT2 #(
		.INIT('h2)
	) name9783 (
		_w3411_,
		_w10244_,
		_w10245_
	);
	LUT2 #(
		.INIT('h8)
	) name9784 (
		_w2040_,
		_w9670_,
		_w10246_
	);
	LUT2 #(
		.INIT('h1)
	) name9785 (
		_w10242_,
		_w10246_,
		_w10247_
	);
	LUT2 #(
		.INIT('h1)
	) name9786 (
		_w3177_,
		_w10247_,
		_w10248_
	);
	LUT2 #(
		.INIT('h8)
	) name9787 (
		_w2495_,
		_w3358_,
		_w10249_
	);
	LUT2 #(
		.INIT('h1)
	) name9788 (
		_w3320_,
		_w9676_,
		_w10250_
	);
	LUT2 #(
		.INIT('h1)
	) name9789 (
		_w9682_,
		_w10249_,
		_w10251_
	);
	LUT2 #(
		.INIT('h4)
	) name9790 (
		_w10250_,
		_w10251_,
		_w10252_
	);
	LUT2 #(
		.INIT('h2)
	) name9791 (
		_w2040_,
		_w10252_,
		_w10253_
	);
	LUT2 #(
		.INIT('h1)
	) name9792 (
		_w10241_,
		_w10253_,
		_w10254_
	);
	LUT2 #(
		.INIT('h4)
	) name9793 (
		_w10248_,
		_w10254_,
		_w10255_
	);
	LUT2 #(
		.INIT('h4)
	) name9794 (
		_w10245_,
		_w10255_,
		_w10256_
	);
	LUT2 #(
		.INIT('h2)
	) name9795 (
		_w2026_,
		_w10256_,
		_w10257_
	);
	LUT2 #(
		.INIT('h1)
	) name9796 (
		_w10240_,
		_w10257_,
		_w10258_
	);
	LUT2 #(
		.INIT('h2)
	) name9797 (
		\P1_state_reg[0]/NET0131 ,
		_w10258_,
		_w10259_
	);
	LUT2 #(
		.INIT('h1)
	) name9798 (
		_w10239_,
		_w10259_,
		_w10260_
	);
	LUT2 #(
		.INIT('h2)
	) name9799 (
		\P2_reg1_reg[3]/NET0131 ,
		_w1983_,
		_w10261_
	);
	LUT2 #(
		.INIT('h8)
	) name9800 (
		\P2_reg1_reg[3]/NET0131 ,
		_w2024_,
		_w10262_
	);
	LUT2 #(
		.INIT('h2)
	) name9801 (
		\P2_reg1_reg[3]/NET0131 ,
		_w9906_,
		_w10263_
	);
	LUT2 #(
		.INIT('h2)
	) name9802 (
		\P2_reg1_reg[3]/NET0131 ,
		_w3733_,
		_w10264_
	);
	LUT2 #(
		.INIT('h8)
	) name9803 (
		_w3733_,
		_w9597_,
		_w10265_
	);
	LUT2 #(
		.INIT('h1)
	) name9804 (
		_w10264_,
		_w10265_,
		_w10266_
	);
	LUT2 #(
		.INIT('h2)
	) name9805 (
		_w3411_,
		_w10266_,
		_w10267_
	);
	LUT2 #(
		.INIT('h2)
	) name9806 (
		_w3733_,
		_w9591_,
		_w10268_
	);
	LUT2 #(
		.INIT('h1)
	) name9807 (
		_w10264_,
		_w10268_,
		_w10269_
	);
	LUT2 #(
		.INIT('h1)
	) name9808 (
		_w3177_,
		_w10269_,
		_w10270_
	);
	LUT2 #(
		.INIT('h2)
	) name9809 (
		_w3733_,
		_w9587_,
		_w10271_
	);
	LUT2 #(
		.INIT('h1)
	) name9810 (
		_w10263_,
		_w10271_,
		_w10272_
	);
	LUT2 #(
		.INIT('h4)
	) name9811 (
		_w10270_,
		_w10272_,
		_w10273_
	);
	LUT2 #(
		.INIT('h4)
	) name9812 (
		_w10267_,
		_w10273_,
		_w10274_
	);
	LUT2 #(
		.INIT('h2)
	) name9813 (
		_w2026_,
		_w10274_,
		_w10275_
	);
	LUT2 #(
		.INIT('h1)
	) name9814 (
		_w10262_,
		_w10275_,
		_w10276_
	);
	LUT2 #(
		.INIT('h2)
	) name9815 (
		\P1_state_reg[0]/NET0131 ,
		_w10276_,
		_w10277_
	);
	LUT2 #(
		.INIT('h1)
	) name9816 (
		_w10261_,
		_w10277_,
		_w10278_
	);
	LUT2 #(
		.INIT('h2)
	) name9817 (
		\P2_reg1_reg[7]/NET0131 ,
		_w1983_,
		_w10279_
	);
	LUT2 #(
		.INIT('h8)
	) name9818 (
		\P2_reg1_reg[7]/NET0131 ,
		_w2024_,
		_w10280_
	);
	LUT2 #(
		.INIT('h2)
	) name9819 (
		\P2_reg1_reg[7]/NET0131 ,
		_w8532_,
		_w10281_
	);
	LUT2 #(
		.INIT('h2)
	) name9820 (
		\P2_reg1_reg[7]/NET0131 ,
		_w3733_,
		_w10282_
	);
	LUT2 #(
		.INIT('h8)
	) name9821 (
		_w3733_,
		_w9664_,
		_w10283_
	);
	LUT2 #(
		.INIT('h1)
	) name9822 (
		_w10282_,
		_w10283_,
		_w10284_
	);
	LUT2 #(
		.INIT('h2)
	) name9823 (
		_w3411_,
		_w10284_,
		_w10285_
	);
	LUT2 #(
		.INIT('h8)
	) name9824 (
		_w3733_,
		_w9670_,
		_w10286_
	);
	LUT2 #(
		.INIT('h1)
	) name9825 (
		_w10282_,
		_w10286_,
		_w10287_
	);
	LUT2 #(
		.INIT('h1)
	) name9826 (
		_w3177_,
		_w10287_,
		_w10288_
	);
	LUT2 #(
		.INIT('h2)
	) name9827 (
		_w3733_,
		_w10252_,
		_w10289_
	);
	LUT2 #(
		.INIT('h1)
	) name9828 (
		_w10281_,
		_w10289_,
		_w10290_
	);
	LUT2 #(
		.INIT('h4)
	) name9829 (
		_w10288_,
		_w10290_,
		_w10291_
	);
	LUT2 #(
		.INIT('h4)
	) name9830 (
		_w10285_,
		_w10291_,
		_w10292_
	);
	LUT2 #(
		.INIT('h2)
	) name9831 (
		_w2026_,
		_w10292_,
		_w10293_
	);
	LUT2 #(
		.INIT('h1)
	) name9832 (
		_w10280_,
		_w10293_,
		_w10294_
	);
	LUT2 #(
		.INIT('h2)
	) name9833 (
		\P1_state_reg[0]/NET0131 ,
		_w10294_,
		_w10295_
	);
	LUT2 #(
		.INIT('h1)
	) name9834 (
		_w10279_,
		_w10295_,
		_w10296_
	);
	LUT2 #(
		.INIT('h2)
	) name9835 (
		\P1_reg2_reg[3]/NET0131 ,
		_w3435_,
		_w10297_
	);
	LUT2 #(
		.INIT('h8)
	) name9836 (
		\P1_reg2_reg[3]/NET0131 ,
		_w3448_,
		_w10298_
	);
	LUT2 #(
		.INIT('h2)
	) name9837 (
		_w3466_,
		_w9702_,
		_w10299_
	);
	LUT2 #(
		.INIT('h2)
	) name9838 (
		\P1_reg2_reg[3]/NET0131 ,
		_w3466_,
		_w10300_
	);
	LUT2 #(
		.INIT('h8)
	) name9839 (
		_w3466_,
		_w9709_,
		_w10301_
	);
	LUT2 #(
		.INIT('h1)
	) name9840 (
		_w10300_,
		_w10301_,
		_w10302_
	);
	LUT2 #(
		.INIT('h2)
	) name9841 (
		_w1936_,
		_w10302_,
		_w10303_
	);
	LUT2 #(
		.INIT('h2)
	) name9842 (
		_w3466_,
		_w9716_,
		_w10304_
	);
	LUT2 #(
		.INIT('h1)
	) name9843 (
		_w10300_,
		_w10304_,
		_w10305_
	);
	LUT2 #(
		.INIT('h1)
	) name9844 (
		_w3563_,
		_w10305_,
		_w10306_
	);
	LUT2 #(
		.INIT('h8)
	) name9845 (
		_w3466_,
		_w9723_,
		_w10307_
	);
	LUT2 #(
		.INIT('h1)
	) name9846 (
		_w10300_,
		_w10307_,
		_w10308_
	);
	LUT2 #(
		.INIT('h1)
	) name9847 (
		_w3677_,
		_w10308_,
		_w10309_
	);
	LUT2 #(
		.INIT('h4)
	) name9848 (
		\P1_reg3_reg[3]/NET0131 ,
		_w1763_,
		_w10310_
	);
	LUT2 #(
		.INIT('h2)
	) name9849 (
		\P1_reg2_reg[3]/NET0131 ,
		_w9954_,
		_w10311_
	);
	LUT2 #(
		.INIT('h1)
	) name9850 (
		_w10310_,
		_w10311_,
		_w10312_
	);
	LUT2 #(
		.INIT('h4)
	) name9851 (
		_w10299_,
		_w10312_,
		_w10313_
	);
	LUT2 #(
		.INIT('h4)
	) name9852 (
		_w10309_,
		_w10313_,
		_w10314_
	);
	LUT2 #(
		.INIT('h4)
	) name9853 (
		_w10306_,
		_w10314_,
		_w10315_
	);
	LUT2 #(
		.INIT('h4)
	) name9854 (
		_w10303_,
		_w10315_,
		_w10316_
	);
	LUT2 #(
		.INIT('h2)
	) name9855 (
		_w3450_,
		_w10316_,
		_w10317_
	);
	LUT2 #(
		.INIT('h1)
	) name9856 (
		_w10298_,
		_w10317_,
		_w10318_
	);
	LUT2 #(
		.INIT('h2)
	) name9857 (
		\P1_state_reg[0]/NET0131 ,
		_w10318_,
		_w10319_
	);
	LUT2 #(
		.INIT('h1)
	) name9858 (
		_w10297_,
		_w10319_,
		_w10320_
	);
	LUT2 #(
		.INIT('h2)
	) name9859 (
		\P1_reg2_reg[6]/NET0131 ,
		_w3435_,
		_w10321_
	);
	LUT2 #(
		.INIT('h8)
	) name9860 (
		\P1_reg2_reg[6]/NET0131 ,
		_w3448_,
		_w10322_
	);
	LUT2 #(
		.INIT('h4)
	) name9861 (
		_w1537_,
		_w1880_,
		_w10323_
	);
	LUT2 #(
		.INIT('h8)
	) name9862 (
		_w3466_,
		_w10323_,
		_w10324_
	);
	LUT2 #(
		.INIT('h2)
	) name9863 (
		\P1_reg2_reg[6]/NET0131 ,
		_w3466_,
		_w10325_
	);
	LUT2 #(
		.INIT('h8)
	) name9864 (
		_w3466_,
		_w9755_,
		_w10326_
	);
	LUT2 #(
		.INIT('h1)
	) name9865 (
		_w10325_,
		_w10326_,
		_w10327_
	);
	LUT2 #(
		.INIT('h1)
	) name9866 (
		_w3677_,
		_w10327_,
		_w10328_
	);
	LUT2 #(
		.INIT('h2)
	) name9867 (
		_w3466_,
		_w9761_,
		_w10329_
	);
	LUT2 #(
		.INIT('h1)
	) name9868 (
		_w10325_,
		_w10329_,
		_w10330_
	);
	LUT2 #(
		.INIT('h1)
	) name9869 (
		_w3563_,
		_w10330_,
		_w10331_
	);
	LUT2 #(
		.INIT('h2)
	) name9870 (
		_w3466_,
		_w9749_,
		_w10332_
	);
	LUT2 #(
		.INIT('h1)
	) name9871 (
		_w10325_,
		_w10332_,
		_w10333_
	);
	LUT2 #(
		.INIT('h2)
	) name9872 (
		_w1936_,
		_w10333_,
		_w10334_
	);
	LUT2 #(
		.INIT('h8)
	) name9873 (
		_w3466_,
		_w9766_,
		_w10335_
	);
	LUT2 #(
		.INIT('h1)
	) name9874 (
		_w10325_,
		_w10335_,
		_w10336_
	);
	LUT2 #(
		.INIT('h2)
	) name9875 (
		_w3712_,
		_w10336_,
		_w10337_
	);
	LUT2 #(
		.INIT('h8)
	) name9876 (
		_w1518_,
		_w1763_,
		_w10338_
	);
	LUT2 #(
		.INIT('h2)
	) name9877 (
		\P1_reg2_reg[6]/NET0131 ,
		_w3718_,
		_w10339_
	);
	LUT2 #(
		.INIT('h1)
	) name9878 (
		_w10324_,
		_w10338_,
		_w10340_
	);
	LUT2 #(
		.INIT('h4)
	) name9879 (
		_w10339_,
		_w10340_,
		_w10341_
	);
	LUT2 #(
		.INIT('h4)
	) name9880 (
		_w10337_,
		_w10341_,
		_w10342_
	);
	LUT2 #(
		.INIT('h4)
	) name9881 (
		_w10328_,
		_w10342_,
		_w10343_
	);
	LUT2 #(
		.INIT('h1)
	) name9882 (
		_w10331_,
		_w10334_,
		_w10344_
	);
	LUT2 #(
		.INIT('h8)
	) name9883 (
		_w10343_,
		_w10344_,
		_w10345_
	);
	LUT2 #(
		.INIT('h2)
	) name9884 (
		_w3450_,
		_w10345_,
		_w10346_
	);
	LUT2 #(
		.INIT('h1)
	) name9885 (
		_w10322_,
		_w10346_,
		_w10347_
	);
	LUT2 #(
		.INIT('h2)
	) name9886 (
		\P1_state_reg[0]/NET0131 ,
		_w10347_,
		_w10348_
	);
	LUT2 #(
		.INIT('h1)
	) name9887 (
		_w10321_,
		_w10348_,
		_w10349_
	);
	LUT2 #(
		.INIT('h2)
	) name9888 (
		\P1_reg2_reg[7]/NET0131 ,
		_w3435_,
		_w10350_
	);
	LUT2 #(
		.INIT('h8)
	) name9889 (
		\P1_reg2_reg[7]/NET0131 ,
		_w3448_,
		_w10351_
	);
	LUT2 #(
		.INIT('h2)
	) name9890 (
		\P1_reg2_reg[7]/NET0131 ,
		_w5914_,
		_w10352_
	);
	LUT2 #(
		.INIT('h2)
	) name9891 (
		\P1_reg2_reg[7]/NET0131 ,
		_w3466_,
		_w10353_
	);
	LUT2 #(
		.INIT('h8)
	) name9892 (
		_w3466_,
		_w9794_,
		_w10354_
	);
	LUT2 #(
		.INIT('h1)
	) name9893 (
		_w10353_,
		_w10354_,
		_w10355_
	);
	LUT2 #(
		.INIT('h1)
	) name9894 (
		_w3563_,
		_w10355_,
		_w10356_
	);
	LUT2 #(
		.INIT('h8)
	) name9895 (
		_w3466_,
		_w9802_,
		_w10357_
	);
	LUT2 #(
		.INIT('h1)
	) name9896 (
		_w10353_,
		_w10357_,
		_w10358_
	);
	LUT2 #(
		.INIT('h2)
	) name9897 (
		_w1936_,
		_w10358_,
		_w10359_
	);
	LUT2 #(
		.INIT('h2)
	) name9898 (
		_w3466_,
		_w9788_,
		_w10360_
	);
	LUT2 #(
		.INIT('h1)
	) name9899 (
		_w10353_,
		_w10360_,
		_w10361_
	);
	LUT2 #(
		.INIT('h1)
	) name9900 (
		_w3677_,
		_w10361_,
		_w10362_
	);
	LUT2 #(
		.INIT('h2)
	) name9901 (
		_w3466_,
		_w10209_,
		_w10363_
	);
	LUT2 #(
		.INIT('h8)
	) name9902 (
		_w1491_,
		_w1763_,
		_w10364_
	);
	LUT2 #(
		.INIT('h1)
	) name9903 (
		_w10352_,
		_w10364_,
		_w10365_
	);
	LUT2 #(
		.INIT('h4)
	) name9904 (
		_w10363_,
		_w10365_,
		_w10366_
	);
	LUT2 #(
		.INIT('h4)
	) name9905 (
		_w10356_,
		_w10366_,
		_w10367_
	);
	LUT2 #(
		.INIT('h1)
	) name9906 (
		_w10359_,
		_w10362_,
		_w10368_
	);
	LUT2 #(
		.INIT('h8)
	) name9907 (
		_w10367_,
		_w10368_,
		_w10369_
	);
	LUT2 #(
		.INIT('h2)
	) name9908 (
		_w3450_,
		_w10369_,
		_w10370_
	);
	LUT2 #(
		.INIT('h1)
	) name9909 (
		_w10351_,
		_w10370_,
		_w10371_
	);
	LUT2 #(
		.INIT('h2)
	) name9910 (
		\P1_state_reg[0]/NET0131 ,
		_w10371_,
		_w10372_
	);
	LUT2 #(
		.INIT('h1)
	) name9911 (
		_w10350_,
		_w10372_,
		_w10373_
	);
	LUT2 #(
		.INIT('h2)
	) name9912 (
		\P2_reg2_reg[3]/NET0131 ,
		_w1983_,
		_w10374_
	);
	LUT2 #(
		.INIT('h8)
	) name9913 (
		\P2_reg2_reg[3]/NET0131 ,
		_w2024_,
		_w10375_
	);
	LUT2 #(
		.INIT('h4)
	) name9914 (
		\P2_reg3_reg[3]/NET0131 ,
		_w3420_,
		_w10376_
	);
	LUT2 #(
		.INIT('h2)
	) name9915 (
		\P2_reg2_reg[3]/NET0131 ,
		_w3758_,
		_w10377_
	);
	LUT2 #(
		.INIT('h8)
	) name9916 (
		_w3758_,
		_w9597_,
		_w10378_
	);
	LUT2 #(
		.INIT('h1)
	) name9917 (
		_w10377_,
		_w10378_,
		_w10379_
	);
	LUT2 #(
		.INIT('h2)
	) name9918 (
		_w3411_,
		_w10379_,
		_w10380_
	);
	LUT2 #(
		.INIT('h2)
	) name9919 (
		_w3758_,
		_w9591_,
		_w10381_
	);
	LUT2 #(
		.INIT('h1)
	) name9920 (
		_w10377_,
		_w10381_,
		_w10382_
	);
	LUT2 #(
		.INIT('h1)
	) name9921 (
		_w3177_,
		_w10382_,
		_w10383_
	);
	LUT2 #(
		.INIT('h2)
	) name9922 (
		_w3758_,
		_w9587_,
		_w10384_
	);
	LUT2 #(
		.INIT('h4)
	) name9923 (
		_w7769_,
		_w10016_,
		_w10385_
	);
	LUT2 #(
		.INIT('h2)
	) name9924 (
		\P2_reg2_reg[3]/NET0131 ,
		_w10385_,
		_w10386_
	);
	LUT2 #(
		.INIT('h1)
	) name9925 (
		_w10376_,
		_w10386_,
		_w10387_
	);
	LUT2 #(
		.INIT('h4)
	) name9926 (
		_w10384_,
		_w10387_,
		_w10388_
	);
	LUT2 #(
		.INIT('h4)
	) name9927 (
		_w10383_,
		_w10388_,
		_w10389_
	);
	LUT2 #(
		.INIT('h4)
	) name9928 (
		_w10380_,
		_w10389_,
		_w10390_
	);
	LUT2 #(
		.INIT('h2)
	) name9929 (
		_w2026_,
		_w10390_,
		_w10391_
	);
	LUT2 #(
		.INIT('h1)
	) name9930 (
		_w10375_,
		_w10391_,
		_w10392_
	);
	LUT2 #(
		.INIT('h2)
	) name9931 (
		\P1_state_reg[0]/NET0131 ,
		_w10392_,
		_w10393_
	);
	LUT2 #(
		.INIT('h1)
	) name9932 (
		_w10374_,
		_w10393_,
		_w10394_
	);
	LUT2 #(
		.INIT('h2)
	) name9933 (
		\P2_reg2_reg[6]/NET0131 ,
		_w1983_,
		_w10395_
	);
	LUT2 #(
		.INIT('h8)
	) name9934 (
		\P2_reg2_reg[6]/NET0131 ,
		_w2024_,
		_w10396_
	);
	LUT2 #(
		.INIT('h4)
	) name9935 (
		_w2521_,
		_w3358_,
		_w10397_
	);
	LUT2 #(
		.INIT('h8)
	) name9936 (
		_w3758_,
		_w10397_,
		_w10398_
	);
	LUT2 #(
		.INIT('h2)
	) name9937 (
		\P2_reg2_reg[6]/NET0131 ,
		_w3758_,
		_w10399_
	);
	LUT2 #(
		.INIT('h8)
	) name9938 (
		_w3758_,
		_w9624_,
		_w10400_
	);
	LUT2 #(
		.INIT('h1)
	) name9939 (
		_w10399_,
		_w10400_,
		_w10401_
	);
	LUT2 #(
		.INIT('h2)
	) name9940 (
		_w3411_,
		_w10401_,
		_w10402_
	);
	LUT2 #(
		.INIT('h2)
	) name9941 (
		_w3758_,
		_w9630_,
		_w10403_
	);
	LUT2 #(
		.INIT('h1)
	) name9942 (
		_w10399_,
		_w10403_,
		_w10404_
	);
	LUT2 #(
		.INIT('h1)
	) name9943 (
		_w3320_,
		_w10404_,
		_w10405_
	);
	LUT2 #(
		.INIT('h8)
	) name9944 (
		_w3758_,
		_w9636_,
		_w10406_
	);
	LUT2 #(
		.INIT('h1)
	) name9945 (
		_w10399_,
		_w10406_,
		_w10407_
	);
	LUT2 #(
		.INIT('h1)
	) name9946 (
		_w3177_,
		_w10407_,
		_w10408_
	);
	LUT2 #(
		.INIT('h8)
	) name9947 (
		_w3758_,
		_w9641_,
		_w10409_
	);
	LUT2 #(
		.INIT('h1)
	) name9948 (
		_w10399_,
		_w10409_,
		_w10410_
	);
	LUT2 #(
		.INIT('h2)
	) name9949 (
		_w3355_,
		_w10410_,
		_w10411_
	);
	LUT2 #(
		.INIT('h8)
	) name9950 (
		_w2499_,
		_w3420_,
		_w10412_
	);
	LUT2 #(
		.INIT('h2)
	) name9951 (
		\P2_reg2_reg[6]/NET0131 ,
		_w3774_,
		_w10413_
	);
	LUT2 #(
		.INIT('h1)
	) name9952 (
		_w10398_,
		_w10412_,
		_w10414_
	);
	LUT2 #(
		.INIT('h4)
	) name9953 (
		_w10413_,
		_w10414_,
		_w10415_
	);
	LUT2 #(
		.INIT('h4)
	) name9954 (
		_w10411_,
		_w10415_,
		_w10416_
	);
	LUT2 #(
		.INIT('h4)
	) name9955 (
		_w10405_,
		_w10416_,
		_w10417_
	);
	LUT2 #(
		.INIT('h4)
	) name9956 (
		_w10408_,
		_w10417_,
		_w10418_
	);
	LUT2 #(
		.INIT('h4)
	) name9957 (
		_w10402_,
		_w10418_,
		_w10419_
	);
	LUT2 #(
		.INIT('h2)
	) name9958 (
		_w2026_,
		_w10419_,
		_w10420_
	);
	LUT2 #(
		.INIT('h1)
	) name9959 (
		_w10396_,
		_w10420_,
		_w10421_
	);
	LUT2 #(
		.INIT('h2)
	) name9960 (
		\P1_state_reg[0]/NET0131 ,
		_w10421_,
		_w10422_
	);
	LUT2 #(
		.INIT('h1)
	) name9961 (
		_w10395_,
		_w10422_,
		_w10423_
	);
	LUT2 #(
		.INIT('h8)
	) name9962 (
		\P2_reg2_reg[7]/NET0131 ,
		_w2024_,
		_w10424_
	);
	LUT2 #(
		.INIT('h2)
	) name9963 (
		\P2_reg2_reg[7]/NET0131 ,
		_w3774_,
		_w10425_
	);
	LUT2 #(
		.INIT('h2)
	) name9964 (
		\P2_reg2_reg[7]/NET0131 ,
		_w3758_,
		_w10426_
	);
	LUT2 #(
		.INIT('h8)
	) name9965 (
		_w3758_,
		_w9664_,
		_w10427_
	);
	LUT2 #(
		.INIT('h1)
	) name9966 (
		_w10426_,
		_w10427_,
		_w10428_
	);
	LUT2 #(
		.INIT('h2)
	) name9967 (
		_w3411_,
		_w10428_,
		_w10429_
	);
	LUT2 #(
		.INIT('h8)
	) name9968 (
		_w3758_,
		_w9670_,
		_w10430_
	);
	LUT2 #(
		.INIT('h1)
	) name9969 (
		_w10426_,
		_w10430_,
		_w10431_
	);
	LUT2 #(
		.INIT('h1)
	) name9970 (
		_w3177_,
		_w10431_,
		_w10432_
	);
	LUT2 #(
		.INIT('h2)
	) name9971 (
		_w3758_,
		_w9676_,
		_w10433_
	);
	LUT2 #(
		.INIT('h1)
	) name9972 (
		_w10426_,
		_w10433_,
		_w10434_
	);
	LUT2 #(
		.INIT('h1)
	) name9973 (
		_w3320_,
		_w10434_,
		_w10435_
	);
	LUT2 #(
		.INIT('h8)
	) name9974 (
		_w3758_,
		_w9681_,
		_w10436_
	);
	LUT2 #(
		.INIT('h1)
	) name9975 (
		_w10426_,
		_w10436_,
		_w10437_
	);
	LUT2 #(
		.INIT('h2)
	) name9976 (
		_w3355_,
		_w10437_,
		_w10438_
	);
	LUT2 #(
		.INIT('h8)
	) name9977 (
		_w2476_,
		_w3420_,
		_w10439_
	);
	LUT2 #(
		.INIT('h8)
	) name9978 (
		_w3758_,
		_w10249_,
		_w10440_
	);
	LUT2 #(
		.INIT('h1)
	) name9979 (
		_w10439_,
		_w10440_,
		_w10441_
	);
	LUT2 #(
		.INIT('h4)
	) name9980 (
		_w10425_,
		_w10441_,
		_w10442_
	);
	LUT2 #(
		.INIT('h4)
	) name9981 (
		_w10435_,
		_w10442_,
		_w10443_
	);
	LUT2 #(
		.INIT('h4)
	) name9982 (
		_w10438_,
		_w10443_,
		_w10444_
	);
	LUT2 #(
		.INIT('h4)
	) name9983 (
		_w10432_,
		_w10444_,
		_w10445_
	);
	LUT2 #(
		.INIT('h4)
	) name9984 (
		_w10429_,
		_w10445_,
		_w10446_
	);
	LUT2 #(
		.INIT('h2)
	) name9985 (
		_w2026_,
		_w10446_,
		_w10447_
	);
	LUT2 #(
		.INIT('h1)
	) name9986 (
		_w10424_,
		_w10447_,
		_w10448_
	);
	LUT2 #(
		.INIT('h2)
	) name9987 (
		\P1_state_reg[0]/NET0131 ,
		_w10448_,
		_w10449_
	);
	LUT2 #(
		.INIT('h2)
	) name9988 (
		\P2_reg2_reg[7]/NET0131 ,
		_w1983_,
		_w10450_
	);
	LUT2 #(
		.INIT('h1)
	) name9989 (
		_w10449_,
		_w10450_,
		_w10451_
	);
	LUT2 #(
		.INIT('h2)
	) name9990 (
		\P1_reg0_reg[3]/NET0131 ,
		_w3435_,
		_w10452_
	);
	LUT2 #(
		.INIT('h8)
	) name9991 (
		\P1_reg0_reg[3]/NET0131 ,
		_w3448_,
		_w10453_
	);
	LUT2 #(
		.INIT('h2)
	) name9992 (
		_w4396_,
		_w10176_,
		_w10454_
	);
	LUT2 #(
		.INIT('h2)
	) name9993 (
		\P1_reg0_reg[3]/NET0131 ,
		_w4396_,
		_w10455_
	);
	LUT2 #(
		.INIT('h8)
	) name9994 (
		_w4396_,
		_w9709_,
		_w10456_
	);
	LUT2 #(
		.INIT('h1)
	) name9995 (
		_w10455_,
		_w10456_,
		_w10457_
	);
	LUT2 #(
		.INIT('h2)
	) name9996 (
		_w1936_,
		_w10457_,
		_w10458_
	);
	LUT2 #(
		.INIT('h2)
	) name9997 (
		_w4396_,
		_w9716_,
		_w10459_
	);
	LUT2 #(
		.INIT('h1)
	) name9998 (
		_w10455_,
		_w10459_,
		_w10460_
	);
	LUT2 #(
		.INIT('h1)
	) name9999 (
		_w3563_,
		_w10460_,
		_w10461_
	);
	LUT2 #(
		.INIT('h1)
	) name10000 (
		_w3677_,
		_w4396_,
		_w10462_
	);
	LUT2 #(
		.INIT('h2)
	) name10001 (
		_w4494_,
		_w10462_,
		_w10463_
	);
	LUT2 #(
		.INIT('h2)
	) name10002 (
		\P1_reg0_reg[3]/NET0131 ,
		_w10463_,
		_w10464_
	);
	LUT2 #(
		.INIT('h1)
	) name10003 (
		_w10454_,
		_w10464_,
		_w10465_
	);
	LUT2 #(
		.INIT('h4)
	) name10004 (
		_w10461_,
		_w10465_,
		_w10466_
	);
	LUT2 #(
		.INIT('h4)
	) name10005 (
		_w10458_,
		_w10466_,
		_w10467_
	);
	LUT2 #(
		.INIT('h2)
	) name10006 (
		_w3450_,
		_w10467_,
		_w10468_
	);
	LUT2 #(
		.INIT('h1)
	) name10007 (
		_w10453_,
		_w10468_,
		_w10469_
	);
	LUT2 #(
		.INIT('h2)
	) name10008 (
		\P1_state_reg[0]/NET0131 ,
		_w10469_,
		_w10470_
	);
	LUT2 #(
		.INIT('h1)
	) name10009 (
		_w10452_,
		_w10470_,
		_w10471_
	);
	LUT2 #(
		.INIT('h2)
	) name10010 (
		\P1_reg0_reg[7]/NET0131 ,
		_w3435_,
		_w10472_
	);
	LUT2 #(
		.INIT('h8)
	) name10011 (
		\P1_reg0_reg[7]/NET0131 ,
		_w3448_,
		_w10473_
	);
	LUT2 #(
		.INIT('h2)
	) name10012 (
		\P1_reg0_reg[7]/NET0131 ,
		_w4491_,
		_w10474_
	);
	LUT2 #(
		.INIT('h2)
	) name10013 (
		\P1_reg0_reg[7]/NET0131 ,
		_w4396_,
		_w10475_
	);
	LUT2 #(
		.INIT('h8)
	) name10014 (
		_w4396_,
		_w9794_,
		_w10476_
	);
	LUT2 #(
		.INIT('h1)
	) name10015 (
		_w10475_,
		_w10476_,
		_w10477_
	);
	LUT2 #(
		.INIT('h1)
	) name10016 (
		_w3563_,
		_w10477_,
		_w10478_
	);
	LUT2 #(
		.INIT('h8)
	) name10017 (
		_w4396_,
		_w9802_,
		_w10479_
	);
	LUT2 #(
		.INIT('h1)
	) name10018 (
		_w10475_,
		_w10479_,
		_w10480_
	);
	LUT2 #(
		.INIT('h2)
	) name10019 (
		_w1936_,
		_w10480_,
		_w10481_
	);
	LUT2 #(
		.INIT('h2)
	) name10020 (
		_w4396_,
		_w9788_,
		_w10482_
	);
	LUT2 #(
		.INIT('h1)
	) name10021 (
		_w10475_,
		_w10482_,
		_w10483_
	);
	LUT2 #(
		.INIT('h1)
	) name10022 (
		_w3677_,
		_w10483_,
		_w10484_
	);
	LUT2 #(
		.INIT('h8)
	) name10023 (
		_w4396_,
		_w9807_,
		_w10485_
	);
	LUT2 #(
		.INIT('h1)
	) name10024 (
		_w10475_,
		_w10485_,
		_w10486_
	);
	LUT2 #(
		.INIT('h2)
	) name10025 (
		_w3712_,
		_w10486_,
		_w10487_
	);
	LUT2 #(
		.INIT('h4)
	) name10026 (
		_w1514_,
		_w4396_,
		_w10488_
	);
	LUT2 #(
		.INIT('h1)
	) name10027 (
		_w10475_,
		_w10488_,
		_w10489_
	);
	LUT2 #(
		.INIT('h2)
	) name10028 (
		_w1880_,
		_w10489_,
		_w10490_
	);
	LUT2 #(
		.INIT('h1)
	) name10029 (
		_w10474_,
		_w10490_,
		_w10491_
	);
	LUT2 #(
		.INIT('h4)
	) name10030 (
		_w10487_,
		_w10491_,
		_w10492_
	);
	LUT2 #(
		.INIT('h4)
	) name10031 (
		_w10478_,
		_w10492_,
		_w10493_
	);
	LUT2 #(
		.INIT('h1)
	) name10032 (
		_w10481_,
		_w10484_,
		_w10494_
	);
	LUT2 #(
		.INIT('h8)
	) name10033 (
		_w10493_,
		_w10494_,
		_w10495_
	);
	LUT2 #(
		.INIT('h2)
	) name10034 (
		_w3450_,
		_w10495_,
		_w10496_
	);
	LUT2 #(
		.INIT('h1)
	) name10035 (
		_w10473_,
		_w10496_,
		_w10497_
	);
	LUT2 #(
		.INIT('h2)
	) name10036 (
		\P1_state_reg[0]/NET0131 ,
		_w10497_,
		_w10498_
	);
	LUT2 #(
		.INIT('h1)
	) name10037 (
		_w10472_,
		_w10498_,
		_w10499_
	);
	LUT2 #(
		.INIT('h2)
	) name10038 (
		\P1_reg1_reg[6]/NET0131 ,
		_w3435_,
		_w10500_
	);
	LUT2 #(
		.INIT('h8)
	) name10039 (
		\P1_reg1_reg[6]/NET0131 ,
		_w3448_,
		_w10501_
	);
	LUT2 #(
		.INIT('h8)
	) name10040 (
		_w4532_,
		_w10323_,
		_w10502_
	);
	LUT2 #(
		.INIT('h2)
	) name10041 (
		\P1_reg1_reg[6]/NET0131 ,
		_w4532_,
		_w10503_
	);
	LUT2 #(
		.INIT('h2)
	) name10042 (
		_w4532_,
		_w9749_,
		_w10504_
	);
	LUT2 #(
		.INIT('h1)
	) name10043 (
		_w10503_,
		_w10504_,
		_w10505_
	);
	LUT2 #(
		.INIT('h2)
	) name10044 (
		_w1936_,
		_w10505_,
		_w10506_
	);
	LUT2 #(
		.INIT('h2)
	) name10045 (
		_w4532_,
		_w9761_,
		_w10507_
	);
	LUT2 #(
		.INIT('h1)
	) name10046 (
		_w10503_,
		_w10507_,
		_w10508_
	);
	LUT2 #(
		.INIT('h1)
	) name10047 (
		_w3563_,
		_w10508_,
		_w10509_
	);
	LUT2 #(
		.INIT('h8)
	) name10048 (
		_w4532_,
		_w9755_,
		_w10510_
	);
	LUT2 #(
		.INIT('h1)
	) name10049 (
		_w10503_,
		_w10510_,
		_w10511_
	);
	LUT2 #(
		.INIT('h1)
	) name10050 (
		_w3677_,
		_w10511_,
		_w10512_
	);
	LUT2 #(
		.INIT('h8)
	) name10051 (
		_w4532_,
		_w9766_,
		_w10513_
	);
	LUT2 #(
		.INIT('h1)
	) name10052 (
		_w10503_,
		_w10513_,
		_w10514_
	);
	LUT2 #(
		.INIT('h2)
	) name10053 (
		_w3712_,
		_w10514_,
		_w10515_
	);
	LUT2 #(
		.INIT('h2)
	) name10054 (
		\P1_reg1_reg[6]/NET0131 ,
		_w4541_,
		_w10516_
	);
	LUT2 #(
		.INIT('h1)
	) name10055 (
		_w10502_,
		_w10516_,
		_w10517_
	);
	LUT2 #(
		.INIT('h4)
	) name10056 (
		_w10515_,
		_w10517_,
		_w10518_
	);
	LUT2 #(
		.INIT('h4)
	) name10057 (
		_w10506_,
		_w10518_,
		_w10519_
	);
	LUT2 #(
		.INIT('h1)
	) name10058 (
		_w10509_,
		_w10512_,
		_w10520_
	);
	LUT2 #(
		.INIT('h8)
	) name10059 (
		_w10519_,
		_w10520_,
		_w10521_
	);
	LUT2 #(
		.INIT('h2)
	) name10060 (
		_w3450_,
		_w10521_,
		_w10522_
	);
	LUT2 #(
		.INIT('h1)
	) name10061 (
		_w10501_,
		_w10522_,
		_w10523_
	);
	LUT2 #(
		.INIT('h2)
	) name10062 (
		\P1_state_reg[0]/NET0131 ,
		_w10523_,
		_w10524_
	);
	LUT2 #(
		.INIT('h1)
	) name10063 (
		_w10500_,
		_w10524_,
		_w10525_
	);
	LUT2 #(
		.INIT('h2)
	) name10064 (
		\P2_reg0_reg[6]/NET0131 ,
		_w1983_,
		_w10526_
	);
	LUT2 #(
		.INIT('h8)
	) name10065 (
		\P2_reg0_reg[6]/NET0131 ,
		_w2024_,
		_w10527_
	);
	LUT2 #(
		.INIT('h2)
	) name10066 (
		\P2_reg0_reg[6]/NET0131 ,
		_w3423_,
		_w10528_
	);
	LUT2 #(
		.INIT('h2)
	) name10067 (
		\P2_reg0_reg[6]/NET0131 ,
		_w2040_,
		_w10529_
	);
	LUT2 #(
		.INIT('h8)
	) name10068 (
		_w2040_,
		_w9624_,
		_w10530_
	);
	LUT2 #(
		.INIT('h1)
	) name10069 (
		_w10529_,
		_w10530_,
		_w10531_
	);
	LUT2 #(
		.INIT('h2)
	) name10070 (
		_w3411_,
		_w10531_,
		_w10532_
	);
	LUT2 #(
		.INIT('h8)
	) name10071 (
		_w2040_,
		_w9636_,
		_w10533_
	);
	LUT2 #(
		.INIT('h1)
	) name10072 (
		_w10529_,
		_w10533_,
		_w10534_
	);
	LUT2 #(
		.INIT('h1)
	) name10073 (
		_w3177_,
		_w10534_,
		_w10535_
	);
	LUT2 #(
		.INIT('h2)
	) name10074 (
		_w2040_,
		_w9630_,
		_w10536_
	);
	LUT2 #(
		.INIT('h1)
	) name10075 (
		_w10529_,
		_w10536_,
		_w10537_
	);
	LUT2 #(
		.INIT('h1)
	) name10076 (
		_w3320_,
		_w10537_,
		_w10538_
	);
	LUT2 #(
		.INIT('h8)
	) name10077 (
		_w2040_,
		_w9641_,
		_w10539_
	);
	LUT2 #(
		.INIT('h1)
	) name10078 (
		_w10529_,
		_w10539_,
		_w10540_
	);
	LUT2 #(
		.INIT('h2)
	) name10079 (
		_w3355_,
		_w10540_,
		_w10541_
	);
	LUT2 #(
		.INIT('h8)
	) name10080 (
		_w2040_,
		_w10397_,
		_w10542_
	);
	LUT2 #(
		.INIT('h1)
	) name10081 (
		_w10528_,
		_w10542_,
		_w10543_
	);
	LUT2 #(
		.INIT('h4)
	) name10082 (
		_w10541_,
		_w10543_,
		_w10544_
	);
	LUT2 #(
		.INIT('h4)
	) name10083 (
		_w10535_,
		_w10544_,
		_w10545_
	);
	LUT2 #(
		.INIT('h4)
	) name10084 (
		_w10538_,
		_w10545_,
		_w10546_
	);
	LUT2 #(
		.INIT('h4)
	) name10085 (
		_w10532_,
		_w10546_,
		_w10547_
	);
	LUT2 #(
		.INIT('h2)
	) name10086 (
		_w2026_,
		_w10547_,
		_w10548_
	);
	LUT2 #(
		.INIT('h1)
	) name10087 (
		_w10527_,
		_w10548_,
		_w10549_
	);
	LUT2 #(
		.INIT('h2)
	) name10088 (
		\P1_state_reg[0]/NET0131 ,
		_w10549_,
		_w10550_
	);
	LUT2 #(
		.INIT('h1)
	) name10089 (
		_w10526_,
		_w10550_,
		_w10551_
	);
	LUT2 #(
		.INIT('h2)
	) name10090 (
		\P2_reg1_reg[6]/NET0131 ,
		_w1983_,
		_w10552_
	);
	LUT2 #(
		.INIT('h8)
	) name10091 (
		\P2_reg1_reg[6]/NET0131 ,
		_w2024_,
		_w10553_
	);
	LUT2 #(
		.INIT('h8)
	) name10092 (
		_w3733_,
		_w10397_,
		_w10554_
	);
	LUT2 #(
		.INIT('h2)
	) name10093 (
		\P2_reg1_reg[6]/NET0131 ,
		_w3733_,
		_w10555_
	);
	LUT2 #(
		.INIT('h8)
	) name10094 (
		_w3733_,
		_w9624_,
		_w10556_
	);
	LUT2 #(
		.INIT('h1)
	) name10095 (
		_w10555_,
		_w10556_,
		_w10557_
	);
	LUT2 #(
		.INIT('h2)
	) name10096 (
		_w3411_,
		_w10557_,
		_w10558_
	);
	LUT2 #(
		.INIT('h8)
	) name10097 (
		_w3733_,
		_w9636_,
		_w10559_
	);
	LUT2 #(
		.INIT('h1)
	) name10098 (
		_w10555_,
		_w10559_,
		_w10560_
	);
	LUT2 #(
		.INIT('h1)
	) name10099 (
		_w3177_,
		_w10560_,
		_w10561_
	);
	LUT2 #(
		.INIT('h2)
	) name10100 (
		_w3733_,
		_w9630_,
		_w10562_
	);
	LUT2 #(
		.INIT('h1)
	) name10101 (
		_w10555_,
		_w10562_,
		_w10563_
	);
	LUT2 #(
		.INIT('h1)
	) name10102 (
		_w3320_,
		_w10563_,
		_w10564_
	);
	LUT2 #(
		.INIT('h8)
	) name10103 (
		_w3733_,
		_w9641_,
		_w10565_
	);
	LUT2 #(
		.INIT('h1)
	) name10104 (
		_w10555_,
		_w10565_,
		_w10566_
	);
	LUT2 #(
		.INIT('h2)
	) name10105 (
		_w3355_,
		_w10566_,
		_w10567_
	);
	LUT2 #(
		.INIT('h2)
	) name10106 (
		\P2_reg1_reg[6]/NET0131 ,
		_w3743_,
		_w10568_
	);
	LUT2 #(
		.INIT('h1)
	) name10107 (
		_w10554_,
		_w10568_,
		_w10569_
	);
	LUT2 #(
		.INIT('h4)
	) name10108 (
		_w10567_,
		_w10569_,
		_w10570_
	);
	LUT2 #(
		.INIT('h4)
	) name10109 (
		_w10561_,
		_w10570_,
		_w10571_
	);
	LUT2 #(
		.INIT('h4)
	) name10110 (
		_w10564_,
		_w10571_,
		_w10572_
	);
	LUT2 #(
		.INIT('h4)
	) name10111 (
		_w10558_,
		_w10572_,
		_w10573_
	);
	LUT2 #(
		.INIT('h2)
	) name10112 (
		_w2026_,
		_w10573_,
		_w10574_
	);
	LUT2 #(
		.INIT('h1)
	) name10113 (
		_w10553_,
		_w10574_,
		_w10575_
	);
	LUT2 #(
		.INIT('h2)
	) name10114 (
		\P1_state_reg[0]/NET0131 ,
		_w10575_,
		_w10576_
	);
	LUT2 #(
		.INIT('h1)
	) name10115 (
		_w10552_,
		_w10576_,
		_w10577_
	);
	LUT2 #(
		.INIT('h2)
	) name10116 (
		\P1_reg0_reg[6]/NET0131 ,
		_w3435_,
		_w10578_
	);
	LUT2 #(
		.INIT('h8)
	) name10117 (
		\P1_reg0_reg[6]/NET0131 ,
		_w3448_,
		_w10579_
	);
	LUT2 #(
		.INIT('h8)
	) name10118 (
		_w4396_,
		_w10323_,
		_w10580_
	);
	LUT2 #(
		.INIT('h2)
	) name10119 (
		\P1_reg0_reg[6]/NET0131 ,
		_w4396_,
		_w10581_
	);
	LUT2 #(
		.INIT('h2)
	) name10120 (
		_w4396_,
		_w9761_,
		_w10582_
	);
	LUT2 #(
		.INIT('h1)
	) name10121 (
		_w10581_,
		_w10582_,
		_w10583_
	);
	LUT2 #(
		.INIT('h1)
	) name10122 (
		_w3563_,
		_w10583_,
		_w10584_
	);
	LUT2 #(
		.INIT('h2)
	) name10123 (
		_w4396_,
		_w9749_,
		_w10585_
	);
	LUT2 #(
		.INIT('h1)
	) name10124 (
		_w10581_,
		_w10585_,
		_w10586_
	);
	LUT2 #(
		.INIT('h2)
	) name10125 (
		_w1936_,
		_w10586_,
		_w10587_
	);
	LUT2 #(
		.INIT('h8)
	) name10126 (
		_w4396_,
		_w9755_,
		_w10588_
	);
	LUT2 #(
		.INIT('h1)
	) name10127 (
		_w10581_,
		_w10588_,
		_w10589_
	);
	LUT2 #(
		.INIT('h1)
	) name10128 (
		_w3677_,
		_w10589_,
		_w10590_
	);
	LUT2 #(
		.INIT('h8)
	) name10129 (
		_w4396_,
		_w9766_,
		_w10591_
	);
	LUT2 #(
		.INIT('h1)
	) name10130 (
		_w10581_,
		_w10591_,
		_w10592_
	);
	LUT2 #(
		.INIT('h2)
	) name10131 (
		_w3712_,
		_w10592_,
		_w10593_
	);
	LUT2 #(
		.INIT('h2)
	) name10132 (
		\P1_reg0_reg[6]/NET0131 ,
		_w4493_,
		_w10594_
	);
	LUT2 #(
		.INIT('h1)
	) name10133 (
		_w10580_,
		_w10594_,
		_w10595_
	);
	LUT2 #(
		.INIT('h4)
	) name10134 (
		_w10593_,
		_w10595_,
		_w10596_
	);
	LUT2 #(
		.INIT('h4)
	) name10135 (
		_w10584_,
		_w10596_,
		_w10597_
	);
	LUT2 #(
		.INIT('h1)
	) name10136 (
		_w10587_,
		_w10590_,
		_w10598_
	);
	LUT2 #(
		.INIT('h8)
	) name10137 (
		_w10597_,
		_w10598_,
		_w10599_
	);
	LUT2 #(
		.INIT('h2)
	) name10138 (
		_w3450_,
		_w10599_,
		_w10600_
	);
	LUT2 #(
		.INIT('h1)
	) name10139 (
		_w10579_,
		_w10600_,
		_w10601_
	);
	LUT2 #(
		.INIT('h2)
	) name10140 (
		\P1_state_reg[0]/NET0131 ,
		_w10601_,
		_w10602_
	);
	LUT2 #(
		.INIT('h1)
	) name10141 (
		_w10578_,
		_w10602_,
		_w10603_
	);
	LUT2 #(
		.INIT('h2)
	) name10142 (
		\P2_reg3_reg[2]/NET0131 ,
		_w1983_,
		_w10604_
	);
	LUT2 #(
		.INIT('h8)
	) name10143 (
		\P2_reg3_reg[2]/NET0131 ,
		_w2024_,
		_w10605_
	);
	LUT2 #(
		.INIT('h1)
	) name10144 (
		_w2566_,
		_w3965_,
		_w10606_
	);
	LUT2 #(
		.INIT('h2)
	) name10145 (
		\P2_reg3_reg[2]/NET0131 ,
		_w3788_,
		_w10607_
	);
	LUT2 #(
		.INIT('h4)
	) name10146 (
		_w2607_,
		_w4202_,
		_w10608_
	);
	LUT2 #(
		.INIT('h2)
	) name10147 (
		_w2607_,
		_w4202_,
		_w10609_
	);
	LUT2 #(
		.INIT('h1)
	) name10148 (
		_w10608_,
		_w10609_,
		_w10610_
	);
	LUT2 #(
		.INIT('h2)
	) name10149 (
		_w3788_,
		_w10610_,
		_w10611_
	);
	LUT2 #(
		.INIT('h1)
	) name10150 (
		_w10607_,
		_w10611_,
		_w10612_
	);
	LUT2 #(
		.INIT('h1)
	) name10151 (
		_w3177_,
		_w10612_,
		_w10613_
	);
	LUT2 #(
		.INIT('h2)
	) name10152 (
		_w3819_,
		_w4202_,
		_w10614_
	);
	LUT2 #(
		.INIT('h4)
	) name10153 (
		_w3819_,
		_w4202_,
		_w10615_
	);
	LUT2 #(
		.INIT('h1)
	) name10154 (
		_w10614_,
		_w10615_,
		_w10616_
	);
	LUT2 #(
		.INIT('h2)
	) name10155 (
		_w3788_,
		_w10616_,
		_w10617_
	);
	LUT2 #(
		.INIT('h1)
	) name10156 (
		_w10607_,
		_w10617_,
		_w10618_
	);
	LUT2 #(
		.INIT('h1)
	) name10157 (
		_w3320_,
		_w10618_,
		_w10619_
	);
	LUT2 #(
		.INIT('h2)
	) name10158 (
		_w2616_,
		_w3375_,
		_w10620_
	);
	LUT2 #(
		.INIT('h1)
	) name10159 (
		_w3376_,
		_w10620_,
		_w10621_
	);
	LUT2 #(
		.INIT('h1)
	) name10160 (
		_w2058_,
		_w10621_,
		_w10622_
	);
	LUT2 #(
		.INIT('h8)
	) name10161 (
		_w2058_,
		_w2574_,
		_w10623_
	);
	LUT2 #(
		.INIT('h1)
	) name10162 (
		_w10622_,
		_w10623_,
		_w10624_
	);
	LUT2 #(
		.INIT('h8)
	) name10163 (
		_w3788_,
		_w10624_,
		_w10625_
	);
	LUT2 #(
		.INIT('h1)
	) name10164 (
		_w10607_,
		_w10625_,
		_w10626_
	);
	LUT2 #(
		.INIT('h2)
	) name10165 (
		_w3411_,
		_w10626_,
		_w10627_
	);
	LUT2 #(
		.INIT('h1)
	) name10166 (
		_w2566_,
		_w3326_,
		_w10628_
	);
	LUT2 #(
		.INIT('h1)
	) name10167 (
		_w3327_,
		_w10628_,
		_w10629_
	);
	LUT2 #(
		.INIT('h8)
	) name10168 (
		_w3788_,
		_w10629_,
		_w10630_
	);
	LUT2 #(
		.INIT('h1)
	) name10169 (
		_w10607_,
		_w10630_,
		_w10631_
	);
	LUT2 #(
		.INIT('h2)
	) name10170 (
		_w3355_,
		_w10631_,
		_w10632_
	);
	LUT2 #(
		.INIT('h2)
	) name10171 (
		\P2_reg3_reg[2]/NET0131 ,
		_w3962_,
		_w10633_
	);
	LUT2 #(
		.INIT('h1)
	) name10172 (
		_w10606_,
		_w10633_,
		_w10634_
	);
	LUT2 #(
		.INIT('h4)
	) name10173 (
		_w10632_,
		_w10634_,
		_w10635_
	);
	LUT2 #(
		.INIT('h4)
	) name10174 (
		_w10613_,
		_w10635_,
		_w10636_
	);
	LUT2 #(
		.INIT('h4)
	) name10175 (
		_w10619_,
		_w10636_,
		_w10637_
	);
	LUT2 #(
		.INIT('h4)
	) name10176 (
		_w10627_,
		_w10637_,
		_w10638_
	);
	LUT2 #(
		.INIT('h2)
	) name10177 (
		_w2026_,
		_w10638_,
		_w10639_
	);
	LUT2 #(
		.INIT('h1)
	) name10178 (
		_w10605_,
		_w10639_,
		_w10640_
	);
	LUT2 #(
		.INIT('h2)
	) name10179 (
		\P1_state_reg[0]/NET0131 ,
		_w10640_,
		_w10641_
	);
	LUT2 #(
		.INIT('h1)
	) name10180 (
		_w10604_,
		_w10641_,
		_w10642_
	);
	LUT2 #(
		.INIT('h2)
	) name10181 (
		\P1_reg3_reg[2]/NET0131 ,
		_w3435_,
		_w10643_
	);
	LUT2 #(
		.INIT('h8)
	) name10182 (
		\P1_reg3_reg[2]/NET0131 ,
		_w3448_,
		_w10644_
	);
	LUT2 #(
		.INIT('h1)
	) name10183 (
		_w1609_,
		_w4067_,
		_w10645_
	);
	LUT2 #(
		.INIT('h2)
	) name10184 (
		\P1_reg3_reg[2]/NET0131 ,
		_w3980_,
		_w10646_
	);
	LUT2 #(
		.INIT('h2)
	) name10185 (
		_w1779_,
		_w3507_,
		_w10647_
	);
	LUT2 #(
		.INIT('h4)
	) name10186 (
		_w1779_,
		_w3507_,
		_w10648_
	);
	LUT2 #(
		.INIT('h1)
	) name10187 (
		_w10647_,
		_w10648_,
		_w10649_
	);
	LUT2 #(
		.INIT('h2)
	) name10188 (
		_w3980_,
		_w10649_,
		_w10650_
	);
	LUT2 #(
		.INIT('h1)
	) name10189 (
		_w10646_,
		_w10650_,
		_w10651_
	);
	LUT2 #(
		.INIT('h1)
	) name10190 (
		_w3563_,
		_w10651_,
		_w10652_
	);
	LUT2 #(
		.INIT('h2)
	) name10191 (
		_w1674_,
		_w1779_,
		_w10653_
	);
	LUT2 #(
		.INIT('h4)
	) name10192 (
		_w1674_,
		_w1779_,
		_w10654_
	);
	LUT2 #(
		.INIT('h1)
	) name10193 (
		_w10653_,
		_w10654_,
		_w10655_
	);
	LUT2 #(
		.INIT('h2)
	) name10194 (
		_w3980_,
		_w10655_,
		_w10656_
	);
	LUT2 #(
		.INIT('h1)
	) name10195 (
		_w10646_,
		_w10656_,
		_w10657_
	);
	LUT2 #(
		.INIT('h1)
	) name10196 (
		_w3677_,
		_w10657_,
		_w10658_
	);
	LUT2 #(
		.INIT('h2)
	) name10197 (
		_w1617_,
		_w3572_,
		_w10659_
	);
	LUT2 #(
		.INIT('h1)
	) name10198 (
		_w3573_,
		_w10659_,
		_w10660_
	);
	LUT2 #(
		.INIT('h1)
	) name10199 (
		_w537_,
		_w10660_,
		_w10661_
	);
	LUT2 #(
		.INIT('h8)
	) name10200 (
		_w537_,
		_w1641_,
		_w10662_
	);
	LUT2 #(
		.INIT('h1)
	) name10201 (
		_w10661_,
		_w10662_,
		_w10663_
	);
	LUT2 #(
		.INIT('h8)
	) name10202 (
		_w3980_,
		_w10663_,
		_w10664_
	);
	LUT2 #(
		.INIT('h1)
	) name10203 (
		_w10646_,
		_w10664_,
		_w10665_
	);
	LUT2 #(
		.INIT('h2)
	) name10204 (
		_w1936_,
		_w10665_,
		_w10666_
	);
	LUT2 #(
		.INIT('h1)
	) name10205 (
		_w1609_,
		_w3679_,
		_w10667_
	);
	LUT2 #(
		.INIT('h1)
	) name10206 (
		_w3680_,
		_w10667_,
		_w10668_
	);
	LUT2 #(
		.INIT('h8)
	) name10207 (
		_w3980_,
		_w10668_,
		_w10669_
	);
	LUT2 #(
		.INIT('h1)
	) name10208 (
		_w10646_,
		_w10669_,
		_w10670_
	);
	LUT2 #(
		.INIT('h2)
	) name10209 (
		_w3712_,
		_w10670_,
		_w10671_
	);
	LUT2 #(
		.INIT('h2)
	) name10210 (
		\P1_reg3_reg[2]/NET0131 ,
		_w4064_,
		_w10672_
	);
	LUT2 #(
		.INIT('h1)
	) name10211 (
		_w10645_,
		_w10672_,
		_w10673_
	);
	LUT2 #(
		.INIT('h4)
	) name10212 (
		_w10671_,
		_w10673_,
		_w10674_
	);
	LUT2 #(
		.INIT('h4)
	) name10213 (
		_w10652_,
		_w10674_,
		_w10675_
	);
	LUT2 #(
		.INIT('h4)
	) name10214 (
		_w10658_,
		_w10675_,
		_w10676_
	);
	LUT2 #(
		.INIT('h4)
	) name10215 (
		_w10666_,
		_w10676_,
		_w10677_
	);
	LUT2 #(
		.INIT('h2)
	) name10216 (
		_w3450_,
		_w10677_,
		_w10678_
	);
	LUT2 #(
		.INIT('h1)
	) name10217 (
		_w10644_,
		_w10678_,
		_w10679_
	);
	LUT2 #(
		.INIT('h2)
	) name10218 (
		\P1_state_reg[0]/NET0131 ,
		_w10679_,
		_w10680_
	);
	LUT2 #(
		.INIT('h1)
	) name10219 (
		_w10643_,
		_w10680_,
		_w10681_
	);
	LUT2 #(
		.INIT('h2)
	) name10220 (
		\P2_reg0_reg[2]/NET0131 ,
		_w1983_,
		_w10682_
	);
	LUT2 #(
		.INIT('h8)
	) name10221 (
		\P2_reg0_reg[2]/NET0131 ,
		_w2024_,
		_w10683_
	);
	LUT2 #(
		.INIT('h4)
	) name10222 (
		_w2566_,
		_w3358_,
		_w10684_
	);
	LUT2 #(
		.INIT('h8)
	) name10223 (
		_w2040_,
		_w10684_,
		_w10685_
	);
	LUT2 #(
		.INIT('h2)
	) name10224 (
		\P2_reg0_reg[2]/NET0131 ,
		_w2040_,
		_w10686_
	);
	LUT2 #(
		.INIT('h2)
	) name10225 (
		_w2040_,
		_w10610_,
		_w10687_
	);
	LUT2 #(
		.INIT('h1)
	) name10226 (
		_w10686_,
		_w10687_,
		_w10688_
	);
	LUT2 #(
		.INIT('h1)
	) name10227 (
		_w3177_,
		_w10688_,
		_w10689_
	);
	LUT2 #(
		.INIT('h2)
	) name10228 (
		_w2040_,
		_w10616_,
		_w10690_
	);
	LUT2 #(
		.INIT('h1)
	) name10229 (
		_w10686_,
		_w10690_,
		_w10691_
	);
	LUT2 #(
		.INIT('h1)
	) name10230 (
		_w3320_,
		_w10691_,
		_w10692_
	);
	LUT2 #(
		.INIT('h8)
	) name10231 (
		_w2040_,
		_w10624_,
		_w10693_
	);
	LUT2 #(
		.INIT('h1)
	) name10232 (
		_w10686_,
		_w10693_,
		_w10694_
	);
	LUT2 #(
		.INIT('h2)
	) name10233 (
		_w3411_,
		_w10694_,
		_w10695_
	);
	LUT2 #(
		.INIT('h8)
	) name10234 (
		_w2040_,
		_w10629_,
		_w10696_
	);
	LUT2 #(
		.INIT('h1)
	) name10235 (
		_w10686_,
		_w10696_,
		_w10697_
	);
	LUT2 #(
		.INIT('h2)
	) name10236 (
		_w3355_,
		_w10697_,
		_w10698_
	);
	LUT2 #(
		.INIT('h2)
	) name10237 (
		\P2_reg0_reg[2]/NET0131 ,
		_w3423_,
		_w10699_
	);
	LUT2 #(
		.INIT('h1)
	) name10238 (
		_w10685_,
		_w10699_,
		_w10700_
	);
	LUT2 #(
		.INIT('h4)
	) name10239 (
		_w10698_,
		_w10700_,
		_w10701_
	);
	LUT2 #(
		.INIT('h4)
	) name10240 (
		_w10689_,
		_w10701_,
		_w10702_
	);
	LUT2 #(
		.INIT('h4)
	) name10241 (
		_w10692_,
		_w10702_,
		_w10703_
	);
	LUT2 #(
		.INIT('h4)
	) name10242 (
		_w10695_,
		_w10703_,
		_w10704_
	);
	LUT2 #(
		.INIT('h2)
	) name10243 (
		_w2026_,
		_w10704_,
		_w10705_
	);
	LUT2 #(
		.INIT('h1)
	) name10244 (
		_w10683_,
		_w10705_,
		_w10706_
	);
	LUT2 #(
		.INIT('h2)
	) name10245 (
		\P1_state_reg[0]/NET0131 ,
		_w10706_,
		_w10707_
	);
	LUT2 #(
		.INIT('h1)
	) name10246 (
		_w10682_,
		_w10707_,
		_w10708_
	);
	LUT2 #(
		.INIT('h2)
	) name10247 (
		\P2_reg1_reg[2]/NET0131 ,
		_w1983_,
		_w10709_
	);
	LUT2 #(
		.INIT('h8)
	) name10248 (
		\P2_reg1_reg[2]/NET0131 ,
		_w2024_,
		_w10710_
	);
	LUT2 #(
		.INIT('h8)
	) name10249 (
		_w3733_,
		_w10684_,
		_w10711_
	);
	LUT2 #(
		.INIT('h2)
	) name10250 (
		\P2_reg1_reg[2]/NET0131 ,
		_w3733_,
		_w10712_
	);
	LUT2 #(
		.INIT('h2)
	) name10251 (
		_w3733_,
		_w10616_,
		_w10713_
	);
	LUT2 #(
		.INIT('h1)
	) name10252 (
		_w10712_,
		_w10713_,
		_w10714_
	);
	LUT2 #(
		.INIT('h1)
	) name10253 (
		_w3320_,
		_w10714_,
		_w10715_
	);
	LUT2 #(
		.INIT('h2)
	) name10254 (
		_w3733_,
		_w10610_,
		_w10716_
	);
	LUT2 #(
		.INIT('h1)
	) name10255 (
		_w10712_,
		_w10716_,
		_w10717_
	);
	LUT2 #(
		.INIT('h1)
	) name10256 (
		_w3177_,
		_w10717_,
		_w10718_
	);
	LUT2 #(
		.INIT('h8)
	) name10257 (
		_w3733_,
		_w10624_,
		_w10719_
	);
	LUT2 #(
		.INIT('h1)
	) name10258 (
		_w10712_,
		_w10719_,
		_w10720_
	);
	LUT2 #(
		.INIT('h2)
	) name10259 (
		_w3411_,
		_w10720_,
		_w10721_
	);
	LUT2 #(
		.INIT('h8)
	) name10260 (
		_w3733_,
		_w10629_,
		_w10722_
	);
	LUT2 #(
		.INIT('h1)
	) name10261 (
		_w10712_,
		_w10722_,
		_w10723_
	);
	LUT2 #(
		.INIT('h2)
	) name10262 (
		_w3355_,
		_w10723_,
		_w10724_
	);
	LUT2 #(
		.INIT('h2)
	) name10263 (
		\P2_reg1_reg[2]/NET0131 ,
		_w3743_,
		_w10725_
	);
	LUT2 #(
		.INIT('h1)
	) name10264 (
		_w10711_,
		_w10725_,
		_w10726_
	);
	LUT2 #(
		.INIT('h4)
	) name10265 (
		_w10724_,
		_w10726_,
		_w10727_
	);
	LUT2 #(
		.INIT('h4)
	) name10266 (
		_w10715_,
		_w10727_,
		_w10728_
	);
	LUT2 #(
		.INIT('h4)
	) name10267 (
		_w10718_,
		_w10728_,
		_w10729_
	);
	LUT2 #(
		.INIT('h4)
	) name10268 (
		_w10721_,
		_w10729_,
		_w10730_
	);
	LUT2 #(
		.INIT('h2)
	) name10269 (
		_w2026_,
		_w10730_,
		_w10731_
	);
	LUT2 #(
		.INIT('h1)
	) name10270 (
		_w10710_,
		_w10731_,
		_w10732_
	);
	LUT2 #(
		.INIT('h2)
	) name10271 (
		\P1_state_reg[0]/NET0131 ,
		_w10732_,
		_w10733_
	);
	LUT2 #(
		.INIT('h1)
	) name10272 (
		_w10709_,
		_w10733_,
		_w10734_
	);
	LUT2 #(
		.INIT('h2)
	) name10273 (
		\P1_reg2_reg[2]/NET0131 ,
		_w3435_,
		_w10735_
	);
	LUT2 #(
		.INIT('h8)
	) name10274 (
		\P1_reg2_reg[2]/NET0131 ,
		_w3448_,
		_w10736_
	);
	LUT2 #(
		.INIT('h4)
	) name10275 (
		_w1609_,
		_w1880_,
		_w10737_
	);
	LUT2 #(
		.INIT('h8)
	) name10276 (
		_w3466_,
		_w10737_,
		_w10738_
	);
	LUT2 #(
		.INIT('h2)
	) name10277 (
		\P1_reg2_reg[2]/NET0131 ,
		_w3466_,
		_w10739_
	);
	LUT2 #(
		.INIT('h2)
	) name10278 (
		_w3466_,
		_w10655_,
		_w10740_
	);
	LUT2 #(
		.INIT('h1)
	) name10279 (
		_w10739_,
		_w10740_,
		_w10741_
	);
	LUT2 #(
		.INIT('h1)
	) name10280 (
		_w3677_,
		_w10741_,
		_w10742_
	);
	LUT2 #(
		.INIT('h2)
	) name10281 (
		_w3466_,
		_w10649_,
		_w10743_
	);
	LUT2 #(
		.INIT('h1)
	) name10282 (
		_w10739_,
		_w10743_,
		_w10744_
	);
	LUT2 #(
		.INIT('h1)
	) name10283 (
		_w3563_,
		_w10744_,
		_w10745_
	);
	LUT2 #(
		.INIT('h8)
	) name10284 (
		_w3466_,
		_w10663_,
		_w10746_
	);
	LUT2 #(
		.INIT('h1)
	) name10285 (
		_w10739_,
		_w10746_,
		_w10747_
	);
	LUT2 #(
		.INIT('h2)
	) name10286 (
		_w1936_,
		_w10747_,
		_w10748_
	);
	LUT2 #(
		.INIT('h8)
	) name10287 (
		_w3466_,
		_w10668_,
		_w10749_
	);
	LUT2 #(
		.INIT('h1)
	) name10288 (
		_w10739_,
		_w10749_,
		_w10750_
	);
	LUT2 #(
		.INIT('h2)
	) name10289 (
		_w3712_,
		_w10750_,
		_w10751_
	);
	LUT2 #(
		.INIT('h8)
	) name10290 (
		\P1_reg3_reg[2]/NET0131 ,
		_w1763_,
		_w10752_
	);
	LUT2 #(
		.INIT('h2)
	) name10291 (
		\P1_reg2_reg[2]/NET0131 ,
		_w3718_,
		_w10753_
	);
	LUT2 #(
		.INIT('h1)
	) name10292 (
		_w10738_,
		_w10752_,
		_w10754_
	);
	LUT2 #(
		.INIT('h4)
	) name10293 (
		_w10753_,
		_w10754_,
		_w10755_
	);
	LUT2 #(
		.INIT('h4)
	) name10294 (
		_w10751_,
		_w10755_,
		_w10756_
	);
	LUT2 #(
		.INIT('h4)
	) name10295 (
		_w10742_,
		_w10756_,
		_w10757_
	);
	LUT2 #(
		.INIT('h4)
	) name10296 (
		_w10745_,
		_w10757_,
		_w10758_
	);
	LUT2 #(
		.INIT('h4)
	) name10297 (
		_w10748_,
		_w10758_,
		_w10759_
	);
	LUT2 #(
		.INIT('h2)
	) name10298 (
		_w3450_,
		_w10759_,
		_w10760_
	);
	LUT2 #(
		.INIT('h1)
	) name10299 (
		_w10736_,
		_w10760_,
		_w10761_
	);
	LUT2 #(
		.INIT('h2)
	) name10300 (
		\P1_state_reg[0]/NET0131 ,
		_w10761_,
		_w10762_
	);
	LUT2 #(
		.INIT('h1)
	) name10301 (
		_w10735_,
		_w10762_,
		_w10763_
	);
	LUT2 #(
		.INIT('h2)
	) name10302 (
		\P1_reg0_reg[2]/NET0131 ,
		_w3435_,
		_w10764_
	);
	LUT2 #(
		.INIT('h8)
	) name10303 (
		\P1_reg0_reg[2]/NET0131 ,
		_w3448_,
		_w10765_
	);
	LUT2 #(
		.INIT('h8)
	) name10304 (
		_w4396_,
		_w10737_,
		_w10766_
	);
	LUT2 #(
		.INIT('h2)
	) name10305 (
		\P1_reg0_reg[2]/NET0131 ,
		_w4396_,
		_w10767_
	);
	LUT2 #(
		.INIT('h2)
	) name10306 (
		_w4396_,
		_w10655_,
		_w10768_
	);
	LUT2 #(
		.INIT('h1)
	) name10307 (
		_w10767_,
		_w10768_,
		_w10769_
	);
	LUT2 #(
		.INIT('h1)
	) name10308 (
		_w3677_,
		_w10769_,
		_w10770_
	);
	LUT2 #(
		.INIT('h2)
	) name10309 (
		_w4396_,
		_w10649_,
		_w10771_
	);
	LUT2 #(
		.INIT('h1)
	) name10310 (
		_w10767_,
		_w10771_,
		_w10772_
	);
	LUT2 #(
		.INIT('h1)
	) name10311 (
		_w3563_,
		_w10772_,
		_w10773_
	);
	LUT2 #(
		.INIT('h8)
	) name10312 (
		_w4396_,
		_w10663_,
		_w10774_
	);
	LUT2 #(
		.INIT('h1)
	) name10313 (
		_w10767_,
		_w10774_,
		_w10775_
	);
	LUT2 #(
		.INIT('h2)
	) name10314 (
		_w1936_,
		_w10775_,
		_w10776_
	);
	LUT2 #(
		.INIT('h8)
	) name10315 (
		_w4396_,
		_w10668_,
		_w10777_
	);
	LUT2 #(
		.INIT('h1)
	) name10316 (
		_w10767_,
		_w10777_,
		_w10778_
	);
	LUT2 #(
		.INIT('h2)
	) name10317 (
		_w3712_,
		_w10778_,
		_w10779_
	);
	LUT2 #(
		.INIT('h2)
	) name10318 (
		\P1_reg0_reg[2]/NET0131 ,
		_w4493_,
		_w10780_
	);
	LUT2 #(
		.INIT('h1)
	) name10319 (
		_w10766_,
		_w10780_,
		_w10781_
	);
	LUT2 #(
		.INIT('h4)
	) name10320 (
		_w10779_,
		_w10781_,
		_w10782_
	);
	LUT2 #(
		.INIT('h4)
	) name10321 (
		_w10770_,
		_w10782_,
		_w10783_
	);
	LUT2 #(
		.INIT('h4)
	) name10322 (
		_w10773_,
		_w10783_,
		_w10784_
	);
	LUT2 #(
		.INIT('h4)
	) name10323 (
		_w10776_,
		_w10784_,
		_w10785_
	);
	LUT2 #(
		.INIT('h2)
	) name10324 (
		_w3450_,
		_w10785_,
		_w10786_
	);
	LUT2 #(
		.INIT('h1)
	) name10325 (
		_w10765_,
		_w10786_,
		_w10787_
	);
	LUT2 #(
		.INIT('h2)
	) name10326 (
		\P1_state_reg[0]/NET0131 ,
		_w10787_,
		_w10788_
	);
	LUT2 #(
		.INIT('h1)
	) name10327 (
		_w10764_,
		_w10788_,
		_w10789_
	);
	LUT2 #(
		.INIT('h2)
	) name10328 (
		\P1_reg1_reg[2]/NET0131 ,
		_w3435_,
		_w10790_
	);
	LUT2 #(
		.INIT('h8)
	) name10329 (
		\P1_reg1_reg[2]/NET0131 ,
		_w3448_,
		_w10791_
	);
	LUT2 #(
		.INIT('h8)
	) name10330 (
		_w4532_,
		_w10737_,
		_w10792_
	);
	LUT2 #(
		.INIT('h2)
	) name10331 (
		\P1_reg1_reg[2]/NET0131 ,
		_w4532_,
		_w10793_
	);
	LUT2 #(
		.INIT('h2)
	) name10332 (
		_w4532_,
		_w10655_,
		_w10794_
	);
	LUT2 #(
		.INIT('h1)
	) name10333 (
		_w10793_,
		_w10794_,
		_w10795_
	);
	LUT2 #(
		.INIT('h1)
	) name10334 (
		_w3677_,
		_w10795_,
		_w10796_
	);
	LUT2 #(
		.INIT('h2)
	) name10335 (
		_w4532_,
		_w10649_,
		_w10797_
	);
	LUT2 #(
		.INIT('h1)
	) name10336 (
		_w10793_,
		_w10797_,
		_w10798_
	);
	LUT2 #(
		.INIT('h1)
	) name10337 (
		_w3563_,
		_w10798_,
		_w10799_
	);
	LUT2 #(
		.INIT('h8)
	) name10338 (
		_w4532_,
		_w10663_,
		_w10800_
	);
	LUT2 #(
		.INIT('h1)
	) name10339 (
		_w10793_,
		_w10800_,
		_w10801_
	);
	LUT2 #(
		.INIT('h2)
	) name10340 (
		_w1936_,
		_w10801_,
		_w10802_
	);
	LUT2 #(
		.INIT('h8)
	) name10341 (
		_w4532_,
		_w10668_,
		_w10803_
	);
	LUT2 #(
		.INIT('h1)
	) name10342 (
		_w10793_,
		_w10803_,
		_w10804_
	);
	LUT2 #(
		.INIT('h2)
	) name10343 (
		_w3712_,
		_w10804_,
		_w10805_
	);
	LUT2 #(
		.INIT('h2)
	) name10344 (
		\P1_reg1_reg[2]/NET0131 ,
		_w4541_,
		_w10806_
	);
	LUT2 #(
		.INIT('h1)
	) name10345 (
		_w10792_,
		_w10806_,
		_w10807_
	);
	LUT2 #(
		.INIT('h4)
	) name10346 (
		_w10805_,
		_w10807_,
		_w10808_
	);
	LUT2 #(
		.INIT('h4)
	) name10347 (
		_w10796_,
		_w10808_,
		_w10809_
	);
	LUT2 #(
		.INIT('h4)
	) name10348 (
		_w10799_,
		_w10809_,
		_w10810_
	);
	LUT2 #(
		.INIT('h4)
	) name10349 (
		_w10802_,
		_w10810_,
		_w10811_
	);
	LUT2 #(
		.INIT('h2)
	) name10350 (
		_w3450_,
		_w10811_,
		_w10812_
	);
	LUT2 #(
		.INIT('h1)
	) name10351 (
		_w10791_,
		_w10812_,
		_w10813_
	);
	LUT2 #(
		.INIT('h2)
	) name10352 (
		\P1_state_reg[0]/NET0131 ,
		_w10813_,
		_w10814_
	);
	LUT2 #(
		.INIT('h1)
	) name10353 (
		_w10790_,
		_w10814_,
		_w10815_
	);
	LUT2 #(
		.INIT('h2)
	) name10354 (
		\P1_reg3_reg[1]/NET0131 ,
		_w3435_,
		_w10816_
	);
	LUT2 #(
		.INIT('h8)
	) name10355 (
		\P1_reg3_reg[1]/NET0131 ,
		_w3448_,
		_w10817_
	);
	LUT2 #(
		.INIT('h1)
	) name10356 (
		_w1655_,
		_w1671_,
		_w10818_
	);
	LUT2 #(
		.INIT('h1)
	) name10357 (
		_w3679_,
		_w10818_,
		_w10819_
	);
	LUT2 #(
		.INIT('h8)
	) name10358 (
		_w3712_,
		_w10819_,
		_w10820_
	);
	LUT2 #(
		.INIT('h8)
	) name10359 (
		_w3980_,
		_w10820_,
		_w10821_
	);
	LUT2 #(
		.INIT('h2)
	) name10360 (
		\P1_reg3_reg[1]/NET0131 ,
		_w3980_,
		_w10822_
	);
	LUT2 #(
		.INIT('h8)
	) name10361 (
		_w1792_,
		_w3505_,
		_w10823_
	);
	LUT2 #(
		.INIT('h1)
	) name10362 (
		_w1792_,
		_w3505_,
		_w10824_
	);
	LUT2 #(
		.INIT('h1)
	) name10363 (
		_w10823_,
		_w10824_,
		_w10825_
	);
	LUT2 #(
		.INIT('h4)
	) name10364 (
		_w1671_,
		_w10825_,
		_w10826_
	);
	LUT2 #(
		.INIT('h2)
	) name10365 (
		_w1671_,
		_w1792_,
		_w10827_
	);
	LUT2 #(
		.INIT('h1)
	) name10366 (
		_w10826_,
		_w10827_,
		_w10828_
	);
	LUT2 #(
		.INIT('h2)
	) name10367 (
		_w3980_,
		_w10828_,
		_w10829_
	);
	LUT2 #(
		.INIT('h1)
	) name10368 (
		_w10822_,
		_w10829_,
		_w10830_
	);
	LUT2 #(
		.INIT('h1)
	) name10369 (
		_w3677_,
		_w10830_,
		_w10831_
	);
	LUT2 #(
		.INIT('h2)
	) name10370 (
		_w1595_,
		_w3571_,
		_w10832_
	);
	LUT2 #(
		.INIT('h1)
	) name10371 (
		_w3572_,
		_w10832_,
		_w10833_
	);
	LUT2 #(
		.INIT('h1)
	) name10372 (
		_w537_,
		_w10833_,
		_w10834_
	);
	LUT2 #(
		.INIT('h8)
	) name10373 (
		_w537_,
		_w1664_,
		_w10835_
	);
	LUT2 #(
		.INIT('h1)
	) name10374 (
		_w10834_,
		_w10835_,
		_w10836_
	);
	LUT2 #(
		.INIT('h8)
	) name10375 (
		_w3980_,
		_w10836_,
		_w10837_
	);
	LUT2 #(
		.INIT('h1)
	) name10376 (
		_w10822_,
		_w10837_,
		_w10838_
	);
	LUT2 #(
		.INIT('h2)
	) name10377 (
		_w1936_,
		_w10838_,
		_w10839_
	);
	LUT2 #(
		.INIT('h2)
	) name10378 (
		_w3980_,
		_w10825_,
		_w10840_
	);
	LUT2 #(
		.INIT('h1)
	) name10379 (
		_w10822_,
		_w10840_,
		_w10841_
	);
	LUT2 #(
		.INIT('h1)
	) name10380 (
		_w3563_,
		_w10841_,
		_w10842_
	);
	LUT2 #(
		.INIT('h1)
	) name10381 (
		_w1655_,
		_w4067_,
		_w10843_
	);
	LUT2 #(
		.INIT('h2)
	) name10382 (
		\P1_reg3_reg[1]/NET0131 ,
		_w4910_,
		_w10844_
	);
	LUT2 #(
		.INIT('h1)
	) name10383 (
		_w10821_,
		_w10843_,
		_w10845_
	);
	LUT2 #(
		.INIT('h4)
	) name10384 (
		_w10844_,
		_w10845_,
		_w10846_
	);
	LUT2 #(
		.INIT('h4)
	) name10385 (
		_w10842_,
		_w10846_,
		_w10847_
	);
	LUT2 #(
		.INIT('h4)
	) name10386 (
		_w10831_,
		_w10847_,
		_w10848_
	);
	LUT2 #(
		.INIT('h4)
	) name10387 (
		_w10839_,
		_w10848_,
		_w10849_
	);
	LUT2 #(
		.INIT('h2)
	) name10388 (
		_w3450_,
		_w10849_,
		_w10850_
	);
	LUT2 #(
		.INIT('h1)
	) name10389 (
		_w10817_,
		_w10850_,
		_w10851_
	);
	LUT2 #(
		.INIT('h2)
	) name10390 (
		\P1_state_reg[0]/NET0131 ,
		_w10851_,
		_w10852_
	);
	LUT2 #(
		.INIT('h1)
	) name10391 (
		_w10816_,
		_w10852_,
		_w10853_
	);
	LUT2 #(
		.INIT('h2)
	) name10392 (
		\P2_reg3_reg[1]/NET0131 ,
		_w1983_,
		_w10854_
	);
	LUT2 #(
		.INIT('h8)
	) name10393 (
		\P2_reg3_reg[1]/NET0131 ,
		_w2024_,
		_w10855_
	);
	LUT2 #(
		.INIT('h2)
	) name10394 (
		\P2_reg3_reg[1]/NET0131 ,
		_w5698_,
		_w10856_
	);
	LUT2 #(
		.INIT('h2)
	) name10395 (
		\P2_reg3_reg[1]/NET0131 ,
		_w3788_,
		_w10857_
	);
	LUT2 #(
		.INIT('h4)
	) name10396 (
		_w2605_,
		_w4199_,
		_w10858_
	);
	LUT2 #(
		.INIT('h2)
	) name10397 (
		_w2605_,
		_w4199_,
		_w10859_
	);
	LUT2 #(
		.INIT('h1)
	) name10398 (
		_w10858_,
		_w10859_,
		_w10860_
	);
	LUT2 #(
		.INIT('h1)
	) name10399 (
		_w2604_,
		_w10860_,
		_w10861_
	);
	LUT2 #(
		.INIT('h2)
	) name10400 (
		_w2604_,
		_w4199_,
		_w10862_
	);
	LUT2 #(
		.INIT('h1)
	) name10401 (
		_w10861_,
		_w10862_,
		_w10863_
	);
	LUT2 #(
		.INIT('h2)
	) name10402 (
		_w3788_,
		_w10863_,
		_w10864_
	);
	LUT2 #(
		.INIT('h1)
	) name10403 (
		_w10857_,
		_w10864_,
		_w10865_
	);
	LUT2 #(
		.INIT('h1)
	) name10404 (
		_w3320_,
		_w10865_,
		_w10866_
	);
	LUT2 #(
		.INIT('h2)
	) name10405 (
		_w2552_,
		_w3374_,
		_w10867_
	);
	LUT2 #(
		.INIT('h1)
	) name10406 (
		_w3375_,
		_w10867_,
		_w10868_
	);
	LUT2 #(
		.INIT('h1)
	) name10407 (
		_w2058_,
		_w10868_,
		_w10869_
	);
	LUT2 #(
		.INIT('h8)
	) name10408 (
		_w2058_,
		_w2597_,
		_w10870_
	);
	LUT2 #(
		.INIT('h1)
	) name10409 (
		_w10869_,
		_w10870_,
		_w10871_
	);
	LUT2 #(
		.INIT('h8)
	) name10410 (
		_w3788_,
		_w10871_,
		_w10872_
	);
	LUT2 #(
		.INIT('h1)
	) name10411 (
		_w10857_,
		_w10872_,
		_w10873_
	);
	LUT2 #(
		.INIT('h2)
	) name10412 (
		_w3411_,
		_w10873_,
		_w10874_
	);
	LUT2 #(
		.INIT('h8)
	) name10413 (
		_w3788_,
		_w10860_,
		_w10875_
	);
	LUT2 #(
		.INIT('h1)
	) name10414 (
		_w10857_,
		_w10875_,
		_w10876_
	);
	LUT2 #(
		.INIT('h1)
	) name10415 (
		_w3177_,
		_w10876_,
		_w10877_
	);
	LUT2 #(
		.INIT('h1)
	) name10416 (
		_w2588_,
		_w3965_,
		_w10878_
	);
	LUT2 #(
		.INIT('h1)
	) name10417 (
		_w2588_,
		_w2604_,
		_w10879_
	);
	LUT2 #(
		.INIT('h4)
	) name10418 (
		_w3326_,
		_w3355_,
		_w10880_
	);
	LUT2 #(
		.INIT('h4)
	) name10419 (
		_w10879_,
		_w10880_,
		_w10881_
	);
	LUT2 #(
		.INIT('h8)
	) name10420 (
		_w3788_,
		_w10881_,
		_w10882_
	);
	LUT2 #(
		.INIT('h1)
	) name10421 (
		_w10878_,
		_w10882_,
		_w10883_
	);
	LUT2 #(
		.INIT('h4)
	) name10422 (
		_w10856_,
		_w10883_,
		_w10884_
	);
	LUT2 #(
		.INIT('h4)
	) name10423 (
		_w10877_,
		_w10884_,
		_w10885_
	);
	LUT2 #(
		.INIT('h4)
	) name10424 (
		_w10866_,
		_w10885_,
		_w10886_
	);
	LUT2 #(
		.INIT('h4)
	) name10425 (
		_w10874_,
		_w10886_,
		_w10887_
	);
	LUT2 #(
		.INIT('h2)
	) name10426 (
		_w2026_,
		_w10887_,
		_w10888_
	);
	LUT2 #(
		.INIT('h1)
	) name10427 (
		_w10855_,
		_w10888_,
		_w10889_
	);
	LUT2 #(
		.INIT('h2)
	) name10428 (
		\P1_state_reg[0]/NET0131 ,
		_w10889_,
		_w10890_
	);
	LUT2 #(
		.INIT('h1)
	) name10429 (
		_w10854_,
		_w10890_,
		_w10891_
	);
	LUT2 #(
		.INIT('h2)
	) name10430 (
		\P2_reg0_reg[1]/NET0131 ,
		_w1983_,
		_w10892_
	);
	LUT2 #(
		.INIT('h8)
	) name10431 (
		\P2_reg0_reg[1]/NET0131 ,
		_w2024_,
		_w10893_
	);
	LUT2 #(
		.INIT('h4)
	) name10432 (
		_w2588_,
		_w3358_,
		_w10894_
	);
	LUT2 #(
		.INIT('h1)
	) name10433 (
		_w10881_,
		_w10894_,
		_w10895_
	);
	LUT2 #(
		.INIT('h2)
	) name10434 (
		_w2040_,
		_w10895_,
		_w10896_
	);
	LUT2 #(
		.INIT('h2)
	) name10435 (
		\P2_reg0_reg[1]/NET0131 ,
		_w2040_,
		_w10897_
	);
	LUT2 #(
		.INIT('h2)
	) name10436 (
		_w2040_,
		_w10863_,
		_w10898_
	);
	LUT2 #(
		.INIT('h1)
	) name10437 (
		_w10897_,
		_w10898_,
		_w10899_
	);
	LUT2 #(
		.INIT('h1)
	) name10438 (
		_w3320_,
		_w10899_,
		_w10900_
	);
	LUT2 #(
		.INIT('h8)
	) name10439 (
		_w2040_,
		_w10871_,
		_w10901_
	);
	LUT2 #(
		.INIT('h1)
	) name10440 (
		_w10897_,
		_w10901_,
		_w10902_
	);
	LUT2 #(
		.INIT('h2)
	) name10441 (
		_w3411_,
		_w10902_,
		_w10903_
	);
	LUT2 #(
		.INIT('h8)
	) name10442 (
		_w2040_,
		_w10860_,
		_w10904_
	);
	LUT2 #(
		.INIT('h1)
	) name10443 (
		_w10897_,
		_w10904_,
		_w10905_
	);
	LUT2 #(
		.INIT('h1)
	) name10444 (
		_w3177_,
		_w10905_,
		_w10906_
	);
	LUT2 #(
		.INIT('h2)
	) name10445 (
		\P2_reg0_reg[1]/NET0131 ,
		_w3425_,
		_w10907_
	);
	LUT2 #(
		.INIT('h1)
	) name10446 (
		_w10896_,
		_w10907_,
		_w10908_
	);
	LUT2 #(
		.INIT('h4)
	) name10447 (
		_w10906_,
		_w10908_,
		_w10909_
	);
	LUT2 #(
		.INIT('h4)
	) name10448 (
		_w10900_,
		_w10909_,
		_w10910_
	);
	LUT2 #(
		.INIT('h4)
	) name10449 (
		_w10903_,
		_w10910_,
		_w10911_
	);
	LUT2 #(
		.INIT('h2)
	) name10450 (
		_w2026_,
		_w10911_,
		_w10912_
	);
	LUT2 #(
		.INIT('h1)
	) name10451 (
		_w10893_,
		_w10912_,
		_w10913_
	);
	LUT2 #(
		.INIT('h2)
	) name10452 (
		\P1_state_reg[0]/NET0131 ,
		_w10913_,
		_w10914_
	);
	LUT2 #(
		.INIT('h1)
	) name10453 (
		_w10892_,
		_w10914_,
		_w10915_
	);
	LUT2 #(
		.INIT('h2)
	) name10454 (
		\P2_reg1_reg[1]/NET0131 ,
		_w1983_,
		_w10916_
	);
	LUT2 #(
		.INIT('h8)
	) name10455 (
		\P2_reg1_reg[1]/NET0131 ,
		_w2024_,
		_w10917_
	);
	LUT2 #(
		.INIT('h2)
	) name10456 (
		_w3733_,
		_w10895_,
		_w10918_
	);
	LUT2 #(
		.INIT('h2)
	) name10457 (
		\P2_reg1_reg[1]/NET0131 ,
		_w3733_,
		_w10919_
	);
	LUT2 #(
		.INIT('h2)
	) name10458 (
		_w3733_,
		_w10863_,
		_w10920_
	);
	LUT2 #(
		.INIT('h1)
	) name10459 (
		_w10919_,
		_w10920_,
		_w10921_
	);
	LUT2 #(
		.INIT('h1)
	) name10460 (
		_w3320_,
		_w10921_,
		_w10922_
	);
	LUT2 #(
		.INIT('h8)
	) name10461 (
		_w3733_,
		_w10871_,
		_w10923_
	);
	LUT2 #(
		.INIT('h1)
	) name10462 (
		_w10919_,
		_w10923_,
		_w10924_
	);
	LUT2 #(
		.INIT('h2)
	) name10463 (
		_w3411_,
		_w10924_,
		_w10925_
	);
	LUT2 #(
		.INIT('h8)
	) name10464 (
		_w3733_,
		_w10860_,
		_w10926_
	);
	LUT2 #(
		.INIT('h1)
	) name10465 (
		_w10919_,
		_w10926_,
		_w10927_
	);
	LUT2 #(
		.INIT('h1)
	) name10466 (
		_w3177_,
		_w10927_,
		_w10928_
	);
	LUT2 #(
		.INIT('h2)
	) name10467 (
		\P2_reg1_reg[1]/NET0131 ,
		_w7598_,
		_w10929_
	);
	LUT2 #(
		.INIT('h1)
	) name10468 (
		_w10918_,
		_w10929_,
		_w10930_
	);
	LUT2 #(
		.INIT('h4)
	) name10469 (
		_w10928_,
		_w10930_,
		_w10931_
	);
	LUT2 #(
		.INIT('h4)
	) name10470 (
		_w10922_,
		_w10931_,
		_w10932_
	);
	LUT2 #(
		.INIT('h4)
	) name10471 (
		_w10925_,
		_w10932_,
		_w10933_
	);
	LUT2 #(
		.INIT('h2)
	) name10472 (
		_w2026_,
		_w10933_,
		_w10934_
	);
	LUT2 #(
		.INIT('h1)
	) name10473 (
		_w10917_,
		_w10934_,
		_w10935_
	);
	LUT2 #(
		.INIT('h2)
	) name10474 (
		\P1_state_reg[0]/NET0131 ,
		_w10935_,
		_w10936_
	);
	LUT2 #(
		.INIT('h1)
	) name10475 (
		_w10916_,
		_w10936_,
		_w10937_
	);
	LUT2 #(
		.INIT('h2)
	) name10476 (
		\P2_reg2_reg[2]/NET0131 ,
		_w1983_,
		_w10938_
	);
	LUT2 #(
		.INIT('h8)
	) name10477 (
		\P2_reg2_reg[2]/NET0131 ,
		_w2024_,
		_w10939_
	);
	LUT2 #(
		.INIT('h8)
	) name10478 (
		_w3758_,
		_w10684_,
		_w10940_
	);
	LUT2 #(
		.INIT('h2)
	) name10479 (
		\P2_reg2_reg[2]/NET0131 ,
		_w3758_,
		_w10941_
	);
	LUT2 #(
		.INIT('h2)
	) name10480 (
		_w3758_,
		_w10616_,
		_w10942_
	);
	LUT2 #(
		.INIT('h1)
	) name10481 (
		_w10941_,
		_w10942_,
		_w10943_
	);
	LUT2 #(
		.INIT('h1)
	) name10482 (
		_w3320_,
		_w10943_,
		_w10944_
	);
	LUT2 #(
		.INIT('h2)
	) name10483 (
		_w3758_,
		_w10610_,
		_w10945_
	);
	LUT2 #(
		.INIT('h1)
	) name10484 (
		_w10941_,
		_w10945_,
		_w10946_
	);
	LUT2 #(
		.INIT('h1)
	) name10485 (
		_w3177_,
		_w10946_,
		_w10947_
	);
	LUT2 #(
		.INIT('h8)
	) name10486 (
		_w3758_,
		_w10624_,
		_w10948_
	);
	LUT2 #(
		.INIT('h1)
	) name10487 (
		_w10941_,
		_w10948_,
		_w10949_
	);
	LUT2 #(
		.INIT('h2)
	) name10488 (
		_w3411_,
		_w10949_,
		_w10950_
	);
	LUT2 #(
		.INIT('h8)
	) name10489 (
		_w3758_,
		_w10629_,
		_w10951_
	);
	LUT2 #(
		.INIT('h1)
	) name10490 (
		_w10941_,
		_w10951_,
		_w10952_
	);
	LUT2 #(
		.INIT('h2)
	) name10491 (
		_w3355_,
		_w10952_,
		_w10953_
	);
	LUT2 #(
		.INIT('h8)
	) name10492 (
		\P2_reg3_reg[2]/NET0131 ,
		_w3420_,
		_w10954_
	);
	LUT2 #(
		.INIT('h2)
	) name10493 (
		\P2_reg2_reg[2]/NET0131 ,
		_w3774_,
		_w10955_
	);
	LUT2 #(
		.INIT('h1)
	) name10494 (
		_w10940_,
		_w10954_,
		_w10956_
	);
	LUT2 #(
		.INIT('h4)
	) name10495 (
		_w10955_,
		_w10956_,
		_w10957_
	);
	LUT2 #(
		.INIT('h4)
	) name10496 (
		_w10953_,
		_w10957_,
		_w10958_
	);
	LUT2 #(
		.INIT('h4)
	) name10497 (
		_w10944_,
		_w10958_,
		_w10959_
	);
	LUT2 #(
		.INIT('h4)
	) name10498 (
		_w10947_,
		_w10959_,
		_w10960_
	);
	LUT2 #(
		.INIT('h4)
	) name10499 (
		_w10950_,
		_w10960_,
		_w10961_
	);
	LUT2 #(
		.INIT('h2)
	) name10500 (
		_w2026_,
		_w10961_,
		_w10962_
	);
	LUT2 #(
		.INIT('h1)
	) name10501 (
		_w10939_,
		_w10962_,
		_w10963_
	);
	LUT2 #(
		.INIT('h2)
	) name10502 (
		\P1_state_reg[0]/NET0131 ,
		_w10963_,
		_w10964_
	);
	LUT2 #(
		.INIT('h1)
	) name10503 (
		_w10938_,
		_w10964_,
		_w10965_
	);
	LUT2 #(
		.INIT('h2)
	) name10504 (
		\P1_reg0_reg[1]/NET0131 ,
		_w3435_,
		_w10966_
	);
	LUT2 #(
		.INIT('h8)
	) name10505 (
		\P1_reg0_reg[1]/NET0131 ,
		_w3448_,
		_w10967_
	);
	LUT2 #(
		.INIT('h2)
	) name10506 (
		\P1_reg0_reg[1]/NET0131 ,
		_w4494_,
		_w10968_
	);
	LUT2 #(
		.INIT('h2)
	) name10507 (
		\P1_reg0_reg[1]/NET0131 ,
		_w4396_,
		_w10969_
	);
	LUT2 #(
		.INIT('h2)
	) name10508 (
		_w4396_,
		_w10828_,
		_w10970_
	);
	LUT2 #(
		.INIT('h1)
	) name10509 (
		_w10969_,
		_w10970_,
		_w10971_
	);
	LUT2 #(
		.INIT('h1)
	) name10510 (
		_w3677_,
		_w10971_,
		_w10972_
	);
	LUT2 #(
		.INIT('h8)
	) name10511 (
		_w4396_,
		_w10836_,
		_w10973_
	);
	LUT2 #(
		.INIT('h1)
	) name10512 (
		_w10969_,
		_w10973_,
		_w10974_
	);
	LUT2 #(
		.INIT('h2)
	) name10513 (
		_w1936_,
		_w10974_,
		_w10975_
	);
	LUT2 #(
		.INIT('h2)
	) name10514 (
		_w4396_,
		_w10825_,
		_w10976_
	);
	LUT2 #(
		.INIT('h1)
	) name10515 (
		_w10969_,
		_w10976_,
		_w10977_
	);
	LUT2 #(
		.INIT('h1)
	) name10516 (
		_w3563_,
		_w10977_,
		_w10978_
	);
	LUT2 #(
		.INIT('h4)
	) name10517 (
		_w1655_,
		_w1880_,
		_w10979_
	);
	LUT2 #(
		.INIT('h1)
	) name10518 (
		_w10820_,
		_w10979_,
		_w10980_
	);
	LUT2 #(
		.INIT('h2)
	) name10519 (
		_w4396_,
		_w10980_,
		_w10981_
	);
	LUT2 #(
		.INIT('h1)
	) name10520 (
		_w10968_,
		_w10981_,
		_w10982_
	);
	LUT2 #(
		.INIT('h4)
	) name10521 (
		_w10978_,
		_w10982_,
		_w10983_
	);
	LUT2 #(
		.INIT('h4)
	) name10522 (
		_w10972_,
		_w10983_,
		_w10984_
	);
	LUT2 #(
		.INIT('h4)
	) name10523 (
		_w10975_,
		_w10984_,
		_w10985_
	);
	LUT2 #(
		.INIT('h2)
	) name10524 (
		_w3450_,
		_w10985_,
		_w10986_
	);
	LUT2 #(
		.INIT('h1)
	) name10525 (
		_w10967_,
		_w10986_,
		_w10987_
	);
	LUT2 #(
		.INIT('h2)
	) name10526 (
		\P1_state_reg[0]/NET0131 ,
		_w10987_,
		_w10988_
	);
	LUT2 #(
		.INIT('h1)
	) name10527 (
		_w10966_,
		_w10988_,
		_w10989_
	);
	LUT2 #(
		.INIT('h2)
	) name10528 (
		\P1_reg1_reg[1]/NET0131 ,
		_w3435_,
		_w10990_
	);
	LUT2 #(
		.INIT('h8)
	) name10529 (
		\P1_reg1_reg[1]/NET0131 ,
		_w3448_,
		_w10991_
	);
	LUT2 #(
		.INIT('h2)
	) name10530 (
		\P1_reg1_reg[1]/NET0131 ,
		_w4573_,
		_w10992_
	);
	LUT2 #(
		.INIT('h2)
	) name10531 (
		\P1_reg1_reg[1]/NET0131 ,
		_w4532_,
		_w10993_
	);
	LUT2 #(
		.INIT('h2)
	) name10532 (
		_w4532_,
		_w10828_,
		_w10994_
	);
	LUT2 #(
		.INIT('h1)
	) name10533 (
		_w10993_,
		_w10994_,
		_w10995_
	);
	LUT2 #(
		.INIT('h1)
	) name10534 (
		_w3677_,
		_w10995_,
		_w10996_
	);
	LUT2 #(
		.INIT('h8)
	) name10535 (
		_w4532_,
		_w10836_,
		_w10997_
	);
	LUT2 #(
		.INIT('h1)
	) name10536 (
		_w10993_,
		_w10997_,
		_w10998_
	);
	LUT2 #(
		.INIT('h2)
	) name10537 (
		_w1936_,
		_w10998_,
		_w10999_
	);
	LUT2 #(
		.INIT('h2)
	) name10538 (
		_w4532_,
		_w10825_,
		_w11000_
	);
	LUT2 #(
		.INIT('h1)
	) name10539 (
		_w10993_,
		_w11000_,
		_w11001_
	);
	LUT2 #(
		.INIT('h1)
	) name10540 (
		_w3563_,
		_w11001_,
		_w11002_
	);
	LUT2 #(
		.INIT('h2)
	) name10541 (
		_w4532_,
		_w10980_,
		_w11003_
	);
	LUT2 #(
		.INIT('h1)
	) name10542 (
		_w10992_,
		_w11003_,
		_w11004_
	);
	LUT2 #(
		.INIT('h4)
	) name10543 (
		_w11002_,
		_w11004_,
		_w11005_
	);
	LUT2 #(
		.INIT('h4)
	) name10544 (
		_w10996_,
		_w11005_,
		_w11006_
	);
	LUT2 #(
		.INIT('h4)
	) name10545 (
		_w10999_,
		_w11006_,
		_w11007_
	);
	LUT2 #(
		.INIT('h2)
	) name10546 (
		_w3450_,
		_w11007_,
		_w11008_
	);
	LUT2 #(
		.INIT('h1)
	) name10547 (
		_w10991_,
		_w11008_,
		_w11009_
	);
	LUT2 #(
		.INIT('h2)
	) name10548 (
		\P1_state_reg[0]/NET0131 ,
		_w11009_,
		_w11010_
	);
	LUT2 #(
		.INIT('h1)
	) name10549 (
		_w10990_,
		_w11010_,
		_w11011_
	);
	LUT2 #(
		.INIT('h2)
	) name10550 (
		\P1_reg2_reg[1]/NET0131 ,
		_w3435_,
		_w11012_
	);
	LUT2 #(
		.INIT('h8)
	) name10551 (
		\P1_reg2_reg[1]/NET0131 ,
		_w3448_,
		_w11013_
	);
	LUT2 #(
		.INIT('h8)
	) name10552 (
		\P1_reg3_reg[1]/NET0131 ,
		_w1763_,
		_w11014_
	);
	LUT2 #(
		.INIT('h2)
	) name10553 (
		\P1_reg2_reg[1]/NET0131 ,
		_w3466_,
		_w11015_
	);
	LUT2 #(
		.INIT('h2)
	) name10554 (
		_w3466_,
		_w10828_,
		_w11016_
	);
	LUT2 #(
		.INIT('h1)
	) name10555 (
		_w11015_,
		_w11016_,
		_w11017_
	);
	LUT2 #(
		.INIT('h1)
	) name10556 (
		_w3677_,
		_w11017_,
		_w11018_
	);
	LUT2 #(
		.INIT('h8)
	) name10557 (
		_w3466_,
		_w10836_,
		_w11019_
	);
	LUT2 #(
		.INIT('h1)
	) name10558 (
		_w11015_,
		_w11019_,
		_w11020_
	);
	LUT2 #(
		.INIT('h2)
	) name10559 (
		_w1936_,
		_w11020_,
		_w11021_
	);
	LUT2 #(
		.INIT('h2)
	) name10560 (
		_w3466_,
		_w10825_,
		_w11022_
	);
	LUT2 #(
		.INIT('h1)
	) name10561 (
		_w11015_,
		_w11022_,
		_w11023_
	);
	LUT2 #(
		.INIT('h1)
	) name10562 (
		_w3563_,
		_w11023_,
		_w11024_
	);
	LUT2 #(
		.INIT('h4)
	) name10563 (
		_w1655_,
		_w3466_,
		_w11025_
	);
	LUT2 #(
		.INIT('h1)
	) name10564 (
		_w11015_,
		_w11025_,
		_w11026_
	);
	LUT2 #(
		.INIT('h2)
	) name10565 (
		_w1880_,
		_w11026_,
		_w11027_
	);
	LUT2 #(
		.INIT('h8)
	) name10566 (
		_w3466_,
		_w10819_,
		_w11028_
	);
	LUT2 #(
		.INIT('h1)
	) name10567 (
		_w11015_,
		_w11028_,
		_w11029_
	);
	LUT2 #(
		.INIT('h2)
	) name10568 (
		_w3712_,
		_w11029_,
		_w11030_
	);
	LUT2 #(
		.INIT('h8)
	) name10569 (
		\P1_reg2_reg[1]/NET0131 ,
		_w3716_,
		_w11031_
	);
	LUT2 #(
		.INIT('h1)
	) name10570 (
		_w11014_,
		_w11031_,
		_w11032_
	);
	LUT2 #(
		.INIT('h4)
	) name10571 (
		_w11027_,
		_w11032_,
		_w11033_
	);
	LUT2 #(
		.INIT('h4)
	) name10572 (
		_w11030_,
		_w11033_,
		_w11034_
	);
	LUT2 #(
		.INIT('h4)
	) name10573 (
		_w11024_,
		_w11034_,
		_w11035_
	);
	LUT2 #(
		.INIT('h4)
	) name10574 (
		_w11018_,
		_w11035_,
		_w11036_
	);
	LUT2 #(
		.INIT('h4)
	) name10575 (
		_w11021_,
		_w11036_,
		_w11037_
	);
	LUT2 #(
		.INIT('h2)
	) name10576 (
		_w3450_,
		_w11037_,
		_w11038_
	);
	LUT2 #(
		.INIT('h1)
	) name10577 (
		_w11013_,
		_w11038_,
		_w11039_
	);
	LUT2 #(
		.INIT('h2)
	) name10578 (
		\P1_state_reg[0]/NET0131 ,
		_w11039_,
		_w11040_
	);
	LUT2 #(
		.INIT('h1)
	) name10579 (
		_w11012_,
		_w11040_,
		_w11041_
	);
	LUT2 #(
		.INIT('h2)
	) name10580 (
		\P2_reg2_reg[1]/NET0131 ,
		_w1983_,
		_w11042_
	);
	LUT2 #(
		.INIT('h8)
	) name10581 (
		\P2_reg2_reg[1]/NET0131 ,
		_w2024_,
		_w11043_
	);
	LUT2 #(
		.INIT('h8)
	) name10582 (
		\P2_reg3_reg[1]/NET0131 ,
		_w3420_,
		_w11044_
	);
	LUT2 #(
		.INIT('h2)
	) name10583 (
		\P2_reg2_reg[1]/NET0131 ,
		_w3758_,
		_w11045_
	);
	LUT2 #(
		.INIT('h2)
	) name10584 (
		_w3758_,
		_w10863_,
		_w11046_
	);
	LUT2 #(
		.INIT('h1)
	) name10585 (
		_w11045_,
		_w11046_,
		_w11047_
	);
	LUT2 #(
		.INIT('h1)
	) name10586 (
		_w3320_,
		_w11047_,
		_w11048_
	);
	LUT2 #(
		.INIT('h8)
	) name10587 (
		_w3758_,
		_w10871_,
		_w11049_
	);
	LUT2 #(
		.INIT('h1)
	) name10588 (
		_w11045_,
		_w11049_,
		_w11050_
	);
	LUT2 #(
		.INIT('h2)
	) name10589 (
		_w3411_,
		_w11050_,
		_w11051_
	);
	LUT2 #(
		.INIT('h8)
	) name10590 (
		_w3758_,
		_w10860_,
		_w11052_
	);
	LUT2 #(
		.INIT('h1)
	) name10591 (
		_w11045_,
		_w11052_,
		_w11053_
	);
	LUT2 #(
		.INIT('h1)
	) name10592 (
		_w3177_,
		_w11053_,
		_w11054_
	);
	LUT2 #(
		.INIT('h2)
	) name10593 (
		\P2_reg2_reg[1]/NET0131 ,
		_w4383_,
		_w11055_
	);
	LUT2 #(
		.INIT('h2)
	) name10594 (
		_w3758_,
		_w10895_,
		_w11056_
	);
	LUT2 #(
		.INIT('h1)
	) name10595 (
		_w11044_,
		_w11056_,
		_w11057_
	);
	LUT2 #(
		.INIT('h4)
	) name10596 (
		_w11055_,
		_w11057_,
		_w11058_
	);
	LUT2 #(
		.INIT('h4)
	) name10597 (
		_w11054_,
		_w11058_,
		_w11059_
	);
	LUT2 #(
		.INIT('h4)
	) name10598 (
		_w11048_,
		_w11059_,
		_w11060_
	);
	LUT2 #(
		.INIT('h4)
	) name10599 (
		_w11051_,
		_w11060_,
		_w11061_
	);
	LUT2 #(
		.INIT('h2)
	) name10600 (
		_w2026_,
		_w11061_,
		_w11062_
	);
	LUT2 #(
		.INIT('h1)
	) name10601 (
		_w11043_,
		_w11062_,
		_w11063_
	);
	LUT2 #(
		.INIT('h2)
	) name10602 (
		\P1_state_reg[0]/NET0131 ,
		_w11063_,
		_w11064_
	);
	LUT2 #(
		.INIT('h1)
	) name10603 (
		_w11042_,
		_w11064_,
		_w11065_
	);
	LUT2 #(
		.INIT('h2)
	) name10604 (
		\P1_reg3_reg[0]/NET0131 ,
		_w3435_,
		_w11066_
	);
	LUT2 #(
		.INIT('h8)
	) name10605 (
		\P1_reg3_reg[0]/NET0131 ,
		_w3448_,
		_w11067_
	);
	LUT2 #(
		.INIT('h1)
	) name10606 (
		_w1765_,
		_w1888_,
		_w11068_
	);
	LUT2 #(
		.INIT('h2)
	) name10607 (
		\P1_reg3_reg[0]/NET0131 ,
		_w3980_,
		_w11069_
	);
	LUT2 #(
		.INIT('h4)
	) name10608 (
		_w1804_,
		_w3980_,
		_w11070_
	);
	LUT2 #(
		.INIT('h1)
	) name10609 (
		_w11069_,
		_w11070_,
		_w11071_
	);
	LUT2 #(
		.INIT('h1)
	) name10610 (
		_w11068_,
		_w11071_,
		_w11072_
	);
	LUT2 #(
		.INIT('h1)
	) name10611 (
		_w1761_,
		_w3980_,
		_w11073_
	);
	LUT2 #(
		.INIT('h4)
	) name10612 (
		_w1671_,
		_w1762_,
		_w11074_
	);
	LUT2 #(
		.INIT('h4)
	) name10613 (
		_w11073_,
		_w11074_,
		_w11075_
	);
	LUT2 #(
		.INIT('h2)
	) name10614 (
		\P1_reg3_reg[0]/NET0131 ,
		_w9092_,
		_w11076_
	);
	LUT2 #(
		.INIT('h2)
	) name10615 (
		_w1641_,
		_w3570_,
		_w11077_
	);
	LUT2 #(
		.INIT('h1)
	) name10616 (
		_w537_,
		_w3571_,
		_w11078_
	);
	LUT2 #(
		.INIT('h4)
	) name10617 (
		_w11077_,
		_w11078_,
		_w11079_
	);
	LUT2 #(
		.INIT('h8)
	) name10618 (
		_w3980_,
		_w11079_,
		_w11080_
	);
	LUT2 #(
		.INIT('h1)
	) name10619 (
		_w11069_,
		_w11080_,
		_w11081_
	);
	LUT2 #(
		.INIT('h2)
	) name10620 (
		_w1936_,
		_w11081_,
		_w11082_
	);
	LUT2 #(
		.INIT('h1)
	) name10621 (
		_w11072_,
		_w11075_,
		_w11083_
	);
	LUT2 #(
		.INIT('h4)
	) name10622 (
		_w11076_,
		_w11083_,
		_w11084_
	);
	LUT2 #(
		.INIT('h4)
	) name10623 (
		_w11082_,
		_w11084_,
		_w11085_
	);
	LUT2 #(
		.INIT('h2)
	) name10624 (
		_w3450_,
		_w11085_,
		_w11086_
	);
	LUT2 #(
		.INIT('h1)
	) name10625 (
		_w11067_,
		_w11086_,
		_w11087_
	);
	LUT2 #(
		.INIT('h2)
	) name10626 (
		\P1_state_reg[0]/NET0131 ,
		_w11087_,
		_w11088_
	);
	LUT2 #(
		.INIT('h1)
	) name10627 (
		_w11066_,
		_w11088_,
		_w11089_
	);
	LUT2 #(
		.INIT('h2)
	) name10628 (
		\P2_reg3_reg[0]/NET0131 ,
		_w1983_,
		_w11090_
	);
	LUT2 #(
		.INIT('h8)
	) name10629 (
		\P2_reg3_reg[0]/NET0131 ,
		_w2024_,
		_w11091_
	);
	LUT2 #(
		.INIT('h8)
	) name10630 (
		\P2_reg3_reg[0]/NET0131 ,
		_w3417_,
		_w11092_
	);
	LUT2 #(
		.INIT('h2)
	) name10631 (
		\P2_reg3_reg[0]/NET0131 ,
		_w3788_,
		_w11093_
	);
	LUT2 #(
		.INIT('h2)
	) name10632 (
		_w3788_,
		_w4204_,
		_w11094_
	);
	LUT2 #(
		.INIT('h1)
	) name10633 (
		_w11093_,
		_w11094_,
		_w11095_
	);
	LUT2 #(
		.INIT('h1)
	) name10634 (
		_w3744_,
		_w11095_,
		_w11096_
	);
	LUT2 #(
		.INIT('h4)
	) name10635 (
		_w2604_,
		_w3788_,
		_w11097_
	);
	LUT2 #(
		.INIT('h1)
	) name10636 (
		_w11093_,
		_w11097_,
		_w11098_
	);
	LUT2 #(
		.INIT('h2)
	) name10637 (
		_w9903_,
		_w11098_,
		_w11099_
	);
	LUT2 #(
		.INIT('h2)
	) name10638 (
		_w2574_,
		_w3373_,
		_w11100_
	);
	LUT2 #(
		.INIT('h1)
	) name10639 (
		_w2058_,
		_w3374_,
		_w11101_
	);
	LUT2 #(
		.INIT('h4)
	) name10640 (
		_w11100_,
		_w11101_,
		_w11102_
	);
	LUT2 #(
		.INIT('h8)
	) name10641 (
		_w3788_,
		_w11102_,
		_w11103_
	);
	LUT2 #(
		.INIT('h1)
	) name10642 (
		_w11093_,
		_w11103_,
		_w11104_
	);
	LUT2 #(
		.INIT('h2)
	) name10643 (
		_w3411_,
		_w11104_,
		_w11105_
	);
	LUT2 #(
		.INIT('h4)
	) name10644 (
		_w2604_,
		_w3420_,
		_w11106_
	);
	LUT2 #(
		.INIT('h1)
	) name10645 (
		_w11092_,
		_w11106_,
		_w11107_
	);
	LUT2 #(
		.INIT('h4)
	) name10646 (
		_w11096_,
		_w11107_,
		_w11108_
	);
	LUT2 #(
		.INIT('h4)
	) name10647 (
		_w11099_,
		_w11108_,
		_w11109_
	);
	LUT2 #(
		.INIT('h4)
	) name10648 (
		_w11105_,
		_w11109_,
		_w11110_
	);
	LUT2 #(
		.INIT('h2)
	) name10649 (
		_w2026_,
		_w11110_,
		_w11111_
	);
	LUT2 #(
		.INIT('h1)
	) name10650 (
		_w11091_,
		_w11111_,
		_w11112_
	);
	LUT2 #(
		.INIT('h2)
	) name10651 (
		\P1_state_reg[0]/NET0131 ,
		_w11112_,
		_w11113_
	);
	LUT2 #(
		.INIT('h1)
	) name10652 (
		_w11090_,
		_w11113_,
		_w11114_
	);
	LUT2 #(
		.INIT('h1)
	) name10653 (
		\P1_reg2_reg[0]/NET0131 ,
		_w5812_,
		_w11115_
	);
	LUT2 #(
		.INIT('h8)
	) name10654 (
		\P1_reg3_reg[0]/NET0131 ,
		_w1763_,
		_w11116_
	);
	LUT2 #(
		.INIT('h8)
	) name10655 (
		_w1936_,
		_w11079_,
		_w11117_
	);
	LUT2 #(
		.INIT('h4)
	) name10656 (
		_w1671_,
		_w9090_,
		_w11118_
	);
	LUT2 #(
		.INIT('h1)
	) name10657 (
		_w1804_,
		_w11068_,
		_w11119_
	);
	LUT2 #(
		.INIT('h1)
	) name10658 (
		_w11118_,
		_w11119_,
		_w11120_
	);
	LUT2 #(
		.INIT('h4)
	) name10659 (
		_w11117_,
		_w11120_,
		_w11121_
	);
	LUT2 #(
		.INIT('h2)
	) name10660 (
		_w3466_,
		_w11121_,
		_w11122_
	);
	LUT2 #(
		.INIT('h4)
	) name10661 (
		_w1936_,
		_w11068_,
		_w11123_
	);
	LUT2 #(
		.INIT('h1)
	) name10662 (
		_w3466_,
		_w11123_,
		_w11124_
	);
	LUT2 #(
		.INIT('h2)
	) name10663 (
		_w5815_,
		_w9953_,
		_w11125_
	);
	LUT2 #(
		.INIT('h4)
	) name10664 (
		_w11124_,
		_w11125_,
		_w11126_
	);
	LUT2 #(
		.INIT('h2)
	) name10665 (
		\P1_reg2_reg[0]/NET0131 ,
		_w11126_,
		_w11127_
	);
	LUT2 #(
		.INIT('h1)
	) name10666 (
		_w11116_,
		_w11127_,
		_w11128_
	);
	LUT2 #(
		.INIT('h4)
	) name10667 (
		_w11122_,
		_w11128_,
		_w11129_
	);
	LUT2 #(
		.INIT('h1)
	) name10668 (
		_w11115_,
		_w11129_,
		_w11130_
	);
	LUT2 #(
		.INIT('h2)
	) name10669 (
		\P2_reg1_reg[0]/NET0131 ,
		_w1983_,
		_w11131_
	);
	LUT2 #(
		.INIT('h8)
	) name10670 (
		\P2_reg1_reg[0]/NET0131 ,
		_w2024_,
		_w11132_
	);
	LUT2 #(
		.INIT('h2)
	) name10671 (
		\P2_reg1_reg[0]/NET0131 ,
		_w3733_,
		_w11133_
	);
	LUT2 #(
		.INIT('h4)
	) name10672 (
		_w2604_,
		_w3733_,
		_w11134_
	);
	LUT2 #(
		.INIT('h1)
	) name10673 (
		_w11133_,
		_w11134_,
		_w11135_
	);
	LUT2 #(
		.INIT('h2)
	) name10674 (
		_w9903_,
		_w11135_,
		_w11136_
	);
	LUT2 #(
		.INIT('h2)
	) name10675 (
		_w3733_,
		_w4204_,
		_w11137_
	);
	LUT2 #(
		.INIT('h1)
	) name10676 (
		_w11133_,
		_w11137_,
		_w11138_
	);
	LUT2 #(
		.INIT('h1)
	) name10677 (
		_w3744_,
		_w11138_,
		_w11139_
	);
	LUT2 #(
		.INIT('h2)
	) name10678 (
		\P2_reg1_reg[0]/NET0131 ,
		_w3421_,
		_w11140_
	);
	LUT2 #(
		.INIT('h8)
	) name10679 (
		_w3733_,
		_w11102_,
		_w11141_
	);
	LUT2 #(
		.INIT('h1)
	) name10680 (
		_w11133_,
		_w11141_,
		_w11142_
	);
	LUT2 #(
		.INIT('h2)
	) name10681 (
		_w3411_,
		_w11142_,
		_w11143_
	);
	LUT2 #(
		.INIT('h1)
	) name10682 (
		_w11136_,
		_w11140_,
		_w11144_
	);
	LUT2 #(
		.INIT('h4)
	) name10683 (
		_w11139_,
		_w11144_,
		_w11145_
	);
	LUT2 #(
		.INIT('h4)
	) name10684 (
		_w11143_,
		_w11145_,
		_w11146_
	);
	LUT2 #(
		.INIT('h2)
	) name10685 (
		_w2026_,
		_w11146_,
		_w11147_
	);
	LUT2 #(
		.INIT('h1)
	) name10686 (
		_w11132_,
		_w11147_,
		_w11148_
	);
	LUT2 #(
		.INIT('h2)
	) name10687 (
		\P1_state_reg[0]/NET0131 ,
		_w11148_,
		_w11149_
	);
	LUT2 #(
		.INIT('h1)
	) name10688 (
		_w11131_,
		_w11149_,
		_w11150_
	);
	LUT2 #(
		.INIT('h8)
	) name10689 (
		\P2_reg3_reg[0]/NET0131 ,
		_w3420_,
		_w11151_
	);
	LUT2 #(
		.INIT('h1)
	) name10690 (
		_w3744_,
		_w4204_,
		_w11152_
	);
	LUT2 #(
		.INIT('h4)
	) name10691 (
		_w2604_,
		_w9903_,
		_w11153_
	);
	LUT2 #(
		.INIT('h8)
	) name10692 (
		_w3411_,
		_w11102_,
		_w11154_
	);
	LUT2 #(
		.INIT('h1)
	) name10693 (
		_w11152_,
		_w11153_,
		_w11155_
	);
	LUT2 #(
		.INIT('h4)
	) name10694 (
		_w11154_,
		_w11155_,
		_w11156_
	);
	LUT2 #(
		.INIT('h2)
	) name10695 (
		_w3758_,
		_w11156_,
		_w11157_
	);
	LUT2 #(
		.INIT('h1)
	) name10696 (
		_w11151_,
		_w11157_,
		_w11158_
	);
	LUT2 #(
		.INIT('h2)
	) name10697 (
		_w5287_,
		_w11158_,
		_w11159_
	);
	LUT2 #(
		.INIT('h2)
	) name10698 (
		\P2_reg2_reg[0]/NET0131 ,
		_w10018_,
		_w11160_
	);
	LUT2 #(
		.INIT('h1)
	) name10699 (
		_w11159_,
		_w11160_,
		_w11161_
	);
	LUT2 #(
		.INIT('h2)
	) name10700 (
		\P1_reg0_reg[0]/NET0131 ,
		_w3435_,
		_w11162_
	);
	LUT2 #(
		.INIT('h8)
	) name10701 (
		\P1_reg0_reg[0]/NET0131 ,
		_w3448_,
		_w11163_
	);
	LUT2 #(
		.INIT('h2)
	) name10702 (
		\P1_reg0_reg[0]/NET0131 ,
		_w4396_,
		_w11164_
	);
	LUT2 #(
		.INIT('h4)
	) name10703 (
		_w1804_,
		_w4396_,
		_w11165_
	);
	LUT2 #(
		.INIT('h1)
	) name10704 (
		_w11164_,
		_w11165_,
		_w11166_
	);
	LUT2 #(
		.INIT('h1)
	) name10705 (
		_w11068_,
		_w11166_,
		_w11167_
	);
	LUT2 #(
		.INIT('h4)
	) name10706 (
		_w1671_,
		_w4396_,
		_w11168_
	);
	LUT2 #(
		.INIT('h1)
	) name10707 (
		_w11164_,
		_w11168_,
		_w11169_
	);
	LUT2 #(
		.INIT('h2)
	) name10708 (
		_w9090_,
		_w11169_,
		_w11170_
	);
	LUT2 #(
		.INIT('h2)
	) name10709 (
		\P1_reg0_reg[0]/NET0131 ,
		_w4491_,
		_w11171_
	);
	LUT2 #(
		.INIT('h8)
	) name10710 (
		_w4396_,
		_w11079_,
		_w11172_
	);
	LUT2 #(
		.INIT('h1)
	) name10711 (
		_w11164_,
		_w11172_,
		_w11173_
	);
	LUT2 #(
		.INIT('h2)
	) name10712 (
		_w1936_,
		_w11173_,
		_w11174_
	);
	LUT2 #(
		.INIT('h1)
	) name10713 (
		_w11167_,
		_w11171_,
		_w11175_
	);
	LUT2 #(
		.INIT('h4)
	) name10714 (
		_w11170_,
		_w11175_,
		_w11176_
	);
	LUT2 #(
		.INIT('h4)
	) name10715 (
		_w11174_,
		_w11176_,
		_w11177_
	);
	LUT2 #(
		.INIT('h2)
	) name10716 (
		_w3450_,
		_w11177_,
		_w11178_
	);
	LUT2 #(
		.INIT('h1)
	) name10717 (
		_w11163_,
		_w11178_,
		_w11179_
	);
	LUT2 #(
		.INIT('h2)
	) name10718 (
		\P1_state_reg[0]/NET0131 ,
		_w11179_,
		_w11180_
	);
	LUT2 #(
		.INIT('h1)
	) name10719 (
		_w11162_,
		_w11180_,
		_w11181_
	);
	LUT2 #(
		.INIT('h2)
	) name10720 (
		_w6368_,
		_w11121_,
		_w11182_
	);
	LUT2 #(
		.INIT('h1)
	) name10721 (
		_w4532_,
		_w11123_,
		_w11183_
	);
	LUT2 #(
		.INIT('h2)
	) name10722 (
		_w5812_,
		_w11183_,
		_w11184_
	);
	LUT2 #(
		.INIT('h8)
	) name10723 (
		_w9835_,
		_w11184_,
		_w11185_
	);
	LUT2 #(
		.INIT('h2)
	) name10724 (
		\P1_reg1_reg[0]/NET0131 ,
		_w11185_,
		_w11186_
	);
	LUT2 #(
		.INIT('h1)
	) name10725 (
		_w11182_,
		_w11186_,
		_w11187_
	);
	LUT2 #(
		.INIT('h2)
	) name10726 (
		\P2_reg0_reg[0]/NET0131 ,
		_w1983_,
		_w11188_
	);
	LUT2 #(
		.INIT('h8)
	) name10727 (
		\P2_reg0_reg[0]/NET0131 ,
		_w2024_,
		_w11189_
	);
	LUT2 #(
		.INIT('h2)
	) name10728 (
		\P2_reg0_reg[0]/NET0131 ,
		_w2040_,
		_w11190_
	);
	LUT2 #(
		.INIT('h2)
	) name10729 (
		_w2040_,
		_w2604_,
		_w11191_
	);
	LUT2 #(
		.INIT('h1)
	) name10730 (
		_w11190_,
		_w11191_,
		_w11192_
	);
	LUT2 #(
		.INIT('h2)
	) name10731 (
		_w9903_,
		_w11192_,
		_w11193_
	);
	LUT2 #(
		.INIT('h2)
	) name10732 (
		_w2040_,
		_w4204_,
		_w11194_
	);
	LUT2 #(
		.INIT('h1)
	) name10733 (
		_w11190_,
		_w11194_,
		_w11195_
	);
	LUT2 #(
		.INIT('h1)
	) name10734 (
		_w3744_,
		_w11195_,
		_w11196_
	);
	LUT2 #(
		.INIT('h2)
	) name10735 (
		\P2_reg0_reg[0]/NET0131 ,
		_w3421_,
		_w11197_
	);
	LUT2 #(
		.INIT('h8)
	) name10736 (
		_w2040_,
		_w11102_,
		_w11198_
	);
	LUT2 #(
		.INIT('h1)
	) name10737 (
		_w11190_,
		_w11198_,
		_w11199_
	);
	LUT2 #(
		.INIT('h2)
	) name10738 (
		_w3411_,
		_w11199_,
		_w11200_
	);
	LUT2 #(
		.INIT('h1)
	) name10739 (
		_w11193_,
		_w11197_,
		_w11201_
	);
	LUT2 #(
		.INIT('h4)
	) name10740 (
		_w11196_,
		_w11201_,
		_w11202_
	);
	LUT2 #(
		.INIT('h4)
	) name10741 (
		_w11200_,
		_w11202_,
		_w11203_
	);
	LUT2 #(
		.INIT('h2)
	) name10742 (
		_w2026_,
		_w11203_,
		_w11204_
	);
	LUT2 #(
		.INIT('h1)
	) name10743 (
		_w11189_,
		_w11204_,
		_w11205_
	);
	LUT2 #(
		.INIT('h2)
	) name10744 (
		\P1_state_reg[0]/NET0131 ,
		_w11205_,
		_w11206_
	);
	LUT2 #(
		.INIT('h1)
	) name10745 (
		_w11188_,
		_w11206_,
		_w11207_
	);
	LUT2 #(
		.INIT('h1)
	) name10746 (
		\P1_state_reg[0]/NET0131 ,
		_w1028_,
		_w11208_
	);
	LUT2 #(
		.INIT('h2)
	) name10747 (
		\P1_state_reg[0]/NET0131 ,
		_w3439_,
		_w11209_
	);
	LUT2 #(
		.INIT('h1)
	) name10748 (
		_w11208_,
		_w11209_,
		_w11210_
	);
	LUT2 #(
		.INIT('h1)
	) name10749 (
		\P1_state_reg[0]/NET0131 ,
		_w996_,
		_w11211_
	);
	LUT2 #(
		.INIT('h2)
	) name10750 (
		\P1_state_reg[0]/NET0131 ,
		_w3442_,
		_w11212_
	);
	LUT2 #(
		.INIT('h1)
	) name10751 (
		_w11211_,
		_w11212_,
		_w11213_
	);
	LUT2 #(
		.INIT('h1)
	) name10752 (
		\P1_state_reg[0]/NET0131 ,
		_w968_,
		_w11214_
	);
	LUT2 #(
		.INIT('h8)
	) name10753 (
		\P1_state_reg[0]/NET0131 ,
		_w527_,
		_w11215_
	);
	LUT2 #(
		.INIT('h1)
	) name10754 (
		_w11214_,
		_w11215_,
		_w11216_
	);
	LUT2 #(
		.INIT('h1)
	) name10755 (
		\P1_state_reg[0]/NET0131 ,
		_w3033_,
		_w11217_
	);
	LUT2 #(
		.INIT('h8)
	) name10756 (
		\P1_state_reg[0]/NET0131 ,
		_w2022_,
		_w11218_
	);
	LUT2 #(
		.INIT('h1)
	) name10757 (
		_w11217_,
		_w11218_,
		_w11219_
	);
	LUT2 #(
		.INIT('h1)
	) name10758 (
		\P1_state_reg[0]/NET0131 ,
		_w3011_,
		_w11220_
	);
	LUT2 #(
		.INIT('h8)
	) name10759 (
		\P1_state_reg[0]/NET0131 ,
		_w2001_,
		_w11221_
	);
	LUT2 #(
		.INIT('h1)
	) name10760 (
		_w11220_,
		_w11221_,
		_w11222_
	);
	LUT2 #(
		.INIT('h1)
	) name10761 (
		\P1_state_reg[0]/NET0131 ,
		_w2981_,
		_w11223_
	);
	LUT2 #(
		.INIT('h8)
	) name10762 (
		\P1_state_reg[0]/NET0131 ,
		_w2051_,
		_w11224_
	);
	LUT2 #(
		.INIT('h1)
	) name10763 (
		_w11223_,
		_w11224_,
		_w11225_
	);
	LUT2 #(
		.INIT('h1)
	) name10764 (
		\P1_state_reg[0]/NET0131 ,
		_w2753_,
		_w11226_
	);
	LUT2 #(
		.INIT('h2)
	) name10765 (
		\P1_state_reg[0]/NET0131 ,
		_w2745_,
		_w11227_
	);
	LUT2 #(
		.INIT('h1)
	) name10766 (
		_w11226_,
		_w11227_,
		_w11228_
	);
	LUT2 #(
		.INIT('h2)
	) name10767 (
		\P1_state_reg[0]/NET0131 ,
		_w2694_,
		_w11229_
	);
	LUT2 #(
		.INIT('h4)
	) name10768 (
		\P1_state_reg[0]/NET0131 ,
		_w2702_,
		_w11230_
	);
	LUT2 #(
		.INIT('h1)
	) name10769 (
		_w11229_,
		_w11230_,
		_w11231_
	);
	LUT2 #(
		.INIT('h2)
	) name10770 (
		\P1_state_reg[0]/NET0131 ,
		_w2720_,
		_w11232_
	);
	LUT2 #(
		.INIT('h4)
	) name10771 (
		\P1_state_reg[0]/NET0131 ,
		_w2729_,
		_w11233_
	);
	LUT2 #(
		.INIT('h1)
	) name10772 (
		_w11232_,
		_w11233_,
		_w11234_
	);
	LUT2 #(
		.INIT('h1)
	) name10773 (
		\P1_state_reg[0]/NET0131 ,
		_w2891_,
		_w11235_
	);
	LUT2 #(
		.INIT('h2)
	) name10774 (
		\P1_state_reg[0]/NET0131 ,
		_w2883_,
		_w11236_
	);
	LUT2 #(
		.INIT('h1)
	) name10775 (
		_w11235_,
		_w11236_,
		_w11237_
	);
	LUT2 #(
		.INIT('h2)
	) name10776 (
		\P1_state_reg[0]/NET0131 ,
		_w2849_,
		_w11238_
	);
	LUT2 #(
		.INIT('h4)
	) name10777 (
		\P1_state_reg[0]/NET0131 ,
		_w2858_,
		_w11239_
	);
	LUT2 #(
		.INIT('h1)
	) name10778 (
		_w11238_,
		_w11239_,
		_w11240_
	);
	LUT2 #(
		.INIT('h1)
	) name10779 (
		\P1_state_reg[0]/NET0131 ,
		_w2841_,
		_w11241_
	);
	LUT2 #(
		.INIT('h8)
	) name10780 (
		\P1_state_reg[0]/NET0131 ,
		_w2832_,
		_w11242_
	);
	LUT2 #(
		.INIT('h1)
	) name10781 (
		_w11241_,
		_w11242_,
		_w11243_
	);
	LUT2 #(
		.INIT('h2)
	) name10782 (
		\P1_state_reg[0]/NET0131 ,
		_w2808_,
		_w11244_
	);
	LUT2 #(
		.INIT('h4)
	) name10783 (
		\P1_state_reg[0]/NET0131 ,
		_w2816_,
		_w11245_
	);
	LUT2 #(
		.INIT('h1)
	) name10784 (
		_w11244_,
		_w11245_,
		_w11246_
	);
	LUT2 #(
		.INIT('h2)
	) name10785 (
		\P1_state_reg[0]/NET0131 ,
		_w2385_,
		_w11247_
	);
	LUT2 #(
		.INIT('h4)
	) name10786 (
		\P1_state_reg[0]/NET0131 ,
		_w2397_,
		_w11248_
	);
	LUT2 #(
		.INIT('h1)
	) name10787 (
		_w11247_,
		_w11248_,
		_w11249_
	);
	LUT2 #(
		.INIT('h2)
	) name10788 (
		\P1_state_reg[0]/NET0131 ,
		_w2404_,
		_w11250_
	);
	LUT2 #(
		.INIT('h4)
	) name10789 (
		\P1_state_reg[0]/NET0131 ,
		_w2431_,
		_w11251_
	);
	LUT2 #(
		.INIT('h1)
	) name10790 (
		_w11250_,
		_w11251_,
		_w11252_
	);
	LUT2 #(
		.INIT('h1)
	) name10791 (
		\P1_state_reg[0]/NET0131 ,
		_w2297_,
		_w11253_
	);
	LUT2 #(
		.INIT('h8)
	) name10792 (
		\P1_state_reg[0]/NET0131 ,
		_w2258_,
		_w11254_
	);
	LUT2 #(
		.INIT('h1)
	) name10793 (
		_w11253_,
		_w11254_,
		_w11255_
	);
	LUT2 #(
		.INIT('h8)
	) name10794 (
		\P1_state_reg[0]/NET0131 ,
		_w2578_,
		_w11256_
	);
	LUT2 #(
		.INIT('h4)
	) name10795 (
		\P1_state_reg[0]/NET0131 ,
		_w2586_,
		_w11257_
	);
	LUT2 #(
		.INIT('h1)
	) name10796 (
		_w11256_,
		_w11257_,
		_w11258_
	);
	LUT2 #(
		.INIT('h1)
	) name10797 (
		\P1_state_reg[0]/NET0131 ,
		_w2357_,
		_w11259_
	);
	LUT2 #(
		.INIT('h2)
	) name10798 (
		\P1_state_reg[0]/NET0131 ,
		_w3175_,
		_w11260_
	);
	LUT2 #(
		.INIT('h1)
	) name10799 (
		_w11259_,
		_w11260_,
		_w11261_
	);
	LUT2 #(
		.INIT('h1)
	) name10800 (
		\P1_state_reg[0]/NET0131 ,
		_w3120_,
		_w11262_
	);
	LUT2 #(
		.INIT('h2)
	) name10801 (
		\P1_state_reg[0]/NET0131 ,
		_w3170_,
		_w11263_
	);
	LUT2 #(
		.INIT('h1)
	) name10802 (
		_w11262_,
		_w11263_,
		_w11264_
	);
	LUT2 #(
		.INIT('h1)
	) name10803 (
		\P1_state_reg[0]/NET0131 ,
		_w3101_,
		_w11265_
	);
	LUT2 #(
		.INIT('h8)
	) name10804 (
		\P1_state_reg[0]/NET0131 ,
		_w3166_,
		_w11266_
	);
	LUT2 #(
		.INIT('h1)
	) name10805 (
		_w11265_,
		_w11266_,
		_w11267_
	);
	LUT2 #(
		.INIT('h1)
	) name10806 (
		\P1_state_reg[0]/NET0131 ,
		_w3078_,
		_w11268_
	);
	LUT2 #(
		.INIT('h1)
	) name10807 (
		_w3976_,
		_w11268_,
		_w11269_
	);
	LUT2 #(
		.INIT('h1)
	) name10808 (
		\P1_state_reg[0]/NET0131 ,
		_w3053_,
		_w11270_
	);
	LUT2 #(
		.INIT('h8)
	) name10809 (
		\P1_state_reg[0]/NET0131 ,
		_w2008_,
		_w11271_
	);
	LUT2 #(
		.INIT('h1)
	) name10810 (
		_w11270_,
		_w11271_,
		_w11272_
	);
	LUT2 #(
		.INIT('h2)
	) name10811 (
		\P1_state_reg[0]/NET0131 ,
		_w2215_,
		_w11273_
	);
	LUT2 #(
		.INIT('h4)
	) name10812 (
		\P1_state_reg[0]/NET0131 ,
		_w2197_,
		_w11274_
	);
	LUT2 #(
		.INIT('h1)
	) name10813 (
		_w11273_,
		_w11274_,
		_w11275_
	);
	LUT2 #(
		.INIT('h1)
	) name10814 (
		\P1_state_reg[0]/NET0131 ,
		_w2559_,
		_w11276_
	);
	LUT2 #(
		.INIT('h8)
	) name10815 (
		\P1_state_reg[0]/NET0131 ,
		_w2564_,
		_w11277_
	);
	LUT2 #(
		.INIT('h1)
	) name10816 (
		_w11276_,
		_w11277_,
		_w11278_
	);
	LUT2 #(
		.INIT('h1)
	) name10817 (
		\P1_state_reg[0]/NET0131 ,
		_w4158_,
		_w11279_
	);
	LUT2 #(
		.INIT('h8)
	) name10818 (
		\P1_state_reg[0]/NET0131 ,
		_w2207_,
		_w11280_
	);
	LUT2 #(
		.INIT('h1)
	) name10819 (
		_w11279_,
		_w11280_,
		_w11281_
	);
	LUT2 #(
		.INIT('h2)
	) name10820 (
		\P1_state_reg[0]/NET0131 ,
		_w2629_,
		_w11282_
	);
	LUT2 #(
		.INIT('h4)
	) name10821 (
		\P1_state_reg[0]/NET0131 ,
		_w2623_,
		_w11283_
	);
	LUT2 #(
		.INIT('h1)
	) name10822 (
		_w11282_,
		_w11283_,
		_w11284_
	);
	LUT2 #(
		.INIT('h8)
	) name10823 (
		\P1_state_reg[0]/NET0131 ,
		_w2646_,
		_w11285_
	);
	LUT2 #(
		.INIT('h4)
	) name10824 (
		\P1_state_reg[0]/NET0131 ,
		_w2654_,
		_w11286_
	);
	LUT2 #(
		.INIT('h1)
	) name10825 (
		_w11285_,
		_w11286_,
		_w11287_
	);
	LUT2 #(
		.INIT('h1)
	) name10826 (
		\P1_state_reg[0]/NET0131 ,
		_w2538_,
		_w11288_
	);
	LUT2 #(
		.INIT('h2)
	) name10827 (
		\P1_state_reg[0]/NET0131 ,
		_w2542_,
		_w11289_
	);
	LUT2 #(
		.INIT('h1)
	) name10828 (
		_w11288_,
		_w11289_,
		_w11290_
	);
	LUT2 #(
		.INIT('h1)
	) name10829 (
		\P1_state_reg[0]/NET0131 ,
		_w2513_,
		_w11291_
	);
	LUT2 #(
		.INIT('h8)
	) name10830 (
		\P1_state_reg[0]/NET0131 ,
		_w2519_,
		_w11292_
	);
	LUT2 #(
		.INIT('h1)
	) name10831 (
		_w11291_,
		_w11292_,
		_w11293_
	);
	LUT2 #(
		.INIT('h2)
	) name10832 (
		\P1_state_reg[0]/NET0131 ,
		_w2485_,
		_w11294_
	);
	LUT2 #(
		.INIT('h4)
	) name10833 (
		\P1_state_reg[0]/NET0131 ,
		_w2493_,
		_w11295_
	);
	LUT2 #(
		.INIT('h1)
	) name10834 (
		_w11294_,
		_w11295_,
		_w11296_
	);
	LUT2 #(
		.INIT('h2)
	) name10835 (
		\P1_state_reg[0]/NET0131 ,
		_w2460_,
		_w11297_
	);
	LUT2 #(
		.INIT('h4)
	) name10836 (
		\P1_state_reg[0]/NET0131 ,
		_w2468_,
		_w11298_
	);
	LUT2 #(
		.INIT('h1)
	) name10837 (
		_w11297_,
		_w11298_,
		_w11299_
	);
	LUT2 #(
		.INIT('h1)
	) name10838 (
		\P1_state_reg[0]/NET0131 ,
		_w2777_,
		_w11300_
	);
	LUT2 #(
		.INIT('h2)
	) name10839 (
		\P1_state_reg[0]/NET0131 ,
		_w2769_,
		_w11301_
	);
	LUT2 #(
		.INIT('h1)
	) name10840 (
		_w11300_,
		_w11301_,
		_w11302_
	);
	LUT2 #(
		.INIT('h1)
	) name10841 (
		\P1_state_reg[0]/NET0131 ,
		_w2948_,
		_w11303_
	);
	LUT2 #(
		.INIT('h8)
	) name10842 (
		\P1_state_reg[0]/NET0131 ,
		_w2058_,
		_w11304_
	);
	LUT2 #(
		.INIT('h1)
	) name10843 (
		_w11303_,
		_w11304_,
		_w11305_
	);
	LUT2 #(
		.INIT('h2)
	) name10844 (
		\P1_state_reg[0]/NET0131 ,
		_w1223_,
		_w11306_
	);
	LUT2 #(
		.INIT('h4)
	) name10845 (
		\P1_state_reg[0]/NET0131 ,
		_w1231_,
		_w11307_
	);
	LUT2 #(
		.INIT('h1)
	) name10846 (
		_w11306_,
		_w11307_,
		_w11308_
	);
	LUT2 #(
		.INIT('h1)
	) name10847 (
		\P1_state_reg[0]/NET0131 ,
		_w1196_,
		_w11309_
	);
	LUT2 #(
		.INIT('h8)
	) name10848 (
		\P1_state_reg[0]/NET0131 ,
		_w1188_,
		_w11310_
	);
	LUT2 #(
		.INIT('h1)
	) name10849 (
		_w11309_,
		_w11310_,
		_w11311_
	);
	LUT2 #(
		.INIT('h2)
	) name10850 (
		\P1_state_reg[0]/NET0131 ,
		_w1154_,
		_w11312_
	);
	LUT2 #(
		.INIT('h4)
	) name10851 (
		\P1_state_reg[0]/NET0131 ,
		_w1163_,
		_w11313_
	);
	LUT2 #(
		.INIT('h1)
	) name10852 (
		_w11312_,
		_w11313_,
		_w11314_
	);
	LUT2 #(
		.INIT('h2)
	) name10853 (
		\P1_state_reg[0]/NET0131 ,
		_w1126_,
		_w11315_
	);
	LUT2 #(
		.INIT('h4)
	) name10854 (
		\P1_state_reg[0]/NET0131 ,
		_w1134_,
		_w11316_
	);
	LUT2 #(
		.INIT('h1)
	) name10855 (
		_w11315_,
		_w11316_,
		_w11317_
	);
	LUT2 #(
		.INIT('h1)
	) name10856 (
		\P1_state_reg[0]/NET0131 ,
		_w1107_,
		_w11318_
	);
	LUT2 #(
		.INIT('h8)
	) name10857 (
		\P1_state_reg[0]/NET0131 ,
		_w1099_,
		_w11319_
	);
	LUT2 #(
		.INIT('h1)
	) name10858 (
		_w11318_,
		_w11319_,
		_w11320_
	);
	LUT2 #(
		.INIT('h1)
	) name10859 (
		\P1_state_reg[0]/NET0131 ,
		_w1081_,
		_w11321_
	);
	LUT2 #(
		.INIT('h8)
	) name10860 (
		\P1_state_reg[0]/NET0131 ,
		_w1073_,
		_w11322_
	);
	LUT2 #(
		.INIT('h1)
	) name10861 (
		_w11321_,
		_w11322_,
		_w11323_
	);
	LUT2 #(
		.INIT('h1)
	) name10862 (
		\P1_state_reg[0]/NET0131 ,
		_w1464_,
		_w11324_
	);
	LUT2 #(
		.INIT('h8)
	) name10863 (
		\P1_state_reg[0]/NET0131 ,
		_w1456_,
		_w11325_
	);
	LUT2 #(
		.INIT('h1)
	) name10864 (
		_w11324_,
		_w11325_,
		_w11326_
	);
	LUT2 #(
		.INIT('h1)
	) name10865 (
		\P1_state_reg[0]/NET0131 ,
		_w1441_,
		_w11327_
	);
	LUT2 #(
		.INIT('h2)
	) name10866 (
		\P1_state_reg[0]/NET0131 ,
		_w1433_,
		_w11328_
	);
	LUT2 #(
		.INIT('h1)
	) name10867 (
		_w11327_,
		_w11328_,
		_w11329_
	);
	LUT2 #(
		.INIT('h2)
	) name10868 (
		\P1_state_reg[0]/NET0131 ,
		_w1384_,
		_w11330_
	);
	LUT2 #(
		.INIT('h4)
	) name10869 (
		\P1_state_reg[0]/NET0131 ,
		_w1392_,
		_w11331_
	);
	LUT2 #(
		.INIT('h1)
	) name10870 (
		_w11330_,
		_w11331_,
		_w11332_
	);
	LUT2 #(
		.INIT('h1)
	) name10871 (
		\P1_state_reg[0]/NET0131 ,
		_w1416_,
		_w11333_
	);
	LUT2 #(
		.INIT('h8)
	) name10872 (
		\P1_state_reg[0]/NET0131 ,
		_w1408_,
		_w11334_
	);
	LUT2 #(
		.INIT('h1)
	) name10873 (
		_w11333_,
		_w11334_,
		_w11335_
	);
	LUT2 #(
		.INIT('h8)
	) name10874 (
		\P1_state_reg[0]/NET0131 ,
		_w1645_,
		_w11336_
	);
	LUT2 #(
		.INIT('h4)
	) name10875 (
		\P1_state_reg[0]/NET0131 ,
		_w1653_,
		_w11337_
	);
	LUT2 #(
		.INIT('h1)
	) name10876 (
		_w11336_,
		_w11337_,
		_w11338_
	);
	LUT2 #(
		.INIT('h2)
	) name10877 (
		\P1_state_reg[0]/NET0131 ,
		_w519_,
		_w11339_
	);
	LUT2 #(
		.INIT('h4)
	) name10878 (
		\P1_state_reg[0]/NET0131 ,
		_w1364_,
		_w11340_
	);
	LUT2 #(
		.INIT('h1)
	) name10879 (
		_w11339_,
		_w11340_,
		_w11341_
	);
	LUT2 #(
		.INIT('h1)
	) name10880 (
		\P1_state_reg[0]/NET0131 ,
		_w1345_,
		_w11342_
	);
	LUT2 #(
		.INIT('h8)
	) name10881 (
		\P1_state_reg[0]/NET0131 ,
		_w501_,
		_w11343_
	);
	LUT2 #(
		.INIT('h1)
	) name10882 (
		_w11342_,
		_w11343_,
		_w11344_
	);
	LUT2 #(
		.INIT('h1)
	) name10883 (
		\P1_state_reg[0]/NET0131 ,
		_w1326_,
		_w11345_
	);
	LUT2 #(
		.INIT('h1)
	) name10884 (
		_w1953_,
		_w11345_,
		_w11346_
	);
	LUT2 #(
		.INIT('h1)
	) name10885 (
		\P1_state_reg[0]/NET0131 ,
		_w1046_,
		_w11347_
	);
	LUT2 #(
		.INIT('h8)
	) name10886 (
		\P1_state_reg[0]/NET0131 ,
		_w3445_,
		_w11348_
	);
	LUT2 #(
		.INIT('h1)
	) name10887 (
		_w11347_,
		_w11348_,
		_w11349_
	);
	LUT2 #(
		.INIT('h1)
	) name10888 (
		\P1_state_reg[0]/NET0131 ,
		_w1308_,
		_w11350_
	);
	LUT2 #(
		.INIT('h8)
	) name10889 (
		\P1_state_reg[0]/NET0131 ,
		_w486_,
		_w11351_
	);
	LUT2 #(
		.INIT('h1)
	) name10890 (
		_w11350_,
		_w11351_,
		_w11352_
	);
	LUT2 #(
		.INIT('h1)
	) name10891 (
		\P1_state_reg[0]/NET0131 ,
		_w932_,
		_w11353_
	);
	LUT2 #(
		.INIT('h8)
	) name10892 (
		\P1_state_reg[0]/NET0131 ,
		_w537_,
		_w11354_
	);
	LUT2 #(
		.INIT('h1)
	) name10893 (
		_w11353_,
		_w11354_,
		_w11355_
	);
	LUT2 #(
		.INIT('h1)
	) name10894 (
		\P1_state_reg[0]/NET0131 ,
		_w880_,
		_w11356_
	);
	LUT2 #(
		.INIT('h8)
	) name10895 (
		\P1_state_reg[0]/NET0131 ,
		_w714_,
		_w11357_
	);
	LUT2 #(
		.INIT('h1)
	) name10896 (
		_w11356_,
		_w11357_,
		_w11358_
	);
	LUT2 #(
		.INIT('h1)
	) name10897 (
		\P1_state_reg[0]/NET0131 ,
		_w1602_,
		_w11359_
	);
	LUT2 #(
		.INIT('h8)
	) name10898 (
		\P1_state_reg[0]/NET0131 ,
		_w1607_,
		_w11360_
	);
	LUT2 #(
		.INIT('h1)
	) name10899 (
		_w11359_,
		_w11360_,
		_w11361_
	);
	LUT2 #(
		.INIT('h1)
	) name10900 (
		\P1_state_reg[0]/NET0131 ,
		_w824_,
		_w11362_
	);
	LUT2 #(
		.INIT('h8)
	) name10901 (
		\P1_state_reg[0]/NET0131 ,
		_w704_,
		_w11363_
	);
	LUT2 #(
		.INIT('h1)
	) name10902 (
		_w11362_,
		_w11363_,
		_w11364_
	);
	LUT2 #(
		.INIT('h4)
	) name10903 (
		\P1_state_reg[0]/NET0131 ,
		_w691_,
		_w11365_
	);
	LUT2 #(
		.INIT('h4)
	) name10904 (
		\P1_IR_reg[30]/NET0131 ,
		\P1_IR_reg[31]/NET0131 ,
		_w11366_
	);
	LUT2 #(
		.INIT('h8)
	) name10905 (
		\P1_state_reg[0]/NET0131 ,
		_w11366_,
		_w11367_
	);
	LUT2 #(
		.INIT('h8)
	) name10906 (
		_w698_,
		_w11367_,
		_w11368_
	);
	LUT2 #(
		.INIT('h8)
	) name10907 (
		_w523_,
		_w11368_,
		_w11369_
	);
	LUT2 #(
		.INIT('h1)
	) name10908 (
		_w11365_,
		_w11369_,
		_w11370_
	);
	LUT2 #(
		.INIT('h2)
	) name10909 (
		\P1_state_reg[0]/NET0131 ,
		_w1621_,
		_w11371_
	);
	LUT2 #(
		.INIT('h4)
	) name10910 (
		\P1_state_reg[0]/NET0131 ,
		_w1630_,
		_w11372_
	);
	LUT2 #(
		.INIT('h1)
	) name10911 (
		_w11371_,
		_w11372_,
		_w11373_
	);
	LUT2 #(
		.INIT('h1)
	) name10912 (
		\P1_state_reg[0]/NET0131 ,
		_w1579_,
		_w11374_
	);
	LUT2 #(
		.INIT('h2)
	) name10913 (
		\P1_state_reg[0]/NET0131 ,
		_w1584_,
		_w11375_
	);
	LUT2 #(
		.INIT('h1)
	) name10914 (
		_w11374_,
		_w11375_,
		_w11376_
	);
	LUT2 #(
		.INIT('h1)
	) name10915 (
		\P1_state_reg[0]/NET0131 ,
		_w1555_,
		_w11377_
	);
	LUT2 #(
		.INIT('h2)
	) name10916 (
		\P1_state_reg[0]/NET0131 ,
		_w1560_,
		_w11378_
	);
	LUT2 #(
		.INIT('h1)
	) name10917 (
		_w11377_,
		_w11378_,
		_w11379_
	);
	LUT2 #(
		.INIT('h1)
	) name10918 (
		\P1_state_reg[0]/NET0131 ,
		_w1531_,
		_w11380_
	);
	LUT2 #(
		.INIT('h2)
	) name10919 (
		\P1_state_reg[0]/NET0131 ,
		_w1535_,
		_w11381_
	);
	LUT2 #(
		.INIT('h1)
	) name10920 (
		_w11380_,
		_w11381_,
		_w11382_
	);
	LUT2 #(
		.INIT('h1)
	) name10921 (
		\P1_state_reg[0]/NET0131 ,
		_w1505_,
		_w11383_
	);
	LUT2 #(
		.INIT('h8)
	) name10922 (
		\P1_state_reg[0]/NET0131 ,
		_w1512_,
		_w11384_
	);
	LUT2 #(
		.INIT('h1)
	) name10923 (
		_w11383_,
		_w11384_,
		_w11385_
	);
	LUT2 #(
		.INIT('h1)
	) name10924 (
		\P1_state_reg[0]/NET0131 ,
		_w1279_,
		_w11386_
	);
	LUT2 #(
		.INIT('h8)
	) name10925 (
		\P1_state_reg[0]/NET0131 ,
		_w1271_,
		_w11387_
	);
	LUT2 #(
		.INIT('h1)
	) name10926 (
		_w11386_,
		_w11387_,
		_w11388_
	);
	LUT2 #(
		.INIT('h1)
	) name10927 (
		\P1_state_reg[0]/NET0131 ,
		_w1255_,
		_w11389_
	);
	LUT2 #(
		.INIT('h8)
	) name10928 (
		\P1_state_reg[0]/NET0131 ,
		_w1247_,
		_w11390_
	);
	LUT2 #(
		.INIT('h1)
	) name10929 (
		_w11389_,
		_w11390_,
		_w11391_
	);
	LUT2 #(
		.INIT('h4)
	) name10930 (
		\P1_state_reg[0]/NET0131 ,
		_w4140_,
		_w11392_
	);
	LUT2 #(
		.INIT('h2)
	) name10931 (
		\P1_state_reg[0]/NET0131 ,
		\P2_IR_reg[30]/NET0131 ,
		_w11393_
	);
	LUT2 #(
		.INIT('h8)
	) name10932 (
		\P2_IR_reg[31]/NET0131 ,
		_w11393_,
		_w11394_
	);
	LUT2 #(
		.INIT('h8)
	) name10933 (
		_w2044_,
		_w11394_,
		_w11395_
	);
	LUT2 #(
		.INIT('h8)
	) name10934 (
		_w2201_,
		_w11395_,
		_w11396_
	);
	LUT2 #(
		.INIT('h8)
	) name10935 (
		_w1978_,
		_w11396_,
		_w11397_
	);
	LUT2 #(
		.INIT('h1)
	) name10936 (
		_w11392_,
		_w11397_,
		_w11398_
	);
	LUT2 #(
		.INIT('h1)
	) name10937 (
		_w527_,
		_w3448_,
		_w11399_
	);
	LUT2 #(
		.INIT('h4)
	) name10938 (
		\P1_addr_reg[7]/NET0131 ,
		_w11399_,
		_w11400_
	);
	LUT2 #(
		.INIT('h1)
	) name10939 (
		_w1512_,
		_w11399_,
		_w11401_
	);
	LUT2 #(
		.INIT('h1)
	) name10940 (
		_w537_,
		_w11400_,
		_w11402_
	);
	LUT2 #(
		.INIT('h4)
	) name10941 (
		_w11401_,
		_w11402_,
		_w11403_
	);
	LUT2 #(
		.INIT('h4)
	) name10942 (
		_w527_,
		_w537_,
		_w11404_
	);
	LUT2 #(
		.INIT('h8)
	) name10943 (
		\P1_reg1_reg[7]/NET0131 ,
		_w1512_,
		_w11405_
	);
	LUT2 #(
		.INIT('h1)
	) name10944 (
		\P1_reg1_reg[7]/NET0131 ,
		_w1512_,
		_w11406_
	);
	LUT2 #(
		.INIT('h1)
	) name10945 (
		_w11405_,
		_w11406_,
		_w11407_
	);
	LUT2 #(
		.INIT('h2)
	) name10946 (
		\P1_reg1_reg[6]/NET0131 ,
		_w1535_,
		_w11408_
	);
	LUT2 #(
		.INIT('h4)
	) name10947 (
		\P1_reg1_reg[6]/NET0131 ,
		_w1535_,
		_w11409_
	);
	LUT2 #(
		.INIT('h2)
	) name10948 (
		\P1_reg1_reg[5]/NET0131 ,
		_w1560_,
		_w11410_
	);
	LUT2 #(
		.INIT('h2)
	) name10949 (
		\P1_reg1_reg[4]/NET0131 ,
		_w1584_,
		_w11411_
	);
	LUT2 #(
		.INIT('h4)
	) name10950 (
		\P1_reg1_reg[3]/NET0131 ,
		_w1621_,
		_w11412_
	);
	LUT2 #(
		.INIT('h2)
	) name10951 (
		\P1_reg1_reg[3]/NET0131 ,
		_w1621_,
		_w11413_
	);
	LUT2 #(
		.INIT('h1)
	) name10952 (
		\P1_reg1_reg[2]/NET0131 ,
		_w1607_,
		_w11414_
	);
	LUT2 #(
		.INIT('h8)
	) name10953 (
		\P1_reg1_reg[2]/NET0131 ,
		_w1607_,
		_w11415_
	);
	LUT2 #(
		.INIT('h1)
	) name10954 (
		\P1_reg1_reg[1]/NET0131 ,
		_w1645_,
		_w11416_
	);
	LUT2 #(
		.INIT('h8)
	) name10955 (
		\P1_reg1_reg[1]/NET0131 ,
		_w1645_,
		_w11417_
	);
	LUT2 #(
		.INIT('h8)
	) name10956 (
		\P1_IR_reg[0]/NET0131 ,
		\P1_reg1_reg[0]/NET0131 ,
		_w11418_
	);
	LUT2 #(
		.INIT('h1)
	) name10957 (
		_w11417_,
		_w11418_,
		_w11419_
	);
	LUT2 #(
		.INIT('h1)
	) name10958 (
		_w11416_,
		_w11419_,
		_w11420_
	);
	LUT2 #(
		.INIT('h1)
	) name10959 (
		_w11415_,
		_w11420_,
		_w11421_
	);
	LUT2 #(
		.INIT('h1)
	) name10960 (
		_w11414_,
		_w11421_,
		_w11422_
	);
	LUT2 #(
		.INIT('h1)
	) name10961 (
		_w11413_,
		_w11422_,
		_w11423_
	);
	LUT2 #(
		.INIT('h1)
	) name10962 (
		_w11412_,
		_w11423_,
		_w11424_
	);
	LUT2 #(
		.INIT('h1)
	) name10963 (
		_w11411_,
		_w11424_,
		_w11425_
	);
	LUT2 #(
		.INIT('h4)
	) name10964 (
		\P1_reg1_reg[5]/NET0131 ,
		_w1560_,
		_w11426_
	);
	LUT2 #(
		.INIT('h4)
	) name10965 (
		\P1_reg1_reg[4]/NET0131 ,
		_w1584_,
		_w11427_
	);
	LUT2 #(
		.INIT('h1)
	) name10966 (
		_w11426_,
		_w11427_,
		_w11428_
	);
	LUT2 #(
		.INIT('h4)
	) name10967 (
		_w11425_,
		_w11428_,
		_w11429_
	);
	LUT2 #(
		.INIT('h1)
	) name10968 (
		_w11410_,
		_w11429_,
		_w11430_
	);
	LUT2 #(
		.INIT('h1)
	) name10969 (
		_w11409_,
		_w11430_,
		_w11431_
	);
	LUT2 #(
		.INIT('h1)
	) name10970 (
		_w11408_,
		_w11431_,
		_w11432_
	);
	LUT2 #(
		.INIT('h4)
	) name10971 (
		_w11407_,
		_w11432_,
		_w11433_
	);
	LUT2 #(
		.INIT('h2)
	) name10972 (
		_w11407_,
		_w11432_,
		_w11434_
	);
	LUT2 #(
		.INIT('h2)
	) name10973 (
		_w11404_,
		_w11433_,
		_w11435_
	);
	LUT2 #(
		.INIT('h4)
	) name10974 (
		_w11434_,
		_w11435_,
		_w11436_
	);
	LUT2 #(
		.INIT('h8)
	) name10975 (
		_w527_,
		_w537_,
		_w11437_
	);
	LUT2 #(
		.INIT('h8)
	) name10976 (
		\P1_reg2_reg[7]/NET0131 ,
		_w1512_,
		_w11438_
	);
	LUT2 #(
		.INIT('h1)
	) name10977 (
		\P1_reg2_reg[7]/NET0131 ,
		_w1512_,
		_w11439_
	);
	LUT2 #(
		.INIT('h1)
	) name10978 (
		_w11438_,
		_w11439_,
		_w11440_
	);
	LUT2 #(
		.INIT('h2)
	) name10979 (
		\P1_reg2_reg[6]/NET0131 ,
		_w1535_,
		_w11441_
	);
	LUT2 #(
		.INIT('h4)
	) name10980 (
		\P1_reg2_reg[6]/NET0131 ,
		_w1535_,
		_w11442_
	);
	LUT2 #(
		.INIT('h2)
	) name10981 (
		\P1_reg2_reg[5]/NET0131 ,
		_w1560_,
		_w11443_
	);
	LUT2 #(
		.INIT('h2)
	) name10982 (
		\P1_reg2_reg[4]/NET0131 ,
		_w1584_,
		_w11444_
	);
	LUT2 #(
		.INIT('h4)
	) name10983 (
		\P1_reg2_reg[3]/NET0131 ,
		_w1621_,
		_w11445_
	);
	LUT2 #(
		.INIT('h2)
	) name10984 (
		\P1_reg2_reg[3]/NET0131 ,
		_w1621_,
		_w11446_
	);
	LUT2 #(
		.INIT('h1)
	) name10985 (
		\P1_reg2_reg[2]/NET0131 ,
		_w1607_,
		_w11447_
	);
	LUT2 #(
		.INIT('h8)
	) name10986 (
		\P1_reg2_reg[2]/NET0131 ,
		_w1607_,
		_w11448_
	);
	LUT2 #(
		.INIT('h1)
	) name10987 (
		\P1_reg2_reg[1]/NET0131 ,
		_w1645_,
		_w11449_
	);
	LUT2 #(
		.INIT('h8)
	) name10988 (
		\P1_reg2_reg[1]/NET0131 ,
		_w1645_,
		_w11450_
	);
	LUT2 #(
		.INIT('h8)
	) name10989 (
		\P1_IR_reg[0]/NET0131 ,
		\P1_reg2_reg[0]/NET0131 ,
		_w11451_
	);
	LUT2 #(
		.INIT('h1)
	) name10990 (
		_w11450_,
		_w11451_,
		_w11452_
	);
	LUT2 #(
		.INIT('h1)
	) name10991 (
		_w11449_,
		_w11452_,
		_w11453_
	);
	LUT2 #(
		.INIT('h1)
	) name10992 (
		_w11448_,
		_w11453_,
		_w11454_
	);
	LUT2 #(
		.INIT('h1)
	) name10993 (
		_w11447_,
		_w11454_,
		_w11455_
	);
	LUT2 #(
		.INIT('h1)
	) name10994 (
		_w11446_,
		_w11455_,
		_w11456_
	);
	LUT2 #(
		.INIT('h1)
	) name10995 (
		_w11445_,
		_w11456_,
		_w11457_
	);
	LUT2 #(
		.INIT('h1)
	) name10996 (
		_w11444_,
		_w11457_,
		_w11458_
	);
	LUT2 #(
		.INIT('h4)
	) name10997 (
		\P1_reg2_reg[5]/NET0131 ,
		_w1560_,
		_w11459_
	);
	LUT2 #(
		.INIT('h4)
	) name10998 (
		\P1_reg2_reg[4]/NET0131 ,
		_w1584_,
		_w11460_
	);
	LUT2 #(
		.INIT('h1)
	) name10999 (
		_w11459_,
		_w11460_,
		_w11461_
	);
	LUT2 #(
		.INIT('h4)
	) name11000 (
		_w11458_,
		_w11461_,
		_w11462_
	);
	LUT2 #(
		.INIT('h1)
	) name11001 (
		_w11443_,
		_w11462_,
		_w11463_
	);
	LUT2 #(
		.INIT('h1)
	) name11002 (
		_w11442_,
		_w11463_,
		_w11464_
	);
	LUT2 #(
		.INIT('h1)
	) name11003 (
		_w11441_,
		_w11464_,
		_w11465_
	);
	LUT2 #(
		.INIT('h4)
	) name11004 (
		_w11440_,
		_w11465_,
		_w11466_
	);
	LUT2 #(
		.INIT('h2)
	) name11005 (
		_w11440_,
		_w11465_,
		_w11467_
	);
	LUT2 #(
		.INIT('h2)
	) name11006 (
		_w11437_,
		_w11466_,
		_w11468_
	);
	LUT2 #(
		.INIT('h4)
	) name11007 (
		_w11467_,
		_w11468_,
		_w11469_
	);
	LUT2 #(
		.INIT('h1)
	) name11008 (
		_w11403_,
		_w11436_,
		_w11470_
	);
	LUT2 #(
		.INIT('h4)
	) name11009 (
		_w11469_,
		_w11470_,
		_w11471_
	);
	LUT2 #(
		.INIT('h2)
	) name11010 (
		\P1_state_reg[0]/NET0131 ,
		_w11471_,
		_w11472_
	);
	LUT2 #(
		.INIT('h1)
	) name11011 (
		_w9781_,
		_w11472_,
		_w11473_
	);
	LUT2 #(
		.INIT('h4)
	) name11012 (
		\P1_addr_reg[9]/NET0131 ,
		_w11399_,
		_w11474_
	);
	LUT2 #(
		.INIT('h1)
	) name11013 (
		_w1247_,
		_w11399_,
		_w11475_
	);
	LUT2 #(
		.INIT('h1)
	) name11014 (
		_w537_,
		_w11474_,
		_w11476_
	);
	LUT2 #(
		.INIT('h4)
	) name11015 (
		_w11475_,
		_w11476_,
		_w11477_
	);
	LUT2 #(
		.INIT('h1)
	) name11016 (
		\P1_reg1_reg[8]/NET0131 ,
		_w1271_,
		_w11478_
	);
	LUT2 #(
		.INIT('h1)
	) name11017 (
		_w11406_,
		_w11432_,
		_w11479_
	);
	LUT2 #(
		.INIT('h8)
	) name11018 (
		\P1_reg1_reg[8]/NET0131 ,
		_w1271_,
		_w11480_
	);
	LUT2 #(
		.INIT('h1)
	) name11019 (
		_w11405_,
		_w11480_,
		_w11481_
	);
	LUT2 #(
		.INIT('h4)
	) name11020 (
		_w11479_,
		_w11481_,
		_w11482_
	);
	LUT2 #(
		.INIT('h1)
	) name11021 (
		_w11478_,
		_w11482_,
		_w11483_
	);
	LUT2 #(
		.INIT('h8)
	) name11022 (
		\P1_reg1_reg[9]/NET0131 ,
		_w1247_,
		_w11484_
	);
	LUT2 #(
		.INIT('h1)
	) name11023 (
		\P1_reg1_reg[9]/NET0131 ,
		_w1247_,
		_w11485_
	);
	LUT2 #(
		.INIT('h1)
	) name11024 (
		_w11484_,
		_w11485_,
		_w11486_
	);
	LUT2 #(
		.INIT('h1)
	) name11025 (
		_w11483_,
		_w11486_,
		_w11487_
	);
	LUT2 #(
		.INIT('h8)
	) name11026 (
		_w11483_,
		_w11486_,
		_w11488_
	);
	LUT2 #(
		.INIT('h2)
	) name11027 (
		_w11404_,
		_w11487_,
		_w11489_
	);
	LUT2 #(
		.INIT('h4)
	) name11028 (
		_w11488_,
		_w11489_,
		_w11490_
	);
	LUT2 #(
		.INIT('h1)
	) name11029 (
		\P1_reg2_reg[9]/NET0131 ,
		_w1247_,
		_w11491_
	);
	LUT2 #(
		.INIT('h8)
	) name11030 (
		\P1_reg2_reg[9]/NET0131 ,
		_w1247_,
		_w11492_
	);
	LUT2 #(
		.INIT('h1)
	) name11031 (
		_w11491_,
		_w11492_,
		_w11493_
	);
	LUT2 #(
		.INIT('h1)
	) name11032 (
		\P1_reg2_reg[8]/NET0131 ,
		_w1271_,
		_w11494_
	);
	LUT2 #(
		.INIT('h1)
	) name11033 (
		_w11439_,
		_w11465_,
		_w11495_
	);
	LUT2 #(
		.INIT('h8)
	) name11034 (
		\P1_reg2_reg[8]/NET0131 ,
		_w1271_,
		_w11496_
	);
	LUT2 #(
		.INIT('h1)
	) name11035 (
		_w11438_,
		_w11496_,
		_w11497_
	);
	LUT2 #(
		.INIT('h4)
	) name11036 (
		_w11495_,
		_w11497_,
		_w11498_
	);
	LUT2 #(
		.INIT('h1)
	) name11037 (
		_w11494_,
		_w11498_,
		_w11499_
	);
	LUT2 #(
		.INIT('h1)
	) name11038 (
		_w11493_,
		_w11499_,
		_w11500_
	);
	LUT2 #(
		.INIT('h8)
	) name11039 (
		_w11493_,
		_w11499_,
		_w11501_
	);
	LUT2 #(
		.INIT('h2)
	) name11040 (
		_w11437_,
		_w11500_,
		_w11502_
	);
	LUT2 #(
		.INIT('h4)
	) name11041 (
		_w11501_,
		_w11502_,
		_w11503_
	);
	LUT2 #(
		.INIT('h1)
	) name11042 (
		_w11477_,
		_w11490_,
		_w11504_
	);
	LUT2 #(
		.INIT('h4)
	) name11043 (
		_w11503_,
		_w11504_,
		_w11505_
	);
	LUT2 #(
		.INIT('h2)
	) name11044 (
		\P1_state_reg[0]/NET0131 ,
		_w11505_,
		_w11506_
	);
	LUT2 #(
		.INIT('h1)
	) name11045 (
		_w7281_,
		_w11506_,
		_w11507_
	);
	LUT2 #(
		.INIT('h1)
	) name11046 (
		_w11408_,
		_w11409_,
		_w11508_
	);
	LUT2 #(
		.INIT('h2)
	) name11047 (
		_w11430_,
		_w11508_,
		_w11509_
	);
	LUT2 #(
		.INIT('h4)
	) name11048 (
		_w11430_,
		_w11508_,
		_w11510_
	);
	LUT2 #(
		.INIT('h2)
	) name11049 (
		_w11404_,
		_w11509_,
		_w11511_
	);
	LUT2 #(
		.INIT('h4)
	) name11050 (
		_w11510_,
		_w11511_,
		_w11512_
	);
	LUT2 #(
		.INIT('h1)
	) name11051 (
		_w11441_,
		_w11442_,
		_w11513_
	);
	LUT2 #(
		.INIT('h2)
	) name11052 (
		_w11463_,
		_w11513_,
		_w11514_
	);
	LUT2 #(
		.INIT('h4)
	) name11053 (
		_w11463_,
		_w11513_,
		_w11515_
	);
	LUT2 #(
		.INIT('h2)
	) name11054 (
		_w11437_,
		_w11514_,
		_w11516_
	);
	LUT2 #(
		.INIT('h4)
	) name11055 (
		_w11515_,
		_w11516_,
		_w11517_
	);
	LUT2 #(
		.INIT('h4)
	) name11056 (
		\P1_addr_reg[6]/NET0131 ,
		_w11399_,
		_w11518_
	);
	LUT2 #(
		.INIT('h2)
	) name11057 (
		_w1535_,
		_w11399_,
		_w11519_
	);
	LUT2 #(
		.INIT('h1)
	) name11058 (
		_w537_,
		_w11518_,
		_w11520_
	);
	LUT2 #(
		.INIT('h4)
	) name11059 (
		_w11519_,
		_w11520_,
		_w11521_
	);
	LUT2 #(
		.INIT('h1)
	) name11060 (
		_w11512_,
		_w11517_,
		_w11522_
	);
	LUT2 #(
		.INIT('h4)
	) name11061 (
		_w11521_,
		_w11522_,
		_w11523_
	);
	LUT2 #(
		.INIT('h2)
	) name11062 (
		\P1_state_reg[0]/NET0131 ,
		_w11523_,
		_w11524_
	);
	LUT2 #(
		.INIT('h1)
	) name11063 (
		_w9740_,
		_w11524_,
		_w11525_
	);
	LUT2 #(
		.INIT('h2)
	) name11064 (
		\P1_reg3_reg[2]/NET0131 ,
		\P1_state_reg[0]/NET0131 ,
		_w11526_
	);
	LUT2 #(
		.INIT('h2)
	) name11065 (
		_w527_,
		_w537_,
		_w11527_
	);
	LUT2 #(
		.INIT('h8)
	) name11066 (
		_w1607_,
		_w11527_,
		_w11528_
	);
	LUT2 #(
		.INIT('h1)
	) name11067 (
		\P1_addr_reg[2]/NET0131 ,
		_w3448_,
		_w11529_
	);
	LUT2 #(
		.INIT('h4)
	) name11068 (
		_w1607_,
		_w3448_,
		_w11530_
	);
	LUT2 #(
		.INIT('h2)
	) name11069 (
		_w538_,
		_w11529_,
		_w11531_
	);
	LUT2 #(
		.INIT('h4)
	) name11070 (
		_w11530_,
		_w11531_,
		_w11532_
	);
	LUT2 #(
		.INIT('h1)
	) name11071 (
		_w11447_,
		_w11448_,
		_w11533_
	);
	LUT2 #(
		.INIT('h1)
	) name11072 (
		_w11453_,
		_w11533_,
		_w11534_
	);
	LUT2 #(
		.INIT('h8)
	) name11073 (
		_w11453_,
		_w11533_,
		_w11535_
	);
	LUT2 #(
		.INIT('h1)
	) name11074 (
		_w11534_,
		_w11535_,
		_w11536_
	);
	LUT2 #(
		.INIT('h8)
	) name11075 (
		_w11437_,
		_w11536_,
		_w11537_
	);
	LUT2 #(
		.INIT('h1)
	) name11076 (
		_w11414_,
		_w11415_,
		_w11538_
	);
	LUT2 #(
		.INIT('h1)
	) name11077 (
		_w11420_,
		_w11538_,
		_w11539_
	);
	LUT2 #(
		.INIT('h8)
	) name11078 (
		_w11420_,
		_w11538_,
		_w11540_
	);
	LUT2 #(
		.INIT('h1)
	) name11079 (
		_w11539_,
		_w11540_,
		_w11541_
	);
	LUT2 #(
		.INIT('h8)
	) name11080 (
		_w11404_,
		_w11541_,
		_w11542_
	);
	LUT2 #(
		.INIT('h1)
	) name11081 (
		_w11528_,
		_w11537_,
		_w11543_
	);
	LUT2 #(
		.INIT('h4)
	) name11082 (
		_w11542_,
		_w11543_,
		_w11544_
	);
	LUT2 #(
		.INIT('h4)
	) name11083 (
		_w11532_,
		_w11544_,
		_w11545_
	);
	LUT2 #(
		.INIT('h2)
	) name11084 (
		\P1_state_reg[0]/NET0131 ,
		_w11545_,
		_w11546_
	);
	LUT2 #(
		.INIT('h1)
	) name11085 (
		_w11526_,
		_w11546_,
		_w11547_
	);
	LUT2 #(
		.INIT('h4)
	) name11086 (
		_w1621_,
		_w11527_,
		_w11548_
	);
	LUT2 #(
		.INIT('h1)
	) name11087 (
		\P1_addr_reg[3]/NET0131 ,
		_w3448_,
		_w11549_
	);
	LUT2 #(
		.INIT('h8)
	) name11088 (
		_w1621_,
		_w3448_,
		_w11550_
	);
	LUT2 #(
		.INIT('h2)
	) name11089 (
		_w538_,
		_w11549_,
		_w11551_
	);
	LUT2 #(
		.INIT('h4)
	) name11090 (
		_w11550_,
		_w11551_,
		_w11552_
	);
	LUT2 #(
		.INIT('h1)
	) name11091 (
		_w11412_,
		_w11413_,
		_w11553_
	);
	LUT2 #(
		.INIT('h1)
	) name11092 (
		_w11422_,
		_w11553_,
		_w11554_
	);
	LUT2 #(
		.INIT('h8)
	) name11093 (
		_w11422_,
		_w11553_,
		_w11555_
	);
	LUT2 #(
		.INIT('h1)
	) name11094 (
		_w11554_,
		_w11555_,
		_w11556_
	);
	LUT2 #(
		.INIT('h8)
	) name11095 (
		_w11404_,
		_w11556_,
		_w11557_
	);
	LUT2 #(
		.INIT('h1)
	) name11096 (
		_w11445_,
		_w11446_,
		_w11558_
	);
	LUT2 #(
		.INIT('h1)
	) name11097 (
		_w11455_,
		_w11558_,
		_w11559_
	);
	LUT2 #(
		.INIT('h8)
	) name11098 (
		_w11455_,
		_w11558_,
		_w11560_
	);
	LUT2 #(
		.INIT('h1)
	) name11099 (
		_w11559_,
		_w11560_,
		_w11561_
	);
	LUT2 #(
		.INIT('h8)
	) name11100 (
		_w11437_,
		_w11561_,
		_w11562_
	);
	LUT2 #(
		.INIT('h1)
	) name11101 (
		_w11548_,
		_w11557_,
		_w11563_
	);
	LUT2 #(
		.INIT('h4)
	) name11102 (
		_w11562_,
		_w11563_,
		_w11564_
	);
	LUT2 #(
		.INIT('h4)
	) name11103 (
		_w11552_,
		_w11564_,
		_w11565_
	);
	LUT2 #(
		.INIT('h2)
	) name11104 (
		\P1_state_reg[0]/NET0131 ,
		_w11565_,
		_w11566_
	);
	LUT2 #(
		.INIT('h1)
	) name11105 (
		_w9696_,
		_w11566_,
		_w11567_
	);
	LUT2 #(
		.INIT('h8)
	) name11106 (
		\P1_reg2_reg[13]/NET0131 ,
		_w1126_,
		_w11568_
	);
	LUT2 #(
		.INIT('h1)
	) name11107 (
		\P1_reg2_reg[13]/NET0131 ,
		_w1126_,
		_w11569_
	);
	LUT2 #(
		.INIT('h1)
	) name11108 (
		_w11568_,
		_w11569_,
		_w11570_
	);
	LUT2 #(
		.INIT('h1)
	) name11109 (
		\P1_reg2_reg[12]/NET0131 ,
		_w1154_,
		_w11571_
	);
	LUT2 #(
		.INIT('h1)
	) name11110 (
		\P1_reg2_reg[11]/NET0131 ,
		_w1188_,
		_w11572_
	);
	LUT2 #(
		.INIT('h1)
	) name11111 (
		\P1_reg2_reg[10]/NET0131 ,
		_w1223_,
		_w11573_
	);
	LUT2 #(
		.INIT('h4)
	) name11112 (
		_w11491_,
		_w11499_,
		_w11574_
	);
	LUT2 #(
		.INIT('h8)
	) name11113 (
		\P1_reg2_reg[10]/NET0131 ,
		_w1223_,
		_w11575_
	);
	LUT2 #(
		.INIT('h1)
	) name11114 (
		_w11492_,
		_w11575_,
		_w11576_
	);
	LUT2 #(
		.INIT('h4)
	) name11115 (
		_w11574_,
		_w11576_,
		_w11577_
	);
	LUT2 #(
		.INIT('h1)
	) name11116 (
		_w11573_,
		_w11577_,
		_w11578_
	);
	LUT2 #(
		.INIT('h4)
	) name11117 (
		_w11572_,
		_w11578_,
		_w11579_
	);
	LUT2 #(
		.INIT('h8)
	) name11118 (
		\P1_reg2_reg[12]/NET0131 ,
		_w1154_,
		_w11580_
	);
	LUT2 #(
		.INIT('h8)
	) name11119 (
		\P1_reg2_reg[11]/NET0131 ,
		_w1188_,
		_w11581_
	);
	LUT2 #(
		.INIT('h1)
	) name11120 (
		_w11580_,
		_w11581_,
		_w11582_
	);
	LUT2 #(
		.INIT('h4)
	) name11121 (
		_w11579_,
		_w11582_,
		_w11583_
	);
	LUT2 #(
		.INIT('h1)
	) name11122 (
		_w11571_,
		_w11583_,
		_w11584_
	);
	LUT2 #(
		.INIT('h1)
	) name11123 (
		_w11570_,
		_w11584_,
		_w11585_
	);
	LUT2 #(
		.INIT('h8)
	) name11124 (
		_w11570_,
		_w11584_,
		_w11586_
	);
	LUT2 #(
		.INIT('h2)
	) name11125 (
		_w11437_,
		_w11585_,
		_w11587_
	);
	LUT2 #(
		.INIT('h4)
	) name11126 (
		_w11586_,
		_w11587_,
		_w11588_
	);
	LUT2 #(
		.INIT('h4)
	) name11127 (
		\P1_addr_reg[13]/NET0131 ,
		_w11399_,
		_w11589_
	);
	LUT2 #(
		.INIT('h1)
	) name11128 (
		_w1126_,
		_w11399_,
		_w11590_
	);
	LUT2 #(
		.INIT('h1)
	) name11129 (
		_w537_,
		_w11589_,
		_w11591_
	);
	LUT2 #(
		.INIT('h4)
	) name11130 (
		_w11590_,
		_w11591_,
		_w11592_
	);
	LUT2 #(
		.INIT('h8)
	) name11131 (
		\P1_reg1_reg[13]/NET0131 ,
		_w1126_,
		_w11593_
	);
	LUT2 #(
		.INIT('h1)
	) name11132 (
		\P1_reg1_reg[13]/NET0131 ,
		_w1126_,
		_w11594_
	);
	LUT2 #(
		.INIT('h1)
	) name11133 (
		_w11593_,
		_w11594_,
		_w11595_
	);
	LUT2 #(
		.INIT('h1)
	) name11134 (
		\P1_reg1_reg[12]/NET0131 ,
		_w1154_,
		_w11596_
	);
	LUT2 #(
		.INIT('h1)
	) name11135 (
		\P1_reg1_reg[11]/NET0131 ,
		_w1188_,
		_w11597_
	);
	LUT2 #(
		.INIT('h1)
	) name11136 (
		\P1_reg1_reg[10]/NET0131 ,
		_w1223_,
		_w11598_
	);
	LUT2 #(
		.INIT('h2)
	) name11137 (
		_w11483_,
		_w11485_,
		_w11599_
	);
	LUT2 #(
		.INIT('h8)
	) name11138 (
		\P1_reg1_reg[10]/NET0131 ,
		_w1223_,
		_w11600_
	);
	LUT2 #(
		.INIT('h1)
	) name11139 (
		_w11484_,
		_w11600_,
		_w11601_
	);
	LUT2 #(
		.INIT('h4)
	) name11140 (
		_w11599_,
		_w11601_,
		_w11602_
	);
	LUT2 #(
		.INIT('h1)
	) name11141 (
		_w11598_,
		_w11602_,
		_w11603_
	);
	LUT2 #(
		.INIT('h4)
	) name11142 (
		_w11597_,
		_w11603_,
		_w11604_
	);
	LUT2 #(
		.INIT('h8)
	) name11143 (
		\P1_reg1_reg[12]/NET0131 ,
		_w1154_,
		_w11605_
	);
	LUT2 #(
		.INIT('h8)
	) name11144 (
		\P1_reg1_reg[11]/NET0131 ,
		_w1188_,
		_w11606_
	);
	LUT2 #(
		.INIT('h1)
	) name11145 (
		_w11605_,
		_w11606_,
		_w11607_
	);
	LUT2 #(
		.INIT('h4)
	) name11146 (
		_w11604_,
		_w11607_,
		_w11608_
	);
	LUT2 #(
		.INIT('h1)
	) name11147 (
		_w11596_,
		_w11608_,
		_w11609_
	);
	LUT2 #(
		.INIT('h1)
	) name11148 (
		_w11595_,
		_w11609_,
		_w11610_
	);
	LUT2 #(
		.INIT('h8)
	) name11149 (
		_w11595_,
		_w11609_,
		_w11611_
	);
	LUT2 #(
		.INIT('h2)
	) name11150 (
		_w11404_,
		_w11610_,
		_w11612_
	);
	LUT2 #(
		.INIT('h4)
	) name11151 (
		_w11611_,
		_w11612_,
		_w11613_
	);
	LUT2 #(
		.INIT('h1)
	) name11152 (
		_w11588_,
		_w11592_,
		_w11614_
	);
	LUT2 #(
		.INIT('h4)
	) name11153 (
		_w11613_,
		_w11614_,
		_w11615_
	);
	LUT2 #(
		.INIT('h2)
	) name11154 (
		\P1_state_reg[0]/NET0131 ,
		_w11615_,
		_w11616_
	);
	LUT2 #(
		.INIT('h1)
	) name11155 (
		_w7113_,
		_w11616_,
		_w11617_
	);
	LUT2 #(
		.INIT('h4)
	) name11156 (
		\P1_state_reg[0]/NET0131 ,
		\P2_reg3_reg[0]/NET0131 ,
		_w11618_
	);
	LUT2 #(
		.INIT('h2)
	) name11157 (
		_w2051_,
		_w2058_,
		_w11619_
	);
	LUT2 #(
		.INIT('h8)
	) name11158 (
		\P2_IR_reg[0]/NET0131 ,
		_w11619_,
		_w11620_
	);
	LUT2 #(
		.INIT('h1)
	) name11159 (
		\P2_addr_reg[0]/NET0131 ,
		_w2024_,
		_w11621_
	);
	LUT2 #(
		.INIT('h4)
	) name11160 (
		\P2_IR_reg[0]/NET0131 ,
		_w2024_,
		_w11622_
	);
	LUT2 #(
		.INIT('h2)
	) name11161 (
		_w2059_,
		_w11621_,
		_w11623_
	);
	LUT2 #(
		.INIT('h4)
	) name11162 (
		_w11622_,
		_w11623_,
		_w11624_
	);
	LUT2 #(
		.INIT('h1)
	) name11163 (
		\P2_IR_reg[0]/NET0131 ,
		\P2_reg1_reg[0]/NET0131 ,
		_w11625_
	);
	LUT2 #(
		.INIT('h4)
	) name11164 (
		_w2051_,
		_w2058_,
		_w11626_
	);
	LUT2 #(
		.INIT('h8)
	) name11165 (
		\P2_IR_reg[0]/NET0131 ,
		\P2_reg1_reg[0]/NET0131 ,
		_w11627_
	);
	LUT2 #(
		.INIT('h1)
	) name11166 (
		_w11625_,
		_w11627_,
		_w11628_
	);
	LUT2 #(
		.INIT('h8)
	) name11167 (
		_w11626_,
		_w11628_,
		_w11629_
	);
	LUT2 #(
		.INIT('h8)
	) name11168 (
		_w2051_,
		_w2058_,
		_w11630_
	);
	LUT2 #(
		.INIT('h1)
	) name11169 (
		\P2_IR_reg[0]/NET0131 ,
		\P2_reg2_reg[0]/NET0131 ,
		_w11631_
	);
	LUT2 #(
		.INIT('h8)
	) name11170 (
		\P2_IR_reg[0]/NET0131 ,
		\P2_reg2_reg[0]/NET0131 ,
		_w11632_
	);
	LUT2 #(
		.INIT('h1)
	) name11171 (
		_w11631_,
		_w11632_,
		_w11633_
	);
	LUT2 #(
		.INIT('h8)
	) name11172 (
		_w11630_,
		_w11633_,
		_w11634_
	);
	LUT2 #(
		.INIT('h1)
	) name11173 (
		_w11620_,
		_w11629_,
		_w11635_
	);
	LUT2 #(
		.INIT('h4)
	) name11174 (
		_w11634_,
		_w11635_,
		_w11636_
	);
	LUT2 #(
		.INIT('h4)
	) name11175 (
		_w11624_,
		_w11636_,
		_w11637_
	);
	LUT2 #(
		.INIT('h2)
	) name11176 (
		\P1_state_reg[0]/NET0131 ,
		_w11637_,
		_w11638_
	);
	LUT2 #(
		.INIT('h1)
	) name11177 (
		_w11618_,
		_w11638_,
		_w11639_
	);
	LUT2 #(
		.INIT('h2)
	) name11178 (
		\P1_reg3_reg[0]/NET0131 ,
		\P1_state_reg[0]/NET0131 ,
		_w11640_
	);
	LUT2 #(
		.INIT('h8)
	) name11179 (
		\P1_IR_reg[0]/NET0131 ,
		_w11527_,
		_w11641_
	);
	LUT2 #(
		.INIT('h1)
	) name11180 (
		\P1_addr_reg[0]/NET0131 ,
		_w3448_,
		_w11642_
	);
	LUT2 #(
		.INIT('h4)
	) name11181 (
		\P1_IR_reg[0]/NET0131 ,
		_w3448_,
		_w11643_
	);
	LUT2 #(
		.INIT('h2)
	) name11182 (
		_w538_,
		_w11642_,
		_w11644_
	);
	LUT2 #(
		.INIT('h4)
	) name11183 (
		_w11643_,
		_w11644_,
		_w11645_
	);
	LUT2 #(
		.INIT('h1)
	) name11184 (
		\P1_IR_reg[0]/NET0131 ,
		\P1_reg1_reg[0]/NET0131 ,
		_w11646_
	);
	LUT2 #(
		.INIT('h1)
	) name11185 (
		_w11418_,
		_w11646_,
		_w11647_
	);
	LUT2 #(
		.INIT('h8)
	) name11186 (
		_w11404_,
		_w11647_,
		_w11648_
	);
	LUT2 #(
		.INIT('h1)
	) name11187 (
		\P1_IR_reg[0]/NET0131 ,
		\P1_reg2_reg[0]/NET0131 ,
		_w11649_
	);
	LUT2 #(
		.INIT('h1)
	) name11188 (
		_w11451_,
		_w11649_,
		_w11650_
	);
	LUT2 #(
		.INIT('h8)
	) name11189 (
		_w11437_,
		_w11650_,
		_w11651_
	);
	LUT2 #(
		.INIT('h1)
	) name11190 (
		_w11641_,
		_w11648_,
		_w11652_
	);
	LUT2 #(
		.INIT('h4)
	) name11191 (
		_w11651_,
		_w11652_,
		_w11653_
	);
	LUT2 #(
		.INIT('h4)
	) name11192 (
		_w11645_,
		_w11653_,
		_w11654_
	);
	LUT2 #(
		.INIT('h2)
	) name11193 (
		\P1_state_reg[0]/NET0131 ,
		_w11654_,
		_w11655_
	);
	LUT2 #(
		.INIT('h1)
	) name11194 (
		_w11640_,
		_w11655_,
		_w11656_
	);
	LUT2 #(
		.INIT('h4)
	) name11195 (
		\P1_addr_reg[10]/NET0131 ,
		_w11399_,
		_w11657_
	);
	LUT2 #(
		.INIT('h1)
	) name11196 (
		_w1223_,
		_w11399_,
		_w11658_
	);
	LUT2 #(
		.INIT('h1)
	) name11197 (
		_w537_,
		_w11657_,
		_w11659_
	);
	LUT2 #(
		.INIT('h4)
	) name11198 (
		_w11658_,
		_w11659_,
		_w11660_
	);
	LUT2 #(
		.INIT('h1)
	) name11199 (
		_w11598_,
		_w11600_,
		_w11661_
	);
	LUT2 #(
		.INIT('h1)
	) name11200 (
		_w11405_,
		_w11479_,
		_w11662_
	);
	LUT2 #(
		.INIT('h1)
	) name11201 (
		_w11478_,
		_w11662_,
		_w11663_
	);
	LUT2 #(
		.INIT('h1)
	) name11202 (
		_w11480_,
		_w11484_,
		_w11664_
	);
	LUT2 #(
		.INIT('h4)
	) name11203 (
		_w11663_,
		_w11664_,
		_w11665_
	);
	LUT2 #(
		.INIT('h1)
	) name11204 (
		_w11485_,
		_w11665_,
		_w11666_
	);
	LUT2 #(
		.INIT('h1)
	) name11205 (
		_w11661_,
		_w11666_,
		_w11667_
	);
	LUT2 #(
		.INIT('h8)
	) name11206 (
		_w11661_,
		_w11666_,
		_w11668_
	);
	LUT2 #(
		.INIT('h2)
	) name11207 (
		_w11404_,
		_w11667_,
		_w11669_
	);
	LUT2 #(
		.INIT('h4)
	) name11208 (
		_w11668_,
		_w11669_,
		_w11670_
	);
	LUT2 #(
		.INIT('h1)
	) name11209 (
		_w11573_,
		_w11575_,
		_w11671_
	);
	LUT2 #(
		.INIT('h1)
	) name11210 (
		_w11438_,
		_w11495_,
		_w11672_
	);
	LUT2 #(
		.INIT('h1)
	) name11211 (
		_w11494_,
		_w11672_,
		_w11673_
	);
	LUT2 #(
		.INIT('h1)
	) name11212 (
		_w11492_,
		_w11496_,
		_w11674_
	);
	LUT2 #(
		.INIT('h4)
	) name11213 (
		_w11673_,
		_w11674_,
		_w11675_
	);
	LUT2 #(
		.INIT('h1)
	) name11214 (
		_w11491_,
		_w11675_,
		_w11676_
	);
	LUT2 #(
		.INIT('h1)
	) name11215 (
		_w11671_,
		_w11676_,
		_w11677_
	);
	LUT2 #(
		.INIT('h8)
	) name11216 (
		_w11671_,
		_w11676_,
		_w11678_
	);
	LUT2 #(
		.INIT('h2)
	) name11217 (
		_w11437_,
		_w11677_,
		_w11679_
	);
	LUT2 #(
		.INIT('h4)
	) name11218 (
		_w11678_,
		_w11679_,
		_w11680_
	);
	LUT2 #(
		.INIT('h1)
	) name11219 (
		_w11660_,
		_w11670_,
		_w11681_
	);
	LUT2 #(
		.INIT('h4)
	) name11220 (
		_w11680_,
		_w11681_,
		_w11682_
	);
	LUT2 #(
		.INIT('h2)
	) name11221 (
		\P1_state_reg[0]/NET0131 ,
		_w11682_,
		_w11683_
	);
	LUT2 #(
		.INIT('h1)
	) name11222 (
		_w7071_,
		_w11683_,
		_w11684_
	);
	LUT2 #(
		.INIT('h4)
	) name11223 (
		\P1_addr_reg[11]/NET0131 ,
		_w11399_,
		_w11685_
	);
	LUT2 #(
		.INIT('h1)
	) name11224 (
		_w1188_,
		_w11399_,
		_w11686_
	);
	LUT2 #(
		.INIT('h1)
	) name11225 (
		_w537_,
		_w11685_,
		_w11687_
	);
	LUT2 #(
		.INIT('h4)
	) name11226 (
		_w11686_,
		_w11687_,
		_w11688_
	);
	LUT2 #(
		.INIT('h1)
	) name11227 (
		_w11597_,
		_w11606_,
		_w11689_
	);
	LUT2 #(
		.INIT('h1)
	) name11228 (
		_w11603_,
		_w11689_,
		_w11690_
	);
	LUT2 #(
		.INIT('h8)
	) name11229 (
		_w11603_,
		_w11689_,
		_w11691_
	);
	LUT2 #(
		.INIT('h2)
	) name11230 (
		_w11404_,
		_w11690_,
		_w11692_
	);
	LUT2 #(
		.INIT('h4)
	) name11231 (
		_w11691_,
		_w11692_,
		_w11693_
	);
	LUT2 #(
		.INIT('h1)
	) name11232 (
		_w11572_,
		_w11581_,
		_w11694_
	);
	LUT2 #(
		.INIT('h1)
	) name11233 (
		_w11578_,
		_w11694_,
		_w11695_
	);
	LUT2 #(
		.INIT('h8)
	) name11234 (
		_w11578_,
		_w11694_,
		_w11696_
	);
	LUT2 #(
		.INIT('h2)
	) name11235 (
		_w11437_,
		_w11695_,
		_w11697_
	);
	LUT2 #(
		.INIT('h4)
	) name11236 (
		_w11696_,
		_w11697_,
		_w11698_
	);
	LUT2 #(
		.INIT('h1)
	) name11237 (
		_w11688_,
		_w11693_,
		_w11699_
	);
	LUT2 #(
		.INIT('h4)
	) name11238 (
		_w11698_,
		_w11699_,
		_w11700_
	);
	LUT2 #(
		.INIT('h2)
	) name11239 (
		\P1_state_reg[0]/NET0131 ,
		_w11700_,
		_w11701_
	);
	LUT2 #(
		.INIT('h1)
	) name11240 (
		_w7997_,
		_w11701_,
		_w11702_
	);
	LUT2 #(
		.INIT('h4)
	) name11241 (
		\P1_addr_reg[12]/NET0131 ,
		_w11399_,
		_w11703_
	);
	LUT2 #(
		.INIT('h1)
	) name11242 (
		_w1154_,
		_w11399_,
		_w11704_
	);
	LUT2 #(
		.INIT('h1)
	) name11243 (
		_w537_,
		_w11703_,
		_w11705_
	);
	LUT2 #(
		.INIT('h4)
	) name11244 (
		_w11704_,
		_w11705_,
		_w11706_
	);
	LUT2 #(
		.INIT('h1)
	) name11245 (
		_w11596_,
		_w11605_,
		_w11707_
	);
	LUT2 #(
		.INIT('h4)
	) name11246 (
		_w11598_,
		_w11666_,
		_w11708_
	);
	LUT2 #(
		.INIT('h1)
	) name11247 (
		_w11600_,
		_w11606_,
		_w11709_
	);
	LUT2 #(
		.INIT('h4)
	) name11248 (
		_w11708_,
		_w11709_,
		_w11710_
	);
	LUT2 #(
		.INIT('h1)
	) name11249 (
		_w11597_,
		_w11710_,
		_w11711_
	);
	LUT2 #(
		.INIT('h1)
	) name11250 (
		_w11707_,
		_w11711_,
		_w11712_
	);
	LUT2 #(
		.INIT('h8)
	) name11251 (
		_w11707_,
		_w11711_,
		_w11713_
	);
	LUT2 #(
		.INIT('h2)
	) name11252 (
		_w11404_,
		_w11712_,
		_w11714_
	);
	LUT2 #(
		.INIT('h4)
	) name11253 (
		_w11713_,
		_w11714_,
		_w11715_
	);
	LUT2 #(
		.INIT('h1)
	) name11254 (
		_w11571_,
		_w11580_,
		_w11716_
	);
	LUT2 #(
		.INIT('h4)
	) name11255 (
		_w11573_,
		_w11676_,
		_w11717_
	);
	LUT2 #(
		.INIT('h1)
	) name11256 (
		_w11575_,
		_w11581_,
		_w11718_
	);
	LUT2 #(
		.INIT('h4)
	) name11257 (
		_w11717_,
		_w11718_,
		_w11719_
	);
	LUT2 #(
		.INIT('h1)
	) name11258 (
		_w11572_,
		_w11719_,
		_w11720_
	);
	LUT2 #(
		.INIT('h1)
	) name11259 (
		_w11716_,
		_w11720_,
		_w11721_
	);
	LUT2 #(
		.INIT('h8)
	) name11260 (
		_w11716_,
		_w11720_,
		_w11722_
	);
	LUT2 #(
		.INIT('h2)
	) name11261 (
		_w11437_,
		_w11721_,
		_w11723_
	);
	LUT2 #(
		.INIT('h4)
	) name11262 (
		_w11722_,
		_w11723_,
		_w11724_
	);
	LUT2 #(
		.INIT('h1)
	) name11263 (
		_w11706_,
		_w11715_,
		_w11725_
	);
	LUT2 #(
		.INIT('h4)
	) name11264 (
		_w11724_,
		_w11725_,
		_w11726_
	);
	LUT2 #(
		.INIT('h2)
	) name11265 (
		\P1_state_reg[0]/NET0131 ,
		_w11726_,
		_w11727_
	);
	LUT2 #(
		.INIT('h1)
	) name11266 (
		_w6089_,
		_w11727_,
		_w11728_
	);
	LUT2 #(
		.INIT('h1)
	) name11267 (
		_w2024_,
		_w2051_,
		_w11729_
	);
	LUT2 #(
		.INIT('h4)
	) name11268 (
		\P2_addr_reg[10]/NET0131 ,
		_w11729_,
		_w11730_
	);
	LUT2 #(
		.INIT('h2)
	) name11269 (
		_w2745_,
		_w11729_,
		_w11731_
	);
	LUT2 #(
		.INIT('h1)
	) name11270 (
		_w2058_,
		_w11730_,
		_w11732_
	);
	LUT2 #(
		.INIT('h4)
	) name11271 (
		_w11731_,
		_w11732_,
		_w11733_
	);
	LUT2 #(
		.INIT('h2)
	) name11272 (
		\P2_reg1_reg[10]/NET0131 ,
		_w2745_,
		_w11734_
	);
	LUT2 #(
		.INIT('h4)
	) name11273 (
		\P2_reg1_reg[10]/NET0131 ,
		_w2745_,
		_w11735_
	);
	LUT2 #(
		.INIT('h1)
	) name11274 (
		_w11734_,
		_w11735_,
		_w11736_
	);
	LUT2 #(
		.INIT('h2)
	) name11275 (
		\P2_reg1_reg[9]/NET0131 ,
		_w2769_,
		_w11737_
	);
	LUT2 #(
		.INIT('h4)
	) name11276 (
		\P2_reg1_reg[9]/NET0131 ,
		_w2769_,
		_w11738_
	);
	LUT2 #(
		.INIT('h1)
	) name11277 (
		\P2_reg1_reg[8]/NET0131 ,
		_w2460_,
		_w11739_
	);
	LUT2 #(
		.INIT('h1)
	) name11278 (
		_w11738_,
		_w11739_,
		_w11740_
	);
	LUT2 #(
		.INIT('h8)
	) name11279 (
		\P2_reg1_reg[8]/NET0131 ,
		_w2460_,
		_w11741_
	);
	LUT2 #(
		.INIT('h1)
	) name11280 (
		\P2_reg1_reg[7]/NET0131 ,
		_w2485_,
		_w11742_
	);
	LUT2 #(
		.INIT('h8)
	) name11281 (
		\P2_reg1_reg[6]/NET0131 ,
		_w2519_,
		_w11743_
	);
	LUT2 #(
		.INIT('h1)
	) name11282 (
		\P2_reg1_reg[6]/NET0131 ,
		_w2519_,
		_w11744_
	);
	LUT2 #(
		.INIT('h2)
	) name11283 (
		\P2_reg1_reg[5]/NET0131 ,
		_w2542_,
		_w11745_
	);
	LUT2 #(
		.INIT('h4)
	) name11284 (
		\P2_reg1_reg[5]/NET0131 ,
		_w2542_,
		_w11746_
	);
	LUT2 #(
		.INIT('h1)
	) name11285 (
		\P2_reg1_reg[4]/NET0131 ,
		_w2646_,
		_w11747_
	);
	LUT2 #(
		.INIT('h1)
	) name11286 (
		\P2_reg1_reg[3]/NET0131 ,
		_w2629_,
		_w11748_
	);
	LUT2 #(
		.INIT('h1)
	) name11287 (
		\P2_reg1_reg[2]/NET0131 ,
		_w2564_,
		_w11749_
	);
	LUT2 #(
		.INIT('h8)
	) name11288 (
		\P2_reg1_reg[2]/NET0131 ,
		_w2564_,
		_w11750_
	);
	LUT2 #(
		.INIT('h1)
	) name11289 (
		\P2_reg1_reg[1]/NET0131 ,
		_w2578_,
		_w11751_
	);
	LUT2 #(
		.INIT('h8)
	) name11290 (
		\P2_reg1_reg[1]/NET0131 ,
		_w2578_,
		_w11752_
	);
	LUT2 #(
		.INIT('h1)
	) name11291 (
		_w11627_,
		_w11752_,
		_w11753_
	);
	LUT2 #(
		.INIT('h1)
	) name11292 (
		_w11751_,
		_w11753_,
		_w11754_
	);
	LUT2 #(
		.INIT('h1)
	) name11293 (
		_w11750_,
		_w11754_,
		_w11755_
	);
	LUT2 #(
		.INIT('h1)
	) name11294 (
		_w11749_,
		_w11755_,
		_w11756_
	);
	LUT2 #(
		.INIT('h4)
	) name11295 (
		_w11748_,
		_w11756_,
		_w11757_
	);
	LUT2 #(
		.INIT('h8)
	) name11296 (
		\P2_reg1_reg[4]/NET0131 ,
		_w2646_,
		_w11758_
	);
	LUT2 #(
		.INIT('h8)
	) name11297 (
		\P2_reg1_reg[3]/NET0131 ,
		_w2629_,
		_w11759_
	);
	LUT2 #(
		.INIT('h1)
	) name11298 (
		_w11758_,
		_w11759_,
		_w11760_
	);
	LUT2 #(
		.INIT('h4)
	) name11299 (
		_w11757_,
		_w11760_,
		_w11761_
	);
	LUT2 #(
		.INIT('h1)
	) name11300 (
		_w11747_,
		_w11761_,
		_w11762_
	);
	LUT2 #(
		.INIT('h4)
	) name11301 (
		_w11746_,
		_w11762_,
		_w11763_
	);
	LUT2 #(
		.INIT('h1)
	) name11302 (
		_w11745_,
		_w11763_,
		_w11764_
	);
	LUT2 #(
		.INIT('h1)
	) name11303 (
		_w11744_,
		_w11764_,
		_w11765_
	);
	LUT2 #(
		.INIT('h8)
	) name11304 (
		\P2_reg1_reg[7]/NET0131 ,
		_w2485_,
		_w11766_
	);
	LUT2 #(
		.INIT('h1)
	) name11305 (
		_w11743_,
		_w11766_,
		_w11767_
	);
	LUT2 #(
		.INIT('h4)
	) name11306 (
		_w11765_,
		_w11767_,
		_w11768_
	);
	LUT2 #(
		.INIT('h1)
	) name11307 (
		_w11742_,
		_w11768_,
		_w11769_
	);
	LUT2 #(
		.INIT('h1)
	) name11308 (
		_w11741_,
		_w11769_,
		_w11770_
	);
	LUT2 #(
		.INIT('h2)
	) name11309 (
		_w11740_,
		_w11770_,
		_w11771_
	);
	LUT2 #(
		.INIT('h1)
	) name11310 (
		_w11737_,
		_w11771_,
		_w11772_
	);
	LUT2 #(
		.INIT('h4)
	) name11311 (
		_w11736_,
		_w11772_,
		_w11773_
	);
	LUT2 #(
		.INIT('h2)
	) name11312 (
		_w11736_,
		_w11772_,
		_w11774_
	);
	LUT2 #(
		.INIT('h2)
	) name11313 (
		_w11626_,
		_w11773_,
		_w11775_
	);
	LUT2 #(
		.INIT('h4)
	) name11314 (
		_w11774_,
		_w11775_,
		_w11776_
	);
	LUT2 #(
		.INIT('h2)
	) name11315 (
		\P2_reg2_reg[10]/NET0131 ,
		_w2745_,
		_w11777_
	);
	LUT2 #(
		.INIT('h4)
	) name11316 (
		\P2_reg2_reg[10]/NET0131 ,
		_w2745_,
		_w11778_
	);
	LUT2 #(
		.INIT('h1)
	) name11317 (
		_w11777_,
		_w11778_,
		_w11779_
	);
	LUT2 #(
		.INIT('h2)
	) name11318 (
		\P2_reg2_reg[9]/NET0131 ,
		_w2769_,
		_w11780_
	);
	LUT2 #(
		.INIT('h4)
	) name11319 (
		\P2_reg2_reg[9]/NET0131 ,
		_w2769_,
		_w11781_
	);
	LUT2 #(
		.INIT('h1)
	) name11320 (
		\P2_reg2_reg[8]/NET0131 ,
		_w2460_,
		_w11782_
	);
	LUT2 #(
		.INIT('h1)
	) name11321 (
		_w11781_,
		_w11782_,
		_w11783_
	);
	LUT2 #(
		.INIT('h8)
	) name11322 (
		\P2_reg2_reg[8]/NET0131 ,
		_w2460_,
		_w11784_
	);
	LUT2 #(
		.INIT('h1)
	) name11323 (
		\P2_reg2_reg[7]/NET0131 ,
		_w2485_,
		_w11785_
	);
	LUT2 #(
		.INIT('h8)
	) name11324 (
		\P2_reg2_reg[6]/NET0131 ,
		_w2519_,
		_w11786_
	);
	LUT2 #(
		.INIT('h1)
	) name11325 (
		\P2_reg2_reg[6]/NET0131 ,
		_w2519_,
		_w11787_
	);
	LUT2 #(
		.INIT('h2)
	) name11326 (
		\P2_reg2_reg[5]/NET0131 ,
		_w2542_,
		_w11788_
	);
	LUT2 #(
		.INIT('h4)
	) name11327 (
		\P2_reg2_reg[5]/NET0131 ,
		_w2542_,
		_w11789_
	);
	LUT2 #(
		.INIT('h1)
	) name11328 (
		\P2_reg2_reg[4]/NET0131 ,
		_w2646_,
		_w11790_
	);
	LUT2 #(
		.INIT('h8)
	) name11329 (
		\P2_reg2_reg[4]/NET0131 ,
		_w2646_,
		_w11791_
	);
	LUT2 #(
		.INIT('h1)
	) name11330 (
		\P2_reg2_reg[3]/NET0131 ,
		_w2629_,
		_w11792_
	);
	LUT2 #(
		.INIT('h8)
	) name11331 (
		\P2_reg2_reg[3]/NET0131 ,
		_w2629_,
		_w11793_
	);
	LUT2 #(
		.INIT('h1)
	) name11332 (
		\P2_reg2_reg[2]/NET0131 ,
		_w2564_,
		_w11794_
	);
	LUT2 #(
		.INIT('h8)
	) name11333 (
		\P2_reg2_reg[2]/NET0131 ,
		_w2564_,
		_w11795_
	);
	LUT2 #(
		.INIT('h1)
	) name11334 (
		\P2_reg2_reg[1]/NET0131 ,
		_w2578_,
		_w11796_
	);
	LUT2 #(
		.INIT('h8)
	) name11335 (
		\P2_reg2_reg[1]/NET0131 ,
		_w2578_,
		_w11797_
	);
	LUT2 #(
		.INIT('h1)
	) name11336 (
		_w11632_,
		_w11797_,
		_w11798_
	);
	LUT2 #(
		.INIT('h1)
	) name11337 (
		_w11796_,
		_w11798_,
		_w11799_
	);
	LUT2 #(
		.INIT('h1)
	) name11338 (
		_w11795_,
		_w11799_,
		_w11800_
	);
	LUT2 #(
		.INIT('h1)
	) name11339 (
		_w11794_,
		_w11800_,
		_w11801_
	);
	LUT2 #(
		.INIT('h1)
	) name11340 (
		_w11793_,
		_w11801_,
		_w11802_
	);
	LUT2 #(
		.INIT('h1)
	) name11341 (
		_w11792_,
		_w11802_,
		_w11803_
	);
	LUT2 #(
		.INIT('h1)
	) name11342 (
		_w11791_,
		_w11803_,
		_w11804_
	);
	LUT2 #(
		.INIT('h1)
	) name11343 (
		_w11790_,
		_w11804_,
		_w11805_
	);
	LUT2 #(
		.INIT('h4)
	) name11344 (
		_w11789_,
		_w11805_,
		_w11806_
	);
	LUT2 #(
		.INIT('h1)
	) name11345 (
		_w11788_,
		_w11806_,
		_w11807_
	);
	LUT2 #(
		.INIT('h1)
	) name11346 (
		_w11787_,
		_w11807_,
		_w11808_
	);
	LUT2 #(
		.INIT('h8)
	) name11347 (
		\P2_reg2_reg[7]/NET0131 ,
		_w2485_,
		_w11809_
	);
	LUT2 #(
		.INIT('h1)
	) name11348 (
		_w11786_,
		_w11809_,
		_w11810_
	);
	LUT2 #(
		.INIT('h4)
	) name11349 (
		_w11808_,
		_w11810_,
		_w11811_
	);
	LUT2 #(
		.INIT('h1)
	) name11350 (
		_w11785_,
		_w11811_,
		_w11812_
	);
	LUT2 #(
		.INIT('h1)
	) name11351 (
		_w11784_,
		_w11812_,
		_w11813_
	);
	LUT2 #(
		.INIT('h2)
	) name11352 (
		_w11783_,
		_w11813_,
		_w11814_
	);
	LUT2 #(
		.INIT('h1)
	) name11353 (
		_w11780_,
		_w11814_,
		_w11815_
	);
	LUT2 #(
		.INIT('h4)
	) name11354 (
		_w11779_,
		_w11815_,
		_w11816_
	);
	LUT2 #(
		.INIT('h2)
	) name11355 (
		_w11779_,
		_w11815_,
		_w11817_
	);
	LUT2 #(
		.INIT('h2)
	) name11356 (
		_w11630_,
		_w11816_,
		_w11818_
	);
	LUT2 #(
		.INIT('h4)
	) name11357 (
		_w11817_,
		_w11818_,
		_w11819_
	);
	LUT2 #(
		.INIT('h1)
	) name11358 (
		_w11733_,
		_w11776_,
		_w11820_
	);
	LUT2 #(
		.INIT('h4)
	) name11359 (
		_w11819_,
		_w11820_,
		_w11821_
	);
	LUT2 #(
		.INIT('h2)
	) name11360 (
		\P1_state_reg[0]/NET0131 ,
		_w11821_,
		_w11822_
	);
	LUT2 #(
		.INIT('h1)
	) name11361 (
		_w7154_,
		_w11822_,
		_w11823_
	);
	LUT2 #(
		.INIT('h4)
	) name11362 (
		\P1_addr_reg[14]/NET0131 ,
		_w11399_,
		_w11824_
	);
	LUT2 #(
		.INIT('h1)
	) name11363 (
		_w1099_,
		_w11399_,
		_w11825_
	);
	LUT2 #(
		.INIT('h1)
	) name11364 (
		_w537_,
		_w11824_,
		_w11826_
	);
	LUT2 #(
		.INIT('h4)
	) name11365 (
		_w11825_,
		_w11826_,
		_w11827_
	);
	LUT2 #(
		.INIT('h8)
	) name11366 (
		\P1_reg1_reg[14]/NET0131 ,
		_w1099_,
		_w11828_
	);
	LUT2 #(
		.INIT('h1)
	) name11367 (
		\P1_reg1_reg[14]/NET0131 ,
		_w1099_,
		_w11829_
	);
	LUT2 #(
		.INIT('h1)
	) name11368 (
		_w11828_,
		_w11829_,
		_w11830_
	);
	LUT2 #(
		.INIT('h4)
	) name11369 (
		_w11596_,
		_w11711_,
		_w11831_
	);
	LUT2 #(
		.INIT('h1)
	) name11370 (
		_w11593_,
		_w11605_,
		_w11832_
	);
	LUT2 #(
		.INIT('h4)
	) name11371 (
		_w11831_,
		_w11832_,
		_w11833_
	);
	LUT2 #(
		.INIT('h1)
	) name11372 (
		_w11594_,
		_w11833_,
		_w11834_
	);
	LUT2 #(
		.INIT('h1)
	) name11373 (
		_w11830_,
		_w11834_,
		_w11835_
	);
	LUT2 #(
		.INIT('h8)
	) name11374 (
		_w11830_,
		_w11834_,
		_w11836_
	);
	LUT2 #(
		.INIT('h2)
	) name11375 (
		_w11404_,
		_w11835_,
		_w11837_
	);
	LUT2 #(
		.INIT('h4)
	) name11376 (
		_w11836_,
		_w11837_,
		_w11838_
	);
	LUT2 #(
		.INIT('h8)
	) name11377 (
		\P1_reg2_reg[14]/NET0131 ,
		_w1099_,
		_w11839_
	);
	LUT2 #(
		.INIT('h1)
	) name11378 (
		\P1_reg2_reg[14]/NET0131 ,
		_w1099_,
		_w11840_
	);
	LUT2 #(
		.INIT('h1)
	) name11379 (
		_w11839_,
		_w11840_,
		_w11841_
	);
	LUT2 #(
		.INIT('h4)
	) name11380 (
		_w11571_,
		_w11720_,
		_w11842_
	);
	LUT2 #(
		.INIT('h1)
	) name11381 (
		_w11568_,
		_w11580_,
		_w11843_
	);
	LUT2 #(
		.INIT('h4)
	) name11382 (
		_w11842_,
		_w11843_,
		_w11844_
	);
	LUT2 #(
		.INIT('h1)
	) name11383 (
		_w11569_,
		_w11844_,
		_w11845_
	);
	LUT2 #(
		.INIT('h1)
	) name11384 (
		_w11841_,
		_w11845_,
		_w11846_
	);
	LUT2 #(
		.INIT('h8)
	) name11385 (
		_w11841_,
		_w11845_,
		_w11847_
	);
	LUT2 #(
		.INIT('h2)
	) name11386 (
		_w11437_,
		_w11846_,
		_w11848_
	);
	LUT2 #(
		.INIT('h4)
	) name11387 (
		_w11847_,
		_w11848_,
		_w11849_
	);
	LUT2 #(
		.INIT('h1)
	) name11388 (
		_w11827_,
		_w11838_,
		_w11850_
	);
	LUT2 #(
		.INIT('h4)
	) name11389 (
		_w11849_,
		_w11850_,
		_w11851_
	);
	LUT2 #(
		.INIT('h2)
	) name11390 (
		\P1_state_reg[0]/NET0131 ,
		_w11851_,
		_w11852_
	);
	LUT2 #(
		.INIT('h1)
	) name11391 (
		_w8038_,
		_w11852_,
		_w11853_
	);
	LUT2 #(
		.INIT('h4)
	) name11392 (
		\P2_addr_reg[11]/NET0131 ,
		_w11729_,
		_w11854_
	);
	LUT2 #(
		.INIT('h1)
	) name11393 (
		_w2694_,
		_w11729_,
		_w11855_
	);
	LUT2 #(
		.INIT('h1)
	) name11394 (
		_w2058_,
		_w11854_,
		_w11856_
	);
	LUT2 #(
		.INIT('h4)
	) name11395 (
		_w11855_,
		_w11856_,
		_w11857_
	);
	LUT2 #(
		.INIT('h1)
	) name11396 (
		\P2_reg1_reg[11]/NET0131 ,
		_w2694_,
		_w11858_
	);
	LUT2 #(
		.INIT('h8)
	) name11397 (
		\P2_reg1_reg[11]/NET0131 ,
		_w2694_,
		_w11859_
	);
	LUT2 #(
		.INIT('h1)
	) name11398 (
		_w11858_,
		_w11859_,
		_w11860_
	);
	LUT2 #(
		.INIT('h1)
	) name11399 (
		_w11743_,
		_w11745_,
		_w11861_
	);
	LUT2 #(
		.INIT('h4)
	) name11400 (
		_w11763_,
		_w11861_,
		_w11862_
	);
	LUT2 #(
		.INIT('h1)
	) name11401 (
		_w11744_,
		_w11862_,
		_w11863_
	);
	LUT2 #(
		.INIT('h4)
	) name11402 (
		_w11742_,
		_w11863_,
		_w11864_
	);
	LUT2 #(
		.INIT('h1)
	) name11403 (
		_w11741_,
		_w11766_,
		_w11865_
	);
	LUT2 #(
		.INIT('h4)
	) name11404 (
		_w11864_,
		_w11865_,
		_w11866_
	);
	LUT2 #(
		.INIT('h2)
	) name11405 (
		_w11740_,
		_w11866_,
		_w11867_
	);
	LUT2 #(
		.INIT('h1)
	) name11406 (
		_w11734_,
		_w11737_,
		_w11868_
	);
	LUT2 #(
		.INIT('h4)
	) name11407 (
		_w11867_,
		_w11868_,
		_w11869_
	);
	LUT2 #(
		.INIT('h1)
	) name11408 (
		_w11735_,
		_w11869_,
		_w11870_
	);
	LUT2 #(
		.INIT('h1)
	) name11409 (
		_w11860_,
		_w11870_,
		_w11871_
	);
	LUT2 #(
		.INIT('h8)
	) name11410 (
		_w11860_,
		_w11870_,
		_w11872_
	);
	LUT2 #(
		.INIT('h2)
	) name11411 (
		_w11626_,
		_w11871_,
		_w11873_
	);
	LUT2 #(
		.INIT('h4)
	) name11412 (
		_w11872_,
		_w11873_,
		_w11874_
	);
	LUT2 #(
		.INIT('h1)
	) name11413 (
		\P2_reg2_reg[11]/NET0131 ,
		_w2694_,
		_w11875_
	);
	LUT2 #(
		.INIT('h8)
	) name11414 (
		\P2_reg2_reg[11]/NET0131 ,
		_w2694_,
		_w11876_
	);
	LUT2 #(
		.INIT('h1)
	) name11415 (
		_w11875_,
		_w11876_,
		_w11877_
	);
	LUT2 #(
		.INIT('h1)
	) name11416 (
		_w11786_,
		_w11788_,
		_w11878_
	);
	LUT2 #(
		.INIT('h4)
	) name11417 (
		_w11806_,
		_w11878_,
		_w11879_
	);
	LUT2 #(
		.INIT('h1)
	) name11418 (
		_w11787_,
		_w11879_,
		_w11880_
	);
	LUT2 #(
		.INIT('h4)
	) name11419 (
		_w11785_,
		_w11880_,
		_w11881_
	);
	LUT2 #(
		.INIT('h1)
	) name11420 (
		_w11784_,
		_w11809_,
		_w11882_
	);
	LUT2 #(
		.INIT('h4)
	) name11421 (
		_w11881_,
		_w11882_,
		_w11883_
	);
	LUT2 #(
		.INIT('h2)
	) name11422 (
		_w11783_,
		_w11883_,
		_w11884_
	);
	LUT2 #(
		.INIT('h1)
	) name11423 (
		_w11777_,
		_w11780_,
		_w11885_
	);
	LUT2 #(
		.INIT('h4)
	) name11424 (
		_w11884_,
		_w11885_,
		_w11886_
	);
	LUT2 #(
		.INIT('h1)
	) name11425 (
		_w11778_,
		_w11886_,
		_w11887_
	);
	LUT2 #(
		.INIT('h1)
	) name11426 (
		_w11877_,
		_w11887_,
		_w11888_
	);
	LUT2 #(
		.INIT('h8)
	) name11427 (
		_w11877_,
		_w11887_,
		_w11889_
	);
	LUT2 #(
		.INIT('h2)
	) name11428 (
		_w11630_,
		_w11888_,
		_w11890_
	);
	LUT2 #(
		.INIT('h4)
	) name11429 (
		_w11889_,
		_w11890_,
		_w11891_
	);
	LUT2 #(
		.INIT('h1)
	) name11430 (
		_w11857_,
		_w11874_,
		_w11892_
	);
	LUT2 #(
		.INIT('h4)
	) name11431 (
		_w11891_,
		_w11892_,
		_w11893_
	);
	LUT2 #(
		.INIT('h2)
	) name11432 (
		\P1_state_reg[0]/NET0131 ,
		_w11893_,
		_w11894_
	);
	LUT2 #(
		.INIT('h1)
	) name11433 (
		_w8121_,
		_w11894_,
		_w11895_
	);
	LUT2 #(
		.INIT('h4)
	) name11434 (
		\P2_addr_reg[12]/NET0131 ,
		_w11729_,
		_w11896_
	);
	LUT2 #(
		.INIT('h1)
	) name11435 (
		_w2720_,
		_w11729_,
		_w11897_
	);
	LUT2 #(
		.INIT('h1)
	) name11436 (
		_w2058_,
		_w11896_,
		_w11898_
	);
	LUT2 #(
		.INIT('h4)
	) name11437 (
		_w11897_,
		_w11898_,
		_w11899_
	);
	LUT2 #(
		.INIT('h8)
	) name11438 (
		\P2_reg1_reg[12]/NET0131 ,
		_w2720_,
		_w11900_
	);
	LUT2 #(
		.INIT('h1)
	) name11439 (
		\P2_reg1_reg[12]/NET0131 ,
		_w2720_,
		_w11901_
	);
	LUT2 #(
		.INIT('h1)
	) name11440 (
		_w11900_,
		_w11901_,
		_w11902_
	);
	LUT2 #(
		.INIT('h1)
	) name11441 (
		_w11735_,
		_w11772_,
		_w11903_
	);
	LUT2 #(
		.INIT('h1)
	) name11442 (
		_w11734_,
		_w11859_,
		_w11904_
	);
	LUT2 #(
		.INIT('h4)
	) name11443 (
		_w11903_,
		_w11904_,
		_w11905_
	);
	LUT2 #(
		.INIT('h1)
	) name11444 (
		_w11858_,
		_w11905_,
		_w11906_
	);
	LUT2 #(
		.INIT('h1)
	) name11445 (
		_w11902_,
		_w11906_,
		_w11907_
	);
	LUT2 #(
		.INIT('h8)
	) name11446 (
		_w11902_,
		_w11906_,
		_w11908_
	);
	LUT2 #(
		.INIT('h2)
	) name11447 (
		_w11626_,
		_w11907_,
		_w11909_
	);
	LUT2 #(
		.INIT('h4)
	) name11448 (
		_w11908_,
		_w11909_,
		_w11910_
	);
	LUT2 #(
		.INIT('h8)
	) name11449 (
		\P2_reg2_reg[12]/NET0131 ,
		_w2720_,
		_w11911_
	);
	LUT2 #(
		.INIT('h1)
	) name11450 (
		\P2_reg2_reg[12]/NET0131 ,
		_w2720_,
		_w11912_
	);
	LUT2 #(
		.INIT('h1)
	) name11451 (
		_w11911_,
		_w11912_,
		_w11913_
	);
	LUT2 #(
		.INIT('h1)
	) name11452 (
		_w11778_,
		_w11815_,
		_w11914_
	);
	LUT2 #(
		.INIT('h1)
	) name11453 (
		_w11777_,
		_w11876_,
		_w11915_
	);
	LUT2 #(
		.INIT('h4)
	) name11454 (
		_w11914_,
		_w11915_,
		_w11916_
	);
	LUT2 #(
		.INIT('h1)
	) name11455 (
		_w11875_,
		_w11916_,
		_w11917_
	);
	LUT2 #(
		.INIT('h1)
	) name11456 (
		_w11913_,
		_w11917_,
		_w11918_
	);
	LUT2 #(
		.INIT('h8)
	) name11457 (
		_w11913_,
		_w11917_,
		_w11919_
	);
	LUT2 #(
		.INIT('h2)
	) name11458 (
		_w11630_,
		_w11918_,
		_w11920_
	);
	LUT2 #(
		.INIT('h4)
	) name11459 (
		_w11919_,
		_w11920_,
		_w11921_
	);
	LUT2 #(
		.INIT('h1)
	) name11460 (
		_w11899_,
		_w11910_,
		_w11922_
	);
	LUT2 #(
		.INIT('h4)
	) name11461 (
		_w11921_,
		_w11922_,
		_w11923_
	);
	LUT2 #(
		.INIT('h2)
	) name11462 (
		\P1_state_reg[0]/NET0131 ,
		_w11923_,
		_w11924_
	);
	LUT2 #(
		.INIT('h1)
	) name11463 (
		_w6174_,
		_w11924_,
		_w11925_
	);
	LUT2 #(
		.INIT('h4)
	) name11464 (
		\P2_addr_reg[13]/NET0131 ,
		_w11729_,
		_w11926_
	);
	LUT2 #(
		.INIT('h2)
	) name11465 (
		_w2883_,
		_w11729_,
		_w11927_
	);
	LUT2 #(
		.INIT('h1)
	) name11466 (
		_w2058_,
		_w11926_,
		_w11928_
	);
	LUT2 #(
		.INIT('h4)
	) name11467 (
		_w11927_,
		_w11928_,
		_w11929_
	);
	LUT2 #(
		.INIT('h2)
	) name11468 (
		\P2_reg1_reg[13]/NET0131 ,
		_w2883_,
		_w11930_
	);
	LUT2 #(
		.INIT('h4)
	) name11469 (
		\P2_reg1_reg[13]/NET0131 ,
		_w2883_,
		_w11931_
	);
	LUT2 #(
		.INIT('h1)
	) name11470 (
		_w11930_,
		_w11931_,
		_w11932_
	);
	LUT2 #(
		.INIT('h4)
	) name11471 (
		_w11858_,
		_w11870_,
		_w11933_
	);
	LUT2 #(
		.INIT('h1)
	) name11472 (
		_w11859_,
		_w11900_,
		_w11934_
	);
	LUT2 #(
		.INIT('h4)
	) name11473 (
		_w11933_,
		_w11934_,
		_w11935_
	);
	LUT2 #(
		.INIT('h1)
	) name11474 (
		_w11901_,
		_w11935_,
		_w11936_
	);
	LUT2 #(
		.INIT('h1)
	) name11475 (
		_w11932_,
		_w11936_,
		_w11937_
	);
	LUT2 #(
		.INIT('h8)
	) name11476 (
		_w11932_,
		_w11936_,
		_w11938_
	);
	LUT2 #(
		.INIT('h2)
	) name11477 (
		_w11626_,
		_w11937_,
		_w11939_
	);
	LUT2 #(
		.INIT('h4)
	) name11478 (
		_w11938_,
		_w11939_,
		_w11940_
	);
	LUT2 #(
		.INIT('h2)
	) name11479 (
		\P2_reg2_reg[13]/NET0131 ,
		_w2883_,
		_w11941_
	);
	LUT2 #(
		.INIT('h4)
	) name11480 (
		\P2_reg2_reg[13]/NET0131 ,
		_w2883_,
		_w11942_
	);
	LUT2 #(
		.INIT('h1)
	) name11481 (
		_w11941_,
		_w11942_,
		_w11943_
	);
	LUT2 #(
		.INIT('h4)
	) name11482 (
		_w11875_,
		_w11887_,
		_w11944_
	);
	LUT2 #(
		.INIT('h1)
	) name11483 (
		_w11876_,
		_w11911_,
		_w11945_
	);
	LUT2 #(
		.INIT('h4)
	) name11484 (
		_w11944_,
		_w11945_,
		_w11946_
	);
	LUT2 #(
		.INIT('h1)
	) name11485 (
		_w11912_,
		_w11946_,
		_w11947_
	);
	LUT2 #(
		.INIT('h1)
	) name11486 (
		_w11943_,
		_w11947_,
		_w11948_
	);
	LUT2 #(
		.INIT('h8)
	) name11487 (
		_w11943_,
		_w11947_,
		_w11949_
	);
	LUT2 #(
		.INIT('h2)
	) name11488 (
		_w11630_,
		_w11948_,
		_w11950_
	);
	LUT2 #(
		.INIT('h4)
	) name11489 (
		_w11949_,
		_w11950_,
		_w11951_
	);
	LUT2 #(
		.INIT('h1)
	) name11490 (
		_w11929_,
		_w11940_,
		_w11952_
	);
	LUT2 #(
		.INIT('h4)
	) name11491 (
		_w11951_,
		_w11952_,
		_w11953_
	);
	LUT2 #(
		.INIT('h2)
	) name11492 (
		\P1_state_reg[0]/NET0131 ,
		_w11953_,
		_w11954_
	);
	LUT2 #(
		.INIT('h1)
	) name11493 (
		_w7197_,
		_w11954_,
		_w11955_
	);
	LUT2 #(
		.INIT('h4)
	) name11494 (
		\P1_addr_reg[15]/NET0131 ,
		_w11399_,
		_w11956_
	);
	LUT2 #(
		.INIT('h1)
	) name11495 (
		_w1073_,
		_w11399_,
		_w11957_
	);
	LUT2 #(
		.INIT('h1)
	) name11496 (
		_w537_,
		_w11956_,
		_w11958_
	);
	LUT2 #(
		.INIT('h4)
	) name11497 (
		_w11957_,
		_w11958_,
		_w11959_
	);
	LUT2 #(
		.INIT('h1)
	) name11498 (
		\P1_reg2_reg[15]/NET0131 ,
		_w1073_,
		_w11960_
	);
	LUT2 #(
		.INIT('h8)
	) name11499 (
		\P1_reg2_reg[15]/NET0131 ,
		_w1073_,
		_w11961_
	);
	LUT2 #(
		.INIT('h1)
	) name11500 (
		_w11960_,
		_w11961_,
		_w11962_
	);
	LUT2 #(
		.INIT('h1)
	) name11501 (
		_w11569_,
		_w11840_,
		_w11963_
	);
	LUT2 #(
		.INIT('h8)
	) name11502 (
		_w11584_,
		_w11963_,
		_w11964_
	);
	LUT2 #(
		.INIT('h2)
	) name11503 (
		_w11568_,
		_w11840_,
		_w11965_
	);
	LUT2 #(
		.INIT('h1)
	) name11504 (
		_w11839_,
		_w11965_,
		_w11966_
	);
	LUT2 #(
		.INIT('h4)
	) name11505 (
		_w11964_,
		_w11966_,
		_w11967_
	);
	LUT2 #(
		.INIT('h4)
	) name11506 (
		_w11962_,
		_w11967_,
		_w11968_
	);
	LUT2 #(
		.INIT('h2)
	) name11507 (
		_w11962_,
		_w11967_,
		_w11969_
	);
	LUT2 #(
		.INIT('h2)
	) name11508 (
		_w11437_,
		_w11968_,
		_w11970_
	);
	LUT2 #(
		.INIT('h4)
	) name11509 (
		_w11969_,
		_w11970_,
		_w11971_
	);
	LUT2 #(
		.INIT('h1)
	) name11510 (
		\P1_reg1_reg[15]/NET0131 ,
		_w1073_,
		_w11972_
	);
	LUT2 #(
		.INIT('h8)
	) name11511 (
		\P1_reg1_reg[15]/NET0131 ,
		_w1073_,
		_w11973_
	);
	LUT2 #(
		.INIT('h1)
	) name11512 (
		_w11972_,
		_w11973_,
		_w11974_
	);
	LUT2 #(
		.INIT('h4)
	) name11513 (
		_w11594_,
		_w11609_,
		_w11975_
	);
	LUT2 #(
		.INIT('h1)
	) name11514 (
		_w11593_,
		_w11828_,
		_w11976_
	);
	LUT2 #(
		.INIT('h4)
	) name11515 (
		_w11975_,
		_w11976_,
		_w11977_
	);
	LUT2 #(
		.INIT('h1)
	) name11516 (
		_w11829_,
		_w11977_,
		_w11978_
	);
	LUT2 #(
		.INIT('h1)
	) name11517 (
		_w11974_,
		_w11978_,
		_w11979_
	);
	LUT2 #(
		.INIT('h8)
	) name11518 (
		_w11974_,
		_w11978_,
		_w11980_
	);
	LUT2 #(
		.INIT('h2)
	) name11519 (
		_w11404_,
		_w11979_,
		_w11981_
	);
	LUT2 #(
		.INIT('h4)
	) name11520 (
		_w11980_,
		_w11981_,
		_w11982_
	);
	LUT2 #(
		.INIT('h1)
	) name11521 (
		_w11959_,
		_w11971_,
		_w11983_
	);
	LUT2 #(
		.INIT('h4)
	) name11522 (
		_w11982_,
		_w11983_,
		_w11984_
	);
	LUT2 #(
		.INIT('h2)
	) name11523 (
		\P1_state_reg[0]/NET0131 ,
		_w11984_,
		_w11985_
	);
	LUT2 #(
		.INIT('h1)
	) name11524 (
		_w8082_,
		_w11985_,
		_w11986_
	);
	LUT2 #(
		.INIT('h4)
	) name11525 (
		\P2_addr_reg[14]/NET0131 ,
		_w11729_,
		_w11987_
	);
	LUT2 #(
		.INIT('h1)
	) name11526 (
		_w2849_,
		_w11729_,
		_w11988_
	);
	LUT2 #(
		.INIT('h1)
	) name11527 (
		_w2058_,
		_w11987_,
		_w11989_
	);
	LUT2 #(
		.INIT('h4)
	) name11528 (
		_w11988_,
		_w11989_,
		_w11990_
	);
	LUT2 #(
		.INIT('h8)
	) name11529 (
		\P2_reg1_reg[14]/NET0131 ,
		_w2849_,
		_w11991_
	);
	LUT2 #(
		.INIT('h1)
	) name11530 (
		\P2_reg1_reg[14]/NET0131 ,
		_w2849_,
		_w11992_
	);
	LUT2 #(
		.INIT('h1)
	) name11531 (
		_w11991_,
		_w11992_,
		_w11993_
	);
	LUT2 #(
		.INIT('h4)
	) name11532 (
		_w11901_,
		_w11906_,
		_w11994_
	);
	LUT2 #(
		.INIT('h1)
	) name11533 (
		_w11900_,
		_w11930_,
		_w11995_
	);
	LUT2 #(
		.INIT('h4)
	) name11534 (
		_w11994_,
		_w11995_,
		_w11996_
	);
	LUT2 #(
		.INIT('h1)
	) name11535 (
		_w11931_,
		_w11996_,
		_w11997_
	);
	LUT2 #(
		.INIT('h1)
	) name11536 (
		_w11993_,
		_w11997_,
		_w11998_
	);
	LUT2 #(
		.INIT('h8)
	) name11537 (
		_w11993_,
		_w11997_,
		_w11999_
	);
	LUT2 #(
		.INIT('h2)
	) name11538 (
		_w11626_,
		_w11998_,
		_w12000_
	);
	LUT2 #(
		.INIT('h4)
	) name11539 (
		_w11999_,
		_w12000_,
		_w12001_
	);
	LUT2 #(
		.INIT('h8)
	) name11540 (
		\P2_reg2_reg[14]/NET0131 ,
		_w2849_,
		_w12002_
	);
	LUT2 #(
		.INIT('h1)
	) name11541 (
		\P2_reg2_reg[14]/NET0131 ,
		_w2849_,
		_w12003_
	);
	LUT2 #(
		.INIT('h1)
	) name11542 (
		_w12002_,
		_w12003_,
		_w12004_
	);
	LUT2 #(
		.INIT('h4)
	) name11543 (
		_w11912_,
		_w11917_,
		_w12005_
	);
	LUT2 #(
		.INIT('h1)
	) name11544 (
		_w11911_,
		_w11941_,
		_w12006_
	);
	LUT2 #(
		.INIT('h4)
	) name11545 (
		_w12005_,
		_w12006_,
		_w12007_
	);
	LUT2 #(
		.INIT('h1)
	) name11546 (
		_w11942_,
		_w12007_,
		_w12008_
	);
	LUT2 #(
		.INIT('h1)
	) name11547 (
		_w12004_,
		_w12008_,
		_w12009_
	);
	LUT2 #(
		.INIT('h8)
	) name11548 (
		_w12004_,
		_w12008_,
		_w12010_
	);
	LUT2 #(
		.INIT('h2)
	) name11549 (
		_w11630_,
		_w12009_,
		_w12011_
	);
	LUT2 #(
		.INIT('h4)
	) name11550 (
		_w12010_,
		_w12011_,
		_w12012_
	);
	LUT2 #(
		.INIT('h1)
	) name11551 (
		_w11990_,
		_w12001_,
		_w12013_
	);
	LUT2 #(
		.INIT('h4)
	) name11552 (
		_w12012_,
		_w12013_,
		_w12014_
	);
	LUT2 #(
		.INIT('h2)
	) name11553 (
		\P1_state_reg[0]/NET0131 ,
		_w12014_,
		_w12015_
	);
	LUT2 #(
		.INIT('h1)
	) name11554 (
		_w8162_,
		_w12015_,
		_w12016_
	);
	LUT2 #(
		.INIT('h4)
	) name11555 (
		\P2_addr_reg[15]/NET0131 ,
		_w11729_,
		_w12017_
	);
	LUT2 #(
		.INIT('h1)
	) name11556 (
		_w2832_,
		_w11729_,
		_w12018_
	);
	LUT2 #(
		.INIT('h1)
	) name11557 (
		_w2058_,
		_w12017_,
		_w12019_
	);
	LUT2 #(
		.INIT('h4)
	) name11558 (
		_w12018_,
		_w12019_,
		_w12020_
	);
	LUT2 #(
		.INIT('h1)
	) name11559 (
		\P2_reg1_reg[15]/NET0131 ,
		_w2832_,
		_w12021_
	);
	LUT2 #(
		.INIT('h8)
	) name11560 (
		\P2_reg1_reg[15]/NET0131 ,
		_w2832_,
		_w12022_
	);
	LUT2 #(
		.INIT('h1)
	) name11561 (
		_w12021_,
		_w12022_,
		_w12023_
	);
	LUT2 #(
		.INIT('h4)
	) name11562 (
		_w11931_,
		_w11936_,
		_w12024_
	);
	LUT2 #(
		.INIT('h1)
	) name11563 (
		_w11930_,
		_w11991_,
		_w12025_
	);
	LUT2 #(
		.INIT('h4)
	) name11564 (
		_w12024_,
		_w12025_,
		_w12026_
	);
	LUT2 #(
		.INIT('h1)
	) name11565 (
		_w11992_,
		_w12026_,
		_w12027_
	);
	LUT2 #(
		.INIT('h1)
	) name11566 (
		_w12023_,
		_w12027_,
		_w12028_
	);
	LUT2 #(
		.INIT('h8)
	) name11567 (
		_w12023_,
		_w12027_,
		_w12029_
	);
	LUT2 #(
		.INIT('h2)
	) name11568 (
		_w11626_,
		_w12028_,
		_w12030_
	);
	LUT2 #(
		.INIT('h4)
	) name11569 (
		_w12029_,
		_w12030_,
		_w12031_
	);
	LUT2 #(
		.INIT('h1)
	) name11570 (
		\P2_reg2_reg[15]/NET0131 ,
		_w2832_,
		_w12032_
	);
	LUT2 #(
		.INIT('h8)
	) name11571 (
		\P2_reg2_reg[15]/NET0131 ,
		_w2832_,
		_w12033_
	);
	LUT2 #(
		.INIT('h1)
	) name11572 (
		_w12032_,
		_w12033_,
		_w12034_
	);
	LUT2 #(
		.INIT('h4)
	) name11573 (
		_w11942_,
		_w11947_,
		_w12035_
	);
	LUT2 #(
		.INIT('h1)
	) name11574 (
		_w11941_,
		_w12002_,
		_w12036_
	);
	LUT2 #(
		.INIT('h4)
	) name11575 (
		_w12035_,
		_w12036_,
		_w12037_
	);
	LUT2 #(
		.INIT('h1)
	) name11576 (
		_w12003_,
		_w12037_,
		_w12038_
	);
	LUT2 #(
		.INIT('h1)
	) name11577 (
		_w12034_,
		_w12038_,
		_w12039_
	);
	LUT2 #(
		.INIT('h8)
	) name11578 (
		_w12034_,
		_w12038_,
		_w12040_
	);
	LUT2 #(
		.INIT('h2)
	) name11579 (
		_w11630_,
		_w12039_,
		_w12041_
	);
	LUT2 #(
		.INIT('h4)
	) name11580 (
		_w12040_,
		_w12041_,
		_w12042_
	);
	LUT2 #(
		.INIT('h1)
	) name11581 (
		_w12020_,
		_w12031_,
		_w12043_
	);
	LUT2 #(
		.INIT('h4)
	) name11582 (
		_w12042_,
		_w12043_,
		_w12044_
	);
	LUT2 #(
		.INIT('h2)
	) name11583 (
		\P1_state_reg[0]/NET0131 ,
		_w12044_,
		_w12045_
	);
	LUT2 #(
		.INIT('h1)
	) name11584 (
		_w8203_,
		_w12045_,
		_w12046_
	);
	LUT2 #(
		.INIT('h4)
	) name11585 (
		\P2_addr_reg[16]/NET0131 ,
		_w11729_,
		_w12047_
	);
	LUT2 #(
		.INIT('h1)
	) name11586 (
		_w2808_,
		_w11729_,
		_w12048_
	);
	LUT2 #(
		.INIT('h1)
	) name11587 (
		_w2058_,
		_w12047_,
		_w12049_
	);
	LUT2 #(
		.INIT('h4)
	) name11588 (
		_w12048_,
		_w12049_,
		_w12050_
	);
	LUT2 #(
		.INIT('h8)
	) name11589 (
		\P2_reg1_reg[16]/NET0131 ,
		_w2808_,
		_w12051_
	);
	LUT2 #(
		.INIT('h1)
	) name11590 (
		\P2_reg1_reg[16]/NET0131 ,
		_w2808_,
		_w12052_
	);
	LUT2 #(
		.INIT('h1)
	) name11591 (
		_w12051_,
		_w12052_,
		_w12053_
	);
	LUT2 #(
		.INIT('h4)
	) name11592 (
		_w11992_,
		_w11997_,
		_w12054_
	);
	LUT2 #(
		.INIT('h1)
	) name11593 (
		_w11991_,
		_w12022_,
		_w12055_
	);
	LUT2 #(
		.INIT('h4)
	) name11594 (
		_w12054_,
		_w12055_,
		_w12056_
	);
	LUT2 #(
		.INIT('h1)
	) name11595 (
		_w12021_,
		_w12056_,
		_w12057_
	);
	LUT2 #(
		.INIT('h1)
	) name11596 (
		_w12053_,
		_w12057_,
		_w12058_
	);
	LUT2 #(
		.INIT('h8)
	) name11597 (
		_w12053_,
		_w12057_,
		_w12059_
	);
	LUT2 #(
		.INIT('h2)
	) name11598 (
		_w11626_,
		_w12058_,
		_w12060_
	);
	LUT2 #(
		.INIT('h4)
	) name11599 (
		_w12059_,
		_w12060_,
		_w12061_
	);
	LUT2 #(
		.INIT('h8)
	) name11600 (
		\P2_reg2_reg[16]/NET0131 ,
		_w2808_,
		_w12062_
	);
	LUT2 #(
		.INIT('h1)
	) name11601 (
		\P2_reg2_reg[16]/NET0131 ,
		_w2808_,
		_w12063_
	);
	LUT2 #(
		.INIT('h1)
	) name11602 (
		_w12062_,
		_w12063_,
		_w12064_
	);
	LUT2 #(
		.INIT('h4)
	) name11603 (
		_w12003_,
		_w12008_,
		_w12065_
	);
	LUT2 #(
		.INIT('h1)
	) name11604 (
		_w12002_,
		_w12033_,
		_w12066_
	);
	LUT2 #(
		.INIT('h4)
	) name11605 (
		_w12065_,
		_w12066_,
		_w12067_
	);
	LUT2 #(
		.INIT('h1)
	) name11606 (
		_w12032_,
		_w12067_,
		_w12068_
	);
	LUT2 #(
		.INIT('h1)
	) name11607 (
		_w12064_,
		_w12068_,
		_w12069_
	);
	LUT2 #(
		.INIT('h8)
	) name11608 (
		_w12064_,
		_w12068_,
		_w12070_
	);
	LUT2 #(
		.INIT('h2)
	) name11609 (
		_w11630_,
		_w12069_,
		_w12071_
	);
	LUT2 #(
		.INIT('h4)
	) name11610 (
		_w12070_,
		_w12071_,
		_w12072_
	);
	LUT2 #(
		.INIT('h1)
	) name11611 (
		_w12050_,
		_w12061_,
		_w12073_
	);
	LUT2 #(
		.INIT('h4)
	) name11612 (
		_w12072_,
		_w12073_,
		_w12074_
	);
	LUT2 #(
		.INIT('h2)
	) name11613 (
		\P1_state_reg[0]/NET0131 ,
		_w12074_,
		_w12075_
	);
	LUT2 #(
		.INIT('h1)
	) name11614 (
		_w6218_,
		_w12075_,
		_w12076_
	);
	LUT2 #(
		.INIT('h4)
	) name11615 (
		\P2_addr_reg[17]/NET0131 ,
		_w11729_,
		_w12077_
	);
	LUT2 #(
		.INIT('h1)
	) name11616 (
		_w2385_,
		_w11729_,
		_w12078_
	);
	LUT2 #(
		.INIT('h1)
	) name11617 (
		_w2058_,
		_w12077_,
		_w12079_
	);
	LUT2 #(
		.INIT('h4)
	) name11618 (
		_w12078_,
		_w12079_,
		_w12080_
	);
	LUT2 #(
		.INIT('h1)
	) name11619 (
		\P2_reg1_reg[17]/NET0131 ,
		_w2385_,
		_w12081_
	);
	LUT2 #(
		.INIT('h8)
	) name11620 (
		\P2_reg1_reg[17]/NET0131 ,
		_w2385_,
		_w12082_
	);
	LUT2 #(
		.INIT('h1)
	) name11621 (
		_w12081_,
		_w12082_,
		_w12083_
	);
	LUT2 #(
		.INIT('h4)
	) name11622 (
		_w12021_,
		_w12027_,
		_w12084_
	);
	LUT2 #(
		.INIT('h1)
	) name11623 (
		_w12022_,
		_w12051_,
		_w12085_
	);
	LUT2 #(
		.INIT('h4)
	) name11624 (
		_w12084_,
		_w12085_,
		_w12086_
	);
	LUT2 #(
		.INIT('h1)
	) name11625 (
		_w12052_,
		_w12086_,
		_w12087_
	);
	LUT2 #(
		.INIT('h1)
	) name11626 (
		_w12083_,
		_w12087_,
		_w12088_
	);
	LUT2 #(
		.INIT('h8)
	) name11627 (
		_w12083_,
		_w12087_,
		_w12089_
	);
	LUT2 #(
		.INIT('h2)
	) name11628 (
		_w11626_,
		_w12088_,
		_w12090_
	);
	LUT2 #(
		.INIT('h4)
	) name11629 (
		_w12089_,
		_w12090_,
		_w12091_
	);
	LUT2 #(
		.INIT('h1)
	) name11630 (
		\P2_reg2_reg[17]/NET0131 ,
		_w2385_,
		_w12092_
	);
	LUT2 #(
		.INIT('h8)
	) name11631 (
		\P2_reg2_reg[17]/NET0131 ,
		_w2385_,
		_w12093_
	);
	LUT2 #(
		.INIT('h1)
	) name11632 (
		_w12092_,
		_w12093_,
		_w12094_
	);
	LUT2 #(
		.INIT('h4)
	) name11633 (
		_w12032_,
		_w12038_,
		_w12095_
	);
	LUT2 #(
		.INIT('h1)
	) name11634 (
		_w12033_,
		_w12062_,
		_w12096_
	);
	LUT2 #(
		.INIT('h4)
	) name11635 (
		_w12095_,
		_w12096_,
		_w12097_
	);
	LUT2 #(
		.INIT('h1)
	) name11636 (
		_w12063_,
		_w12097_,
		_w12098_
	);
	LUT2 #(
		.INIT('h1)
	) name11637 (
		_w12094_,
		_w12098_,
		_w12099_
	);
	LUT2 #(
		.INIT('h8)
	) name11638 (
		_w12094_,
		_w12098_,
		_w12100_
	);
	LUT2 #(
		.INIT('h2)
	) name11639 (
		_w11630_,
		_w12099_,
		_w12101_
	);
	LUT2 #(
		.INIT('h4)
	) name11640 (
		_w12100_,
		_w12101_,
		_w12102_
	);
	LUT2 #(
		.INIT('h1)
	) name11641 (
		_w12080_,
		_w12091_,
		_w12103_
	);
	LUT2 #(
		.INIT('h4)
	) name11642 (
		_w12102_,
		_w12103_,
		_w12104_
	);
	LUT2 #(
		.INIT('h2)
	) name11643 (
		\P1_state_reg[0]/NET0131 ,
		_w12104_,
		_w12105_
	);
	LUT2 #(
		.INIT('h1)
	) name11644 (
		_w5551_,
		_w12105_,
		_w12106_
	);
	LUT2 #(
		.INIT('h4)
	) name11645 (
		\P1_addr_reg[16]/NET0131 ,
		_w11399_,
		_w12107_
	);
	LUT2 #(
		.INIT('h1)
	) name11646 (
		_w1456_,
		_w11399_,
		_w12108_
	);
	LUT2 #(
		.INIT('h1)
	) name11647 (
		_w537_,
		_w12107_,
		_w12109_
	);
	LUT2 #(
		.INIT('h4)
	) name11648 (
		_w12108_,
		_w12109_,
		_w12110_
	);
	LUT2 #(
		.INIT('h8)
	) name11649 (
		\P1_reg1_reg[16]/NET0131 ,
		_w1456_,
		_w12111_
	);
	LUT2 #(
		.INIT('h1)
	) name11650 (
		\P1_reg1_reg[16]/NET0131 ,
		_w1456_,
		_w12112_
	);
	LUT2 #(
		.INIT('h1)
	) name11651 (
		_w12111_,
		_w12112_,
		_w12113_
	);
	LUT2 #(
		.INIT('h4)
	) name11652 (
		_w11829_,
		_w11834_,
		_w12114_
	);
	LUT2 #(
		.INIT('h1)
	) name11653 (
		_w11828_,
		_w11973_,
		_w12115_
	);
	LUT2 #(
		.INIT('h4)
	) name11654 (
		_w12114_,
		_w12115_,
		_w12116_
	);
	LUT2 #(
		.INIT('h1)
	) name11655 (
		_w11972_,
		_w12116_,
		_w12117_
	);
	LUT2 #(
		.INIT('h1)
	) name11656 (
		_w12113_,
		_w12117_,
		_w12118_
	);
	LUT2 #(
		.INIT('h8)
	) name11657 (
		_w12113_,
		_w12117_,
		_w12119_
	);
	LUT2 #(
		.INIT('h2)
	) name11658 (
		_w11404_,
		_w12118_,
		_w12120_
	);
	LUT2 #(
		.INIT('h4)
	) name11659 (
		_w12119_,
		_w12120_,
		_w12121_
	);
	LUT2 #(
		.INIT('h8)
	) name11660 (
		\P1_reg2_reg[16]/NET0131 ,
		_w1456_,
		_w12122_
	);
	LUT2 #(
		.INIT('h1)
	) name11661 (
		\P1_reg2_reg[16]/NET0131 ,
		_w1456_,
		_w12123_
	);
	LUT2 #(
		.INIT('h1)
	) name11662 (
		_w12122_,
		_w12123_,
		_w12124_
	);
	LUT2 #(
		.INIT('h4)
	) name11663 (
		_w11840_,
		_w11845_,
		_w12125_
	);
	LUT2 #(
		.INIT('h1)
	) name11664 (
		_w11839_,
		_w11961_,
		_w12126_
	);
	LUT2 #(
		.INIT('h4)
	) name11665 (
		_w12125_,
		_w12126_,
		_w12127_
	);
	LUT2 #(
		.INIT('h1)
	) name11666 (
		_w11960_,
		_w12127_,
		_w12128_
	);
	LUT2 #(
		.INIT('h1)
	) name11667 (
		_w12124_,
		_w12128_,
		_w12129_
	);
	LUT2 #(
		.INIT('h8)
	) name11668 (
		_w12124_,
		_w12128_,
		_w12130_
	);
	LUT2 #(
		.INIT('h2)
	) name11669 (
		_w11437_,
		_w12129_,
		_w12131_
	);
	LUT2 #(
		.INIT('h4)
	) name11670 (
		_w12130_,
		_w12131_,
		_w12132_
	);
	LUT2 #(
		.INIT('h1)
	) name11671 (
		_w12110_,
		_w12121_,
		_w12133_
	);
	LUT2 #(
		.INIT('h4)
	) name11672 (
		_w12132_,
		_w12133_,
		_w12134_
	);
	LUT2 #(
		.INIT('h2)
	) name11673 (
		\P1_state_reg[0]/NET0131 ,
		_w12134_,
		_w12135_
	);
	LUT2 #(
		.INIT('h1)
	) name11674 (
		_w6132_,
		_w12135_,
		_w12136_
	);
	LUT2 #(
		.INIT('h4)
	) name11675 (
		\P1_state_reg[0]/NET0131 ,
		\P2_reg3_reg[1]/NET0131 ,
		_w12137_
	);
	LUT2 #(
		.INIT('h8)
	) name11676 (
		_w2578_,
		_w11619_,
		_w12138_
	);
	LUT2 #(
		.INIT('h1)
	) name11677 (
		\P2_addr_reg[1]/NET0131 ,
		_w2024_,
		_w12139_
	);
	LUT2 #(
		.INIT('h2)
	) name11678 (
		_w2024_,
		_w2578_,
		_w12140_
	);
	LUT2 #(
		.INIT('h2)
	) name11679 (
		_w2059_,
		_w12139_,
		_w12141_
	);
	LUT2 #(
		.INIT('h4)
	) name11680 (
		_w12140_,
		_w12141_,
		_w12142_
	);
	LUT2 #(
		.INIT('h1)
	) name11681 (
		_w11796_,
		_w11797_,
		_w12143_
	);
	LUT2 #(
		.INIT('h1)
	) name11682 (
		_w11632_,
		_w12143_,
		_w12144_
	);
	LUT2 #(
		.INIT('h8)
	) name11683 (
		_w11632_,
		_w12143_,
		_w12145_
	);
	LUT2 #(
		.INIT('h1)
	) name11684 (
		_w12144_,
		_w12145_,
		_w12146_
	);
	LUT2 #(
		.INIT('h8)
	) name11685 (
		_w11630_,
		_w12146_,
		_w12147_
	);
	LUT2 #(
		.INIT('h1)
	) name11686 (
		_w11751_,
		_w11752_,
		_w12148_
	);
	LUT2 #(
		.INIT('h1)
	) name11687 (
		_w11627_,
		_w12148_,
		_w12149_
	);
	LUT2 #(
		.INIT('h8)
	) name11688 (
		_w11627_,
		_w12148_,
		_w12150_
	);
	LUT2 #(
		.INIT('h1)
	) name11689 (
		_w12149_,
		_w12150_,
		_w12151_
	);
	LUT2 #(
		.INIT('h8)
	) name11690 (
		_w11626_,
		_w12151_,
		_w12152_
	);
	LUT2 #(
		.INIT('h1)
	) name11691 (
		_w12138_,
		_w12147_,
		_w12153_
	);
	LUT2 #(
		.INIT('h4)
	) name11692 (
		_w12152_,
		_w12153_,
		_w12154_
	);
	LUT2 #(
		.INIT('h4)
	) name11693 (
		_w12142_,
		_w12154_,
		_w12155_
	);
	LUT2 #(
		.INIT('h2)
	) name11694 (
		\P1_state_reg[0]/NET0131 ,
		_w12155_,
		_w12156_
	);
	LUT2 #(
		.INIT('h1)
	) name11695 (
		_w12137_,
		_w12156_,
		_w12157_
	);
	LUT2 #(
		.INIT('h4)
	) name11696 (
		\P1_addr_reg[17]/NET0131 ,
		_w11399_,
		_w12158_
	);
	LUT2 #(
		.INIT('h2)
	) name11697 (
		_w1433_,
		_w11399_,
		_w12159_
	);
	LUT2 #(
		.INIT('h1)
	) name11698 (
		_w537_,
		_w12158_,
		_w12160_
	);
	LUT2 #(
		.INIT('h4)
	) name11699 (
		_w12159_,
		_w12160_,
		_w12161_
	);
	LUT2 #(
		.INIT('h4)
	) name11700 (
		\P1_reg2_reg[17]/NET0131 ,
		_w1433_,
		_w12162_
	);
	LUT2 #(
		.INIT('h2)
	) name11701 (
		\P1_reg2_reg[17]/NET0131 ,
		_w1433_,
		_w12163_
	);
	LUT2 #(
		.INIT('h1)
	) name11702 (
		_w12162_,
		_w12163_,
		_w12164_
	);
	LUT2 #(
		.INIT('h1)
	) name11703 (
		_w11960_,
		_w11967_,
		_w12165_
	);
	LUT2 #(
		.INIT('h1)
	) name11704 (
		_w11961_,
		_w12122_,
		_w12166_
	);
	LUT2 #(
		.INIT('h4)
	) name11705 (
		_w12165_,
		_w12166_,
		_w12167_
	);
	LUT2 #(
		.INIT('h1)
	) name11706 (
		_w12123_,
		_w12167_,
		_w12168_
	);
	LUT2 #(
		.INIT('h1)
	) name11707 (
		_w12164_,
		_w12168_,
		_w12169_
	);
	LUT2 #(
		.INIT('h8)
	) name11708 (
		_w12164_,
		_w12168_,
		_w12170_
	);
	LUT2 #(
		.INIT('h2)
	) name11709 (
		_w11437_,
		_w12169_,
		_w12171_
	);
	LUT2 #(
		.INIT('h4)
	) name11710 (
		_w12170_,
		_w12171_,
		_w12172_
	);
	LUT2 #(
		.INIT('h4)
	) name11711 (
		\P1_reg1_reg[17]/NET0131 ,
		_w1433_,
		_w12173_
	);
	LUT2 #(
		.INIT('h2)
	) name11712 (
		\P1_reg1_reg[17]/NET0131 ,
		_w1433_,
		_w12174_
	);
	LUT2 #(
		.INIT('h1)
	) name11713 (
		_w12173_,
		_w12174_,
		_w12175_
	);
	LUT2 #(
		.INIT('h4)
	) name11714 (
		_w11972_,
		_w11978_,
		_w12176_
	);
	LUT2 #(
		.INIT('h1)
	) name11715 (
		_w11973_,
		_w12111_,
		_w12177_
	);
	LUT2 #(
		.INIT('h4)
	) name11716 (
		_w12176_,
		_w12177_,
		_w12178_
	);
	LUT2 #(
		.INIT('h1)
	) name11717 (
		_w12112_,
		_w12178_,
		_w12179_
	);
	LUT2 #(
		.INIT('h1)
	) name11718 (
		_w12175_,
		_w12179_,
		_w12180_
	);
	LUT2 #(
		.INIT('h8)
	) name11719 (
		_w12175_,
		_w12179_,
		_w12181_
	);
	LUT2 #(
		.INIT('h2)
	) name11720 (
		_w11404_,
		_w12180_,
		_w12182_
	);
	LUT2 #(
		.INIT('h4)
	) name11721 (
		_w12181_,
		_w12182_,
		_w12183_
	);
	LUT2 #(
		.INIT('h1)
	) name11722 (
		_w12161_,
		_w12172_,
		_w12184_
	);
	LUT2 #(
		.INIT('h4)
	) name11723 (
		_w12183_,
		_w12184_,
		_w12185_
	);
	LUT2 #(
		.INIT('h2)
	) name11724 (
		\P1_state_reg[0]/NET0131 ,
		_w12185_,
		_w12186_
	);
	LUT2 #(
		.INIT('h1)
	) name11725 (
		_w5426_,
		_w12186_,
		_w12187_
	);
	LUT2 #(
		.INIT('h4)
	) name11726 (
		\P1_state_reg[0]/NET0131 ,
		\P2_reg3_reg[2]/NET0131 ,
		_w12188_
	);
	LUT2 #(
		.INIT('h8)
	) name11727 (
		_w2564_,
		_w11619_,
		_w12189_
	);
	LUT2 #(
		.INIT('h1)
	) name11728 (
		\P2_addr_reg[2]/NET0131 ,
		_w2024_,
		_w12190_
	);
	LUT2 #(
		.INIT('h2)
	) name11729 (
		_w2024_,
		_w2564_,
		_w12191_
	);
	LUT2 #(
		.INIT('h2)
	) name11730 (
		_w2059_,
		_w12190_,
		_w12192_
	);
	LUT2 #(
		.INIT('h4)
	) name11731 (
		_w12191_,
		_w12192_,
		_w12193_
	);
	LUT2 #(
		.INIT('h1)
	) name11732 (
		_w11794_,
		_w11795_,
		_w12194_
	);
	LUT2 #(
		.INIT('h1)
	) name11733 (
		_w11799_,
		_w12194_,
		_w12195_
	);
	LUT2 #(
		.INIT('h8)
	) name11734 (
		_w11799_,
		_w12194_,
		_w12196_
	);
	LUT2 #(
		.INIT('h1)
	) name11735 (
		_w12195_,
		_w12196_,
		_w12197_
	);
	LUT2 #(
		.INIT('h8)
	) name11736 (
		_w11630_,
		_w12197_,
		_w12198_
	);
	LUT2 #(
		.INIT('h1)
	) name11737 (
		_w11749_,
		_w11750_,
		_w12199_
	);
	LUT2 #(
		.INIT('h1)
	) name11738 (
		_w11754_,
		_w12199_,
		_w12200_
	);
	LUT2 #(
		.INIT('h8)
	) name11739 (
		_w11754_,
		_w12199_,
		_w12201_
	);
	LUT2 #(
		.INIT('h1)
	) name11740 (
		_w12200_,
		_w12201_,
		_w12202_
	);
	LUT2 #(
		.INIT('h8)
	) name11741 (
		_w11626_,
		_w12202_,
		_w12203_
	);
	LUT2 #(
		.INIT('h1)
	) name11742 (
		_w12189_,
		_w12198_,
		_w12204_
	);
	LUT2 #(
		.INIT('h4)
	) name11743 (
		_w12203_,
		_w12204_,
		_w12205_
	);
	LUT2 #(
		.INIT('h4)
	) name11744 (
		_w12193_,
		_w12205_,
		_w12206_
	);
	LUT2 #(
		.INIT('h2)
	) name11745 (
		\P1_state_reg[0]/NET0131 ,
		_w12206_,
		_w12207_
	);
	LUT2 #(
		.INIT('h1)
	) name11746 (
		_w12188_,
		_w12207_,
		_w12208_
	);
	LUT2 #(
		.INIT('h8)
	) name11747 (
		_w2629_,
		_w11619_,
		_w12209_
	);
	LUT2 #(
		.INIT('h1)
	) name11748 (
		\P2_addr_reg[3]/NET0131 ,
		_w2024_,
		_w12210_
	);
	LUT2 #(
		.INIT('h2)
	) name11749 (
		_w2024_,
		_w2629_,
		_w12211_
	);
	LUT2 #(
		.INIT('h2)
	) name11750 (
		_w2059_,
		_w12210_,
		_w12212_
	);
	LUT2 #(
		.INIT('h4)
	) name11751 (
		_w12211_,
		_w12212_,
		_w12213_
	);
	LUT2 #(
		.INIT('h1)
	) name11752 (
		_w11748_,
		_w11759_,
		_w12214_
	);
	LUT2 #(
		.INIT('h1)
	) name11753 (
		_w11756_,
		_w12214_,
		_w12215_
	);
	LUT2 #(
		.INIT('h8)
	) name11754 (
		_w11756_,
		_w12214_,
		_w12216_
	);
	LUT2 #(
		.INIT('h1)
	) name11755 (
		_w12215_,
		_w12216_,
		_w12217_
	);
	LUT2 #(
		.INIT('h8)
	) name11756 (
		_w11626_,
		_w12217_,
		_w12218_
	);
	LUT2 #(
		.INIT('h1)
	) name11757 (
		_w11792_,
		_w11793_,
		_w12219_
	);
	LUT2 #(
		.INIT('h1)
	) name11758 (
		_w11801_,
		_w12219_,
		_w12220_
	);
	LUT2 #(
		.INIT('h8)
	) name11759 (
		_w11801_,
		_w12219_,
		_w12221_
	);
	LUT2 #(
		.INIT('h1)
	) name11760 (
		_w12220_,
		_w12221_,
		_w12222_
	);
	LUT2 #(
		.INIT('h8)
	) name11761 (
		_w11630_,
		_w12222_,
		_w12223_
	);
	LUT2 #(
		.INIT('h1)
	) name11762 (
		_w12209_,
		_w12218_,
		_w12224_
	);
	LUT2 #(
		.INIT('h4)
	) name11763 (
		_w12223_,
		_w12224_,
		_w12225_
	);
	LUT2 #(
		.INIT('h4)
	) name11764 (
		_w12213_,
		_w12225_,
		_w12226_
	);
	LUT2 #(
		.INIT('h2)
	) name11765 (
		\P1_state_reg[0]/NET0131 ,
		_w12226_,
		_w12227_
	);
	LUT2 #(
		.INIT('h1)
	) name11766 (
		_w9575_,
		_w12227_,
		_w12228_
	);
	LUT2 #(
		.INIT('h8)
	) name11767 (
		_w2646_,
		_w11619_,
		_w12229_
	);
	LUT2 #(
		.INIT('h1)
	) name11768 (
		\P2_addr_reg[4]/NET0131 ,
		_w2024_,
		_w12230_
	);
	LUT2 #(
		.INIT('h2)
	) name11769 (
		_w2024_,
		_w2646_,
		_w12231_
	);
	LUT2 #(
		.INIT('h2)
	) name11770 (
		_w2059_,
		_w12230_,
		_w12232_
	);
	LUT2 #(
		.INIT('h4)
	) name11771 (
		_w12231_,
		_w12232_,
		_w12233_
	);
	LUT2 #(
		.INIT('h1)
	) name11772 (
		_w11790_,
		_w11791_,
		_w12234_
	);
	LUT2 #(
		.INIT('h1)
	) name11773 (
		_w11803_,
		_w12234_,
		_w12235_
	);
	LUT2 #(
		.INIT('h8)
	) name11774 (
		_w11803_,
		_w12234_,
		_w12236_
	);
	LUT2 #(
		.INIT('h1)
	) name11775 (
		_w12235_,
		_w12236_,
		_w12237_
	);
	LUT2 #(
		.INIT('h8)
	) name11776 (
		_w11630_,
		_w12237_,
		_w12238_
	);
	LUT2 #(
		.INIT('h1)
	) name11777 (
		_w11757_,
		_w11759_,
		_w12239_
	);
	LUT2 #(
		.INIT('h1)
	) name11778 (
		_w11747_,
		_w11758_,
		_w12240_
	);
	LUT2 #(
		.INIT('h2)
	) name11779 (
		_w12239_,
		_w12240_,
		_w12241_
	);
	LUT2 #(
		.INIT('h4)
	) name11780 (
		_w12239_,
		_w12240_,
		_w12242_
	);
	LUT2 #(
		.INIT('h1)
	) name11781 (
		_w12241_,
		_w12242_,
		_w12243_
	);
	LUT2 #(
		.INIT('h8)
	) name11782 (
		_w11626_,
		_w12243_,
		_w12244_
	);
	LUT2 #(
		.INIT('h1)
	) name11783 (
		_w12229_,
		_w12238_,
		_w12245_
	);
	LUT2 #(
		.INIT('h4)
	) name11784 (
		_w12244_,
		_w12245_,
		_w12246_
	);
	LUT2 #(
		.INIT('h4)
	) name11785 (
		_w12233_,
		_w12246_,
		_w12247_
	);
	LUT2 #(
		.INIT('h2)
	) name11786 (
		\P1_state_reg[0]/NET0131 ,
		_w12247_,
		_w12248_
	);
	LUT2 #(
		.INIT('h1)
	) name11787 (
		_w8935_,
		_w12248_,
		_w12249_
	);
	LUT2 #(
		.INIT('h4)
	) name11788 (
		_w2542_,
		_w11619_,
		_w12250_
	);
	LUT2 #(
		.INIT('h1)
	) name11789 (
		\P2_addr_reg[5]/NET0131 ,
		_w2024_,
		_w12251_
	);
	LUT2 #(
		.INIT('h8)
	) name11790 (
		_w2024_,
		_w2542_,
		_w12252_
	);
	LUT2 #(
		.INIT('h2)
	) name11791 (
		_w2059_,
		_w12251_,
		_w12253_
	);
	LUT2 #(
		.INIT('h4)
	) name11792 (
		_w12252_,
		_w12253_,
		_w12254_
	);
	LUT2 #(
		.INIT('h1)
	) name11793 (
		_w11745_,
		_w11746_,
		_w12255_
	);
	LUT2 #(
		.INIT('h1)
	) name11794 (
		_w11762_,
		_w12255_,
		_w12256_
	);
	LUT2 #(
		.INIT('h4)
	) name11795 (
		_w11745_,
		_w11763_,
		_w12257_
	);
	LUT2 #(
		.INIT('h2)
	) name11796 (
		_w11626_,
		_w12256_,
		_w12258_
	);
	LUT2 #(
		.INIT('h4)
	) name11797 (
		_w12257_,
		_w12258_,
		_w12259_
	);
	LUT2 #(
		.INIT('h1)
	) name11798 (
		_w11788_,
		_w11789_,
		_w12260_
	);
	LUT2 #(
		.INIT('h1)
	) name11799 (
		_w11805_,
		_w12260_,
		_w12261_
	);
	LUT2 #(
		.INIT('h8)
	) name11800 (
		_w11805_,
		_w12260_,
		_w12262_
	);
	LUT2 #(
		.INIT('h2)
	) name11801 (
		_w11630_,
		_w12261_,
		_w12263_
	);
	LUT2 #(
		.INIT('h4)
	) name11802 (
		_w12262_,
		_w12263_,
		_w12264_
	);
	LUT2 #(
		.INIT('h1)
	) name11803 (
		_w12250_,
		_w12259_,
		_w12265_
	);
	LUT2 #(
		.INIT('h4)
	) name11804 (
		_w12264_,
		_w12265_,
		_w12266_
	);
	LUT2 #(
		.INIT('h4)
	) name11805 (
		_w12254_,
		_w12266_,
		_w12267_
	);
	LUT2 #(
		.INIT('h2)
	) name11806 (
		\P1_state_reg[0]/NET0131 ,
		_w12267_,
		_w12268_
	);
	LUT2 #(
		.INIT('h1)
	) name11807 (
		_w8977_,
		_w12268_,
		_w12269_
	);
	LUT2 #(
		.INIT('h4)
	) name11808 (
		\P2_addr_reg[6]/NET0131 ,
		_w11729_,
		_w12270_
	);
	LUT2 #(
		.INIT('h1)
	) name11809 (
		_w2519_,
		_w11729_,
		_w12271_
	);
	LUT2 #(
		.INIT('h1)
	) name11810 (
		_w2058_,
		_w12270_,
		_w12272_
	);
	LUT2 #(
		.INIT('h4)
	) name11811 (
		_w12271_,
		_w12272_,
		_w12273_
	);
	LUT2 #(
		.INIT('h1)
	) name11812 (
		_w11743_,
		_w11744_,
		_w12274_
	);
	LUT2 #(
		.INIT('h2)
	) name11813 (
		_w11764_,
		_w12274_,
		_w12275_
	);
	LUT2 #(
		.INIT('h4)
	) name11814 (
		_w11764_,
		_w12274_,
		_w12276_
	);
	LUT2 #(
		.INIT('h2)
	) name11815 (
		_w11626_,
		_w12275_,
		_w12277_
	);
	LUT2 #(
		.INIT('h4)
	) name11816 (
		_w12276_,
		_w12277_,
		_w12278_
	);
	LUT2 #(
		.INIT('h1)
	) name11817 (
		_w11786_,
		_w11787_,
		_w12279_
	);
	LUT2 #(
		.INIT('h2)
	) name11818 (
		_w11807_,
		_w12279_,
		_w12280_
	);
	LUT2 #(
		.INIT('h4)
	) name11819 (
		_w11807_,
		_w12279_,
		_w12281_
	);
	LUT2 #(
		.INIT('h2)
	) name11820 (
		_w11630_,
		_w12280_,
		_w12282_
	);
	LUT2 #(
		.INIT('h4)
	) name11821 (
		_w12281_,
		_w12282_,
		_w12283_
	);
	LUT2 #(
		.INIT('h1)
	) name11822 (
		_w12273_,
		_w12278_,
		_w12284_
	);
	LUT2 #(
		.INIT('h4)
	) name11823 (
		_w12283_,
		_w12284_,
		_w12285_
	);
	LUT2 #(
		.INIT('h2)
	) name11824 (
		\P1_state_reg[0]/NET0131 ,
		_w12285_,
		_w12286_
	);
	LUT2 #(
		.INIT('h1)
	) name11825 (
		_w9615_,
		_w12286_,
		_w12287_
	);
	LUT2 #(
		.INIT('h1)
	) name11826 (
		_w11742_,
		_w11766_,
		_w12288_
	);
	LUT2 #(
		.INIT('h1)
	) name11827 (
		_w11863_,
		_w12288_,
		_w12289_
	);
	LUT2 #(
		.INIT('h4)
	) name11828 (
		_w11766_,
		_w11864_,
		_w12290_
	);
	LUT2 #(
		.INIT('h2)
	) name11829 (
		_w11626_,
		_w12289_,
		_w12291_
	);
	LUT2 #(
		.INIT('h4)
	) name11830 (
		_w12290_,
		_w12291_,
		_w12292_
	);
	LUT2 #(
		.INIT('h4)
	) name11831 (
		\P2_addr_reg[7]/NET0131 ,
		_w11729_,
		_w12293_
	);
	LUT2 #(
		.INIT('h1)
	) name11832 (
		_w2485_,
		_w11729_,
		_w12294_
	);
	LUT2 #(
		.INIT('h1)
	) name11833 (
		_w2058_,
		_w12293_,
		_w12295_
	);
	LUT2 #(
		.INIT('h4)
	) name11834 (
		_w12294_,
		_w12295_,
		_w12296_
	);
	LUT2 #(
		.INIT('h1)
	) name11835 (
		_w11785_,
		_w11809_,
		_w12297_
	);
	LUT2 #(
		.INIT('h1)
	) name11836 (
		_w11880_,
		_w12297_,
		_w12298_
	);
	LUT2 #(
		.INIT('h4)
	) name11837 (
		_w11809_,
		_w11881_,
		_w12299_
	);
	LUT2 #(
		.INIT('h2)
	) name11838 (
		_w11630_,
		_w12298_,
		_w12300_
	);
	LUT2 #(
		.INIT('h4)
	) name11839 (
		_w12299_,
		_w12300_,
		_w12301_
	);
	LUT2 #(
		.INIT('h1)
	) name11840 (
		_w12292_,
		_w12296_,
		_w12302_
	);
	LUT2 #(
		.INIT('h4)
	) name11841 (
		_w12301_,
		_w12302_,
		_w12303_
	);
	LUT2 #(
		.INIT('h2)
	) name11842 (
		\P1_state_reg[0]/NET0131 ,
		_w12303_,
		_w12304_
	);
	LUT2 #(
		.INIT('h1)
	) name11843 (
		_w9656_,
		_w12304_,
		_w12305_
	);
	LUT2 #(
		.INIT('h1)
	) name11844 (
		_w11739_,
		_w11741_,
		_w12306_
	);
	LUT2 #(
		.INIT('h1)
	) name11845 (
		_w11769_,
		_w12306_,
		_w12307_
	);
	LUT2 #(
		.INIT('h8)
	) name11846 (
		_w11769_,
		_w12306_,
		_w12308_
	);
	LUT2 #(
		.INIT('h2)
	) name11847 (
		_w11626_,
		_w12307_,
		_w12309_
	);
	LUT2 #(
		.INIT('h4)
	) name11848 (
		_w12308_,
		_w12309_,
		_w12310_
	);
	LUT2 #(
		.INIT('h4)
	) name11849 (
		\P2_addr_reg[8]/NET0131 ,
		_w11729_,
		_w12311_
	);
	LUT2 #(
		.INIT('h1)
	) name11850 (
		_w2460_,
		_w11729_,
		_w12312_
	);
	LUT2 #(
		.INIT('h1)
	) name11851 (
		_w2058_,
		_w12311_,
		_w12313_
	);
	LUT2 #(
		.INIT('h4)
	) name11852 (
		_w12312_,
		_w12313_,
		_w12314_
	);
	LUT2 #(
		.INIT('h1)
	) name11853 (
		_w11782_,
		_w11784_,
		_w12315_
	);
	LUT2 #(
		.INIT('h1)
	) name11854 (
		_w11812_,
		_w12315_,
		_w12316_
	);
	LUT2 #(
		.INIT('h8)
	) name11855 (
		_w11812_,
		_w12315_,
		_w12317_
	);
	LUT2 #(
		.INIT('h2)
	) name11856 (
		_w11630_,
		_w12316_,
		_w12318_
	);
	LUT2 #(
		.INIT('h4)
	) name11857 (
		_w12317_,
		_w12318_,
		_w12319_
	);
	LUT2 #(
		.INIT('h1)
	) name11858 (
		_w12310_,
		_w12314_,
		_w12320_
	);
	LUT2 #(
		.INIT('h4)
	) name11859 (
		_w12319_,
		_w12320_,
		_w12321_
	);
	LUT2 #(
		.INIT('h2)
	) name11860 (
		\P1_state_reg[0]/NET0131 ,
		_w12321_,
		_w12322_
	);
	LUT2 #(
		.INIT('h1)
	) name11861 (
		_w8243_,
		_w12322_,
		_w12323_
	);
	LUT2 #(
		.INIT('h1)
	) name11862 (
		_w11737_,
		_w11738_,
		_w12324_
	);
	LUT2 #(
		.INIT('h1)
	) name11863 (
		_w11739_,
		_w11866_,
		_w12325_
	);
	LUT2 #(
		.INIT('h1)
	) name11864 (
		_w12324_,
		_w12325_,
		_w12326_
	);
	LUT2 #(
		.INIT('h4)
	) name11865 (
		_w11737_,
		_w11867_,
		_w12327_
	);
	LUT2 #(
		.INIT('h2)
	) name11866 (
		_w11626_,
		_w12326_,
		_w12328_
	);
	LUT2 #(
		.INIT('h4)
	) name11867 (
		_w12327_,
		_w12328_,
		_w12329_
	);
	LUT2 #(
		.INIT('h4)
	) name11868 (
		\P2_addr_reg[9]/NET0131 ,
		_w11729_,
		_w12330_
	);
	LUT2 #(
		.INIT('h2)
	) name11869 (
		_w2769_,
		_w11729_,
		_w12331_
	);
	LUT2 #(
		.INIT('h1)
	) name11870 (
		_w2058_,
		_w12330_,
		_w12332_
	);
	LUT2 #(
		.INIT('h4)
	) name11871 (
		_w12331_,
		_w12332_,
		_w12333_
	);
	LUT2 #(
		.INIT('h1)
	) name11872 (
		_w11780_,
		_w11781_,
		_w12334_
	);
	LUT2 #(
		.INIT('h1)
	) name11873 (
		_w11782_,
		_w11883_,
		_w12335_
	);
	LUT2 #(
		.INIT('h1)
	) name11874 (
		_w12334_,
		_w12335_,
		_w12336_
	);
	LUT2 #(
		.INIT('h4)
	) name11875 (
		_w11780_,
		_w11884_,
		_w12337_
	);
	LUT2 #(
		.INIT('h2)
	) name11876 (
		_w11630_,
		_w12336_,
		_w12338_
	);
	LUT2 #(
		.INIT('h4)
	) name11877 (
		_w12337_,
		_w12338_,
		_w12339_
	);
	LUT2 #(
		.INIT('h1)
	) name11878 (
		_w12329_,
		_w12333_,
		_w12340_
	);
	LUT2 #(
		.INIT('h4)
	) name11879 (
		_w12339_,
		_w12340_,
		_w12341_
	);
	LUT2 #(
		.INIT('h2)
	) name11880 (
		\P1_state_reg[0]/NET0131 ,
		_w12341_,
		_w12342_
	);
	LUT2 #(
		.INIT('h1)
	) name11881 (
		_w7238_,
		_w12342_,
		_w12343_
	);
	LUT2 #(
		.INIT('h4)
	) name11882 (
		\P1_addr_reg[8]/NET0131 ,
		_w11399_,
		_w12344_
	);
	LUT2 #(
		.INIT('h1)
	) name11883 (
		_w1271_,
		_w11399_,
		_w12345_
	);
	LUT2 #(
		.INIT('h1)
	) name11884 (
		_w537_,
		_w12344_,
		_w12346_
	);
	LUT2 #(
		.INIT('h4)
	) name11885 (
		_w12345_,
		_w12346_,
		_w12347_
	);
	LUT2 #(
		.INIT('h1)
	) name11886 (
		_w11494_,
		_w11496_,
		_w12348_
	);
	LUT2 #(
		.INIT('h2)
	) name11887 (
		_w11672_,
		_w12348_,
		_w12349_
	);
	LUT2 #(
		.INIT('h4)
	) name11888 (
		_w11672_,
		_w12348_,
		_w12350_
	);
	LUT2 #(
		.INIT('h2)
	) name11889 (
		_w11437_,
		_w12349_,
		_w12351_
	);
	LUT2 #(
		.INIT('h4)
	) name11890 (
		_w12350_,
		_w12351_,
		_w12352_
	);
	LUT2 #(
		.INIT('h1)
	) name11891 (
		_w11478_,
		_w11480_,
		_w12353_
	);
	LUT2 #(
		.INIT('h2)
	) name11892 (
		_w11662_,
		_w12353_,
		_w12354_
	);
	LUT2 #(
		.INIT('h4)
	) name11893 (
		_w11662_,
		_w12353_,
		_w12355_
	);
	LUT2 #(
		.INIT('h2)
	) name11894 (
		_w11404_,
		_w12354_,
		_w12356_
	);
	LUT2 #(
		.INIT('h4)
	) name11895 (
		_w12355_,
		_w12356_,
		_w12357_
	);
	LUT2 #(
		.INIT('h1)
	) name11896 (
		_w12347_,
		_w12352_,
		_w12358_
	);
	LUT2 #(
		.INIT('h4)
	) name11897 (
		_w12357_,
		_w12358_,
		_w12359_
	);
	LUT2 #(
		.INIT('h2)
	) name11898 (
		\P1_state_reg[0]/NET0131 ,
		_w12359_,
		_w12360_
	);
	LUT2 #(
		.INIT('h1)
	) name11899 (
		_w8283_,
		_w12360_,
		_w12361_
	);
	LUT2 #(
		.INIT('h2)
	) name11900 (
		\P1_reg3_reg[1]/NET0131 ,
		\P1_state_reg[0]/NET0131 ,
		_w12362_
	);
	LUT2 #(
		.INIT('h8)
	) name11901 (
		_w1645_,
		_w11527_,
		_w12363_
	);
	LUT2 #(
		.INIT('h1)
	) name11902 (
		\P1_addr_reg[1]/NET0131 ,
		_w3448_,
		_w12364_
	);
	LUT2 #(
		.INIT('h4)
	) name11903 (
		_w1645_,
		_w3448_,
		_w12365_
	);
	LUT2 #(
		.INIT('h2)
	) name11904 (
		_w538_,
		_w12364_,
		_w12366_
	);
	LUT2 #(
		.INIT('h4)
	) name11905 (
		_w12365_,
		_w12366_,
		_w12367_
	);
	LUT2 #(
		.INIT('h1)
	) name11906 (
		_w11416_,
		_w11417_,
		_w12368_
	);
	LUT2 #(
		.INIT('h1)
	) name11907 (
		_w11418_,
		_w12368_,
		_w12369_
	);
	LUT2 #(
		.INIT('h8)
	) name11908 (
		_w11418_,
		_w12368_,
		_w12370_
	);
	LUT2 #(
		.INIT('h1)
	) name11909 (
		_w12369_,
		_w12370_,
		_w12371_
	);
	LUT2 #(
		.INIT('h8)
	) name11910 (
		_w11404_,
		_w12371_,
		_w12372_
	);
	LUT2 #(
		.INIT('h1)
	) name11911 (
		_w11449_,
		_w11450_,
		_w12373_
	);
	LUT2 #(
		.INIT('h1)
	) name11912 (
		_w11451_,
		_w12373_,
		_w12374_
	);
	LUT2 #(
		.INIT('h8)
	) name11913 (
		_w11451_,
		_w12373_,
		_w12375_
	);
	LUT2 #(
		.INIT('h1)
	) name11914 (
		_w12374_,
		_w12375_,
		_w12376_
	);
	LUT2 #(
		.INIT('h8)
	) name11915 (
		_w11437_,
		_w12376_,
		_w12377_
	);
	LUT2 #(
		.INIT('h1)
	) name11916 (
		_w12363_,
		_w12372_,
		_w12378_
	);
	LUT2 #(
		.INIT('h4)
	) name11917 (
		_w12377_,
		_w12378_,
		_w12379_
	);
	LUT2 #(
		.INIT('h4)
	) name11918 (
		_w12367_,
		_w12379_,
		_w12380_
	);
	LUT2 #(
		.INIT('h2)
	) name11919 (
		\P1_state_reg[0]/NET0131 ,
		_w12380_,
		_w12381_
	);
	LUT2 #(
		.INIT('h1)
	) name11920 (
		_w12362_,
		_w12381_,
		_w12382_
	);
	LUT2 #(
		.INIT('h4)
	) name11921 (
		_w1584_,
		_w11527_,
		_w12383_
	);
	LUT2 #(
		.INIT('h1)
	) name11922 (
		\P1_addr_reg[4]/NET0131 ,
		_w3448_,
		_w12384_
	);
	LUT2 #(
		.INIT('h8)
	) name11923 (
		_w1584_,
		_w3448_,
		_w12385_
	);
	LUT2 #(
		.INIT('h2)
	) name11924 (
		_w538_,
		_w12384_,
		_w12386_
	);
	LUT2 #(
		.INIT('h4)
	) name11925 (
		_w12385_,
		_w12386_,
		_w12387_
	);
	LUT2 #(
		.INIT('h1)
	) name11926 (
		_w11444_,
		_w11460_,
		_w12388_
	);
	LUT2 #(
		.INIT('h1)
	) name11927 (
		_w11457_,
		_w12388_,
		_w12389_
	);
	LUT2 #(
		.INIT('h8)
	) name11928 (
		_w11457_,
		_w12388_,
		_w12390_
	);
	LUT2 #(
		.INIT('h1)
	) name11929 (
		_w12389_,
		_w12390_,
		_w12391_
	);
	LUT2 #(
		.INIT('h8)
	) name11930 (
		_w11437_,
		_w12391_,
		_w12392_
	);
	LUT2 #(
		.INIT('h1)
	) name11931 (
		_w11411_,
		_w11427_,
		_w12393_
	);
	LUT2 #(
		.INIT('h1)
	) name11932 (
		_w11424_,
		_w12393_,
		_w12394_
	);
	LUT2 #(
		.INIT('h8)
	) name11933 (
		_w11424_,
		_w12393_,
		_w12395_
	);
	LUT2 #(
		.INIT('h1)
	) name11934 (
		_w12394_,
		_w12395_,
		_w12396_
	);
	LUT2 #(
		.INIT('h8)
	) name11935 (
		_w11404_,
		_w12396_,
		_w12397_
	);
	LUT2 #(
		.INIT('h1)
	) name11936 (
		_w12383_,
		_w12392_,
		_w12398_
	);
	LUT2 #(
		.INIT('h4)
	) name11937 (
		_w12397_,
		_w12398_,
		_w12399_
	);
	LUT2 #(
		.INIT('h4)
	) name11938 (
		_w12387_,
		_w12399_,
		_w12400_
	);
	LUT2 #(
		.INIT('h2)
	) name11939 (
		\P1_state_reg[0]/NET0131 ,
		_w12400_,
		_w12401_
	);
	LUT2 #(
		.INIT('h1)
	) name11940 (
		_w9016_,
		_w12401_,
		_w12402_
	);
	LUT2 #(
		.INIT('h1)
	) name11941 (
		_w11425_,
		_w11427_,
		_w12403_
	);
	LUT2 #(
		.INIT('h1)
	) name11942 (
		_w11410_,
		_w11426_,
		_w12404_
	);
	LUT2 #(
		.INIT('h1)
	) name11943 (
		_w12403_,
		_w12404_,
		_w12405_
	);
	LUT2 #(
		.INIT('h4)
	) name11944 (
		_w11410_,
		_w11429_,
		_w12406_
	);
	LUT2 #(
		.INIT('h2)
	) name11945 (
		_w11404_,
		_w12405_,
		_w12407_
	);
	LUT2 #(
		.INIT('h4)
	) name11946 (
		_w12406_,
		_w12407_,
		_w12408_
	);
	LUT2 #(
		.INIT('h1)
	) name11947 (
		_w11458_,
		_w11460_,
		_w12409_
	);
	LUT2 #(
		.INIT('h1)
	) name11948 (
		_w11443_,
		_w11459_,
		_w12410_
	);
	LUT2 #(
		.INIT('h1)
	) name11949 (
		_w12409_,
		_w12410_,
		_w12411_
	);
	LUT2 #(
		.INIT('h4)
	) name11950 (
		_w11443_,
		_w11462_,
		_w12412_
	);
	LUT2 #(
		.INIT('h2)
	) name11951 (
		_w11437_,
		_w12411_,
		_w12413_
	);
	LUT2 #(
		.INIT('h4)
	) name11952 (
		_w12412_,
		_w12413_,
		_w12414_
	);
	LUT2 #(
		.INIT('h4)
	) name11953 (
		\P1_addr_reg[5]/NET0131 ,
		_w11399_,
		_w12415_
	);
	LUT2 #(
		.INIT('h2)
	) name11954 (
		_w1560_,
		_w11399_,
		_w12416_
	);
	LUT2 #(
		.INIT('h1)
	) name11955 (
		_w537_,
		_w12415_,
		_w12417_
	);
	LUT2 #(
		.INIT('h4)
	) name11956 (
		_w12416_,
		_w12417_,
		_w12418_
	);
	LUT2 #(
		.INIT('h1)
	) name11957 (
		_w12408_,
		_w12414_,
		_w12419_
	);
	LUT2 #(
		.INIT('h4)
	) name11958 (
		_w12418_,
		_w12419_,
		_w12420_
	);
	LUT2 #(
		.INIT('h2)
	) name11959 (
		\P1_state_reg[0]/NET0131 ,
		_w12420_,
		_w12421_
	);
	LUT2 #(
		.INIT('h1)
	) name11960 (
		_w9058_,
		_w12421_,
		_w12422_
	);
	LUT2 #(
		.INIT('h4)
	) name11961 (
		\P1_state_reg[0]/NET0131 ,
		\P2_reg3_reg[18]/NET0131 ,
		_w12423_
	);
	LUT2 #(
		.INIT('h8)
	) name11962 (
		\P2_reg1_reg[18]/NET0131 ,
		_w2404_,
		_w12424_
	);
	LUT2 #(
		.INIT('h1)
	) name11963 (
		\P2_reg1_reg[18]/NET0131 ,
		_w2404_,
		_w12425_
	);
	LUT2 #(
		.INIT('h1)
	) name11964 (
		_w12424_,
		_w12425_,
		_w12426_
	);
	LUT2 #(
		.INIT('h4)
	) name11965 (
		_w12052_,
		_w12057_,
		_w12427_
	);
	LUT2 #(
		.INIT('h1)
	) name11966 (
		_w12051_,
		_w12082_,
		_w12428_
	);
	LUT2 #(
		.INIT('h4)
	) name11967 (
		_w12427_,
		_w12428_,
		_w12429_
	);
	LUT2 #(
		.INIT('h1)
	) name11968 (
		_w12081_,
		_w12429_,
		_w12430_
	);
	LUT2 #(
		.INIT('h1)
	) name11969 (
		_w12426_,
		_w12430_,
		_w12431_
	);
	LUT2 #(
		.INIT('h8)
	) name11970 (
		_w12426_,
		_w12430_,
		_w12432_
	);
	LUT2 #(
		.INIT('h2)
	) name11971 (
		_w11626_,
		_w12431_,
		_w12433_
	);
	LUT2 #(
		.INIT('h4)
	) name11972 (
		_w12432_,
		_w12433_,
		_w12434_
	);
	LUT2 #(
		.INIT('h4)
	) name11973 (
		\P2_addr_reg[18]/NET0131 ,
		_w11729_,
		_w12435_
	);
	LUT2 #(
		.INIT('h1)
	) name11974 (
		_w2404_,
		_w11729_,
		_w12436_
	);
	LUT2 #(
		.INIT('h1)
	) name11975 (
		_w2058_,
		_w12435_,
		_w12437_
	);
	LUT2 #(
		.INIT('h4)
	) name11976 (
		_w12436_,
		_w12437_,
		_w12438_
	);
	LUT2 #(
		.INIT('h8)
	) name11977 (
		\P2_reg2_reg[18]/NET0131 ,
		_w2404_,
		_w12439_
	);
	LUT2 #(
		.INIT('h1)
	) name11978 (
		\P2_reg2_reg[18]/NET0131 ,
		_w2404_,
		_w12440_
	);
	LUT2 #(
		.INIT('h1)
	) name11979 (
		_w12439_,
		_w12440_,
		_w12441_
	);
	LUT2 #(
		.INIT('h4)
	) name11980 (
		_w12063_,
		_w12068_,
		_w12442_
	);
	LUT2 #(
		.INIT('h1)
	) name11981 (
		_w12062_,
		_w12093_,
		_w12443_
	);
	LUT2 #(
		.INIT('h4)
	) name11982 (
		_w12442_,
		_w12443_,
		_w12444_
	);
	LUT2 #(
		.INIT('h1)
	) name11983 (
		_w12092_,
		_w12444_,
		_w12445_
	);
	LUT2 #(
		.INIT('h1)
	) name11984 (
		_w12441_,
		_w12445_,
		_w12446_
	);
	LUT2 #(
		.INIT('h8)
	) name11985 (
		_w12441_,
		_w12445_,
		_w12447_
	);
	LUT2 #(
		.INIT('h2)
	) name11986 (
		_w11630_,
		_w12446_,
		_w12448_
	);
	LUT2 #(
		.INIT('h4)
	) name11987 (
		_w12447_,
		_w12448_,
		_w12449_
	);
	LUT2 #(
		.INIT('h1)
	) name11988 (
		_w12434_,
		_w12438_,
		_w12450_
	);
	LUT2 #(
		.INIT('h4)
	) name11989 (
		_w12449_,
		_w12450_,
		_w12451_
	);
	LUT2 #(
		.INIT('h2)
	) name11990 (
		\P1_state_reg[0]/NET0131 ,
		_w12451_,
		_w12452_
	);
	LUT2 #(
		.INIT('h1)
	) name11991 (
		_w12423_,
		_w12452_,
		_w12453_
	);
	LUT2 #(
		.INIT('h4)
	) name11992 (
		_w12081_,
		_w12087_,
		_w12454_
	);
	LUT2 #(
		.INIT('h1)
	) name11993 (
		_w12082_,
		_w12424_,
		_w12455_
	);
	LUT2 #(
		.INIT('h4)
	) name11994 (
		_w12454_,
		_w12455_,
		_w12456_
	);
	LUT2 #(
		.INIT('h1)
	) name11995 (
		_w12425_,
		_w12456_,
		_w12457_
	);
	LUT2 #(
		.INIT('h2)
	) name11996 (
		\P2_reg1_reg[19]/NET0131 ,
		_w12457_,
		_w12458_
	);
	LUT2 #(
		.INIT('h4)
	) name11997 (
		\P2_reg1_reg[19]/NET0131 ,
		_w12457_,
		_w12459_
	);
	LUT2 #(
		.INIT('h1)
	) name11998 (
		_w12458_,
		_w12459_,
		_w12460_
	);
	LUT2 #(
		.INIT('h2)
	) name11999 (
		_w2258_,
		_w12460_,
		_w12461_
	);
	LUT2 #(
		.INIT('h4)
	) name12000 (
		_w2258_,
		_w12460_,
		_w12462_
	);
	LUT2 #(
		.INIT('h2)
	) name12001 (
		_w11626_,
		_w12461_,
		_w12463_
	);
	LUT2 #(
		.INIT('h4)
	) name12002 (
		_w12462_,
		_w12463_,
		_w12464_
	);
	LUT2 #(
		.INIT('h4)
	) name12003 (
		\P2_addr_reg[19]/NET0131 ,
		_w11729_,
		_w12465_
	);
	LUT2 #(
		.INIT('h1)
	) name12004 (
		_w2258_,
		_w11729_,
		_w12466_
	);
	LUT2 #(
		.INIT('h1)
	) name12005 (
		_w2058_,
		_w12465_,
		_w12467_
	);
	LUT2 #(
		.INIT('h4)
	) name12006 (
		_w12466_,
		_w12467_,
		_w12468_
	);
	LUT2 #(
		.INIT('h4)
	) name12007 (
		_w12092_,
		_w12098_,
		_w12469_
	);
	LUT2 #(
		.INIT('h1)
	) name12008 (
		_w12093_,
		_w12439_,
		_w12470_
	);
	LUT2 #(
		.INIT('h4)
	) name12009 (
		_w12469_,
		_w12470_,
		_w12471_
	);
	LUT2 #(
		.INIT('h1)
	) name12010 (
		_w12440_,
		_w12471_,
		_w12472_
	);
	LUT2 #(
		.INIT('h8)
	) name12011 (
		\P2_reg2_reg[19]/NET0131 ,
		_w12472_,
		_w12473_
	);
	LUT2 #(
		.INIT('h1)
	) name12012 (
		\P2_reg2_reg[19]/NET0131 ,
		_w12472_,
		_w12474_
	);
	LUT2 #(
		.INIT('h1)
	) name12013 (
		_w12473_,
		_w12474_,
		_w12475_
	);
	LUT2 #(
		.INIT('h8)
	) name12014 (
		_w2258_,
		_w12475_,
		_w12476_
	);
	LUT2 #(
		.INIT('h1)
	) name12015 (
		_w2258_,
		_w12475_,
		_w12477_
	);
	LUT2 #(
		.INIT('h2)
	) name12016 (
		_w11630_,
		_w12476_,
		_w12478_
	);
	LUT2 #(
		.INIT('h4)
	) name12017 (
		_w12477_,
		_w12478_,
		_w12479_
	);
	LUT2 #(
		.INIT('h1)
	) name12018 (
		_w12464_,
		_w12468_,
		_w12480_
	);
	LUT2 #(
		.INIT('h4)
	) name12019 (
		_w12479_,
		_w12480_,
		_w12481_
	);
	LUT2 #(
		.INIT('h2)
	) name12020 (
		\P1_state_reg[0]/NET0131 ,
		_w12481_,
		_w12482_
	);
	LUT2 #(
		.INIT('h1)
	) name12021 (
		_w5602_,
		_w12482_,
		_w12483_
	);
	LUT2 #(
		.INIT('h8)
	) name12022 (
		\P1_reg1_reg[18]/NET0131 ,
		_w1384_,
		_w12484_
	);
	LUT2 #(
		.INIT('h1)
	) name12023 (
		\P1_reg1_reg[18]/NET0131 ,
		_w1384_,
		_w12485_
	);
	LUT2 #(
		.INIT('h1)
	) name12024 (
		_w12484_,
		_w12485_,
		_w12486_
	);
	LUT2 #(
		.INIT('h4)
	) name12025 (
		_w12112_,
		_w12117_,
		_w12487_
	);
	LUT2 #(
		.INIT('h1)
	) name12026 (
		_w12111_,
		_w12174_,
		_w12488_
	);
	LUT2 #(
		.INIT('h4)
	) name12027 (
		_w12487_,
		_w12488_,
		_w12489_
	);
	LUT2 #(
		.INIT('h1)
	) name12028 (
		_w12173_,
		_w12489_,
		_w12490_
	);
	LUT2 #(
		.INIT('h1)
	) name12029 (
		_w12486_,
		_w12490_,
		_w12491_
	);
	LUT2 #(
		.INIT('h8)
	) name12030 (
		_w12486_,
		_w12490_,
		_w12492_
	);
	LUT2 #(
		.INIT('h2)
	) name12031 (
		_w11404_,
		_w12491_,
		_w12493_
	);
	LUT2 #(
		.INIT('h4)
	) name12032 (
		_w12492_,
		_w12493_,
		_w12494_
	);
	LUT2 #(
		.INIT('h4)
	) name12033 (
		\P1_addr_reg[18]/NET0131 ,
		_w11399_,
		_w12495_
	);
	LUT2 #(
		.INIT('h1)
	) name12034 (
		_w1384_,
		_w11399_,
		_w12496_
	);
	LUT2 #(
		.INIT('h1)
	) name12035 (
		_w537_,
		_w12495_,
		_w12497_
	);
	LUT2 #(
		.INIT('h4)
	) name12036 (
		_w12496_,
		_w12497_,
		_w12498_
	);
	LUT2 #(
		.INIT('h8)
	) name12037 (
		\P1_reg2_reg[18]/NET0131 ,
		_w1384_,
		_w12499_
	);
	LUT2 #(
		.INIT('h1)
	) name12038 (
		\P1_reg2_reg[18]/NET0131 ,
		_w1384_,
		_w12500_
	);
	LUT2 #(
		.INIT('h1)
	) name12039 (
		_w12499_,
		_w12500_,
		_w12501_
	);
	LUT2 #(
		.INIT('h4)
	) name12040 (
		_w12123_,
		_w12128_,
		_w12502_
	);
	LUT2 #(
		.INIT('h1)
	) name12041 (
		_w12122_,
		_w12163_,
		_w12503_
	);
	LUT2 #(
		.INIT('h4)
	) name12042 (
		_w12502_,
		_w12503_,
		_w12504_
	);
	LUT2 #(
		.INIT('h1)
	) name12043 (
		_w12162_,
		_w12504_,
		_w12505_
	);
	LUT2 #(
		.INIT('h1)
	) name12044 (
		_w12501_,
		_w12505_,
		_w12506_
	);
	LUT2 #(
		.INIT('h8)
	) name12045 (
		_w12501_,
		_w12505_,
		_w12507_
	);
	LUT2 #(
		.INIT('h2)
	) name12046 (
		_w11437_,
		_w12506_,
		_w12508_
	);
	LUT2 #(
		.INIT('h4)
	) name12047 (
		_w12507_,
		_w12508_,
		_w12509_
	);
	LUT2 #(
		.INIT('h1)
	) name12048 (
		_w12494_,
		_w12498_,
		_w12510_
	);
	LUT2 #(
		.INIT('h4)
	) name12049 (
		_w12509_,
		_w12510_,
		_w12511_
	);
	LUT2 #(
		.INIT('h2)
	) name12050 (
		\P1_state_reg[0]/NET0131 ,
		_w12511_,
		_w12512_
	);
	LUT2 #(
		.INIT('h1)
	) name12051 (
		_w5477_,
		_w12512_,
		_w12513_
	);
	LUT2 #(
		.INIT('h4)
	) name12052 (
		_w12173_,
		_w12179_,
		_w12514_
	);
	LUT2 #(
		.INIT('h1)
	) name12053 (
		_w12174_,
		_w12484_,
		_w12515_
	);
	LUT2 #(
		.INIT('h4)
	) name12054 (
		_w12514_,
		_w12515_,
		_w12516_
	);
	LUT2 #(
		.INIT('h1)
	) name12055 (
		_w12485_,
		_w12516_,
		_w12517_
	);
	LUT2 #(
		.INIT('h1)
	) name12056 (
		\P1_reg1_reg[19]/NET0131 ,
		_w1408_,
		_w12518_
	);
	LUT2 #(
		.INIT('h8)
	) name12057 (
		\P1_reg1_reg[19]/NET0131 ,
		_w1408_,
		_w12519_
	);
	LUT2 #(
		.INIT('h1)
	) name12058 (
		_w12518_,
		_w12519_,
		_w12520_
	);
	LUT2 #(
		.INIT('h1)
	) name12059 (
		_w12517_,
		_w12520_,
		_w12521_
	);
	LUT2 #(
		.INIT('h8)
	) name12060 (
		_w12517_,
		_w12520_,
		_w12522_
	);
	LUT2 #(
		.INIT('h2)
	) name12061 (
		_w11404_,
		_w12521_,
		_w12523_
	);
	LUT2 #(
		.INIT('h4)
	) name12062 (
		_w12522_,
		_w12523_,
		_w12524_
	);
	LUT2 #(
		.INIT('h4)
	) name12063 (
		\P1_addr_reg[19]/NET0131 ,
		_w11399_,
		_w12525_
	);
	LUT2 #(
		.INIT('h1)
	) name12064 (
		_w1408_,
		_w11399_,
		_w12526_
	);
	LUT2 #(
		.INIT('h1)
	) name12065 (
		_w537_,
		_w12525_,
		_w12527_
	);
	LUT2 #(
		.INIT('h4)
	) name12066 (
		_w12526_,
		_w12527_,
		_w12528_
	);
	LUT2 #(
		.INIT('h4)
	) name12067 (
		_w12162_,
		_w12168_,
		_w12529_
	);
	LUT2 #(
		.INIT('h1)
	) name12068 (
		_w12163_,
		_w12499_,
		_w12530_
	);
	LUT2 #(
		.INIT('h4)
	) name12069 (
		_w12529_,
		_w12530_,
		_w12531_
	);
	LUT2 #(
		.INIT('h1)
	) name12070 (
		_w12500_,
		_w12531_,
		_w12532_
	);
	LUT2 #(
		.INIT('h8)
	) name12071 (
		\P1_reg2_reg[19]/NET0131 ,
		_w12532_,
		_w12533_
	);
	LUT2 #(
		.INIT('h1)
	) name12072 (
		\P1_reg2_reg[19]/NET0131 ,
		_w12532_,
		_w12534_
	);
	LUT2 #(
		.INIT('h1)
	) name12073 (
		_w12533_,
		_w12534_,
		_w12535_
	);
	LUT2 #(
		.INIT('h8)
	) name12074 (
		_w1408_,
		_w12535_,
		_w12536_
	);
	LUT2 #(
		.INIT('h1)
	) name12075 (
		_w1408_,
		_w12535_,
		_w12537_
	);
	LUT2 #(
		.INIT('h2)
	) name12076 (
		_w11437_,
		_w12536_,
		_w12538_
	);
	LUT2 #(
		.INIT('h4)
	) name12077 (
		_w12537_,
		_w12538_,
		_w12539_
	);
	LUT2 #(
		.INIT('h1)
	) name12078 (
		_w12524_,
		_w12528_,
		_w12540_
	);
	LUT2 #(
		.INIT('h4)
	) name12079 (
		_w12539_,
		_w12540_,
		_w12541_
	);
	LUT2 #(
		.INIT('h2)
	) name12080 (
		\P1_state_reg[0]/NET0131 ,
		_w12541_,
		_w12542_
	);
	LUT2 #(
		.INIT('h1)
	) name12081 (
		_w5685_,
		_w12542_,
		_w12543_
	);
	LUT2 #(
		.INIT('h1)
	) name12082 (
		_w538_,
		_w3448_,
		_w12544_
	);
	LUT2 #(
		.INIT('h2)
	) name12083 (
		\P1_state_reg[0]/NET0131 ,
		_w12544_,
		_w12545_
	);
	LUT2 #(
		.INIT('h1)
	) name12084 (
		_w2024_,
		_w2059_,
		_w12546_
	);
	LUT2 #(
		.INIT('h2)
	) name12085 (
		\P1_state_reg[0]/NET0131 ,
		_w12546_,
		_w12547_
	);
	LUT2 #(
		.INIT('h8)
	) name12086 (
		\P1_state_reg[0]/NET0131 ,
		_w3448_,
		_w12548_
	);
	LUT2 #(
		.INIT('h8)
	) name12087 (
		\P1_state_reg[0]/NET0131 ,
		_w2024_,
		_w12549_
	);
	LUT2 #(
		.INIT('h2)
	) name12088 (
		_w2023_,
		_w3043_,
		_w12550_
	);
	LUT2 #(
		.INIT('h2)
	) name12089 (
		\P2_datao_reg[25]/NET0131 ,
		_w2023_,
		_w12551_
	);
	LUT2 #(
		.INIT('h1)
	) name12090 (
		_w12550_,
		_w12551_,
		_w12552_
	);
	LUT2 #(
		.INIT('h4)
	) name12091 (
		_w1038_,
		_w3447_,
		_w12553_
	);
	LUT2 #(
		.INIT('h2)
	) name12092 (
		\P1_datao_reg[25]/NET0131 ,
		_w3447_,
		_w12554_
	);
	LUT2 #(
		.INIT('h1)
	) name12093 (
		_w12553_,
		_w12554_,
		_w12555_
	);
	LUT2 #(
		.INIT('h2)
	) name12094 (
		\P2_reg1_reg[16]/NET0131 ,
		_w5961_,
		_w12556_
	);
	LUT2 #(
		.INIT('h8)
	) name12095 (
		\P2_reg1_reg[16]/NET0131 ,
		_w6642_,
		_w12557_
	);
	LUT2 #(
		.INIT('h8)
	) name12096 (
		_w3355_,
		_w6240_,
		_w12558_
	);
	LUT2 #(
		.INIT('h1)
	) name12097 (
		_w3177_,
		_w6226_,
		_w12559_
	);
	LUT2 #(
		.INIT('h8)
	) name12098 (
		_w3411_,
		_w6234_,
		_w12560_
	);
	LUT2 #(
		.INIT('h2)
	) name12099 (
		_w7983_,
		_w12558_,
		_w12561_
	);
	LUT2 #(
		.INIT('h1)
	) name12100 (
		_w12559_,
		_w12560_,
		_w12562_
	);
	LUT2 #(
		.INIT('h8)
	) name12101 (
		_w12561_,
		_w12562_,
		_w12563_
	);
	LUT2 #(
		.INIT('h2)
	) name12102 (
		_w3733_,
		_w12563_,
		_w12564_
	);
	LUT2 #(
		.INIT('h1)
	) name12103 (
		_w12557_,
		_w12564_,
		_w12565_
	);
	LUT2 #(
		.INIT('h2)
	) name12104 (
		_w5287_,
		_w12565_,
		_w12566_
	);
	LUT2 #(
		.INIT('h1)
	) name12105 (
		_w12556_,
		_w12566_,
		_w12567_
	);
	LUT2 #(
		.INIT('h8)
	) name12106 (
		_w2438_,
		_w3976_,
		_w12568_
	);
	LUT2 #(
		.INIT('h8)
	) name12107 (
		_w2024_,
		_w2438_,
		_w12569_
	);
	LUT2 #(
		.INIT('h2)
	) name12108 (
		_w2438_,
		_w3962_,
		_w12570_
	);
	LUT2 #(
		.INIT('h2)
	) name12109 (
		_w2438_,
		_w3788_,
		_w12571_
	);
	LUT2 #(
		.INIT('h8)
	) name12110 (
		_w3788_,
		_w6331_,
		_w12572_
	);
	LUT2 #(
		.INIT('h1)
	) name12111 (
		_w12571_,
		_w12572_,
		_w12573_
	);
	LUT2 #(
		.INIT('h2)
	) name12112 (
		_w3355_,
		_w12573_,
		_w12574_
	);
	LUT2 #(
		.INIT('h8)
	) name12113 (
		_w3788_,
		_w6337_,
		_w12575_
	);
	LUT2 #(
		.INIT('h1)
	) name12114 (
		_w12571_,
		_w12575_,
		_w12576_
	);
	LUT2 #(
		.INIT('h1)
	) name12115 (
		_w3177_,
		_w12576_,
		_w12577_
	);
	LUT2 #(
		.INIT('h2)
	) name12116 (
		_w3788_,
		_w6343_,
		_w12578_
	);
	LUT2 #(
		.INIT('h1)
	) name12117 (
		_w12571_,
		_w12578_,
		_w12579_
	);
	LUT2 #(
		.INIT('h1)
	) name12118 (
		_w3320_,
		_w12579_,
		_w12580_
	);
	LUT2 #(
		.INIT('h8)
	) name12119 (
		_w3788_,
		_w6351_,
		_w12581_
	);
	LUT2 #(
		.INIT('h1)
	) name12120 (
		_w12571_,
		_w12581_,
		_w12582_
	);
	LUT2 #(
		.INIT('h2)
	) name12121 (
		_w3411_,
		_w12582_,
		_w12583_
	);
	LUT2 #(
		.INIT('h2)
	) name12122 (
		_w2433_,
		_w3965_,
		_w12584_
	);
	LUT2 #(
		.INIT('h1)
	) name12123 (
		_w12570_,
		_w12584_,
		_w12585_
	);
	LUT2 #(
		.INIT('h4)
	) name12124 (
		_w12583_,
		_w12585_,
		_w12586_
	);
	LUT2 #(
		.INIT('h4)
	) name12125 (
		_w12577_,
		_w12586_,
		_w12587_
	);
	LUT2 #(
		.INIT('h4)
	) name12126 (
		_w12580_,
		_w12587_,
		_w12588_
	);
	LUT2 #(
		.INIT('h4)
	) name12127 (
		_w12574_,
		_w12588_,
		_w12589_
	);
	LUT2 #(
		.INIT('h2)
	) name12128 (
		_w2026_,
		_w12589_,
		_w12590_
	);
	LUT2 #(
		.INIT('h1)
	) name12129 (
		_w12569_,
		_w12590_,
		_w12591_
	);
	LUT2 #(
		.INIT('h2)
	) name12130 (
		\P1_state_reg[0]/NET0131 ,
		_w12591_,
		_w12592_
	);
	LUT2 #(
		.INIT('h1)
	) name12131 (
		_w12423_,
		_w12568_,
		_w12593_
	);
	LUT2 #(
		.INIT('h4)
	) name12132 (
		_w12592_,
		_w12593_,
		_w12594_
	);
	LUT2 #(
		.INIT('h2)
	) name12133 (
		_w997_,
		_w4067_,
		_w12595_
	);
	LUT2 #(
		.INIT('h2)
	) name12134 (
		_w1002_,
		_w3980_,
		_w12596_
	);
	LUT2 #(
		.INIT('h2)
	) name12135 (
		_w3980_,
		_w5948_,
		_w12597_
	);
	LUT2 #(
		.INIT('h1)
	) name12136 (
		_w12596_,
		_w12597_,
		_w12598_
	);
	LUT2 #(
		.INIT('h1)
	) name12137 (
		_w3563_,
		_w12598_,
		_w12599_
	);
	LUT2 #(
		.INIT('h2)
	) name12138 (
		_w3980_,
		_w5930_,
		_w12600_
	);
	LUT2 #(
		.INIT('h1)
	) name12139 (
		_w12596_,
		_w12600_,
		_w12601_
	);
	LUT2 #(
		.INIT('h1)
	) name12140 (
		_w3677_,
		_w12601_,
		_w12602_
	);
	LUT2 #(
		.INIT('h2)
	) name12141 (
		_w3980_,
		_w5903_,
		_w12603_
	);
	LUT2 #(
		.INIT('h1)
	) name12142 (
		_w12596_,
		_w12603_,
		_w12604_
	);
	LUT2 #(
		.INIT('h2)
	) name12143 (
		_w1936_,
		_w12604_,
		_w12605_
	);
	LUT2 #(
		.INIT('h8)
	) name12144 (
		_w3980_,
		_w5908_,
		_w12606_
	);
	LUT2 #(
		.INIT('h1)
	) name12145 (
		_w12596_,
		_w12606_,
		_w12607_
	);
	LUT2 #(
		.INIT('h2)
	) name12146 (
		_w3712_,
		_w12607_,
		_w12608_
	);
	LUT2 #(
		.INIT('h2)
	) name12147 (
		_w1002_,
		_w4064_,
		_w12609_
	);
	LUT2 #(
		.INIT('h1)
	) name12148 (
		_w12595_,
		_w12609_,
		_w12610_
	);
	LUT2 #(
		.INIT('h4)
	) name12149 (
		_w12608_,
		_w12610_,
		_w12611_
	);
	LUT2 #(
		.INIT('h4)
	) name12150 (
		_w12599_,
		_w12611_,
		_w12612_
	);
	LUT2 #(
		.INIT('h1)
	) name12151 (
		_w12602_,
		_w12605_,
		_w12613_
	);
	LUT2 #(
		.INIT('h8)
	) name12152 (
		_w12612_,
		_w12613_,
		_w12614_
	);
	LUT2 #(
		.INIT('h2)
	) name12153 (
		_w5812_,
		_w12614_,
		_w12615_
	);
	LUT2 #(
		.INIT('h2)
	) name12154 (
		\P1_reg3_reg[26]/NET0131 ,
		\P1_state_reg[0]/NET0131 ,
		_w12616_
	);
	LUT2 #(
		.INIT('h2)
	) name12155 (
		\P1_state_reg[0]/NET0131 ,
		_w3450_,
		_w12617_
	);
	LUT2 #(
		.INIT('h8)
	) name12156 (
		_w1002_,
		_w12617_,
		_w12618_
	);
	LUT2 #(
		.INIT('h1)
	) name12157 (
		_w12616_,
		_w12618_,
		_w12619_
	);
	LUT2 #(
		.INIT('h4)
	) name12158 (
		_w12615_,
		_w12619_,
		_w12620_
	);
	LUT2 #(
		.INIT('h2)
	) name12159 (
		\P2_reg2_reg[15]/NET0131 ,
		_w1983_,
		_w12621_
	);
	LUT2 #(
		.INIT('h8)
	) name12160 (
		\P2_reg2_reg[15]/NET0131 ,
		_w2024_,
		_w12622_
	);
	LUT2 #(
		.INIT('h8)
	) name12161 (
		_w2822_,
		_w3420_,
		_w12623_
	);
	LUT2 #(
		.INIT('h2)
	) name12162 (
		\P2_reg2_reg[15]/NET0131 ,
		_w3758_,
		_w12624_
	);
	LUT2 #(
		.INIT('h8)
	) name12163 (
		_w3758_,
		_w8211_,
		_w12625_
	);
	LUT2 #(
		.INIT('h1)
	) name12164 (
		_w12624_,
		_w12625_,
		_w12626_
	);
	LUT2 #(
		.INIT('h2)
	) name12165 (
		_w3411_,
		_w12626_,
		_w12627_
	);
	LUT2 #(
		.INIT('h8)
	) name12166 (
		_w3758_,
		_w8217_,
		_w12628_
	);
	LUT2 #(
		.INIT('h1)
	) name12167 (
		_w12624_,
		_w12628_,
		_w12629_
	);
	LUT2 #(
		.INIT('h1)
	) name12168 (
		_w3177_,
		_w12629_,
		_w12630_
	);
	LUT2 #(
		.INIT('h2)
	) name12169 (
		\P2_reg2_reg[15]/NET0131 ,
		_w7770_,
		_w12631_
	);
	LUT2 #(
		.INIT('h2)
	) name12170 (
		_w3758_,
		_w9361_,
		_w12632_
	);
	LUT2 #(
		.INIT('h8)
	) name12171 (
		_w3758_,
		_w8222_,
		_w12633_
	);
	LUT2 #(
		.INIT('h1)
	) name12172 (
		_w12624_,
		_w12633_,
		_w12634_
	);
	LUT2 #(
		.INIT('h2)
	) name12173 (
		_w3355_,
		_w12634_,
		_w12635_
	);
	LUT2 #(
		.INIT('h1)
	) name12174 (
		_w12623_,
		_w12631_,
		_w12636_
	);
	LUT2 #(
		.INIT('h4)
	) name12175 (
		_w12632_,
		_w12636_,
		_w12637_
	);
	LUT2 #(
		.INIT('h4)
	) name12176 (
		_w12635_,
		_w12637_,
		_w12638_
	);
	LUT2 #(
		.INIT('h4)
	) name12177 (
		_w12627_,
		_w12638_,
		_w12639_
	);
	LUT2 #(
		.INIT('h4)
	) name12178 (
		_w12630_,
		_w12639_,
		_w12640_
	);
	LUT2 #(
		.INIT('h2)
	) name12179 (
		_w2026_,
		_w12640_,
		_w12641_
	);
	LUT2 #(
		.INIT('h1)
	) name12180 (
		_w12622_,
		_w12641_,
		_w12642_
	);
	LUT2 #(
		.INIT('h2)
	) name12181 (
		\P1_state_reg[0]/NET0131 ,
		_w12642_,
		_w12643_
	);
	LUT2 #(
		.INIT('h1)
	) name12182 (
		_w12621_,
		_w12643_,
		_w12644_
	);
	LUT2 #(
		.INIT('h2)
	) name12183 (
		\P2_reg2_reg[24]/NET0131 ,
		_w1983_,
		_w12645_
	);
	LUT2 #(
		.INIT('h8)
	) name12184 (
		\P2_reg2_reg[24]/NET0131 ,
		_w2024_,
		_w12646_
	);
	LUT2 #(
		.INIT('h2)
	) name12185 (
		\P2_reg2_reg[24]/NET0131 ,
		_w3758_,
		_w12647_
	);
	LUT2 #(
		.INIT('h2)
	) name12186 (
		_w3758_,
		_w4983_,
		_w12648_
	);
	LUT2 #(
		.INIT('h1)
	) name12187 (
		_w12647_,
		_w12648_,
		_w12649_
	);
	LUT2 #(
		.INIT('h1)
	) name12188 (
		_w3320_,
		_w12649_,
		_w12650_
	);
	LUT2 #(
		.INIT('h2)
	) name12189 (
		_w3758_,
		_w4997_,
		_w12651_
	);
	LUT2 #(
		.INIT('h1)
	) name12190 (
		_w12647_,
		_w12651_,
		_w12652_
	);
	LUT2 #(
		.INIT('h1)
	) name12191 (
		_w3177_,
		_w12652_,
		_w12653_
	);
	LUT2 #(
		.INIT('h8)
	) name12192 (
		_w3758_,
		_w5002_,
		_w12654_
	);
	LUT2 #(
		.INIT('h1)
	) name12193 (
		_w12647_,
		_w12654_,
		_w12655_
	);
	LUT2 #(
		.INIT('h2)
	) name12194 (
		_w3355_,
		_w12655_,
		_w12656_
	);
	LUT2 #(
		.INIT('h8)
	) name12195 (
		_w3758_,
		_w5008_,
		_w12657_
	);
	LUT2 #(
		.INIT('h1)
	) name12196 (
		_w12647_,
		_w12657_,
		_w12658_
	);
	LUT2 #(
		.INIT('h2)
	) name12197 (
		_w3411_,
		_w12658_,
		_w12659_
	);
	LUT2 #(
		.INIT('h8)
	) name12198 (
		_w3758_,
		_w5010_,
		_w12660_
	);
	LUT2 #(
		.INIT('h8)
	) name12199 (
		_w3058_,
		_w3420_,
		_w12661_
	);
	LUT2 #(
		.INIT('h2)
	) name12200 (
		\P2_reg2_reg[24]/NET0131 ,
		_w3774_,
		_w12662_
	);
	LUT2 #(
		.INIT('h1)
	) name12201 (
		_w12661_,
		_w12662_,
		_w12663_
	);
	LUT2 #(
		.INIT('h4)
	) name12202 (
		_w12660_,
		_w12663_,
		_w12664_
	);
	LUT2 #(
		.INIT('h4)
	) name12203 (
		_w12656_,
		_w12664_,
		_w12665_
	);
	LUT2 #(
		.INIT('h4)
	) name12204 (
		_w12659_,
		_w12665_,
		_w12666_
	);
	LUT2 #(
		.INIT('h4)
	) name12205 (
		_w12653_,
		_w12666_,
		_w12667_
	);
	LUT2 #(
		.INIT('h4)
	) name12206 (
		_w12650_,
		_w12667_,
		_w12668_
	);
	LUT2 #(
		.INIT('h2)
	) name12207 (
		_w2026_,
		_w12668_,
		_w12669_
	);
	LUT2 #(
		.INIT('h1)
	) name12208 (
		_w12646_,
		_w12669_,
		_w12670_
	);
	LUT2 #(
		.INIT('h2)
	) name12209 (
		\P1_state_reg[0]/NET0131 ,
		_w12670_,
		_w12671_
	);
	LUT2 #(
		.INIT('h1)
	) name12210 (
		_w12645_,
		_w12671_,
		_w12672_
	);
	LUT2 #(
		.INIT('h1)
	) name12211 (
		\P1_rd_reg/NET0131 ,
		\P2_rd_reg/NET0131 ,
		_w12673_
	);
	LUT2 #(
		.INIT('h8)
	) name12212 (
		\P1_rd_reg/NET0131 ,
		\P2_rd_reg/NET0131 ,
		_w12674_
	);
	LUT2 #(
		.INIT('h1)
	) name12213 (
		_w12673_,
		_w12674_,
		_w12675_
	);
	LUT2 #(
		.INIT('h8)
	) name12214 (
		\P1_addr_reg[0]/NET0131 ,
		\P2_addr_reg[0]/NET0131 ,
		_w12676_
	);
	LUT2 #(
		.INIT('h1)
	) name12215 (
		\P1_addr_reg[0]/NET0131 ,
		\P2_addr_reg[0]/NET0131 ,
		_w12677_
	);
	LUT2 #(
		.INIT('h1)
	) name12216 (
		_w12676_,
		_w12677_,
		_w12678_
	);
	LUT2 #(
		.INIT('h8)
	) name12217 (
		\P1_addr_reg[10]/NET0131 ,
		\P2_addr_reg[10]/NET0131 ,
		_w12679_
	);
	LUT2 #(
		.INIT('h1)
	) name12218 (
		\P1_addr_reg[10]/NET0131 ,
		\P2_addr_reg[10]/NET0131 ,
		_w12680_
	);
	LUT2 #(
		.INIT('h1)
	) name12219 (
		_w12679_,
		_w12680_,
		_w12681_
	);
	LUT2 #(
		.INIT('h1)
	) name12220 (
		\P1_addr_reg[9]/NET0131 ,
		\P2_addr_reg[9]/NET0131 ,
		_w12682_
	);
	LUT2 #(
		.INIT('h8)
	) name12221 (
		\P1_addr_reg[9]/NET0131 ,
		\P2_addr_reg[9]/NET0131 ,
		_w12683_
	);
	LUT2 #(
		.INIT('h1)
	) name12222 (
		\P1_addr_reg[8]/NET0131 ,
		\P2_addr_reg[8]/NET0131 ,
		_w12684_
	);
	LUT2 #(
		.INIT('h8)
	) name12223 (
		\P1_addr_reg[8]/NET0131 ,
		\P2_addr_reg[8]/NET0131 ,
		_w12685_
	);
	LUT2 #(
		.INIT('h1)
	) name12224 (
		\P1_addr_reg[7]/NET0131 ,
		\P2_addr_reg[7]/NET0131 ,
		_w12686_
	);
	LUT2 #(
		.INIT('h8)
	) name12225 (
		\P1_addr_reg[7]/NET0131 ,
		\P2_addr_reg[7]/NET0131 ,
		_w12687_
	);
	LUT2 #(
		.INIT('h1)
	) name12226 (
		\P1_addr_reg[6]/NET0131 ,
		\P2_addr_reg[6]/NET0131 ,
		_w12688_
	);
	LUT2 #(
		.INIT('h8)
	) name12227 (
		\P1_addr_reg[6]/NET0131 ,
		\P2_addr_reg[6]/NET0131 ,
		_w12689_
	);
	LUT2 #(
		.INIT('h1)
	) name12228 (
		\P1_addr_reg[5]/NET0131 ,
		\P2_addr_reg[5]/NET0131 ,
		_w12690_
	);
	LUT2 #(
		.INIT('h8)
	) name12229 (
		\P1_addr_reg[5]/NET0131 ,
		\P2_addr_reg[5]/NET0131 ,
		_w12691_
	);
	LUT2 #(
		.INIT('h1)
	) name12230 (
		\P1_addr_reg[4]/NET0131 ,
		\P2_addr_reg[4]/NET0131 ,
		_w12692_
	);
	LUT2 #(
		.INIT('h8)
	) name12231 (
		\P1_addr_reg[4]/NET0131 ,
		\P2_addr_reg[4]/NET0131 ,
		_w12693_
	);
	LUT2 #(
		.INIT('h1)
	) name12232 (
		\P1_addr_reg[3]/NET0131 ,
		\P2_addr_reg[3]/NET0131 ,
		_w12694_
	);
	LUT2 #(
		.INIT('h8)
	) name12233 (
		\P1_addr_reg[3]/NET0131 ,
		\P2_addr_reg[3]/NET0131 ,
		_w12695_
	);
	LUT2 #(
		.INIT('h1)
	) name12234 (
		\P1_addr_reg[2]/NET0131 ,
		\P2_addr_reg[2]/NET0131 ,
		_w12696_
	);
	LUT2 #(
		.INIT('h8)
	) name12235 (
		\P1_addr_reg[2]/NET0131 ,
		\P2_addr_reg[2]/NET0131 ,
		_w12697_
	);
	LUT2 #(
		.INIT('h1)
	) name12236 (
		\P1_addr_reg[1]/NET0131 ,
		\P2_addr_reg[1]/NET0131 ,
		_w12698_
	);
	LUT2 #(
		.INIT('h8)
	) name12237 (
		\P1_addr_reg[1]/NET0131 ,
		\P2_addr_reg[1]/NET0131 ,
		_w12699_
	);
	LUT2 #(
		.INIT('h1)
	) name12238 (
		_w12676_,
		_w12699_,
		_w12700_
	);
	LUT2 #(
		.INIT('h1)
	) name12239 (
		_w12698_,
		_w12700_,
		_w12701_
	);
	LUT2 #(
		.INIT('h1)
	) name12240 (
		_w12697_,
		_w12701_,
		_w12702_
	);
	LUT2 #(
		.INIT('h1)
	) name12241 (
		_w12696_,
		_w12702_,
		_w12703_
	);
	LUT2 #(
		.INIT('h1)
	) name12242 (
		_w12695_,
		_w12703_,
		_w12704_
	);
	LUT2 #(
		.INIT('h1)
	) name12243 (
		_w12694_,
		_w12704_,
		_w12705_
	);
	LUT2 #(
		.INIT('h1)
	) name12244 (
		_w12693_,
		_w12705_,
		_w12706_
	);
	LUT2 #(
		.INIT('h1)
	) name12245 (
		_w12692_,
		_w12706_,
		_w12707_
	);
	LUT2 #(
		.INIT('h1)
	) name12246 (
		_w12691_,
		_w12707_,
		_w12708_
	);
	LUT2 #(
		.INIT('h1)
	) name12247 (
		_w12690_,
		_w12708_,
		_w12709_
	);
	LUT2 #(
		.INIT('h1)
	) name12248 (
		_w12689_,
		_w12709_,
		_w12710_
	);
	LUT2 #(
		.INIT('h1)
	) name12249 (
		_w12688_,
		_w12710_,
		_w12711_
	);
	LUT2 #(
		.INIT('h1)
	) name12250 (
		_w12687_,
		_w12711_,
		_w12712_
	);
	LUT2 #(
		.INIT('h1)
	) name12251 (
		_w12686_,
		_w12712_,
		_w12713_
	);
	LUT2 #(
		.INIT('h1)
	) name12252 (
		_w12685_,
		_w12713_,
		_w12714_
	);
	LUT2 #(
		.INIT('h1)
	) name12253 (
		_w12684_,
		_w12714_,
		_w12715_
	);
	LUT2 #(
		.INIT('h1)
	) name12254 (
		_w12683_,
		_w12715_,
		_w12716_
	);
	LUT2 #(
		.INIT('h1)
	) name12255 (
		_w12682_,
		_w12716_,
		_w12717_
	);
	LUT2 #(
		.INIT('h4)
	) name12256 (
		_w12681_,
		_w12717_,
		_w12718_
	);
	LUT2 #(
		.INIT('h2)
	) name12257 (
		_w12681_,
		_w12717_,
		_w12719_
	);
	LUT2 #(
		.INIT('h1)
	) name12258 (
		_w12718_,
		_w12719_,
		_w12720_
	);
	LUT2 #(
		.INIT('h8)
	) name12259 (
		\P1_addr_reg[11]/NET0131 ,
		\P2_addr_reg[11]/NET0131 ,
		_w12721_
	);
	LUT2 #(
		.INIT('h1)
	) name12260 (
		\P1_addr_reg[11]/NET0131 ,
		\P2_addr_reg[11]/NET0131 ,
		_w12722_
	);
	LUT2 #(
		.INIT('h1)
	) name12261 (
		_w12721_,
		_w12722_,
		_w12723_
	);
	LUT2 #(
		.INIT('h1)
	) name12262 (
		_w12679_,
		_w12717_,
		_w12724_
	);
	LUT2 #(
		.INIT('h1)
	) name12263 (
		_w12680_,
		_w12724_,
		_w12725_
	);
	LUT2 #(
		.INIT('h4)
	) name12264 (
		_w12723_,
		_w12725_,
		_w12726_
	);
	LUT2 #(
		.INIT('h2)
	) name12265 (
		_w12723_,
		_w12725_,
		_w12727_
	);
	LUT2 #(
		.INIT('h1)
	) name12266 (
		_w12726_,
		_w12727_,
		_w12728_
	);
	LUT2 #(
		.INIT('h8)
	) name12267 (
		\P1_addr_reg[12]/NET0131 ,
		\P2_addr_reg[12]/NET0131 ,
		_w12729_
	);
	LUT2 #(
		.INIT('h1)
	) name12268 (
		\P1_addr_reg[12]/NET0131 ,
		\P2_addr_reg[12]/NET0131 ,
		_w12730_
	);
	LUT2 #(
		.INIT('h1)
	) name12269 (
		_w12729_,
		_w12730_,
		_w12731_
	);
	LUT2 #(
		.INIT('h1)
	) name12270 (
		_w12721_,
		_w12725_,
		_w12732_
	);
	LUT2 #(
		.INIT('h1)
	) name12271 (
		_w12722_,
		_w12732_,
		_w12733_
	);
	LUT2 #(
		.INIT('h4)
	) name12272 (
		_w12731_,
		_w12733_,
		_w12734_
	);
	LUT2 #(
		.INIT('h2)
	) name12273 (
		_w12731_,
		_w12733_,
		_w12735_
	);
	LUT2 #(
		.INIT('h1)
	) name12274 (
		_w12734_,
		_w12735_,
		_w12736_
	);
	LUT2 #(
		.INIT('h8)
	) name12275 (
		\P1_addr_reg[13]/NET0131 ,
		\P2_addr_reg[13]/NET0131 ,
		_w12737_
	);
	LUT2 #(
		.INIT('h1)
	) name12276 (
		\P1_addr_reg[13]/NET0131 ,
		\P2_addr_reg[13]/NET0131 ,
		_w12738_
	);
	LUT2 #(
		.INIT('h1)
	) name12277 (
		_w12737_,
		_w12738_,
		_w12739_
	);
	LUT2 #(
		.INIT('h1)
	) name12278 (
		_w12729_,
		_w12733_,
		_w12740_
	);
	LUT2 #(
		.INIT('h1)
	) name12279 (
		_w12730_,
		_w12740_,
		_w12741_
	);
	LUT2 #(
		.INIT('h4)
	) name12280 (
		_w12739_,
		_w12741_,
		_w12742_
	);
	LUT2 #(
		.INIT('h2)
	) name12281 (
		_w12739_,
		_w12741_,
		_w12743_
	);
	LUT2 #(
		.INIT('h1)
	) name12282 (
		_w12742_,
		_w12743_,
		_w12744_
	);
	LUT2 #(
		.INIT('h8)
	) name12283 (
		\P1_addr_reg[14]/NET0131 ,
		\P2_addr_reg[14]/NET0131 ,
		_w12745_
	);
	LUT2 #(
		.INIT('h1)
	) name12284 (
		\P1_addr_reg[14]/NET0131 ,
		\P2_addr_reg[14]/NET0131 ,
		_w12746_
	);
	LUT2 #(
		.INIT('h1)
	) name12285 (
		_w12745_,
		_w12746_,
		_w12747_
	);
	LUT2 #(
		.INIT('h1)
	) name12286 (
		_w12737_,
		_w12741_,
		_w12748_
	);
	LUT2 #(
		.INIT('h1)
	) name12287 (
		_w12738_,
		_w12748_,
		_w12749_
	);
	LUT2 #(
		.INIT('h4)
	) name12288 (
		_w12747_,
		_w12749_,
		_w12750_
	);
	LUT2 #(
		.INIT('h2)
	) name12289 (
		_w12747_,
		_w12749_,
		_w12751_
	);
	LUT2 #(
		.INIT('h1)
	) name12290 (
		_w12750_,
		_w12751_,
		_w12752_
	);
	LUT2 #(
		.INIT('h8)
	) name12291 (
		\P1_addr_reg[15]/NET0131 ,
		\P2_addr_reg[15]/NET0131 ,
		_w12753_
	);
	LUT2 #(
		.INIT('h1)
	) name12292 (
		\P1_addr_reg[15]/NET0131 ,
		\P2_addr_reg[15]/NET0131 ,
		_w12754_
	);
	LUT2 #(
		.INIT('h1)
	) name12293 (
		_w12753_,
		_w12754_,
		_w12755_
	);
	LUT2 #(
		.INIT('h1)
	) name12294 (
		_w12745_,
		_w12749_,
		_w12756_
	);
	LUT2 #(
		.INIT('h1)
	) name12295 (
		_w12746_,
		_w12756_,
		_w12757_
	);
	LUT2 #(
		.INIT('h4)
	) name12296 (
		_w12755_,
		_w12757_,
		_w12758_
	);
	LUT2 #(
		.INIT('h2)
	) name12297 (
		_w12755_,
		_w12757_,
		_w12759_
	);
	LUT2 #(
		.INIT('h1)
	) name12298 (
		_w12758_,
		_w12759_,
		_w12760_
	);
	LUT2 #(
		.INIT('h8)
	) name12299 (
		\P1_addr_reg[16]/NET0131 ,
		\P2_addr_reg[16]/NET0131 ,
		_w12761_
	);
	LUT2 #(
		.INIT('h1)
	) name12300 (
		\P1_addr_reg[16]/NET0131 ,
		\P2_addr_reg[16]/NET0131 ,
		_w12762_
	);
	LUT2 #(
		.INIT('h1)
	) name12301 (
		_w12761_,
		_w12762_,
		_w12763_
	);
	LUT2 #(
		.INIT('h1)
	) name12302 (
		_w12753_,
		_w12757_,
		_w12764_
	);
	LUT2 #(
		.INIT('h1)
	) name12303 (
		_w12754_,
		_w12764_,
		_w12765_
	);
	LUT2 #(
		.INIT('h4)
	) name12304 (
		_w12763_,
		_w12765_,
		_w12766_
	);
	LUT2 #(
		.INIT('h2)
	) name12305 (
		_w12763_,
		_w12765_,
		_w12767_
	);
	LUT2 #(
		.INIT('h1)
	) name12306 (
		_w12766_,
		_w12767_,
		_w12768_
	);
	LUT2 #(
		.INIT('h8)
	) name12307 (
		\P1_addr_reg[17]/NET0131 ,
		\P2_addr_reg[17]/NET0131 ,
		_w12769_
	);
	LUT2 #(
		.INIT('h1)
	) name12308 (
		\P1_addr_reg[17]/NET0131 ,
		\P2_addr_reg[17]/NET0131 ,
		_w12770_
	);
	LUT2 #(
		.INIT('h1)
	) name12309 (
		_w12769_,
		_w12770_,
		_w12771_
	);
	LUT2 #(
		.INIT('h1)
	) name12310 (
		_w12761_,
		_w12765_,
		_w12772_
	);
	LUT2 #(
		.INIT('h1)
	) name12311 (
		_w12762_,
		_w12772_,
		_w12773_
	);
	LUT2 #(
		.INIT('h4)
	) name12312 (
		_w12771_,
		_w12773_,
		_w12774_
	);
	LUT2 #(
		.INIT('h2)
	) name12313 (
		_w12771_,
		_w12773_,
		_w12775_
	);
	LUT2 #(
		.INIT('h1)
	) name12314 (
		_w12774_,
		_w12775_,
		_w12776_
	);
	LUT2 #(
		.INIT('h8)
	) name12315 (
		\P1_addr_reg[18]/NET0131 ,
		\P2_addr_reg[18]/NET0131 ,
		_w12777_
	);
	LUT2 #(
		.INIT('h1)
	) name12316 (
		\P1_addr_reg[18]/NET0131 ,
		\P2_addr_reg[18]/NET0131 ,
		_w12778_
	);
	LUT2 #(
		.INIT('h1)
	) name12317 (
		_w12777_,
		_w12778_,
		_w12779_
	);
	LUT2 #(
		.INIT('h1)
	) name12318 (
		_w12769_,
		_w12773_,
		_w12780_
	);
	LUT2 #(
		.INIT('h1)
	) name12319 (
		_w12770_,
		_w12780_,
		_w12781_
	);
	LUT2 #(
		.INIT('h4)
	) name12320 (
		_w12779_,
		_w12781_,
		_w12782_
	);
	LUT2 #(
		.INIT('h2)
	) name12321 (
		_w12779_,
		_w12781_,
		_w12783_
	);
	LUT2 #(
		.INIT('h1)
	) name12322 (
		_w12782_,
		_w12783_,
		_w12784_
	);
	LUT2 #(
		.INIT('h1)
	) name12323 (
		_w539_,
		_w541_,
		_w12785_
	);
	LUT2 #(
		.INIT('h1)
	) name12324 (
		_w12777_,
		_w12781_,
		_w12786_
	);
	LUT2 #(
		.INIT('h1)
	) name12325 (
		_w12778_,
		_w12786_,
		_w12787_
	);
	LUT2 #(
		.INIT('h2)
	) name12326 (
		_w12785_,
		_w12787_,
		_w12788_
	);
	LUT2 #(
		.INIT('h4)
	) name12327 (
		_w12785_,
		_w12787_,
		_w12789_
	);
	LUT2 #(
		.INIT('h1)
	) name12328 (
		_w12788_,
		_w12789_,
		_w12790_
	);
	LUT2 #(
		.INIT('h1)
	) name12329 (
		_w12698_,
		_w12699_,
		_w12791_
	);
	LUT2 #(
		.INIT('h2)
	) name12330 (
		_w12676_,
		_w12791_,
		_w12792_
	);
	LUT2 #(
		.INIT('h4)
	) name12331 (
		_w12676_,
		_w12791_,
		_w12793_
	);
	LUT2 #(
		.INIT('h1)
	) name12332 (
		_w12792_,
		_w12793_,
		_w12794_
	);
	LUT2 #(
		.INIT('h1)
	) name12333 (
		_w12696_,
		_w12697_,
		_w12795_
	);
	LUT2 #(
		.INIT('h2)
	) name12334 (
		_w12701_,
		_w12795_,
		_w12796_
	);
	LUT2 #(
		.INIT('h4)
	) name12335 (
		_w12701_,
		_w12795_,
		_w12797_
	);
	LUT2 #(
		.INIT('h1)
	) name12336 (
		_w12796_,
		_w12797_,
		_w12798_
	);
	LUT2 #(
		.INIT('h1)
	) name12337 (
		_w12694_,
		_w12695_,
		_w12799_
	);
	LUT2 #(
		.INIT('h2)
	) name12338 (
		_w12703_,
		_w12799_,
		_w12800_
	);
	LUT2 #(
		.INIT('h4)
	) name12339 (
		_w12703_,
		_w12799_,
		_w12801_
	);
	LUT2 #(
		.INIT('h1)
	) name12340 (
		_w12800_,
		_w12801_,
		_w12802_
	);
	LUT2 #(
		.INIT('h1)
	) name12341 (
		_w12692_,
		_w12693_,
		_w12803_
	);
	LUT2 #(
		.INIT('h2)
	) name12342 (
		_w12705_,
		_w12803_,
		_w12804_
	);
	LUT2 #(
		.INIT('h4)
	) name12343 (
		_w12705_,
		_w12803_,
		_w12805_
	);
	LUT2 #(
		.INIT('h1)
	) name12344 (
		_w12804_,
		_w12805_,
		_w12806_
	);
	LUT2 #(
		.INIT('h1)
	) name12345 (
		_w12690_,
		_w12691_,
		_w12807_
	);
	LUT2 #(
		.INIT('h2)
	) name12346 (
		_w12707_,
		_w12807_,
		_w12808_
	);
	LUT2 #(
		.INIT('h4)
	) name12347 (
		_w12707_,
		_w12807_,
		_w12809_
	);
	LUT2 #(
		.INIT('h1)
	) name12348 (
		_w12808_,
		_w12809_,
		_w12810_
	);
	LUT2 #(
		.INIT('h1)
	) name12349 (
		_w12688_,
		_w12689_,
		_w12811_
	);
	LUT2 #(
		.INIT('h2)
	) name12350 (
		_w12709_,
		_w12811_,
		_w12812_
	);
	LUT2 #(
		.INIT('h4)
	) name12351 (
		_w12709_,
		_w12811_,
		_w12813_
	);
	LUT2 #(
		.INIT('h1)
	) name12352 (
		_w12812_,
		_w12813_,
		_w12814_
	);
	LUT2 #(
		.INIT('h1)
	) name12353 (
		_w12686_,
		_w12687_,
		_w12815_
	);
	LUT2 #(
		.INIT('h2)
	) name12354 (
		_w12711_,
		_w12815_,
		_w12816_
	);
	LUT2 #(
		.INIT('h4)
	) name12355 (
		_w12711_,
		_w12815_,
		_w12817_
	);
	LUT2 #(
		.INIT('h1)
	) name12356 (
		_w12816_,
		_w12817_,
		_w12818_
	);
	LUT2 #(
		.INIT('h1)
	) name12357 (
		_w12684_,
		_w12685_,
		_w12819_
	);
	LUT2 #(
		.INIT('h2)
	) name12358 (
		_w12713_,
		_w12819_,
		_w12820_
	);
	LUT2 #(
		.INIT('h4)
	) name12359 (
		_w12713_,
		_w12819_,
		_w12821_
	);
	LUT2 #(
		.INIT('h1)
	) name12360 (
		_w12820_,
		_w12821_,
		_w12822_
	);
	LUT2 #(
		.INIT('h1)
	) name12361 (
		_w12682_,
		_w12683_,
		_w12823_
	);
	LUT2 #(
		.INIT('h2)
	) name12362 (
		_w12715_,
		_w12823_,
		_w12824_
	);
	LUT2 #(
		.INIT('h4)
	) name12363 (
		_w12715_,
		_w12823_,
		_w12825_
	);
	LUT2 #(
		.INIT('h1)
	) name12364 (
		_w12824_,
		_w12825_,
		_w12826_
	);
	LUT2 #(
		.INIT('h1)
	) name12365 (
		\P1_wr_reg/NET0131 ,
		\P2_wr_reg/NET0131 ,
		_w12827_
	);
	LUT2 #(
		.INIT('h8)
	) name12366 (
		\P1_wr_reg/NET0131 ,
		\P2_wr_reg/NET0131 ,
		_w12828_
	);
	LUT2 #(
		.INIT('h1)
	) name12367 (
		_w12827_,
		_w12828_,
		_w12829_
	);
	assign \P1_state_reg[0]/NET0131_syn_2  = \P1_state_reg[0]/NET0131 ;
	assign \_al_n0  = 1'b0;
	assign \_al_n1  = 1'b0;
	assign \g73521/_0_  = _w1956_ ;
	assign \g73537/_0_  = _w3434_ ;
	assign \g73538/_0_  = _w3730_ ;
	assign \g73539/_0_  = _w3755_ ;
	assign \g73540/_0_  = _w3786_ ;
	assign \g73570/_0_  = _w3979_ ;
	assign \g73571/_0_  = _w4117_ ;
	assign \g73572/_0_  = _w4327_ ;
	assign \g73573/_0_  = _w4350_ ;
	assign \g73574/_0_  = _w4368_ ;
	assign \g73575/_0_  = _w4393_ ;
	assign \g73576/_0_  = _w4503_ ;
	assign \g73577/_0_  = _w4529_ ;
	assign \g73578/_0_  = _w4558_ ;
	assign \g73579/_0_  = _w4582_ ;
	assign \g73609/_0_  = _w4643_ ;
	assign \g73610/_0_  = _w4702_ ;
	assign \g73611/_0_  = _w4797_ ;
	assign \g73613/_0_  = _w4895_ ;
	assign \g73614/_0_  = _w4923_ ;
	assign \g73615/_0_  = _w4949_ ;
	assign \g73617/_0_  = _w4974_ ;
	assign \g73618/_0_  = _w5021_ ;
	assign \g73619/_0_  = _w5048_ ;
	assign \g73620/_0_  = _w5078_ ;
	assign \g73621/_0_  = _w5096_ ;
	assign \g73622/_0_  = _w5114_ ;
	assign \g73623/_0_  = _w5132_ ;
	assign \g73624/_0_  = _w5158_ ;
	assign \g73625/_0_  = _w5217_ ;
	assign \g73626/_0_  = _w5246_ ;
	assign \g73627/_0_  = _w5274_ ;
	assign \g73628/_0_  = _w5294_ ;
	assign \g73629/_0_  = _w5321_ ;
	assign \g73630/_0_  = _w5347_ ;
	assign \g73631/_0_  = _w5373_ ;
	assign \g73632/_0_  = _w5399_ ;
	assign \g73633/_0_  = _w5425_ ;
	assign \g73692/_0_  = _w5475_ ;
	assign \g73693/_0_  = _w5550_ ;
	assign \g73694/_0_  = _w5600_ ;
	assign \g73696/_0_  = _w5644_ ;
	assign \g73697/_0_  = _w5688_ ;
	assign \g73703/_0_  = _w5716_ ;
	assign \g73704/_0_  = _w5744_ ;
	assign \g73709/_0_  = _w5793_ ;
	assign \g73710/_0_  = _w5818_ ;
	assign \g73711/_0_  = _w5841_ ;
	assign \g73712/_0_  = _w5859_ ;
	assign \g73713/_0_  = _w5866_ ;
	assign \g73714/_0_  = _w5894_ ;
	assign \g73715/_0_  = _w5960_ ;
	assign \g73716/_0_  = _w5966_ ;
	assign \g73717/_0_  = _w5992_ ;
	assign \g73718/_0_  = _w6014_ ;
	assign \g73719/_0_  = _w6066_ ;
	assign \g73720/_0_  = _w6088_ ;
	assign \g73774/_0_  = _w6131_ ;
	assign \g73775/_0_  = _w6173_ ;
	assign \g73776/_0_  = _w6216_ ;
	assign \g73777/_0_  = _w6259_ ;
	assign \g73806/_0_  = _w6285_ ;
	assign \g73807/_0_  = _w6325_ ;
	assign \g73808/_0_  = _w6367_ ;
	assign \g73809/_0_  = _w6372_ ;
	assign \g73810/_0_  = _w6395_ ;
	assign \g73811/_0_  = _w6424_ ;
	assign \g73812/_0_  = _w6453_ ;
	assign \g73813/_0_  = _w6483_ ;
	assign \g73814/_0_  = _w6526_ ;
	assign \g73815/_0_  = _w6553_ ;
	assign \g73816/_0_  = _w6583_ ;
	assign \g73817/_0_  = _w6609_ ;
	assign \g73818/_0_  = _w6636_ ;
	assign \g73819/_0_  = _w6654_ ;
	assign \g73820/_0_  = _w6672_ ;
	assign \g73821/_0_  = _w6700_ ;
	assign \g73822/_0_  = _w6728_ ;
	assign \g73823/_0_  = _w6770_ ;
	assign \g73824/_0_  = _w6790_ ;
	assign \g73825/_0_  = _w6816_ ;
	assign \g73826/_0_  = _w6842_ ;
	assign \g73827/_0_  = _w6863_ ;
	assign \g73828/_0_  = _w6885_ ;
	assign \g73829/_0_  = _w6890_ ;
	assign \g73830/_0_  = _w6916_ ;
	assign \g73831/_0_  = _w6942_ ;
	assign \g73832/_0_  = _w6952_ ;
	assign \g73833/_0_  = _w6992_ ;
	assign \g73834/_0_  = _w7018_ ;
	assign \g73835/_0_  = _w7044_ ;
	assign \g73836/_0_  = _w7070_ ;
	assign \g73908/_0_  = _w7111_ ;
	assign \g73909/_0_  = _w7153_ ;
	assign \g73911/_0_  = _w7195_ ;
	assign \g73912/_0_  = _w7237_ ;
	assign \g73915/_0_  = _w7280_ ;
	assign \g73916/_0_  = _w7324_ ;
	assign \g73946/_0_  = _w7352_ ;
	assign \g73950/_0_  = _w7380_ ;
	assign \g73957/_0_  = _w7408_ ;
	assign \g73958/_0_  = _w7462_ ;
	assign \g73959/_0_  = _w7488_ ;
	assign \g73960/_0_  = _w7503_ ;
	assign \g73961/_0_  = _w7514_ ;
	assign \g73962/_0_  = _w7543_ ;
	assign \g73963/_0_  = _w7552_ ;
	assign \g73964/_0_  = _w7581_ ;
	assign \g73965/_0_  = _w7607_ ;
	assign \g73966/_0_  = _w7635_ ;
	assign \g73968/_0_  = _w7664_ ;
	assign \g73969/_0_  = _w7690_ ;
	assign \g73970/_0_  = _w7693_ ;
	assign \g73971/_0_  = _w7707_ ;
	assign \g73972/_0_  = _w7735_ ;
	assign \g73973/_0_  = _w7764_ ;
	assign \g73974/_0_  = _w7775_ ;
	assign \g73975/_0_  = _w7790_ ;
	assign \g73976/_0_  = _w7816_ ;
	assign \g73977/_0_  = _w7832_ ;
	assign \g73978/_0_  = _w7858_ ;
	assign \g73979/_0_  = _w7884_ ;
	assign \g73980/_0_  = _w7887_ ;
	assign \g73981/_0_  = _w7913_ ;
	assign \g73982/_0_  = _w7924_ ;
	assign \g73983/_0_  = _w7950_ ;
	assign \g73984/_0_  = _w7972_ ;
	assign \g73985/_0_  = _w7996_ ;
	assign \g74044/_0_  = _w8036_ ;
	assign \g74045/_0_  = _w8080_ ;
	assign \g74046/_0_  = _w8120_ ;
	assign \g74047/_0_  = _w8160_ ;
	assign \g74048/_0_  = _w8201_ ;
	assign \g74049/_0_  = _w8242_ ;
	assign \g74051/_0_  = _w8282_ ;
	assign \g74052/_0_  = _w8324_ ;
	assign \g74099/_0_  = _w8369_ ;
	assign \g74100/_0_  = _w8393_ ;
	assign \g74101/_0_  = _w8420_ ;
	assign \g74102/_0_  = _w8449_ ;
	assign \g74103/_0_  = _w8478_ ;
	assign \g74104/_0_  = _w8500_ ;
	assign \g74105/_0_  = _w8527_ ;
	assign \g74106/_0_  = _w8550_ ;
	assign \g74107/_0_  = _w8568_ ;
	assign \g74108/_0_  = _w8594_ ;
	assign \g74109/_0_  = _w8612_ ;
	assign \g74110/_0_  = _w8640_ ;
	assign \g74111/_0_  = _w8664_ ;
	assign \g74112/_0_  = _w8692_ ;
	assign \g74113/_0_  = _w8713_ ;
	assign \g74114/_0_  = _w8741_ ;
	assign \g74115/_0_  = _w8767_ ;
	assign \g74116/_0_  = _w8790_ ;
	assign \g74117/_0_  = _w8816_ ;
	assign \g74118/_0_  = _w8842_ ;
	assign \g74119/_0_  = _w8868_ ;
	assign \g74120/_0_  = _w8894_ ;
	assign \g74121/_0_  = _w8912_ ;
	assign \g74122/_0_  = _w8934_ ;
	assign \g74199/_0_  = _w8976_ ;
	assign \g74200/_0_  = _w9015_ ;
	assign \g74201/_0_  = _w9057_ ;
	assign \g74202/_0_  = _w9103_ ;
	assign \g74279/_0_  = _w9130_ ;
	assign \g74280/_0_  = _w9156_ ;
	assign \g74284/_0_  = _w9183_ ;
	assign \g74285/_0_  = _w9209_ ;
	assign \g74287/_0_  = _w9238_ ;
	assign \g74288/_0_  = _w9264_ ;
	assign \g74289/_0_  = _w9290_ ;
	assign \g74290/_0_  = _w9317_ ;
	assign \g74291/_0_  = _w9343_ ;
	assign \g74292/_0_  = _w9356_ ;
	assign \g74293/_0_  = _w9381_ ;
	assign \g74294/_0_  = _w9390_ ;
	assign \g74295/_0_  = _w9419_ ;
	assign \g74296/_0_  = _w9448_ ;
	assign \g74298/_0_  = _w9476_ ;
	assign \g74299/_0_  = _w9498_ ;
	assign \g74300/_0_  = _w9524_ ;
	assign \g74301/_0_  = _w9552_ ;
	assign \g74302/_0_  = _w9574_ ;
	assign \g74382/_0_  = _w9614_ ;
	assign \g74383/_0_  = _w9655_ ;
	assign \g74384/_0_  = _w9695_ ;
	assign \g74385/_0_  = _w9739_ ;
	assign \g74386/_0_  = _w9780_ ;
	assign \g74387/_0_  = _w9820_ ;
	assign \g74456/_0_  = _w9844_ ;
	assign \g74457/_0_  = _w9854_ ;
	assign \g74458/_0_  = _w9875_ ;
	assign \g74459/_0_  = _w9901_ ;
	assign \g74460/_0_  = _w9910_ ;
	assign \g74461/_0_  = _w9938_ ;
	assign \g74462/_0_  = _w9964_ ;
	assign \g74463/_0_  = _w9986_ ;
	assign \g74464/_0_  = _w10014_ ;
	assign \g74465/_0_  = _w10024_ ;
	assign \g74466/_0_  = _w10048_ ;
	assign \g74467/_0_  = _w10076_ ;
	assign \g74468/_0_  = _w10104_ ;
	assign \g74469/_0_  = _w10128_ ;
	assign \g74470/_0_  = _w10146_ ;
	assign \g74471/_0_  = _w10172_ ;
	assign \g74661/_0_  = _w10194_ ;
	assign \g74662/_0_  = _w10218_ ;
	assign \g74663/_0_  = _w10238_ ;
	assign \g74664/_0_  = _w10260_ ;
	assign \g74665/_0_  = _w10278_ ;
	assign \g74666/_0_  = _w10296_ ;
	assign \g74667/_0_  = _w10320_ ;
	assign \g74668/_0_  = _w10349_ ;
	assign \g74669/_0_  = _w10373_ ;
	assign \g74670/_0_  = _w10394_ ;
	assign \g74671/_0_  = _w10423_ ;
	assign \g74672/_0_  = _w10451_ ;
	assign \g74673/_0_  = _w10471_ ;
	assign \g74674/_0_  = _w10499_ ;
	assign \g74899/_0_  = _w10525_ ;
	assign \g74900/_0_  = _w10551_ ;
	assign \g74901/_0_  = _w10577_ ;
	assign \g74902/_0_  = _w10603_ ;
	assign \g75002/_0_  = _w10642_ ;
	assign \g75005/_0_  = _w10681_ ;
	assign \g75191/_0_  = _w10708_ ;
	assign \g75192/_0_  = _w10734_ ;
	assign \g75193/_0_  = _w10763_ ;
	assign \g75194/_0_  = _w10789_ ;
	assign \g75195/_0_  = _w10815_ ;
	assign \g75392/_0_  = _w10853_ ;
	assign \g75399/_0_  = _w10891_ ;
	assign \g75606/_0_  = _w10915_ ;
	assign \g75607/_0_  = _w10937_ ;
	assign \g75608/_0_  = _w10965_ ;
	assign \g75609/_0_  = _w10989_ ;
	assign \g75610/_0_  = _w11011_ ;
	assign \g76007/_0_  = _w11041_ ;
	assign \g76008/_0_  = _w11065_ ;
	assign \g76685/_0_  = _w11089_ ;
	assign \g76696/_0_  = _w11114_ ;
	assign \g77574/_0_  = _w11130_ ;
	assign \g77575/_0_  = _w11150_ ;
	assign \g77576/_0_  = _w11161_ ;
	assign \g77577/_0_  = _w11181_ ;
	assign \g77578/_0_  = _w11187_ ;
	assign \g77579/_0_  = _w11207_ ;
	assign \g82699/_3_  = _w11210_ ;
	assign \g82700/_3_  = _w11213_ ;
	assign \g82701/_3_  = _w11216_ ;
	assign \g82702/_3_  = _w11219_ ;
	assign \g82703/_3_  = _w11222_ ;
	assign \g82704/_3_  = _w11225_ ;
	assign \g83319/_0_  = _w11228_ ;
	assign \g83320/_0_  = _w11231_ ;
	assign \g83321/_0_  = _w11234_ ;
	assign \g83322/_0_  = _w11237_ ;
	assign \g83323/_3_  = _w11240_ ;
	assign \g83324/_0_  = _w11243_ ;
	assign \g83325/_0_  = _w11246_ ;
	assign \g83326/_0_  = _w11249_ ;
	assign \g83327/_0_  = _w11252_ ;
	assign \g83328/_0_  = _w11255_ ;
	assign \g83329/_0_  = _w11258_ ;
	assign \g83330/_0_  = _w11261_ ;
	assign \g83331/_0_  = _w11264_ ;
	assign \g83332/_0_  = _w11267_ ;
	assign \g83333/_0_  = _w11269_ ;
	assign \g83334/_0_  = _w11272_ ;
	assign \g83335/_0_  = _w11275_ ;
	assign \g83336/_3_  = _w11278_ ;
	assign \g83337/_0_  = _w11281_ ;
	assign \g83338/_0_  = _w11284_ ;
	assign \g83339/_0_  = _w11287_ ;
	assign \g83340/_0_  = _w11290_ ;
	assign \g83341/_0_  = _w11293_ ;
	assign \g83342/_0_  = _w11296_ ;
	assign \g83343/_0_  = _w11299_ ;
	assign \g83344/_0_  = _w11302_ ;
	assign \g83345/_0_  = _w11305_ ;
	assign \g83347/_3_  = _w11308_ ;
	assign \g83348/_3_  = _w11311_ ;
	assign \g83349/_3_  = _w11314_ ;
	assign \g83350/_3_  = _w11317_ ;
	assign \g83351/_3_  = _w11320_ ;
	assign \g83352/_3_  = _w11323_ ;
	assign \g83353/_3_  = _w11326_ ;
	assign \g83354/_3_  = _w11329_ ;
	assign \g83355/_3_  = _w11332_ ;
	assign \g83356/_3_  = _w11335_ ;
	assign \g83357/_0_  = _w11338_ ;
	assign \g83358/_3_  = _w11341_ ;
	assign \g83359/_3_  = _w11344_ ;
	assign \g83360/_3_  = _w11346_ ;
	assign \g83361/_3_  = _w11349_ ;
	assign \g83362/_3_  = _w11352_ ;
	assign \g83363/_3_  = _w11355_ ;
	assign \g83364/_3_  = _w11358_ ;
	assign \g83365/_0_  = _w11361_ ;
	assign \g83366/_3_  = _w11364_ ;
	assign \g83367/_0_  = _w11370_ ;
	assign \g83368/_3_  = _w11373_ ;
	assign \g83369/_3_  = _w11376_ ;
	assign \g83370/_0_  = _w11379_ ;
	assign \g83371/_3_  = _w11382_ ;
	assign \g83372/_3_  = _w11385_ ;
	assign \g83373/_3_  = _w11388_ ;
	assign \g83374/_3_  = _w11391_ ;
	assign \g83376/_0_  = _w11398_ ;
	assign \g83778/_0_  = _w1668_ ;
	assign \g83784/_0_  = _w2601_ ;
	assign \g84388/_0_  = _w11473_ ;
	assign \g84389/_0_  = _w11507_ ;
	assign \g84391/_0_  = _w11525_ ;
	assign \g84395/_0_  = _w11547_ ;
	assign \g84397/_0_  = _w11567_ ;
	assign \g84398/_0_  = _w11617_ ;
	assign \g84399/_0_  = _w11639_ ;
	assign \g84400/_0_  = _w11656_ ;
	assign \g84401/_0_  = _w11684_ ;
	assign \g84402/_0_  = _w11702_ ;
	assign \g84403/_0_  = _w11728_ ;
	assign \g84405/_0_  = _w11823_ ;
	assign \g84406/_0_  = _w11853_ ;
	assign \g84407/_0_  = _w11895_ ;
	assign \g84408/_0_  = _w11925_ ;
	assign \g84409/_0_  = _w11955_ ;
	assign \g84410/_0_  = _w11986_ ;
	assign \g84411/_0_  = _w12016_ ;
	assign \g84412/_0_  = _w12046_ ;
	assign \g84413/_0_  = _w12076_ ;
	assign \g84414/_0_  = _w12106_ ;
	assign \g84415/_0_  = _w12136_ ;
	assign \g84416/_0_  = _w12157_ ;
	assign \g84417/_0_  = _w12187_ ;
	assign \g84418/_0_  = _w12208_ ;
	assign \g84419/_0_  = _w12228_ ;
	assign \g84420/_0_  = _w12249_ ;
	assign \g84421/_0_  = _w12269_ ;
	assign \g84422/_0_  = _w12287_ ;
	assign \g84423/_0_  = _w12305_ ;
	assign \g84424/_0_  = _w12323_ ;
	assign \g84425/_0_  = _w12343_ ;
	assign \g84426/_0_  = _w12361_ ;
	assign \g84427/_0_  = _w12382_ ;
	assign \g84429/_0_  = _w12402_ ;
	assign \g84430/_0_  = _w12422_ ;
	assign \g84442/_0_  = _w12453_ ;
	assign \g84443/_0_  = _w12483_ ;
	assign \g84444/_0_  = _w12513_ ;
	assign \g84445/_0_  = _w12543_ ;
	assign \g84908/_0_  = _w12545_ ;
	assign \g84961/_0_  = _w12547_ ;
	assign \g84984/u3_syn_4  = _w5812_ ;
	assign \g84985/u3_syn_4  = _w5287_ ;
	assign \g85802/_0_  = _w3460_ ;
	assign \g86055/_1_  = _w2035_ ;
	assign \g86073/_0_  = _w3465_ ;
	assign \g86298/u3_syn_4  = _w12548_ ;
	assign \g86300/u3_syn_4  = _w12549_ ;
	assign \g87397/_0_  = _w12552_ ;
	assign \g87409/_0_  = _w12555_ ;
	assign \g87480/_0_  = _w887_ ;
	assign \g87494/_0_  = _w831_ ;
	assign \g87544/_0_  = _w750_ ;
	assign \g87555/_0_  = _w2251_ ;
	assign \g87567/_0_  = _w3372_ ;
	assign \g87576/_0_  = _w3402_ ;
	assign \g87894/_0_  = _w1475_ ;
	assign \g87905/_0_  = _w3021_ ;
	assign \g87914/_0_  = _w978_ ;
	assign \g87955/_1_  = _w1062_ ;
	assign \g88030/_0_  = _w1524_ ;
	assign \g88039/_0_  = _w1244_ ;
	assign \g88054/_0_  = _w1267_ ;
	assign \g88079/_0_  = _w2828_ ;
	assign \g88094/_0_  = _w945_ ;
	assign \g88111/_0_  = _w1498_ ;
	assign \g88122/_0_  = _w1664_ ;
	assign \g88129/_0_  = _w1427_ ;
	assign \g88162/_0_  = _w1174_ ;
	assign \g88185/_0_  = _w2715_ ;
	assign \g88196/_0_  = _w2880_ ;
	assign \g88204/_0_  = _w1118_ ;
	assign \g88220/_0_  = _w1218_ ;
	assign \g88226/_0_  = _w2597_ ;
	assign \g88243/_0_  = _w1548_ ;
	assign \g88252/_0_  = _w2531_ ;
	assign \g88261/_0_  = _w2506_ ;
	assign \g88269/_0_  = _w2742_ ;
	assign \g88288/_0_  = _w2379_ ;
	assign \g88299/_0_  = _w2442_ ;
	assign \g88310/_0_  = _w2962_ ;
	assign \g88321/_0_  = _w3130_ ;
	assign \g88328/_0_  = _w3112_ ;
	assign \g88335/_0_  = _w3088_ ;
	assign \g88356/_0_  = _w2454_ ;
	assign \g88366/_0_  = _w2688_ ;
	assign \g88372/_0_  = _w2552_ ;
	assign \g88380/_0_  = _w2311_ ;
	assign \g88395_dup/_0_  = _w2574_ ;
	assign \g88403/_0_  = _w2991_ ;
	assign \g88414/_0_  = _w2368_ ;
	assign \g88425/_0_  = _w1146_ ;
	assign \g88443/_0_  = _w1374_ ;
	assign \g88453/_0_  = _w1318_ ;
	assign \g88471/_0_  = _w1336_ ;
	assign \g88524/_0_  = _w1356_ ;
	assign \g88546/_0_  = _w1006_ ;
	assign \g88556/_0_  = _w2765_ ;
	assign \g88563/_0_  = _w1207_ ;
	assign \g89966/_1_  = _w3435_ ;
	assign \g89999/_1_  = _w1983_ ;
	assign \g95209/_0_  = _w12567_ ;
	assign \g95269/_0_  = _w2642_ ;
	assign \g95319/_0_  = _w12594_ ;
	assign \g95354/_0_  = _w2804_ ;
	assign \g95786/_0_  = _w2616_ ;
	assign \g95909/_0_  = _w1595_ ;
	assign \g95914/_0_  = _w1572_ ;
	assign \g95918/_0_  = _w1617_ ;
	assign \g95984/_0_  = _w2870_ ;
	assign \g96009/_0_  = _w3065_ ;
	assign \g96124/_0_  = _w1094_ ;
	assign \g96218/_0_  = _w1452_ ;
	assign \g96286/_0_  = _w1641_ ;
	assign \g96335/_0_  = _w2480_ ;
	assign \g96465/_0_  = _w2039_ ;
	assign \g96694/_0_  = _w12620_ ;
	assign \g96713/_0_  = _w1403_ ;
	assign \g96830/_0_  = _w12644_ ;
	assign \g96875/_0_  = _w12672_ ;
	assign rd_pad = _w12675_ ;
	assign \so[0]_pad  = _w12678_ ;
	assign \so[10]_pad  = _w12720_ ;
	assign \so[11]_pad  = _w12728_ ;
	assign \so[12]_pad  = _w12736_ ;
	assign \so[13]_pad  = _w12744_ ;
	assign \so[14]_pad  = _w12752_ ;
	assign \so[15]_pad  = _w12760_ ;
	assign \so[16]_pad  = _w12768_ ;
	assign \so[17]_pad  = _w12776_ ;
	assign \so[18]_pad  = _w12784_ ;
	assign \so[19]_pad  = _w12790_ ;
	assign \so[1]_pad  = _w12794_ ;
	assign \so[2]_pad  = _w12798_ ;
	assign \so[3]_pad  = _w12802_ ;
	assign \so[4]_pad  = _w12806_ ;
	assign \so[5]_pad  = _w12810_ ;
	assign \so[6]_pad  = _w12814_ ;
	assign \so[7]_pad  = _w12818_ ;
	assign \so[8]_pad  = _w12822_ ;
	assign \so[9]_pad  = _w12826_ ;
	assign wr_pad = _w12829_ ;
endmodule;