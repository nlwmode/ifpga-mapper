module top (\G0_pad , \G10_reg/NET0131 , \G11_reg/NET0131 , \G12_reg/NET0131 , \G13_reg/NET0131 , \G147_pad , \G148_pad , \G14_reg/NET0131 , \G15_reg/NET0131 , \G16_reg/NET0131 , \G17_reg/NET0131 , \G18_reg/NET0131 , \G198_pad , \G199_pad , \G19_reg/NET0131 , \G1_pad , \G20_reg/NET0131 , \G213_pad , \G214_pad , \G21_reg/NET0131 , \G22_reg/NET0131 , \G29_reg/NET0131 , \G2_pad , \G30_reg/NET0131 , \_al_n0 , \_al_n1 , \g1001/_0_ , \g1006/_0_ , \g1008/_0_ , \g1012/_0_ , \g1020/_0_ , \g1036/_0_ , \g1056/_0_ , \g1068/_0_ , \g1070/_0_ , \g1152/_0_ , \g1298/_0_ , \g1331/_2_ , \g971/_2_ , \g973/_2_ , \g975/_2_ , \g983/_0_ , \g984/_0_ , \g985/_0_ , \g991/_2_ , \g993/_0_ , \g997/_0_ );
	input \G0_pad  ;
	input \G10_reg/NET0131  ;
	input \G11_reg/NET0131  ;
	input \G12_reg/NET0131  ;
	input \G13_reg/NET0131  ;
	input \G147_pad  ;
	input \G148_pad  ;
	input \G14_reg/NET0131  ;
	input \G15_reg/NET0131  ;
	input \G16_reg/NET0131  ;
	input \G17_reg/NET0131  ;
	input \G18_reg/NET0131  ;
	input \G198_pad  ;
	input \G199_pad  ;
	input \G19_reg/NET0131  ;
	input \G1_pad  ;
	input \G20_reg/NET0131  ;
	input \G213_pad  ;
	input \G214_pad  ;
	input \G21_reg/NET0131  ;
	input \G22_reg/NET0131  ;
	input \G29_reg/NET0131  ;
	input \G2_pad  ;
	input \G30_reg/NET0131  ;
	output \_al_n0  ;
	output \_al_n1  ;
	output \g1001/_0_  ;
	output \g1006/_0_  ;
	output \g1008/_0_  ;
	output \g1012/_0_  ;
	output \g1020/_0_  ;
	output \g1036/_0_  ;
	output \g1056/_0_  ;
	output \g1068/_0_  ;
	output \g1070/_0_  ;
	output \g1152/_0_  ;
	output \g1298/_0_  ;
	output \g1331/_2_  ;
	output \g971/_2_  ;
	output \g973/_2_  ;
	output \g975/_2_  ;
	output \g983/_0_  ;
	output \g984/_0_  ;
	output \g985/_0_  ;
	output \g991/_2_  ;
	output \g993/_0_  ;
	output \g997/_0_  ;
	wire _w94_ ;
	wire _w93_ ;
	wire _w92_ ;
	wire _w91_ ;
	wire _w90_ ;
	wire _w89_ ;
	wire _w88_ ;
	wire _w87_ ;
	wire _w86_ ;
	wire _w85_ ;
	wire _w54_ ;
	wire _w53_ ;
	wire _w52_ ;
	wire _w51_ ;
	wire _w50_ ;
	wire _w49_ ;
	wire _w48_ ;
	wire _w47_ ;
	wire _w46_ ;
	wire _w45_ ;
	wire _w44_ ;
	wire _w43_ ;
	wire _w42_ ;
	wire _w41_ ;
	wire _w40_ ;
	wire _w39_ ;
	wire _w26_ ;
	wire _w27_ ;
	wire _w28_ ;
	wire _w29_ ;
	wire _w30_ ;
	wire _w31_ ;
	wire _w32_ ;
	wire _w33_ ;
	wire _w34_ ;
	wire _w35_ ;
	wire _w36_ ;
	wire _w37_ ;
	wire _w38_ ;
	wire _w55_ ;
	wire _w56_ ;
	wire _w57_ ;
	wire _w58_ ;
	wire _w59_ ;
	wire _w60_ ;
	wire _w61_ ;
	wire _w62_ ;
	wire _w63_ ;
	wire _w64_ ;
	wire _w65_ ;
	wire _w66_ ;
	wire _w67_ ;
	wire _w68_ ;
	wire _w69_ ;
	wire _w70_ ;
	wire _w71_ ;
	wire _w72_ ;
	wire _w73_ ;
	wire _w74_ ;
	wire _w75_ ;
	wire _w76_ ;
	wire _w77_ ;
	wire _w78_ ;
	wire _w79_ ;
	wire _w80_ ;
	wire _w81_ ;
	wire _w82_ ;
	wire _w83_ ;
	wire _w84_ ;
	LUT4 #(
		.INIT('h0200)
	) name0 (
		\G10_reg/NET0131 ,
		\G11_reg/NET0131 ,
		\G14_reg/NET0131 ,
		\G15_reg/NET0131 ,
		_w26_
	);
	LUT3 #(
		.INIT('ha8)
	) name1 (
		\G16_reg/NET0131 ,
		\G30_reg/NET0131 ,
		_w26_,
		_w27_
	);
	LUT4 #(
		.INIT('h8880)
	) name2 (
		\G16_reg/NET0131 ,
		\G17_reg/NET0131 ,
		\G30_reg/NET0131 ,
		_w26_,
		_w28_
	);
	LUT3 #(
		.INIT('h14)
	) name3 (
		\G0_pad ,
		\G18_reg/NET0131 ,
		_w28_,
		_w29_
	);
	LUT4 #(
		.INIT('h0200)
	) name4 (
		\G16_reg/NET0131 ,
		\G17_reg/NET0131 ,
		\G18_reg/NET0131 ,
		\G19_reg/NET0131 ,
		_w30_
	);
	LUT3 #(
		.INIT('he0)
	) name5 (
		\G30_reg/NET0131 ,
		_w26_,
		_w30_,
		_w31_
	);
	LUT4 #(
		.INIT('ha800)
	) name6 (
		\G20_reg/NET0131 ,
		\G30_reg/NET0131 ,
		_w26_,
		_w30_,
		_w32_
	);
	LUT3 #(
		.INIT('h14)
	) name7 (
		\G0_pad ,
		\G20_reg/NET0131 ,
		_w31_,
		_w33_
	);
	LUT2 #(
		.INIT('h2)
	) name8 (
		\G12_reg/NET0131 ,
		\G13_reg/NET0131 ,
		_w34_
	);
	LUT3 #(
		.INIT('h02)
	) name9 (
		\G20_reg/NET0131 ,
		\G21_reg/NET0131 ,
		\G29_reg/NET0131 ,
		_w35_
	);
	LUT3 #(
		.INIT('h10)
	) name10 (
		\G20_reg/NET0131 ,
		\G21_reg/NET0131 ,
		\G29_reg/NET0131 ,
		_w36_
	);
	LUT4 #(
		.INIT('h11d5)
	) name11 (
		\G22_reg/NET0131 ,
		_w34_,
		_w35_,
		_w36_,
		_w37_
	);
	LUT2 #(
		.INIT('h1)
	) name12 (
		\G0_pad ,
		_w37_,
		_w38_
	);
	LUT4 #(
		.INIT('h1114)
	) name13 (
		\G0_pad ,
		\G16_reg/NET0131 ,
		\G30_reg/NET0131 ,
		_w26_,
		_w39_
	);
	LUT3 #(
		.INIT('h80)
	) name14 (
		\G10_reg/NET0131 ,
		\G11_reg/NET0131 ,
		\G14_reg/NET0131 ,
		_w40_
	);
	LUT4 #(
		.INIT('h1540)
	) name15 (
		\G0_pad ,
		\G10_reg/NET0131 ,
		\G11_reg/NET0131 ,
		\G14_reg/NET0131 ,
		_w41_
	);
	LUT4 #(
		.INIT('h5551)
	) name16 (
		\G0_pad ,
		\G10_reg/NET0131 ,
		\G11_reg/NET0131 ,
		\G14_reg/NET0131 ,
		_w42_
	);
	LUT3 #(
		.INIT('h60)
	) name17 (
		\G15_reg/NET0131 ,
		_w40_,
		_w42_,
		_w43_
	);
	LUT4 #(
		.INIT('h1311)
	) name18 (
		\G10_reg/NET0131 ,
		\G11_reg/NET0131 ,
		\G14_reg/NET0131 ,
		\G15_reg/NET0131 ,
		_w44_
	);
	LUT3 #(
		.INIT('h15)
	) name19 (
		\G0_pad ,
		\G10_reg/NET0131 ,
		\G11_reg/NET0131 ,
		_w45_
	);
	LUT2 #(
		.INIT('h4)
	) name20 (
		_w44_,
		_w45_,
		_w46_
	);
	LUT3 #(
		.INIT('h14)
	) name21 (
		\G0_pad ,
		\G1_pad ,
		\G30_reg/NET0131 ,
		_w47_
	);
	LUT3 #(
		.INIT('h14)
	) name22 (
		\G0_pad ,
		\G29_reg/NET0131 ,
		\G2_pad ,
		_w48_
	);
	LUT2 #(
		.INIT('h1)
	) name23 (
		\G0_pad ,
		\G10_reg/NET0131 ,
		_w49_
	);
	LUT2 #(
		.INIT('h6)
	) name24 (
		\G12_reg/NET0131 ,
		\G21_reg/NET0131 ,
		_w50_
	);
	LUT2 #(
		.INIT('h4)
	) name25 (
		\G0_pad ,
		\G13_reg/NET0131 ,
		_w51_
	);
	LUT3 #(
		.INIT('hd0)
	) name26 (
		_w32_,
		_w50_,
		_w51_,
		_w52_
	);
	LUT2 #(
		.INIT('h4)
	) name27 (
		\G0_pad ,
		\G12_reg/NET0131 ,
		_w53_
	);
	LUT3 #(
		.INIT('h40)
	) name28 (
		\G13_reg/NET0131 ,
		\G20_reg/NET0131 ,
		\G21_reg/NET0131 ,
		_w54_
	);
	LUT2 #(
		.INIT('h8)
	) name29 (
		_w53_,
		_w54_,
		_w55_
	);
	LUT2 #(
		.INIT('h8)
	) name30 (
		_w31_,
		_w55_,
		_w56_
	);
	LUT2 #(
		.INIT('he)
	) name31 (
		_w52_,
		_w56_,
		_w57_
	);
	LUT3 #(
		.INIT('h02)
	) name32 (
		\G13_reg/NET0131 ,
		\G20_reg/NET0131 ,
		\G21_reg/NET0131 ,
		_w58_
	);
	LUT4 #(
		.INIT('h1555)
	) name33 (
		\G12_reg/NET0131 ,
		\G13_reg/NET0131 ,
		\G199_pad ,
		\G21_reg/NET0131 ,
		_w59_
	);
	LUT2 #(
		.INIT('h4)
	) name34 (
		_w58_,
		_w59_,
		_w60_
	);
	LUT2 #(
		.INIT('h2)
	) name35 (
		\G13_reg/NET0131 ,
		\G22_reg/NET0131 ,
		_w61_
	);
	LUT4 #(
		.INIT('h0008)
	) name36 (
		\G12_reg/NET0131 ,
		\G13_reg/NET0131 ,
		\G199_pad ,
		\G22_reg/NET0131 ,
		_w62_
	);
	LUT4 #(
		.INIT('h001d)
	) name37 (
		\G18_reg/NET0131 ,
		_w37_,
		_w60_,
		_w62_,
		_w63_
	);
	LUT4 #(
		.INIT('hddd9)
	) name38 (
		\G12_reg/NET0131 ,
		\G13_reg/NET0131 ,
		\G20_reg/NET0131 ,
		\G21_reg/NET0131 ,
		_w64_
	);
	LUT4 #(
		.INIT('h0e0a)
	) name39 (
		\G12_reg/NET0131 ,
		\G13_reg/NET0131 ,
		\G148_pad ,
		\G21_reg/NET0131 ,
		_w65_
	);
	LUT3 #(
		.INIT('h10)
	) name40 (
		_w54_,
		_w65_,
		_w64_,
		_w66_
	);
	LUT2 #(
		.INIT('h8)
	) name41 (
		_w37_,
		_w66_,
		_w67_
	);
	LUT4 #(
		.INIT('h0e0a)
	) name42 (
		\G12_reg/NET0131 ,
		\G13_reg/NET0131 ,
		\G198_pad ,
		\G21_reg/NET0131 ,
		_w68_
	);
	LUT2 #(
		.INIT('h2)
	) name43 (
		_w64_,
		_w68_,
		_w69_
	);
	LUT2 #(
		.INIT('h8)
	) name44 (
		_w37_,
		_w69_,
		_w70_
	);
	LUT3 #(
		.INIT('h1b)
	) name45 (
		\G13_reg/NET0131 ,
		\G20_reg/NET0131 ,
		\G214_pad ,
		_w71_
	);
	LUT3 #(
		.INIT('hd8)
	) name46 (
		\G12_reg/NET0131 ,
		\G13_reg/NET0131 ,
		\G21_reg/NET0131 ,
		_w72_
	);
	LUT2 #(
		.INIT('h4)
	) name47 (
		_w71_,
		_w72_,
		_w73_
	);
	LUT2 #(
		.INIT('h8)
	) name48 (
		_w37_,
		_w73_,
		_w74_
	);
	LUT3 #(
		.INIT('h04)
	) name49 (
		\G0_pad ,
		\G21_reg/NET0131 ,
		_w32_,
		_w75_
	);
	LUT2 #(
		.INIT('h4)
	) name50 (
		\G12_reg/NET0131 ,
		\G13_reg/NET0131 ,
		_w76_
	);
	LUT3 #(
		.INIT('h04)
	) name51 (
		\G0_pad ,
		\G20_reg/NET0131 ,
		\G21_reg/NET0131 ,
		_w77_
	);
	LUT2 #(
		.INIT('h4)
	) name52 (
		_w76_,
		_w77_,
		_w78_
	);
	LUT2 #(
		.INIT('h8)
	) name53 (
		_w31_,
		_w78_,
		_w79_
	);
	LUT2 #(
		.INIT('he)
	) name54 (
		_w75_,
		_w79_,
		_w80_
	);
	LUT3 #(
		.INIT('h04)
	) name55 (
		\G12_reg/NET0131 ,
		\G20_reg/NET0131 ,
		\G21_reg/NET0131 ,
		_w81_
	);
	LUT3 #(
		.INIT('h32)
	) name56 (
		\G12_reg/NET0131 ,
		\G213_pad ,
		\G21_reg/NET0131 ,
		_w82_
	);
	LUT3 #(
		.INIT('h02)
	) name57 (
		_w61_,
		_w82_,
		_w81_,
		_w83_
	);
	LUT3 #(
		.INIT('hf1)
	) name58 (
		\G18_reg/NET0131 ,
		_w37_,
		_w83_,
		_w84_
	);
	LUT4 #(
		.INIT('h1444)
	) name59 (
		\G0_pad ,
		\G12_reg/NET0131 ,
		\G21_reg/NET0131 ,
		_w32_,
		_w85_
	);
	LUT3 #(
		.INIT('h13)
	) name60 (
		\G18_reg/NET0131 ,
		\G19_reg/NET0131 ,
		_w28_,
		_w86_
	);
	LUT3 #(
		.INIT('h6e)
	) name61 (
		\G17_reg/NET0131 ,
		\G18_reg/NET0131 ,
		\G19_reg/NET0131 ,
		_w87_
	);
	LUT4 #(
		.INIT('h00a8)
	) name62 (
		\G16_reg/NET0131 ,
		\G30_reg/NET0131 ,
		_w26_,
		_w87_,
		_w88_
	);
	LUT2 #(
		.INIT('h1)
	) name63 (
		\G0_pad ,
		_w88_,
		_w89_
	);
	LUT2 #(
		.INIT('h4)
	) name64 (
		_w86_,
		_w89_,
		_w90_
	);
	LUT4 #(
		.INIT('he2a2)
	) name65 (
		\G12_reg/NET0131 ,
		\G13_reg/NET0131 ,
		\G147_pad ,
		\G21_reg/NET0131 ,
		_w91_
	);
	LUT2 #(
		.INIT('h8)
	) name66 (
		_w37_,
		_w91_,
		_w92_
	);
	LUT2 #(
		.INIT('h4)
	) name67 (
		\G18_reg/NET0131 ,
		\G19_reg/NET0131 ,
		_w93_
	);
	LUT4 #(
		.INIT('h0414)
	) name68 (
		\G0_pad ,
		\G17_reg/NET0131 ,
		_w27_,
		_w93_,
		_w94_
	);
	assign \_al_n0  = 1'b0;
	assign \_al_n1  = 1'b1;
	assign \g1001/_0_  = _w29_ ;
	assign \g1006/_0_  = _w33_ ;
	assign \g1008/_0_  = _w38_ ;
	assign \g1012/_0_  = _w39_ ;
	assign \g1020/_0_  = _w41_ ;
	assign \g1036/_0_  = _w43_ ;
	assign \g1056/_0_  = _w46_ ;
	assign \g1068/_0_  = _w47_ ;
	assign \g1070/_0_  = _w48_ ;
	assign \g1152/_0_  = _w49_ ;
	assign \g1298/_0_  = _w57_ ;
	assign \g1331/_2_  = _w63_ ;
	assign \g971/_2_  = _w67_ ;
	assign \g973/_2_  = _w70_ ;
	assign \g975/_2_  = _w74_ ;
	assign \g983/_0_  = _w80_ ;
	assign \g984/_0_  = _w84_ ;
	assign \g985/_0_  = _w85_ ;
	assign \g991/_2_  = _w90_ ;
	assign \g993/_0_  = _w92_ ;
	assign \g997/_0_  = _w94_ ;
endmodule;