module top (\v0_pad , \v10_reg/NET0131 , \v11_reg/NET0131 , \v12_reg/NET0131 , \v1_pad , \v2_pad , \v3_pad , \v4_pad , \v5_pad , \v6_pad , \v7_reg/NET0131 , \v8_reg/NET0131 , \v9_reg/NET0131 , \_al_n0 , \_al_n1 , \g528/_2_ , \g534/_0_ , \g535/_0_ , \g537/_0_ , \g560/_3_ , \g722/_0_ , \g754/_0_ , \v13_D_10_pad , \v13_D_11_pad , \v13_D_12_pad , \v13_D_6_pad , \v13_D_7_pad , \v13_D_9_pad );
	input \v0_pad  ;
	input \v10_reg/NET0131  ;
	input \v11_reg/NET0131  ;
	input \v12_reg/NET0131  ;
	input \v1_pad  ;
	input \v2_pad  ;
	input \v3_pad  ;
	input \v4_pad  ;
	input \v5_pad  ;
	input \v6_pad  ;
	input \v7_reg/NET0131  ;
	input \v8_reg/NET0131  ;
	input \v9_reg/NET0131  ;
	output \_al_n0  ;
	output \_al_n1  ;
	output \g528/_2_  ;
	output \g534/_0_  ;
	output \g535/_0_  ;
	output \g537/_0_  ;
	output \g560/_3_  ;
	output \g722/_0_  ;
	output \g754/_0_  ;
	output \v13_D_10_pad  ;
	output \v13_D_11_pad  ;
	output \v13_D_12_pad  ;
	output \v13_D_6_pad  ;
	output \v13_D_7_pad  ;
	output \v13_D_9_pad  ;
	wire _w138_ ;
	wire _w137_ ;
	wire _w136_ ;
	wire _w135_ ;
	wire _w134_ ;
	wire _w133_ ;
	wire _w132_ ;
	wire _w131_ ;
	wire _w130_ ;
	wire _w129_ ;
	wire _w128_ ;
	wire _w127_ ;
	wire _w126_ ;
	wire _w125_ ;
	wire _w124_ ;
	wire _w123_ ;
	wire _w122_ ;
	wire _w121_ ;
	wire _w120_ ;
	wire _w119_ ;
	wire _w118_ ;
	wire _w117_ ;
	wire _w116_ ;
	wire _w115_ ;
	wire _w114_ ;
	wire _w113_ ;
	wire _w112_ ;
	wire _w111_ ;
	wire _w110_ ;
	wire _w109_ ;
	wire _w108_ ;
	wire _w107_ ;
	wire _w106_ ;
	wire _w105_ ;
	wire _w104_ ;
	wire _w103_ ;
	wire _w102_ ;
	wire _w101_ ;
	wire _w100_ ;
	wire _w99_ ;
	wire _w98_ ;
	wire _w97_ ;
	wire _w96_ ;
	wire _w95_ ;
	wire _w94_ ;
	wire _w93_ ;
	wire _w92_ ;
	wire _w91_ ;
	wire _w90_ ;
	wire _w89_ ;
	wire _w88_ ;
	wire _w87_ ;
	wire _w86_ ;
	wire _w85_ ;
	wire _w84_ ;
	wire _w83_ ;
	wire _w82_ ;
	wire _w81_ ;
	wire _w80_ ;
	wire _w79_ ;
	wire _w78_ ;
	wire _w77_ ;
	wire _w76_ ;
	wire _w75_ ;
	wire _w74_ ;
	wire _w73_ ;
	wire _w42_ ;
	wire _w41_ ;
	wire _w40_ ;
	wire _w39_ ;
	wire _w38_ ;
	wire _w37_ ;
	wire _w36_ ;
	wire _w35_ ;
	wire _w34_ ;
	wire _w33_ ;
	wire _w32_ ;
	wire _w31_ ;
	wire _w30_ ;
	wire _w29_ ;
	wire _w28_ ;
	wire _w27_ ;
	wire _w14_ ;
	wire _w15_ ;
	wire _w16_ ;
	wire _w17_ ;
	wire _w18_ ;
	wire _w19_ ;
	wire _w20_ ;
	wire _w21_ ;
	wire _w22_ ;
	wire _w23_ ;
	wire _w24_ ;
	wire _w25_ ;
	wire _w26_ ;
	wire _w43_ ;
	wire _w44_ ;
	wire _w45_ ;
	wire _w46_ ;
	wire _w47_ ;
	wire _w48_ ;
	wire _w49_ ;
	wire _w50_ ;
	wire _w51_ ;
	wire _w52_ ;
	wire _w53_ ;
	wire _w54_ ;
	wire _w55_ ;
	wire _w56_ ;
	wire _w57_ ;
	wire _w58_ ;
	wire _w59_ ;
	wire _w60_ ;
	wire _w61_ ;
	wire _w62_ ;
	wire _w63_ ;
	wire _w64_ ;
	wire _w65_ ;
	wire _w66_ ;
	wire _w67_ ;
	wire _w68_ ;
	wire _w69_ ;
	wire _w70_ ;
	wire _w71_ ;
	wire _w72_ ;
	LUT2 #(
		.INIT('h1)
	) name0 (
		\v12_reg/NET0131 ,
		\v9_reg/NET0131 ,
		_w14_
	);
	LUT2 #(
		.INIT('h1)
	) name1 (
		\v0_pad ,
		\v10_reg/NET0131 ,
		_w15_
	);
	LUT2 #(
		.INIT('h8)
	) name2 (
		_w14_,
		_w15_,
		_w16_
	);
	LUT2 #(
		.INIT('h1)
	) name3 (
		\v7_reg/NET0131 ,
		\v8_reg/NET0131 ,
		_w17_
	);
	LUT2 #(
		.INIT('h8)
	) name4 (
		\v1_pad ,
		_w17_,
		_w18_
	);
	LUT2 #(
		.INIT('h1)
	) name5 (
		\v10_reg/NET0131 ,
		\v9_reg/NET0131 ,
		_w19_
	);
	LUT2 #(
		.INIT('h2)
	) name6 (
		\v0_pad ,
		\v11_reg/NET0131 ,
		_w20_
	);
	LUT2 #(
		.INIT('h4)
	) name7 (
		\v12_reg/NET0131 ,
		_w20_,
		_w21_
	);
	LUT2 #(
		.INIT('h1)
	) name8 (
		_w19_,
		_w21_,
		_w22_
	);
	LUT2 #(
		.INIT('h2)
	) name9 (
		_w18_,
		_w22_,
		_w23_
	);
	LUT2 #(
		.INIT('h4)
	) name10 (
		\v12_reg/NET0131 ,
		\v1_pad ,
		_w24_
	);
	LUT2 #(
		.INIT('h8)
	) name11 (
		_w19_,
		_w24_,
		_w25_
	);
	LUT2 #(
		.INIT('h1)
	) name12 (
		\v11_reg/NET0131 ,
		\v12_reg/NET0131 ,
		_w26_
	);
	LUT2 #(
		.INIT('h8)
	) name13 (
		\v9_reg/NET0131 ,
		_w26_,
		_w27_
	);
	LUT2 #(
		.INIT('h4)
	) name14 (
		\v5_pad ,
		_w27_,
		_w28_
	);
	LUT2 #(
		.INIT('h2)
	) name15 (
		\v10_reg/NET0131 ,
		_w28_,
		_w29_
	);
	LUT2 #(
		.INIT('h4)
	) name16 (
		\v0_pad ,
		_w17_,
		_w30_
	);
	LUT2 #(
		.INIT('h4)
	) name17 (
		_w29_,
		_w30_,
		_w31_
	);
	LUT2 #(
		.INIT('h1)
	) name18 (
		_w16_,
		_w25_,
		_w32_
	);
	LUT2 #(
		.INIT('h4)
	) name19 (
		_w23_,
		_w32_,
		_w33_
	);
	LUT2 #(
		.INIT('h4)
	) name20 (
		_w31_,
		_w33_,
		_w34_
	);
	LUT2 #(
		.INIT('h2)
	) name21 (
		\v1_pad ,
		\v9_reg/NET0131 ,
		_w35_
	);
	LUT2 #(
		.INIT('h2)
	) name22 (
		\v0_pad ,
		_w35_,
		_w36_
	);
	LUT2 #(
		.INIT('h2)
	) name23 (
		\v10_reg/NET0131 ,
		_w26_,
		_w37_
	);
	LUT2 #(
		.INIT('h2)
	) name24 (
		_w17_,
		_w36_,
		_w38_
	);
	LUT2 #(
		.INIT('h4)
	) name25 (
		_w37_,
		_w38_,
		_w39_
	);
	LUT2 #(
		.INIT('h8)
	) name26 (
		\v10_reg/NET0131 ,
		_w17_,
		_w40_
	);
	LUT2 #(
		.INIT('h1)
	) name27 (
		\v11_reg/NET0131 ,
		\v5_pad ,
		_w41_
	);
	LUT2 #(
		.INIT('h8)
	) name28 (
		_w40_,
		_w41_,
		_w42_
	);
	LUT2 #(
		.INIT('h1)
	) name29 (
		_w19_,
		_w42_,
		_w43_
	);
	LUT2 #(
		.INIT('h2)
	) name30 (
		_w24_,
		_w43_,
		_w44_
	);
	LUT2 #(
		.INIT('h1)
	) name31 (
		_w16_,
		_w39_,
		_w45_
	);
	LUT2 #(
		.INIT('h4)
	) name32 (
		_w44_,
		_w45_,
		_w46_
	);
	LUT2 #(
		.INIT('h2)
	) name33 (
		\v11_reg/NET0131 ,
		\v8_reg/NET0131 ,
		_w47_
	);
	LUT2 #(
		.INIT('h8)
	) name34 (
		\v12_reg/NET0131 ,
		_w47_,
		_w48_
	);
	LUT2 #(
		.INIT('h8)
	) name35 (
		\v3_pad ,
		\v8_reg/NET0131 ,
		_w49_
	);
	LUT2 #(
		.INIT('h8)
	) name36 (
		\v2_pad ,
		_w26_,
		_w50_
	);
	LUT2 #(
		.INIT('h8)
	) name37 (
		_w49_,
		_w50_,
		_w51_
	);
	LUT2 #(
		.INIT('h1)
	) name38 (
		_w48_,
		_w51_,
		_w52_
	);
	LUT2 #(
		.INIT('h1)
	) name39 (
		\v7_reg/NET0131 ,
		_w52_,
		_w53_
	);
	LUT2 #(
		.INIT('h8)
	) name40 (
		\v11_reg/NET0131 ,
		\v7_reg/NET0131 ,
		_w54_
	);
	LUT2 #(
		.INIT('h4)
	) name41 (
		\v12_reg/NET0131 ,
		\v8_reg/NET0131 ,
		_w55_
	);
	LUT2 #(
		.INIT('h8)
	) name42 (
		_w54_,
		_w55_,
		_w56_
	);
	LUT2 #(
		.INIT('h1)
	) name43 (
		_w53_,
		_w56_,
		_w57_
	);
	LUT2 #(
		.INIT('h1)
	) name44 (
		\v10_reg/NET0131 ,
		\v1_pad ,
		_w58_
	);
	LUT2 #(
		.INIT('h2)
	) name45 (
		\v0_pad ,
		\v9_reg/NET0131 ,
		_w59_
	);
	LUT2 #(
		.INIT('h8)
	) name46 (
		_w58_,
		_w59_,
		_w60_
	);
	LUT2 #(
		.INIT('h4)
	) name47 (
		_w57_,
		_w60_,
		_w61_
	);
	LUT2 #(
		.INIT('h4)
	) name48 (
		\v12_reg/NET0131 ,
		_w60_,
		_w62_
	);
	LUT2 #(
		.INIT('h1)
	) name49 (
		\v11_reg/NET0131 ,
		\v3_pad ,
		_w63_
	);
	LUT2 #(
		.INIT('h4)
	) name50 (
		\v4_pad ,
		_w63_,
		_w64_
	);
	LUT2 #(
		.INIT('h8)
	) name51 (
		\v8_reg/NET0131 ,
		_w64_,
		_w65_
	);
	LUT2 #(
		.INIT('h8)
	) name52 (
		\v7_reg/NET0131 ,
		\v8_reg/NET0131 ,
		_w66_
	);
	LUT2 #(
		.INIT('h2)
	) name53 (
		\v11_reg/NET0131 ,
		_w66_,
		_w67_
	);
	LUT2 #(
		.INIT('h1)
	) name54 (
		_w65_,
		_w67_,
		_w68_
	);
	LUT2 #(
		.INIT('h2)
	) name55 (
		_w62_,
		_w68_,
		_w69_
	);
	LUT2 #(
		.INIT('h1)
	) name56 (
		\v11_reg/NET0131 ,
		\v7_reg/NET0131 ,
		_w70_
	);
	LUT2 #(
		.INIT('h4)
	) name57 (
		\v8_reg/NET0131 ,
		_w70_,
		_w71_
	);
	LUT2 #(
		.INIT('h4)
	) name58 (
		\v12_reg/NET0131 ,
		_w71_,
		_w72_
	);
	LUT2 #(
		.INIT('h2)
	) name59 (
		\v10_reg/NET0131 ,
		\v6_pad ,
		_w73_
	);
	LUT2 #(
		.INIT('h8)
	) name60 (
		_w59_,
		_w73_,
		_w74_
	);
	LUT2 #(
		.INIT('h8)
	) name61 (
		_w72_,
		_w74_,
		_w75_
	);
	LUT2 #(
		.INIT('h2)
	) name62 (
		\v2_pad ,
		\v8_reg/NET0131 ,
		_w76_
	);
	LUT2 #(
		.INIT('h1)
	) name63 (
		\v7_reg/NET0131 ,
		_w76_,
		_w77_
	);
	LUT2 #(
		.INIT('h2)
	) name64 (
		\v4_pad ,
		_w77_,
		_w78_
	);
	LUT2 #(
		.INIT('h8)
	) name65 (
		\v3_pad ,
		_w66_,
		_w79_
	);
	LUT2 #(
		.INIT('h1)
	) name66 (
		_w78_,
		_w79_,
		_w80_
	);
	LUT2 #(
		.INIT('h1)
	) name67 (
		\v11_reg/NET0131 ,
		_w80_,
		_w81_
	);
	LUT2 #(
		.INIT('h8)
	) name68 (
		\v7_reg/NET0131 ,
		_w47_,
		_w82_
	);
	LUT2 #(
		.INIT('h8)
	) name69 (
		\v5_pad ,
		_w82_,
		_w83_
	);
	LUT2 #(
		.INIT('h1)
	) name70 (
		\v2_pad ,
		\v7_reg/NET0131 ,
		_w84_
	);
	LUT2 #(
		.INIT('h8)
	) name71 (
		_w49_,
		_w84_,
		_w85_
	);
	LUT2 #(
		.INIT('h1)
	) name72 (
		\v7_reg/NET0131 ,
		_w26_,
		_w86_
	);
	LUT2 #(
		.INIT('h4)
	) name73 (
		_w47_,
		_w86_,
		_w87_
	);
	LUT2 #(
		.INIT('h1)
	) name74 (
		_w83_,
		_w85_,
		_w88_
	);
	LUT2 #(
		.INIT('h4)
	) name75 (
		_w87_,
		_w88_,
		_w89_
	);
	LUT2 #(
		.INIT('h4)
	) name76 (
		_w81_,
		_w89_,
		_w90_
	);
	LUT2 #(
		.INIT('h2)
	) name77 (
		\v12_reg/NET0131 ,
		_w71_,
		_w91_
	);
	LUT2 #(
		.INIT('h2)
	) name78 (
		_w60_,
		_w91_,
		_w92_
	);
	LUT2 #(
		.INIT('h4)
	) name79 (
		_w90_,
		_w92_,
		_w93_
	);
	LUT2 #(
		.INIT('h8)
	) name80 (
		_w26_,
		_w76_,
		_w94_
	);
	LUT2 #(
		.INIT('h1)
	) name81 (
		\v7_reg/NET0131 ,
		_w65_,
		_w95_
	);
	LUT2 #(
		.INIT('h1)
	) name82 (
		\v12_reg/NET0131 ,
		_w95_,
		_w96_
	);
	LUT2 #(
		.INIT('h4)
	) name83 (
		\v7_reg/NET0131 ,
		_w48_,
		_w97_
	);
	LUT2 #(
		.INIT('h4)
	) name84 (
		\v5_pad ,
		_w97_,
		_w98_
	);
	LUT2 #(
		.INIT('h1)
	) name85 (
		_w94_,
		_w98_,
		_w99_
	);
	LUT2 #(
		.INIT('h4)
	) name86 (
		_w96_,
		_w99_,
		_w100_
	);
	LUT2 #(
		.INIT('h2)
	) name87 (
		_w60_,
		_w100_,
		_w101_
	);
	LUT2 #(
		.INIT('h8)
	) name88 (
		\v0_pad ,
		\v5_pad ,
		_w102_
	);
	LUT2 #(
		.INIT('h2)
	) name89 (
		\v10_reg/NET0131 ,
		_w102_,
		_w103_
	);
	LUT2 #(
		.INIT('h8)
	) name90 (
		_w18_,
		_w27_,
		_w104_
	);
	LUT2 #(
		.INIT('h4)
	) name91 (
		_w103_,
		_w104_,
		_w105_
	);
	LUT2 #(
		.INIT('h2)
	) name92 (
		\v12_reg/NET0131 ,
		_w17_,
		_w106_
	);
	LUT2 #(
		.INIT('h2)
	) name93 (
		\v1_pad ,
		_w106_,
		_w107_
	);
	LUT2 #(
		.INIT('h1)
	) name94 (
		_w54_,
		_w64_,
		_w108_
	);
	LUT2 #(
		.INIT('h2)
	) name95 (
		_w55_,
		_w108_,
		_w109_
	);
	LUT2 #(
		.INIT('h1)
	) name96 (
		_w107_,
		_w109_,
		_w110_
	);
	LUT2 #(
		.INIT('h1)
	) name97 (
		\v10_reg/NET0131 ,
		_w110_,
		_w111_
	);
	LUT2 #(
		.INIT('h8)
	) name98 (
		_w21_,
		_w40_,
		_w112_
	);
	LUT2 #(
		.INIT('h1)
	) name99 (
		_w111_,
		_w112_,
		_w113_
	);
	LUT2 #(
		.INIT('h1)
	) name100 (
		\v9_reg/NET0131 ,
		_w113_,
		_w114_
	);
	LUT2 #(
		.INIT('h1)
	) name101 (
		_w14_,
		_w17_,
		_w115_
	);
	LUT2 #(
		.INIT('h2)
	) name102 (
		_w15_,
		_w115_,
		_w116_
	);
	LUT2 #(
		.INIT('h1)
	) name103 (
		_w114_,
		_w116_,
		_w117_
	);
	LUT2 #(
		.INIT('h4)
	) name104 (
		\v0_pad ,
		\v10_reg/NET0131 ,
		_w118_
	);
	LUT2 #(
		.INIT('h8)
	) name105 (
		\v5_pad ,
		\v9_reg/NET0131 ,
		_w119_
	);
	LUT2 #(
		.INIT('h8)
	) name106 (
		_w118_,
		_w119_,
		_w120_
	);
	LUT2 #(
		.INIT('h8)
	) name107 (
		_w72_,
		_w120_,
		_w121_
	);
	LUT2 #(
		.INIT('h4)
	) name108 (
		\v3_pad ,
		\v8_reg/NET0131 ,
		_w122_
	);
	LUT2 #(
		.INIT('h1)
	) name109 (
		_w84_,
		_w122_,
		_w123_
	);
	LUT2 #(
		.INIT('h8)
	) name110 (
		\v4_pad ,
		\v7_reg/NET0131 ,
		_w124_
	);
	LUT2 #(
		.INIT('h1)
	) name111 (
		_w123_,
		_w124_,
		_w125_
	);
	LUT2 #(
		.INIT('h2)
	) name112 (
		_w26_,
		_w125_,
		_w126_
	);
	LUT2 #(
		.INIT('h8)
	) name113 (
		\v5_pad ,
		_w97_,
		_w127_
	);
	LUT2 #(
		.INIT('h1)
	) name114 (
		_w126_,
		_w127_,
		_w128_
	);
	LUT2 #(
		.INIT('h2)
	) name115 (
		_w60_,
		_w128_,
		_w129_
	);
	LUT2 #(
		.INIT('h1)
	) name116 (
		_w65_,
		_w82_,
		_w130_
	);
	LUT2 #(
		.INIT('h2)
	) name117 (
		_w62_,
		_w130_,
		_w131_
	);
	LUT2 #(
		.INIT('h8)
	) name118 (
		\v0_pad ,
		\v10_reg/NET0131 ,
		_w132_
	);
	LUT2 #(
		.INIT('h4)
	) name119 (
		\v8_reg/NET0131 ,
		_w132_,
		_w133_
	);
	LUT2 #(
		.INIT('h8)
	) name120 (
		\v4_pad ,
		_w58_,
		_w134_
	);
	LUT2 #(
		.INIT('h8)
	) name121 (
		_w122_,
		_w134_,
		_w135_
	);
	LUT2 #(
		.INIT('h1)
	) name122 (
		_w133_,
		_w135_,
		_w136_
	);
	LUT2 #(
		.INIT('h8)
	) name123 (
		_w14_,
		_w70_,
		_w137_
	);
	LUT2 #(
		.INIT('h4)
	) name124 (
		_w136_,
		_w137_,
		_w138_
	);
	assign \_al_n0  = 1'b0;
	assign \_al_n1  = 1'b0;
	assign \g528/_2_  = _w34_ ;
	assign \g534/_0_  = _w46_ ;
	assign \g535/_0_  = _w61_ ;
	assign \g537/_0_  = _w69_ ;
	assign \g560/_3_  = _w75_ ;
	assign \g722/_0_  = _w93_ ;
	assign \g754/_0_  = _w101_ ;
	assign \v13_D_10_pad  = _w105_ ;
	assign \v13_D_11_pad  = _w117_ ;
	assign \v13_D_12_pad  = _w121_ ;
	assign \v13_D_6_pad  = _w129_ ;
	assign \v13_D_7_pad  = _w131_ ;
	assign \v13_D_9_pad  = _w138_ ;
endmodule;