module top( \A[0]  , \A[1]  , \A[2]  , \A[3]  , \A[4]  , \A[5]  , \A[6]  , \A[7]  , \A[8]  , \A[9]  , \A[10]  , \A[11]  , \A[12]  , \A[13]  , \A[14]  , \A[15]  , \A[16]  , \A[17]  , \A[18]  , \A[19]  , \A[20]  , \A[21]  , \A[22]  , \A[23]  , \A[24]  , \A[25]  , \A[26]  , \A[27]  , \A[28]  , \A[29]  , \A[30]  , \A[31]  , \A[32]  , \A[33]  , \A[34]  , \A[35]  , \A[36]  , \A[37]  , \A[38]  , \A[39]  , \A[40]  , \A[41]  , \A[42]  , \A[43]  , \A[44]  , \A[45]  , \A[46]  , \A[47]  , \A[48]  , \A[49]  , \A[50]  , \A[51]  , \A[52]  , \A[53]  , \A[54]  , \A[55]  , \A[56]  , \A[57]  , \A[58]  , \A[59]  , \A[60]  , \A[61]  , \A[62]  , \A[63]  , \A[64]  , \A[65]  , \A[66]  , \A[67]  , \A[68]  , \A[69]  , \A[70]  , \A[71]  , \A[72]  , \A[73]  , \A[74]  , \A[75]  , \A[76]  , \A[77]  , \A[78]  , \A[79]  , \A[80]  , \A[81]  , \A[82]  , \A[83]  , \A[84]  , \A[85]  , \A[86]  , \A[87]  , \A[88]  , \A[89]  , \A[90]  , \A[91]  , \A[92]  , \A[93]  , \A[94]  , \A[95]  , \A[96]  , \A[97]  , \A[98]  , \A[99]  , \A[100]  , \A[101]  , \A[102]  , \A[103]  , \A[104]  , \A[105]  , \A[106]  , \A[107]  , \A[108]  , \A[109]  , \A[110]  , \A[111]  , \A[112]  , \A[113]  , \A[114]  , \A[115]  , \A[116]  , \A[117]  , \A[118]  , \A[119]  , \A[120]  , \A[121]  , \A[122]  , \A[123]  , \A[124]  , \A[125]  , \A[126]  , \A[127]  , \A[128]  , \A[129]  , \A[130]  , \A[131]  , \A[132]  , \A[133]  , \A[134]  , \A[135]  , \A[136]  , \A[137]  , \A[138]  , \A[139]  , \A[140]  , \A[141]  , \A[142]  , \A[143]  , \A[144]  , \A[145]  , \A[146]  , \A[147]  , \A[148]  , \A[149]  , \A[150]  , \A[151]  , \A[152]  , \A[153]  , \A[154]  , \A[155]  , \A[156]  , \A[157]  , \A[158]  , \A[159]  , \A[160]  , \A[161]  , \A[162]  , \A[163]  , \A[164]  , \A[165]  , \A[166]  , \A[167]  , \A[168]  , \A[169]  , \A[170]  , \A[171]  , \A[172]  , \A[173]  , \A[174]  , \A[175]  , \A[176]  , \A[177]  , \A[178]  , \A[179]  , \A[180]  , \A[181]  , \A[182]  , \A[183]  , \A[184]  , \A[185]  , \A[186]  , \A[187]  , \A[188]  , \A[189]  , \A[190]  , \A[191]  , \A[192]  , \A[193]  , \A[194]  , \A[195]  , \A[196]  , \A[197]  , \A[198]  , \A[199]  , \A[200]  , \A[201]  , \A[202]  , \A[203]  , \A[204]  , \A[205]  , \A[206]  , \A[207]  , \A[208]  , \A[209]  , \A[210]  , \A[211]  , \A[212]  , \A[213]  , \A[214]  , \A[215]  , \A[216]  , \A[217]  , \A[218]  , \A[219]  , \A[220]  , \A[221]  , \A[222]  , \A[223]  , \A[224]  , \A[225]  , \A[226]  , \A[227]  , \A[228]  , \A[229]  , \A[230]  , \A[231]  , \A[232]  , \A[233]  , \A[234]  , \A[235]  , \A[236]  , \A[237]  , \A[238]  , \A[239]  , \A[240]  , \A[241]  , \A[242]  , \A[243]  , \A[244]  , \A[245]  , \A[246]  , \A[247]  , \A[248]  , \A[249]  , \A[250]  , \A[251]  , \A[252]  , \A[253]  , \A[254]  , \A[255]  , \A[256]  , \A[257]  , \A[258]  , \A[259]  , \A[260]  , \A[261]  , \A[262]  , \A[263]  , \A[264]  , \A[265]  , \A[266]  , \A[267]  , \A[268]  , \A[269]  , \A[270]  , \A[271]  , \A[272]  , \A[273]  , \A[274]  , \A[275]  , \A[276]  , \A[277]  , \A[278]  , \A[279]  , \A[280]  , \A[281]  , \A[282]  , \A[283]  , \A[284]  , \A[285]  , \A[286]  , \A[287]  , \A[288]  , \A[289]  , \A[290]  , \A[291]  , \A[292]  , \A[293]  , \A[294]  , \A[295]  , \A[296]  , \A[297]  , \A[298]  , \A[299]  , \A[300]  , \A[301]  , \A[302]  , \A[303]  , \A[304]  , \A[305]  , \A[306]  , \A[307]  , \A[308]  , \A[309]  , \A[310]  , \A[311]  , \A[312]  , \A[313]  , \A[314]  , \A[315]  , \A[316]  , \A[317]  , \A[318]  , \A[319]  , \A[320]  , \A[321]  , \A[322]  , \A[323]  , \A[324]  , \A[325]  , \A[326]  , \A[327]  , \A[328]  , \A[329]  , \A[330]  , \A[331]  , \A[332]  , \A[333]  , \A[334]  , \A[335]  , \A[336]  , \A[337]  , \A[338]  , \A[339]  , \A[340]  , \A[341]  , \A[342]  , \A[343]  , \A[344]  , \A[345]  , \A[346]  , \A[347]  , \A[348]  , \A[349]  , \A[350]  , \A[351]  , \A[352]  , \A[353]  , \A[354]  , \A[355]  , \A[356]  , \A[357]  , \A[358]  , \A[359]  , \A[360]  , \A[361]  , \A[362]  , \A[363]  , \A[364]  , \A[365]  , \A[366]  , \A[367]  , \A[368]  , \A[369]  , \A[370]  , \A[371]  , \A[372]  , \A[373]  , \A[374]  , \A[375]  , \A[376]  , \A[377]  , \A[378]  , \A[379]  , \A[380]  , \A[381]  , \A[382]  , \A[383]  , \A[384]  , \A[385]  , \A[386]  , \A[387]  , \A[388]  , \A[389]  , \A[390]  , \A[391]  , \A[392]  , \A[393]  , \A[394]  , \A[395]  , \A[396]  , \A[397]  , \A[398]  , \A[399]  , \A[400]  , \A[401]  , \A[402]  , \A[403]  , \A[404]  , \A[405]  , \A[406]  , \A[407]  , \A[408]  , \A[409]  , \A[410]  , \A[411]  , \A[412]  , \A[413]  , \A[414]  , \A[415]  , \A[416]  , \A[417]  , \A[418]  , \A[419]  , \A[420]  , \A[421]  , \A[422]  , \A[423]  , \A[424]  , \A[425]  , \A[426]  , \A[427]  , \A[428]  , \A[429]  , \A[430]  , \A[431]  , \A[432]  , \A[433]  , \A[434]  , \A[435]  , \A[436]  , \A[437]  , \A[438]  , \A[439]  , \A[440]  , \A[441]  , \A[442]  , \A[443]  , \A[444]  , \A[445]  , \A[446]  , \A[447]  , \A[448]  , \A[449]  , \A[450]  , \A[451]  , \A[452]  , \A[453]  , \A[454]  , \A[455]  , \A[456]  , \A[457]  , \A[458]  , \A[459]  , \A[460]  , \A[461]  , \A[462]  , \A[463]  , \A[464]  , \A[465]  , \A[466]  , \A[467]  , \A[468]  , \A[469]  , \A[470]  , \A[471]  , \A[472]  , \A[473]  , \A[474]  , \A[475]  , \A[476]  , \A[477]  , \A[478]  , \A[479]  , \A[480]  , \A[481]  , \A[482]  , \A[483]  , \A[484]  , \A[485]  , \A[486]  , \A[487]  , \A[488]  , \A[489]  , \A[490]  , \A[491]  , \A[492]  , \A[493]  , \A[494]  , \A[495]  , \A[496]  , \A[497]  , \A[498]  , \A[499]  , \A[500]  , \A[501]  , \A[502]  , \A[503]  , \A[504]  , \A[505]  , \A[506]  , \A[507]  , \A[508]  , \A[509]  , \A[510]  , \A[511]  , \A[512]  , \A[513]  , \A[514]  , \A[515]  , \A[516]  , \A[517]  , \A[518]  , \A[519]  , \A[520]  , \A[521]  , \A[522]  , \A[523]  , \A[524]  , \A[525]  , \A[526]  , \A[527]  , \A[528]  , \A[529]  , \A[530]  , \A[531]  , \A[532]  , \A[533]  , \A[534]  , \A[535]  , \A[536]  , \A[537]  , \A[538]  , \A[539]  , \A[540]  , \A[541]  , \A[542]  , \A[543]  , \A[544]  , \A[545]  , \A[546]  , \A[547]  , \A[548]  , \A[549]  , \A[550]  , \A[551]  , \A[552]  , \A[553]  , \A[554]  , \A[555]  , \A[556]  , \A[557]  , \A[558]  , \A[559]  , \A[560]  , \A[561]  , \A[562]  , \A[563]  , \A[564]  , \A[565]  , \A[566]  , \A[567]  , \A[568]  , \A[569]  , \A[570]  , \A[571]  , \A[572]  , \A[573]  , \A[574]  , \A[575]  , \A[576]  , \A[577]  , \A[578]  , \A[579]  , \A[580]  , \A[581]  , \A[582]  , \A[583]  , \A[584]  , \A[585]  , \A[586]  , \A[587]  , \A[588]  , \A[589]  , \A[590]  , \A[591]  , \A[592]  , \A[593]  , \A[594]  , \A[595]  , \A[596]  , \A[597]  , \A[598]  , \A[599]  , \A[600]  , \A[601]  , \A[602]  , \A[603]  , \A[604]  , \A[605]  , \A[606]  , \A[607]  , \A[608]  , \A[609]  , \A[610]  , \A[611]  , \A[612]  , \A[613]  , \A[614]  , \A[615]  , \A[616]  , \A[617]  , \A[618]  , \A[619]  , \A[620]  , \A[621]  , \A[622]  , \A[623]  , \A[624]  , \A[625]  , \A[626]  , \A[627]  , \A[628]  , \A[629]  , \A[630]  , \A[631]  , \A[632]  , \A[633]  , \A[634]  , \A[635]  , \A[636]  , \A[637]  , \A[638]  , \A[639]  , \A[640]  , \A[641]  , \A[642]  , \A[643]  , \A[644]  , \A[645]  , \A[646]  , \A[647]  , \A[648]  , \A[649]  , \A[650]  , \A[651]  , \A[652]  , \A[653]  , \A[654]  , \A[655]  , \A[656]  , \A[657]  , \A[658]  , \A[659]  , \A[660]  , \A[661]  , \A[662]  , \A[663]  , \A[664]  , \A[665]  , \A[666]  , \A[667]  , \A[668]  , \A[669]  , \A[670]  , \A[671]  , \A[672]  , \A[673]  , \A[674]  , \A[675]  , \A[676]  , \A[677]  , \A[678]  , \A[679]  , \A[680]  , \A[681]  , \A[682]  , \A[683]  , \A[684]  , \A[685]  , \A[686]  , \A[687]  , \A[688]  , \A[689]  , \A[690]  , \A[691]  , \A[692]  , \A[693]  , \A[694]  , \A[695]  , \A[696]  , \A[697]  , \A[698]  , \A[699]  , \A[700]  , \A[701]  , \A[702]  , \A[703]  , \A[704]  , \A[705]  , \A[706]  , \A[707]  , \A[708]  , \A[709]  , \A[710]  , \A[711]  , \A[712]  , \A[713]  , \A[714]  , \A[715]  , \A[716]  , \A[717]  , \A[718]  , \A[719]  , \A[720]  , \A[721]  , \A[722]  , \A[723]  , \A[724]  , \A[725]  , \A[726]  , \A[727]  , \A[728]  , \A[729]  , \A[730]  , \A[731]  , \A[732]  , \A[733]  , \A[734]  , \A[735]  , \A[736]  , \A[737]  , \A[738]  , \A[739]  , \A[740]  , \A[741]  , \A[742]  , \A[743]  , \A[744]  , \A[745]  , \A[746]  , \A[747]  , \A[748]  , \A[749]  , \A[750]  , \A[751]  , \A[752]  , \A[753]  , \A[754]  , \A[755]  , \A[756]  , \A[757]  , \A[758]  , \A[759]  , \A[760]  , \A[761]  , \A[762]  , \A[763]  , \A[764]  , \A[765]  , \A[766]  , \A[767]  , \A[768]  , \A[769]  , \A[770]  , \A[771]  , \A[772]  , \A[773]  , \A[774]  , \A[775]  , \A[776]  , \A[777]  , \A[778]  , \A[779]  , \A[780]  , \A[781]  , \A[782]  , \A[783]  , \A[784]  , \A[785]  , \A[786]  , \A[787]  , \A[788]  , \A[789]  , \A[790]  , \A[791]  , \A[792]  , \A[793]  , \A[794]  , \A[795]  , \A[796]  , \A[797]  , \A[798]  , \A[799]  , \A[800]  , \A[801]  , \A[802]  , \A[803]  , \A[804]  , \A[805]  , \A[806]  , \A[807]  , \A[808]  , \A[809]  , \A[810]  , \A[811]  , \A[812]  , \A[813]  , \A[814]  , \A[815]  , \A[816]  , \A[817]  , \A[818]  , \A[819]  , \A[820]  , \A[821]  , \A[822]  , \A[823]  , \A[824]  , \A[825]  , \A[826]  , \A[827]  , \A[828]  , \A[829]  , \A[830]  , \A[831]  , \A[832]  , \A[833]  , \A[834]  , \A[835]  , \A[836]  , \A[837]  , \A[838]  , \A[839]  , \A[840]  , \A[841]  , \A[842]  , \A[843]  , \A[844]  , \A[845]  , \A[846]  , \A[847]  , \A[848]  , \A[849]  , \A[850]  , \A[851]  , \A[852]  , \A[853]  , \A[854]  , \A[855]  , \A[856]  , \A[857]  , \A[858]  , \A[859]  , \A[860]  , \A[861]  , \A[862]  , \A[863]  , \A[864]  , \A[865]  , \A[866]  , \A[867]  , \A[868]  , \A[869]  , \A[870]  , \A[871]  , \A[872]  , \A[873]  , \A[874]  , \A[875]  , \A[876]  , \A[877]  , \A[878]  , \A[879]  , \A[880]  , \A[881]  , \A[882]  , \A[883]  , \A[884]  , \A[885]  , \A[886]  , \A[887]  , \A[888]  , \A[889]  , \A[890]  , \A[891]  , \A[892]  , \A[893]  , \A[894]  , \A[895]  , \A[896]  , \A[897]  , \A[898]  , \A[899]  , \A[900]  , \A[901]  , \A[902]  , \A[903]  , \A[904]  , \A[905]  , \A[906]  , \A[907]  , \A[908]  , \A[909]  , \A[910]  , \A[911]  , \A[912]  , \A[913]  , \A[914]  , \A[915]  , \A[916]  , \A[917]  , \A[918]  , \A[919]  , \A[920]  , \A[921]  , \A[922]  , \A[923]  , \A[924]  , \A[925]  , \A[926]  , \A[927]  , \A[928]  , \A[929]  , \A[930]  , \A[931]  , \A[932]  , \A[933]  , \A[934]  , \A[935]  , \A[936]  , \A[937]  , \A[938]  , \A[939]  , \A[940]  , \A[941]  , \A[942]  , \A[943]  , \A[944]  , \A[945]  , \A[946]  , \A[947]  , \A[948]  , \A[949]  , \A[950]  , \A[951]  , \A[952]  , \A[953]  , \A[954]  , \A[955]  , \A[956]  , \A[957]  , \A[958]  , \A[959]  , \A[960]  , \A[961]  , \A[962]  , \A[963]  , \A[964]  , \A[965]  , \A[966]  , \A[967]  , \A[968]  , \A[969]  , \A[970]  , \A[971]  , \A[972]  , \A[973]  , \A[974]  , \A[975]  , \A[976]  , \A[977]  , \A[978]  , \A[979]  , \A[980]  , \A[981]  , \A[982]  , \A[983]  , \A[984]  , \A[985]  , \A[986]  , \A[987]  , \A[988]  , \A[989]  , \A[990]  , \A[991]  , \A[992]  , \A[993]  , \A[994]  , \A[995]  , \A[996]  , \A[997]  , \A[998]  , \A[999]  , \A[1000]  , maj );
  input \A[0]  ;
  input \A[1]  ;
  input \A[2]  ;
  input \A[3]  ;
  input \A[4]  ;
  input \A[5]  ;
  input \A[6]  ;
  input \A[7]  ;
  input \A[8]  ;
  input \A[9]  ;
  input \A[10]  ;
  input \A[11]  ;
  input \A[12]  ;
  input \A[13]  ;
  input \A[14]  ;
  input \A[15]  ;
  input \A[16]  ;
  input \A[17]  ;
  input \A[18]  ;
  input \A[19]  ;
  input \A[20]  ;
  input \A[21]  ;
  input \A[22]  ;
  input \A[23]  ;
  input \A[24]  ;
  input \A[25]  ;
  input \A[26]  ;
  input \A[27]  ;
  input \A[28]  ;
  input \A[29]  ;
  input \A[30]  ;
  input \A[31]  ;
  input \A[32]  ;
  input \A[33]  ;
  input \A[34]  ;
  input \A[35]  ;
  input \A[36]  ;
  input \A[37]  ;
  input \A[38]  ;
  input \A[39]  ;
  input \A[40]  ;
  input \A[41]  ;
  input \A[42]  ;
  input \A[43]  ;
  input \A[44]  ;
  input \A[45]  ;
  input \A[46]  ;
  input \A[47]  ;
  input \A[48]  ;
  input \A[49]  ;
  input \A[50]  ;
  input \A[51]  ;
  input \A[52]  ;
  input \A[53]  ;
  input \A[54]  ;
  input \A[55]  ;
  input \A[56]  ;
  input \A[57]  ;
  input \A[58]  ;
  input \A[59]  ;
  input \A[60]  ;
  input \A[61]  ;
  input \A[62]  ;
  input \A[63]  ;
  input \A[64]  ;
  input \A[65]  ;
  input \A[66]  ;
  input \A[67]  ;
  input \A[68]  ;
  input \A[69]  ;
  input \A[70]  ;
  input \A[71]  ;
  input \A[72]  ;
  input \A[73]  ;
  input \A[74]  ;
  input \A[75]  ;
  input \A[76]  ;
  input \A[77]  ;
  input \A[78]  ;
  input \A[79]  ;
  input \A[80]  ;
  input \A[81]  ;
  input \A[82]  ;
  input \A[83]  ;
  input \A[84]  ;
  input \A[85]  ;
  input \A[86]  ;
  input \A[87]  ;
  input \A[88]  ;
  input \A[89]  ;
  input \A[90]  ;
  input \A[91]  ;
  input \A[92]  ;
  input \A[93]  ;
  input \A[94]  ;
  input \A[95]  ;
  input \A[96]  ;
  input \A[97]  ;
  input \A[98]  ;
  input \A[99]  ;
  input \A[100]  ;
  input \A[101]  ;
  input \A[102]  ;
  input \A[103]  ;
  input \A[104]  ;
  input \A[105]  ;
  input \A[106]  ;
  input \A[107]  ;
  input \A[108]  ;
  input \A[109]  ;
  input \A[110]  ;
  input \A[111]  ;
  input \A[112]  ;
  input \A[113]  ;
  input \A[114]  ;
  input \A[115]  ;
  input \A[116]  ;
  input \A[117]  ;
  input \A[118]  ;
  input \A[119]  ;
  input \A[120]  ;
  input \A[121]  ;
  input \A[122]  ;
  input \A[123]  ;
  input \A[124]  ;
  input \A[125]  ;
  input \A[126]  ;
  input \A[127]  ;
  input \A[128]  ;
  input \A[129]  ;
  input \A[130]  ;
  input \A[131]  ;
  input \A[132]  ;
  input \A[133]  ;
  input \A[134]  ;
  input \A[135]  ;
  input \A[136]  ;
  input \A[137]  ;
  input \A[138]  ;
  input \A[139]  ;
  input \A[140]  ;
  input \A[141]  ;
  input \A[142]  ;
  input \A[143]  ;
  input \A[144]  ;
  input \A[145]  ;
  input \A[146]  ;
  input \A[147]  ;
  input \A[148]  ;
  input \A[149]  ;
  input \A[150]  ;
  input \A[151]  ;
  input \A[152]  ;
  input \A[153]  ;
  input \A[154]  ;
  input \A[155]  ;
  input \A[156]  ;
  input \A[157]  ;
  input \A[158]  ;
  input \A[159]  ;
  input \A[160]  ;
  input \A[161]  ;
  input \A[162]  ;
  input \A[163]  ;
  input \A[164]  ;
  input \A[165]  ;
  input \A[166]  ;
  input \A[167]  ;
  input \A[168]  ;
  input \A[169]  ;
  input \A[170]  ;
  input \A[171]  ;
  input \A[172]  ;
  input \A[173]  ;
  input \A[174]  ;
  input \A[175]  ;
  input \A[176]  ;
  input \A[177]  ;
  input \A[178]  ;
  input \A[179]  ;
  input \A[180]  ;
  input \A[181]  ;
  input \A[182]  ;
  input \A[183]  ;
  input \A[184]  ;
  input \A[185]  ;
  input \A[186]  ;
  input \A[187]  ;
  input \A[188]  ;
  input \A[189]  ;
  input \A[190]  ;
  input \A[191]  ;
  input \A[192]  ;
  input \A[193]  ;
  input \A[194]  ;
  input \A[195]  ;
  input \A[196]  ;
  input \A[197]  ;
  input \A[198]  ;
  input \A[199]  ;
  input \A[200]  ;
  input \A[201]  ;
  input \A[202]  ;
  input \A[203]  ;
  input \A[204]  ;
  input \A[205]  ;
  input \A[206]  ;
  input \A[207]  ;
  input \A[208]  ;
  input \A[209]  ;
  input \A[210]  ;
  input \A[211]  ;
  input \A[212]  ;
  input \A[213]  ;
  input \A[214]  ;
  input \A[215]  ;
  input \A[216]  ;
  input \A[217]  ;
  input \A[218]  ;
  input \A[219]  ;
  input \A[220]  ;
  input \A[221]  ;
  input \A[222]  ;
  input \A[223]  ;
  input \A[224]  ;
  input \A[225]  ;
  input \A[226]  ;
  input \A[227]  ;
  input \A[228]  ;
  input \A[229]  ;
  input \A[230]  ;
  input \A[231]  ;
  input \A[232]  ;
  input \A[233]  ;
  input \A[234]  ;
  input \A[235]  ;
  input \A[236]  ;
  input \A[237]  ;
  input \A[238]  ;
  input \A[239]  ;
  input \A[240]  ;
  input \A[241]  ;
  input \A[242]  ;
  input \A[243]  ;
  input \A[244]  ;
  input \A[245]  ;
  input \A[246]  ;
  input \A[247]  ;
  input \A[248]  ;
  input \A[249]  ;
  input \A[250]  ;
  input \A[251]  ;
  input \A[252]  ;
  input \A[253]  ;
  input \A[254]  ;
  input \A[255]  ;
  input \A[256]  ;
  input \A[257]  ;
  input \A[258]  ;
  input \A[259]  ;
  input \A[260]  ;
  input \A[261]  ;
  input \A[262]  ;
  input \A[263]  ;
  input \A[264]  ;
  input \A[265]  ;
  input \A[266]  ;
  input \A[267]  ;
  input \A[268]  ;
  input \A[269]  ;
  input \A[270]  ;
  input \A[271]  ;
  input \A[272]  ;
  input \A[273]  ;
  input \A[274]  ;
  input \A[275]  ;
  input \A[276]  ;
  input \A[277]  ;
  input \A[278]  ;
  input \A[279]  ;
  input \A[280]  ;
  input \A[281]  ;
  input \A[282]  ;
  input \A[283]  ;
  input \A[284]  ;
  input \A[285]  ;
  input \A[286]  ;
  input \A[287]  ;
  input \A[288]  ;
  input \A[289]  ;
  input \A[290]  ;
  input \A[291]  ;
  input \A[292]  ;
  input \A[293]  ;
  input \A[294]  ;
  input \A[295]  ;
  input \A[296]  ;
  input \A[297]  ;
  input \A[298]  ;
  input \A[299]  ;
  input \A[300]  ;
  input \A[301]  ;
  input \A[302]  ;
  input \A[303]  ;
  input \A[304]  ;
  input \A[305]  ;
  input \A[306]  ;
  input \A[307]  ;
  input \A[308]  ;
  input \A[309]  ;
  input \A[310]  ;
  input \A[311]  ;
  input \A[312]  ;
  input \A[313]  ;
  input \A[314]  ;
  input \A[315]  ;
  input \A[316]  ;
  input \A[317]  ;
  input \A[318]  ;
  input \A[319]  ;
  input \A[320]  ;
  input \A[321]  ;
  input \A[322]  ;
  input \A[323]  ;
  input \A[324]  ;
  input \A[325]  ;
  input \A[326]  ;
  input \A[327]  ;
  input \A[328]  ;
  input \A[329]  ;
  input \A[330]  ;
  input \A[331]  ;
  input \A[332]  ;
  input \A[333]  ;
  input \A[334]  ;
  input \A[335]  ;
  input \A[336]  ;
  input \A[337]  ;
  input \A[338]  ;
  input \A[339]  ;
  input \A[340]  ;
  input \A[341]  ;
  input \A[342]  ;
  input \A[343]  ;
  input \A[344]  ;
  input \A[345]  ;
  input \A[346]  ;
  input \A[347]  ;
  input \A[348]  ;
  input \A[349]  ;
  input \A[350]  ;
  input \A[351]  ;
  input \A[352]  ;
  input \A[353]  ;
  input \A[354]  ;
  input \A[355]  ;
  input \A[356]  ;
  input \A[357]  ;
  input \A[358]  ;
  input \A[359]  ;
  input \A[360]  ;
  input \A[361]  ;
  input \A[362]  ;
  input \A[363]  ;
  input \A[364]  ;
  input \A[365]  ;
  input \A[366]  ;
  input \A[367]  ;
  input \A[368]  ;
  input \A[369]  ;
  input \A[370]  ;
  input \A[371]  ;
  input \A[372]  ;
  input \A[373]  ;
  input \A[374]  ;
  input \A[375]  ;
  input \A[376]  ;
  input \A[377]  ;
  input \A[378]  ;
  input \A[379]  ;
  input \A[380]  ;
  input \A[381]  ;
  input \A[382]  ;
  input \A[383]  ;
  input \A[384]  ;
  input \A[385]  ;
  input \A[386]  ;
  input \A[387]  ;
  input \A[388]  ;
  input \A[389]  ;
  input \A[390]  ;
  input \A[391]  ;
  input \A[392]  ;
  input \A[393]  ;
  input \A[394]  ;
  input \A[395]  ;
  input \A[396]  ;
  input \A[397]  ;
  input \A[398]  ;
  input \A[399]  ;
  input \A[400]  ;
  input \A[401]  ;
  input \A[402]  ;
  input \A[403]  ;
  input \A[404]  ;
  input \A[405]  ;
  input \A[406]  ;
  input \A[407]  ;
  input \A[408]  ;
  input \A[409]  ;
  input \A[410]  ;
  input \A[411]  ;
  input \A[412]  ;
  input \A[413]  ;
  input \A[414]  ;
  input \A[415]  ;
  input \A[416]  ;
  input \A[417]  ;
  input \A[418]  ;
  input \A[419]  ;
  input \A[420]  ;
  input \A[421]  ;
  input \A[422]  ;
  input \A[423]  ;
  input \A[424]  ;
  input \A[425]  ;
  input \A[426]  ;
  input \A[427]  ;
  input \A[428]  ;
  input \A[429]  ;
  input \A[430]  ;
  input \A[431]  ;
  input \A[432]  ;
  input \A[433]  ;
  input \A[434]  ;
  input \A[435]  ;
  input \A[436]  ;
  input \A[437]  ;
  input \A[438]  ;
  input \A[439]  ;
  input \A[440]  ;
  input \A[441]  ;
  input \A[442]  ;
  input \A[443]  ;
  input \A[444]  ;
  input \A[445]  ;
  input \A[446]  ;
  input \A[447]  ;
  input \A[448]  ;
  input \A[449]  ;
  input \A[450]  ;
  input \A[451]  ;
  input \A[452]  ;
  input \A[453]  ;
  input \A[454]  ;
  input \A[455]  ;
  input \A[456]  ;
  input \A[457]  ;
  input \A[458]  ;
  input \A[459]  ;
  input \A[460]  ;
  input \A[461]  ;
  input \A[462]  ;
  input \A[463]  ;
  input \A[464]  ;
  input \A[465]  ;
  input \A[466]  ;
  input \A[467]  ;
  input \A[468]  ;
  input \A[469]  ;
  input \A[470]  ;
  input \A[471]  ;
  input \A[472]  ;
  input \A[473]  ;
  input \A[474]  ;
  input \A[475]  ;
  input \A[476]  ;
  input \A[477]  ;
  input \A[478]  ;
  input \A[479]  ;
  input \A[480]  ;
  input \A[481]  ;
  input \A[482]  ;
  input \A[483]  ;
  input \A[484]  ;
  input \A[485]  ;
  input \A[486]  ;
  input \A[487]  ;
  input \A[488]  ;
  input \A[489]  ;
  input \A[490]  ;
  input \A[491]  ;
  input \A[492]  ;
  input \A[493]  ;
  input \A[494]  ;
  input \A[495]  ;
  input \A[496]  ;
  input \A[497]  ;
  input \A[498]  ;
  input \A[499]  ;
  input \A[500]  ;
  input \A[501]  ;
  input \A[502]  ;
  input \A[503]  ;
  input \A[504]  ;
  input \A[505]  ;
  input \A[506]  ;
  input \A[507]  ;
  input \A[508]  ;
  input \A[509]  ;
  input \A[510]  ;
  input \A[511]  ;
  input \A[512]  ;
  input \A[513]  ;
  input \A[514]  ;
  input \A[515]  ;
  input \A[516]  ;
  input \A[517]  ;
  input \A[518]  ;
  input \A[519]  ;
  input \A[520]  ;
  input \A[521]  ;
  input \A[522]  ;
  input \A[523]  ;
  input \A[524]  ;
  input \A[525]  ;
  input \A[526]  ;
  input \A[527]  ;
  input \A[528]  ;
  input \A[529]  ;
  input \A[530]  ;
  input \A[531]  ;
  input \A[532]  ;
  input \A[533]  ;
  input \A[534]  ;
  input \A[535]  ;
  input \A[536]  ;
  input \A[537]  ;
  input \A[538]  ;
  input \A[539]  ;
  input \A[540]  ;
  input \A[541]  ;
  input \A[542]  ;
  input \A[543]  ;
  input \A[544]  ;
  input \A[545]  ;
  input \A[546]  ;
  input \A[547]  ;
  input \A[548]  ;
  input \A[549]  ;
  input \A[550]  ;
  input \A[551]  ;
  input \A[552]  ;
  input \A[553]  ;
  input \A[554]  ;
  input \A[555]  ;
  input \A[556]  ;
  input \A[557]  ;
  input \A[558]  ;
  input \A[559]  ;
  input \A[560]  ;
  input \A[561]  ;
  input \A[562]  ;
  input \A[563]  ;
  input \A[564]  ;
  input \A[565]  ;
  input \A[566]  ;
  input \A[567]  ;
  input \A[568]  ;
  input \A[569]  ;
  input \A[570]  ;
  input \A[571]  ;
  input \A[572]  ;
  input \A[573]  ;
  input \A[574]  ;
  input \A[575]  ;
  input \A[576]  ;
  input \A[577]  ;
  input \A[578]  ;
  input \A[579]  ;
  input \A[580]  ;
  input \A[581]  ;
  input \A[582]  ;
  input \A[583]  ;
  input \A[584]  ;
  input \A[585]  ;
  input \A[586]  ;
  input \A[587]  ;
  input \A[588]  ;
  input \A[589]  ;
  input \A[590]  ;
  input \A[591]  ;
  input \A[592]  ;
  input \A[593]  ;
  input \A[594]  ;
  input \A[595]  ;
  input \A[596]  ;
  input \A[597]  ;
  input \A[598]  ;
  input \A[599]  ;
  input \A[600]  ;
  input \A[601]  ;
  input \A[602]  ;
  input \A[603]  ;
  input \A[604]  ;
  input \A[605]  ;
  input \A[606]  ;
  input \A[607]  ;
  input \A[608]  ;
  input \A[609]  ;
  input \A[610]  ;
  input \A[611]  ;
  input \A[612]  ;
  input \A[613]  ;
  input \A[614]  ;
  input \A[615]  ;
  input \A[616]  ;
  input \A[617]  ;
  input \A[618]  ;
  input \A[619]  ;
  input \A[620]  ;
  input \A[621]  ;
  input \A[622]  ;
  input \A[623]  ;
  input \A[624]  ;
  input \A[625]  ;
  input \A[626]  ;
  input \A[627]  ;
  input \A[628]  ;
  input \A[629]  ;
  input \A[630]  ;
  input \A[631]  ;
  input \A[632]  ;
  input \A[633]  ;
  input \A[634]  ;
  input \A[635]  ;
  input \A[636]  ;
  input \A[637]  ;
  input \A[638]  ;
  input \A[639]  ;
  input \A[640]  ;
  input \A[641]  ;
  input \A[642]  ;
  input \A[643]  ;
  input \A[644]  ;
  input \A[645]  ;
  input \A[646]  ;
  input \A[647]  ;
  input \A[648]  ;
  input \A[649]  ;
  input \A[650]  ;
  input \A[651]  ;
  input \A[652]  ;
  input \A[653]  ;
  input \A[654]  ;
  input \A[655]  ;
  input \A[656]  ;
  input \A[657]  ;
  input \A[658]  ;
  input \A[659]  ;
  input \A[660]  ;
  input \A[661]  ;
  input \A[662]  ;
  input \A[663]  ;
  input \A[664]  ;
  input \A[665]  ;
  input \A[666]  ;
  input \A[667]  ;
  input \A[668]  ;
  input \A[669]  ;
  input \A[670]  ;
  input \A[671]  ;
  input \A[672]  ;
  input \A[673]  ;
  input \A[674]  ;
  input \A[675]  ;
  input \A[676]  ;
  input \A[677]  ;
  input \A[678]  ;
  input \A[679]  ;
  input \A[680]  ;
  input \A[681]  ;
  input \A[682]  ;
  input \A[683]  ;
  input \A[684]  ;
  input \A[685]  ;
  input \A[686]  ;
  input \A[687]  ;
  input \A[688]  ;
  input \A[689]  ;
  input \A[690]  ;
  input \A[691]  ;
  input \A[692]  ;
  input \A[693]  ;
  input \A[694]  ;
  input \A[695]  ;
  input \A[696]  ;
  input \A[697]  ;
  input \A[698]  ;
  input \A[699]  ;
  input \A[700]  ;
  input \A[701]  ;
  input \A[702]  ;
  input \A[703]  ;
  input \A[704]  ;
  input \A[705]  ;
  input \A[706]  ;
  input \A[707]  ;
  input \A[708]  ;
  input \A[709]  ;
  input \A[710]  ;
  input \A[711]  ;
  input \A[712]  ;
  input \A[713]  ;
  input \A[714]  ;
  input \A[715]  ;
  input \A[716]  ;
  input \A[717]  ;
  input \A[718]  ;
  input \A[719]  ;
  input \A[720]  ;
  input \A[721]  ;
  input \A[722]  ;
  input \A[723]  ;
  input \A[724]  ;
  input \A[725]  ;
  input \A[726]  ;
  input \A[727]  ;
  input \A[728]  ;
  input \A[729]  ;
  input \A[730]  ;
  input \A[731]  ;
  input \A[732]  ;
  input \A[733]  ;
  input \A[734]  ;
  input \A[735]  ;
  input \A[736]  ;
  input \A[737]  ;
  input \A[738]  ;
  input \A[739]  ;
  input \A[740]  ;
  input \A[741]  ;
  input \A[742]  ;
  input \A[743]  ;
  input \A[744]  ;
  input \A[745]  ;
  input \A[746]  ;
  input \A[747]  ;
  input \A[748]  ;
  input \A[749]  ;
  input \A[750]  ;
  input \A[751]  ;
  input \A[752]  ;
  input \A[753]  ;
  input \A[754]  ;
  input \A[755]  ;
  input \A[756]  ;
  input \A[757]  ;
  input \A[758]  ;
  input \A[759]  ;
  input \A[760]  ;
  input \A[761]  ;
  input \A[762]  ;
  input \A[763]  ;
  input \A[764]  ;
  input \A[765]  ;
  input \A[766]  ;
  input \A[767]  ;
  input \A[768]  ;
  input \A[769]  ;
  input \A[770]  ;
  input \A[771]  ;
  input \A[772]  ;
  input \A[773]  ;
  input \A[774]  ;
  input \A[775]  ;
  input \A[776]  ;
  input \A[777]  ;
  input \A[778]  ;
  input \A[779]  ;
  input \A[780]  ;
  input \A[781]  ;
  input \A[782]  ;
  input \A[783]  ;
  input \A[784]  ;
  input \A[785]  ;
  input \A[786]  ;
  input \A[787]  ;
  input \A[788]  ;
  input \A[789]  ;
  input \A[790]  ;
  input \A[791]  ;
  input \A[792]  ;
  input \A[793]  ;
  input \A[794]  ;
  input \A[795]  ;
  input \A[796]  ;
  input \A[797]  ;
  input \A[798]  ;
  input \A[799]  ;
  input \A[800]  ;
  input \A[801]  ;
  input \A[802]  ;
  input \A[803]  ;
  input \A[804]  ;
  input \A[805]  ;
  input \A[806]  ;
  input \A[807]  ;
  input \A[808]  ;
  input \A[809]  ;
  input \A[810]  ;
  input \A[811]  ;
  input \A[812]  ;
  input \A[813]  ;
  input \A[814]  ;
  input \A[815]  ;
  input \A[816]  ;
  input \A[817]  ;
  input \A[818]  ;
  input \A[819]  ;
  input \A[820]  ;
  input \A[821]  ;
  input \A[822]  ;
  input \A[823]  ;
  input \A[824]  ;
  input \A[825]  ;
  input \A[826]  ;
  input \A[827]  ;
  input \A[828]  ;
  input \A[829]  ;
  input \A[830]  ;
  input \A[831]  ;
  input \A[832]  ;
  input \A[833]  ;
  input \A[834]  ;
  input \A[835]  ;
  input \A[836]  ;
  input \A[837]  ;
  input \A[838]  ;
  input \A[839]  ;
  input \A[840]  ;
  input \A[841]  ;
  input \A[842]  ;
  input \A[843]  ;
  input \A[844]  ;
  input \A[845]  ;
  input \A[846]  ;
  input \A[847]  ;
  input \A[848]  ;
  input \A[849]  ;
  input \A[850]  ;
  input \A[851]  ;
  input \A[852]  ;
  input \A[853]  ;
  input \A[854]  ;
  input \A[855]  ;
  input \A[856]  ;
  input \A[857]  ;
  input \A[858]  ;
  input \A[859]  ;
  input \A[860]  ;
  input \A[861]  ;
  input \A[862]  ;
  input \A[863]  ;
  input \A[864]  ;
  input \A[865]  ;
  input \A[866]  ;
  input \A[867]  ;
  input \A[868]  ;
  input \A[869]  ;
  input \A[870]  ;
  input \A[871]  ;
  input \A[872]  ;
  input \A[873]  ;
  input \A[874]  ;
  input \A[875]  ;
  input \A[876]  ;
  input \A[877]  ;
  input \A[878]  ;
  input \A[879]  ;
  input \A[880]  ;
  input \A[881]  ;
  input \A[882]  ;
  input \A[883]  ;
  input \A[884]  ;
  input \A[885]  ;
  input \A[886]  ;
  input \A[887]  ;
  input \A[888]  ;
  input \A[889]  ;
  input \A[890]  ;
  input \A[891]  ;
  input \A[892]  ;
  input \A[893]  ;
  input \A[894]  ;
  input \A[895]  ;
  input \A[896]  ;
  input \A[897]  ;
  input \A[898]  ;
  input \A[899]  ;
  input \A[900]  ;
  input \A[901]  ;
  input \A[902]  ;
  input \A[903]  ;
  input \A[904]  ;
  input \A[905]  ;
  input \A[906]  ;
  input \A[907]  ;
  input \A[908]  ;
  input \A[909]  ;
  input \A[910]  ;
  input \A[911]  ;
  input \A[912]  ;
  input \A[913]  ;
  input \A[914]  ;
  input \A[915]  ;
  input \A[916]  ;
  input \A[917]  ;
  input \A[918]  ;
  input \A[919]  ;
  input \A[920]  ;
  input \A[921]  ;
  input \A[922]  ;
  input \A[923]  ;
  input \A[924]  ;
  input \A[925]  ;
  input \A[926]  ;
  input \A[927]  ;
  input \A[928]  ;
  input \A[929]  ;
  input \A[930]  ;
  input \A[931]  ;
  input \A[932]  ;
  input \A[933]  ;
  input \A[934]  ;
  input \A[935]  ;
  input \A[936]  ;
  input \A[937]  ;
  input \A[938]  ;
  input \A[939]  ;
  input \A[940]  ;
  input \A[941]  ;
  input \A[942]  ;
  input \A[943]  ;
  input \A[944]  ;
  input \A[945]  ;
  input \A[946]  ;
  input \A[947]  ;
  input \A[948]  ;
  input \A[949]  ;
  input \A[950]  ;
  input \A[951]  ;
  input \A[952]  ;
  input \A[953]  ;
  input \A[954]  ;
  input \A[955]  ;
  input \A[956]  ;
  input \A[957]  ;
  input \A[958]  ;
  input \A[959]  ;
  input \A[960]  ;
  input \A[961]  ;
  input \A[962]  ;
  input \A[963]  ;
  input \A[964]  ;
  input \A[965]  ;
  input \A[966]  ;
  input \A[967]  ;
  input \A[968]  ;
  input \A[969]  ;
  input \A[970]  ;
  input \A[971]  ;
  input \A[972]  ;
  input \A[973]  ;
  input \A[974]  ;
  input \A[975]  ;
  input \A[976]  ;
  input \A[977]  ;
  input \A[978]  ;
  input \A[979]  ;
  input \A[980]  ;
  input \A[981]  ;
  input \A[982]  ;
  input \A[983]  ;
  input \A[984]  ;
  input \A[985]  ;
  input \A[986]  ;
  input \A[987]  ;
  input \A[988]  ;
  input \A[989]  ;
  input \A[990]  ;
  input \A[991]  ;
  input \A[992]  ;
  input \A[993]  ;
  input \A[994]  ;
  input \A[995]  ;
  input \A[996]  ;
  input \A[997]  ;
  input \A[998]  ;
  input \A[999]  ;
  input \A[1000]  ;
  output maj ;
  wire n1002 , n1003 , n1004 , n1005 , n1006 , n1007 , n1008 , n1009 , n1010 , n1011 , n1012 , n1013 , n1014 , n1015 , n1016 , n1017 , n1018 , n1019 , n1020 , n1021 , n1022 , n1023 , n1024 , n1025 , n1026 , n1027 , n1028 , n1029 , n1030 , n1031 , n1032 , n1033 , n1034 , n1035 , n1036 , n1037 , n1038 , n1039 , n1040 , n1041 , n1042 , n1043 , n1044 , n1045 , n1046 , n1047 , n1048 , n1049 , n1050 , n1051 , n1052 , n1053 , n1054 , n1055 , n1056 , n1057 , n1058 , n1059 , n1060 , n1061 , n1062 , n1063 , n1064 , n1065 , n1066 , n1067 , n1068 , n1069 , n1070 , n1071 , n1072 , n1073 , n1074 , n1075 , n1076 , n1077 , n1078 , n1079 , n1080 , n1081 , n1082 , n1083 , n1084 , n1085 , n1086 , n1087 , n1088 , n1089 , n1090 , n1091 , n1092 , n1093 , n1094 , n1095 , n1096 , n1097 , n1098 , n1099 , n1100 , n1101 , n1102 , n1103 , n1104 , n1105 , n1106 , n1107 , n1108 , n1109 , n1110 , n1111 , n1112 , n1113 , n1114 , n1115 , n1116 , n1117 , n1118 , n1119 , n1120 , n1121 , n1122 , n1123 , n1124 , n1125 , n1126 , n1127 , n1128 , n1129 , n1130 , n1131 , n1132 , n1133 , n1134 , n1135 , n1136 , n1137 , n1138 , n1139 , n1140 , n1141 , n1142 , n1143 , n1144 , n1145 , n1146 , n1147 , n1148 , n1149 , n1150 , n1151 , n1152 , n1153 , n1154 , n1155 , n1156 , n1157 , n1158 , n1159 , n1160 , n1161 , n1162 , n1163 , n1164 , n1165 , n1166 , n1167 , n1168 , n1169 , n1170 , n1171 , n1172 , n1173 , n1174 , n1175 , n1176 , n1177 , n1178 , n1179 , n1180 , n1181 , n1182 , n1183 , n1184 , n1185 , n1186 , n1187 , n1188 , n1189 , n1190 , n1191 , n1192 , n1193 , n1194 , n1195 , n1196 , n1197 , n1198 , n1199 , n1200 , n1201 , n1202 , n1203 , n1204 , n1205 , n1206 , n1207 , n1208 , n1209 , n1210 , n1211 , n1212 , n1213 , n1214 , n1215 , n1216 , n1217 , n1218 , n1219 , n1220 , n1221 , n1222 , n1223 , n1224 , n1225 , n1226 , n1227 , n1228 , n1229 , n1230 , n1231 , n1232 , n1233 , n1234 , n1235 , n1236 , n1237 , n1238 , n1239 , n1240 , n1241 , n1242 , n1243 , n1244 , n1245 , n1246 , n1247 , n1248 , n1249 , n1250 , n1251 , n1252 , n1253 , n1254 , n1255 , n1256 , n1257 , n1258 , n1259 , n1260 , n1261 , n1262 , n1263 , n1264 , n1265 , n1266 , n1267 , n1268 , n1269 , n1270 , n1271 , n1272 , n1273 , n1274 , n1275 , n1276 , n1277 , n1278 , n1279 , n1280 , n1281 , n1282 , n1283 , n1284 , n1285 , n1286 , n1287 , n1288 , n1289 , n1290 , n1291 , n1292 , n1293 , n1294 , n1295 , n1296 , n1297 , n1298 , n1299 , n1300 , n1301 , n1302 , n1303 , n1304 , n1305 , n1306 , n1307 , n1308 , n1309 , n1310 , n1311 , n1312 , n1313 , n1314 , n1315 , n1316 , n1317 , n1318 , n1319 , n1320 , n1321 , n1322 , n1323 , n1324 , n1325 , n1326 , n1327 , n1328 , n1329 , n1330 , n1331 , n1332 , n1333 , n1334 , n1335 , n1336 , n1337 , n1338 , n1339 , n1340 , n1341 , n1342 , n1343 , n1344 , n1345 , n1346 , n1347 , n1348 , n1349 , n1350 , n1351 , n1352 , n1353 , n1354 , n1355 , n1356 , n1357 , n1358 , n1359 , n1360 , n1361 , n1362 , n1363 , n1364 , n1365 , n1366 , n1367 , n1368 , n1369 , n1370 , n1371 , n1372 , n1373 , n1374 , n1375 , n1376 , n1377 , n1378 , n1379 , n1380 , n1381 , n1382 , n1383 , n1384 , n1385 , n1386 , n1387 , n1388 , n1389 , n1390 , n1391 , n1392 , n1393 , n1394 , n1395 , n1396 , n1397 , n1398 , n1399 , n1400 , n1401 , n1402 , n1403 , n1404 , n1405 , n1406 , n1407 , n1408 , n1409 , n1410 , n1411 , n1412 , n1413 , n1414 , n1415 , n1416 , n1417 , n1418 , n1419 , n1420 , n1421 , n1422 , n1423 , n1424 , n1425 , n1426 , n1427 , n1428 , n1429 , n1430 , n1431 , n1432 , n1433 , n1434 , n1435 , n1436 , n1437 , n1438 , n1439 , n1440 , n1441 , n1442 , n1443 , n1444 , n1445 , n1446 , n1447 , n1448 , n1449 , n1450 , n1451 , n1452 , n1453 , n1454 , n1455 , n1456 , n1457 , n1458 , n1459 , n1460 , n1461 , n1462 , n1463 , n1464 , n1465 , n1466 , n1467 , n1468 , n1469 , n1470 , n1471 , n1472 , n1473 , n1474 , n1475 , n1476 , n1477 , n1478 , n1479 , n1480 , n1481 , n1482 , n1483 , n1484 , n1485 , n1486 , n1487 , n1488 , n1489 , n1490 , n1491 , n1492 , n1493 , n1494 , n1495 , n1496 , n1497 , n1498 , n1499 , n1500 , n1501 , n1502 , n1503 , n1504 , n1505 , n1506 , n1507 , n1508 , n1509 , n1510 , n1511 , n1512 , n1513 , n1514 , n1515 , n1516 , n1517 , n1518 , n1519 , n1520 , n1521 , n1522 , n1523 , n1524 , n1525 , n1526 , n1527 , n1528 , n1529 , n1530 , n1531 , n1532 , n1533 , n1534 , n1535 , n1536 , n1537 , n1538 , n1539 , n1540 , n1541 , n1542 , n1543 , n1544 , n1545 , n1546 , n1547 , n1548 , n1549 , n1550 , n1551 , n1552 , n1553 , n1554 , n1555 , n1556 , n1557 , n1558 , n1559 , n1560 , n1561 , n1562 , n1563 , n1564 , n1565 , n1566 , n1567 , n1568 , n1569 , n1570 , n1571 , n1572 , n1573 , n1574 , n1575 , n1576 , n1577 , n1578 , n1579 , n1580 , n1581 , n1582 , n1583 , n1584 , n1585 , n1586 , n1587 , n1588 , n1589 , n1590 , n1591 , n1592 , n1593 , n1594 , n1595 , n1596 , n1597 , n1598 , n1599 , n1600 , n1601 , n1602 , n1603 , n1604 , n1605 , n1606 , n1607 , n1608 , n1609 , n1610 , n1611 , n1612 , n1613 , n1614 , n1615 , n1616 , n1617 , n1618 , n1619 , n1620 , n1621 , n1622 , n1623 , n1624 , n1625 , n1626 , n1627 , n1628 , n1629 , n1630 , n1631 , n1632 , n1633 , n1634 , n1635 , n1636 , n1637 , n1638 , n1639 , n1640 , n1641 , n1642 , n1643 , n1644 , n1645 , n1646 , n1647 , n1648 , n1649 , n1650 , n1651 , n1652 , n1653 , n1654 , n1655 , n1656 , n1657 , n1658 , n1659 , n1660 , n1661 , n1662 , n1663 , n1664 , n1665 , n1666 , n1667 , n1668 , n1669 , n1670 , n1671 , n1672 , n1673 , n1674 , n1675 , n1676 , n1677 , n1678 , n1679 , n1680 , n1681 , n1682 , n1683 , n1684 , n1685 , n1686 , n1687 , n1688 , n1689 , n1690 , n1691 , n1692 , n1693 , n1694 , n1695 , n1696 , n1697 , n1698 , n1699 , n1700 , n1701 , n1702 , n1703 , n1704 , n1705 , n1706 , n1707 , n1708 , n1709 , n1710 , n1711 , n1712 , n1713 , n1714 , n1715 , n1716 , n1717 , n1718 , n1719 , n1720 , n1721 , n1722 , n1723 , n1724 , n1725 , n1726 , n1727 , n1728 , n1729 , n1730 , n1731 , n1732 , n1733 , n1734 , n1735 , n1736 , n1737 , n1738 , n1739 , n1740 , n1741 , n1742 , n1743 , n1744 , n1745 , n1746 , n1747 , n1748 , n1749 , n1750 , n1751 , n1752 , n1753 , n1754 , n1755 , n1756 , n1757 , n1758 , n1759 , n1760 , n1761 , n1762 , n1763 , n1764 , n1765 , n1766 , n1767 , n1768 , n1769 , n1770 , n1771 , n1772 , n1773 , n1774 , n1775 , n1776 , n1777 , n1778 , n1779 , n1780 , n1781 , n1782 , n1783 , n1784 , n1785 , n1786 , n1787 , n1788 , n1789 , n1790 , n1791 , n1792 , n1793 , n1794 , n1795 , n1796 , n1797 , n1798 , n1799 , n1800 , n1801 , n1802 , n1803 , n1804 , n1805 , n1806 , n1807 , n1808 , n1809 , n1810 , n1811 , n1812 , n1813 , n1814 , n1815 , n1816 , n1817 , n1818 , n1819 , n1820 , n1821 , n1822 , n1823 , n1824 , n1825 , n1826 , n1827 , n1828 , n1829 , n1830 , n1831 , n1832 , n1833 , n1834 , n1835 , n1836 , n1837 , n1838 , n1839 , n1840 , n1841 , n1842 , n1843 , n1844 , n1845 , n1846 , n1847 , n1848 , n1849 , n1850 , n1851 , n1852 , n1853 , n1854 , n1855 , n1856 , n1857 , n1858 , n1859 , n1860 , n1861 , n1862 , n1863 , n1864 , n1865 , n1866 , n1867 , n1868 , n1869 , n1870 , n1871 , n1872 , n1873 , n1874 , n1875 , n1876 , n1877 , n1878 , n1879 , n1880 , n1881 , n1882 , n1883 , n1884 , n1885 , n1886 , n1887 , n1888 , n1889 , n1890 , n1891 , n1892 , n1893 , n1894 , n1895 , n1896 , n1897 , n1898 , n1899 , n1900 , n1901 , n1902 , n1903 , n1904 , n1905 , n1906 , n1907 , n1908 , n1909 , n1910 , n1911 , n1912 , n1913 , n1914 , n1915 , n1916 , n1917 , n1918 , n1919 , n1920 , n1921 , n1922 , n1923 , n1924 , n1925 , n1926 , n1927 , n1928 , n1929 , n1930 , n1931 , n1932 , n1933 , n1934 , n1935 , n1936 , n1937 , n1938 , n1939 , n1940 , n1941 , n1942 , n1943 , n1944 , n1945 , n1946 , n1947 , n1948 , n1949 , n1950 , n1951 , n1952 , n1953 , n1954 , n1955 , n1956 , n1957 , n1958 , n1959 , n1960 , n1961 , n1962 , n1963 , n1964 , n1965 , n1966 , n1967 , n1968 , n1969 , n1970 , n1971 , n1972 , n1973 , n1974 , n1975 , n1976 , n1977 , n1978 , n1979 , n1980 , n1981 , n1982 , n1983 , n1984 , n1985 , n1986 , n1987 , n1988 , n1989 , n1990 , n1991 , n1992 , n1993 , n1994 , n1995 , n1996 , n1997 , n1998 , n1999 , n2000 , n2001 , n2002 , n2003 , n2004 , n2005 , n2006 , n2007 , n2008 , n2009 , n2010 , n2011 , n2012 , n2013 , n2014 , n2015 , n2016 , n2017 , n2018 , n2019 , n2020 , n2021 , n2022 , n2023 , n2024 , n2025 , n2026 , n2027 , n2028 , n2029 , n2030 , n2031 , n2032 , n2033 , n2034 , n2035 , n2036 , n2037 , n2038 , n2039 , n2040 , n2041 , n2042 , n2043 , n2044 , n2045 , n2046 , n2047 , n2048 , n2049 , n2050 , n2051 , n2052 , n2053 , n2054 , n2055 , n2056 , n2057 , n2058 , n2059 , n2060 , n2061 , n2062 , n2063 , n2064 , n2065 , n2066 , n2067 , n2068 , n2069 , n2070 , n2071 , n2072 , n2073 , n2074 , n2075 , n2076 , n2077 , n2078 , n2079 , n2080 , n2081 , n2082 , n2083 , n2084 , n2085 , n2086 , n2087 , n2088 , n2089 , n2090 , n2091 , n2092 , n2093 , n2094 , n2095 , n2096 , n2097 , n2098 , n2099 , n2100 , n2101 , n2102 , n2103 , n2104 , n2105 , n2106 , n2107 , n2108 , n2109 , n2110 , n2111 , n2112 , n2113 , n2114 , n2115 , n2116 , n2117 , n2118 , n2119 , n2120 , n2121 , n2122 , n2123 , n2124 , n2125 , n2126 , n2127 , n2128 , n2129 , n2130 , n2131 , n2132 , n2133 , n2134 , n2135 , n2136 , n2137 , n2138 , n2139 , n2140 , n2141 , n2142 , n2143 , n2144 , n2145 , n2146 , n2147 , n2148 , n2149 , n2150 , n2151 , n2152 , n2153 , n2154 , n2155 , n2156 , n2157 , n2158 , n2159 , n2160 , n2161 , n2162 , n2163 , n2164 , n2165 , n2166 , n2167 , n2168 , n2169 , n2170 , n2171 , n2172 , n2173 , n2174 , n2175 , n2176 , n2177 , n2178 , n2179 , n2180 , n2181 , n2182 , n2183 , n2184 , n2185 , n2186 , n2187 , n2188 , n2189 , n2190 , n2191 , n2192 , n2193 , n2194 , n2195 , n2196 , n2197 , n2198 , n2199 , n2200 , n2201 , n2202 , n2203 , n2204 , n2205 , n2206 , n2207 , n2208 , n2209 , n2210 , n2211 , n2212 , n2213 , n2214 , n2215 , n2216 , n2217 , n2218 , n2219 , n2220 , n2221 , n2222 , n2223 , n2224 , n2225 , n2226 , n2227 , n2228 , n2229 , n2230 , n2231 , n2232 , n2233 , n2234 , n2235 , n2236 , n2237 , n2238 , n2239 , n2240 , n2241 , n2242 , n2243 , n2244 , n2245 , n2246 , n2247 , n2248 , n2249 , n2250 , n2251 , n2252 , n2253 , n2254 , n2255 , n2256 , n2257 , n2258 , n2259 , n2260 , n2261 , n2262 , n2263 , n2264 , n2265 , n2266 , n2267 , n2268 , n2269 , n2270 , n2271 , n2272 , n2273 , n2274 , n2275 , n2276 , n2277 , n2278 , n2279 , n2280 , n2281 , n2282 , n2283 , n2284 , n2285 , n2286 , n2287 , n2288 , n2289 , n2290 , n2291 , n2292 , n2293 , n2294 , n2295 , n2296 , n2297 , n2298 , n2299 , n2300 , n2301 , n2302 , n2303 , n2304 , n2305 , n2306 , n2307 , n2308 , n2309 , n2310 , n2311 , n2312 , n2313 , n2314 , n2315 , n2316 , n2317 , n2318 , n2319 , n2320 , n2321 , n2322 , n2323 , n2324 , n2325 , n2326 , n2327 , n2328 , n2329 , n2330 , n2331 , n2332 , n2333 , n2334 , n2335 , n2336 , n2337 , n2338 , n2339 , n2340 , n2341 , n2342 , n2343 , n2344 , n2345 , n2346 , n2347 , n2348 , n2349 , n2350 , n2351 , n2352 , n2353 , n2354 , n2355 , n2356 , n2357 , n2358 , n2359 , n2360 , n2361 , n2362 , n2363 , n2364 , n2365 , n2366 , n2367 , n2368 , n2369 , n2370 , n2371 , n2372 , n2373 , n2374 , n2375 , n2376 , n2377 , n2378 , n2379 , n2380 , n2381 , n2382 , n2383 , n2384 , n2385 , n2386 , n2387 , n2388 , n2389 , n2390 , n2391 , n2392 , n2393 , n2394 , n2395 , n2396 , n2397 , n2398 , n2399 , n2400 , n2401 , n2402 , n2403 , n2404 , n2405 , n2406 , n2407 , n2408 , n2409 , n2410 , n2411 , n2412 , n2413 , n2414 , n2415 , n2416 , n2417 , n2418 , n2419 , n2420 , n2421 , n2422 , n2423 , n2424 , n2425 , n2426 , n2427 , n2428 , n2429 , n2430 , n2431 , n2432 , n2433 , n2434 , n2435 , n2436 , n2437 , n2438 , n2439 , n2440 , n2441 , n2442 , n2443 , n2444 , n2445 , n2446 , n2447 , n2448 , n2449 , n2450 , n2451 , n2452 , n2453 , n2454 , n2455 , n2456 , n2457 , n2458 , n2459 , n2460 , n2461 , n2462 , n2463 , n2464 , n2465 , n2466 , n2467 , n2468 , n2469 , n2470 , n2471 , n2472 , n2473 , n2474 , n2475 , n2476 , n2477 , n2478 , n2479 , n2480 , n2481 , n2482 , n2483 , n2484 , n2485 , n2486 , n2487 , n2488 , n2489 , n2490 , n2491 , n2492 , n2493 , n2494 , n2495 , n2496 , n2497 , n2498 , n2499 , n2500 , n2501 , n2502 , n2503 , n2504 , n2505 , n2506 , n2507 , n2508 , n2509 , n2510 , n2511 , n2512 , n2513 , n2514 , n2515 , n2516 , n2517 , n2518 , n2519 , n2520 , n2521 , n2522 , n2523 , n2524 , n2525 , n2526 , n2527 , n2528 , n2529 , n2530 , n2531 , n2532 , n2533 , n2534 , n2535 , n2536 , n2537 , n2538 , n2539 , n2540 , n2541 , n2542 , n2543 , n2544 , n2545 , n2546 , n2547 , n2548 , n2549 , n2550 , n2551 , n2552 , n2553 , n2554 , n2555 , n2556 , n2557 , n2558 , n2559 , n2560 , n2561 , n2562 , n2563 , n2564 , n2565 , n2566 , n2567 , n2568 , n2569 , n2570 , n2571 , n2572 , n2573 , n2574 , n2575 , n2576 , n2577 , n2578 , n2579 , n2580 , n2581 , n2582 , n2583 , n2584 , n2585 , n2586 , n2587 , n2588 , n2589 , n2590 , n2591 , n2592 , n2593 , n2594 , n2595 , n2596 , n2597 , n2598 , n2599 , n2600 , n2601 , n2602 , n2603 , n2604 , n2605 , n2606 , n2607 , n2608 , n2609 , n2610 , n2611 , n2612 , n2613 , n2614 , n2615 , n2616 , n2617 , n2618 , n2619 , n2620 , n2621 , n2622 , n2623 , n2624 , n2625 , n2626 , n2627 , n2628 , n2629 , n2630 , n2631 , n2632 , n2633 , n2634 , n2635 , n2636 , n2637 , n2638 , n2639 , n2640 , n2641 , n2642 , n2643 , n2644 , n2645 , n2646 , n2647 , n2648 , n2649 , n2650 , n2651 , n2652 , n2653 , n2654 , n2655 , n2656 , n2657 , n2658 , n2659 , n2660 , n2661 , n2662 , n2663 , n2664 , n2665 , n2666 , n2667 , n2668 , n2669 , n2670 , n2671 , n2672 , n2673 , n2674 , n2675 , n2676 , n2677 , n2678 , n2679 , n2680 , n2681 , n2682 , n2683 , n2684 , n2685 , n2686 , n2687 , n2688 , n2689 , n2690 , n2691 , n2692 , n2693 , n2694 , n2695 , n2696 , n2697 , n2698 , n2699 , n2700 , n2701 , n2702 , n2703 , n2704 , n2705 , n2706 , n2707 , n2708 , n2709 , n2710 , n2711 , n2712 , n2713 , n2714 , n2715 , n2716 , n2717 , n2718 , n2719 , n2720 , n2721 , n2722 , n2723 , n2724 , n2725 , n2726 , n2727 , n2728 , n2729 , n2730 , n2731 , n2732 , n2733 , n2734 , n2735 , n2736 , n2737 , n2738 , n2739 , n2740 , n2741 , n2742 , n2743 , n2744 , n2745 , n2746 , n2747 , n2748 , n2749 , n2750 , n2751 , n2752 , n2753 , n2754 , n2755 , n2756 , n2757 , n2758 , n2759 , n2760 , n2761 , n2762 , n2763 , n2764 , n2765 , n2766 , n2767 , n2768 , n2769 , n2770 , n2771 , n2772 , n2773 , n2774 , n2775 , n2776 , n2777 , n2778 , n2779 , n2780 , n2781 , n2782 , n2783 , n2784 , n2785 , n2786 , n2787 , n2788 , n2789 , n2790 , n2791 , n2792 , n2793 , n2794 , n2795 , n2796 , n2797 , n2798 , n2799 , n2800 , n2801 , n2802 , n2803 , n2804 , n2805 , n2806 , n2807 , n2808 , n2809 , n2810 , n2811 , n2812 , n2813 , n2814 , n2815 , n2816 , n2817 , n2818 , n2819 , n2820 , n2821 , n2822 , n2823 , n2824 , n2825 , n2826 , n2827 , n2828 , n2829 , n2830 , n2831 , n2832 , n2833 , n2834 , n2835 , n2836 , n2837 , n2838 , n2839 , n2840 , n2841 , n2842 , n2843 , n2844 , n2845 , n2846 , n2847 , n2848 , n2849 , n2850 , n2851 , n2852 , n2853 , n2854 , n2855 , n2856 , n2857 , n2858 , n2859 , n2860 , n2861 , n2862 , n2863 , n2864 , n2865 , n2866 , n2867 , n2868 , n2869 , n2870 , n2871 , n2872 , n2873 , n2874 , n2875 , n2876 , n2877 , n2878 , n2879 , n2880 , n2881 , n2882 , n2883 , n2884 , n2885 , n2886 , n2887 , n2888 , n2889 , n2890 , n2891 , n2892 , n2893 , n2894 , n2895 , n2896 , n2897 , n2898 , n2899 , n2900 , n2901 , n2902 , n2903 , n2904 , n2905 , n2906 , n2907 , n2908 , n2909 , n2910 , n2911 , n2912 , n2913 , n2914 , n2915 , n2916 , n2917 , n2918 , n2919 , n2920 , n2921 , n2922 , n2923 , n2924 , n2925 , n2926 , n2927 , n2928 , n2929 , n2930 , n2931 , n2932 , n2933 , n2934 , n2935 , n2936 , n2937 , n2938 , n2939 , n2940 , n2941 , n2942 , n2943 , n2944 , n2945 , n2946 , n2947 , n2948 , n2949 , n2950 , n2951 , n2952 , n2953 , n2954 , n2955 , n2956 , n2957 , n2958 , n2959 , n2960 , n2961 , n2962 , n2963 , n2964 , n2965 , n2966 , n2967 , n2968 , n2969 , n2970 , n2971 , n2972 , n2973 , n2974 , n2975 , n2976 , n2977 , n2978 , n2979 , n2980 , n2981 , n2982 , n2983 , n2984 , n2985 , n2986 , n2987 , n2988 , n2989 , n2990 , n2991 , n2992 , n2993 , n2994 , n2995 , n2996 , n2997 , n2998 , n2999 , n3000 , n3001 , n3002 , n3003 , n3004 , n3005 , n3006 , n3007 , n3008 , n3009 , n3010 , n3011 , n3012 , n3013 , n3014 , n3015 , n3016 , n3017 , n3018 , n3019 , n3020 , n3021 , n3022 , n3023 , n3024 , n3025 , n3026 , n3027 , n3028 , n3029 , n3030 , n3031 , n3032 , n3033 , n3034 , n3035 , n3036 , n3037 , n3038 , n3039 , n3040 , n3041 , n3042 , n3043 , n3044 , n3045 , n3046 , n3047 , n3048 , n3049 , n3050 , n3051 , n3052 , n3053 , n3054 , n3055 , n3056 , n3057 , n3058 , n3059 , n3060 , n3061 , n3062 , n3063 , n3064 , n3065 , n3066 , n3067 , n3068 , n3069 , n3070 , n3071 , n3072 , n3073 , n3074 , n3075 , n3076 , n3077 , n3078 , n3079 , n3080 , n3081 , n3082 , n3083 , n3084 , n3085 , n3086 , n3087 , n3088 , n3089 , n3090 , n3091 , n3092 , n3093 , n3094 , n3095 , n3096 , n3097 , n3098 , n3099 , n3100 , n3101 , n3102 , n3103 , n3104 , n3105 , n3106 , n3107 , n3108 , n3109 , n3110 , n3111 , n3112 , n3113 , n3114 , n3115 , n3116 , n3117 , n3118 , n3119 , n3120 , n3121 , n3122 , n3123 , n3124 , n3125 , n3126 , n3127 , n3128 , n3129 , n3130 , n3131 , n3132 , n3133 , n3134 , n3135 , n3136 , n3137 , n3138 , n3139 , n3140 , n3141 , n3142 , n3143 , n3144 , n3145 , n3146 , n3147 , n3148 , n3149 , n3150 , n3151 , n3152 , n3153 , n3154 , n3155 , n3156 , n3157 , n3158 , n3159 , n3160 , n3161 , n3162 , n3163 , n3164 , n3165 , n3166 , n3167 , n3168 , n3169 , n3170 , n3171 , n3172 , n3173 , n3174 , n3175 , n3176 , n3177 , n3178 , n3179 , n3180 , n3181 , n3182 , n3183 , n3184 , n3185 , n3186 , n3187 , n3188 , n3189 , n3190 , n3191 , n3192 , n3193 , n3194 , n3195 , n3196 , n3197 , n3198 , n3199 , n3200 , n3201 , n3202 , n3203 , n3204 , n3205 , n3206 , n3207 , n3208 , n3209 , n3210 , n3211 , n3212 , n3213 , n3214 , n3215 , n3216 , n3217 , n3218 , n3219 , n3220 , n3221 , n3222 , n3223 , n3224 , n3225 , n3226 , n3227 , n3228 , n3229 , n3230 , n3231 , n3232 , n3233 , n3234 , n3235 , n3236 , n3237 , n3238 , n3239 , n3240 , n3241 , n3242 , n3243 , n3244 , n3245 , n3246 , n3247 , n3248 , n3249 , n3250 , n3251 , n3252 , n3253 , n3254 , n3255 , n3256 , n3257 , n3258 , n3259 , n3260 , n3261 , n3262 , n3263 , n3264 , n3265 , n3266 , n3267 , n3268 , n3269 , n3270 , n3271 , n3272 , n3273 , n3274 , n3275 , n3276 , n3277 , n3278 , n3279 , n3280 , n3281 , n3282 , n3283 , n3284 , n3285 , n3286 , n3287 , n3288 , n3289 , n3290 , n3291 , n3292 , n3293 , n3294 , n3295 , n3296 , n3297 , n3298 , n3299 , n3300 , n3301 , n3302 , n3303 , n3304 , n3305 , n3306 , n3307 , n3308 , n3309 , n3310 , n3311 , n3312 , n3313 , n3314 , n3315 , n3316 , n3317 , n3318 , n3319 , n3320 , n3321 , n3322 , n3323 , n3324 , n3325 , n3326 , n3327 , n3328 , n3329 , n3330 , n3331 , n3332 , n3333 , n3334 , n3335 , n3336 , n3337 , n3338 , n3339 , n3340 , n3341 , n3342 , n3343 , n3344 , n3345 , n3346 , n3347 , n3348 , n3349 , n3350 , n3351 , n3352 , n3353 , n3354 , n3355 , n3356 , n3357 , n3358 , n3359 , n3360 , n3361 , n3362 , n3363 , n3364 , n3365 , n3366 , n3367 , n3368 , n3369 , n3370 , n3371 , n3372 , n3373 , n3374 , n3375 , n3376 , n3377 , n3378 , n3379 , n3380 , n3381 , n3382 , n3383 , n3384 , n3385 , n3386 , n3387 , n3388 , n3389 , n3390 , n3391 , n3392 , n3393 , n3394 , n3395 , n3396 , n3397 , n3398 , n3399 , n3400 , n3401 , n3402 , n3403 , n3404 , n3405 , n3406 , n3407 , n3408 , n3409 , n3410 , n3411 , n3412 , n3413 , n3414 , n3415 , n3416 , n3417 , n3418 , n3419 , n3420 , n3421 , n3422 , n3423 , n3424 , n3425 , n3426 , n3427 , n3428 , n3429 , n3430 , n3431 , n3432 , n3433 , n3434 , n3435 , n3436 , n3437 , n3438 , n3439 , n3440 , n3441 , n3442 , n3443 , n3444 , n3445 , n3446 , n3447 , n3448 , n3449 , n3450 , n3451 , n3452 , n3453 , n3454 , n3455 , n3456 , n3457 , n3458 , n3459 , n3460 , n3461 , n3462 , n3463 , n3464 , n3465 , n3466 , n3467 , n3468 , n3469 , n3470 , n3471 , n3472 , n3473 , n3474 , n3475 , n3476 , n3477 , n3478 , n3479 , n3480 , n3481 , n3482 , n3483 , n3484 , n3485 , n3486 , n3487 , n3488 , n3489 , n3490 , n3491 , n3492 , n3493 , n3494 , n3495 , n3496 , n3497 , n3498 , n3499 , n3500 , n3501 , n3502 , n3503 , n3504 , n3505 , n3506 , n3507 , n3508 , n3509 , n3510 , n3511 , n3512 , n3513 , n3514 , n3515 , n3516 , n3517 , n3518 , n3519 , n3520 , n3521 , n3522 , n3523 , n3524 , n3525 , n3526 , n3527 , n3528 , n3529 , n3530 , n3531 , n3532 , n3533 , n3534 , n3535 , n3536 , n3537 , n3538 , n3539 , n3540 , n3541 , n3542 , n3543 , n3544 , n3545 , n3546 , n3547 , n3548 , n3549 , n3550 , n3551 , n3552 , n3553 , n3554 , n3555 , n3556 , n3557 , n3558 , n3559 , n3560 , n3561 , n3562 , n3563 , n3564 , n3565 , n3566 , n3567 , n3568 , n3569 , n3570 , n3571 , n3572 , n3573 , n3574 , n3575 , n3576 , n3577 , n3578 , n3579 , n3580 , n3581 , n3582 , n3583 , n3584 , n3585 , n3586 , n3587 , n3588 , n3589 , n3590 , n3591 , n3592 , n3593 , n3594 , n3595 , n3596 , n3597 , n3598 , n3599 , n3600 , n3601 , n3602 , n3603 , n3604 , n3605 , n3606 , n3607 , n3608 , n3609 , n3610 , n3611 , n3612 , n3613 , n3614 , n3615 , n3616 , n3617 , n3618 , n3619 , n3620 , n3621 , n3622 , n3623 , n3624 , n3625 , n3626 , n3627 , n3628 , n3629 , n3630 , n3631 , n3632 , n3633 , n3634 , n3635 , n3636 , n3637 , n3638 , n3639 , n3640 , n3641 , n3642 , n3643 , n3644 , n3645 , n3646 , n3647 , n3648 , n3649 , n3650 , n3651 , n3652 , n3653 , n3654 , n3655 , n3656 , n3657 , n3658 , n3659 , n3660 , n3661 , n3662 , n3663 , n3664 , n3665 , n3666 , n3667 , n3668 , n3669 , n3670 , n3671 , n3672 , n3673 , n3674 , n3675 , n3676 , n3677 , n3678 , n3679 , n3680 , n3681 , n3682 , n3683 , n3684 , n3685 , n3686 , n3687 , n3688 , n3689 , n3690 , n3691 , n3692 , n3693 , n3694 , n3695 , n3696 , n3697 , n3698 , n3699 , n3700 , n3701 , n3702 , n3703 , n3704 , n3705 , n3706 , n3707 , n3708 , n3709 , n3710 , n3711 , n3712 , n3713 , n3714 , n3715 , n3716 , n3717 , n3718 , n3719 , n3720 , n3721 , n3722 , n3723 , n3724 , n3725 , n3726 , n3727 , n3728 , n3729 , n3730 , n3731 , n3732 , n3733 , n3734 , n3735 , n3736 , n3737 , n3738 , n3739 , n3740 , n3741 , n3742 , n3743 , n3744 , n3745 , n3746 , n3747 , n3748 , n3749 , n3750 , n3751 , n3752 , n3753 , n3754 , n3755 , n3756 , n3757 , n3758 , n3759 , n3760 , n3761 , n3762 , n3763 , n3764 , n3765 , n3766 , n3767 , n3768 , n3769 , n3770 , n3771 , n3772 , n3773 , n3774 , n3775 , n3776 , n3777 , n3778 , n3779 , n3780 , n3781 , n3782 , n3783 , n3784 , n3785 , n3786 , n3787 , n3788 , n3789 , n3790 , n3791 , n3792 , n3793 , n3794 , n3795 , n3796 , n3797 , n3798 , n3799 , n3800 , n3801 , n3802 , n3803 , n3804 , n3805 , n3806 , n3807 , n3808 , n3809 , n3810 , n3811 , n3812 , n3813 , n3814 , n3815 , n3816 , n3817 , n3818 , n3819 , n3820 , n3821 , n3822 , n3823 , n3824 , n3825 , n3826 , n3827 , n3828 , n3829 , n3830 , n3831 , n3832 , n3833 , n3834 , n3835 , n3836 , n3837 , n3838 , n3839 , n3840 , n3841 , n3842 , n3843 , n3844 , n3845 , n3846 , n3847 , n3848 , n3849 , n3850 , n3851 , n3852 , n3853 , n3854 , n3855 , n3856 , n3857 , n3858 , n3859 , n3860 , n3861 , n3862 , n3863 , n3864 , n3865 , n3866 , n3867 , n3868 , n3869 , n3870 , n3871 , n3872 , n3873 , n3874 , n3875 , n3876 , n3877 , n3878 , n3879 , n3880 , n3881 , n3882 , n3883 , n3884 , n3885 , n3886 , n3887 , n3888 , n3889 , n3890 , n3891 , n3892 , n3893 , n3894 , n3895 , n3896 , n3897 , n3898 , n3899 , n3900 , n3901 , n3902 , n3903 , n3904 , n3905 , n3906 , n3907 , n3908 , n3909 , n3910 , n3911 , n3912 , n3913 , n3914 , n3915 , n3916 , n3917 , n3918 , n3919 , n3920 , n3921 , n3922 , n3923 , n3924 , n3925 , n3926 , n3927 , n3928 , n3929 , n3930 , n3931 , n3932 , n3933 , n3934 , n3935 , n3936 , n3937 , n3938 , n3939 , n3940 , n3941 , n3942 , n3943 , n3944 , n3945 , n3946 , n3947 , n3948 , n3949 , n3950 , n3951 , n3952 , n3953 , n3954 , n3955 , n3956 , n3957 , n3958 , n3959 , n3960 , n3961 , n3962 , n3963 , n3964 , n3965 , n3966 , n3967 , n3968 , n3969 , n3970 , n3971 , n3972 , n3973 , n3974 , n3975 , n3976 , n3977 , n3978 , n3979 , n3980 , n3981 , n3982 , n3983 , n3984 , n3985 , n3986 , n3987 , n3988 , n3989 , n3990 , n3991 , n3992 , n3993 , n3994 , n3995 , n3996 , n3997 , n3998 , n3999 , n4000 , n4001 , n4002 , n4003 , n4004 , n4005 , n4006 , n4007 , n4008 , n4009 , n4010 , n4011 , n4012 , n4013 , n4014 , n4015 , n4016 , n4017 , n4018 , n4019 , n4020 , n4021 , n4022 , n4023 , n4024 , n4025 , n4026 , n4027 , n4028 , n4029 , n4030 , n4031 , n4032 , n4033 , n4034 , n4035 , n4036 , n4037 , n4038 , n4039 , n4040 , n4041 , n4042 , n4043 , n4044 , n4045 , n4046 , n4047 , n4048 , n4049 , n4050 , n4051 , n4052 , n4053 , n4054 , n4055 , n4056 , n4057 , n4058 , n4059 , n4060 , n4061 , n4062 , n4063 , n4064 , n4065 , n4066 , n4067 , n4068 , n4069 , n4070 , n4071 , n4072 , n4073 , n4074 , n4075 , n4076 , n4077 , n4078 , n4079 , n4080 , n4081 , n4082 , n4083 , n4084 , n4085 , n4086 , n4087 , n4088 , n4089 , n4090 , n4091 , n4092 , n4093 , n4094 , n4095 , n4096 , n4097 , n4098 , n4099 , n4100 , n4101 , n4102 , n4103 , n4104 , n4105 , n4106 , n4107 , n4108 , n4109 , n4110 , n4111 , n4112 , n4113 , n4114 , n4115 , n4116 , n4117 , n4118 , n4119 , n4120 , n4121 , n4122 , n4123 , n4124 , n4125 , n4126 , n4127 , n4128 , n4129 , n4130 , n4131 , n4132 , n4133 , n4134 , n4135 , n4136 , n4137 , n4138 , n4139 , n4140 , n4141 , n4142 , n4143 , n4144 , n4145 , n4146 , n4147 , n4148 , n4149 , n4150 , n4151 , n4152 , n4153 , n4154 , n4155 , n4156 , n4157 , n4158 , n4159 , n4160 , n4161 , n4162 , n4163 , n4164 , n4165 , n4166 , n4167 , n4168 , n4169 , n4170 , n4171 , n4172 , n4173 , n4174 , n4175 , n4176 , n4177 , n4178 , n4179 , n4180 , n4181 , n4182 , n4183 , n4184 , n4185 , n4186 , n4187 , n4188 , n4189 , n4190 , n4191 , n4192 , n4193 , n4194 , n4195 , n4196 , n4197 , n4198 , n4199 , n4200 , n4201 , n4202 , n4203 , n4204 , n4205 , n4206 , n4207 , n4208 , n4209 , n4210 , n4211 , n4212 , n4213 , n4214 , n4215 , n4216 , n4217 , n4218 , n4219 , n4220 , n4221 , n4222 , n4223 , n4224 , n4225 , n4226 , n4227 , n4228 , n4229 , n4230 , n4231 , n4232 , n4233 , n4234 , n4235 , n4236 , n4237 , n4238 , n4239 , n4240 , n4241 , n4242 , n4243 , n4244 , n4245 , n4246 , n4247 , n4248 , n4249 , n4250 , n4251 , n4252 , n4253 , n4254 , n4255 , n4256 , n4257 , n4258 , n4259 , n4260 , n4261 , n4262 , n4263 , n4264 , n4265 , n4266 , n4267 , n4268 , n4269 , n4270 , n4271 , n4272 , n4273 , n4274 , n4275 , n4276 , n4277 , n4278 , n4279 , n4280 , n4281 , n4282 , n4283 , n4284 , n4285 , n4286 , n4287 , n4288 , n4289 , n4290 , n4291 , n4292 , n4293 , n4294 , n4295 , n4296 , n4297 , n4298 , n4299 , n4300 , n4301 , n4302 , n4303 , n4304 , n4305 , n4306 , n4307 , n4308 , n4309 , n4310 , n4311 , n4312 , n4313 , n4314 , n4315 , n4316 , n4317 , n4318 , n4319 , n4320 , n4321 , n4322 , n4323 , n4324 , n4325 , n4326 , n4327 , n4328 , n4329 , n4330 , n4331 , n4332 , n4333 , n4334 , n4335 , n4336 , n4337 , n4338 , n4339 , n4340 , n4341 , n4342 , n4343 , n4344 , n4345 , n4346 , n4347 , n4348 , n4349 , n4350 , n4351 , n4352 , n4353 , n4354 , n4355 , n4356 , n4357 , n4358 , n4359 , n4360 , n4361 , n4362 , n4363 , n4364 , n4365 , n4366 , n4367 , n4368 , n4369 , n4370 , n4371 , n4372 , n4373 , n4374 , n4375 , n4376 , n4377 , n4378 , n4379 , n4380 , n4381 , n4382 , n4383 , n4384 , n4385 , n4386 , n4387 , n4388 , n4389 , n4390 , n4391 , n4392 , n4393 , n4394 , n4395 , n4396 , n4397 , n4398 , n4399 , n4400 , n4401 , n4402 , n4403 , n4404 , n4405 , n4406 , n4407 , n4408 , n4409 , n4410 , n4411 , n4412 , n4413 , n4414 , n4415 , n4416 , n4417 , n4418 , n4419 , n4420 , n4421 , n4422 , n4423 , n4424 , n4425 , n4426 , n4427 , n4428 , n4429 , n4430 , n4431 , n4432 , n4433 , n4434 , n4435 , n4436 , n4437 , n4438 , n4439 , n4440 , n4441 , n4442 , n4443 , n4444 , n4445 , n4446 , n4447 , n4448 , n4449 , n4450 , n4451 , n4452 , n4453 , n4454 , n4455 , n4456 , n4457 , n4458 , n4459 , n4460 , n4461 , n4462 , n4463 , n4464 , n4465 , n4466 , n4467 , n4468 , n4469 , n4470 , n4471 , n4472 , n4473 , n4474 , n4475 , n4476 , n4477 , n4478 , n4479 , n4480 , n4481 , n4482 , n4483 , n4484 , n4485 , n4486 , n4487 , n4488 , n4489 , n4490 , n4491 , n4492 , n4493 , n4494 , n4495 , n4496 , n4497 , n4498 , n4499 , n4500 , n4501 , n4502 , n4503 , n4504 , n4505 , n4506 , n4507 , n4508 , n4509 , n4510 , n4511 , n4512 , n4513 , n4514 , n4515 , n4516 , n4517 , n4518 , n4519 , n4520 , n4521 , n4522 , n4523 , n4524 , n4525 , n4526 , n4527 , n4528 , n4529 , n4530 , n4531 , n4532 , n4533 , n4534 , n4535 , n4536 , n4537 , n4538 , n4539 , n4540 , n4541 , n4542 , n4543 , n4544 , n4545 , n4546 , n4547 , n4548 , n4549 , n4550 , n4551 , n4552 , n4553 , n4554 , n4555 , n4556 , n4557 , n4558 , n4559 , n4560 , n4561 , n4562 , n4563 , n4564 , n4565 , n4566 , n4567 , n4568 , n4569 , n4570 , n4571 , n4572 , n4573 , n4574 , n4575 , n4576 , n4577 , n4578 , n4579 , n4580 , n4581 , n4582 , n4583 , n4584 , n4585 , n4586 , n4587 , n4588 , n4589 , n4590 , n4591 , n4592 , n4593 , n4594 , n4595 , n4596 , n4597 , n4598 , n4599 , n4600 , n4601 , n4602 , n4603 , n4604 , n4605 , n4606 , n4607 , n4608 , n4609 , n4610 , n4611 , n4612 , n4613 , n4614 , n4615 , n4616 , n4617 , n4618 , n4619 , n4620 , n4621 , n4622 , n4623 , n4624 , n4625 , n4626 , n4627 , n4628 , n4629 , n4630 , n4631 , n4632 , n4633 , n4634 , n4635 , n4636 , n4637 , n4638 , n4639 , n4640 , n4641 , n4642 , n4643 , n4644 , n4645 , n4646 , n4647 , n4648 , n4649 , n4650 , n4651 , n4652 , n4653 , n4654 , n4655 , n4656 , n4657 , n4658 , n4659 , n4660 , n4661 , n4662 , n4663 , n4664 , n4665 , n4666 , n4667 , n4668 , n4669 , n4670 , n4671 , n4672 , n4673 , n4674 , n4675 , n4676 , n4677 , n4678 , n4679 , n4680 , n4681 , n4682 , n4683 , n4684 , n4685 , n4686 , n4687 , n4688 , n4689 , n4690 , n4691 , n4692 , n4693 , n4694 , n4695 , n4696 , n4697 , n4698 , n4699 , n4700 , n4701 , n4702 , n4703 , n4704 , n4705 , n4706 , n4707 , n4708 , n4709 , n4710 , n4711 , n4712 , n4713 , n4714 , n4715 , n4716 , n4717 , n4718 , n4719 , n4720 , n4721 , n4722 , n4723 , n4724 , n4725 , n4726 , n4727 , n4728 , n4729 , n4730 , n4731 , n4732 , n4733 , n4734 , n4735 , n4736 , n4737 , n4738 , n4739 , n4740 , n4741 , n4742 , n4743 , n4744 , n4745 , n4746 , n4747 , n4748 , n4749 , n4750 , n4751 , n4752 , n4753 , n4754 , n4755 , n4756 , n4757 , n4758 , n4759 , n4760 , n4761 , n4762 , n4763 , n4764 , n4765 , n4766 , n4767 , n4768 , n4769 , n4770 , n4771 , n4772 , n4773 , n4774 , n4775 , n4776 , n4777 , n4778 , n4779 , n4780 , n4781 , n4782 , n4783 , n4784 , n4785 , n4786 , n4787 , n4788 , n4789 , n4790 , n4791 , n4792 , n4793 , n4794 , n4795 , n4796 , n4797 , n4798 , n4799 , n4800 , n4801 , n4802 , n4803 , n4804 , n4805 , n4806 , n4807 , n4808 , n4809 , n4810 , n4811 , n4812 , n4813 , n4814 , n4815 , n4816 , n4817 , n4818 , n4819 , n4820 , n4821 , n4822 , n4823 , n4824 , n4825 , n4826 , n4827 , n4828 , n4829 , n4830 , n4831 , n4832 , n4833 , n4834 , n4835 , n4836 , n4837 , n4838 , n4839 , n4840 , n4841 , n4842 , n4843 , n4844 , n4845 , n4846 , n4847 , n4848 , n4849 , n4850 , n4851 , n4852 , n4853 , n4854 , n4855 , n4856 , n4857 , n4858 , n4859 , n4860 , n4861 , n4862 , n4863 , n4864 , n4865 , n4866 , n4867 , n4868 , n4869 , n4870 , n4871 , n4872 , n4873 , n4874 , n4875 , n4876 , n4877 , n4878 , n4879 , n4880 , n4881 , n4882 , n4883 , n4884 , n4885 , n4886 , n4887 , n4888 , n4889 , n4890 , n4891 , n4892 , n4893 , n4894 , n4895 , n4896 , n4897 , n4898 , n4899 , n4900 , n4901 , n4902 , n4903 , n4904 , n4905 , n4906 , n4907 , n4908 , n4909 , n4910 , n4911 , n4912 , n4913 , n4914 , n4915 , n4916 , n4917 , n4918 , n4919 , n4920 , n4921 , n4922 , n4923 , n4924 , n4925 , n4926 , n4927 , n4928 , n4929 , n4930 , n4931 , n4932 , n4933 , n4934 , n4935 , n4936 , n4937 , n4938 , n4939 , n4940 , n4941 , n4942 , n4943 , n4944 , n4945 , n4946 , n4947 , n4948 , n4949 , n4950 , n4951 , n4952 , n4953 , n4954 , n4955 , n4956 , n4957 , n4958 , n4959 , n4960 , n4961 , n4962 , n4963 , n4964 , n4965 , n4966 , n4967 , n4968 , n4969 , n4970 , n4971 , n4972 , n4973 , n4974 , n4975 , n4976 , n4977 , n4978 , n4979 , n4980 , n4981 , n4982 , n4983 , n4984 , n4985 , n4986 , n4987 , n4988 , n4989 , n4990 , n4991 , n4992 , n4993 , n4994 , n4995 , n4996 , n4997 , n4998 , n4999 , n5000 , n5001 , n5002 , n5003 , n5004 , n5005 , n5006 , n5007 , n5008 , n5009 , n5010 , n5011 , n5012 , n5013 , n5014 , n5015 , n5016 , n5017 , n5018 , n5019 , n5020 , n5021 , n5022 , n5023 , n5024 , n5025 , n5026 , n5027 , n5028 , n5029 , n5030 , n5031 , n5032 , n5033 , n5034 , n5035 , n5036 , n5037 , n5038 , n5039 , n5040 , n5041 , n5042 , n5043 , n5044 , n5045 , n5046 , n5047 , n5048 , n5049 , n5050 , n5051 , n5052 , n5053 , n5054 , n5055 , n5056 , n5057 , n5058 , n5059 , n5060 , n5061 , n5062 , n5063 , n5064 , n5065 , n5066 , n5067 , n5068 , n5069 , n5070 , n5071 , n5072 , n5073 , n5074 , n5075 , n5076 , n5077 , n5078 , n5079 , n5080 , n5081 , n5082 , n5083 , n5084 , n5085 , n5086 , n5087 , n5088 , n5089 , n5090 , n5091 , n5092 , n5093 , n5094 , n5095 , n5096 , n5097 , n5098 , n5099 , n5100 , n5101 , n5102 , n5103 , n5104 , n5105 , n5106 , n5107 , n5108 , n5109 , n5110 , n5111 , n5112 , n5113 , n5114 , n5115 , n5116 , n5117 , n5118 , n5119 , n5120 , n5121 , n5122 , n5123 , n5124 , n5125 , n5126 , n5127 , n5128 , n5129 , n5130 , n5131 , n5132 , n5133 , n5134 , n5135 , n5136 , n5137 , n5138 , n5139 , n5140 , n5141 , n5142 , n5143 , n5144 , n5145 , n5146 , n5147 , n5148 , n5149 , n5150 , n5151 , n5152 , n5153 , n5154 , n5155 , n5156 , n5157 , n5158 , n5159 , n5160 , n5161 , n5162 , n5163 , n5164 , n5165 , n5166 , n5167 , n5168 , n5169 , n5170 , n5171 , n5172 , n5173 , n5174 , n5175 , n5176 , n5177 , n5178 , n5179 , n5180 , n5181 , n5182 , n5183 , n5184 , n5185 , n5186 , n5187 , n5188 , n5189 , n5190 , n5191 , n5192 , n5193 , n5194 , n5195 , n5196 , n5197 , n5198 , n5199 , n5200 , n5201 , n5202 , n5203 , n5204 , n5205 , n5206 , n5207 , n5208 , n5209 , n5210 , n5211 , n5212 , n5213 , n5214 , n5215 , n5216 , n5217 , n5218 , n5219 , n5220 , n5221 , n5222 , n5223 , n5224 , n5225 , n5226 , n5227 , n5228 , n5229 , n5230 , n5231 , n5232 , n5233 , n5234 , n5235 , n5236 , n5237 , n5238 , n5239 , n5240 , n5241 , n5242 , n5243 , n5244 , n5245 , n5246 , n5247 , n5248 , n5249 , n5250 , n5251 , n5252 , n5253 , n5254 , n5255 , n5256 , n5257 , n5258 , n5259 , n5260 , n5261 , n5262 , n5263 , n5264 , n5265 , n5266 , n5267 , n5268 , n5269 , n5270 , n5271 , n5272 , n5273 , n5274 , n5275 , n5276 , n5277 , n5278 , n5279 , n5280 , n5281 , n5282 , n5283 , n5284 , n5285 , n5286 , n5287 , n5288 , n5289 , n5290 , n5291 , n5292 , n5293 , n5294 , n5295 , n5296 , n5297 , n5298 , n5299 , n5300 , n5301 , n5302 , n5303 , n5304 , n5305 , n5306 , n5307 , n5308 , n5309 , n5310 , n5311 , n5312 , n5313 , n5314 , n5315 , n5316 , n5317 , n5318 , n5319 , n5320 , n5321 , n5322 , n5323 , n5324 , n5325 , n5326 , n5327 , n5328 , n5329 , n5330 , n5331 , n5332 , n5333 , n5334 , n5335 , n5336 , n5337 , n5338 , n5339 , n5340 , n5341 , n5342 , n5343 , n5344 , n5345 , n5346 , n5347 , n5348 , n5349 , n5350 , n5351 , n5352 , n5353 , n5354 , n5355 , n5356 , n5357 , n5358 , n5359 , n5360 , n5361 , n5362 , n5363 , n5364 , n5365 , n5366 , n5367 , n5368 , n5369 , n5370 , n5371 , n5372 , n5373 , n5374 , n5375 , n5376 , n5377 , n5378 , n5379 , n5380 , n5381 , n5382 , n5383 , n5384 , n5385 , n5386 , n5387 , n5388 , n5389 , n5390 , n5391 , n5392 , n5393 , n5394 , n5395 , n5396 , n5397 , n5398 , n5399 , n5400 , n5401 , n5402 , n5403 , n5404 , n5405 , n5406 , n5407 , n5408 , n5409 , n5410 , n5411 , n5412 , n5413 , n5414 , n5415 , n5416 , n5417 , n5418 , n5419 , n5420 , n5421 , n5422 , n5423 , n5424 , n5425 , n5426 , n5427 , n5428 , n5429 , n5430 , n5431 , n5432 , n5433 , n5434 , n5435 , n5436 , n5437 , n5438 , n5439 , n5440 , n5441 , n5442 , n5443 , n5444 , n5445 , n5446 , n5447 , n5448 , n5449 , n5450 , n5451 , n5452 , n5453 , n5454 , n5455 , n5456 , n5457 , n5458 , n5459 , n5460 , n5461 , n5462 , n5463 , n5464 , n5465 , n5466 , n5467 , n5468 , n5469 , n5470 , n5471 , n5472 , n5473 , n5474 , n5475 , n5476 , n5477 , n5478 , n5479 , n5480 , n5481 , n5482 , n5483 , n5484 , n5485 , n5486 , n5487 , n5488 , n5489 , n5490 , n5491 , n5492 , n5493 , n5494 , n5495 , n5496 , n5497 , n5498 , n5499 , n5500 , n5501 , n5502 , n5503 , n5504 , n5505 , n5506 , n5507 , n5508 , n5509 , n5510 , n5511 , n5512 , n5513 , n5514 , n5515 , n5516 , n5517 , n5518 , n5519 , n5520 , n5521 , n5522 , n5523 , n5524 , n5525 , n5526 , n5527 , n5528 , n5529 , n5530 , n5531 , n5532 , n5533 , n5534 , n5535 , n5536 , n5537 , n5538 , n5539 , n5540 , n5541 , n5542 , n5543 , n5544 , n5545 , n5546 , n5547 , n5548 , n5549 , n5550 , n5551 , n5552 , n5553 , n5554 , n5555 , n5556 , n5557 , n5558 , n5559 , n5560 , n5561 , n5562 , n5563 , n5564 , n5565 , n5566 , n5567 , n5568 , n5569 , n5570 , n5571 , n5572 , n5573 , n5574 , n5575 , n5576 , n5577 , n5578 , n5579 , n5580 , n5581 , n5582 , n5583 , n5584 , n5585 , n5586 , n5587 , n5588 , n5589 , n5590 , n5591 , n5592 , n5593 , n5594 , n5595 , n5596 , n5597 , n5598 , n5599 , n5600 , n5601 , n5602 , n5603 , n5604 , n5605 , n5606 , n5607 , n5608 , n5609 , n5610 , n5611 , n5612 , n5613 , n5614 , n5615 , n5616 , n5617 , n5618 , n5619 , n5620 , n5621 , n5622 , n5623 , n5624 , n5625 , n5626 , n5627 , n5628 , n5629 , n5630 , n5631 , n5632 , n5633 , n5634 , n5635 , n5636 , n5637 , n5638 , n5639 , n5640 , n5641 , n5642 , n5643 , n5644 , n5645 , n5646 , n5647 , n5648 , n5649 , n5650 , n5651 , n5652 , n5653 , n5654 , n5655 , n5656 , n5657 , n5658 , n5659 , n5660 , n5661 , n5662 , n5663 , n5664 , n5665 , n5666 , n5667 , n5668 , n5669 , n5670 , n5671 , n5672 , n5673 , n5674 , n5675 , n5676 , n5677 , n5678 , n5679 , n5680 , n5681 , n5682 , n5683 , n5684 , n5685 , n5686 , n5687 , n5688 , n5689 , n5690 , n5691 , n5692 , n5693 , n5694 , n5695 , n5696 , n5697 , n5698 , n5699 , n5700 , n5701 , n5702 , n5703 , n5704 , n5705 , n5706 , n5707 , n5708 , n5709 , n5710 , n5711 , n5712 , n5713 , n5714 , n5715 , n5716 , n5717 , n5718 , n5719 , n5720 , n5721 , n5722 , n5723 , n5724 , n5725 , n5726 , n5727 , n5728 , n5729 , n5730 , n5731 , n5732 , n5733 , n5734 , n5735 , n5736 , n5737 , n5738 , n5739 , n5740 , n5741 , n5742 , n5743 , n5744 , n5745 , n5746 , n5747 , n5748 , n5749 , n5750 , n5751 , n5752 , n5753 , n5754 , n5755 , n5756 , n5757 , n5758 , n5759 , n5760 , n5761 , n5762 , n5763 , n5764 , n5765 , n5766 , n5767 , n5768 , n5769 , n5770 , n5771 , n5772 , n5773 , n5774 , n5775 , n5776 , n5777 , n5778 , n5779 , n5780 , n5781 , n5782 , n5783 , n5784 , n5785 , n5786 , n5787 , n5788 , n5789 , n5790 , n5791 , n5792 , n5793 , n5794 , n5795 , n5796 , n5797 , n5798 , n5799 , n5800 , n5801 , n5802 , n5803 , n5804 , n5805 , n5806 , n5807 , n5808 , n5809 , n5810 , n5811 , n5812 , n5813 , n5814 , n5815 , n5816 , n5817 , n5818 , n5819 , n5820 , n5821 , n5822 , n5823 , n5824 , n5825 , n5826 , n5827 , n5828 , n5829 , n5830 , n5831 , n5832 , n5833 , n5834 , n5835 , n5836 , n5837 , n5838 , n5839 , n5840 , n5841 , n5842 , n5843 , n5844 , n5845 , n5846 , n5847 , n5848 , n5849 , n5850 , n5851 , n5852 , n5853 , n5854 , n5855 , n5856 , n5857 , n5858 , n5859 , n5860 , n5861 , n5862 , n5863 , n5864 , n5865 , n5866 , n5867 , n5868 , n5869 , n5870 , n5871 , n5872 , n5873 , n5874 , n5875 , n5876 , n5877 , n5878 , n5879 , n5880 , n5881 , n5882 , n5883 , n5884 , n5885 , n5886 , n5887 , n5888 , n5889 , n5890 , n5891 , n5892 , n5893 , n5894 , n5895 , n5896 , n5897 , n5898 , n5899 , n5900 , n5901 , n5902 , n5903 , n5904 , n5905 , n5906 , n5907 , n5908 , n5909 , n5910 , n5911 , n5912 , n5913 , n5914 , n5915 , n5916 , n5917 , n5918 , n5919 , n5920 , n5921 , n5922 , n5923 , n5924 , n5925 , n5926 , n5927 , n5928 , n5929 , n5930 , n5931 , n5932 , n5933 , n5934 , n5935 , n5936 , n5937 , n5938 , n5939 , n5940 , n5941 , n5942 , n5943 , n5944 , n5945 , n5946 , n5947 , n5948 , n5949 , n5950 , n5951 , n5952 , n5953 , n5954 , n5955 , n5956 , n5957 , n5958 , n5959 , n5960 , n5961 , n5962 , n5963 , n5964 , n5965 , n5966 , n5967 , n5968 , n5969 , n5970 , n5971 , n5972 , n5973 , n5974 , n5975 , n5976 , n5977 , n5978 , n5979 , n5980 , n5981 , n5982 , n5983 , n5984 , n5985 , n5986 , n5987 , n5988 , n5989 , n5990 , n5991 , n5992 , n5993 , n5994 , n5995 , n5996 , n5997 , n5998 , n5999 , n6000 , n6001 , n6002 , n6003 , n6004 , n6005 , n6006 , n6007 , n6008 , n6009 , n6010 , n6011 , n6012 , n6013 , n6014 , n6015 , n6016 , n6017 , n6018 , n6019 , n6020 , n6021 , n6022 , n6023 , n6024 , n6025 , n6026 , n6027 , n6028 , n6029 , n6030 , n6031 , n6032 , n6033 , n6034 , n6035 , n6036 , n6037 , n6038 , n6039 , n6040 , n6041 , n6042 , n6043 , n6044 , n6045 , n6046 , n6047 , n6048 , n6049 , n6050 , n6051 , n6052 , n6053 , n6054 , n6055 , n6056 , n6057 , n6058 , n6059 , n6060 , n6061 , n6062 , n6063 , n6064 , n6065 , n6066 , n6067 , n6068 , n6069 , n6070 , n6071 , n6072 , n6073 , n6074 , n6075 , n6076 , n6077 , n6078 , n6079 , n6080 , n6081 , n6082 , n6083 , n6084 , n6085 , n6086 , n6087 , n6088 , n6089 , n6090 , n6091 , n6092 , n6093 , n6094 , n6095 , n6096 , n6097 , n6098 , n6099 , n6100 , n6101 , n6102 , n6103 , n6104 , n6105 , n6106 , n6107 , n6108 , n6109 , n6110 , n6111 , n6112 , n6113 , n6114 , n6115 , n6116 , n6117 , n6118 , n6119 , n6120 , n6121 , n6122 , n6123 , n6124 , n6125 , n6126 , n6127 , n6128 , n6129 , n6130 , n6131 , n6132 , n6133 , n6134 , n6135 , n6136 , n6137 , n6138 , n6139 , n6140 , n6141 , n6142 , n6143 , n6144 , n6145 , n6146 , n6147 , n6148 , n6149 , n6150 , n6151 , n6152 , n6153 , n6154 , n6155 , n6156 , n6157 , n6158 , n6159 , n6160 , n6161 , n6162 , n6163 , n6164 , n6165 , n6166 , n6167 , n6168 , n6169 , n6170 , n6171 , n6172 , n6173 , n6174 , n6175 , n6176 , n6177 , n6178 , n6179 , n6180 , n6181 , n6182 , n6183 , n6184 , n6185 , n6186 , n6187 , n6188 , n6189 , n6190 , n6191 , n6192 , n6193 , n6194 , n6195 , n6196 , n6197 , n6198 , n6199 , n6200 , n6201 , n6202 , n6203 , n6204 , n6205 , n6206 , n6207 , n6208 , n6209 , n6210 , n6211 , n6212 , n6213 , n6214 , n6215 , n6216 , n6217 , n6218 , n6219 , n6220 , n6221 , n6222 , n6223 , n6224 , n6225 , n6226 , n6227 , n6228 , n6229 , n6230 , n6231 , n6232 , n6233 , n6234 , n6235 , n6236 , n6237 , n6238 , n6239 , n6240 , n6241 , n6242 , n6243 , n6244 , n6245 , n6246 , n6247 , n6248 , n6249 , n6250 , n6251 , n6252 , n6253 , n6254 , n6255 , n6256 , n6257 , n6258 , n6259 , n6260 , n6261 , n6262 , n6263 , n6264 , n6265 , n6266 , n6267 , n6268 , n6269 , n6270 , n6271 , n6272 , n6273 , n6274 , n6275 , n6276 , n6277 , n6278 , n6279 , n6280 , n6281 , n6282 , n6283 , n6284 , n6285 , n6286 , n6287 , n6288 , n6289 , n6290 , n6291 , n6292 , n6293 , n6294 , n6295 , n6296 , n6297 , n6298 , n6299 , n6300 , n6301 , n6302 , n6303 , n6304 , n6305 , n6306 , n6307 , n6308 , n6309 , n6310 , n6311 , n6312 , n6313 , n6314 , n6315 , n6316 , n6317 , n6318 , n6319 , n6320 , n6321 , n6322 , n6323 , n6324 , n6325 , n6326 , n6327 , n6328 , n6329 , n6330 , n6331 , n6332 , n6333 , n6334 , n6335 , n6336 , n6337 , n6338 , n6339 , n6340 , n6341 , n6342 , n6343 , n6344 , n6345 , n6346 , n6347 , n6348 , n6349 , n6350 , n6351 , n6352 , n6353 , n6354 , n6355 , n6356 , n6357 , n6358 , n6359 , n6360 , n6361 , n6362 , n6363 , n6364 , n6365 , n6366 , n6367 , n6368 , n6369 , n6370 , n6371 , n6372 , n6373 , n6374 , n6375 , n6376 , n6377 , n6378 , n6379 , n6380 , n6381 , n6382 , n6383 , n6384 , n6385 , n6386 , n6387 , n6388 , n6389 , n6390 , n6391 , n6392 , n6393 , n6394 , n6395 , n6396 , n6397 , n6398 , n6399 , n6400 , n6401 , n6402 , n6403 , n6404 , n6405 , n6406 , n6407 , n6408 , n6409 , n6410 , n6411 , n6412 , n6413 , n6414 , n6415 , n6416 , n6417 , n6418 , n6419 , n6420 , n6421 , n6422 , n6423 , n6424 , n6425 , n6426 , n6427 , n6428 , n6429 , n6430 , n6431 , n6432 , n6433 , n6434 , n6435 , n6436 , n6437 , n6438 , n6439 , n6440 , n6441 , n6442 , n6443 , n6444 , n6445 , n6446 , n6447 , n6448 , n6449 , n6450 , n6451 , n6452 , n6453 , n6454 , n6455 , n6456 , n6457 , n6458 , n6459 , n6460 , n6461 , n6462 , n6463 , n6464 , n6465 , n6466 , n6467 , n6468 , n6469 , n6470 , n6471 , n6472 , n6473 , n6474 , n6475 , n6476 , n6477 , n6478 , n6479 , n6480 , n6481 , n6482 , n6483 , n6484 , n6485 , n6486 , n6487 , n6488 , n6489 , n6490 , n6491 , n6492 , n6493 , n6494 , n6495 , n6496 , n6497 , n6498 , n6499 , n6500 , n6501 , n6502 , n6503 , n6504 , n6505 , n6506 , n6507 , n6508 , n6509 , n6510 , n6511 , n6512 , n6513 , n6514 , n6515 , n6516 , n6517 , n6518 , n6519 , n6520 , n6521 , n6522 , n6523 , n6524 , n6525 , n6526 , n6527 , n6528 , n6529 , n6530 , n6531 , n6532 , n6533 , n6534 , n6535 , n6536 , n6537 , n6538 , n6539 , n6540 , n6541 , n6542 , n6543 , n6544 , n6545 , n6546 , n6547 , n6548 , n6549 , n6550 , n6551 , n6552 , n6553 , n6554 , n6555 , n6556 , n6557 , n6558 , n6559 , n6560 , n6561 , n6562 , n6563 , n6564 , n6565 , n6566 , n6567 , n6568 , n6569 , n6570 , n6571 , n6572 , n6573 , n6574 , n6575 , n6576 , n6577 , n6578 , n6579 , n6580 , n6581 , n6582 , n6583 , n6584 , n6585 , n6586 , n6587 , n6588 , n6589 , n6590 , n6591 , n6592 , n6593 , n6594 , n6595 , n6596 , n6597 , n6598 , n6599 , n6600 , n6601 , n6602 , n6603 , n6604 , n6605 , n6606 , n6607 , n6608 , n6609 , n6610 , n6611 , n6612 , n6613 , n6614 , n6615 , n6616 , n6617 , n6618 , n6619 , n6620 , n6621 , n6622 , n6623 , n6624 , n6625 , n6626 , n6627 , n6628 , n6629 , n6630 , n6631 , n6632 , n6633 , n6634 , n6635 , n6636 , n6637 , n6638 , n6639 , n6640 , n6641 , n6642 , n6643 , n6644 , n6645 , n6646 , n6647 , n6648 , n6649 , n6650 , n6651 , n6652 , n6653 , n6654 , n6655 , n6656 , n6657 , n6658 , n6659 , n6660 , n6661 , n6662 , n6663 , n6664 , n6665 , n6666 , n6667 , n6668 , n6669 , n6670 , n6671 , n6672 , n6673 , n6674 , n6675 , n6676 , n6677 , n6678 , n6679 , n6680 , n6681 , n6682 , n6683 , n6684 , n6685 , n6686 , n6687 , n6688 , n6689 , n6690 , n6691 , n6692 , n6693 , n6694 , n6695 , n6696 , n6697 , n6698 , n6699 , n6700 , n6701 , n6702 , n6703 , n6704 , n6705 , n6706 , n6707 , n6708 , n6709 , n6710 , n6711 , n6712 , n6713 , n6714 , n6715 , n6716 , n6717 , n6718 , n6719 , n6720 , n6721 , n6722 , n6723 , n6724 , n6725 , n6726 , n6727 , n6728 , n6729 , n6730 , n6731 , n6732 , n6733 , n6734 , n6735 , n6736 , n6737 , n6738 , n6739 , n6740 , n6741 , n6742 , n6743 , n6744 , n6745 , n6746 , n6747 , n6748 , n6749 , n6750 , n6751 , n6752 , n6753 , n6754 , n6755 , n6756 , n6757 , n6758 , n6759 , n6760 , n6761 , n6762 , n6763 , n6764 , n6765 , n6766 , n6767 , n6768 , n6769 , n6770 , n6771 , n6772 , n6773 , n6774 , n6775 , n6776 , n6777 , n6778 , n6779 , n6780 , n6781 , n6782 , n6783 , n6784 , n6785 , n6786 , n6787 , n6788 , n6789 , n6790 , n6791 , n6792 , n6793 , n6794 , n6795 , n6796 , n6797 , n6798 , n6799 , n6800 , n6801 , n6802 , n6803 , n6804 , n6805 , n6806 , n6807 , n6808 , n6809 , n6810 , n6811 , n6812 , n6813 , n6814 , n6815 , n6816 , n6817 , n6818 , n6819 , n6820 , n6821 , n6822 , n6823 , n6824 , n6825 , n6826 , n6827 , n6828 , n6829 , n6830 , n6831 , n6832 , n6833 , n6834 , n6835 , n6836 , n6837 , n6838 , n6839 , n6840 , n6841 , n6842 , n6843 , n6844 , n6845 , n6846 , n6847 , n6848 , n6849 , n6850 , n6851 , n6852 , n6853 , n6854 , n6855 , n6856 , n6857 , n6858 , n6859 , n6860 , n6861 , n6862 , n6863 , n6864 , n6865 , n6866 , n6867 , n6868 , n6869 , n6870 , n6871 , n6872 , n6873 , n6874 , n6875 , n6876 , n6877 , n6878 , n6879 , n6880 , n6881 , n6882 , n6883 , n6884 , n6885 , n6886 , n6887 , n6888 , n6889 , n6890 , n6891 , n6892 , n6893 , n6894 , n6895 , n6896 , n6897 , n6898 , n6899 , n6900 , n6901 , n6902 , n6903 , n6904 , n6905 , n6906 , n6907 , n6908 , n6909 , n6910 , n6911 , n6912 , n6913 , n6914 , n6915 , n6916 , n6917 , n6918 , n6919 , n6920 , n6921 , n6922 , n6923 , n6924 , n6925 , n6926 , n6927 , n6928 , n6929 , n6930 , n6931 , n6932 , n6933 , n6934 , n6935 , n6936 , n6937 , n6938 , n6939 , n6940 , n6941 , n6942 , n6943 , n6944 , n6945 , n6946 , n6947 , n6948 , n6949 , n6950 , n6951 , n6952 , n6953 , n6954 , n6955 , n6956 , n6957 , n6958 , n6959 , n6960 , n6961 , n6962 , n6963 , n6964 , n6965 , n6966 , n6967 , n6968 , n6969 , n6970 , n6971 , n6972 , n6973 , n6974 , n6975 , n6976 , n6977 , n6978 , n6979 , n6980 , n6981 , n6982 , n6983 , n6984 , n6985 , n6986 , n6987 , n6988 , n6989 , n6990 , n6991 , n6992 , n6993 , n6994 , n6995 , n6996 , n6997 , n6998 , n6999 , n7000 , n7001 , n7002 , n7003 , n7004 , n7005 , n7006 , n7007 , n7008 , n7009 , n7010 , n7011 , n7012 , n7013 , n7014 , n7015 , n7016 , n7017 , n7018 , n7019 , n7020 , n7021 , n7022 , n7023 , n7024 , n7025 , n7026 , n7027 , n7028 , n7029 , n7030 , n7031 , n7032 , n7033 , n7034 , n7035 , n7036 , n7037 , n7038 , n7039 , n7040 , n7041 , n7042 , n7043 , n7044 , n7045 , n7046 , n7047 , n7048 , n7049 , n7050 , n7051 , n7052 , n7053 , n7054 , n7055 , n7056 , n7057 , n7058 , n7059 , n7060 , n7061 , n7062 , n7063 , n7064 , n7065 , n7066 , n7067 , n7068 , n7069 , n7070 , n7071 , n7072 , n7073 , n7074 , n7075 , n7076 , n7077 , n7078 , n7079 , n7080 , n7081 , n7082 , n7083 , n7084 , n7085 , n7086 , n7087 , n7088 , n7089 , n7090 , n7091 , n7092 , n7093 , n7094 , n7095 , n7096 , n7097 , n7098 , n7099 , n7100 , n7101 , n7102 , n7103 , n7104 , n7105 , n7106 , n7107 , n7108 , n7109 , n7110 , n7111 , n7112 , n7113 , n7114 , n7115 , n7116 , n7117 , n7118 , n7119 , n7120 , n7121 , n7122 , n7123 , n7124 , n7125 , n7126 , n7127 , n7128 , n7129 , n7130 , n7131 , n7132 , n7133 , n7134 , n7135 , n7136 , n7137 , n7138 , n7139 , n7140 , n7141 , n7142 , n7143 , n7144 , n7145 , n7146 , n7147 , n7148 , n7149 , n7150 , n7151 , n7152 , n7153 , n7154 , n7155 , n7156 , n7157 , n7158 , n7159 , n7160 , n7161 , n7162 , n7163 , n7164 , n7165 , n7166 , n7167 , n7168 , n7169 , n7170 , n7171 , n7172 , n7173 , n7174 , n7175 , n7176 , n7177 , n7178 , n7179 , n7180 , n7181 , n7182 , n7183 , n7184 , n7185 , n7186 , n7187 , n7188 , n7189 , n7190 , n7191 , n7192 , n7193 , n7194 , n7195 , n7196 , n7197 , n7198 , n7199 , n7200 , n7201 , n7202 , n7203 , n7204 , n7205 , n7206 , n7207 , n7208 , n7209 , n7210 , n7211 , n7212 , n7213 , n7214 , n7215 , n7216 , n7217 , n7218 , n7219 , n7220 , n7221 , n7222 , n7223 , n7224 , n7225 , n7226 , n7227 , n7228 , n7229 , n7230 , n7231 , n7232 , n7233 , n7234 , n7235 , n7236 , n7237 , n7238 , n7239 , n7240 , n7241 , n7242 , n7243 , n7244 , n7245 , n7246 , n7247 , n7248 , n7249 , n7250 , n7251 , n7252 , n7253 , n7254 , n7255 , n7256 , n7257 , n7258 , n7259 , n7260 , n7261 , n7262 , n7263 , n7264 , n7265 , n7266 , n7267 , n7268 , n7269 , n7270 , n7271 , n7272 , n7273 , n7274 , n7275 , n7276 , n7277 , n7278 , n7279 , n7280 , n7281 , n7282 , n7283 , n7284 , n7285 , n7286 , n7287 , n7288 , n7289 , n7290 , n7291 , n7292 , n7293 , n7294 , n7295 , n7296 , n7297 , n7298 , n7299 , n7300 , n7301 , n7302 , n7303 , n7304 , n7305 , n7306 , n7307 , n7308 , n7309 , n7310 , n7311 , n7312 , n7313 , n7314 , n7315 , n7316 , n7317 , n7318 , n7319 , n7320 , n7321 , n7322 , n7323 , n7324 , n7325 , n7326 , n7327 , n7328 , n7329 , n7330 , n7331 , n7332 , n7333 , n7334 , n7335 , n7336 , n7337 , n7338 , n7339 , n7340 , n7341 , n7342 , n7343 , n7344 , n7345 , n7346 , n7347 , n7348 , n7349 , n7350 , n7351 , n7352 , n7353 , n7354 , n7355 , n7356 , n7357 , n7358 , n7359 , n7360 , n7361 , n7362 , n7363 , n7364 , n7365 , n7366 , n7367 , n7368 , n7369 , n7370 , n7371 , n7372 , n7373 , n7374 , n7375 , n7376 , n7377 , n7378 , n7379 , n7380 , n7381 , n7382 , n7383 , n7384 , n7385 , n7386 , n7387 , n7388 , n7389 , n7390 , n7391 , n7392 , n7393 , n7394 , n7395 , n7396 , n7397 , n7398 , n7399 , n7400 , n7401 , n7402 , n7403 , n7404 , n7405 , n7406 , n7407 , n7408 , n7409 , n7410 , n7411 , n7412 , n7413 , n7414 , n7415 , n7416 , n7417 , n7418 , n7419 , n7420 , n7421 , n7422 , n7423 , n7424 , n7425 , n7426 , n7427 , n7428 , n7429 , n7430 , n7431 , n7432 , n7433 , n7434 , n7435 , n7436 , n7437 , n7438 , n7439 , n7440 , n7441 , n7442 , n7443 , n7444 , n7445 , n7446 , n7447 , n7448 , n7449 , n7450 , n7451 , n7452 , n7453 , n7454 , n7455 , n7456 , n7457 , n7458 , n7459 , n7460 , n7461 , n7462 , n7463 , n7464 , n7465 , n7466 , n7467 , n7468 , n7469 , n7470 , n7471 , n7472 , n7473 , n7474 , n7475 , n7476 , n7477 , n7478 , n7479 , n7480 , n7481 , n7482 , n7483 , n7484 , n7485 , n7486 , n7487 , n7488 , n7489 , n7490 , n7491 , n7492 , n7493 , n7494 , n7495 , n7496 , n7497 , n7498 , n7499 , n7500 , n7501 , n7502 , n7503 , n7504 , n7505 , n7506 , n7507 , n7508 , n7509 , n7510 , n7511 , n7512 , n7513 , n7514 , n7515 , n7516 , n7517 , n7518 , n7519 , n7520 , n7521 , n7522 , n7523 , n7524 , n7525 , n7526 , n7527 , n7528 , n7529 , n7530 , n7531 , n7532 , n7533 , n7534 , n7535 , n7536 , n7537 , n7538 , n7539 , n7540 , n7541 , n7542 , n7543 , n7544 , n7545 , n7546 , n7547 , n7548 , n7549 , n7550 , n7551 , n7552 , n7553 , n7554 , n7555 , n7556 , n7557 , n7558 , n7559 , n7560 , n7561 , n7562 , n7563 , n7564 , n7565 , n7566 , n7567 , n7568 , n7569 , n7570 , n7571 , n7572 , n7573 , n7574 , n7575 , n7576 , n7577 , n7578 , n7579 , n7580 , n7581 , n7582 , n7583 , n7584 , n7585 , n7586 , n7587 , n7588 , n7589 , n7590 , n7591 , n7592 , n7593 , n7594 , n7595 , n7596 , n7597 , n7598 , n7599 , n7600 , n7601 , n7602 , n7603 , n7604 , n7605 , n7606 , n7607 , n7608 , n7609 , n7610 , n7611 , n7612 , n7613 , n7614 , n7615 , n7616 , n7617 , n7618 , n7619 , n7620 , n7621 , n7622 , n7623 , n7624 , n7625 , n7626 , n7627 , n7628 , n7629 , n7630 , n7631 , n7632 , n7633 , n7634 , n7635 , n7636 , n7637 , n7638 , n7639 , n7640 , n7641 , n7642 , n7643 , n7644 , n7645 , n7646 , n7647 , n7648 , n7649 , n7650 , n7651 , n7652 , n7653 , n7654 , n7655 , n7656 , n7657 , n7658 , n7659 , n7660 , n7661 , n7662 , n7663 , n7664 , n7665 , n7666 , n7667 , n7668 , n7669 , n7670 , n7671 , n7672 , n7673 , n7674 , n7675 , n7676 , n7677 , n7678 , n7679 , n7680 , n7681 , n7682 , n7683 , n7684 , n7685 , n7686 , n7687 , n7688 , n7689 , n7690 , n7691 , n7692 , n7693 , n7694 , n7695 , n7696 , n7697 , n7698 , n7699 , n7700 , n7701 , n7702 , n7703 , n7704 , n7705 , n7706 , n7707 , n7708 , n7709 , n7710 , n7711 , n7712 , n7713 , n7714 , n7715 , n7716 , n7717 , n7718 , n7719 , n7720 , n7721 , n7722 , n7723 , n7724 , n7725 , n7726 , n7727 , n7728 , n7729 , n7730 , n7731 , n7732 , n7733 , n7734 , n7735 , n7736 , n7737 , n7738 , n7739 , n7740 , n7741 , n7742 , n7743 , n7744 , n7745 , n7746 , n7747 , n7748 , n7749 , n7750 , n7751 , n7752 , n7753 , n7754 , n7755 , n7756 , n7757 , n7758 , n7759 , n7760 , n7761 , n7762 , n7763 , n7764 , n7765 , n7766 , n7767 , n7768 , n7769 , n7770 , n7771 , n7772 , n7773 , n7774 , n7775 , n7776 , n7777 , n7778 , n7779 , n7780 , n7781 , n7782 , n7783 , n7784 , n7785 , n7786 , n7787 , n7788 , n7789 , n7790 , n7791 , n7792 , n7793 , n7794 , n7795 , n7796 , n7797 , n7798 , n7799 , n7800 , n7801 , n7802 , n7803 , n7804 , n7805 , n7806 , n7807 , n7808 , n7809 , n7810 , n7811 , n7812 , n7813 , n7814 , n7815 , n7816 , n7817 , n7818 , n7819 , n7820 , n7821 , n7822 , n7823 , n7824 , n7825 , n7826 , n7827 , n7828 , n7829 , n7830 , n7831 , n7832 , n7833 , n7834 , n7835 , n7836 , n7837 , n7838 , n7839 , n7840 , n7841 , n7842 , n7843 , n7844 , n7845 , n7846 , n7847 , n7848 , n7849 , n7850 , n7851 , n7852 , n7853 , n7854 , n7855 , n7856 , n7857 , n7858 , n7859 , n7860 , n7861 , n7862 , n7863 , n7864 , n7865 , n7866 , n7867 , n7868 , n7869 , n7870 , n7871 , n7872 , n7873 , n7874 , n7875 , n7876 , n7877 , n7878 , n7879 , n7880 , n7881 , n7882 , n7883 , n7884 , n7885 , n7886 , n7887 , n7888 , n7889 , n7890 , n7891 , n7892 , n7893 , n7894 , n7895 , n7896 , n7897 , n7898 , n7899 , n7900 , n7901 , n7902 , n7903 , n7904 , n7905 , n7906 , n7907 , n7908 , n7909 , n7910 , n7911 , n7912 , n7913 , n7914 , n7915 , n7916 , n7917 , n7918 , n7919 , n7920 , n7921 , n7922 , n7923 , n7924 , n7925 , n7926 , n7927 , n7928 , n7929 , n7930 , n7931 , n7932 , n7933 , n7934 , n7935 , n7936 , n7937 , n7938 , n7939 , n7940 , n7941 , n7942 , n7943 , n7944 , n7945 , n7946 , n7947 , n7948 , n7949 , n7950 , n7951 , n7952 , n7953 , n7954 , n7955 , n7956 , n7957 , n7958 , n7959 , n7960 , n7961 , n7962 , n7963 , n7964 , n7965 , n7966 , n7967 , n7968 , n7969 , n7970 , n7971 , n7972 , n7973 , n7974 , n7975 , n7976 , n7977 , n7978 , n7979 , n7980 , n7981 , n7982 , n7983 , n7984 , n7985 , n7986 , n7987 , n7988 , n7989 , n7990 , n7991 , n7992 , n7993 , n7994 , n7995 , n7996 , n7997 , n7998 , n7999 , n8000 , n8001 , n8002 , n8003 , n8004 , n8005 , n8006 , n8007 , n8008 , n8009 , n8010 , n8011 , n8012 , n8013 , n8014 , n8015 , n8016 , n8017 , n8018 , n8019 , n8020 , n8021 , n8022 , n8023 , n8024 , n8025 , n8026 , n8027 , n8028 , n8029 , n8030 , n8031 , n8032 , n8033 , n8034 , n8035 , n8036 , n8037 , n8038 , n8039 , n8040 , n8041 , n8042 , n8043 , n8044 , n8045 , n8046 , n8047 , n8048 , n8049 , n8050 , n8051 , n8052 , n8053 , n8054 , n8055 , n8056 , n8057 , n8058 , n8059 , n8060 , n8061 , n8062 , n8063 , n8064 , n8065 , n8066 , n8067 , n8068 , n8069 , n8070 , n8071 , n8072 , n8073 , n8074 , n8075 , n8076 , n8077 , n8078 , n8079 , n8080 , n8081 , n8082 , n8083 , n8084 , n8085 , n8086 , n8087 , n8088 , n8089 , n8090 , n8091 , n8092 , n8093 , n8094 , n8095 , n8096 , n8097 , n8098 , n8099 , n8100 , n8101 , n8102 , n8103 , n8104 , n8105 , n8106 , n8107 , n8108 , n8109 , n8110 , n8111 , n8112 , n8113 , n8114 , n8115 , n8116 , n8117 , n8118 , n8119 , n8120 , n8121 , n8122 , n8123 , n8124 , n8125 , n8126 , n8127 , n8128 , n8129 , n8130 , n8131 , n8132 , n8133 , n8134 , n8135 , n8136 , n8137 , n8138 , n8139 , n8140 , n8141 , n8142 , n8143 , n8144 , n8145 , n8146 , n8147 , n8148 , n8149 , n8150 , n8151 , n8152 , n8153 , n8154 , n8155 , n8156 , n8157 , n8158 , n8159 , n8160 , n8161 , n8162 , n8163 , n8164 , n8165 , n8166 , n8167 , n8168 , n8169 , n8170 , n8171 , n8172 , n8173 , n8174 , n8175 , n8176 , n8177 , n8178 , n8179 , n8180 , n8181 , n8182 , n8183 , n8184 , n8185 , n8186 , n8187 , n8188 , n8189 , n8190 , n8191 , n8192 , n8193 , n8194 , n8195 , n8196 , n8197 , n8198 , n8199 , n8200 , n8201 , n8202 , n8203 , n8204 , n8205 , n8206 , n8207 , n8208 , n8209 , n8210 , n8211 , n8212 , n8213 , n8214 , n8215 , n8216 , n8217 , n8218 , n8219 , n8220 , n8221 , n8222 , n8223 , n8224 , n8225 , n8226 , n8227 , n8228 , n8229 , n8230 , n8231 , n8232 , n8233 , n8234 , n8235 , n8236 , n8237 , n8238 , n8239 , n8240 , n8241 , n8242 , n8243 , n8244 , n8245 , n8246 , n8247 , n8248 , n8249 , n8250 , n8251 , n8252 , n8253 , n8254 , n8255 , n8256 , n8257 , n8258 , n8259 , n8260 , n8261 , n8262 , n8263 , n8264 , n8265 , n8266 , n8267 , n8268 , n8269 , n8270 , n8271 , n8272 , n8273 , n8274 , n8275 , n8276 , n8277 , n8278 , n8279 , n8280 , n8281 , n8282 , n8283 , n8284 , n8285 , n8286 , n8287 , n8288 , n8289 , n8290 , n8291 , n8292 , n8293 , n8294 , n8295 , n8296 , n8297 , n8298 , n8299 , n8300 , n8301 , n8302 , n8303 , n8304 , n8305 , n8306 , n8307 , n8308 , n8309 , n8310 , n8311 , n8312 , n8313 , n8314 , n8315 , n8316 , n8317 , n8318 , n8319 , n8320 , n8321 , n8322 , n8323 , n8324 , n8325 , n8326 , n8327 , n8328 , n8329 , n8330 , n8331 , n8332 , n8333 , n8334 , n8335 , n8336 , n8337 , n8338 , n8339 , n8340 , n8341 , n8342 , n8343 , n8344 , n8345 , n8346 , n8347 , n8348 , n8349 , n8350 , n8351 , n8352 , n8353 , n8354 , n8355 , n8356 , n8357 , n8358 , n8359 , n8360 , n8361 , n8362 , n8363 , n8364 , n8365 , n8366 , n8367 , n8368 , n8369 , n8370 , n8371 , n8372 , n8373 , n8374 , n8375 , n8376 , n8377 , n8378 , n8379 , n8380 , n8381 , n8382 , n8383 , n8384 , n8385 , n8386 , n8387 , n8388 , n8389 , n8390 , n8391 , n8392 , n8393 , n8394 , n8395 , n8396 , n8397 , n8398 , n8399 , n8400 , n8401 , n8402 , n8403 , n8404 , n8405 , n8406 , n8407 , n8408 , n8409 , n8410 , n8411 , n8412 , n8413 , n8414 , n8415 , n8416 , n8417 , n8418 , n8419 , n8420 , n8421 , n8422 , n8423 , n8424 , n8425 , n8426 , n8427 , n8428 , n8429 , n8430 , n8431 , n8432 , n8433 , n8434 , n8435 , n8436 , n8437 , n8438 , n8439 , n8440 , n8441 , n8442 , n8443 , n8444 , n8445 , n8446 , n8447 , n8448 , n8449 , n8450 , n8451 , n8452 , n8453 , n8454 , n8455 , n8456 , n8457 , n8458 , n8459 , n8460 , n8461 , n8462 , n8463 , n8464 , n8465 , n8466 , n8467 , n8468 , n8469 , n8470 , n8471 , n8472 , n8473 , n8474 , n8475 , n8476 , n8477 , n8478 , n8479 , n8480 , n8481 , n8482 , n8483 , n8484 , n8485 , n8486 , n8487 , n8488 , n8489 , n8490 , n8491 , n8492 , n8493 , n8494 , n8495 , n8496 , n8497 , n8498 , n8499 , n8500 , n8501 , n8502 , n8503 , n8504 , n8505 , n8506 , n8507 , n8508 , n8509 , n8510 , n8511 , n8512 , n8513 , n8514 , n8515 , n8516 , n8517 , n8518 , n8519 , n8520 , n8521 , n8522 , n8523 , n8524 , n8525 , n8526 , n8527 , n8528 , n8529 , n8530 , n8531 , n8532 , n8533 , n8534 , n8535 , n8536 , n8537 , n8538 , n8539 , n8540 , n8541 , n8542 , n8543 , n8544 , n8545 , n8546 , n8547 , n8548 , n8549 , n8550 , n8551 , n8552 , n8553 , n8554 , n8555 , n8556 , n8557 , n8558 , n8559 , n8560 , n8561 , n8562 , n8563 , n8564 , n8565 , n8566 , n8567 , n8568 , n8569 , n8570 , n8571 , n8572 , n8573 , n8574 , n8575 , n8576 , n8577 , n8578 , n8579 , n8580 , n8581 , n8582 , n8583 , n8584 , n8585 , n8586 , n8587 , n8588 , n8589 , n8590 , n8591 , n8592 , n8593 , n8594 , n8595 , n8596 , n8597 , n8598 , n8599 , n8600 , n8601 , n8602 , n8603 , n8604 , n8605 , n8606 , n8607 , n8608 , n8609 , n8610 , n8611 , n8612 , n8613 , n8614 , n8615 , n8616 , n8617 , n8618 , n8619 , n8620 , n8621 , n8622 , n8623 , n8624 , n8625 , n8626 , n8627 , n8628 , n8629 , n8630 , n8631 , n8632 , n8633 , n8634 , n8635 , n8636 , n8637 , n8638 , n8639 , n8640 , n8641 , n8642 , n8643 , n8644 , n8645 , n8646 , n8647 , n8648 , n8649 , n8650 , n8651 , n8652 , n8653 , n8654 , n8655 , n8656 , n8657 , n8658 , n8659 , n8660 , n8661 , n8662 , n8663 , n8664 , n8665 , n8666 , n8667 , n8668 , n8669 , n8670 , n8671 , n8672 , n8673 , n8674 , n8675 , n8676 , n8677 , n8678 , n8679 , n8680 , n8681 , n8682 , n8683 , n8684 , n8685 , n8686 , n8687 , n8688 , n8689 , n8690 , n8691 , n8692 , n8693 , n8694 , n8695 , n8696 , n8697 , n8698 , n8699 , n8700 , n8701 , n8702 , n8703 , n8704 , n8705 , n8706 , n8707 , n8708 , n8709 , n8710 , n8711 , n8712 , n8713 , n8714 , n8715 , n8716 , n8717 , n8718 , n8719 , n8720 , n8721 , n8722 , n8723 , n8724 , n8725 , n8726 , n8727 , n8728 , n8729 , n8730 , n8731 , n8732 , n8733 , n8734 , n8735 , n8736 , n8737 , n8738 , n8739 , n8740 , n8741 , n8742 , n8743 , n8744 , n8745 , n8746 , n8747 , n8748 , n8749 , n8750 , n8751 , n8752 , n8753 , n8754 , n8755 , n8756 , n8757 , n8758 , n8759 , n8760 , n8761 , n8762 , n8763 , n8764 , n8765 , n8766 , n8767 , n8768 , n8769 , n8770 , n8771 , n8772 , n8773 , n8774 , n8775 , n8776 , n8777 , n8778 , n8779 , n8780 , n8781 , n8782 , n8783 , n8784 , n8785 , n8786 , n8787 , n8788 , n8789 , n8790 , n8791 , n8792 , n8793 , n8794 , n8795 , n8796 , n8797 , n8798 , n8799 , n8800 , n8801 , n8802 , n8803 , n8804 , n8805 , n8806 , n8807 , n8808 , n8809 , n8810 , n8811 , n8812 , n8813 , n8814 , n8815 , n8816 , n8817 , n8818 , n8819 , n8820 , n8821 , n8822 , n8823 , n8824 , n8825 , n8826 , n8827 , n8828 , n8829 , n8830 , n8831 , n8832 , n8833 , n8834 , n8835 , n8836 , n8837 , n8838 , n8839 , n8840 , n8841 , n8842 , n8843 , n8844 , n8845 , n8846 , n8847 , n8848 , n8849 , n8850 , n8851 , n8852 , n8853 , n8854 , n8855 , n8856 , n8857 , n8858 , n8859 , n8860 , n8861 , n8862 , n8863 , n8864 , n8865 , n8866 , n8867 , n8868 , n8869 , n8870 , n8871 , n8872 , n8873 , n8874 , n8875 , n8876 , n8877 , n8878 , n8879 , n8880 , n8881 , n8882 , n8883 , n8884 , n8885 , n8886 , n8887 , n8888 , n8889 , n8890 , n8891 , n8892 , n8893 , n8894 , n8895 , n8896 , n8897 , n8898 , n8899 , n8900 , n8901 , n8902 , n8903 , n8904 , n8905 , n8906 , n8907 , n8908 , n8909 , n8910 , n8911 , n8912 , n8913 , n8914 , n8915 , n8916 , n8917 , n8918 , n8919 , n8920 , n8921 , n8922 , n8923 , n8924 , n8925 , n8926 , n8927 , n8928 , n8929 , n8930 , n8931 , n8932 , n8933 , n8934 , n8935 , n8936 , n8937 , n8938 , n8939 , n8940 , n8941 , n8942 , n8943 , n8944 , n8945 , n8946 , n8947 , n8948 , n8949 , n8950 , n8951 , n8952 , n8953 , n8954 , n8955 , n8956 , n8957 , n8958 , n8959 , n8960 , n8961 , n8962 , n8963 , n8964 , n8965 , n8966 , n8967 , n8968 , n8969 , n8970 , n8971 , n8972 , n8973 , n8974 , n8975 , n8976 , n8977 , n8978 , n8979 , n8980 , n8981 , n8982 , n8983 , n8984 , n8985 , n8986 , n8987 , n8988 , n8989 , n8990 , n8991 , n8992 , n8993 , n8994 , n8995 , n8996 , n8997 , n8998 , n8999 , n9000 , n9001 , n9002 , n9003 , n9004 , n9005 , n9006 , n9007 , n9008 , n9009 , n9010 , n9011 , n9012 , n9013 , n9014 , n9015 , n9016 , n9017 , n9018 , n9019 , n9020 , n9021 , n9022 , n9023 , n9024 , n9025 , n9026 , n9027 , n9028 , n9029 , n9030 , n9031 , n9032 , n9033 , n9034 , n9035 , n9036 , n9037 , n9038 , n9039 , n9040 , n9041 , n9042 , n9043 , n9044 , n9045 , n9046 , n9047 , n9048 , n9049 , n9050 , n9051 , n9052 , n9053 , n9054 , n9055 , n9056 , n9057 , n9058 , n9059 , n9060 , n9061 , n9062 , n9063 , n9064 , n9065 , n9066 , n9067 , n9068 , n9069 , n9070 , n9071 , n9072 , n9073 , n9074 , n9075 , n9076 , n9077 , n9078 , n9079 , n9080 , n9081 , n9082 , n9083 , n9084 , n9085 , n9086 , n9087 , n9088 , n9089 , n9090 , n9091 , n9092 , n9093 , n9094 , n9095 , n9096 , n9097 , n9098 , n9099 , n9100 , n9101 , n9102 , n9103 , n9104 , n9105 , n9106 , n9107 , n9108 , n9109 , n9110 , n9111 , n9112 , n9113 , n9114 , n9115 , n9116 , n9117 , n9118 , n9119 , n9120 , n9121 , n9122 , n9123 , n9124 , n9125 , n9126 , n9127 , n9128 , n9129 , n9130 , n9131 , n9132 , n9133 , n9134 , n9135 , n9136 , n9137 , n9138 , n9139 , n9140 , n9141 , n9142 , n9143 , n9144 , n9145 , n9146 , n9147 , n9148 , n9149 , n9150 , n9151 , n9152 , n9153 , n9154 , n9155 , n9156 , n9157 , n9158 , n9159 , n9160 , n9161 , n9162 , n9163 , n9164 , n9165 , n9166 , n9167 , n9168 , n9169 , n9170 , n9171 , n9172 , n9173 , n9174 , n9175 , n9176 , n9177 , n9178 , n9179 , n9180 , n9181 , n9182 , n9183 , n9184 , n9185 , n9186 , n9187 , n9188 , n9189 , n9190 , n9191 , n9192 , n9193 , n9194 , n9195 , n9196 , n9197 , n9198 , n9199 , n9200 , n9201 , n9202 , n9203 , n9204 , n9205 , n9206 , n9207 , n9208 , n9209 , n9210 , n9211 , n9212 , n9213 , n9214 , n9215 , n9216 , n9217 , n9218 , n9219 , n9220 , n9221 , n9222 , n9223 , n9224 , n9225 , n9226 , n9227 , n9228 , n9229 , n9230 , n9231 , n9232 , n9233 , n9234 , n9235 , n9236 , n9237 , n9238 , n9239 , n9240 , n9241 , n9242 , n9243 , n9244 , n9245 , n9246 , n9247 , n9248 , n9249 , n9250 , n9251 , n9252 , n9253 , n9254 , n9255 , n9256 , n9257 , n9258 , n9259 , n9260 , n9261 , n9262 , n9263 , n9264 , n9265 , n9266 , n9267 , n9268 , n9269 , n9270 , n9271 , n9272 , n9273 , n9274 , n9275 , n9276 , n9277 , n9278 , n9279 , n9280 , n9281 , n9282 , n9283 , n9284 , n9285 , n9286 , n9287 , n9288 , n9289 , n9290 , n9291 , n9292 , n9293 , n9294 , n9295 , n9296 , n9297 , n9298 , n9299 , n9300 , n9301 , n9302 , n9303 , n9304 , n9305 , n9306 , n9307 , n9308 , n9309 , n9310 , n9311 , n9312 , n9313 , n9314 , n9315 , n9316 , n9317 , n9318 , n9319 , n9320 , n9321 , n9322 , n9323 , n9324 , n9325 , n9326 , n9327 , n9328 , n9329 , n9330 , n9331 , n9332 , n9333 , n9334 , n9335 , n9336 , n9337 , n9338 , n9339 , n9340 , n9341 , n9342 , n9343 , n9344 , n9345 , n9346 , n9347 , n9348 , n9349 , n9350 , n9351 , n9352 , n9353 , n9354 , n9355 , n9356 , n9357 , n9358 , n9359 , n9360 , n9361 , n9362 , n9363 , n9364 , n9365 , n9366 , n9367 , n9368 , n9369 , n9370 , n9371 , n9372 , n9373 , n9374 , n9375 , n9376 , n9377 , n9378 , n9379 , n9380 , n9381 , n9382 , n9383 , n9384 , n9385 , n9386 , n9387 , n9388 , n9389 , n9390 , n9391 , n9392 , n9393 , n9394 , n9395 , n9396 , n9397 , n9398 , n9399 , n9400 , n9401 , n9402 , n9403 , n9404 , n9405 , n9406 , n9407 , n9408 , n9409 , n9410 , n9411 , n9412 , n9413 , n9414 , n9415 , n9416 , n9417 , n9418 , n9419 , n9420 , n9421 , n9422 , n9423 , n9424 , n9425 , n9426 , n9427 , n9428 , n9429 , n9430 , n9431 , n9432 , n9433 , n9434 , n9435 , n9436 , n9437 , n9438 , n9439 , n9440 , n9441 , n9442 , n9443 , n9444 , n9445 , n9446 , n9447 , n9448 , n9449 , n9450 , n9451 , n9452 , n9453 , n9454 , n9455 , n9456 , n9457 , n9458 , n9459 , n9460 , n9461 , n9462 , n9463 , n9464 , n9465 , n9466 , n9467 , n9468 , n9469 , n9470 , n9471 , n9472 , n9473 , n9474 , n9475 , n9476 , n9477 , n9478 , n9479 , n9480 , n9481 , n9482 , n9483 , n9484 , n9485 , n9486 , n9487 , n9488 , n9489 , n9490 , n9491 , n9492 , n9493 , n9494 , n9495 , n9496 , n9497 , n9498 , n9499 , n9500 , n9501 , n9502 , n9503 , n9504 , n9505 , n9506 , n9507 , n9508 , n9509 , n9510 , n9511 , n9512 , n9513 , n9514 , n9515 , n9516 , n9517 , n9518 , n9519 , n9520 , n9521 , n9522 , n9523 , n9524 , n9525 , n9526 , n9527 , n9528 , n9529 , n9530 , n9531 , n9532 , n9533 , n9534 , n9535 , n9536 , n9537 , n9538 , n9539 , n9540 , n9541 , n9542 , n9543 , n9544 , n9545 , n9546 , n9547 , n9548 , n9549 , n9550 , n9551 , n9552 , n9553 , n9554 , n9555 , n9556 , n9557 , n9558 , n9559 , n9560 , n9561 , n9562 , n9563 , n9564 , n9565 , n9566 , n9567 , n9568 , n9569 , n9570 , n9571 , n9572 , n9573 , n9574 , n9575 , n9576 , n9577 , n9578 , n9579 , n9580 , n9581 , n9582 , n9583 , n9584 , n9585 , n9586 , n9587 , n9588 , n9589 , n9590 , n9591 , n9592 , n9593 , n9594 , n9595 , n9596 , n9597 , n9598 , n9599 , n9600 , n9601 , n9602 , n9603 , n9604 , n9605 , n9606 , n9607 , n9608 , n9609 , n9610 , n9611 , n9612 , n9613 , n9614 , n9615 , n9616 , n9617 , n9618 , n9619 , n9620 , n9621 , n9622 , n9623 , n9624 , n9625 , n9626 , n9627 , n9628 , n9629 , n9630 , n9631 , n9632 , n9633 , n9634 , n9635 , n9636 , n9637 , n9638 , n9639 , n9640 , n9641 , n9642 , n9643 , n9644 , n9645 , n9646 , n9647 , n9648 , n9649 , n9650 , n9651 , n9652 , n9653 , n9654 , n9655 , n9656 , n9657 , n9658 , n9659 , n9660 , n9661 , n9662 , n9663 , n9664 , n9665 , n9666 , n9667 , n9668 , n9669 , n9670 , n9671 , n9672 , n9673 , n9674 , n9675 , n9676 , n9677 , n9678 , n9679 , n9680 , n9681 , n9682 , n9683 , n9684 , n9685 , n9686 , n9687 , n9688 , n9689 , n9690 , n9691 , n9692 , n9693 , n9694 , n9695 , n9696 , n9697 , n9698 , n9699 , n9700 , n9701 , n9702 , n9703 , n9704 , n9705 , n9706 , n9707 , n9708 , n9709 ;
  assign n1002 = \A[67]  & \A[68]  ;
  assign n1003 = ~\A[67]  & ~\A[68]  ;
  assign n1004 = ~n1002 & ~n1003 ;
  assign n1005 = \A[69]  & n1004 ;
  assign n1006 = ~n1002 & ~n1005 ;
  assign n1007 = \A[70]  & \A[71]  ;
  assign n1008 = ~\A[69]  & ~n1004 ;
  assign n1009 = ~n1005 & ~n1008 ;
  assign n1010 = ~\A[70]  & ~\A[71]  ;
  assign n1011 = ~n1007 & ~n1010 ;
  assign n1012 = \A[72]  & n1011 ;
  assign n1013 = ~\A[72]  & ~n1011 ;
  assign n1014 = ~n1012 & ~n1013 ;
  assign n1015 = n1009 & n1014 ;
  assign n1016 = n1007 & n1015 ;
  assign n1017 = ~n1007 & ~n1012 ;
  assign n1018 = ~n1015 & n1017 ;
  assign n1019 = ~n1016 & ~n1018 ;
  assign n1020 = n1006 & ~n1019 ;
  assign n1021 = ~n1006 & n1019 ;
  assign n1022 = ~n1020 & ~n1021 ;
  assign n1023 = \A[73]  & \A[74]  ;
  assign n1024 = ~\A[73]  & ~\A[74]  ;
  assign n1025 = ~n1023 & ~n1024 ;
  assign n1026 = \A[75]  & n1025 ;
  assign n1027 = ~\A[75]  & ~n1025 ;
  assign n1028 = ~n1026 & ~n1027 ;
  assign n1029 = \A[76]  & \A[77]  ;
  assign n1030 = ~\A[76]  & ~\A[77]  ;
  assign n1031 = ~n1029 & ~n1030 ;
  assign n1032 = \A[78]  & n1031 ;
  assign n1033 = ~\A[78]  & ~n1031 ;
  assign n1034 = ~n1032 & ~n1033 ;
  assign n1035 = n1028 & n1034 ;
  assign n1036 = ~n1029 & ~n1032 ;
  assign n1037 = ~n1023 & ~n1026 ;
  assign n1038 = ~n1036 & ~n1037 ;
  assign n1039 = n1036 & n1037 ;
  assign n1040 = ~n1038 & ~n1039 ;
  assign n1047 = n1035 & ~n1040 ;
  assign n1041 = ~n1035 & n1040 ;
  assign n1042 = ~n1009 & ~n1014 ;
  assign n1043 = ~n1015 & ~n1042 ;
  assign n1044 = ~n1028 & ~n1034 ;
  assign n1045 = ~n1035 & ~n1044 ;
  assign n1046 = n1043 & n1045 ;
  assign n1048 = ~n1041 & ~n1046 ;
  assign n1049 = ~n1047 & n1048 ;
  assign n1050 = n1022 & ~n1049 ;
  assign n1051 = n1040 & n1046 ;
  assign n1052 = ~n1006 & n1016 ;
  assign n1053 = n1051 & ~n1052 ;
  assign n1054 = ~n1050 & ~n1053 ;
  assign n1055 = ~n1029 & n1037 ;
  assign n1056 = n1035 & ~n1055 ;
  assign n1057 = ~n1038 & ~n1056 ;
  assign n1058 = ~n1054 & ~n1057 ;
  assign n1059 = ~n1006 & ~n1018 ;
  assign n1060 = ~n1016 & ~n1059 ;
  assign n1061 = n1054 & n1057 ;
  assign n1062 = ~n1060 & ~n1061 ;
  assign n1063 = ~n1058 & ~n1062 ;
  assign n1064 = \A[61]  & \A[62]  ;
  assign n1065 = ~\A[61]  & ~\A[62]  ;
  assign n1066 = ~n1064 & ~n1065 ;
  assign n1067 = \A[63]  & n1066 ;
  assign n1068 = ~\A[63]  & ~n1066 ;
  assign n1069 = ~n1067 & ~n1068 ;
  assign n1070 = \A[64]  & \A[65]  ;
  assign n1071 = ~\A[64]  & ~\A[65]  ;
  assign n1072 = ~n1070 & ~n1071 ;
  assign n1073 = \A[66]  & n1072 ;
  assign n1074 = ~\A[66]  & ~n1072 ;
  assign n1075 = ~n1073 & ~n1074 ;
  assign n1076 = n1069 & n1075 ;
  assign n1077 = ~n1069 & ~n1075 ;
  assign n1078 = ~n1076 & ~n1077 ;
  assign n1079 = \A[55]  & \A[56]  ;
  assign n1080 = ~\A[55]  & ~\A[56]  ;
  assign n1081 = ~n1079 & ~n1080 ;
  assign n1082 = \A[57]  & n1081 ;
  assign n1083 = ~\A[57]  & ~n1081 ;
  assign n1084 = ~n1082 & ~n1083 ;
  assign n1085 = \A[58]  & \A[59]  ;
  assign n1086 = ~\A[58]  & ~\A[59]  ;
  assign n1087 = ~n1085 & ~n1086 ;
  assign n1088 = \A[60]  & n1087 ;
  assign n1089 = ~\A[60]  & ~n1087 ;
  assign n1090 = ~n1088 & ~n1089 ;
  assign n1091 = n1084 & n1090 ;
  assign n1092 = ~n1084 & ~n1090 ;
  assign n1093 = ~n1091 & ~n1092 ;
  assign n1094 = n1078 & n1093 ;
  assign n1095 = ~n1064 & ~n1067 ;
  assign n1096 = ~n1070 & ~n1073 ;
  assign n1097 = ~n1076 & n1096 ;
  assign n1098 = n1070 & n1076 ;
  assign n1099 = ~n1097 & ~n1098 ;
  assign n1100 = n1095 & ~n1099 ;
  assign n1101 = ~n1095 & n1099 ;
  assign n1102 = ~n1100 & ~n1101 ;
  assign n1103 = ~n1094 & ~n1102 ;
  assign n1104 = ~n1079 & ~n1082 ;
  assign n1105 = n1085 & n1091 ;
  assign n1106 = ~n1085 & ~n1088 ;
  assign n1107 = ~n1091 & n1106 ;
  assign n1108 = ~n1105 & ~n1107 ;
  assign n1109 = n1104 & ~n1108 ;
  assign n1110 = ~n1104 & n1108 ;
  assign n1111 = ~n1109 & ~n1110 ;
  assign n1112 = ~n1103 & n1111 ;
  assign n1113 = n1094 & n1102 ;
  assign n1114 = ~n1095 & ~n1096 ;
  assign n1115 = ~n1104 & n1105 ;
  assign n1116 = ~n1114 & ~n1115 ;
  assign n1117 = n1113 & n1116 ;
  assign n1118 = ~n1112 & ~n1117 ;
  assign n1119 = ~n1095 & ~n1097 ;
  assign n1120 = ~n1098 & ~n1119 ;
  assign n1121 = ~n1118 & ~n1120 ;
  assign n1122 = ~n1104 & ~n1107 ;
  assign n1123 = ~n1105 & ~n1122 ;
  assign n1124 = n1118 & n1120 ;
  assign n1125 = ~n1123 & ~n1124 ;
  assign n1126 = ~n1121 & ~n1125 ;
  assign n1127 = n1063 & n1126 ;
  assign n1128 = ~n1063 & ~n1126 ;
  assign n1129 = ~n1121 & ~n1124 ;
  assign n1130 = n1123 & ~n1129 ;
  assign n1131 = ~n1123 & n1129 ;
  assign n1132 = ~n1130 & ~n1131 ;
  assign n1133 = ~n1058 & ~n1061 ;
  assign n1134 = n1060 & ~n1133 ;
  assign n1135 = ~n1060 & n1133 ;
  assign n1136 = ~n1134 & ~n1135 ;
  assign n1137 = ~n1132 & ~n1136 ;
  assign n1138 = ~n1043 & ~n1045 ;
  assign n1139 = ~n1046 & ~n1138 ;
  assign n1140 = ~n1078 & ~n1093 ;
  assign n1141 = ~n1094 & ~n1140 ;
  assign n1142 = n1139 & n1141 ;
  assign n1143 = n1050 & ~n1053 ;
  assign n1144 = ~n1049 & ~n1051 ;
  assign n1145 = ~n1022 & ~n1144 ;
  assign n1146 = ~n1143 & ~n1145 ;
  assign n1147 = ~n1142 & ~n1146 ;
  assign n1148 = n1112 & ~n1117 ;
  assign n1149 = ~n1103 & ~n1113 ;
  assign n1150 = ~n1111 & ~n1149 ;
  assign n1151 = ~n1148 & ~n1150 ;
  assign n1152 = n1142 & n1146 ;
  assign n1153 = ~n1151 & ~n1152 ;
  assign n1154 = ~n1147 & ~n1153 ;
  assign n1155 = n1132 & n1136 ;
  assign n1156 = ~n1154 & ~n1155 ;
  assign n1157 = ~n1137 & ~n1156 ;
  assign n1158 = ~n1128 & ~n1157 ;
  assign n1159 = ~n1127 & ~n1158 ;
  assign n1160 = \A[43]  & \A[44]  ;
  assign n1161 = ~\A[43]  & ~\A[44]  ;
  assign n1162 = ~n1160 & ~n1161 ;
  assign n1163 = \A[45]  & n1162 ;
  assign n1164 = ~n1160 & ~n1163 ;
  assign n1165 = \A[46]  & \A[47]  ;
  assign n1166 = ~\A[45]  & ~n1162 ;
  assign n1167 = ~n1163 & ~n1166 ;
  assign n1168 = ~\A[46]  & ~\A[47]  ;
  assign n1169 = ~n1165 & ~n1168 ;
  assign n1170 = \A[48]  & n1169 ;
  assign n1171 = ~\A[48]  & ~n1169 ;
  assign n1172 = ~n1170 & ~n1171 ;
  assign n1173 = n1167 & n1172 ;
  assign n1174 = n1165 & n1173 ;
  assign n1175 = ~n1165 & ~n1170 ;
  assign n1176 = ~n1173 & n1175 ;
  assign n1177 = ~n1174 & ~n1176 ;
  assign n1178 = n1164 & ~n1177 ;
  assign n1179 = ~n1164 & n1177 ;
  assign n1180 = ~n1178 & ~n1179 ;
  assign n1181 = \A[49]  & \A[50]  ;
  assign n1182 = ~\A[49]  & ~\A[50]  ;
  assign n1183 = ~n1181 & ~n1182 ;
  assign n1184 = \A[51]  & n1183 ;
  assign n1185 = ~\A[51]  & ~n1183 ;
  assign n1186 = ~n1184 & ~n1185 ;
  assign n1187 = \A[52]  & \A[53]  ;
  assign n1188 = ~\A[52]  & ~\A[53]  ;
  assign n1189 = ~n1187 & ~n1188 ;
  assign n1190 = \A[54]  & n1189 ;
  assign n1191 = ~\A[54]  & ~n1189 ;
  assign n1192 = ~n1190 & ~n1191 ;
  assign n1193 = n1186 & n1192 ;
  assign n1194 = ~n1187 & ~n1190 ;
  assign n1195 = ~n1181 & ~n1184 ;
  assign n1196 = ~n1194 & ~n1195 ;
  assign n1197 = n1194 & n1195 ;
  assign n1198 = ~n1196 & ~n1197 ;
  assign n1205 = n1193 & ~n1198 ;
  assign n1199 = ~n1193 & n1198 ;
  assign n1200 = ~n1167 & ~n1172 ;
  assign n1201 = ~n1173 & ~n1200 ;
  assign n1202 = ~n1186 & ~n1192 ;
  assign n1203 = ~n1193 & ~n1202 ;
  assign n1204 = n1201 & n1203 ;
  assign n1206 = ~n1199 & ~n1204 ;
  assign n1207 = ~n1205 & n1206 ;
  assign n1208 = n1180 & ~n1207 ;
  assign n1209 = n1198 & n1204 ;
  assign n1210 = ~n1164 & n1174 ;
  assign n1211 = n1209 & ~n1210 ;
  assign n1212 = ~n1208 & ~n1211 ;
  assign n1213 = ~n1187 & n1195 ;
  assign n1214 = n1193 & ~n1213 ;
  assign n1215 = ~n1196 & ~n1214 ;
  assign n1216 = ~n1212 & ~n1215 ;
  assign n1217 = ~n1164 & ~n1176 ;
  assign n1218 = ~n1174 & ~n1217 ;
  assign n1219 = n1212 & n1215 ;
  assign n1220 = ~n1218 & ~n1219 ;
  assign n1221 = ~n1216 & ~n1220 ;
  assign n1222 = \A[37]  & \A[38]  ;
  assign n1223 = ~\A[37]  & ~\A[38]  ;
  assign n1224 = ~n1222 & ~n1223 ;
  assign n1225 = \A[39]  & n1224 ;
  assign n1226 = ~\A[39]  & ~n1224 ;
  assign n1227 = ~n1225 & ~n1226 ;
  assign n1228 = \A[40]  & \A[41]  ;
  assign n1229 = ~\A[40]  & ~\A[41]  ;
  assign n1230 = ~n1228 & ~n1229 ;
  assign n1231 = \A[42]  & n1230 ;
  assign n1232 = ~\A[42]  & ~n1230 ;
  assign n1233 = ~n1231 & ~n1232 ;
  assign n1234 = n1227 & n1233 ;
  assign n1235 = ~n1227 & ~n1233 ;
  assign n1236 = ~n1234 & ~n1235 ;
  assign n1237 = \A[31]  & \A[32]  ;
  assign n1238 = ~\A[31]  & ~\A[32]  ;
  assign n1239 = ~n1237 & ~n1238 ;
  assign n1240 = \A[33]  & n1239 ;
  assign n1241 = ~\A[33]  & ~n1239 ;
  assign n1242 = ~n1240 & ~n1241 ;
  assign n1243 = \A[34]  & \A[35]  ;
  assign n1244 = ~\A[34]  & ~\A[35]  ;
  assign n1245 = ~n1243 & ~n1244 ;
  assign n1246 = \A[36]  & n1245 ;
  assign n1247 = ~\A[36]  & ~n1245 ;
  assign n1248 = ~n1246 & ~n1247 ;
  assign n1249 = n1242 & n1248 ;
  assign n1250 = ~n1242 & ~n1248 ;
  assign n1251 = ~n1249 & ~n1250 ;
  assign n1252 = n1236 & n1251 ;
  assign n1253 = ~n1228 & ~n1231 ;
  assign n1254 = ~n1222 & ~n1225 ;
  assign n1255 = ~n1253 & ~n1254 ;
  assign n1256 = n1253 & n1254 ;
  assign n1257 = ~n1255 & ~n1256 ;
  assign n1258 = n1252 & n1257 ;
  assign n1259 = ~n1243 & ~n1246 ;
  assign n1260 = ~n1237 & ~n1240 ;
  assign n1261 = ~n1259 & ~n1260 ;
  assign n1262 = n1259 & n1260 ;
  assign n1263 = ~n1261 & ~n1262 ;
  assign n1264 = n1249 & ~n1263 ;
  assign n1265 = ~n1249 & n1263 ;
  assign n1266 = ~n1264 & ~n1265 ;
  assign n1267 = ~n1258 & n1266 ;
  assign n1269 = n1234 & ~n1257 ;
  assign n1268 = ~n1234 & n1257 ;
  assign n1270 = ~n1252 & ~n1268 ;
  assign n1271 = ~n1269 & n1270 ;
  assign n1272 = ~n1267 & ~n1271 ;
  assign n1273 = ~n1234 & ~n1255 ;
  assign n1274 = ~n1256 & ~n1273 ;
  assign n1275 = ~n1272 & ~n1274 ;
  assign n1276 = n1272 & n1274 ;
  assign n1277 = ~n1249 & ~n1261 ;
  assign n1278 = ~n1262 & ~n1277 ;
  assign n1279 = ~n1276 & ~n1278 ;
  assign n1280 = ~n1275 & ~n1279 ;
  assign n1281 = ~n1221 & n1280 ;
  assign n1282 = n1221 & ~n1280 ;
  assign n1283 = ~n1216 & ~n1219 ;
  assign n1284 = n1218 & ~n1283 ;
  assign n1285 = ~n1218 & n1283 ;
  assign n1286 = ~n1284 & ~n1285 ;
  assign n1287 = ~n1275 & ~n1276 ;
  assign n1288 = ~n1278 & n1287 ;
  assign n1289 = n1278 & ~n1287 ;
  assign n1290 = ~n1288 & ~n1289 ;
  assign n1291 = n1286 & ~n1290 ;
  assign n1292 = ~n1286 & n1290 ;
  assign n1293 = ~n1201 & ~n1203 ;
  assign n1294 = ~n1204 & ~n1293 ;
  assign n1295 = ~n1236 & ~n1251 ;
  assign n1296 = ~n1252 & ~n1295 ;
  assign n1297 = n1294 & n1296 ;
  assign n1298 = n1208 & ~n1211 ;
  assign n1299 = ~n1207 & ~n1209 ;
  assign n1300 = ~n1180 & ~n1299 ;
  assign n1301 = ~n1298 & ~n1300 ;
  assign n1302 = n1297 & n1301 ;
  assign n1303 = ~n1297 & ~n1301 ;
  assign n1304 = ~n1258 & ~n1271 ;
  assign n1305 = n1266 & n1304 ;
  assign n1306 = ~n1266 & ~n1304 ;
  assign n1307 = ~n1305 & ~n1306 ;
  assign n1308 = ~n1303 & ~n1307 ;
  assign n1309 = ~n1302 & ~n1308 ;
  assign n1310 = ~n1292 & ~n1309 ;
  assign n1311 = ~n1291 & ~n1310 ;
  assign n1312 = ~n1282 & ~n1311 ;
  assign n1313 = ~n1281 & ~n1312 ;
  assign n1314 = n1159 & ~n1313 ;
  assign n1315 = ~n1159 & n1313 ;
  assign n1316 = ~n1127 & ~n1128 ;
  assign n1317 = n1157 & ~n1316 ;
  assign n1318 = ~n1157 & n1316 ;
  assign n1319 = ~n1317 & ~n1318 ;
  assign n1320 = ~n1281 & ~n1282 ;
  assign n1321 = ~n1311 & n1320 ;
  assign n1322 = n1311 & ~n1320 ;
  assign n1323 = ~n1321 & ~n1322 ;
  assign n1324 = n1319 & ~n1323 ;
  assign n1325 = ~n1319 & n1323 ;
  assign n1326 = ~n1137 & ~n1155 ;
  assign n1327 = n1154 & n1326 ;
  assign n1328 = ~n1154 & ~n1326 ;
  assign n1329 = ~n1327 & ~n1328 ;
  assign n1330 = ~n1291 & ~n1292 ;
  assign n1331 = ~n1309 & n1330 ;
  assign n1332 = n1309 & ~n1330 ;
  assign n1333 = ~n1331 & ~n1332 ;
  assign n1334 = n1329 & n1333 ;
  assign n1335 = ~n1329 & ~n1333 ;
  assign n1336 = ~n1139 & ~n1141 ;
  assign n1337 = ~n1142 & ~n1336 ;
  assign n1338 = ~n1294 & ~n1296 ;
  assign n1339 = ~n1297 & ~n1338 ;
  assign n1340 = n1337 & n1339 ;
  assign n1341 = ~n1147 & ~n1152 ;
  assign n1342 = n1151 & ~n1341 ;
  assign n1343 = ~n1151 & n1341 ;
  assign n1344 = ~n1342 & ~n1343 ;
  assign n1345 = n1340 & ~n1344 ;
  assign n1346 = ~n1340 & n1344 ;
  assign n1347 = ~n1302 & ~n1303 ;
  assign n1348 = ~n1307 & n1347 ;
  assign n1349 = n1307 & ~n1347 ;
  assign n1350 = ~n1348 & ~n1349 ;
  assign n1351 = ~n1346 & n1350 ;
  assign n1352 = ~n1345 & ~n1351 ;
  assign n1353 = ~n1335 & ~n1352 ;
  assign n1354 = ~n1334 & ~n1353 ;
  assign n1355 = ~n1325 & n1354 ;
  assign n1356 = ~n1324 & ~n1355 ;
  assign n1357 = ~n1315 & n1356 ;
  assign n1358 = ~n1314 & ~n1357 ;
  assign n1359 = \A[3]  & \A[4]  ;
  assign n1360 = ~\A[3]  & ~\A[4]  ;
  assign n1361 = ~n1359 & ~n1360 ;
  assign n1362 = \A[5]  & n1361 ;
  assign n1363 = ~n1359 & ~n1362 ;
  assign n1364 = \A[0]  & \A[1]  ;
  assign n1365 = ~\A[0]  & ~\A[1]  ;
  assign n1366 = ~n1364 & ~n1365 ;
  assign n1367 = \A[2]  & n1366 ;
  assign n1368 = ~n1364 & ~n1367 ;
  assign n1369 = ~n1363 & ~n1368 ;
  assign n1370 = ~\A[2]  & ~n1366 ;
  assign n1371 = ~n1367 & ~n1370 ;
  assign n1372 = \A[6]  & n1371 ;
  assign n1373 = ~\A[6]  & ~n1371 ;
  assign n1374 = ~n1372 & ~n1373 ;
  assign n1375 = ~\A[5]  & ~n1361 ;
  assign n1376 = ~n1362 & ~n1375 ;
  assign n1377 = n1374 & n1376 ;
  assign n1378 = ~n1372 & ~n1377 ;
  assign n1379 = n1363 & n1368 ;
  assign n1380 = ~n1369 & ~n1379 ;
  assign n1381 = ~n1378 & n1380 ;
  assign n1382 = ~n1369 & ~n1381 ;
  assign n1383 = ~n1374 & ~n1376 ;
  assign n1384 = ~n1377 & ~n1383 ;
  assign n1385 = \A[997]  & \A[998]  ;
  assign n1386 = ~\A[997]  & ~\A[998]  ;
  assign n1387 = ~n1385 & ~n1386 ;
  assign n1388 = \A[999]  & n1387 ;
  assign n1389 = ~\A[999]  & ~n1387 ;
  assign n1390 = ~n1388 & ~n1389 ;
  assign n1391 = n1384 & n1390 ;
  assign n1392 = n1378 & ~n1380 ;
  assign n1393 = ~n1381 & ~n1392 ;
  assign n1394 = ~n1391 & ~n1393 ;
  assign n1395 = ~n1385 & ~n1388 ;
  assign n1396 = n1391 & n1393 ;
  assign n1397 = n1395 & ~n1396 ;
  assign n1398 = ~n1394 & ~n1397 ;
  assign n1399 = ~n1382 & n1398 ;
  assign n1400 = ~n1384 & ~n1390 ;
  assign n1401 = ~n1391 & ~n1400 ;
  assign n1402 = \A[991]  & \A[992]  ;
  assign n1403 = ~\A[991]  & ~\A[992]  ;
  assign n1404 = ~n1402 & ~n1403 ;
  assign n1405 = \A[993]  & n1404 ;
  assign n1406 = ~\A[993]  & ~n1404 ;
  assign n1407 = ~n1405 & ~n1406 ;
  assign n1408 = \A[994]  & \A[995]  ;
  assign n1409 = ~\A[994]  & ~\A[995]  ;
  assign n1410 = ~n1408 & ~n1409 ;
  assign n1411 = \A[996]  & n1410 ;
  assign n1412 = ~\A[996]  & ~n1410 ;
  assign n1413 = ~n1411 & ~n1412 ;
  assign n1414 = n1407 & n1413 ;
  assign n1415 = ~n1407 & ~n1413 ;
  assign n1416 = ~n1414 & ~n1415 ;
  assign n1417 = n1401 & n1416 ;
  assign n1418 = ~n1394 & ~n1396 ;
  assign n1419 = n1395 & ~n1418 ;
  assign n1420 = ~n1395 & n1418 ;
  assign n1421 = ~n1419 & ~n1420 ;
  assign n1422 = ~n1417 & ~n1421 ;
  assign n1423 = n1417 & n1421 ;
  assign n1424 = ~n1408 & ~n1411 ;
  assign n1425 = ~n1402 & ~n1405 ;
  assign n1426 = ~n1424 & ~n1425 ;
  assign n1427 = n1424 & n1425 ;
  assign n1428 = ~n1426 & ~n1427 ;
  assign n1429 = n1414 & ~n1428 ;
  assign n1430 = ~n1414 & n1428 ;
  assign n1431 = ~n1429 & ~n1430 ;
  assign n1432 = ~n1423 & n1431 ;
  assign n1433 = ~n1422 & ~n1432 ;
  assign n1434 = ~n1414 & ~n1426 ;
  assign n1435 = ~n1427 & ~n1434 ;
  assign n1436 = n1433 & n1435 ;
  assign n1437 = n1399 & n1436 ;
  assign n1438 = \A[19]  & \A[20]  ;
  assign n1439 = ~\A[19]  & ~\A[20]  ;
  assign n1440 = ~n1438 & ~n1439 ;
  assign n1441 = \A[21]  & n1440 ;
  assign n1442 = ~\A[21]  & ~n1440 ;
  assign n1443 = ~n1441 & ~n1442 ;
  assign n1444 = \A[22]  & \A[23]  ;
  assign n1445 = ~\A[22]  & ~\A[23]  ;
  assign n1446 = ~n1444 & ~n1445 ;
  assign n1447 = \A[24]  & n1446 ;
  assign n1448 = ~\A[24]  & ~n1446 ;
  assign n1449 = ~n1447 & ~n1448 ;
  assign n1450 = n1443 & n1449 ;
  assign n1451 = ~n1443 & ~n1449 ;
  assign n1452 = ~n1450 & ~n1451 ;
  assign n1453 = \A[25]  & \A[26]  ;
  assign n1454 = ~\A[25]  & ~\A[26]  ;
  assign n1455 = ~n1453 & ~n1454 ;
  assign n1456 = \A[27]  & n1455 ;
  assign n1457 = ~\A[27]  & ~n1455 ;
  assign n1458 = ~n1456 & ~n1457 ;
  assign n1459 = \A[28]  & \A[29]  ;
  assign n1460 = ~\A[28]  & ~\A[29]  ;
  assign n1461 = ~n1459 & ~n1460 ;
  assign n1462 = \A[30]  & n1461 ;
  assign n1463 = ~\A[30]  & ~n1461 ;
  assign n1464 = ~n1462 & ~n1463 ;
  assign n1465 = n1458 & n1464 ;
  assign n1466 = ~n1458 & ~n1464 ;
  assign n1467 = ~n1465 & ~n1466 ;
  assign n1468 = n1452 & n1467 ;
  assign n1469 = ~n1459 & ~n1462 ;
  assign n1470 = ~n1453 & ~n1456 ;
  assign n1471 = n1469 & n1470 ;
  assign n1472 = ~n1469 & ~n1470 ;
  assign n1473 = ~n1471 & ~n1472 ;
  assign n1474 = n1468 & n1473 ;
  assign n1475 = ~n1444 & ~n1447 ;
  assign n1476 = ~n1438 & ~n1441 ;
  assign n1477 = ~n1475 & ~n1476 ;
  assign n1478 = n1475 & n1476 ;
  assign n1479 = ~n1477 & ~n1478 ;
  assign n1480 = n1450 & ~n1479 ;
  assign n1481 = ~n1450 & n1479 ;
  assign n1482 = ~n1480 & ~n1481 ;
  assign n1483 = ~n1474 & n1482 ;
  assign n1485 = n1465 & ~n1473 ;
  assign n1484 = ~n1465 & n1473 ;
  assign n1486 = ~n1468 & ~n1484 ;
  assign n1487 = ~n1485 & n1486 ;
  assign n1488 = ~n1483 & ~n1487 ;
  assign n1489 = n1465 & ~n1471 ;
  assign n1490 = ~n1472 & ~n1489 ;
  assign n1491 = ~n1488 & n1490 ;
  assign n1492 = n1488 & ~n1490 ;
  assign n1493 = ~n1450 & ~n1477 ;
  assign n1494 = ~n1478 & ~n1493 ;
  assign n1495 = ~n1492 & ~n1494 ;
  assign n1496 = ~n1491 & ~n1495 ;
  assign n1497 = \A[7]  & \A[8]  ;
  assign n1498 = ~\A[7]  & ~\A[8]  ;
  assign n1499 = ~n1497 & ~n1498 ;
  assign n1500 = \A[9]  & n1499 ;
  assign n1501 = ~\A[9]  & ~n1499 ;
  assign n1502 = ~n1500 & ~n1501 ;
  assign n1503 = \A[10]  & \A[11]  ;
  assign n1504 = ~\A[10]  & ~\A[11]  ;
  assign n1505 = ~n1503 & ~n1504 ;
  assign n1506 = \A[12]  & n1505 ;
  assign n1507 = ~\A[12]  & ~n1505 ;
  assign n1508 = ~n1506 & ~n1507 ;
  assign n1509 = n1502 & n1508 ;
  assign n1510 = ~n1502 & ~n1508 ;
  assign n1511 = ~n1509 & ~n1510 ;
  assign n1512 = \A[13]  & \A[14]  ;
  assign n1513 = ~\A[13]  & ~\A[14]  ;
  assign n1514 = ~n1512 & ~n1513 ;
  assign n1515 = \A[15]  & n1514 ;
  assign n1516 = ~\A[15]  & ~n1514 ;
  assign n1517 = ~n1515 & ~n1516 ;
  assign n1518 = \A[16]  & \A[17]  ;
  assign n1519 = ~\A[16]  & ~\A[17]  ;
  assign n1520 = ~n1518 & ~n1519 ;
  assign n1521 = \A[18]  & n1520 ;
  assign n1522 = ~\A[18]  & ~n1520 ;
  assign n1523 = ~n1521 & ~n1522 ;
  assign n1524 = n1517 & n1523 ;
  assign n1525 = ~n1517 & ~n1523 ;
  assign n1526 = ~n1524 & ~n1525 ;
  assign n1527 = n1511 & n1526 ;
  assign n1528 = ~n1518 & ~n1521 ;
  assign n1529 = ~n1512 & ~n1515 ;
  assign n1530 = n1528 & n1529 ;
  assign n1531 = ~n1528 & ~n1529 ;
  assign n1532 = ~n1530 & ~n1531 ;
  assign n1533 = n1527 & n1532 ;
  assign n1534 = ~n1503 & ~n1506 ;
  assign n1535 = ~n1497 & ~n1500 ;
  assign n1536 = ~n1534 & ~n1535 ;
  assign n1537 = n1534 & n1535 ;
  assign n1538 = ~n1536 & ~n1537 ;
  assign n1539 = n1509 & ~n1538 ;
  assign n1540 = ~n1509 & n1538 ;
  assign n1541 = ~n1539 & ~n1540 ;
  assign n1542 = ~n1533 & n1541 ;
  assign n1544 = n1524 & ~n1532 ;
  assign n1543 = ~n1524 & n1532 ;
  assign n1545 = ~n1527 & ~n1543 ;
  assign n1546 = ~n1544 & n1545 ;
  assign n1547 = ~n1542 & ~n1546 ;
  assign n1548 = n1524 & ~n1530 ;
  assign n1549 = ~n1531 & ~n1548 ;
  assign n1550 = ~n1547 & n1549 ;
  assign n1551 = n1547 & ~n1549 ;
  assign n1552 = ~n1509 & ~n1536 ;
  assign n1553 = ~n1537 & ~n1552 ;
  assign n1554 = ~n1551 & ~n1553 ;
  assign n1555 = ~n1550 & ~n1554 ;
  assign n1556 = n1496 & n1555 ;
  assign n1557 = ~n1496 & ~n1555 ;
  assign n1558 = ~n1550 & ~n1551 ;
  assign n1559 = ~n1553 & n1558 ;
  assign n1560 = n1553 & ~n1558 ;
  assign n1561 = ~n1559 & ~n1560 ;
  assign n1562 = ~n1491 & ~n1492 ;
  assign n1563 = ~n1494 & n1562 ;
  assign n1564 = n1494 & ~n1562 ;
  assign n1565 = ~n1563 & ~n1564 ;
  assign n1566 = ~n1561 & ~n1565 ;
  assign n1567 = n1561 & n1565 ;
  assign n1568 = ~n1452 & ~n1467 ;
  assign n1569 = ~n1468 & ~n1568 ;
  assign n1570 = ~n1511 & ~n1526 ;
  assign n1571 = ~n1527 & ~n1570 ;
  assign n1572 = n1569 & n1571 ;
  assign n1573 = ~n1474 & ~n1487 ;
  assign n1574 = n1482 & n1573 ;
  assign n1575 = ~n1482 & ~n1573 ;
  assign n1576 = ~n1574 & ~n1575 ;
  assign n1577 = n1572 & ~n1576 ;
  assign n1578 = ~n1572 & n1576 ;
  assign n1579 = ~n1533 & ~n1546 ;
  assign n1580 = n1541 & n1579 ;
  assign n1581 = ~n1541 & ~n1579 ;
  assign n1582 = ~n1580 & ~n1581 ;
  assign n1583 = ~n1578 & ~n1582 ;
  assign n1584 = ~n1577 & ~n1583 ;
  assign n1585 = ~n1567 & ~n1584 ;
  assign n1586 = ~n1566 & ~n1585 ;
  assign n1587 = ~n1557 & ~n1586 ;
  assign n1588 = ~n1556 & ~n1587 ;
  assign n1589 = n1437 & ~n1588 ;
  assign n1590 = ~n1437 & n1588 ;
  assign n1591 = ~n1399 & ~n1436 ;
  assign n1592 = ~n1437 & ~n1591 ;
  assign n1593 = n1382 & ~n1398 ;
  assign n1594 = ~n1399 & ~n1593 ;
  assign n1595 = ~n1433 & ~n1435 ;
  assign n1596 = n1594 & ~n1595 ;
  assign n1597 = ~n1592 & ~n1596 ;
  assign n1598 = ~n1556 & ~n1557 ;
  assign n1599 = ~n1586 & n1598 ;
  assign n1600 = n1586 & ~n1598 ;
  assign n1601 = ~n1599 & ~n1600 ;
  assign n1602 = n1597 & ~n1601 ;
  assign n1603 = ~n1597 & n1601 ;
  assign n1604 = ~n1435 & n1594 ;
  assign n1605 = n1435 & ~n1594 ;
  assign n1606 = ~n1604 & ~n1605 ;
  assign n1607 = n1433 & n1606 ;
  assign n1608 = ~n1433 & ~n1606 ;
  assign n1609 = ~n1607 & ~n1608 ;
  assign n1610 = ~n1566 & ~n1567 ;
  assign n1611 = ~n1584 & n1610 ;
  assign n1612 = n1584 & ~n1610 ;
  assign n1613 = ~n1611 & ~n1612 ;
  assign n1614 = ~n1609 & n1613 ;
  assign n1615 = n1609 & ~n1613 ;
  assign n1616 = ~n1569 & ~n1571 ;
  assign n1617 = ~n1572 & ~n1616 ;
  assign n1618 = ~n1401 & ~n1416 ;
  assign n1619 = ~n1417 & ~n1618 ;
  assign n1620 = n1617 & n1619 ;
  assign n1621 = ~n1577 & ~n1578 ;
  assign n1622 = ~n1582 & n1621 ;
  assign n1623 = n1582 & ~n1621 ;
  assign n1624 = ~n1622 & ~n1623 ;
  assign n1625 = n1620 & n1624 ;
  assign n1626 = ~n1620 & ~n1624 ;
  assign n1627 = ~n1422 & ~n1423 ;
  assign n1628 = n1431 & n1627 ;
  assign n1629 = ~n1431 & ~n1627 ;
  assign n1630 = ~n1628 & ~n1629 ;
  assign n1631 = ~n1626 & ~n1630 ;
  assign n1632 = ~n1625 & ~n1631 ;
  assign n1633 = ~n1615 & ~n1632 ;
  assign n1634 = ~n1614 & ~n1633 ;
  assign n1635 = ~n1603 & n1634 ;
  assign n1636 = ~n1602 & ~n1635 ;
  assign n1637 = ~n1590 & n1636 ;
  assign n1638 = ~n1589 & ~n1637 ;
  assign n1639 = n1358 & n1638 ;
  assign n1640 = ~n1358 & ~n1638 ;
  assign n1641 = ~n1639 & ~n1640 ;
  assign n1642 = ~n1314 & ~n1315 ;
  assign n1643 = ~n1356 & n1642 ;
  assign n1644 = n1356 & ~n1642 ;
  assign n1645 = ~n1643 & ~n1644 ;
  assign n1646 = ~n1589 & ~n1590 ;
  assign n1647 = ~n1636 & n1646 ;
  assign n1648 = n1636 & ~n1646 ;
  assign n1649 = ~n1647 & ~n1648 ;
  assign n1650 = ~n1645 & ~n1649 ;
  assign n1651 = n1645 & n1649 ;
  assign n1652 = ~n1324 & ~n1325 ;
  assign n1653 = ~n1354 & n1652 ;
  assign n1654 = n1354 & ~n1652 ;
  assign n1655 = ~n1653 & ~n1654 ;
  assign n1656 = ~n1602 & ~n1603 ;
  assign n1657 = n1634 & n1656 ;
  assign n1658 = ~n1634 & ~n1656 ;
  assign n1659 = ~n1657 & ~n1658 ;
  assign n1660 = n1655 & ~n1659 ;
  assign n1661 = ~n1655 & n1659 ;
  assign n1662 = ~n1614 & ~n1615 ;
  assign n1663 = ~n1632 & n1662 ;
  assign n1664 = n1632 & ~n1662 ;
  assign n1665 = ~n1663 & ~n1664 ;
  assign n1666 = ~n1334 & ~n1335 ;
  assign n1667 = ~n1352 & n1666 ;
  assign n1668 = n1352 & ~n1666 ;
  assign n1669 = ~n1667 & ~n1668 ;
  assign n1670 = ~n1665 & ~n1669 ;
  assign n1671 = n1665 & n1669 ;
  assign n1672 = ~n1617 & ~n1619 ;
  assign n1673 = ~n1620 & ~n1672 ;
  assign n1674 = ~n1337 & ~n1339 ;
  assign n1675 = ~n1340 & ~n1674 ;
  assign n1676 = n1673 & n1675 ;
  assign n1677 = ~n1345 & ~n1346 ;
  assign n1678 = ~n1350 & n1677 ;
  assign n1679 = n1350 & ~n1677 ;
  assign n1680 = ~n1678 & ~n1679 ;
  assign n1681 = n1676 & ~n1680 ;
  assign n1682 = ~n1676 & n1680 ;
  assign n1683 = ~n1625 & ~n1626 ;
  assign n1684 = ~n1630 & n1683 ;
  assign n1685 = n1630 & ~n1683 ;
  assign n1686 = ~n1684 & ~n1685 ;
  assign n1687 = ~n1682 & n1686 ;
  assign n1688 = ~n1681 & ~n1687 ;
  assign n1689 = ~n1671 & n1688 ;
  assign n1690 = ~n1670 & ~n1689 ;
  assign n1691 = ~n1661 & n1690 ;
  assign n1692 = ~n1660 & ~n1691 ;
  assign n1693 = ~n1651 & ~n1692 ;
  assign n1694 = ~n1650 & ~n1693 ;
  assign n1695 = n1641 & ~n1694 ;
  assign n1696 = ~n1641 & n1694 ;
  assign n1697 = ~n1695 & ~n1696 ;
  assign n1698 = \A[946]  & \A[947]  ;
  assign n1699 = \A[943]  & \A[944]  ;
  assign n1700 = ~\A[943]  & ~\A[944]  ;
  assign n1701 = ~n1699 & ~n1700 ;
  assign n1702 = \A[945]  & n1701 ;
  assign n1703 = ~\A[945]  & ~n1701 ;
  assign n1704 = ~n1702 & ~n1703 ;
  assign n1705 = ~\A[946]  & ~\A[947]  ;
  assign n1706 = ~n1698 & ~n1705 ;
  assign n1707 = \A[948]  & n1706 ;
  assign n1708 = ~\A[948]  & ~n1706 ;
  assign n1709 = ~n1707 & ~n1708 ;
  assign n1710 = n1704 & n1709 ;
  assign n1711 = n1698 & n1710 ;
  assign n1712 = ~n1699 & ~n1702 ;
  assign n1713 = ~n1698 & ~n1707 ;
  assign n1714 = ~n1710 & n1713 ;
  assign n1715 = ~n1712 & ~n1714 ;
  assign n1716 = ~n1711 & ~n1715 ;
  assign n1717 = \A[952]  & \A[953]  ;
  assign n1718 = ~\A[952]  & ~\A[953]  ;
  assign n1719 = ~n1717 & ~n1718 ;
  assign n1720 = \A[954]  & n1719 ;
  assign n1721 = ~n1717 & ~n1720 ;
  assign n1722 = \A[949]  & \A[950]  ;
  assign n1723 = ~\A[949]  & ~\A[950]  ;
  assign n1724 = ~n1722 & ~n1723 ;
  assign n1725 = \A[951]  & n1724 ;
  assign n1726 = ~n1722 & ~n1725 ;
  assign n1727 = n1721 & n1726 ;
  assign n1728 = ~n1721 & ~n1726 ;
  assign n1729 = ~\A[951]  & ~n1724 ;
  assign n1730 = ~n1725 & ~n1729 ;
  assign n1731 = ~\A[954]  & ~n1719 ;
  assign n1732 = ~n1720 & ~n1731 ;
  assign n1733 = n1730 & n1732 ;
  assign n1734 = ~n1728 & ~n1733 ;
  assign n1735 = ~n1727 & ~n1734 ;
  assign n1736 = ~n1730 & ~n1732 ;
  assign n1737 = ~n1733 & ~n1736 ;
  assign n1738 = ~n1704 & ~n1709 ;
  assign n1739 = ~n1710 & ~n1738 ;
  assign n1740 = n1737 & n1739 ;
  assign n1741 = n1711 & ~n1712 ;
  assign n1742 = n1740 & ~n1741 ;
  assign n1743 = ~n1727 & ~n1728 ;
  assign n1744 = n1733 & ~n1743 ;
  assign n1745 = ~n1733 & n1743 ;
  assign n1746 = ~n1744 & ~n1745 ;
  assign n1747 = n1742 & ~n1746 ;
  assign n1748 = ~n1742 & n1746 ;
  assign n1749 = ~n1711 & ~n1714 ;
  assign n1750 = n1712 & ~n1749 ;
  assign n1751 = ~n1712 & n1749 ;
  assign n1752 = ~n1750 & ~n1751 ;
  assign n1753 = ~n1748 & n1752 ;
  assign n1754 = ~n1747 & ~n1753 ;
  assign n1755 = n1735 & ~n1754 ;
  assign n1756 = ~n1735 & n1754 ;
  assign n1757 = ~n1755 & ~n1756 ;
  assign n1758 = n1716 & n1757 ;
  assign n1759 = ~n1716 & ~n1757 ;
  assign n1760 = ~n1758 & ~n1759 ;
  assign n1761 = \A[958]  & \A[959]  ;
  assign n1762 = \A[955]  & \A[956]  ;
  assign n1763 = ~\A[955]  & ~\A[956]  ;
  assign n1764 = ~n1762 & ~n1763 ;
  assign n1765 = \A[957]  & n1764 ;
  assign n1766 = ~\A[957]  & ~n1764 ;
  assign n1767 = ~n1765 & ~n1766 ;
  assign n1768 = ~\A[958]  & ~\A[959]  ;
  assign n1769 = ~n1761 & ~n1768 ;
  assign n1770 = \A[960]  & n1769 ;
  assign n1771 = ~\A[960]  & ~n1769 ;
  assign n1772 = ~n1770 & ~n1771 ;
  assign n1773 = n1767 & n1772 ;
  assign n1774 = n1761 & n1773 ;
  assign n1775 = ~n1762 & ~n1765 ;
  assign n1776 = ~n1761 & ~n1770 ;
  assign n1777 = ~n1773 & n1776 ;
  assign n1778 = ~n1775 & ~n1777 ;
  assign n1779 = ~n1774 & ~n1778 ;
  assign n1780 = \A[964]  & \A[965]  ;
  assign n1781 = ~\A[964]  & ~\A[965]  ;
  assign n1782 = ~n1780 & ~n1781 ;
  assign n1783 = \A[966]  & n1782 ;
  assign n1784 = ~n1780 & ~n1783 ;
  assign n1785 = \A[961]  & \A[962]  ;
  assign n1786 = ~\A[961]  & ~\A[962]  ;
  assign n1787 = ~n1785 & ~n1786 ;
  assign n1788 = \A[963]  & n1787 ;
  assign n1789 = ~n1785 & ~n1788 ;
  assign n1790 = n1784 & n1789 ;
  assign n1791 = ~n1784 & ~n1789 ;
  assign n1792 = ~\A[963]  & ~n1787 ;
  assign n1793 = ~n1788 & ~n1792 ;
  assign n1794 = ~\A[966]  & ~n1782 ;
  assign n1795 = ~n1783 & ~n1794 ;
  assign n1796 = n1793 & n1795 ;
  assign n1797 = ~n1791 & ~n1796 ;
  assign n1798 = ~n1790 & ~n1797 ;
  assign n1799 = ~n1793 & ~n1795 ;
  assign n1800 = ~n1796 & ~n1799 ;
  assign n1801 = ~n1767 & ~n1772 ;
  assign n1802 = ~n1773 & ~n1801 ;
  assign n1803 = n1800 & n1802 ;
  assign n1804 = n1774 & ~n1775 ;
  assign n1805 = n1803 & ~n1804 ;
  assign n1806 = ~n1790 & ~n1791 ;
  assign n1807 = n1796 & ~n1806 ;
  assign n1808 = ~n1796 & n1806 ;
  assign n1809 = ~n1807 & ~n1808 ;
  assign n1810 = n1805 & ~n1809 ;
  assign n1811 = ~n1805 & n1809 ;
  assign n1812 = ~n1774 & ~n1777 ;
  assign n1813 = n1775 & ~n1812 ;
  assign n1814 = ~n1775 & n1812 ;
  assign n1815 = ~n1813 & ~n1814 ;
  assign n1816 = ~n1811 & n1815 ;
  assign n1817 = ~n1810 & ~n1816 ;
  assign n1818 = n1798 & ~n1817 ;
  assign n1819 = ~n1798 & n1817 ;
  assign n1820 = ~n1818 & ~n1819 ;
  assign n1821 = n1779 & n1820 ;
  assign n1822 = ~n1779 & ~n1820 ;
  assign n1823 = ~n1821 & ~n1822 ;
  assign n1824 = ~n1760 & ~n1823 ;
  assign n1825 = n1760 & n1823 ;
  assign n1826 = ~n1800 & ~n1802 ;
  assign n1827 = ~n1803 & ~n1826 ;
  assign n1828 = ~n1737 & ~n1739 ;
  assign n1829 = ~n1740 & ~n1828 ;
  assign n1830 = n1827 & n1829 ;
  assign n1831 = ~n1810 & ~n1811 ;
  assign n1832 = n1815 & n1831 ;
  assign n1833 = ~n1815 & ~n1831 ;
  assign n1834 = ~n1832 & ~n1833 ;
  assign n1835 = n1830 & n1834 ;
  assign n1836 = ~n1830 & ~n1834 ;
  assign n1837 = ~n1747 & ~n1748 ;
  assign n1838 = n1752 & n1837 ;
  assign n1839 = ~n1752 & ~n1837 ;
  assign n1840 = ~n1838 & ~n1839 ;
  assign n1841 = ~n1836 & n1840 ;
  assign n1842 = ~n1835 & ~n1841 ;
  assign n1843 = ~n1825 & ~n1842 ;
  assign n1844 = ~n1824 & ~n1843 ;
  assign n1845 = ~n1779 & ~n1819 ;
  assign n1846 = ~n1818 & ~n1845 ;
  assign n1847 = ~n1844 & ~n1846 ;
  assign n1848 = n1844 & n1846 ;
  assign n1849 = ~n1716 & ~n1756 ;
  assign n1850 = ~n1755 & ~n1849 ;
  assign n1851 = ~n1848 & ~n1850 ;
  assign n1852 = ~n1847 & ~n1851 ;
  assign n1853 = \A[979]  & \A[980]  ;
  assign n1854 = ~\A[979]  & ~\A[980]  ;
  assign n1855 = ~n1853 & ~n1854 ;
  assign n1856 = \A[981]  & n1855 ;
  assign n1857 = ~\A[981]  & ~n1855 ;
  assign n1858 = ~n1856 & ~n1857 ;
  assign n1859 = \A[982]  & \A[983]  ;
  assign n1860 = ~\A[982]  & ~\A[983]  ;
  assign n1861 = ~n1859 & ~n1860 ;
  assign n1862 = \A[984]  & n1861 ;
  assign n1863 = ~\A[984]  & ~n1861 ;
  assign n1864 = ~n1862 & ~n1863 ;
  assign n1865 = n1858 & n1864 ;
  assign n1866 = ~n1858 & ~n1864 ;
  assign n1867 = ~n1865 & ~n1866 ;
  assign n1868 = \A[985]  & \A[986]  ;
  assign n1869 = ~\A[985]  & ~\A[986]  ;
  assign n1870 = ~n1868 & ~n1869 ;
  assign n1871 = \A[987]  & n1870 ;
  assign n1872 = ~\A[987]  & ~n1870 ;
  assign n1873 = ~n1871 & ~n1872 ;
  assign n1874 = \A[988]  & \A[989]  ;
  assign n1875 = ~\A[988]  & ~\A[989]  ;
  assign n1876 = ~n1874 & ~n1875 ;
  assign n1877 = \A[990]  & n1876 ;
  assign n1878 = ~\A[990]  & ~n1876 ;
  assign n1879 = ~n1877 & ~n1878 ;
  assign n1880 = n1873 & n1879 ;
  assign n1881 = ~n1873 & ~n1879 ;
  assign n1882 = ~n1880 & ~n1881 ;
  assign n1883 = n1867 & n1882 ;
  assign n1884 = ~n1874 & ~n1877 ;
  assign n1885 = ~n1868 & ~n1871 ;
  assign n1886 = n1884 & n1885 ;
  assign n1887 = ~n1884 & ~n1885 ;
  assign n1888 = ~n1886 & ~n1887 ;
  assign n1889 = n1883 & n1888 ;
  assign n1890 = ~n1859 & ~n1862 ;
  assign n1891 = ~n1853 & ~n1856 ;
  assign n1892 = ~n1890 & ~n1891 ;
  assign n1893 = n1890 & n1891 ;
  assign n1894 = ~n1892 & ~n1893 ;
  assign n1895 = n1865 & ~n1894 ;
  assign n1896 = ~n1865 & n1894 ;
  assign n1897 = ~n1895 & ~n1896 ;
  assign n1898 = ~n1889 & n1897 ;
  assign n1900 = n1880 & ~n1888 ;
  assign n1899 = ~n1880 & n1888 ;
  assign n1901 = ~n1883 & ~n1899 ;
  assign n1902 = ~n1900 & n1901 ;
  assign n1903 = ~n1898 & ~n1902 ;
  assign n1904 = n1880 & ~n1886 ;
  assign n1905 = ~n1887 & ~n1904 ;
  assign n1906 = ~n1903 & n1905 ;
  assign n1907 = n1903 & ~n1905 ;
  assign n1908 = ~n1865 & ~n1892 ;
  assign n1909 = ~n1893 & ~n1908 ;
  assign n1910 = ~n1907 & ~n1909 ;
  assign n1911 = ~n1906 & ~n1910 ;
  assign n1912 = \A[967]  & \A[968]  ;
  assign n1913 = ~\A[967]  & ~\A[968]  ;
  assign n1914 = ~n1912 & ~n1913 ;
  assign n1915 = \A[969]  & n1914 ;
  assign n1916 = ~\A[969]  & ~n1914 ;
  assign n1917 = ~n1915 & ~n1916 ;
  assign n1918 = \A[970]  & \A[971]  ;
  assign n1919 = ~\A[970]  & ~\A[971]  ;
  assign n1920 = ~n1918 & ~n1919 ;
  assign n1921 = \A[972]  & n1920 ;
  assign n1922 = ~\A[972]  & ~n1920 ;
  assign n1923 = ~n1921 & ~n1922 ;
  assign n1924 = n1917 & n1923 ;
  assign n1925 = ~n1917 & ~n1923 ;
  assign n1926 = ~n1924 & ~n1925 ;
  assign n1927 = \A[973]  & \A[974]  ;
  assign n1928 = ~\A[973]  & ~\A[974]  ;
  assign n1929 = ~n1927 & ~n1928 ;
  assign n1930 = \A[975]  & n1929 ;
  assign n1931 = ~\A[975]  & ~n1929 ;
  assign n1932 = ~n1930 & ~n1931 ;
  assign n1933 = \A[976]  & \A[977]  ;
  assign n1934 = ~\A[976]  & ~\A[977]  ;
  assign n1935 = ~n1933 & ~n1934 ;
  assign n1936 = \A[978]  & n1935 ;
  assign n1937 = ~\A[978]  & ~n1935 ;
  assign n1938 = ~n1936 & ~n1937 ;
  assign n1939 = n1932 & n1938 ;
  assign n1940 = ~n1932 & ~n1938 ;
  assign n1941 = ~n1939 & ~n1940 ;
  assign n1942 = n1926 & n1941 ;
  assign n1943 = ~n1933 & ~n1936 ;
  assign n1944 = ~n1927 & ~n1930 ;
  assign n1945 = n1943 & n1944 ;
  assign n1946 = ~n1943 & ~n1944 ;
  assign n1947 = ~n1945 & ~n1946 ;
  assign n1948 = n1942 & n1947 ;
  assign n1949 = ~n1918 & ~n1921 ;
  assign n1950 = ~n1912 & ~n1915 ;
  assign n1951 = ~n1949 & ~n1950 ;
  assign n1952 = n1949 & n1950 ;
  assign n1953 = ~n1951 & ~n1952 ;
  assign n1954 = n1924 & ~n1953 ;
  assign n1955 = ~n1924 & n1953 ;
  assign n1956 = ~n1954 & ~n1955 ;
  assign n1957 = ~n1948 & n1956 ;
  assign n1959 = n1939 & ~n1947 ;
  assign n1958 = ~n1939 & n1947 ;
  assign n1960 = ~n1942 & ~n1958 ;
  assign n1961 = ~n1959 & n1960 ;
  assign n1962 = ~n1957 & ~n1961 ;
  assign n1963 = n1939 & ~n1945 ;
  assign n1964 = ~n1946 & ~n1963 ;
  assign n1965 = ~n1962 & n1964 ;
  assign n1966 = n1962 & ~n1964 ;
  assign n1967 = ~n1924 & ~n1951 ;
  assign n1968 = ~n1952 & ~n1967 ;
  assign n1969 = ~n1966 & ~n1968 ;
  assign n1970 = ~n1965 & ~n1969 ;
  assign n1971 = n1911 & n1970 ;
  assign n1972 = ~n1911 & ~n1970 ;
  assign n1973 = ~n1965 & ~n1966 ;
  assign n1974 = ~n1968 & n1973 ;
  assign n1975 = n1968 & ~n1973 ;
  assign n1976 = ~n1974 & ~n1975 ;
  assign n1977 = ~n1906 & ~n1907 ;
  assign n1978 = ~n1909 & n1977 ;
  assign n1979 = n1909 & ~n1977 ;
  assign n1980 = ~n1978 & ~n1979 ;
  assign n1981 = ~n1976 & ~n1980 ;
  assign n1982 = n1976 & n1980 ;
  assign n1983 = ~n1867 & ~n1882 ;
  assign n1984 = ~n1883 & ~n1983 ;
  assign n1985 = ~n1926 & ~n1941 ;
  assign n1986 = ~n1942 & ~n1985 ;
  assign n1987 = n1984 & n1986 ;
  assign n1988 = ~n1889 & ~n1902 ;
  assign n1989 = n1897 & n1988 ;
  assign n1990 = ~n1897 & ~n1988 ;
  assign n1991 = ~n1989 & ~n1990 ;
  assign n1992 = n1987 & ~n1991 ;
  assign n1993 = ~n1987 & n1991 ;
  assign n1994 = ~n1948 & ~n1961 ;
  assign n1995 = n1956 & n1994 ;
  assign n1996 = ~n1956 & ~n1994 ;
  assign n1997 = ~n1995 & ~n1996 ;
  assign n1998 = ~n1993 & ~n1997 ;
  assign n1999 = ~n1992 & ~n1998 ;
  assign n2000 = ~n1982 & ~n1999 ;
  assign n2001 = ~n1981 & ~n2000 ;
  assign n2002 = ~n1972 & ~n2001 ;
  assign n2003 = ~n1971 & ~n2002 ;
  assign n2004 = ~n1852 & ~n2003 ;
  assign n2005 = n1852 & n2003 ;
  assign n2006 = ~n1847 & ~n1848 ;
  assign n2007 = ~n1850 & n2006 ;
  assign n2008 = n1850 & ~n2006 ;
  assign n2009 = ~n2007 & ~n2008 ;
  assign n2010 = ~n1971 & ~n1972 ;
  assign n2011 = ~n2001 & n2010 ;
  assign n2012 = n2001 & ~n2010 ;
  assign n2013 = ~n2011 & ~n2012 ;
  assign n2014 = n2009 & n2013 ;
  assign n2015 = ~n2009 & ~n2013 ;
  assign n2016 = ~n1824 & ~n1825 ;
  assign n2017 = ~n1842 & n2016 ;
  assign n2018 = n1842 & ~n2016 ;
  assign n2019 = ~n2017 & ~n2018 ;
  assign n2020 = ~n1981 & ~n1982 ;
  assign n2021 = ~n1999 & n2020 ;
  assign n2022 = n1999 & ~n2020 ;
  assign n2023 = ~n2021 & ~n2022 ;
  assign n2024 = n2019 & n2023 ;
  assign n2025 = ~n2019 & ~n2023 ;
  assign n2026 = ~n1984 & ~n1986 ;
  assign n2027 = ~n1987 & ~n2026 ;
  assign n2028 = ~n1827 & ~n1829 ;
  assign n2029 = ~n1830 & ~n2028 ;
  assign n2030 = n2027 & n2029 ;
  assign n2031 = ~n1992 & ~n1993 ;
  assign n2032 = ~n1997 & n2031 ;
  assign n2033 = n1997 & ~n2031 ;
  assign n2034 = ~n2032 & ~n2033 ;
  assign n2035 = n2030 & n2034 ;
  assign n2036 = ~n2030 & ~n2034 ;
  assign n2037 = ~n1835 & ~n1836 ;
  assign n2038 = ~n1840 & n2037 ;
  assign n2039 = n1840 & ~n2037 ;
  assign n2040 = ~n2038 & ~n2039 ;
  assign n2041 = ~n2036 & ~n2040 ;
  assign n2042 = ~n2035 & ~n2041 ;
  assign n2043 = ~n2025 & ~n2042 ;
  assign n2044 = ~n2024 & ~n2043 ;
  assign n2045 = ~n2015 & ~n2044 ;
  assign n2046 = ~n2014 & ~n2045 ;
  assign n2047 = ~n2005 & ~n2046 ;
  assign n2048 = ~n2004 & ~n2047 ;
  assign n2049 = n1697 & ~n2048 ;
  assign n2050 = ~n1697 & n2048 ;
  assign n2051 = ~n2004 & ~n2005 ;
  assign n2052 = ~n2046 & n2051 ;
  assign n2053 = n2046 & ~n2051 ;
  assign n2054 = ~n2052 & ~n2053 ;
  assign n2055 = ~n1650 & ~n1651 ;
  assign n2056 = ~n1692 & n2055 ;
  assign n2057 = n1692 & ~n2055 ;
  assign n2058 = ~n2056 & ~n2057 ;
  assign n2059 = ~n2054 & ~n2058 ;
  assign n2060 = n2054 & n2058 ;
  assign n2061 = ~n1660 & ~n1661 ;
  assign n2062 = n1690 & n2061 ;
  assign n2063 = ~n1690 & ~n2061 ;
  assign n2064 = ~n2062 & ~n2063 ;
  assign n2065 = ~n2014 & ~n2015 ;
  assign n2066 = ~n2044 & n2065 ;
  assign n2067 = n2044 & ~n2065 ;
  assign n2068 = ~n2066 & ~n2067 ;
  assign n2069 = ~n2064 & ~n2068 ;
  assign n2070 = n2064 & n2068 ;
  assign n2071 = ~n2024 & ~n2025 ;
  assign n2072 = ~n2042 & n2071 ;
  assign n2073 = n2042 & ~n2071 ;
  assign n2074 = ~n2072 & ~n2073 ;
  assign n2075 = ~n1670 & ~n1671 ;
  assign n2076 = ~n1688 & n2075 ;
  assign n2077 = n1688 & ~n2075 ;
  assign n2078 = ~n2076 & ~n2077 ;
  assign n2079 = ~n2074 & ~n2078 ;
  assign n2080 = n2074 & n2078 ;
  assign n2081 = ~n1673 & ~n1675 ;
  assign n2082 = ~n1676 & ~n2081 ;
  assign n2083 = ~n2027 & ~n2029 ;
  assign n2084 = ~n2030 & ~n2083 ;
  assign n2085 = n2082 & n2084 ;
  assign n2086 = ~n1681 & ~n1682 ;
  assign n2087 = ~n1686 & n2086 ;
  assign n2088 = n1686 & ~n2086 ;
  assign n2089 = ~n2087 & ~n2088 ;
  assign n2090 = n2085 & ~n2089 ;
  assign n2091 = ~n2085 & n2089 ;
  assign n2092 = ~n2035 & ~n2036 ;
  assign n2093 = ~n2040 & n2092 ;
  assign n2094 = n2040 & ~n2092 ;
  assign n2095 = ~n2093 & ~n2094 ;
  assign n2096 = ~n2091 & n2095 ;
  assign n2097 = ~n2090 & ~n2096 ;
  assign n2098 = ~n2080 & n2097 ;
  assign n2099 = ~n2079 & ~n2098 ;
  assign n2100 = ~n2070 & ~n2099 ;
  assign n2101 = ~n2069 & ~n2100 ;
  assign n2102 = ~n2060 & ~n2101 ;
  assign n2103 = ~n2059 & ~n2102 ;
  assign n2104 = ~n2050 & n2103 ;
  assign n2105 = ~n2049 & ~n2104 ;
  assign n2106 = ~n1639 & ~n1694 ;
  assign n2107 = ~n1640 & ~n2106 ;
  assign n2108 = ~n2105 & ~n2107 ;
  assign n2109 = n2105 & n2107 ;
  assign n2110 = ~n2108 & ~n2109 ;
  assign n2111 = \A[874]  & \A[875]  ;
  assign n2112 = \A[871]  & \A[872]  ;
  assign n2113 = ~\A[871]  & ~\A[872]  ;
  assign n2114 = ~n2112 & ~n2113 ;
  assign n2115 = \A[873]  & n2114 ;
  assign n2116 = ~\A[873]  & ~n2114 ;
  assign n2117 = ~n2115 & ~n2116 ;
  assign n2118 = ~\A[874]  & ~\A[875]  ;
  assign n2119 = ~n2111 & ~n2118 ;
  assign n2120 = \A[876]  & n2119 ;
  assign n2121 = ~\A[876]  & ~n2119 ;
  assign n2122 = ~n2120 & ~n2121 ;
  assign n2123 = n2117 & n2122 ;
  assign n2124 = n2111 & n2123 ;
  assign n2125 = ~n2112 & ~n2115 ;
  assign n2126 = ~n2111 & ~n2120 ;
  assign n2127 = ~n2123 & n2126 ;
  assign n2128 = ~n2125 & ~n2127 ;
  assign n2129 = ~n2124 & ~n2128 ;
  assign n2130 = \A[880]  & \A[881]  ;
  assign n2131 = ~\A[880]  & ~\A[881]  ;
  assign n2132 = ~n2130 & ~n2131 ;
  assign n2133 = \A[882]  & n2132 ;
  assign n2134 = ~n2130 & ~n2133 ;
  assign n2135 = \A[877]  & \A[878]  ;
  assign n2136 = ~\A[877]  & ~\A[878]  ;
  assign n2137 = ~n2135 & ~n2136 ;
  assign n2138 = \A[879]  & n2137 ;
  assign n2139 = ~n2135 & ~n2138 ;
  assign n2140 = n2134 & n2139 ;
  assign n2141 = ~n2134 & ~n2139 ;
  assign n2142 = ~\A[879]  & ~n2137 ;
  assign n2143 = ~n2138 & ~n2142 ;
  assign n2144 = ~\A[882]  & ~n2132 ;
  assign n2145 = ~n2133 & ~n2144 ;
  assign n2146 = n2143 & n2145 ;
  assign n2147 = ~n2141 & ~n2146 ;
  assign n2148 = ~n2140 & ~n2147 ;
  assign n2149 = ~n2143 & ~n2145 ;
  assign n2150 = ~n2146 & ~n2149 ;
  assign n2151 = ~n2117 & ~n2122 ;
  assign n2152 = ~n2123 & ~n2151 ;
  assign n2153 = n2150 & n2152 ;
  assign n2154 = n2124 & ~n2125 ;
  assign n2155 = n2153 & ~n2154 ;
  assign n2156 = ~n2140 & ~n2141 ;
  assign n2157 = n2146 & ~n2156 ;
  assign n2158 = ~n2146 & n2156 ;
  assign n2159 = ~n2157 & ~n2158 ;
  assign n2160 = n2155 & ~n2159 ;
  assign n2161 = ~n2155 & n2159 ;
  assign n2162 = ~n2124 & ~n2127 ;
  assign n2163 = n2125 & ~n2162 ;
  assign n2164 = ~n2125 & n2162 ;
  assign n2165 = ~n2163 & ~n2164 ;
  assign n2166 = ~n2161 & n2165 ;
  assign n2167 = ~n2160 & ~n2166 ;
  assign n2168 = n2148 & ~n2167 ;
  assign n2169 = ~n2148 & n2167 ;
  assign n2170 = ~n2168 & ~n2169 ;
  assign n2171 = n2129 & n2170 ;
  assign n2172 = ~n2129 & ~n2170 ;
  assign n2173 = ~n2171 & ~n2172 ;
  assign n2174 = \A[886]  & \A[887]  ;
  assign n2175 = \A[883]  & \A[884]  ;
  assign n2176 = ~\A[883]  & ~\A[884]  ;
  assign n2177 = ~n2175 & ~n2176 ;
  assign n2178 = \A[885]  & n2177 ;
  assign n2179 = ~\A[885]  & ~n2177 ;
  assign n2180 = ~n2178 & ~n2179 ;
  assign n2181 = ~\A[886]  & ~\A[887]  ;
  assign n2182 = ~n2174 & ~n2181 ;
  assign n2183 = \A[888]  & n2182 ;
  assign n2184 = ~\A[888]  & ~n2182 ;
  assign n2185 = ~n2183 & ~n2184 ;
  assign n2186 = n2180 & n2185 ;
  assign n2187 = n2174 & n2186 ;
  assign n2188 = ~n2175 & ~n2178 ;
  assign n2189 = ~n2174 & ~n2183 ;
  assign n2190 = ~n2186 & n2189 ;
  assign n2191 = ~n2188 & ~n2190 ;
  assign n2192 = ~n2187 & ~n2191 ;
  assign n2193 = \A[892]  & \A[893]  ;
  assign n2194 = ~\A[892]  & ~\A[893]  ;
  assign n2195 = ~n2193 & ~n2194 ;
  assign n2196 = \A[894]  & n2195 ;
  assign n2197 = ~n2193 & ~n2196 ;
  assign n2198 = \A[889]  & \A[890]  ;
  assign n2199 = ~\A[889]  & ~\A[890]  ;
  assign n2200 = ~n2198 & ~n2199 ;
  assign n2201 = \A[891]  & n2200 ;
  assign n2202 = ~n2198 & ~n2201 ;
  assign n2203 = n2197 & n2202 ;
  assign n2204 = ~n2197 & ~n2202 ;
  assign n2205 = ~\A[891]  & ~n2200 ;
  assign n2206 = ~n2201 & ~n2205 ;
  assign n2207 = ~\A[894]  & ~n2195 ;
  assign n2208 = ~n2196 & ~n2207 ;
  assign n2209 = n2206 & n2208 ;
  assign n2210 = ~n2204 & ~n2209 ;
  assign n2211 = ~n2203 & ~n2210 ;
  assign n2212 = ~n2206 & ~n2208 ;
  assign n2213 = ~n2209 & ~n2212 ;
  assign n2214 = ~n2180 & ~n2185 ;
  assign n2215 = ~n2186 & ~n2214 ;
  assign n2216 = n2213 & n2215 ;
  assign n2217 = n2187 & ~n2188 ;
  assign n2218 = n2216 & ~n2217 ;
  assign n2219 = ~n2203 & ~n2204 ;
  assign n2220 = n2209 & ~n2219 ;
  assign n2221 = ~n2209 & n2219 ;
  assign n2222 = ~n2220 & ~n2221 ;
  assign n2223 = n2218 & ~n2222 ;
  assign n2224 = ~n2218 & n2222 ;
  assign n2225 = ~n2187 & ~n2190 ;
  assign n2226 = n2188 & ~n2225 ;
  assign n2227 = ~n2188 & n2225 ;
  assign n2228 = ~n2226 & ~n2227 ;
  assign n2229 = ~n2224 & n2228 ;
  assign n2230 = ~n2223 & ~n2229 ;
  assign n2231 = n2211 & ~n2230 ;
  assign n2232 = ~n2211 & n2230 ;
  assign n2233 = ~n2231 & ~n2232 ;
  assign n2234 = n2192 & n2233 ;
  assign n2235 = ~n2192 & ~n2233 ;
  assign n2236 = ~n2234 & ~n2235 ;
  assign n2237 = ~n2173 & ~n2236 ;
  assign n2238 = n2173 & n2236 ;
  assign n2239 = ~n2213 & ~n2215 ;
  assign n2240 = ~n2216 & ~n2239 ;
  assign n2241 = ~n2150 & ~n2152 ;
  assign n2242 = ~n2153 & ~n2241 ;
  assign n2243 = n2240 & n2242 ;
  assign n2244 = ~n2223 & ~n2224 ;
  assign n2245 = n2228 & n2244 ;
  assign n2246 = ~n2228 & ~n2244 ;
  assign n2247 = ~n2245 & ~n2246 ;
  assign n2248 = n2243 & n2247 ;
  assign n2249 = ~n2243 & ~n2247 ;
  assign n2250 = ~n2160 & ~n2161 ;
  assign n2251 = n2165 & n2250 ;
  assign n2252 = ~n2165 & ~n2250 ;
  assign n2253 = ~n2251 & ~n2252 ;
  assign n2254 = ~n2249 & n2253 ;
  assign n2255 = ~n2248 & ~n2254 ;
  assign n2256 = ~n2238 & ~n2255 ;
  assign n2257 = ~n2237 & ~n2256 ;
  assign n2258 = ~n2192 & ~n2232 ;
  assign n2259 = ~n2231 & ~n2258 ;
  assign n2260 = ~n2257 & ~n2259 ;
  assign n2261 = n2257 & n2259 ;
  assign n2262 = ~n2129 & ~n2169 ;
  assign n2263 = ~n2168 & ~n2262 ;
  assign n2264 = ~n2261 & ~n2263 ;
  assign n2265 = ~n2260 & ~n2264 ;
  assign n2266 = ~n2260 & ~n2261 ;
  assign n2267 = ~n2263 & n2266 ;
  assign n2268 = n2263 & ~n2266 ;
  assign n2269 = ~n2267 & ~n2268 ;
  assign n2270 = \A[850]  & \A[851]  ;
  assign n2271 = \A[847]  & \A[848]  ;
  assign n2272 = ~\A[847]  & ~\A[848]  ;
  assign n2273 = ~n2271 & ~n2272 ;
  assign n2274 = \A[849]  & n2273 ;
  assign n2275 = ~\A[849]  & ~n2273 ;
  assign n2276 = ~n2274 & ~n2275 ;
  assign n2277 = ~\A[850]  & ~\A[851]  ;
  assign n2278 = ~n2270 & ~n2277 ;
  assign n2279 = \A[852]  & n2278 ;
  assign n2280 = ~\A[852]  & ~n2278 ;
  assign n2281 = ~n2279 & ~n2280 ;
  assign n2282 = n2276 & n2281 ;
  assign n2283 = n2270 & n2282 ;
  assign n2284 = ~n2271 & ~n2274 ;
  assign n2285 = ~n2270 & ~n2279 ;
  assign n2286 = ~n2282 & n2285 ;
  assign n2287 = ~n2284 & ~n2286 ;
  assign n2288 = ~n2283 & ~n2287 ;
  assign n2289 = \A[856]  & \A[857]  ;
  assign n2290 = ~\A[856]  & ~\A[857]  ;
  assign n2291 = ~n2289 & ~n2290 ;
  assign n2292 = \A[858]  & n2291 ;
  assign n2293 = ~n2289 & ~n2292 ;
  assign n2294 = \A[853]  & \A[854]  ;
  assign n2295 = ~\A[853]  & ~\A[854]  ;
  assign n2296 = ~n2294 & ~n2295 ;
  assign n2297 = \A[855]  & n2296 ;
  assign n2298 = ~n2294 & ~n2297 ;
  assign n2299 = n2293 & n2298 ;
  assign n2300 = ~n2293 & ~n2298 ;
  assign n2301 = ~\A[855]  & ~n2296 ;
  assign n2302 = ~n2297 & ~n2301 ;
  assign n2303 = ~\A[858]  & ~n2291 ;
  assign n2304 = ~n2292 & ~n2303 ;
  assign n2305 = n2302 & n2304 ;
  assign n2306 = ~n2300 & ~n2305 ;
  assign n2307 = ~n2299 & ~n2306 ;
  assign n2308 = ~n2302 & ~n2304 ;
  assign n2309 = ~n2305 & ~n2308 ;
  assign n2310 = ~n2276 & ~n2281 ;
  assign n2311 = ~n2282 & ~n2310 ;
  assign n2312 = n2309 & n2311 ;
  assign n2313 = n2283 & ~n2284 ;
  assign n2314 = n2312 & ~n2313 ;
  assign n2315 = ~n2299 & ~n2300 ;
  assign n2316 = n2305 & ~n2315 ;
  assign n2317 = ~n2305 & n2315 ;
  assign n2318 = ~n2316 & ~n2317 ;
  assign n2319 = n2314 & ~n2318 ;
  assign n2320 = ~n2314 & n2318 ;
  assign n2321 = ~n2283 & ~n2286 ;
  assign n2322 = n2284 & ~n2321 ;
  assign n2323 = ~n2284 & n2321 ;
  assign n2324 = ~n2322 & ~n2323 ;
  assign n2325 = ~n2320 & n2324 ;
  assign n2326 = ~n2319 & ~n2325 ;
  assign n2327 = n2307 & ~n2326 ;
  assign n2328 = ~n2307 & n2326 ;
  assign n2329 = ~n2327 & ~n2328 ;
  assign n2330 = n2288 & n2329 ;
  assign n2331 = ~n2288 & ~n2329 ;
  assign n2332 = ~n2330 & ~n2331 ;
  assign n2333 = \A[862]  & \A[863]  ;
  assign n2334 = \A[859]  & \A[860]  ;
  assign n2335 = ~\A[859]  & ~\A[860]  ;
  assign n2336 = ~n2334 & ~n2335 ;
  assign n2337 = \A[861]  & n2336 ;
  assign n2338 = ~\A[861]  & ~n2336 ;
  assign n2339 = ~n2337 & ~n2338 ;
  assign n2340 = ~\A[862]  & ~\A[863]  ;
  assign n2341 = ~n2333 & ~n2340 ;
  assign n2342 = \A[864]  & n2341 ;
  assign n2343 = ~\A[864]  & ~n2341 ;
  assign n2344 = ~n2342 & ~n2343 ;
  assign n2345 = n2339 & n2344 ;
  assign n2346 = n2333 & n2345 ;
  assign n2347 = ~n2334 & ~n2337 ;
  assign n2348 = ~n2333 & ~n2342 ;
  assign n2349 = ~n2345 & n2348 ;
  assign n2350 = ~n2347 & ~n2349 ;
  assign n2351 = ~n2346 & ~n2350 ;
  assign n2352 = \A[868]  & \A[869]  ;
  assign n2353 = ~\A[868]  & ~\A[869]  ;
  assign n2354 = ~n2352 & ~n2353 ;
  assign n2355 = \A[870]  & n2354 ;
  assign n2356 = ~n2352 & ~n2355 ;
  assign n2357 = \A[865]  & \A[866]  ;
  assign n2358 = ~\A[865]  & ~\A[866]  ;
  assign n2359 = ~n2357 & ~n2358 ;
  assign n2360 = \A[867]  & n2359 ;
  assign n2361 = ~n2357 & ~n2360 ;
  assign n2362 = n2356 & n2361 ;
  assign n2363 = ~n2356 & ~n2361 ;
  assign n2364 = ~\A[867]  & ~n2359 ;
  assign n2365 = ~n2360 & ~n2364 ;
  assign n2366 = ~\A[870]  & ~n2354 ;
  assign n2367 = ~n2355 & ~n2366 ;
  assign n2368 = n2365 & n2367 ;
  assign n2369 = ~n2363 & ~n2368 ;
  assign n2370 = ~n2362 & ~n2369 ;
  assign n2371 = ~n2365 & ~n2367 ;
  assign n2372 = ~n2368 & ~n2371 ;
  assign n2373 = ~n2339 & ~n2344 ;
  assign n2374 = ~n2345 & ~n2373 ;
  assign n2375 = n2372 & n2374 ;
  assign n2376 = n2346 & ~n2347 ;
  assign n2377 = n2375 & ~n2376 ;
  assign n2378 = ~n2362 & ~n2363 ;
  assign n2379 = n2368 & ~n2378 ;
  assign n2380 = ~n2368 & n2378 ;
  assign n2381 = ~n2379 & ~n2380 ;
  assign n2382 = n2377 & ~n2381 ;
  assign n2383 = ~n2377 & n2381 ;
  assign n2384 = ~n2346 & ~n2349 ;
  assign n2385 = n2347 & ~n2384 ;
  assign n2386 = ~n2347 & n2384 ;
  assign n2387 = ~n2385 & ~n2386 ;
  assign n2388 = ~n2383 & n2387 ;
  assign n2389 = ~n2382 & ~n2388 ;
  assign n2390 = n2370 & ~n2389 ;
  assign n2391 = ~n2370 & n2389 ;
  assign n2392 = ~n2390 & ~n2391 ;
  assign n2393 = n2351 & n2392 ;
  assign n2394 = ~n2351 & ~n2392 ;
  assign n2395 = ~n2393 & ~n2394 ;
  assign n2396 = ~n2332 & ~n2395 ;
  assign n2397 = n2332 & n2395 ;
  assign n2398 = ~n2372 & ~n2374 ;
  assign n2399 = ~n2375 & ~n2398 ;
  assign n2400 = ~n2309 & ~n2311 ;
  assign n2401 = ~n2312 & ~n2400 ;
  assign n2402 = n2399 & n2401 ;
  assign n2403 = ~n2382 & ~n2383 ;
  assign n2404 = n2387 & n2403 ;
  assign n2405 = ~n2387 & ~n2403 ;
  assign n2406 = ~n2404 & ~n2405 ;
  assign n2407 = n2402 & n2406 ;
  assign n2408 = ~n2402 & ~n2406 ;
  assign n2409 = ~n2319 & ~n2320 ;
  assign n2410 = n2324 & n2409 ;
  assign n2411 = ~n2324 & ~n2409 ;
  assign n2412 = ~n2410 & ~n2411 ;
  assign n2413 = ~n2408 & n2412 ;
  assign n2414 = ~n2407 & ~n2413 ;
  assign n2415 = ~n2397 & ~n2414 ;
  assign n2416 = ~n2396 & ~n2415 ;
  assign n2417 = ~n2351 & ~n2391 ;
  assign n2418 = ~n2390 & ~n2417 ;
  assign n2419 = ~n2416 & ~n2418 ;
  assign n2420 = n2416 & n2418 ;
  assign n2421 = ~n2419 & ~n2420 ;
  assign n2422 = ~n2288 & ~n2328 ;
  assign n2423 = ~n2327 & ~n2422 ;
  assign n2424 = n2421 & ~n2423 ;
  assign n2425 = ~n2421 & n2423 ;
  assign n2426 = ~n2424 & ~n2425 ;
  assign n2427 = ~n2269 & ~n2426 ;
  assign n2428 = n2269 & n2426 ;
  assign n2429 = ~n2396 & ~n2397 ;
  assign n2430 = ~n2414 & n2429 ;
  assign n2431 = n2414 & ~n2429 ;
  assign n2432 = ~n2430 & ~n2431 ;
  assign n2433 = ~n2237 & ~n2238 ;
  assign n2434 = ~n2255 & n2433 ;
  assign n2435 = n2255 & ~n2433 ;
  assign n2436 = ~n2434 & ~n2435 ;
  assign n2437 = ~n2432 & ~n2436 ;
  assign n2438 = n2432 & n2436 ;
  assign n2439 = ~n2240 & ~n2242 ;
  assign n2440 = ~n2243 & ~n2439 ;
  assign n2441 = ~n2399 & ~n2401 ;
  assign n2442 = ~n2402 & ~n2441 ;
  assign n2443 = n2440 & n2442 ;
  assign n2444 = ~n2248 & ~n2249 ;
  assign n2445 = ~n2253 & n2444 ;
  assign n2446 = n2253 & ~n2444 ;
  assign n2447 = ~n2445 & ~n2446 ;
  assign n2448 = n2443 & ~n2447 ;
  assign n2449 = ~n2443 & n2447 ;
  assign n2450 = ~n2407 & ~n2408 ;
  assign n2451 = ~n2412 & n2450 ;
  assign n2452 = n2412 & ~n2450 ;
  assign n2453 = ~n2451 & ~n2452 ;
  assign n2454 = ~n2449 & ~n2453 ;
  assign n2455 = ~n2448 & ~n2454 ;
  assign n2456 = ~n2438 & n2455 ;
  assign n2457 = ~n2437 & ~n2456 ;
  assign n2458 = ~n2428 & ~n2457 ;
  assign n2459 = ~n2427 & ~n2458 ;
  assign n2460 = n2265 & ~n2459 ;
  assign n2461 = ~n2265 & n2459 ;
  assign n2462 = ~n2460 & ~n2461 ;
  assign n2463 = ~n2420 & ~n2423 ;
  assign n2464 = ~n2419 & ~n2463 ;
  assign n2465 = n2462 & n2464 ;
  assign n2466 = ~n2462 & ~n2464 ;
  assign n2467 = ~n2465 & ~n2466 ;
  assign n2468 = \A[922]  & \A[923]  ;
  assign n2469 = \A[919]  & \A[920]  ;
  assign n2470 = ~\A[919]  & ~\A[920]  ;
  assign n2471 = ~n2469 & ~n2470 ;
  assign n2472 = \A[921]  & n2471 ;
  assign n2473 = ~\A[921]  & ~n2471 ;
  assign n2474 = ~n2472 & ~n2473 ;
  assign n2475 = ~\A[922]  & ~\A[923]  ;
  assign n2476 = ~n2468 & ~n2475 ;
  assign n2477 = \A[924]  & n2476 ;
  assign n2478 = ~\A[924]  & ~n2476 ;
  assign n2479 = ~n2477 & ~n2478 ;
  assign n2480 = n2474 & n2479 ;
  assign n2481 = n2468 & n2480 ;
  assign n2482 = ~n2469 & ~n2472 ;
  assign n2483 = ~n2468 & ~n2477 ;
  assign n2484 = ~n2480 & n2483 ;
  assign n2485 = ~n2482 & ~n2484 ;
  assign n2486 = ~n2481 & ~n2485 ;
  assign n2487 = \A[928]  & \A[929]  ;
  assign n2488 = ~\A[928]  & ~\A[929]  ;
  assign n2489 = ~n2487 & ~n2488 ;
  assign n2490 = \A[930]  & n2489 ;
  assign n2491 = ~n2487 & ~n2490 ;
  assign n2492 = \A[925]  & \A[926]  ;
  assign n2493 = ~\A[925]  & ~\A[926]  ;
  assign n2494 = ~n2492 & ~n2493 ;
  assign n2495 = \A[927]  & n2494 ;
  assign n2496 = ~n2492 & ~n2495 ;
  assign n2497 = n2491 & n2496 ;
  assign n2498 = ~n2491 & ~n2496 ;
  assign n2499 = ~\A[927]  & ~n2494 ;
  assign n2500 = ~n2495 & ~n2499 ;
  assign n2501 = ~\A[930]  & ~n2489 ;
  assign n2502 = ~n2490 & ~n2501 ;
  assign n2503 = n2500 & n2502 ;
  assign n2504 = ~n2498 & ~n2503 ;
  assign n2505 = ~n2497 & ~n2504 ;
  assign n2506 = ~n2500 & ~n2502 ;
  assign n2507 = ~n2503 & ~n2506 ;
  assign n2508 = ~n2474 & ~n2479 ;
  assign n2509 = ~n2480 & ~n2508 ;
  assign n2510 = n2507 & n2509 ;
  assign n2511 = n2481 & ~n2482 ;
  assign n2512 = n2510 & ~n2511 ;
  assign n2513 = ~n2497 & ~n2498 ;
  assign n2514 = n2503 & ~n2513 ;
  assign n2515 = ~n2503 & n2513 ;
  assign n2516 = ~n2514 & ~n2515 ;
  assign n2517 = n2512 & ~n2516 ;
  assign n2518 = ~n2512 & n2516 ;
  assign n2519 = ~n2481 & ~n2484 ;
  assign n2520 = n2482 & ~n2519 ;
  assign n2521 = ~n2482 & n2519 ;
  assign n2522 = ~n2520 & ~n2521 ;
  assign n2523 = ~n2518 & n2522 ;
  assign n2524 = ~n2517 & ~n2523 ;
  assign n2525 = n2505 & ~n2524 ;
  assign n2526 = ~n2505 & n2524 ;
  assign n2527 = ~n2525 & ~n2526 ;
  assign n2528 = n2486 & n2527 ;
  assign n2529 = ~n2486 & ~n2527 ;
  assign n2530 = ~n2528 & ~n2529 ;
  assign n2531 = \A[934]  & \A[935]  ;
  assign n2532 = \A[931]  & \A[932]  ;
  assign n2533 = ~\A[931]  & ~\A[932]  ;
  assign n2534 = ~n2532 & ~n2533 ;
  assign n2535 = \A[933]  & n2534 ;
  assign n2536 = ~\A[933]  & ~n2534 ;
  assign n2537 = ~n2535 & ~n2536 ;
  assign n2538 = ~\A[934]  & ~\A[935]  ;
  assign n2539 = ~n2531 & ~n2538 ;
  assign n2540 = \A[936]  & n2539 ;
  assign n2541 = ~\A[936]  & ~n2539 ;
  assign n2542 = ~n2540 & ~n2541 ;
  assign n2543 = n2537 & n2542 ;
  assign n2544 = n2531 & n2543 ;
  assign n2545 = ~n2532 & ~n2535 ;
  assign n2546 = ~n2531 & ~n2540 ;
  assign n2547 = ~n2543 & n2546 ;
  assign n2548 = ~n2545 & ~n2547 ;
  assign n2549 = ~n2544 & ~n2548 ;
  assign n2550 = \A[940]  & \A[941]  ;
  assign n2551 = ~\A[940]  & ~\A[941]  ;
  assign n2552 = ~n2550 & ~n2551 ;
  assign n2553 = \A[942]  & n2552 ;
  assign n2554 = ~n2550 & ~n2553 ;
  assign n2555 = \A[937]  & \A[938]  ;
  assign n2556 = ~\A[937]  & ~\A[938]  ;
  assign n2557 = ~n2555 & ~n2556 ;
  assign n2558 = \A[939]  & n2557 ;
  assign n2559 = ~n2555 & ~n2558 ;
  assign n2560 = n2554 & n2559 ;
  assign n2561 = ~n2554 & ~n2559 ;
  assign n2562 = ~\A[939]  & ~n2557 ;
  assign n2563 = ~n2558 & ~n2562 ;
  assign n2564 = ~\A[942]  & ~n2552 ;
  assign n2565 = ~n2553 & ~n2564 ;
  assign n2566 = n2563 & n2565 ;
  assign n2567 = ~n2561 & ~n2566 ;
  assign n2568 = ~n2560 & ~n2567 ;
  assign n2569 = ~n2563 & ~n2565 ;
  assign n2570 = ~n2566 & ~n2569 ;
  assign n2571 = ~n2537 & ~n2542 ;
  assign n2572 = ~n2543 & ~n2571 ;
  assign n2573 = n2570 & n2572 ;
  assign n2574 = n2544 & ~n2545 ;
  assign n2575 = n2573 & ~n2574 ;
  assign n2576 = ~n2560 & ~n2561 ;
  assign n2577 = n2566 & ~n2576 ;
  assign n2578 = ~n2566 & n2576 ;
  assign n2579 = ~n2577 & ~n2578 ;
  assign n2580 = n2575 & ~n2579 ;
  assign n2581 = ~n2575 & n2579 ;
  assign n2582 = ~n2544 & ~n2547 ;
  assign n2583 = n2545 & ~n2582 ;
  assign n2584 = ~n2545 & n2582 ;
  assign n2585 = ~n2583 & ~n2584 ;
  assign n2586 = ~n2581 & n2585 ;
  assign n2587 = ~n2580 & ~n2586 ;
  assign n2588 = n2568 & ~n2587 ;
  assign n2589 = ~n2568 & n2587 ;
  assign n2590 = ~n2588 & ~n2589 ;
  assign n2591 = n2549 & n2590 ;
  assign n2592 = ~n2549 & ~n2590 ;
  assign n2593 = ~n2591 & ~n2592 ;
  assign n2594 = ~n2530 & ~n2593 ;
  assign n2595 = n2530 & n2593 ;
  assign n2596 = ~n2570 & ~n2572 ;
  assign n2597 = ~n2573 & ~n2596 ;
  assign n2598 = ~n2507 & ~n2509 ;
  assign n2599 = ~n2510 & ~n2598 ;
  assign n2600 = n2597 & n2599 ;
  assign n2601 = ~n2580 & ~n2581 ;
  assign n2602 = n2585 & n2601 ;
  assign n2603 = ~n2585 & ~n2601 ;
  assign n2604 = ~n2602 & ~n2603 ;
  assign n2605 = n2600 & n2604 ;
  assign n2606 = ~n2600 & ~n2604 ;
  assign n2607 = ~n2517 & ~n2518 ;
  assign n2608 = n2522 & n2607 ;
  assign n2609 = ~n2522 & ~n2607 ;
  assign n2610 = ~n2608 & ~n2609 ;
  assign n2611 = ~n2606 & n2610 ;
  assign n2612 = ~n2605 & ~n2611 ;
  assign n2613 = ~n2595 & ~n2612 ;
  assign n2614 = ~n2594 & ~n2613 ;
  assign n2615 = ~n2549 & ~n2589 ;
  assign n2616 = ~n2588 & ~n2615 ;
  assign n2617 = ~n2614 & ~n2616 ;
  assign n2618 = n2614 & n2616 ;
  assign n2619 = ~n2486 & ~n2526 ;
  assign n2620 = ~n2525 & ~n2619 ;
  assign n2621 = ~n2618 & ~n2620 ;
  assign n2622 = ~n2617 & ~n2621 ;
  assign n2623 = ~n2617 & ~n2618 ;
  assign n2624 = ~n2620 & n2623 ;
  assign n2625 = n2620 & ~n2623 ;
  assign n2626 = ~n2624 & ~n2625 ;
  assign n2627 = \A[898]  & \A[899]  ;
  assign n2628 = \A[895]  & \A[896]  ;
  assign n2629 = ~\A[895]  & ~\A[896]  ;
  assign n2630 = ~n2628 & ~n2629 ;
  assign n2631 = \A[897]  & n2630 ;
  assign n2632 = ~\A[897]  & ~n2630 ;
  assign n2633 = ~n2631 & ~n2632 ;
  assign n2634 = ~\A[898]  & ~\A[899]  ;
  assign n2635 = ~n2627 & ~n2634 ;
  assign n2636 = \A[900]  & n2635 ;
  assign n2637 = ~\A[900]  & ~n2635 ;
  assign n2638 = ~n2636 & ~n2637 ;
  assign n2639 = n2633 & n2638 ;
  assign n2640 = n2627 & n2639 ;
  assign n2641 = ~n2628 & ~n2631 ;
  assign n2642 = ~n2627 & ~n2636 ;
  assign n2643 = ~n2639 & n2642 ;
  assign n2644 = ~n2641 & ~n2643 ;
  assign n2645 = ~n2640 & ~n2644 ;
  assign n2646 = \A[904]  & \A[905]  ;
  assign n2647 = ~\A[904]  & ~\A[905]  ;
  assign n2648 = ~n2646 & ~n2647 ;
  assign n2649 = \A[906]  & n2648 ;
  assign n2650 = ~n2646 & ~n2649 ;
  assign n2651 = \A[901]  & \A[902]  ;
  assign n2652 = ~\A[901]  & ~\A[902]  ;
  assign n2653 = ~n2651 & ~n2652 ;
  assign n2654 = \A[903]  & n2653 ;
  assign n2655 = ~n2651 & ~n2654 ;
  assign n2656 = n2650 & n2655 ;
  assign n2657 = ~n2650 & ~n2655 ;
  assign n2658 = ~\A[903]  & ~n2653 ;
  assign n2659 = ~n2654 & ~n2658 ;
  assign n2660 = ~\A[906]  & ~n2648 ;
  assign n2661 = ~n2649 & ~n2660 ;
  assign n2662 = n2659 & n2661 ;
  assign n2663 = ~n2657 & ~n2662 ;
  assign n2664 = ~n2656 & ~n2663 ;
  assign n2665 = ~n2659 & ~n2661 ;
  assign n2666 = ~n2662 & ~n2665 ;
  assign n2667 = ~n2633 & ~n2638 ;
  assign n2668 = ~n2639 & ~n2667 ;
  assign n2669 = n2666 & n2668 ;
  assign n2670 = n2640 & ~n2641 ;
  assign n2671 = n2669 & ~n2670 ;
  assign n2672 = ~n2656 & ~n2657 ;
  assign n2673 = n2662 & ~n2672 ;
  assign n2674 = ~n2662 & n2672 ;
  assign n2675 = ~n2673 & ~n2674 ;
  assign n2676 = n2671 & ~n2675 ;
  assign n2677 = ~n2671 & n2675 ;
  assign n2678 = ~n2640 & ~n2643 ;
  assign n2679 = n2641 & ~n2678 ;
  assign n2680 = ~n2641 & n2678 ;
  assign n2681 = ~n2679 & ~n2680 ;
  assign n2682 = ~n2677 & n2681 ;
  assign n2683 = ~n2676 & ~n2682 ;
  assign n2684 = n2664 & ~n2683 ;
  assign n2685 = ~n2664 & n2683 ;
  assign n2686 = ~n2684 & ~n2685 ;
  assign n2687 = n2645 & n2686 ;
  assign n2688 = ~n2645 & ~n2686 ;
  assign n2689 = ~n2687 & ~n2688 ;
  assign n2690 = \A[910]  & \A[911]  ;
  assign n2691 = \A[907]  & \A[908]  ;
  assign n2692 = ~\A[907]  & ~\A[908]  ;
  assign n2693 = ~n2691 & ~n2692 ;
  assign n2694 = \A[909]  & n2693 ;
  assign n2695 = ~\A[909]  & ~n2693 ;
  assign n2696 = ~n2694 & ~n2695 ;
  assign n2697 = ~\A[910]  & ~\A[911]  ;
  assign n2698 = ~n2690 & ~n2697 ;
  assign n2699 = \A[912]  & n2698 ;
  assign n2700 = ~\A[912]  & ~n2698 ;
  assign n2701 = ~n2699 & ~n2700 ;
  assign n2702 = n2696 & n2701 ;
  assign n2703 = n2690 & n2702 ;
  assign n2704 = ~n2691 & ~n2694 ;
  assign n2705 = ~n2690 & ~n2699 ;
  assign n2706 = ~n2702 & n2705 ;
  assign n2707 = ~n2704 & ~n2706 ;
  assign n2708 = ~n2703 & ~n2707 ;
  assign n2709 = \A[916]  & \A[917]  ;
  assign n2710 = ~\A[916]  & ~\A[917]  ;
  assign n2711 = ~n2709 & ~n2710 ;
  assign n2712 = \A[918]  & n2711 ;
  assign n2713 = ~n2709 & ~n2712 ;
  assign n2714 = \A[913]  & \A[914]  ;
  assign n2715 = ~\A[913]  & ~\A[914]  ;
  assign n2716 = ~n2714 & ~n2715 ;
  assign n2717 = \A[915]  & n2716 ;
  assign n2718 = ~n2714 & ~n2717 ;
  assign n2719 = n2713 & n2718 ;
  assign n2720 = ~n2713 & ~n2718 ;
  assign n2721 = ~\A[915]  & ~n2716 ;
  assign n2722 = ~n2717 & ~n2721 ;
  assign n2723 = ~\A[918]  & ~n2711 ;
  assign n2724 = ~n2712 & ~n2723 ;
  assign n2725 = n2722 & n2724 ;
  assign n2726 = ~n2720 & ~n2725 ;
  assign n2727 = ~n2719 & ~n2726 ;
  assign n2728 = ~n2722 & ~n2724 ;
  assign n2729 = ~n2725 & ~n2728 ;
  assign n2730 = ~n2696 & ~n2701 ;
  assign n2731 = ~n2702 & ~n2730 ;
  assign n2732 = n2729 & n2731 ;
  assign n2733 = n2703 & ~n2704 ;
  assign n2734 = n2732 & ~n2733 ;
  assign n2735 = ~n2719 & ~n2720 ;
  assign n2736 = n2725 & ~n2735 ;
  assign n2737 = ~n2725 & n2735 ;
  assign n2738 = ~n2736 & ~n2737 ;
  assign n2739 = n2734 & ~n2738 ;
  assign n2740 = ~n2734 & n2738 ;
  assign n2741 = ~n2703 & ~n2706 ;
  assign n2742 = n2704 & ~n2741 ;
  assign n2743 = ~n2704 & n2741 ;
  assign n2744 = ~n2742 & ~n2743 ;
  assign n2745 = ~n2740 & n2744 ;
  assign n2746 = ~n2739 & ~n2745 ;
  assign n2747 = n2727 & ~n2746 ;
  assign n2748 = ~n2727 & n2746 ;
  assign n2749 = ~n2747 & ~n2748 ;
  assign n2750 = n2708 & n2749 ;
  assign n2751 = ~n2708 & ~n2749 ;
  assign n2752 = ~n2750 & ~n2751 ;
  assign n2753 = ~n2689 & ~n2752 ;
  assign n2754 = n2689 & n2752 ;
  assign n2755 = ~n2729 & ~n2731 ;
  assign n2756 = ~n2732 & ~n2755 ;
  assign n2757 = ~n2666 & ~n2668 ;
  assign n2758 = ~n2669 & ~n2757 ;
  assign n2759 = n2756 & n2758 ;
  assign n2760 = ~n2739 & ~n2740 ;
  assign n2761 = n2744 & n2760 ;
  assign n2762 = ~n2744 & ~n2760 ;
  assign n2763 = ~n2761 & ~n2762 ;
  assign n2764 = n2759 & n2763 ;
  assign n2765 = ~n2759 & ~n2763 ;
  assign n2766 = ~n2676 & ~n2677 ;
  assign n2767 = n2681 & n2766 ;
  assign n2768 = ~n2681 & ~n2766 ;
  assign n2769 = ~n2767 & ~n2768 ;
  assign n2770 = ~n2765 & n2769 ;
  assign n2771 = ~n2764 & ~n2770 ;
  assign n2772 = ~n2754 & ~n2771 ;
  assign n2773 = ~n2753 & ~n2772 ;
  assign n2774 = ~n2708 & ~n2748 ;
  assign n2775 = ~n2747 & ~n2774 ;
  assign n2776 = ~n2773 & ~n2775 ;
  assign n2777 = n2773 & n2775 ;
  assign n2778 = ~n2776 & ~n2777 ;
  assign n2779 = ~n2645 & ~n2685 ;
  assign n2780 = ~n2684 & ~n2779 ;
  assign n2781 = n2778 & ~n2780 ;
  assign n2782 = ~n2778 & n2780 ;
  assign n2783 = ~n2781 & ~n2782 ;
  assign n2784 = ~n2626 & ~n2783 ;
  assign n2785 = n2626 & n2783 ;
  assign n2786 = ~n2753 & ~n2754 ;
  assign n2787 = ~n2771 & n2786 ;
  assign n2788 = n2771 & ~n2786 ;
  assign n2789 = ~n2787 & ~n2788 ;
  assign n2790 = ~n2594 & ~n2595 ;
  assign n2791 = ~n2612 & n2790 ;
  assign n2792 = n2612 & ~n2790 ;
  assign n2793 = ~n2791 & ~n2792 ;
  assign n2794 = ~n2789 & ~n2793 ;
  assign n2795 = n2789 & n2793 ;
  assign n2796 = ~n2597 & ~n2599 ;
  assign n2797 = ~n2600 & ~n2796 ;
  assign n2798 = ~n2756 & ~n2758 ;
  assign n2799 = ~n2759 & ~n2798 ;
  assign n2800 = n2797 & n2799 ;
  assign n2801 = ~n2605 & ~n2606 ;
  assign n2802 = ~n2610 & n2801 ;
  assign n2803 = n2610 & ~n2801 ;
  assign n2804 = ~n2802 & ~n2803 ;
  assign n2805 = n2800 & ~n2804 ;
  assign n2806 = ~n2800 & n2804 ;
  assign n2807 = ~n2764 & ~n2765 ;
  assign n2808 = ~n2769 & n2807 ;
  assign n2809 = n2769 & ~n2807 ;
  assign n2810 = ~n2808 & ~n2809 ;
  assign n2811 = ~n2806 & ~n2810 ;
  assign n2812 = ~n2805 & ~n2811 ;
  assign n2813 = ~n2795 & n2812 ;
  assign n2814 = ~n2794 & ~n2813 ;
  assign n2815 = ~n2785 & ~n2814 ;
  assign n2816 = ~n2784 & ~n2815 ;
  assign n2817 = n2622 & ~n2816 ;
  assign n2818 = ~n2622 & n2816 ;
  assign n2819 = ~n2817 & ~n2818 ;
  assign n2820 = ~n2777 & ~n2780 ;
  assign n2821 = ~n2776 & ~n2820 ;
  assign n2822 = n2819 & n2821 ;
  assign n2823 = ~n2819 & ~n2821 ;
  assign n2824 = ~n2822 & ~n2823 ;
  assign n2825 = ~n2467 & ~n2824 ;
  assign n2826 = n2467 & n2824 ;
  assign n2827 = ~n2784 & ~n2785 ;
  assign n2828 = ~n2814 & n2827 ;
  assign n2829 = n2814 & ~n2827 ;
  assign n2830 = ~n2828 & ~n2829 ;
  assign n2831 = ~n2427 & ~n2428 ;
  assign n2832 = ~n2457 & n2831 ;
  assign n2833 = n2457 & ~n2831 ;
  assign n2834 = ~n2832 & ~n2833 ;
  assign n2835 = ~n2830 & ~n2834 ;
  assign n2836 = n2830 & n2834 ;
  assign n2837 = ~n2437 & ~n2438 ;
  assign n2838 = ~n2455 & n2837 ;
  assign n2839 = n2455 & ~n2837 ;
  assign n2840 = ~n2838 & ~n2839 ;
  assign n2841 = ~n2794 & ~n2795 ;
  assign n2842 = ~n2812 & n2841 ;
  assign n2843 = n2812 & ~n2841 ;
  assign n2844 = ~n2842 & ~n2843 ;
  assign n2845 = ~n2840 & ~n2844 ;
  assign n2846 = n2840 & n2844 ;
  assign n2847 = ~n2797 & ~n2799 ;
  assign n2848 = ~n2800 & ~n2847 ;
  assign n2849 = ~n2440 & ~n2442 ;
  assign n2850 = ~n2443 & ~n2849 ;
  assign n2851 = n2848 & n2850 ;
  assign n2852 = ~n2805 & ~n2806 ;
  assign n2853 = ~n2810 & n2852 ;
  assign n2854 = n2810 & ~n2852 ;
  assign n2855 = ~n2853 & ~n2854 ;
  assign n2856 = n2851 & n2855 ;
  assign n2857 = ~n2851 & ~n2855 ;
  assign n2858 = ~n2448 & ~n2449 ;
  assign n2859 = ~n2453 & n2858 ;
  assign n2860 = n2453 & ~n2858 ;
  assign n2861 = ~n2859 & ~n2860 ;
  assign n2862 = ~n2857 & n2861 ;
  assign n2863 = ~n2856 & ~n2862 ;
  assign n2864 = ~n2846 & n2863 ;
  assign n2865 = ~n2845 & ~n2864 ;
  assign n2866 = ~n2836 & n2865 ;
  assign n2867 = ~n2835 & ~n2866 ;
  assign n2868 = ~n2826 & ~n2867 ;
  assign n2869 = ~n2825 & ~n2868 ;
  assign n2870 = ~n2818 & n2821 ;
  assign n2871 = ~n2817 & ~n2870 ;
  assign n2872 = n2869 & ~n2871 ;
  assign n2873 = ~n2869 & n2871 ;
  assign n2874 = ~n2461 & n2464 ;
  assign n2875 = ~n2460 & ~n2874 ;
  assign n2876 = ~n2873 & ~n2875 ;
  assign n2877 = ~n2872 & ~n2876 ;
  assign n2878 = ~n2110 & ~n2877 ;
  assign n2879 = ~n2049 & ~n2050 ;
  assign n2880 = n2103 & n2879 ;
  assign n2881 = ~n2103 & ~n2879 ;
  assign n2882 = ~n2880 & ~n2881 ;
  assign n2883 = ~n2872 & ~n2873 ;
  assign n2884 = n2875 & n2883 ;
  assign n2885 = ~n2875 & ~n2883 ;
  assign n2886 = ~n2884 & ~n2885 ;
  assign n2887 = ~n2882 & ~n2886 ;
  assign n2888 = n2882 & n2886 ;
  assign n2889 = ~n2825 & ~n2826 ;
  assign n2890 = ~n2867 & n2889 ;
  assign n2891 = n2867 & ~n2889 ;
  assign n2892 = ~n2890 & ~n2891 ;
  assign n2893 = ~n2059 & ~n2060 ;
  assign n2894 = ~n2101 & n2893 ;
  assign n2895 = n2101 & ~n2893 ;
  assign n2896 = ~n2894 & ~n2895 ;
  assign n2897 = ~n2892 & n2896 ;
  assign n2898 = n2892 & ~n2896 ;
  assign n2899 = ~n2069 & ~n2070 ;
  assign n2900 = ~n2099 & n2899 ;
  assign n2901 = n2099 & ~n2899 ;
  assign n2902 = ~n2900 & ~n2901 ;
  assign n2903 = ~n2835 & ~n2836 ;
  assign n2904 = n2865 & n2903 ;
  assign n2905 = ~n2865 & ~n2903 ;
  assign n2906 = ~n2904 & ~n2905 ;
  assign n2907 = n2902 & ~n2906 ;
  assign n2908 = ~n2902 & n2906 ;
  assign n2909 = ~n2845 & ~n2846 ;
  assign n2910 = ~n2863 & n2909 ;
  assign n2911 = n2863 & ~n2909 ;
  assign n2912 = ~n2910 & ~n2911 ;
  assign n2913 = ~n2079 & ~n2080 ;
  assign n2914 = ~n2097 & n2913 ;
  assign n2915 = n2097 & ~n2913 ;
  assign n2916 = ~n2914 & ~n2915 ;
  assign n2917 = ~n2912 & ~n2916 ;
  assign n2918 = n2912 & n2916 ;
  assign n2919 = ~n2848 & ~n2850 ;
  assign n2920 = ~n2851 & ~n2919 ;
  assign n2921 = ~n2082 & ~n2084 ;
  assign n2922 = ~n2085 & ~n2921 ;
  assign n2923 = n2920 & n2922 ;
  assign n2924 = ~n2090 & ~n2091 ;
  assign n2925 = ~n2095 & n2924 ;
  assign n2926 = n2095 & ~n2924 ;
  assign n2927 = ~n2925 & ~n2926 ;
  assign n2928 = n2923 & ~n2927 ;
  assign n2929 = ~n2923 & n2927 ;
  assign n2930 = ~n2856 & ~n2857 ;
  assign n2931 = ~n2861 & n2930 ;
  assign n2932 = n2861 & ~n2930 ;
  assign n2933 = ~n2931 & ~n2932 ;
  assign n2934 = ~n2929 & ~n2933 ;
  assign n2935 = ~n2928 & ~n2934 ;
  assign n2936 = ~n2918 & n2935 ;
  assign n2937 = ~n2917 & ~n2936 ;
  assign n2938 = ~n2908 & ~n2937 ;
  assign n2939 = ~n2907 & ~n2938 ;
  assign n2940 = ~n2898 & ~n2939 ;
  assign n2941 = ~n2897 & ~n2940 ;
  assign n2942 = ~n2888 & ~n2941 ;
  assign n2943 = ~n2887 & ~n2942 ;
  assign n2944 = ~n2878 & n2943 ;
  assign n2945 = n2108 & n2944 ;
  assign n2946 = \A[403]  & \A[404]  ;
  assign n2947 = ~\A[403]  & ~\A[404]  ;
  assign n2948 = ~n2946 & ~n2947 ;
  assign n2949 = \A[405]  & n2948 ;
  assign n2950 = ~n2946 & ~n2949 ;
  assign n2951 = \A[406]  & \A[407]  ;
  assign n2952 = ~\A[405]  & ~n2948 ;
  assign n2953 = ~n2949 & ~n2952 ;
  assign n2954 = ~\A[406]  & ~\A[407]  ;
  assign n2955 = ~n2951 & ~n2954 ;
  assign n2956 = \A[408]  & n2955 ;
  assign n2957 = ~\A[408]  & ~n2955 ;
  assign n2958 = ~n2956 & ~n2957 ;
  assign n2959 = n2953 & n2958 ;
  assign n2960 = n2951 & n2959 ;
  assign n2961 = ~n2951 & ~n2956 ;
  assign n2962 = ~n2959 & n2961 ;
  assign n2963 = ~n2960 & ~n2962 ;
  assign n2964 = n2950 & ~n2963 ;
  assign n2965 = ~n2950 & n2963 ;
  assign n2966 = ~n2964 & ~n2965 ;
  assign n2967 = \A[409]  & \A[410]  ;
  assign n2968 = ~\A[409]  & ~\A[410]  ;
  assign n2969 = ~n2967 & ~n2968 ;
  assign n2970 = \A[411]  & n2969 ;
  assign n2971 = ~\A[411]  & ~n2969 ;
  assign n2972 = ~n2970 & ~n2971 ;
  assign n2973 = \A[412]  & \A[413]  ;
  assign n2974 = ~\A[412]  & ~\A[413]  ;
  assign n2975 = ~n2973 & ~n2974 ;
  assign n2976 = \A[414]  & n2975 ;
  assign n2977 = ~\A[414]  & ~n2975 ;
  assign n2978 = ~n2976 & ~n2977 ;
  assign n2979 = n2972 & n2978 ;
  assign n2980 = ~n2973 & ~n2976 ;
  assign n2981 = ~n2967 & ~n2970 ;
  assign n2982 = ~n2980 & ~n2981 ;
  assign n2983 = n2980 & n2981 ;
  assign n2984 = ~n2982 & ~n2983 ;
  assign n2991 = n2979 & ~n2984 ;
  assign n2985 = ~n2979 & n2984 ;
  assign n2986 = ~n2953 & ~n2958 ;
  assign n2987 = ~n2959 & ~n2986 ;
  assign n2988 = ~n2972 & ~n2978 ;
  assign n2989 = ~n2979 & ~n2988 ;
  assign n2990 = n2987 & n2989 ;
  assign n2992 = ~n2985 & ~n2990 ;
  assign n2993 = ~n2991 & n2992 ;
  assign n2994 = n2966 & ~n2993 ;
  assign n2995 = n2984 & n2990 ;
  assign n2996 = ~n2950 & n2960 ;
  assign n2997 = n2995 & ~n2996 ;
  assign n2998 = ~n2994 & ~n2997 ;
  assign n2999 = ~n2973 & n2981 ;
  assign n3000 = n2979 & ~n2999 ;
  assign n3001 = ~n2982 & ~n3000 ;
  assign n3002 = ~n2998 & ~n3001 ;
  assign n3003 = ~n2950 & ~n2962 ;
  assign n3004 = ~n2960 & ~n3003 ;
  assign n3005 = n2998 & n3001 ;
  assign n3006 = ~n3004 & ~n3005 ;
  assign n3007 = ~n3002 & ~n3006 ;
  assign n3008 = \A[397]  & \A[398]  ;
  assign n3009 = ~\A[397]  & ~\A[398]  ;
  assign n3010 = ~n3008 & ~n3009 ;
  assign n3011 = \A[399]  & n3010 ;
  assign n3012 = ~\A[399]  & ~n3010 ;
  assign n3013 = ~n3011 & ~n3012 ;
  assign n3014 = \A[400]  & \A[401]  ;
  assign n3015 = ~\A[400]  & ~\A[401]  ;
  assign n3016 = ~n3014 & ~n3015 ;
  assign n3017 = \A[402]  & n3016 ;
  assign n3018 = ~\A[402]  & ~n3016 ;
  assign n3019 = ~n3017 & ~n3018 ;
  assign n3020 = n3013 & n3019 ;
  assign n3021 = ~n3013 & ~n3019 ;
  assign n3022 = ~n3020 & ~n3021 ;
  assign n3023 = \A[391]  & \A[392]  ;
  assign n3024 = ~\A[391]  & ~\A[392]  ;
  assign n3025 = ~n3023 & ~n3024 ;
  assign n3026 = \A[393]  & n3025 ;
  assign n3027 = ~\A[393]  & ~n3025 ;
  assign n3028 = ~n3026 & ~n3027 ;
  assign n3029 = \A[394]  & \A[395]  ;
  assign n3030 = ~\A[394]  & ~\A[395]  ;
  assign n3031 = ~n3029 & ~n3030 ;
  assign n3032 = \A[396]  & n3031 ;
  assign n3033 = ~\A[396]  & ~n3031 ;
  assign n3034 = ~n3032 & ~n3033 ;
  assign n3035 = n3028 & n3034 ;
  assign n3036 = ~n3028 & ~n3034 ;
  assign n3037 = ~n3035 & ~n3036 ;
  assign n3038 = n3022 & n3037 ;
  assign n3039 = ~n3008 & ~n3011 ;
  assign n3040 = ~n3014 & ~n3017 ;
  assign n3041 = ~n3020 & n3040 ;
  assign n3042 = n3014 & n3020 ;
  assign n3043 = ~n3041 & ~n3042 ;
  assign n3044 = n3039 & ~n3043 ;
  assign n3045 = ~n3039 & n3043 ;
  assign n3046 = ~n3044 & ~n3045 ;
  assign n3047 = ~n3038 & ~n3046 ;
  assign n3048 = ~n3023 & ~n3026 ;
  assign n3049 = n3029 & n3035 ;
  assign n3050 = ~n3029 & ~n3032 ;
  assign n3051 = ~n3035 & n3050 ;
  assign n3052 = ~n3049 & ~n3051 ;
  assign n3053 = n3048 & ~n3052 ;
  assign n3054 = ~n3048 & n3052 ;
  assign n3055 = ~n3053 & ~n3054 ;
  assign n3056 = ~n3047 & n3055 ;
  assign n3057 = n3038 & n3046 ;
  assign n3058 = ~n3039 & ~n3040 ;
  assign n3059 = ~n3048 & n3049 ;
  assign n3060 = ~n3058 & ~n3059 ;
  assign n3061 = n3057 & n3060 ;
  assign n3062 = ~n3056 & ~n3061 ;
  assign n3063 = ~n3039 & ~n3041 ;
  assign n3064 = ~n3042 & ~n3063 ;
  assign n3065 = ~n3062 & ~n3064 ;
  assign n3066 = ~n3048 & ~n3051 ;
  assign n3067 = ~n3049 & ~n3066 ;
  assign n3068 = n3062 & n3064 ;
  assign n3069 = ~n3067 & ~n3068 ;
  assign n3070 = ~n3065 & ~n3069 ;
  assign n3071 = ~n3007 & ~n3070 ;
  assign n3072 = n3007 & n3070 ;
  assign n3073 = ~n3065 & ~n3068 ;
  assign n3074 = n3067 & ~n3073 ;
  assign n3075 = ~n3067 & n3073 ;
  assign n3076 = ~n3074 & ~n3075 ;
  assign n3077 = ~n3002 & ~n3005 ;
  assign n3078 = n3004 & ~n3077 ;
  assign n3079 = ~n3004 & n3077 ;
  assign n3080 = ~n3078 & ~n3079 ;
  assign n3081 = ~n3076 & ~n3080 ;
  assign n3082 = ~n2987 & ~n2989 ;
  assign n3083 = ~n2990 & ~n3082 ;
  assign n3084 = ~n3022 & ~n3037 ;
  assign n3085 = ~n3038 & ~n3084 ;
  assign n3086 = n3083 & n3085 ;
  assign n3087 = n2994 & ~n2997 ;
  assign n3088 = ~n2993 & ~n2995 ;
  assign n3089 = ~n2966 & ~n3088 ;
  assign n3090 = ~n3087 & ~n3089 ;
  assign n3091 = ~n3086 & ~n3090 ;
  assign n3092 = n3056 & ~n3061 ;
  assign n3093 = ~n3047 & ~n3057 ;
  assign n3094 = ~n3055 & ~n3093 ;
  assign n3095 = ~n3092 & ~n3094 ;
  assign n3096 = n3086 & n3090 ;
  assign n3097 = ~n3095 & ~n3096 ;
  assign n3098 = ~n3091 & ~n3097 ;
  assign n3099 = n3076 & n3080 ;
  assign n3100 = ~n3098 & ~n3099 ;
  assign n3101 = ~n3081 & ~n3100 ;
  assign n3102 = ~n3072 & n3101 ;
  assign n3103 = ~n3071 & ~n3102 ;
  assign n3104 = \A[385]  & \A[386]  ;
  assign n3105 = ~\A[385]  & ~\A[386]  ;
  assign n3106 = ~n3104 & ~n3105 ;
  assign n3107 = \A[387]  & n3106 ;
  assign n3108 = ~\A[387]  & ~n3106 ;
  assign n3109 = ~n3107 & ~n3108 ;
  assign n3110 = \A[388]  & \A[389]  ;
  assign n3111 = ~\A[388]  & ~\A[389]  ;
  assign n3112 = ~n3110 & ~n3111 ;
  assign n3113 = \A[390]  & n3112 ;
  assign n3114 = ~\A[390]  & ~n3112 ;
  assign n3115 = ~n3113 & ~n3114 ;
  assign n3116 = n3109 & n3115 ;
  assign n3117 = ~n3109 & ~n3115 ;
  assign n3118 = ~n3116 & ~n3117 ;
  assign n3119 = \A[379]  & \A[380]  ;
  assign n3120 = ~\A[379]  & ~\A[380]  ;
  assign n3121 = ~n3119 & ~n3120 ;
  assign n3122 = \A[381]  & n3121 ;
  assign n3123 = ~\A[381]  & ~n3121 ;
  assign n3124 = ~n3122 & ~n3123 ;
  assign n3125 = \A[382]  & \A[383]  ;
  assign n3126 = ~\A[382]  & ~\A[383]  ;
  assign n3127 = ~n3125 & ~n3126 ;
  assign n3128 = \A[384]  & n3127 ;
  assign n3129 = ~\A[384]  & ~n3127 ;
  assign n3130 = ~n3128 & ~n3129 ;
  assign n3131 = n3124 & n3130 ;
  assign n3132 = ~n3124 & ~n3130 ;
  assign n3133 = ~n3131 & ~n3132 ;
  assign n3134 = n3118 & n3133 ;
  assign n3135 = ~n3110 & ~n3113 ;
  assign n3136 = ~n3104 & ~n3107 ;
  assign n3137 = ~n3135 & ~n3136 ;
  assign n3138 = n3135 & n3136 ;
  assign n3139 = ~n3137 & ~n3138 ;
  assign n3140 = n3134 & n3139 ;
  assign n3141 = ~n3119 & ~n3122 ;
  assign n3142 = ~n3125 & ~n3128 ;
  assign n3143 = ~n3131 & n3142 ;
  assign n3144 = n3125 & n3131 ;
  assign n3145 = ~n3143 & ~n3144 ;
  assign n3146 = n3141 & ~n3145 ;
  assign n3147 = ~n3141 & n3145 ;
  assign n3148 = ~n3146 & ~n3147 ;
  assign n3149 = ~n3140 & ~n3148 ;
  assign n3151 = n3116 & ~n3139 ;
  assign n3150 = ~n3116 & n3139 ;
  assign n3152 = ~n3134 & ~n3150 ;
  assign n3153 = ~n3151 & n3152 ;
  assign n3154 = ~n3149 & ~n3153 ;
  assign n3155 = ~n3116 & ~n3137 ;
  assign n3156 = ~n3138 & ~n3155 ;
  assign n3157 = ~n3154 & ~n3156 ;
  assign n3158 = n3154 & n3156 ;
  assign n3159 = ~n3141 & ~n3143 ;
  assign n3160 = ~n3144 & ~n3159 ;
  assign n3161 = ~n3158 & n3160 ;
  assign n3162 = ~n3157 & ~n3161 ;
  assign n3163 = ~n3157 & ~n3158 ;
  assign n3164 = ~n3160 & n3163 ;
  assign n3165 = n3160 & ~n3163 ;
  assign n3166 = ~n3164 & ~n3165 ;
  assign n3167 = \A[370]  & \A[371]  ;
  assign n3168 = \A[367]  & \A[368]  ;
  assign n3169 = ~\A[367]  & ~\A[368]  ;
  assign n3170 = ~n3168 & ~n3169 ;
  assign n3171 = \A[369]  & n3170 ;
  assign n3172 = ~\A[369]  & ~n3170 ;
  assign n3173 = ~n3171 & ~n3172 ;
  assign n3174 = ~\A[370]  & ~\A[371]  ;
  assign n3175 = ~n3167 & ~n3174 ;
  assign n3176 = \A[372]  & n3175 ;
  assign n3177 = ~\A[372]  & ~n3175 ;
  assign n3178 = ~n3176 & ~n3177 ;
  assign n3179 = n3173 & n3178 ;
  assign n3180 = n3167 & n3179 ;
  assign n3181 = ~n3168 & ~n3171 ;
  assign n3182 = ~n3167 & ~n3176 ;
  assign n3183 = ~n3179 & n3182 ;
  assign n3184 = ~n3181 & ~n3183 ;
  assign n3185 = ~n3180 & ~n3184 ;
  assign n3186 = \A[373]  & \A[374]  ;
  assign n3187 = ~\A[373]  & ~\A[374]  ;
  assign n3188 = ~n3186 & ~n3187 ;
  assign n3189 = \A[375]  & n3188 ;
  assign n3190 = ~\A[375]  & ~n3188 ;
  assign n3191 = ~n3189 & ~n3190 ;
  assign n3192 = \A[376]  & \A[377]  ;
  assign n3193 = ~\A[376]  & ~\A[377]  ;
  assign n3194 = ~n3192 & ~n3193 ;
  assign n3195 = \A[378]  & n3194 ;
  assign n3196 = ~\A[378]  & ~n3194 ;
  assign n3197 = ~n3195 & ~n3196 ;
  assign n3198 = n3191 & n3197 ;
  assign n3199 = ~n3191 & ~n3197 ;
  assign n3200 = ~n3198 & ~n3199 ;
  assign n3201 = ~n3173 & ~n3178 ;
  assign n3202 = ~n3179 & ~n3201 ;
  assign n3203 = n3200 & n3202 ;
  assign n3204 = ~n3192 & ~n3195 ;
  assign n3205 = ~n3186 & ~n3189 ;
  assign n3206 = ~n3204 & ~n3205 ;
  assign n3207 = n3204 & n3205 ;
  assign n3208 = ~n3206 & ~n3207 ;
  assign n3209 = n3203 & n3208 ;
  assign n3210 = ~n3180 & ~n3183 ;
  assign n3211 = n3181 & ~n3210 ;
  assign n3212 = ~n3181 & n3210 ;
  assign n3213 = ~n3211 & ~n3212 ;
  assign n3214 = ~n3209 & ~n3213 ;
  assign n3216 = n3198 & ~n3208 ;
  assign n3215 = ~n3198 & n3208 ;
  assign n3217 = ~n3203 & ~n3215 ;
  assign n3218 = ~n3216 & n3217 ;
  assign n3219 = ~n3214 & ~n3218 ;
  assign n3220 = ~n3198 & ~n3206 ;
  assign n3221 = ~n3207 & ~n3220 ;
  assign n3222 = n3219 & n3221 ;
  assign n3223 = ~n3219 & ~n3221 ;
  assign n3224 = ~n3222 & ~n3223 ;
  assign n3225 = n3185 & ~n3224 ;
  assign n3226 = ~n3185 & n3224 ;
  assign n3227 = ~n3225 & ~n3226 ;
  assign n3228 = n3166 & n3227 ;
  assign n3229 = ~n3166 & ~n3227 ;
  assign n3230 = ~n3118 & ~n3133 ;
  assign n3231 = ~n3134 & ~n3230 ;
  assign n3232 = ~n3200 & ~n3202 ;
  assign n3233 = ~n3203 & ~n3232 ;
  assign n3234 = n3231 & n3233 ;
  assign n3235 = ~n3140 & ~n3153 ;
  assign n3236 = ~n3148 & n3235 ;
  assign n3237 = n3148 & ~n3235 ;
  assign n3238 = ~n3236 & ~n3237 ;
  assign n3239 = n3234 & ~n3238 ;
  assign n3240 = ~n3234 & n3238 ;
  assign n3241 = ~n3209 & ~n3218 ;
  assign n3242 = ~n3213 & n3241 ;
  assign n3243 = n3213 & ~n3241 ;
  assign n3244 = ~n3242 & ~n3243 ;
  assign n3245 = ~n3240 & ~n3244 ;
  assign n3246 = ~n3239 & ~n3245 ;
  assign n3247 = ~n3229 & ~n3246 ;
  assign n3248 = ~n3228 & ~n3247 ;
  assign n3249 = n3162 & ~n3248 ;
  assign n3250 = ~n3162 & n3248 ;
  assign n3251 = n3185 & ~n3222 ;
  assign n3252 = ~n3223 & ~n3251 ;
  assign n3253 = ~n3250 & n3252 ;
  assign n3254 = ~n3249 & ~n3253 ;
  assign n3255 = ~n3103 & ~n3254 ;
  assign n3256 = n3103 & n3254 ;
  assign n3257 = ~n3071 & ~n3072 ;
  assign n3258 = n3101 & ~n3257 ;
  assign n3259 = ~n3101 & n3257 ;
  assign n3260 = ~n3258 & ~n3259 ;
  assign n3261 = ~n3249 & ~n3250 ;
  assign n3262 = n3252 & n3261 ;
  assign n3263 = ~n3252 & ~n3261 ;
  assign n3264 = ~n3262 & ~n3263 ;
  assign n3265 = ~n3260 & n3264 ;
  assign n3266 = n3260 & ~n3264 ;
  assign n3267 = ~n3081 & ~n3099 ;
  assign n3268 = n3098 & n3267 ;
  assign n3269 = ~n3098 & ~n3267 ;
  assign n3270 = ~n3268 & ~n3269 ;
  assign n3271 = ~n3228 & ~n3229 ;
  assign n3272 = ~n3246 & n3271 ;
  assign n3273 = n3246 & ~n3271 ;
  assign n3274 = ~n3272 & ~n3273 ;
  assign n3275 = n3270 & n3274 ;
  assign n3276 = ~n3270 & ~n3274 ;
  assign n3277 = ~n3083 & ~n3085 ;
  assign n3278 = ~n3086 & ~n3277 ;
  assign n3279 = ~n3231 & ~n3233 ;
  assign n3280 = ~n3234 & ~n3279 ;
  assign n3281 = n3278 & n3280 ;
  assign n3282 = ~n3091 & ~n3096 ;
  assign n3283 = n3095 & ~n3282 ;
  assign n3284 = ~n3095 & n3282 ;
  assign n3285 = ~n3283 & ~n3284 ;
  assign n3286 = n3281 & ~n3285 ;
  assign n3287 = ~n3281 & n3285 ;
  assign n3288 = ~n3239 & ~n3240 ;
  assign n3289 = ~n3244 & n3288 ;
  assign n3290 = n3244 & ~n3288 ;
  assign n3291 = ~n3289 & ~n3290 ;
  assign n3292 = ~n3287 & n3291 ;
  assign n3293 = ~n3286 & ~n3292 ;
  assign n3294 = ~n3276 & ~n3293 ;
  assign n3295 = ~n3275 & ~n3294 ;
  assign n3296 = ~n3266 & ~n3295 ;
  assign n3297 = ~n3265 & ~n3296 ;
  assign n3298 = ~n3256 & ~n3297 ;
  assign n3299 = ~n3255 & ~n3298 ;
  assign n3300 = \A[445]  & \A[446]  ;
  assign n3301 = ~\A[445]  & ~\A[446]  ;
  assign n3302 = ~n3300 & ~n3301 ;
  assign n3303 = \A[447]  & n3302 ;
  assign n3304 = ~\A[447]  & ~n3302 ;
  assign n3305 = ~n3303 & ~n3304 ;
  assign n3306 = \A[448]  & \A[449]  ;
  assign n3307 = ~\A[448]  & ~\A[449]  ;
  assign n3308 = ~n3306 & ~n3307 ;
  assign n3309 = \A[450]  & n3308 ;
  assign n3310 = ~\A[450]  & ~n3308 ;
  assign n3311 = ~n3309 & ~n3310 ;
  assign n3312 = n3305 & n3311 ;
  assign n3313 = ~n3305 & ~n3311 ;
  assign n3314 = ~n3312 & ~n3313 ;
  assign n3315 = \A[439]  & \A[440]  ;
  assign n3316 = ~\A[439]  & ~\A[440]  ;
  assign n3317 = ~n3315 & ~n3316 ;
  assign n3318 = \A[441]  & n3317 ;
  assign n3319 = ~\A[441]  & ~n3317 ;
  assign n3320 = ~n3318 & ~n3319 ;
  assign n3321 = \A[442]  & \A[443]  ;
  assign n3322 = ~\A[442]  & ~\A[443]  ;
  assign n3323 = ~n3321 & ~n3322 ;
  assign n3324 = \A[444]  & n3323 ;
  assign n3325 = ~\A[444]  & ~n3323 ;
  assign n3326 = ~n3324 & ~n3325 ;
  assign n3327 = n3320 & n3326 ;
  assign n3328 = ~n3320 & ~n3326 ;
  assign n3329 = ~n3327 & ~n3328 ;
  assign n3330 = n3314 & n3329 ;
  assign n3331 = ~n3300 & ~n3303 ;
  assign n3332 = ~n3306 & ~n3309 ;
  assign n3333 = ~n3312 & n3332 ;
  assign n3334 = n3306 & n3312 ;
  assign n3335 = ~n3333 & ~n3334 ;
  assign n3336 = n3331 & ~n3335 ;
  assign n3337 = ~n3331 & n3335 ;
  assign n3338 = ~n3336 & ~n3337 ;
  assign n3339 = ~n3330 & ~n3338 ;
  assign n3340 = ~n3315 & ~n3318 ;
  assign n3341 = n3321 & n3327 ;
  assign n3342 = ~n3321 & ~n3324 ;
  assign n3343 = ~n3327 & n3342 ;
  assign n3344 = ~n3341 & ~n3343 ;
  assign n3345 = n3340 & ~n3344 ;
  assign n3346 = ~n3340 & n3344 ;
  assign n3347 = ~n3345 & ~n3346 ;
  assign n3348 = ~n3339 & n3347 ;
  assign n3349 = n3330 & n3338 ;
  assign n3350 = ~n3331 & ~n3332 ;
  assign n3351 = ~n3340 & n3341 ;
  assign n3352 = ~n3350 & ~n3351 ;
  assign n3353 = n3349 & n3352 ;
  assign n3354 = ~n3348 & ~n3353 ;
  assign n3355 = ~n3331 & ~n3333 ;
  assign n3356 = ~n3334 & ~n3355 ;
  assign n3357 = ~n3354 & ~n3356 ;
  assign n3358 = ~n3340 & ~n3343 ;
  assign n3359 = ~n3341 & ~n3358 ;
  assign n3360 = n3354 & n3356 ;
  assign n3361 = ~n3359 & ~n3360 ;
  assign n3362 = ~n3357 & ~n3361 ;
  assign n3363 = \A[451]  & \A[452]  ;
  assign n3364 = ~\A[451]  & ~\A[452]  ;
  assign n3365 = ~n3363 & ~n3364 ;
  assign n3366 = \A[453]  & n3365 ;
  assign n3367 = ~\A[453]  & ~n3365 ;
  assign n3368 = ~n3366 & ~n3367 ;
  assign n3369 = \A[454]  & \A[455]  ;
  assign n3370 = ~\A[454]  & ~\A[455]  ;
  assign n3371 = ~n3369 & ~n3370 ;
  assign n3372 = \A[456]  & n3371 ;
  assign n3373 = ~\A[456]  & ~n3371 ;
  assign n3374 = ~n3372 & ~n3373 ;
  assign n3375 = n3368 & n3374 ;
  assign n3376 = ~n3369 & ~n3372 ;
  assign n3377 = ~n3363 & ~n3366 ;
  assign n3378 = n3376 & n3377 ;
  assign n3379 = ~n3376 & ~n3377 ;
  assign n3380 = ~n3378 & ~n3379 ;
  assign n3381 = n3375 & ~n3380 ;
  assign n3382 = ~n3375 & n3380 ;
  assign n3383 = ~n3381 & ~n3382 ;
  assign n3384 = \A[457]  & \A[458]  ;
  assign n3385 = ~\A[457]  & ~\A[458]  ;
  assign n3386 = ~n3384 & ~n3385 ;
  assign n3387 = \A[459]  & n3386 ;
  assign n3388 = ~\A[459]  & ~n3386 ;
  assign n3389 = ~n3387 & ~n3388 ;
  assign n3390 = \A[460]  & \A[461]  ;
  assign n3391 = ~\A[460]  & ~\A[461]  ;
  assign n3392 = ~n3390 & ~n3391 ;
  assign n3393 = \A[462]  & n3392 ;
  assign n3394 = ~\A[462]  & ~n3392 ;
  assign n3395 = ~n3393 & ~n3394 ;
  assign n3396 = n3389 & n3395 ;
  assign n3397 = ~n3390 & ~n3393 ;
  assign n3398 = ~n3384 & ~n3387 ;
  assign n3399 = ~n3397 & ~n3398 ;
  assign n3400 = n3397 & n3398 ;
  assign n3401 = ~n3399 & ~n3400 ;
  assign n3408 = n3396 & ~n3401 ;
  assign n3402 = ~n3396 & n3401 ;
  assign n3403 = ~n3389 & ~n3395 ;
  assign n3404 = ~n3396 & ~n3403 ;
  assign n3405 = ~n3368 & ~n3374 ;
  assign n3406 = ~n3375 & ~n3405 ;
  assign n3407 = n3404 & n3406 ;
  assign n3409 = ~n3402 & ~n3407 ;
  assign n3410 = ~n3408 & n3409 ;
  assign n3411 = ~n3383 & ~n3410 ;
  assign n3412 = n3375 & n3379 ;
  assign n3413 = n3401 & n3407 ;
  assign n3414 = ~n3412 & n3413 ;
  assign n3415 = ~n3411 & ~n3414 ;
  assign n3416 = ~n3390 & n3398 ;
  assign n3417 = n3396 & ~n3416 ;
  assign n3418 = ~n3399 & ~n3417 ;
  assign n3419 = n3415 & n3418 ;
  assign n3420 = ~n3415 & ~n3418 ;
  assign n3421 = ~n3375 & ~n3379 ;
  assign n3422 = ~n3378 & ~n3421 ;
  assign n3423 = ~n3420 & ~n3422 ;
  assign n3424 = ~n3419 & ~n3423 ;
  assign n3425 = ~n3362 & n3424 ;
  assign n3426 = n3362 & ~n3424 ;
  assign n3427 = ~n3357 & ~n3360 ;
  assign n3428 = n3359 & ~n3427 ;
  assign n3429 = ~n3359 & n3427 ;
  assign n3430 = ~n3428 & ~n3429 ;
  assign n3431 = ~n3419 & ~n3420 ;
  assign n3432 = ~n3422 & n3431 ;
  assign n3433 = n3422 & ~n3431 ;
  assign n3434 = ~n3432 & ~n3433 ;
  assign n3435 = n3430 & ~n3434 ;
  assign n3436 = ~n3430 & n3434 ;
  assign n3437 = ~n3404 & ~n3406 ;
  assign n3438 = ~n3407 & ~n3437 ;
  assign n3439 = ~n3314 & ~n3329 ;
  assign n3440 = ~n3330 & ~n3439 ;
  assign n3441 = n3438 & n3440 ;
  assign n3442 = n3411 & ~n3414 ;
  assign n3443 = ~n3410 & ~n3413 ;
  assign n3444 = n3383 & ~n3443 ;
  assign n3445 = ~n3442 & ~n3444 ;
  assign n3446 = ~n3441 & ~n3445 ;
  assign n3447 = n3348 & ~n3353 ;
  assign n3448 = ~n3339 & ~n3349 ;
  assign n3449 = ~n3347 & ~n3448 ;
  assign n3450 = ~n3447 & ~n3449 ;
  assign n3451 = n3441 & n3445 ;
  assign n3452 = ~n3450 & ~n3451 ;
  assign n3453 = ~n3446 & ~n3452 ;
  assign n3454 = ~n3436 & n3453 ;
  assign n3455 = ~n3435 & ~n3454 ;
  assign n3456 = ~n3426 & ~n3455 ;
  assign n3457 = ~n3425 & ~n3456 ;
  assign n3458 = \A[427]  & \A[428]  ;
  assign n3459 = ~\A[427]  & ~\A[428]  ;
  assign n3460 = ~n3458 & ~n3459 ;
  assign n3461 = \A[429]  & n3460 ;
  assign n3462 = ~n3458 & ~n3461 ;
  assign n3463 = \A[430]  & \A[431]  ;
  assign n3464 = ~\A[429]  & ~n3460 ;
  assign n3465 = ~n3461 & ~n3464 ;
  assign n3466 = ~\A[430]  & ~\A[431]  ;
  assign n3467 = ~n3463 & ~n3466 ;
  assign n3468 = \A[432]  & n3467 ;
  assign n3469 = ~\A[432]  & ~n3467 ;
  assign n3470 = ~n3468 & ~n3469 ;
  assign n3471 = n3465 & n3470 ;
  assign n3472 = n3463 & n3471 ;
  assign n3473 = ~n3463 & ~n3468 ;
  assign n3474 = ~n3471 & n3473 ;
  assign n3475 = ~n3472 & ~n3474 ;
  assign n3476 = n3462 & ~n3475 ;
  assign n3477 = ~n3462 & n3475 ;
  assign n3478 = ~n3476 & ~n3477 ;
  assign n3479 = \A[433]  & \A[434]  ;
  assign n3480 = ~\A[433]  & ~\A[434]  ;
  assign n3481 = ~n3479 & ~n3480 ;
  assign n3482 = \A[435]  & n3481 ;
  assign n3483 = ~\A[435]  & ~n3481 ;
  assign n3484 = ~n3482 & ~n3483 ;
  assign n3485 = \A[436]  & \A[437]  ;
  assign n3486 = ~\A[436]  & ~\A[437]  ;
  assign n3487 = ~n3485 & ~n3486 ;
  assign n3488 = \A[438]  & n3487 ;
  assign n3489 = ~\A[438]  & ~n3487 ;
  assign n3490 = ~n3488 & ~n3489 ;
  assign n3491 = n3484 & n3490 ;
  assign n3492 = ~n3485 & ~n3488 ;
  assign n3493 = ~n3479 & ~n3482 ;
  assign n3494 = ~n3492 & ~n3493 ;
  assign n3495 = n3492 & n3493 ;
  assign n3496 = ~n3494 & ~n3495 ;
  assign n3503 = n3491 & ~n3496 ;
  assign n3497 = ~n3491 & n3496 ;
  assign n3498 = ~n3465 & ~n3470 ;
  assign n3499 = ~n3471 & ~n3498 ;
  assign n3500 = ~n3484 & ~n3490 ;
  assign n3501 = ~n3491 & ~n3500 ;
  assign n3502 = n3499 & n3501 ;
  assign n3504 = ~n3497 & ~n3502 ;
  assign n3505 = ~n3503 & n3504 ;
  assign n3506 = n3478 & ~n3505 ;
  assign n3507 = n3496 & n3502 ;
  assign n3508 = ~n3462 & n3472 ;
  assign n3509 = n3507 & ~n3508 ;
  assign n3510 = ~n3506 & ~n3509 ;
  assign n3511 = ~n3485 & n3493 ;
  assign n3512 = n3491 & ~n3511 ;
  assign n3513 = ~n3494 & ~n3512 ;
  assign n3514 = ~n3510 & ~n3513 ;
  assign n3515 = ~n3462 & ~n3474 ;
  assign n3516 = ~n3472 & ~n3515 ;
  assign n3517 = n3510 & n3513 ;
  assign n3518 = ~n3516 & ~n3517 ;
  assign n3519 = ~n3514 & ~n3518 ;
  assign n3520 = \A[421]  & \A[422]  ;
  assign n3521 = ~\A[421]  & ~\A[422]  ;
  assign n3522 = ~n3520 & ~n3521 ;
  assign n3523 = \A[423]  & n3522 ;
  assign n3524 = ~\A[423]  & ~n3522 ;
  assign n3525 = ~n3523 & ~n3524 ;
  assign n3526 = \A[424]  & \A[425]  ;
  assign n3527 = ~\A[424]  & ~\A[425]  ;
  assign n3528 = ~n3526 & ~n3527 ;
  assign n3529 = \A[426]  & n3528 ;
  assign n3530 = ~\A[426]  & ~n3528 ;
  assign n3531 = ~n3529 & ~n3530 ;
  assign n3532 = n3525 & n3531 ;
  assign n3533 = ~n3525 & ~n3531 ;
  assign n3534 = ~n3532 & ~n3533 ;
  assign n3535 = \A[415]  & \A[416]  ;
  assign n3536 = ~\A[415]  & ~\A[416]  ;
  assign n3537 = ~n3535 & ~n3536 ;
  assign n3538 = \A[417]  & n3537 ;
  assign n3539 = ~\A[417]  & ~n3537 ;
  assign n3540 = ~n3538 & ~n3539 ;
  assign n3541 = \A[418]  & \A[419]  ;
  assign n3542 = ~\A[418]  & ~\A[419]  ;
  assign n3543 = ~n3541 & ~n3542 ;
  assign n3544 = \A[420]  & n3543 ;
  assign n3545 = ~\A[420]  & ~n3543 ;
  assign n3546 = ~n3544 & ~n3545 ;
  assign n3547 = n3540 & n3546 ;
  assign n3548 = ~n3540 & ~n3546 ;
  assign n3549 = ~n3547 & ~n3548 ;
  assign n3550 = n3534 & n3549 ;
  assign n3551 = ~n3526 & ~n3529 ;
  assign n3552 = ~n3520 & ~n3523 ;
  assign n3553 = ~n3551 & ~n3552 ;
  assign n3554 = n3551 & n3552 ;
  assign n3555 = ~n3553 & ~n3554 ;
  assign n3556 = n3550 & n3555 ;
  assign n3557 = ~n3541 & ~n3544 ;
  assign n3558 = ~n3535 & ~n3538 ;
  assign n3559 = n3557 & n3558 ;
  assign n3560 = ~n3557 & ~n3558 ;
  assign n3561 = ~n3559 & ~n3560 ;
  assign n3562 = n3547 & ~n3561 ;
  assign n3563 = ~n3547 & n3561 ;
  assign n3564 = ~n3562 & ~n3563 ;
  assign n3565 = ~n3556 & n3564 ;
  assign n3567 = n3532 & ~n3555 ;
  assign n3566 = ~n3532 & n3555 ;
  assign n3568 = ~n3550 & ~n3566 ;
  assign n3569 = ~n3567 & n3568 ;
  assign n3570 = ~n3565 & ~n3569 ;
  assign n3571 = ~n3532 & ~n3553 ;
  assign n3572 = ~n3554 & ~n3571 ;
  assign n3573 = ~n3570 & ~n3572 ;
  assign n3574 = n3570 & n3572 ;
  assign n3575 = ~n3547 & ~n3560 ;
  assign n3576 = ~n3559 & ~n3575 ;
  assign n3577 = ~n3574 & ~n3576 ;
  assign n3578 = ~n3573 & ~n3577 ;
  assign n3579 = ~n3519 & n3578 ;
  assign n3580 = n3519 & ~n3578 ;
  assign n3581 = ~n3514 & ~n3517 ;
  assign n3582 = n3516 & ~n3581 ;
  assign n3583 = ~n3516 & n3581 ;
  assign n3584 = ~n3582 & ~n3583 ;
  assign n3585 = ~n3573 & ~n3574 ;
  assign n3586 = ~n3576 & n3585 ;
  assign n3587 = n3576 & ~n3585 ;
  assign n3588 = ~n3586 & ~n3587 ;
  assign n3589 = n3584 & ~n3588 ;
  assign n3590 = ~n3584 & n3588 ;
  assign n3591 = ~n3499 & ~n3501 ;
  assign n3592 = ~n3502 & ~n3591 ;
  assign n3593 = ~n3534 & ~n3549 ;
  assign n3594 = ~n3550 & ~n3593 ;
  assign n3595 = n3592 & n3594 ;
  assign n3596 = n3506 & ~n3509 ;
  assign n3597 = ~n3505 & ~n3507 ;
  assign n3598 = ~n3478 & ~n3597 ;
  assign n3599 = ~n3596 & ~n3598 ;
  assign n3600 = n3595 & n3599 ;
  assign n3601 = ~n3595 & ~n3599 ;
  assign n3602 = ~n3556 & ~n3569 ;
  assign n3603 = n3564 & n3602 ;
  assign n3604 = ~n3564 & ~n3602 ;
  assign n3605 = ~n3603 & ~n3604 ;
  assign n3606 = ~n3601 & ~n3605 ;
  assign n3607 = ~n3600 & ~n3606 ;
  assign n3608 = ~n3590 & ~n3607 ;
  assign n3609 = ~n3589 & ~n3608 ;
  assign n3610 = ~n3580 & ~n3609 ;
  assign n3611 = ~n3579 & ~n3610 ;
  assign n3612 = ~n3457 & ~n3611 ;
  assign n3613 = n3457 & n3611 ;
  assign n3614 = ~n3425 & ~n3426 ;
  assign n3615 = ~n3455 & n3614 ;
  assign n3616 = n3455 & ~n3614 ;
  assign n3617 = ~n3615 & ~n3616 ;
  assign n3618 = ~n3579 & ~n3580 ;
  assign n3619 = ~n3609 & n3618 ;
  assign n3620 = n3609 & ~n3618 ;
  assign n3621 = ~n3619 & ~n3620 ;
  assign n3622 = ~n3617 & ~n3621 ;
  assign n3623 = n3617 & n3621 ;
  assign n3624 = ~n3589 & ~n3590 ;
  assign n3625 = ~n3607 & n3624 ;
  assign n3626 = n3607 & ~n3624 ;
  assign n3627 = ~n3625 & ~n3626 ;
  assign n3628 = ~n3435 & ~n3436 ;
  assign n3629 = n3453 & n3628 ;
  assign n3630 = ~n3453 & ~n3628 ;
  assign n3631 = ~n3629 & ~n3630 ;
  assign n3632 = n3627 & n3631 ;
  assign n3633 = ~n3627 & ~n3631 ;
  assign n3634 = ~n3438 & ~n3440 ;
  assign n3635 = ~n3441 & ~n3634 ;
  assign n3636 = ~n3592 & ~n3594 ;
  assign n3637 = ~n3595 & ~n3636 ;
  assign n3638 = n3635 & n3637 ;
  assign n3639 = ~n3446 & ~n3451 ;
  assign n3640 = n3450 & ~n3639 ;
  assign n3641 = ~n3450 & n3639 ;
  assign n3642 = ~n3640 & ~n3641 ;
  assign n3643 = n3638 & ~n3642 ;
  assign n3644 = ~n3638 & n3642 ;
  assign n3645 = ~n3600 & ~n3601 ;
  assign n3646 = ~n3605 & n3645 ;
  assign n3647 = n3605 & ~n3645 ;
  assign n3648 = ~n3646 & ~n3647 ;
  assign n3649 = ~n3644 & n3648 ;
  assign n3650 = ~n3643 & ~n3649 ;
  assign n3651 = ~n3633 & ~n3650 ;
  assign n3652 = ~n3632 & ~n3651 ;
  assign n3653 = ~n3623 & n3652 ;
  assign n3654 = ~n3622 & ~n3653 ;
  assign n3655 = ~n3613 & n3654 ;
  assign n3656 = ~n3612 & ~n3655 ;
  assign n3657 = ~n3299 & ~n3656 ;
  assign n3658 = n3299 & n3656 ;
  assign n3659 = ~n3612 & ~n3613 ;
  assign n3660 = ~n3654 & n3659 ;
  assign n3661 = n3654 & ~n3659 ;
  assign n3662 = ~n3660 & ~n3661 ;
  assign n3663 = ~n3255 & ~n3256 ;
  assign n3664 = ~n3297 & n3663 ;
  assign n3665 = n3297 & ~n3663 ;
  assign n3666 = ~n3664 & ~n3665 ;
  assign n3667 = n3662 & ~n3666 ;
  assign n3668 = ~n3662 & n3666 ;
  assign n3669 = ~n3265 & ~n3266 ;
  assign n3670 = ~n3295 & n3669 ;
  assign n3671 = n3295 & ~n3669 ;
  assign n3672 = ~n3670 & ~n3671 ;
  assign n3673 = ~n3622 & ~n3623 ;
  assign n3674 = ~n3652 & n3673 ;
  assign n3675 = n3652 & ~n3673 ;
  assign n3676 = ~n3674 & ~n3675 ;
  assign n3677 = ~n3672 & ~n3676 ;
  assign n3678 = n3672 & n3676 ;
  assign n3679 = ~n3275 & ~n3276 ;
  assign n3680 = ~n3293 & n3679 ;
  assign n3681 = n3293 & ~n3679 ;
  assign n3682 = ~n3680 & ~n3681 ;
  assign n3683 = ~n3632 & ~n3633 ;
  assign n3684 = ~n3650 & n3683 ;
  assign n3685 = n3650 & ~n3683 ;
  assign n3686 = ~n3684 & ~n3685 ;
  assign n3687 = ~n3682 & ~n3686 ;
  assign n3688 = n3682 & n3686 ;
  assign n3689 = ~n3635 & ~n3637 ;
  assign n3690 = ~n3638 & ~n3689 ;
  assign n3691 = ~n3278 & ~n3280 ;
  assign n3692 = ~n3281 & ~n3691 ;
  assign n3693 = n3690 & n3692 ;
  assign n3694 = ~n3643 & ~n3644 ;
  assign n3695 = ~n3648 & n3694 ;
  assign n3696 = n3648 & ~n3694 ;
  assign n3697 = ~n3695 & ~n3696 ;
  assign n3698 = n3693 & ~n3697 ;
  assign n3699 = ~n3693 & n3697 ;
  assign n3700 = ~n3286 & ~n3287 ;
  assign n3701 = ~n3291 & n3700 ;
  assign n3702 = n3291 & ~n3700 ;
  assign n3703 = ~n3701 & ~n3702 ;
  assign n3704 = ~n3699 & ~n3703 ;
  assign n3705 = ~n3698 & ~n3704 ;
  assign n3706 = ~n3688 & n3705 ;
  assign n3707 = ~n3687 & ~n3706 ;
  assign n3708 = ~n3678 & ~n3707 ;
  assign n3709 = ~n3677 & ~n3708 ;
  assign n3710 = ~n3668 & ~n3709 ;
  assign n3711 = ~n3667 & ~n3710 ;
  assign n3712 = ~n3658 & n3711 ;
  assign n3713 = ~n3657 & ~n3712 ;
  assign n3714 = \A[355]  & \A[356]  ;
  assign n3715 = ~\A[355]  & ~\A[356]  ;
  assign n3716 = ~n3714 & ~n3715 ;
  assign n3717 = \A[357]  & n3716 ;
  assign n3718 = ~n3714 & ~n3717 ;
  assign n3719 = \A[358]  & \A[359]  ;
  assign n3720 = ~\A[357]  & ~n3716 ;
  assign n3721 = ~n3717 & ~n3720 ;
  assign n3722 = ~\A[358]  & ~\A[359]  ;
  assign n3723 = ~n3719 & ~n3722 ;
  assign n3724 = \A[360]  & n3723 ;
  assign n3725 = ~\A[360]  & ~n3723 ;
  assign n3726 = ~n3724 & ~n3725 ;
  assign n3727 = n3721 & n3726 ;
  assign n3728 = n3719 & n3727 ;
  assign n3729 = ~n3719 & ~n3724 ;
  assign n3730 = ~n3727 & n3729 ;
  assign n3731 = ~n3728 & ~n3730 ;
  assign n3732 = n3718 & ~n3731 ;
  assign n3733 = ~n3718 & n3731 ;
  assign n3734 = ~n3732 & ~n3733 ;
  assign n3735 = \A[361]  & \A[362]  ;
  assign n3736 = ~\A[361]  & ~\A[362]  ;
  assign n3737 = ~n3735 & ~n3736 ;
  assign n3738 = \A[363]  & n3737 ;
  assign n3739 = ~\A[363]  & ~n3737 ;
  assign n3740 = ~n3738 & ~n3739 ;
  assign n3741 = \A[364]  & \A[365]  ;
  assign n3742 = ~\A[364]  & ~\A[365]  ;
  assign n3743 = ~n3741 & ~n3742 ;
  assign n3744 = \A[366]  & n3743 ;
  assign n3745 = ~\A[366]  & ~n3743 ;
  assign n3746 = ~n3744 & ~n3745 ;
  assign n3747 = n3740 & n3746 ;
  assign n3748 = ~n3741 & ~n3744 ;
  assign n3749 = ~n3735 & ~n3738 ;
  assign n3750 = ~n3748 & ~n3749 ;
  assign n3751 = n3748 & n3749 ;
  assign n3752 = ~n3750 & ~n3751 ;
  assign n3759 = n3747 & ~n3752 ;
  assign n3753 = ~n3747 & n3752 ;
  assign n3754 = ~n3721 & ~n3726 ;
  assign n3755 = ~n3727 & ~n3754 ;
  assign n3756 = ~n3740 & ~n3746 ;
  assign n3757 = ~n3747 & ~n3756 ;
  assign n3758 = n3755 & n3757 ;
  assign n3760 = ~n3753 & ~n3758 ;
  assign n3761 = ~n3759 & n3760 ;
  assign n3762 = n3734 & ~n3761 ;
  assign n3763 = n3752 & n3758 ;
  assign n3764 = ~n3718 & n3728 ;
  assign n3765 = n3763 & ~n3764 ;
  assign n3766 = ~n3762 & ~n3765 ;
  assign n3767 = ~n3741 & n3749 ;
  assign n3768 = n3747 & ~n3767 ;
  assign n3769 = ~n3750 & ~n3768 ;
  assign n3770 = ~n3766 & ~n3769 ;
  assign n3771 = ~n3718 & ~n3730 ;
  assign n3772 = ~n3728 & ~n3771 ;
  assign n3773 = n3766 & n3769 ;
  assign n3774 = ~n3772 & ~n3773 ;
  assign n3775 = ~n3770 & ~n3774 ;
  assign n3776 = \A[349]  & \A[350]  ;
  assign n3777 = ~\A[349]  & ~\A[350]  ;
  assign n3778 = ~n3776 & ~n3777 ;
  assign n3779 = \A[351]  & n3778 ;
  assign n3780 = ~\A[351]  & ~n3778 ;
  assign n3781 = ~n3779 & ~n3780 ;
  assign n3782 = \A[352]  & \A[353]  ;
  assign n3783 = ~\A[352]  & ~\A[353]  ;
  assign n3784 = ~n3782 & ~n3783 ;
  assign n3785 = \A[354]  & n3784 ;
  assign n3786 = ~\A[354]  & ~n3784 ;
  assign n3787 = ~n3785 & ~n3786 ;
  assign n3788 = n3781 & n3787 ;
  assign n3789 = ~n3781 & ~n3787 ;
  assign n3790 = ~n3788 & ~n3789 ;
  assign n3791 = \A[343]  & \A[344]  ;
  assign n3792 = ~\A[343]  & ~\A[344]  ;
  assign n3793 = ~n3791 & ~n3792 ;
  assign n3794 = \A[345]  & n3793 ;
  assign n3795 = ~\A[345]  & ~n3793 ;
  assign n3796 = ~n3794 & ~n3795 ;
  assign n3797 = \A[346]  & \A[347]  ;
  assign n3798 = ~\A[346]  & ~\A[347]  ;
  assign n3799 = ~n3797 & ~n3798 ;
  assign n3800 = \A[348]  & n3799 ;
  assign n3801 = ~\A[348]  & ~n3799 ;
  assign n3802 = ~n3800 & ~n3801 ;
  assign n3803 = n3796 & n3802 ;
  assign n3804 = ~n3796 & ~n3802 ;
  assign n3805 = ~n3803 & ~n3804 ;
  assign n3806 = n3790 & n3805 ;
  assign n3807 = ~n3776 & ~n3779 ;
  assign n3808 = ~n3782 & ~n3785 ;
  assign n3809 = ~n3788 & n3808 ;
  assign n3810 = n3782 & n3788 ;
  assign n3811 = ~n3809 & ~n3810 ;
  assign n3812 = n3807 & ~n3811 ;
  assign n3813 = ~n3807 & n3811 ;
  assign n3814 = ~n3812 & ~n3813 ;
  assign n3815 = ~n3806 & ~n3814 ;
  assign n3816 = ~n3791 & ~n3794 ;
  assign n3817 = n3797 & n3803 ;
  assign n3818 = ~n3797 & ~n3800 ;
  assign n3819 = ~n3803 & n3818 ;
  assign n3820 = ~n3817 & ~n3819 ;
  assign n3821 = n3816 & ~n3820 ;
  assign n3822 = ~n3816 & n3820 ;
  assign n3823 = ~n3821 & ~n3822 ;
  assign n3824 = ~n3815 & n3823 ;
  assign n3825 = n3806 & n3814 ;
  assign n3826 = ~n3807 & ~n3808 ;
  assign n3827 = ~n3816 & n3817 ;
  assign n3828 = ~n3826 & ~n3827 ;
  assign n3829 = n3825 & n3828 ;
  assign n3830 = ~n3824 & ~n3829 ;
  assign n3831 = ~n3807 & ~n3809 ;
  assign n3832 = ~n3810 & ~n3831 ;
  assign n3833 = ~n3830 & ~n3832 ;
  assign n3834 = ~n3816 & ~n3819 ;
  assign n3835 = ~n3817 & ~n3834 ;
  assign n3836 = n3830 & n3832 ;
  assign n3837 = ~n3835 & ~n3836 ;
  assign n3838 = ~n3833 & ~n3837 ;
  assign n3839 = ~n3775 & ~n3838 ;
  assign n3840 = n3775 & n3838 ;
  assign n3841 = ~n3833 & ~n3836 ;
  assign n3842 = n3835 & ~n3841 ;
  assign n3843 = ~n3835 & n3841 ;
  assign n3844 = ~n3842 & ~n3843 ;
  assign n3845 = ~n3770 & ~n3773 ;
  assign n3846 = n3772 & ~n3845 ;
  assign n3847 = ~n3772 & n3845 ;
  assign n3848 = ~n3846 & ~n3847 ;
  assign n3849 = ~n3844 & ~n3848 ;
  assign n3850 = ~n3755 & ~n3757 ;
  assign n3851 = ~n3758 & ~n3850 ;
  assign n3852 = ~n3790 & ~n3805 ;
  assign n3853 = ~n3806 & ~n3852 ;
  assign n3854 = n3851 & n3853 ;
  assign n3855 = n3762 & ~n3765 ;
  assign n3856 = ~n3761 & ~n3763 ;
  assign n3857 = ~n3734 & ~n3856 ;
  assign n3858 = ~n3855 & ~n3857 ;
  assign n3859 = ~n3854 & ~n3858 ;
  assign n3860 = n3824 & ~n3829 ;
  assign n3861 = ~n3815 & ~n3825 ;
  assign n3862 = ~n3823 & ~n3861 ;
  assign n3863 = ~n3860 & ~n3862 ;
  assign n3864 = n3854 & n3858 ;
  assign n3865 = ~n3863 & ~n3864 ;
  assign n3866 = ~n3859 & ~n3865 ;
  assign n3867 = n3844 & n3848 ;
  assign n3868 = ~n3866 & ~n3867 ;
  assign n3869 = ~n3849 & ~n3868 ;
  assign n3870 = ~n3840 & n3869 ;
  assign n3871 = ~n3839 & ~n3870 ;
  assign n3872 = \A[331]  & \A[332]  ;
  assign n3873 = ~\A[331]  & ~\A[332]  ;
  assign n3874 = ~n3872 & ~n3873 ;
  assign n3875 = \A[333]  & n3874 ;
  assign n3876 = ~n3872 & ~n3875 ;
  assign n3877 = \A[334]  & \A[335]  ;
  assign n3878 = ~\A[333]  & ~n3874 ;
  assign n3879 = ~n3875 & ~n3878 ;
  assign n3880 = ~\A[334]  & ~\A[335]  ;
  assign n3881 = ~n3877 & ~n3880 ;
  assign n3882 = \A[336]  & n3881 ;
  assign n3883 = ~\A[336]  & ~n3881 ;
  assign n3884 = ~n3882 & ~n3883 ;
  assign n3885 = n3879 & n3884 ;
  assign n3886 = n3877 & n3885 ;
  assign n3887 = ~n3877 & ~n3882 ;
  assign n3888 = ~n3885 & n3887 ;
  assign n3889 = ~n3886 & ~n3888 ;
  assign n3890 = n3876 & ~n3889 ;
  assign n3891 = ~n3876 & n3889 ;
  assign n3892 = ~n3890 & ~n3891 ;
  assign n3893 = \A[337]  & \A[338]  ;
  assign n3894 = ~\A[337]  & ~\A[338]  ;
  assign n3895 = ~n3893 & ~n3894 ;
  assign n3896 = \A[339]  & n3895 ;
  assign n3897 = ~\A[339]  & ~n3895 ;
  assign n3898 = ~n3896 & ~n3897 ;
  assign n3899 = \A[340]  & \A[341]  ;
  assign n3900 = ~\A[340]  & ~\A[341]  ;
  assign n3901 = ~n3899 & ~n3900 ;
  assign n3902 = \A[342]  & n3901 ;
  assign n3903 = ~\A[342]  & ~n3901 ;
  assign n3904 = ~n3902 & ~n3903 ;
  assign n3905 = n3898 & n3904 ;
  assign n3906 = ~n3899 & ~n3902 ;
  assign n3907 = ~n3893 & ~n3896 ;
  assign n3908 = ~n3906 & ~n3907 ;
  assign n3909 = n3906 & n3907 ;
  assign n3910 = ~n3908 & ~n3909 ;
  assign n3917 = n3905 & ~n3910 ;
  assign n3911 = ~n3905 & n3910 ;
  assign n3912 = ~n3879 & ~n3884 ;
  assign n3913 = ~n3885 & ~n3912 ;
  assign n3914 = ~n3898 & ~n3904 ;
  assign n3915 = ~n3905 & ~n3914 ;
  assign n3916 = n3913 & n3915 ;
  assign n3918 = ~n3911 & ~n3916 ;
  assign n3919 = ~n3917 & n3918 ;
  assign n3920 = n3892 & ~n3919 ;
  assign n3921 = n3910 & n3916 ;
  assign n3922 = ~n3876 & n3886 ;
  assign n3923 = n3921 & ~n3922 ;
  assign n3924 = ~n3920 & ~n3923 ;
  assign n3925 = ~n3899 & n3907 ;
  assign n3926 = n3905 & ~n3925 ;
  assign n3927 = ~n3908 & ~n3926 ;
  assign n3928 = ~n3924 & ~n3927 ;
  assign n3929 = ~n3876 & ~n3888 ;
  assign n3930 = ~n3886 & ~n3929 ;
  assign n3931 = n3924 & n3927 ;
  assign n3932 = ~n3930 & ~n3931 ;
  assign n3933 = ~n3928 & ~n3932 ;
  assign n3934 = \A[325]  & \A[326]  ;
  assign n3935 = ~\A[325]  & ~\A[326]  ;
  assign n3936 = ~n3934 & ~n3935 ;
  assign n3937 = \A[327]  & n3936 ;
  assign n3938 = ~\A[327]  & ~n3936 ;
  assign n3939 = ~n3937 & ~n3938 ;
  assign n3940 = \A[328]  & \A[329]  ;
  assign n3941 = ~\A[328]  & ~\A[329]  ;
  assign n3942 = ~n3940 & ~n3941 ;
  assign n3943 = \A[330]  & n3942 ;
  assign n3944 = ~\A[330]  & ~n3942 ;
  assign n3945 = ~n3943 & ~n3944 ;
  assign n3946 = n3939 & n3945 ;
  assign n3947 = ~n3939 & ~n3945 ;
  assign n3948 = ~n3946 & ~n3947 ;
  assign n3949 = \A[319]  & \A[320]  ;
  assign n3950 = ~\A[319]  & ~\A[320]  ;
  assign n3951 = ~n3949 & ~n3950 ;
  assign n3952 = \A[321]  & n3951 ;
  assign n3953 = ~\A[321]  & ~n3951 ;
  assign n3954 = ~n3952 & ~n3953 ;
  assign n3955 = \A[322]  & \A[323]  ;
  assign n3956 = ~\A[322]  & ~\A[323]  ;
  assign n3957 = ~n3955 & ~n3956 ;
  assign n3958 = \A[324]  & n3957 ;
  assign n3959 = ~\A[324]  & ~n3957 ;
  assign n3960 = ~n3958 & ~n3959 ;
  assign n3961 = n3954 & n3960 ;
  assign n3962 = ~n3954 & ~n3960 ;
  assign n3963 = ~n3961 & ~n3962 ;
  assign n3964 = n3948 & n3963 ;
  assign n3965 = ~n3940 & ~n3943 ;
  assign n3966 = ~n3934 & ~n3937 ;
  assign n3967 = ~n3965 & ~n3966 ;
  assign n3968 = n3965 & n3966 ;
  assign n3969 = ~n3967 & ~n3968 ;
  assign n3970 = n3964 & n3969 ;
  assign n3971 = ~n3955 & ~n3958 ;
  assign n3972 = ~n3949 & ~n3952 ;
  assign n3973 = n3971 & n3972 ;
  assign n3974 = ~n3971 & ~n3972 ;
  assign n3975 = ~n3973 & ~n3974 ;
  assign n3976 = n3961 & ~n3975 ;
  assign n3977 = ~n3961 & n3975 ;
  assign n3978 = ~n3976 & ~n3977 ;
  assign n3979 = ~n3970 & n3978 ;
  assign n3981 = n3946 & ~n3969 ;
  assign n3980 = ~n3946 & n3969 ;
  assign n3982 = ~n3964 & ~n3980 ;
  assign n3983 = ~n3981 & n3982 ;
  assign n3984 = ~n3979 & ~n3983 ;
  assign n3985 = ~n3946 & ~n3967 ;
  assign n3986 = ~n3968 & ~n3985 ;
  assign n3987 = ~n3984 & ~n3986 ;
  assign n3988 = n3984 & n3986 ;
  assign n3989 = ~n3961 & ~n3974 ;
  assign n3990 = ~n3973 & ~n3989 ;
  assign n3991 = ~n3988 & ~n3990 ;
  assign n3992 = ~n3987 & ~n3991 ;
  assign n3993 = ~n3933 & n3992 ;
  assign n3994 = n3933 & ~n3992 ;
  assign n3995 = ~n3928 & ~n3931 ;
  assign n3996 = n3930 & ~n3995 ;
  assign n3997 = ~n3930 & n3995 ;
  assign n3998 = ~n3996 & ~n3997 ;
  assign n3999 = ~n3987 & ~n3988 ;
  assign n4000 = ~n3990 & n3999 ;
  assign n4001 = n3990 & ~n3999 ;
  assign n4002 = ~n4000 & ~n4001 ;
  assign n4003 = n3998 & ~n4002 ;
  assign n4004 = ~n3998 & n4002 ;
  assign n4005 = ~n3913 & ~n3915 ;
  assign n4006 = ~n3916 & ~n4005 ;
  assign n4007 = ~n3948 & ~n3963 ;
  assign n4008 = ~n3964 & ~n4007 ;
  assign n4009 = n4006 & n4008 ;
  assign n4010 = n3920 & ~n3923 ;
  assign n4011 = ~n3919 & ~n3921 ;
  assign n4012 = ~n3892 & ~n4011 ;
  assign n4013 = ~n4010 & ~n4012 ;
  assign n4014 = n4009 & n4013 ;
  assign n4015 = ~n4009 & ~n4013 ;
  assign n4016 = ~n3970 & ~n3983 ;
  assign n4017 = n3978 & n4016 ;
  assign n4018 = ~n3978 & ~n4016 ;
  assign n4019 = ~n4017 & ~n4018 ;
  assign n4020 = ~n4015 & ~n4019 ;
  assign n4021 = ~n4014 & ~n4020 ;
  assign n4022 = ~n4004 & ~n4021 ;
  assign n4023 = ~n4003 & ~n4022 ;
  assign n4024 = ~n3994 & ~n4023 ;
  assign n4025 = ~n3993 & ~n4024 ;
  assign n4026 = ~n3871 & ~n4025 ;
  assign n4027 = n3871 & n4025 ;
  assign n4028 = ~n3839 & ~n3840 ;
  assign n4029 = n3869 & ~n4028 ;
  assign n4030 = ~n3869 & n4028 ;
  assign n4031 = ~n4029 & ~n4030 ;
  assign n4032 = ~n3993 & ~n3994 ;
  assign n4033 = ~n4023 & n4032 ;
  assign n4034 = n4023 & ~n4032 ;
  assign n4035 = ~n4033 & ~n4034 ;
  assign n4036 = n4031 & ~n4035 ;
  assign n4037 = ~n4031 & n4035 ;
  assign n4038 = ~n3849 & ~n3867 ;
  assign n4039 = n3866 & n4038 ;
  assign n4040 = ~n3866 & ~n4038 ;
  assign n4041 = ~n4039 & ~n4040 ;
  assign n4042 = ~n4003 & ~n4004 ;
  assign n4043 = ~n4021 & n4042 ;
  assign n4044 = n4021 & ~n4042 ;
  assign n4045 = ~n4043 & ~n4044 ;
  assign n4046 = n4041 & n4045 ;
  assign n4047 = ~n4041 & ~n4045 ;
  assign n4048 = ~n3851 & ~n3853 ;
  assign n4049 = ~n3854 & ~n4048 ;
  assign n4050 = ~n4006 & ~n4008 ;
  assign n4051 = ~n4009 & ~n4050 ;
  assign n4052 = n4049 & n4051 ;
  assign n4053 = ~n3859 & ~n3864 ;
  assign n4054 = n3863 & ~n4053 ;
  assign n4055 = ~n3863 & n4053 ;
  assign n4056 = ~n4054 & ~n4055 ;
  assign n4057 = n4052 & ~n4056 ;
  assign n4058 = ~n4052 & n4056 ;
  assign n4059 = ~n4014 & ~n4015 ;
  assign n4060 = ~n4019 & n4059 ;
  assign n4061 = n4019 & ~n4059 ;
  assign n4062 = ~n4060 & ~n4061 ;
  assign n4063 = ~n4058 & n4062 ;
  assign n4064 = ~n4057 & ~n4063 ;
  assign n4065 = ~n4047 & ~n4064 ;
  assign n4066 = ~n4046 & ~n4065 ;
  assign n4067 = ~n4037 & n4066 ;
  assign n4068 = ~n4036 & ~n4067 ;
  assign n4069 = ~n4027 & n4068 ;
  assign n4070 = ~n4026 & ~n4069 ;
  assign n4071 = \A[301]  & \A[302]  ;
  assign n4072 = ~\A[301]  & ~\A[302]  ;
  assign n4073 = ~n4071 & ~n4072 ;
  assign n4074 = \A[303]  & n4073 ;
  assign n4075 = ~\A[303]  & ~n4073 ;
  assign n4076 = ~n4074 & ~n4075 ;
  assign n4077 = \A[304]  & \A[305]  ;
  assign n4078 = ~\A[304]  & ~\A[305]  ;
  assign n4079 = ~n4077 & ~n4078 ;
  assign n4080 = \A[306]  & n4079 ;
  assign n4081 = ~\A[306]  & ~n4079 ;
  assign n4082 = ~n4080 & ~n4081 ;
  assign n4083 = n4076 & n4082 ;
  assign n4084 = ~n4076 & ~n4082 ;
  assign n4085 = ~n4083 & ~n4084 ;
  assign n4086 = \A[295]  & \A[296]  ;
  assign n4087 = ~\A[295]  & ~\A[296]  ;
  assign n4088 = ~n4086 & ~n4087 ;
  assign n4089 = \A[297]  & n4088 ;
  assign n4090 = ~\A[297]  & ~n4088 ;
  assign n4091 = ~n4089 & ~n4090 ;
  assign n4092 = \A[298]  & \A[299]  ;
  assign n4093 = ~\A[298]  & ~\A[299]  ;
  assign n4094 = ~n4092 & ~n4093 ;
  assign n4095 = \A[300]  & n4094 ;
  assign n4096 = ~\A[300]  & ~n4094 ;
  assign n4097 = ~n4095 & ~n4096 ;
  assign n4098 = n4091 & n4097 ;
  assign n4099 = ~n4091 & ~n4097 ;
  assign n4100 = ~n4098 & ~n4099 ;
  assign n4101 = n4085 & n4100 ;
  assign n4102 = ~n4077 & ~n4080 ;
  assign n4103 = ~n4071 & ~n4074 ;
  assign n4104 = ~n4102 & ~n4103 ;
  assign n4105 = n4102 & n4103 ;
  assign n4106 = ~n4104 & ~n4105 ;
  assign n4107 = n4101 & n4106 ;
  assign n4108 = ~n4092 & ~n4095 ;
  assign n4109 = ~n4086 & ~n4089 ;
  assign n4110 = ~n4108 & ~n4109 ;
  assign n4111 = n4108 & n4109 ;
  assign n4112 = ~n4110 & ~n4111 ;
  assign n4113 = n4098 & ~n4112 ;
  assign n4114 = ~n4098 & n4112 ;
  assign n4115 = ~n4113 & ~n4114 ;
  assign n4116 = ~n4107 & n4115 ;
  assign n4118 = n4083 & ~n4106 ;
  assign n4117 = ~n4083 & n4106 ;
  assign n4119 = ~n4101 & ~n4117 ;
  assign n4120 = ~n4118 & n4119 ;
  assign n4121 = ~n4116 & ~n4120 ;
  assign n4122 = ~n4083 & ~n4104 ;
  assign n4123 = ~n4105 & ~n4122 ;
  assign n4124 = ~n4121 & ~n4123 ;
  assign n4125 = n4121 & n4123 ;
  assign n4126 = ~n4098 & ~n4110 ;
  assign n4127 = ~n4111 & ~n4126 ;
  assign n4128 = ~n4125 & ~n4127 ;
  assign n4129 = ~n4124 & ~n4128 ;
  assign n4130 = ~n4124 & ~n4125 ;
  assign n4131 = ~n4127 & n4130 ;
  assign n4132 = n4127 & ~n4130 ;
  assign n4133 = ~n4131 & ~n4132 ;
  assign n4134 = \A[313]  & \A[314]  ;
  assign n4135 = ~\A[313]  & ~\A[314]  ;
  assign n4136 = ~n4134 & ~n4135 ;
  assign n4137 = \A[315]  & n4136 ;
  assign n4138 = ~\A[315]  & ~n4136 ;
  assign n4139 = ~n4137 & ~n4138 ;
  assign n4140 = \A[316]  & \A[317]  ;
  assign n4141 = ~\A[316]  & ~\A[317]  ;
  assign n4142 = ~n4140 & ~n4141 ;
  assign n4143 = \A[318]  & n4142 ;
  assign n4144 = ~\A[318]  & ~n4142 ;
  assign n4145 = ~n4143 & ~n4144 ;
  assign n4146 = n4139 & n4145 ;
  assign n4147 = ~n4139 & ~n4145 ;
  assign n4148 = ~n4146 & ~n4147 ;
  assign n4149 = \A[307]  & \A[308]  ;
  assign n4150 = ~\A[307]  & ~\A[308]  ;
  assign n4151 = ~n4149 & ~n4150 ;
  assign n4152 = \A[309]  & n4151 ;
  assign n4153 = ~\A[309]  & ~n4151 ;
  assign n4154 = ~n4152 & ~n4153 ;
  assign n4155 = \A[310]  & \A[311]  ;
  assign n4156 = ~\A[310]  & ~\A[311]  ;
  assign n4157 = ~n4155 & ~n4156 ;
  assign n4158 = \A[312]  & n4157 ;
  assign n4159 = ~\A[312]  & ~n4157 ;
  assign n4160 = ~n4158 & ~n4159 ;
  assign n4161 = n4154 & n4160 ;
  assign n4162 = ~n4154 & ~n4160 ;
  assign n4163 = ~n4161 & ~n4162 ;
  assign n4164 = n4148 & n4163 ;
  assign n4165 = ~n4140 & ~n4143 ;
  assign n4166 = ~n4134 & ~n4137 ;
  assign n4167 = ~n4165 & ~n4166 ;
  assign n4168 = n4165 & n4166 ;
  assign n4169 = ~n4167 & ~n4168 ;
  assign n4170 = n4164 & n4169 ;
  assign n4171 = ~n4155 & ~n4158 ;
  assign n4172 = ~n4149 & ~n4152 ;
  assign n4173 = ~n4171 & ~n4172 ;
  assign n4174 = n4171 & n4172 ;
  assign n4175 = ~n4173 & ~n4174 ;
  assign n4176 = n4161 & ~n4175 ;
  assign n4177 = ~n4161 & n4175 ;
  assign n4178 = ~n4176 & ~n4177 ;
  assign n4179 = ~n4170 & n4178 ;
  assign n4181 = n4146 & ~n4169 ;
  assign n4180 = ~n4146 & n4169 ;
  assign n4182 = ~n4164 & ~n4180 ;
  assign n4183 = ~n4181 & n4182 ;
  assign n4184 = ~n4179 & ~n4183 ;
  assign n4185 = ~n4146 & ~n4167 ;
  assign n4186 = ~n4168 & ~n4185 ;
  assign n4187 = ~n4184 & ~n4186 ;
  assign n4188 = n4184 & n4186 ;
  assign n4189 = ~n4187 & ~n4188 ;
  assign n4190 = ~n4161 & ~n4173 ;
  assign n4191 = ~n4174 & ~n4190 ;
  assign n4192 = n4189 & ~n4191 ;
  assign n4193 = ~n4189 & n4191 ;
  assign n4194 = ~n4192 & ~n4193 ;
  assign n4195 = ~n4133 & ~n4194 ;
  assign n4196 = n4133 & n4194 ;
  assign n4197 = ~n4148 & ~n4163 ;
  assign n4198 = ~n4164 & ~n4197 ;
  assign n4199 = ~n4085 & ~n4100 ;
  assign n4200 = ~n4101 & ~n4199 ;
  assign n4201 = n4198 & n4200 ;
  assign n4202 = ~n4170 & ~n4183 ;
  assign n4203 = n4178 & n4202 ;
  assign n4204 = ~n4178 & ~n4202 ;
  assign n4205 = ~n4203 & ~n4204 ;
  assign n4206 = n4201 & ~n4205 ;
  assign n4207 = ~n4201 & n4205 ;
  assign n4208 = ~n4107 & ~n4120 ;
  assign n4209 = n4115 & n4208 ;
  assign n4210 = ~n4115 & ~n4208 ;
  assign n4211 = ~n4209 & ~n4210 ;
  assign n4212 = ~n4207 & ~n4211 ;
  assign n4213 = ~n4206 & ~n4212 ;
  assign n4214 = ~n4196 & ~n4213 ;
  assign n4215 = ~n4195 & ~n4214 ;
  assign n4216 = n4129 & ~n4215 ;
  assign n4217 = ~n4129 & n4215 ;
  assign n4218 = ~n4188 & ~n4191 ;
  assign n4219 = ~n4187 & ~n4218 ;
  assign n4220 = ~n4217 & n4219 ;
  assign n4221 = ~n4216 & ~n4220 ;
  assign n4222 = \A[277]  & \A[278]  ;
  assign n4223 = ~\A[277]  & ~\A[278]  ;
  assign n4224 = ~n4222 & ~n4223 ;
  assign n4225 = \A[279]  & n4224 ;
  assign n4226 = ~\A[279]  & ~n4224 ;
  assign n4227 = ~n4225 & ~n4226 ;
  assign n4228 = \A[280]  & \A[281]  ;
  assign n4229 = ~\A[280]  & ~\A[281]  ;
  assign n4230 = ~n4228 & ~n4229 ;
  assign n4231 = \A[282]  & n4230 ;
  assign n4232 = ~\A[282]  & ~n4230 ;
  assign n4233 = ~n4231 & ~n4232 ;
  assign n4234 = n4227 & n4233 ;
  assign n4235 = ~n4227 & ~n4233 ;
  assign n4236 = ~n4234 & ~n4235 ;
  assign n4237 = \A[271]  & \A[272]  ;
  assign n4238 = ~\A[271]  & ~\A[272]  ;
  assign n4239 = ~n4237 & ~n4238 ;
  assign n4240 = \A[273]  & n4239 ;
  assign n4241 = ~\A[273]  & ~n4239 ;
  assign n4242 = ~n4240 & ~n4241 ;
  assign n4243 = \A[274]  & \A[275]  ;
  assign n4244 = ~\A[274]  & ~\A[275]  ;
  assign n4245 = ~n4243 & ~n4244 ;
  assign n4246 = \A[276]  & n4245 ;
  assign n4247 = ~\A[276]  & ~n4245 ;
  assign n4248 = ~n4246 & ~n4247 ;
  assign n4249 = n4242 & n4248 ;
  assign n4250 = ~n4242 & ~n4248 ;
  assign n4251 = ~n4249 & ~n4250 ;
  assign n4252 = n4236 & n4251 ;
  assign n4253 = ~n4228 & ~n4231 ;
  assign n4254 = ~n4222 & ~n4225 ;
  assign n4255 = ~n4253 & ~n4254 ;
  assign n4256 = n4253 & n4254 ;
  assign n4257 = ~n4255 & ~n4256 ;
  assign n4258 = n4252 & n4257 ;
  assign n4259 = ~n4243 & ~n4246 ;
  assign n4260 = ~n4237 & ~n4240 ;
  assign n4261 = ~n4259 & ~n4260 ;
  assign n4262 = n4259 & n4260 ;
  assign n4263 = ~n4261 & ~n4262 ;
  assign n4264 = n4249 & ~n4263 ;
  assign n4265 = ~n4249 & n4263 ;
  assign n4266 = ~n4264 & ~n4265 ;
  assign n4267 = ~n4258 & n4266 ;
  assign n4269 = n4234 & ~n4257 ;
  assign n4268 = ~n4234 & n4257 ;
  assign n4270 = ~n4252 & ~n4268 ;
  assign n4271 = ~n4269 & n4270 ;
  assign n4272 = ~n4267 & ~n4271 ;
  assign n4273 = ~n4234 & ~n4255 ;
  assign n4274 = ~n4256 & ~n4273 ;
  assign n4275 = ~n4272 & ~n4274 ;
  assign n4276 = n4272 & n4274 ;
  assign n4277 = ~n4249 & ~n4261 ;
  assign n4278 = ~n4262 & ~n4277 ;
  assign n4279 = ~n4276 & ~n4278 ;
  assign n4280 = ~n4275 & ~n4279 ;
  assign n4281 = ~n4275 & ~n4276 ;
  assign n4282 = ~n4278 & n4281 ;
  assign n4283 = n4278 & ~n4281 ;
  assign n4284 = ~n4282 & ~n4283 ;
  assign n4285 = \A[289]  & \A[290]  ;
  assign n4286 = ~\A[289]  & ~\A[290]  ;
  assign n4287 = ~n4285 & ~n4286 ;
  assign n4288 = \A[291]  & n4287 ;
  assign n4289 = ~\A[291]  & ~n4287 ;
  assign n4290 = ~n4288 & ~n4289 ;
  assign n4291 = \A[292]  & \A[293]  ;
  assign n4292 = ~\A[292]  & ~\A[293]  ;
  assign n4293 = ~n4291 & ~n4292 ;
  assign n4294 = \A[294]  & n4293 ;
  assign n4295 = ~\A[294]  & ~n4293 ;
  assign n4296 = ~n4294 & ~n4295 ;
  assign n4297 = n4290 & n4296 ;
  assign n4298 = ~n4290 & ~n4296 ;
  assign n4299 = ~n4297 & ~n4298 ;
  assign n4300 = \A[283]  & \A[284]  ;
  assign n4301 = ~\A[283]  & ~\A[284]  ;
  assign n4302 = ~n4300 & ~n4301 ;
  assign n4303 = \A[285]  & n4302 ;
  assign n4304 = ~\A[285]  & ~n4302 ;
  assign n4305 = ~n4303 & ~n4304 ;
  assign n4306 = \A[286]  & \A[287]  ;
  assign n4307 = ~\A[286]  & ~\A[287]  ;
  assign n4308 = ~n4306 & ~n4307 ;
  assign n4309 = \A[288]  & n4308 ;
  assign n4310 = ~\A[288]  & ~n4308 ;
  assign n4311 = ~n4309 & ~n4310 ;
  assign n4312 = n4305 & n4311 ;
  assign n4313 = ~n4305 & ~n4311 ;
  assign n4314 = ~n4312 & ~n4313 ;
  assign n4315 = n4299 & n4314 ;
  assign n4316 = ~n4291 & ~n4294 ;
  assign n4317 = ~n4285 & ~n4288 ;
  assign n4318 = ~n4316 & ~n4317 ;
  assign n4319 = n4316 & n4317 ;
  assign n4320 = ~n4318 & ~n4319 ;
  assign n4321 = n4315 & n4320 ;
  assign n4322 = ~n4306 & ~n4309 ;
  assign n4323 = ~n4300 & ~n4303 ;
  assign n4324 = ~n4322 & ~n4323 ;
  assign n4325 = n4322 & n4323 ;
  assign n4326 = ~n4324 & ~n4325 ;
  assign n4327 = n4312 & ~n4326 ;
  assign n4328 = ~n4312 & n4326 ;
  assign n4329 = ~n4327 & ~n4328 ;
  assign n4330 = ~n4321 & n4329 ;
  assign n4332 = n4297 & ~n4320 ;
  assign n4331 = ~n4297 & n4320 ;
  assign n4333 = ~n4315 & ~n4331 ;
  assign n4334 = ~n4332 & n4333 ;
  assign n4335 = ~n4330 & ~n4334 ;
  assign n4336 = ~n4297 & ~n4318 ;
  assign n4337 = ~n4319 & ~n4336 ;
  assign n4338 = ~n4335 & ~n4337 ;
  assign n4339 = n4335 & n4337 ;
  assign n4340 = ~n4338 & ~n4339 ;
  assign n4341 = ~n4312 & ~n4324 ;
  assign n4342 = ~n4325 & ~n4341 ;
  assign n4343 = n4340 & ~n4342 ;
  assign n4344 = ~n4340 & n4342 ;
  assign n4345 = ~n4343 & ~n4344 ;
  assign n4346 = ~n4284 & ~n4345 ;
  assign n4347 = n4284 & n4345 ;
  assign n4348 = ~n4299 & ~n4314 ;
  assign n4349 = ~n4315 & ~n4348 ;
  assign n4350 = ~n4236 & ~n4251 ;
  assign n4351 = ~n4252 & ~n4350 ;
  assign n4352 = n4349 & n4351 ;
  assign n4353 = ~n4321 & ~n4334 ;
  assign n4354 = n4329 & n4353 ;
  assign n4355 = ~n4329 & ~n4353 ;
  assign n4356 = ~n4354 & ~n4355 ;
  assign n4357 = n4352 & ~n4356 ;
  assign n4358 = ~n4352 & n4356 ;
  assign n4359 = ~n4258 & ~n4271 ;
  assign n4360 = n4266 & n4359 ;
  assign n4361 = ~n4266 & ~n4359 ;
  assign n4362 = ~n4360 & ~n4361 ;
  assign n4363 = ~n4358 & ~n4362 ;
  assign n4364 = ~n4357 & ~n4363 ;
  assign n4365 = ~n4347 & ~n4364 ;
  assign n4366 = ~n4346 & ~n4365 ;
  assign n4367 = n4280 & ~n4366 ;
  assign n4368 = ~n4280 & n4366 ;
  assign n4369 = ~n4339 & ~n4342 ;
  assign n4370 = ~n4338 & ~n4369 ;
  assign n4371 = ~n4368 & n4370 ;
  assign n4372 = ~n4367 & ~n4371 ;
  assign n4373 = ~n4221 & ~n4372 ;
  assign n4374 = n4221 & n4372 ;
  assign n4375 = ~n4216 & ~n4217 ;
  assign n4376 = n4219 & n4375 ;
  assign n4377 = ~n4219 & ~n4375 ;
  assign n4378 = ~n4376 & ~n4377 ;
  assign n4379 = ~n4367 & ~n4368 ;
  assign n4380 = n4370 & n4379 ;
  assign n4381 = ~n4370 & ~n4379 ;
  assign n4382 = ~n4380 & ~n4381 ;
  assign n4383 = ~n4378 & ~n4382 ;
  assign n4384 = n4378 & n4382 ;
  assign n4385 = ~n4346 & ~n4347 ;
  assign n4386 = ~n4364 & n4385 ;
  assign n4387 = n4364 & ~n4385 ;
  assign n4388 = ~n4386 & ~n4387 ;
  assign n4389 = ~n4195 & ~n4196 ;
  assign n4390 = ~n4213 & n4389 ;
  assign n4391 = n4213 & ~n4389 ;
  assign n4392 = ~n4390 & ~n4391 ;
  assign n4393 = ~n4388 & ~n4392 ;
  assign n4394 = n4388 & n4392 ;
  assign n4395 = ~n4198 & ~n4200 ;
  assign n4396 = ~n4201 & ~n4395 ;
  assign n4397 = ~n4349 & ~n4351 ;
  assign n4398 = ~n4352 & ~n4397 ;
  assign n4399 = n4396 & n4398 ;
  assign n4400 = ~n4206 & ~n4207 ;
  assign n4401 = ~n4211 & n4400 ;
  assign n4402 = n4211 & ~n4400 ;
  assign n4403 = ~n4401 & ~n4402 ;
  assign n4404 = n4399 & n4403 ;
  assign n4405 = ~n4399 & ~n4403 ;
  assign n4406 = ~n4357 & ~n4358 ;
  assign n4407 = ~n4362 & n4406 ;
  assign n4408 = n4362 & ~n4406 ;
  assign n4409 = ~n4407 & ~n4408 ;
  assign n4410 = ~n4405 & n4409 ;
  assign n4411 = ~n4404 & ~n4410 ;
  assign n4412 = ~n4394 & n4411 ;
  assign n4413 = ~n4393 & ~n4412 ;
  assign n4414 = ~n4384 & ~n4413 ;
  assign n4415 = ~n4383 & ~n4414 ;
  assign n4416 = ~n4374 & n4415 ;
  assign n4417 = ~n4373 & ~n4416 ;
  assign n4418 = ~n4070 & ~n4417 ;
  assign n4419 = n4070 & n4417 ;
  assign n4420 = ~n4026 & ~n4027 ;
  assign n4421 = ~n4068 & n4420 ;
  assign n4422 = n4068 & ~n4420 ;
  assign n4423 = ~n4421 & ~n4422 ;
  assign n4424 = ~n4373 & ~n4374 ;
  assign n4425 = ~n4415 & n4424 ;
  assign n4426 = n4415 & ~n4424 ;
  assign n4427 = ~n4425 & ~n4426 ;
  assign n4428 = ~n4423 & ~n4427 ;
  assign n4429 = n4423 & n4427 ;
  assign n4430 = ~n4383 & ~n4384 ;
  assign n4431 = ~n4413 & n4430 ;
  assign n4432 = n4413 & ~n4430 ;
  assign n4433 = ~n4431 & ~n4432 ;
  assign n4434 = ~n4036 & ~n4037 ;
  assign n4435 = n4066 & n4434 ;
  assign n4436 = ~n4066 & ~n4434 ;
  assign n4437 = ~n4435 & ~n4436 ;
  assign n4438 = ~n4433 & ~n4437 ;
  assign n4439 = n4433 & n4437 ;
  assign n4440 = ~n4393 & ~n4394 ;
  assign n4441 = ~n4411 & n4440 ;
  assign n4442 = n4411 & ~n4440 ;
  assign n4443 = ~n4441 & ~n4442 ;
  assign n4444 = ~n4046 & ~n4047 ;
  assign n4445 = ~n4064 & n4444 ;
  assign n4446 = n4064 & ~n4444 ;
  assign n4447 = ~n4445 & ~n4446 ;
  assign n4448 = ~n4443 & ~n4447 ;
  assign n4449 = n4443 & n4447 ;
  assign n4450 = ~n4049 & ~n4051 ;
  assign n4451 = ~n4052 & ~n4450 ;
  assign n4452 = ~n4396 & ~n4398 ;
  assign n4453 = ~n4399 & ~n4452 ;
  assign n4454 = n4451 & n4453 ;
  assign n4455 = ~n4057 & ~n4058 ;
  assign n4456 = ~n4062 & n4455 ;
  assign n4457 = n4062 & ~n4455 ;
  assign n4458 = ~n4456 & ~n4457 ;
  assign n4459 = n4454 & ~n4458 ;
  assign n4460 = ~n4454 & n4458 ;
  assign n4461 = ~n4404 & ~n4405 ;
  assign n4462 = ~n4409 & n4461 ;
  assign n4463 = n4409 & ~n4461 ;
  assign n4464 = ~n4462 & ~n4463 ;
  assign n4465 = ~n4460 & ~n4464 ;
  assign n4466 = ~n4459 & ~n4465 ;
  assign n4467 = ~n4449 & n4466 ;
  assign n4468 = ~n4448 & ~n4467 ;
  assign n4469 = ~n4439 & n4468 ;
  assign n4470 = ~n4438 & ~n4469 ;
  assign n4471 = ~n4429 & ~n4470 ;
  assign n4472 = ~n4428 & ~n4471 ;
  assign n4473 = ~n4419 & ~n4472 ;
  assign n4474 = ~n4418 & ~n4473 ;
  assign n4475 = ~n3713 & ~n4474 ;
  assign n4476 = n3713 & n4474 ;
  assign n4477 = ~n3657 & ~n3658 ;
  assign n4478 = ~n3711 & n4477 ;
  assign n4479 = n3711 & ~n4477 ;
  assign n4480 = ~n4478 & ~n4479 ;
  assign n4481 = ~n4418 & ~n4419 ;
  assign n4482 = ~n4472 & n4481 ;
  assign n4483 = n4472 & ~n4481 ;
  assign n4484 = ~n4482 & ~n4483 ;
  assign n4485 = n4480 & ~n4484 ;
  assign n4486 = ~n4480 & n4484 ;
  assign n4487 = ~n4428 & ~n4429 ;
  assign n4488 = ~n4470 & n4487 ;
  assign n4489 = n4470 & ~n4487 ;
  assign n4490 = ~n4488 & ~n4489 ;
  assign n4491 = ~n3667 & ~n3668 ;
  assign n4492 = ~n3709 & n4491 ;
  assign n4493 = n3709 & ~n4491 ;
  assign n4494 = ~n4492 & ~n4493 ;
  assign n4495 = ~n4490 & n4494 ;
  assign n4496 = n4490 & ~n4494 ;
  assign n4497 = ~n3677 & ~n3678 ;
  assign n4498 = ~n3707 & n4497 ;
  assign n4499 = n3707 & ~n4497 ;
  assign n4500 = ~n4498 & ~n4499 ;
  assign n4501 = ~n4438 & ~n4439 ;
  assign n4502 = n4468 & n4501 ;
  assign n4503 = ~n4468 & ~n4501 ;
  assign n4504 = ~n4502 & ~n4503 ;
  assign n4505 = n4500 & ~n4504 ;
  assign n4506 = ~n4500 & n4504 ;
  assign n4507 = ~n4448 & ~n4449 ;
  assign n4508 = ~n4466 & n4507 ;
  assign n4509 = n4466 & ~n4507 ;
  assign n4510 = ~n4508 & ~n4509 ;
  assign n4511 = ~n3687 & ~n3688 ;
  assign n4512 = ~n3705 & n4511 ;
  assign n4513 = n3705 & ~n4511 ;
  assign n4514 = ~n4512 & ~n4513 ;
  assign n4515 = ~n4510 & ~n4514 ;
  assign n4516 = n4510 & n4514 ;
  assign n4517 = ~n3690 & ~n3692 ;
  assign n4518 = ~n3693 & ~n4517 ;
  assign n4519 = ~n4451 & ~n4453 ;
  assign n4520 = ~n4454 & ~n4519 ;
  assign n4521 = n4518 & n4520 ;
  assign n4522 = ~n3698 & ~n3699 ;
  assign n4523 = ~n3703 & n4522 ;
  assign n4524 = n3703 & ~n4522 ;
  assign n4525 = ~n4523 & ~n4524 ;
  assign n4526 = n4521 & n4525 ;
  assign n4527 = ~n4521 & ~n4525 ;
  assign n4528 = ~n4459 & ~n4460 ;
  assign n4529 = ~n4464 & n4528 ;
  assign n4530 = n4464 & ~n4528 ;
  assign n4531 = ~n4529 & ~n4530 ;
  assign n4532 = ~n4527 & n4531 ;
  assign n4533 = ~n4526 & ~n4532 ;
  assign n4534 = ~n4516 & n4533 ;
  assign n4535 = ~n4515 & ~n4534 ;
  assign n4536 = ~n4506 & ~n4535 ;
  assign n4537 = ~n4505 & ~n4536 ;
  assign n4538 = ~n4496 & ~n4537 ;
  assign n4539 = ~n4495 & ~n4538 ;
  assign n4540 = ~n4486 & ~n4539 ;
  assign n4541 = ~n4485 & ~n4540 ;
  assign n4542 = ~n4476 & n4541 ;
  assign n4543 = ~n4475 & ~n4542 ;
  assign n4544 = \A[211]  & \A[212]  ;
  assign n4545 = ~\A[211]  & ~\A[212]  ;
  assign n4546 = ~n4544 & ~n4545 ;
  assign n4547 = \A[213]  & n4546 ;
  assign n4548 = ~n4544 & ~n4547 ;
  assign n4549 = \A[214]  & \A[215]  ;
  assign n4550 = ~\A[213]  & ~n4546 ;
  assign n4551 = ~n4547 & ~n4550 ;
  assign n4552 = ~\A[214]  & ~\A[215]  ;
  assign n4553 = ~n4549 & ~n4552 ;
  assign n4554 = \A[216]  & n4553 ;
  assign n4555 = ~\A[216]  & ~n4553 ;
  assign n4556 = ~n4554 & ~n4555 ;
  assign n4557 = n4551 & n4556 ;
  assign n4558 = n4549 & n4557 ;
  assign n4559 = ~n4549 & ~n4554 ;
  assign n4560 = ~n4557 & n4559 ;
  assign n4561 = ~n4558 & ~n4560 ;
  assign n4562 = n4548 & ~n4561 ;
  assign n4563 = ~n4548 & n4561 ;
  assign n4564 = ~n4562 & ~n4563 ;
  assign n4565 = \A[217]  & \A[218]  ;
  assign n4566 = ~\A[217]  & ~\A[218]  ;
  assign n4567 = ~n4565 & ~n4566 ;
  assign n4568 = \A[219]  & n4567 ;
  assign n4569 = ~\A[219]  & ~n4567 ;
  assign n4570 = ~n4568 & ~n4569 ;
  assign n4571 = \A[220]  & \A[221]  ;
  assign n4572 = ~\A[220]  & ~\A[221]  ;
  assign n4573 = ~n4571 & ~n4572 ;
  assign n4574 = \A[222]  & n4573 ;
  assign n4575 = ~\A[222]  & ~n4573 ;
  assign n4576 = ~n4574 & ~n4575 ;
  assign n4577 = n4570 & n4576 ;
  assign n4578 = ~n4571 & ~n4574 ;
  assign n4579 = ~n4565 & ~n4568 ;
  assign n4580 = ~n4578 & ~n4579 ;
  assign n4581 = n4578 & n4579 ;
  assign n4582 = ~n4580 & ~n4581 ;
  assign n4589 = n4577 & ~n4582 ;
  assign n4583 = ~n4577 & n4582 ;
  assign n4584 = ~n4551 & ~n4556 ;
  assign n4585 = ~n4557 & ~n4584 ;
  assign n4586 = ~n4570 & ~n4576 ;
  assign n4587 = ~n4577 & ~n4586 ;
  assign n4588 = n4585 & n4587 ;
  assign n4590 = ~n4583 & ~n4588 ;
  assign n4591 = ~n4589 & n4590 ;
  assign n4592 = n4564 & ~n4591 ;
  assign n4593 = n4582 & n4588 ;
  assign n4594 = ~n4548 & n4558 ;
  assign n4595 = n4593 & ~n4594 ;
  assign n4596 = ~n4592 & ~n4595 ;
  assign n4597 = ~n4571 & n4579 ;
  assign n4598 = n4577 & ~n4597 ;
  assign n4599 = ~n4580 & ~n4598 ;
  assign n4600 = ~n4596 & ~n4599 ;
  assign n4601 = ~n4548 & ~n4560 ;
  assign n4602 = ~n4558 & ~n4601 ;
  assign n4603 = n4596 & n4599 ;
  assign n4604 = ~n4602 & ~n4603 ;
  assign n4605 = ~n4600 & ~n4604 ;
  assign n4606 = \A[205]  & \A[206]  ;
  assign n4607 = ~\A[205]  & ~\A[206]  ;
  assign n4608 = ~n4606 & ~n4607 ;
  assign n4609 = \A[207]  & n4608 ;
  assign n4610 = ~\A[207]  & ~n4608 ;
  assign n4611 = ~n4609 & ~n4610 ;
  assign n4612 = \A[208]  & \A[209]  ;
  assign n4613 = ~\A[208]  & ~\A[209]  ;
  assign n4614 = ~n4612 & ~n4613 ;
  assign n4615 = \A[210]  & n4614 ;
  assign n4616 = ~\A[210]  & ~n4614 ;
  assign n4617 = ~n4615 & ~n4616 ;
  assign n4618 = n4611 & n4617 ;
  assign n4619 = ~n4611 & ~n4617 ;
  assign n4620 = ~n4618 & ~n4619 ;
  assign n4621 = \A[199]  & \A[200]  ;
  assign n4622 = ~\A[199]  & ~\A[200]  ;
  assign n4623 = ~n4621 & ~n4622 ;
  assign n4624 = \A[201]  & n4623 ;
  assign n4625 = ~\A[201]  & ~n4623 ;
  assign n4626 = ~n4624 & ~n4625 ;
  assign n4627 = \A[202]  & \A[203]  ;
  assign n4628 = ~\A[202]  & ~\A[203]  ;
  assign n4629 = ~n4627 & ~n4628 ;
  assign n4630 = \A[204]  & n4629 ;
  assign n4631 = ~\A[204]  & ~n4629 ;
  assign n4632 = ~n4630 & ~n4631 ;
  assign n4633 = n4626 & n4632 ;
  assign n4634 = ~n4626 & ~n4632 ;
  assign n4635 = ~n4633 & ~n4634 ;
  assign n4636 = n4620 & n4635 ;
  assign n4637 = ~n4606 & ~n4609 ;
  assign n4638 = ~n4612 & ~n4615 ;
  assign n4639 = ~n4618 & n4638 ;
  assign n4640 = n4612 & n4618 ;
  assign n4641 = ~n4639 & ~n4640 ;
  assign n4642 = n4637 & ~n4641 ;
  assign n4643 = ~n4637 & n4641 ;
  assign n4644 = ~n4642 & ~n4643 ;
  assign n4645 = ~n4636 & ~n4644 ;
  assign n4646 = ~n4621 & ~n4624 ;
  assign n4647 = n4627 & n4633 ;
  assign n4648 = ~n4627 & ~n4630 ;
  assign n4649 = ~n4633 & n4648 ;
  assign n4650 = ~n4647 & ~n4649 ;
  assign n4651 = n4646 & ~n4650 ;
  assign n4652 = ~n4646 & n4650 ;
  assign n4653 = ~n4651 & ~n4652 ;
  assign n4654 = ~n4645 & n4653 ;
  assign n4655 = n4636 & n4644 ;
  assign n4656 = ~n4637 & ~n4638 ;
  assign n4657 = ~n4646 & n4647 ;
  assign n4658 = ~n4656 & ~n4657 ;
  assign n4659 = n4655 & n4658 ;
  assign n4660 = ~n4654 & ~n4659 ;
  assign n4661 = ~n4637 & ~n4639 ;
  assign n4662 = ~n4640 & ~n4661 ;
  assign n4663 = ~n4660 & ~n4662 ;
  assign n4664 = ~n4646 & ~n4649 ;
  assign n4665 = ~n4647 & ~n4664 ;
  assign n4666 = n4660 & n4662 ;
  assign n4667 = ~n4665 & ~n4666 ;
  assign n4668 = ~n4663 & ~n4667 ;
  assign n4669 = ~n4605 & ~n4668 ;
  assign n4670 = n4605 & n4668 ;
  assign n4671 = ~n4663 & ~n4666 ;
  assign n4672 = n4665 & ~n4671 ;
  assign n4673 = ~n4665 & n4671 ;
  assign n4674 = ~n4672 & ~n4673 ;
  assign n4675 = ~n4600 & ~n4603 ;
  assign n4676 = n4602 & ~n4675 ;
  assign n4677 = ~n4602 & n4675 ;
  assign n4678 = ~n4676 & ~n4677 ;
  assign n4679 = ~n4674 & ~n4678 ;
  assign n4680 = ~n4585 & ~n4587 ;
  assign n4681 = ~n4588 & ~n4680 ;
  assign n4682 = ~n4620 & ~n4635 ;
  assign n4683 = ~n4636 & ~n4682 ;
  assign n4684 = n4681 & n4683 ;
  assign n4685 = n4592 & ~n4595 ;
  assign n4686 = ~n4591 & ~n4593 ;
  assign n4687 = ~n4564 & ~n4686 ;
  assign n4688 = ~n4685 & ~n4687 ;
  assign n4689 = ~n4684 & ~n4688 ;
  assign n4690 = n4654 & ~n4659 ;
  assign n4691 = ~n4645 & ~n4655 ;
  assign n4692 = ~n4653 & ~n4691 ;
  assign n4693 = ~n4690 & ~n4692 ;
  assign n4694 = n4684 & n4688 ;
  assign n4695 = ~n4693 & ~n4694 ;
  assign n4696 = ~n4689 & ~n4695 ;
  assign n4697 = n4674 & n4678 ;
  assign n4698 = ~n4696 & ~n4697 ;
  assign n4699 = ~n4679 & ~n4698 ;
  assign n4700 = ~n4670 & n4699 ;
  assign n4701 = ~n4669 & ~n4700 ;
  assign n4702 = \A[193]  & \A[194]  ;
  assign n4703 = ~\A[193]  & ~\A[194]  ;
  assign n4704 = ~n4702 & ~n4703 ;
  assign n4705 = \A[195]  & n4704 ;
  assign n4706 = ~\A[195]  & ~n4704 ;
  assign n4707 = ~n4705 & ~n4706 ;
  assign n4708 = \A[196]  & \A[197]  ;
  assign n4709 = ~\A[196]  & ~\A[197]  ;
  assign n4710 = ~n4708 & ~n4709 ;
  assign n4711 = \A[198]  & n4710 ;
  assign n4712 = ~\A[198]  & ~n4710 ;
  assign n4713 = ~n4711 & ~n4712 ;
  assign n4714 = n4707 & n4713 ;
  assign n4715 = ~n4707 & ~n4713 ;
  assign n4716 = ~n4714 & ~n4715 ;
  assign n4717 = \A[187]  & \A[188]  ;
  assign n4718 = ~\A[187]  & ~\A[188]  ;
  assign n4719 = ~n4717 & ~n4718 ;
  assign n4720 = \A[189]  & n4719 ;
  assign n4721 = ~\A[189]  & ~n4719 ;
  assign n4722 = ~n4720 & ~n4721 ;
  assign n4723 = \A[190]  & \A[191]  ;
  assign n4724 = ~\A[190]  & ~\A[191]  ;
  assign n4725 = ~n4723 & ~n4724 ;
  assign n4726 = \A[192]  & n4725 ;
  assign n4727 = ~\A[192]  & ~n4725 ;
  assign n4728 = ~n4726 & ~n4727 ;
  assign n4729 = n4722 & n4728 ;
  assign n4730 = ~n4722 & ~n4728 ;
  assign n4731 = ~n4729 & ~n4730 ;
  assign n4732 = n4716 & n4731 ;
  assign n4733 = ~n4708 & ~n4711 ;
  assign n4734 = ~n4702 & ~n4705 ;
  assign n4735 = ~n4733 & ~n4734 ;
  assign n4736 = n4733 & n4734 ;
  assign n4737 = ~n4735 & ~n4736 ;
  assign n4738 = n4732 & n4737 ;
  assign n4739 = ~n4717 & ~n4720 ;
  assign n4740 = ~n4723 & ~n4726 ;
  assign n4741 = ~n4729 & n4740 ;
  assign n4742 = n4723 & n4729 ;
  assign n4743 = ~n4741 & ~n4742 ;
  assign n4744 = n4739 & ~n4743 ;
  assign n4745 = ~n4739 & n4743 ;
  assign n4746 = ~n4744 & ~n4745 ;
  assign n4747 = ~n4738 & ~n4746 ;
  assign n4749 = n4714 & ~n4737 ;
  assign n4748 = ~n4714 & n4737 ;
  assign n4750 = ~n4732 & ~n4748 ;
  assign n4751 = ~n4749 & n4750 ;
  assign n4752 = ~n4747 & ~n4751 ;
  assign n4753 = ~n4714 & ~n4735 ;
  assign n4754 = ~n4736 & ~n4753 ;
  assign n4755 = ~n4752 & ~n4754 ;
  assign n4756 = n4752 & n4754 ;
  assign n4757 = ~n4739 & ~n4741 ;
  assign n4758 = ~n4742 & ~n4757 ;
  assign n4759 = ~n4756 & n4758 ;
  assign n4760 = ~n4755 & ~n4759 ;
  assign n4761 = ~n4755 & ~n4756 ;
  assign n4762 = ~n4758 & n4761 ;
  assign n4763 = n4758 & ~n4761 ;
  assign n4764 = ~n4762 & ~n4763 ;
  assign n4765 = \A[178]  & \A[179]  ;
  assign n4766 = \A[175]  & \A[176]  ;
  assign n4767 = ~\A[175]  & ~\A[176]  ;
  assign n4768 = ~n4766 & ~n4767 ;
  assign n4769 = \A[177]  & n4768 ;
  assign n4770 = ~\A[177]  & ~n4768 ;
  assign n4771 = ~n4769 & ~n4770 ;
  assign n4772 = ~\A[178]  & ~\A[179]  ;
  assign n4773 = ~n4765 & ~n4772 ;
  assign n4774 = \A[180]  & n4773 ;
  assign n4775 = ~\A[180]  & ~n4773 ;
  assign n4776 = ~n4774 & ~n4775 ;
  assign n4777 = n4771 & n4776 ;
  assign n4778 = n4765 & n4777 ;
  assign n4779 = ~n4766 & ~n4769 ;
  assign n4780 = ~n4765 & ~n4774 ;
  assign n4781 = ~n4777 & n4780 ;
  assign n4782 = ~n4779 & ~n4781 ;
  assign n4783 = ~n4778 & ~n4782 ;
  assign n4784 = \A[181]  & \A[182]  ;
  assign n4785 = ~\A[181]  & ~\A[182]  ;
  assign n4786 = ~n4784 & ~n4785 ;
  assign n4787 = \A[183]  & n4786 ;
  assign n4788 = ~\A[183]  & ~n4786 ;
  assign n4789 = ~n4787 & ~n4788 ;
  assign n4790 = \A[184]  & \A[185]  ;
  assign n4791 = ~\A[184]  & ~\A[185]  ;
  assign n4792 = ~n4790 & ~n4791 ;
  assign n4793 = \A[186]  & n4792 ;
  assign n4794 = ~\A[186]  & ~n4792 ;
  assign n4795 = ~n4793 & ~n4794 ;
  assign n4796 = n4789 & n4795 ;
  assign n4797 = ~n4789 & ~n4795 ;
  assign n4798 = ~n4796 & ~n4797 ;
  assign n4799 = ~n4771 & ~n4776 ;
  assign n4800 = ~n4777 & ~n4799 ;
  assign n4801 = n4798 & n4800 ;
  assign n4802 = ~n4790 & ~n4793 ;
  assign n4803 = ~n4784 & ~n4787 ;
  assign n4804 = ~n4802 & ~n4803 ;
  assign n4805 = n4802 & n4803 ;
  assign n4806 = ~n4804 & ~n4805 ;
  assign n4807 = n4801 & n4806 ;
  assign n4808 = ~n4778 & ~n4781 ;
  assign n4809 = n4779 & ~n4808 ;
  assign n4810 = ~n4779 & n4808 ;
  assign n4811 = ~n4809 & ~n4810 ;
  assign n4812 = ~n4807 & ~n4811 ;
  assign n4814 = n4796 & ~n4806 ;
  assign n4813 = ~n4796 & n4806 ;
  assign n4815 = ~n4801 & ~n4813 ;
  assign n4816 = ~n4814 & n4815 ;
  assign n4817 = ~n4812 & ~n4816 ;
  assign n4818 = ~n4796 & ~n4804 ;
  assign n4819 = ~n4805 & ~n4818 ;
  assign n4820 = n4817 & n4819 ;
  assign n4821 = ~n4817 & ~n4819 ;
  assign n4822 = ~n4820 & ~n4821 ;
  assign n4823 = n4783 & ~n4822 ;
  assign n4824 = ~n4783 & n4822 ;
  assign n4825 = ~n4823 & ~n4824 ;
  assign n4826 = n4764 & n4825 ;
  assign n4827 = ~n4764 & ~n4825 ;
  assign n4828 = ~n4716 & ~n4731 ;
  assign n4829 = ~n4732 & ~n4828 ;
  assign n4830 = ~n4798 & ~n4800 ;
  assign n4831 = ~n4801 & ~n4830 ;
  assign n4832 = n4829 & n4831 ;
  assign n4833 = ~n4738 & ~n4751 ;
  assign n4834 = ~n4746 & n4833 ;
  assign n4835 = n4746 & ~n4833 ;
  assign n4836 = ~n4834 & ~n4835 ;
  assign n4837 = n4832 & ~n4836 ;
  assign n4838 = ~n4832 & n4836 ;
  assign n4839 = ~n4807 & ~n4816 ;
  assign n4840 = ~n4811 & n4839 ;
  assign n4841 = n4811 & ~n4839 ;
  assign n4842 = ~n4840 & ~n4841 ;
  assign n4843 = ~n4838 & ~n4842 ;
  assign n4844 = ~n4837 & ~n4843 ;
  assign n4845 = ~n4827 & ~n4844 ;
  assign n4846 = ~n4826 & ~n4845 ;
  assign n4847 = n4760 & ~n4846 ;
  assign n4848 = ~n4760 & n4846 ;
  assign n4849 = n4783 & ~n4820 ;
  assign n4850 = ~n4821 & ~n4849 ;
  assign n4851 = ~n4848 & n4850 ;
  assign n4852 = ~n4847 & ~n4851 ;
  assign n4853 = ~n4701 & ~n4852 ;
  assign n4854 = n4701 & n4852 ;
  assign n4855 = ~n4669 & ~n4670 ;
  assign n4856 = n4699 & ~n4855 ;
  assign n4857 = ~n4699 & n4855 ;
  assign n4858 = ~n4856 & ~n4857 ;
  assign n4859 = ~n4847 & ~n4848 ;
  assign n4860 = n4850 & n4859 ;
  assign n4861 = ~n4850 & ~n4859 ;
  assign n4862 = ~n4860 & ~n4861 ;
  assign n4863 = ~n4858 & n4862 ;
  assign n4864 = n4858 & ~n4862 ;
  assign n4865 = ~n4679 & ~n4697 ;
  assign n4866 = n4696 & n4865 ;
  assign n4867 = ~n4696 & ~n4865 ;
  assign n4868 = ~n4866 & ~n4867 ;
  assign n4869 = ~n4826 & ~n4827 ;
  assign n4870 = ~n4844 & n4869 ;
  assign n4871 = n4844 & ~n4869 ;
  assign n4872 = ~n4870 & ~n4871 ;
  assign n4873 = n4868 & n4872 ;
  assign n4874 = ~n4868 & ~n4872 ;
  assign n4875 = ~n4681 & ~n4683 ;
  assign n4876 = ~n4684 & ~n4875 ;
  assign n4877 = ~n4829 & ~n4831 ;
  assign n4878 = ~n4832 & ~n4877 ;
  assign n4879 = n4876 & n4878 ;
  assign n4880 = ~n4689 & ~n4694 ;
  assign n4881 = n4693 & ~n4880 ;
  assign n4882 = ~n4693 & n4880 ;
  assign n4883 = ~n4881 & ~n4882 ;
  assign n4884 = n4879 & ~n4883 ;
  assign n4885 = ~n4879 & n4883 ;
  assign n4886 = ~n4837 & ~n4838 ;
  assign n4887 = ~n4842 & n4886 ;
  assign n4888 = n4842 & ~n4886 ;
  assign n4889 = ~n4887 & ~n4888 ;
  assign n4890 = ~n4885 & n4889 ;
  assign n4891 = ~n4884 & ~n4890 ;
  assign n4892 = ~n4874 & ~n4891 ;
  assign n4893 = ~n4873 & ~n4892 ;
  assign n4894 = ~n4864 & ~n4893 ;
  assign n4895 = ~n4863 & ~n4894 ;
  assign n4896 = ~n4854 & ~n4895 ;
  assign n4897 = ~n4853 & ~n4896 ;
  assign n4898 = \A[259]  & \A[260]  ;
  assign n4899 = ~\A[259]  & ~\A[260]  ;
  assign n4900 = ~n4898 & ~n4899 ;
  assign n4901 = \A[261]  & n4900 ;
  assign n4902 = ~n4898 & ~n4901 ;
  assign n4903 = \A[262]  & \A[263]  ;
  assign n4904 = ~\A[261]  & ~n4900 ;
  assign n4905 = ~n4901 & ~n4904 ;
  assign n4906 = ~\A[262]  & ~\A[263]  ;
  assign n4907 = ~n4903 & ~n4906 ;
  assign n4908 = \A[264]  & n4907 ;
  assign n4909 = ~\A[264]  & ~n4907 ;
  assign n4910 = ~n4908 & ~n4909 ;
  assign n4911 = n4905 & n4910 ;
  assign n4912 = n4903 & n4911 ;
  assign n4913 = ~n4903 & ~n4908 ;
  assign n4914 = ~n4911 & n4913 ;
  assign n4915 = ~n4912 & ~n4914 ;
  assign n4916 = n4902 & ~n4915 ;
  assign n4917 = ~n4902 & n4915 ;
  assign n4918 = ~n4916 & ~n4917 ;
  assign n4919 = \A[265]  & \A[266]  ;
  assign n4920 = ~\A[265]  & ~\A[266]  ;
  assign n4921 = ~n4919 & ~n4920 ;
  assign n4922 = \A[267]  & n4921 ;
  assign n4923 = ~\A[267]  & ~n4921 ;
  assign n4924 = ~n4922 & ~n4923 ;
  assign n4925 = \A[268]  & \A[269]  ;
  assign n4926 = ~\A[268]  & ~\A[269]  ;
  assign n4927 = ~n4925 & ~n4926 ;
  assign n4928 = \A[270]  & n4927 ;
  assign n4929 = ~\A[270]  & ~n4927 ;
  assign n4930 = ~n4928 & ~n4929 ;
  assign n4931 = n4924 & n4930 ;
  assign n4932 = ~n4925 & ~n4928 ;
  assign n4933 = ~n4919 & ~n4922 ;
  assign n4934 = ~n4932 & ~n4933 ;
  assign n4935 = n4932 & n4933 ;
  assign n4936 = ~n4934 & ~n4935 ;
  assign n4943 = n4931 & ~n4936 ;
  assign n4937 = ~n4931 & n4936 ;
  assign n4938 = ~n4905 & ~n4910 ;
  assign n4939 = ~n4911 & ~n4938 ;
  assign n4940 = ~n4924 & ~n4930 ;
  assign n4941 = ~n4931 & ~n4940 ;
  assign n4942 = n4939 & n4941 ;
  assign n4944 = ~n4937 & ~n4942 ;
  assign n4945 = ~n4943 & n4944 ;
  assign n4946 = n4918 & ~n4945 ;
  assign n4947 = n4936 & n4942 ;
  assign n4948 = ~n4902 & n4912 ;
  assign n4949 = n4947 & ~n4948 ;
  assign n4950 = ~n4946 & ~n4949 ;
  assign n4951 = ~n4925 & n4933 ;
  assign n4952 = n4931 & ~n4951 ;
  assign n4953 = ~n4934 & ~n4952 ;
  assign n4954 = ~n4950 & ~n4953 ;
  assign n4955 = ~n4902 & ~n4914 ;
  assign n4956 = ~n4912 & ~n4955 ;
  assign n4957 = n4950 & n4953 ;
  assign n4958 = ~n4956 & ~n4957 ;
  assign n4959 = ~n4954 & ~n4958 ;
  assign n4960 = \A[253]  & \A[254]  ;
  assign n4961 = ~\A[253]  & ~\A[254]  ;
  assign n4962 = ~n4960 & ~n4961 ;
  assign n4963 = \A[255]  & n4962 ;
  assign n4964 = ~\A[255]  & ~n4962 ;
  assign n4965 = ~n4963 & ~n4964 ;
  assign n4966 = \A[256]  & \A[257]  ;
  assign n4967 = ~\A[256]  & ~\A[257]  ;
  assign n4968 = ~n4966 & ~n4967 ;
  assign n4969 = \A[258]  & n4968 ;
  assign n4970 = ~\A[258]  & ~n4968 ;
  assign n4971 = ~n4969 & ~n4970 ;
  assign n4972 = n4965 & n4971 ;
  assign n4973 = ~n4965 & ~n4971 ;
  assign n4974 = ~n4972 & ~n4973 ;
  assign n4975 = \A[247]  & \A[248]  ;
  assign n4976 = ~\A[247]  & ~\A[248]  ;
  assign n4977 = ~n4975 & ~n4976 ;
  assign n4978 = \A[249]  & n4977 ;
  assign n4979 = ~\A[249]  & ~n4977 ;
  assign n4980 = ~n4978 & ~n4979 ;
  assign n4981 = \A[250]  & \A[251]  ;
  assign n4982 = ~\A[250]  & ~\A[251]  ;
  assign n4983 = ~n4981 & ~n4982 ;
  assign n4984 = \A[252]  & n4983 ;
  assign n4985 = ~\A[252]  & ~n4983 ;
  assign n4986 = ~n4984 & ~n4985 ;
  assign n4987 = n4980 & n4986 ;
  assign n4988 = ~n4980 & ~n4986 ;
  assign n4989 = ~n4987 & ~n4988 ;
  assign n4990 = n4974 & n4989 ;
  assign n4991 = ~n4960 & ~n4963 ;
  assign n4992 = ~n4966 & ~n4969 ;
  assign n4993 = ~n4972 & n4992 ;
  assign n4994 = n4966 & n4972 ;
  assign n4995 = ~n4993 & ~n4994 ;
  assign n4996 = n4991 & ~n4995 ;
  assign n4997 = ~n4991 & n4995 ;
  assign n4998 = ~n4996 & ~n4997 ;
  assign n4999 = ~n4990 & ~n4998 ;
  assign n5000 = ~n4975 & ~n4978 ;
  assign n5001 = n4981 & n4987 ;
  assign n5002 = ~n4981 & ~n4984 ;
  assign n5003 = ~n4987 & n5002 ;
  assign n5004 = ~n5001 & ~n5003 ;
  assign n5005 = n5000 & ~n5004 ;
  assign n5006 = ~n5000 & n5004 ;
  assign n5007 = ~n5005 & ~n5006 ;
  assign n5008 = ~n4999 & n5007 ;
  assign n5009 = n4990 & n4998 ;
  assign n5010 = ~n4991 & ~n4992 ;
  assign n5011 = ~n5000 & n5001 ;
  assign n5012 = ~n5010 & ~n5011 ;
  assign n5013 = n5009 & n5012 ;
  assign n5014 = ~n5008 & ~n5013 ;
  assign n5015 = ~n4991 & ~n4993 ;
  assign n5016 = ~n4994 & ~n5015 ;
  assign n5017 = ~n5014 & ~n5016 ;
  assign n5018 = ~n5000 & ~n5003 ;
  assign n5019 = ~n5001 & ~n5018 ;
  assign n5020 = n5014 & n5016 ;
  assign n5021 = ~n5019 & ~n5020 ;
  assign n5022 = ~n5017 & ~n5021 ;
  assign n5023 = ~n4959 & ~n5022 ;
  assign n5024 = n4959 & n5022 ;
  assign n5025 = ~n5017 & ~n5020 ;
  assign n5026 = n5019 & ~n5025 ;
  assign n5027 = ~n5019 & n5025 ;
  assign n5028 = ~n5026 & ~n5027 ;
  assign n5029 = ~n4954 & ~n4957 ;
  assign n5030 = n4956 & ~n5029 ;
  assign n5031 = ~n4956 & n5029 ;
  assign n5032 = ~n5030 & ~n5031 ;
  assign n5033 = ~n5028 & ~n5032 ;
  assign n5034 = ~n4939 & ~n4941 ;
  assign n5035 = ~n4942 & ~n5034 ;
  assign n5036 = ~n4974 & ~n4989 ;
  assign n5037 = ~n4990 & ~n5036 ;
  assign n5038 = n5035 & n5037 ;
  assign n5039 = n4946 & ~n4949 ;
  assign n5040 = ~n4945 & ~n4947 ;
  assign n5041 = ~n4918 & ~n5040 ;
  assign n5042 = ~n5039 & ~n5041 ;
  assign n5043 = ~n5038 & ~n5042 ;
  assign n5044 = n5008 & ~n5013 ;
  assign n5045 = ~n4999 & ~n5009 ;
  assign n5046 = ~n5007 & ~n5045 ;
  assign n5047 = ~n5044 & ~n5046 ;
  assign n5048 = n5038 & n5042 ;
  assign n5049 = ~n5047 & ~n5048 ;
  assign n5050 = ~n5043 & ~n5049 ;
  assign n5051 = n5028 & n5032 ;
  assign n5052 = ~n5050 & ~n5051 ;
  assign n5053 = ~n5033 & ~n5052 ;
  assign n5054 = ~n5024 & n5053 ;
  assign n5055 = ~n5023 & ~n5054 ;
  assign n5056 = \A[235]  & \A[236]  ;
  assign n5057 = ~\A[235]  & ~\A[236]  ;
  assign n5058 = ~n5056 & ~n5057 ;
  assign n5059 = \A[237]  & n5058 ;
  assign n5060 = ~n5056 & ~n5059 ;
  assign n5061 = \A[238]  & \A[239]  ;
  assign n5062 = ~\A[237]  & ~n5058 ;
  assign n5063 = ~n5059 & ~n5062 ;
  assign n5064 = ~\A[238]  & ~\A[239]  ;
  assign n5065 = ~n5061 & ~n5064 ;
  assign n5066 = \A[240]  & n5065 ;
  assign n5067 = ~\A[240]  & ~n5065 ;
  assign n5068 = ~n5066 & ~n5067 ;
  assign n5069 = n5063 & n5068 ;
  assign n5070 = n5061 & n5069 ;
  assign n5071 = ~n5061 & ~n5066 ;
  assign n5072 = ~n5069 & n5071 ;
  assign n5073 = ~n5070 & ~n5072 ;
  assign n5074 = n5060 & ~n5073 ;
  assign n5075 = ~n5060 & n5073 ;
  assign n5076 = ~n5074 & ~n5075 ;
  assign n5077 = \A[241]  & \A[242]  ;
  assign n5078 = ~\A[241]  & ~\A[242]  ;
  assign n5079 = ~n5077 & ~n5078 ;
  assign n5080 = \A[243]  & n5079 ;
  assign n5081 = ~\A[243]  & ~n5079 ;
  assign n5082 = ~n5080 & ~n5081 ;
  assign n5083 = \A[244]  & \A[245]  ;
  assign n5084 = ~\A[244]  & ~\A[245]  ;
  assign n5085 = ~n5083 & ~n5084 ;
  assign n5086 = \A[246]  & n5085 ;
  assign n5087 = ~\A[246]  & ~n5085 ;
  assign n5088 = ~n5086 & ~n5087 ;
  assign n5089 = n5082 & n5088 ;
  assign n5090 = ~n5083 & ~n5086 ;
  assign n5091 = ~n5077 & ~n5080 ;
  assign n5092 = ~n5090 & ~n5091 ;
  assign n5093 = n5090 & n5091 ;
  assign n5094 = ~n5092 & ~n5093 ;
  assign n5101 = n5089 & ~n5094 ;
  assign n5095 = ~n5089 & n5094 ;
  assign n5096 = ~n5063 & ~n5068 ;
  assign n5097 = ~n5069 & ~n5096 ;
  assign n5098 = ~n5082 & ~n5088 ;
  assign n5099 = ~n5089 & ~n5098 ;
  assign n5100 = n5097 & n5099 ;
  assign n5102 = ~n5095 & ~n5100 ;
  assign n5103 = ~n5101 & n5102 ;
  assign n5104 = n5076 & ~n5103 ;
  assign n5105 = n5094 & n5100 ;
  assign n5106 = ~n5060 & n5070 ;
  assign n5107 = n5105 & ~n5106 ;
  assign n5108 = ~n5104 & ~n5107 ;
  assign n5109 = ~n5083 & n5091 ;
  assign n5110 = n5089 & ~n5109 ;
  assign n5111 = ~n5092 & ~n5110 ;
  assign n5112 = ~n5108 & ~n5111 ;
  assign n5113 = ~n5060 & ~n5072 ;
  assign n5114 = ~n5070 & ~n5113 ;
  assign n5115 = n5108 & n5111 ;
  assign n5116 = ~n5114 & ~n5115 ;
  assign n5117 = ~n5112 & ~n5116 ;
  assign n5118 = \A[229]  & \A[230]  ;
  assign n5119 = ~\A[229]  & ~\A[230]  ;
  assign n5120 = ~n5118 & ~n5119 ;
  assign n5121 = \A[231]  & n5120 ;
  assign n5122 = ~\A[231]  & ~n5120 ;
  assign n5123 = ~n5121 & ~n5122 ;
  assign n5124 = \A[232]  & \A[233]  ;
  assign n5125 = ~\A[232]  & ~\A[233]  ;
  assign n5126 = ~n5124 & ~n5125 ;
  assign n5127 = \A[234]  & n5126 ;
  assign n5128 = ~\A[234]  & ~n5126 ;
  assign n5129 = ~n5127 & ~n5128 ;
  assign n5130 = n5123 & n5129 ;
  assign n5131 = ~n5123 & ~n5129 ;
  assign n5132 = ~n5130 & ~n5131 ;
  assign n5133 = \A[223]  & \A[224]  ;
  assign n5134 = ~\A[223]  & ~\A[224]  ;
  assign n5135 = ~n5133 & ~n5134 ;
  assign n5136 = \A[225]  & n5135 ;
  assign n5137 = ~\A[225]  & ~n5135 ;
  assign n5138 = ~n5136 & ~n5137 ;
  assign n5139 = \A[226]  & \A[227]  ;
  assign n5140 = ~\A[226]  & ~\A[227]  ;
  assign n5141 = ~n5139 & ~n5140 ;
  assign n5142 = \A[228]  & n5141 ;
  assign n5143 = ~\A[228]  & ~n5141 ;
  assign n5144 = ~n5142 & ~n5143 ;
  assign n5145 = n5138 & n5144 ;
  assign n5146 = ~n5138 & ~n5144 ;
  assign n5147 = ~n5145 & ~n5146 ;
  assign n5148 = n5132 & n5147 ;
  assign n5149 = ~n5124 & ~n5127 ;
  assign n5150 = ~n5118 & ~n5121 ;
  assign n5151 = ~n5149 & ~n5150 ;
  assign n5152 = n5149 & n5150 ;
  assign n5153 = ~n5151 & ~n5152 ;
  assign n5154 = n5148 & n5153 ;
  assign n5155 = ~n5139 & ~n5142 ;
  assign n5156 = ~n5133 & ~n5136 ;
  assign n5157 = n5155 & n5156 ;
  assign n5158 = ~n5155 & ~n5156 ;
  assign n5159 = ~n5157 & ~n5158 ;
  assign n5160 = n5145 & ~n5159 ;
  assign n5161 = ~n5145 & n5159 ;
  assign n5162 = ~n5160 & ~n5161 ;
  assign n5163 = ~n5154 & n5162 ;
  assign n5165 = n5130 & ~n5153 ;
  assign n5164 = ~n5130 & n5153 ;
  assign n5166 = ~n5148 & ~n5164 ;
  assign n5167 = ~n5165 & n5166 ;
  assign n5168 = ~n5163 & ~n5167 ;
  assign n5169 = ~n5130 & ~n5151 ;
  assign n5170 = ~n5152 & ~n5169 ;
  assign n5171 = ~n5168 & ~n5170 ;
  assign n5172 = n5168 & n5170 ;
  assign n5173 = ~n5145 & ~n5158 ;
  assign n5174 = ~n5157 & ~n5173 ;
  assign n5175 = ~n5172 & ~n5174 ;
  assign n5176 = ~n5171 & ~n5175 ;
  assign n5177 = ~n5117 & n5176 ;
  assign n5178 = n5117 & ~n5176 ;
  assign n5179 = ~n5112 & ~n5115 ;
  assign n5180 = n5114 & ~n5179 ;
  assign n5181 = ~n5114 & n5179 ;
  assign n5182 = ~n5180 & ~n5181 ;
  assign n5183 = ~n5171 & ~n5172 ;
  assign n5184 = ~n5174 & n5183 ;
  assign n5185 = n5174 & ~n5183 ;
  assign n5186 = ~n5184 & ~n5185 ;
  assign n5187 = n5182 & ~n5186 ;
  assign n5188 = ~n5182 & n5186 ;
  assign n5189 = ~n5097 & ~n5099 ;
  assign n5190 = ~n5100 & ~n5189 ;
  assign n5191 = ~n5132 & ~n5147 ;
  assign n5192 = ~n5148 & ~n5191 ;
  assign n5193 = n5190 & n5192 ;
  assign n5194 = n5104 & ~n5107 ;
  assign n5195 = ~n5103 & ~n5105 ;
  assign n5196 = ~n5076 & ~n5195 ;
  assign n5197 = ~n5194 & ~n5196 ;
  assign n5198 = n5193 & n5197 ;
  assign n5199 = ~n5193 & ~n5197 ;
  assign n5200 = ~n5154 & ~n5167 ;
  assign n5201 = n5162 & n5200 ;
  assign n5202 = ~n5162 & ~n5200 ;
  assign n5203 = ~n5201 & ~n5202 ;
  assign n5204 = ~n5199 & ~n5203 ;
  assign n5205 = ~n5198 & ~n5204 ;
  assign n5206 = ~n5188 & ~n5205 ;
  assign n5207 = ~n5187 & ~n5206 ;
  assign n5208 = ~n5178 & ~n5207 ;
  assign n5209 = ~n5177 & ~n5208 ;
  assign n5210 = ~n5055 & ~n5209 ;
  assign n5211 = n5055 & n5209 ;
  assign n5212 = ~n5023 & ~n5024 ;
  assign n5213 = n5053 & ~n5212 ;
  assign n5214 = ~n5053 & n5212 ;
  assign n5215 = ~n5213 & ~n5214 ;
  assign n5216 = ~n5177 & ~n5178 ;
  assign n5217 = ~n5207 & n5216 ;
  assign n5218 = n5207 & ~n5216 ;
  assign n5219 = ~n5217 & ~n5218 ;
  assign n5220 = n5215 & ~n5219 ;
  assign n5221 = ~n5215 & n5219 ;
  assign n5222 = ~n5033 & ~n5051 ;
  assign n5223 = n5050 & n5222 ;
  assign n5224 = ~n5050 & ~n5222 ;
  assign n5225 = ~n5223 & ~n5224 ;
  assign n5226 = ~n5187 & ~n5188 ;
  assign n5227 = ~n5205 & n5226 ;
  assign n5228 = n5205 & ~n5226 ;
  assign n5229 = ~n5227 & ~n5228 ;
  assign n5230 = n5225 & n5229 ;
  assign n5231 = ~n5225 & ~n5229 ;
  assign n5232 = ~n5035 & ~n5037 ;
  assign n5233 = ~n5038 & ~n5232 ;
  assign n5234 = ~n5190 & ~n5192 ;
  assign n5235 = ~n5193 & ~n5234 ;
  assign n5236 = n5233 & n5235 ;
  assign n5237 = ~n5043 & ~n5048 ;
  assign n5238 = n5047 & ~n5237 ;
  assign n5239 = ~n5047 & n5237 ;
  assign n5240 = ~n5238 & ~n5239 ;
  assign n5241 = n5236 & ~n5240 ;
  assign n5242 = ~n5236 & n5240 ;
  assign n5243 = ~n5198 & ~n5199 ;
  assign n5244 = ~n5203 & n5243 ;
  assign n5245 = n5203 & ~n5243 ;
  assign n5246 = ~n5244 & ~n5245 ;
  assign n5247 = ~n5242 & n5246 ;
  assign n5248 = ~n5241 & ~n5247 ;
  assign n5249 = ~n5231 & ~n5248 ;
  assign n5250 = ~n5230 & ~n5249 ;
  assign n5251 = ~n5221 & n5250 ;
  assign n5252 = ~n5220 & ~n5251 ;
  assign n5253 = ~n5211 & n5252 ;
  assign n5254 = ~n5210 & ~n5253 ;
  assign n5255 = ~n4897 & ~n5254 ;
  assign n5256 = n4897 & n5254 ;
  assign n5257 = ~n5210 & ~n5211 ;
  assign n5258 = ~n5252 & n5257 ;
  assign n5259 = n5252 & ~n5257 ;
  assign n5260 = ~n5258 & ~n5259 ;
  assign n5261 = ~n4853 & ~n4854 ;
  assign n5262 = ~n4895 & n5261 ;
  assign n5263 = n4895 & ~n5261 ;
  assign n5264 = ~n5262 & ~n5263 ;
  assign n5265 = n5260 & ~n5264 ;
  assign n5266 = ~n5260 & n5264 ;
  assign n5267 = ~n4863 & ~n4864 ;
  assign n5268 = ~n4893 & n5267 ;
  assign n5269 = n4893 & ~n5267 ;
  assign n5270 = ~n5268 & ~n5269 ;
  assign n5271 = ~n5220 & ~n5221 ;
  assign n5272 = ~n5250 & n5271 ;
  assign n5273 = n5250 & ~n5271 ;
  assign n5274 = ~n5272 & ~n5273 ;
  assign n5275 = ~n5270 & ~n5274 ;
  assign n5276 = n5270 & n5274 ;
  assign n5277 = ~n4873 & ~n4874 ;
  assign n5278 = ~n4891 & n5277 ;
  assign n5279 = n4891 & ~n5277 ;
  assign n5280 = ~n5278 & ~n5279 ;
  assign n5281 = ~n5230 & ~n5231 ;
  assign n5282 = ~n5248 & n5281 ;
  assign n5283 = n5248 & ~n5281 ;
  assign n5284 = ~n5282 & ~n5283 ;
  assign n5285 = ~n5280 & ~n5284 ;
  assign n5286 = n5280 & n5284 ;
  assign n5287 = ~n5233 & ~n5235 ;
  assign n5288 = ~n5236 & ~n5287 ;
  assign n5289 = ~n4876 & ~n4878 ;
  assign n5290 = ~n4879 & ~n5289 ;
  assign n5291 = n5288 & n5290 ;
  assign n5292 = ~n5241 & ~n5242 ;
  assign n5293 = ~n5246 & n5292 ;
  assign n5294 = n5246 & ~n5292 ;
  assign n5295 = ~n5293 & ~n5294 ;
  assign n5296 = n5291 & ~n5295 ;
  assign n5297 = ~n5291 & n5295 ;
  assign n5298 = ~n4884 & ~n4885 ;
  assign n5299 = ~n4889 & n5298 ;
  assign n5300 = n4889 & ~n5298 ;
  assign n5301 = ~n5299 & ~n5300 ;
  assign n5302 = ~n5297 & ~n5301 ;
  assign n5303 = ~n5296 & ~n5302 ;
  assign n5304 = ~n5286 & n5303 ;
  assign n5305 = ~n5285 & ~n5304 ;
  assign n5306 = ~n5276 & ~n5305 ;
  assign n5307 = ~n5275 & ~n5306 ;
  assign n5308 = ~n5266 & ~n5307 ;
  assign n5309 = ~n5265 & ~n5308 ;
  assign n5310 = ~n5256 & n5309 ;
  assign n5311 = ~n5255 & ~n5310 ;
  assign n5312 = \A[145]  & \A[146]  ;
  assign n5313 = ~\A[145]  & ~\A[146]  ;
  assign n5314 = ~n5312 & ~n5313 ;
  assign n5315 = \A[147]  & n5314 ;
  assign n5316 = ~\A[147]  & ~n5314 ;
  assign n5317 = ~n5315 & ~n5316 ;
  assign n5318 = \A[148]  & \A[149]  ;
  assign n5319 = ~\A[148]  & ~\A[149]  ;
  assign n5320 = ~n5318 & ~n5319 ;
  assign n5321 = \A[150]  & n5320 ;
  assign n5322 = ~\A[150]  & ~n5320 ;
  assign n5323 = ~n5321 & ~n5322 ;
  assign n5324 = n5317 & n5323 ;
  assign n5325 = ~n5317 & ~n5323 ;
  assign n5326 = ~n5324 & ~n5325 ;
  assign n5327 = \A[139]  & \A[140]  ;
  assign n5328 = ~\A[139]  & ~\A[140]  ;
  assign n5329 = ~n5327 & ~n5328 ;
  assign n5330 = \A[141]  & n5329 ;
  assign n5331 = ~\A[141]  & ~n5329 ;
  assign n5332 = ~n5330 & ~n5331 ;
  assign n5333 = \A[142]  & \A[143]  ;
  assign n5334 = ~\A[142]  & ~\A[143]  ;
  assign n5335 = ~n5333 & ~n5334 ;
  assign n5336 = \A[144]  & n5335 ;
  assign n5337 = ~\A[144]  & ~n5335 ;
  assign n5338 = ~n5336 & ~n5337 ;
  assign n5339 = n5332 & n5338 ;
  assign n5340 = ~n5332 & ~n5338 ;
  assign n5341 = ~n5339 & ~n5340 ;
  assign n5342 = n5326 & n5341 ;
  assign n5343 = ~n5318 & ~n5321 ;
  assign n5344 = ~n5312 & ~n5315 ;
  assign n5345 = ~n5343 & ~n5344 ;
  assign n5346 = n5343 & n5344 ;
  assign n5347 = ~n5345 & ~n5346 ;
  assign n5348 = n5342 & n5347 ;
  assign n5349 = ~n5327 & ~n5330 ;
  assign n5350 = ~n5333 & ~n5336 ;
  assign n5351 = ~n5339 & n5350 ;
  assign n5352 = n5333 & n5339 ;
  assign n5353 = ~n5351 & ~n5352 ;
  assign n5354 = n5349 & ~n5353 ;
  assign n5355 = ~n5349 & n5353 ;
  assign n5356 = ~n5354 & ~n5355 ;
  assign n5357 = ~n5348 & ~n5356 ;
  assign n5359 = n5324 & ~n5347 ;
  assign n5358 = ~n5324 & n5347 ;
  assign n5360 = ~n5342 & ~n5358 ;
  assign n5361 = ~n5359 & n5360 ;
  assign n5362 = ~n5357 & ~n5361 ;
  assign n5363 = ~n5324 & ~n5345 ;
  assign n5364 = ~n5346 & ~n5363 ;
  assign n5365 = ~n5362 & ~n5364 ;
  assign n5366 = n5362 & n5364 ;
  assign n5367 = ~n5349 & ~n5351 ;
  assign n5368 = ~n5352 & ~n5367 ;
  assign n5369 = ~n5366 & n5368 ;
  assign n5370 = ~n5365 & ~n5369 ;
  assign n5371 = ~n5365 & ~n5366 ;
  assign n5372 = ~n5368 & n5371 ;
  assign n5373 = n5368 & ~n5371 ;
  assign n5374 = ~n5372 & ~n5373 ;
  assign n5375 = \A[130]  & \A[131]  ;
  assign n5376 = \A[127]  & \A[128]  ;
  assign n5377 = ~\A[127]  & ~\A[128]  ;
  assign n5378 = ~n5376 & ~n5377 ;
  assign n5379 = \A[129]  & n5378 ;
  assign n5380 = ~\A[129]  & ~n5378 ;
  assign n5381 = ~n5379 & ~n5380 ;
  assign n5382 = ~\A[130]  & ~\A[131]  ;
  assign n5383 = ~n5375 & ~n5382 ;
  assign n5384 = \A[132]  & n5383 ;
  assign n5385 = ~\A[132]  & ~n5383 ;
  assign n5386 = ~n5384 & ~n5385 ;
  assign n5387 = n5381 & n5386 ;
  assign n5388 = n5375 & n5387 ;
  assign n5389 = ~n5376 & ~n5379 ;
  assign n5390 = ~n5375 & ~n5384 ;
  assign n5391 = ~n5387 & n5390 ;
  assign n5392 = ~n5389 & ~n5391 ;
  assign n5393 = ~n5388 & ~n5392 ;
  assign n5394 = \A[133]  & \A[134]  ;
  assign n5395 = ~\A[133]  & ~\A[134]  ;
  assign n5396 = ~n5394 & ~n5395 ;
  assign n5397 = \A[135]  & n5396 ;
  assign n5398 = ~\A[135]  & ~n5396 ;
  assign n5399 = ~n5397 & ~n5398 ;
  assign n5400 = \A[136]  & \A[137]  ;
  assign n5401 = ~\A[136]  & ~\A[137]  ;
  assign n5402 = ~n5400 & ~n5401 ;
  assign n5403 = \A[138]  & n5402 ;
  assign n5404 = ~\A[138]  & ~n5402 ;
  assign n5405 = ~n5403 & ~n5404 ;
  assign n5406 = n5399 & n5405 ;
  assign n5407 = ~n5399 & ~n5405 ;
  assign n5408 = ~n5406 & ~n5407 ;
  assign n5409 = ~n5381 & ~n5386 ;
  assign n5410 = ~n5387 & ~n5409 ;
  assign n5411 = n5408 & n5410 ;
  assign n5412 = ~n5400 & ~n5403 ;
  assign n5413 = ~n5394 & ~n5397 ;
  assign n5414 = ~n5412 & ~n5413 ;
  assign n5415 = n5412 & n5413 ;
  assign n5416 = ~n5414 & ~n5415 ;
  assign n5417 = n5411 & n5416 ;
  assign n5418 = ~n5388 & ~n5391 ;
  assign n5419 = n5389 & ~n5418 ;
  assign n5420 = ~n5389 & n5418 ;
  assign n5421 = ~n5419 & ~n5420 ;
  assign n5422 = ~n5417 & ~n5421 ;
  assign n5424 = n5406 & ~n5416 ;
  assign n5423 = ~n5406 & n5416 ;
  assign n5425 = ~n5411 & ~n5423 ;
  assign n5426 = ~n5424 & n5425 ;
  assign n5427 = ~n5422 & ~n5426 ;
  assign n5428 = ~n5406 & ~n5414 ;
  assign n5429 = ~n5415 & ~n5428 ;
  assign n5430 = ~n5427 & ~n5429 ;
  assign n5431 = n5427 & n5429 ;
  assign n5432 = ~n5430 & ~n5431 ;
  assign n5433 = n5393 & ~n5432 ;
  assign n5434 = ~n5393 & n5432 ;
  assign n5435 = ~n5433 & ~n5434 ;
  assign n5436 = n5374 & n5435 ;
  assign n5437 = ~n5374 & ~n5435 ;
  assign n5438 = ~n5326 & ~n5341 ;
  assign n5439 = ~n5342 & ~n5438 ;
  assign n5440 = ~n5408 & ~n5410 ;
  assign n5441 = ~n5411 & ~n5440 ;
  assign n5442 = n5439 & n5441 ;
  assign n5443 = ~n5348 & ~n5361 ;
  assign n5444 = ~n5356 & n5443 ;
  assign n5445 = n5356 & ~n5443 ;
  assign n5446 = ~n5444 & ~n5445 ;
  assign n5447 = n5442 & ~n5446 ;
  assign n5448 = ~n5442 & n5446 ;
  assign n5449 = ~n5417 & ~n5426 ;
  assign n5450 = ~n5421 & n5449 ;
  assign n5451 = n5421 & ~n5449 ;
  assign n5452 = ~n5450 & ~n5451 ;
  assign n5453 = ~n5448 & ~n5452 ;
  assign n5454 = ~n5447 & ~n5453 ;
  assign n5455 = ~n5437 & ~n5454 ;
  assign n5456 = ~n5436 & ~n5455 ;
  assign n5457 = ~n5370 & n5456 ;
  assign n5458 = n5370 & ~n5456 ;
  assign n5459 = n5393 & ~n5431 ;
  assign n5460 = ~n5430 & ~n5459 ;
  assign n5461 = ~n5458 & ~n5460 ;
  assign n5462 = ~n5457 & ~n5461 ;
  assign n5463 = \A[169]  & \A[170]  ;
  assign n5464 = ~\A[169]  & ~\A[170]  ;
  assign n5465 = ~n5463 & ~n5464 ;
  assign n5466 = \A[171]  & n5465 ;
  assign n5467 = ~\A[171]  & ~n5465 ;
  assign n5468 = ~n5466 & ~n5467 ;
  assign n5469 = \A[172]  & \A[173]  ;
  assign n5470 = ~\A[172]  & ~\A[173]  ;
  assign n5471 = ~n5469 & ~n5470 ;
  assign n5472 = \A[174]  & n5471 ;
  assign n5473 = ~\A[174]  & ~n5471 ;
  assign n5474 = ~n5472 & ~n5473 ;
  assign n5475 = n5468 & n5474 ;
  assign n5476 = ~n5468 & ~n5474 ;
  assign n5477 = ~n5475 & ~n5476 ;
  assign n5478 = \A[163]  & \A[164]  ;
  assign n5479 = ~\A[163]  & ~\A[164]  ;
  assign n5480 = ~n5478 & ~n5479 ;
  assign n5481 = \A[165]  & n5480 ;
  assign n5482 = ~\A[165]  & ~n5480 ;
  assign n5483 = ~n5481 & ~n5482 ;
  assign n5484 = \A[166]  & \A[167]  ;
  assign n5485 = ~\A[166]  & ~\A[167]  ;
  assign n5486 = ~n5484 & ~n5485 ;
  assign n5487 = \A[168]  & n5486 ;
  assign n5488 = ~\A[168]  & ~n5486 ;
  assign n5489 = ~n5487 & ~n5488 ;
  assign n5490 = n5483 & n5489 ;
  assign n5491 = ~n5483 & ~n5489 ;
  assign n5492 = ~n5490 & ~n5491 ;
  assign n5493 = n5477 & n5492 ;
  assign n5494 = ~n5469 & ~n5472 ;
  assign n5495 = ~n5463 & ~n5466 ;
  assign n5496 = ~n5494 & ~n5495 ;
  assign n5497 = n5494 & n5495 ;
  assign n5498 = ~n5496 & ~n5497 ;
  assign n5499 = n5493 & n5498 ;
  assign n5500 = ~n5478 & ~n5481 ;
  assign n5501 = ~n5484 & ~n5487 ;
  assign n5502 = ~n5490 & n5501 ;
  assign n5503 = n5484 & n5490 ;
  assign n5504 = ~n5502 & ~n5503 ;
  assign n5505 = n5500 & ~n5504 ;
  assign n5506 = ~n5500 & n5504 ;
  assign n5507 = ~n5505 & ~n5506 ;
  assign n5508 = ~n5499 & ~n5507 ;
  assign n5510 = n5475 & ~n5498 ;
  assign n5509 = ~n5475 & n5498 ;
  assign n5511 = ~n5493 & ~n5509 ;
  assign n5512 = ~n5510 & n5511 ;
  assign n5513 = ~n5508 & ~n5512 ;
  assign n5514 = ~n5475 & ~n5496 ;
  assign n5515 = ~n5497 & ~n5514 ;
  assign n5516 = ~n5513 & ~n5515 ;
  assign n5517 = n5513 & n5515 ;
  assign n5518 = ~n5500 & ~n5502 ;
  assign n5519 = ~n5503 & ~n5518 ;
  assign n5520 = ~n5517 & n5519 ;
  assign n5521 = ~n5516 & ~n5520 ;
  assign n5522 = ~n5516 & ~n5517 ;
  assign n5523 = ~n5519 & n5522 ;
  assign n5524 = n5519 & ~n5522 ;
  assign n5525 = ~n5523 & ~n5524 ;
  assign n5526 = \A[154]  & \A[155]  ;
  assign n5527 = \A[151]  & \A[152]  ;
  assign n5528 = ~\A[151]  & ~\A[152]  ;
  assign n5529 = ~n5527 & ~n5528 ;
  assign n5530 = \A[153]  & n5529 ;
  assign n5531 = ~\A[153]  & ~n5529 ;
  assign n5532 = ~n5530 & ~n5531 ;
  assign n5533 = ~\A[154]  & ~\A[155]  ;
  assign n5534 = ~n5526 & ~n5533 ;
  assign n5535 = \A[156]  & n5534 ;
  assign n5536 = ~\A[156]  & ~n5534 ;
  assign n5537 = ~n5535 & ~n5536 ;
  assign n5538 = n5532 & n5537 ;
  assign n5539 = n5526 & n5538 ;
  assign n5540 = ~n5527 & ~n5530 ;
  assign n5541 = ~n5526 & ~n5535 ;
  assign n5542 = ~n5538 & n5541 ;
  assign n5543 = ~n5540 & ~n5542 ;
  assign n5544 = ~n5539 & ~n5543 ;
  assign n5545 = \A[157]  & \A[158]  ;
  assign n5546 = ~\A[157]  & ~\A[158]  ;
  assign n5547 = ~n5545 & ~n5546 ;
  assign n5548 = \A[159]  & n5547 ;
  assign n5549 = ~\A[159]  & ~n5547 ;
  assign n5550 = ~n5548 & ~n5549 ;
  assign n5551 = \A[160]  & \A[161]  ;
  assign n5552 = ~\A[160]  & ~\A[161]  ;
  assign n5553 = ~n5551 & ~n5552 ;
  assign n5554 = \A[162]  & n5553 ;
  assign n5555 = ~\A[162]  & ~n5553 ;
  assign n5556 = ~n5554 & ~n5555 ;
  assign n5557 = n5550 & n5556 ;
  assign n5558 = ~n5550 & ~n5556 ;
  assign n5559 = ~n5557 & ~n5558 ;
  assign n5560 = ~n5532 & ~n5537 ;
  assign n5561 = ~n5538 & ~n5560 ;
  assign n5562 = n5559 & n5561 ;
  assign n5563 = ~n5551 & ~n5554 ;
  assign n5564 = ~n5545 & ~n5548 ;
  assign n5565 = ~n5563 & ~n5564 ;
  assign n5566 = n5563 & n5564 ;
  assign n5567 = ~n5565 & ~n5566 ;
  assign n5568 = n5562 & n5567 ;
  assign n5569 = ~n5539 & ~n5542 ;
  assign n5570 = n5540 & ~n5569 ;
  assign n5571 = ~n5540 & n5569 ;
  assign n5572 = ~n5570 & ~n5571 ;
  assign n5573 = ~n5568 & ~n5572 ;
  assign n5575 = n5557 & ~n5567 ;
  assign n5574 = ~n5557 & n5567 ;
  assign n5576 = ~n5562 & ~n5574 ;
  assign n5577 = ~n5575 & n5576 ;
  assign n5578 = ~n5573 & ~n5577 ;
  assign n5579 = ~n5557 & ~n5565 ;
  assign n5580 = ~n5566 & ~n5579 ;
  assign n5581 = ~n5578 & ~n5580 ;
  assign n5582 = n5578 & n5580 ;
  assign n5583 = ~n5581 & ~n5582 ;
  assign n5584 = n5544 & ~n5583 ;
  assign n5585 = ~n5544 & n5583 ;
  assign n5586 = ~n5584 & ~n5585 ;
  assign n5587 = n5525 & n5586 ;
  assign n5588 = ~n5525 & ~n5586 ;
  assign n5589 = ~n5477 & ~n5492 ;
  assign n5590 = ~n5493 & ~n5589 ;
  assign n5591 = ~n5559 & ~n5561 ;
  assign n5592 = ~n5562 & ~n5591 ;
  assign n5593 = n5590 & n5592 ;
  assign n5594 = ~n5499 & ~n5512 ;
  assign n5595 = ~n5507 & n5594 ;
  assign n5596 = n5507 & ~n5594 ;
  assign n5597 = ~n5595 & ~n5596 ;
  assign n5598 = n5593 & ~n5597 ;
  assign n5599 = ~n5593 & n5597 ;
  assign n5600 = ~n5568 & ~n5577 ;
  assign n5601 = ~n5572 & n5600 ;
  assign n5602 = n5572 & ~n5600 ;
  assign n5603 = ~n5601 & ~n5602 ;
  assign n5604 = ~n5599 & ~n5603 ;
  assign n5605 = ~n5598 & ~n5604 ;
  assign n5606 = ~n5588 & ~n5605 ;
  assign n5607 = ~n5587 & ~n5606 ;
  assign n5608 = ~n5521 & n5607 ;
  assign n5609 = n5521 & ~n5607 ;
  assign n5610 = n5544 & ~n5582 ;
  assign n5611 = ~n5581 & ~n5610 ;
  assign n5612 = ~n5609 & ~n5611 ;
  assign n5613 = ~n5608 & ~n5612 ;
  assign n5614 = ~n5462 & ~n5613 ;
  assign n5615 = n5462 & n5613 ;
  assign n5616 = ~n5608 & ~n5609 ;
  assign n5617 = ~n5611 & n5616 ;
  assign n5618 = n5611 & ~n5616 ;
  assign n5619 = ~n5617 & ~n5618 ;
  assign n5620 = ~n5457 & ~n5458 ;
  assign n5621 = ~n5460 & n5620 ;
  assign n5622 = n5460 & ~n5620 ;
  assign n5623 = ~n5621 & ~n5622 ;
  assign n5624 = n5619 & n5623 ;
  assign n5625 = ~n5619 & ~n5623 ;
  assign n5626 = ~n5436 & ~n5437 ;
  assign n5627 = ~n5454 & n5626 ;
  assign n5628 = n5454 & ~n5626 ;
  assign n5629 = ~n5627 & ~n5628 ;
  assign n5630 = ~n5587 & ~n5588 ;
  assign n5631 = ~n5605 & n5630 ;
  assign n5632 = n5605 & ~n5630 ;
  assign n5633 = ~n5631 & ~n5632 ;
  assign n5634 = ~n5629 & ~n5633 ;
  assign n5635 = n5629 & n5633 ;
  assign n5636 = ~n5590 & ~n5592 ;
  assign n5637 = ~n5593 & ~n5636 ;
  assign n5638 = ~n5439 & ~n5441 ;
  assign n5639 = ~n5442 & ~n5638 ;
  assign n5640 = n5637 & n5639 ;
  assign n5641 = ~n5598 & ~n5599 ;
  assign n5642 = ~n5603 & n5641 ;
  assign n5643 = n5603 & ~n5641 ;
  assign n5644 = ~n5642 & ~n5643 ;
  assign n5645 = n5640 & n5644 ;
  assign n5646 = ~n5640 & ~n5644 ;
  assign n5647 = ~n5447 & ~n5448 ;
  assign n5648 = ~n5452 & n5647 ;
  assign n5649 = n5452 & ~n5647 ;
  assign n5650 = ~n5648 & ~n5649 ;
  assign n5651 = ~n5646 & n5650 ;
  assign n5652 = ~n5645 & ~n5651 ;
  assign n5653 = ~n5635 & n5652 ;
  assign n5654 = ~n5634 & ~n5653 ;
  assign n5655 = ~n5625 & ~n5654 ;
  assign n5656 = ~n5624 & ~n5655 ;
  assign n5657 = ~n5615 & ~n5656 ;
  assign n5658 = ~n5614 & ~n5657 ;
  assign n5659 = \A[97]  & \A[98]  ;
  assign n5660 = ~\A[97]  & ~\A[98]  ;
  assign n5661 = ~n5659 & ~n5660 ;
  assign n5662 = \A[99]  & n5661 ;
  assign n5663 = ~\A[99]  & ~n5661 ;
  assign n5664 = ~n5662 & ~n5663 ;
  assign n5665 = \A[100]  & \A[101]  ;
  assign n5666 = ~\A[100]  & ~\A[101]  ;
  assign n5667 = ~n5665 & ~n5666 ;
  assign n5668 = \A[102]  & n5667 ;
  assign n5669 = ~\A[102]  & ~n5667 ;
  assign n5670 = ~n5668 & ~n5669 ;
  assign n5671 = n5664 & n5670 ;
  assign n5672 = ~n5664 & ~n5670 ;
  assign n5673 = ~n5671 & ~n5672 ;
  assign n5674 = \A[91]  & \A[92]  ;
  assign n5675 = ~\A[91]  & ~\A[92]  ;
  assign n5676 = ~n5674 & ~n5675 ;
  assign n5677 = \A[93]  & n5676 ;
  assign n5678 = ~\A[93]  & ~n5676 ;
  assign n5679 = ~n5677 & ~n5678 ;
  assign n5680 = \A[94]  & \A[95]  ;
  assign n5681 = ~\A[94]  & ~\A[95]  ;
  assign n5682 = ~n5680 & ~n5681 ;
  assign n5683 = \A[96]  & n5682 ;
  assign n5684 = ~\A[96]  & ~n5682 ;
  assign n5685 = ~n5683 & ~n5684 ;
  assign n5686 = n5679 & n5685 ;
  assign n5687 = ~n5679 & ~n5685 ;
  assign n5688 = ~n5686 & ~n5687 ;
  assign n5689 = n5673 & n5688 ;
  assign n5690 = ~n5665 & ~n5668 ;
  assign n5691 = ~n5659 & ~n5662 ;
  assign n5692 = ~n5690 & ~n5691 ;
  assign n5693 = n5690 & n5691 ;
  assign n5694 = ~n5692 & ~n5693 ;
  assign n5695 = n5689 & n5694 ;
  assign n5696 = ~n5674 & ~n5677 ;
  assign n5697 = ~n5680 & ~n5683 ;
  assign n5698 = ~n5686 & n5697 ;
  assign n5699 = n5680 & n5686 ;
  assign n5700 = ~n5698 & ~n5699 ;
  assign n5701 = n5696 & ~n5700 ;
  assign n5702 = ~n5696 & n5700 ;
  assign n5703 = ~n5701 & ~n5702 ;
  assign n5704 = ~n5695 & ~n5703 ;
  assign n5706 = n5671 & ~n5694 ;
  assign n5705 = ~n5671 & n5694 ;
  assign n5707 = ~n5689 & ~n5705 ;
  assign n5708 = ~n5706 & n5707 ;
  assign n5709 = ~n5704 & ~n5708 ;
  assign n5710 = ~n5671 & ~n5692 ;
  assign n5711 = ~n5693 & ~n5710 ;
  assign n5712 = ~n5709 & ~n5711 ;
  assign n5713 = n5709 & n5711 ;
  assign n5714 = ~n5696 & ~n5698 ;
  assign n5715 = ~n5699 & ~n5714 ;
  assign n5716 = ~n5713 & n5715 ;
  assign n5717 = ~n5712 & ~n5716 ;
  assign n5718 = ~n5712 & ~n5713 ;
  assign n5719 = ~n5715 & n5718 ;
  assign n5720 = n5715 & ~n5718 ;
  assign n5721 = ~n5719 & ~n5720 ;
  assign n5722 = \A[82]  & \A[83]  ;
  assign n5723 = \A[79]  & \A[80]  ;
  assign n5724 = ~\A[79]  & ~\A[80]  ;
  assign n5725 = ~n5723 & ~n5724 ;
  assign n5726 = \A[81]  & n5725 ;
  assign n5727 = ~\A[81]  & ~n5725 ;
  assign n5728 = ~n5726 & ~n5727 ;
  assign n5729 = ~\A[82]  & ~\A[83]  ;
  assign n5730 = ~n5722 & ~n5729 ;
  assign n5731 = \A[84]  & n5730 ;
  assign n5732 = ~\A[84]  & ~n5730 ;
  assign n5733 = ~n5731 & ~n5732 ;
  assign n5734 = n5728 & n5733 ;
  assign n5735 = n5722 & n5734 ;
  assign n5736 = ~n5723 & ~n5726 ;
  assign n5737 = ~n5722 & ~n5731 ;
  assign n5738 = ~n5734 & n5737 ;
  assign n5739 = ~n5736 & ~n5738 ;
  assign n5740 = ~n5735 & ~n5739 ;
  assign n5741 = \A[85]  & \A[86]  ;
  assign n5742 = ~\A[85]  & ~\A[86]  ;
  assign n5743 = ~n5741 & ~n5742 ;
  assign n5744 = \A[87]  & n5743 ;
  assign n5745 = ~\A[87]  & ~n5743 ;
  assign n5746 = ~n5744 & ~n5745 ;
  assign n5747 = \A[88]  & \A[89]  ;
  assign n5748 = ~\A[88]  & ~\A[89]  ;
  assign n5749 = ~n5747 & ~n5748 ;
  assign n5750 = \A[90]  & n5749 ;
  assign n5751 = ~\A[90]  & ~n5749 ;
  assign n5752 = ~n5750 & ~n5751 ;
  assign n5753 = n5746 & n5752 ;
  assign n5754 = ~n5746 & ~n5752 ;
  assign n5755 = ~n5753 & ~n5754 ;
  assign n5756 = ~n5728 & ~n5733 ;
  assign n5757 = ~n5734 & ~n5756 ;
  assign n5758 = n5755 & n5757 ;
  assign n5759 = ~n5747 & ~n5750 ;
  assign n5760 = ~n5741 & ~n5744 ;
  assign n5761 = ~n5759 & ~n5760 ;
  assign n5762 = n5759 & n5760 ;
  assign n5763 = ~n5761 & ~n5762 ;
  assign n5764 = n5758 & n5763 ;
  assign n5765 = ~n5735 & ~n5738 ;
  assign n5766 = n5736 & ~n5765 ;
  assign n5767 = ~n5736 & n5765 ;
  assign n5768 = ~n5766 & ~n5767 ;
  assign n5769 = ~n5764 & ~n5768 ;
  assign n5771 = n5753 & ~n5763 ;
  assign n5770 = ~n5753 & n5763 ;
  assign n5772 = ~n5758 & ~n5770 ;
  assign n5773 = ~n5771 & n5772 ;
  assign n5774 = ~n5769 & ~n5773 ;
  assign n5775 = ~n5753 & ~n5761 ;
  assign n5776 = ~n5762 & ~n5775 ;
  assign n5777 = ~n5774 & ~n5776 ;
  assign n5778 = n5774 & n5776 ;
  assign n5779 = ~n5777 & ~n5778 ;
  assign n5780 = n5740 & ~n5779 ;
  assign n5781 = ~n5740 & n5779 ;
  assign n5782 = ~n5780 & ~n5781 ;
  assign n5783 = n5721 & n5782 ;
  assign n5784 = ~n5721 & ~n5782 ;
  assign n5785 = ~n5673 & ~n5688 ;
  assign n5786 = ~n5689 & ~n5785 ;
  assign n5787 = ~n5755 & ~n5757 ;
  assign n5788 = ~n5758 & ~n5787 ;
  assign n5789 = n5786 & n5788 ;
  assign n5790 = ~n5695 & ~n5708 ;
  assign n5791 = ~n5703 & n5790 ;
  assign n5792 = n5703 & ~n5790 ;
  assign n5793 = ~n5791 & ~n5792 ;
  assign n5794 = n5789 & ~n5793 ;
  assign n5795 = ~n5789 & n5793 ;
  assign n5796 = ~n5764 & ~n5773 ;
  assign n5797 = ~n5768 & n5796 ;
  assign n5798 = n5768 & ~n5796 ;
  assign n5799 = ~n5797 & ~n5798 ;
  assign n5800 = ~n5795 & ~n5799 ;
  assign n5801 = ~n5794 & ~n5800 ;
  assign n5802 = ~n5784 & ~n5801 ;
  assign n5803 = ~n5783 & ~n5802 ;
  assign n5804 = ~n5717 & n5803 ;
  assign n5805 = n5717 & ~n5803 ;
  assign n5806 = n5740 & ~n5778 ;
  assign n5807 = ~n5777 & ~n5806 ;
  assign n5808 = ~n5805 & ~n5807 ;
  assign n5809 = ~n5804 & ~n5808 ;
  assign n5810 = \A[121]  & \A[122]  ;
  assign n5811 = ~\A[121]  & ~\A[122]  ;
  assign n5812 = ~n5810 & ~n5811 ;
  assign n5813 = \A[123]  & n5812 ;
  assign n5814 = ~\A[123]  & ~n5812 ;
  assign n5815 = ~n5813 & ~n5814 ;
  assign n5816 = \A[124]  & \A[125]  ;
  assign n5817 = ~\A[124]  & ~\A[125]  ;
  assign n5818 = ~n5816 & ~n5817 ;
  assign n5819 = \A[126]  & n5818 ;
  assign n5820 = ~\A[126]  & ~n5818 ;
  assign n5821 = ~n5819 & ~n5820 ;
  assign n5822 = n5815 & n5821 ;
  assign n5823 = ~n5815 & ~n5821 ;
  assign n5824 = ~n5822 & ~n5823 ;
  assign n5825 = \A[115]  & \A[116]  ;
  assign n5826 = ~\A[115]  & ~\A[116]  ;
  assign n5827 = ~n5825 & ~n5826 ;
  assign n5828 = \A[117]  & n5827 ;
  assign n5829 = ~\A[117]  & ~n5827 ;
  assign n5830 = ~n5828 & ~n5829 ;
  assign n5831 = \A[118]  & \A[119]  ;
  assign n5832 = ~\A[118]  & ~\A[119]  ;
  assign n5833 = ~n5831 & ~n5832 ;
  assign n5834 = \A[120]  & n5833 ;
  assign n5835 = ~\A[120]  & ~n5833 ;
  assign n5836 = ~n5834 & ~n5835 ;
  assign n5837 = n5830 & n5836 ;
  assign n5838 = ~n5830 & ~n5836 ;
  assign n5839 = ~n5837 & ~n5838 ;
  assign n5840 = n5824 & n5839 ;
  assign n5841 = ~n5816 & ~n5819 ;
  assign n5842 = ~n5810 & ~n5813 ;
  assign n5843 = ~n5841 & ~n5842 ;
  assign n5844 = n5841 & n5842 ;
  assign n5845 = ~n5843 & ~n5844 ;
  assign n5846 = n5840 & n5845 ;
  assign n5847 = ~n5825 & ~n5828 ;
  assign n5848 = ~n5831 & ~n5834 ;
  assign n5849 = ~n5837 & n5848 ;
  assign n5850 = n5831 & n5837 ;
  assign n5851 = ~n5849 & ~n5850 ;
  assign n5852 = n5847 & ~n5851 ;
  assign n5853 = ~n5847 & n5851 ;
  assign n5854 = ~n5852 & ~n5853 ;
  assign n5855 = ~n5846 & ~n5854 ;
  assign n5857 = n5822 & ~n5845 ;
  assign n5856 = ~n5822 & n5845 ;
  assign n5858 = ~n5840 & ~n5856 ;
  assign n5859 = ~n5857 & n5858 ;
  assign n5860 = ~n5855 & ~n5859 ;
  assign n5861 = ~n5822 & ~n5843 ;
  assign n5862 = ~n5844 & ~n5861 ;
  assign n5863 = ~n5860 & ~n5862 ;
  assign n5864 = n5860 & n5862 ;
  assign n5865 = ~n5847 & ~n5849 ;
  assign n5866 = ~n5850 & ~n5865 ;
  assign n5867 = ~n5864 & n5866 ;
  assign n5868 = ~n5863 & ~n5867 ;
  assign n5869 = ~n5863 & ~n5864 ;
  assign n5870 = ~n5866 & n5869 ;
  assign n5871 = n5866 & ~n5869 ;
  assign n5872 = ~n5870 & ~n5871 ;
  assign n5873 = \A[106]  & \A[107]  ;
  assign n5874 = \A[103]  & \A[104]  ;
  assign n5875 = ~\A[103]  & ~\A[104]  ;
  assign n5876 = ~n5874 & ~n5875 ;
  assign n5877 = \A[105]  & n5876 ;
  assign n5878 = ~\A[105]  & ~n5876 ;
  assign n5879 = ~n5877 & ~n5878 ;
  assign n5880 = ~\A[106]  & ~\A[107]  ;
  assign n5881 = ~n5873 & ~n5880 ;
  assign n5882 = \A[108]  & n5881 ;
  assign n5883 = ~\A[108]  & ~n5881 ;
  assign n5884 = ~n5882 & ~n5883 ;
  assign n5885 = n5879 & n5884 ;
  assign n5886 = n5873 & n5885 ;
  assign n5887 = ~n5874 & ~n5877 ;
  assign n5888 = ~n5873 & ~n5882 ;
  assign n5889 = ~n5885 & n5888 ;
  assign n5890 = ~n5887 & ~n5889 ;
  assign n5891 = ~n5886 & ~n5890 ;
  assign n5892 = \A[109]  & \A[110]  ;
  assign n5893 = ~\A[109]  & ~\A[110]  ;
  assign n5894 = ~n5892 & ~n5893 ;
  assign n5895 = \A[111]  & n5894 ;
  assign n5896 = ~\A[111]  & ~n5894 ;
  assign n5897 = ~n5895 & ~n5896 ;
  assign n5898 = \A[112]  & \A[113]  ;
  assign n5899 = ~\A[112]  & ~\A[113]  ;
  assign n5900 = ~n5898 & ~n5899 ;
  assign n5901 = \A[114]  & n5900 ;
  assign n5902 = ~\A[114]  & ~n5900 ;
  assign n5903 = ~n5901 & ~n5902 ;
  assign n5904 = n5897 & n5903 ;
  assign n5905 = ~n5897 & ~n5903 ;
  assign n5906 = ~n5904 & ~n5905 ;
  assign n5907 = ~n5879 & ~n5884 ;
  assign n5908 = ~n5885 & ~n5907 ;
  assign n5909 = n5906 & n5908 ;
  assign n5910 = ~n5898 & ~n5901 ;
  assign n5911 = ~n5892 & ~n5895 ;
  assign n5912 = ~n5910 & ~n5911 ;
  assign n5913 = n5910 & n5911 ;
  assign n5914 = ~n5912 & ~n5913 ;
  assign n5915 = n5909 & n5914 ;
  assign n5916 = ~n5886 & ~n5889 ;
  assign n5917 = n5887 & ~n5916 ;
  assign n5918 = ~n5887 & n5916 ;
  assign n5919 = ~n5917 & ~n5918 ;
  assign n5920 = ~n5915 & ~n5919 ;
  assign n5922 = n5904 & ~n5914 ;
  assign n5921 = ~n5904 & n5914 ;
  assign n5923 = ~n5909 & ~n5921 ;
  assign n5924 = ~n5922 & n5923 ;
  assign n5925 = ~n5920 & ~n5924 ;
  assign n5926 = ~n5904 & ~n5912 ;
  assign n5927 = ~n5913 & ~n5926 ;
  assign n5928 = ~n5925 & ~n5927 ;
  assign n5929 = n5925 & n5927 ;
  assign n5930 = ~n5928 & ~n5929 ;
  assign n5931 = n5891 & ~n5930 ;
  assign n5932 = ~n5891 & n5930 ;
  assign n5933 = ~n5931 & ~n5932 ;
  assign n5934 = n5872 & n5933 ;
  assign n5935 = ~n5872 & ~n5933 ;
  assign n5936 = ~n5824 & ~n5839 ;
  assign n5937 = ~n5840 & ~n5936 ;
  assign n5938 = ~n5906 & ~n5908 ;
  assign n5939 = ~n5909 & ~n5938 ;
  assign n5940 = n5937 & n5939 ;
  assign n5941 = ~n5846 & ~n5859 ;
  assign n5942 = ~n5854 & n5941 ;
  assign n5943 = n5854 & ~n5941 ;
  assign n5944 = ~n5942 & ~n5943 ;
  assign n5945 = n5940 & ~n5944 ;
  assign n5946 = ~n5940 & n5944 ;
  assign n5947 = ~n5915 & ~n5924 ;
  assign n5948 = ~n5919 & n5947 ;
  assign n5949 = n5919 & ~n5947 ;
  assign n5950 = ~n5948 & ~n5949 ;
  assign n5951 = ~n5946 & ~n5950 ;
  assign n5952 = ~n5945 & ~n5951 ;
  assign n5953 = ~n5935 & ~n5952 ;
  assign n5954 = ~n5934 & ~n5953 ;
  assign n5955 = ~n5868 & n5954 ;
  assign n5956 = n5868 & ~n5954 ;
  assign n5957 = n5891 & ~n5929 ;
  assign n5958 = ~n5928 & ~n5957 ;
  assign n5959 = ~n5956 & ~n5958 ;
  assign n5960 = ~n5955 & ~n5959 ;
  assign n5961 = ~n5809 & ~n5960 ;
  assign n5962 = n5809 & n5960 ;
  assign n5963 = ~n5955 & ~n5956 ;
  assign n5964 = ~n5958 & n5963 ;
  assign n5965 = n5958 & ~n5963 ;
  assign n5966 = ~n5964 & ~n5965 ;
  assign n5967 = ~n5804 & ~n5805 ;
  assign n5968 = ~n5807 & n5967 ;
  assign n5969 = n5807 & ~n5967 ;
  assign n5970 = ~n5968 & ~n5969 ;
  assign n5971 = n5966 & n5970 ;
  assign n5972 = ~n5966 & ~n5970 ;
  assign n5973 = ~n5783 & ~n5784 ;
  assign n5974 = ~n5801 & n5973 ;
  assign n5975 = n5801 & ~n5973 ;
  assign n5976 = ~n5974 & ~n5975 ;
  assign n5977 = ~n5934 & ~n5935 ;
  assign n5978 = ~n5952 & n5977 ;
  assign n5979 = n5952 & ~n5977 ;
  assign n5980 = ~n5978 & ~n5979 ;
  assign n5981 = ~n5976 & ~n5980 ;
  assign n5982 = n5976 & n5980 ;
  assign n5983 = ~n5937 & ~n5939 ;
  assign n5984 = ~n5940 & ~n5983 ;
  assign n5985 = ~n5786 & ~n5788 ;
  assign n5986 = ~n5789 & ~n5985 ;
  assign n5987 = n5984 & n5986 ;
  assign n5988 = ~n5945 & ~n5946 ;
  assign n5989 = ~n5950 & n5988 ;
  assign n5990 = n5950 & ~n5988 ;
  assign n5991 = ~n5989 & ~n5990 ;
  assign n5992 = n5987 & n5991 ;
  assign n5993 = ~n5987 & ~n5991 ;
  assign n5994 = ~n5794 & ~n5795 ;
  assign n5995 = ~n5799 & n5994 ;
  assign n5996 = n5799 & ~n5994 ;
  assign n5997 = ~n5995 & ~n5996 ;
  assign n5998 = ~n5993 & n5997 ;
  assign n5999 = ~n5992 & ~n5998 ;
  assign n6000 = ~n5982 & n5999 ;
  assign n6001 = ~n5981 & ~n6000 ;
  assign n6002 = ~n5972 & ~n6001 ;
  assign n6003 = ~n5971 & ~n6002 ;
  assign n6004 = ~n5962 & ~n6003 ;
  assign n6005 = ~n5961 & ~n6004 ;
  assign n6006 = ~n5658 & ~n6005 ;
  assign n6007 = n5658 & n6005 ;
  assign n6008 = ~n5961 & ~n5962 ;
  assign n6009 = ~n6003 & n6008 ;
  assign n6010 = n6003 & ~n6008 ;
  assign n6011 = ~n6009 & ~n6010 ;
  assign n6012 = ~n5614 & ~n5615 ;
  assign n6013 = ~n5656 & n6012 ;
  assign n6014 = n5656 & ~n6012 ;
  assign n6015 = ~n6013 & ~n6014 ;
  assign n6016 = ~n6011 & ~n6015 ;
  assign n6017 = n6011 & n6015 ;
  assign n6018 = ~n5624 & ~n5625 ;
  assign n6019 = ~n5654 & n6018 ;
  assign n6020 = n5654 & ~n6018 ;
  assign n6021 = ~n6019 & ~n6020 ;
  assign n6022 = ~n5971 & ~n5972 ;
  assign n6023 = ~n6001 & n6022 ;
  assign n6024 = n6001 & ~n6022 ;
  assign n6025 = ~n6023 & ~n6024 ;
  assign n6026 = ~n6021 & ~n6025 ;
  assign n6027 = n6021 & n6025 ;
  assign n6028 = ~n5981 & ~n5982 ;
  assign n6029 = ~n5999 & n6028 ;
  assign n6030 = n5999 & ~n6028 ;
  assign n6031 = ~n6029 & ~n6030 ;
  assign n6032 = ~n5634 & ~n5635 ;
  assign n6033 = ~n5652 & n6032 ;
  assign n6034 = n5652 & ~n6032 ;
  assign n6035 = ~n6033 & ~n6034 ;
  assign n6036 = ~n6031 & ~n6035 ;
  assign n6037 = n6031 & n6035 ;
  assign n6038 = ~n5637 & ~n5639 ;
  assign n6039 = ~n5640 & ~n6038 ;
  assign n6040 = ~n5984 & ~n5986 ;
  assign n6041 = ~n5987 & ~n6040 ;
  assign n6042 = n6039 & n6041 ;
  assign n6043 = ~n5645 & ~n5646 ;
  assign n6044 = ~n5650 & n6043 ;
  assign n6045 = n5650 & ~n6043 ;
  assign n6046 = ~n6044 & ~n6045 ;
  assign n6047 = n6042 & ~n6046 ;
  assign n6048 = ~n6042 & n6046 ;
  assign n6049 = ~n5992 & ~n5993 ;
  assign n6050 = ~n5997 & n6049 ;
  assign n6051 = n5997 & ~n6049 ;
  assign n6052 = ~n6050 & ~n6051 ;
  assign n6053 = ~n6048 & ~n6052 ;
  assign n6054 = ~n6047 & ~n6053 ;
  assign n6055 = ~n6037 & n6054 ;
  assign n6056 = ~n6036 & ~n6055 ;
  assign n6057 = ~n6027 & n6056 ;
  assign n6058 = ~n6026 & ~n6057 ;
  assign n6059 = ~n6017 & ~n6058 ;
  assign n6060 = ~n6016 & ~n6059 ;
  assign n6061 = ~n6007 & n6060 ;
  assign n6062 = ~n6006 & ~n6061 ;
  assign n6063 = ~n5311 & n6062 ;
  assign n6064 = n5311 & ~n6062 ;
  assign n6065 = ~n6006 & ~n6007 ;
  assign n6066 = ~n6060 & n6065 ;
  assign n6067 = n6060 & ~n6065 ;
  assign n6068 = ~n6066 & ~n6067 ;
  assign n6069 = ~n5255 & ~n5256 ;
  assign n6070 = ~n5309 & n6069 ;
  assign n6071 = n5309 & ~n6069 ;
  assign n6072 = ~n6070 & ~n6071 ;
  assign n6073 = n6068 & ~n6072 ;
  assign n6074 = ~n6068 & n6072 ;
  assign n6075 = ~n6016 & ~n6017 ;
  assign n6076 = ~n6058 & n6075 ;
  assign n6077 = n6058 & ~n6075 ;
  assign n6078 = ~n6076 & ~n6077 ;
  assign n6079 = ~n5265 & ~n5266 ;
  assign n6080 = ~n5307 & n6079 ;
  assign n6081 = n5307 & ~n6079 ;
  assign n6082 = ~n6080 & ~n6081 ;
  assign n6083 = ~n6078 & n6082 ;
  assign n6084 = n6078 & ~n6082 ;
  assign n6085 = ~n5275 & ~n5276 ;
  assign n6086 = ~n5305 & n6085 ;
  assign n6087 = n5305 & ~n6085 ;
  assign n6088 = ~n6086 & ~n6087 ;
  assign n6089 = ~n6026 & ~n6027 ;
  assign n6090 = n6056 & n6089 ;
  assign n6091 = ~n6056 & ~n6089 ;
  assign n6092 = ~n6090 & ~n6091 ;
  assign n6093 = n6088 & ~n6092 ;
  assign n6094 = ~n6088 & n6092 ;
  assign n6095 = ~n6036 & ~n6037 ;
  assign n6096 = ~n6054 & n6095 ;
  assign n6097 = n6054 & ~n6095 ;
  assign n6098 = ~n6096 & ~n6097 ;
  assign n6099 = ~n5285 & ~n5286 ;
  assign n6100 = ~n5303 & n6099 ;
  assign n6101 = n5303 & ~n6099 ;
  assign n6102 = ~n6100 & ~n6101 ;
  assign n6103 = ~n6098 & ~n6102 ;
  assign n6104 = n6098 & n6102 ;
  assign n6105 = ~n5288 & ~n5290 ;
  assign n6106 = ~n5291 & ~n6105 ;
  assign n6107 = ~n6039 & ~n6041 ;
  assign n6108 = ~n6042 & ~n6107 ;
  assign n6109 = n6106 & n6108 ;
  assign n6110 = ~n5296 & ~n5297 ;
  assign n6111 = ~n5301 & n6110 ;
  assign n6112 = n5301 & ~n6110 ;
  assign n6113 = ~n6111 & ~n6112 ;
  assign n6114 = n6109 & n6113 ;
  assign n6115 = ~n6109 & ~n6113 ;
  assign n6116 = ~n6047 & ~n6048 ;
  assign n6117 = ~n6052 & n6116 ;
  assign n6118 = n6052 & ~n6116 ;
  assign n6119 = ~n6117 & ~n6118 ;
  assign n6120 = ~n6115 & n6119 ;
  assign n6121 = ~n6114 & ~n6120 ;
  assign n6122 = ~n6104 & n6121 ;
  assign n6123 = ~n6103 & ~n6122 ;
  assign n6124 = ~n6094 & ~n6123 ;
  assign n6125 = ~n6093 & ~n6124 ;
  assign n6126 = ~n6084 & ~n6125 ;
  assign n6127 = ~n6083 & ~n6126 ;
  assign n6128 = ~n6074 & n6127 ;
  assign n6129 = ~n6073 & ~n6128 ;
  assign n6130 = ~n6064 & ~n6129 ;
  assign n6131 = ~n6063 & ~n6130 ;
  assign n6132 = ~n4543 & ~n6131 ;
  assign n6133 = n4543 & n6131 ;
  assign n6134 = ~n4475 & ~n4476 ;
  assign n6135 = ~n4541 & n6134 ;
  assign n6136 = n4541 & ~n6134 ;
  assign n6137 = ~n6135 & ~n6136 ;
  assign n6138 = ~n6063 & ~n6064 ;
  assign n6139 = ~n6129 & n6138 ;
  assign n6140 = n6129 & ~n6138 ;
  assign n6141 = ~n6139 & ~n6140 ;
  assign n6142 = n6137 & ~n6141 ;
  assign n6143 = ~n6137 & n6141 ;
  assign n6144 = ~n6073 & ~n6074 ;
  assign n6145 = ~n6127 & n6144 ;
  assign n6146 = n6127 & ~n6144 ;
  assign n6147 = ~n6145 & ~n6146 ;
  assign n6148 = ~n4485 & ~n4486 ;
  assign n6149 = ~n4539 & n6148 ;
  assign n6150 = n4539 & ~n6148 ;
  assign n6151 = ~n6149 & ~n6150 ;
  assign n6152 = ~n6147 & ~n6151 ;
  assign n6153 = n6147 & n6151 ;
  assign n6154 = ~n6083 & ~n6084 ;
  assign n6155 = ~n6125 & n6154 ;
  assign n6156 = n6125 & ~n6154 ;
  assign n6157 = ~n6155 & ~n6156 ;
  assign n6158 = ~n4495 & ~n4496 ;
  assign n6159 = ~n4537 & n6158 ;
  assign n6160 = n4537 & ~n6158 ;
  assign n6161 = ~n6159 & ~n6160 ;
  assign n6162 = ~n6157 & ~n6161 ;
  assign n6163 = n6157 & n6161 ;
  assign n6164 = ~n4505 & ~n4506 ;
  assign n6165 = ~n4535 & n6164 ;
  assign n6166 = n4535 & ~n6164 ;
  assign n6167 = ~n6165 & ~n6166 ;
  assign n6168 = ~n6093 & ~n6094 ;
  assign n6169 = ~n6123 & n6168 ;
  assign n6170 = n6123 & ~n6168 ;
  assign n6171 = ~n6169 & ~n6170 ;
  assign n6172 = ~n6167 & ~n6171 ;
  assign n6173 = n6167 & n6171 ;
  assign n6174 = ~n6103 & ~n6104 ;
  assign n6175 = ~n6121 & n6174 ;
  assign n6176 = n6121 & ~n6174 ;
  assign n6177 = ~n6175 & ~n6176 ;
  assign n6178 = ~n4515 & ~n4516 ;
  assign n6179 = ~n4533 & n6178 ;
  assign n6180 = n4533 & ~n6178 ;
  assign n6181 = ~n6179 & ~n6180 ;
  assign n6182 = ~n6177 & ~n6181 ;
  assign n6183 = n6177 & n6181 ;
  assign n6184 = ~n4518 & ~n4520 ;
  assign n6185 = ~n4521 & ~n6184 ;
  assign n6186 = ~n6106 & ~n6108 ;
  assign n6187 = ~n6109 & ~n6186 ;
  assign n6188 = n6185 & n6187 ;
  assign n6189 = ~n4526 & ~n4527 ;
  assign n6190 = ~n4531 & n6189 ;
  assign n6191 = n4531 & ~n6189 ;
  assign n6192 = ~n6190 & ~n6191 ;
  assign n6193 = n6188 & ~n6192 ;
  assign n6194 = ~n6188 & n6192 ;
  assign n6195 = ~n6114 & ~n6115 ;
  assign n6196 = n6119 & n6195 ;
  assign n6197 = ~n6119 & ~n6195 ;
  assign n6198 = ~n6196 & ~n6197 ;
  assign n6199 = ~n6194 & n6198 ;
  assign n6200 = ~n6193 & ~n6199 ;
  assign n6201 = ~n6183 & n6200 ;
  assign n6202 = ~n6182 & ~n6201 ;
  assign n6203 = ~n6173 & n6202 ;
  assign n6204 = ~n6172 & ~n6203 ;
  assign n6205 = ~n6163 & ~n6204 ;
  assign n6206 = ~n6162 & ~n6205 ;
  assign n6207 = ~n6153 & ~n6206 ;
  assign n6208 = ~n6152 & ~n6207 ;
  assign n6209 = ~n6143 & n6208 ;
  assign n6210 = ~n6142 & ~n6209 ;
  assign n6211 = ~n6133 & n6210 ;
  assign n6212 = ~n6132 & ~n6211 ;
  assign n6213 = ~n2945 & n6212 ;
  assign n6214 = n2945 & ~n6212 ;
  assign n6215 = ~n6213 & ~n6214 ;
  assign n6216 = n2110 & n2877 ;
  assign n6217 = ~n2108 & ~n2944 ;
  assign n6218 = ~n2945 & ~n6217 ;
  assign n6219 = ~n6216 & ~n6218 ;
  assign n6220 = ~n6132 & ~n6133 ;
  assign n6221 = ~n6210 & n6220 ;
  assign n6222 = n6210 & ~n6220 ;
  assign n6223 = ~n6221 & ~n6222 ;
  assign n6224 = n6219 & n6223 ;
  assign n6225 = ~n6219 & ~n6223 ;
  assign n6226 = ~n2878 & ~n6216 ;
  assign n6227 = ~n2943 & n6226 ;
  assign n6228 = n2943 & ~n6226 ;
  assign n6229 = ~n6227 & ~n6228 ;
  assign n6230 = ~n6142 & ~n6143 ;
  assign n6231 = ~n6208 & n6230 ;
  assign n6232 = n6208 & ~n6230 ;
  assign n6233 = ~n6231 & ~n6232 ;
  assign n6234 = n6229 & ~n6233 ;
  assign n6235 = ~n6229 & n6233 ;
  assign n6236 = ~n2887 & ~n2888 ;
  assign n6237 = ~n2941 & n6236 ;
  assign n6238 = n2941 & ~n6236 ;
  assign n6239 = ~n6237 & ~n6238 ;
  assign n6240 = ~n6152 & ~n6153 ;
  assign n6241 = ~n6206 & n6240 ;
  assign n6242 = n6206 & ~n6240 ;
  assign n6243 = ~n6241 & ~n6242 ;
  assign n6244 = n6239 & ~n6243 ;
  assign n6245 = ~n6239 & n6243 ;
  assign n6246 = ~n2897 & ~n2898 ;
  assign n6247 = ~n2939 & n6246 ;
  assign n6248 = n2939 & ~n6246 ;
  assign n6249 = ~n6247 & ~n6248 ;
  assign n6250 = ~n6162 & ~n6163 ;
  assign n6251 = ~n6204 & n6250 ;
  assign n6252 = n6204 & ~n6250 ;
  assign n6253 = ~n6251 & ~n6252 ;
  assign n6254 = n6249 & ~n6253 ;
  assign n6255 = ~n6249 & n6253 ;
  assign n6256 = ~n6172 & ~n6173 ;
  assign n6257 = ~n6202 & n6256 ;
  assign n6258 = n6202 & ~n6256 ;
  assign n6259 = ~n6257 & ~n6258 ;
  assign n6260 = ~n2907 & ~n2908 ;
  assign n6261 = ~n2937 & n6260 ;
  assign n6262 = n2937 & ~n6260 ;
  assign n6263 = ~n6261 & ~n6262 ;
  assign n6264 = ~n6259 & ~n6263 ;
  assign n6265 = n6259 & n6263 ;
  assign n6266 = ~n2917 & ~n2918 ;
  assign n6267 = ~n2935 & n6266 ;
  assign n6268 = n2935 & ~n6266 ;
  assign n6269 = ~n6267 & ~n6268 ;
  assign n6270 = ~n6182 & ~n6183 ;
  assign n6271 = ~n6200 & n6270 ;
  assign n6272 = n6200 & ~n6270 ;
  assign n6273 = ~n6271 & ~n6272 ;
  assign n6274 = ~n6269 & ~n6273 ;
  assign n6275 = n6269 & n6273 ;
  assign n6276 = ~n2920 & ~n2922 ;
  assign n6277 = ~n2923 & ~n6276 ;
  assign n6278 = ~n6185 & ~n6187 ;
  assign n6279 = ~n6188 & ~n6278 ;
  assign n6280 = n6277 & n6279 ;
  assign n6281 = ~n6193 & ~n6194 ;
  assign n6282 = ~n6198 & n6281 ;
  assign n6283 = n6198 & ~n6281 ;
  assign n6284 = ~n6282 & ~n6283 ;
  assign n6285 = n6280 & ~n6284 ;
  assign n6286 = ~n6280 & n6284 ;
  assign n6287 = ~n2928 & ~n2929 ;
  assign n6288 = ~n2933 & n6287 ;
  assign n6289 = n2933 & ~n6287 ;
  assign n6290 = ~n6288 & ~n6289 ;
  assign n6291 = ~n6286 & n6290 ;
  assign n6292 = ~n6285 & ~n6291 ;
  assign n6293 = ~n6275 & n6292 ;
  assign n6294 = ~n6274 & ~n6293 ;
  assign n6295 = ~n6265 & n6294 ;
  assign n6296 = ~n6264 & ~n6295 ;
  assign n6297 = ~n6255 & n6296 ;
  assign n6298 = ~n6254 & ~n6297 ;
  assign n6299 = ~n6245 & ~n6298 ;
  assign n6300 = ~n6244 & ~n6299 ;
  assign n6301 = ~n6235 & ~n6300 ;
  assign n6302 = ~n6234 & ~n6301 ;
  assign n6303 = ~n6225 & ~n6302 ;
  assign n6304 = ~n6224 & ~n6303 ;
  assign n6305 = n6215 & ~n6304 ;
  assign n6306 = ~n6215 & n6304 ;
  assign n6307 = ~n6305 & ~n6306 ;
  assign n6308 = \A[835]  & \A[836]  ;
  assign n6309 = ~\A[835]  & ~\A[836]  ;
  assign n6310 = ~n6308 & ~n6309 ;
  assign n6311 = \A[837]  & n6310 ;
  assign n6312 = ~\A[837]  & ~n6310 ;
  assign n6313 = ~n6311 & ~n6312 ;
  assign n6314 = \A[838]  & \A[839]  ;
  assign n6315 = ~\A[838]  & ~\A[839]  ;
  assign n6316 = ~n6314 & ~n6315 ;
  assign n6317 = \A[840]  & n6316 ;
  assign n6318 = ~\A[840]  & ~n6316 ;
  assign n6319 = ~n6317 & ~n6318 ;
  assign n6320 = n6313 & n6319 ;
  assign n6321 = ~n6313 & ~n6319 ;
  assign n6322 = ~n6320 & ~n6321 ;
  assign n6323 = \A[841]  & \A[842]  ;
  assign n6324 = ~\A[841]  & ~\A[842]  ;
  assign n6325 = ~n6323 & ~n6324 ;
  assign n6326 = \A[843]  & n6325 ;
  assign n6327 = ~\A[843]  & ~n6325 ;
  assign n6328 = ~n6326 & ~n6327 ;
  assign n6329 = \A[844]  & \A[845]  ;
  assign n6330 = ~\A[844]  & ~\A[845]  ;
  assign n6331 = ~n6329 & ~n6330 ;
  assign n6332 = \A[846]  & n6331 ;
  assign n6333 = ~\A[846]  & ~n6331 ;
  assign n6334 = ~n6332 & ~n6333 ;
  assign n6335 = n6328 & n6334 ;
  assign n6336 = ~n6328 & ~n6334 ;
  assign n6337 = ~n6335 & ~n6336 ;
  assign n6338 = n6322 & n6337 ;
  assign n6339 = ~n6329 & ~n6332 ;
  assign n6340 = ~n6323 & ~n6326 ;
  assign n6341 = n6339 & n6340 ;
  assign n6342 = ~n6339 & ~n6340 ;
  assign n6343 = ~n6341 & ~n6342 ;
  assign n6344 = n6338 & n6343 ;
  assign n6345 = ~n6308 & ~n6311 ;
  assign n6346 = n6314 & n6320 ;
  assign n6347 = ~n6314 & ~n6317 ;
  assign n6348 = ~n6320 & n6347 ;
  assign n6349 = ~n6346 & ~n6348 ;
  assign n6350 = n6345 & ~n6349 ;
  assign n6351 = ~n6345 & n6349 ;
  assign n6352 = ~n6350 & ~n6351 ;
  assign n6353 = ~n6344 & ~n6352 ;
  assign n6355 = n6335 & ~n6343 ;
  assign n6354 = ~n6335 & n6343 ;
  assign n6356 = ~n6338 & ~n6354 ;
  assign n6357 = ~n6355 & n6356 ;
  assign n6358 = ~n6353 & ~n6357 ;
  assign n6359 = n6335 & ~n6341 ;
  assign n6360 = ~n6342 & ~n6359 ;
  assign n6361 = n6358 & ~n6360 ;
  assign n6362 = ~n6358 & n6360 ;
  assign n6363 = ~n6345 & ~n6348 ;
  assign n6364 = ~n6346 & ~n6363 ;
  assign n6365 = ~n6362 & ~n6364 ;
  assign n6366 = ~n6361 & ~n6365 ;
  assign n6367 = \A[823]  & \A[824]  ;
  assign n6368 = ~\A[823]  & ~\A[824]  ;
  assign n6369 = ~n6367 & ~n6368 ;
  assign n6370 = \A[825]  & n6369 ;
  assign n6371 = ~\A[825]  & ~n6369 ;
  assign n6372 = ~n6370 & ~n6371 ;
  assign n6373 = \A[826]  & \A[827]  ;
  assign n6374 = ~\A[826]  & ~\A[827]  ;
  assign n6375 = ~n6373 & ~n6374 ;
  assign n6376 = \A[828]  & n6375 ;
  assign n6377 = ~\A[828]  & ~n6375 ;
  assign n6378 = ~n6376 & ~n6377 ;
  assign n6379 = n6372 & n6378 ;
  assign n6380 = ~n6372 & ~n6378 ;
  assign n6381 = ~n6379 & ~n6380 ;
  assign n6382 = \A[829]  & \A[830]  ;
  assign n6383 = ~\A[829]  & ~\A[830]  ;
  assign n6384 = ~n6382 & ~n6383 ;
  assign n6385 = \A[831]  & n6384 ;
  assign n6386 = ~\A[831]  & ~n6384 ;
  assign n6387 = ~n6385 & ~n6386 ;
  assign n6388 = \A[832]  & \A[833]  ;
  assign n6389 = ~\A[832]  & ~\A[833]  ;
  assign n6390 = ~n6388 & ~n6389 ;
  assign n6391 = \A[834]  & n6390 ;
  assign n6392 = ~\A[834]  & ~n6390 ;
  assign n6393 = ~n6391 & ~n6392 ;
  assign n6394 = n6387 & n6393 ;
  assign n6395 = ~n6387 & ~n6393 ;
  assign n6396 = ~n6394 & ~n6395 ;
  assign n6397 = n6381 & n6396 ;
  assign n6398 = ~n6388 & ~n6391 ;
  assign n6399 = ~n6382 & ~n6385 ;
  assign n6400 = n6398 & n6399 ;
  assign n6401 = ~n6398 & ~n6399 ;
  assign n6402 = ~n6400 & ~n6401 ;
  assign n6403 = n6397 & n6402 ;
  assign n6404 = ~n6367 & ~n6370 ;
  assign n6405 = n6373 & n6379 ;
  assign n6406 = ~n6373 & ~n6376 ;
  assign n6407 = ~n6379 & n6406 ;
  assign n6408 = ~n6405 & ~n6407 ;
  assign n6409 = n6404 & ~n6408 ;
  assign n6410 = ~n6404 & n6408 ;
  assign n6411 = ~n6409 & ~n6410 ;
  assign n6412 = ~n6403 & ~n6411 ;
  assign n6414 = n6394 & ~n6402 ;
  assign n6413 = ~n6394 & n6402 ;
  assign n6415 = ~n6397 & ~n6413 ;
  assign n6416 = ~n6414 & n6415 ;
  assign n6417 = ~n6412 & ~n6416 ;
  assign n6418 = n6394 & ~n6400 ;
  assign n6419 = ~n6401 & ~n6418 ;
  assign n6420 = n6417 & ~n6419 ;
  assign n6421 = ~n6417 & n6419 ;
  assign n6422 = ~n6404 & ~n6407 ;
  assign n6423 = ~n6405 & ~n6422 ;
  assign n6424 = ~n6421 & ~n6423 ;
  assign n6425 = ~n6420 & ~n6424 ;
  assign n6426 = ~n6366 & ~n6425 ;
  assign n6427 = n6366 & n6425 ;
  assign n6428 = ~n6426 & ~n6427 ;
  assign n6429 = ~n6420 & ~n6421 ;
  assign n6430 = ~n6423 & n6429 ;
  assign n6431 = n6423 & ~n6429 ;
  assign n6432 = ~n6430 & ~n6431 ;
  assign n6433 = ~n6361 & ~n6362 ;
  assign n6434 = ~n6364 & n6433 ;
  assign n6435 = n6364 & ~n6433 ;
  assign n6436 = ~n6434 & ~n6435 ;
  assign n6437 = ~n6432 & ~n6436 ;
  assign n6438 = n6432 & n6436 ;
  assign n6439 = ~n6322 & ~n6337 ;
  assign n6440 = ~n6338 & ~n6439 ;
  assign n6441 = ~n6381 & ~n6396 ;
  assign n6442 = ~n6397 & ~n6441 ;
  assign n6443 = n6440 & n6442 ;
  assign n6444 = ~n6344 & ~n6357 ;
  assign n6445 = ~n6352 & n6444 ;
  assign n6446 = n6352 & ~n6444 ;
  assign n6447 = ~n6445 & ~n6446 ;
  assign n6448 = n6443 & ~n6447 ;
  assign n6449 = ~n6443 & n6447 ;
  assign n6450 = ~n6403 & ~n6416 ;
  assign n6451 = ~n6411 & n6450 ;
  assign n6452 = n6411 & ~n6450 ;
  assign n6453 = ~n6451 & ~n6452 ;
  assign n6454 = ~n6449 & ~n6453 ;
  assign n6455 = ~n6448 & ~n6454 ;
  assign n6456 = ~n6438 & n6455 ;
  assign n6457 = ~n6437 & ~n6456 ;
  assign n6458 = n6428 & ~n6457 ;
  assign n6459 = ~n6428 & n6457 ;
  assign n6460 = ~n6458 & ~n6459 ;
  assign n6461 = \A[811]  & \A[812]  ;
  assign n6462 = ~\A[811]  & ~\A[812]  ;
  assign n6463 = ~n6461 & ~n6462 ;
  assign n6464 = \A[813]  & n6463 ;
  assign n6465 = ~\A[813]  & ~n6463 ;
  assign n6466 = ~n6464 & ~n6465 ;
  assign n6467 = \A[814]  & \A[815]  ;
  assign n6468 = ~\A[814]  & ~\A[815]  ;
  assign n6469 = ~n6467 & ~n6468 ;
  assign n6470 = \A[816]  & n6469 ;
  assign n6471 = ~\A[816]  & ~n6469 ;
  assign n6472 = ~n6470 & ~n6471 ;
  assign n6473 = n6466 & n6472 ;
  assign n6474 = ~n6466 & ~n6472 ;
  assign n6475 = ~n6473 & ~n6474 ;
  assign n6476 = \A[817]  & \A[818]  ;
  assign n6477 = ~\A[817]  & ~\A[818]  ;
  assign n6478 = ~n6476 & ~n6477 ;
  assign n6479 = \A[819]  & n6478 ;
  assign n6480 = ~\A[819]  & ~n6478 ;
  assign n6481 = ~n6479 & ~n6480 ;
  assign n6482 = \A[820]  & \A[821]  ;
  assign n6483 = ~\A[820]  & ~\A[821]  ;
  assign n6484 = ~n6482 & ~n6483 ;
  assign n6485 = \A[822]  & n6484 ;
  assign n6486 = ~\A[822]  & ~n6484 ;
  assign n6487 = ~n6485 & ~n6486 ;
  assign n6488 = n6481 & n6487 ;
  assign n6489 = ~n6481 & ~n6487 ;
  assign n6490 = ~n6488 & ~n6489 ;
  assign n6491 = n6475 & n6490 ;
  assign n6492 = ~n6482 & ~n6485 ;
  assign n6493 = ~n6476 & ~n6479 ;
  assign n6494 = n6492 & n6493 ;
  assign n6495 = ~n6492 & ~n6493 ;
  assign n6496 = ~n6494 & ~n6495 ;
  assign n6497 = n6491 & n6496 ;
  assign n6498 = ~n6461 & ~n6464 ;
  assign n6499 = n6467 & n6473 ;
  assign n6500 = ~n6467 & ~n6470 ;
  assign n6501 = ~n6473 & n6500 ;
  assign n6502 = ~n6499 & ~n6501 ;
  assign n6503 = n6498 & ~n6502 ;
  assign n6504 = ~n6498 & n6502 ;
  assign n6505 = ~n6503 & ~n6504 ;
  assign n6506 = ~n6497 & ~n6505 ;
  assign n6508 = n6488 & ~n6496 ;
  assign n6507 = ~n6488 & n6496 ;
  assign n6509 = ~n6491 & ~n6507 ;
  assign n6510 = ~n6508 & n6509 ;
  assign n6511 = ~n6506 & ~n6510 ;
  assign n6512 = n6488 & ~n6494 ;
  assign n6513 = ~n6495 & ~n6512 ;
  assign n6514 = n6511 & ~n6513 ;
  assign n6515 = ~n6511 & n6513 ;
  assign n6516 = ~n6498 & ~n6501 ;
  assign n6517 = ~n6499 & ~n6516 ;
  assign n6518 = ~n6515 & ~n6517 ;
  assign n6519 = ~n6514 & ~n6518 ;
  assign n6520 = \A[805]  & \A[806]  ;
  assign n6521 = ~\A[805]  & ~\A[806]  ;
  assign n6522 = ~n6520 & ~n6521 ;
  assign n6523 = \A[807]  & n6522 ;
  assign n6524 = ~\A[807]  & ~n6522 ;
  assign n6525 = ~n6523 & ~n6524 ;
  assign n6526 = \A[808]  & \A[809]  ;
  assign n6527 = ~\A[808]  & ~\A[809]  ;
  assign n6528 = ~n6526 & ~n6527 ;
  assign n6529 = \A[810]  & n6528 ;
  assign n6530 = ~\A[810]  & ~n6528 ;
  assign n6531 = ~n6529 & ~n6530 ;
  assign n6532 = n6525 & n6531 ;
  assign n6533 = ~n6525 & ~n6531 ;
  assign n6534 = ~n6532 & ~n6533 ;
  assign n6535 = \A[799]  & \A[800]  ;
  assign n6536 = ~\A[799]  & ~\A[800]  ;
  assign n6537 = ~n6535 & ~n6536 ;
  assign n6538 = \A[801]  & n6537 ;
  assign n6539 = ~\A[801]  & ~n6537 ;
  assign n6540 = ~n6538 & ~n6539 ;
  assign n6541 = \A[802]  & \A[803]  ;
  assign n6542 = ~\A[802]  & ~\A[803]  ;
  assign n6543 = ~n6541 & ~n6542 ;
  assign n6544 = \A[804]  & n6543 ;
  assign n6545 = ~\A[804]  & ~n6543 ;
  assign n6546 = ~n6544 & ~n6545 ;
  assign n6547 = n6540 & n6546 ;
  assign n6548 = ~n6540 & ~n6546 ;
  assign n6549 = ~n6547 & ~n6548 ;
  assign n6550 = n6534 & n6549 ;
  assign n6551 = ~n6526 & ~n6529 ;
  assign n6552 = ~n6520 & ~n6523 ;
  assign n6553 = ~n6551 & ~n6552 ;
  assign n6554 = n6551 & n6552 ;
  assign n6555 = ~n6553 & ~n6554 ;
  assign n6556 = n6550 & n6555 ;
  assign n6557 = ~n6541 & ~n6544 ;
  assign n6558 = ~n6535 & ~n6538 ;
  assign n6559 = ~n6557 & ~n6558 ;
  assign n6560 = n6557 & n6558 ;
  assign n6561 = ~n6559 & ~n6560 ;
  assign n6562 = n6547 & ~n6561 ;
  assign n6563 = ~n6547 & n6561 ;
  assign n6564 = ~n6562 & ~n6563 ;
  assign n6565 = ~n6556 & n6564 ;
  assign n6567 = n6532 & ~n6555 ;
  assign n6566 = ~n6532 & n6555 ;
  assign n6568 = ~n6550 & ~n6566 ;
  assign n6569 = ~n6567 & n6568 ;
  assign n6570 = ~n6565 & ~n6569 ;
  assign n6571 = ~n6532 & ~n6553 ;
  assign n6572 = ~n6554 & ~n6571 ;
  assign n6573 = ~n6570 & ~n6572 ;
  assign n6574 = n6570 & n6572 ;
  assign n6575 = ~n6547 & ~n6559 ;
  assign n6576 = ~n6560 & ~n6575 ;
  assign n6577 = ~n6574 & ~n6576 ;
  assign n6578 = ~n6573 & ~n6577 ;
  assign n6579 = ~n6519 & n6578 ;
  assign n6580 = n6519 & ~n6578 ;
  assign n6581 = ~n6579 & ~n6580 ;
  assign n6582 = ~n6573 & ~n6574 ;
  assign n6583 = ~n6576 & n6582 ;
  assign n6584 = n6576 & ~n6582 ;
  assign n6585 = ~n6583 & ~n6584 ;
  assign n6586 = ~n6514 & ~n6515 ;
  assign n6587 = ~n6517 & n6586 ;
  assign n6588 = n6517 & ~n6586 ;
  assign n6589 = ~n6587 & ~n6588 ;
  assign n6590 = ~n6585 & n6589 ;
  assign n6591 = n6585 & ~n6589 ;
  assign n6592 = ~n6475 & ~n6490 ;
  assign n6593 = ~n6491 & ~n6592 ;
  assign n6594 = ~n6534 & ~n6549 ;
  assign n6595 = ~n6550 & ~n6594 ;
  assign n6596 = n6593 & n6595 ;
  assign n6597 = ~n6497 & ~n6510 ;
  assign n6598 = ~n6505 & n6597 ;
  assign n6599 = n6505 & ~n6597 ;
  assign n6600 = ~n6598 & ~n6599 ;
  assign n6601 = n6596 & ~n6600 ;
  assign n6602 = ~n6596 & n6600 ;
  assign n6603 = ~n6556 & ~n6569 ;
  assign n6604 = n6564 & n6603 ;
  assign n6605 = ~n6564 & ~n6603 ;
  assign n6606 = ~n6604 & ~n6605 ;
  assign n6607 = ~n6602 & ~n6606 ;
  assign n6608 = ~n6601 & ~n6607 ;
  assign n6609 = ~n6591 & ~n6608 ;
  assign n6610 = ~n6590 & ~n6609 ;
  assign n6611 = n6581 & ~n6610 ;
  assign n6612 = ~n6581 & n6610 ;
  assign n6613 = ~n6611 & ~n6612 ;
  assign n6614 = n6460 & ~n6613 ;
  assign n6615 = ~n6460 & n6613 ;
  assign n6616 = ~n6590 & ~n6591 ;
  assign n6617 = ~n6608 & n6616 ;
  assign n6618 = n6608 & ~n6616 ;
  assign n6619 = ~n6617 & ~n6618 ;
  assign n6620 = ~n6437 & ~n6438 ;
  assign n6621 = ~n6455 & n6620 ;
  assign n6622 = n6455 & ~n6620 ;
  assign n6623 = ~n6621 & ~n6622 ;
  assign n6624 = ~n6619 & ~n6623 ;
  assign n6625 = n6619 & n6623 ;
  assign n6626 = ~n6440 & ~n6442 ;
  assign n6627 = ~n6443 & ~n6626 ;
  assign n6628 = ~n6593 & ~n6595 ;
  assign n6629 = ~n6596 & ~n6628 ;
  assign n6630 = n6627 & n6629 ;
  assign n6631 = ~n6448 & ~n6449 ;
  assign n6632 = ~n6453 & n6631 ;
  assign n6633 = n6453 & ~n6631 ;
  assign n6634 = ~n6632 & ~n6633 ;
  assign n6635 = n6630 & n6634 ;
  assign n6636 = ~n6630 & ~n6634 ;
  assign n6637 = ~n6601 & ~n6602 ;
  assign n6638 = ~n6606 & n6637 ;
  assign n6639 = n6606 & ~n6637 ;
  assign n6640 = ~n6638 & ~n6639 ;
  assign n6641 = ~n6636 & n6640 ;
  assign n6642 = ~n6635 & ~n6641 ;
  assign n6643 = ~n6625 & n6642 ;
  assign n6644 = ~n6624 & ~n6643 ;
  assign n6645 = ~n6615 & ~n6644 ;
  assign n6646 = ~n6614 & ~n6645 ;
  assign n6647 = ~n6427 & n6457 ;
  assign n6648 = ~n6426 & ~n6647 ;
  assign n6649 = n6646 & ~n6648 ;
  assign n6650 = ~n6646 & n6648 ;
  assign n6651 = ~n6580 & ~n6610 ;
  assign n6652 = ~n6579 & ~n6651 ;
  assign n6653 = ~n6650 & ~n6652 ;
  assign n6654 = ~n6649 & ~n6653 ;
  assign n6655 = \A[787]  & \A[788]  ;
  assign n6656 = ~\A[787]  & ~\A[788]  ;
  assign n6657 = ~n6655 & ~n6656 ;
  assign n6658 = \A[789]  & n6657 ;
  assign n6659 = ~\A[789]  & ~n6657 ;
  assign n6660 = ~n6658 & ~n6659 ;
  assign n6661 = \A[790]  & \A[791]  ;
  assign n6662 = ~\A[790]  & ~\A[791]  ;
  assign n6663 = ~n6661 & ~n6662 ;
  assign n6664 = \A[792]  & n6663 ;
  assign n6665 = ~\A[792]  & ~n6663 ;
  assign n6666 = ~n6664 & ~n6665 ;
  assign n6667 = n6660 & n6666 ;
  assign n6668 = ~n6660 & ~n6666 ;
  assign n6669 = ~n6667 & ~n6668 ;
  assign n6670 = \A[793]  & \A[794]  ;
  assign n6671 = ~\A[793]  & ~\A[794]  ;
  assign n6672 = ~n6670 & ~n6671 ;
  assign n6673 = \A[795]  & n6672 ;
  assign n6674 = ~\A[795]  & ~n6672 ;
  assign n6675 = ~n6673 & ~n6674 ;
  assign n6676 = \A[796]  & \A[797]  ;
  assign n6677 = ~\A[796]  & ~\A[797]  ;
  assign n6678 = ~n6676 & ~n6677 ;
  assign n6679 = \A[798]  & n6678 ;
  assign n6680 = ~\A[798]  & ~n6678 ;
  assign n6681 = ~n6679 & ~n6680 ;
  assign n6682 = n6675 & n6681 ;
  assign n6683 = ~n6675 & ~n6681 ;
  assign n6684 = ~n6682 & ~n6683 ;
  assign n6685 = n6669 & n6684 ;
  assign n6686 = ~n6676 & ~n6679 ;
  assign n6687 = ~n6670 & ~n6673 ;
  assign n6688 = n6686 & n6687 ;
  assign n6689 = ~n6686 & ~n6687 ;
  assign n6690 = ~n6688 & ~n6689 ;
  assign n6691 = n6685 & n6690 ;
  assign n6692 = ~n6655 & ~n6658 ;
  assign n6693 = n6661 & n6667 ;
  assign n6694 = ~n6661 & ~n6664 ;
  assign n6695 = ~n6667 & n6694 ;
  assign n6696 = ~n6693 & ~n6695 ;
  assign n6697 = n6692 & ~n6696 ;
  assign n6698 = ~n6692 & n6696 ;
  assign n6699 = ~n6697 & ~n6698 ;
  assign n6700 = ~n6691 & ~n6699 ;
  assign n6702 = n6682 & ~n6690 ;
  assign n6701 = ~n6682 & n6690 ;
  assign n6703 = ~n6685 & ~n6701 ;
  assign n6704 = ~n6702 & n6703 ;
  assign n6705 = ~n6700 & ~n6704 ;
  assign n6706 = n6682 & ~n6688 ;
  assign n6707 = ~n6689 & ~n6706 ;
  assign n6708 = n6705 & ~n6707 ;
  assign n6709 = ~n6705 & n6707 ;
  assign n6710 = ~n6692 & ~n6695 ;
  assign n6711 = ~n6693 & ~n6710 ;
  assign n6712 = ~n6709 & ~n6711 ;
  assign n6713 = ~n6708 & ~n6712 ;
  assign n6714 = \A[775]  & \A[776]  ;
  assign n6715 = ~\A[775]  & ~\A[776]  ;
  assign n6716 = ~n6714 & ~n6715 ;
  assign n6717 = \A[777]  & n6716 ;
  assign n6718 = ~\A[777]  & ~n6716 ;
  assign n6719 = ~n6717 & ~n6718 ;
  assign n6720 = \A[778]  & \A[779]  ;
  assign n6721 = ~\A[778]  & ~\A[779]  ;
  assign n6722 = ~n6720 & ~n6721 ;
  assign n6723 = \A[780]  & n6722 ;
  assign n6724 = ~\A[780]  & ~n6722 ;
  assign n6725 = ~n6723 & ~n6724 ;
  assign n6726 = n6719 & n6725 ;
  assign n6727 = ~n6719 & ~n6725 ;
  assign n6728 = ~n6726 & ~n6727 ;
  assign n6729 = \A[781]  & \A[782]  ;
  assign n6730 = ~\A[781]  & ~\A[782]  ;
  assign n6731 = ~n6729 & ~n6730 ;
  assign n6732 = \A[783]  & n6731 ;
  assign n6733 = ~\A[783]  & ~n6731 ;
  assign n6734 = ~n6732 & ~n6733 ;
  assign n6735 = \A[784]  & \A[785]  ;
  assign n6736 = ~\A[784]  & ~\A[785]  ;
  assign n6737 = ~n6735 & ~n6736 ;
  assign n6738 = \A[786]  & n6737 ;
  assign n6739 = ~\A[786]  & ~n6737 ;
  assign n6740 = ~n6738 & ~n6739 ;
  assign n6741 = n6734 & n6740 ;
  assign n6742 = ~n6734 & ~n6740 ;
  assign n6743 = ~n6741 & ~n6742 ;
  assign n6744 = n6728 & n6743 ;
  assign n6745 = ~n6735 & ~n6738 ;
  assign n6746 = ~n6729 & ~n6732 ;
  assign n6747 = n6745 & n6746 ;
  assign n6748 = ~n6745 & ~n6746 ;
  assign n6749 = ~n6747 & ~n6748 ;
  assign n6750 = n6744 & n6749 ;
  assign n6751 = ~n6714 & ~n6717 ;
  assign n6752 = n6720 & n6726 ;
  assign n6753 = ~n6720 & ~n6723 ;
  assign n6754 = ~n6726 & n6753 ;
  assign n6755 = ~n6752 & ~n6754 ;
  assign n6756 = n6751 & ~n6755 ;
  assign n6757 = ~n6751 & n6755 ;
  assign n6758 = ~n6756 & ~n6757 ;
  assign n6759 = ~n6750 & ~n6758 ;
  assign n6761 = n6741 & ~n6749 ;
  assign n6760 = ~n6741 & n6749 ;
  assign n6762 = ~n6744 & ~n6760 ;
  assign n6763 = ~n6761 & n6762 ;
  assign n6764 = ~n6759 & ~n6763 ;
  assign n6765 = n6741 & ~n6747 ;
  assign n6766 = ~n6748 & ~n6765 ;
  assign n6767 = n6764 & ~n6766 ;
  assign n6768 = ~n6764 & n6766 ;
  assign n6769 = ~n6751 & ~n6754 ;
  assign n6770 = ~n6752 & ~n6769 ;
  assign n6771 = ~n6768 & ~n6770 ;
  assign n6772 = ~n6767 & ~n6771 ;
  assign n6773 = ~n6713 & ~n6772 ;
  assign n6774 = n6713 & n6772 ;
  assign n6775 = ~n6767 & ~n6768 ;
  assign n6776 = ~n6770 & n6775 ;
  assign n6777 = n6770 & ~n6775 ;
  assign n6778 = ~n6776 & ~n6777 ;
  assign n6779 = ~n6708 & ~n6709 ;
  assign n6780 = ~n6711 & n6779 ;
  assign n6781 = n6711 & ~n6779 ;
  assign n6782 = ~n6780 & ~n6781 ;
  assign n6783 = ~n6778 & ~n6782 ;
  assign n6784 = n6778 & n6782 ;
  assign n6785 = ~n6669 & ~n6684 ;
  assign n6786 = ~n6685 & ~n6785 ;
  assign n6787 = ~n6728 & ~n6743 ;
  assign n6788 = ~n6744 & ~n6787 ;
  assign n6789 = n6786 & n6788 ;
  assign n6790 = ~n6691 & ~n6704 ;
  assign n6791 = ~n6699 & n6790 ;
  assign n6792 = n6699 & ~n6790 ;
  assign n6793 = ~n6791 & ~n6792 ;
  assign n6794 = n6789 & ~n6793 ;
  assign n6795 = ~n6789 & n6793 ;
  assign n6796 = ~n6750 & ~n6763 ;
  assign n6797 = ~n6758 & n6796 ;
  assign n6798 = n6758 & ~n6796 ;
  assign n6799 = ~n6797 & ~n6798 ;
  assign n6800 = ~n6795 & ~n6799 ;
  assign n6801 = ~n6794 & ~n6800 ;
  assign n6802 = ~n6784 & n6801 ;
  assign n6803 = ~n6783 & ~n6802 ;
  assign n6804 = ~n6774 & n6803 ;
  assign n6805 = ~n6773 & ~n6804 ;
  assign n6806 = \A[757]  & \A[758]  ;
  assign n6807 = ~\A[757]  & ~\A[758]  ;
  assign n6808 = ~n6806 & ~n6807 ;
  assign n6809 = \A[759]  & n6808 ;
  assign n6810 = ~\A[759]  & ~n6808 ;
  assign n6811 = ~n6809 & ~n6810 ;
  assign n6812 = \A[760]  & \A[761]  ;
  assign n6813 = ~\A[760]  & ~\A[761]  ;
  assign n6814 = ~n6812 & ~n6813 ;
  assign n6815 = \A[762]  & n6814 ;
  assign n6816 = ~\A[762]  & ~n6814 ;
  assign n6817 = ~n6815 & ~n6816 ;
  assign n6818 = n6811 & n6817 ;
  assign n6819 = ~n6811 & ~n6817 ;
  assign n6820 = ~n6818 & ~n6819 ;
  assign n6821 = \A[751]  & \A[752]  ;
  assign n6822 = ~\A[751]  & ~\A[752]  ;
  assign n6823 = ~n6821 & ~n6822 ;
  assign n6824 = \A[753]  & n6823 ;
  assign n6825 = ~\A[753]  & ~n6823 ;
  assign n6826 = ~n6824 & ~n6825 ;
  assign n6827 = \A[754]  & \A[755]  ;
  assign n6828 = ~\A[754]  & ~\A[755]  ;
  assign n6829 = ~n6827 & ~n6828 ;
  assign n6830 = \A[756]  & n6829 ;
  assign n6831 = ~\A[756]  & ~n6829 ;
  assign n6832 = ~n6830 & ~n6831 ;
  assign n6833 = n6826 & n6832 ;
  assign n6834 = ~n6826 & ~n6832 ;
  assign n6835 = ~n6833 & ~n6834 ;
  assign n6836 = n6820 & n6835 ;
  assign n6837 = ~n6812 & ~n6815 ;
  assign n6838 = ~n6806 & ~n6809 ;
  assign n6839 = n6837 & n6838 ;
  assign n6840 = ~n6837 & ~n6838 ;
  assign n6841 = ~n6839 & ~n6840 ;
  assign n6842 = n6836 & n6841 ;
  assign n6843 = ~n6827 & ~n6830 ;
  assign n6844 = ~n6821 & ~n6824 ;
  assign n6845 = ~n6843 & ~n6844 ;
  assign n6846 = n6843 & n6844 ;
  assign n6847 = ~n6845 & ~n6846 ;
  assign n6848 = n6833 & ~n6847 ;
  assign n6849 = ~n6833 & n6847 ;
  assign n6850 = ~n6848 & ~n6849 ;
  assign n6851 = ~n6842 & n6850 ;
  assign n6853 = n6818 & ~n6841 ;
  assign n6852 = ~n6818 & n6841 ;
  assign n6854 = ~n6836 & ~n6852 ;
  assign n6855 = ~n6853 & n6854 ;
  assign n6856 = ~n6851 & ~n6855 ;
  assign n6857 = ~n6833 & ~n6845 ;
  assign n6858 = ~n6846 & ~n6857 ;
  assign n6859 = n6856 & n6858 ;
  assign n6860 = ~n6856 & ~n6858 ;
  assign n6861 = ~n6859 & ~n6860 ;
  assign n6862 = ~n6818 & ~n6840 ;
  assign n6863 = ~n6839 & ~n6862 ;
  assign n6864 = n6861 & ~n6863 ;
  assign n6865 = ~n6861 & n6863 ;
  assign n6866 = ~n6864 & ~n6865 ;
  assign n6867 = \A[766]  & \A[767]  ;
  assign n6868 = \A[763]  & \A[764]  ;
  assign n6869 = ~\A[763]  & ~\A[764]  ;
  assign n6870 = ~n6868 & ~n6869 ;
  assign n6871 = \A[765]  & n6870 ;
  assign n6872 = ~\A[765]  & ~n6870 ;
  assign n6873 = ~n6871 & ~n6872 ;
  assign n6874 = ~\A[766]  & ~\A[767]  ;
  assign n6875 = ~n6867 & ~n6874 ;
  assign n6876 = \A[768]  & n6875 ;
  assign n6877 = ~\A[768]  & ~n6875 ;
  assign n6878 = ~n6876 & ~n6877 ;
  assign n6879 = n6873 & n6878 ;
  assign n6880 = n6867 & n6879 ;
  assign n6881 = ~n6868 & ~n6871 ;
  assign n6882 = ~n6867 & ~n6876 ;
  assign n6883 = ~n6879 & n6882 ;
  assign n6884 = ~n6881 & ~n6883 ;
  assign n6885 = ~n6880 & ~n6884 ;
  assign n6886 = \A[772]  & \A[773]  ;
  assign n6887 = ~\A[772]  & ~\A[773]  ;
  assign n6888 = ~n6886 & ~n6887 ;
  assign n6889 = \A[774]  & n6888 ;
  assign n6890 = ~n6886 & ~n6889 ;
  assign n6891 = \A[769]  & \A[770]  ;
  assign n6892 = ~\A[769]  & ~\A[770]  ;
  assign n6893 = ~n6891 & ~n6892 ;
  assign n6894 = \A[771]  & n6893 ;
  assign n6895 = ~n6891 & ~n6894 ;
  assign n6896 = n6890 & n6895 ;
  assign n6897 = ~n6890 & ~n6895 ;
  assign n6898 = ~\A[771]  & ~n6893 ;
  assign n6899 = ~n6894 & ~n6898 ;
  assign n6900 = ~\A[774]  & ~n6888 ;
  assign n6901 = ~n6889 & ~n6900 ;
  assign n6902 = n6899 & n6901 ;
  assign n6903 = ~n6897 & ~n6902 ;
  assign n6904 = ~n6896 & ~n6903 ;
  assign n6905 = ~n6899 & ~n6901 ;
  assign n6906 = ~n6902 & ~n6905 ;
  assign n6907 = ~n6873 & ~n6878 ;
  assign n6908 = ~n6879 & ~n6907 ;
  assign n6909 = n6906 & n6908 ;
  assign n6910 = n6880 & ~n6881 ;
  assign n6911 = n6909 & ~n6910 ;
  assign n6912 = ~n6896 & ~n6897 ;
  assign n6913 = n6902 & ~n6912 ;
  assign n6914 = ~n6902 & n6912 ;
  assign n6915 = ~n6913 & ~n6914 ;
  assign n6916 = n6911 & ~n6915 ;
  assign n6917 = ~n6911 & n6915 ;
  assign n6918 = ~n6880 & ~n6883 ;
  assign n6919 = n6881 & ~n6918 ;
  assign n6920 = ~n6881 & n6918 ;
  assign n6921 = ~n6919 & ~n6920 ;
  assign n6922 = ~n6917 & n6921 ;
  assign n6923 = ~n6916 & ~n6922 ;
  assign n6924 = n6904 & ~n6923 ;
  assign n6925 = ~n6904 & n6923 ;
  assign n6926 = ~n6924 & ~n6925 ;
  assign n6927 = n6885 & n6926 ;
  assign n6928 = ~n6885 & ~n6926 ;
  assign n6929 = ~n6927 & ~n6928 ;
  assign n6930 = ~n6866 & ~n6929 ;
  assign n6931 = n6866 & n6929 ;
  assign n6932 = ~n6906 & ~n6908 ;
  assign n6933 = ~n6909 & ~n6932 ;
  assign n6934 = ~n6820 & ~n6835 ;
  assign n6935 = ~n6836 & ~n6934 ;
  assign n6936 = n6933 & n6935 ;
  assign n6937 = ~n6916 & ~n6917 ;
  assign n6938 = n6921 & n6937 ;
  assign n6939 = ~n6921 & ~n6937 ;
  assign n6940 = ~n6938 & ~n6939 ;
  assign n6941 = n6936 & n6940 ;
  assign n6942 = ~n6936 & ~n6940 ;
  assign n6943 = ~n6842 & ~n6855 ;
  assign n6944 = n6850 & n6943 ;
  assign n6945 = ~n6850 & ~n6943 ;
  assign n6946 = ~n6944 & ~n6945 ;
  assign n6947 = ~n6942 & ~n6946 ;
  assign n6948 = ~n6941 & ~n6947 ;
  assign n6949 = ~n6931 & ~n6948 ;
  assign n6950 = ~n6930 & ~n6949 ;
  assign n6951 = ~n6885 & ~n6925 ;
  assign n6952 = ~n6924 & ~n6951 ;
  assign n6953 = n6950 & n6952 ;
  assign n6954 = ~n6950 & ~n6952 ;
  assign n6955 = ~n6859 & ~n6863 ;
  assign n6956 = ~n6860 & ~n6955 ;
  assign n6957 = ~n6954 & ~n6956 ;
  assign n6958 = ~n6953 & ~n6957 ;
  assign n6959 = ~n6805 & n6958 ;
  assign n6960 = n6805 & ~n6958 ;
  assign n6961 = ~n6773 & ~n6774 ;
  assign n6962 = ~n6803 & n6961 ;
  assign n6963 = n6803 & ~n6961 ;
  assign n6964 = ~n6962 & ~n6963 ;
  assign n6965 = ~n6953 & ~n6954 ;
  assign n6966 = ~n6956 & n6965 ;
  assign n6967 = n6956 & ~n6965 ;
  assign n6968 = ~n6966 & ~n6967 ;
  assign n6969 = ~n6964 & ~n6968 ;
  assign n6970 = n6964 & n6968 ;
  assign n6971 = ~n6930 & ~n6931 ;
  assign n6972 = ~n6948 & n6971 ;
  assign n6973 = n6948 & ~n6971 ;
  assign n6974 = ~n6972 & ~n6973 ;
  assign n6975 = ~n6783 & ~n6784 ;
  assign n6976 = ~n6801 & n6975 ;
  assign n6977 = n6801 & ~n6975 ;
  assign n6978 = ~n6976 & ~n6977 ;
  assign n6979 = ~n6974 & ~n6978 ;
  assign n6980 = n6974 & n6978 ;
  assign n6981 = ~n6786 & ~n6788 ;
  assign n6982 = ~n6789 & ~n6981 ;
  assign n6983 = ~n6933 & ~n6935 ;
  assign n6984 = ~n6936 & ~n6983 ;
  assign n6985 = n6982 & n6984 ;
  assign n6986 = ~n6794 & ~n6795 ;
  assign n6987 = ~n6799 & n6986 ;
  assign n6988 = n6799 & ~n6986 ;
  assign n6989 = ~n6987 & ~n6988 ;
  assign n6990 = n6985 & n6989 ;
  assign n6991 = ~n6985 & ~n6989 ;
  assign n6992 = ~n6941 & ~n6942 ;
  assign n6993 = ~n6946 & n6992 ;
  assign n6994 = n6946 & ~n6992 ;
  assign n6995 = ~n6993 & ~n6994 ;
  assign n6996 = ~n6991 & n6995 ;
  assign n6997 = ~n6990 & ~n6996 ;
  assign n6998 = ~n6980 & n6997 ;
  assign n6999 = ~n6979 & ~n6998 ;
  assign n7000 = ~n6970 & n6999 ;
  assign n7001 = ~n6969 & ~n7000 ;
  assign n7002 = ~n6960 & ~n7001 ;
  assign n7003 = ~n6959 & ~n7002 ;
  assign n7004 = ~n6654 & ~n7003 ;
  assign n7005 = n6654 & n7003 ;
  assign n7006 = ~n6959 & ~n6960 ;
  assign n7007 = ~n7001 & n7006 ;
  assign n7008 = n7001 & ~n7006 ;
  assign n7009 = ~n7007 & ~n7008 ;
  assign n7010 = ~n6649 & ~n6650 ;
  assign n7011 = n6652 & n7010 ;
  assign n7012 = ~n6652 & ~n7010 ;
  assign n7013 = ~n7011 & ~n7012 ;
  assign n7014 = n7009 & ~n7013 ;
  assign n7015 = ~n7009 & n7013 ;
  assign n7016 = ~n6614 & ~n6615 ;
  assign n7017 = ~n6644 & n7016 ;
  assign n7018 = n6644 & ~n7016 ;
  assign n7019 = ~n7017 & ~n7018 ;
  assign n7020 = ~n6969 & ~n6970 ;
  assign n7021 = n6999 & n7020 ;
  assign n7022 = ~n6999 & ~n7020 ;
  assign n7023 = ~n7021 & ~n7022 ;
  assign n7024 = n7019 & ~n7023 ;
  assign n7025 = ~n7019 & n7023 ;
  assign n7026 = ~n6979 & ~n6980 ;
  assign n7027 = ~n6997 & n7026 ;
  assign n7028 = n6997 & ~n7026 ;
  assign n7029 = ~n7027 & ~n7028 ;
  assign n7030 = ~n6624 & ~n6625 ;
  assign n7031 = ~n6642 & n7030 ;
  assign n7032 = n6642 & ~n7030 ;
  assign n7033 = ~n7031 & ~n7032 ;
  assign n7034 = ~n7029 & ~n7033 ;
  assign n7035 = n7029 & n7033 ;
  assign n7036 = ~n6627 & ~n6629 ;
  assign n7037 = ~n6630 & ~n7036 ;
  assign n7038 = ~n6982 & ~n6984 ;
  assign n7039 = ~n6985 & ~n7038 ;
  assign n7040 = n7037 & n7039 ;
  assign n7041 = ~n6635 & ~n6636 ;
  assign n7042 = ~n6640 & n7041 ;
  assign n7043 = n6640 & ~n7041 ;
  assign n7044 = ~n7042 & ~n7043 ;
  assign n7045 = n7040 & ~n7044 ;
  assign n7046 = ~n7040 & n7044 ;
  assign n7047 = ~n6990 & ~n6991 ;
  assign n7048 = ~n6995 & n7047 ;
  assign n7049 = n6995 & ~n7047 ;
  assign n7050 = ~n7048 & ~n7049 ;
  assign n7051 = ~n7046 & ~n7050 ;
  assign n7052 = ~n7045 & ~n7051 ;
  assign n7053 = ~n7035 & n7052 ;
  assign n7054 = ~n7034 & ~n7053 ;
  assign n7055 = ~n7025 & ~n7054 ;
  assign n7056 = ~n7024 & ~n7055 ;
  assign n7057 = ~n7015 & n7056 ;
  assign n7058 = ~n7014 & ~n7057 ;
  assign n7059 = ~n7005 & ~n7058 ;
  assign n7060 = ~n7004 & ~n7059 ;
  assign n7061 = \A[739]  & \A[740]  ;
  assign n7062 = ~\A[739]  & ~\A[740]  ;
  assign n7063 = ~n7061 & ~n7062 ;
  assign n7064 = \A[741]  & n7063 ;
  assign n7065 = ~\A[741]  & ~n7063 ;
  assign n7066 = ~n7064 & ~n7065 ;
  assign n7067 = \A[742]  & \A[743]  ;
  assign n7068 = ~\A[742]  & ~\A[743]  ;
  assign n7069 = ~n7067 & ~n7068 ;
  assign n7070 = \A[744]  & n7069 ;
  assign n7071 = ~\A[744]  & ~n7069 ;
  assign n7072 = ~n7070 & ~n7071 ;
  assign n7073 = n7066 & n7072 ;
  assign n7074 = ~n7066 & ~n7072 ;
  assign n7075 = ~n7073 & ~n7074 ;
  assign n7076 = \A[745]  & \A[746]  ;
  assign n7077 = ~\A[745]  & ~\A[746]  ;
  assign n7078 = ~n7076 & ~n7077 ;
  assign n7079 = \A[747]  & n7078 ;
  assign n7080 = ~\A[747]  & ~n7078 ;
  assign n7081 = ~n7079 & ~n7080 ;
  assign n7082 = \A[748]  & \A[749]  ;
  assign n7083 = ~\A[748]  & ~\A[749]  ;
  assign n7084 = ~n7082 & ~n7083 ;
  assign n7085 = \A[750]  & n7084 ;
  assign n7086 = ~\A[750]  & ~n7084 ;
  assign n7087 = ~n7085 & ~n7086 ;
  assign n7088 = n7081 & n7087 ;
  assign n7089 = ~n7081 & ~n7087 ;
  assign n7090 = ~n7088 & ~n7089 ;
  assign n7091 = n7075 & n7090 ;
  assign n7092 = ~n7082 & ~n7085 ;
  assign n7093 = ~n7076 & ~n7079 ;
  assign n7094 = n7092 & n7093 ;
  assign n7095 = ~n7092 & ~n7093 ;
  assign n7096 = ~n7094 & ~n7095 ;
  assign n7097 = n7091 & n7096 ;
  assign n7098 = ~n7061 & ~n7064 ;
  assign n7099 = n7067 & n7073 ;
  assign n7100 = ~n7067 & ~n7070 ;
  assign n7101 = ~n7073 & n7100 ;
  assign n7102 = ~n7099 & ~n7101 ;
  assign n7103 = n7098 & ~n7102 ;
  assign n7104 = ~n7098 & n7102 ;
  assign n7105 = ~n7103 & ~n7104 ;
  assign n7106 = ~n7097 & ~n7105 ;
  assign n7108 = n7088 & ~n7096 ;
  assign n7107 = ~n7088 & n7096 ;
  assign n7109 = ~n7091 & ~n7107 ;
  assign n7110 = ~n7108 & n7109 ;
  assign n7111 = ~n7106 & ~n7110 ;
  assign n7112 = n7088 & ~n7094 ;
  assign n7113 = ~n7095 & ~n7112 ;
  assign n7114 = n7111 & ~n7113 ;
  assign n7115 = ~n7111 & n7113 ;
  assign n7116 = ~n7098 & ~n7101 ;
  assign n7117 = ~n7099 & ~n7116 ;
  assign n7118 = ~n7115 & ~n7117 ;
  assign n7119 = ~n7114 & ~n7118 ;
  assign n7120 = \A[727]  & \A[728]  ;
  assign n7121 = ~\A[727]  & ~\A[728]  ;
  assign n7122 = ~n7120 & ~n7121 ;
  assign n7123 = \A[729]  & n7122 ;
  assign n7124 = ~\A[729]  & ~n7122 ;
  assign n7125 = ~n7123 & ~n7124 ;
  assign n7126 = \A[730]  & \A[731]  ;
  assign n7127 = ~\A[730]  & ~\A[731]  ;
  assign n7128 = ~n7126 & ~n7127 ;
  assign n7129 = \A[732]  & n7128 ;
  assign n7130 = ~\A[732]  & ~n7128 ;
  assign n7131 = ~n7129 & ~n7130 ;
  assign n7132 = n7125 & n7131 ;
  assign n7133 = ~n7125 & ~n7131 ;
  assign n7134 = ~n7132 & ~n7133 ;
  assign n7135 = \A[733]  & \A[734]  ;
  assign n7136 = ~\A[733]  & ~\A[734]  ;
  assign n7137 = ~n7135 & ~n7136 ;
  assign n7138 = \A[735]  & n7137 ;
  assign n7139 = ~\A[735]  & ~n7137 ;
  assign n7140 = ~n7138 & ~n7139 ;
  assign n7141 = \A[736]  & \A[737]  ;
  assign n7142 = ~\A[736]  & ~\A[737]  ;
  assign n7143 = ~n7141 & ~n7142 ;
  assign n7144 = \A[738]  & n7143 ;
  assign n7145 = ~\A[738]  & ~n7143 ;
  assign n7146 = ~n7144 & ~n7145 ;
  assign n7147 = n7140 & n7146 ;
  assign n7148 = ~n7140 & ~n7146 ;
  assign n7149 = ~n7147 & ~n7148 ;
  assign n7150 = n7134 & n7149 ;
  assign n7151 = ~n7141 & ~n7144 ;
  assign n7152 = ~n7135 & ~n7138 ;
  assign n7153 = n7151 & n7152 ;
  assign n7154 = ~n7151 & ~n7152 ;
  assign n7155 = ~n7153 & ~n7154 ;
  assign n7156 = n7150 & n7155 ;
  assign n7157 = ~n7120 & ~n7123 ;
  assign n7158 = n7126 & n7132 ;
  assign n7159 = ~n7126 & ~n7129 ;
  assign n7160 = ~n7132 & n7159 ;
  assign n7161 = ~n7158 & ~n7160 ;
  assign n7162 = n7157 & ~n7161 ;
  assign n7163 = ~n7157 & n7161 ;
  assign n7164 = ~n7162 & ~n7163 ;
  assign n7165 = ~n7156 & ~n7164 ;
  assign n7167 = n7147 & ~n7155 ;
  assign n7166 = ~n7147 & n7155 ;
  assign n7168 = ~n7150 & ~n7166 ;
  assign n7169 = ~n7167 & n7168 ;
  assign n7170 = ~n7165 & ~n7169 ;
  assign n7171 = n7147 & ~n7153 ;
  assign n7172 = ~n7154 & ~n7171 ;
  assign n7173 = n7170 & ~n7172 ;
  assign n7174 = ~n7170 & n7172 ;
  assign n7175 = ~n7157 & ~n7160 ;
  assign n7176 = ~n7158 & ~n7175 ;
  assign n7177 = ~n7174 & ~n7176 ;
  assign n7178 = ~n7173 & ~n7177 ;
  assign n7179 = ~n7119 & ~n7178 ;
  assign n7180 = n7119 & n7178 ;
  assign n7181 = ~n7179 & ~n7180 ;
  assign n7182 = ~n7173 & ~n7174 ;
  assign n7183 = ~n7176 & n7182 ;
  assign n7184 = n7176 & ~n7182 ;
  assign n7185 = ~n7183 & ~n7184 ;
  assign n7186 = ~n7114 & ~n7115 ;
  assign n7187 = ~n7117 & n7186 ;
  assign n7188 = n7117 & ~n7186 ;
  assign n7189 = ~n7187 & ~n7188 ;
  assign n7190 = ~n7185 & ~n7189 ;
  assign n7191 = n7185 & n7189 ;
  assign n7192 = ~n7075 & ~n7090 ;
  assign n7193 = ~n7091 & ~n7192 ;
  assign n7194 = ~n7134 & ~n7149 ;
  assign n7195 = ~n7150 & ~n7194 ;
  assign n7196 = n7193 & n7195 ;
  assign n7197 = ~n7097 & ~n7110 ;
  assign n7198 = ~n7105 & n7197 ;
  assign n7199 = n7105 & ~n7197 ;
  assign n7200 = ~n7198 & ~n7199 ;
  assign n7201 = n7196 & ~n7200 ;
  assign n7202 = ~n7196 & n7200 ;
  assign n7203 = ~n7156 & ~n7169 ;
  assign n7204 = ~n7164 & n7203 ;
  assign n7205 = n7164 & ~n7203 ;
  assign n7206 = ~n7204 & ~n7205 ;
  assign n7207 = ~n7202 & ~n7206 ;
  assign n7208 = ~n7201 & ~n7207 ;
  assign n7209 = ~n7191 & n7208 ;
  assign n7210 = ~n7190 & ~n7209 ;
  assign n7211 = n7181 & ~n7210 ;
  assign n7212 = ~n7181 & n7210 ;
  assign n7213 = ~n7211 & ~n7212 ;
  assign n7214 = \A[715]  & \A[716]  ;
  assign n7215 = ~\A[715]  & ~\A[716]  ;
  assign n7216 = ~n7214 & ~n7215 ;
  assign n7217 = \A[717]  & n7216 ;
  assign n7218 = ~\A[717]  & ~n7216 ;
  assign n7219 = ~n7217 & ~n7218 ;
  assign n7220 = \A[718]  & \A[719]  ;
  assign n7221 = ~\A[718]  & ~\A[719]  ;
  assign n7222 = ~n7220 & ~n7221 ;
  assign n7223 = \A[720]  & n7222 ;
  assign n7224 = ~\A[720]  & ~n7222 ;
  assign n7225 = ~n7223 & ~n7224 ;
  assign n7226 = n7219 & n7225 ;
  assign n7227 = ~n7219 & ~n7225 ;
  assign n7228 = ~n7226 & ~n7227 ;
  assign n7229 = \A[721]  & \A[722]  ;
  assign n7230 = ~\A[721]  & ~\A[722]  ;
  assign n7231 = ~n7229 & ~n7230 ;
  assign n7232 = \A[723]  & n7231 ;
  assign n7233 = ~\A[723]  & ~n7231 ;
  assign n7234 = ~n7232 & ~n7233 ;
  assign n7235 = \A[724]  & \A[725]  ;
  assign n7236 = ~\A[724]  & ~\A[725]  ;
  assign n7237 = ~n7235 & ~n7236 ;
  assign n7238 = \A[726]  & n7237 ;
  assign n7239 = ~\A[726]  & ~n7237 ;
  assign n7240 = ~n7238 & ~n7239 ;
  assign n7241 = n7234 & n7240 ;
  assign n7242 = ~n7234 & ~n7240 ;
  assign n7243 = ~n7241 & ~n7242 ;
  assign n7244 = n7228 & n7243 ;
  assign n7245 = ~n7235 & ~n7238 ;
  assign n7246 = ~n7229 & ~n7232 ;
  assign n7247 = n7245 & n7246 ;
  assign n7248 = ~n7245 & ~n7246 ;
  assign n7249 = ~n7247 & ~n7248 ;
  assign n7250 = n7244 & n7249 ;
  assign n7251 = ~n7214 & ~n7217 ;
  assign n7252 = n7220 & n7226 ;
  assign n7253 = ~n7220 & ~n7223 ;
  assign n7254 = ~n7226 & n7253 ;
  assign n7255 = ~n7252 & ~n7254 ;
  assign n7256 = n7251 & ~n7255 ;
  assign n7257 = ~n7251 & n7255 ;
  assign n7258 = ~n7256 & ~n7257 ;
  assign n7259 = ~n7250 & ~n7258 ;
  assign n7261 = n7241 & ~n7249 ;
  assign n7260 = ~n7241 & n7249 ;
  assign n7262 = ~n7244 & ~n7260 ;
  assign n7263 = ~n7261 & n7262 ;
  assign n7264 = ~n7259 & ~n7263 ;
  assign n7265 = n7241 & ~n7247 ;
  assign n7266 = ~n7248 & ~n7265 ;
  assign n7267 = n7264 & ~n7266 ;
  assign n7268 = ~n7264 & n7266 ;
  assign n7269 = ~n7251 & ~n7254 ;
  assign n7270 = ~n7252 & ~n7269 ;
  assign n7271 = ~n7268 & ~n7270 ;
  assign n7272 = ~n7267 & ~n7271 ;
  assign n7273 = \A[709]  & \A[710]  ;
  assign n7274 = ~\A[709]  & ~\A[710]  ;
  assign n7275 = ~n7273 & ~n7274 ;
  assign n7276 = \A[711]  & n7275 ;
  assign n7277 = ~\A[711]  & ~n7275 ;
  assign n7278 = ~n7276 & ~n7277 ;
  assign n7279 = \A[712]  & \A[713]  ;
  assign n7280 = ~\A[712]  & ~\A[713]  ;
  assign n7281 = ~n7279 & ~n7280 ;
  assign n7282 = \A[714]  & n7281 ;
  assign n7283 = ~\A[714]  & ~n7281 ;
  assign n7284 = ~n7282 & ~n7283 ;
  assign n7285 = n7278 & n7284 ;
  assign n7286 = ~n7278 & ~n7284 ;
  assign n7287 = ~n7285 & ~n7286 ;
  assign n7288 = \A[703]  & \A[704]  ;
  assign n7289 = ~\A[703]  & ~\A[704]  ;
  assign n7290 = ~n7288 & ~n7289 ;
  assign n7291 = \A[705]  & n7290 ;
  assign n7292 = ~\A[705]  & ~n7290 ;
  assign n7293 = ~n7291 & ~n7292 ;
  assign n7294 = \A[706]  & \A[707]  ;
  assign n7295 = ~\A[706]  & ~\A[707]  ;
  assign n7296 = ~n7294 & ~n7295 ;
  assign n7297 = \A[708]  & n7296 ;
  assign n7298 = ~\A[708]  & ~n7296 ;
  assign n7299 = ~n7297 & ~n7298 ;
  assign n7300 = n7293 & n7299 ;
  assign n7301 = ~n7293 & ~n7299 ;
  assign n7302 = ~n7300 & ~n7301 ;
  assign n7303 = n7287 & n7302 ;
  assign n7304 = ~n7279 & ~n7282 ;
  assign n7305 = ~n7273 & ~n7276 ;
  assign n7306 = ~n7304 & ~n7305 ;
  assign n7307 = n7304 & n7305 ;
  assign n7308 = ~n7306 & ~n7307 ;
  assign n7309 = n7303 & n7308 ;
  assign n7310 = ~n7294 & ~n7297 ;
  assign n7311 = ~n7288 & ~n7291 ;
  assign n7312 = ~n7310 & ~n7311 ;
  assign n7313 = n7310 & n7311 ;
  assign n7314 = ~n7312 & ~n7313 ;
  assign n7315 = n7300 & ~n7314 ;
  assign n7316 = ~n7300 & n7314 ;
  assign n7317 = ~n7315 & ~n7316 ;
  assign n7318 = ~n7309 & n7317 ;
  assign n7320 = n7285 & ~n7308 ;
  assign n7319 = ~n7285 & n7308 ;
  assign n7321 = ~n7303 & ~n7319 ;
  assign n7322 = ~n7320 & n7321 ;
  assign n7323 = ~n7318 & ~n7322 ;
  assign n7324 = ~n7285 & ~n7306 ;
  assign n7325 = ~n7307 & ~n7324 ;
  assign n7326 = ~n7323 & ~n7325 ;
  assign n7327 = n7323 & n7325 ;
  assign n7328 = ~n7300 & ~n7312 ;
  assign n7329 = ~n7313 & ~n7328 ;
  assign n7330 = ~n7327 & ~n7329 ;
  assign n7331 = ~n7326 & ~n7330 ;
  assign n7332 = ~n7272 & n7331 ;
  assign n7333 = n7272 & ~n7331 ;
  assign n7334 = ~n7332 & ~n7333 ;
  assign n7335 = ~n7326 & ~n7327 ;
  assign n7336 = ~n7329 & n7335 ;
  assign n7337 = n7329 & ~n7335 ;
  assign n7338 = ~n7336 & ~n7337 ;
  assign n7339 = ~n7267 & ~n7268 ;
  assign n7340 = ~n7270 & n7339 ;
  assign n7341 = n7270 & ~n7339 ;
  assign n7342 = ~n7340 & ~n7341 ;
  assign n7343 = ~n7338 & n7342 ;
  assign n7344 = n7338 & ~n7342 ;
  assign n7345 = ~n7228 & ~n7243 ;
  assign n7346 = ~n7244 & ~n7345 ;
  assign n7347 = ~n7287 & ~n7302 ;
  assign n7348 = ~n7303 & ~n7347 ;
  assign n7349 = n7346 & n7348 ;
  assign n7350 = ~n7250 & ~n7263 ;
  assign n7351 = ~n7258 & n7350 ;
  assign n7352 = n7258 & ~n7350 ;
  assign n7353 = ~n7351 & ~n7352 ;
  assign n7354 = n7349 & ~n7353 ;
  assign n7355 = ~n7349 & n7353 ;
  assign n7356 = ~n7309 & ~n7322 ;
  assign n7357 = n7317 & n7356 ;
  assign n7358 = ~n7317 & ~n7356 ;
  assign n7359 = ~n7357 & ~n7358 ;
  assign n7360 = ~n7355 & ~n7359 ;
  assign n7361 = ~n7354 & ~n7360 ;
  assign n7362 = ~n7344 & ~n7361 ;
  assign n7363 = ~n7343 & ~n7362 ;
  assign n7364 = n7334 & ~n7363 ;
  assign n7365 = ~n7334 & n7363 ;
  assign n7366 = ~n7364 & ~n7365 ;
  assign n7367 = n7213 & ~n7366 ;
  assign n7368 = ~n7213 & n7366 ;
  assign n7369 = ~n7343 & ~n7344 ;
  assign n7370 = ~n7361 & n7369 ;
  assign n7371 = n7361 & ~n7369 ;
  assign n7372 = ~n7370 & ~n7371 ;
  assign n7373 = ~n7190 & ~n7191 ;
  assign n7374 = ~n7208 & n7373 ;
  assign n7375 = n7208 & ~n7373 ;
  assign n7376 = ~n7374 & ~n7375 ;
  assign n7377 = ~n7372 & ~n7376 ;
  assign n7378 = n7372 & n7376 ;
  assign n7379 = ~n7193 & ~n7195 ;
  assign n7380 = ~n7196 & ~n7379 ;
  assign n7381 = ~n7346 & ~n7348 ;
  assign n7382 = ~n7349 & ~n7381 ;
  assign n7383 = n7380 & n7382 ;
  assign n7384 = ~n7201 & ~n7202 ;
  assign n7385 = ~n7206 & n7384 ;
  assign n7386 = n7206 & ~n7384 ;
  assign n7387 = ~n7385 & ~n7386 ;
  assign n7388 = n7383 & n7387 ;
  assign n7389 = ~n7383 & ~n7387 ;
  assign n7390 = ~n7354 & ~n7355 ;
  assign n7391 = ~n7359 & n7390 ;
  assign n7392 = n7359 & ~n7390 ;
  assign n7393 = ~n7391 & ~n7392 ;
  assign n7394 = ~n7389 & n7393 ;
  assign n7395 = ~n7388 & ~n7394 ;
  assign n7396 = ~n7378 & n7395 ;
  assign n7397 = ~n7377 & ~n7396 ;
  assign n7398 = ~n7368 & ~n7397 ;
  assign n7399 = ~n7367 & ~n7398 ;
  assign n7400 = ~n7180 & n7210 ;
  assign n7401 = ~n7179 & ~n7400 ;
  assign n7402 = n7399 & ~n7401 ;
  assign n7403 = ~n7399 & n7401 ;
  assign n7404 = ~n7333 & ~n7363 ;
  assign n7405 = ~n7332 & ~n7404 ;
  assign n7406 = ~n7403 & ~n7405 ;
  assign n7407 = ~n7402 & ~n7406 ;
  assign n7408 = \A[658]  & \A[659]  ;
  assign n7409 = \A[655]  & \A[656]  ;
  assign n7410 = ~\A[655]  & ~\A[656]  ;
  assign n7411 = ~n7409 & ~n7410 ;
  assign n7412 = \A[657]  & n7411 ;
  assign n7413 = ~\A[657]  & ~n7411 ;
  assign n7414 = ~n7412 & ~n7413 ;
  assign n7415 = ~\A[658]  & ~\A[659]  ;
  assign n7416 = ~n7408 & ~n7415 ;
  assign n7417 = \A[660]  & n7416 ;
  assign n7418 = ~\A[660]  & ~n7416 ;
  assign n7419 = ~n7417 & ~n7418 ;
  assign n7420 = n7414 & n7419 ;
  assign n7421 = n7408 & n7420 ;
  assign n7422 = ~n7409 & ~n7412 ;
  assign n7423 = ~n7408 & ~n7417 ;
  assign n7424 = ~n7420 & n7423 ;
  assign n7425 = ~n7422 & ~n7424 ;
  assign n7426 = ~n7421 & ~n7425 ;
  assign n7427 = \A[664]  & \A[665]  ;
  assign n7428 = ~\A[664]  & ~\A[665]  ;
  assign n7429 = ~n7427 & ~n7428 ;
  assign n7430 = \A[666]  & n7429 ;
  assign n7431 = ~n7427 & ~n7430 ;
  assign n7432 = \A[661]  & \A[662]  ;
  assign n7433 = ~\A[661]  & ~\A[662]  ;
  assign n7434 = ~n7432 & ~n7433 ;
  assign n7435 = \A[663]  & n7434 ;
  assign n7436 = ~n7432 & ~n7435 ;
  assign n7437 = n7431 & n7436 ;
  assign n7438 = ~n7431 & ~n7436 ;
  assign n7439 = ~\A[663]  & ~n7434 ;
  assign n7440 = ~n7435 & ~n7439 ;
  assign n7441 = ~\A[666]  & ~n7429 ;
  assign n7442 = ~n7430 & ~n7441 ;
  assign n7443 = n7440 & n7442 ;
  assign n7444 = ~n7438 & ~n7443 ;
  assign n7445 = ~n7437 & ~n7444 ;
  assign n7446 = ~n7440 & ~n7442 ;
  assign n7447 = ~n7443 & ~n7446 ;
  assign n7448 = ~n7414 & ~n7419 ;
  assign n7449 = ~n7420 & ~n7448 ;
  assign n7450 = n7447 & n7449 ;
  assign n7451 = n7421 & ~n7422 ;
  assign n7452 = n7450 & ~n7451 ;
  assign n7453 = ~n7437 & ~n7438 ;
  assign n7454 = n7443 & ~n7453 ;
  assign n7455 = ~n7443 & n7453 ;
  assign n7456 = ~n7454 & ~n7455 ;
  assign n7457 = n7452 & ~n7456 ;
  assign n7458 = ~n7452 & n7456 ;
  assign n7459 = ~n7421 & ~n7424 ;
  assign n7460 = n7422 & ~n7459 ;
  assign n7461 = ~n7422 & n7459 ;
  assign n7462 = ~n7460 & ~n7461 ;
  assign n7463 = ~n7458 & n7462 ;
  assign n7464 = ~n7457 & ~n7463 ;
  assign n7465 = n7445 & ~n7464 ;
  assign n7466 = ~n7445 & n7464 ;
  assign n7467 = ~n7465 & ~n7466 ;
  assign n7468 = n7426 & n7467 ;
  assign n7469 = ~n7426 & ~n7467 ;
  assign n7470 = ~n7468 & ~n7469 ;
  assign n7471 = \A[670]  & \A[671]  ;
  assign n7472 = \A[667]  & \A[668]  ;
  assign n7473 = ~\A[667]  & ~\A[668]  ;
  assign n7474 = ~n7472 & ~n7473 ;
  assign n7475 = \A[669]  & n7474 ;
  assign n7476 = ~\A[669]  & ~n7474 ;
  assign n7477 = ~n7475 & ~n7476 ;
  assign n7478 = ~\A[670]  & ~\A[671]  ;
  assign n7479 = ~n7471 & ~n7478 ;
  assign n7480 = \A[672]  & n7479 ;
  assign n7481 = ~\A[672]  & ~n7479 ;
  assign n7482 = ~n7480 & ~n7481 ;
  assign n7483 = n7477 & n7482 ;
  assign n7484 = n7471 & n7483 ;
  assign n7485 = ~n7472 & ~n7475 ;
  assign n7486 = ~n7471 & ~n7480 ;
  assign n7487 = ~n7483 & n7486 ;
  assign n7488 = ~n7485 & ~n7487 ;
  assign n7489 = ~n7484 & ~n7488 ;
  assign n7490 = \A[676]  & \A[677]  ;
  assign n7491 = ~\A[676]  & ~\A[677]  ;
  assign n7492 = ~n7490 & ~n7491 ;
  assign n7493 = \A[678]  & n7492 ;
  assign n7494 = ~n7490 & ~n7493 ;
  assign n7495 = \A[673]  & \A[674]  ;
  assign n7496 = ~\A[673]  & ~\A[674]  ;
  assign n7497 = ~n7495 & ~n7496 ;
  assign n7498 = \A[675]  & n7497 ;
  assign n7499 = ~n7495 & ~n7498 ;
  assign n7500 = n7494 & n7499 ;
  assign n7501 = ~n7494 & ~n7499 ;
  assign n7502 = ~\A[675]  & ~n7497 ;
  assign n7503 = ~n7498 & ~n7502 ;
  assign n7504 = ~\A[678]  & ~n7492 ;
  assign n7505 = ~n7493 & ~n7504 ;
  assign n7506 = n7503 & n7505 ;
  assign n7507 = ~n7501 & ~n7506 ;
  assign n7508 = ~n7500 & ~n7507 ;
  assign n7509 = ~n7503 & ~n7505 ;
  assign n7510 = ~n7506 & ~n7509 ;
  assign n7511 = ~n7477 & ~n7482 ;
  assign n7512 = ~n7483 & ~n7511 ;
  assign n7513 = n7510 & n7512 ;
  assign n7514 = n7484 & ~n7485 ;
  assign n7515 = n7513 & ~n7514 ;
  assign n7516 = ~n7500 & ~n7501 ;
  assign n7517 = n7506 & ~n7516 ;
  assign n7518 = ~n7506 & n7516 ;
  assign n7519 = ~n7517 & ~n7518 ;
  assign n7520 = n7515 & ~n7519 ;
  assign n7521 = ~n7515 & n7519 ;
  assign n7522 = ~n7484 & ~n7487 ;
  assign n7523 = n7485 & ~n7522 ;
  assign n7524 = ~n7485 & n7522 ;
  assign n7525 = ~n7523 & ~n7524 ;
  assign n7526 = ~n7521 & n7525 ;
  assign n7527 = ~n7520 & ~n7526 ;
  assign n7528 = n7508 & ~n7527 ;
  assign n7529 = ~n7508 & n7527 ;
  assign n7530 = ~n7528 & ~n7529 ;
  assign n7531 = n7489 & n7530 ;
  assign n7532 = ~n7489 & ~n7530 ;
  assign n7533 = ~n7531 & ~n7532 ;
  assign n7534 = ~n7470 & ~n7533 ;
  assign n7535 = n7470 & n7533 ;
  assign n7536 = ~n7510 & ~n7512 ;
  assign n7537 = ~n7513 & ~n7536 ;
  assign n7538 = ~n7447 & ~n7449 ;
  assign n7539 = ~n7450 & ~n7538 ;
  assign n7540 = n7537 & n7539 ;
  assign n7541 = ~n7520 & ~n7521 ;
  assign n7542 = n7525 & n7541 ;
  assign n7543 = ~n7525 & ~n7541 ;
  assign n7544 = ~n7542 & ~n7543 ;
  assign n7545 = n7540 & n7544 ;
  assign n7546 = ~n7540 & ~n7544 ;
  assign n7547 = ~n7457 & ~n7458 ;
  assign n7548 = n7462 & n7547 ;
  assign n7549 = ~n7462 & ~n7547 ;
  assign n7550 = ~n7548 & ~n7549 ;
  assign n7551 = ~n7546 & n7550 ;
  assign n7552 = ~n7545 & ~n7551 ;
  assign n7553 = ~n7535 & ~n7552 ;
  assign n7554 = ~n7534 & ~n7553 ;
  assign n7555 = ~n7489 & ~n7529 ;
  assign n7556 = ~n7528 & ~n7555 ;
  assign n7557 = ~n7554 & ~n7556 ;
  assign n7558 = n7554 & n7556 ;
  assign n7559 = ~n7426 & ~n7466 ;
  assign n7560 = ~n7465 & ~n7559 ;
  assign n7561 = ~n7558 & ~n7560 ;
  assign n7562 = ~n7557 & ~n7561 ;
  assign n7563 = \A[682]  & \A[683]  ;
  assign n7564 = \A[679]  & \A[680]  ;
  assign n7565 = ~\A[679]  & ~\A[680]  ;
  assign n7566 = ~n7564 & ~n7565 ;
  assign n7567 = \A[681]  & n7566 ;
  assign n7568 = ~\A[681]  & ~n7566 ;
  assign n7569 = ~n7567 & ~n7568 ;
  assign n7570 = ~\A[682]  & ~\A[683]  ;
  assign n7571 = ~n7563 & ~n7570 ;
  assign n7572 = \A[684]  & n7571 ;
  assign n7573 = ~\A[684]  & ~n7571 ;
  assign n7574 = ~n7572 & ~n7573 ;
  assign n7575 = n7569 & n7574 ;
  assign n7576 = n7563 & n7575 ;
  assign n7577 = ~n7564 & ~n7567 ;
  assign n7578 = ~n7563 & ~n7572 ;
  assign n7579 = ~n7575 & n7578 ;
  assign n7580 = ~n7577 & ~n7579 ;
  assign n7581 = ~n7576 & ~n7580 ;
  assign n7582 = \A[688]  & \A[689]  ;
  assign n7583 = ~\A[688]  & ~\A[689]  ;
  assign n7584 = ~n7582 & ~n7583 ;
  assign n7585 = \A[690]  & n7584 ;
  assign n7586 = ~n7582 & ~n7585 ;
  assign n7587 = \A[685]  & \A[686]  ;
  assign n7588 = ~\A[685]  & ~\A[686]  ;
  assign n7589 = ~n7587 & ~n7588 ;
  assign n7590 = \A[687]  & n7589 ;
  assign n7591 = ~n7587 & ~n7590 ;
  assign n7592 = n7586 & n7591 ;
  assign n7593 = ~n7586 & ~n7591 ;
  assign n7594 = ~\A[687]  & ~n7589 ;
  assign n7595 = ~n7590 & ~n7594 ;
  assign n7596 = ~\A[690]  & ~n7584 ;
  assign n7597 = ~n7585 & ~n7596 ;
  assign n7598 = n7595 & n7597 ;
  assign n7599 = ~n7593 & ~n7598 ;
  assign n7600 = ~n7592 & ~n7599 ;
  assign n7601 = ~n7595 & ~n7597 ;
  assign n7602 = ~n7598 & ~n7601 ;
  assign n7603 = ~n7569 & ~n7574 ;
  assign n7604 = ~n7575 & ~n7603 ;
  assign n7605 = n7602 & n7604 ;
  assign n7606 = n7576 & ~n7577 ;
  assign n7607 = n7605 & ~n7606 ;
  assign n7608 = ~n7592 & ~n7593 ;
  assign n7609 = n7598 & ~n7608 ;
  assign n7610 = ~n7598 & n7608 ;
  assign n7611 = ~n7609 & ~n7610 ;
  assign n7612 = n7607 & ~n7611 ;
  assign n7613 = ~n7607 & n7611 ;
  assign n7614 = ~n7576 & ~n7579 ;
  assign n7615 = n7577 & ~n7614 ;
  assign n7616 = ~n7577 & n7614 ;
  assign n7617 = ~n7615 & ~n7616 ;
  assign n7618 = ~n7613 & n7617 ;
  assign n7619 = ~n7612 & ~n7618 ;
  assign n7620 = n7600 & ~n7619 ;
  assign n7621 = ~n7600 & n7619 ;
  assign n7622 = ~n7620 & ~n7621 ;
  assign n7623 = n7581 & n7622 ;
  assign n7624 = ~n7581 & ~n7622 ;
  assign n7625 = ~n7623 & ~n7624 ;
  assign n7626 = \A[694]  & \A[695]  ;
  assign n7627 = \A[691]  & \A[692]  ;
  assign n7628 = ~\A[691]  & ~\A[692]  ;
  assign n7629 = ~n7627 & ~n7628 ;
  assign n7630 = \A[693]  & n7629 ;
  assign n7631 = ~\A[693]  & ~n7629 ;
  assign n7632 = ~n7630 & ~n7631 ;
  assign n7633 = ~\A[694]  & ~\A[695]  ;
  assign n7634 = ~n7626 & ~n7633 ;
  assign n7635 = \A[696]  & n7634 ;
  assign n7636 = ~\A[696]  & ~n7634 ;
  assign n7637 = ~n7635 & ~n7636 ;
  assign n7638 = n7632 & n7637 ;
  assign n7639 = n7626 & n7638 ;
  assign n7640 = ~n7627 & ~n7630 ;
  assign n7641 = ~n7626 & ~n7635 ;
  assign n7642 = ~n7638 & n7641 ;
  assign n7643 = ~n7640 & ~n7642 ;
  assign n7644 = ~n7639 & ~n7643 ;
  assign n7645 = \A[700]  & \A[701]  ;
  assign n7646 = ~\A[700]  & ~\A[701]  ;
  assign n7647 = ~n7645 & ~n7646 ;
  assign n7648 = \A[702]  & n7647 ;
  assign n7649 = ~n7645 & ~n7648 ;
  assign n7650 = \A[697]  & \A[698]  ;
  assign n7651 = ~\A[697]  & ~\A[698]  ;
  assign n7652 = ~n7650 & ~n7651 ;
  assign n7653 = \A[699]  & n7652 ;
  assign n7654 = ~n7650 & ~n7653 ;
  assign n7655 = n7649 & n7654 ;
  assign n7656 = ~n7649 & ~n7654 ;
  assign n7657 = ~\A[699]  & ~n7652 ;
  assign n7658 = ~n7653 & ~n7657 ;
  assign n7659 = ~\A[702]  & ~n7647 ;
  assign n7660 = ~n7648 & ~n7659 ;
  assign n7661 = n7658 & n7660 ;
  assign n7662 = ~n7656 & ~n7661 ;
  assign n7663 = ~n7655 & ~n7662 ;
  assign n7664 = ~n7658 & ~n7660 ;
  assign n7665 = ~n7661 & ~n7664 ;
  assign n7666 = ~n7632 & ~n7637 ;
  assign n7667 = ~n7638 & ~n7666 ;
  assign n7668 = n7665 & n7667 ;
  assign n7669 = n7639 & ~n7640 ;
  assign n7670 = n7668 & ~n7669 ;
  assign n7671 = ~n7655 & ~n7656 ;
  assign n7672 = n7661 & ~n7671 ;
  assign n7673 = ~n7661 & n7671 ;
  assign n7674 = ~n7672 & ~n7673 ;
  assign n7675 = n7670 & ~n7674 ;
  assign n7676 = ~n7670 & n7674 ;
  assign n7677 = ~n7639 & ~n7642 ;
  assign n7678 = n7640 & ~n7677 ;
  assign n7679 = ~n7640 & n7677 ;
  assign n7680 = ~n7678 & ~n7679 ;
  assign n7681 = ~n7676 & n7680 ;
  assign n7682 = ~n7675 & ~n7681 ;
  assign n7683 = n7663 & ~n7682 ;
  assign n7684 = ~n7663 & n7682 ;
  assign n7685 = ~n7683 & ~n7684 ;
  assign n7686 = n7644 & n7685 ;
  assign n7687 = ~n7644 & ~n7685 ;
  assign n7688 = ~n7686 & ~n7687 ;
  assign n7689 = ~n7625 & ~n7688 ;
  assign n7690 = n7625 & n7688 ;
  assign n7691 = ~n7665 & ~n7667 ;
  assign n7692 = ~n7668 & ~n7691 ;
  assign n7693 = ~n7602 & ~n7604 ;
  assign n7694 = ~n7605 & ~n7693 ;
  assign n7695 = n7692 & n7694 ;
  assign n7696 = ~n7675 & ~n7676 ;
  assign n7697 = n7680 & n7696 ;
  assign n7698 = ~n7680 & ~n7696 ;
  assign n7699 = ~n7697 & ~n7698 ;
  assign n7700 = n7695 & n7699 ;
  assign n7701 = ~n7695 & ~n7699 ;
  assign n7702 = ~n7612 & ~n7613 ;
  assign n7703 = n7617 & n7702 ;
  assign n7704 = ~n7617 & ~n7702 ;
  assign n7705 = ~n7703 & ~n7704 ;
  assign n7706 = ~n7701 & n7705 ;
  assign n7707 = ~n7700 & ~n7706 ;
  assign n7708 = ~n7690 & ~n7707 ;
  assign n7709 = ~n7689 & ~n7708 ;
  assign n7710 = ~n7644 & ~n7684 ;
  assign n7711 = ~n7683 & ~n7710 ;
  assign n7712 = ~n7709 & ~n7711 ;
  assign n7713 = n7709 & n7711 ;
  assign n7714 = ~n7712 & ~n7713 ;
  assign n7715 = ~n7581 & ~n7621 ;
  assign n7716 = ~n7620 & ~n7715 ;
  assign n7717 = n7714 & ~n7716 ;
  assign n7718 = ~n7714 & n7716 ;
  assign n7719 = ~n7717 & ~n7718 ;
  assign n7720 = ~n7557 & ~n7558 ;
  assign n7721 = ~n7560 & n7720 ;
  assign n7722 = n7560 & ~n7720 ;
  assign n7723 = ~n7721 & ~n7722 ;
  assign n7724 = ~n7719 & ~n7723 ;
  assign n7725 = n7719 & n7723 ;
  assign n7726 = ~n7534 & ~n7535 ;
  assign n7727 = ~n7552 & n7726 ;
  assign n7728 = n7552 & ~n7726 ;
  assign n7729 = ~n7727 & ~n7728 ;
  assign n7730 = ~n7689 & ~n7690 ;
  assign n7731 = ~n7707 & n7730 ;
  assign n7732 = n7707 & ~n7730 ;
  assign n7733 = ~n7731 & ~n7732 ;
  assign n7734 = ~n7729 & ~n7733 ;
  assign n7735 = n7729 & n7733 ;
  assign n7736 = ~n7692 & ~n7694 ;
  assign n7737 = ~n7695 & ~n7736 ;
  assign n7738 = ~n7537 & ~n7539 ;
  assign n7739 = ~n7540 & ~n7738 ;
  assign n7740 = n7737 & n7739 ;
  assign n7741 = ~n7700 & ~n7701 ;
  assign n7742 = ~n7705 & n7741 ;
  assign n7743 = n7705 & ~n7741 ;
  assign n7744 = ~n7742 & ~n7743 ;
  assign n7745 = n7740 & ~n7744 ;
  assign n7746 = ~n7740 & n7744 ;
  assign n7747 = ~n7545 & ~n7546 ;
  assign n7748 = ~n7550 & n7747 ;
  assign n7749 = n7550 & ~n7747 ;
  assign n7750 = ~n7748 & ~n7749 ;
  assign n7751 = ~n7746 & ~n7750 ;
  assign n7752 = ~n7745 & ~n7751 ;
  assign n7753 = ~n7735 & n7752 ;
  assign n7754 = ~n7734 & ~n7753 ;
  assign n7755 = ~n7725 & ~n7754 ;
  assign n7756 = ~n7724 & ~n7755 ;
  assign n7757 = n7562 & ~n7756 ;
  assign n7758 = ~n7562 & n7756 ;
  assign n7759 = ~n7713 & ~n7716 ;
  assign n7760 = ~n7712 & ~n7759 ;
  assign n7761 = ~n7758 & n7760 ;
  assign n7762 = ~n7757 & ~n7761 ;
  assign n7763 = ~n7407 & n7762 ;
  assign n7764 = n7407 & ~n7762 ;
  assign n7765 = ~n7757 & ~n7758 ;
  assign n7766 = n7760 & n7765 ;
  assign n7767 = ~n7760 & ~n7765 ;
  assign n7768 = ~n7766 & ~n7767 ;
  assign n7769 = ~n7402 & ~n7403 ;
  assign n7770 = ~n7405 & n7769 ;
  assign n7771 = n7405 & ~n7769 ;
  assign n7772 = ~n7770 & ~n7771 ;
  assign n7773 = ~n7768 & n7772 ;
  assign n7774 = n7768 & ~n7772 ;
  assign n7775 = ~n7367 & ~n7368 ;
  assign n7776 = ~n7397 & n7775 ;
  assign n7777 = n7397 & ~n7775 ;
  assign n7778 = ~n7776 & ~n7777 ;
  assign n7779 = ~n7724 & ~n7725 ;
  assign n7780 = ~n7754 & n7779 ;
  assign n7781 = n7754 & ~n7779 ;
  assign n7782 = ~n7780 & ~n7781 ;
  assign n7783 = ~n7778 & ~n7782 ;
  assign n7784 = n7778 & n7782 ;
  assign n7785 = ~n7734 & ~n7735 ;
  assign n7786 = ~n7752 & n7785 ;
  assign n7787 = n7752 & ~n7785 ;
  assign n7788 = ~n7786 & ~n7787 ;
  assign n7789 = ~n7377 & ~n7378 ;
  assign n7790 = ~n7395 & n7789 ;
  assign n7791 = n7395 & ~n7789 ;
  assign n7792 = ~n7790 & ~n7791 ;
  assign n7793 = ~n7788 & ~n7792 ;
  assign n7794 = n7788 & n7792 ;
  assign n7795 = ~n7380 & ~n7382 ;
  assign n7796 = ~n7383 & ~n7795 ;
  assign n7797 = ~n7737 & ~n7739 ;
  assign n7798 = ~n7740 & ~n7797 ;
  assign n7799 = n7796 & n7798 ;
  assign n7800 = ~n7388 & ~n7389 ;
  assign n7801 = ~n7393 & n7800 ;
  assign n7802 = n7393 & ~n7800 ;
  assign n7803 = ~n7801 & ~n7802 ;
  assign n7804 = n7799 & ~n7803 ;
  assign n7805 = ~n7799 & n7803 ;
  assign n7806 = ~n7745 & ~n7746 ;
  assign n7807 = ~n7750 & n7806 ;
  assign n7808 = n7750 & ~n7806 ;
  assign n7809 = ~n7807 & ~n7808 ;
  assign n7810 = ~n7805 & n7809 ;
  assign n7811 = ~n7804 & ~n7810 ;
  assign n7812 = ~n7794 & n7811 ;
  assign n7813 = ~n7793 & ~n7812 ;
  assign n7814 = ~n7784 & n7813 ;
  assign n7815 = ~n7783 & ~n7814 ;
  assign n7816 = ~n7774 & ~n7815 ;
  assign n7817 = ~n7773 & ~n7816 ;
  assign n7818 = ~n7764 & ~n7817 ;
  assign n7819 = ~n7763 & ~n7818 ;
  assign n7820 = ~n7060 & ~n7819 ;
  assign n7821 = n7060 & n7819 ;
  assign n7822 = ~n7004 & ~n7005 ;
  assign n7823 = ~n7058 & n7822 ;
  assign n7824 = n7058 & ~n7822 ;
  assign n7825 = ~n7823 & ~n7824 ;
  assign n7826 = ~n7763 & ~n7764 ;
  assign n7827 = ~n7817 & n7826 ;
  assign n7828 = n7817 & ~n7826 ;
  assign n7829 = ~n7827 & ~n7828 ;
  assign n7830 = ~n7825 & ~n7829 ;
  assign n7831 = n7825 & n7829 ;
  assign n7832 = ~n7014 & ~n7015 ;
  assign n7833 = ~n7056 & n7832 ;
  assign n7834 = n7056 & ~n7832 ;
  assign n7835 = ~n7833 & ~n7834 ;
  assign n7836 = ~n7773 & ~n7774 ;
  assign n7837 = ~n7815 & n7836 ;
  assign n7838 = n7815 & ~n7836 ;
  assign n7839 = ~n7837 & ~n7838 ;
  assign n7840 = n7835 & ~n7839 ;
  assign n7841 = ~n7835 & n7839 ;
  assign n7842 = ~n7024 & ~n7025 ;
  assign n7843 = ~n7054 & n7842 ;
  assign n7844 = n7054 & ~n7842 ;
  assign n7845 = ~n7843 & ~n7844 ;
  assign n7846 = ~n7783 & ~n7784 ;
  assign n7847 = n7813 & n7846 ;
  assign n7848 = ~n7813 & ~n7846 ;
  assign n7849 = ~n7847 & ~n7848 ;
  assign n7850 = n7845 & ~n7849 ;
  assign n7851 = ~n7845 & n7849 ;
  assign n7852 = ~n7793 & ~n7794 ;
  assign n7853 = ~n7811 & n7852 ;
  assign n7854 = n7811 & ~n7852 ;
  assign n7855 = ~n7853 & ~n7854 ;
  assign n7856 = ~n7034 & ~n7035 ;
  assign n7857 = ~n7052 & n7856 ;
  assign n7858 = n7052 & ~n7856 ;
  assign n7859 = ~n7857 & ~n7858 ;
  assign n7860 = ~n7855 & ~n7859 ;
  assign n7861 = n7855 & n7859 ;
  assign n7862 = ~n7037 & ~n7039 ;
  assign n7863 = ~n7040 & ~n7862 ;
  assign n7864 = ~n7796 & ~n7798 ;
  assign n7865 = ~n7799 & ~n7864 ;
  assign n7866 = n7863 & n7865 ;
  assign n7867 = ~n7045 & ~n7046 ;
  assign n7868 = ~n7050 & n7867 ;
  assign n7869 = n7050 & ~n7867 ;
  assign n7870 = ~n7868 & ~n7869 ;
  assign n7871 = n7866 & n7870 ;
  assign n7872 = ~n7866 & ~n7870 ;
  assign n7873 = ~n7804 & ~n7805 ;
  assign n7874 = ~n7809 & n7873 ;
  assign n7875 = n7809 & ~n7873 ;
  assign n7876 = ~n7874 & ~n7875 ;
  assign n7877 = ~n7872 & ~n7876 ;
  assign n7878 = ~n7871 & ~n7877 ;
  assign n7879 = ~n7861 & n7878 ;
  assign n7880 = ~n7860 & ~n7879 ;
  assign n7881 = ~n7851 & ~n7880 ;
  assign n7882 = ~n7850 & ~n7881 ;
  assign n7883 = ~n7841 & ~n7882 ;
  assign n7884 = ~n7840 & ~n7883 ;
  assign n7885 = ~n7831 & ~n7884 ;
  assign n7886 = ~n7830 & ~n7885 ;
  assign n7887 = ~n7821 & n7886 ;
  assign n7888 = ~n7820 & ~n7887 ;
  assign n7889 = \A[562]  & \A[563]  ;
  assign n7890 = \A[559]  & \A[560]  ;
  assign n7891 = ~\A[559]  & ~\A[560]  ;
  assign n7892 = ~n7890 & ~n7891 ;
  assign n7893 = \A[561]  & n7892 ;
  assign n7894 = ~\A[561]  & ~n7892 ;
  assign n7895 = ~n7893 & ~n7894 ;
  assign n7896 = ~\A[562]  & ~\A[563]  ;
  assign n7897 = ~n7889 & ~n7896 ;
  assign n7898 = \A[564]  & n7897 ;
  assign n7899 = ~\A[564]  & ~n7897 ;
  assign n7900 = ~n7898 & ~n7899 ;
  assign n7901 = n7895 & n7900 ;
  assign n7902 = n7889 & n7901 ;
  assign n7903 = ~n7890 & ~n7893 ;
  assign n7904 = ~n7889 & ~n7898 ;
  assign n7905 = ~n7901 & n7904 ;
  assign n7906 = ~n7903 & ~n7905 ;
  assign n7907 = ~n7902 & ~n7906 ;
  assign n7908 = \A[568]  & \A[569]  ;
  assign n7909 = ~\A[568]  & ~\A[569]  ;
  assign n7910 = ~n7908 & ~n7909 ;
  assign n7911 = \A[570]  & n7910 ;
  assign n7912 = ~n7908 & ~n7911 ;
  assign n7913 = \A[565]  & \A[566]  ;
  assign n7914 = ~\A[565]  & ~\A[566]  ;
  assign n7915 = ~n7913 & ~n7914 ;
  assign n7916 = \A[567]  & n7915 ;
  assign n7917 = ~n7913 & ~n7916 ;
  assign n7918 = n7912 & n7917 ;
  assign n7919 = ~n7912 & ~n7917 ;
  assign n7920 = ~\A[567]  & ~n7915 ;
  assign n7921 = ~n7916 & ~n7920 ;
  assign n7922 = ~\A[570]  & ~n7910 ;
  assign n7923 = ~n7911 & ~n7922 ;
  assign n7924 = n7921 & n7923 ;
  assign n7925 = ~n7919 & ~n7924 ;
  assign n7926 = ~n7918 & ~n7925 ;
  assign n7927 = ~n7921 & ~n7923 ;
  assign n7928 = ~n7924 & ~n7927 ;
  assign n7929 = ~n7895 & ~n7900 ;
  assign n7930 = ~n7901 & ~n7929 ;
  assign n7931 = n7928 & n7930 ;
  assign n7932 = n7902 & ~n7903 ;
  assign n7933 = n7931 & ~n7932 ;
  assign n7934 = ~n7918 & ~n7919 ;
  assign n7935 = n7924 & ~n7934 ;
  assign n7936 = ~n7924 & n7934 ;
  assign n7937 = ~n7935 & ~n7936 ;
  assign n7938 = n7933 & ~n7937 ;
  assign n7939 = ~n7933 & n7937 ;
  assign n7940 = ~n7902 & ~n7905 ;
  assign n7941 = n7903 & ~n7940 ;
  assign n7942 = ~n7903 & n7940 ;
  assign n7943 = ~n7941 & ~n7942 ;
  assign n7944 = ~n7939 & n7943 ;
  assign n7945 = ~n7938 & ~n7944 ;
  assign n7946 = n7926 & ~n7945 ;
  assign n7947 = ~n7926 & n7945 ;
  assign n7948 = ~n7946 & ~n7947 ;
  assign n7949 = n7907 & n7948 ;
  assign n7950 = ~n7907 & ~n7948 ;
  assign n7951 = ~n7949 & ~n7950 ;
  assign n7952 = \A[574]  & \A[575]  ;
  assign n7953 = \A[571]  & \A[572]  ;
  assign n7954 = ~\A[571]  & ~\A[572]  ;
  assign n7955 = ~n7953 & ~n7954 ;
  assign n7956 = \A[573]  & n7955 ;
  assign n7957 = ~\A[573]  & ~n7955 ;
  assign n7958 = ~n7956 & ~n7957 ;
  assign n7959 = ~\A[574]  & ~\A[575]  ;
  assign n7960 = ~n7952 & ~n7959 ;
  assign n7961 = \A[576]  & n7960 ;
  assign n7962 = ~\A[576]  & ~n7960 ;
  assign n7963 = ~n7961 & ~n7962 ;
  assign n7964 = n7958 & n7963 ;
  assign n7965 = n7952 & n7964 ;
  assign n7966 = ~n7953 & ~n7956 ;
  assign n7967 = ~n7952 & ~n7961 ;
  assign n7968 = ~n7964 & n7967 ;
  assign n7969 = ~n7966 & ~n7968 ;
  assign n7970 = ~n7965 & ~n7969 ;
  assign n7971 = \A[580]  & \A[581]  ;
  assign n7972 = ~\A[580]  & ~\A[581]  ;
  assign n7973 = ~n7971 & ~n7972 ;
  assign n7974 = \A[582]  & n7973 ;
  assign n7975 = ~n7971 & ~n7974 ;
  assign n7976 = \A[577]  & \A[578]  ;
  assign n7977 = ~\A[577]  & ~\A[578]  ;
  assign n7978 = ~n7976 & ~n7977 ;
  assign n7979 = \A[579]  & n7978 ;
  assign n7980 = ~n7976 & ~n7979 ;
  assign n7981 = n7975 & n7980 ;
  assign n7982 = ~n7975 & ~n7980 ;
  assign n7983 = ~\A[579]  & ~n7978 ;
  assign n7984 = ~n7979 & ~n7983 ;
  assign n7985 = ~\A[582]  & ~n7973 ;
  assign n7986 = ~n7974 & ~n7985 ;
  assign n7987 = n7984 & n7986 ;
  assign n7988 = ~n7982 & ~n7987 ;
  assign n7989 = ~n7981 & ~n7988 ;
  assign n7990 = ~n7984 & ~n7986 ;
  assign n7991 = ~n7987 & ~n7990 ;
  assign n7992 = ~n7958 & ~n7963 ;
  assign n7993 = ~n7964 & ~n7992 ;
  assign n7994 = n7991 & n7993 ;
  assign n7995 = n7965 & ~n7966 ;
  assign n7996 = n7994 & ~n7995 ;
  assign n7997 = ~n7981 & ~n7982 ;
  assign n7998 = n7987 & ~n7997 ;
  assign n7999 = ~n7987 & n7997 ;
  assign n8000 = ~n7998 & ~n7999 ;
  assign n8001 = n7996 & ~n8000 ;
  assign n8002 = ~n7996 & n8000 ;
  assign n8003 = ~n7965 & ~n7968 ;
  assign n8004 = n7966 & ~n8003 ;
  assign n8005 = ~n7966 & n8003 ;
  assign n8006 = ~n8004 & ~n8005 ;
  assign n8007 = ~n8002 & n8006 ;
  assign n8008 = ~n8001 & ~n8007 ;
  assign n8009 = n7989 & ~n8008 ;
  assign n8010 = ~n7989 & n8008 ;
  assign n8011 = ~n8009 & ~n8010 ;
  assign n8012 = n7970 & n8011 ;
  assign n8013 = ~n7970 & ~n8011 ;
  assign n8014 = ~n8012 & ~n8013 ;
  assign n8015 = ~n7951 & ~n8014 ;
  assign n8016 = n7951 & n8014 ;
  assign n8017 = ~n7991 & ~n7993 ;
  assign n8018 = ~n7994 & ~n8017 ;
  assign n8019 = ~n7928 & ~n7930 ;
  assign n8020 = ~n7931 & ~n8019 ;
  assign n8021 = n8018 & n8020 ;
  assign n8022 = ~n8001 & ~n8002 ;
  assign n8023 = n8006 & n8022 ;
  assign n8024 = ~n8006 & ~n8022 ;
  assign n8025 = ~n8023 & ~n8024 ;
  assign n8026 = n8021 & n8025 ;
  assign n8027 = ~n8021 & ~n8025 ;
  assign n8028 = ~n7938 & ~n7939 ;
  assign n8029 = n7943 & n8028 ;
  assign n8030 = ~n7943 & ~n8028 ;
  assign n8031 = ~n8029 & ~n8030 ;
  assign n8032 = ~n8027 & n8031 ;
  assign n8033 = ~n8026 & ~n8032 ;
  assign n8034 = ~n8016 & ~n8033 ;
  assign n8035 = ~n8015 & ~n8034 ;
  assign n8036 = ~n7970 & ~n8010 ;
  assign n8037 = ~n8009 & ~n8036 ;
  assign n8038 = ~n8035 & ~n8037 ;
  assign n8039 = n8035 & n8037 ;
  assign n8040 = ~n7907 & ~n7947 ;
  assign n8041 = ~n7946 & ~n8040 ;
  assign n8042 = ~n8039 & ~n8041 ;
  assign n8043 = ~n8038 & ~n8042 ;
  assign n8044 = \A[586]  & \A[587]  ;
  assign n8045 = \A[583]  & \A[584]  ;
  assign n8046 = ~\A[583]  & ~\A[584]  ;
  assign n8047 = ~n8045 & ~n8046 ;
  assign n8048 = \A[585]  & n8047 ;
  assign n8049 = ~\A[585]  & ~n8047 ;
  assign n8050 = ~n8048 & ~n8049 ;
  assign n8051 = ~\A[586]  & ~\A[587]  ;
  assign n8052 = ~n8044 & ~n8051 ;
  assign n8053 = \A[588]  & n8052 ;
  assign n8054 = ~\A[588]  & ~n8052 ;
  assign n8055 = ~n8053 & ~n8054 ;
  assign n8056 = n8050 & n8055 ;
  assign n8057 = n8044 & n8056 ;
  assign n8058 = ~n8045 & ~n8048 ;
  assign n8059 = ~n8044 & ~n8053 ;
  assign n8060 = ~n8056 & n8059 ;
  assign n8061 = ~n8058 & ~n8060 ;
  assign n8062 = ~n8057 & ~n8061 ;
  assign n8063 = \A[592]  & \A[593]  ;
  assign n8064 = ~\A[592]  & ~\A[593]  ;
  assign n8065 = ~n8063 & ~n8064 ;
  assign n8066 = \A[594]  & n8065 ;
  assign n8067 = ~n8063 & ~n8066 ;
  assign n8068 = \A[589]  & \A[590]  ;
  assign n8069 = ~\A[589]  & ~\A[590]  ;
  assign n8070 = ~n8068 & ~n8069 ;
  assign n8071 = \A[591]  & n8070 ;
  assign n8072 = ~n8068 & ~n8071 ;
  assign n8073 = n8067 & n8072 ;
  assign n8074 = ~n8067 & ~n8072 ;
  assign n8075 = ~\A[591]  & ~n8070 ;
  assign n8076 = ~n8071 & ~n8075 ;
  assign n8077 = ~\A[594]  & ~n8065 ;
  assign n8078 = ~n8066 & ~n8077 ;
  assign n8079 = n8076 & n8078 ;
  assign n8080 = ~n8074 & ~n8079 ;
  assign n8081 = ~n8073 & ~n8080 ;
  assign n8082 = ~n8076 & ~n8078 ;
  assign n8083 = ~n8079 & ~n8082 ;
  assign n8084 = ~n8050 & ~n8055 ;
  assign n8085 = ~n8056 & ~n8084 ;
  assign n8086 = n8083 & n8085 ;
  assign n8087 = n8057 & ~n8058 ;
  assign n8088 = n8086 & ~n8087 ;
  assign n8089 = ~n8073 & ~n8074 ;
  assign n8090 = n8079 & ~n8089 ;
  assign n8091 = ~n8079 & n8089 ;
  assign n8092 = ~n8090 & ~n8091 ;
  assign n8093 = n8088 & ~n8092 ;
  assign n8094 = ~n8088 & n8092 ;
  assign n8095 = ~n8057 & ~n8060 ;
  assign n8096 = n8058 & ~n8095 ;
  assign n8097 = ~n8058 & n8095 ;
  assign n8098 = ~n8096 & ~n8097 ;
  assign n8099 = ~n8094 & n8098 ;
  assign n8100 = ~n8093 & ~n8099 ;
  assign n8101 = n8081 & ~n8100 ;
  assign n8102 = ~n8081 & n8100 ;
  assign n8103 = ~n8101 & ~n8102 ;
  assign n8104 = n8062 & n8103 ;
  assign n8105 = ~n8062 & ~n8103 ;
  assign n8106 = ~n8104 & ~n8105 ;
  assign n8107 = \A[598]  & \A[599]  ;
  assign n8108 = \A[595]  & \A[596]  ;
  assign n8109 = ~\A[595]  & ~\A[596]  ;
  assign n8110 = ~n8108 & ~n8109 ;
  assign n8111 = \A[597]  & n8110 ;
  assign n8112 = ~\A[597]  & ~n8110 ;
  assign n8113 = ~n8111 & ~n8112 ;
  assign n8114 = ~\A[598]  & ~\A[599]  ;
  assign n8115 = ~n8107 & ~n8114 ;
  assign n8116 = \A[600]  & n8115 ;
  assign n8117 = ~\A[600]  & ~n8115 ;
  assign n8118 = ~n8116 & ~n8117 ;
  assign n8119 = n8113 & n8118 ;
  assign n8120 = n8107 & n8119 ;
  assign n8121 = ~n8108 & ~n8111 ;
  assign n8122 = ~n8107 & ~n8116 ;
  assign n8123 = ~n8119 & n8122 ;
  assign n8124 = ~n8121 & ~n8123 ;
  assign n8125 = ~n8120 & ~n8124 ;
  assign n8126 = \A[604]  & \A[605]  ;
  assign n8127 = ~\A[604]  & ~\A[605]  ;
  assign n8128 = ~n8126 & ~n8127 ;
  assign n8129 = \A[606]  & n8128 ;
  assign n8130 = ~n8126 & ~n8129 ;
  assign n8131 = \A[601]  & \A[602]  ;
  assign n8132 = ~\A[601]  & ~\A[602]  ;
  assign n8133 = ~n8131 & ~n8132 ;
  assign n8134 = \A[603]  & n8133 ;
  assign n8135 = ~n8131 & ~n8134 ;
  assign n8136 = n8130 & n8135 ;
  assign n8137 = ~n8130 & ~n8135 ;
  assign n8138 = ~\A[603]  & ~n8133 ;
  assign n8139 = ~n8134 & ~n8138 ;
  assign n8140 = ~\A[606]  & ~n8128 ;
  assign n8141 = ~n8129 & ~n8140 ;
  assign n8142 = n8139 & n8141 ;
  assign n8143 = ~n8137 & ~n8142 ;
  assign n8144 = ~n8136 & ~n8143 ;
  assign n8145 = ~n8139 & ~n8141 ;
  assign n8146 = ~n8142 & ~n8145 ;
  assign n8147 = ~n8113 & ~n8118 ;
  assign n8148 = ~n8119 & ~n8147 ;
  assign n8149 = n8146 & n8148 ;
  assign n8150 = n8120 & ~n8121 ;
  assign n8151 = n8149 & ~n8150 ;
  assign n8152 = ~n8136 & ~n8137 ;
  assign n8153 = n8142 & ~n8152 ;
  assign n8154 = ~n8142 & n8152 ;
  assign n8155 = ~n8153 & ~n8154 ;
  assign n8156 = n8151 & ~n8155 ;
  assign n8157 = ~n8151 & n8155 ;
  assign n8158 = ~n8120 & ~n8123 ;
  assign n8159 = n8121 & ~n8158 ;
  assign n8160 = ~n8121 & n8158 ;
  assign n8161 = ~n8159 & ~n8160 ;
  assign n8162 = ~n8157 & n8161 ;
  assign n8163 = ~n8156 & ~n8162 ;
  assign n8164 = n8144 & ~n8163 ;
  assign n8165 = ~n8144 & n8163 ;
  assign n8166 = ~n8164 & ~n8165 ;
  assign n8167 = n8125 & n8166 ;
  assign n8168 = ~n8125 & ~n8166 ;
  assign n8169 = ~n8167 & ~n8168 ;
  assign n8170 = ~n8106 & ~n8169 ;
  assign n8171 = n8106 & n8169 ;
  assign n8172 = ~n8146 & ~n8148 ;
  assign n8173 = ~n8149 & ~n8172 ;
  assign n8174 = ~n8083 & ~n8085 ;
  assign n8175 = ~n8086 & ~n8174 ;
  assign n8176 = n8173 & n8175 ;
  assign n8177 = ~n8156 & ~n8157 ;
  assign n8178 = n8161 & n8177 ;
  assign n8179 = ~n8161 & ~n8177 ;
  assign n8180 = ~n8178 & ~n8179 ;
  assign n8181 = n8176 & n8180 ;
  assign n8182 = ~n8176 & ~n8180 ;
  assign n8183 = ~n8093 & ~n8094 ;
  assign n8184 = n8098 & n8183 ;
  assign n8185 = ~n8098 & ~n8183 ;
  assign n8186 = ~n8184 & ~n8185 ;
  assign n8187 = ~n8182 & n8186 ;
  assign n8188 = ~n8181 & ~n8187 ;
  assign n8189 = ~n8171 & ~n8188 ;
  assign n8190 = ~n8170 & ~n8189 ;
  assign n8191 = ~n8125 & ~n8165 ;
  assign n8192 = ~n8164 & ~n8191 ;
  assign n8193 = ~n8190 & ~n8192 ;
  assign n8194 = n8190 & n8192 ;
  assign n8195 = ~n8193 & ~n8194 ;
  assign n8196 = ~n8062 & ~n8102 ;
  assign n8197 = ~n8101 & ~n8196 ;
  assign n8198 = n8195 & ~n8197 ;
  assign n8199 = ~n8195 & n8197 ;
  assign n8200 = ~n8198 & ~n8199 ;
  assign n8201 = ~n8038 & ~n8039 ;
  assign n8202 = ~n8041 & n8201 ;
  assign n8203 = n8041 & ~n8201 ;
  assign n8204 = ~n8202 & ~n8203 ;
  assign n8205 = ~n8200 & ~n8204 ;
  assign n8206 = n8200 & n8204 ;
  assign n8207 = ~n8015 & ~n8016 ;
  assign n8208 = ~n8033 & n8207 ;
  assign n8209 = n8033 & ~n8207 ;
  assign n8210 = ~n8208 & ~n8209 ;
  assign n8211 = ~n8170 & ~n8171 ;
  assign n8212 = ~n8188 & n8211 ;
  assign n8213 = n8188 & ~n8211 ;
  assign n8214 = ~n8212 & ~n8213 ;
  assign n8215 = ~n8210 & ~n8214 ;
  assign n8216 = n8210 & n8214 ;
  assign n8217 = ~n8173 & ~n8175 ;
  assign n8218 = ~n8176 & ~n8217 ;
  assign n8219 = ~n8018 & ~n8020 ;
  assign n8220 = ~n8021 & ~n8219 ;
  assign n8221 = n8218 & n8220 ;
  assign n8222 = ~n8181 & ~n8182 ;
  assign n8223 = ~n8186 & n8222 ;
  assign n8224 = n8186 & ~n8222 ;
  assign n8225 = ~n8223 & ~n8224 ;
  assign n8226 = n8221 & ~n8225 ;
  assign n8227 = ~n8221 & n8225 ;
  assign n8228 = ~n8026 & ~n8027 ;
  assign n8229 = ~n8031 & n8228 ;
  assign n8230 = n8031 & ~n8228 ;
  assign n8231 = ~n8229 & ~n8230 ;
  assign n8232 = ~n8227 & ~n8231 ;
  assign n8233 = ~n8226 & ~n8232 ;
  assign n8234 = ~n8216 & n8233 ;
  assign n8235 = ~n8215 & ~n8234 ;
  assign n8236 = ~n8206 & ~n8235 ;
  assign n8237 = ~n8205 & ~n8236 ;
  assign n8238 = n8043 & ~n8237 ;
  assign n8239 = ~n8043 & n8237 ;
  assign n8240 = ~n8238 & ~n8239 ;
  assign n8241 = ~n8194 & ~n8197 ;
  assign n8242 = ~n8193 & ~n8241 ;
  assign n8243 = n8240 & n8242 ;
  assign n8244 = ~n8240 & ~n8242 ;
  assign n8245 = ~n8243 & ~n8244 ;
  assign n8246 = \A[634]  & \A[635]  ;
  assign n8247 = \A[631]  & \A[632]  ;
  assign n8248 = ~\A[631]  & ~\A[632]  ;
  assign n8249 = ~n8247 & ~n8248 ;
  assign n8250 = \A[633]  & n8249 ;
  assign n8251 = ~\A[633]  & ~n8249 ;
  assign n8252 = ~n8250 & ~n8251 ;
  assign n8253 = ~\A[634]  & ~\A[635]  ;
  assign n8254 = ~n8246 & ~n8253 ;
  assign n8255 = \A[636]  & n8254 ;
  assign n8256 = ~\A[636]  & ~n8254 ;
  assign n8257 = ~n8255 & ~n8256 ;
  assign n8258 = n8252 & n8257 ;
  assign n8259 = n8246 & n8258 ;
  assign n8260 = ~n8247 & ~n8250 ;
  assign n8261 = ~n8246 & ~n8255 ;
  assign n8262 = ~n8258 & n8261 ;
  assign n8263 = ~n8260 & ~n8262 ;
  assign n8264 = ~n8259 & ~n8263 ;
  assign n8265 = \A[640]  & \A[641]  ;
  assign n8266 = ~\A[640]  & ~\A[641]  ;
  assign n8267 = ~n8265 & ~n8266 ;
  assign n8268 = \A[642]  & n8267 ;
  assign n8269 = ~n8265 & ~n8268 ;
  assign n8270 = \A[637]  & \A[638]  ;
  assign n8271 = ~\A[637]  & ~\A[638]  ;
  assign n8272 = ~n8270 & ~n8271 ;
  assign n8273 = \A[639]  & n8272 ;
  assign n8274 = ~n8270 & ~n8273 ;
  assign n8275 = n8269 & n8274 ;
  assign n8276 = ~n8269 & ~n8274 ;
  assign n8277 = ~\A[639]  & ~n8272 ;
  assign n8278 = ~n8273 & ~n8277 ;
  assign n8279 = ~\A[642]  & ~n8267 ;
  assign n8280 = ~n8268 & ~n8279 ;
  assign n8281 = n8278 & n8280 ;
  assign n8282 = ~n8276 & ~n8281 ;
  assign n8283 = ~n8275 & ~n8282 ;
  assign n8284 = ~n8278 & ~n8280 ;
  assign n8285 = ~n8281 & ~n8284 ;
  assign n8286 = ~n8252 & ~n8257 ;
  assign n8287 = ~n8258 & ~n8286 ;
  assign n8288 = n8285 & n8287 ;
  assign n8289 = n8259 & ~n8260 ;
  assign n8290 = n8288 & ~n8289 ;
  assign n8291 = ~n8275 & ~n8276 ;
  assign n8292 = n8281 & ~n8291 ;
  assign n8293 = ~n8281 & n8291 ;
  assign n8294 = ~n8292 & ~n8293 ;
  assign n8295 = n8290 & ~n8294 ;
  assign n8296 = ~n8290 & n8294 ;
  assign n8297 = ~n8259 & ~n8262 ;
  assign n8298 = n8260 & ~n8297 ;
  assign n8299 = ~n8260 & n8297 ;
  assign n8300 = ~n8298 & ~n8299 ;
  assign n8301 = ~n8296 & n8300 ;
  assign n8302 = ~n8295 & ~n8301 ;
  assign n8303 = n8283 & ~n8302 ;
  assign n8304 = ~n8283 & n8302 ;
  assign n8305 = ~n8303 & ~n8304 ;
  assign n8306 = n8264 & n8305 ;
  assign n8307 = ~n8264 & ~n8305 ;
  assign n8308 = ~n8306 & ~n8307 ;
  assign n8309 = \A[646]  & \A[647]  ;
  assign n8310 = \A[643]  & \A[644]  ;
  assign n8311 = ~\A[643]  & ~\A[644]  ;
  assign n8312 = ~n8310 & ~n8311 ;
  assign n8313 = \A[645]  & n8312 ;
  assign n8314 = ~\A[645]  & ~n8312 ;
  assign n8315 = ~n8313 & ~n8314 ;
  assign n8316 = ~\A[646]  & ~\A[647]  ;
  assign n8317 = ~n8309 & ~n8316 ;
  assign n8318 = \A[648]  & n8317 ;
  assign n8319 = ~\A[648]  & ~n8317 ;
  assign n8320 = ~n8318 & ~n8319 ;
  assign n8321 = n8315 & n8320 ;
  assign n8322 = n8309 & n8321 ;
  assign n8323 = ~n8310 & ~n8313 ;
  assign n8324 = ~n8309 & ~n8318 ;
  assign n8325 = ~n8321 & n8324 ;
  assign n8326 = ~n8323 & ~n8325 ;
  assign n8327 = ~n8322 & ~n8326 ;
  assign n8328 = \A[652]  & \A[653]  ;
  assign n8329 = ~\A[652]  & ~\A[653]  ;
  assign n8330 = ~n8328 & ~n8329 ;
  assign n8331 = \A[654]  & n8330 ;
  assign n8332 = ~n8328 & ~n8331 ;
  assign n8333 = \A[649]  & \A[650]  ;
  assign n8334 = ~\A[649]  & ~\A[650]  ;
  assign n8335 = ~n8333 & ~n8334 ;
  assign n8336 = \A[651]  & n8335 ;
  assign n8337 = ~n8333 & ~n8336 ;
  assign n8338 = n8332 & n8337 ;
  assign n8339 = ~n8332 & ~n8337 ;
  assign n8340 = ~\A[651]  & ~n8335 ;
  assign n8341 = ~n8336 & ~n8340 ;
  assign n8342 = ~\A[654]  & ~n8330 ;
  assign n8343 = ~n8331 & ~n8342 ;
  assign n8344 = n8341 & n8343 ;
  assign n8345 = ~n8339 & ~n8344 ;
  assign n8346 = ~n8338 & ~n8345 ;
  assign n8347 = ~n8341 & ~n8343 ;
  assign n8348 = ~n8344 & ~n8347 ;
  assign n8349 = ~n8315 & ~n8320 ;
  assign n8350 = ~n8321 & ~n8349 ;
  assign n8351 = n8348 & n8350 ;
  assign n8352 = n8322 & ~n8323 ;
  assign n8353 = n8351 & ~n8352 ;
  assign n8354 = ~n8338 & ~n8339 ;
  assign n8355 = n8344 & ~n8354 ;
  assign n8356 = ~n8344 & n8354 ;
  assign n8357 = ~n8355 & ~n8356 ;
  assign n8358 = n8353 & ~n8357 ;
  assign n8359 = ~n8353 & n8357 ;
  assign n8360 = ~n8322 & ~n8325 ;
  assign n8361 = n8323 & ~n8360 ;
  assign n8362 = ~n8323 & n8360 ;
  assign n8363 = ~n8361 & ~n8362 ;
  assign n8364 = ~n8359 & n8363 ;
  assign n8365 = ~n8358 & ~n8364 ;
  assign n8366 = n8346 & ~n8365 ;
  assign n8367 = ~n8346 & n8365 ;
  assign n8368 = ~n8366 & ~n8367 ;
  assign n8369 = n8327 & n8368 ;
  assign n8370 = ~n8327 & ~n8368 ;
  assign n8371 = ~n8369 & ~n8370 ;
  assign n8372 = ~n8308 & ~n8371 ;
  assign n8373 = n8308 & n8371 ;
  assign n8374 = ~n8348 & ~n8350 ;
  assign n8375 = ~n8351 & ~n8374 ;
  assign n8376 = ~n8285 & ~n8287 ;
  assign n8377 = ~n8288 & ~n8376 ;
  assign n8378 = n8375 & n8377 ;
  assign n8379 = ~n8358 & ~n8359 ;
  assign n8380 = n8363 & n8379 ;
  assign n8381 = ~n8363 & ~n8379 ;
  assign n8382 = ~n8380 & ~n8381 ;
  assign n8383 = n8378 & n8382 ;
  assign n8384 = ~n8378 & ~n8382 ;
  assign n8385 = ~n8295 & ~n8296 ;
  assign n8386 = n8300 & n8385 ;
  assign n8387 = ~n8300 & ~n8385 ;
  assign n8388 = ~n8386 & ~n8387 ;
  assign n8389 = ~n8384 & n8388 ;
  assign n8390 = ~n8383 & ~n8389 ;
  assign n8391 = ~n8373 & ~n8390 ;
  assign n8392 = ~n8372 & ~n8391 ;
  assign n8393 = ~n8327 & ~n8367 ;
  assign n8394 = ~n8366 & ~n8393 ;
  assign n8395 = ~n8392 & ~n8394 ;
  assign n8396 = n8392 & n8394 ;
  assign n8397 = ~n8264 & ~n8304 ;
  assign n8398 = ~n8303 & ~n8397 ;
  assign n8399 = ~n8396 & ~n8398 ;
  assign n8400 = ~n8395 & ~n8399 ;
  assign n8401 = ~n8395 & ~n8396 ;
  assign n8402 = ~n8398 & n8401 ;
  assign n8403 = n8398 & ~n8401 ;
  assign n8404 = ~n8402 & ~n8403 ;
  assign n8405 = \A[610]  & \A[611]  ;
  assign n8406 = \A[607]  & \A[608]  ;
  assign n8407 = ~\A[607]  & ~\A[608]  ;
  assign n8408 = ~n8406 & ~n8407 ;
  assign n8409 = \A[609]  & n8408 ;
  assign n8410 = ~\A[609]  & ~n8408 ;
  assign n8411 = ~n8409 & ~n8410 ;
  assign n8412 = ~\A[610]  & ~\A[611]  ;
  assign n8413 = ~n8405 & ~n8412 ;
  assign n8414 = \A[612]  & n8413 ;
  assign n8415 = ~\A[612]  & ~n8413 ;
  assign n8416 = ~n8414 & ~n8415 ;
  assign n8417 = n8411 & n8416 ;
  assign n8418 = n8405 & n8417 ;
  assign n8419 = ~n8406 & ~n8409 ;
  assign n8420 = ~n8405 & ~n8414 ;
  assign n8421 = ~n8417 & n8420 ;
  assign n8422 = ~n8419 & ~n8421 ;
  assign n8423 = ~n8418 & ~n8422 ;
  assign n8424 = \A[616]  & \A[617]  ;
  assign n8425 = ~\A[616]  & ~\A[617]  ;
  assign n8426 = ~n8424 & ~n8425 ;
  assign n8427 = \A[618]  & n8426 ;
  assign n8428 = ~n8424 & ~n8427 ;
  assign n8429 = \A[613]  & \A[614]  ;
  assign n8430 = ~\A[613]  & ~\A[614]  ;
  assign n8431 = ~n8429 & ~n8430 ;
  assign n8432 = \A[615]  & n8431 ;
  assign n8433 = ~n8429 & ~n8432 ;
  assign n8434 = n8428 & n8433 ;
  assign n8435 = ~n8428 & ~n8433 ;
  assign n8436 = ~\A[615]  & ~n8431 ;
  assign n8437 = ~n8432 & ~n8436 ;
  assign n8438 = ~\A[618]  & ~n8426 ;
  assign n8439 = ~n8427 & ~n8438 ;
  assign n8440 = n8437 & n8439 ;
  assign n8441 = ~n8435 & ~n8440 ;
  assign n8442 = ~n8434 & ~n8441 ;
  assign n8443 = ~n8437 & ~n8439 ;
  assign n8444 = ~n8440 & ~n8443 ;
  assign n8445 = ~n8411 & ~n8416 ;
  assign n8446 = ~n8417 & ~n8445 ;
  assign n8447 = n8444 & n8446 ;
  assign n8448 = n8418 & ~n8419 ;
  assign n8449 = n8447 & ~n8448 ;
  assign n8450 = ~n8434 & ~n8435 ;
  assign n8451 = n8440 & ~n8450 ;
  assign n8452 = ~n8440 & n8450 ;
  assign n8453 = ~n8451 & ~n8452 ;
  assign n8454 = n8449 & ~n8453 ;
  assign n8455 = ~n8449 & n8453 ;
  assign n8456 = ~n8418 & ~n8421 ;
  assign n8457 = n8419 & ~n8456 ;
  assign n8458 = ~n8419 & n8456 ;
  assign n8459 = ~n8457 & ~n8458 ;
  assign n8460 = ~n8455 & n8459 ;
  assign n8461 = ~n8454 & ~n8460 ;
  assign n8462 = n8442 & ~n8461 ;
  assign n8463 = ~n8442 & n8461 ;
  assign n8464 = ~n8462 & ~n8463 ;
  assign n8465 = n8423 & n8464 ;
  assign n8466 = ~n8423 & ~n8464 ;
  assign n8467 = ~n8465 & ~n8466 ;
  assign n8468 = \A[622]  & \A[623]  ;
  assign n8469 = \A[619]  & \A[620]  ;
  assign n8470 = ~\A[619]  & ~\A[620]  ;
  assign n8471 = ~n8469 & ~n8470 ;
  assign n8472 = \A[621]  & n8471 ;
  assign n8473 = ~\A[621]  & ~n8471 ;
  assign n8474 = ~n8472 & ~n8473 ;
  assign n8475 = ~\A[622]  & ~\A[623]  ;
  assign n8476 = ~n8468 & ~n8475 ;
  assign n8477 = \A[624]  & n8476 ;
  assign n8478 = ~\A[624]  & ~n8476 ;
  assign n8479 = ~n8477 & ~n8478 ;
  assign n8480 = n8474 & n8479 ;
  assign n8481 = n8468 & n8480 ;
  assign n8482 = ~n8469 & ~n8472 ;
  assign n8483 = ~n8468 & ~n8477 ;
  assign n8484 = ~n8480 & n8483 ;
  assign n8485 = ~n8482 & ~n8484 ;
  assign n8486 = ~n8481 & ~n8485 ;
  assign n8487 = \A[628]  & \A[629]  ;
  assign n8488 = ~\A[628]  & ~\A[629]  ;
  assign n8489 = ~n8487 & ~n8488 ;
  assign n8490 = \A[630]  & n8489 ;
  assign n8491 = ~n8487 & ~n8490 ;
  assign n8492 = \A[625]  & \A[626]  ;
  assign n8493 = ~\A[625]  & ~\A[626]  ;
  assign n8494 = ~n8492 & ~n8493 ;
  assign n8495 = \A[627]  & n8494 ;
  assign n8496 = ~n8492 & ~n8495 ;
  assign n8497 = n8491 & n8496 ;
  assign n8498 = ~n8491 & ~n8496 ;
  assign n8499 = ~\A[627]  & ~n8494 ;
  assign n8500 = ~n8495 & ~n8499 ;
  assign n8501 = ~\A[630]  & ~n8489 ;
  assign n8502 = ~n8490 & ~n8501 ;
  assign n8503 = n8500 & n8502 ;
  assign n8504 = ~n8498 & ~n8503 ;
  assign n8505 = ~n8497 & ~n8504 ;
  assign n8506 = ~n8500 & ~n8502 ;
  assign n8507 = ~n8503 & ~n8506 ;
  assign n8508 = ~n8474 & ~n8479 ;
  assign n8509 = ~n8480 & ~n8508 ;
  assign n8510 = n8507 & n8509 ;
  assign n8511 = n8481 & ~n8482 ;
  assign n8512 = n8510 & ~n8511 ;
  assign n8513 = ~n8497 & ~n8498 ;
  assign n8514 = n8503 & ~n8513 ;
  assign n8515 = ~n8503 & n8513 ;
  assign n8516 = ~n8514 & ~n8515 ;
  assign n8517 = n8512 & ~n8516 ;
  assign n8518 = ~n8512 & n8516 ;
  assign n8519 = ~n8481 & ~n8484 ;
  assign n8520 = n8482 & ~n8519 ;
  assign n8521 = ~n8482 & n8519 ;
  assign n8522 = ~n8520 & ~n8521 ;
  assign n8523 = ~n8518 & n8522 ;
  assign n8524 = ~n8517 & ~n8523 ;
  assign n8525 = n8505 & ~n8524 ;
  assign n8526 = ~n8505 & n8524 ;
  assign n8527 = ~n8525 & ~n8526 ;
  assign n8528 = n8486 & n8527 ;
  assign n8529 = ~n8486 & ~n8527 ;
  assign n8530 = ~n8528 & ~n8529 ;
  assign n8531 = ~n8467 & ~n8530 ;
  assign n8532 = n8467 & n8530 ;
  assign n8533 = ~n8507 & ~n8509 ;
  assign n8534 = ~n8510 & ~n8533 ;
  assign n8535 = ~n8444 & ~n8446 ;
  assign n8536 = ~n8447 & ~n8535 ;
  assign n8537 = n8534 & n8536 ;
  assign n8538 = ~n8517 & ~n8518 ;
  assign n8539 = n8522 & n8538 ;
  assign n8540 = ~n8522 & ~n8538 ;
  assign n8541 = ~n8539 & ~n8540 ;
  assign n8542 = n8537 & n8541 ;
  assign n8543 = ~n8537 & ~n8541 ;
  assign n8544 = ~n8454 & ~n8455 ;
  assign n8545 = n8459 & n8544 ;
  assign n8546 = ~n8459 & ~n8544 ;
  assign n8547 = ~n8545 & ~n8546 ;
  assign n8548 = ~n8543 & n8547 ;
  assign n8549 = ~n8542 & ~n8548 ;
  assign n8550 = ~n8532 & ~n8549 ;
  assign n8551 = ~n8531 & ~n8550 ;
  assign n8552 = ~n8486 & ~n8526 ;
  assign n8553 = ~n8525 & ~n8552 ;
  assign n8554 = ~n8551 & ~n8553 ;
  assign n8555 = n8551 & n8553 ;
  assign n8556 = ~n8554 & ~n8555 ;
  assign n8557 = ~n8423 & ~n8463 ;
  assign n8558 = ~n8462 & ~n8557 ;
  assign n8559 = n8556 & ~n8558 ;
  assign n8560 = ~n8556 & n8558 ;
  assign n8561 = ~n8559 & ~n8560 ;
  assign n8562 = ~n8404 & ~n8561 ;
  assign n8563 = n8404 & n8561 ;
  assign n8564 = ~n8531 & ~n8532 ;
  assign n8565 = ~n8549 & n8564 ;
  assign n8566 = n8549 & ~n8564 ;
  assign n8567 = ~n8565 & ~n8566 ;
  assign n8568 = ~n8372 & ~n8373 ;
  assign n8569 = ~n8390 & n8568 ;
  assign n8570 = n8390 & ~n8568 ;
  assign n8571 = ~n8569 & ~n8570 ;
  assign n8572 = ~n8567 & ~n8571 ;
  assign n8573 = n8567 & n8571 ;
  assign n8574 = ~n8375 & ~n8377 ;
  assign n8575 = ~n8378 & ~n8574 ;
  assign n8576 = ~n8534 & ~n8536 ;
  assign n8577 = ~n8537 & ~n8576 ;
  assign n8578 = n8575 & n8577 ;
  assign n8579 = ~n8383 & ~n8384 ;
  assign n8580 = ~n8388 & n8579 ;
  assign n8581 = n8388 & ~n8579 ;
  assign n8582 = ~n8580 & ~n8581 ;
  assign n8583 = n8578 & ~n8582 ;
  assign n8584 = ~n8578 & n8582 ;
  assign n8585 = ~n8542 & ~n8543 ;
  assign n8586 = ~n8547 & n8585 ;
  assign n8587 = n8547 & ~n8585 ;
  assign n8588 = ~n8586 & ~n8587 ;
  assign n8589 = ~n8584 & ~n8588 ;
  assign n8590 = ~n8583 & ~n8589 ;
  assign n8591 = ~n8573 & n8590 ;
  assign n8592 = ~n8572 & ~n8591 ;
  assign n8593 = ~n8563 & ~n8592 ;
  assign n8594 = ~n8562 & ~n8593 ;
  assign n8595 = n8400 & ~n8594 ;
  assign n8596 = ~n8400 & n8594 ;
  assign n8597 = ~n8595 & ~n8596 ;
  assign n8598 = ~n8555 & ~n8558 ;
  assign n8599 = ~n8554 & ~n8598 ;
  assign n8600 = n8597 & n8599 ;
  assign n8601 = ~n8597 & ~n8599 ;
  assign n8602 = ~n8600 & ~n8601 ;
  assign n8603 = ~n8245 & ~n8602 ;
  assign n8604 = n8245 & n8602 ;
  assign n8605 = ~n8562 & ~n8563 ;
  assign n8606 = ~n8592 & n8605 ;
  assign n8607 = n8592 & ~n8605 ;
  assign n8608 = ~n8606 & ~n8607 ;
  assign n8609 = ~n8205 & ~n8206 ;
  assign n8610 = ~n8235 & n8609 ;
  assign n8611 = n8235 & ~n8609 ;
  assign n8612 = ~n8610 & ~n8611 ;
  assign n8613 = ~n8608 & ~n8612 ;
  assign n8614 = n8608 & n8612 ;
  assign n8615 = ~n8215 & ~n8216 ;
  assign n8616 = ~n8233 & n8615 ;
  assign n8617 = n8233 & ~n8615 ;
  assign n8618 = ~n8616 & ~n8617 ;
  assign n8619 = ~n8572 & ~n8573 ;
  assign n8620 = ~n8590 & n8619 ;
  assign n8621 = n8590 & ~n8619 ;
  assign n8622 = ~n8620 & ~n8621 ;
  assign n8623 = ~n8618 & ~n8622 ;
  assign n8624 = n8618 & n8622 ;
  assign n8625 = ~n8575 & ~n8577 ;
  assign n8626 = ~n8578 & ~n8625 ;
  assign n8627 = ~n8218 & ~n8220 ;
  assign n8628 = ~n8221 & ~n8627 ;
  assign n8629 = n8626 & n8628 ;
  assign n8630 = ~n8583 & ~n8584 ;
  assign n8631 = ~n8588 & n8630 ;
  assign n8632 = n8588 & ~n8630 ;
  assign n8633 = ~n8631 & ~n8632 ;
  assign n8634 = n8629 & n8633 ;
  assign n8635 = ~n8629 & ~n8633 ;
  assign n8636 = ~n8226 & ~n8227 ;
  assign n8637 = ~n8231 & n8636 ;
  assign n8638 = n8231 & ~n8636 ;
  assign n8639 = ~n8637 & ~n8638 ;
  assign n8640 = ~n8635 & n8639 ;
  assign n8641 = ~n8634 & ~n8640 ;
  assign n8642 = ~n8624 & n8641 ;
  assign n8643 = ~n8623 & ~n8642 ;
  assign n8644 = ~n8614 & n8643 ;
  assign n8645 = ~n8613 & ~n8644 ;
  assign n8646 = ~n8604 & ~n8645 ;
  assign n8647 = ~n8603 & ~n8646 ;
  assign n8648 = ~n8239 & n8242 ;
  assign n8649 = ~n8238 & ~n8648 ;
  assign n8650 = n8647 & ~n8649 ;
  assign n8651 = ~n8647 & n8649 ;
  assign n8652 = ~n8596 & n8599 ;
  assign n8653 = ~n8595 & ~n8652 ;
  assign n8654 = ~n8651 & ~n8653 ;
  assign n8655 = ~n8650 & ~n8654 ;
  assign n8656 = \A[466]  & \A[467]  ;
  assign n8657 = ~\A[466]  & ~\A[467]  ;
  assign n8658 = ~n8656 & ~n8657 ;
  assign n8659 = \A[468]  & n8658 ;
  assign n8660 = ~\A[468]  & ~n8658 ;
  assign n8661 = ~n8659 & ~n8660 ;
  assign n8662 = \A[463]  & \A[464]  ;
  assign n8663 = ~\A[463]  & ~\A[464]  ;
  assign n8664 = ~n8662 & ~n8663 ;
  assign n8665 = \A[465]  & n8664 ;
  assign n8666 = ~\A[465]  & ~n8664 ;
  assign n8667 = ~n8665 & ~n8666 ;
  assign n8668 = n8661 & n8667 ;
  assign n8669 = n8656 & n8668 ;
  assign n8670 = ~n8662 & ~n8665 ;
  assign n8671 = ~n8656 & ~n8659 ;
  assign n8672 = ~n8668 & n8671 ;
  assign n8673 = ~n8670 & ~n8672 ;
  assign n8674 = ~n8669 & ~n8673 ;
  assign n8675 = \A[472]  & \A[473]  ;
  assign n8676 = ~\A[472]  & ~\A[473]  ;
  assign n8677 = ~n8675 & ~n8676 ;
  assign n8678 = \A[474]  & n8677 ;
  assign n8679 = ~n8675 & ~n8678 ;
  assign n8680 = \A[469]  & \A[470]  ;
  assign n8681 = ~\A[469]  & ~\A[470]  ;
  assign n8682 = ~n8680 & ~n8681 ;
  assign n8683 = \A[471]  & n8682 ;
  assign n8684 = ~n8680 & ~n8683 ;
  assign n8685 = n8679 & n8684 ;
  assign n8686 = ~n8679 & ~n8684 ;
  assign n8687 = ~\A[471]  & ~n8682 ;
  assign n8688 = ~n8683 & ~n8687 ;
  assign n8689 = ~\A[474]  & ~n8677 ;
  assign n8690 = ~n8678 & ~n8689 ;
  assign n8691 = n8688 & n8690 ;
  assign n8692 = ~n8686 & ~n8691 ;
  assign n8693 = ~n8685 & ~n8692 ;
  assign n8694 = ~n8688 & ~n8690 ;
  assign n8695 = ~n8691 & ~n8694 ;
  assign n8696 = ~n8661 & ~n8667 ;
  assign n8697 = ~n8668 & ~n8696 ;
  assign n8698 = n8695 & n8697 ;
  assign n8699 = n8669 & ~n8670 ;
  assign n8700 = n8698 & ~n8699 ;
  assign n8701 = ~n8685 & ~n8686 ;
  assign n8702 = n8691 & ~n8701 ;
  assign n8703 = ~n8691 & n8701 ;
  assign n8704 = ~n8702 & ~n8703 ;
  assign n8705 = n8700 & ~n8704 ;
  assign n8706 = ~n8700 & n8704 ;
  assign n8707 = ~n8669 & ~n8672 ;
  assign n8708 = n8670 & ~n8707 ;
  assign n8709 = ~n8670 & n8707 ;
  assign n8710 = ~n8708 & ~n8709 ;
  assign n8711 = ~n8706 & n8710 ;
  assign n8712 = ~n8705 & ~n8711 ;
  assign n8713 = n8693 & ~n8712 ;
  assign n8714 = ~n8693 & n8712 ;
  assign n8715 = ~n8713 & ~n8714 ;
  assign n8716 = n8674 & n8715 ;
  assign n8717 = ~n8674 & ~n8715 ;
  assign n8718 = ~n8716 & ~n8717 ;
  assign n8719 = \A[478]  & \A[479]  ;
  assign n8720 = \A[475]  & \A[476]  ;
  assign n8721 = ~\A[475]  & ~\A[476]  ;
  assign n8722 = ~n8720 & ~n8721 ;
  assign n8723 = \A[477]  & n8722 ;
  assign n8724 = ~\A[477]  & ~n8722 ;
  assign n8725 = ~n8723 & ~n8724 ;
  assign n8726 = ~\A[478]  & ~\A[479]  ;
  assign n8727 = ~n8719 & ~n8726 ;
  assign n8728 = \A[480]  & n8727 ;
  assign n8729 = ~\A[480]  & ~n8727 ;
  assign n8730 = ~n8728 & ~n8729 ;
  assign n8731 = n8725 & n8730 ;
  assign n8732 = n8719 & n8731 ;
  assign n8733 = ~n8720 & ~n8723 ;
  assign n8734 = ~n8719 & ~n8728 ;
  assign n8735 = ~n8731 & n8734 ;
  assign n8736 = ~n8733 & ~n8735 ;
  assign n8737 = ~n8732 & ~n8736 ;
  assign n8738 = \A[484]  & \A[485]  ;
  assign n8739 = ~\A[484]  & ~\A[485]  ;
  assign n8740 = ~n8738 & ~n8739 ;
  assign n8741 = \A[486]  & n8740 ;
  assign n8742 = ~n8738 & ~n8741 ;
  assign n8743 = \A[481]  & \A[482]  ;
  assign n8744 = ~\A[481]  & ~\A[482]  ;
  assign n8745 = ~n8743 & ~n8744 ;
  assign n8746 = \A[483]  & n8745 ;
  assign n8747 = ~n8743 & ~n8746 ;
  assign n8748 = n8742 & n8747 ;
  assign n8749 = ~n8742 & ~n8747 ;
  assign n8750 = ~\A[483]  & ~n8745 ;
  assign n8751 = ~n8746 & ~n8750 ;
  assign n8752 = ~\A[486]  & ~n8740 ;
  assign n8753 = ~n8741 & ~n8752 ;
  assign n8754 = n8751 & n8753 ;
  assign n8755 = ~n8749 & ~n8754 ;
  assign n8756 = ~n8748 & ~n8755 ;
  assign n8757 = ~n8751 & ~n8753 ;
  assign n8758 = ~n8754 & ~n8757 ;
  assign n8759 = ~n8725 & ~n8730 ;
  assign n8760 = ~n8731 & ~n8759 ;
  assign n8761 = n8758 & n8760 ;
  assign n8762 = n8732 & ~n8733 ;
  assign n8763 = n8761 & ~n8762 ;
  assign n8764 = ~n8748 & ~n8749 ;
  assign n8765 = n8754 & ~n8764 ;
  assign n8766 = ~n8754 & n8764 ;
  assign n8767 = ~n8765 & ~n8766 ;
  assign n8768 = n8763 & ~n8767 ;
  assign n8769 = ~n8763 & n8767 ;
  assign n8770 = ~n8732 & ~n8735 ;
  assign n8771 = n8733 & ~n8770 ;
  assign n8772 = ~n8733 & n8770 ;
  assign n8773 = ~n8771 & ~n8772 ;
  assign n8774 = ~n8769 & n8773 ;
  assign n8775 = ~n8768 & ~n8774 ;
  assign n8776 = n8756 & ~n8775 ;
  assign n8777 = ~n8756 & n8775 ;
  assign n8778 = ~n8776 & ~n8777 ;
  assign n8779 = n8737 & n8778 ;
  assign n8780 = ~n8737 & ~n8778 ;
  assign n8781 = ~n8779 & ~n8780 ;
  assign n8782 = ~n8718 & ~n8781 ;
  assign n8783 = n8718 & n8781 ;
  assign n8784 = ~n8695 & ~n8697 ;
  assign n8785 = ~n8698 & ~n8784 ;
  assign n8786 = ~n8758 & ~n8760 ;
  assign n8787 = ~n8761 & ~n8786 ;
  assign n8788 = n8785 & n8787 ;
  assign n8789 = ~n8768 & ~n8769 ;
  assign n8790 = n8773 & n8789 ;
  assign n8791 = ~n8773 & ~n8789 ;
  assign n8792 = ~n8790 & ~n8791 ;
  assign n8793 = n8788 & n8792 ;
  assign n8794 = ~n8788 & ~n8792 ;
  assign n8795 = ~n8705 & ~n8706 ;
  assign n8796 = n8710 & n8795 ;
  assign n8797 = ~n8710 & ~n8795 ;
  assign n8798 = ~n8796 & ~n8797 ;
  assign n8799 = ~n8794 & n8798 ;
  assign n8800 = ~n8793 & ~n8799 ;
  assign n8801 = ~n8783 & ~n8800 ;
  assign n8802 = ~n8782 & ~n8801 ;
  assign n8803 = ~n8737 & ~n8777 ;
  assign n8804 = ~n8776 & ~n8803 ;
  assign n8805 = ~n8802 & ~n8804 ;
  assign n8806 = n8802 & n8804 ;
  assign n8807 = ~n8674 & ~n8714 ;
  assign n8808 = ~n8713 & ~n8807 ;
  assign n8809 = ~n8806 & ~n8808 ;
  assign n8810 = ~n8805 & ~n8809 ;
  assign n8811 = \A[490]  & \A[491]  ;
  assign n8812 = \A[487]  & \A[488]  ;
  assign n8813 = ~\A[487]  & ~\A[488]  ;
  assign n8814 = ~n8812 & ~n8813 ;
  assign n8815 = \A[489]  & n8814 ;
  assign n8816 = ~\A[489]  & ~n8814 ;
  assign n8817 = ~n8815 & ~n8816 ;
  assign n8818 = ~\A[490]  & ~\A[491]  ;
  assign n8819 = ~n8811 & ~n8818 ;
  assign n8820 = \A[492]  & n8819 ;
  assign n8821 = ~\A[492]  & ~n8819 ;
  assign n8822 = ~n8820 & ~n8821 ;
  assign n8823 = n8817 & n8822 ;
  assign n8824 = n8811 & n8823 ;
  assign n8825 = ~n8812 & ~n8815 ;
  assign n8826 = ~n8811 & ~n8820 ;
  assign n8827 = ~n8823 & n8826 ;
  assign n8828 = ~n8825 & ~n8827 ;
  assign n8829 = ~n8824 & ~n8828 ;
  assign n8830 = \A[496]  & \A[497]  ;
  assign n8831 = ~\A[496]  & ~\A[497]  ;
  assign n8832 = ~n8830 & ~n8831 ;
  assign n8833 = \A[498]  & n8832 ;
  assign n8834 = ~n8830 & ~n8833 ;
  assign n8835 = \A[493]  & \A[494]  ;
  assign n8836 = ~\A[493]  & ~\A[494]  ;
  assign n8837 = ~n8835 & ~n8836 ;
  assign n8838 = \A[495]  & n8837 ;
  assign n8839 = ~n8835 & ~n8838 ;
  assign n8840 = n8834 & n8839 ;
  assign n8841 = ~n8834 & ~n8839 ;
  assign n8842 = ~\A[495]  & ~n8837 ;
  assign n8843 = ~n8838 & ~n8842 ;
  assign n8844 = ~\A[498]  & ~n8832 ;
  assign n8845 = ~n8833 & ~n8844 ;
  assign n8846 = n8843 & n8845 ;
  assign n8847 = ~n8841 & ~n8846 ;
  assign n8848 = ~n8840 & ~n8847 ;
  assign n8849 = ~n8843 & ~n8845 ;
  assign n8850 = ~n8846 & ~n8849 ;
  assign n8851 = ~n8817 & ~n8822 ;
  assign n8852 = ~n8823 & ~n8851 ;
  assign n8853 = n8850 & n8852 ;
  assign n8854 = n8824 & ~n8825 ;
  assign n8855 = n8853 & ~n8854 ;
  assign n8856 = ~n8840 & ~n8841 ;
  assign n8857 = n8846 & ~n8856 ;
  assign n8858 = ~n8846 & n8856 ;
  assign n8859 = ~n8857 & ~n8858 ;
  assign n8860 = n8855 & ~n8859 ;
  assign n8861 = ~n8855 & n8859 ;
  assign n8862 = ~n8824 & ~n8827 ;
  assign n8863 = n8825 & ~n8862 ;
  assign n8864 = ~n8825 & n8862 ;
  assign n8865 = ~n8863 & ~n8864 ;
  assign n8866 = ~n8861 & n8865 ;
  assign n8867 = ~n8860 & ~n8866 ;
  assign n8868 = n8848 & ~n8867 ;
  assign n8869 = ~n8848 & n8867 ;
  assign n8870 = ~n8868 & ~n8869 ;
  assign n8871 = n8829 & n8870 ;
  assign n8872 = ~n8829 & ~n8870 ;
  assign n8873 = ~n8871 & ~n8872 ;
  assign n8874 = \A[502]  & \A[503]  ;
  assign n8875 = \A[499]  & \A[500]  ;
  assign n8876 = ~\A[499]  & ~\A[500]  ;
  assign n8877 = ~n8875 & ~n8876 ;
  assign n8878 = \A[501]  & n8877 ;
  assign n8879 = ~\A[501]  & ~n8877 ;
  assign n8880 = ~n8878 & ~n8879 ;
  assign n8881 = ~\A[502]  & ~\A[503]  ;
  assign n8882 = ~n8874 & ~n8881 ;
  assign n8883 = \A[504]  & n8882 ;
  assign n8884 = ~\A[504]  & ~n8882 ;
  assign n8885 = ~n8883 & ~n8884 ;
  assign n8886 = n8880 & n8885 ;
  assign n8887 = n8874 & n8886 ;
  assign n8888 = ~n8875 & ~n8878 ;
  assign n8889 = ~n8874 & ~n8883 ;
  assign n8890 = ~n8886 & n8889 ;
  assign n8891 = ~n8888 & ~n8890 ;
  assign n8892 = ~n8887 & ~n8891 ;
  assign n8893 = \A[508]  & \A[509]  ;
  assign n8894 = ~\A[508]  & ~\A[509]  ;
  assign n8895 = ~n8893 & ~n8894 ;
  assign n8896 = \A[510]  & n8895 ;
  assign n8897 = ~n8893 & ~n8896 ;
  assign n8898 = \A[505]  & \A[506]  ;
  assign n8899 = ~\A[505]  & ~\A[506]  ;
  assign n8900 = ~n8898 & ~n8899 ;
  assign n8901 = \A[507]  & n8900 ;
  assign n8902 = ~n8898 & ~n8901 ;
  assign n8903 = n8897 & n8902 ;
  assign n8904 = ~n8897 & ~n8902 ;
  assign n8905 = ~\A[507]  & ~n8900 ;
  assign n8906 = ~n8901 & ~n8905 ;
  assign n8907 = ~\A[510]  & ~n8895 ;
  assign n8908 = ~n8896 & ~n8907 ;
  assign n8909 = n8906 & n8908 ;
  assign n8910 = ~n8904 & ~n8909 ;
  assign n8911 = ~n8903 & ~n8910 ;
  assign n8912 = ~n8906 & ~n8908 ;
  assign n8913 = ~n8909 & ~n8912 ;
  assign n8914 = ~n8880 & ~n8885 ;
  assign n8915 = ~n8886 & ~n8914 ;
  assign n8916 = n8913 & n8915 ;
  assign n8917 = n8887 & ~n8888 ;
  assign n8918 = n8916 & ~n8917 ;
  assign n8919 = ~n8903 & ~n8904 ;
  assign n8920 = n8909 & ~n8919 ;
  assign n8921 = ~n8909 & n8919 ;
  assign n8922 = ~n8920 & ~n8921 ;
  assign n8923 = n8918 & ~n8922 ;
  assign n8924 = ~n8918 & n8922 ;
  assign n8925 = ~n8887 & ~n8890 ;
  assign n8926 = n8888 & ~n8925 ;
  assign n8927 = ~n8888 & n8925 ;
  assign n8928 = ~n8926 & ~n8927 ;
  assign n8929 = ~n8924 & n8928 ;
  assign n8930 = ~n8923 & ~n8929 ;
  assign n8931 = n8911 & ~n8930 ;
  assign n8932 = ~n8911 & n8930 ;
  assign n8933 = ~n8931 & ~n8932 ;
  assign n8934 = n8892 & n8933 ;
  assign n8935 = ~n8892 & ~n8933 ;
  assign n8936 = ~n8934 & ~n8935 ;
  assign n8937 = ~n8873 & ~n8936 ;
  assign n8938 = n8873 & n8936 ;
  assign n8939 = ~n8913 & ~n8915 ;
  assign n8940 = ~n8916 & ~n8939 ;
  assign n8941 = ~n8850 & ~n8852 ;
  assign n8942 = ~n8853 & ~n8941 ;
  assign n8943 = n8940 & n8942 ;
  assign n8944 = ~n8923 & ~n8924 ;
  assign n8945 = n8928 & n8944 ;
  assign n8946 = ~n8928 & ~n8944 ;
  assign n8947 = ~n8945 & ~n8946 ;
  assign n8948 = n8943 & n8947 ;
  assign n8949 = ~n8943 & ~n8947 ;
  assign n8950 = ~n8860 & ~n8861 ;
  assign n8951 = n8865 & n8950 ;
  assign n8952 = ~n8865 & ~n8950 ;
  assign n8953 = ~n8951 & ~n8952 ;
  assign n8954 = ~n8949 & n8953 ;
  assign n8955 = ~n8948 & ~n8954 ;
  assign n8956 = ~n8938 & ~n8955 ;
  assign n8957 = ~n8937 & ~n8956 ;
  assign n8958 = ~n8892 & ~n8932 ;
  assign n8959 = ~n8931 & ~n8958 ;
  assign n8960 = ~n8957 & ~n8959 ;
  assign n8961 = n8957 & n8959 ;
  assign n8962 = ~n8960 & ~n8961 ;
  assign n8963 = ~n8829 & ~n8869 ;
  assign n8964 = ~n8868 & ~n8963 ;
  assign n8965 = n8962 & ~n8964 ;
  assign n8966 = ~n8962 & n8964 ;
  assign n8967 = ~n8965 & ~n8966 ;
  assign n8968 = ~n8805 & ~n8806 ;
  assign n8969 = ~n8808 & n8968 ;
  assign n8970 = n8808 & ~n8968 ;
  assign n8971 = ~n8969 & ~n8970 ;
  assign n8972 = ~n8967 & ~n8971 ;
  assign n8973 = n8967 & n8971 ;
  assign n8974 = ~n8782 & ~n8783 ;
  assign n8975 = ~n8800 & n8974 ;
  assign n8976 = n8800 & ~n8974 ;
  assign n8977 = ~n8975 & ~n8976 ;
  assign n8978 = ~n8937 & ~n8938 ;
  assign n8979 = ~n8955 & n8978 ;
  assign n8980 = n8955 & ~n8978 ;
  assign n8981 = ~n8979 & ~n8980 ;
  assign n8982 = ~n8977 & ~n8981 ;
  assign n8983 = n8977 & n8981 ;
  assign n8984 = ~n8785 & ~n8787 ;
  assign n8985 = ~n8788 & ~n8984 ;
  assign n8986 = ~n8940 & ~n8942 ;
  assign n8987 = ~n8943 & ~n8986 ;
  assign n8988 = n8985 & n8987 ;
  assign n8989 = ~n8948 & ~n8949 ;
  assign n8990 = ~n8953 & n8989 ;
  assign n8991 = n8953 & ~n8989 ;
  assign n8992 = ~n8990 & ~n8991 ;
  assign n8993 = n8988 & ~n8992 ;
  assign n8994 = ~n8988 & n8992 ;
  assign n8995 = ~n8793 & ~n8794 ;
  assign n8996 = ~n8798 & n8995 ;
  assign n8997 = n8798 & ~n8995 ;
  assign n8998 = ~n8996 & ~n8997 ;
  assign n8999 = ~n8994 & ~n8998 ;
  assign n9000 = ~n8993 & ~n8999 ;
  assign n9001 = ~n8983 & n9000 ;
  assign n9002 = ~n8982 & ~n9001 ;
  assign n9003 = ~n8973 & ~n9002 ;
  assign n9004 = ~n8972 & ~n9003 ;
  assign n9005 = n8810 & ~n9004 ;
  assign n9006 = ~n8810 & n9004 ;
  assign n9007 = ~n9005 & ~n9006 ;
  assign n9008 = ~n8961 & ~n8964 ;
  assign n9009 = ~n8960 & ~n9008 ;
  assign n9010 = n9007 & n9009 ;
  assign n9011 = ~n9007 & ~n9009 ;
  assign n9012 = ~n9010 & ~n9011 ;
  assign n9013 = \A[538]  & \A[539]  ;
  assign n9014 = \A[535]  & \A[536]  ;
  assign n9015 = ~\A[535]  & ~\A[536]  ;
  assign n9016 = ~n9014 & ~n9015 ;
  assign n9017 = \A[537]  & n9016 ;
  assign n9018 = ~\A[537]  & ~n9016 ;
  assign n9019 = ~n9017 & ~n9018 ;
  assign n9020 = ~\A[538]  & ~\A[539]  ;
  assign n9021 = ~n9013 & ~n9020 ;
  assign n9022 = \A[540]  & n9021 ;
  assign n9023 = ~\A[540]  & ~n9021 ;
  assign n9024 = ~n9022 & ~n9023 ;
  assign n9025 = n9019 & n9024 ;
  assign n9026 = n9013 & n9025 ;
  assign n9027 = ~n9014 & ~n9017 ;
  assign n9028 = ~n9013 & ~n9022 ;
  assign n9029 = ~n9025 & n9028 ;
  assign n9030 = ~n9027 & ~n9029 ;
  assign n9031 = ~n9026 & ~n9030 ;
  assign n9032 = \A[544]  & \A[545]  ;
  assign n9033 = ~\A[544]  & ~\A[545]  ;
  assign n9034 = ~n9032 & ~n9033 ;
  assign n9035 = \A[546]  & n9034 ;
  assign n9036 = ~n9032 & ~n9035 ;
  assign n9037 = \A[541]  & \A[542]  ;
  assign n9038 = ~\A[541]  & ~\A[542]  ;
  assign n9039 = ~n9037 & ~n9038 ;
  assign n9040 = \A[543]  & n9039 ;
  assign n9041 = ~n9037 & ~n9040 ;
  assign n9042 = n9036 & n9041 ;
  assign n9043 = ~n9036 & ~n9041 ;
  assign n9044 = ~\A[543]  & ~n9039 ;
  assign n9045 = ~n9040 & ~n9044 ;
  assign n9046 = ~\A[546]  & ~n9034 ;
  assign n9047 = ~n9035 & ~n9046 ;
  assign n9048 = n9045 & n9047 ;
  assign n9049 = ~n9043 & ~n9048 ;
  assign n9050 = ~n9042 & ~n9049 ;
  assign n9051 = ~n9045 & ~n9047 ;
  assign n9052 = ~n9048 & ~n9051 ;
  assign n9053 = ~n9019 & ~n9024 ;
  assign n9054 = ~n9025 & ~n9053 ;
  assign n9055 = n9052 & n9054 ;
  assign n9056 = n9026 & ~n9027 ;
  assign n9057 = n9055 & ~n9056 ;
  assign n9058 = ~n9042 & ~n9043 ;
  assign n9059 = n9048 & ~n9058 ;
  assign n9060 = ~n9048 & n9058 ;
  assign n9061 = ~n9059 & ~n9060 ;
  assign n9062 = n9057 & ~n9061 ;
  assign n9063 = ~n9057 & n9061 ;
  assign n9064 = ~n9026 & ~n9029 ;
  assign n9065 = n9027 & ~n9064 ;
  assign n9066 = ~n9027 & n9064 ;
  assign n9067 = ~n9065 & ~n9066 ;
  assign n9068 = ~n9063 & n9067 ;
  assign n9069 = ~n9062 & ~n9068 ;
  assign n9070 = n9050 & ~n9069 ;
  assign n9071 = ~n9050 & n9069 ;
  assign n9072 = ~n9070 & ~n9071 ;
  assign n9073 = n9031 & n9072 ;
  assign n9074 = ~n9031 & ~n9072 ;
  assign n9075 = ~n9073 & ~n9074 ;
  assign n9076 = \A[550]  & \A[551]  ;
  assign n9077 = \A[547]  & \A[548]  ;
  assign n9078 = ~\A[547]  & ~\A[548]  ;
  assign n9079 = ~n9077 & ~n9078 ;
  assign n9080 = \A[549]  & n9079 ;
  assign n9081 = ~\A[549]  & ~n9079 ;
  assign n9082 = ~n9080 & ~n9081 ;
  assign n9083 = ~\A[550]  & ~\A[551]  ;
  assign n9084 = ~n9076 & ~n9083 ;
  assign n9085 = \A[552]  & n9084 ;
  assign n9086 = ~\A[552]  & ~n9084 ;
  assign n9087 = ~n9085 & ~n9086 ;
  assign n9088 = n9082 & n9087 ;
  assign n9089 = n9076 & n9088 ;
  assign n9090 = ~n9077 & ~n9080 ;
  assign n9091 = ~n9076 & ~n9085 ;
  assign n9092 = ~n9088 & n9091 ;
  assign n9093 = ~n9090 & ~n9092 ;
  assign n9094 = ~n9089 & ~n9093 ;
  assign n9095 = \A[556]  & \A[557]  ;
  assign n9096 = ~\A[556]  & ~\A[557]  ;
  assign n9097 = ~n9095 & ~n9096 ;
  assign n9098 = \A[558]  & n9097 ;
  assign n9099 = ~n9095 & ~n9098 ;
  assign n9100 = \A[553]  & \A[554]  ;
  assign n9101 = ~\A[553]  & ~\A[554]  ;
  assign n9102 = ~n9100 & ~n9101 ;
  assign n9103 = \A[555]  & n9102 ;
  assign n9104 = ~n9100 & ~n9103 ;
  assign n9105 = n9099 & n9104 ;
  assign n9106 = ~n9099 & ~n9104 ;
  assign n9107 = ~\A[555]  & ~n9102 ;
  assign n9108 = ~n9103 & ~n9107 ;
  assign n9109 = ~\A[558]  & ~n9097 ;
  assign n9110 = ~n9098 & ~n9109 ;
  assign n9111 = n9108 & n9110 ;
  assign n9112 = ~n9106 & ~n9111 ;
  assign n9113 = ~n9105 & ~n9112 ;
  assign n9114 = ~n9108 & ~n9110 ;
  assign n9115 = ~n9111 & ~n9114 ;
  assign n9116 = ~n9082 & ~n9087 ;
  assign n9117 = ~n9088 & ~n9116 ;
  assign n9118 = n9115 & n9117 ;
  assign n9119 = n9089 & ~n9090 ;
  assign n9120 = n9118 & ~n9119 ;
  assign n9121 = ~n9105 & ~n9106 ;
  assign n9122 = n9111 & ~n9121 ;
  assign n9123 = ~n9111 & n9121 ;
  assign n9124 = ~n9122 & ~n9123 ;
  assign n9125 = n9120 & ~n9124 ;
  assign n9126 = ~n9120 & n9124 ;
  assign n9127 = ~n9089 & ~n9092 ;
  assign n9128 = n9090 & ~n9127 ;
  assign n9129 = ~n9090 & n9127 ;
  assign n9130 = ~n9128 & ~n9129 ;
  assign n9131 = ~n9126 & n9130 ;
  assign n9132 = ~n9125 & ~n9131 ;
  assign n9133 = n9113 & ~n9132 ;
  assign n9134 = ~n9113 & n9132 ;
  assign n9135 = ~n9133 & ~n9134 ;
  assign n9136 = n9094 & n9135 ;
  assign n9137 = ~n9094 & ~n9135 ;
  assign n9138 = ~n9136 & ~n9137 ;
  assign n9139 = ~n9075 & ~n9138 ;
  assign n9140 = n9075 & n9138 ;
  assign n9141 = ~n9115 & ~n9117 ;
  assign n9142 = ~n9118 & ~n9141 ;
  assign n9143 = ~n9052 & ~n9054 ;
  assign n9144 = ~n9055 & ~n9143 ;
  assign n9145 = n9142 & n9144 ;
  assign n9146 = ~n9125 & ~n9126 ;
  assign n9147 = n9130 & n9146 ;
  assign n9148 = ~n9130 & ~n9146 ;
  assign n9149 = ~n9147 & ~n9148 ;
  assign n9150 = n9145 & n9149 ;
  assign n9151 = ~n9145 & ~n9149 ;
  assign n9152 = ~n9062 & ~n9063 ;
  assign n9153 = n9067 & n9152 ;
  assign n9154 = ~n9067 & ~n9152 ;
  assign n9155 = ~n9153 & ~n9154 ;
  assign n9156 = ~n9151 & n9155 ;
  assign n9157 = ~n9150 & ~n9156 ;
  assign n9158 = ~n9140 & ~n9157 ;
  assign n9159 = ~n9139 & ~n9158 ;
  assign n9160 = ~n9094 & ~n9134 ;
  assign n9161 = ~n9133 & ~n9160 ;
  assign n9162 = ~n9159 & ~n9161 ;
  assign n9163 = n9159 & n9161 ;
  assign n9164 = ~n9031 & ~n9071 ;
  assign n9165 = ~n9070 & ~n9164 ;
  assign n9166 = ~n9163 & ~n9165 ;
  assign n9167 = ~n9162 & ~n9166 ;
  assign n9168 = ~n9162 & ~n9163 ;
  assign n9169 = ~n9165 & n9168 ;
  assign n9170 = n9165 & ~n9168 ;
  assign n9171 = ~n9169 & ~n9170 ;
  assign n9172 = \A[514]  & \A[515]  ;
  assign n9173 = \A[511]  & \A[512]  ;
  assign n9174 = ~\A[511]  & ~\A[512]  ;
  assign n9175 = ~n9173 & ~n9174 ;
  assign n9176 = \A[513]  & n9175 ;
  assign n9177 = ~\A[513]  & ~n9175 ;
  assign n9178 = ~n9176 & ~n9177 ;
  assign n9179 = ~\A[514]  & ~\A[515]  ;
  assign n9180 = ~n9172 & ~n9179 ;
  assign n9181 = \A[516]  & n9180 ;
  assign n9182 = ~\A[516]  & ~n9180 ;
  assign n9183 = ~n9181 & ~n9182 ;
  assign n9184 = n9178 & n9183 ;
  assign n9185 = n9172 & n9184 ;
  assign n9186 = ~n9173 & ~n9176 ;
  assign n9187 = ~n9172 & ~n9181 ;
  assign n9188 = ~n9184 & n9187 ;
  assign n9189 = ~n9186 & ~n9188 ;
  assign n9190 = ~n9185 & ~n9189 ;
  assign n9191 = \A[520]  & \A[521]  ;
  assign n9192 = ~\A[520]  & ~\A[521]  ;
  assign n9193 = ~n9191 & ~n9192 ;
  assign n9194 = \A[522]  & n9193 ;
  assign n9195 = ~n9191 & ~n9194 ;
  assign n9196 = \A[517]  & \A[518]  ;
  assign n9197 = ~\A[517]  & ~\A[518]  ;
  assign n9198 = ~n9196 & ~n9197 ;
  assign n9199 = \A[519]  & n9198 ;
  assign n9200 = ~n9196 & ~n9199 ;
  assign n9201 = n9195 & n9200 ;
  assign n9202 = ~n9195 & ~n9200 ;
  assign n9203 = ~\A[519]  & ~n9198 ;
  assign n9204 = ~n9199 & ~n9203 ;
  assign n9205 = ~\A[522]  & ~n9193 ;
  assign n9206 = ~n9194 & ~n9205 ;
  assign n9207 = n9204 & n9206 ;
  assign n9208 = ~n9202 & ~n9207 ;
  assign n9209 = ~n9201 & ~n9208 ;
  assign n9210 = ~n9204 & ~n9206 ;
  assign n9211 = ~n9207 & ~n9210 ;
  assign n9212 = ~n9178 & ~n9183 ;
  assign n9213 = ~n9184 & ~n9212 ;
  assign n9214 = n9211 & n9213 ;
  assign n9215 = n9185 & ~n9186 ;
  assign n9216 = n9214 & ~n9215 ;
  assign n9217 = ~n9201 & ~n9202 ;
  assign n9218 = n9207 & ~n9217 ;
  assign n9219 = ~n9207 & n9217 ;
  assign n9220 = ~n9218 & ~n9219 ;
  assign n9221 = n9216 & ~n9220 ;
  assign n9222 = ~n9216 & n9220 ;
  assign n9223 = ~n9185 & ~n9188 ;
  assign n9224 = n9186 & ~n9223 ;
  assign n9225 = ~n9186 & n9223 ;
  assign n9226 = ~n9224 & ~n9225 ;
  assign n9227 = ~n9222 & n9226 ;
  assign n9228 = ~n9221 & ~n9227 ;
  assign n9229 = n9209 & ~n9228 ;
  assign n9230 = ~n9209 & n9228 ;
  assign n9231 = ~n9229 & ~n9230 ;
  assign n9232 = n9190 & n9231 ;
  assign n9233 = ~n9190 & ~n9231 ;
  assign n9234 = ~n9232 & ~n9233 ;
  assign n9235 = \A[526]  & \A[527]  ;
  assign n9236 = \A[523]  & \A[524]  ;
  assign n9237 = ~\A[523]  & ~\A[524]  ;
  assign n9238 = ~n9236 & ~n9237 ;
  assign n9239 = \A[525]  & n9238 ;
  assign n9240 = ~\A[525]  & ~n9238 ;
  assign n9241 = ~n9239 & ~n9240 ;
  assign n9242 = ~\A[526]  & ~\A[527]  ;
  assign n9243 = ~n9235 & ~n9242 ;
  assign n9244 = \A[528]  & n9243 ;
  assign n9245 = ~\A[528]  & ~n9243 ;
  assign n9246 = ~n9244 & ~n9245 ;
  assign n9247 = n9241 & n9246 ;
  assign n9248 = n9235 & n9247 ;
  assign n9249 = ~n9236 & ~n9239 ;
  assign n9250 = ~n9235 & ~n9244 ;
  assign n9251 = ~n9247 & n9250 ;
  assign n9252 = ~n9249 & ~n9251 ;
  assign n9253 = ~n9248 & ~n9252 ;
  assign n9254 = \A[532]  & \A[533]  ;
  assign n9255 = ~\A[532]  & ~\A[533]  ;
  assign n9256 = ~n9254 & ~n9255 ;
  assign n9257 = \A[534]  & n9256 ;
  assign n9258 = ~n9254 & ~n9257 ;
  assign n9259 = \A[529]  & \A[530]  ;
  assign n9260 = ~\A[529]  & ~\A[530]  ;
  assign n9261 = ~n9259 & ~n9260 ;
  assign n9262 = \A[531]  & n9261 ;
  assign n9263 = ~n9259 & ~n9262 ;
  assign n9264 = n9258 & n9263 ;
  assign n9265 = ~n9258 & ~n9263 ;
  assign n9266 = ~\A[531]  & ~n9261 ;
  assign n9267 = ~n9262 & ~n9266 ;
  assign n9268 = ~\A[534]  & ~n9256 ;
  assign n9269 = ~n9257 & ~n9268 ;
  assign n9270 = n9267 & n9269 ;
  assign n9271 = ~n9265 & ~n9270 ;
  assign n9272 = ~n9264 & ~n9271 ;
  assign n9273 = ~n9267 & ~n9269 ;
  assign n9274 = ~n9270 & ~n9273 ;
  assign n9275 = ~n9241 & ~n9246 ;
  assign n9276 = ~n9247 & ~n9275 ;
  assign n9277 = n9274 & n9276 ;
  assign n9278 = n9248 & ~n9249 ;
  assign n9279 = n9277 & ~n9278 ;
  assign n9280 = ~n9264 & ~n9265 ;
  assign n9281 = n9270 & ~n9280 ;
  assign n9282 = ~n9270 & n9280 ;
  assign n9283 = ~n9281 & ~n9282 ;
  assign n9284 = n9279 & ~n9283 ;
  assign n9285 = ~n9279 & n9283 ;
  assign n9286 = ~n9248 & ~n9251 ;
  assign n9287 = n9249 & ~n9286 ;
  assign n9288 = ~n9249 & n9286 ;
  assign n9289 = ~n9287 & ~n9288 ;
  assign n9290 = ~n9285 & n9289 ;
  assign n9291 = ~n9284 & ~n9290 ;
  assign n9292 = n9272 & ~n9291 ;
  assign n9293 = ~n9272 & n9291 ;
  assign n9294 = ~n9292 & ~n9293 ;
  assign n9295 = n9253 & n9294 ;
  assign n9296 = ~n9253 & ~n9294 ;
  assign n9297 = ~n9295 & ~n9296 ;
  assign n9298 = ~n9234 & ~n9297 ;
  assign n9299 = n9234 & n9297 ;
  assign n9300 = ~n9274 & ~n9276 ;
  assign n9301 = ~n9277 & ~n9300 ;
  assign n9302 = ~n9211 & ~n9213 ;
  assign n9303 = ~n9214 & ~n9302 ;
  assign n9304 = n9301 & n9303 ;
  assign n9305 = ~n9284 & ~n9285 ;
  assign n9306 = n9289 & n9305 ;
  assign n9307 = ~n9289 & ~n9305 ;
  assign n9308 = ~n9306 & ~n9307 ;
  assign n9309 = n9304 & n9308 ;
  assign n9310 = ~n9304 & ~n9308 ;
  assign n9311 = ~n9221 & ~n9222 ;
  assign n9312 = n9226 & n9311 ;
  assign n9313 = ~n9226 & ~n9311 ;
  assign n9314 = ~n9312 & ~n9313 ;
  assign n9315 = ~n9310 & n9314 ;
  assign n9316 = ~n9309 & ~n9315 ;
  assign n9317 = ~n9299 & ~n9316 ;
  assign n9318 = ~n9298 & ~n9317 ;
  assign n9319 = ~n9253 & ~n9293 ;
  assign n9320 = ~n9292 & ~n9319 ;
  assign n9321 = ~n9318 & ~n9320 ;
  assign n9322 = n9318 & n9320 ;
  assign n9323 = ~n9321 & ~n9322 ;
  assign n9324 = ~n9190 & ~n9230 ;
  assign n9325 = ~n9229 & ~n9324 ;
  assign n9326 = n9323 & ~n9325 ;
  assign n9327 = ~n9323 & n9325 ;
  assign n9328 = ~n9326 & ~n9327 ;
  assign n9329 = ~n9171 & ~n9328 ;
  assign n9330 = n9171 & n9328 ;
  assign n9331 = ~n9298 & ~n9299 ;
  assign n9332 = ~n9316 & n9331 ;
  assign n9333 = n9316 & ~n9331 ;
  assign n9334 = ~n9332 & ~n9333 ;
  assign n9335 = ~n9139 & ~n9140 ;
  assign n9336 = ~n9157 & n9335 ;
  assign n9337 = n9157 & ~n9335 ;
  assign n9338 = ~n9336 & ~n9337 ;
  assign n9339 = ~n9334 & ~n9338 ;
  assign n9340 = n9334 & n9338 ;
  assign n9341 = ~n9142 & ~n9144 ;
  assign n9342 = ~n9145 & ~n9341 ;
  assign n9343 = ~n9301 & ~n9303 ;
  assign n9344 = ~n9304 & ~n9343 ;
  assign n9345 = n9342 & n9344 ;
  assign n9346 = ~n9150 & ~n9151 ;
  assign n9347 = ~n9155 & n9346 ;
  assign n9348 = n9155 & ~n9346 ;
  assign n9349 = ~n9347 & ~n9348 ;
  assign n9350 = n9345 & ~n9349 ;
  assign n9351 = ~n9345 & n9349 ;
  assign n9352 = ~n9309 & ~n9310 ;
  assign n9353 = ~n9314 & n9352 ;
  assign n9354 = n9314 & ~n9352 ;
  assign n9355 = ~n9353 & ~n9354 ;
  assign n9356 = ~n9351 & ~n9355 ;
  assign n9357 = ~n9350 & ~n9356 ;
  assign n9358 = ~n9340 & n9357 ;
  assign n9359 = ~n9339 & ~n9358 ;
  assign n9360 = ~n9330 & ~n9359 ;
  assign n9361 = ~n9329 & ~n9360 ;
  assign n9362 = n9167 & ~n9361 ;
  assign n9363 = ~n9167 & n9361 ;
  assign n9364 = ~n9362 & ~n9363 ;
  assign n9365 = ~n9322 & ~n9325 ;
  assign n9366 = ~n9321 & ~n9365 ;
  assign n9367 = n9364 & n9366 ;
  assign n9368 = ~n9364 & ~n9366 ;
  assign n9369 = ~n9367 & ~n9368 ;
  assign n9370 = ~n9012 & ~n9369 ;
  assign n9371 = n9012 & n9369 ;
  assign n9372 = ~n9329 & ~n9330 ;
  assign n9373 = ~n9359 & n9372 ;
  assign n9374 = n9359 & ~n9372 ;
  assign n9375 = ~n9373 & ~n9374 ;
  assign n9376 = ~n8972 & ~n8973 ;
  assign n9377 = ~n9002 & n9376 ;
  assign n9378 = n9002 & ~n9376 ;
  assign n9379 = ~n9377 & ~n9378 ;
  assign n9380 = ~n9375 & ~n9379 ;
  assign n9381 = n9375 & n9379 ;
  assign n9382 = ~n8982 & ~n8983 ;
  assign n9383 = ~n9000 & n9382 ;
  assign n9384 = n9000 & ~n9382 ;
  assign n9385 = ~n9383 & ~n9384 ;
  assign n9386 = ~n9339 & ~n9340 ;
  assign n9387 = ~n9357 & n9386 ;
  assign n9388 = n9357 & ~n9386 ;
  assign n9389 = ~n9387 & ~n9388 ;
  assign n9390 = ~n9385 & ~n9389 ;
  assign n9391 = n9385 & n9389 ;
  assign n9392 = ~n8985 & ~n8987 ;
  assign n9393 = ~n8988 & ~n9392 ;
  assign n9394 = ~n9342 & ~n9344 ;
  assign n9395 = ~n9345 & ~n9394 ;
  assign n9396 = n9393 & n9395 ;
  assign n9397 = ~n9350 & ~n9351 ;
  assign n9398 = ~n9355 & n9397 ;
  assign n9399 = n9355 & ~n9397 ;
  assign n9400 = ~n9398 & ~n9399 ;
  assign n9401 = n9396 & n9400 ;
  assign n9402 = ~n9396 & ~n9400 ;
  assign n9403 = ~n8993 & ~n8994 ;
  assign n9404 = ~n8998 & n9403 ;
  assign n9405 = n8998 & ~n9403 ;
  assign n9406 = ~n9404 & ~n9405 ;
  assign n9407 = ~n9402 & n9406 ;
  assign n9408 = ~n9401 & ~n9407 ;
  assign n9409 = ~n9391 & n9408 ;
  assign n9410 = ~n9390 & ~n9409 ;
  assign n9411 = ~n9381 & n9410 ;
  assign n9412 = ~n9380 & ~n9411 ;
  assign n9413 = ~n9371 & ~n9412 ;
  assign n9414 = ~n9370 & ~n9413 ;
  assign n9415 = ~n9006 & n9009 ;
  assign n9416 = ~n9005 & ~n9415 ;
  assign n9417 = n9414 & ~n9416 ;
  assign n9418 = ~n9414 & n9416 ;
  assign n9419 = ~n9363 & n9366 ;
  assign n9420 = ~n9362 & ~n9419 ;
  assign n9421 = ~n9418 & ~n9420 ;
  assign n9422 = ~n9417 & ~n9421 ;
  assign n9423 = n8655 & n9422 ;
  assign n9424 = ~n8655 & ~n9422 ;
  assign n9425 = ~n8650 & ~n8651 ;
  assign n9426 = ~n8653 & n9425 ;
  assign n9427 = n8653 & ~n9425 ;
  assign n9428 = ~n9426 & ~n9427 ;
  assign n9429 = ~n9417 & ~n9418 ;
  assign n9430 = ~n9420 & n9429 ;
  assign n9431 = n9420 & ~n9429 ;
  assign n9432 = ~n9430 & ~n9431 ;
  assign n9433 = ~n9428 & ~n9432 ;
  assign n9434 = n9428 & n9432 ;
  assign n9435 = ~n9370 & ~n9371 ;
  assign n9436 = ~n9412 & n9435 ;
  assign n9437 = n9412 & ~n9435 ;
  assign n9438 = ~n9436 & ~n9437 ;
  assign n9439 = ~n8603 & ~n8604 ;
  assign n9440 = ~n8645 & n9439 ;
  assign n9441 = n8645 & ~n9439 ;
  assign n9442 = ~n9440 & ~n9441 ;
  assign n9443 = ~n9438 & ~n9442 ;
  assign n9444 = n9438 & n9442 ;
  assign n9445 = ~n8613 & ~n8614 ;
  assign n9446 = n8643 & n9445 ;
  assign n9447 = ~n8643 & ~n9445 ;
  assign n9448 = ~n9446 & ~n9447 ;
  assign n9449 = ~n9380 & ~n9381 ;
  assign n9450 = n9410 & n9449 ;
  assign n9451 = ~n9410 & ~n9449 ;
  assign n9452 = ~n9450 & ~n9451 ;
  assign n9453 = ~n9448 & ~n9452 ;
  assign n9454 = n9448 & n9452 ;
  assign n9455 = ~n9390 & ~n9391 ;
  assign n9456 = ~n9408 & n9455 ;
  assign n9457 = n9408 & ~n9455 ;
  assign n9458 = ~n9456 & ~n9457 ;
  assign n9459 = ~n8623 & ~n8624 ;
  assign n9460 = ~n8641 & n9459 ;
  assign n9461 = n8641 & ~n9459 ;
  assign n9462 = ~n9460 & ~n9461 ;
  assign n9463 = ~n9458 & ~n9462 ;
  assign n9464 = n9458 & n9462 ;
  assign n9465 = ~n9393 & ~n9395 ;
  assign n9466 = ~n9396 & ~n9465 ;
  assign n9467 = ~n8626 & ~n8628 ;
  assign n9468 = ~n8629 & ~n9467 ;
  assign n9469 = n9466 & n9468 ;
  assign n9470 = ~n8634 & ~n8635 ;
  assign n9471 = ~n8639 & n9470 ;
  assign n9472 = n8639 & ~n9470 ;
  assign n9473 = ~n9471 & ~n9472 ;
  assign n9474 = n9469 & ~n9473 ;
  assign n9475 = ~n9469 & n9473 ;
  assign n9476 = ~n9401 & ~n9402 ;
  assign n9477 = ~n9406 & n9476 ;
  assign n9478 = n9406 & ~n9476 ;
  assign n9479 = ~n9477 & ~n9478 ;
  assign n9480 = ~n9475 & ~n9479 ;
  assign n9481 = ~n9474 & ~n9480 ;
  assign n9482 = ~n9464 & n9481 ;
  assign n9483 = ~n9463 & ~n9482 ;
  assign n9484 = ~n9454 & ~n9483 ;
  assign n9485 = ~n9453 & ~n9484 ;
  assign n9486 = ~n9444 & ~n9485 ;
  assign n9487 = ~n9443 & ~n9486 ;
  assign n9488 = ~n9434 & n9487 ;
  assign n9489 = ~n9433 & ~n9488 ;
  assign n9490 = ~n9424 & ~n9489 ;
  assign n9491 = ~n9423 & ~n9490 ;
  assign n9492 = ~n7888 & ~n9491 ;
  assign n9493 = n7888 & n9491 ;
  assign n9494 = ~n9423 & ~n9424 ;
  assign n9495 = ~n9489 & n9494 ;
  assign n9496 = n9489 & ~n9494 ;
  assign n9497 = ~n9495 & ~n9496 ;
  assign n9498 = ~n7820 & ~n7821 ;
  assign n9499 = ~n7886 & n9498 ;
  assign n9500 = n7886 & ~n9498 ;
  assign n9501 = ~n9499 & ~n9500 ;
  assign n9502 = n9497 & ~n9501 ;
  assign n9503 = ~n9497 & n9501 ;
  assign n9504 = ~n7830 & ~n7831 ;
  assign n9505 = ~n7884 & n9504 ;
  assign n9506 = n7884 & ~n9504 ;
  assign n9507 = ~n9505 & ~n9506 ;
  assign n9508 = ~n9433 & ~n9434 ;
  assign n9509 = ~n9487 & n9508 ;
  assign n9510 = n9487 & ~n9508 ;
  assign n9511 = ~n9509 & ~n9510 ;
  assign n9512 = ~n9507 & ~n9511 ;
  assign n9513 = n9507 & n9511 ;
  assign n9514 = ~n9443 & ~n9444 ;
  assign n9515 = ~n9485 & n9514 ;
  assign n9516 = n9485 & ~n9514 ;
  assign n9517 = ~n9515 & ~n9516 ;
  assign n9518 = ~n7840 & ~n7841 ;
  assign n9519 = ~n7882 & n9518 ;
  assign n9520 = n7882 & ~n9518 ;
  assign n9521 = ~n9519 & ~n9520 ;
  assign n9522 = ~n9517 & ~n9521 ;
  assign n9523 = n9517 & n9521 ;
  assign n9524 = ~n7850 & ~n7851 ;
  assign n9525 = ~n7880 & n9524 ;
  assign n9526 = n7880 & ~n9524 ;
  assign n9527 = ~n9525 & ~n9526 ;
  assign n9528 = ~n9453 & ~n9454 ;
  assign n9529 = ~n9483 & n9528 ;
  assign n9530 = n9483 & ~n9528 ;
  assign n9531 = ~n9529 & ~n9530 ;
  assign n9532 = ~n9527 & ~n9531 ;
  assign n9533 = n9527 & n9531 ;
  assign n9534 = ~n9463 & ~n9464 ;
  assign n9535 = ~n9481 & n9534 ;
  assign n9536 = n9481 & ~n9534 ;
  assign n9537 = ~n9535 & ~n9536 ;
  assign n9538 = ~n7860 & ~n7861 ;
  assign n9539 = ~n7878 & n9538 ;
  assign n9540 = n7878 & ~n9538 ;
  assign n9541 = ~n9539 & ~n9540 ;
  assign n9542 = ~n9537 & ~n9541 ;
  assign n9543 = n9537 & n9541 ;
  assign n9544 = ~n9466 & ~n9468 ;
  assign n9545 = ~n9469 & ~n9544 ;
  assign n9546 = ~n7863 & ~n7865 ;
  assign n9547 = ~n7866 & ~n9546 ;
  assign n9548 = n9545 & n9547 ;
  assign n9549 = ~n7871 & ~n7872 ;
  assign n9550 = ~n7876 & n9549 ;
  assign n9551 = n7876 & ~n9549 ;
  assign n9552 = ~n9550 & ~n9551 ;
  assign n9553 = n9548 & n9552 ;
  assign n9554 = ~n9548 & ~n9552 ;
  assign n9555 = ~n9474 & ~n9475 ;
  assign n9556 = ~n9479 & n9555 ;
  assign n9557 = n9479 & ~n9555 ;
  assign n9558 = ~n9556 & ~n9557 ;
  assign n9559 = ~n9554 & n9558 ;
  assign n9560 = ~n9553 & ~n9559 ;
  assign n9561 = ~n9543 & n9560 ;
  assign n9562 = ~n9542 & ~n9561 ;
  assign n9563 = ~n9533 & n9562 ;
  assign n9564 = ~n9532 & ~n9563 ;
  assign n9565 = ~n9523 & ~n9564 ;
  assign n9566 = ~n9522 & ~n9565 ;
  assign n9567 = ~n9513 & ~n9566 ;
  assign n9568 = ~n9512 & ~n9567 ;
  assign n9569 = ~n9503 & ~n9568 ;
  assign n9570 = ~n9502 & ~n9569 ;
  assign n9571 = ~n9493 & ~n9570 ;
  assign n9572 = ~n9492 & ~n9571 ;
  assign n9573 = n6307 & n9572 ;
  assign n9574 = ~n6224 & ~n6225 ;
  assign n9575 = ~n6302 & n9574 ;
  assign n9576 = n6302 & ~n9574 ;
  assign n9577 = ~n9575 & ~n9576 ;
  assign n9578 = ~n9492 & ~n9493 ;
  assign n9579 = ~n9570 & n9578 ;
  assign n9580 = n9570 & ~n9578 ;
  assign n9581 = ~n9579 & ~n9580 ;
  assign n9582 = n9577 & ~n9581 ;
  assign n9583 = ~n9577 & n9581 ;
  assign n9584 = ~n6234 & ~n6235 ;
  assign n9585 = ~n6300 & n9584 ;
  assign n9586 = n6300 & ~n9584 ;
  assign n9587 = ~n9585 & ~n9586 ;
  assign n9588 = ~n9502 & ~n9503 ;
  assign n9589 = ~n9568 & n9588 ;
  assign n9590 = n9568 & ~n9588 ;
  assign n9591 = ~n9589 & ~n9590 ;
  assign n9592 = n9587 & ~n9591 ;
  assign n9593 = ~n9587 & n9591 ;
  assign n9594 = ~n6244 & ~n6245 ;
  assign n9595 = ~n6298 & n9594 ;
  assign n9596 = n6298 & ~n9594 ;
  assign n9597 = ~n9595 & ~n9596 ;
  assign n9598 = ~n9512 & ~n9513 ;
  assign n9599 = ~n9566 & n9598 ;
  assign n9600 = n9566 & ~n9598 ;
  assign n9601 = ~n9599 & ~n9600 ;
  assign n9602 = ~n9597 & n9601 ;
  assign n9603 = n9597 & ~n9601 ;
  assign n9604 = ~n6254 & ~n6255 ;
  assign n9605 = ~n6296 & n9604 ;
  assign n9606 = n6296 & ~n9604 ;
  assign n9607 = ~n9605 & ~n9606 ;
  assign n9608 = ~n9522 & ~n9523 ;
  assign n9609 = ~n9564 & n9608 ;
  assign n9610 = n9564 & ~n9608 ;
  assign n9611 = ~n9609 & ~n9610 ;
  assign n9612 = ~n9607 & ~n9611 ;
  assign n9613 = n9607 & n9611 ;
  assign n9614 = ~n6264 & ~n6265 ;
  assign n9615 = n6294 & n9614 ;
  assign n9616 = ~n6294 & ~n9614 ;
  assign n9617 = ~n9615 & ~n9616 ;
  assign n9618 = ~n9532 & ~n9533 ;
  assign n9619 = n9562 & n9618 ;
  assign n9620 = ~n9562 & ~n9618 ;
  assign n9621 = ~n9619 & ~n9620 ;
  assign n9622 = ~n9617 & ~n9621 ;
  assign n9623 = n9617 & n9621 ;
  assign n9624 = ~n6274 & ~n6275 ;
  assign n9625 = ~n6292 & n9624 ;
  assign n9626 = n6292 & ~n9624 ;
  assign n9627 = ~n9625 & ~n9626 ;
  assign n9628 = ~n9542 & ~n9543 ;
  assign n9629 = ~n9560 & n9628 ;
  assign n9630 = n9560 & ~n9628 ;
  assign n9631 = ~n9629 & ~n9630 ;
  assign n9632 = n9627 & n9631 ;
  assign n9633 = ~n9627 & ~n9631 ;
  assign n9634 = ~n9545 & ~n9547 ;
  assign n9635 = ~n9548 & ~n9634 ;
  assign n9636 = ~n6277 & ~n6279 ;
  assign n9637 = ~n6280 & ~n9636 ;
  assign n9638 = n9635 & n9637 ;
  assign n9639 = ~n6285 & ~n6286 ;
  assign n9640 = ~n6290 & n9639 ;
  assign n9641 = n6290 & ~n9639 ;
  assign n9642 = ~n9640 & ~n9641 ;
  assign n9643 = ~n9638 & n9642 ;
  assign n9644 = n9638 & ~n9642 ;
  assign n9645 = ~n9553 & ~n9554 ;
  assign n9646 = ~n9558 & n9645 ;
  assign n9647 = n9558 & ~n9645 ;
  assign n9648 = ~n9646 & ~n9647 ;
  assign n9649 = ~n9644 & n9648 ;
  assign n9650 = ~n9643 & ~n9649 ;
  assign n9651 = ~n9633 & n9650 ;
  assign n9652 = ~n9632 & ~n9651 ;
  assign n9653 = ~n9623 & n9652 ;
  assign n9654 = ~n9622 & ~n9653 ;
  assign n9655 = ~n9613 & ~n9654 ;
  assign n9656 = ~n9612 & ~n9655 ;
  assign n9657 = ~n9603 & n9656 ;
  assign n9658 = ~n9602 & ~n9657 ;
  assign n9659 = ~n9593 & n9658 ;
  assign n9660 = ~n9592 & ~n9659 ;
  assign n9661 = ~n9583 & ~n9660 ;
  assign n9662 = ~n9582 & ~n9661 ;
  assign n9663 = n9573 & ~n9662 ;
  assign n9692 = ~n9582 & ~n9583 ;
  assign n9693 = ~n9660 & n9692 ;
  assign n9694 = n9660 & ~n9692 ;
  assign n9695 = ~n9693 & ~n9694 ;
  assign n9668 = ~n9592 & ~n9593 ;
  assign n9670 = ~n9658 & n9668 ;
  assign n9669 = n9658 & ~n9668 ;
  assign n9671 = ~n9602 & ~n9603 ;
  assign n9673 = ~n9656 & ~n9671 ;
  assign n9672 = n9656 & n9671 ;
  assign n9664 = ~n9612 & ~n9613 ;
  assign n9665 = n9654 & ~n9664 ;
  assign n9666 = ~n9654 & n9664 ;
  assign n9667 = ~n9665 & ~n9666 ;
  assign n9687 = ~n9622 & ~n9623 ;
  assign n9689 = n9652 & n9687 ;
  assign n9684 = ~n9632 & n9651 ;
  assign n9674 = ~n9632 & ~n9633 ;
  assign n9675 = ~n9650 & ~n9674 ;
  assign n9677 = ~n9643 & ~n9644 ;
  assign n9678 = ~n9648 & ~n9677 ;
  assign n9676 = ~n9643 & n9649 ;
  assign n9679 = ~n9635 & ~n9637 ;
  assign n9680 = ~n9638 & ~n9679 ;
  assign n9681 = ~\A[1000]  & ~n9680 ;
  assign n9682 = ~n9676 & n9681 ;
  assign n9683 = ~n9678 & n9682 ;
  assign n9685 = ~n9675 & ~n9683 ;
  assign n9686 = ~n9684 & n9685 ;
  assign n9688 = ~n9652 & ~n9687 ;
  assign n9690 = ~n9686 & ~n9688 ;
  assign n9691 = ~n9689 & n9690 ;
  assign n9696 = ~n9667 & ~n9691 ;
  assign n9697 = ~n9672 & n9696 ;
  assign n9698 = ~n9673 & n9697 ;
  assign n9699 = ~n9669 & n9698 ;
  assign n9700 = ~n9670 & n9699 ;
  assign n9701 = ~n9695 & n9700 ;
  assign n9702 = ~n9663 & n9701 ;
  assign n9703 = ~n9573 & n9662 ;
  assign n9705 = ~n6307 & ~n9572 ;
  assign n9704 = ~n6213 & n6304 ;
  assign n9706 = ~n6214 & ~n9704 ;
  assign n9707 = ~n9705 & n9706 ;
  assign n9708 = ~n9703 & n9707 ;
  assign n9709 = ~n9702 & n9708 ;
  assign maj = ~n9709 ;
endmodule
