module top( a_pad , b_pad , c_pad , d_pad , e_pad , f_pad , g_pad , h_pad , i_pad , j_pad , k_pad , l_pad , m_pad , n_pad , o_pad , p_pad , q_pad , r_pad , s_pad , t_pad , u_pad , v_pad );
  input a_pad ;
  input b_pad ;
  input c_pad ;
  input d_pad ;
  input e_pad ;
  input f_pad ;
  input g_pad ;
  input h_pad ;
  input i_pad ;
  input j_pad ;
  input k_pad ;
  input l_pad ;
  input m_pad ;
  input n_pad ;
  input o_pad ;
  input p_pad ;
  input q_pad ;
  input r_pad ;
  input s_pad ;
  input t_pad ;
  input u_pad ;
  output v_pad ;
  wire n22 , n23 , n24 , n25 , n26 , n27 , n28 , n29 , n30 , n31 , n32 , n33 , n34 , n35 , n36 , n37 , n38 , n39 , n40 , n41 , n42 , n43 , n44 , n45 , n46 , n47 , n48 , n49 , n50 , n51 , n52 , n53 , n54 , n55 , n56 , n57 , n58 , n59 , n60 , n61 , n62 , n63 , n64 , n65 , n66 , n67 ;
  assign n33 = o_pad & ~q_pad ;
  assign n32 = p_pad & q_pad ;
  assign n34 = r_pad & ~n32 ;
  assign n35 = ~n33 & n34 ;
  assign n37 = m_pad & ~q_pad ;
  assign n36 = n_pad & q_pad ;
  assign n38 = ~r_pad & ~n36 ;
  assign n39 = ~n37 & n38 ;
  assign n40 = ~n35 & ~n39 ;
  assign n41 = s_pad & ~n40 ;
  assign n23 = i_pad & ~q_pad ;
  assign n22 = j_pad & q_pad ;
  assign n24 = ~r_pad & ~n22 ;
  assign n25 = ~n23 & n24 ;
  assign n27 = k_pad & ~q_pad ;
  assign n26 = l_pad & q_pad ;
  assign n28 = r_pad & ~n26 ;
  assign n29 = ~n27 & n28 ;
  assign n30 = ~n25 & ~n29 ;
  assign n31 = ~s_pad & ~n30 ;
  assign n42 = t_pad & ~n31 ;
  assign n43 = ~n41 & n42 ;
  assign n55 = g_pad & ~q_pad ;
  assign n54 = h_pad & q_pad ;
  assign n56 = r_pad & ~n54 ;
  assign n57 = ~n55 & n56 ;
  assign n59 = e_pad & ~q_pad ;
  assign n58 = f_pad & q_pad ;
  assign n60 = ~r_pad & ~n58 ;
  assign n61 = ~n59 & n60 ;
  assign n62 = ~n57 & ~n61 ;
  assign n63 = s_pad & ~n62 ;
  assign n45 = a_pad & ~q_pad ;
  assign n44 = b_pad & q_pad ;
  assign n46 = ~r_pad & ~n44 ;
  assign n47 = ~n45 & n46 ;
  assign n49 = c_pad & ~q_pad ;
  assign n48 = d_pad & q_pad ;
  assign n50 = r_pad & ~n48 ;
  assign n51 = ~n49 & n50 ;
  assign n52 = ~n47 & ~n51 ;
  assign n53 = ~s_pad & ~n52 ;
  assign n64 = ~t_pad & ~n53 ;
  assign n65 = ~n63 & n64 ;
  assign n66 = ~n43 & ~n65 ;
  assign n67 = ~u_pad & ~n66 ;
  assign v_pad = ~n67 ;
endmodule
