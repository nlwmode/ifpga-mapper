module top( \pi000  , \pi001  , \pi002  , \pi003  , \pi004  , \pi005  , \pi006  , \pi007  , \pi008  , \pi009  , \pi010  , \pi011  , \pi012  , \pi013  , \pi014  , \pi015  , \pi016  , \pi017  , \pi018  , \pi019  , \pi020  , \pi021  , \pi022  , \pi023  , \pi024  , \pi025  , \pi026  , \pi027  , \pi028  , \pi029  , \pi030  , \pi031  , \pi032  , \pi033  , \pi034  , \pi035  , \pi036  , \pi037  , \pi038  , \pi039  , \pi040  , \pi041  , \pi042  , \pi043  , \pi044  , \pi045  , \pi046  , \pi047  , \pi048  , \pi049  , \pi050  , \pi051  , \pi052  , \pi053  , \pi054  , \pi055  , \pi056  , \pi057  , \pi058  , \pi059  , \pi060  , \pi061  , \pi062  , \pi063  , \pi064  , \pi065  , \pi066  , \pi067  , \pi068  , \pi069  , \pi070  , \pi071  , \pi072  , \pi073  , \pi074  , \pi075  , \pi076  , \pi077  , \pi078  , \pi079  , \pi080  , \pi081  , \pi082  , \pi083  , \pi084  , \pi085  , \pi086  , \pi087  , \pi088  , \pi089  , \pi090  , \pi091  , \pi092  , \pi093  , \pi094  , \pi095  , \pi096  , \pi097  , \pi098  , \pi099  , \pi100  , \pi101  , \pi102  , \pi103  , \pi104  , \pi105  , \pi106  , \pi107  , \pi108  , \pi109  , \pi110  , \pi111  , \pi112  , \pi113  , \pi114  , \pi115  , \pi116  , \pi117  , \pi118  , \pi119  , \pi120  , \pi121  , \pi122  , \pi123  , \pi124  , \pi125  , \pi126  , \pi127  , \pi128  , \pi129  , \pi130  , \pi131  , \pi132  , \pi133  , \pi134  , \pi135  , \pi136  , \pi137  , \pi138  , \pi139  , \pi140  , \pi141  , \pi142  , \pi143  , \pi144  , \pi145  , \pi146  , \po000  , \po001  , \po002  , \po003  , \po004  , \po005  , \po006  , \po007  , \po008  , \po009  , \po010  , \po011  , \po012  , \po013  , \po014  , \po015  , \po016  , \po017  , \po018  , \po019  , \po020  , \po021  , \po022  , \po023  , \po024  , \po025  , \po026  , \po027  , \po028  , \po029  , \po030  , \po031  , \po032  , \po033  , \po034  , \po035  , \po036  , \po037  , \po038  , \po039  , \po040  , \po041  , \po042  , \po043  , \po044  , \po045  , \po046  , \po047  , \po048  , \po049  , \po050  , \po051  , \po052  , \po053  , \po054  , \po055  , \po056  , \po057  , \po058  , \po059  , \po060  , \po061  , \po062  , \po063  , \po064  , \po065  , \po066  , \po067  , \po068  , \po069  , \po070  , \po071  , \po072  , \po073  , \po074  , \po075  , \po076  , \po077  , \po078  , \po079  , \po080  , \po081  , \po082  , \po083  , \po084  , \po085  , \po086  , \po087  , \po088  , \po089  , \po090  , \po091  , \po092  , \po093  , \po094  , \po095  , \po096  , \po097  , \po098  , \po099  , \po100  , \po101  , \po102  , \po103  , \po104  , \po105  , \po106  , \po107  , \po108  , \po109  , \po110  , \po111  , \po112  , \po113  , \po114  , \po115  , \po116  , \po117  , \po118  , \po119  , \po120  , \po121  , \po122  , \po123  , \po124  , \po125  , \po126  , \po127  , \po128  , \po129  , \po130  , \po131  , \po132  , \po133  , \po134  , \po135  , \po136  , \po137  , \po138  , \po139  , \po140  , \po141  );
  input \pi000  ;
  input \pi001  ;
  input \pi002  ;
  input \pi003  ;
  input \pi004  ;
  input \pi005  ;
  input \pi006  ;
  input \pi007  ;
  input \pi008  ;
  input \pi009  ;
  input \pi010  ;
  input \pi011  ;
  input \pi012  ;
  input \pi013  ;
  input \pi014  ;
  input \pi015  ;
  input \pi016  ;
  input \pi017  ;
  input \pi018  ;
  input \pi019  ;
  input \pi020  ;
  input \pi021  ;
  input \pi022  ;
  input \pi023  ;
  input \pi024  ;
  input \pi025  ;
  input \pi026  ;
  input \pi027  ;
  input \pi028  ;
  input \pi029  ;
  input \pi030  ;
  input \pi031  ;
  input \pi032  ;
  input \pi033  ;
  input \pi034  ;
  input \pi035  ;
  input \pi036  ;
  input \pi037  ;
  input \pi038  ;
  input \pi039  ;
  input \pi040  ;
  input \pi041  ;
  input \pi042  ;
  input \pi043  ;
  input \pi044  ;
  input \pi045  ;
  input \pi046  ;
  input \pi047  ;
  input \pi048  ;
  input \pi049  ;
  input \pi050  ;
  input \pi051  ;
  input \pi052  ;
  input \pi053  ;
  input \pi054  ;
  input \pi055  ;
  input \pi056  ;
  input \pi057  ;
  input \pi058  ;
  input \pi059  ;
  input \pi060  ;
  input \pi061  ;
  input \pi062  ;
  input \pi063  ;
  input \pi064  ;
  input \pi065  ;
  input \pi066  ;
  input \pi067  ;
  input \pi068  ;
  input \pi069  ;
  input \pi070  ;
  input \pi071  ;
  input \pi072  ;
  input \pi073  ;
  input \pi074  ;
  input \pi075  ;
  input \pi076  ;
  input \pi077  ;
  input \pi078  ;
  input \pi079  ;
  input \pi080  ;
  input \pi081  ;
  input \pi082  ;
  input \pi083  ;
  input \pi084  ;
  input \pi085  ;
  input \pi086  ;
  input \pi087  ;
  input \pi088  ;
  input \pi089  ;
  input \pi090  ;
  input \pi091  ;
  input \pi092  ;
  input \pi093  ;
  input \pi094  ;
  input \pi095  ;
  input \pi096  ;
  input \pi097  ;
  input \pi098  ;
  input \pi099  ;
  input \pi100  ;
  input \pi101  ;
  input \pi102  ;
  input \pi103  ;
  input \pi104  ;
  input \pi105  ;
  input \pi106  ;
  input \pi107  ;
  input \pi108  ;
  input \pi109  ;
  input \pi110  ;
  input \pi111  ;
  input \pi112  ;
  input \pi113  ;
  input \pi114  ;
  input \pi115  ;
  input \pi116  ;
  input \pi117  ;
  input \pi118  ;
  input \pi119  ;
  input \pi120  ;
  input \pi121  ;
  input \pi122  ;
  input \pi123  ;
  input \pi124  ;
  input \pi125  ;
  input \pi126  ;
  input \pi127  ;
  input \pi128  ;
  input \pi129  ;
  input \pi130  ;
  input \pi131  ;
  input \pi132  ;
  input \pi133  ;
  input \pi134  ;
  input \pi135  ;
  input \pi136  ;
  input \pi137  ;
  input \pi138  ;
  input \pi139  ;
  input \pi140  ;
  input \pi141  ;
  input \pi142  ;
  input \pi143  ;
  input \pi144  ;
  input \pi145  ;
  input \pi146  ;
  output \po000  ;
  output \po001  ;
  output \po002  ;
  output \po003  ;
  output \po004  ;
  output \po005  ;
  output \po006  ;
  output \po007  ;
  output \po008  ;
  output \po009  ;
  output \po010  ;
  output \po011  ;
  output \po012  ;
  output \po013  ;
  output \po014  ;
  output \po015  ;
  output \po016  ;
  output \po017  ;
  output \po018  ;
  output \po019  ;
  output \po020  ;
  output \po021  ;
  output \po022  ;
  output \po023  ;
  output \po024  ;
  output \po025  ;
  output \po026  ;
  output \po027  ;
  output \po028  ;
  output \po029  ;
  output \po030  ;
  output \po031  ;
  output \po032  ;
  output \po033  ;
  output \po034  ;
  output \po035  ;
  output \po036  ;
  output \po037  ;
  output \po038  ;
  output \po039  ;
  output \po040  ;
  output \po041  ;
  output \po042  ;
  output \po043  ;
  output \po044  ;
  output \po045  ;
  output \po046  ;
  output \po047  ;
  output \po048  ;
  output \po049  ;
  output \po050  ;
  output \po051  ;
  output \po052  ;
  output \po053  ;
  output \po054  ;
  output \po055  ;
  output \po056  ;
  output \po057  ;
  output \po058  ;
  output \po059  ;
  output \po060  ;
  output \po061  ;
  output \po062  ;
  output \po063  ;
  output \po064  ;
  output \po065  ;
  output \po066  ;
  output \po067  ;
  output \po068  ;
  output \po069  ;
  output \po070  ;
  output \po071  ;
  output \po072  ;
  output \po073  ;
  output \po074  ;
  output \po075  ;
  output \po076  ;
  output \po077  ;
  output \po078  ;
  output \po079  ;
  output \po080  ;
  output \po081  ;
  output \po082  ;
  output \po083  ;
  output \po084  ;
  output \po085  ;
  output \po086  ;
  output \po087  ;
  output \po088  ;
  output \po089  ;
  output \po090  ;
  output \po091  ;
  output \po092  ;
  output \po093  ;
  output \po094  ;
  output \po095  ;
  output \po096  ;
  output \po097  ;
  output \po098  ;
  output \po099  ;
  output \po100  ;
  output \po101  ;
  output \po102  ;
  output \po103  ;
  output \po104  ;
  output \po105  ;
  output \po106  ;
  output \po107  ;
  output \po108  ;
  output \po109  ;
  output \po110  ;
  output \po111  ;
  output \po112  ;
  output \po113  ;
  output \po114  ;
  output \po115  ;
  output \po116  ;
  output \po117  ;
  output \po118  ;
  output \po119  ;
  output \po120  ;
  output \po121  ;
  output \po122  ;
  output \po123  ;
  output \po124  ;
  output \po125  ;
  output \po126  ;
  output \po127  ;
  output \po128  ;
  output \po129  ;
  output \po130  ;
  output \po131  ;
  output \po132  ;
  output \po133  ;
  output \po134  ;
  output \po135  ;
  output \po136  ;
  output \po137  ;
  output \po138  ;
  output \po139  ;
  output \po140  ;
  output \po141  ;
  wire n148 , n149 , n150 , n151 , n152 , n153 , n154 , n155 , n156 , n157 , n158 , n159 , n160 , n161 , n162 , n163 , n164 , n165 , n166 , n167 , n168 , n169 , n170 , n171 , n172 , n173 , n174 , n175 , n176 , n177 , n178 , n179 , n180 , n181 , n182 , n183 , n184 , n185 , n186 , n187 , n188 , n189 , n190 , n191 , n192 , n193 , n194 , n195 , n196 , n197 , n198 , n199 , n200 , n201 , n202 , n203 , n204 , n205 , n206 , n207 , n208 , n209 , n210 , n211 , n212 , n213 , n214 , n215 , n216 , n217 , n218 , n219 , n220 , n221 , n222 , n223 , n224 , n225 , n226 , n227 , n228 , n229 , n230 , n231 , n232 , n233 , n234 , n235 , n236 , n237 , n238 , n239 , n240 , n241 , n242 , n243 , n244 , n245 , n246 , n247 , n248 , n249 , n250 , n251 , n252 , n253 , n254 , n255 , n256 , n257 , n258 , n259 , n260 , n261 , n262 , n263 , n264 , n265 , n266 , n267 , n268 , n269 , n270 , n271 , n272 , n273 , n274 , n275 , n276 , n277 , n278 , n279 , n280 , n281 , n282 , n283 , n284 , n285 , n286 , n287 , n288 , n289 , n290 , n291 , n292 , n293 , n294 , n295 , n296 , n297 , n298 , n299 , n300 , n301 , n302 , n303 , n304 , n305 , n306 , n307 , n308 , n309 , n310 , n311 , n312 , n313 , n314 , n315 , n316 , n317 , n318 , n319 , n320 , n321 , n322 , n323 , n324 , n325 , n326 , n327 , n328 , n329 , n330 , n331 , n332 , n333 , n334 , n335 , n336 , n337 , n338 , n339 , n340 , n341 , n342 , n343 , n344 , n345 , n346 , n347 , n348 , n349 , n350 , n351 , n352 , n353 , n354 , n355 , n356 , n357 , n358 , n359 , n360 , n361 , n362 , n363 , n364 , n365 , n366 , n367 , n368 , n369 , n370 , n371 , n372 , n373 , n374 , n375 , n376 , n377 , n378 , n379 , n380 , n381 , n382 , n383 , n384 , n385 , n386 , n387 , n388 , n389 , n390 , n391 , n392 , n393 , n394 , n395 , n396 , n397 , n398 , n399 , n400 , n401 , n402 , n403 , n404 , n405 , n406 , n407 , n408 , n409 , n410 , n411 , n412 , n413 , n414 , n415 , n416 , n417 , n418 , n419 , n420 , n421 , n422 , n423 , n424 , n425 , n426 , n427 , n428 , n429 , n430 , n431 , n432 , n433 , n434 , n435 , n436 , n437 , n438 , n439 , n440 , n441 , n442 , n443 , n444 , n445 , n446 , n447 , n448 , n449 , n450 , n451 , n452 , n453 , n454 , n455 , n456 , n457 , n458 , n459 , n460 , n461 , n462 , n463 , n464 , n465 , n466 , n467 , n468 , n469 , n470 , n471 , n472 , n473 , n474 , n475 , n476 , n477 , n478 , n479 , n480 , n481 , n482 , n483 , n484 , n485 , n486 , n487 , n488 , n489 , n490 , n491 , n492 , n493 , n494 , n495 , n496 , n497 , n498 , n499 , n500 , n501 , n502 , n503 , n504 , n505 , n506 , n507 , n508 , n509 , n510 , n511 , n512 , n513 , n514 , n515 , n516 , n517 , n518 , n519 , n520 , n521 , n522 , n523 , n524 , n525 , n526 , n527 , n528 , n529 , n530 , n531 , n532 , n533 , n534 , n535 , n536 , n537 , n538 , n539 , n540 , n541 , n542 , n543 , n544 , n545 , n546 , n547 , n548 , n549 , n550 , n551 , n552 , n553 , n554 , n555 , n556 , n557 , n558 , n559 , n560 , n561 , n562 , n563 , n564 , n565 , n566 , n567 , n568 , n569 , n570 , n571 , n572 , n573 , n574 , n575 , n576 , n577 , n578 , n579 , n580 , n581 , n582 , n583 , n584 , n585 , n586 , n587 , n588 , n589 , n590 , n591 , n592 , n593 , n594 , n595 , n596 , n597 , n598 , n599 , n600 , n601 , n602 , n603 , n604 , n605 , n606 , n607 , n608 , n609 , n610 , n611 , n612 , n613 , n614 , n615 , n616 , n617 , n618 , n619 , n620 , n621 , n622 , n623 , n624 , n625 , n626 , n627 , n628 , n629 , n630 , n631 , n632 , n633 , n634 , n635 , n636 , n637 , n638 , n639 , n640 , n641 , n642 , n643 , n644 , n645 , n646 , n647 , n648 , n649 , n650 , n651 , n652 , n653 , n654 , n655 , n656 , n657 , n658 , n659 , n660 , n661 , n662 , n663 , n664 , n665 , n666 , n667 , n668 , n669 , n670 , n671 , n672 , n673 , n674 , n675 , n676 , n677 , n678 , n679 , n680 , n681 , n682 , n683 , n684 , n685 , n686 , n687 , n688 , n689 , n690 , n691 , n692 , n693 , n694 , n695 , n696 , n697 , n698 , n699 , n700 , n701 , n702 , n703 , n704 , n705 , n706 , n707 , n708 , n709 , n710 , n711 , n712 , n713 , n714 , n715 , n716 , n717 , n718 , n719 , n720 , n721 , n722 , n723 , n724 , n725 , n726 , n727 , n728 , n729 , n730 , n731 , n732 , n733 , n734 , n735 , n736 , n737 , n738 , n739 , n740 , n741 , n742 , n743 , n744 , n745 , n746 , n747 , n748 , n749 , n750 , n751 , n752 , n753 , n754 , n755 , n756 , n757 , n758 , n759 , n760 , n761 , n762 , n763 , n764 , n765 , n766 , n767 , n768 , n769 , n770 , n771 , n772 , n773 , n774 , n775 , n776 , n777 , n778 , n779 , n780 , n781 , n782 , n783 , n784 , n785 , n786 , n787 , n788 , n789 , n790 , n791 , n792 , n793 , n794 , n795 , n796 , n797 , n798 , n799 , n800 , n801 , n802 , n803 , n804 , n805 , n806 , n807 , n808 , n809 , n810 , n811 , n812 , n813 , n814 , n815 , n816 , n817 , n818 , n819 , n820 , n821 , n822 , n823 , n824 , n825 , n826 , n827 , n828 , n829 , n830 , n831 , n832 , n833 , n834 , n835 , n836 , n837 , n838 , n839 , n840 , n841 , n842 , n843 , n844 , n845 , n846 , n847 , n848 , n849 , n850 , n851 , n852 , n853 , n854 , n855 , n856 , n857 , n858 , n859 , n860 , n861 , n862 , n863 , n864 , n865 , n866 , n867 , n868 , n869 , n870 , n871 , n872 , n873 , n874 , n875 , n876 , n877 , n878 , n879 , n880 , n881 , n882 , n883 , n884 , n885 , n886 , n887 , n888 , n889 , n890 , n891 , n892 , n893 , n894 , n895 , n896 , n897 , n898 , n899 , n900 , n901 , n902 , n903 , n904 , n905 , n906 , n907 , n908 , n909 , n910 , n911 , n912 , n913 , n914 , n915 , n916 , n917 , n918 , n919 , n920 , n921 , n922 , n923 , n924 , n925 , n926 , n927 , n928 , n929 , n930 , n931 , n932 , n933 , n934 , n935 , n936 , n937 , n938 , n939 , n940 , n941 , n942 , n943 , n944 , n945 , n946 , n947 , n948 , n949 , n950 , n951 , n952 , n953 , n954 , n955 , n956 , n957 , n958 , n959 , n960 , n961 , n962 , n963 , n964 , n965 , n966 , n967 , n968 , n969 , n970 , n971 , n972 , n973 , n974 , n975 , n976 , n977 , n978 , n979 , n980 , n981 , n982 , n983 , n984 , n985 , n986 , n987 , n988 , n989 , n990 , n991 , n992 , n993 , n994 , n995 , n996 , n997 , n998 , n999 , n1000 , n1001 , n1002 , n1003 , n1004 , n1005 , n1006 , n1007 , n1008 , n1009 , n1010 , n1011 , n1012 , n1013 , n1014 , n1015 , n1016 , n1017 , n1018 , n1019 , n1020 , n1021 , n1022 , n1023 , n1024 , n1025 , n1026 , n1027 , n1028 , n1029 , n1030 , n1031 , n1032 , n1033 , n1034 , n1035 , n1036 , n1037 , n1038 , n1039 , n1040 , n1041 , n1042 , n1043 , n1044 , n1045 , n1046 , n1047 , n1048 , n1049 , n1050 , n1051 , n1052 , n1053 , n1054 , n1055 , n1056 , n1057 , n1058 , n1059 , n1060 , n1061 , n1062 , n1063 , n1064 , n1065 , n1066 , n1067 , n1068 , n1069 , n1070 , n1071 , n1072 , n1073 , n1074 , n1075 , n1076 , n1077 , n1078 , n1079 , n1080 , n1081 , n1082 , n1083 , n1084 , n1085 , n1086 , n1087 , n1088 , n1089 , n1090 , n1091 , n1092 , n1093 , n1094 , n1095 , n1096 , n1097 , n1098 , n1099 , n1100 , n1101 , n1102 , n1103 , n1104 , n1105 , n1106 , n1107 , n1108 , n1109 , n1110 , n1111 , n1112 , n1113 , n1114 , n1115 , n1116 , n1117 , n1118 , n1119 , n1120 , n1121 , n1122 , n1123 , n1124 , n1125 , n1126 , n1127 , n1128 , n1129 , n1130 , n1131 , n1132 , n1133 , n1134 , n1135 , n1136 , n1137 , n1138 , n1139 , n1140 , n1141 , n1142 , n1143 , n1144 , n1145 , n1146 , n1147 , n1148 , n1149 , n1150 , n1151 , n1152 , n1153 , n1154 , n1155 , n1156 , n1157 , n1158 , n1159 , n1160 , n1161 , n1162 , n1163 , n1164 , n1165 , n1166 , n1167 , n1168 , n1169 , n1170 , n1171 , n1172 , n1173 , n1174 , n1175 , n1176 , n1177 , n1178 , n1179 , n1180 , n1181 , n1182 , n1183 , n1184 , n1185 , n1186 , n1187 , n1188 , n1189 , n1190 , n1191 , n1192 , n1193 , n1194 , n1195 , n1196 , n1197 , n1198 , n1199 , n1200 , n1201 , n1202 , n1203 , n1204 , n1205 , n1206 , n1207 , n1208 , n1209 , n1210 , n1211 , n1212 , n1213 , n1214 , n1215 , n1216 , n1217 , n1218 , n1219 , n1220 , n1221 , n1222 , n1223 , n1224 , n1225 , n1226 , n1227 , n1228 , n1229 , n1230 , n1231 , n1232 , n1233 , n1234 , n1235 , n1236 , n1237 , n1238 , n1239 , n1240 , n1241 , n1242 , n1243 , n1244 , n1245 , n1246 , n1247 , n1248 , n1249 , n1250 , n1251 , n1252 , n1253 , n1254 , n1255 , n1256 , n1257 , n1258 , n1259 , n1260 , n1261 , n1262 , n1263 , n1264 , n1265 , n1266 , n1267 , n1268 , n1269 , n1270 , n1271 , n1272 , n1273 , n1274 , n1275 , n1276 , n1277 , n1278 , n1279 , n1280 , n1281 , n1282 , n1283 , n1284 , n1285 , n1286 , n1287 , n1288 , n1289 , n1290 , n1291 , n1292 , n1293 , n1294 , n1295 , n1296 , n1297 , n1298 , n1299 , n1300 , n1301 , n1302 , n1303 , n1304 , n1305 , n1306 , n1307 , n1308 , n1309 , n1310 , n1311 , n1312 , n1313 , n1314 , n1315 , n1316 , n1317 , n1318 , n1319 , n1320 , n1321 , n1322 , n1323 , n1324 , n1325 , n1326 , n1327 , n1328 , n1329 , n1330 , n1331 , n1332 , n1333 , n1334 , n1335 , n1336 , n1337 , n1338 , n1339 , n1340 , n1341 , n1342 , n1343 , n1344 , n1345 , n1346 , n1347 , n1348 , n1349 , n1350 , n1351 , n1352 , n1353 , n1354 , n1355 , n1356 , n1357 , n1358 , n1359 , n1360 , n1361 , n1362 , n1363 , n1364 , n1365 , n1366 , n1367 , n1368 , n1369 , n1370 , n1371 , n1372 , n1373 , n1374 , n1375 ;
  assign n148 = ~\pi003  & ~\pi129  ;
  assign n149 = ~\pi000  & ~\pi054  ;
  assign n150 = ~\pi004  & ~\pi019  ;
  assign n151 = ~\pi016  & n150 ;
  assign n152 = ~\pi017  & ~\pi018  ;
  assign n153 = n151 & n152 ;
  assign n154 = ~\pi006  & ~\pi012  ;
  assign n155 = ~\pi005  & ~\pi022  ;
  assign n156 = n154 & n155 ;
  assign n157 = n153 & n156 ;
  assign n158 = ~\pi007  & ~\pi013  ;
  assign n159 = ~\pi014  & n158 ;
  assign n160 = ~\pi008  & ~\pi021  ;
  assign n161 = ~\pi009  & ~\pi011  ;
  assign n162 = n160 & n161 ;
  assign n163 = n159 & n162 ;
  assign n164 = ~\pi000  & n163 ;
  assign n165 = n157 & n164 ;
  assign n166 = ~n149 & ~n165 ;
  assign n167 = \pi054  & n161 ;
  assign n168 = \pi054  & ~\pi056  ;
  assign n169 = n155 & n168 ;
  assign n170 = ~n167 & ~n169 ;
  assign n171 = n166 & n170 ;
  assign n172 = n158 & n160 ;
  assign n173 = \pi010  & ~\pi014  ;
  assign n174 = n172 & n173 ;
  assign n175 = n157 & n174 ;
  assign n176 = \pi014  & ~n172 ;
  assign n177 = ~\pi007  & n160 ;
  assign n178 = \pi008  & \pi021  ;
  assign n179 = ~\pi013  & ~n178 ;
  assign n180 = ~n177 & ~n179 ;
  assign n181 = ~\pi010  & ~n180 ;
  assign n182 = ~n176 & n181 ;
  assign n183 = \pi007  & ~n160 ;
  assign n184 = ~n172 & ~n183 ;
  assign n185 = ~\pi014  & ~n184 ;
  assign n186 = n157 & ~n185 ;
  assign n187 = n182 & n186 ;
  assign n188 = ~n175 & ~n187 ;
  assign n189 = ~\pi056  & ~n155 ;
  assign n190 = n161 & ~n189 ;
  assign n191 = n166 & n190 ;
  assign n192 = n188 & n191 ;
  assign n193 = ~n171 & ~n192 ;
  assign n194 = n148 & n193 ;
  assign n195 = ~\pi017  & \pi054  ;
  assign n196 = ~\pi001  & ~n195 ;
  assign n197 = ~\pi010  & ~\pi022  ;
  assign n198 = ~\pi013  & n197 ;
  assign n199 = ~\pi011  & n160 ;
  assign n200 = ~\pi014  & ~\pi018  ;
  assign n201 = n199 & n200 ;
  assign n202 = n198 & n201 ;
  assign n203 = ~\pi005  & ~\pi006  ;
  assign n204 = ~\pi007  & ~\pi012  ;
  assign n205 = n203 & n204 ;
  assign n206 = n151 & n205 ;
  assign n207 = ~\pi001  & n206 ;
  assign n208 = n202 & n207 ;
  assign n209 = ~n196 & ~n208 ;
  assign n210 = n148 & ~n209 ;
  assign n211 = ~\pi009  & ~\pi013  ;
  assign n212 = n205 & n211 ;
  assign n213 = n153 & n199 ;
  assign n214 = \pi013  & ~n205 ;
  assign n215 = ~\pi022  & \pi054  ;
  assign n216 = ~\pi010  & ~\pi014  ;
  assign n217 = n215 & n216 ;
  assign n218 = ~n214 & n217 ;
  assign n219 = n213 & n218 ;
  assign n220 = ~n212 & n219 ;
  assign n221 = ~\pi013  & n205 ;
  assign n222 = ~\pi005  & ~\pi007  ;
  assign n223 = ~n154 & ~n222 ;
  assign n224 = ~n203 & ~n204 ;
  assign n225 = ~\pi009  & ~n224 ;
  assign n226 = ~n223 & n225 ;
  assign n227 = ~n221 & ~n226 ;
  assign n228 = n148 & ~n227 ;
  assign n229 = n220 & n228 ;
  assign n230 = ~n210 & ~n229 ;
  assign n231 = \pi122  & \pi127  ;
  assign n232 = ~\pi082  & ~n231 ;
  assign n233 = ~\pi065  & n232 ;
  assign n234 = ~\pi042  & ~\pi044  ;
  assign n235 = ~\pi038  & ~\pi040  ;
  assign n236 = n234 & n235 ;
  assign n237 = ~\pi046  & ~\pi050  ;
  assign n238 = n236 & n237 ;
  assign n239 = ~\pi041  & ~\pi043  ;
  assign n240 = ~\pi047  & n239 ;
  assign n241 = ~\pi048  & n240 ;
  assign n242 = n238 & n241 ;
  assign n243 = ~\pi002  & ~\pi020  ;
  assign n244 = ~\pi015  & ~\pi049  ;
  assign n245 = n243 & n244 ;
  assign n246 = ~\pi024  & ~\pi045  ;
  assign n247 = ~n231 & n246 ;
  assign n248 = n245 & n247 ;
  assign n249 = ~\pi065  & n248 ;
  assign n250 = n242 & n249 ;
  assign n251 = ~n233 & ~n250 ;
  assign n252 = ~\pi082  & n231 ;
  assign n253 = \pi002  & n252 ;
  assign n254 = ~\pi045  & ~\pi048  ;
  assign n255 = n240 & n254 ;
  assign n256 = n238 & n255 ;
  assign n257 = ~\pi020  & ~\pi024  ;
  assign n258 = n244 & n257 ;
  assign n259 = n256 & n258 ;
  assign n260 = \pi002  & \pi082  ;
  assign n261 = ~n259 & n260 ;
  assign n262 = ~n253 & ~n261 ;
  assign n263 = n251 & n262 ;
  assign n264 = ~\pi129  & ~n263 ;
  assign n265 = \pi000  & ~\pi113  ;
  assign n266 = ~\pi123  & n265 ;
  assign n267 = ~\pi129  & n266 ;
  assign n268 = ~\pi009  & ~\pi014  ;
  assign n269 = n204 & n268 ;
  assign n270 = n198 & n269 ;
  assign n271 = n203 & n270 ;
  assign n272 = n213 & n271 ;
  assign n273 = ~\pi061  & ~\pi118  ;
  assign n274 = ~\pi129  & n273 ;
  assign n275 = ~n272 & n274 ;
  assign n276 = ~n267 & ~n275 ;
  assign n277 = \pi004  & ~\pi054  ;
  assign n278 = \pi054  & n199 ;
  assign n279 = n153 & n278 ;
  assign n280 = ~\pi022  & n173 ;
  assign n281 = n212 & n280 ;
  assign n282 = n279 & n281 ;
  assign n283 = ~n277 & ~n282 ;
  assign n284 = n148 & ~n283 ;
  assign n285 = \pi005  & ~\pi054  ;
  assign n286 = n198 & n268 ;
  assign n287 = ~\pi011  & ~\pi017  ;
  assign n288 = n160 & n287 ;
  assign n289 = ~\pi059  & n288 ;
  assign n290 = n286 & n289 ;
  assign n291 = ~\pi016  & \pi054  ;
  assign n292 = n205 & n291 ;
  assign n293 = ~\pi018  & ~\pi029  ;
  assign n294 = n150 & n293 ;
  assign n295 = ~\pi025  & \pi028  ;
  assign n296 = n294 & n295 ;
  assign n297 = n292 & n296 ;
  assign n298 = n290 & n297 ;
  assign n299 = ~n285 & ~n298 ;
  assign n300 = n148 & ~n299 ;
  assign n301 = \pi006  & ~\pi054  ;
  assign n302 = \pi025  & ~\pi028  ;
  assign n303 = n294 & n302 ;
  assign n304 = n292 & n303 ;
  assign n305 = n290 & n304 ;
  assign n306 = ~n301 & ~n305 ;
  assign n307 = n148 & ~n306 ;
  assign n308 = \pi007  & ~\pi054  ;
  assign n309 = n150 & n291 ;
  assign n310 = n203 & n309 ;
  assign n311 = n270 & n310 ;
  assign n312 = ~\pi011  & n152 ;
  assign n313 = \pi008  & ~\pi021  ;
  assign n314 = n312 & n313 ;
  assign n315 = n311 & n314 ;
  assign n316 = ~n308 & ~n315 ;
  assign n317 = n148 & ~n316 ;
  assign n318 = \pi008  & ~\pi054  ;
  assign n319 = ~\pi008  & \pi021  ;
  assign n320 = n312 & n319 ;
  assign n321 = n311 & n320 ;
  assign n322 = ~n318 & ~n321 ;
  assign n323 = n148 & ~n322 ;
  assign n324 = \pi009  & ~\pi054  ;
  assign n325 = n152 & n160 ;
  assign n326 = n221 & n325 ;
  assign n327 = n197 & n309 ;
  assign n328 = \pi011  & n268 ;
  assign n329 = n327 & n328 ;
  assign n330 = n326 & n329 ;
  assign n331 = ~n324 & ~n330 ;
  assign n332 = n148 & ~n331 ;
  assign n333 = \pi010  & ~\pi054  ;
  assign n334 = n148 & n333 ;
  assign n335 = ~\pi009  & n325 ;
  assign n336 = n327 & n335 ;
  assign n337 = ~\pi011  & \pi014  ;
  assign n338 = ~\pi013  & n337 ;
  assign n339 = n205 & n338 ;
  assign n340 = n148 & n339 ;
  assign n341 = n336 & n340 ;
  assign n342 = ~n334 & ~n341 ;
  assign n343 = \pi011  & ~\pi054  ;
  assign n344 = \pi022  & n161 ;
  assign n345 = n216 & n344 ;
  assign n346 = n309 & n345 ;
  assign n347 = n326 & n346 ;
  assign n348 = ~n343 & ~n347 ;
  assign n349 = n148 & ~n348 ;
  assign n350 = \pi012  & ~\pi054  ;
  assign n351 = n148 & n350 ;
  assign n352 = \pi018  & n288 ;
  assign n353 = n148 & n352 ;
  assign n354 = n311 & n353 ;
  assign n355 = ~n351 & ~n354 ;
  assign n356 = \pi013  & ~\pi054  ;
  assign n357 = n148 & n356 ;
  assign n358 = ~\pi018  & n203 ;
  assign n359 = n309 & n358 ;
  assign n360 = n270 & n359 ;
  assign n361 = ~\pi025  & ~\pi028  ;
  assign n362 = \pi029  & ~\pi059  ;
  assign n363 = n361 & n362 ;
  assign n364 = n288 & n363 ;
  assign n365 = n148 & n364 ;
  assign n366 = n360 & n365 ;
  assign n367 = ~n357 & ~n366 ;
  assign n368 = \pi014  & ~\pi054  ;
  assign n369 = n148 & n368 ;
  assign n370 = ~\pi011  & \pi013  ;
  assign n371 = n217 & n370 ;
  assign n372 = n206 & n371 ;
  assign n373 = n148 & n335 ;
  assign n374 = n372 & n373 ;
  assign n375 = ~n369 & ~n374 ;
  assign n376 = ~\pi024  & n244 ;
  assign n377 = ~n243 & n376 ;
  assign n378 = n256 & n377 ;
  assign n379 = \pi082  & n378 ;
  assign n380 = ~\pi024  & ~\pi049  ;
  assign n381 = n256 & n380 ;
  assign n382 = \pi015  & \pi082  ;
  assign n383 = ~n381 & n382 ;
  assign n384 = ~n379 & ~n383 ;
  assign n385 = \pi015  & ~\pi082  ;
  assign n386 = n231 & n385 ;
  assign n387 = ~\pi070  & ~n231 ;
  assign n388 = ~n386 & ~n387 ;
  assign n389 = n256 & n376 ;
  assign n390 = \pi082  & ~n386 ;
  assign n391 = ~n389 & n390 ;
  assign n392 = ~n388 & ~n391 ;
  assign n393 = n384 & ~n392 ;
  assign n394 = ~\pi129  & ~n393 ;
  assign n395 = \pi016  & ~\pi054  ;
  assign n396 = ~\pi005  & \pi006  ;
  assign n397 = n270 & n396 ;
  assign n398 = n279 & n397 ;
  assign n399 = ~n395 & ~n398 ;
  assign n400 = n148 & ~n399 ;
  assign n401 = \pi017  & ~\pi054  ;
  assign n402 = n148 & n401 ;
  assign n403 = ~\pi029  & \pi054  ;
  assign n404 = \pi059  & n403 ;
  assign n405 = n361 & n404 ;
  assign n406 = n148 & n405 ;
  assign n407 = n272 & n406 ;
  assign n408 = ~n402 & ~n407 ;
  assign n409 = \pi018  & ~\pi054  ;
  assign n410 = n286 & n288 ;
  assign n411 = \pi054  & n205 ;
  assign n412 = \pi016  & ~\pi018  ;
  assign n413 = n150 & n412 ;
  assign n414 = n411 & n413 ;
  assign n415 = n410 & n414 ;
  assign n416 = ~n409 & ~n415 ;
  assign n417 = n148 & ~n416 ;
  assign n418 = \pi019  & ~\pi054  ;
  assign n419 = n148 & n418 ;
  assign n420 = ~\pi011  & \pi017  ;
  assign n421 = n160 & n420 ;
  assign n422 = n148 & n421 ;
  assign n423 = n360 & n422 ;
  assign n424 = ~n419 & ~n423 ;
  assign n425 = \pi020  & \pi082  ;
  assign n426 = ~n389 & n425 ;
  assign n427 = ~\pi020  & n260 ;
  assign n428 = n389 & n427 ;
  assign n429 = ~n426 & ~n428 ;
  assign n430 = \pi020  & ~\pi082  ;
  assign n431 = n231 & n430 ;
  assign n432 = ~\pi071  & ~n231 ;
  assign n433 = ~n431 & ~n432 ;
  assign n434 = \pi082  & ~n431 ;
  assign n435 = ~n259 & n434 ;
  assign n436 = ~n433 & ~n435 ;
  assign n437 = n429 & ~n436 ;
  assign n438 = ~\pi129  & ~n437 ;
  assign n439 = \pi021  & ~\pi054  ;
  assign n440 = ~\pi004  & ~\pi016  ;
  assign n441 = ~\pi018  & \pi019  ;
  assign n442 = n440 & n441 ;
  assign n443 = n411 & n442 ;
  assign n444 = n410 & n443 ;
  assign n445 = ~n439 & ~n444 ;
  assign n446 = n148 & ~n445 ;
  assign n447 = \pi022  & ~\pi054  ;
  assign n448 = n148 & n447 ;
  assign n449 = \pi005  & ~\pi011  ;
  assign n450 = n154 & n449 ;
  assign n451 = n159 & n450 ;
  assign n452 = n148 & n451 ;
  assign n453 = n336 & n452 ;
  assign n454 = ~n448 & ~n453 ;
  assign n455 = ~\pi023  & \pi055  ;
  assign n456 = \pi061  & ~\pi129  ;
  assign n457 = ~n455 & n456 ;
  assign n458 = \pi063  & ~n231 ;
  assign n459 = ~\pi082  & n458 ;
  assign n460 = n245 & n458 ;
  assign n461 = n256 & n460 ;
  assign n462 = ~n459 & ~n461 ;
  assign n463 = \pi082  & ~n245 ;
  assign n464 = n231 & ~n463 ;
  assign n465 = ~\pi024  & n464 ;
  assign n466 = ~\pi024  & \pi082  ;
  assign n467 = ~n256 & n466 ;
  assign n468 = ~n465 & ~n467 ;
  assign n469 = \pi082  & n237 ;
  assign n470 = n236 & n469 ;
  assign n471 = \pi024  & ~\pi045  ;
  assign n472 = ~\pi048  & n471 ;
  assign n473 = n240 & n472 ;
  assign n474 = n470 & n473 ;
  assign n475 = ~\pi129  & ~n474 ;
  assign n476 = n468 & n475 ;
  assign n477 = n462 & n476 ;
  assign n478 = ~\pi053  & \pi058  ;
  assign n479 = \pi053  & ~\pi058  ;
  assign n480 = ~n478 & ~n479 ;
  assign n481 = \pi053  & n480 ;
  assign n482 = ~\pi096  & ~\pi110  ;
  assign n483 = ~\pi085  & ~n482 ;
  assign n484 = \pi085  & ~\pi116  ;
  assign n485 = \pi100  & ~n484 ;
  assign n486 = ~n483 & n485 ;
  assign n487 = \pi025  & n484 ;
  assign n488 = ~n486 & ~n487 ;
  assign n489 = ~\pi027  & ~n488 ;
  assign n490 = ~\pi026  & n489 ;
  assign n491 = \pi025  & ~\pi116  ;
  assign n492 = ~\pi039  & ~\pi052  ;
  assign n493 = ~\pi051  & \pi116  ;
  assign n494 = n492 & n493 ;
  assign n495 = ~n491 & ~n494 ;
  assign n496 = \pi027  & ~n495 ;
  assign n497 = ~\pi051  & ~\pi052  ;
  assign n498 = ~\pi039  & n497 ;
  assign n499 = \pi027  & ~n498 ;
  assign n500 = \pi025  & \pi110  ;
  assign n501 = ~\pi095  & ~\pi100  ;
  assign n502 = \pi025  & ~\pi097  ;
  assign n503 = n501 & n502 ;
  assign n504 = ~n500 & ~n503 ;
  assign n505 = ~n499 & ~n504 ;
  assign n506 = ~n496 & ~n505 ;
  assign n507 = ~\pi026  & ~\pi085  ;
  assign n508 = ~n506 & n507 ;
  assign n509 = ~n490 & ~n508 ;
  assign n510 = \pi026  & ~\pi085  ;
  assign n511 = ~n494 & n510 ;
  assign n512 = ~\pi025  & ~\pi116  ;
  assign n513 = ~\pi027  & ~n512 ;
  assign n514 = n511 & n513 ;
  assign n515 = n480 & ~n514 ;
  assign n516 = n509 & n515 ;
  assign n517 = ~n481 & ~n516 ;
  assign n518 = ~\pi053  & ~\pi058  ;
  assign n519 = n148 & n518 ;
  assign n520 = ~\pi026  & ~\pi027  ;
  assign n521 = ~\pi085  & n520 ;
  assign n522 = n148 & n491 ;
  assign n523 = n521 & n522 ;
  assign n524 = ~n519 & ~n523 ;
  assign n525 = n517 & ~n524 ;
  assign n526 = \pi026  & \pi116  ;
  assign n527 = n486 & ~n526 ;
  assign n528 = ~n511 & ~n527 ;
  assign n529 = ~\pi027  & n518 ;
  assign n530 = n148 & n529 ;
  assign n531 = ~n528 & n530 ;
  assign n532 = \pi027  & ~\pi085  ;
  assign n533 = ~n494 & n532 ;
  assign n534 = \pi085  & \pi116  ;
  assign n535 = ~\pi085  & \pi095  ;
  assign n536 = n482 & n535 ;
  assign n537 = ~n534 & ~n536 ;
  assign n538 = \pi027  & \pi116  ;
  assign n539 = ~\pi100  & ~n538 ;
  assign n540 = ~n537 & n539 ;
  assign n541 = ~n533 & ~n540 ;
  assign n542 = ~\pi026  & n148 ;
  assign n543 = n518 & n542 ;
  assign n544 = ~n541 & n543 ;
  assign n545 = \pi053  & ~\pi116  ;
  assign n546 = \pi028  & n545 ;
  assign n547 = n521 & n546 ;
  assign n548 = ~\pi058  & n547 ;
  assign n549 = \pi026  & \pi027  ;
  assign n550 = ~n520 & ~n549 ;
  assign n551 = ~\pi116  & n550 ;
  assign n552 = \pi028  & n551 ;
  assign n553 = ~\pi026  & ~n498 ;
  assign n554 = ~\pi027  & ~\pi051  ;
  assign n555 = n492 & n554 ;
  assign n556 = ~n553 & ~n555 ;
  assign n557 = ~\pi097  & n501 ;
  assign n558 = ~\pi110  & ~n557 ;
  assign n559 = \pi028  & ~n558 ;
  assign n560 = ~n556 & n559 ;
  assign n561 = ~n552 & ~n560 ;
  assign n562 = ~\pi026  & \pi095  ;
  assign n563 = ~\pi100  & n562 ;
  assign n564 = n482 & n563 ;
  assign n565 = \pi026  & n494 ;
  assign n566 = ~n564 & ~n565 ;
  assign n567 = ~\pi027  & ~n566 ;
  assign n568 = ~\pi026  & n538 ;
  assign n569 = ~n498 & n568 ;
  assign n570 = ~\pi085  & ~n569 ;
  assign n571 = ~n567 & n570 ;
  assign n572 = n561 & n571 ;
  assign n573 = ~\pi053  & ~\pi085  ;
  assign n574 = ~\pi028  & ~\pi116  ;
  assign n575 = n520 & ~n574 ;
  assign n576 = \pi100  & \pi116  ;
  assign n577 = ~\pi053  & ~n576 ;
  assign n578 = n575 & n577 ;
  assign n579 = ~n573 & ~n578 ;
  assign n580 = ~\pi058  & ~n579 ;
  assign n581 = ~n572 & n580 ;
  assign n582 = ~n548 & ~n581 ;
  assign n583 = ~\pi026  & ~\pi053  ;
  assign n584 = ~\pi085  & n583 ;
  assign n585 = \pi058  & ~\pi116  ;
  assign n586 = ~\pi027  & \pi028  ;
  assign n587 = n585 & n586 ;
  assign n588 = n584 & n587 ;
  assign n589 = n582 & ~n588 ;
  assign n590 = n148 & ~n589 ;
  assign n591 = \pi029  & ~\pi116  ;
  assign n592 = n510 & n591 ;
  assign n593 = n529 & n592 ;
  assign n594 = \pi026  & ~n593 ;
  assign n595 = \pi027  & n518 ;
  assign n596 = n591 & n595 ;
  assign n597 = ~\pi085  & n596 ;
  assign n598 = \pi097  & \pi116  ;
  assign n599 = \pi058  & ~n591 ;
  assign n600 = ~n598 & n599 ;
  assign n601 = ~\pi053  & ~n600 ;
  assign n602 = n479 & n591 ;
  assign n603 = ~n601 & ~n602 ;
  assign n604 = n482 & n501 ;
  assign n605 = \pi097  & n604 ;
  assign n606 = ~\pi058  & ~n605 ;
  assign n607 = \pi029  & \pi110  ;
  assign n608 = \pi029  & ~\pi097  ;
  assign n609 = n501 & n608 ;
  assign n610 = ~n607 & ~n609 ;
  assign n611 = ~n602 & n610 ;
  assign n612 = n606 & n611 ;
  assign n613 = ~n603 & ~n612 ;
  assign n614 = ~\pi027  & ~\pi085  ;
  assign n615 = n613 & n614 ;
  assign n616 = ~n597 & ~n615 ;
  assign n617 = \pi085  & n591 ;
  assign n618 = n529 & n617 ;
  assign n619 = ~n593 & ~n618 ;
  assign n620 = n616 & n619 ;
  assign n621 = ~n594 & ~n620 ;
  assign n622 = n148 & n621 ;
  assign n623 = ~\pi030  & ~\pi109  ;
  assign n624 = ~\pi060  & \pi109  ;
  assign n625 = ~n623 & ~n624 ;
  assign n626 = ~\pi106  & ~n625 ;
  assign n627 = ~\pi088  & \pi106  ;
  assign n628 = ~\pi129  & ~n627 ;
  assign n629 = ~n626 & n628 ;
  assign n630 = ~\pi031  & ~\pi109  ;
  assign n631 = ~\pi030  & \pi109  ;
  assign n632 = ~n630 & ~n631 ;
  assign n633 = ~\pi106  & ~n632 ;
  assign n634 = ~\pi089  & \pi106  ;
  assign n635 = ~\pi129  & ~n634 ;
  assign n636 = ~n633 & n635 ;
  assign n637 = ~\pi032  & ~\pi109  ;
  assign n638 = ~\pi031  & \pi109  ;
  assign n639 = ~n637 & ~n638 ;
  assign n640 = ~\pi106  & ~n639 ;
  assign n641 = ~\pi099  & \pi106  ;
  assign n642 = ~\pi129  & ~n641 ;
  assign n643 = ~n640 & n642 ;
  assign n644 = ~\pi033  & ~\pi109  ;
  assign n645 = ~\pi032  & \pi109  ;
  assign n646 = ~n644 & ~n645 ;
  assign n647 = ~\pi106  & ~n646 ;
  assign n648 = ~\pi090  & \pi106  ;
  assign n649 = ~\pi129  & ~n648 ;
  assign n650 = ~n647 & n649 ;
  assign n651 = ~\pi034  & ~\pi109  ;
  assign n652 = ~\pi033  & \pi109  ;
  assign n653 = ~n651 & ~n652 ;
  assign n654 = ~\pi106  & ~n653 ;
  assign n655 = ~\pi091  & \pi106  ;
  assign n656 = ~\pi129  & ~n655 ;
  assign n657 = ~n654 & n656 ;
  assign n658 = ~\pi035  & ~\pi109  ;
  assign n659 = ~\pi034  & \pi109  ;
  assign n660 = ~n658 & ~n659 ;
  assign n661 = ~\pi106  & ~n660 ;
  assign n662 = ~\pi092  & \pi106  ;
  assign n663 = ~\pi129  & ~n662 ;
  assign n664 = ~n661 & n663 ;
  assign n665 = ~\pi036  & ~\pi109  ;
  assign n666 = ~\pi035  & \pi109  ;
  assign n667 = ~n665 & ~n666 ;
  assign n668 = ~\pi106  & ~n667 ;
  assign n669 = ~\pi098  & \pi106  ;
  assign n670 = ~\pi129  & ~n669 ;
  assign n671 = ~n668 & n670 ;
  assign n672 = ~\pi037  & ~\pi109  ;
  assign n673 = ~\pi036  & \pi109  ;
  assign n674 = ~n672 & ~n673 ;
  assign n675 = ~\pi106  & ~n674 ;
  assign n676 = ~\pi093  & \pi106  ;
  assign n677 = ~\pi129  & ~n676 ;
  assign n678 = ~n675 & n677 ;
  assign n679 = ~\pi024  & ~\pi048  ;
  assign n680 = ~\pi045  & n679 ;
  assign n681 = n245 & n680 ;
  assign n682 = n237 & n240 ;
  assign n683 = n681 & n682 ;
  assign n684 = \pi082  & n236 ;
  assign n685 = ~n683 & n684 ;
  assign n686 = ~\pi044  & \pi082  ;
  assign n687 = ~\pi040  & ~\pi042  ;
  assign n688 = n686 & n687 ;
  assign n689 = \pi038  & ~n232 ;
  assign n690 = ~n688 & n689 ;
  assign n691 = \pi082  & ~n236 ;
  assign n692 = ~\pi074  & ~n231 ;
  assign n693 = ~n691 & n692 ;
  assign n694 = ~n690 & ~n693 ;
  assign n695 = ~n685 & n694 ;
  assign n696 = ~\pi129  & ~n695 ;
  assign n697 = \pi109  & n497 ;
  assign n698 = \pi039  & ~n697 ;
  assign n699 = ~\pi051  & \pi109  ;
  assign n700 = n492 & n699 ;
  assign n701 = ~\pi106  & ~n700 ;
  assign n702 = ~n698 & n701 ;
  assign n703 = ~\pi129  & ~n702 ;
  assign n704 = \pi082  & ~n234 ;
  assign n705 = ~n231 & ~n704 ;
  assign n706 = ~\pi038  & n237 ;
  assign n707 = n240 & n706 ;
  assign n708 = n681 & n707 ;
  assign n709 = \pi082  & ~n704 ;
  assign n710 = ~n708 & n709 ;
  assign n711 = ~n705 & ~n710 ;
  assign n712 = ~\pi040  & n711 ;
  assign n713 = \pi073  & ~n231 ;
  assign n714 = ~\pi082  & n713 ;
  assign n715 = n234 & n713 ;
  assign n716 = n708 & n715 ;
  assign n717 = ~n714 & ~n716 ;
  assign n718 = \pi040  & ~\pi042  ;
  assign n719 = n686 & n718 ;
  assign n720 = ~\pi129  & ~n719 ;
  assign n721 = n717 & n720 ;
  assign n722 = ~n712 & n721 ;
  assign n723 = ~\pi043  & ~\pi047  ;
  assign n724 = n681 & n723 ;
  assign n725 = ~\pi041  & \pi082  ;
  assign n726 = n237 & n725 ;
  assign n727 = n236 & n726 ;
  assign n728 = ~n724 & n727 ;
  assign n729 = \pi041  & ~n232 ;
  assign n730 = ~n470 & n729 ;
  assign n731 = ~\pi041  & n237 ;
  assign n732 = n236 & n731 ;
  assign n733 = \pi082  & ~n732 ;
  assign n734 = ~\pi076  & ~n231 ;
  assign n735 = ~n733 & n734 ;
  assign n736 = ~n730 & ~n735 ;
  assign n737 = ~n728 & n736 ;
  assign n738 = ~\pi129  & ~n737 ;
  assign n739 = ~\pi072  & ~n231 ;
  assign n740 = ~n704 & n739 ;
  assign n741 = n235 & n237 ;
  assign n742 = n240 & n741 ;
  assign n743 = n681 & n742 ;
  assign n744 = n709 & ~n743 ;
  assign n745 = ~n740 & ~n744 ;
  assign n746 = \pi042  & ~n686 ;
  assign n747 = ~n232 & n746 ;
  assign n748 = n745 & ~n747 ;
  assign n749 = ~\pi129  & ~n748 ;
  assign n750 = ~\pi047  & n681 ;
  assign n751 = n237 & n239 ;
  assign n752 = n236 & n751 ;
  assign n753 = \pi082  & n752 ;
  assign n754 = ~n750 & n753 ;
  assign n755 = \pi043  & ~n232 ;
  assign n756 = ~n727 & n755 ;
  assign n757 = \pi082  & ~n752 ;
  assign n758 = ~\pi077  & ~n231 ;
  assign n759 = ~n757 & n758 ;
  assign n760 = ~n756 & ~n759 ;
  assign n761 = ~n754 & n760 ;
  assign n762 = ~\pi129  & ~n761 ;
  assign n763 = ~\pi067  & ~n231 ;
  assign n764 = \pi044  & n231 ;
  assign n765 = ~n763 & ~n764 ;
  assign n766 = ~\pi082  & n765 ;
  assign n767 = ~\pi042  & n765 ;
  assign n768 = n743 & n767 ;
  assign n769 = ~n766 & ~n768 ;
  assign n770 = \pi044  & \pi082  ;
  assign n771 = ~\pi129  & ~n770 ;
  assign n772 = n769 & n771 ;
  assign n773 = \pi045  & n252 ;
  assign n774 = \pi045  & \pi082  ;
  assign n775 = ~n242 & n774 ;
  assign n776 = ~n773 & ~n775 ;
  assign n777 = \pi082  & ~n256 ;
  assign n778 = ~\pi024  & n245 ;
  assign n779 = \pi082  & ~n778 ;
  assign n780 = ~\pi068  & ~n231 ;
  assign n781 = ~n779 & ~n780 ;
  assign n782 = ~n777 & ~n781 ;
  assign n783 = n776 & ~n782 ;
  assign n784 = ~\pi129  & ~n783 ;
  assign n785 = ~\pi075  & ~\pi082  ;
  assign n786 = ~n231 & n785 ;
  assign n787 = ~\pi050  & \pi082  ;
  assign n788 = n236 & n787 ;
  assign n789 = \pi046  & ~n232 ;
  assign n790 = ~n788 & n789 ;
  assign n791 = ~n786 & ~n790 ;
  assign n792 = ~\pi129  & ~n791 ;
  assign n793 = ~\pi075  & ~n231 ;
  assign n794 = ~\pi082  & ~n793 ;
  assign n795 = n240 & ~n793 ;
  assign n796 = n681 & n795 ;
  assign n797 = ~n794 & ~n796 ;
  assign n798 = ~\pi129  & n238 ;
  assign n799 = n797 & n798 ;
  assign n800 = ~n792 & ~n799 ;
  assign n801 = \pi082  & ~n681 ;
  assign n802 = ~\pi064  & ~n231 ;
  assign n803 = ~n801 & ~n802 ;
  assign n804 = n238 & n240 ;
  assign n805 = \pi082  & ~n804 ;
  assign n806 = ~n803 & ~n805 ;
  assign n807 = \pi047  & n252 ;
  assign n808 = \pi047  & \pi082  ;
  assign n809 = ~n752 & n808 ;
  assign n810 = ~n807 & ~n809 ;
  assign n811 = ~n806 & n810 ;
  assign n812 = ~\pi129  & ~n811 ;
  assign n813 = ~\pi082  & ~n252 ;
  assign n814 = n240 & ~n252 ;
  assign n815 = n238 & n814 ;
  assign n816 = ~n813 & ~n815 ;
  assign n817 = \pi048  & n816 ;
  assign n818 = \pi082  & ~n242 ;
  assign n819 = n245 & n246 ;
  assign n820 = \pi082  & ~n819 ;
  assign n821 = ~\pi062  & ~n231 ;
  assign n822 = ~n820 & ~n821 ;
  assign n823 = ~n818 & ~n822 ;
  assign n824 = ~n817 & ~n823 ;
  assign n825 = ~\pi129  & ~n824 ;
  assign n826 = ~n252 & ~n463 ;
  assign n827 = ~\pi024  & ~n252 ;
  assign n828 = n256 & n827 ;
  assign n829 = ~n826 & ~n828 ;
  assign n830 = \pi049  & n829 ;
  assign n831 = \pi082  & ~n381 ;
  assign n832 = ~\pi069  & ~n231 ;
  assign n833 = ~n463 & ~n832 ;
  assign n834 = ~n831 & ~n833 ;
  assign n835 = ~n830 & ~n834 ;
  assign n836 = ~\pi129  & ~n835 ;
  assign n837 = ~n231 & ~n691 ;
  assign n838 = ~\pi046  & n240 ;
  assign n839 = n681 & n838 ;
  assign n840 = \pi082  & ~n691 ;
  assign n841 = ~n839 & n840 ;
  assign n842 = ~n837 & ~n841 ;
  assign n843 = ~\pi050  & n842 ;
  assign n844 = \pi066  & ~n231 ;
  assign n845 = ~\pi082  & n844 ;
  assign n846 = n236 & n844 ;
  assign n847 = n839 & n846 ;
  assign n848 = ~n845 & ~n847 ;
  assign n849 = \pi050  & \pi082  ;
  assign n850 = n236 & n849 ;
  assign n851 = ~\pi129  & ~n850 ;
  assign n852 = n848 & n851 ;
  assign n853 = ~n843 & n852 ;
  assign n854 = \pi051  & ~\pi109  ;
  assign n855 = ~\pi106  & ~n699 ;
  assign n856 = ~n854 & n855 ;
  assign n857 = ~\pi129  & ~n856 ;
  assign n858 = \pi052  & ~n699 ;
  assign n859 = ~\pi106  & ~n697 ;
  assign n860 = ~n858 & n859 ;
  assign n861 = ~\pi129  & ~n860 ;
  assign n862 = ~\pi053  & \pi097  ;
  assign n863 = ~n545 & ~n862 ;
  assign n864 = ~\pi058  & ~n545 ;
  assign n865 = ~n604 & n864 ;
  assign n866 = ~n863 & ~n865 ;
  assign n867 = n148 & ~n585 ;
  assign n868 = n521 & n867 ;
  assign n869 = n866 & n868 ;
  assign n870 = n242 & n248 ;
  assign n871 = ~\pi129  & ~n232 ;
  assign n872 = ~n870 & n871 ;
  assign n873 = ~\pi123  & ~\pi129  ;
  assign n874 = \pi114  & ~\pi122  ;
  assign n875 = n873 & n874 ;
  assign n876 = ~\pi026  & \pi037  ;
  assign n877 = ~\pi058  & n876 ;
  assign n878 = ~\pi026  & \pi058  ;
  assign n879 = \pi094  & n878 ;
  assign n880 = ~\pi058  & \pi094  ;
  assign n881 = n526 & n880 ;
  assign n882 = ~n879 & ~n881 ;
  assign n883 = \pi037  & ~\pi116  ;
  assign n884 = ~n878 & ~n883 ;
  assign n885 = ~n585 & ~n884 ;
  assign n886 = n882 & ~n885 ;
  assign n887 = ~\pi053  & ~n886 ;
  assign n888 = ~n877 & ~n887 ;
  assign n889 = n518 & n876 ;
  assign n890 = \pi085  & ~n889 ;
  assign n891 = ~\pi027  & n148 ;
  assign n892 = n148 & n573 ;
  assign n893 = n877 & n892 ;
  assign n894 = ~n891 & ~n893 ;
  assign n895 = ~n890 & ~n894 ;
  assign n896 = ~n888 & n895 ;
  assign n897 = \pi058  & \pi060  ;
  assign n898 = \pi116  & n897 ;
  assign n899 = n584 & n898 ;
  assign n900 = ~\pi027  & n899 ;
  assign n901 = ~\pi085  & ~\pi116  ;
  assign n902 = n583 & n901 ;
  assign n903 = \pi085  & ~n583 ;
  assign n904 = \pi026  & \pi053  ;
  assign n905 = ~\pi058  & ~n904 ;
  assign n906 = ~n903 & n905 ;
  assign n907 = ~n902 & ~n906 ;
  assign n908 = ~\pi027  & \pi057  ;
  assign n909 = ~n907 & n908 ;
  assign n910 = ~n900 & ~n909 ;
  assign n911 = \pi057  & ~\pi058  ;
  assign n912 = n584 & n911 ;
  assign n913 = n910 & ~n912 ;
  assign n914 = n148 & ~n913 ;
  assign n915 = n520 & n585 ;
  assign n916 = n892 & n915 ;
  assign n917 = ~\pi058  & n550 ;
  assign n918 = n494 & n892 ;
  assign n919 = n917 & n918 ;
  assign n920 = ~n916 & ~n919 ;
  assign n921 = \pi059  & ~\pi116  ;
  assign n922 = n510 & n921 ;
  assign n923 = n529 & n922 ;
  assign n924 = n148 & n923 ;
  assign n925 = ~\pi085  & n921 ;
  assign n926 = n595 & n925 ;
  assign n927 = \pi027  & ~n926 ;
  assign n928 = ~n480 & n921 ;
  assign n929 = ~\pi085  & n928 ;
  assign n930 = ~\pi059  & \pi110  ;
  assign n931 = ~\pi059  & ~\pi097  ;
  assign n932 = n501 & n931 ;
  assign n933 = ~n930 & ~n932 ;
  assign n934 = n518 & n933 ;
  assign n935 = n482 & ~n557 ;
  assign n936 = ~\pi085  & ~n935 ;
  assign n937 = n934 & n936 ;
  assign n938 = ~n929 & ~n937 ;
  assign n939 = \pi085  & n518 ;
  assign n940 = n921 & n939 ;
  assign n941 = ~n926 & ~n940 ;
  assign n942 = n938 & n941 ;
  assign n943 = ~n927 & ~n942 ;
  assign n944 = n542 & n943 ;
  assign n945 = ~n924 & ~n944 ;
  assign n946 = ~\pi117  & ~\pi122  ;
  assign n947 = \pi060  & ~n946 ;
  assign n948 = \pi123  & n946 ;
  assign n949 = ~n947 & ~n948 ;
  assign n950 = ~\pi114  & ~\pi122  ;
  assign n951 = \pi123  & ~\pi129  ;
  assign n952 = n950 & n951 ;
  assign n953 = \pi131  & \pi132  ;
  assign n954 = \pi133  & ~\pi138  ;
  assign n955 = n953 & n954 ;
  assign n956 = \pi136  & ~\pi137  ;
  assign n957 = \pi140  & n956 ;
  assign n958 = n955 & n957 ;
  assign n959 = \pi062  & ~\pi129  ;
  assign n960 = ~\pi129  & n956 ;
  assign n961 = n955 & n960 ;
  assign n962 = ~n959 & ~n961 ;
  assign n963 = ~n958 & ~n962 ;
  assign n964 = \pi142  & n956 ;
  assign n965 = n955 & n964 ;
  assign n966 = \pi063  & ~\pi129  ;
  assign n967 = ~n961 & ~n966 ;
  assign n968 = ~n965 & ~n967 ;
  assign n969 = \pi139  & n956 ;
  assign n970 = n955 & n969 ;
  assign n971 = \pi064  & ~\pi129  ;
  assign n972 = ~n961 & ~n971 ;
  assign n973 = ~n970 & ~n972 ;
  assign n974 = \pi146  & n956 ;
  assign n975 = n955 & n974 ;
  assign n976 = \pi065  & ~\pi129  ;
  assign n977 = ~n961 & ~n976 ;
  assign n978 = ~n975 & ~n977 ;
  assign n979 = ~\pi136  & ~\pi137  ;
  assign n980 = \pi143  & n979 ;
  assign n981 = n955 & n980 ;
  assign n982 = \pi066  & ~\pi129  ;
  assign n983 = ~\pi129  & n979 ;
  assign n984 = n955 & n983 ;
  assign n985 = ~n982 & ~n984 ;
  assign n986 = ~n981 & ~n985 ;
  assign n987 = \pi139  & n979 ;
  assign n988 = n955 & n987 ;
  assign n989 = \pi067  & ~\pi129  ;
  assign n990 = ~n984 & ~n989 ;
  assign n991 = ~n988 & ~n990 ;
  assign n992 = \pi141  & n956 ;
  assign n993 = n955 & n992 ;
  assign n994 = \pi068  & ~\pi129  ;
  assign n995 = ~n961 & ~n994 ;
  assign n996 = ~n993 & ~n995 ;
  assign n997 = \pi143  & n956 ;
  assign n998 = n955 & n997 ;
  assign n999 = \pi069  & ~\pi129  ;
  assign n1000 = ~n961 & ~n999 ;
  assign n1001 = ~n998 & ~n1000 ;
  assign n1002 = \pi144  & n956 ;
  assign n1003 = n955 & n1002 ;
  assign n1004 = \pi070  & ~\pi129  ;
  assign n1005 = ~n961 & ~n1004 ;
  assign n1006 = ~n1003 & ~n1005 ;
  assign n1007 = \pi145  & n956 ;
  assign n1008 = n955 & n1007 ;
  assign n1009 = \pi071  & ~\pi129  ;
  assign n1010 = ~n961 & ~n1009 ;
  assign n1011 = ~n1008 & ~n1010 ;
  assign n1012 = \pi140  & n979 ;
  assign n1013 = n955 & n1012 ;
  assign n1014 = \pi072  & ~\pi129  ;
  assign n1015 = ~n984 & ~n1014 ;
  assign n1016 = ~n1013 & ~n1015 ;
  assign n1017 = \pi141  & n979 ;
  assign n1018 = n955 & n1017 ;
  assign n1019 = \pi073  & ~\pi129  ;
  assign n1020 = ~n984 & ~n1019 ;
  assign n1021 = ~n1018 & ~n1020 ;
  assign n1022 = \pi142  & n979 ;
  assign n1023 = n955 & n1022 ;
  assign n1024 = \pi074  & ~\pi129  ;
  assign n1025 = ~n984 & ~n1024 ;
  assign n1026 = ~n1023 & ~n1025 ;
  assign n1027 = \pi144  & n979 ;
  assign n1028 = n955 & n1027 ;
  assign n1029 = \pi075  & ~\pi129  ;
  assign n1030 = ~n984 & ~n1029 ;
  assign n1031 = ~n1028 & ~n1030 ;
  assign n1032 = \pi145  & n979 ;
  assign n1033 = n955 & n1032 ;
  assign n1034 = \pi076  & ~\pi129  ;
  assign n1035 = ~n984 & ~n1034 ;
  assign n1036 = ~n1033 & ~n1035 ;
  assign n1037 = \pi146  & n979 ;
  assign n1038 = n955 & n1037 ;
  assign n1039 = \pi077  & ~\pi129  ;
  assign n1040 = ~n984 & ~n1039 ;
  assign n1041 = ~n1038 & ~n1040 ;
  assign n1042 = ~\pi136  & \pi137  ;
  assign n1043 = ~\pi142  & n1042 ;
  assign n1044 = n955 & n1043 ;
  assign n1045 = \pi078  & ~\pi129  ;
  assign n1046 = ~\pi129  & n1042 ;
  assign n1047 = n955 & n1046 ;
  assign n1048 = ~n1045 & ~n1047 ;
  assign n1049 = ~n1044 & ~n1048 ;
  assign n1050 = ~\pi143  & n1042 ;
  assign n1051 = n955 & n1050 ;
  assign n1052 = \pi079  & ~\pi129  ;
  assign n1053 = ~n1047 & ~n1052 ;
  assign n1054 = ~n1051 & ~n1053 ;
  assign n1055 = ~\pi144  & n1042 ;
  assign n1056 = n955 & n1055 ;
  assign n1057 = \pi080  & ~\pi129  ;
  assign n1058 = ~n1047 & ~n1057 ;
  assign n1059 = ~n1056 & ~n1058 ;
  assign n1060 = ~\pi145  & n1042 ;
  assign n1061 = n955 & n1060 ;
  assign n1062 = \pi081  & ~\pi129  ;
  assign n1063 = ~n1047 & ~n1062 ;
  assign n1064 = ~n1061 & ~n1063 ;
  assign n1065 = ~\pi146  & n1042 ;
  assign n1066 = n955 & n1065 ;
  assign n1067 = \pi082  & ~\pi129  ;
  assign n1068 = ~n1047 & ~n1067 ;
  assign n1069 = ~n1066 & ~n1068 ;
  assign n1070 = \pi136  & ~\pi138  ;
  assign n1071 = \pi031  & n1070 ;
  assign n1072 = \pi137  & n1071 ;
  assign n1073 = ~\pi087  & ~\pi138  ;
  assign n1074 = ~\pi136  & ~n1073 ;
  assign n1075 = \pi115  & \pi138  ;
  assign n1076 = \pi137  & ~n1075 ;
  assign n1077 = n1074 & n1076 ;
  assign n1078 = ~n1072 & ~n1077 ;
  assign n1079 = \pi062  & ~\pi138  ;
  assign n1080 = ~\pi089  & \pi138  ;
  assign n1081 = \pi136  & ~n1080 ;
  assign n1082 = ~n1079 & n1081 ;
  assign n1083 = \pi072  & ~\pi138  ;
  assign n1084 = ~\pi119  & \pi138  ;
  assign n1085 = ~\pi136  & ~n1084 ;
  assign n1086 = ~n1083 & n1085 ;
  assign n1087 = ~n1082 & ~n1086 ;
  assign n1088 = ~\pi137  & ~n1087 ;
  assign n1089 = n1078 & ~n1088 ;
  assign n1090 = ~\pi141  & n1042 ;
  assign n1091 = n955 & n1090 ;
  assign n1092 = \pi084  & ~\pi129  ;
  assign n1093 = ~n1047 & ~n1092 ;
  assign n1094 = ~n1091 & ~n1093 ;
  assign n1095 = ~\pi085  & ~\pi110  ;
  assign n1096 = \pi096  & n1095 ;
  assign n1097 = ~n557 & n1096 ;
  assign n1098 = ~n484 & ~n1097 ;
  assign n1099 = n529 & n542 ;
  assign n1100 = ~n1098 & n1099 ;
  assign n1101 = ~\pi139  & n1042 ;
  assign n1102 = n955 & n1101 ;
  assign n1103 = \pi086  & ~\pi129  ;
  assign n1104 = ~n1047 & ~n1103 ;
  assign n1105 = ~n1102 & ~n1104 ;
  assign n1106 = ~\pi140  & n1042 ;
  assign n1107 = n955 & n1106 ;
  assign n1108 = \pi087  & ~\pi129  ;
  assign n1109 = ~n1047 & ~n1108 ;
  assign n1110 = ~n1107 & ~n1109 ;
  assign n1111 = \pi133  & n953 ;
  assign n1112 = \pi137  & n1070 ;
  assign n1113 = n1111 & n1112 ;
  assign n1114 = ~\pi088  & ~n1113 ;
  assign n1115 = \pi133  & ~\pi139  ;
  assign n1116 = n953 & n1115 ;
  assign n1117 = n1112 & n1116 ;
  assign n1118 = ~\pi129  & ~n1117 ;
  assign n1119 = ~n1114 & n1118 ;
  assign n1120 = ~\pi089  & ~n1113 ;
  assign n1121 = \pi133  & ~\pi140  ;
  assign n1122 = n953 & n1121 ;
  assign n1123 = n1112 & n1122 ;
  assign n1124 = ~\pi129  & ~n1123 ;
  assign n1125 = ~n1120 & n1124 ;
  assign n1126 = ~\pi090  & ~n1113 ;
  assign n1127 = \pi133  & ~\pi142  ;
  assign n1128 = n953 & n1127 ;
  assign n1129 = n1112 & n1128 ;
  assign n1130 = ~\pi129  & ~n1129 ;
  assign n1131 = ~n1126 & n1130 ;
  assign n1132 = ~\pi091  & ~n1113 ;
  assign n1133 = \pi133  & ~\pi143  ;
  assign n1134 = n953 & n1133 ;
  assign n1135 = n1112 & n1134 ;
  assign n1136 = ~\pi129  & ~n1135 ;
  assign n1137 = ~n1132 & n1136 ;
  assign n1138 = ~\pi092  & ~n1113 ;
  assign n1139 = \pi133  & ~\pi144  ;
  assign n1140 = n953 & n1139 ;
  assign n1141 = n1112 & n1140 ;
  assign n1142 = ~\pi129  & ~n1141 ;
  assign n1143 = ~n1138 & n1142 ;
  assign n1144 = ~\pi093  & ~n1113 ;
  assign n1145 = \pi133  & ~\pi146  ;
  assign n1146 = n953 & n1145 ;
  assign n1147 = n1112 & n1146 ;
  assign n1148 = ~\pi129  & ~n1147 ;
  assign n1149 = ~n1144 & n1148 ;
  assign n1150 = \pi082  & \pi138  ;
  assign n1151 = n979 & n1150 ;
  assign n1152 = n1111 & n1151 ;
  assign n1153 = ~\pi094  & ~n1152 ;
  assign n1154 = n1128 & n1151 ;
  assign n1155 = ~\pi129  & ~n1154 ;
  assign n1156 = ~n1153 & n1155 ;
  assign n1157 = \pi133  & \pi143  ;
  assign n1158 = n953 & n1157 ;
  assign n1159 = n1151 & n1158 ;
  assign n1160 = ~\pi129  & n1159 ;
  assign n1161 = ~\pi003  & ~\pi110  ;
  assign n1162 = ~n1111 & ~n1161 ;
  assign n1163 = ~n1152 & ~n1162 ;
  assign n1164 = \pi095  & ~\pi129  ;
  assign n1165 = n1163 & n1164 ;
  assign n1166 = ~n1160 & ~n1165 ;
  assign n1167 = \pi133  & \pi146  ;
  assign n1168 = n953 & n1167 ;
  assign n1169 = n1151 & n1168 ;
  assign n1170 = ~\pi129  & n1169 ;
  assign n1171 = \pi096  & ~\pi129  ;
  assign n1172 = n1163 & n1171 ;
  assign n1173 = ~n1170 & ~n1172 ;
  assign n1174 = \pi133  & \pi145  ;
  assign n1175 = n953 & n1174 ;
  assign n1176 = n1151 & n1175 ;
  assign n1177 = ~\pi129  & n1176 ;
  assign n1178 = \pi097  & ~\pi129  ;
  assign n1179 = n1163 & n1178 ;
  assign n1180 = ~n1177 & ~n1179 ;
  assign n1181 = ~\pi098  & ~n1113 ;
  assign n1182 = \pi133  & ~\pi145  ;
  assign n1183 = n953 & n1182 ;
  assign n1184 = n1112 & n1183 ;
  assign n1185 = ~\pi129  & ~n1184 ;
  assign n1186 = ~n1181 & n1185 ;
  assign n1187 = ~\pi099  & ~n1113 ;
  assign n1188 = \pi133  & ~\pi141  ;
  assign n1189 = n953 & n1188 ;
  assign n1190 = n1112 & n1189 ;
  assign n1191 = ~\pi129  & ~n1190 ;
  assign n1192 = ~n1187 & n1191 ;
  assign n1193 = \pi133  & \pi144  ;
  assign n1194 = n953 & n1193 ;
  assign n1195 = n1151 & n1194 ;
  assign n1196 = ~\pi129  & n1195 ;
  assign n1197 = \pi100  & ~\pi129  ;
  assign n1198 = n1163 & n1197 ;
  assign n1199 = ~n1196 & ~n1198 ;
  assign n1200 = \pi037  & n1070 ;
  assign n1201 = \pi137  & n1200 ;
  assign n1202 = ~\pi082  & ~\pi138  ;
  assign n1203 = ~\pi136  & ~n1202 ;
  assign n1204 = ~\pi096  & \pi138  ;
  assign n1205 = \pi137  & ~n1204 ;
  assign n1206 = n1203 & n1205 ;
  assign n1207 = ~n1201 & ~n1206 ;
  assign n1208 = \pi065  & ~\pi138  ;
  assign n1209 = ~\pi093  & \pi138  ;
  assign n1210 = \pi136  & ~n1209 ;
  assign n1211 = ~n1208 & n1210 ;
  assign n1212 = \pi077  & ~\pi138  ;
  assign n1213 = ~\pi124  & \pi138  ;
  assign n1214 = ~\pi136  & ~n1213 ;
  assign n1215 = ~n1212 & n1214 ;
  assign n1216 = ~n1211 & ~n1215 ;
  assign n1217 = ~\pi137  & ~n1216 ;
  assign n1218 = n1207 & ~n1217 ;
  assign n1219 = \pi091  & n956 ;
  assign n1220 = \pi095  & n1042 ;
  assign n1221 = ~n1219 & ~n1220 ;
  assign n1222 = \pi138  & ~n1221 ;
  assign n1223 = ~\pi034  & \pi136  ;
  assign n1224 = ~\pi079  & ~\pi136  ;
  assign n1225 = \pi137  & ~n1224 ;
  assign n1226 = ~n1223 & n1225 ;
  assign n1227 = \pi069  & \pi136  ;
  assign n1228 = \pi066  & ~\pi136  ;
  assign n1229 = ~\pi137  & ~n1228 ;
  assign n1230 = ~n1227 & n1229 ;
  assign n1231 = ~n1226 & ~n1230 ;
  assign n1232 = ~\pi138  & ~n1231 ;
  assign n1233 = ~n1222 & ~n1232 ;
  assign n1234 = \pi090  & n956 ;
  assign n1235 = \pi094  & n1042 ;
  assign n1236 = ~n1234 & ~n1235 ;
  assign n1237 = \pi138  & ~n1236 ;
  assign n1238 = ~\pi033  & \pi136  ;
  assign n1239 = ~\pi078  & ~\pi136  ;
  assign n1240 = \pi137  & ~n1239 ;
  assign n1241 = ~n1238 & n1240 ;
  assign n1242 = \pi063  & \pi136  ;
  assign n1243 = \pi074  & ~\pi136  ;
  assign n1244 = ~\pi137  & ~n1243 ;
  assign n1245 = ~n1242 & n1244 ;
  assign n1246 = ~n1241 & ~n1245 ;
  assign n1247 = ~\pi138  & ~n1246 ;
  assign n1248 = ~n1237 & ~n1247 ;
  assign n1249 = \pi099  & n956 ;
  assign n1250 = ~\pi112  & n1042 ;
  assign n1251 = ~n1249 & ~n1250 ;
  assign n1252 = \pi138  & ~n1251 ;
  assign n1253 = ~\pi032  & \pi136  ;
  assign n1254 = ~\pi084  & ~\pi136  ;
  assign n1255 = \pi137  & ~n1254 ;
  assign n1256 = ~n1253 & n1255 ;
  assign n1257 = \pi068  & \pi136  ;
  assign n1258 = \pi073  & ~\pi136  ;
  assign n1259 = ~\pi137  & ~n1258 ;
  assign n1260 = ~n1257 & n1259 ;
  assign n1261 = ~n1256 & ~n1260 ;
  assign n1262 = ~\pi138  & ~n1261 ;
  assign n1263 = ~n1252 & ~n1262 ;
  assign n1264 = \pi035  & n1070 ;
  assign n1265 = \pi137  & n1264 ;
  assign n1266 = ~\pi080  & ~\pi138  ;
  assign n1267 = ~\pi136  & ~n1266 ;
  assign n1268 = ~\pi100  & \pi138  ;
  assign n1269 = \pi137  & ~n1268 ;
  assign n1270 = n1267 & n1269 ;
  assign n1271 = ~n1265 & ~n1270 ;
  assign n1272 = \pi070  & ~\pi138  ;
  assign n1273 = ~\pi092  & \pi138  ;
  assign n1274 = \pi136  & ~n1273 ;
  assign n1275 = ~n1272 & n1274 ;
  assign n1276 = \pi075  & ~\pi138  ;
  assign n1277 = ~\pi125  & \pi138  ;
  assign n1278 = ~\pi136  & ~n1277 ;
  assign n1279 = ~n1276 & n1278 ;
  assign n1280 = ~n1275 & ~n1279 ;
  assign n1281 = ~\pi137  & ~n1280 ;
  assign n1282 = n1271 & ~n1281 ;
  assign n1283 = n148 & n534 ;
  assign n1284 = ~n557 & n1095 ;
  assign n1285 = n518 & n520 ;
  assign n1286 = n148 & n1285 ;
  assign n1287 = n1284 & n1286 ;
  assign n1288 = ~n1283 & ~n1287 ;
  assign n1289 = \pi036  & n1070 ;
  assign n1290 = \pi137  & n1289 ;
  assign n1291 = ~\pi081  & ~\pi138  ;
  assign n1292 = ~\pi136  & ~n1291 ;
  assign n1293 = ~\pi097  & \pi138  ;
  assign n1294 = \pi137  & ~n1293 ;
  assign n1295 = n1292 & n1294 ;
  assign n1296 = ~n1290 & ~n1295 ;
  assign n1297 = \pi071  & ~\pi138  ;
  assign n1298 = ~\pi098  & \pi138  ;
  assign n1299 = \pi136  & ~n1298 ;
  assign n1300 = ~n1297 & n1299 ;
  assign n1301 = \pi076  & ~\pi138  ;
  assign n1302 = ~\pi023  & \pi138  ;
  assign n1303 = ~\pi136  & ~n1302 ;
  assign n1304 = ~n1301 & n1303 ;
  assign n1305 = ~n1300 & ~n1304 ;
  assign n1306 = ~\pi137  & ~n1305 ;
  assign n1307 = n1296 & ~n1306 ;
  assign n1308 = \pi030  & n1070 ;
  assign n1309 = \pi137  & n1308 ;
  assign n1310 = ~\pi086  & ~\pi138  ;
  assign n1311 = ~\pi136  & ~n1310 ;
  assign n1312 = ~\pi111  & \pi138  ;
  assign n1313 = \pi137  & ~n1312 ;
  assign n1314 = n1311 & n1313 ;
  assign n1315 = ~n1309 & ~n1314 ;
  assign n1316 = \pi064  & ~\pi138  ;
  assign n1317 = ~\pi088  & \pi138  ;
  assign n1318 = \pi136  & ~n1317 ;
  assign n1319 = ~n1316 & n1318 ;
  assign n1320 = \pi067  & ~\pi138  ;
  assign n1321 = ~\pi120  & \pi138  ;
  assign n1322 = ~\pi136  & ~n1321 ;
  assign n1323 = ~n1320 & n1322 ;
  assign n1324 = ~n1319 & ~n1323 ;
  assign n1325 = ~\pi137  & ~n1324 ;
  assign n1326 = n1315 & ~n1325 ;
  assign n1327 = ~\pi026  & ~\pi039  ;
  assign n1328 = n497 & n1327 ;
  assign n1329 = \pi116  & n148 ;
  assign n1330 = n550 & n1329 ;
  assign n1331 = ~n1328 & n1330 ;
  assign n1332 = ~\pi097  & n478 ;
  assign n1333 = ~n479 & ~n1332 ;
  assign n1334 = n1329 & ~n1333 ;
  assign n1335 = ~\pi139  & n1151 ;
  assign n1336 = ~\pi129  & \pi133  ;
  assign n1337 = n953 & n1336 ;
  assign n1338 = ~\pi111  & ~n1151 ;
  assign n1339 = n1337 & ~n1338 ;
  assign n1340 = ~n1335 & n1339 ;
  assign n1341 = \pi112  & ~n1151 ;
  assign n1342 = ~\pi141  & n1151 ;
  assign n1343 = n1337 & ~n1342 ;
  assign n1344 = ~n1341 & n1343 ;
  assign n1345 = ~\pi011  & n215 ;
  assign n1346 = ~\pi054  & \pi113  ;
  assign n1347 = n148 & ~n1346 ;
  assign n1348 = ~n1345 & n1347 ;
  assign n1349 = \pi115  & ~n1151 ;
  assign n1350 = ~\pi140  & n1151 ;
  assign n1351 = n1337 & ~n1350 ;
  assign n1352 = ~n1349 & n1351 ;
  assign n1353 = ~\pi004  & ~\pi009  ;
  assign n1354 = n204 & n1353 ;
  assign n1355 = \pi054  & n148 ;
  assign n1356 = ~n1354 & n1355 ;
  assign n1357 = \pi122  & ~\pi129  ;
  assign n1358 = \pi054  & ~n363 ;
  assign n1359 = ~\pi054  & ~\pi118  ;
  assign n1360 = ~\pi129  & ~n1359 ;
  assign n1361 = ~n1358 & n1360 ;
  assign n1362 = ~\pi129  & ~n501 ;
  assign n1363 = ~\pi120  & n1161 ;
  assign n1364 = ~\pi111  & ~\pi129  ;
  assign n1365 = ~n1363 & n1364 ;
  assign n1366 = \pi081  & \pi120  ;
  assign n1367 = ~\pi129  & n1366 ;
  assign n1368 = ~\pi129  & ~\pi134  ;
  assign n1369 = ~\pi129  & ~\pi135  ;
  assign n1370 = \pi057  & ~\pi129  ;
  assign n1371 = ~\pi096  & \pi125  ;
  assign n1372 = ~\pi003  & ~n1371 ;
  assign n1373 = ~\pi129  & ~n1372 ;
  assign n1374 = ~\pi126  & \pi132  ;
  assign n1375 = \pi133  & n1374 ;
  assign \po000  = \pi108  ;
  assign \po001  = \pi083  ;
  assign \po002  = \pi104  ;
  assign \po003  = \pi103  ;
  assign \po004  = \pi102  ;
  assign \po005  = \pi105  ;
  assign \po006  = \pi107  ;
  assign \po007  = \pi101  ;
  assign \po008  = \pi126  ;
  assign \po009  = \pi121  ;
  assign \po010  = \pi001  ;
  assign \po011  = \pi000  ;
  assign \po012  = ~1'b0 ;
  assign \po013  = \pi130  ;
  assign \po014  = \pi128  ;
  assign \po015  = ~n194 ;
  assign \po016  = n230 ;
  assign \po017  = n264 ;
  assign \po018  = ~n276 ;
  assign \po019  = n284 ;
  assign \po020  = n300 ;
  assign \po021  = n307 ;
  assign \po022  = n317 ;
  assign \po023  = n323 ;
  assign \po024  = n332 ;
  assign \po025  = ~n342 ;
  assign \po026  = n349 ;
  assign \po027  = ~n355 ;
  assign \po028  = ~n367 ;
  assign \po029  = ~n375 ;
  assign \po030  = n394 ;
  assign \po031  = n400 ;
  assign \po032  = ~n408 ;
  assign \po033  = n417 ;
  assign \po034  = ~n424 ;
  assign \po035  = n438 ;
  assign \po036  = n446 ;
  assign \po037  = ~n454 ;
  assign \po038  = n457 ;
  assign \po039  = n477 ;
  assign \po040  = n525 ;
  assign \po041  = n531 ;
  assign \po042  = n544 ;
  assign \po043  = n590 ;
  assign \po044  = n622 ;
  assign \po045  = n629 ;
  assign \po046  = n636 ;
  assign \po047  = n643 ;
  assign \po048  = n650 ;
  assign \po049  = n657 ;
  assign \po050  = n664 ;
  assign \po051  = n671 ;
  assign \po052  = n678 ;
  assign \po053  = n696 ;
  assign \po054  = n703 ;
  assign \po055  = n722 ;
  assign \po056  = n738 ;
  assign \po057  = n749 ;
  assign \po058  = n762 ;
  assign \po059  = n772 ;
  assign \po060  = n784 ;
  assign \po061  = ~n800 ;
  assign \po062  = n812 ;
  assign \po063  = n825 ;
  assign \po064  = n836 ;
  assign \po065  = n853 ;
  assign \po066  = n857 ;
  assign \po067  = n861 ;
  assign \po068  = n869 ;
  assign \po069  = ~n872 ;
  assign \po070  = n875 ;
  assign \po071  = n896 ;
  assign \po072  = n914 ;
  assign \po073  = ~n920 ;
  assign \po074  = ~n945 ;
  assign \po075  = ~n949 ;
  assign \po076  = n952 ;
  assign \po077  = ~n963 ;
  assign \po078  = ~n968 ;
  assign \po079  = ~n973 ;
  assign \po080  = ~n978 ;
  assign \po081  = ~n986 ;
  assign \po082  = ~n991 ;
  assign \po083  = ~n996 ;
  assign \po084  = ~n1001 ;
  assign \po085  = ~n1006 ;
  assign \po086  = ~n1011 ;
  assign \po087  = ~n1016 ;
  assign \po088  = ~n1021 ;
  assign \po089  = ~n1026 ;
  assign \po090  = ~n1031 ;
  assign \po091  = ~n1036 ;
  assign \po092  = ~n1041 ;
  assign \po093  = n1049 ;
  assign \po094  = n1054 ;
  assign \po095  = n1059 ;
  assign \po096  = n1064 ;
  assign \po097  = n1069 ;
  assign \po098  = ~n1089 ;
  assign \po099  = n1094 ;
  assign \po100  = n1100 ;
  assign \po101  = n1105 ;
  assign \po102  = n1110 ;
  assign \po103  = n1119 ;
  assign \po104  = n1125 ;
  assign \po105  = n1131 ;
  assign \po106  = n1137 ;
  assign \po107  = n1143 ;
  assign \po108  = n1149 ;
  assign \po109  = n1156 ;
  assign \po110  = ~n1166 ;
  assign \po111  = ~n1173 ;
  assign \po112  = ~n1180 ;
  assign \po113  = n1186 ;
  assign \po114  = n1192 ;
  assign \po115  = ~n1199 ;
  assign \po116  = ~n1218 ;
  assign \po117  = ~n1233 ;
  assign \po118  = ~n1248 ;
  assign \po119  = ~n1263 ;
  assign \po120  = ~n1282 ;
  assign \po121  = ~n1288 ;
  assign \po122  = ~n1307 ;
  assign \po123  = ~n1326 ;
  assign \po124  = n1331 ;
  assign \po125  = n1334 ;
  assign \po126  = n1340 ;
  assign \po127  = n1344 ;
  assign \po128  = n1348 ;
  assign \po129  = ~n873 ;
  assign \po130  = n1352 ;
  assign \po131  = n1356 ;
  assign \po132  = ~n1357 ;
  assign \po133  = n1361 ;
  assign \po134  = n1362 ;
  assign \po135  = n1365 ;
  assign \po136  = n1367 ;
  assign \po137  = ~n1368 ;
  assign \po138  = ~n1369 ;
  assign \po139  = n1370 ;
  assign \po140  = n1373 ;
  assign \po141  = n1375 ;
endmodule
