module top (\P1_B_reg/NET0131 , \P1_IR_reg[0]/NET0131 , \P1_IR_reg[10]/NET0131 , \P1_IR_reg[11]/NET0131 , \P1_IR_reg[12]/NET0131 , \P1_IR_reg[13]/NET0131 , \P1_IR_reg[14]/NET0131 , \P1_IR_reg[15]/NET0131 , \P1_IR_reg[16]/NET0131 , \P1_IR_reg[17]/NET0131 , \P1_IR_reg[18]/NET0131 , \P1_IR_reg[19]/NET0131 , \P1_IR_reg[1]/NET0131 , \P1_IR_reg[20]/NET0131 , \P1_IR_reg[21]/NET0131 , \P1_IR_reg[22]/NET0131 , \P1_IR_reg[23]/NET0131 , \P1_IR_reg[24]/NET0131 , \P1_IR_reg[25]/NET0131 , \P1_IR_reg[26]/NET0131 , \P1_IR_reg[27]/NET0131 , \P1_IR_reg[28]/NET0131 , \P1_IR_reg[29]/NET0131 , \P1_IR_reg[2]/NET0131 , \P1_IR_reg[30]/NET0131 , \P1_IR_reg[31]/NET0131 , \P1_IR_reg[3]/NET0131 , \P1_IR_reg[4]/NET0131 , \P1_IR_reg[5]/NET0131 , \P1_IR_reg[6]/NET0131 , \P1_IR_reg[7]/NET0131 , \P1_IR_reg[8]/NET0131 , \P1_IR_reg[9]/NET0131 , \P1_addr_reg[0]/NET0131 , \P1_addr_reg[10]/NET0131 , \P1_addr_reg[11]/NET0131 , \P1_addr_reg[12]/NET0131 , \P1_addr_reg[13]/NET0131 , \P1_addr_reg[14]/NET0131 , \P1_addr_reg[15]/NET0131 , \P1_addr_reg[16]/NET0131 , \P1_addr_reg[17]/NET0131 , \P1_addr_reg[18]/NET0131 , \P1_addr_reg[19]/NET0131 , \P1_addr_reg[1]/NET0131 , \P1_addr_reg[2]/NET0131 , \P1_addr_reg[3]/NET0131 , \P1_addr_reg[4]/NET0131 , \P1_addr_reg[5]/NET0131 , \P1_addr_reg[6]/NET0131 , \P1_addr_reg[7]/NET0131 , \P1_addr_reg[8]/NET0131 , \P1_addr_reg[9]/NET0131 , \P1_d_reg[0]/NET0131 , \P1_d_reg[1]/NET0131 , \P1_datao_reg[0]/NET0131 , \P1_datao_reg[10]/NET0131 , \P1_datao_reg[11]/NET0131 , \P1_datao_reg[12]/NET0131 , \P1_datao_reg[13]/NET0131 , \P1_datao_reg[14]/NET0131 , \P1_datao_reg[15]/NET0131 , \P1_datao_reg[16]/NET0131 , \P1_datao_reg[17]/NET0131 , \P1_datao_reg[18]/NET0131 , \P1_datao_reg[19]/NET0131 , \P1_datao_reg[1]/NET0131 , \P1_datao_reg[20]/NET0131 , \P1_datao_reg[21]/NET0131 , \P1_datao_reg[22]/NET0131 , \P1_datao_reg[23]/NET0131 , \P1_datao_reg[24]/NET0131 , \P1_datao_reg[25]/NET0131 , \P1_datao_reg[26]/NET0131 , \P1_datao_reg[27]/NET0131 , \P1_datao_reg[28]/NET0131 , \P1_datao_reg[29]/NET0131 , \P1_datao_reg[2]/NET0131 , \P1_datao_reg[30]/NET0131 , \P1_datao_reg[31]/NET0131 , \P1_datao_reg[3]/NET0131 , \P1_datao_reg[4]/NET0131 , \P1_datao_reg[5]/NET0131 , \P1_datao_reg[6]/NET0131 , \P1_datao_reg[7]/NET0131 , \P1_datao_reg[8]/NET0131 , \P1_datao_reg[9]/NET0131 , \P1_rd_reg/NET0131 , \P1_reg0_reg[0]/NET0131 , \P1_reg0_reg[10]/NET0131 , \P1_reg0_reg[11]/NET0131 , \P1_reg0_reg[12]/NET0131 , \P1_reg0_reg[13]/NET0131 , \P1_reg0_reg[14]/NET0131 , \P1_reg0_reg[15]/NET0131 , \P1_reg0_reg[16]/NET0131 , \P1_reg0_reg[17]/NET0131 , \P1_reg0_reg[18]/NET0131 , \P1_reg0_reg[19]/NET0131 , \P1_reg0_reg[1]/NET0131 , \P1_reg0_reg[20]/NET0131 , \P1_reg0_reg[21]/NET0131 , \P1_reg0_reg[22]/NET0131 , \P1_reg0_reg[23]/NET0131 , \P1_reg0_reg[24]/NET0131 , \P1_reg0_reg[25]/NET0131 , \P1_reg0_reg[26]/NET0131 , \P1_reg0_reg[27]/NET0131 , \P1_reg0_reg[28]/NET0131 , \P1_reg0_reg[29]/NET0131 , \P1_reg0_reg[2]/NET0131 , \P1_reg0_reg[30]/NET0131 , \P1_reg0_reg[31]/NET0131 , \P1_reg0_reg[3]/NET0131 , \P1_reg0_reg[4]/NET0131 , \P1_reg0_reg[5]/NET0131 , \P1_reg0_reg[6]/NET0131 , \P1_reg0_reg[7]/NET0131 , \P1_reg0_reg[8]/NET0131 , \P1_reg0_reg[9]/NET0131 , \P1_reg1_reg[0]/NET0131 , \P1_reg1_reg[10]/NET0131 , \P1_reg1_reg[11]/NET0131 , \P1_reg1_reg[12]/NET0131 , \P1_reg1_reg[13]/NET0131 , \P1_reg1_reg[14]/NET0131 , \P1_reg1_reg[15]/NET0131 , \P1_reg1_reg[16]/NET0131 , \P1_reg1_reg[17]/NET0131 , \P1_reg1_reg[18]/NET0131 , \P1_reg1_reg[19]/NET0131 , \P1_reg1_reg[1]/NET0131 , \P1_reg1_reg[20]/NET0131 , \P1_reg1_reg[21]/NET0131 , \P1_reg1_reg[22]/NET0131 , \P1_reg1_reg[23]/NET0131 , \P1_reg1_reg[24]/NET0131 , \P1_reg1_reg[25]/NET0131 , \P1_reg1_reg[26]/NET0131 , \P1_reg1_reg[27]/NET0131 , \P1_reg1_reg[28]/NET0131 , \P1_reg1_reg[29]/NET0131 , \P1_reg1_reg[2]/NET0131 , \P1_reg1_reg[30]/NET0131 , \P1_reg1_reg[31]/NET0131 , \P1_reg1_reg[3]/NET0131 , \P1_reg1_reg[4]/NET0131 , \P1_reg1_reg[5]/NET0131 , \P1_reg1_reg[6]/NET0131 , \P1_reg1_reg[7]/NET0131 , \P1_reg1_reg[8]/NET0131 , \P1_reg1_reg[9]/NET0131 , \P1_reg2_reg[0]/NET0131 , \P1_reg2_reg[10]/NET0131 , \P1_reg2_reg[11]/NET0131 , \P1_reg2_reg[12]/NET0131 , \P1_reg2_reg[13]/NET0131 , \P1_reg2_reg[14]/NET0131 , \P1_reg2_reg[15]/NET0131 , \P1_reg2_reg[16]/NET0131 , \P1_reg2_reg[17]/NET0131 , \P1_reg2_reg[18]/NET0131 , \P1_reg2_reg[19]/NET0131 , \P1_reg2_reg[1]/NET0131 , \P1_reg2_reg[20]/NET0131 , \P1_reg2_reg[21]/NET0131 , \P1_reg2_reg[22]/NET0131 , \P1_reg2_reg[23]/NET0131 , \P1_reg2_reg[24]/NET0131 , \P1_reg2_reg[25]/NET0131 , \P1_reg2_reg[26]/NET0131 , \P1_reg2_reg[27]/NET0131 , \P1_reg2_reg[28]/NET0131 , \P1_reg2_reg[29]/NET0131 , \P1_reg2_reg[2]/NET0131 , \P1_reg2_reg[30]/NET0131 , \P1_reg2_reg[31]/NET0131 , \P1_reg2_reg[3]/NET0131 , \P1_reg2_reg[4]/NET0131 , \P1_reg2_reg[5]/NET0131 , \P1_reg2_reg[6]/NET0131 , \P1_reg2_reg[7]/NET0131 , \P1_reg2_reg[8]/NET0131 , \P1_reg2_reg[9]/NET0131 , \P1_reg3_reg[0]/NET0131 , \P1_reg3_reg[10]/NET0131 , \P1_reg3_reg[11]/NET0131 , \P1_reg3_reg[12]/NET0131 , \P1_reg3_reg[13]/NET0131 , \P1_reg3_reg[14]/NET0131 , \P1_reg3_reg[15]/NET0131 , \P1_reg3_reg[16]/NET0131 , \P1_reg3_reg[17]/NET0131 , \P1_reg3_reg[18]/NET0131 , \P1_reg3_reg[19]/NET0131 , \P1_reg3_reg[1]/NET0131 , \P1_reg3_reg[20]/NET0131 , \P1_reg3_reg[21]/NET0131 , \P1_reg3_reg[22]/NET0131 , \P1_reg3_reg[23]/NET0131 , \P1_reg3_reg[24]/NET0131 , \P1_reg3_reg[25]/NET0131 , \P1_reg3_reg[26]/NET0131 , \P1_reg3_reg[27]/NET0131 , \P1_reg3_reg[28]/NET0131 , \P1_reg3_reg[2]/NET0131 , \P1_reg3_reg[3]/NET0131 , \P1_reg3_reg[4]/NET0131 , \P1_reg3_reg[5]/NET0131 , \P1_reg3_reg[6]/NET0131 , \P1_reg3_reg[7]/NET0131 , \P1_reg3_reg[8]/NET0131 , \P1_reg3_reg[9]/NET0131 , \P1_state_reg[0]/NET0131 , \P1_wr_reg/NET0131 , \P2_B_reg/NET0131 , \P2_IR_reg[0]/NET0131 , \P2_IR_reg[10]/NET0131 , \P2_IR_reg[11]/NET0131 , \P2_IR_reg[12]/NET0131 , \P2_IR_reg[13]/NET0131 , \P2_IR_reg[14]/NET0131 , \P2_IR_reg[15]/NET0131 , \P2_IR_reg[16]/NET0131 , \P2_IR_reg[17]/NET0131 , \P2_IR_reg[18]/NET0131 , \P2_IR_reg[19]/NET0131 , \P2_IR_reg[1]/NET0131 , \P2_IR_reg[20]/NET0131 , \P2_IR_reg[21]/NET0131 , \P2_IR_reg[22]/NET0131 , \P2_IR_reg[23]/NET0131 , \P2_IR_reg[24]/NET0131 , \P2_IR_reg[25]/NET0131 , \P2_IR_reg[26]/NET0131 , \P2_IR_reg[27]/NET0131 , \P2_IR_reg[28]/NET0131 , \P2_IR_reg[29]/NET0131 , \P2_IR_reg[2]/NET0131 , \P2_IR_reg[30]/NET0131 , \P2_IR_reg[31]/NET0131 , \P2_IR_reg[3]/NET0131 , \P2_IR_reg[4]/NET0131 , \P2_IR_reg[5]/NET0131 , \P2_IR_reg[6]/NET0131 , \P2_IR_reg[7]/NET0131 , \P2_IR_reg[8]/NET0131 , \P2_IR_reg[9]/NET0131 , \P2_addr_reg[0]/NET0131 , \P2_addr_reg[10]/NET0131 , \P2_addr_reg[11]/NET0131 , \P2_addr_reg[12]/NET0131 , \P2_addr_reg[13]/NET0131 , \P2_addr_reg[14]/NET0131 , \P2_addr_reg[15]/NET0131 , \P2_addr_reg[16]/NET0131 , \P2_addr_reg[17]/NET0131 , \P2_addr_reg[18]/NET0131 , \P2_addr_reg[19]/NET0131 , \P2_addr_reg[1]/NET0131 , \P2_addr_reg[2]/NET0131 , \P2_addr_reg[3]/NET0131 , \P2_addr_reg[4]/NET0131 , \P2_addr_reg[5]/NET0131 , \P2_addr_reg[6]/NET0131 , \P2_addr_reg[7]/NET0131 , \P2_addr_reg[8]/NET0131 , \P2_addr_reg[9]/NET0131 , \P2_d_reg[0]/NET0131 , \P2_d_reg[1]/NET0131 , \P2_datao_reg[0]/NET0131 , \P2_datao_reg[10]/NET0131 , \P2_datao_reg[11]/NET0131 , \P2_datao_reg[12]/NET0131 , \P2_datao_reg[13]/NET0131 , \P2_datao_reg[14]/NET0131 , \P2_datao_reg[15]/NET0131 , \P2_datao_reg[16]/NET0131 , \P2_datao_reg[17]/NET0131 , \P2_datao_reg[18]/NET0131 , \P2_datao_reg[19]/NET0131 , \P2_datao_reg[1]/NET0131 , \P2_datao_reg[20]/NET0131 , \P2_datao_reg[21]/NET0131 , \P2_datao_reg[22]/NET0131 , \P2_datao_reg[23]/NET0131 , \P2_datao_reg[24]/NET0131 , \P2_datao_reg[25]/NET0131 , \P2_datao_reg[26]/NET0131 , \P2_datao_reg[27]/NET0131 , \P2_datao_reg[28]/NET0131 , \P2_datao_reg[29]/NET0131 , \P2_datao_reg[2]/NET0131 , \P2_datao_reg[30]/NET0131 , \P2_datao_reg[31]/NET0131 , \P2_datao_reg[3]/NET0131 , \P2_datao_reg[4]/NET0131 , \P2_datao_reg[5]/NET0131 , \P2_datao_reg[6]/NET0131 , \P2_datao_reg[7]/NET0131 , \P2_datao_reg[8]/NET0131 , \P2_datao_reg[9]/NET0131 , \P2_rd_reg/NET0131 , \P2_reg0_reg[0]/NET0131 , \P2_reg0_reg[10]/NET0131 , \P2_reg0_reg[11]/NET0131 , \P2_reg0_reg[12]/NET0131 , \P2_reg0_reg[13]/NET0131 , \P2_reg0_reg[14]/NET0131 , \P2_reg0_reg[15]/NET0131 , \P2_reg0_reg[16]/NET0131 , \P2_reg0_reg[17]/NET0131 , \P2_reg0_reg[18]/NET0131 , \P2_reg0_reg[19]/NET0131 , \P2_reg0_reg[1]/NET0131 , \P2_reg0_reg[20]/NET0131 , \P2_reg0_reg[21]/NET0131 , \P2_reg0_reg[22]/NET0131 , \P2_reg0_reg[23]/NET0131 , \P2_reg0_reg[24]/NET0131 , \P2_reg0_reg[25]/NET0131 , \P2_reg0_reg[26]/NET0131 , \P2_reg0_reg[27]/NET0131 , \P2_reg0_reg[28]/NET0131 , \P2_reg0_reg[29]/NET0131 , \P2_reg0_reg[2]/NET0131 , \P2_reg0_reg[30]/NET0131 , \P2_reg0_reg[31]/NET0131 , \P2_reg0_reg[3]/NET0131 , \P2_reg0_reg[4]/NET0131 , \P2_reg0_reg[5]/NET0131 , \P2_reg0_reg[6]/NET0131 , \P2_reg0_reg[7]/NET0131 , \P2_reg0_reg[8]/NET0131 , \P2_reg0_reg[9]/NET0131 , \P2_reg1_reg[0]/NET0131 , \P2_reg1_reg[10]/NET0131 , \P2_reg1_reg[11]/NET0131 , \P2_reg1_reg[12]/NET0131 , \P2_reg1_reg[13]/NET0131 , \P2_reg1_reg[14]/NET0131 , \P2_reg1_reg[15]/NET0131 , \P2_reg1_reg[16]/NET0131 , \P2_reg1_reg[17]/NET0131 , \P2_reg1_reg[18]/NET0131 , \P2_reg1_reg[19]/NET0131 , \P2_reg1_reg[1]/NET0131 , \P2_reg1_reg[20]/NET0131 , \P2_reg1_reg[21]/NET0131 , \P2_reg1_reg[22]/NET0131 , \P2_reg1_reg[23]/NET0131 , \P2_reg1_reg[24]/NET0131 , \P2_reg1_reg[25]/NET0131 , \P2_reg1_reg[26]/NET0131 , \P2_reg1_reg[27]/NET0131 , \P2_reg1_reg[28]/NET0131 , \P2_reg1_reg[29]/NET0131 , \P2_reg1_reg[2]/NET0131 , \P2_reg1_reg[30]/NET0131 , \P2_reg1_reg[31]/NET0131 , \P2_reg1_reg[3]/NET0131 , \P2_reg1_reg[4]/NET0131 , \P2_reg1_reg[5]/NET0131 , \P2_reg1_reg[6]/NET0131 , \P2_reg1_reg[7]/NET0131 , \P2_reg1_reg[8]/NET0131 , \P2_reg1_reg[9]/NET0131 , \P2_reg2_reg[0]/NET0131 , \P2_reg2_reg[10]/NET0131 , \P2_reg2_reg[11]/NET0131 , \P2_reg2_reg[12]/NET0131 , \P2_reg2_reg[13]/NET0131 , \P2_reg2_reg[14]/NET0131 , \P2_reg2_reg[15]/NET0131 , \P2_reg2_reg[16]/NET0131 , \P2_reg2_reg[17]/NET0131 , \P2_reg2_reg[18]/NET0131 , \P2_reg2_reg[19]/NET0131 , \P2_reg2_reg[1]/NET0131 , \P2_reg2_reg[20]/NET0131 , \P2_reg2_reg[21]/NET0131 , \P2_reg2_reg[22]/NET0131 , \P2_reg2_reg[23]/NET0131 , \P2_reg2_reg[24]/NET0131 , \P2_reg2_reg[25]/NET0131 , \P2_reg2_reg[26]/NET0131 , \P2_reg2_reg[27]/NET0131 , \P2_reg2_reg[28]/NET0131 , \P2_reg2_reg[29]/NET0131 , \P2_reg2_reg[2]/NET0131 , \P2_reg2_reg[30]/NET0131 , \P2_reg2_reg[31]/NET0131 , \P2_reg2_reg[3]/NET0131 , \P2_reg2_reg[4]/NET0131 , \P2_reg2_reg[5]/NET0131 , \P2_reg2_reg[6]/NET0131 , \P2_reg2_reg[7]/NET0131 , \P2_reg2_reg[8]/NET0131 , \P2_reg2_reg[9]/NET0131 , \P2_reg3_reg[0]/NET0131 , \P2_reg3_reg[10]/NET0131 , \P2_reg3_reg[11]/NET0131 , \P2_reg3_reg[12]/NET0131 , \P2_reg3_reg[13]/NET0131 , \P2_reg3_reg[14]/NET0131 , \P2_reg3_reg[15]/NET0131 , \P2_reg3_reg[16]/NET0131 , \P2_reg3_reg[17]/NET0131 , \P2_reg3_reg[18]/NET0131 , \P2_reg3_reg[19]/NET0131 , \P2_reg3_reg[1]/NET0131 , \P2_reg3_reg[20]/NET0131 , \P2_reg3_reg[21]/NET0131 , \P2_reg3_reg[22]/NET0131 , \P2_reg3_reg[23]/NET0131 , \P2_reg3_reg[24]/NET0131 , \P2_reg3_reg[25]/NET0131 , \P2_reg3_reg[26]/NET0131 , \P2_reg3_reg[27]/NET0131 , \P2_reg3_reg[28]/NET0131 , \P2_reg3_reg[2]/NET0131 , \P2_reg3_reg[3]/NET0131 , \P2_reg3_reg[4]/NET0131 , \P2_reg3_reg[5]/NET0131 , \P2_reg3_reg[6]/NET0131 , \P2_reg3_reg[7]/NET0131 , \P2_reg3_reg[8]/NET0131 , \P2_reg3_reg[9]/NET0131 , \P2_wr_reg/NET0131 , \si[0]_pad , \si[10]_pad , \si[11]_pad , \si[12]_pad , \si[13]_pad , \si[14]_pad , \si[15]_pad , \si[16]_pad , \si[17]_pad , \si[18]_pad , \si[19]_pad , \si[1]_pad , \si[20]_pad , \si[21]_pad , \si[22]_pad , \si[23]_pad , \si[24]_pad , \si[25]_pad , \si[26]_pad , \si[27]_pad , \si[28]_pad , \si[29]_pad , \si[2]_pad , \si[30]_pad , \si[31]_pad , \si[3]_pad , \si[4]_pad , \si[5]_pad , \si[6]_pad , \si[7]_pad , \si[8]_pad , \si[9]_pad , \P1_state_reg[0]/NET0131_syn_2 , \_al_n0 , \_al_n1 , \g35/_0_ , \g73637/_0_ , \g73647/_0_ , \g73648/_0_ , \g73649/_0_ , \g73650/_0_ , \g73667/_0_ , \g73668/_0_ , \g73669/_0_ , \g73670/_0_ , \g73671/_0_ , \g73672/_0_ , \g73674/_0_ , \g73675/_0_ , \g73709/_0_ , \g73710/_0_ , \g73711/_0_ , \g73716/_0_ , \g73717/_0_ , \g73718/_0_ , \g73719/_0_ , \g73720/_0_ , \g73721/_0_ , \g73722/_0_ , \g73723/_0_ , \g73724/_0_ , \g73765/_0_ , \g73769/_0_ , \g73770/_0_ , \g73771/_0_ , \g73772/_0_ , \g73773/_0_ , \g73774/_0_ , \g73775/_0_ , \g73776/_0_ , \g73777/_0_ , \g73778/_0_ , \g73779/_0_ , \g73780/_0_ , \g73781/_0_ , \g73782/_0_ , \g73783/_0_ , \g73784/_0_ , \g73785/_0_ , \g73786/_0_ , \g73787/_0_ , \g73788/_0_ , \g73789/_0_ , \g73790/_0_ , \g73791/_0_ , \g73792/_0_ , \g73845/_0_ , \g73846/_0_ , \g73847/_0_ , \g73848/_0_ , \g73860/_0_ , \g73863/_0_ , \g73864/_0_ , \g73867/_0_ , \g73870/_0_ , \g73871/_0_ , \g73872/_0_ , \g73873/_0_ , \g73874/_0_ , \g73875/_0_ , \g73876/_0_ , \g73877/_0_ , \g73878/_0_ , \g73879/_0_ , \g73880/_0_ , \g73924/_0_ , \g73925/_0_ , \g73949/_0_ , \g73950/_0_ , \g73953/_0_ , \g73954/_0_ , \g73955/_0_ , \g73956/_0_ , \g73957/_0_ , \g73958/_0_ , \g73960/_0_ , \g73961/_0_ , \g73962/_0_ , \g73963/_0_ , \g73964/_0_ , \g73965/_0_ , \g73966/_0_ , \g73967/_0_ , \g73968/_0_ , \g73969/_0_ , \g73970/_0_ , \g73971/_0_ , \g73972/_0_ , \g73973/_0_ , \g73974/_0_ , \g73975/_0_ , \g73976/_0_ , \g73977/_0_ , \g73978/_0_ , \g73979/_0_ , \g73980/_0_ , \g74062/_0_ , \g74063/_0_ , \g74064/_0_ , \g74065/_0_ , \g74066/_0_ , \g74071/_0_ , \g74072/_0_ , \g74105/_0_ , \g74106/_0_ , \g74107/_0_ , \g74108/_0_ , \g74109/_0_ , \g74110/_0_ , \g74111/_0_ , \g74112/_0_ , \g74113/_0_ , \g74114/_0_ , \g74115/_0_ , \g74167/_0_ , \g74168/_0_ , \g74169/_0_ , \g74170/_0_ , \g74172/_0_ , \g74173/_0_ , \g74174/_0_ , \g74175/_0_ , \g74225/_0_ , \g74226/_0_ , \g74227/_0_ , \g74229/_0_ , \g74230/_0_ , \g74231/_0_ , \g74232/_0_ , \g74233/_0_ , \g74234/_0_ , \g74235/_0_ , \g74236/_0_ , \g74237/_0_ , \g74238/_0_ , \g74239/_0_ , \g74240/_0_ , \g74241/_0_ , \g74242/_0_ , \g74243/_0_ , \g74244/_0_ , \g74245/_0_ , \g74246/_0_ , \g74247/_0_ , \g74248/_0_ , \g74249/_0_ , \g74250/_0_ , \g74251/_0_ , \g74252/_0_ , \g74253/_0_ , \g74254/_0_ , \g74255/_0_ , \g74330/_0_ , \g74331/_0_ , \g74333/_0_ , \g74334/_0_ , \g74335/_0_ , \g74390/_0_ , \g74391/_0_ , \g74405/_0_ , \g74407/_0_ , \g74408/_0_ , \g74409/_0_ , \g74410/_0_ , \g74411/_0_ , \g74412/_0_ , \g74413/_0_ , \g74414/_0_ , \g74415/_0_ , \g74416/_0_ , \g74417/_0_ , \g74418/_0_ , \g74419/_0_ , \g74420/_0_ , \g74421/_0_ , \g74422/_0_ , \g74483/_0_ , \g74485/_0_ , \g74486/_0_ , \g74487/_0_ , \g74576/_0_ , \g74578/_0_ , \g74581/_0_ , \g74582/_0_ , \g74583/_0_ , \g74584/_0_ , \g74585/_0_ , \g74588/_0_ , \g74589/_0_ , \g74590/_0_ , \g74591/_0_ , \g74592/_0_ , \g74595/_0_ , \g74596/_0_ , \g74597/_0_ , \g74598/_0_ , \g74599/_0_ , \g74600/_0_ , \g74601/_0_ , \g74602/_0_ , \g74711/_0_ , \g74835/_0_ , \g74836/_0_ , \g74838/_0_ , \g74840/_0_ , \g74841/_0_ , \g74843/_0_ , \g74844/_0_ , \g74963/_0_ , \g75075/_0_ , \g75078/_0_ , \g75079/_0_ , \g75083/_0_ , \g75084/_0_ , \g75089/_0_ , \g75090/_0_ , \g75091/_0_ , \g75224/_0_ , \g75233/_0_ , \g75234/_0_ , \g75427/_0_ , \g75430/_0_ , \g75434/_0_ , \g75436/_0_ , \g75438/_0_ , \g75844/_0_ , \g75850/_0_ , \g75851/_0_ , \g75860/_0_ , \g75865/_0_ , \g75867/_0_ , \g76076/_0_ , \g76375/_0_ , \g76896/_0_ , \g76901/_0_ , \g76905/_0_ , \g77085/_0_ , \g77892/_0_ , \g77897/_0_ , \g77902/_0_ , \g78635/_0_ , \g78636/_0_ , \g78640/_0_ , \g78642/_0_ , \g78645/_0_ , \g78964/_0_ , \g83163/_3_ , \g83164/_3_ , \g83165/_3_ , \g83166/_3_ , \g83167/_3_ , \g83168/_3_ , \g83644/_0_ , \g83645/_0_ , \g83646/_0_ , \g83647/_0_ , \g83648/_0_ , \g83649/_0_ , \g83650/_0_ , \g83651/_0_ , \g83652/_0_ , \g83653/_0_ , \g83654/_0_ , \g83655/_0_ , \g83656/_0_ , \g83657/_0_ , \g83658/_0_ , \g83659/_0_ , \g83660/_0_ , \g83661/_0_ , \g83662/_0_ , \g83663/_0_ , \g83664/_0_ , \g83665/_0_ , \g83666/_0_ , \g83667/_3_ , \g83668/_0_ , \g83669/_0_ , \g83670/_0_ , \g83671/_0_ , \g83715/_3_ , \g83716/_3_ , \g83717/_3_ , \g83718/_3_ , \g83719/_3_ , \g83720/_3_ , \g83721/_3_ , \g83722/_3_ , \g83723/_3_ , \g83724/_3_ , \g83725/_0_ , \g83726/_3_ , \g83727/_3_ , \g83728/_3_ , \g83729/_3_ , \g83730/_3_ , \g83731/_3_ , \g83732/_3_ , \g83733/_3_ , \g83734/_3_ , \g83735/_0_ , \g83736/_0_ , \g83737/_0_ , \g83738/_3_ , \g83739/_3_ , \g83740/_0_ , \g83741/_3_ , \g83742/_3_ , \g84164/_0_ , \g84181/_0_ , \g85146/_0_ , \g85147/_0_ , \g85148/_0_ , \g85149/_0_ , \g85151/_0_ , \g85152/_0_ , \g85154/_0_ , \g85155/_0_ , \g85156/_0_ , \g85157/_0_ , \g85158/_0_ , \g85159/_0_ , \g85160/_0_ , \g85161/_0_ , \g85162/_0_ , \g85163/_0_ , \g85164/_0_ , \g85165/_0_ , \g85166/_0_ , \g85167/_0_ , \g85168/_0_ , \g85169/_0_ , \g85171/_0_ , \g85173/_0_ , \g85174/_0_ , \g85175/_0_ , \g85176/_0_ , \g85178/_0_ , \g85179/_0_ , \g85180/_0_ , \g85181/_0_ , \g85182/_0_ , \g85183/_0_ , \g85184/_0_ , \g85185/_0_ , \g85186/_0_ , \g85187/_0_ , \g85188/_0_ , \g85189/_0_ , \g85190/_0_ , \g85510/_0_ , \g85711/u3_syn_4 , \g85972/_0_ , \g86107/_0_ , \g86200/u3_syn_4 , \g86477/_0_ , \g86548/_0_ , \g86652/u3_syn_4 , \g86807/u3_syn_4 , \g87581/_0_ , \g88104/_0_ , \g88112/_0_ , \g88136/_0_ , \g88148/_0_ , \g88157/_0_ , \g88171/_0_ , \g88179/_0_ , \g88208/_0_ , \g88217/_0_ , \g88222/_0_ , \g88228/_0_ , \g88236/_0_ , \g88242/_0_ , \g88252_dup/_0_ , \g88253/_2_ , \g88259/_0_ , \g88274/_0_ , \g88286/_0_ , \g88296/_0_ , \g88306/_0_ , \g88319/_0_ , \g88330/_0_ , \g88370/_0_ , \g88375/_0_ , \g88388/_0_ , \g88397/_0_ , \g88404/_0_ , \g88793/_0_ , \g88834/_0_ , \g88905/_0_ , \g88910/_0_ , \g88936_dup/_0_ , \g88953/_0_ , \g88962/_0_ , \g89007/_0_ , \g89018/_0_ , \g89024/_0_ , \g89031/_0_ , \g89066/_0_ , \g89082/_0_ , \g89097/_0_ , \g90677/_1__syn_2 , \g96226/_0_ , \g96236/_0_ , \g96261/_0_ , \g96339/_0_ , \g96380/_1_ , \g96418/_0_ , \g96566/_1_ , \g96574/_0_ , \g96620/_0_ , \g96629/_0_ , \g96735/_0_ , \g96866/_0_ , \g96875/_0_ , \g96910/_0_ , \g96946/_0_ , \g96965/_0_ , \g97098/_0_ , \g97228/_0_ , \g97231/_0_ , \g97242/_0_ , \g97384/_0_ , \g97409/_0_ , \g97506/_0_ , \g97626/_0_ , rd_pad, \so[0]_pad , \so[10]_pad , \so[11]_pad , \so[12]_pad , \so[13]_pad , \so[14]_pad , \so[15]_pad , \so[16]_pad , \so[17]_pad , \so[18]_pad , \so[19]_pad , \so[1]_pad , \so[2]_pad , \so[3]_pad , \so[4]_pad , \so[5]_pad , \so[6]_pad , \so[7]_pad , \so[8]_pad , \so[9]_pad , wr_pad);
	input \P1_B_reg/NET0131  ;
	input \P1_IR_reg[0]/NET0131  ;
	input \P1_IR_reg[10]/NET0131  ;
	input \P1_IR_reg[11]/NET0131  ;
	input \P1_IR_reg[12]/NET0131  ;
	input \P1_IR_reg[13]/NET0131  ;
	input \P1_IR_reg[14]/NET0131  ;
	input \P1_IR_reg[15]/NET0131  ;
	input \P1_IR_reg[16]/NET0131  ;
	input \P1_IR_reg[17]/NET0131  ;
	input \P1_IR_reg[18]/NET0131  ;
	input \P1_IR_reg[19]/NET0131  ;
	input \P1_IR_reg[1]/NET0131  ;
	input \P1_IR_reg[20]/NET0131  ;
	input \P1_IR_reg[21]/NET0131  ;
	input \P1_IR_reg[22]/NET0131  ;
	input \P1_IR_reg[23]/NET0131  ;
	input \P1_IR_reg[24]/NET0131  ;
	input \P1_IR_reg[25]/NET0131  ;
	input \P1_IR_reg[26]/NET0131  ;
	input \P1_IR_reg[27]/NET0131  ;
	input \P1_IR_reg[28]/NET0131  ;
	input \P1_IR_reg[29]/NET0131  ;
	input \P1_IR_reg[2]/NET0131  ;
	input \P1_IR_reg[30]/NET0131  ;
	input \P1_IR_reg[31]/NET0131  ;
	input \P1_IR_reg[3]/NET0131  ;
	input \P1_IR_reg[4]/NET0131  ;
	input \P1_IR_reg[5]/NET0131  ;
	input \P1_IR_reg[6]/NET0131  ;
	input \P1_IR_reg[7]/NET0131  ;
	input \P1_IR_reg[8]/NET0131  ;
	input \P1_IR_reg[9]/NET0131  ;
	input \P1_addr_reg[0]/NET0131  ;
	input \P1_addr_reg[10]/NET0131  ;
	input \P1_addr_reg[11]/NET0131  ;
	input \P1_addr_reg[12]/NET0131  ;
	input \P1_addr_reg[13]/NET0131  ;
	input \P1_addr_reg[14]/NET0131  ;
	input \P1_addr_reg[15]/NET0131  ;
	input \P1_addr_reg[16]/NET0131  ;
	input \P1_addr_reg[17]/NET0131  ;
	input \P1_addr_reg[18]/NET0131  ;
	input \P1_addr_reg[19]/NET0131  ;
	input \P1_addr_reg[1]/NET0131  ;
	input \P1_addr_reg[2]/NET0131  ;
	input \P1_addr_reg[3]/NET0131  ;
	input \P1_addr_reg[4]/NET0131  ;
	input \P1_addr_reg[5]/NET0131  ;
	input \P1_addr_reg[6]/NET0131  ;
	input \P1_addr_reg[7]/NET0131  ;
	input \P1_addr_reg[8]/NET0131  ;
	input \P1_addr_reg[9]/NET0131  ;
	input \P1_d_reg[0]/NET0131  ;
	input \P1_d_reg[1]/NET0131  ;
	input \P1_datao_reg[0]/NET0131  ;
	input \P1_datao_reg[10]/NET0131  ;
	input \P1_datao_reg[11]/NET0131  ;
	input \P1_datao_reg[12]/NET0131  ;
	input \P1_datao_reg[13]/NET0131  ;
	input \P1_datao_reg[14]/NET0131  ;
	input \P1_datao_reg[15]/NET0131  ;
	input \P1_datao_reg[16]/NET0131  ;
	input \P1_datao_reg[17]/NET0131  ;
	input \P1_datao_reg[18]/NET0131  ;
	input \P1_datao_reg[19]/NET0131  ;
	input \P1_datao_reg[1]/NET0131  ;
	input \P1_datao_reg[20]/NET0131  ;
	input \P1_datao_reg[21]/NET0131  ;
	input \P1_datao_reg[22]/NET0131  ;
	input \P1_datao_reg[23]/NET0131  ;
	input \P1_datao_reg[24]/NET0131  ;
	input \P1_datao_reg[25]/NET0131  ;
	input \P1_datao_reg[26]/NET0131  ;
	input \P1_datao_reg[27]/NET0131  ;
	input \P1_datao_reg[28]/NET0131  ;
	input \P1_datao_reg[29]/NET0131  ;
	input \P1_datao_reg[2]/NET0131  ;
	input \P1_datao_reg[30]/NET0131  ;
	input \P1_datao_reg[31]/NET0131  ;
	input \P1_datao_reg[3]/NET0131  ;
	input \P1_datao_reg[4]/NET0131  ;
	input \P1_datao_reg[5]/NET0131  ;
	input \P1_datao_reg[6]/NET0131  ;
	input \P1_datao_reg[7]/NET0131  ;
	input \P1_datao_reg[8]/NET0131  ;
	input \P1_datao_reg[9]/NET0131  ;
	input \P1_rd_reg/NET0131  ;
	input \P1_reg0_reg[0]/NET0131  ;
	input \P1_reg0_reg[10]/NET0131  ;
	input \P1_reg0_reg[11]/NET0131  ;
	input \P1_reg0_reg[12]/NET0131  ;
	input \P1_reg0_reg[13]/NET0131  ;
	input \P1_reg0_reg[14]/NET0131  ;
	input \P1_reg0_reg[15]/NET0131  ;
	input \P1_reg0_reg[16]/NET0131  ;
	input \P1_reg0_reg[17]/NET0131  ;
	input \P1_reg0_reg[18]/NET0131  ;
	input \P1_reg0_reg[19]/NET0131  ;
	input \P1_reg0_reg[1]/NET0131  ;
	input \P1_reg0_reg[20]/NET0131  ;
	input \P1_reg0_reg[21]/NET0131  ;
	input \P1_reg0_reg[22]/NET0131  ;
	input \P1_reg0_reg[23]/NET0131  ;
	input \P1_reg0_reg[24]/NET0131  ;
	input \P1_reg0_reg[25]/NET0131  ;
	input \P1_reg0_reg[26]/NET0131  ;
	input \P1_reg0_reg[27]/NET0131  ;
	input \P1_reg0_reg[28]/NET0131  ;
	input \P1_reg0_reg[29]/NET0131  ;
	input \P1_reg0_reg[2]/NET0131  ;
	input \P1_reg0_reg[30]/NET0131  ;
	input \P1_reg0_reg[31]/NET0131  ;
	input \P1_reg0_reg[3]/NET0131  ;
	input \P1_reg0_reg[4]/NET0131  ;
	input \P1_reg0_reg[5]/NET0131  ;
	input \P1_reg0_reg[6]/NET0131  ;
	input \P1_reg0_reg[7]/NET0131  ;
	input \P1_reg0_reg[8]/NET0131  ;
	input \P1_reg0_reg[9]/NET0131  ;
	input \P1_reg1_reg[0]/NET0131  ;
	input \P1_reg1_reg[10]/NET0131  ;
	input \P1_reg1_reg[11]/NET0131  ;
	input \P1_reg1_reg[12]/NET0131  ;
	input \P1_reg1_reg[13]/NET0131  ;
	input \P1_reg1_reg[14]/NET0131  ;
	input \P1_reg1_reg[15]/NET0131  ;
	input \P1_reg1_reg[16]/NET0131  ;
	input \P1_reg1_reg[17]/NET0131  ;
	input \P1_reg1_reg[18]/NET0131  ;
	input \P1_reg1_reg[19]/NET0131  ;
	input \P1_reg1_reg[1]/NET0131  ;
	input \P1_reg1_reg[20]/NET0131  ;
	input \P1_reg1_reg[21]/NET0131  ;
	input \P1_reg1_reg[22]/NET0131  ;
	input \P1_reg1_reg[23]/NET0131  ;
	input \P1_reg1_reg[24]/NET0131  ;
	input \P1_reg1_reg[25]/NET0131  ;
	input \P1_reg1_reg[26]/NET0131  ;
	input \P1_reg1_reg[27]/NET0131  ;
	input \P1_reg1_reg[28]/NET0131  ;
	input \P1_reg1_reg[29]/NET0131  ;
	input \P1_reg1_reg[2]/NET0131  ;
	input \P1_reg1_reg[30]/NET0131  ;
	input \P1_reg1_reg[31]/NET0131  ;
	input \P1_reg1_reg[3]/NET0131  ;
	input \P1_reg1_reg[4]/NET0131  ;
	input \P1_reg1_reg[5]/NET0131  ;
	input \P1_reg1_reg[6]/NET0131  ;
	input \P1_reg1_reg[7]/NET0131  ;
	input \P1_reg1_reg[8]/NET0131  ;
	input \P1_reg1_reg[9]/NET0131  ;
	input \P1_reg2_reg[0]/NET0131  ;
	input \P1_reg2_reg[10]/NET0131  ;
	input \P1_reg2_reg[11]/NET0131  ;
	input \P1_reg2_reg[12]/NET0131  ;
	input \P1_reg2_reg[13]/NET0131  ;
	input \P1_reg2_reg[14]/NET0131  ;
	input \P1_reg2_reg[15]/NET0131  ;
	input \P1_reg2_reg[16]/NET0131  ;
	input \P1_reg2_reg[17]/NET0131  ;
	input \P1_reg2_reg[18]/NET0131  ;
	input \P1_reg2_reg[19]/NET0131  ;
	input \P1_reg2_reg[1]/NET0131  ;
	input \P1_reg2_reg[20]/NET0131  ;
	input \P1_reg2_reg[21]/NET0131  ;
	input \P1_reg2_reg[22]/NET0131  ;
	input \P1_reg2_reg[23]/NET0131  ;
	input \P1_reg2_reg[24]/NET0131  ;
	input \P1_reg2_reg[25]/NET0131  ;
	input \P1_reg2_reg[26]/NET0131  ;
	input \P1_reg2_reg[27]/NET0131  ;
	input \P1_reg2_reg[28]/NET0131  ;
	input \P1_reg2_reg[29]/NET0131  ;
	input \P1_reg2_reg[2]/NET0131  ;
	input \P1_reg2_reg[30]/NET0131  ;
	input \P1_reg2_reg[31]/NET0131  ;
	input \P1_reg2_reg[3]/NET0131  ;
	input \P1_reg2_reg[4]/NET0131  ;
	input \P1_reg2_reg[5]/NET0131  ;
	input \P1_reg2_reg[6]/NET0131  ;
	input \P1_reg2_reg[7]/NET0131  ;
	input \P1_reg2_reg[8]/NET0131  ;
	input \P1_reg2_reg[9]/NET0131  ;
	input \P1_reg3_reg[0]/NET0131  ;
	input \P1_reg3_reg[10]/NET0131  ;
	input \P1_reg3_reg[11]/NET0131  ;
	input \P1_reg3_reg[12]/NET0131  ;
	input \P1_reg3_reg[13]/NET0131  ;
	input \P1_reg3_reg[14]/NET0131  ;
	input \P1_reg3_reg[15]/NET0131  ;
	input \P1_reg3_reg[16]/NET0131  ;
	input \P1_reg3_reg[17]/NET0131  ;
	input \P1_reg3_reg[18]/NET0131  ;
	input \P1_reg3_reg[19]/NET0131  ;
	input \P1_reg3_reg[1]/NET0131  ;
	input \P1_reg3_reg[20]/NET0131  ;
	input \P1_reg3_reg[21]/NET0131  ;
	input \P1_reg3_reg[22]/NET0131  ;
	input \P1_reg3_reg[23]/NET0131  ;
	input \P1_reg3_reg[24]/NET0131  ;
	input \P1_reg3_reg[25]/NET0131  ;
	input \P1_reg3_reg[26]/NET0131  ;
	input \P1_reg3_reg[27]/NET0131  ;
	input \P1_reg3_reg[28]/NET0131  ;
	input \P1_reg3_reg[2]/NET0131  ;
	input \P1_reg3_reg[3]/NET0131  ;
	input \P1_reg3_reg[4]/NET0131  ;
	input \P1_reg3_reg[5]/NET0131  ;
	input \P1_reg3_reg[6]/NET0131  ;
	input \P1_reg3_reg[7]/NET0131  ;
	input \P1_reg3_reg[8]/NET0131  ;
	input \P1_reg3_reg[9]/NET0131  ;
	input \P1_state_reg[0]/NET0131  ;
	input \P1_wr_reg/NET0131  ;
	input \P2_B_reg/NET0131  ;
	input \P2_IR_reg[0]/NET0131  ;
	input \P2_IR_reg[10]/NET0131  ;
	input \P2_IR_reg[11]/NET0131  ;
	input \P2_IR_reg[12]/NET0131  ;
	input \P2_IR_reg[13]/NET0131  ;
	input \P2_IR_reg[14]/NET0131  ;
	input \P2_IR_reg[15]/NET0131  ;
	input \P2_IR_reg[16]/NET0131  ;
	input \P2_IR_reg[17]/NET0131  ;
	input \P2_IR_reg[18]/NET0131  ;
	input \P2_IR_reg[19]/NET0131  ;
	input \P2_IR_reg[1]/NET0131  ;
	input \P2_IR_reg[20]/NET0131  ;
	input \P2_IR_reg[21]/NET0131  ;
	input \P2_IR_reg[22]/NET0131  ;
	input \P2_IR_reg[23]/NET0131  ;
	input \P2_IR_reg[24]/NET0131  ;
	input \P2_IR_reg[25]/NET0131  ;
	input \P2_IR_reg[26]/NET0131  ;
	input \P2_IR_reg[27]/NET0131  ;
	input \P2_IR_reg[28]/NET0131  ;
	input \P2_IR_reg[29]/NET0131  ;
	input \P2_IR_reg[2]/NET0131  ;
	input \P2_IR_reg[30]/NET0131  ;
	input \P2_IR_reg[31]/NET0131  ;
	input \P2_IR_reg[3]/NET0131  ;
	input \P2_IR_reg[4]/NET0131  ;
	input \P2_IR_reg[5]/NET0131  ;
	input \P2_IR_reg[6]/NET0131  ;
	input \P2_IR_reg[7]/NET0131  ;
	input \P2_IR_reg[8]/NET0131  ;
	input \P2_IR_reg[9]/NET0131  ;
	input \P2_addr_reg[0]/NET0131  ;
	input \P2_addr_reg[10]/NET0131  ;
	input \P2_addr_reg[11]/NET0131  ;
	input \P2_addr_reg[12]/NET0131  ;
	input \P2_addr_reg[13]/NET0131  ;
	input \P2_addr_reg[14]/NET0131  ;
	input \P2_addr_reg[15]/NET0131  ;
	input \P2_addr_reg[16]/NET0131  ;
	input \P2_addr_reg[17]/NET0131  ;
	input \P2_addr_reg[18]/NET0131  ;
	input \P2_addr_reg[19]/NET0131  ;
	input \P2_addr_reg[1]/NET0131  ;
	input \P2_addr_reg[2]/NET0131  ;
	input \P2_addr_reg[3]/NET0131  ;
	input \P2_addr_reg[4]/NET0131  ;
	input \P2_addr_reg[5]/NET0131  ;
	input \P2_addr_reg[6]/NET0131  ;
	input \P2_addr_reg[7]/NET0131  ;
	input \P2_addr_reg[8]/NET0131  ;
	input \P2_addr_reg[9]/NET0131  ;
	input \P2_d_reg[0]/NET0131  ;
	input \P2_d_reg[1]/NET0131  ;
	input \P2_datao_reg[0]/NET0131  ;
	input \P2_datao_reg[10]/NET0131  ;
	input \P2_datao_reg[11]/NET0131  ;
	input \P2_datao_reg[12]/NET0131  ;
	input \P2_datao_reg[13]/NET0131  ;
	input \P2_datao_reg[14]/NET0131  ;
	input \P2_datao_reg[15]/NET0131  ;
	input \P2_datao_reg[16]/NET0131  ;
	input \P2_datao_reg[17]/NET0131  ;
	input \P2_datao_reg[18]/NET0131  ;
	input \P2_datao_reg[19]/NET0131  ;
	input \P2_datao_reg[1]/NET0131  ;
	input \P2_datao_reg[20]/NET0131  ;
	input \P2_datao_reg[21]/NET0131  ;
	input \P2_datao_reg[22]/NET0131  ;
	input \P2_datao_reg[23]/NET0131  ;
	input \P2_datao_reg[24]/NET0131  ;
	input \P2_datao_reg[25]/NET0131  ;
	input \P2_datao_reg[26]/NET0131  ;
	input \P2_datao_reg[27]/NET0131  ;
	input \P2_datao_reg[28]/NET0131  ;
	input \P2_datao_reg[29]/NET0131  ;
	input \P2_datao_reg[2]/NET0131  ;
	input \P2_datao_reg[30]/NET0131  ;
	input \P2_datao_reg[31]/NET0131  ;
	input \P2_datao_reg[3]/NET0131  ;
	input \P2_datao_reg[4]/NET0131  ;
	input \P2_datao_reg[5]/NET0131  ;
	input \P2_datao_reg[6]/NET0131  ;
	input \P2_datao_reg[7]/NET0131  ;
	input \P2_datao_reg[8]/NET0131  ;
	input \P2_datao_reg[9]/NET0131  ;
	input \P2_rd_reg/NET0131  ;
	input \P2_reg0_reg[0]/NET0131  ;
	input \P2_reg0_reg[10]/NET0131  ;
	input \P2_reg0_reg[11]/NET0131  ;
	input \P2_reg0_reg[12]/NET0131  ;
	input \P2_reg0_reg[13]/NET0131  ;
	input \P2_reg0_reg[14]/NET0131  ;
	input \P2_reg0_reg[15]/NET0131  ;
	input \P2_reg0_reg[16]/NET0131  ;
	input \P2_reg0_reg[17]/NET0131  ;
	input \P2_reg0_reg[18]/NET0131  ;
	input \P2_reg0_reg[19]/NET0131  ;
	input \P2_reg0_reg[1]/NET0131  ;
	input \P2_reg0_reg[20]/NET0131  ;
	input \P2_reg0_reg[21]/NET0131  ;
	input \P2_reg0_reg[22]/NET0131  ;
	input \P2_reg0_reg[23]/NET0131  ;
	input \P2_reg0_reg[24]/NET0131  ;
	input \P2_reg0_reg[25]/NET0131  ;
	input \P2_reg0_reg[26]/NET0131  ;
	input \P2_reg0_reg[27]/NET0131  ;
	input \P2_reg0_reg[28]/NET0131  ;
	input \P2_reg0_reg[29]/NET0131  ;
	input \P2_reg0_reg[2]/NET0131  ;
	input \P2_reg0_reg[30]/NET0131  ;
	input \P2_reg0_reg[31]/NET0131  ;
	input \P2_reg0_reg[3]/NET0131  ;
	input \P2_reg0_reg[4]/NET0131  ;
	input \P2_reg0_reg[5]/NET0131  ;
	input \P2_reg0_reg[6]/NET0131  ;
	input \P2_reg0_reg[7]/NET0131  ;
	input \P2_reg0_reg[8]/NET0131  ;
	input \P2_reg0_reg[9]/NET0131  ;
	input \P2_reg1_reg[0]/NET0131  ;
	input \P2_reg1_reg[10]/NET0131  ;
	input \P2_reg1_reg[11]/NET0131  ;
	input \P2_reg1_reg[12]/NET0131  ;
	input \P2_reg1_reg[13]/NET0131  ;
	input \P2_reg1_reg[14]/NET0131  ;
	input \P2_reg1_reg[15]/NET0131  ;
	input \P2_reg1_reg[16]/NET0131  ;
	input \P2_reg1_reg[17]/NET0131  ;
	input \P2_reg1_reg[18]/NET0131  ;
	input \P2_reg1_reg[19]/NET0131  ;
	input \P2_reg1_reg[1]/NET0131  ;
	input \P2_reg1_reg[20]/NET0131  ;
	input \P2_reg1_reg[21]/NET0131  ;
	input \P2_reg1_reg[22]/NET0131  ;
	input \P2_reg1_reg[23]/NET0131  ;
	input \P2_reg1_reg[24]/NET0131  ;
	input \P2_reg1_reg[25]/NET0131  ;
	input \P2_reg1_reg[26]/NET0131  ;
	input \P2_reg1_reg[27]/NET0131  ;
	input \P2_reg1_reg[28]/NET0131  ;
	input \P2_reg1_reg[29]/NET0131  ;
	input \P2_reg1_reg[2]/NET0131  ;
	input \P2_reg1_reg[30]/NET0131  ;
	input \P2_reg1_reg[31]/NET0131  ;
	input \P2_reg1_reg[3]/NET0131  ;
	input \P2_reg1_reg[4]/NET0131  ;
	input \P2_reg1_reg[5]/NET0131  ;
	input \P2_reg1_reg[6]/NET0131  ;
	input \P2_reg1_reg[7]/NET0131  ;
	input \P2_reg1_reg[8]/NET0131  ;
	input \P2_reg1_reg[9]/NET0131  ;
	input \P2_reg2_reg[0]/NET0131  ;
	input \P2_reg2_reg[10]/NET0131  ;
	input \P2_reg2_reg[11]/NET0131  ;
	input \P2_reg2_reg[12]/NET0131  ;
	input \P2_reg2_reg[13]/NET0131  ;
	input \P2_reg2_reg[14]/NET0131  ;
	input \P2_reg2_reg[15]/NET0131  ;
	input \P2_reg2_reg[16]/NET0131  ;
	input \P2_reg2_reg[17]/NET0131  ;
	input \P2_reg2_reg[18]/NET0131  ;
	input \P2_reg2_reg[19]/NET0131  ;
	input \P2_reg2_reg[1]/NET0131  ;
	input \P2_reg2_reg[20]/NET0131  ;
	input \P2_reg2_reg[21]/NET0131  ;
	input \P2_reg2_reg[22]/NET0131  ;
	input \P2_reg2_reg[23]/NET0131  ;
	input \P2_reg2_reg[24]/NET0131  ;
	input \P2_reg2_reg[25]/NET0131  ;
	input \P2_reg2_reg[26]/NET0131  ;
	input \P2_reg2_reg[27]/NET0131  ;
	input \P2_reg2_reg[28]/NET0131  ;
	input \P2_reg2_reg[29]/NET0131  ;
	input \P2_reg2_reg[2]/NET0131  ;
	input \P2_reg2_reg[30]/NET0131  ;
	input \P2_reg2_reg[31]/NET0131  ;
	input \P2_reg2_reg[3]/NET0131  ;
	input \P2_reg2_reg[4]/NET0131  ;
	input \P2_reg2_reg[5]/NET0131  ;
	input \P2_reg2_reg[6]/NET0131  ;
	input \P2_reg2_reg[7]/NET0131  ;
	input \P2_reg2_reg[8]/NET0131  ;
	input \P2_reg2_reg[9]/NET0131  ;
	input \P2_reg3_reg[0]/NET0131  ;
	input \P2_reg3_reg[10]/NET0131  ;
	input \P2_reg3_reg[11]/NET0131  ;
	input \P2_reg3_reg[12]/NET0131  ;
	input \P2_reg3_reg[13]/NET0131  ;
	input \P2_reg3_reg[14]/NET0131  ;
	input \P2_reg3_reg[15]/NET0131  ;
	input \P2_reg3_reg[16]/NET0131  ;
	input \P2_reg3_reg[17]/NET0131  ;
	input \P2_reg3_reg[18]/NET0131  ;
	input \P2_reg3_reg[19]/NET0131  ;
	input \P2_reg3_reg[1]/NET0131  ;
	input \P2_reg3_reg[20]/NET0131  ;
	input \P2_reg3_reg[21]/NET0131  ;
	input \P2_reg3_reg[22]/NET0131  ;
	input \P2_reg3_reg[23]/NET0131  ;
	input \P2_reg3_reg[24]/NET0131  ;
	input \P2_reg3_reg[25]/NET0131  ;
	input \P2_reg3_reg[26]/NET0131  ;
	input \P2_reg3_reg[27]/NET0131  ;
	input \P2_reg3_reg[28]/NET0131  ;
	input \P2_reg3_reg[2]/NET0131  ;
	input \P2_reg3_reg[3]/NET0131  ;
	input \P2_reg3_reg[4]/NET0131  ;
	input \P2_reg3_reg[5]/NET0131  ;
	input \P2_reg3_reg[6]/NET0131  ;
	input \P2_reg3_reg[7]/NET0131  ;
	input \P2_reg3_reg[8]/NET0131  ;
	input \P2_reg3_reg[9]/NET0131  ;
	input \P2_wr_reg/NET0131  ;
	input \si[0]_pad  ;
	input \si[10]_pad  ;
	input \si[11]_pad  ;
	input \si[12]_pad  ;
	input \si[13]_pad  ;
	input \si[14]_pad  ;
	input \si[15]_pad  ;
	input \si[16]_pad  ;
	input \si[17]_pad  ;
	input \si[18]_pad  ;
	input \si[19]_pad  ;
	input \si[1]_pad  ;
	input \si[20]_pad  ;
	input \si[21]_pad  ;
	input \si[22]_pad  ;
	input \si[23]_pad  ;
	input \si[24]_pad  ;
	input \si[25]_pad  ;
	input \si[26]_pad  ;
	input \si[27]_pad  ;
	input \si[28]_pad  ;
	input \si[29]_pad  ;
	input \si[2]_pad  ;
	input \si[30]_pad  ;
	input \si[31]_pad  ;
	input \si[3]_pad  ;
	input \si[4]_pad  ;
	input \si[5]_pad  ;
	input \si[6]_pad  ;
	input \si[7]_pad  ;
	input \si[8]_pad  ;
	input \si[9]_pad  ;
	output \P1_state_reg[0]/NET0131_syn_2  ;
	output \_al_n0  ;
	output \_al_n1  ;
	output \g35/_0_  ;
	output \g73637/_0_  ;
	output \g73647/_0_  ;
	output \g73648/_0_  ;
	output \g73649/_0_  ;
	output \g73650/_0_  ;
	output \g73667/_0_  ;
	output \g73668/_0_  ;
	output \g73669/_0_  ;
	output \g73670/_0_  ;
	output \g73671/_0_  ;
	output \g73672/_0_  ;
	output \g73674/_0_  ;
	output \g73675/_0_  ;
	output \g73709/_0_  ;
	output \g73710/_0_  ;
	output \g73711/_0_  ;
	output \g73716/_0_  ;
	output \g73717/_0_  ;
	output \g73718/_0_  ;
	output \g73719/_0_  ;
	output \g73720/_0_  ;
	output \g73721/_0_  ;
	output \g73722/_0_  ;
	output \g73723/_0_  ;
	output \g73724/_0_  ;
	output \g73765/_0_  ;
	output \g73769/_0_  ;
	output \g73770/_0_  ;
	output \g73771/_0_  ;
	output \g73772/_0_  ;
	output \g73773/_0_  ;
	output \g73774/_0_  ;
	output \g73775/_0_  ;
	output \g73776/_0_  ;
	output \g73777/_0_  ;
	output \g73778/_0_  ;
	output \g73779/_0_  ;
	output \g73780/_0_  ;
	output \g73781/_0_  ;
	output \g73782/_0_  ;
	output \g73783/_0_  ;
	output \g73784/_0_  ;
	output \g73785/_0_  ;
	output \g73786/_0_  ;
	output \g73787/_0_  ;
	output \g73788/_0_  ;
	output \g73789/_0_  ;
	output \g73790/_0_  ;
	output \g73791/_0_  ;
	output \g73792/_0_  ;
	output \g73845/_0_  ;
	output \g73846/_0_  ;
	output \g73847/_0_  ;
	output \g73848/_0_  ;
	output \g73860/_0_  ;
	output \g73863/_0_  ;
	output \g73864/_0_  ;
	output \g73867/_0_  ;
	output \g73870/_0_  ;
	output \g73871/_0_  ;
	output \g73872/_0_  ;
	output \g73873/_0_  ;
	output \g73874/_0_  ;
	output \g73875/_0_  ;
	output \g73876/_0_  ;
	output \g73877/_0_  ;
	output \g73878/_0_  ;
	output \g73879/_0_  ;
	output \g73880/_0_  ;
	output \g73924/_0_  ;
	output \g73925/_0_  ;
	output \g73949/_0_  ;
	output \g73950/_0_  ;
	output \g73953/_0_  ;
	output \g73954/_0_  ;
	output \g73955/_0_  ;
	output \g73956/_0_  ;
	output \g73957/_0_  ;
	output \g73958/_0_  ;
	output \g73960/_0_  ;
	output \g73961/_0_  ;
	output \g73962/_0_  ;
	output \g73963/_0_  ;
	output \g73964/_0_  ;
	output \g73965/_0_  ;
	output \g73966/_0_  ;
	output \g73967/_0_  ;
	output \g73968/_0_  ;
	output \g73969/_0_  ;
	output \g73970/_0_  ;
	output \g73971/_0_  ;
	output \g73972/_0_  ;
	output \g73973/_0_  ;
	output \g73974/_0_  ;
	output \g73975/_0_  ;
	output \g73976/_0_  ;
	output \g73977/_0_  ;
	output \g73978/_0_  ;
	output \g73979/_0_  ;
	output \g73980/_0_  ;
	output \g74062/_0_  ;
	output \g74063/_0_  ;
	output \g74064/_0_  ;
	output \g74065/_0_  ;
	output \g74066/_0_  ;
	output \g74071/_0_  ;
	output \g74072/_0_  ;
	output \g74105/_0_  ;
	output \g74106/_0_  ;
	output \g74107/_0_  ;
	output \g74108/_0_  ;
	output \g74109/_0_  ;
	output \g74110/_0_  ;
	output \g74111/_0_  ;
	output \g74112/_0_  ;
	output \g74113/_0_  ;
	output \g74114/_0_  ;
	output \g74115/_0_  ;
	output \g74167/_0_  ;
	output \g74168/_0_  ;
	output \g74169/_0_  ;
	output \g74170/_0_  ;
	output \g74172/_0_  ;
	output \g74173/_0_  ;
	output \g74174/_0_  ;
	output \g74175/_0_  ;
	output \g74225/_0_  ;
	output \g74226/_0_  ;
	output \g74227/_0_  ;
	output \g74229/_0_  ;
	output \g74230/_0_  ;
	output \g74231/_0_  ;
	output \g74232/_0_  ;
	output \g74233/_0_  ;
	output \g74234/_0_  ;
	output \g74235/_0_  ;
	output \g74236/_0_  ;
	output \g74237/_0_  ;
	output \g74238/_0_  ;
	output \g74239/_0_  ;
	output \g74240/_0_  ;
	output \g74241/_0_  ;
	output \g74242/_0_  ;
	output \g74243/_0_  ;
	output \g74244/_0_  ;
	output \g74245/_0_  ;
	output \g74246/_0_  ;
	output \g74247/_0_  ;
	output \g74248/_0_  ;
	output \g74249/_0_  ;
	output \g74250/_0_  ;
	output \g74251/_0_  ;
	output \g74252/_0_  ;
	output \g74253/_0_  ;
	output \g74254/_0_  ;
	output \g74255/_0_  ;
	output \g74330/_0_  ;
	output \g74331/_0_  ;
	output \g74333/_0_  ;
	output \g74334/_0_  ;
	output \g74335/_0_  ;
	output \g74390/_0_  ;
	output \g74391/_0_  ;
	output \g74405/_0_  ;
	output \g74407/_0_  ;
	output \g74408/_0_  ;
	output \g74409/_0_  ;
	output \g74410/_0_  ;
	output \g74411/_0_  ;
	output \g74412/_0_  ;
	output \g74413/_0_  ;
	output \g74414/_0_  ;
	output \g74415/_0_  ;
	output \g74416/_0_  ;
	output \g74417/_0_  ;
	output \g74418/_0_  ;
	output \g74419/_0_  ;
	output \g74420/_0_  ;
	output \g74421/_0_  ;
	output \g74422/_0_  ;
	output \g74483/_0_  ;
	output \g74485/_0_  ;
	output \g74486/_0_  ;
	output \g74487/_0_  ;
	output \g74576/_0_  ;
	output \g74578/_0_  ;
	output \g74581/_0_  ;
	output \g74582/_0_  ;
	output \g74583/_0_  ;
	output \g74584/_0_  ;
	output \g74585/_0_  ;
	output \g74588/_0_  ;
	output \g74589/_0_  ;
	output \g74590/_0_  ;
	output \g74591/_0_  ;
	output \g74592/_0_  ;
	output \g74595/_0_  ;
	output \g74596/_0_  ;
	output \g74597/_0_  ;
	output \g74598/_0_  ;
	output \g74599/_0_  ;
	output \g74600/_0_  ;
	output \g74601/_0_  ;
	output \g74602/_0_  ;
	output \g74711/_0_  ;
	output \g74835/_0_  ;
	output \g74836/_0_  ;
	output \g74838/_0_  ;
	output \g74840/_0_  ;
	output \g74841/_0_  ;
	output \g74843/_0_  ;
	output \g74844/_0_  ;
	output \g74963/_0_  ;
	output \g75075/_0_  ;
	output \g75078/_0_  ;
	output \g75079/_0_  ;
	output \g75083/_0_  ;
	output \g75084/_0_  ;
	output \g75089/_0_  ;
	output \g75090/_0_  ;
	output \g75091/_0_  ;
	output \g75224/_0_  ;
	output \g75233/_0_  ;
	output \g75234/_0_  ;
	output \g75427/_0_  ;
	output \g75430/_0_  ;
	output \g75434/_0_  ;
	output \g75436/_0_  ;
	output \g75438/_0_  ;
	output \g75844/_0_  ;
	output \g75850/_0_  ;
	output \g75851/_0_  ;
	output \g75860/_0_  ;
	output \g75865/_0_  ;
	output \g75867/_0_  ;
	output \g76076/_0_  ;
	output \g76375/_0_  ;
	output \g76896/_0_  ;
	output \g76901/_0_  ;
	output \g76905/_0_  ;
	output \g77085/_0_  ;
	output \g77892/_0_  ;
	output \g77897/_0_  ;
	output \g77902/_0_  ;
	output \g78635/_0_  ;
	output \g78636/_0_  ;
	output \g78640/_0_  ;
	output \g78642/_0_  ;
	output \g78645/_0_  ;
	output \g78964/_0_  ;
	output \g83163/_3_  ;
	output \g83164/_3_  ;
	output \g83165/_3_  ;
	output \g83166/_3_  ;
	output \g83167/_3_  ;
	output \g83168/_3_  ;
	output \g83644/_0_  ;
	output \g83645/_0_  ;
	output \g83646/_0_  ;
	output \g83647/_0_  ;
	output \g83648/_0_  ;
	output \g83649/_0_  ;
	output \g83650/_0_  ;
	output \g83651/_0_  ;
	output \g83652/_0_  ;
	output \g83653/_0_  ;
	output \g83654/_0_  ;
	output \g83655/_0_  ;
	output \g83656/_0_  ;
	output \g83657/_0_  ;
	output \g83658/_0_  ;
	output \g83659/_0_  ;
	output \g83660/_0_  ;
	output \g83661/_0_  ;
	output \g83662/_0_  ;
	output \g83663/_0_  ;
	output \g83664/_0_  ;
	output \g83665/_0_  ;
	output \g83666/_0_  ;
	output \g83667/_3_  ;
	output \g83668/_0_  ;
	output \g83669/_0_  ;
	output \g83670/_0_  ;
	output \g83671/_0_  ;
	output \g83715/_3_  ;
	output \g83716/_3_  ;
	output \g83717/_3_  ;
	output \g83718/_3_  ;
	output \g83719/_3_  ;
	output \g83720/_3_  ;
	output \g83721/_3_  ;
	output \g83722/_3_  ;
	output \g83723/_3_  ;
	output \g83724/_3_  ;
	output \g83725/_0_  ;
	output \g83726/_3_  ;
	output \g83727/_3_  ;
	output \g83728/_3_  ;
	output \g83729/_3_  ;
	output \g83730/_3_  ;
	output \g83731/_3_  ;
	output \g83732/_3_  ;
	output \g83733/_3_  ;
	output \g83734/_3_  ;
	output \g83735/_0_  ;
	output \g83736/_0_  ;
	output \g83737/_0_  ;
	output \g83738/_3_  ;
	output \g83739/_3_  ;
	output \g83740/_0_  ;
	output \g83741/_3_  ;
	output \g83742/_3_  ;
	output \g84164/_0_  ;
	output \g84181/_0_  ;
	output \g85146/_0_  ;
	output \g85147/_0_  ;
	output \g85148/_0_  ;
	output \g85149/_0_  ;
	output \g85151/_0_  ;
	output \g85152/_0_  ;
	output \g85154/_0_  ;
	output \g85155/_0_  ;
	output \g85156/_0_  ;
	output \g85157/_0_  ;
	output \g85158/_0_  ;
	output \g85159/_0_  ;
	output \g85160/_0_  ;
	output \g85161/_0_  ;
	output \g85162/_0_  ;
	output \g85163/_0_  ;
	output \g85164/_0_  ;
	output \g85165/_0_  ;
	output \g85166/_0_  ;
	output \g85167/_0_  ;
	output \g85168/_0_  ;
	output \g85169/_0_  ;
	output \g85171/_0_  ;
	output \g85173/_0_  ;
	output \g85174/_0_  ;
	output \g85175/_0_  ;
	output \g85176/_0_  ;
	output \g85178/_0_  ;
	output \g85179/_0_  ;
	output \g85180/_0_  ;
	output \g85181/_0_  ;
	output \g85182/_0_  ;
	output \g85183/_0_  ;
	output \g85184/_0_  ;
	output \g85185/_0_  ;
	output \g85186/_0_  ;
	output \g85187/_0_  ;
	output \g85188/_0_  ;
	output \g85189/_0_  ;
	output \g85190/_0_  ;
	output \g85510/_0_  ;
	output \g85711/u3_syn_4  ;
	output \g85972/_0_  ;
	output \g86107/_0_  ;
	output \g86200/u3_syn_4  ;
	output \g86477/_0_  ;
	output \g86548/_0_  ;
	output \g86652/u3_syn_4  ;
	output \g86807/u3_syn_4  ;
	output \g87581/_0_  ;
	output \g88104/_0_  ;
	output \g88112/_0_  ;
	output \g88136/_0_  ;
	output \g88148/_0_  ;
	output \g88157/_0_  ;
	output \g88171/_0_  ;
	output \g88179/_0_  ;
	output \g88208/_0_  ;
	output \g88217/_0_  ;
	output \g88222/_0_  ;
	output \g88228/_0_  ;
	output \g88236/_0_  ;
	output \g88242/_0_  ;
	output \g88252_dup/_0_  ;
	output \g88253/_2_  ;
	output \g88259/_0_  ;
	output \g88274/_0_  ;
	output \g88286/_0_  ;
	output \g88296/_0_  ;
	output \g88306/_0_  ;
	output \g88319/_0_  ;
	output \g88330/_0_  ;
	output \g88370/_0_  ;
	output \g88375/_0_  ;
	output \g88388/_0_  ;
	output \g88397/_0_  ;
	output \g88404/_0_  ;
	output \g88793/_0_  ;
	output \g88834/_0_  ;
	output \g88905/_0_  ;
	output \g88910/_0_  ;
	output \g88936_dup/_0_  ;
	output \g88953/_0_  ;
	output \g88962/_0_  ;
	output \g89007/_0_  ;
	output \g89018/_0_  ;
	output \g89024/_0_  ;
	output \g89031/_0_  ;
	output \g89066/_0_  ;
	output \g89082/_0_  ;
	output \g89097/_0_  ;
	output \g90677/_1__syn_2  ;
	output \g96226/_0_  ;
	output \g96236/_0_  ;
	output \g96261/_0_  ;
	output \g96339/_0_  ;
	output \g96380/_1_  ;
	output \g96418/_0_  ;
	output \g96566/_1_  ;
	output \g96574/_0_  ;
	output \g96620/_0_  ;
	output \g96629/_0_  ;
	output \g96735/_0_  ;
	output \g96866/_0_  ;
	output \g96875/_0_  ;
	output \g96910/_0_  ;
	output \g96946/_0_  ;
	output \g96965/_0_  ;
	output \g97098/_0_  ;
	output \g97228/_0_  ;
	output \g97231/_0_  ;
	output \g97242/_0_  ;
	output \g97384/_0_  ;
	output \g97409/_0_  ;
	output \g97506/_0_  ;
	output \g97626/_0_  ;
	output rd_pad ;
	output \so[0]_pad  ;
	output \so[10]_pad  ;
	output \so[11]_pad  ;
	output \so[12]_pad  ;
	output \so[13]_pad  ;
	output \so[14]_pad  ;
	output \so[15]_pad  ;
	output \so[16]_pad  ;
	output \so[17]_pad  ;
	output \so[18]_pad  ;
	output \so[19]_pad  ;
	output \so[1]_pad  ;
	output \so[2]_pad  ;
	output \so[3]_pad  ;
	output \so[4]_pad  ;
	output \so[5]_pad  ;
	output \so[6]_pad  ;
	output \so[7]_pad  ;
	output \so[8]_pad  ;
	output \so[9]_pad  ;
	output wr_pad ;
	wire _w7356_ ;
	wire _w7355_ ;
	wire _w7354_ ;
	wire _w7353_ ;
	wire _w7352_ ;
	wire _w7351_ ;
	wire _w7350_ ;
	wire _w7349_ ;
	wire _w7348_ ;
	wire _w7347_ ;
	wire _w7346_ ;
	wire _w7345_ ;
	wire _w7344_ ;
	wire _w7343_ ;
	wire _w7342_ ;
	wire _w7341_ ;
	wire _w7340_ ;
	wire _w7339_ ;
	wire _w7338_ ;
	wire _w7337_ ;
	wire _w7336_ ;
	wire _w7335_ ;
	wire _w7334_ ;
	wire _w7333_ ;
	wire _w7332_ ;
	wire _w7331_ ;
	wire _w7330_ ;
	wire _w7329_ ;
	wire _w7328_ ;
	wire _w7327_ ;
	wire _w7326_ ;
	wire _w7325_ ;
	wire _w7324_ ;
	wire _w7323_ ;
	wire _w7322_ ;
	wire _w7321_ ;
	wire _w7320_ ;
	wire _w7319_ ;
	wire _w7318_ ;
	wire _w7317_ ;
	wire _w7316_ ;
	wire _w7315_ ;
	wire _w7314_ ;
	wire _w7313_ ;
	wire _w7312_ ;
	wire _w7311_ ;
	wire _w7310_ ;
	wire _w7309_ ;
	wire _w7308_ ;
	wire _w7307_ ;
	wire _w7306_ ;
	wire _w7305_ ;
	wire _w7304_ ;
	wire _w7303_ ;
	wire _w7302_ ;
	wire _w7301_ ;
	wire _w7300_ ;
	wire _w7299_ ;
	wire _w7298_ ;
	wire _w7297_ ;
	wire _w7296_ ;
	wire _w7295_ ;
	wire _w7294_ ;
	wire _w7293_ ;
	wire _w7292_ ;
	wire _w7291_ ;
	wire _w7290_ ;
	wire _w7289_ ;
	wire _w7288_ ;
	wire _w7287_ ;
	wire _w7286_ ;
	wire _w7285_ ;
	wire _w7284_ ;
	wire _w7283_ ;
	wire _w7282_ ;
	wire _w7281_ ;
	wire _w7280_ ;
	wire _w7279_ ;
	wire _w7278_ ;
	wire _w7277_ ;
	wire _w7276_ ;
	wire _w7275_ ;
	wire _w7274_ ;
	wire _w7273_ ;
	wire _w7272_ ;
	wire _w7271_ ;
	wire _w7270_ ;
	wire _w7269_ ;
	wire _w7268_ ;
	wire _w7267_ ;
	wire _w7266_ ;
	wire _w7265_ ;
	wire _w7264_ ;
	wire _w7263_ ;
	wire _w7262_ ;
	wire _w7261_ ;
	wire _w7260_ ;
	wire _w7259_ ;
	wire _w7258_ ;
	wire _w7257_ ;
	wire _w7256_ ;
	wire _w7255_ ;
	wire _w7254_ ;
	wire _w7253_ ;
	wire _w7252_ ;
	wire _w7251_ ;
	wire _w7250_ ;
	wire _w7249_ ;
	wire _w7248_ ;
	wire _w7247_ ;
	wire _w7246_ ;
	wire _w7245_ ;
	wire _w7244_ ;
	wire _w7243_ ;
	wire _w7242_ ;
	wire _w7241_ ;
	wire _w7240_ ;
	wire _w7239_ ;
	wire _w7238_ ;
	wire _w7237_ ;
	wire _w7236_ ;
	wire _w7235_ ;
	wire _w7234_ ;
	wire _w7233_ ;
	wire _w7232_ ;
	wire _w7231_ ;
	wire _w7230_ ;
	wire _w7229_ ;
	wire _w7228_ ;
	wire _w7227_ ;
	wire _w7226_ ;
	wire _w7225_ ;
	wire _w7224_ ;
	wire _w7223_ ;
	wire _w7222_ ;
	wire _w7221_ ;
	wire _w7220_ ;
	wire _w7219_ ;
	wire _w7218_ ;
	wire _w7217_ ;
	wire _w7216_ ;
	wire _w7215_ ;
	wire _w7214_ ;
	wire _w7213_ ;
	wire _w7212_ ;
	wire _w7211_ ;
	wire _w7210_ ;
	wire _w7209_ ;
	wire _w7208_ ;
	wire _w7207_ ;
	wire _w7206_ ;
	wire _w7205_ ;
	wire _w7204_ ;
	wire _w7203_ ;
	wire _w7202_ ;
	wire _w7201_ ;
	wire _w7200_ ;
	wire _w7199_ ;
	wire _w7198_ ;
	wire _w7197_ ;
	wire _w7196_ ;
	wire _w7195_ ;
	wire _w7194_ ;
	wire _w7193_ ;
	wire _w7192_ ;
	wire _w7191_ ;
	wire _w7190_ ;
	wire _w7189_ ;
	wire _w7188_ ;
	wire _w7187_ ;
	wire _w7186_ ;
	wire _w7185_ ;
	wire _w7184_ ;
	wire _w7183_ ;
	wire _w7182_ ;
	wire _w7181_ ;
	wire _w7180_ ;
	wire _w7179_ ;
	wire _w7178_ ;
	wire _w7177_ ;
	wire _w7176_ ;
	wire _w7175_ ;
	wire _w7174_ ;
	wire _w7173_ ;
	wire _w7172_ ;
	wire _w7171_ ;
	wire _w7170_ ;
	wire _w7169_ ;
	wire _w7168_ ;
	wire _w7167_ ;
	wire _w7166_ ;
	wire _w7165_ ;
	wire _w7164_ ;
	wire _w7163_ ;
	wire _w7162_ ;
	wire _w7161_ ;
	wire _w7160_ ;
	wire _w7159_ ;
	wire _w7158_ ;
	wire _w7157_ ;
	wire _w7156_ ;
	wire _w7155_ ;
	wire _w7154_ ;
	wire _w7153_ ;
	wire _w7152_ ;
	wire _w7151_ ;
	wire _w7150_ ;
	wire _w7149_ ;
	wire _w7148_ ;
	wire _w7147_ ;
	wire _w7146_ ;
	wire _w7145_ ;
	wire _w7144_ ;
	wire _w7143_ ;
	wire _w7142_ ;
	wire _w7141_ ;
	wire _w7140_ ;
	wire _w7139_ ;
	wire _w7138_ ;
	wire _w7137_ ;
	wire _w7136_ ;
	wire _w7135_ ;
	wire _w7134_ ;
	wire _w7133_ ;
	wire _w7132_ ;
	wire _w7131_ ;
	wire _w7130_ ;
	wire _w7129_ ;
	wire _w7128_ ;
	wire _w7127_ ;
	wire _w7126_ ;
	wire _w7125_ ;
	wire _w7124_ ;
	wire _w7123_ ;
	wire _w7122_ ;
	wire _w7121_ ;
	wire _w7120_ ;
	wire _w7119_ ;
	wire _w7118_ ;
	wire _w7117_ ;
	wire _w7116_ ;
	wire _w7115_ ;
	wire _w7114_ ;
	wire _w7113_ ;
	wire _w7112_ ;
	wire _w7111_ ;
	wire _w7110_ ;
	wire _w7109_ ;
	wire _w7108_ ;
	wire _w7107_ ;
	wire _w7106_ ;
	wire _w7105_ ;
	wire _w7104_ ;
	wire _w7103_ ;
	wire _w7102_ ;
	wire _w7101_ ;
	wire _w7100_ ;
	wire _w7099_ ;
	wire _w7098_ ;
	wire _w7097_ ;
	wire _w7096_ ;
	wire _w7095_ ;
	wire _w7094_ ;
	wire _w7093_ ;
	wire _w7092_ ;
	wire _w7091_ ;
	wire _w7090_ ;
	wire _w7089_ ;
	wire _w7088_ ;
	wire _w7087_ ;
	wire _w7086_ ;
	wire _w7085_ ;
	wire _w7084_ ;
	wire _w7083_ ;
	wire _w7082_ ;
	wire _w7081_ ;
	wire _w7080_ ;
	wire _w7079_ ;
	wire _w7078_ ;
	wire _w7077_ ;
	wire _w7076_ ;
	wire _w7075_ ;
	wire _w7074_ ;
	wire _w7073_ ;
	wire _w7072_ ;
	wire _w7071_ ;
	wire _w7070_ ;
	wire _w7069_ ;
	wire _w7068_ ;
	wire _w7067_ ;
	wire _w7066_ ;
	wire _w7065_ ;
	wire _w7064_ ;
	wire _w7063_ ;
	wire _w7062_ ;
	wire _w7061_ ;
	wire _w7060_ ;
	wire _w7059_ ;
	wire _w7058_ ;
	wire _w7057_ ;
	wire _w7056_ ;
	wire _w7055_ ;
	wire _w7054_ ;
	wire _w7053_ ;
	wire _w7052_ ;
	wire _w7051_ ;
	wire _w7050_ ;
	wire _w7049_ ;
	wire _w7048_ ;
	wire _w7047_ ;
	wire _w7046_ ;
	wire _w7045_ ;
	wire _w7044_ ;
	wire _w7043_ ;
	wire _w7042_ ;
	wire _w7041_ ;
	wire _w7040_ ;
	wire _w7039_ ;
	wire _w7038_ ;
	wire _w7037_ ;
	wire _w7036_ ;
	wire _w7035_ ;
	wire _w7034_ ;
	wire _w7033_ ;
	wire _w7032_ ;
	wire _w7031_ ;
	wire _w7030_ ;
	wire _w7029_ ;
	wire _w7028_ ;
	wire _w7027_ ;
	wire _w7026_ ;
	wire _w7025_ ;
	wire _w7024_ ;
	wire _w7023_ ;
	wire _w7022_ ;
	wire _w7021_ ;
	wire _w7020_ ;
	wire _w7019_ ;
	wire _w7018_ ;
	wire _w7017_ ;
	wire _w7016_ ;
	wire _w7015_ ;
	wire _w7014_ ;
	wire _w7013_ ;
	wire _w7012_ ;
	wire _w7011_ ;
	wire _w7010_ ;
	wire _w7009_ ;
	wire _w7008_ ;
	wire _w7007_ ;
	wire _w7006_ ;
	wire _w7005_ ;
	wire _w7004_ ;
	wire _w7003_ ;
	wire _w7002_ ;
	wire _w7001_ ;
	wire _w7000_ ;
	wire _w6999_ ;
	wire _w6998_ ;
	wire _w6997_ ;
	wire _w6996_ ;
	wire _w6995_ ;
	wire _w6994_ ;
	wire _w6993_ ;
	wire _w6992_ ;
	wire _w6991_ ;
	wire _w6990_ ;
	wire _w6989_ ;
	wire _w6988_ ;
	wire _w6987_ ;
	wire _w6986_ ;
	wire _w6985_ ;
	wire _w6984_ ;
	wire _w6983_ ;
	wire _w6982_ ;
	wire _w6981_ ;
	wire _w6980_ ;
	wire _w6979_ ;
	wire _w6978_ ;
	wire _w6977_ ;
	wire _w6976_ ;
	wire _w6975_ ;
	wire _w6974_ ;
	wire _w6973_ ;
	wire _w6972_ ;
	wire _w6971_ ;
	wire _w6970_ ;
	wire _w6969_ ;
	wire _w6968_ ;
	wire _w6967_ ;
	wire _w6966_ ;
	wire _w6965_ ;
	wire _w6964_ ;
	wire _w6963_ ;
	wire _w6962_ ;
	wire _w6961_ ;
	wire _w6960_ ;
	wire _w6959_ ;
	wire _w6958_ ;
	wire _w6957_ ;
	wire _w6956_ ;
	wire _w6955_ ;
	wire _w6954_ ;
	wire _w6953_ ;
	wire _w6952_ ;
	wire _w6951_ ;
	wire _w6950_ ;
	wire _w6949_ ;
	wire _w6948_ ;
	wire _w6947_ ;
	wire _w6946_ ;
	wire _w6945_ ;
	wire _w6944_ ;
	wire _w6943_ ;
	wire _w6942_ ;
	wire _w6941_ ;
	wire _w6940_ ;
	wire _w6939_ ;
	wire _w6938_ ;
	wire _w6937_ ;
	wire _w6936_ ;
	wire _w6935_ ;
	wire _w6934_ ;
	wire _w6933_ ;
	wire _w6932_ ;
	wire _w6931_ ;
	wire _w6930_ ;
	wire _w6929_ ;
	wire _w6928_ ;
	wire _w6927_ ;
	wire _w6926_ ;
	wire _w6925_ ;
	wire _w6924_ ;
	wire _w6923_ ;
	wire _w6922_ ;
	wire _w6921_ ;
	wire _w6920_ ;
	wire _w6919_ ;
	wire _w6918_ ;
	wire _w6917_ ;
	wire _w6916_ ;
	wire _w6915_ ;
	wire _w6914_ ;
	wire _w6913_ ;
	wire _w6912_ ;
	wire _w6911_ ;
	wire _w6910_ ;
	wire _w6909_ ;
	wire _w6908_ ;
	wire _w6907_ ;
	wire _w6906_ ;
	wire _w6905_ ;
	wire _w6904_ ;
	wire _w6903_ ;
	wire _w6902_ ;
	wire _w6901_ ;
	wire _w6900_ ;
	wire _w6899_ ;
	wire _w6898_ ;
	wire _w6897_ ;
	wire _w6896_ ;
	wire _w6895_ ;
	wire _w6894_ ;
	wire _w6893_ ;
	wire _w6892_ ;
	wire _w6891_ ;
	wire _w6890_ ;
	wire _w6889_ ;
	wire _w6888_ ;
	wire _w6887_ ;
	wire _w6886_ ;
	wire _w6885_ ;
	wire _w6884_ ;
	wire _w6883_ ;
	wire _w6882_ ;
	wire _w6881_ ;
	wire _w6880_ ;
	wire _w6879_ ;
	wire _w6878_ ;
	wire _w6877_ ;
	wire _w6876_ ;
	wire _w6875_ ;
	wire _w6874_ ;
	wire _w6873_ ;
	wire _w6872_ ;
	wire _w6871_ ;
	wire _w6870_ ;
	wire _w6869_ ;
	wire _w6868_ ;
	wire _w6867_ ;
	wire _w6866_ ;
	wire _w6865_ ;
	wire _w6864_ ;
	wire _w6863_ ;
	wire _w6862_ ;
	wire _w6861_ ;
	wire _w6860_ ;
	wire _w6859_ ;
	wire _w6858_ ;
	wire _w6857_ ;
	wire _w6856_ ;
	wire _w6855_ ;
	wire _w6854_ ;
	wire _w6853_ ;
	wire _w6852_ ;
	wire _w6851_ ;
	wire _w6850_ ;
	wire _w6849_ ;
	wire _w6848_ ;
	wire _w6847_ ;
	wire _w6846_ ;
	wire _w6845_ ;
	wire _w6844_ ;
	wire _w6843_ ;
	wire _w6842_ ;
	wire _w6841_ ;
	wire _w6840_ ;
	wire _w6839_ ;
	wire _w6838_ ;
	wire _w6837_ ;
	wire _w6836_ ;
	wire _w6835_ ;
	wire _w6834_ ;
	wire _w6833_ ;
	wire _w6832_ ;
	wire _w6831_ ;
	wire _w6830_ ;
	wire _w6829_ ;
	wire _w6828_ ;
	wire _w6827_ ;
	wire _w6826_ ;
	wire _w6825_ ;
	wire _w6824_ ;
	wire _w6823_ ;
	wire _w6822_ ;
	wire _w6821_ ;
	wire _w6820_ ;
	wire _w6819_ ;
	wire _w6818_ ;
	wire _w6817_ ;
	wire _w6816_ ;
	wire _w6815_ ;
	wire _w6814_ ;
	wire _w6813_ ;
	wire _w6812_ ;
	wire _w6811_ ;
	wire _w6810_ ;
	wire _w6809_ ;
	wire _w6808_ ;
	wire _w6807_ ;
	wire _w6806_ ;
	wire _w6805_ ;
	wire _w6804_ ;
	wire _w6803_ ;
	wire _w6802_ ;
	wire _w6801_ ;
	wire _w6800_ ;
	wire _w6799_ ;
	wire _w6798_ ;
	wire _w6797_ ;
	wire _w6796_ ;
	wire _w6795_ ;
	wire _w6794_ ;
	wire _w6793_ ;
	wire _w6792_ ;
	wire _w6791_ ;
	wire _w6790_ ;
	wire _w6789_ ;
	wire _w6788_ ;
	wire _w6787_ ;
	wire _w6786_ ;
	wire _w6785_ ;
	wire _w6784_ ;
	wire _w6783_ ;
	wire _w6782_ ;
	wire _w6781_ ;
	wire _w6780_ ;
	wire _w6779_ ;
	wire _w6778_ ;
	wire _w6777_ ;
	wire _w6776_ ;
	wire _w6775_ ;
	wire _w6774_ ;
	wire _w6773_ ;
	wire _w6772_ ;
	wire _w6771_ ;
	wire _w6770_ ;
	wire _w6769_ ;
	wire _w6768_ ;
	wire _w6767_ ;
	wire _w6766_ ;
	wire _w6765_ ;
	wire _w6764_ ;
	wire _w6763_ ;
	wire _w6762_ ;
	wire _w6761_ ;
	wire _w6760_ ;
	wire _w6759_ ;
	wire _w6758_ ;
	wire _w6757_ ;
	wire _w6756_ ;
	wire _w6755_ ;
	wire _w6754_ ;
	wire _w6753_ ;
	wire _w6752_ ;
	wire _w6751_ ;
	wire _w6750_ ;
	wire _w6749_ ;
	wire _w6748_ ;
	wire _w6747_ ;
	wire _w6746_ ;
	wire _w6745_ ;
	wire _w6744_ ;
	wire _w6743_ ;
	wire _w6742_ ;
	wire _w6741_ ;
	wire _w6740_ ;
	wire _w6739_ ;
	wire _w6738_ ;
	wire _w6737_ ;
	wire _w6736_ ;
	wire _w6735_ ;
	wire _w6734_ ;
	wire _w6733_ ;
	wire _w6732_ ;
	wire _w6731_ ;
	wire _w6730_ ;
	wire _w6729_ ;
	wire _w6728_ ;
	wire _w6727_ ;
	wire _w6726_ ;
	wire _w6725_ ;
	wire _w6724_ ;
	wire _w6723_ ;
	wire _w6722_ ;
	wire _w6721_ ;
	wire _w6720_ ;
	wire _w6719_ ;
	wire _w6718_ ;
	wire _w6717_ ;
	wire _w6716_ ;
	wire _w6715_ ;
	wire _w6714_ ;
	wire _w6713_ ;
	wire _w6712_ ;
	wire _w6711_ ;
	wire _w6710_ ;
	wire _w6709_ ;
	wire _w6708_ ;
	wire _w6707_ ;
	wire _w6706_ ;
	wire _w6705_ ;
	wire _w6704_ ;
	wire _w6703_ ;
	wire _w6702_ ;
	wire _w6701_ ;
	wire _w6700_ ;
	wire _w6699_ ;
	wire _w6698_ ;
	wire _w6697_ ;
	wire _w6696_ ;
	wire _w6695_ ;
	wire _w6694_ ;
	wire _w6693_ ;
	wire _w6692_ ;
	wire _w6691_ ;
	wire _w6690_ ;
	wire _w6689_ ;
	wire _w6688_ ;
	wire _w6687_ ;
	wire _w6686_ ;
	wire _w6685_ ;
	wire _w6684_ ;
	wire _w6683_ ;
	wire _w6682_ ;
	wire _w6681_ ;
	wire _w6680_ ;
	wire _w6679_ ;
	wire _w6678_ ;
	wire _w6677_ ;
	wire _w6676_ ;
	wire _w6675_ ;
	wire _w6674_ ;
	wire _w6673_ ;
	wire _w6672_ ;
	wire _w6671_ ;
	wire _w6670_ ;
	wire _w6669_ ;
	wire _w6668_ ;
	wire _w6667_ ;
	wire _w6666_ ;
	wire _w6665_ ;
	wire _w6664_ ;
	wire _w6663_ ;
	wire _w6662_ ;
	wire _w6661_ ;
	wire _w6660_ ;
	wire _w6659_ ;
	wire _w6658_ ;
	wire _w6657_ ;
	wire _w6656_ ;
	wire _w6655_ ;
	wire _w6654_ ;
	wire _w6653_ ;
	wire _w6652_ ;
	wire _w6651_ ;
	wire _w6650_ ;
	wire _w6649_ ;
	wire _w6648_ ;
	wire _w6647_ ;
	wire _w6646_ ;
	wire _w6645_ ;
	wire _w6644_ ;
	wire _w6643_ ;
	wire _w6642_ ;
	wire _w6641_ ;
	wire _w6640_ ;
	wire _w6639_ ;
	wire _w6638_ ;
	wire _w6637_ ;
	wire _w6636_ ;
	wire _w6635_ ;
	wire _w6634_ ;
	wire _w6633_ ;
	wire _w6632_ ;
	wire _w6631_ ;
	wire _w6630_ ;
	wire _w6629_ ;
	wire _w6628_ ;
	wire _w6627_ ;
	wire _w6626_ ;
	wire _w6625_ ;
	wire _w6624_ ;
	wire _w6623_ ;
	wire _w6622_ ;
	wire _w6621_ ;
	wire _w6620_ ;
	wire _w6619_ ;
	wire _w6618_ ;
	wire _w6617_ ;
	wire _w6616_ ;
	wire _w6615_ ;
	wire _w6614_ ;
	wire _w6613_ ;
	wire _w6612_ ;
	wire _w6611_ ;
	wire _w6610_ ;
	wire _w6609_ ;
	wire _w6608_ ;
	wire _w6607_ ;
	wire _w6606_ ;
	wire _w6605_ ;
	wire _w6604_ ;
	wire _w6603_ ;
	wire _w6602_ ;
	wire _w6601_ ;
	wire _w6600_ ;
	wire _w6599_ ;
	wire _w6598_ ;
	wire _w6597_ ;
	wire _w6596_ ;
	wire _w6595_ ;
	wire _w6594_ ;
	wire _w6593_ ;
	wire _w6592_ ;
	wire _w6591_ ;
	wire _w6590_ ;
	wire _w6589_ ;
	wire _w6588_ ;
	wire _w6587_ ;
	wire _w6586_ ;
	wire _w6585_ ;
	wire _w6584_ ;
	wire _w6583_ ;
	wire _w6582_ ;
	wire _w6581_ ;
	wire _w6580_ ;
	wire _w6579_ ;
	wire _w6578_ ;
	wire _w6577_ ;
	wire _w6576_ ;
	wire _w6575_ ;
	wire _w6574_ ;
	wire _w6573_ ;
	wire _w6572_ ;
	wire _w6571_ ;
	wire _w6570_ ;
	wire _w6569_ ;
	wire _w6568_ ;
	wire _w6567_ ;
	wire _w6566_ ;
	wire _w6565_ ;
	wire _w6564_ ;
	wire _w6563_ ;
	wire _w6562_ ;
	wire _w6561_ ;
	wire _w6560_ ;
	wire _w6559_ ;
	wire _w6558_ ;
	wire _w6557_ ;
	wire _w6556_ ;
	wire _w6555_ ;
	wire _w6554_ ;
	wire _w6553_ ;
	wire _w6552_ ;
	wire _w6551_ ;
	wire _w6550_ ;
	wire _w6549_ ;
	wire _w6548_ ;
	wire _w6547_ ;
	wire _w6546_ ;
	wire _w6545_ ;
	wire _w6544_ ;
	wire _w6543_ ;
	wire _w6542_ ;
	wire _w6541_ ;
	wire _w6540_ ;
	wire _w6539_ ;
	wire _w6538_ ;
	wire _w6537_ ;
	wire _w6536_ ;
	wire _w6535_ ;
	wire _w6534_ ;
	wire _w6533_ ;
	wire _w6532_ ;
	wire _w6531_ ;
	wire _w6530_ ;
	wire _w6529_ ;
	wire _w6528_ ;
	wire _w6527_ ;
	wire _w6526_ ;
	wire _w6525_ ;
	wire _w6524_ ;
	wire _w6523_ ;
	wire _w6522_ ;
	wire _w6521_ ;
	wire _w6520_ ;
	wire _w6519_ ;
	wire _w6518_ ;
	wire _w6517_ ;
	wire _w6516_ ;
	wire _w6515_ ;
	wire _w6514_ ;
	wire _w6513_ ;
	wire _w6512_ ;
	wire _w6511_ ;
	wire _w6510_ ;
	wire _w6509_ ;
	wire _w6508_ ;
	wire _w6507_ ;
	wire _w6506_ ;
	wire _w6505_ ;
	wire _w6504_ ;
	wire _w6503_ ;
	wire _w6502_ ;
	wire _w6501_ ;
	wire _w6500_ ;
	wire _w6499_ ;
	wire _w6498_ ;
	wire _w6497_ ;
	wire _w6496_ ;
	wire _w6495_ ;
	wire _w6494_ ;
	wire _w6493_ ;
	wire _w6492_ ;
	wire _w6491_ ;
	wire _w6490_ ;
	wire _w6489_ ;
	wire _w6488_ ;
	wire _w6487_ ;
	wire _w6486_ ;
	wire _w6485_ ;
	wire _w6484_ ;
	wire _w6483_ ;
	wire _w6482_ ;
	wire _w6481_ ;
	wire _w6480_ ;
	wire _w6479_ ;
	wire _w6478_ ;
	wire _w6477_ ;
	wire _w6476_ ;
	wire _w6475_ ;
	wire _w6474_ ;
	wire _w6473_ ;
	wire _w6472_ ;
	wire _w6471_ ;
	wire _w6470_ ;
	wire _w6469_ ;
	wire _w6468_ ;
	wire _w6467_ ;
	wire _w6466_ ;
	wire _w6465_ ;
	wire _w6464_ ;
	wire _w6463_ ;
	wire _w6462_ ;
	wire _w6461_ ;
	wire _w6460_ ;
	wire _w6459_ ;
	wire _w6458_ ;
	wire _w6457_ ;
	wire _w6456_ ;
	wire _w6455_ ;
	wire _w6454_ ;
	wire _w6453_ ;
	wire _w6452_ ;
	wire _w6451_ ;
	wire _w6450_ ;
	wire _w6449_ ;
	wire _w6448_ ;
	wire _w6447_ ;
	wire _w6446_ ;
	wire _w6445_ ;
	wire _w6444_ ;
	wire _w6443_ ;
	wire _w6442_ ;
	wire _w6441_ ;
	wire _w6440_ ;
	wire _w6439_ ;
	wire _w6438_ ;
	wire _w6437_ ;
	wire _w6436_ ;
	wire _w6435_ ;
	wire _w6434_ ;
	wire _w6433_ ;
	wire _w6432_ ;
	wire _w6431_ ;
	wire _w6430_ ;
	wire _w6429_ ;
	wire _w6428_ ;
	wire _w6427_ ;
	wire _w6426_ ;
	wire _w6425_ ;
	wire _w6424_ ;
	wire _w6423_ ;
	wire _w6422_ ;
	wire _w6421_ ;
	wire _w6420_ ;
	wire _w6419_ ;
	wire _w6418_ ;
	wire _w6417_ ;
	wire _w6416_ ;
	wire _w6415_ ;
	wire _w6414_ ;
	wire _w6413_ ;
	wire _w6412_ ;
	wire _w6411_ ;
	wire _w6410_ ;
	wire _w6409_ ;
	wire _w6408_ ;
	wire _w6407_ ;
	wire _w6406_ ;
	wire _w6405_ ;
	wire _w6404_ ;
	wire _w6403_ ;
	wire _w6402_ ;
	wire _w6401_ ;
	wire _w6400_ ;
	wire _w6399_ ;
	wire _w6398_ ;
	wire _w6397_ ;
	wire _w6396_ ;
	wire _w6395_ ;
	wire _w6394_ ;
	wire _w6393_ ;
	wire _w6392_ ;
	wire _w6391_ ;
	wire _w6390_ ;
	wire _w6389_ ;
	wire _w6388_ ;
	wire _w6387_ ;
	wire _w6386_ ;
	wire _w6385_ ;
	wire _w6384_ ;
	wire _w6383_ ;
	wire _w6382_ ;
	wire _w6381_ ;
	wire _w6380_ ;
	wire _w6379_ ;
	wire _w6378_ ;
	wire _w6377_ ;
	wire _w6376_ ;
	wire _w6375_ ;
	wire _w6374_ ;
	wire _w6373_ ;
	wire _w6372_ ;
	wire _w6371_ ;
	wire _w6370_ ;
	wire _w6369_ ;
	wire _w6368_ ;
	wire _w6367_ ;
	wire _w6366_ ;
	wire _w6365_ ;
	wire _w6364_ ;
	wire _w6363_ ;
	wire _w6362_ ;
	wire _w6361_ ;
	wire _w6360_ ;
	wire _w6359_ ;
	wire _w6358_ ;
	wire _w6357_ ;
	wire _w6356_ ;
	wire _w6355_ ;
	wire _w6354_ ;
	wire _w6353_ ;
	wire _w6352_ ;
	wire _w6351_ ;
	wire _w6350_ ;
	wire _w6349_ ;
	wire _w6348_ ;
	wire _w6347_ ;
	wire _w6346_ ;
	wire _w6345_ ;
	wire _w6344_ ;
	wire _w6343_ ;
	wire _w6342_ ;
	wire _w6341_ ;
	wire _w6340_ ;
	wire _w6339_ ;
	wire _w6338_ ;
	wire _w6337_ ;
	wire _w6336_ ;
	wire _w6335_ ;
	wire _w6334_ ;
	wire _w6333_ ;
	wire _w6332_ ;
	wire _w6331_ ;
	wire _w6330_ ;
	wire _w6329_ ;
	wire _w6328_ ;
	wire _w6327_ ;
	wire _w6326_ ;
	wire _w6325_ ;
	wire _w6324_ ;
	wire _w6323_ ;
	wire _w6322_ ;
	wire _w6321_ ;
	wire _w6320_ ;
	wire _w6319_ ;
	wire _w6318_ ;
	wire _w6317_ ;
	wire _w6316_ ;
	wire _w6315_ ;
	wire _w6314_ ;
	wire _w6313_ ;
	wire _w6312_ ;
	wire _w6311_ ;
	wire _w6310_ ;
	wire _w6309_ ;
	wire _w6308_ ;
	wire _w6307_ ;
	wire _w6306_ ;
	wire _w6305_ ;
	wire _w6304_ ;
	wire _w6303_ ;
	wire _w6302_ ;
	wire _w6301_ ;
	wire _w6300_ ;
	wire _w6299_ ;
	wire _w6298_ ;
	wire _w6297_ ;
	wire _w6296_ ;
	wire _w6295_ ;
	wire _w6294_ ;
	wire _w6293_ ;
	wire _w6292_ ;
	wire _w6291_ ;
	wire _w6290_ ;
	wire _w6289_ ;
	wire _w6288_ ;
	wire _w6287_ ;
	wire _w6286_ ;
	wire _w6285_ ;
	wire _w6284_ ;
	wire _w6283_ ;
	wire _w6282_ ;
	wire _w6281_ ;
	wire _w6280_ ;
	wire _w6279_ ;
	wire _w6278_ ;
	wire _w6277_ ;
	wire _w6276_ ;
	wire _w6275_ ;
	wire _w6274_ ;
	wire _w6273_ ;
	wire _w6272_ ;
	wire _w6271_ ;
	wire _w6270_ ;
	wire _w6269_ ;
	wire _w6268_ ;
	wire _w6267_ ;
	wire _w6266_ ;
	wire _w6265_ ;
	wire _w6264_ ;
	wire _w6263_ ;
	wire _w6262_ ;
	wire _w6261_ ;
	wire _w6260_ ;
	wire _w6259_ ;
	wire _w6258_ ;
	wire _w6257_ ;
	wire _w6256_ ;
	wire _w6255_ ;
	wire _w6254_ ;
	wire _w6253_ ;
	wire _w6252_ ;
	wire _w6251_ ;
	wire _w6250_ ;
	wire _w6249_ ;
	wire _w6248_ ;
	wire _w6247_ ;
	wire _w6246_ ;
	wire _w6245_ ;
	wire _w6244_ ;
	wire _w6243_ ;
	wire _w6242_ ;
	wire _w6241_ ;
	wire _w6240_ ;
	wire _w6239_ ;
	wire _w6238_ ;
	wire _w6237_ ;
	wire _w6236_ ;
	wire _w6235_ ;
	wire _w6234_ ;
	wire _w6233_ ;
	wire _w6232_ ;
	wire _w6231_ ;
	wire _w6230_ ;
	wire _w6229_ ;
	wire _w6228_ ;
	wire _w6227_ ;
	wire _w6226_ ;
	wire _w6225_ ;
	wire _w6224_ ;
	wire _w6223_ ;
	wire _w6222_ ;
	wire _w6221_ ;
	wire _w6220_ ;
	wire _w6219_ ;
	wire _w6218_ ;
	wire _w6217_ ;
	wire _w6216_ ;
	wire _w6215_ ;
	wire _w6214_ ;
	wire _w6213_ ;
	wire _w6212_ ;
	wire _w6211_ ;
	wire _w6210_ ;
	wire _w6209_ ;
	wire _w6208_ ;
	wire _w6207_ ;
	wire _w6206_ ;
	wire _w6205_ ;
	wire _w6204_ ;
	wire _w6203_ ;
	wire _w6202_ ;
	wire _w6201_ ;
	wire _w6200_ ;
	wire _w6199_ ;
	wire _w6198_ ;
	wire _w6197_ ;
	wire _w6196_ ;
	wire _w6195_ ;
	wire _w6194_ ;
	wire _w6193_ ;
	wire _w6192_ ;
	wire _w6191_ ;
	wire _w6190_ ;
	wire _w6189_ ;
	wire _w6188_ ;
	wire _w6187_ ;
	wire _w6186_ ;
	wire _w6185_ ;
	wire _w6184_ ;
	wire _w6183_ ;
	wire _w6182_ ;
	wire _w6181_ ;
	wire _w6180_ ;
	wire _w6179_ ;
	wire _w6178_ ;
	wire _w6177_ ;
	wire _w6176_ ;
	wire _w6175_ ;
	wire _w6174_ ;
	wire _w6173_ ;
	wire _w6172_ ;
	wire _w6171_ ;
	wire _w6170_ ;
	wire _w6169_ ;
	wire _w6168_ ;
	wire _w6167_ ;
	wire _w6166_ ;
	wire _w6165_ ;
	wire _w6164_ ;
	wire _w6163_ ;
	wire _w6162_ ;
	wire _w6161_ ;
	wire _w6160_ ;
	wire _w6159_ ;
	wire _w6158_ ;
	wire _w6157_ ;
	wire _w6156_ ;
	wire _w6155_ ;
	wire _w6154_ ;
	wire _w6153_ ;
	wire _w6152_ ;
	wire _w6151_ ;
	wire _w6150_ ;
	wire _w6149_ ;
	wire _w6148_ ;
	wire _w6147_ ;
	wire _w6146_ ;
	wire _w6145_ ;
	wire _w6144_ ;
	wire _w6143_ ;
	wire _w6142_ ;
	wire _w6141_ ;
	wire _w6140_ ;
	wire _w6139_ ;
	wire _w6138_ ;
	wire _w6137_ ;
	wire _w6136_ ;
	wire _w6135_ ;
	wire _w6134_ ;
	wire _w6133_ ;
	wire _w6132_ ;
	wire _w6131_ ;
	wire _w6130_ ;
	wire _w6129_ ;
	wire _w6128_ ;
	wire _w6127_ ;
	wire _w6126_ ;
	wire _w6125_ ;
	wire _w6124_ ;
	wire _w6123_ ;
	wire _w6122_ ;
	wire _w6121_ ;
	wire _w6120_ ;
	wire _w6119_ ;
	wire _w6118_ ;
	wire _w6117_ ;
	wire _w6116_ ;
	wire _w6115_ ;
	wire _w6114_ ;
	wire _w6113_ ;
	wire _w6112_ ;
	wire _w6111_ ;
	wire _w6110_ ;
	wire _w6109_ ;
	wire _w6108_ ;
	wire _w6107_ ;
	wire _w6106_ ;
	wire _w6105_ ;
	wire _w6104_ ;
	wire _w6103_ ;
	wire _w6102_ ;
	wire _w6101_ ;
	wire _w6100_ ;
	wire _w6099_ ;
	wire _w6098_ ;
	wire _w6097_ ;
	wire _w6096_ ;
	wire _w6095_ ;
	wire _w6094_ ;
	wire _w6093_ ;
	wire _w6092_ ;
	wire _w6091_ ;
	wire _w6090_ ;
	wire _w6089_ ;
	wire _w6088_ ;
	wire _w6087_ ;
	wire _w6086_ ;
	wire _w6085_ ;
	wire _w6084_ ;
	wire _w6083_ ;
	wire _w6082_ ;
	wire _w6081_ ;
	wire _w6080_ ;
	wire _w6079_ ;
	wire _w6078_ ;
	wire _w6077_ ;
	wire _w6076_ ;
	wire _w6075_ ;
	wire _w6074_ ;
	wire _w6073_ ;
	wire _w6072_ ;
	wire _w6071_ ;
	wire _w6070_ ;
	wire _w6069_ ;
	wire _w6068_ ;
	wire _w6067_ ;
	wire _w6066_ ;
	wire _w6065_ ;
	wire _w6064_ ;
	wire _w6063_ ;
	wire _w6062_ ;
	wire _w6061_ ;
	wire _w6060_ ;
	wire _w6059_ ;
	wire _w6058_ ;
	wire _w6057_ ;
	wire _w6056_ ;
	wire _w6055_ ;
	wire _w6054_ ;
	wire _w6053_ ;
	wire _w6052_ ;
	wire _w6051_ ;
	wire _w6050_ ;
	wire _w6049_ ;
	wire _w6048_ ;
	wire _w6047_ ;
	wire _w6046_ ;
	wire _w6045_ ;
	wire _w6044_ ;
	wire _w6043_ ;
	wire _w6042_ ;
	wire _w6041_ ;
	wire _w6040_ ;
	wire _w6039_ ;
	wire _w6038_ ;
	wire _w6037_ ;
	wire _w6036_ ;
	wire _w6035_ ;
	wire _w6034_ ;
	wire _w6033_ ;
	wire _w6032_ ;
	wire _w6031_ ;
	wire _w6030_ ;
	wire _w6029_ ;
	wire _w6028_ ;
	wire _w6027_ ;
	wire _w6026_ ;
	wire _w6025_ ;
	wire _w6024_ ;
	wire _w6023_ ;
	wire _w6022_ ;
	wire _w6021_ ;
	wire _w6020_ ;
	wire _w6019_ ;
	wire _w6018_ ;
	wire _w6017_ ;
	wire _w6016_ ;
	wire _w6015_ ;
	wire _w6014_ ;
	wire _w6013_ ;
	wire _w6012_ ;
	wire _w6011_ ;
	wire _w6010_ ;
	wire _w6009_ ;
	wire _w6008_ ;
	wire _w6007_ ;
	wire _w6006_ ;
	wire _w6005_ ;
	wire _w6004_ ;
	wire _w6003_ ;
	wire _w6002_ ;
	wire _w6001_ ;
	wire _w6000_ ;
	wire _w5999_ ;
	wire _w5998_ ;
	wire _w5997_ ;
	wire _w5996_ ;
	wire _w5995_ ;
	wire _w5994_ ;
	wire _w5993_ ;
	wire _w5992_ ;
	wire _w5991_ ;
	wire _w5990_ ;
	wire _w5989_ ;
	wire _w5988_ ;
	wire _w5987_ ;
	wire _w5986_ ;
	wire _w5985_ ;
	wire _w5984_ ;
	wire _w5983_ ;
	wire _w5982_ ;
	wire _w5981_ ;
	wire _w5980_ ;
	wire _w5979_ ;
	wire _w5978_ ;
	wire _w5977_ ;
	wire _w5976_ ;
	wire _w5975_ ;
	wire _w5974_ ;
	wire _w5973_ ;
	wire _w5972_ ;
	wire _w5971_ ;
	wire _w5970_ ;
	wire _w5969_ ;
	wire _w5968_ ;
	wire _w5967_ ;
	wire _w5966_ ;
	wire _w5965_ ;
	wire _w5964_ ;
	wire _w5963_ ;
	wire _w5962_ ;
	wire _w5961_ ;
	wire _w5960_ ;
	wire _w5959_ ;
	wire _w5958_ ;
	wire _w5957_ ;
	wire _w5956_ ;
	wire _w5955_ ;
	wire _w5954_ ;
	wire _w5953_ ;
	wire _w5952_ ;
	wire _w5951_ ;
	wire _w5950_ ;
	wire _w5949_ ;
	wire _w5948_ ;
	wire _w5947_ ;
	wire _w5946_ ;
	wire _w5945_ ;
	wire _w5944_ ;
	wire _w5943_ ;
	wire _w5942_ ;
	wire _w5941_ ;
	wire _w5940_ ;
	wire _w5939_ ;
	wire _w5938_ ;
	wire _w5937_ ;
	wire _w5936_ ;
	wire _w5935_ ;
	wire _w5934_ ;
	wire _w5933_ ;
	wire _w5932_ ;
	wire _w5931_ ;
	wire _w5930_ ;
	wire _w5929_ ;
	wire _w5928_ ;
	wire _w5927_ ;
	wire _w5926_ ;
	wire _w5925_ ;
	wire _w5924_ ;
	wire _w5923_ ;
	wire _w5922_ ;
	wire _w5921_ ;
	wire _w5920_ ;
	wire _w5919_ ;
	wire _w5918_ ;
	wire _w5917_ ;
	wire _w5916_ ;
	wire _w5915_ ;
	wire _w5914_ ;
	wire _w5913_ ;
	wire _w5912_ ;
	wire _w5911_ ;
	wire _w5910_ ;
	wire _w5909_ ;
	wire _w5908_ ;
	wire _w5907_ ;
	wire _w5906_ ;
	wire _w5905_ ;
	wire _w5904_ ;
	wire _w5903_ ;
	wire _w5902_ ;
	wire _w5901_ ;
	wire _w5900_ ;
	wire _w5899_ ;
	wire _w5898_ ;
	wire _w5897_ ;
	wire _w5896_ ;
	wire _w5895_ ;
	wire _w5894_ ;
	wire _w5893_ ;
	wire _w5892_ ;
	wire _w5891_ ;
	wire _w5890_ ;
	wire _w5889_ ;
	wire _w5888_ ;
	wire _w5887_ ;
	wire _w5886_ ;
	wire _w5885_ ;
	wire _w5884_ ;
	wire _w5883_ ;
	wire _w5882_ ;
	wire _w5881_ ;
	wire _w5880_ ;
	wire _w5879_ ;
	wire _w5878_ ;
	wire _w5877_ ;
	wire _w5876_ ;
	wire _w5875_ ;
	wire _w5874_ ;
	wire _w5873_ ;
	wire _w5872_ ;
	wire _w5871_ ;
	wire _w5870_ ;
	wire _w5869_ ;
	wire _w5868_ ;
	wire _w5867_ ;
	wire _w5866_ ;
	wire _w5865_ ;
	wire _w5864_ ;
	wire _w5863_ ;
	wire _w5862_ ;
	wire _w5861_ ;
	wire _w5860_ ;
	wire _w5859_ ;
	wire _w5858_ ;
	wire _w5857_ ;
	wire _w5856_ ;
	wire _w5855_ ;
	wire _w5854_ ;
	wire _w5853_ ;
	wire _w5852_ ;
	wire _w5851_ ;
	wire _w5850_ ;
	wire _w5849_ ;
	wire _w5848_ ;
	wire _w5847_ ;
	wire _w5846_ ;
	wire _w5845_ ;
	wire _w5844_ ;
	wire _w5843_ ;
	wire _w5842_ ;
	wire _w5841_ ;
	wire _w5840_ ;
	wire _w5839_ ;
	wire _w5838_ ;
	wire _w5837_ ;
	wire _w5836_ ;
	wire _w5835_ ;
	wire _w5834_ ;
	wire _w5833_ ;
	wire _w5832_ ;
	wire _w5831_ ;
	wire _w5830_ ;
	wire _w5829_ ;
	wire _w5828_ ;
	wire _w5827_ ;
	wire _w5826_ ;
	wire _w5825_ ;
	wire _w5824_ ;
	wire _w5823_ ;
	wire _w5822_ ;
	wire _w5821_ ;
	wire _w5820_ ;
	wire _w5819_ ;
	wire _w5818_ ;
	wire _w5817_ ;
	wire _w5816_ ;
	wire _w5815_ ;
	wire _w5814_ ;
	wire _w5813_ ;
	wire _w5812_ ;
	wire _w5811_ ;
	wire _w5810_ ;
	wire _w5809_ ;
	wire _w5808_ ;
	wire _w5807_ ;
	wire _w5806_ ;
	wire _w5805_ ;
	wire _w5804_ ;
	wire _w5803_ ;
	wire _w5802_ ;
	wire _w5801_ ;
	wire _w5800_ ;
	wire _w5799_ ;
	wire _w5798_ ;
	wire _w5797_ ;
	wire _w5796_ ;
	wire _w5795_ ;
	wire _w5794_ ;
	wire _w5793_ ;
	wire _w5792_ ;
	wire _w5791_ ;
	wire _w5790_ ;
	wire _w5789_ ;
	wire _w5788_ ;
	wire _w5787_ ;
	wire _w5786_ ;
	wire _w5785_ ;
	wire _w5784_ ;
	wire _w5783_ ;
	wire _w5782_ ;
	wire _w5781_ ;
	wire _w5780_ ;
	wire _w5779_ ;
	wire _w5778_ ;
	wire _w5777_ ;
	wire _w5776_ ;
	wire _w5775_ ;
	wire _w5774_ ;
	wire _w5773_ ;
	wire _w5772_ ;
	wire _w5771_ ;
	wire _w5770_ ;
	wire _w5769_ ;
	wire _w5768_ ;
	wire _w5767_ ;
	wire _w5766_ ;
	wire _w5765_ ;
	wire _w5764_ ;
	wire _w5763_ ;
	wire _w5762_ ;
	wire _w5761_ ;
	wire _w5760_ ;
	wire _w5759_ ;
	wire _w5758_ ;
	wire _w5757_ ;
	wire _w5756_ ;
	wire _w5755_ ;
	wire _w5754_ ;
	wire _w5753_ ;
	wire _w5752_ ;
	wire _w5751_ ;
	wire _w5750_ ;
	wire _w5749_ ;
	wire _w5748_ ;
	wire _w5747_ ;
	wire _w5746_ ;
	wire _w5745_ ;
	wire _w5744_ ;
	wire _w5743_ ;
	wire _w5742_ ;
	wire _w5741_ ;
	wire _w5740_ ;
	wire _w5739_ ;
	wire _w5738_ ;
	wire _w5737_ ;
	wire _w5736_ ;
	wire _w5735_ ;
	wire _w5734_ ;
	wire _w5733_ ;
	wire _w5732_ ;
	wire _w5731_ ;
	wire _w5730_ ;
	wire _w5729_ ;
	wire _w5728_ ;
	wire _w5727_ ;
	wire _w5726_ ;
	wire _w5725_ ;
	wire _w5724_ ;
	wire _w5723_ ;
	wire _w5722_ ;
	wire _w5721_ ;
	wire _w5720_ ;
	wire _w5719_ ;
	wire _w5718_ ;
	wire _w5717_ ;
	wire _w5716_ ;
	wire _w5715_ ;
	wire _w5714_ ;
	wire _w5713_ ;
	wire _w5712_ ;
	wire _w5711_ ;
	wire _w5710_ ;
	wire _w5709_ ;
	wire _w5708_ ;
	wire _w5707_ ;
	wire _w5706_ ;
	wire _w5705_ ;
	wire _w5704_ ;
	wire _w5703_ ;
	wire _w5702_ ;
	wire _w5701_ ;
	wire _w5700_ ;
	wire _w5699_ ;
	wire _w5698_ ;
	wire _w5697_ ;
	wire _w5696_ ;
	wire _w5695_ ;
	wire _w5694_ ;
	wire _w5693_ ;
	wire _w5692_ ;
	wire _w5691_ ;
	wire _w5690_ ;
	wire _w5689_ ;
	wire _w5688_ ;
	wire _w5687_ ;
	wire _w5686_ ;
	wire _w5685_ ;
	wire _w5684_ ;
	wire _w5683_ ;
	wire _w5682_ ;
	wire _w5681_ ;
	wire _w5680_ ;
	wire _w5679_ ;
	wire _w5678_ ;
	wire _w5677_ ;
	wire _w5676_ ;
	wire _w5675_ ;
	wire _w5674_ ;
	wire _w5673_ ;
	wire _w5672_ ;
	wire _w5671_ ;
	wire _w5670_ ;
	wire _w5669_ ;
	wire _w5668_ ;
	wire _w5667_ ;
	wire _w5666_ ;
	wire _w5665_ ;
	wire _w5664_ ;
	wire _w5663_ ;
	wire _w5662_ ;
	wire _w5661_ ;
	wire _w5660_ ;
	wire _w5659_ ;
	wire _w5658_ ;
	wire _w5657_ ;
	wire _w5656_ ;
	wire _w5655_ ;
	wire _w5654_ ;
	wire _w5653_ ;
	wire _w5652_ ;
	wire _w5651_ ;
	wire _w5650_ ;
	wire _w5649_ ;
	wire _w5648_ ;
	wire _w5647_ ;
	wire _w5646_ ;
	wire _w5645_ ;
	wire _w5644_ ;
	wire _w5643_ ;
	wire _w5642_ ;
	wire _w5641_ ;
	wire _w5640_ ;
	wire _w5639_ ;
	wire _w5638_ ;
	wire _w5637_ ;
	wire _w5636_ ;
	wire _w5635_ ;
	wire _w5634_ ;
	wire _w5633_ ;
	wire _w5632_ ;
	wire _w5631_ ;
	wire _w5630_ ;
	wire _w5629_ ;
	wire _w5628_ ;
	wire _w5627_ ;
	wire _w5626_ ;
	wire _w5625_ ;
	wire _w5624_ ;
	wire _w5623_ ;
	wire _w5622_ ;
	wire _w5621_ ;
	wire _w5620_ ;
	wire _w5619_ ;
	wire _w5618_ ;
	wire _w5617_ ;
	wire _w5616_ ;
	wire _w5615_ ;
	wire _w5614_ ;
	wire _w5613_ ;
	wire _w5612_ ;
	wire _w5611_ ;
	wire _w5610_ ;
	wire _w5609_ ;
	wire _w5608_ ;
	wire _w5607_ ;
	wire _w5606_ ;
	wire _w5605_ ;
	wire _w5604_ ;
	wire _w5603_ ;
	wire _w5602_ ;
	wire _w5601_ ;
	wire _w5600_ ;
	wire _w5599_ ;
	wire _w5598_ ;
	wire _w5597_ ;
	wire _w5596_ ;
	wire _w5595_ ;
	wire _w5594_ ;
	wire _w5593_ ;
	wire _w5592_ ;
	wire _w5591_ ;
	wire _w5590_ ;
	wire _w5589_ ;
	wire _w5588_ ;
	wire _w5587_ ;
	wire _w5586_ ;
	wire _w5585_ ;
	wire _w5584_ ;
	wire _w5583_ ;
	wire _w5582_ ;
	wire _w5581_ ;
	wire _w5580_ ;
	wire _w5579_ ;
	wire _w5578_ ;
	wire _w5577_ ;
	wire _w5576_ ;
	wire _w5575_ ;
	wire _w5574_ ;
	wire _w5573_ ;
	wire _w5572_ ;
	wire _w5571_ ;
	wire _w5570_ ;
	wire _w5569_ ;
	wire _w5568_ ;
	wire _w5567_ ;
	wire _w5566_ ;
	wire _w5565_ ;
	wire _w5564_ ;
	wire _w5563_ ;
	wire _w5562_ ;
	wire _w5561_ ;
	wire _w5560_ ;
	wire _w5559_ ;
	wire _w5558_ ;
	wire _w5557_ ;
	wire _w5556_ ;
	wire _w5555_ ;
	wire _w5554_ ;
	wire _w5553_ ;
	wire _w5552_ ;
	wire _w5551_ ;
	wire _w5550_ ;
	wire _w2819_ ;
	wire _w2818_ ;
	wire _w2817_ ;
	wire _w2816_ ;
	wire _w2815_ ;
	wire _w2814_ ;
	wire _w2813_ ;
	wire _w2812_ ;
	wire _w2811_ ;
	wire _w2810_ ;
	wire _w2809_ ;
	wire _w2808_ ;
	wire _w2807_ ;
	wire _w2806_ ;
	wire _w2805_ ;
	wire _w2804_ ;
	wire _w2803_ ;
	wire _w2802_ ;
	wire _w2801_ ;
	wire _w2800_ ;
	wire _w2799_ ;
	wire _w2798_ ;
	wire _w2797_ ;
	wire _w2796_ ;
	wire _w2795_ ;
	wire _w2794_ ;
	wire _w2793_ ;
	wire _w2792_ ;
	wire _w2791_ ;
	wire _w2790_ ;
	wire _w2789_ ;
	wire _w2788_ ;
	wire _w2787_ ;
	wire _w2786_ ;
	wire _w2785_ ;
	wire _w2784_ ;
	wire _w2783_ ;
	wire _w2782_ ;
	wire _w2781_ ;
	wire _w2780_ ;
	wire _w2779_ ;
	wire _w2778_ ;
	wire _w2777_ ;
	wire _w2776_ ;
	wire _w2775_ ;
	wire _w2774_ ;
	wire _w2773_ ;
	wire _w2772_ ;
	wire _w2771_ ;
	wire _w2770_ ;
	wire _w2769_ ;
	wire _w2768_ ;
	wire _w2767_ ;
	wire _w2766_ ;
	wire _w2765_ ;
	wire _w2764_ ;
	wire _w2763_ ;
	wire _w2762_ ;
	wire _w2761_ ;
	wire _w2760_ ;
	wire _w2759_ ;
	wire _w2758_ ;
	wire _w2757_ ;
	wire _w2756_ ;
	wire _w2755_ ;
	wire _w2754_ ;
	wire _w2753_ ;
	wire _w2752_ ;
	wire _w2751_ ;
	wire _w2750_ ;
	wire _w2749_ ;
	wire _w2748_ ;
	wire _w2747_ ;
	wire _w2746_ ;
	wire _w2745_ ;
	wire _w2744_ ;
	wire _w2743_ ;
	wire _w2742_ ;
	wire _w2741_ ;
	wire _w2740_ ;
	wire _w2739_ ;
	wire _w2738_ ;
	wire _w2737_ ;
	wire _w2736_ ;
	wire _w2735_ ;
	wire _w2734_ ;
	wire _w2733_ ;
	wire _w2732_ ;
	wire _w2731_ ;
	wire _w2730_ ;
	wire _w2729_ ;
	wire _w2728_ ;
	wire _w2727_ ;
	wire _w2726_ ;
	wire _w2725_ ;
	wire _w2724_ ;
	wire _w2723_ ;
	wire _w2722_ ;
	wire _w2721_ ;
	wire _w2720_ ;
	wire _w2719_ ;
	wire _w2718_ ;
	wire _w2717_ ;
	wire _w2716_ ;
	wire _w2715_ ;
	wire _w2714_ ;
	wire _w2713_ ;
	wire _w2712_ ;
	wire _w2711_ ;
	wire _w2710_ ;
	wire _w2709_ ;
	wire _w2708_ ;
	wire _w2707_ ;
	wire _w2706_ ;
	wire _w2705_ ;
	wire _w2704_ ;
	wire _w2703_ ;
	wire _w2702_ ;
	wire _w2701_ ;
	wire _w2700_ ;
	wire _w2699_ ;
	wire _w2698_ ;
	wire _w2697_ ;
	wire _w2696_ ;
	wire _w2695_ ;
	wire _w2694_ ;
	wire _w2693_ ;
	wire _w2692_ ;
	wire _w2691_ ;
	wire _w2690_ ;
	wire _w2689_ ;
	wire _w2688_ ;
	wire _w2687_ ;
	wire _w2686_ ;
	wire _w2685_ ;
	wire _w2684_ ;
	wire _w2683_ ;
	wire _w2682_ ;
	wire _w2681_ ;
	wire _w2680_ ;
	wire _w2679_ ;
	wire _w2678_ ;
	wire _w2677_ ;
	wire _w2676_ ;
	wire _w2675_ ;
	wire _w2674_ ;
	wire _w2673_ ;
	wire _w2672_ ;
	wire _w2671_ ;
	wire _w2670_ ;
	wire _w2669_ ;
	wire _w2668_ ;
	wire _w2667_ ;
	wire _w2666_ ;
	wire _w2665_ ;
	wire _w2664_ ;
	wire _w2663_ ;
	wire _w2662_ ;
	wire _w2661_ ;
	wire _w2660_ ;
	wire _w2659_ ;
	wire _w2658_ ;
	wire _w2657_ ;
	wire _w2656_ ;
	wire _w2655_ ;
	wire _w2654_ ;
	wire _w2653_ ;
	wire _w2652_ ;
	wire _w2651_ ;
	wire _w2650_ ;
	wire _w2649_ ;
	wire _w2648_ ;
	wire _w2647_ ;
	wire _w2646_ ;
	wire _w2645_ ;
	wire _w2644_ ;
	wire _w2643_ ;
	wire _w2642_ ;
	wire _w2641_ ;
	wire _w2640_ ;
	wire _w2639_ ;
	wire _w2638_ ;
	wire _w2637_ ;
	wire _w2636_ ;
	wire _w2635_ ;
	wire _w2634_ ;
	wire _w2633_ ;
	wire _w2632_ ;
	wire _w2631_ ;
	wire _w2630_ ;
	wire _w2629_ ;
	wire _w2628_ ;
	wire _w2627_ ;
	wire _w2626_ ;
	wire _w2625_ ;
	wire _w2624_ ;
	wire _w2623_ ;
	wire _w2622_ ;
	wire _w2621_ ;
	wire _w2620_ ;
	wire _w2619_ ;
	wire _w2618_ ;
	wire _w2617_ ;
	wire _w2616_ ;
	wire _w2615_ ;
	wire _w2614_ ;
	wire _w2613_ ;
	wire _w2612_ ;
	wire _w2611_ ;
	wire _w2610_ ;
	wire _w2609_ ;
	wire _w2608_ ;
	wire _w2607_ ;
	wire _w2606_ ;
	wire _w2605_ ;
	wire _w2604_ ;
	wire _w2603_ ;
	wire _w2602_ ;
	wire _w2601_ ;
	wire _w2600_ ;
	wire _w2599_ ;
	wire _w2598_ ;
	wire _w2597_ ;
	wire _w2596_ ;
	wire _w2595_ ;
	wire _w2594_ ;
	wire _w2593_ ;
	wire _w2592_ ;
	wire _w2591_ ;
	wire _w2590_ ;
	wire _w2589_ ;
	wire _w2588_ ;
	wire _w2587_ ;
	wire _w2586_ ;
	wire _w2585_ ;
	wire _w2584_ ;
	wire _w2583_ ;
	wire _w2582_ ;
	wire _w2581_ ;
	wire _w2580_ ;
	wire _w2579_ ;
	wire _w2578_ ;
	wire _w2577_ ;
	wire _w2576_ ;
	wire _w2575_ ;
	wire _w2574_ ;
	wire _w2572_ ;
	wire _w2571_ ;
	wire _w2570_ ;
	wire _w2569_ ;
	wire _w2568_ ;
	wire _w2567_ ;
	wire _w2566_ ;
	wire _w2565_ ;
	wire _w2564_ ;
	wire _w2563_ ;
	wire _w2562_ ;
	wire _w2561_ ;
	wire _w2560_ ;
	wire _w2559_ ;
	wire _w2558_ ;
	wire _w2557_ ;
	wire _w2556_ ;
	wire _w2555_ ;
	wire _w2554_ ;
	wire _w2553_ ;
	wire _w2552_ ;
	wire _w2551_ ;
	wire _w2550_ ;
	wire _w2549_ ;
	wire _w2548_ ;
	wire _w2547_ ;
	wire _w2546_ ;
	wire _w2545_ ;
	wire _w2544_ ;
	wire _w2543_ ;
	wire _w2542_ ;
	wire _w2541_ ;
	wire _w2540_ ;
	wire _w2539_ ;
	wire _w2538_ ;
	wire _w2537_ ;
	wire _w2536_ ;
	wire _w2535_ ;
	wire _w2534_ ;
	wire _w2533_ ;
	wire _w2532_ ;
	wire _w2531_ ;
	wire _w2530_ ;
	wire _w2529_ ;
	wire _w2528_ ;
	wire _w2527_ ;
	wire _w2526_ ;
	wire _w2525_ ;
	wire _w2524_ ;
	wire _w2523_ ;
	wire _w2522_ ;
	wire _w2521_ ;
	wire _w2520_ ;
	wire _w2519_ ;
	wire _w2518_ ;
	wire _w2517_ ;
	wire _w2516_ ;
	wire _w2515_ ;
	wire _w2514_ ;
	wire _w2513_ ;
	wire _w2512_ ;
	wire _w2511_ ;
	wire _w2510_ ;
	wire _w2509_ ;
	wire _w2508_ ;
	wire _w2507_ ;
	wire _w2506_ ;
	wire _w2505_ ;
	wire _w2504_ ;
	wire _w2503_ ;
	wire _w2502_ ;
	wire _w2501_ ;
	wire _w2500_ ;
	wire _w2499_ ;
	wire _w2498_ ;
	wire _w2497_ ;
	wire _w2496_ ;
	wire _w2495_ ;
	wire _w2494_ ;
	wire _w2493_ ;
	wire _w2492_ ;
	wire _w2491_ ;
	wire _w2490_ ;
	wire _w2489_ ;
	wire _w2488_ ;
	wire _w2487_ ;
	wire _w2486_ ;
	wire _w2485_ ;
	wire _w2484_ ;
	wire _w2483_ ;
	wire _w2482_ ;
	wire _w2481_ ;
	wire _w2480_ ;
	wire _w2479_ ;
	wire _w2478_ ;
	wire _w2477_ ;
	wire _w2476_ ;
	wire _w2475_ ;
	wire _w2474_ ;
	wire _w2473_ ;
	wire _w2472_ ;
	wire _w2471_ ;
	wire _w2470_ ;
	wire _w2469_ ;
	wire _w2468_ ;
	wire _w2467_ ;
	wire _w2466_ ;
	wire _w2465_ ;
	wire _w2464_ ;
	wire _w2463_ ;
	wire _w2462_ ;
	wire _w2461_ ;
	wire _w2460_ ;
	wire _w2459_ ;
	wire _w2458_ ;
	wire _w2457_ ;
	wire _w2456_ ;
	wire _w2455_ ;
	wire _w2454_ ;
	wire _w2453_ ;
	wire _w2452_ ;
	wire _w2451_ ;
	wire _w2450_ ;
	wire _w2449_ ;
	wire _w2448_ ;
	wire _w2447_ ;
	wire _w2446_ ;
	wire _w2445_ ;
	wire _w2444_ ;
	wire _w2443_ ;
	wire _w2442_ ;
	wire _w2441_ ;
	wire _w2440_ ;
	wire _w2439_ ;
	wire _w2438_ ;
	wire _w2437_ ;
	wire _w2436_ ;
	wire _w2435_ ;
	wire _w2434_ ;
	wire _w2433_ ;
	wire _w2432_ ;
	wire _w2431_ ;
	wire _w2430_ ;
	wire _w2429_ ;
	wire _w2428_ ;
	wire _w2427_ ;
	wire _w2426_ ;
	wire _w2425_ ;
	wire _w2424_ ;
	wire _w2423_ ;
	wire _w2422_ ;
	wire _w2421_ ;
	wire _w2420_ ;
	wire _w2419_ ;
	wire _w2418_ ;
	wire _w2417_ ;
	wire _w2416_ ;
	wire _w2415_ ;
	wire _w2414_ ;
	wire _w2413_ ;
	wire _w2412_ ;
	wire _w2411_ ;
	wire _w2410_ ;
	wire _w2409_ ;
	wire _w2408_ ;
	wire _w2407_ ;
	wire _w2406_ ;
	wire _w2405_ ;
	wire _w2404_ ;
	wire _w2403_ ;
	wire _w2402_ ;
	wire _w2401_ ;
	wire _w2400_ ;
	wire _w2399_ ;
	wire _w2398_ ;
	wire _w2397_ ;
	wire _w2396_ ;
	wire _w2395_ ;
	wire _w2394_ ;
	wire _w2393_ ;
	wire _w2392_ ;
	wire _w2391_ ;
	wire _w2390_ ;
	wire _w2389_ ;
	wire _w2388_ ;
	wire _w2387_ ;
	wire _w2386_ ;
	wire _w2385_ ;
	wire _w2384_ ;
	wire _w2383_ ;
	wire _w2382_ ;
	wire _w2381_ ;
	wire _w2380_ ;
	wire _w2379_ ;
	wire _w2378_ ;
	wire _w2377_ ;
	wire _w2376_ ;
	wire _w2375_ ;
	wire _w2374_ ;
	wire _w2373_ ;
	wire _w2372_ ;
	wire _w2371_ ;
	wire _w2370_ ;
	wire _w2369_ ;
	wire _w2368_ ;
	wire _w2367_ ;
	wire _w2366_ ;
	wire _w2365_ ;
	wire _w2364_ ;
	wire _w2363_ ;
	wire _w2362_ ;
	wire _w2361_ ;
	wire _w2360_ ;
	wire _w2359_ ;
	wire _w2358_ ;
	wire _w2357_ ;
	wire _w2356_ ;
	wire _w2355_ ;
	wire _w2354_ ;
	wire _w2353_ ;
	wire _w2352_ ;
	wire _w2351_ ;
	wire _w2350_ ;
	wire _w2349_ ;
	wire _w2348_ ;
	wire _w2347_ ;
	wire _w2346_ ;
	wire _w2345_ ;
	wire _w2344_ ;
	wire _w2343_ ;
	wire _w2342_ ;
	wire _w2341_ ;
	wire _w2340_ ;
	wire _w2339_ ;
	wire _w2338_ ;
	wire _w2337_ ;
	wire _w2336_ ;
	wire _w2335_ ;
	wire _w2334_ ;
	wire _w2333_ ;
	wire _w2332_ ;
	wire _w2331_ ;
	wire _w2330_ ;
	wire _w2329_ ;
	wire _w2328_ ;
	wire _w2327_ ;
	wire _w2326_ ;
	wire _w2325_ ;
	wire _w2324_ ;
	wire _w2323_ ;
	wire _w2322_ ;
	wire _w2321_ ;
	wire _w2320_ ;
	wire _w2319_ ;
	wire _w2318_ ;
	wire _w2317_ ;
	wire _w2316_ ;
	wire _w2315_ ;
	wire _w2314_ ;
	wire _w2313_ ;
	wire _w2312_ ;
	wire _w2311_ ;
	wire _w2310_ ;
	wire _w2309_ ;
	wire _w2308_ ;
	wire _w2307_ ;
	wire _w2306_ ;
	wire _w2305_ ;
	wire _w2304_ ;
	wire _w2303_ ;
	wire _w2302_ ;
	wire _w2301_ ;
	wire _w2300_ ;
	wire _w2299_ ;
	wire _w2298_ ;
	wire _w2297_ ;
	wire _w2296_ ;
	wire _w2295_ ;
	wire _w2294_ ;
	wire _w2293_ ;
	wire _w2292_ ;
	wire _w2291_ ;
	wire _w2290_ ;
	wire _w2289_ ;
	wire _w2288_ ;
	wire _w2287_ ;
	wire _w2286_ ;
	wire _w2285_ ;
	wire _w2284_ ;
	wire _w2283_ ;
	wire _w2282_ ;
	wire _w2281_ ;
	wire _w2280_ ;
	wire _w2279_ ;
	wire _w2278_ ;
	wire _w2277_ ;
	wire _w2276_ ;
	wire _w2275_ ;
	wire _w2274_ ;
	wire _w2273_ ;
	wire _w2272_ ;
	wire _w2271_ ;
	wire _w2270_ ;
	wire _w2269_ ;
	wire _w2268_ ;
	wire _w2267_ ;
	wire _w2266_ ;
	wire _w2265_ ;
	wire _w2264_ ;
	wire _w2263_ ;
	wire _w2262_ ;
	wire _w2261_ ;
	wire _w2260_ ;
	wire _w2259_ ;
	wire _w2258_ ;
	wire _w2257_ ;
	wire _w2256_ ;
	wire _w2255_ ;
	wire _w2254_ ;
	wire _w2253_ ;
	wire _w2252_ ;
	wire _w2251_ ;
	wire _w2250_ ;
	wire _w2249_ ;
	wire _w2248_ ;
	wire _w2247_ ;
	wire _w2246_ ;
	wire _w2245_ ;
	wire _w2244_ ;
	wire _w2243_ ;
	wire _w2242_ ;
	wire _w2241_ ;
	wire _w2240_ ;
	wire _w2239_ ;
	wire _w2238_ ;
	wire _w2237_ ;
	wire _w2236_ ;
	wire _w2235_ ;
	wire _w2234_ ;
	wire _w2233_ ;
	wire _w2232_ ;
	wire _w2231_ ;
	wire _w2230_ ;
	wire _w2229_ ;
	wire _w2228_ ;
	wire _w2227_ ;
	wire _w2226_ ;
	wire _w2225_ ;
	wire _w2224_ ;
	wire _w2223_ ;
	wire _w2222_ ;
	wire _w2221_ ;
	wire _w2220_ ;
	wire _w2219_ ;
	wire _w2218_ ;
	wire _w2217_ ;
	wire _w2216_ ;
	wire _w2215_ ;
	wire _w2214_ ;
	wire _w2213_ ;
	wire _w2212_ ;
	wire _w2211_ ;
	wire _w2210_ ;
	wire _w2209_ ;
	wire _w2208_ ;
	wire _w2207_ ;
	wire _w2206_ ;
	wire _w2205_ ;
	wire _w2204_ ;
	wire _w2203_ ;
	wire _w2202_ ;
	wire _w2201_ ;
	wire _w2200_ ;
	wire _w2199_ ;
	wire _w2198_ ;
	wire _w2197_ ;
	wire _w2196_ ;
	wire _w2195_ ;
	wire _w2194_ ;
	wire _w2193_ ;
	wire _w2192_ ;
	wire _w2191_ ;
	wire _w2190_ ;
	wire _w2189_ ;
	wire _w2188_ ;
	wire _w2187_ ;
	wire _w2186_ ;
	wire _w2185_ ;
	wire _w2184_ ;
	wire _w2183_ ;
	wire _w2182_ ;
	wire _w2181_ ;
	wire _w2180_ ;
	wire _w2179_ ;
	wire _w2178_ ;
	wire _w2177_ ;
	wire _w2176_ ;
	wire _w2175_ ;
	wire _w2174_ ;
	wire _w2173_ ;
	wire _w2172_ ;
	wire _w2171_ ;
	wire _w2170_ ;
	wire _w2169_ ;
	wire _w2168_ ;
	wire _w2167_ ;
	wire _w2166_ ;
	wire _w2165_ ;
	wire _w2164_ ;
	wire _w2163_ ;
	wire _w2162_ ;
	wire _w2161_ ;
	wire _w2160_ ;
	wire _w2159_ ;
	wire _w2158_ ;
	wire _w2157_ ;
	wire _w2156_ ;
	wire _w2155_ ;
	wire _w2154_ ;
	wire _w2153_ ;
	wire _w2152_ ;
	wire _w2151_ ;
	wire _w2150_ ;
	wire _w2149_ ;
	wire _w2148_ ;
	wire _w2147_ ;
	wire _w2146_ ;
	wire _w2145_ ;
	wire _w2144_ ;
	wire _w2143_ ;
	wire _w2142_ ;
	wire _w2141_ ;
	wire _w2140_ ;
	wire _w2139_ ;
	wire _w2138_ ;
	wire _w2137_ ;
	wire _w2136_ ;
	wire _w2135_ ;
	wire _w2134_ ;
	wire _w2133_ ;
	wire _w2132_ ;
	wire _w2131_ ;
	wire _w2130_ ;
	wire _w2129_ ;
	wire _w2128_ ;
	wire _w2127_ ;
	wire _w2126_ ;
	wire _w2125_ ;
	wire _w2124_ ;
	wire _w2123_ ;
	wire _w2122_ ;
	wire _w2121_ ;
	wire _w2120_ ;
	wire _w2119_ ;
	wire _w2118_ ;
	wire _w2117_ ;
	wire _w2116_ ;
	wire _w2115_ ;
	wire _w2114_ ;
	wire _w2113_ ;
	wire _w2112_ ;
	wire _w2111_ ;
	wire _w2110_ ;
	wire _w2109_ ;
	wire _w2108_ ;
	wire _w2107_ ;
	wire _w2106_ ;
	wire _w2105_ ;
	wire _w2104_ ;
	wire _w2103_ ;
	wire _w2102_ ;
	wire _w2101_ ;
	wire _w2100_ ;
	wire _w2099_ ;
	wire _w2098_ ;
	wire _w2097_ ;
	wire _w2096_ ;
	wire _w2095_ ;
	wire _w2094_ ;
	wire _w2093_ ;
	wire _w2092_ ;
	wire _w2091_ ;
	wire _w2090_ ;
	wire _w2089_ ;
	wire _w2088_ ;
	wire _w2087_ ;
	wire _w2086_ ;
	wire _w2085_ ;
	wire _w2084_ ;
	wire _w2083_ ;
	wire _w2082_ ;
	wire _w2081_ ;
	wire _w2080_ ;
	wire _w2079_ ;
	wire _w2078_ ;
	wire _w2077_ ;
	wire _w2076_ ;
	wire _w2075_ ;
	wire _w2074_ ;
	wire _w2073_ ;
	wire _w2072_ ;
	wire _w2071_ ;
	wire _w2070_ ;
	wire _w2069_ ;
	wire _w2068_ ;
	wire _w2067_ ;
	wire _w2066_ ;
	wire _w2065_ ;
	wire _w2064_ ;
	wire _w2063_ ;
	wire _w2062_ ;
	wire _w2061_ ;
	wire _w2060_ ;
	wire _w2059_ ;
	wire _w2058_ ;
	wire _w2057_ ;
	wire _w2056_ ;
	wire _w2055_ ;
	wire _w2054_ ;
	wire _w2053_ ;
	wire _w2052_ ;
	wire _w2051_ ;
	wire _w2050_ ;
	wire _w2049_ ;
	wire _w2048_ ;
	wire _w2047_ ;
	wire _w2046_ ;
	wire _w2045_ ;
	wire _w2044_ ;
	wire _w2043_ ;
	wire _w2042_ ;
	wire _w2041_ ;
	wire _w2040_ ;
	wire _w2039_ ;
	wire _w2038_ ;
	wire _w2037_ ;
	wire _w2036_ ;
	wire _w2035_ ;
	wire _w2034_ ;
	wire _w2033_ ;
	wire _w2032_ ;
	wire _w2031_ ;
	wire _w2030_ ;
	wire _w2029_ ;
	wire _w2028_ ;
	wire _w2027_ ;
	wire _w2026_ ;
	wire _w2025_ ;
	wire _w2024_ ;
	wire _w2023_ ;
	wire _w2022_ ;
	wire _w2021_ ;
	wire _w2020_ ;
	wire _w2019_ ;
	wire _w2018_ ;
	wire _w2017_ ;
	wire _w2016_ ;
	wire _w2015_ ;
	wire _w2014_ ;
	wire _w2013_ ;
	wire _w2012_ ;
	wire _w2011_ ;
	wire _w2010_ ;
	wire _w2009_ ;
	wire _w2008_ ;
	wire _w2007_ ;
	wire _w2006_ ;
	wire _w2005_ ;
	wire _w2004_ ;
	wire _w2003_ ;
	wire _w2002_ ;
	wire _w2001_ ;
	wire _w2000_ ;
	wire _w1999_ ;
	wire _w1998_ ;
	wire _w1997_ ;
	wire _w1996_ ;
	wire _w1995_ ;
	wire _w1994_ ;
	wire _w1993_ ;
	wire _w1992_ ;
	wire _w1991_ ;
	wire _w1990_ ;
	wire _w1989_ ;
	wire _w1988_ ;
	wire _w1987_ ;
	wire _w1986_ ;
	wire _w1985_ ;
	wire _w1984_ ;
	wire _w1983_ ;
	wire _w1982_ ;
	wire _w1981_ ;
	wire _w1980_ ;
	wire _w1979_ ;
	wire _w1978_ ;
	wire _w1977_ ;
	wire _w1976_ ;
	wire _w1975_ ;
	wire _w1974_ ;
	wire _w1973_ ;
	wire _w1972_ ;
	wire _w1971_ ;
	wire _w1970_ ;
	wire _w1969_ ;
	wire _w1968_ ;
	wire _w1967_ ;
	wire _w1966_ ;
	wire _w1965_ ;
	wire _w1964_ ;
	wire _w1963_ ;
	wire _w1962_ ;
	wire _w1961_ ;
	wire _w1960_ ;
	wire _w1959_ ;
	wire _w1958_ ;
	wire _w1957_ ;
	wire _w1956_ ;
	wire _w1955_ ;
	wire _w1954_ ;
	wire _w1953_ ;
	wire _w1952_ ;
	wire _w1951_ ;
	wire _w1950_ ;
	wire _w1949_ ;
	wire _w1948_ ;
	wire _w1947_ ;
	wire _w1946_ ;
	wire _w1945_ ;
	wire _w1944_ ;
	wire _w1943_ ;
	wire _w1942_ ;
	wire _w1941_ ;
	wire _w1940_ ;
	wire _w1939_ ;
	wire _w1938_ ;
	wire _w1937_ ;
	wire _w1936_ ;
	wire _w1935_ ;
	wire _w1934_ ;
	wire _w1933_ ;
	wire _w1932_ ;
	wire _w1931_ ;
	wire _w1930_ ;
	wire _w1929_ ;
	wire _w1928_ ;
	wire _w1927_ ;
	wire _w1926_ ;
	wire _w1925_ ;
	wire _w1924_ ;
	wire _w1923_ ;
	wire _w1922_ ;
	wire _w1921_ ;
	wire _w1920_ ;
	wire _w1919_ ;
	wire _w1918_ ;
	wire _w1917_ ;
	wire _w1916_ ;
	wire _w1915_ ;
	wire _w1914_ ;
	wire _w1913_ ;
	wire _w1912_ ;
	wire _w1911_ ;
	wire _w1910_ ;
	wire _w1909_ ;
	wire _w1908_ ;
	wire _w1907_ ;
	wire _w1906_ ;
	wire _w1905_ ;
	wire _w1904_ ;
	wire _w1903_ ;
	wire _w1902_ ;
	wire _w1901_ ;
	wire _w1900_ ;
	wire _w1899_ ;
	wire _w1898_ ;
	wire _w1897_ ;
	wire _w1896_ ;
	wire _w1895_ ;
	wire _w1894_ ;
	wire _w1893_ ;
	wire _w1892_ ;
	wire _w1891_ ;
	wire _w1890_ ;
	wire _w1889_ ;
	wire _w1888_ ;
	wire _w1887_ ;
	wire _w1886_ ;
	wire _w1885_ ;
	wire _w1884_ ;
	wire _w1883_ ;
	wire _w1882_ ;
	wire _w1881_ ;
	wire _w1880_ ;
	wire _w1879_ ;
	wire _w1878_ ;
	wire _w1877_ ;
	wire _w1876_ ;
	wire _w1875_ ;
	wire _w1874_ ;
	wire _w1873_ ;
	wire _w1872_ ;
	wire _w1871_ ;
	wire _w1870_ ;
	wire _w1869_ ;
	wire _w1868_ ;
	wire _w1867_ ;
	wire _w1866_ ;
	wire _w1865_ ;
	wire _w1864_ ;
	wire _w1863_ ;
	wire _w1862_ ;
	wire _w1861_ ;
	wire _w1860_ ;
	wire _w1859_ ;
	wire _w1858_ ;
	wire _w1857_ ;
	wire _w1856_ ;
	wire _w1855_ ;
	wire _w1854_ ;
	wire _w1853_ ;
	wire _w1852_ ;
	wire _w1851_ ;
	wire _w1850_ ;
	wire _w1849_ ;
	wire _w1848_ ;
	wire _w1847_ ;
	wire _w1846_ ;
	wire _w1845_ ;
	wire _w1844_ ;
	wire _w1843_ ;
	wire _w1842_ ;
	wire _w1841_ ;
	wire _w1840_ ;
	wire _w1839_ ;
	wire _w1838_ ;
	wire _w1837_ ;
	wire _w1836_ ;
	wire _w1835_ ;
	wire _w1834_ ;
	wire _w1833_ ;
	wire _w1832_ ;
	wire _w1831_ ;
	wire _w1830_ ;
	wire _w1829_ ;
	wire _w1828_ ;
	wire _w1827_ ;
	wire _w1826_ ;
	wire _w1825_ ;
	wire _w1824_ ;
	wire _w1823_ ;
	wire _w1822_ ;
	wire _w1821_ ;
	wire _w1820_ ;
	wire _w1819_ ;
	wire _w1818_ ;
	wire _w1817_ ;
	wire _w1816_ ;
	wire _w1815_ ;
	wire _w1814_ ;
	wire _w1813_ ;
	wire _w1812_ ;
	wire _w1811_ ;
	wire _w1810_ ;
	wire _w1809_ ;
	wire _w1808_ ;
	wire _w1807_ ;
	wire _w1806_ ;
	wire _w1805_ ;
	wire _w1804_ ;
	wire _w1803_ ;
	wire _w1802_ ;
	wire _w1801_ ;
	wire _w1800_ ;
	wire _w1799_ ;
	wire _w1798_ ;
	wire _w1797_ ;
	wire _w1796_ ;
	wire _w1795_ ;
	wire _w1794_ ;
	wire _w1793_ ;
	wire _w1792_ ;
	wire _w1791_ ;
	wire _w1790_ ;
	wire _w1789_ ;
	wire _w1788_ ;
	wire _w1787_ ;
	wire _w1786_ ;
	wire _w1785_ ;
	wire _w1784_ ;
	wire _w1783_ ;
	wire _w1782_ ;
	wire _w1781_ ;
	wire _w1780_ ;
	wire _w1779_ ;
	wire _w1778_ ;
	wire _w1777_ ;
	wire _w1776_ ;
	wire _w1775_ ;
	wire _w1774_ ;
	wire _w1773_ ;
	wire _w1772_ ;
	wire _w1771_ ;
	wire _w1770_ ;
	wire _w1769_ ;
	wire _w1768_ ;
	wire _w1767_ ;
	wire _w1766_ ;
	wire _w1765_ ;
	wire _w1764_ ;
	wire _w1763_ ;
	wire _w1762_ ;
	wire _w1761_ ;
	wire _w1760_ ;
	wire _w1759_ ;
	wire _w1758_ ;
	wire _w1757_ ;
	wire _w1756_ ;
	wire _w1755_ ;
	wire _w1754_ ;
	wire _w1753_ ;
	wire _w1752_ ;
	wire _w1751_ ;
	wire _w1750_ ;
	wire _w1749_ ;
	wire _w1748_ ;
	wire _w1747_ ;
	wire _w1746_ ;
	wire _w1745_ ;
	wire _w1744_ ;
	wire _w1743_ ;
	wire _w1742_ ;
	wire _w1741_ ;
	wire _w1740_ ;
	wire _w1739_ ;
	wire _w1738_ ;
	wire _w1737_ ;
	wire _w1736_ ;
	wire _w1735_ ;
	wire _w1734_ ;
	wire _w1733_ ;
	wire _w1732_ ;
	wire _w1731_ ;
	wire _w1730_ ;
	wire _w1729_ ;
	wire _w1728_ ;
	wire _w1727_ ;
	wire _w1726_ ;
	wire _w1725_ ;
	wire _w1724_ ;
	wire _w1723_ ;
	wire _w1722_ ;
	wire _w1721_ ;
	wire _w1720_ ;
	wire _w1719_ ;
	wire _w1718_ ;
	wire _w1717_ ;
	wire _w1716_ ;
	wire _w1715_ ;
	wire _w1714_ ;
	wire _w1713_ ;
	wire _w1712_ ;
	wire _w1711_ ;
	wire _w1710_ ;
	wire _w1709_ ;
	wire _w1708_ ;
	wire _w1707_ ;
	wire _w1706_ ;
	wire _w1705_ ;
	wire _w1704_ ;
	wire _w1703_ ;
	wire _w1702_ ;
	wire _w1701_ ;
	wire _w1700_ ;
	wire _w1699_ ;
	wire _w1698_ ;
	wire _w1697_ ;
	wire _w1696_ ;
	wire _w1695_ ;
	wire _w1694_ ;
	wire _w1693_ ;
	wire _w1692_ ;
	wire _w1691_ ;
	wire _w1690_ ;
	wire _w1689_ ;
	wire _w1688_ ;
	wire _w1687_ ;
	wire _w1686_ ;
	wire _w1685_ ;
	wire _w1684_ ;
	wire _w1683_ ;
	wire _w1682_ ;
	wire _w1681_ ;
	wire _w1680_ ;
	wire _w1679_ ;
	wire _w1678_ ;
	wire _w1677_ ;
	wire _w1676_ ;
	wire _w1675_ ;
	wire _w1674_ ;
	wire _w1673_ ;
	wire _w1672_ ;
	wire _w1671_ ;
	wire _w1670_ ;
	wire _w1669_ ;
	wire _w1668_ ;
	wire _w1667_ ;
	wire _w1666_ ;
	wire _w1665_ ;
	wire _w1664_ ;
	wire _w1663_ ;
	wire _w1662_ ;
	wire _w1661_ ;
	wire _w1660_ ;
	wire _w1659_ ;
	wire _w1658_ ;
	wire _w1657_ ;
	wire _w1656_ ;
	wire _w1655_ ;
	wire _w1654_ ;
	wire _w1653_ ;
	wire _w1652_ ;
	wire _w1651_ ;
	wire _w1650_ ;
	wire _w1649_ ;
	wire _w1648_ ;
	wire _w1647_ ;
	wire _w1646_ ;
	wire _w1645_ ;
	wire _w1644_ ;
	wire _w1643_ ;
	wire _w1642_ ;
	wire _w1641_ ;
	wire _w1640_ ;
	wire _w1639_ ;
	wire _w1638_ ;
	wire _w1637_ ;
	wire _w1636_ ;
	wire _w1635_ ;
	wire _w1634_ ;
	wire _w1633_ ;
	wire _w1632_ ;
	wire _w1631_ ;
	wire _w1630_ ;
	wire _w1629_ ;
	wire _w1628_ ;
	wire _w1627_ ;
	wire _w1626_ ;
	wire _w1625_ ;
	wire _w1624_ ;
	wire _w1623_ ;
	wire _w1622_ ;
	wire _w1621_ ;
	wire _w1620_ ;
	wire _w1619_ ;
	wire _w1618_ ;
	wire _w1617_ ;
	wire _w1616_ ;
	wire _w1615_ ;
	wire _w1614_ ;
	wire _w1613_ ;
	wire _w1612_ ;
	wire _w1611_ ;
	wire _w1610_ ;
	wire _w1609_ ;
	wire _w1608_ ;
	wire _w1607_ ;
	wire _w1606_ ;
	wire _w1605_ ;
	wire _w1604_ ;
	wire _w1603_ ;
	wire _w1602_ ;
	wire _w1601_ ;
	wire _w1600_ ;
	wire _w1599_ ;
	wire _w1598_ ;
	wire _w1597_ ;
	wire _w1596_ ;
	wire _w1595_ ;
	wire _w1594_ ;
	wire _w1593_ ;
	wire _w1592_ ;
	wire _w1591_ ;
	wire _w1590_ ;
	wire _w1589_ ;
	wire _w1588_ ;
	wire _w1587_ ;
	wire _w1586_ ;
	wire _w1585_ ;
	wire _w1584_ ;
	wire _w1583_ ;
	wire _w1582_ ;
	wire _w1581_ ;
	wire _w1580_ ;
	wire _w1579_ ;
	wire _w1578_ ;
	wire _w1577_ ;
	wire _w1576_ ;
	wire _w1575_ ;
	wire _w1574_ ;
	wire _w1573_ ;
	wire _w1572_ ;
	wire _w1003_ ;
	wire _w1002_ ;
	wire _w1001_ ;
	wire _w1000_ ;
	wire _w999_ ;
	wire _w998_ ;
	wire _w997_ ;
	wire _w996_ ;
	wire _w995_ ;
	wire _w994_ ;
	wire _w993_ ;
	wire _w992_ ;
	wire _w991_ ;
	wire _w990_ ;
	wire _w989_ ;
	wire _w988_ ;
	wire _w987_ ;
	wire _w986_ ;
	wire _w985_ ;
	wire _w984_ ;
	wire _w983_ ;
	wire _w982_ ;
	wire _w981_ ;
	wire _w980_ ;
	wire _w979_ ;
	wire _w978_ ;
	wire _w977_ ;
	wire _w976_ ;
	wire _w975_ ;
	wire _w974_ ;
	wire _w973_ ;
	wire _w972_ ;
	wire _w971_ ;
	wire _w970_ ;
	wire _w969_ ;
	wire _w968_ ;
	wire _w967_ ;
	wire _w966_ ;
	wire _w965_ ;
	wire _w964_ ;
	wire _w963_ ;
	wire _w962_ ;
	wire _w961_ ;
	wire _w960_ ;
	wire _w959_ ;
	wire _w958_ ;
	wire _w957_ ;
	wire _w956_ ;
	wire _w955_ ;
	wire _w954_ ;
	wire _w953_ ;
	wire _w952_ ;
	wire _w951_ ;
	wire _w950_ ;
	wire _w949_ ;
	wire _w948_ ;
	wire _w947_ ;
	wire _w946_ ;
	wire _w945_ ;
	wire _w944_ ;
	wire _w943_ ;
	wire _w942_ ;
	wire _w941_ ;
	wire _w940_ ;
	wire _w939_ ;
	wire _w938_ ;
	wire _w937_ ;
	wire _w936_ ;
	wire _w935_ ;
	wire _w934_ ;
	wire _w933_ ;
	wire _w932_ ;
	wire _w931_ ;
	wire _w930_ ;
	wire _w929_ ;
	wire _w928_ ;
	wire _w927_ ;
	wire _w926_ ;
	wire _w925_ ;
	wire _w924_ ;
	wire _w923_ ;
	wire _w922_ ;
	wire _w921_ ;
	wire _w920_ ;
	wire _w919_ ;
	wire _w918_ ;
	wire _w917_ ;
	wire _w916_ ;
	wire _w915_ ;
	wire _w914_ ;
	wire _w913_ ;
	wire _w912_ ;
	wire _w911_ ;
	wire _w910_ ;
	wire _w909_ ;
	wire _w908_ ;
	wire _w907_ ;
	wire _w906_ ;
	wire _w905_ ;
	wire _w904_ ;
	wire _w903_ ;
	wire _w902_ ;
	wire _w901_ ;
	wire _w900_ ;
	wire _w899_ ;
	wire _w898_ ;
	wire _w897_ ;
	wire _w896_ ;
	wire _w895_ ;
	wire _w894_ ;
	wire _w893_ ;
	wire _w892_ ;
	wire _w891_ ;
	wire _w890_ ;
	wire _w889_ ;
	wire _w888_ ;
	wire _w887_ ;
	wire _w886_ ;
	wire _w885_ ;
	wire _w884_ ;
	wire _w883_ ;
	wire _w882_ ;
	wire _w881_ ;
	wire _w880_ ;
	wire _w879_ ;
	wire _w878_ ;
	wire _w877_ ;
	wire _w876_ ;
	wire _w875_ ;
	wire _w874_ ;
	wire _w873_ ;
	wire _w872_ ;
	wire _w871_ ;
	wire _w870_ ;
	wire _w869_ ;
	wire _w868_ ;
	wire _w867_ ;
	wire _w866_ ;
	wire _w865_ ;
	wire _w864_ ;
	wire _w863_ ;
	wire _w862_ ;
	wire _w861_ ;
	wire _w860_ ;
	wire _w859_ ;
	wire _w858_ ;
	wire _w857_ ;
	wire _w856_ ;
	wire _w855_ ;
	wire _w854_ ;
	wire _w853_ ;
	wire _w852_ ;
	wire _w851_ ;
	wire _w850_ ;
	wire _w849_ ;
	wire _w848_ ;
	wire _w847_ ;
	wire _w846_ ;
	wire _w845_ ;
	wire _w844_ ;
	wire _w843_ ;
	wire _w842_ ;
	wire _w841_ ;
	wire _w840_ ;
	wire _w839_ ;
	wire _w838_ ;
	wire _w837_ ;
	wire _w836_ ;
	wire _w835_ ;
	wire _w834_ ;
	wire _w833_ ;
	wire _w832_ ;
	wire _w831_ ;
	wire _w830_ ;
	wire _w829_ ;
	wire _w828_ ;
	wire _w827_ ;
	wire _w826_ ;
	wire _w825_ ;
	wire _w824_ ;
	wire _w823_ ;
	wire _w822_ ;
	wire _w821_ ;
	wire _w820_ ;
	wire _w819_ ;
	wire _w818_ ;
	wire _w817_ ;
	wire _w816_ ;
	wire _w815_ ;
	wire _w814_ ;
	wire _w813_ ;
	wire _w812_ ;
	wire _w811_ ;
	wire _w810_ ;
	wire _w809_ ;
	wire _w808_ ;
	wire _w807_ ;
	wire _w806_ ;
	wire _w805_ ;
	wire _w804_ ;
	wire _w803_ ;
	wire _w802_ ;
	wire _w801_ ;
	wire _w800_ ;
	wire _w799_ ;
	wire _w798_ ;
	wire _w797_ ;
	wire _w796_ ;
	wire _w795_ ;
	wire _w794_ ;
	wire _w793_ ;
	wire _w792_ ;
	wire _w791_ ;
	wire _w790_ ;
	wire _w789_ ;
	wire _w788_ ;
	wire _w787_ ;
	wire _w786_ ;
	wire _w785_ ;
	wire _w784_ ;
	wire _w783_ ;
	wire _w782_ ;
	wire _w781_ ;
	wire _w780_ ;
	wire _w779_ ;
	wire _w778_ ;
	wire _w777_ ;
	wire _w776_ ;
	wire _w775_ ;
	wire _w774_ ;
	wire _w773_ ;
	wire _w772_ ;
	wire _w771_ ;
	wire _w770_ ;
	wire _w769_ ;
	wire _w768_ ;
	wire _w767_ ;
	wire _w766_ ;
	wire _w765_ ;
	wire _w764_ ;
	wire _w763_ ;
	wire _w762_ ;
	wire _w761_ ;
	wire _w760_ ;
	wire _w759_ ;
	wire _w758_ ;
	wire _w756_ ;
	wire _w755_ ;
	wire _w754_ ;
	wire _w753_ ;
	wire _w752_ ;
	wire _w751_ ;
	wire _w750_ ;
	wire _w749_ ;
	wire _w748_ ;
	wire _w747_ ;
	wire _w746_ ;
	wire _w745_ ;
	wire _w744_ ;
	wire _w743_ ;
	wire _w742_ ;
	wire _w741_ ;
	wire _w740_ ;
	wire _w739_ ;
	wire _w738_ ;
	wire _w737_ ;
	wire _w736_ ;
	wire _w735_ ;
	wire _w734_ ;
	wire _w733_ ;
	wire _w732_ ;
	wire _w731_ ;
	wire _w730_ ;
	wire _w729_ ;
	wire _w728_ ;
	wire _w727_ ;
	wire _w726_ ;
	wire _w725_ ;
	wire _w724_ ;
	wire _w723_ ;
	wire _w722_ ;
	wire _w721_ ;
	wire _w720_ ;
	wire _w589_ ;
	wire _w588_ ;
	wire _w587_ ;
	wire _w586_ ;
	wire _w585_ ;
	wire _w584_ ;
	wire _w583_ ;
	wire _w582_ ;
	wire _w581_ ;
	wire _w580_ ;
	wire _w579_ ;
	wire _w578_ ;
	wire _w577_ ;
	wire _w576_ ;
	wire _w575_ ;
	wire _w574_ ;
	wire _w573_ ;
	wire _w572_ ;
	wire _w571_ ;
	wire _w570_ ;
	wire _w569_ ;
	wire _w568_ ;
	wire _w567_ ;
	wire _w566_ ;
	wire _w565_ ;
	wire _w564_ ;
	wire _w563_ ;
	wire _w562_ ;
	wire _w561_ ;
	wire _w560_ ;
	wire _w559_ ;
	wire _w558_ ;
	wire _w557_ ;
	wire _w556_ ;
	wire _w555_ ;
	wire _w554_ ;
	wire _w553_ ;
	wire _w552_ ;
	wire _w551_ ;
	wire _w550_ ;
	wire _w549_ ;
	wire _w548_ ;
	wire _w547_ ;
	wire _w546_ ;
	wire _w545_ ;
	wire _w544_ ;
	wire _w543_ ;
	wire _w542_ ;
	wire _w541_ ;
	wire _w540_ ;
	wire _w539_ ;
	wire _w538_ ;
	wire _w537_ ;
	wire _w536_ ;
	wire _w535_ ;
	wire _w534_ ;
	wire _w533_ ;
	wire _w532_ ;
	wire _w531_ ;
	wire _w530_ ;
	wire _w529_ ;
	wire _w528_ ;
	wire _w527_ ;
	wire _w526_ ;
	wire _w525_ ;
	wire _w524_ ;
	wire _w523_ ;
	wire _w522_ ;
	wire _w491_ ;
	wire _w490_ ;
	wire _w489_ ;
	wire _w488_ ;
	wire _w487_ ;
	wire _w486_ ;
	wire _w485_ ;
	wire _w484_ ;
	wire _w483_ ;
	wire _w482_ ;
	wire _w481_ ;
	wire _w480_ ;
	wire _w479_ ;
	wire _w478_ ;
	wire _w476_ ;
	wire _w477_ ;
	wire _w511_ ;
	wire _w464_ ;
	wire _w465_ ;
	wire _w466_ ;
	wire _w467_ ;
	wire _w468_ ;
	wire _w469_ ;
	wire _w757_ ;
	wire _w2573_ ;
	wire _w216_ ;
	wire _w5303_ ;
	wire _w1325_ ;
	wire _w473_ ;
	wire _w470_ ;
	wire _w471_ ;
	wire _w472_ ;
	wire _w474_ ;
	wire _w475_ ;
	wire _w492_ ;
	wire _w493_ ;
	wire _w494_ ;
	wire _w495_ ;
	wire _w496_ ;
	wire _w497_ ;
	wire _w498_ ;
	wire _w499_ ;
	wire _w500_ ;
	wire _w501_ ;
	wire _w502_ ;
	wire _w503_ ;
	wire _w504_ ;
	wire _w505_ ;
	wire _w506_ ;
	wire _w507_ ;
	wire _w508_ ;
	wire _w509_ ;
	wire _w510_ ;
	wire _w512_ ;
	wire _w513_ ;
	wire _w514_ ;
	wire _w515_ ;
	wire _w516_ ;
	wire _w517_ ;
	wire _w518_ ;
	wire _w519_ ;
	wire _w520_ ;
	wire _w521_ ;
	wire _w590_ ;
	wire _w591_ ;
	wire _w592_ ;
	wire _w593_ ;
	wire _w594_ ;
	wire _w595_ ;
	wire _w596_ ;
	wire _w597_ ;
	wire _w598_ ;
	wire _w599_ ;
	wire _w600_ ;
	wire _w601_ ;
	wire _w602_ ;
	wire _w603_ ;
	wire _w604_ ;
	wire _w605_ ;
	wire _w606_ ;
	wire _w607_ ;
	wire _w608_ ;
	wire _w609_ ;
	wire _w610_ ;
	wire _w611_ ;
	wire _w612_ ;
	wire _w613_ ;
	wire _w614_ ;
	wire _w615_ ;
	wire _w616_ ;
	wire _w617_ ;
	wire _w618_ ;
	wire _w619_ ;
	wire _w620_ ;
	wire _w621_ ;
	wire _w622_ ;
	wire _w623_ ;
	wire _w624_ ;
	wire _w625_ ;
	wire _w626_ ;
	wire _w627_ ;
	wire _w628_ ;
	wire _w629_ ;
	wire _w630_ ;
	wire _w631_ ;
	wire _w632_ ;
	wire _w633_ ;
	wire _w634_ ;
	wire _w635_ ;
	wire _w636_ ;
	wire _w637_ ;
	wire _w638_ ;
	wire _w639_ ;
	wire _w640_ ;
	wire _w641_ ;
	wire _w642_ ;
	wire _w643_ ;
	wire _w644_ ;
	wire _w645_ ;
	wire _w646_ ;
	wire _w647_ ;
	wire _w648_ ;
	wire _w649_ ;
	wire _w650_ ;
	wire _w651_ ;
	wire _w652_ ;
	wire _w653_ ;
	wire _w654_ ;
	wire _w655_ ;
	wire _w656_ ;
	wire _w657_ ;
	wire _w658_ ;
	wire _w659_ ;
	wire _w660_ ;
	wire _w661_ ;
	wire _w662_ ;
	wire _w663_ ;
	wire _w664_ ;
	wire _w665_ ;
	wire _w666_ ;
	wire _w667_ ;
	wire _w668_ ;
	wire _w669_ ;
	wire _w670_ ;
	wire _w671_ ;
	wire _w672_ ;
	wire _w673_ ;
	wire _w674_ ;
	wire _w675_ ;
	wire _w676_ ;
	wire _w677_ ;
	wire _w678_ ;
	wire _w679_ ;
	wire _w680_ ;
	wire _w681_ ;
	wire _w682_ ;
	wire _w683_ ;
	wire _w684_ ;
	wire _w685_ ;
	wire _w686_ ;
	wire _w687_ ;
	wire _w688_ ;
	wire _w689_ ;
	wire _w690_ ;
	wire _w691_ ;
	wire _w692_ ;
	wire _w693_ ;
	wire _w694_ ;
	wire _w695_ ;
	wire _w696_ ;
	wire _w697_ ;
	wire _w698_ ;
	wire _w699_ ;
	wire _w700_ ;
	wire _w701_ ;
	wire _w702_ ;
	wire _w703_ ;
	wire _w704_ ;
	wire _w705_ ;
	wire _w706_ ;
	wire _w707_ ;
	wire _w708_ ;
	wire _w709_ ;
	wire _w710_ ;
	wire _w711_ ;
	wire _w712_ ;
	wire _w713_ ;
	wire _w714_ ;
	wire _w715_ ;
	wire _w716_ ;
	wire _w717_ ;
	wire _w718_ ;
	wire _w719_ ;
	wire _w1004_ ;
	wire _w1005_ ;
	wire _w1006_ ;
	wire _w1007_ ;
	wire _w1008_ ;
	wire _w1009_ ;
	wire _w1010_ ;
	wire _w1011_ ;
	wire _w1012_ ;
	wire _w1013_ ;
	wire _w1014_ ;
	wire _w1015_ ;
	wire _w1016_ ;
	wire _w1017_ ;
	wire _w1018_ ;
	wire _w1019_ ;
	wire _w1020_ ;
	wire _w1021_ ;
	wire _w1022_ ;
	wire _w1023_ ;
	wire _w1024_ ;
	wire _w1025_ ;
	wire _w1026_ ;
	wire _w1027_ ;
	wire _w1028_ ;
	wire _w1029_ ;
	wire _w1030_ ;
	wire _w1031_ ;
	wire _w1032_ ;
	wire _w1033_ ;
	wire _w1034_ ;
	wire _w1035_ ;
	wire _w1036_ ;
	wire _w1037_ ;
	wire _w1038_ ;
	wire _w1039_ ;
	wire _w1040_ ;
	wire _w1041_ ;
	wire _w1042_ ;
	wire _w1043_ ;
	wire _w1044_ ;
	wire _w1045_ ;
	wire _w1046_ ;
	wire _w1047_ ;
	wire _w1048_ ;
	wire _w1049_ ;
	wire _w1050_ ;
	wire _w1051_ ;
	wire _w1052_ ;
	wire _w1053_ ;
	wire _w1054_ ;
	wire _w1055_ ;
	wire _w1056_ ;
	wire _w1057_ ;
	wire _w1058_ ;
	wire _w1059_ ;
	wire _w1060_ ;
	wire _w1061_ ;
	wire _w1062_ ;
	wire _w1063_ ;
	wire _w1064_ ;
	wire _w1065_ ;
	wire _w1066_ ;
	wire _w1067_ ;
	wire _w1068_ ;
	wire _w1069_ ;
	wire _w1070_ ;
	wire _w1071_ ;
	wire _w1072_ ;
	wire _w1073_ ;
	wire _w1074_ ;
	wire _w1075_ ;
	wire _w1076_ ;
	wire _w1077_ ;
	wire _w1078_ ;
	wire _w1079_ ;
	wire _w1080_ ;
	wire _w1081_ ;
	wire _w1082_ ;
	wire _w1083_ ;
	wire _w1084_ ;
	wire _w1085_ ;
	wire _w1086_ ;
	wire _w1087_ ;
	wire _w1088_ ;
	wire _w1089_ ;
	wire _w1090_ ;
	wire _w1091_ ;
	wire _w1092_ ;
	wire _w1093_ ;
	wire _w1094_ ;
	wire _w1095_ ;
	wire _w1096_ ;
	wire _w1097_ ;
	wire _w1098_ ;
	wire _w1099_ ;
	wire _w1100_ ;
	wire _w1101_ ;
	wire _w1102_ ;
	wire _w1103_ ;
	wire _w1104_ ;
	wire _w1105_ ;
	wire _w1106_ ;
	wire _w1107_ ;
	wire _w1108_ ;
	wire _w1109_ ;
	wire _w1110_ ;
	wire _w1111_ ;
	wire _w1112_ ;
	wire _w1113_ ;
	wire _w1114_ ;
	wire _w1115_ ;
	wire _w1116_ ;
	wire _w1117_ ;
	wire _w1118_ ;
	wire _w1119_ ;
	wire _w1120_ ;
	wire _w1121_ ;
	wire _w1122_ ;
	wire _w1123_ ;
	wire _w1124_ ;
	wire _w1125_ ;
	wire _w1126_ ;
	wire _w1127_ ;
	wire _w1128_ ;
	wire _w1129_ ;
	wire _w1130_ ;
	wire _w1131_ ;
	wire _w1132_ ;
	wire _w1133_ ;
	wire _w1134_ ;
	wire _w1135_ ;
	wire _w1136_ ;
	wire _w1137_ ;
	wire _w1138_ ;
	wire _w1139_ ;
	wire _w1140_ ;
	wire _w1141_ ;
	wire _w1142_ ;
	wire _w1143_ ;
	wire _w1144_ ;
	wire _w1145_ ;
	wire _w1146_ ;
	wire _w1147_ ;
	wire _w1148_ ;
	wire _w1149_ ;
	wire _w1150_ ;
	wire _w1151_ ;
	wire _w1152_ ;
	wire _w1153_ ;
	wire _w1154_ ;
	wire _w1155_ ;
	wire _w1156_ ;
	wire _w1157_ ;
	wire _w1158_ ;
	wire _w1159_ ;
	wire _w1160_ ;
	wire _w1161_ ;
	wire _w1162_ ;
	wire _w1163_ ;
	wire _w1164_ ;
	wire _w1165_ ;
	wire _w1166_ ;
	wire _w1167_ ;
	wire _w1168_ ;
	wire _w1169_ ;
	wire _w1170_ ;
	wire _w1171_ ;
	wire _w1172_ ;
	wire _w1173_ ;
	wire _w1174_ ;
	wire _w1175_ ;
	wire _w1176_ ;
	wire _w1177_ ;
	wire _w1178_ ;
	wire _w1179_ ;
	wire _w1180_ ;
	wire _w1181_ ;
	wire _w1182_ ;
	wire _w1183_ ;
	wire _w1184_ ;
	wire _w1185_ ;
	wire _w1186_ ;
	wire _w1187_ ;
	wire _w1188_ ;
	wire _w1189_ ;
	wire _w1190_ ;
	wire _w1191_ ;
	wire _w1192_ ;
	wire _w1193_ ;
	wire _w1194_ ;
	wire _w1195_ ;
	wire _w1196_ ;
	wire _w1197_ ;
	wire _w1198_ ;
	wire _w1199_ ;
	wire _w1200_ ;
	wire _w1201_ ;
	wire _w1202_ ;
	wire _w1203_ ;
	wire _w1204_ ;
	wire _w1205_ ;
	wire _w1206_ ;
	wire _w1207_ ;
	wire _w1208_ ;
	wire _w1209_ ;
	wire _w1210_ ;
	wire _w1211_ ;
	wire _w1212_ ;
	wire _w1213_ ;
	wire _w1214_ ;
	wire _w1215_ ;
	wire _w1216_ ;
	wire _w1217_ ;
	wire _w1218_ ;
	wire _w1219_ ;
	wire _w1220_ ;
	wire _w1221_ ;
	wire _w1222_ ;
	wire _w1223_ ;
	wire _w1224_ ;
	wire _w1225_ ;
	wire _w1226_ ;
	wire _w1227_ ;
	wire _w1228_ ;
	wire _w1229_ ;
	wire _w1230_ ;
	wire _w1231_ ;
	wire _w1232_ ;
	wire _w1233_ ;
	wire _w1234_ ;
	wire _w1235_ ;
	wire _w1236_ ;
	wire _w1237_ ;
	wire _w1238_ ;
	wire _w1239_ ;
	wire _w1240_ ;
	wire _w1241_ ;
	wire _w1242_ ;
	wire _w1243_ ;
	wire _w1244_ ;
	wire _w1245_ ;
	wire _w1246_ ;
	wire _w1247_ ;
	wire _w1248_ ;
	wire _w1249_ ;
	wire _w1250_ ;
	wire _w1251_ ;
	wire _w1252_ ;
	wire _w1253_ ;
	wire _w1254_ ;
	wire _w1255_ ;
	wire _w1256_ ;
	wire _w1257_ ;
	wire _w1258_ ;
	wire _w1259_ ;
	wire _w1260_ ;
	wire _w1261_ ;
	wire _w1262_ ;
	wire _w1263_ ;
	wire _w1264_ ;
	wire _w1265_ ;
	wire _w1266_ ;
	wire _w1267_ ;
	wire _w1268_ ;
	wire _w1269_ ;
	wire _w1270_ ;
	wire _w1271_ ;
	wire _w1272_ ;
	wire _w1273_ ;
	wire _w1274_ ;
	wire _w1275_ ;
	wire _w1276_ ;
	wire _w1277_ ;
	wire _w1278_ ;
	wire _w1279_ ;
	wire _w1280_ ;
	wire _w1281_ ;
	wire _w1282_ ;
	wire _w1283_ ;
	wire _w1284_ ;
	wire _w1285_ ;
	wire _w1286_ ;
	wire _w1287_ ;
	wire _w1288_ ;
	wire _w1289_ ;
	wire _w1290_ ;
	wire _w1291_ ;
	wire _w1292_ ;
	wire _w1293_ ;
	wire _w1294_ ;
	wire _w1295_ ;
	wire _w1296_ ;
	wire _w1297_ ;
	wire _w1298_ ;
	wire _w1299_ ;
	wire _w1300_ ;
	wire _w1301_ ;
	wire _w1302_ ;
	wire _w1303_ ;
	wire _w1304_ ;
	wire _w1305_ ;
	wire _w1306_ ;
	wire _w1307_ ;
	wire _w1308_ ;
	wire _w1309_ ;
	wire _w1310_ ;
	wire _w1311_ ;
	wire _w1312_ ;
	wire _w1313_ ;
	wire _w1314_ ;
	wire _w1315_ ;
	wire _w1316_ ;
	wire _w1317_ ;
	wire _w1318_ ;
	wire _w1319_ ;
	wire _w1320_ ;
	wire _w1321_ ;
	wire _w1322_ ;
	wire _w1323_ ;
	wire _w1324_ ;
	wire _w1326_ ;
	wire _w1327_ ;
	wire _w1328_ ;
	wire _w1329_ ;
	wire _w1330_ ;
	wire _w1331_ ;
	wire _w1332_ ;
	wire _w1333_ ;
	wire _w1334_ ;
	wire _w1335_ ;
	wire _w1336_ ;
	wire _w1337_ ;
	wire _w1338_ ;
	wire _w1339_ ;
	wire _w1340_ ;
	wire _w1341_ ;
	wire _w1342_ ;
	wire _w1343_ ;
	wire _w1344_ ;
	wire _w1345_ ;
	wire _w1346_ ;
	wire _w1347_ ;
	wire _w1348_ ;
	wire _w1349_ ;
	wire _w1350_ ;
	wire _w1351_ ;
	wire _w1352_ ;
	wire _w1353_ ;
	wire _w1354_ ;
	wire _w1355_ ;
	wire _w1356_ ;
	wire _w1357_ ;
	wire _w1358_ ;
	wire _w1359_ ;
	wire _w1360_ ;
	wire _w1361_ ;
	wire _w1362_ ;
	wire _w1363_ ;
	wire _w1364_ ;
	wire _w1365_ ;
	wire _w1366_ ;
	wire _w1367_ ;
	wire _w1368_ ;
	wire _w1369_ ;
	wire _w1370_ ;
	wire _w1371_ ;
	wire _w1372_ ;
	wire _w1373_ ;
	wire _w1374_ ;
	wire _w1375_ ;
	wire _w1376_ ;
	wire _w1377_ ;
	wire _w1378_ ;
	wire _w1379_ ;
	wire _w1380_ ;
	wire _w1381_ ;
	wire _w1382_ ;
	wire _w1383_ ;
	wire _w1384_ ;
	wire _w1385_ ;
	wire _w1386_ ;
	wire _w1387_ ;
	wire _w1388_ ;
	wire _w1389_ ;
	wire _w1390_ ;
	wire _w1391_ ;
	wire _w1392_ ;
	wire _w1393_ ;
	wire _w1394_ ;
	wire _w1395_ ;
	wire _w1396_ ;
	wire _w1397_ ;
	wire _w1398_ ;
	wire _w1399_ ;
	wire _w1400_ ;
	wire _w1401_ ;
	wire _w1402_ ;
	wire _w1403_ ;
	wire _w1404_ ;
	wire _w1405_ ;
	wire _w1406_ ;
	wire _w1407_ ;
	wire _w1408_ ;
	wire _w1409_ ;
	wire _w1410_ ;
	wire _w1411_ ;
	wire _w1412_ ;
	wire _w1413_ ;
	wire _w1414_ ;
	wire _w1415_ ;
	wire _w1416_ ;
	wire _w1417_ ;
	wire _w1418_ ;
	wire _w1419_ ;
	wire _w1420_ ;
	wire _w1421_ ;
	wire _w1422_ ;
	wire _w1423_ ;
	wire _w1424_ ;
	wire _w1425_ ;
	wire _w1426_ ;
	wire _w1427_ ;
	wire _w1428_ ;
	wire _w1429_ ;
	wire _w1430_ ;
	wire _w1431_ ;
	wire _w1432_ ;
	wire _w1433_ ;
	wire _w1434_ ;
	wire _w1435_ ;
	wire _w1436_ ;
	wire _w1437_ ;
	wire _w1438_ ;
	wire _w1439_ ;
	wire _w1440_ ;
	wire _w1441_ ;
	wire _w1442_ ;
	wire _w1443_ ;
	wire _w1444_ ;
	wire _w1445_ ;
	wire _w1446_ ;
	wire _w1447_ ;
	wire _w1448_ ;
	wire _w1449_ ;
	wire _w1450_ ;
	wire _w1451_ ;
	wire _w1452_ ;
	wire _w1453_ ;
	wire _w1454_ ;
	wire _w1455_ ;
	wire _w1456_ ;
	wire _w1457_ ;
	wire _w1458_ ;
	wire _w1459_ ;
	wire _w1460_ ;
	wire _w1461_ ;
	wire _w1462_ ;
	wire _w1463_ ;
	wire _w1464_ ;
	wire _w1465_ ;
	wire _w1466_ ;
	wire _w1467_ ;
	wire _w1468_ ;
	wire _w1469_ ;
	wire _w1470_ ;
	wire _w1471_ ;
	wire _w1472_ ;
	wire _w1473_ ;
	wire _w1474_ ;
	wire _w1475_ ;
	wire _w1476_ ;
	wire _w1477_ ;
	wire _w1478_ ;
	wire _w1479_ ;
	wire _w1480_ ;
	wire _w1481_ ;
	wire _w1482_ ;
	wire _w1483_ ;
	wire _w1484_ ;
	wire _w1485_ ;
	wire _w1486_ ;
	wire _w1487_ ;
	wire _w1488_ ;
	wire _w1489_ ;
	wire _w1490_ ;
	wire _w1491_ ;
	wire _w1492_ ;
	wire _w1493_ ;
	wire _w1494_ ;
	wire _w1495_ ;
	wire _w1496_ ;
	wire _w1497_ ;
	wire _w1498_ ;
	wire _w1499_ ;
	wire _w1500_ ;
	wire _w1501_ ;
	wire _w1502_ ;
	wire _w1503_ ;
	wire _w1504_ ;
	wire _w1505_ ;
	wire _w1506_ ;
	wire _w1507_ ;
	wire _w1508_ ;
	wire _w1509_ ;
	wire _w1510_ ;
	wire _w1511_ ;
	wire _w1512_ ;
	wire _w1513_ ;
	wire _w1514_ ;
	wire _w1515_ ;
	wire _w1516_ ;
	wire _w1517_ ;
	wire _w1518_ ;
	wire _w1519_ ;
	wire _w1520_ ;
	wire _w1521_ ;
	wire _w1522_ ;
	wire _w1523_ ;
	wire _w1524_ ;
	wire _w1525_ ;
	wire _w1526_ ;
	wire _w1527_ ;
	wire _w1528_ ;
	wire _w1529_ ;
	wire _w1530_ ;
	wire _w1531_ ;
	wire _w1532_ ;
	wire _w1533_ ;
	wire _w1534_ ;
	wire _w1535_ ;
	wire _w1536_ ;
	wire _w1537_ ;
	wire _w1538_ ;
	wire _w1539_ ;
	wire _w1540_ ;
	wire _w1541_ ;
	wire _w1542_ ;
	wire _w1543_ ;
	wire _w1544_ ;
	wire _w1545_ ;
	wire _w1546_ ;
	wire _w1547_ ;
	wire _w1548_ ;
	wire _w1549_ ;
	wire _w1550_ ;
	wire _w1551_ ;
	wire _w1552_ ;
	wire _w1553_ ;
	wire _w1554_ ;
	wire _w1555_ ;
	wire _w1556_ ;
	wire _w1557_ ;
	wire _w1558_ ;
	wire _w1559_ ;
	wire _w1560_ ;
	wire _w1561_ ;
	wire _w1562_ ;
	wire _w1563_ ;
	wire _w1564_ ;
	wire _w1565_ ;
	wire _w1566_ ;
	wire _w1567_ ;
	wire _w1568_ ;
	wire _w1569_ ;
	wire _w1570_ ;
	wire _w1571_ ;
	wire _w2820_ ;
	wire _w2821_ ;
	wire _w2822_ ;
	wire _w2823_ ;
	wire _w2824_ ;
	wire _w2825_ ;
	wire _w2826_ ;
	wire _w2827_ ;
	wire _w2828_ ;
	wire _w2829_ ;
	wire _w2830_ ;
	wire _w2831_ ;
	wire _w2832_ ;
	wire _w2833_ ;
	wire _w2834_ ;
	wire _w2835_ ;
	wire _w2836_ ;
	wire _w2837_ ;
	wire _w2838_ ;
	wire _w2839_ ;
	wire _w2840_ ;
	wire _w2841_ ;
	wire _w2842_ ;
	wire _w2843_ ;
	wire _w2844_ ;
	wire _w2845_ ;
	wire _w2846_ ;
	wire _w2847_ ;
	wire _w2848_ ;
	wire _w2849_ ;
	wire _w2850_ ;
	wire _w2851_ ;
	wire _w2852_ ;
	wire _w2853_ ;
	wire _w2854_ ;
	wire _w2855_ ;
	wire _w2856_ ;
	wire _w2857_ ;
	wire _w2858_ ;
	wire _w2859_ ;
	wire _w2860_ ;
	wire _w2861_ ;
	wire _w2862_ ;
	wire _w2863_ ;
	wire _w2864_ ;
	wire _w2865_ ;
	wire _w2866_ ;
	wire _w2867_ ;
	wire _w2868_ ;
	wire _w2869_ ;
	wire _w2870_ ;
	wire _w2871_ ;
	wire _w2872_ ;
	wire _w2873_ ;
	wire _w2874_ ;
	wire _w2875_ ;
	wire _w2876_ ;
	wire _w2877_ ;
	wire _w2878_ ;
	wire _w2879_ ;
	wire _w2880_ ;
	wire _w2881_ ;
	wire _w2882_ ;
	wire _w2883_ ;
	wire _w2884_ ;
	wire _w2885_ ;
	wire _w2886_ ;
	wire _w2887_ ;
	wire _w2888_ ;
	wire _w2889_ ;
	wire _w2890_ ;
	wire _w2891_ ;
	wire _w2892_ ;
	wire _w2893_ ;
	wire _w2894_ ;
	wire _w2895_ ;
	wire _w2896_ ;
	wire _w2897_ ;
	wire _w2898_ ;
	wire _w2899_ ;
	wire _w2900_ ;
	wire _w2901_ ;
	wire _w2902_ ;
	wire _w2903_ ;
	wire _w2904_ ;
	wire _w2905_ ;
	wire _w2906_ ;
	wire _w2907_ ;
	wire _w2908_ ;
	wire _w2909_ ;
	wire _w2910_ ;
	wire _w2911_ ;
	wire _w2912_ ;
	wire _w2913_ ;
	wire _w2914_ ;
	wire _w2915_ ;
	wire _w2916_ ;
	wire _w2917_ ;
	wire _w2918_ ;
	wire _w2919_ ;
	wire _w2920_ ;
	wire _w2921_ ;
	wire _w2922_ ;
	wire _w2923_ ;
	wire _w2924_ ;
	wire _w2925_ ;
	wire _w2926_ ;
	wire _w2927_ ;
	wire _w2928_ ;
	wire _w2929_ ;
	wire _w2930_ ;
	wire _w2931_ ;
	wire _w2932_ ;
	wire _w2933_ ;
	wire _w2934_ ;
	wire _w2935_ ;
	wire _w2936_ ;
	wire _w2937_ ;
	wire _w2938_ ;
	wire _w2939_ ;
	wire _w2940_ ;
	wire _w2941_ ;
	wire _w2942_ ;
	wire _w2943_ ;
	wire _w2944_ ;
	wire _w2945_ ;
	wire _w2946_ ;
	wire _w2947_ ;
	wire _w2948_ ;
	wire _w2949_ ;
	wire _w2950_ ;
	wire _w2951_ ;
	wire _w2952_ ;
	wire _w2953_ ;
	wire _w2954_ ;
	wire _w2955_ ;
	wire _w2956_ ;
	wire _w2957_ ;
	wire _w2958_ ;
	wire _w2959_ ;
	wire _w2960_ ;
	wire _w2961_ ;
	wire _w2962_ ;
	wire _w2963_ ;
	wire _w2964_ ;
	wire _w2965_ ;
	wire _w2966_ ;
	wire _w2967_ ;
	wire _w2968_ ;
	wire _w2969_ ;
	wire _w2970_ ;
	wire _w2971_ ;
	wire _w2972_ ;
	wire _w2973_ ;
	wire _w2974_ ;
	wire _w2975_ ;
	wire _w2976_ ;
	wire _w2977_ ;
	wire _w2978_ ;
	wire _w2979_ ;
	wire _w2980_ ;
	wire _w2981_ ;
	wire _w2982_ ;
	wire _w2983_ ;
	wire _w2984_ ;
	wire _w2985_ ;
	wire _w2986_ ;
	wire _w2987_ ;
	wire _w2988_ ;
	wire _w2989_ ;
	wire _w2990_ ;
	wire _w2991_ ;
	wire _w2992_ ;
	wire _w2993_ ;
	wire _w2994_ ;
	wire _w2995_ ;
	wire _w2996_ ;
	wire _w2997_ ;
	wire _w2998_ ;
	wire _w2999_ ;
	wire _w3000_ ;
	wire _w3001_ ;
	wire _w3002_ ;
	wire _w3003_ ;
	wire _w3004_ ;
	wire _w3005_ ;
	wire _w3006_ ;
	wire _w3007_ ;
	wire _w3008_ ;
	wire _w3009_ ;
	wire _w3010_ ;
	wire _w3011_ ;
	wire _w3012_ ;
	wire _w3013_ ;
	wire _w3014_ ;
	wire _w3015_ ;
	wire _w3016_ ;
	wire _w3017_ ;
	wire _w3018_ ;
	wire _w3019_ ;
	wire _w3020_ ;
	wire _w3021_ ;
	wire _w3022_ ;
	wire _w3023_ ;
	wire _w3024_ ;
	wire _w3025_ ;
	wire _w3026_ ;
	wire _w3027_ ;
	wire _w3028_ ;
	wire _w3029_ ;
	wire _w3030_ ;
	wire _w3031_ ;
	wire _w3032_ ;
	wire _w3033_ ;
	wire _w3034_ ;
	wire _w3035_ ;
	wire _w3036_ ;
	wire _w3037_ ;
	wire _w3038_ ;
	wire _w3039_ ;
	wire _w3040_ ;
	wire _w3041_ ;
	wire _w3042_ ;
	wire _w3043_ ;
	wire _w3044_ ;
	wire _w3045_ ;
	wire _w3046_ ;
	wire _w3047_ ;
	wire _w3048_ ;
	wire _w3049_ ;
	wire _w3050_ ;
	wire _w3051_ ;
	wire _w3052_ ;
	wire _w3053_ ;
	wire _w3054_ ;
	wire _w3055_ ;
	wire _w3056_ ;
	wire _w3057_ ;
	wire _w3058_ ;
	wire _w3059_ ;
	wire _w3060_ ;
	wire _w3061_ ;
	wire _w3062_ ;
	wire _w3063_ ;
	wire _w3064_ ;
	wire _w3065_ ;
	wire _w3066_ ;
	wire _w3067_ ;
	wire _w3068_ ;
	wire _w3069_ ;
	wire _w3070_ ;
	wire _w3071_ ;
	wire _w3072_ ;
	wire _w3073_ ;
	wire _w3074_ ;
	wire _w3075_ ;
	wire _w3076_ ;
	wire _w3077_ ;
	wire _w3078_ ;
	wire _w3079_ ;
	wire _w3080_ ;
	wire _w3081_ ;
	wire _w3082_ ;
	wire _w3083_ ;
	wire _w3084_ ;
	wire _w3085_ ;
	wire _w3086_ ;
	wire _w3087_ ;
	wire _w3088_ ;
	wire _w3089_ ;
	wire _w3090_ ;
	wire _w3091_ ;
	wire _w3092_ ;
	wire _w3093_ ;
	wire _w3094_ ;
	wire _w3095_ ;
	wire _w3096_ ;
	wire _w3097_ ;
	wire _w3098_ ;
	wire _w3099_ ;
	wire _w3100_ ;
	wire _w3101_ ;
	wire _w3102_ ;
	wire _w3103_ ;
	wire _w3104_ ;
	wire _w3105_ ;
	wire _w3106_ ;
	wire _w3107_ ;
	wire _w3108_ ;
	wire _w3109_ ;
	wire _w3110_ ;
	wire _w3111_ ;
	wire _w3112_ ;
	wire _w3113_ ;
	wire _w3114_ ;
	wire _w3115_ ;
	wire _w3116_ ;
	wire _w3117_ ;
	wire _w3118_ ;
	wire _w3119_ ;
	wire _w3120_ ;
	wire _w3121_ ;
	wire _w3122_ ;
	wire _w3123_ ;
	wire _w3124_ ;
	wire _w3125_ ;
	wire _w3126_ ;
	wire _w3127_ ;
	wire _w3128_ ;
	wire _w3129_ ;
	wire _w3130_ ;
	wire _w3131_ ;
	wire _w3132_ ;
	wire _w3133_ ;
	wire _w3134_ ;
	wire _w3135_ ;
	wire _w3136_ ;
	wire _w3137_ ;
	wire _w3138_ ;
	wire _w3139_ ;
	wire _w3140_ ;
	wire _w3141_ ;
	wire _w3142_ ;
	wire _w3143_ ;
	wire _w3144_ ;
	wire _w3145_ ;
	wire _w3146_ ;
	wire _w3147_ ;
	wire _w3148_ ;
	wire _w3149_ ;
	wire _w3150_ ;
	wire _w3151_ ;
	wire _w3152_ ;
	wire _w3153_ ;
	wire _w3154_ ;
	wire _w3155_ ;
	wire _w3156_ ;
	wire _w3157_ ;
	wire _w3158_ ;
	wire _w3159_ ;
	wire _w3160_ ;
	wire _w3161_ ;
	wire _w3162_ ;
	wire _w3163_ ;
	wire _w3164_ ;
	wire _w3165_ ;
	wire _w3166_ ;
	wire _w3167_ ;
	wire _w3168_ ;
	wire _w3169_ ;
	wire _w3170_ ;
	wire _w3171_ ;
	wire _w3172_ ;
	wire _w3173_ ;
	wire _w3174_ ;
	wire _w3175_ ;
	wire _w3176_ ;
	wire _w3177_ ;
	wire _w3178_ ;
	wire _w3179_ ;
	wire _w3180_ ;
	wire _w3181_ ;
	wire _w3182_ ;
	wire _w3183_ ;
	wire _w3184_ ;
	wire _w3185_ ;
	wire _w3186_ ;
	wire _w3187_ ;
	wire _w3188_ ;
	wire _w3189_ ;
	wire _w3190_ ;
	wire _w3191_ ;
	wire _w3192_ ;
	wire _w3193_ ;
	wire _w3194_ ;
	wire _w3195_ ;
	wire _w3196_ ;
	wire _w3197_ ;
	wire _w3198_ ;
	wire _w3199_ ;
	wire _w3200_ ;
	wire _w3201_ ;
	wire _w3202_ ;
	wire _w3203_ ;
	wire _w3204_ ;
	wire _w3205_ ;
	wire _w3206_ ;
	wire _w3207_ ;
	wire _w3208_ ;
	wire _w3209_ ;
	wire _w3210_ ;
	wire _w3211_ ;
	wire _w3212_ ;
	wire _w3213_ ;
	wire _w3214_ ;
	wire _w3215_ ;
	wire _w3216_ ;
	wire _w3217_ ;
	wire _w3218_ ;
	wire _w3219_ ;
	wire _w3220_ ;
	wire _w3221_ ;
	wire _w3222_ ;
	wire _w3223_ ;
	wire _w3224_ ;
	wire _w3225_ ;
	wire _w3226_ ;
	wire _w3227_ ;
	wire _w3228_ ;
	wire _w3229_ ;
	wire _w3230_ ;
	wire _w3231_ ;
	wire _w3232_ ;
	wire _w3233_ ;
	wire _w3234_ ;
	wire _w3235_ ;
	wire _w3236_ ;
	wire _w3237_ ;
	wire _w3238_ ;
	wire _w3239_ ;
	wire _w3240_ ;
	wire _w3241_ ;
	wire _w3242_ ;
	wire _w3243_ ;
	wire _w3244_ ;
	wire _w3245_ ;
	wire _w3246_ ;
	wire _w3247_ ;
	wire _w3248_ ;
	wire _w3249_ ;
	wire _w3250_ ;
	wire _w3251_ ;
	wire _w3252_ ;
	wire _w3253_ ;
	wire _w3254_ ;
	wire _w3255_ ;
	wire _w3256_ ;
	wire _w3257_ ;
	wire _w3258_ ;
	wire _w3259_ ;
	wire _w3260_ ;
	wire _w3261_ ;
	wire _w3262_ ;
	wire _w3263_ ;
	wire _w3264_ ;
	wire _w3265_ ;
	wire _w3266_ ;
	wire _w3267_ ;
	wire _w3268_ ;
	wire _w3269_ ;
	wire _w3270_ ;
	wire _w3271_ ;
	wire _w3272_ ;
	wire _w3273_ ;
	wire _w3274_ ;
	wire _w3275_ ;
	wire _w3276_ ;
	wire _w3277_ ;
	wire _w3278_ ;
	wire _w3279_ ;
	wire _w3280_ ;
	wire _w3281_ ;
	wire _w3282_ ;
	wire _w3283_ ;
	wire _w3284_ ;
	wire _w3285_ ;
	wire _w3286_ ;
	wire _w3287_ ;
	wire _w3288_ ;
	wire _w3289_ ;
	wire _w3290_ ;
	wire _w3291_ ;
	wire _w3292_ ;
	wire _w3293_ ;
	wire _w3294_ ;
	wire _w3295_ ;
	wire _w3296_ ;
	wire _w3297_ ;
	wire _w3298_ ;
	wire _w3299_ ;
	wire _w3300_ ;
	wire _w3301_ ;
	wire _w3302_ ;
	wire _w3303_ ;
	wire _w3304_ ;
	wire _w3305_ ;
	wire _w3306_ ;
	wire _w3307_ ;
	wire _w3308_ ;
	wire _w3309_ ;
	wire _w3310_ ;
	wire _w3311_ ;
	wire _w3312_ ;
	wire _w3313_ ;
	wire _w3314_ ;
	wire _w3315_ ;
	wire _w3316_ ;
	wire _w3317_ ;
	wire _w3318_ ;
	wire _w3319_ ;
	wire _w3320_ ;
	wire _w3321_ ;
	wire _w3322_ ;
	wire _w3323_ ;
	wire _w3324_ ;
	wire _w3325_ ;
	wire _w3326_ ;
	wire _w3327_ ;
	wire _w3328_ ;
	wire _w3329_ ;
	wire _w3330_ ;
	wire _w3331_ ;
	wire _w3332_ ;
	wire _w3333_ ;
	wire _w3334_ ;
	wire _w3335_ ;
	wire _w3336_ ;
	wire _w3337_ ;
	wire _w3338_ ;
	wire _w3339_ ;
	wire _w3340_ ;
	wire _w3341_ ;
	wire _w3342_ ;
	wire _w3343_ ;
	wire _w3344_ ;
	wire _w3345_ ;
	wire _w3346_ ;
	wire _w3347_ ;
	wire _w3348_ ;
	wire _w3349_ ;
	wire _w3350_ ;
	wire _w3351_ ;
	wire _w3352_ ;
	wire _w3353_ ;
	wire _w3354_ ;
	wire _w3355_ ;
	wire _w3356_ ;
	wire _w3357_ ;
	wire _w3358_ ;
	wire _w3359_ ;
	wire _w3360_ ;
	wire _w3361_ ;
	wire _w3362_ ;
	wire _w3363_ ;
	wire _w3364_ ;
	wire _w3365_ ;
	wire _w3366_ ;
	wire _w3367_ ;
	wire _w3368_ ;
	wire _w3369_ ;
	wire _w3370_ ;
	wire _w3371_ ;
	wire _w3372_ ;
	wire _w3373_ ;
	wire _w3374_ ;
	wire _w3375_ ;
	wire _w3376_ ;
	wire _w3377_ ;
	wire _w3378_ ;
	wire _w3379_ ;
	wire _w3380_ ;
	wire _w3381_ ;
	wire _w3382_ ;
	wire _w3383_ ;
	wire _w3384_ ;
	wire _w3385_ ;
	wire _w3386_ ;
	wire _w3387_ ;
	wire _w3388_ ;
	wire _w3389_ ;
	wire _w3390_ ;
	wire _w3391_ ;
	wire _w3392_ ;
	wire _w3393_ ;
	wire _w3394_ ;
	wire _w3395_ ;
	wire _w3396_ ;
	wire _w3397_ ;
	wire _w3398_ ;
	wire _w3399_ ;
	wire _w3400_ ;
	wire _w3401_ ;
	wire _w3402_ ;
	wire _w3403_ ;
	wire _w3404_ ;
	wire _w3405_ ;
	wire _w3406_ ;
	wire _w3407_ ;
	wire _w3408_ ;
	wire _w3409_ ;
	wire _w3410_ ;
	wire _w3411_ ;
	wire _w3412_ ;
	wire _w3413_ ;
	wire _w3414_ ;
	wire _w3415_ ;
	wire _w3416_ ;
	wire _w3417_ ;
	wire _w3418_ ;
	wire _w3419_ ;
	wire _w3420_ ;
	wire _w3421_ ;
	wire _w3422_ ;
	wire _w3423_ ;
	wire _w3424_ ;
	wire _w3425_ ;
	wire _w3426_ ;
	wire _w3427_ ;
	wire _w3428_ ;
	wire _w3429_ ;
	wire _w3430_ ;
	wire _w3431_ ;
	wire _w3432_ ;
	wire _w3433_ ;
	wire _w3434_ ;
	wire _w3435_ ;
	wire _w3436_ ;
	wire _w3437_ ;
	wire _w3438_ ;
	wire _w3439_ ;
	wire _w3440_ ;
	wire _w3441_ ;
	wire _w3442_ ;
	wire _w3443_ ;
	wire _w3444_ ;
	wire _w3445_ ;
	wire _w3446_ ;
	wire _w3447_ ;
	wire _w3448_ ;
	wire _w3449_ ;
	wire _w3450_ ;
	wire _w3451_ ;
	wire _w3452_ ;
	wire _w3453_ ;
	wire _w3454_ ;
	wire _w3455_ ;
	wire _w3456_ ;
	wire _w3457_ ;
	wire _w3458_ ;
	wire _w3459_ ;
	wire _w3460_ ;
	wire _w3461_ ;
	wire _w3462_ ;
	wire _w3463_ ;
	wire _w3464_ ;
	wire _w3465_ ;
	wire _w3466_ ;
	wire _w3467_ ;
	wire _w3468_ ;
	wire _w3469_ ;
	wire _w3470_ ;
	wire _w3471_ ;
	wire _w3472_ ;
	wire _w3473_ ;
	wire _w3474_ ;
	wire _w3475_ ;
	wire _w3476_ ;
	wire _w3477_ ;
	wire _w3478_ ;
	wire _w3479_ ;
	wire _w3480_ ;
	wire _w3481_ ;
	wire _w3482_ ;
	wire _w3483_ ;
	wire _w3484_ ;
	wire _w3485_ ;
	wire _w3486_ ;
	wire _w3487_ ;
	wire _w3488_ ;
	wire _w3489_ ;
	wire _w3490_ ;
	wire _w3491_ ;
	wire _w3492_ ;
	wire _w3493_ ;
	wire _w3494_ ;
	wire _w3495_ ;
	wire _w3496_ ;
	wire _w3497_ ;
	wire _w3498_ ;
	wire _w3499_ ;
	wire _w3500_ ;
	wire _w3501_ ;
	wire _w3502_ ;
	wire _w3503_ ;
	wire _w3504_ ;
	wire _w3505_ ;
	wire _w3506_ ;
	wire _w3507_ ;
	wire _w3508_ ;
	wire _w3509_ ;
	wire _w3510_ ;
	wire _w3511_ ;
	wire _w3512_ ;
	wire _w3513_ ;
	wire _w3514_ ;
	wire _w3515_ ;
	wire _w3516_ ;
	wire _w3517_ ;
	wire _w3518_ ;
	wire _w3519_ ;
	wire _w3520_ ;
	wire _w3521_ ;
	wire _w3522_ ;
	wire _w3523_ ;
	wire _w3524_ ;
	wire _w3525_ ;
	wire _w3526_ ;
	wire _w3527_ ;
	wire _w3528_ ;
	wire _w3529_ ;
	wire _w3530_ ;
	wire _w3531_ ;
	wire _w3532_ ;
	wire _w3533_ ;
	wire _w3534_ ;
	wire _w3535_ ;
	wire _w3536_ ;
	wire _w3537_ ;
	wire _w3538_ ;
	wire _w3539_ ;
	wire _w3540_ ;
	wire _w3541_ ;
	wire _w3542_ ;
	wire _w3543_ ;
	wire _w3544_ ;
	wire _w3545_ ;
	wire _w3546_ ;
	wire _w3547_ ;
	wire _w3548_ ;
	wire _w3549_ ;
	wire _w3550_ ;
	wire _w3551_ ;
	wire _w3552_ ;
	wire _w3553_ ;
	wire _w3554_ ;
	wire _w3555_ ;
	wire _w3556_ ;
	wire _w3557_ ;
	wire _w3558_ ;
	wire _w3559_ ;
	wire _w3560_ ;
	wire _w3561_ ;
	wire _w3562_ ;
	wire _w3563_ ;
	wire _w3564_ ;
	wire _w3565_ ;
	wire _w3566_ ;
	wire _w3567_ ;
	wire _w3568_ ;
	wire _w3569_ ;
	wire _w3570_ ;
	wire _w3571_ ;
	wire _w3572_ ;
	wire _w3573_ ;
	wire _w3574_ ;
	wire _w3575_ ;
	wire _w3576_ ;
	wire _w3577_ ;
	wire _w3578_ ;
	wire _w3579_ ;
	wire _w3580_ ;
	wire _w3581_ ;
	wire _w3582_ ;
	wire _w3583_ ;
	wire _w3584_ ;
	wire _w3585_ ;
	wire _w3586_ ;
	wire _w3587_ ;
	wire _w3588_ ;
	wire _w3589_ ;
	wire _w3590_ ;
	wire _w3591_ ;
	wire _w3592_ ;
	wire _w3593_ ;
	wire _w3594_ ;
	wire _w3595_ ;
	wire _w3596_ ;
	wire _w3597_ ;
	wire _w3598_ ;
	wire _w3599_ ;
	wire _w3600_ ;
	wire _w3601_ ;
	wire _w3602_ ;
	wire _w3603_ ;
	wire _w3604_ ;
	wire _w3605_ ;
	wire _w3606_ ;
	wire _w3607_ ;
	wire _w3608_ ;
	wire _w3609_ ;
	wire _w3610_ ;
	wire _w3611_ ;
	wire _w3612_ ;
	wire _w3613_ ;
	wire _w3614_ ;
	wire _w3615_ ;
	wire _w3616_ ;
	wire _w3617_ ;
	wire _w3618_ ;
	wire _w3619_ ;
	wire _w3620_ ;
	wire _w3621_ ;
	wire _w3622_ ;
	wire _w3623_ ;
	wire _w3624_ ;
	wire _w3625_ ;
	wire _w3626_ ;
	wire _w3627_ ;
	wire _w3628_ ;
	wire _w3629_ ;
	wire _w3630_ ;
	wire _w3631_ ;
	wire _w3632_ ;
	wire _w3633_ ;
	wire _w3634_ ;
	wire _w3635_ ;
	wire _w3636_ ;
	wire _w3637_ ;
	wire _w3638_ ;
	wire _w3639_ ;
	wire _w3640_ ;
	wire _w3641_ ;
	wire _w3642_ ;
	wire _w3643_ ;
	wire _w3644_ ;
	wire _w3645_ ;
	wire _w3646_ ;
	wire _w3647_ ;
	wire _w3648_ ;
	wire _w3649_ ;
	wire _w3650_ ;
	wire _w3651_ ;
	wire _w3652_ ;
	wire _w3653_ ;
	wire _w3654_ ;
	wire _w3655_ ;
	wire _w3656_ ;
	wire _w3657_ ;
	wire _w3658_ ;
	wire _w3659_ ;
	wire _w3660_ ;
	wire _w3661_ ;
	wire _w3662_ ;
	wire _w3663_ ;
	wire _w3664_ ;
	wire _w3665_ ;
	wire _w3666_ ;
	wire _w3667_ ;
	wire _w3668_ ;
	wire _w3669_ ;
	wire _w3670_ ;
	wire _w3671_ ;
	wire _w3672_ ;
	wire _w3673_ ;
	wire _w3674_ ;
	wire _w3675_ ;
	wire _w3676_ ;
	wire _w3677_ ;
	wire _w3678_ ;
	wire _w3679_ ;
	wire _w3680_ ;
	wire _w3681_ ;
	wire _w3682_ ;
	wire _w3683_ ;
	wire _w3684_ ;
	wire _w3685_ ;
	wire _w3686_ ;
	wire _w3687_ ;
	wire _w3688_ ;
	wire _w3689_ ;
	wire _w3690_ ;
	wire _w3691_ ;
	wire _w3692_ ;
	wire _w3693_ ;
	wire _w3694_ ;
	wire _w3695_ ;
	wire _w3696_ ;
	wire _w3697_ ;
	wire _w3698_ ;
	wire _w3699_ ;
	wire _w3700_ ;
	wire _w3701_ ;
	wire _w3702_ ;
	wire _w3703_ ;
	wire _w3704_ ;
	wire _w3705_ ;
	wire _w3706_ ;
	wire _w3707_ ;
	wire _w3708_ ;
	wire _w3709_ ;
	wire _w3710_ ;
	wire _w3711_ ;
	wire _w3712_ ;
	wire _w3713_ ;
	wire _w3714_ ;
	wire _w3715_ ;
	wire _w3716_ ;
	wire _w3717_ ;
	wire _w3718_ ;
	wire _w3719_ ;
	wire _w3720_ ;
	wire _w3721_ ;
	wire _w3722_ ;
	wire _w3723_ ;
	wire _w3724_ ;
	wire _w3725_ ;
	wire _w3726_ ;
	wire _w3727_ ;
	wire _w3728_ ;
	wire _w3729_ ;
	wire _w3730_ ;
	wire _w3731_ ;
	wire _w3732_ ;
	wire _w3733_ ;
	wire _w3734_ ;
	wire _w3735_ ;
	wire _w3736_ ;
	wire _w3737_ ;
	wire _w3738_ ;
	wire _w3739_ ;
	wire _w3740_ ;
	wire _w3741_ ;
	wire _w3742_ ;
	wire _w3743_ ;
	wire _w3744_ ;
	wire _w3745_ ;
	wire _w3746_ ;
	wire _w3747_ ;
	wire _w3748_ ;
	wire _w3749_ ;
	wire _w3750_ ;
	wire _w3751_ ;
	wire _w3752_ ;
	wire _w3753_ ;
	wire _w3754_ ;
	wire _w3755_ ;
	wire _w3756_ ;
	wire _w3757_ ;
	wire _w3758_ ;
	wire _w3759_ ;
	wire _w3760_ ;
	wire _w3761_ ;
	wire _w3762_ ;
	wire _w3763_ ;
	wire _w3764_ ;
	wire _w3765_ ;
	wire _w3766_ ;
	wire _w3767_ ;
	wire _w3768_ ;
	wire _w3769_ ;
	wire _w3770_ ;
	wire _w3771_ ;
	wire _w3772_ ;
	wire _w3773_ ;
	wire _w3774_ ;
	wire _w3775_ ;
	wire _w3776_ ;
	wire _w3777_ ;
	wire _w3778_ ;
	wire _w3779_ ;
	wire _w3780_ ;
	wire _w3781_ ;
	wire _w3782_ ;
	wire _w3783_ ;
	wire _w3784_ ;
	wire _w3785_ ;
	wire _w3786_ ;
	wire _w3787_ ;
	wire _w3788_ ;
	wire _w3789_ ;
	wire _w3790_ ;
	wire _w3791_ ;
	wire _w3792_ ;
	wire _w3793_ ;
	wire _w3794_ ;
	wire _w3795_ ;
	wire _w3796_ ;
	wire _w3797_ ;
	wire _w3798_ ;
	wire _w3799_ ;
	wire _w3800_ ;
	wire _w3801_ ;
	wire _w3802_ ;
	wire _w3803_ ;
	wire _w3804_ ;
	wire _w3805_ ;
	wire _w3806_ ;
	wire _w3807_ ;
	wire _w3808_ ;
	wire _w3809_ ;
	wire _w3810_ ;
	wire _w3811_ ;
	wire _w3812_ ;
	wire _w3813_ ;
	wire _w3814_ ;
	wire _w3815_ ;
	wire _w3816_ ;
	wire _w3817_ ;
	wire _w3818_ ;
	wire _w3819_ ;
	wire _w3820_ ;
	wire _w3821_ ;
	wire _w3822_ ;
	wire _w3823_ ;
	wire _w3824_ ;
	wire _w3825_ ;
	wire _w3826_ ;
	wire _w3827_ ;
	wire _w3828_ ;
	wire _w3829_ ;
	wire _w3830_ ;
	wire _w3831_ ;
	wire _w3832_ ;
	wire _w3833_ ;
	wire _w3834_ ;
	wire _w3835_ ;
	wire _w3836_ ;
	wire _w3837_ ;
	wire _w3838_ ;
	wire _w3839_ ;
	wire _w3840_ ;
	wire _w3841_ ;
	wire _w3842_ ;
	wire _w3843_ ;
	wire _w3844_ ;
	wire _w3845_ ;
	wire _w3846_ ;
	wire _w3847_ ;
	wire _w3848_ ;
	wire _w3849_ ;
	wire _w3850_ ;
	wire _w3851_ ;
	wire _w3852_ ;
	wire _w3853_ ;
	wire _w3854_ ;
	wire _w3855_ ;
	wire _w3856_ ;
	wire _w3857_ ;
	wire _w3858_ ;
	wire _w3859_ ;
	wire _w3860_ ;
	wire _w3861_ ;
	wire _w3862_ ;
	wire _w3863_ ;
	wire _w3864_ ;
	wire _w3865_ ;
	wire _w3866_ ;
	wire _w3867_ ;
	wire _w3868_ ;
	wire _w3869_ ;
	wire _w3870_ ;
	wire _w3871_ ;
	wire _w3872_ ;
	wire _w3873_ ;
	wire _w3874_ ;
	wire _w3875_ ;
	wire _w3876_ ;
	wire _w3877_ ;
	wire _w3878_ ;
	wire _w3879_ ;
	wire _w3880_ ;
	wire _w3881_ ;
	wire _w3882_ ;
	wire _w3883_ ;
	wire _w3884_ ;
	wire _w3885_ ;
	wire _w3886_ ;
	wire _w3887_ ;
	wire _w3888_ ;
	wire _w3889_ ;
	wire _w3890_ ;
	wire _w3891_ ;
	wire _w3892_ ;
	wire _w3893_ ;
	wire _w3894_ ;
	wire _w3895_ ;
	wire _w3896_ ;
	wire _w3897_ ;
	wire _w3898_ ;
	wire _w3899_ ;
	wire _w3900_ ;
	wire _w3901_ ;
	wire _w3902_ ;
	wire _w3903_ ;
	wire _w3904_ ;
	wire _w3905_ ;
	wire _w3906_ ;
	wire _w3907_ ;
	wire _w3908_ ;
	wire _w3909_ ;
	wire _w3910_ ;
	wire _w3911_ ;
	wire _w3912_ ;
	wire _w3913_ ;
	wire _w3914_ ;
	wire _w3915_ ;
	wire _w3916_ ;
	wire _w3917_ ;
	wire _w3918_ ;
	wire _w3919_ ;
	wire _w3920_ ;
	wire _w3921_ ;
	wire _w3922_ ;
	wire _w3923_ ;
	wire _w3924_ ;
	wire _w3925_ ;
	wire _w3926_ ;
	wire _w3927_ ;
	wire _w3928_ ;
	wire _w3929_ ;
	wire _w3930_ ;
	wire _w3931_ ;
	wire _w3932_ ;
	wire _w3933_ ;
	wire _w3934_ ;
	wire _w3935_ ;
	wire _w3936_ ;
	wire _w3937_ ;
	wire _w3938_ ;
	wire _w3939_ ;
	wire _w3940_ ;
	wire _w3941_ ;
	wire _w3942_ ;
	wire _w3943_ ;
	wire _w3944_ ;
	wire _w3945_ ;
	wire _w3946_ ;
	wire _w3947_ ;
	wire _w3948_ ;
	wire _w3949_ ;
	wire _w3950_ ;
	wire _w3951_ ;
	wire _w3952_ ;
	wire _w3953_ ;
	wire _w3954_ ;
	wire _w3955_ ;
	wire _w3956_ ;
	wire _w3957_ ;
	wire _w3958_ ;
	wire _w3959_ ;
	wire _w3960_ ;
	wire _w3961_ ;
	wire _w3962_ ;
	wire _w3963_ ;
	wire _w3964_ ;
	wire _w3965_ ;
	wire _w3966_ ;
	wire _w3967_ ;
	wire _w3968_ ;
	wire _w3969_ ;
	wire _w3970_ ;
	wire _w3971_ ;
	wire _w3972_ ;
	wire _w3973_ ;
	wire _w3974_ ;
	wire _w3975_ ;
	wire _w3976_ ;
	wire _w3977_ ;
	wire _w3978_ ;
	wire _w3979_ ;
	wire _w3980_ ;
	wire _w3981_ ;
	wire _w3982_ ;
	wire _w3983_ ;
	wire _w3984_ ;
	wire _w3985_ ;
	wire _w3986_ ;
	wire _w3987_ ;
	wire _w3988_ ;
	wire _w3989_ ;
	wire _w3990_ ;
	wire _w3991_ ;
	wire _w3992_ ;
	wire _w3993_ ;
	wire _w3994_ ;
	wire _w3995_ ;
	wire _w3996_ ;
	wire _w3997_ ;
	wire _w3998_ ;
	wire _w3999_ ;
	wire _w4000_ ;
	wire _w4001_ ;
	wire _w4002_ ;
	wire _w4003_ ;
	wire _w4004_ ;
	wire _w4005_ ;
	wire _w4006_ ;
	wire _w4007_ ;
	wire _w4008_ ;
	wire _w4009_ ;
	wire _w4010_ ;
	wire _w4011_ ;
	wire _w4012_ ;
	wire _w4013_ ;
	wire _w4014_ ;
	wire _w4015_ ;
	wire _w4016_ ;
	wire _w4017_ ;
	wire _w4018_ ;
	wire _w4019_ ;
	wire _w4020_ ;
	wire _w4021_ ;
	wire _w4022_ ;
	wire _w4023_ ;
	wire _w4024_ ;
	wire _w4025_ ;
	wire _w4026_ ;
	wire _w4027_ ;
	wire _w4028_ ;
	wire _w4029_ ;
	wire _w4030_ ;
	wire _w4031_ ;
	wire _w4032_ ;
	wire _w4033_ ;
	wire _w4034_ ;
	wire _w4035_ ;
	wire _w4036_ ;
	wire _w4037_ ;
	wire _w4038_ ;
	wire _w4039_ ;
	wire _w4040_ ;
	wire _w4041_ ;
	wire _w4042_ ;
	wire _w4043_ ;
	wire _w4044_ ;
	wire _w4045_ ;
	wire _w4046_ ;
	wire _w4047_ ;
	wire _w4048_ ;
	wire _w4049_ ;
	wire _w4050_ ;
	wire _w4051_ ;
	wire _w4052_ ;
	wire _w4053_ ;
	wire _w4054_ ;
	wire _w4055_ ;
	wire _w4056_ ;
	wire _w4057_ ;
	wire _w4058_ ;
	wire _w4059_ ;
	wire _w4060_ ;
	wire _w4061_ ;
	wire _w4062_ ;
	wire _w4063_ ;
	wire _w4064_ ;
	wire _w4065_ ;
	wire _w4066_ ;
	wire _w4067_ ;
	wire _w4068_ ;
	wire _w4069_ ;
	wire _w4070_ ;
	wire _w4071_ ;
	wire _w4072_ ;
	wire _w4073_ ;
	wire _w4074_ ;
	wire _w4075_ ;
	wire _w4076_ ;
	wire _w4077_ ;
	wire _w4078_ ;
	wire _w4079_ ;
	wire _w4080_ ;
	wire _w4081_ ;
	wire _w4082_ ;
	wire _w4083_ ;
	wire _w4084_ ;
	wire _w4085_ ;
	wire _w4086_ ;
	wire _w4087_ ;
	wire _w4088_ ;
	wire _w4089_ ;
	wire _w4090_ ;
	wire _w4091_ ;
	wire _w4092_ ;
	wire _w4093_ ;
	wire _w4094_ ;
	wire _w4095_ ;
	wire _w4096_ ;
	wire _w4097_ ;
	wire _w4098_ ;
	wire _w4099_ ;
	wire _w4100_ ;
	wire _w4101_ ;
	wire _w4102_ ;
	wire _w4103_ ;
	wire _w4104_ ;
	wire _w4105_ ;
	wire _w4106_ ;
	wire _w4107_ ;
	wire _w4108_ ;
	wire _w4109_ ;
	wire _w4110_ ;
	wire _w4111_ ;
	wire _w4112_ ;
	wire _w4113_ ;
	wire _w4114_ ;
	wire _w4115_ ;
	wire _w4116_ ;
	wire _w4117_ ;
	wire _w4118_ ;
	wire _w4119_ ;
	wire _w4120_ ;
	wire _w4121_ ;
	wire _w4122_ ;
	wire _w4123_ ;
	wire _w4124_ ;
	wire _w4125_ ;
	wire _w4126_ ;
	wire _w4127_ ;
	wire _w4128_ ;
	wire _w4129_ ;
	wire _w4130_ ;
	wire _w4131_ ;
	wire _w4132_ ;
	wire _w4133_ ;
	wire _w4134_ ;
	wire _w4135_ ;
	wire _w4136_ ;
	wire _w4137_ ;
	wire _w4138_ ;
	wire _w4139_ ;
	wire _w4140_ ;
	wire _w4141_ ;
	wire _w4142_ ;
	wire _w4143_ ;
	wire _w4144_ ;
	wire _w4145_ ;
	wire _w4146_ ;
	wire _w4147_ ;
	wire _w4148_ ;
	wire _w4149_ ;
	wire _w4150_ ;
	wire _w4151_ ;
	wire _w4152_ ;
	wire _w4153_ ;
	wire _w4154_ ;
	wire _w4155_ ;
	wire _w4156_ ;
	wire _w4157_ ;
	wire _w4158_ ;
	wire _w4159_ ;
	wire _w4160_ ;
	wire _w4161_ ;
	wire _w4162_ ;
	wire _w4163_ ;
	wire _w4164_ ;
	wire _w4165_ ;
	wire _w4166_ ;
	wire _w4167_ ;
	wire _w4168_ ;
	wire _w4169_ ;
	wire _w4170_ ;
	wire _w4171_ ;
	wire _w4172_ ;
	wire _w4173_ ;
	wire _w4174_ ;
	wire _w4175_ ;
	wire _w4176_ ;
	wire _w4177_ ;
	wire _w4178_ ;
	wire _w4179_ ;
	wire _w4180_ ;
	wire _w4181_ ;
	wire _w4182_ ;
	wire _w4183_ ;
	wire _w4184_ ;
	wire _w4185_ ;
	wire _w4186_ ;
	wire _w4187_ ;
	wire _w4188_ ;
	wire _w4189_ ;
	wire _w4190_ ;
	wire _w4191_ ;
	wire _w4192_ ;
	wire _w4193_ ;
	wire _w4194_ ;
	wire _w4195_ ;
	wire _w4196_ ;
	wire _w4197_ ;
	wire _w4198_ ;
	wire _w4199_ ;
	wire _w4200_ ;
	wire _w4201_ ;
	wire _w4202_ ;
	wire _w4203_ ;
	wire _w4204_ ;
	wire _w4205_ ;
	wire _w4206_ ;
	wire _w4207_ ;
	wire _w4208_ ;
	wire _w4209_ ;
	wire _w4210_ ;
	wire _w4211_ ;
	wire _w4212_ ;
	wire _w4213_ ;
	wire _w4214_ ;
	wire _w4215_ ;
	wire _w4216_ ;
	wire _w4217_ ;
	wire _w4218_ ;
	wire _w4219_ ;
	wire _w4220_ ;
	wire _w4221_ ;
	wire _w4222_ ;
	wire _w4223_ ;
	wire _w4224_ ;
	wire _w4225_ ;
	wire _w4226_ ;
	wire _w4227_ ;
	wire _w4228_ ;
	wire _w4229_ ;
	wire _w4230_ ;
	wire _w4231_ ;
	wire _w4232_ ;
	wire _w4233_ ;
	wire _w4234_ ;
	wire _w4235_ ;
	wire _w4236_ ;
	wire _w4237_ ;
	wire _w4238_ ;
	wire _w4239_ ;
	wire _w4240_ ;
	wire _w4241_ ;
	wire _w4242_ ;
	wire _w4243_ ;
	wire _w4244_ ;
	wire _w4245_ ;
	wire _w4246_ ;
	wire _w4247_ ;
	wire _w4248_ ;
	wire _w4249_ ;
	wire _w4250_ ;
	wire _w4251_ ;
	wire _w4252_ ;
	wire _w4253_ ;
	wire _w4254_ ;
	wire _w4255_ ;
	wire _w4256_ ;
	wire _w4257_ ;
	wire _w4258_ ;
	wire _w4259_ ;
	wire _w4260_ ;
	wire _w4261_ ;
	wire _w4262_ ;
	wire _w4263_ ;
	wire _w4264_ ;
	wire _w4265_ ;
	wire _w4266_ ;
	wire _w4267_ ;
	wire _w4268_ ;
	wire _w4269_ ;
	wire _w4270_ ;
	wire _w4271_ ;
	wire _w4272_ ;
	wire _w4273_ ;
	wire _w4274_ ;
	wire _w4275_ ;
	wire _w4276_ ;
	wire _w4277_ ;
	wire _w4278_ ;
	wire _w4279_ ;
	wire _w4280_ ;
	wire _w4281_ ;
	wire _w4282_ ;
	wire _w4283_ ;
	wire _w4284_ ;
	wire _w4285_ ;
	wire _w4286_ ;
	wire _w4287_ ;
	wire _w4288_ ;
	wire _w4289_ ;
	wire _w4290_ ;
	wire _w4291_ ;
	wire _w4292_ ;
	wire _w4293_ ;
	wire _w4294_ ;
	wire _w4295_ ;
	wire _w4296_ ;
	wire _w4297_ ;
	wire _w4298_ ;
	wire _w4299_ ;
	wire _w4300_ ;
	wire _w4301_ ;
	wire _w4302_ ;
	wire _w4303_ ;
	wire _w4304_ ;
	wire _w4305_ ;
	wire _w4306_ ;
	wire _w4307_ ;
	wire _w4308_ ;
	wire _w4309_ ;
	wire _w4310_ ;
	wire _w4311_ ;
	wire _w4312_ ;
	wire _w4313_ ;
	wire _w4314_ ;
	wire _w4315_ ;
	wire _w4316_ ;
	wire _w4317_ ;
	wire _w4318_ ;
	wire _w4319_ ;
	wire _w4320_ ;
	wire _w4321_ ;
	wire _w4322_ ;
	wire _w4323_ ;
	wire _w4324_ ;
	wire _w4325_ ;
	wire _w4326_ ;
	wire _w4327_ ;
	wire _w4328_ ;
	wire _w4329_ ;
	wire _w4330_ ;
	wire _w4331_ ;
	wire _w4332_ ;
	wire _w4333_ ;
	wire _w4334_ ;
	wire _w4335_ ;
	wire _w4336_ ;
	wire _w4337_ ;
	wire _w4338_ ;
	wire _w4339_ ;
	wire _w4340_ ;
	wire _w4341_ ;
	wire _w4342_ ;
	wire _w4343_ ;
	wire _w4344_ ;
	wire _w4345_ ;
	wire _w4346_ ;
	wire _w4347_ ;
	wire _w4348_ ;
	wire _w4349_ ;
	wire _w4350_ ;
	wire _w4351_ ;
	wire _w4352_ ;
	wire _w4353_ ;
	wire _w4354_ ;
	wire _w4355_ ;
	wire _w4356_ ;
	wire _w4357_ ;
	wire _w4358_ ;
	wire _w4359_ ;
	wire _w4360_ ;
	wire _w4361_ ;
	wire _w4362_ ;
	wire _w4363_ ;
	wire _w4364_ ;
	wire _w4365_ ;
	wire _w4366_ ;
	wire _w4367_ ;
	wire _w4368_ ;
	wire _w4369_ ;
	wire _w4370_ ;
	wire _w4371_ ;
	wire _w4372_ ;
	wire _w4373_ ;
	wire _w4374_ ;
	wire _w4375_ ;
	wire _w4376_ ;
	wire _w4377_ ;
	wire _w4378_ ;
	wire _w4379_ ;
	wire _w4380_ ;
	wire _w4381_ ;
	wire _w4382_ ;
	wire _w4383_ ;
	wire _w4384_ ;
	wire _w4385_ ;
	wire _w4386_ ;
	wire _w4387_ ;
	wire _w4388_ ;
	wire _w4389_ ;
	wire _w4390_ ;
	wire _w4391_ ;
	wire _w4392_ ;
	wire _w4393_ ;
	wire _w4394_ ;
	wire _w4395_ ;
	wire _w4396_ ;
	wire _w4397_ ;
	wire _w4398_ ;
	wire _w4399_ ;
	wire _w4400_ ;
	wire _w4401_ ;
	wire _w4402_ ;
	wire _w4403_ ;
	wire _w4404_ ;
	wire _w4405_ ;
	wire _w4406_ ;
	wire _w4407_ ;
	wire _w4408_ ;
	wire _w4409_ ;
	wire _w4410_ ;
	wire _w4411_ ;
	wire _w4412_ ;
	wire _w4413_ ;
	wire _w4414_ ;
	wire _w4415_ ;
	wire _w4416_ ;
	wire _w4417_ ;
	wire _w4418_ ;
	wire _w4419_ ;
	wire _w4420_ ;
	wire _w4421_ ;
	wire _w4422_ ;
	wire _w4423_ ;
	wire _w4424_ ;
	wire _w4425_ ;
	wire _w4426_ ;
	wire _w4427_ ;
	wire _w4428_ ;
	wire _w4429_ ;
	wire _w4430_ ;
	wire _w4431_ ;
	wire _w4432_ ;
	wire _w4433_ ;
	wire _w4434_ ;
	wire _w4435_ ;
	wire _w4436_ ;
	wire _w4437_ ;
	wire _w4438_ ;
	wire _w4439_ ;
	wire _w4440_ ;
	wire _w4441_ ;
	wire _w4442_ ;
	wire _w4443_ ;
	wire _w4444_ ;
	wire _w4445_ ;
	wire _w4446_ ;
	wire _w4447_ ;
	wire _w4448_ ;
	wire _w4449_ ;
	wire _w4450_ ;
	wire _w4451_ ;
	wire _w4452_ ;
	wire _w4453_ ;
	wire _w4454_ ;
	wire _w4455_ ;
	wire _w4456_ ;
	wire _w4457_ ;
	wire _w4458_ ;
	wire _w4459_ ;
	wire _w4460_ ;
	wire _w4461_ ;
	wire _w4462_ ;
	wire _w4463_ ;
	wire _w4464_ ;
	wire _w4465_ ;
	wire _w4466_ ;
	wire _w4467_ ;
	wire _w4468_ ;
	wire _w4469_ ;
	wire _w4470_ ;
	wire _w4471_ ;
	wire _w4472_ ;
	wire _w4473_ ;
	wire _w4474_ ;
	wire _w4475_ ;
	wire _w4476_ ;
	wire _w4477_ ;
	wire _w4478_ ;
	wire _w4479_ ;
	wire _w4480_ ;
	wire _w4481_ ;
	wire _w4482_ ;
	wire _w4483_ ;
	wire _w4484_ ;
	wire _w4485_ ;
	wire _w4486_ ;
	wire _w4487_ ;
	wire _w4488_ ;
	wire _w4489_ ;
	wire _w4490_ ;
	wire _w4491_ ;
	wire _w4492_ ;
	wire _w4493_ ;
	wire _w4494_ ;
	wire _w4495_ ;
	wire _w4496_ ;
	wire _w4497_ ;
	wire _w4498_ ;
	wire _w4499_ ;
	wire _w4500_ ;
	wire _w4501_ ;
	wire _w4502_ ;
	wire _w4503_ ;
	wire _w4504_ ;
	wire _w4505_ ;
	wire _w4506_ ;
	wire _w4507_ ;
	wire _w4508_ ;
	wire _w4509_ ;
	wire _w4510_ ;
	wire _w4511_ ;
	wire _w4512_ ;
	wire _w4513_ ;
	wire _w4514_ ;
	wire _w4515_ ;
	wire _w4516_ ;
	wire _w4517_ ;
	wire _w4518_ ;
	wire _w4519_ ;
	wire _w4520_ ;
	wire _w4521_ ;
	wire _w4522_ ;
	wire _w4523_ ;
	wire _w4524_ ;
	wire _w4525_ ;
	wire _w4526_ ;
	wire _w4527_ ;
	wire _w4528_ ;
	wire _w4529_ ;
	wire _w4530_ ;
	wire _w4531_ ;
	wire _w4532_ ;
	wire _w4533_ ;
	wire _w4534_ ;
	wire _w4535_ ;
	wire _w4536_ ;
	wire _w4537_ ;
	wire _w4538_ ;
	wire _w4539_ ;
	wire _w4540_ ;
	wire _w4541_ ;
	wire _w4542_ ;
	wire _w4543_ ;
	wire _w4544_ ;
	wire _w4545_ ;
	wire _w4546_ ;
	wire _w4547_ ;
	wire _w4548_ ;
	wire _w4549_ ;
	wire _w4550_ ;
	wire _w4551_ ;
	wire _w4552_ ;
	wire _w4553_ ;
	wire _w4554_ ;
	wire _w4555_ ;
	wire _w4556_ ;
	wire _w4557_ ;
	wire _w4558_ ;
	wire _w4559_ ;
	wire _w4560_ ;
	wire _w4561_ ;
	wire _w4562_ ;
	wire _w4563_ ;
	wire _w4564_ ;
	wire _w4565_ ;
	wire _w4566_ ;
	wire _w4567_ ;
	wire _w4568_ ;
	wire _w4569_ ;
	wire _w4570_ ;
	wire _w4571_ ;
	wire _w4572_ ;
	wire _w4573_ ;
	wire _w4574_ ;
	wire _w4575_ ;
	wire _w4576_ ;
	wire _w4577_ ;
	wire _w4578_ ;
	wire _w4579_ ;
	wire _w4580_ ;
	wire _w4581_ ;
	wire _w4582_ ;
	wire _w4583_ ;
	wire _w4584_ ;
	wire _w4585_ ;
	wire _w4586_ ;
	wire _w4587_ ;
	wire _w4588_ ;
	wire _w4589_ ;
	wire _w4590_ ;
	wire _w4591_ ;
	wire _w4592_ ;
	wire _w4593_ ;
	wire _w4594_ ;
	wire _w4595_ ;
	wire _w4596_ ;
	wire _w4597_ ;
	wire _w4598_ ;
	wire _w4599_ ;
	wire _w4600_ ;
	wire _w4601_ ;
	wire _w4602_ ;
	wire _w4603_ ;
	wire _w4604_ ;
	wire _w4605_ ;
	wire _w4606_ ;
	wire _w4607_ ;
	wire _w4608_ ;
	wire _w4609_ ;
	wire _w4610_ ;
	wire _w4611_ ;
	wire _w4612_ ;
	wire _w4613_ ;
	wire _w4614_ ;
	wire _w4615_ ;
	wire _w4616_ ;
	wire _w4617_ ;
	wire _w4618_ ;
	wire _w4619_ ;
	wire _w4620_ ;
	wire _w4621_ ;
	wire _w4622_ ;
	wire _w4623_ ;
	wire _w4624_ ;
	wire _w4625_ ;
	wire _w4626_ ;
	wire _w4627_ ;
	wire _w4628_ ;
	wire _w4629_ ;
	wire _w4630_ ;
	wire _w4631_ ;
	wire _w4632_ ;
	wire _w4633_ ;
	wire _w4634_ ;
	wire _w4635_ ;
	wire _w4636_ ;
	wire _w4637_ ;
	wire _w4638_ ;
	wire _w4639_ ;
	wire _w4640_ ;
	wire _w4641_ ;
	wire _w4642_ ;
	wire _w4643_ ;
	wire _w4644_ ;
	wire _w4645_ ;
	wire _w4646_ ;
	wire _w4647_ ;
	wire _w4648_ ;
	wire _w4649_ ;
	wire _w4650_ ;
	wire _w4651_ ;
	wire _w4652_ ;
	wire _w4653_ ;
	wire _w4654_ ;
	wire _w4655_ ;
	wire _w4656_ ;
	wire _w4657_ ;
	wire _w4658_ ;
	wire _w4659_ ;
	wire _w4660_ ;
	wire _w4661_ ;
	wire _w4662_ ;
	wire _w4663_ ;
	wire _w4664_ ;
	wire _w4665_ ;
	wire _w4666_ ;
	wire _w4667_ ;
	wire _w4668_ ;
	wire _w4669_ ;
	wire _w4670_ ;
	wire _w4671_ ;
	wire _w4672_ ;
	wire _w4673_ ;
	wire _w4674_ ;
	wire _w4675_ ;
	wire _w4676_ ;
	wire _w4677_ ;
	wire _w4678_ ;
	wire _w4679_ ;
	wire _w4680_ ;
	wire _w4681_ ;
	wire _w4682_ ;
	wire _w4683_ ;
	wire _w4684_ ;
	wire _w4685_ ;
	wire _w4686_ ;
	wire _w4687_ ;
	wire _w4688_ ;
	wire _w4689_ ;
	wire _w4690_ ;
	wire _w4691_ ;
	wire _w4692_ ;
	wire _w4693_ ;
	wire _w4694_ ;
	wire _w4695_ ;
	wire _w4696_ ;
	wire _w4697_ ;
	wire _w4698_ ;
	wire _w4699_ ;
	wire _w4700_ ;
	wire _w4701_ ;
	wire _w4702_ ;
	wire _w4703_ ;
	wire _w4704_ ;
	wire _w4705_ ;
	wire _w4706_ ;
	wire _w4707_ ;
	wire _w4708_ ;
	wire _w4709_ ;
	wire _w4710_ ;
	wire _w4711_ ;
	wire _w4712_ ;
	wire _w4713_ ;
	wire _w4714_ ;
	wire _w4715_ ;
	wire _w4716_ ;
	wire _w4717_ ;
	wire _w4718_ ;
	wire _w4719_ ;
	wire _w4720_ ;
	wire _w4721_ ;
	wire _w4722_ ;
	wire _w4723_ ;
	wire _w4724_ ;
	wire _w4725_ ;
	wire _w4726_ ;
	wire _w4727_ ;
	wire _w4728_ ;
	wire _w4729_ ;
	wire _w4730_ ;
	wire _w4731_ ;
	wire _w4732_ ;
	wire _w4733_ ;
	wire _w4734_ ;
	wire _w4735_ ;
	wire _w4736_ ;
	wire _w4737_ ;
	wire _w4738_ ;
	wire _w4739_ ;
	wire _w4740_ ;
	wire _w4741_ ;
	wire _w4742_ ;
	wire _w4743_ ;
	wire _w4744_ ;
	wire _w4745_ ;
	wire _w4746_ ;
	wire _w4747_ ;
	wire _w4748_ ;
	wire _w4749_ ;
	wire _w4750_ ;
	wire _w4751_ ;
	wire _w4752_ ;
	wire _w4753_ ;
	wire _w4754_ ;
	wire _w4755_ ;
	wire _w4756_ ;
	wire _w4757_ ;
	wire _w4758_ ;
	wire _w4759_ ;
	wire _w4760_ ;
	wire _w4761_ ;
	wire _w4762_ ;
	wire _w4763_ ;
	wire _w4764_ ;
	wire _w4765_ ;
	wire _w4766_ ;
	wire _w4767_ ;
	wire _w4768_ ;
	wire _w4769_ ;
	wire _w4770_ ;
	wire _w4771_ ;
	wire _w4772_ ;
	wire _w4773_ ;
	wire _w4774_ ;
	wire _w4775_ ;
	wire _w4776_ ;
	wire _w4777_ ;
	wire _w4778_ ;
	wire _w4779_ ;
	wire _w4780_ ;
	wire _w4781_ ;
	wire _w4782_ ;
	wire _w4783_ ;
	wire _w4784_ ;
	wire _w4785_ ;
	wire _w4786_ ;
	wire _w4787_ ;
	wire _w4788_ ;
	wire _w4789_ ;
	wire _w4790_ ;
	wire _w4791_ ;
	wire _w4792_ ;
	wire _w4793_ ;
	wire _w4794_ ;
	wire _w4795_ ;
	wire _w4796_ ;
	wire _w4797_ ;
	wire _w4798_ ;
	wire _w4799_ ;
	wire _w4800_ ;
	wire _w4801_ ;
	wire _w4802_ ;
	wire _w4803_ ;
	wire _w4804_ ;
	wire _w4805_ ;
	wire _w4806_ ;
	wire _w4807_ ;
	wire _w4808_ ;
	wire _w4809_ ;
	wire _w4810_ ;
	wire _w4811_ ;
	wire _w4812_ ;
	wire _w4813_ ;
	wire _w4814_ ;
	wire _w4815_ ;
	wire _w4816_ ;
	wire _w4817_ ;
	wire _w4818_ ;
	wire _w4819_ ;
	wire _w4820_ ;
	wire _w4821_ ;
	wire _w4822_ ;
	wire _w4823_ ;
	wire _w4824_ ;
	wire _w4825_ ;
	wire _w4826_ ;
	wire _w4827_ ;
	wire _w4828_ ;
	wire _w4829_ ;
	wire _w4830_ ;
	wire _w4831_ ;
	wire _w4832_ ;
	wire _w4833_ ;
	wire _w4834_ ;
	wire _w4835_ ;
	wire _w4836_ ;
	wire _w4837_ ;
	wire _w4838_ ;
	wire _w4839_ ;
	wire _w4840_ ;
	wire _w4841_ ;
	wire _w4842_ ;
	wire _w4843_ ;
	wire _w4844_ ;
	wire _w4845_ ;
	wire _w4846_ ;
	wire _w4847_ ;
	wire _w4848_ ;
	wire _w4849_ ;
	wire _w4850_ ;
	wire _w4851_ ;
	wire _w4852_ ;
	wire _w4853_ ;
	wire _w4854_ ;
	wire _w4855_ ;
	wire _w4856_ ;
	wire _w4857_ ;
	wire _w4858_ ;
	wire _w4859_ ;
	wire _w4860_ ;
	wire _w4861_ ;
	wire _w4862_ ;
	wire _w4863_ ;
	wire _w4864_ ;
	wire _w4865_ ;
	wire _w4866_ ;
	wire _w4867_ ;
	wire _w4868_ ;
	wire _w4869_ ;
	wire _w4870_ ;
	wire _w4871_ ;
	wire _w4872_ ;
	wire _w4873_ ;
	wire _w4874_ ;
	wire _w4875_ ;
	wire _w4876_ ;
	wire _w4877_ ;
	wire _w4878_ ;
	wire _w4879_ ;
	wire _w4880_ ;
	wire _w4881_ ;
	wire _w4882_ ;
	wire _w4883_ ;
	wire _w4884_ ;
	wire _w4885_ ;
	wire _w4886_ ;
	wire _w4887_ ;
	wire _w4888_ ;
	wire _w4889_ ;
	wire _w4890_ ;
	wire _w4891_ ;
	wire _w4892_ ;
	wire _w4893_ ;
	wire _w4894_ ;
	wire _w4895_ ;
	wire _w4896_ ;
	wire _w4897_ ;
	wire _w4898_ ;
	wire _w4899_ ;
	wire _w4900_ ;
	wire _w4901_ ;
	wire _w4902_ ;
	wire _w4903_ ;
	wire _w4904_ ;
	wire _w4905_ ;
	wire _w4906_ ;
	wire _w4907_ ;
	wire _w4908_ ;
	wire _w4909_ ;
	wire _w4910_ ;
	wire _w4911_ ;
	wire _w4912_ ;
	wire _w4913_ ;
	wire _w4914_ ;
	wire _w4915_ ;
	wire _w4916_ ;
	wire _w4917_ ;
	wire _w4918_ ;
	wire _w4919_ ;
	wire _w4920_ ;
	wire _w4921_ ;
	wire _w4922_ ;
	wire _w4923_ ;
	wire _w4924_ ;
	wire _w4925_ ;
	wire _w4926_ ;
	wire _w4927_ ;
	wire _w4928_ ;
	wire _w4929_ ;
	wire _w4930_ ;
	wire _w4931_ ;
	wire _w4932_ ;
	wire _w4933_ ;
	wire _w4934_ ;
	wire _w4935_ ;
	wire _w4936_ ;
	wire _w4937_ ;
	wire _w4938_ ;
	wire _w4939_ ;
	wire _w4940_ ;
	wire _w4941_ ;
	wire _w4942_ ;
	wire _w4943_ ;
	wire _w4944_ ;
	wire _w4945_ ;
	wire _w4946_ ;
	wire _w4947_ ;
	wire _w4948_ ;
	wire _w4949_ ;
	wire _w4950_ ;
	wire _w4951_ ;
	wire _w4952_ ;
	wire _w4953_ ;
	wire _w4954_ ;
	wire _w4955_ ;
	wire _w4956_ ;
	wire _w4957_ ;
	wire _w4958_ ;
	wire _w4959_ ;
	wire _w4960_ ;
	wire _w4961_ ;
	wire _w4962_ ;
	wire _w4963_ ;
	wire _w4964_ ;
	wire _w4965_ ;
	wire _w4966_ ;
	wire _w4967_ ;
	wire _w4968_ ;
	wire _w4969_ ;
	wire _w4970_ ;
	wire _w4971_ ;
	wire _w4972_ ;
	wire _w4973_ ;
	wire _w4974_ ;
	wire _w4975_ ;
	wire _w4976_ ;
	wire _w4977_ ;
	wire _w4978_ ;
	wire _w4979_ ;
	wire _w4980_ ;
	wire _w4981_ ;
	wire _w4982_ ;
	wire _w4983_ ;
	wire _w4984_ ;
	wire _w4985_ ;
	wire _w4986_ ;
	wire _w4987_ ;
	wire _w4988_ ;
	wire _w4989_ ;
	wire _w4990_ ;
	wire _w4991_ ;
	wire _w4992_ ;
	wire _w4993_ ;
	wire _w4994_ ;
	wire _w4995_ ;
	wire _w4996_ ;
	wire _w4997_ ;
	wire _w4998_ ;
	wire _w4999_ ;
	wire _w5000_ ;
	wire _w5001_ ;
	wire _w5002_ ;
	wire _w5003_ ;
	wire _w5004_ ;
	wire _w5005_ ;
	wire _w5006_ ;
	wire _w5007_ ;
	wire _w5008_ ;
	wire _w5009_ ;
	wire _w5010_ ;
	wire _w5011_ ;
	wire _w5012_ ;
	wire _w5013_ ;
	wire _w5014_ ;
	wire _w5015_ ;
	wire _w5016_ ;
	wire _w5017_ ;
	wire _w5018_ ;
	wire _w5019_ ;
	wire _w5020_ ;
	wire _w5021_ ;
	wire _w5022_ ;
	wire _w5023_ ;
	wire _w5024_ ;
	wire _w5025_ ;
	wire _w5026_ ;
	wire _w5027_ ;
	wire _w5028_ ;
	wire _w5029_ ;
	wire _w5030_ ;
	wire _w5031_ ;
	wire _w5032_ ;
	wire _w5033_ ;
	wire _w5034_ ;
	wire _w5035_ ;
	wire _w5036_ ;
	wire _w5037_ ;
	wire _w5038_ ;
	wire _w5039_ ;
	wire _w5040_ ;
	wire _w5041_ ;
	wire _w5042_ ;
	wire _w5043_ ;
	wire _w5044_ ;
	wire _w5045_ ;
	wire _w5046_ ;
	wire _w5047_ ;
	wire _w5048_ ;
	wire _w5049_ ;
	wire _w5050_ ;
	wire _w5051_ ;
	wire _w5052_ ;
	wire _w5053_ ;
	wire _w5054_ ;
	wire _w5055_ ;
	wire _w5056_ ;
	wire _w5057_ ;
	wire _w5058_ ;
	wire _w5059_ ;
	wire _w5060_ ;
	wire _w5061_ ;
	wire _w5062_ ;
	wire _w5063_ ;
	wire _w5064_ ;
	wire _w5065_ ;
	wire _w5066_ ;
	wire _w5067_ ;
	wire _w5068_ ;
	wire _w5069_ ;
	wire _w5070_ ;
	wire _w5071_ ;
	wire _w5072_ ;
	wire _w5073_ ;
	wire _w5074_ ;
	wire _w5075_ ;
	wire _w5076_ ;
	wire _w5077_ ;
	wire _w5078_ ;
	wire _w5079_ ;
	wire _w5080_ ;
	wire _w5081_ ;
	wire _w5082_ ;
	wire _w5083_ ;
	wire _w5084_ ;
	wire _w5085_ ;
	wire _w5086_ ;
	wire _w5087_ ;
	wire _w5088_ ;
	wire _w5089_ ;
	wire _w5090_ ;
	wire _w5091_ ;
	wire _w5092_ ;
	wire _w5093_ ;
	wire _w5094_ ;
	wire _w5095_ ;
	wire _w5096_ ;
	wire _w5097_ ;
	wire _w5098_ ;
	wire _w5099_ ;
	wire _w5100_ ;
	wire _w5101_ ;
	wire _w5102_ ;
	wire _w5103_ ;
	wire _w5104_ ;
	wire _w5105_ ;
	wire _w5106_ ;
	wire _w5107_ ;
	wire _w5108_ ;
	wire _w5109_ ;
	wire _w5110_ ;
	wire _w5111_ ;
	wire _w5112_ ;
	wire _w5113_ ;
	wire _w5114_ ;
	wire _w5115_ ;
	wire _w5116_ ;
	wire _w5117_ ;
	wire _w5118_ ;
	wire _w5119_ ;
	wire _w5120_ ;
	wire _w5121_ ;
	wire _w5122_ ;
	wire _w5123_ ;
	wire _w5124_ ;
	wire _w5125_ ;
	wire _w5126_ ;
	wire _w5127_ ;
	wire _w5128_ ;
	wire _w5129_ ;
	wire _w5130_ ;
	wire _w5131_ ;
	wire _w5132_ ;
	wire _w5133_ ;
	wire _w5134_ ;
	wire _w5135_ ;
	wire _w5136_ ;
	wire _w5137_ ;
	wire _w5138_ ;
	wire _w5139_ ;
	wire _w5140_ ;
	wire _w5141_ ;
	wire _w5142_ ;
	wire _w5143_ ;
	wire _w5144_ ;
	wire _w5145_ ;
	wire _w5146_ ;
	wire _w5147_ ;
	wire _w5148_ ;
	wire _w5149_ ;
	wire _w5150_ ;
	wire _w5151_ ;
	wire _w5152_ ;
	wire _w5153_ ;
	wire _w5154_ ;
	wire _w5155_ ;
	wire _w5156_ ;
	wire _w5157_ ;
	wire _w5158_ ;
	wire _w5159_ ;
	wire _w5160_ ;
	wire _w5161_ ;
	wire _w5162_ ;
	wire _w5163_ ;
	wire _w5164_ ;
	wire _w5165_ ;
	wire _w5166_ ;
	wire _w5167_ ;
	wire _w5168_ ;
	wire _w5169_ ;
	wire _w5170_ ;
	wire _w5171_ ;
	wire _w5172_ ;
	wire _w5173_ ;
	wire _w5174_ ;
	wire _w5175_ ;
	wire _w5176_ ;
	wire _w5177_ ;
	wire _w5178_ ;
	wire _w5179_ ;
	wire _w5180_ ;
	wire _w5181_ ;
	wire _w5182_ ;
	wire _w5183_ ;
	wire _w5184_ ;
	wire _w5185_ ;
	wire _w5186_ ;
	wire _w5187_ ;
	wire _w5188_ ;
	wire _w5189_ ;
	wire _w5190_ ;
	wire _w5191_ ;
	wire _w5192_ ;
	wire _w5193_ ;
	wire _w5194_ ;
	wire _w5195_ ;
	wire _w5196_ ;
	wire _w5197_ ;
	wire _w5198_ ;
	wire _w5199_ ;
	wire _w5200_ ;
	wire _w5201_ ;
	wire _w5202_ ;
	wire _w5203_ ;
	wire _w5204_ ;
	wire _w5205_ ;
	wire _w5206_ ;
	wire _w5207_ ;
	wire _w5208_ ;
	wire _w5209_ ;
	wire _w5210_ ;
	wire _w5211_ ;
	wire _w5212_ ;
	wire _w5213_ ;
	wire _w5214_ ;
	wire _w5215_ ;
	wire _w5216_ ;
	wire _w5217_ ;
	wire _w5218_ ;
	wire _w5219_ ;
	wire _w5220_ ;
	wire _w5221_ ;
	wire _w5222_ ;
	wire _w5223_ ;
	wire _w5224_ ;
	wire _w5225_ ;
	wire _w5226_ ;
	wire _w5227_ ;
	wire _w5228_ ;
	wire _w5229_ ;
	wire _w5230_ ;
	wire _w5231_ ;
	wire _w5232_ ;
	wire _w5233_ ;
	wire _w5234_ ;
	wire _w5235_ ;
	wire _w5236_ ;
	wire _w5237_ ;
	wire _w5238_ ;
	wire _w5239_ ;
	wire _w5240_ ;
	wire _w5241_ ;
	wire _w5242_ ;
	wire _w5243_ ;
	wire _w5244_ ;
	wire _w5245_ ;
	wire _w5246_ ;
	wire _w5247_ ;
	wire _w5248_ ;
	wire _w5249_ ;
	wire _w5250_ ;
	wire _w5251_ ;
	wire _w5252_ ;
	wire _w5253_ ;
	wire _w5254_ ;
	wire _w5255_ ;
	wire _w5256_ ;
	wire _w5257_ ;
	wire _w5258_ ;
	wire _w5259_ ;
	wire _w5260_ ;
	wire _w5261_ ;
	wire _w5262_ ;
	wire _w5263_ ;
	wire _w5264_ ;
	wire _w5265_ ;
	wire _w5266_ ;
	wire _w5267_ ;
	wire _w5268_ ;
	wire _w5269_ ;
	wire _w5270_ ;
	wire _w5271_ ;
	wire _w5272_ ;
	wire _w5273_ ;
	wire _w5274_ ;
	wire _w5275_ ;
	wire _w5276_ ;
	wire _w5277_ ;
	wire _w5278_ ;
	wire _w5279_ ;
	wire _w5280_ ;
	wire _w5281_ ;
	wire _w5282_ ;
	wire _w5283_ ;
	wire _w5284_ ;
	wire _w5285_ ;
	wire _w5286_ ;
	wire _w5287_ ;
	wire _w5288_ ;
	wire _w5289_ ;
	wire _w5290_ ;
	wire _w5291_ ;
	wire _w5292_ ;
	wire _w5293_ ;
	wire _w5294_ ;
	wire _w5295_ ;
	wire _w5296_ ;
	wire _w5297_ ;
	wire _w5298_ ;
	wire _w5299_ ;
	wire _w5300_ ;
	wire _w5301_ ;
	wire _w5302_ ;
	wire _w5304_ ;
	wire _w5305_ ;
	wire _w5306_ ;
	wire _w5307_ ;
	wire _w5308_ ;
	wire _w5309_ ;
	wire _w5310_ ;
	wire _w5311_ ;
	wire _w5312_ ;
	wire _w5313_ ;
	wire _w5314_ ;
	wire _w5315_ ;
	wire _w5316_ ;
	wire _w5317_ ;
	wire _w5318_ ;
	wire _w5319_ ;
	wire _w5320_ ;
	wire _w5321_ ;
	wire _w5322_ ;
	wire _w5323_ ;
	wire _w5324_ ;
	wire _w5325_ ;
	wire _w5326_ ;
	wire _w5327_ ;
	wire _w5328_ ;
	wire _w5329_ ;
	wire _w5330_ ;
	wire _w5331_ ;
	wire _w5332_ ;
	wire _w5333_ ;
	wire _w5334_ ;
	wire _w5335_ ;
	wire _w5336_ ;
	wire _w5337_ ;
	wire _w5338_ ;
	wire _w5339_ ;
	wire _w5340_ ;
	wire _w5341_ ;
	wire _w5342_ ;
	wire _w5343_ ;
	wire _w5344_ ;
	wire _w5345_ ;
	wire _w5346_ ;
	wire _w5347_ ;
	wire _w5348_ ;
	wire _w5349_ ;
	wire _w5350_ ;
	wire _w5351_ ;
	wire _w5352_ ;
	wire _w5353_ ;
	wire _w5354_ ;
	wire _w5355_ ;
	wire _w5356_ ;
	wire _w5357_ ;
	wire _w5358_ ;
	wire _w5359_ ;
	wire _w5360_ ;
	wire _w5361_ ;
	wire _w5362_ ;
	wire _w5363_ ;
	wire _w5364_ ;
	wire _w5365_ ;
	wire _w5366_ ;
	wire _w5367_ ;
	wire _w5368_ ;
	wire _w5369_ ;
	wire _w5370_ ;
	wire _w5371_ ;
	wire _w5372_ ;
	wire _w5373_ ;
	wire _w5374_ ;
	wire _w5375_ ;
	wire _w5376_ ;
	wire _w5377_ ;
	wire _w5378_ ;
	wire _w5379_ ;
	wire _w5380_ ;
	wire _w5381_ ;
	wire _w5382_ ;
	wire _w5383_ ;
	wire _w5384_ ;
	wire _w5385_ ;
	wire _w5386_ ;
	wire _w5387_ ;
	wire _w5388_ ;
	wire _w5389_ ;
	wire _w5390_ ;
	wire _w5391_ ;
	wire _w5392_ ;
	wire _w5393_ ;
	wire _w5394_ ;
	wire _w5395_ ;
	wire _w5396_ ;
	wire _w5397_ ;
	wire _w5398_ ;
	wire _w5399_ ;
	wire _w5400_ ;
	wire _w5401_ ;
	wire _w5402_ ;
	wire _w5403_ ;
	wire _w5404_ ;
	wire _w5405_ ;
	wire _w5406_ ;
	wire _w5407_ ;
	wire _w5408_ ;
	wire _w5409_ ;
	wire _w5410_ ;
	wire _w5411_ ;
	wire _w5412_ ;
	wire _w5413_ ;
	wire _w5414_ ;
	wire _w5415_ ;
	wire _w5416_ ;
	wire _w5417_ ;
	wire _w5418_ ;
	wire _w5419_ ;
	wire _w5420_ ;
	wire _w5421_ ;
	wire _w5422_ ;
	wire _w5423_ ;
	wire _w5424_ ;
	wire _w5425_ ;
	wire _w5426_ ;
	wire _w5427_ ;
	wire _w5428_ ;
	wire _w5429_ ;
	wire _w5430_ ;
	wire _w5431_ ;
	wire _w5432_ ;
	wire _w5433_ ;
	wire _w5434_ ;
	wire _w5435_ ;
	wire _w5436_ ;
	wire _w5437_ ;
	wire _w5438_ ;
	wire _w5439_ ;
	wire _w5440_ ;
	wire _w5441_ ;
	wire _w5442_ ;
	wire _w5443_ ;
	wire _w5444_ ;
	wire _w5445_ ;
	wire _w5446_ ;
	wire _w5447_ ;
	wire _w5448_ ;
	wire _w5449_ ;
	wire _w5450_ ;
	wire _w5451_ ;
	wire _w5452_ ;
	wire _w5453_ ;
	wire _w5454_ ;
	wire _w5455_ ;
	wire _w5456_ ;
	wire _w5457_ ;
	wire _w5458_ ;
	wire _w5459_ ;
	wire _w5460_ ;
	wire _w5461_ ;
	wire _w5462_ ;
	wire _w5463_ ;
	wire _w5464_ ;
	wire _w5465_ ;
	wire _w5466_ ;
	wire _w5467_ ;
	wire _w5468_ ;
	wire _w5469_ ;
	wire _w5470_ ;
	wire _w5471_ ;
	wire _w5472_ ;
	wire _w5473_ ;
	wire _w5474_ ;
	wire _w5475_ ;
	wire _w5476_ ;
	wire _w5477_ ;
	wire _w5478_ ;
	wire _w5479_ ;
	wire _w5480_ ;
	wire _w5481_ ;
	wire _w5482_ ;
	wire _w5483_ ;
	wire _w5484_ ;
	wire _w5485_ ;
	wire _w5486_ ;
	wire _w5487_ ;
	wire _w5488_ ;
	wire _w5489_ ;
	wire _w5490_ ;
	wire _w5491_ ;
	wire _w5492_ ;
	wire _w5493_ ;
	wire _w5494_ ;
	wire _w5495_ ;
	wire _w5496_ ;
	wire _w5497_ ;
	wire _w5498_ ;
	wire _w5499_ ;
	wire _w5500_ ;
	wire _w5501_ ;
	wire _w5502_ ;
	wire _w5503_ ;
	wire _w5504_ ;
	wire _w5505_ ;
	wire _w5506_ ;
	wire _w5507_ ;
	wire _w5508_ ;
	wire _w5509_ ;
	wire _w5510_ ;
	wire _w5511_ ;
	wire _w5512_ ;
	wire _w5513_ ;
	wire _w5514_ ;
	wire _w5515_ ;
	wire _w5516_ ;
	wire _w5517_ ;
	wire _w5518_ ;
	wire _w5519_ ;
	wire _w5520_ ;
	wire _w5521_ ;
	wire _w5522_ ;
	wire _w5523_ ;
	wire _w5524_ ;
	wire _w5525_ ;
	wire _w5526_ ;
	wire _w5527_ ;
	wire _w5528_ ;
	wire _w5529_ ;
	wire _w5530_ ;
	wire _w5531_ ;
	wire _w5532_ ;
	wire _w5533_ ;
	wire _w5534_ ;
	wire _w5535_ ;
	wire _w5536_ ;
	wire _w5537_ ;
	wire _w5538_ ;
	wire _w5539_ ;
	wire _w5540_ ;
	wire _w5541_ ;
	wire _w5542_ ;
	wire _w5543_ ;
	wire _w5544_ ;
	wire _w5545_ ;
	wire _w5546_ ;
	wire _w5547_ ;
	wire _w5548_ ;
	wire _w5549_ ;
	LUT1 #(
		.INIT('h1)
	) name0 (
		\P1_state_reg[0]/NET0131 ,
		_w216_
	);
	LUT2 #(
		.INIT('h1)
	) name1 (
		\P1_IR_reg[6]/NET0131 ,
		\P1_IR_reg[7]/NET0131 ,
		_w464_
	);
	LUT4 #(
		.INIT('h0001)
	) name2 (
		\P1_IR_reg[0]/NET0131 ,
		\P1_IR_reg[1]/NET0131 ,
		\P1_IR_reg[2]/NET0131 ,
		\P1_IR_reg[3]/NET0131 ,
		_w465_
	);
	LUT2 #(
		.INIT('h1)
	) name3 (
		\P1_IR_reg[4]/NET0131 ,
		\P1_IR_reg[5]/NET0131 ,
		_w466_
	);
	LUT4 #(
		.INIT('h4000)
	) name4 (
		\P1_IR_reg[8]/NET0131 ,
		_w464_,
		_w465_,
		_w466_,
		_w467_
	);
	LUT2 #(
		.INIT('h1)
	) name5 (
		\P1_IR_reg[14]/NET0131 ,
		\P1_IR_reg[15]/NET0131 ,
		_w468_
	);
	LUT3 #(
		.INIT('h01)
	) name6 (
		\P1_IR_reg[14]/NET0131 ,
		\P1_IR_reg[15]/NET0131 ,
		\P1_IR_reg[16]/NET0131 ,
		_w469_
	);
	LUT4 #(
		.INIT('h0001)
	) name7 (
		\P1_IR_reg[10]/NET0131 ,
		\P1_IR_reg[11]/NET0131 ,
		\P1_IR_reg[12]/NET0131 ,
		\P1_IR_reg[13]/NET0131 ,
		_w470_
	);
	LUT3 #(
		.INIT('h40)
	) name8 (
		\P1_IR_reg[9]/NET0131 ,
		_w470_,
		_w469_,
		_w471_
	);
	LUT4 #(
		.INIT('h0001)
	) name9 (
		\P1_IR_reg[17]/NET0131 ,
		\P1_IR_reg[18]/NET0131 ,
		\P1_IR_reg[19]/NET0131 ,
		\P1_IR_reg[20]/NET0131 ,
		_w472_
	);
	LUT4 #(
		.INIT('h0001)
	) name10 (
		\P1_IR_reg[21]/NET0131 ,
		\P1_IR_reg[22]/NET0131 ,
		\P1_IR_reg[23]/NET0131 ,
		\P1_IR_reg[24]/NET0131 ,
		_w473_
	);
	LUT2 #(
		.INIT('h8)
	) name11 (
		_w472_,
		_w473_,
		_w474_
	);
	LUT4 #(
		.INIT('h2aaa)
	) name12 (
		\P1_IR_reg[31]/NET0131 ,
		_w467_,
		_w471_,
		_w474_,
		_w475_
	);
	LUT4 #(
		.INIT('h0001)
	) name13 (
		\P1_IR_reg[25]/NET0131 ,
		\P1_IR_reg[26]/NET0131 ,
		\P1_IR_reg[27]/NET0131 ,
		\P1_IR_reg[28]/NET0131 ,
		_w476_
	);
	LUT2 #(
		.INIT('h2)
	) name14 (
		\P1_IR_reg[31]/NET0131 ,
		_w476_,
		_w477_
	);
	LUT3 #(
		.INIT('h56)
	) name15 (
		\P1_IR_reg[29]/NET0131 ,
		_w475_,
		_w477_,
		_w478_
	);
	LUT4 #(
		.INIT('h0001)
	) name16 (
		\P1_IR_reg[6]/NET0131 ,
		\P1_IR_reg[7]/NET0131 ,
		\P1_IR_reg[8]/NET0131 ,
		\P1_IR_reg[9]/NET0131 ,
		_w479_
	);
	LUT4 #(
		.INIT('h8000)
	) name17 (
		_w465_,
		_w466_,
		_w470_,
		_w479_,
		_w480_
	);
	LUT4 #(
		.INIT('h0001)
	) name18 (
		\P1_IR_reg[14]/NET0131 ,
		\P1_IR_reg[15]/NET0131 ,
		\P1_IR_reg[16]/NET0131 ,
		\P1_IR_reg[21]/NET0131 ,
		_w481_
	);
	LUT2 #(
		.INIT('h8)
	) name19 (
		_w472_,
		_w481_,
		_w482_
	);
	LUT4 #(
		.INIT('h0001)
	) name20 (
		\P1_IR_reg[22]/NET0131 ,
		\P1_IR_reg[23]/NET0131 ,
		\P1_IR_reg[24]/NET0131 ,
		\P1_IR_reg[25]/NET0131 ,
		_w483_
	);
	LUT4 #(
		.INIT('h2aaa)
	) name21 (
		\P1_IR_reg[31]/NET0131 ,
		_w480_,
		_w482_,
		_w483_,
		_w484_
	);
	LUT3 #(
		.INIT('h01)
	) name22 (
		\P1_IR_reg[27]/NET0131 ,
		\P1_IR_reg[28]/NET0131 ,
		\P1_IR_reg[29]/NET0131 ,
		_w485_
	);
	LUT4 #(
		.INIT('h0001)
	) name23 (
		\P1_IR_reg[26]/NET0131 ,
		\P1_IR_reg[27]/NET0131 ,
		\P1_IR_reg[28]/NET0131 ,
		\P1_IR_reg[29]/NET0131 ,
		_w486_
	);
	LUT2 #(
		.INIT('h2)
	) name24 (
		\P1_IR_reg[31]/NET0131 ,
		_w486_,
		_w487_
	);
	LUT3 #(
		.INIT('h56)
	) name25 (
		\P1_IR_reg[30]/NET0131 ,
		_w484_,
		_w487_,
		_w488_
	);
	LUT4 #(
		.INIT('hf35f)
	) name26 (
		\P1_reg1_reg[3]/NET0131 ,
		\P1_reg2_reg[3]/NET0131 ,
		_w478_,
		_w488_,
		_w489_
	);
	LUT2 #(
		.INIT('h8)
	) name27 (
		_w478_,
		_w488_,
		_w490_
	);
	LUT4 #(
		.INIT('hcff5)
	) name28 (
		\P1_reg0_reg[3]/NET0131 ,
		\P1_reg3_reg[3]/NET0131 ,
		_w478_,
		_w488_,
		_w491_
	);
	LUT2 #(
		.INIT('h8)
	) name29 (
		_w489_,
		_w491_,
		_w492_
	);
	LUT2 #(
		.INIT('h7)
	) name30 (
		_w489_,
		_w491_,
		_w493_
	);
	LUT4 #(
		.INIT('h0001)
	) name31 (
		\P2_IR_reg[10]/NET0131 ,
		\P2_IR_reg[11]/NET0131 ,
		\P2_IR_reg[12]/NET0131 ,
		\P2_IR_reg[9]/NET0131 ,
		_w494_
	);
	LUT2 #(
		.INIT('h1)
	) name32 (
		\P2_IR_reg[7]/NET0131 ,
		\P2_IR_reg[8]/NET0131 ,
		_w495_
	);
	LUT4 #(
		.INIT('h0001)
	) name33 (
		\P2_IR_reg[0]/NET0131 ,
		\P2_IR_reg[1]/NET0131 ,
		\P2_IR_reg[2]/NET0131 ,
		\P2_IR_reg[3]/NET0131 ,
		_w496_
	);
	LUT3 #(
		.INIT('h01)
	) name34 (
		\P2_IR_reg[4]/NET0131 ,
		\P2_IR_reg[5]/NET0131 ,
		\P2_IR_reg[6]/NET0131 ,
		_w497_
	);
	LUT4 #(
		.INIT('h8000)
	) name35 (
		_w494_,
		_w495_,
		_w496_,
		_w497_,
		_w498_
	);
	LUT2 #(
		.INIT('h1)
	) name36 (
		\P2_IR_reg[14]/NET0131 ,
		\P2_IR_reg[15]/NET0131 ,
		_w499_
	);
	LUT4 #(
		.INIT('h0001)
	) name37 (
		\P2_IR_reg[13]/NET0131 ,
		\P2_IR_reg[14]/NET0131 ,
		\P2_IR_reg[15]/NET0131 ,
		\P2_IR_reg[16]/NET0131 ,
		_w500_
	);
	LUT4 #(
		.INIT('h0001)
	) name38 (
		\P2_IR_reg[17]/NET0131 ,
		\P2_IR_reg[18]/NET0131 ,
		\P2_IR_reg[19]/NET0131 ,
		\P2_IR_reg[20]/NET0131 ,
		_w501_
	);
	LUT4 #(
		.INIT('h0001)
	) name39 (
		\P2_IR_reg[21]/NET0131 ,
		\P2_IR_reg[22]/NET0131 ,
		\P2_IR_reg[23]/NET0131 ,
		\P2_IR_reg[24]/NET0131 ,
		_w502_
	);
	LUT4 #(
		.INIT('h0001)
	) name40 (
		\P2_IR_reg[25]/NET0131 ,
		\P2_IR_reg[26]/NET0131 ,
		\P2_IR_reg[27]/NET0131 ,
		\P2_IR_reg[28]/NET0131 ,
		_w503_
	);
	LUT4 #(
		.INIT('h8000)
	) name41 (
		_w500_,
		_w501_,
		_w502_,
		_w503_,
		_w504_
	);
	LUT4 #(
		.INIT('ha666)
	) name42 (
		\P2_IR_reg[29]/NET0131 ,
		\P2_IR_reg[31]/NET0131 ,
		_w498_,
		_w504_,
		_w505_
	);
	LUT3 #(
		.INIT('h40)
	) name43 (
		\P2_IR_reg[7]/NET0131 ,
		_w496_,
		_w497_,
		_w506_
	);
	LUT2 #(
		.INIT('h1)
	) name44 (
		\P2_IR_reg[13]/NET0131 ,
		\P2_IR_reg[8]/NET0131 ,
		_w507_
	);
	LUT2 #(
		.INIT('h8)
	) name45 (
		_w494_,
		_w507_,
		_w508_
	);
	LUT4 #(
		.INIT('h0001)
	) name46 (
		\P2_IR_reg[14]/NET0131 ,
		\P2_IR_reg[15]/NET0131 ,
		\P2_IR_reg[16]/NET0131 ,
		\P2_IR_reg[17]/NET0131 ,
		_w509_
	);
	LUT4 #(
		.INIT('h0001)
	) name47 (
		\P2_IR_reg[18]/NET0131 ,
		\P2_IR_reg[19]/NET0131 ,
		\P2_IR_reg[20]/NET0131 ,
		\P2_IR_reg[21]/NET0131 ,
		_w510_
	);
	LUT2 #(
		.INIT('h8)
	) name48 (
		_w509_,
		_w510_,
		_w511_
	);
	LUT4 #(
		.INIT('h0001)
	) name49 (
		\P2_IR_reg[22]/NET0131 ,
		\P2_IR_reg[23]/NET0131 ,
		\P2_IR_reg[24]/NET0131 ,
		\P2_IR_reg[25]/NET0131 ,
		_w512_
	);
	LUT2 #(
		.INIT('h1)
	) name50 (
		\P2_IR_reg[28]/NET0131 ,
		\P2_IR_reg[29]/NET0131 ,
		_w513_
	);
	LUT4 #(
		.INIT('h0001)
	) name51 (
		\P2_IR_reg[26]/NET0131 ,
		\P2_IR_reg[27]/NET0131 ,
		\P2_IR_reg[28]/NET0131 ,
		\P2_IR_reg[29]/NET0131 ,
		_w514_
	);
	LUT4 #(
		.INIT('h8000)
	) name52 (
		_w509_,
		_w510_,
		_w512_,
		_w514_,
		_w515_
	);
	LUT4 #(
		.INIT('hd555)
	) name53 (
		\P2_IR_reg[31]/NET0131 ,
		_w506_,
		_w508_,
		_w515_,
		_w516_
	);
	LUT4 #(
		.INIT('h4080)
	) name54 (
		\P2_IR_reg[30]/NET0131 ,
		\P2_reg1_reg[15]/NET0131 ,
		_w505_,
		_w516_,
		_w517_
	);
	LUT4 #(
		.INIT('h0408)
	) name55 (
		\P2_IR_reg[30]/NET0131 ,
		\P2_reg0_reg[15]/NET0131 ,
		_w505_,
		_w516_,
		_w518_
	);
	LUT3 #(
		.INIT('h84)
	) name56 (
		\P2_IR_reg[30]/NET0131 ,
		_w505_,
		_w516_,
		_w519_
	);
	LUT4 #(
		.INIT('h0001)
	) name57 (
		\P2_reg3_reg[3]/NET0131 ,
		\P2_reg3_reg[4]/NET0131 ,
		\P2_reg3_reg[5]/NET0131 ,
		\P2_reg3_reg[6]/NET0131 ,
		_w520_
	);
	LUT2 #(
		.INIT('h1)
	) name58 (
		\P2_reg3_reg[8]/NET0131 ,
		\P2_reg3_reg[9]/NET0131 ,
		_w521_
	);
	LUT4 #(
		.INIT('h1000)
	) name59 (
		\P2_reg3_reg[10]/NET0131 ,
		\P2_reg3_reg[7]/NET0131 ,
		_w520_,
		_w521_,
		_w522_
	);
	LUT4 #(
		.INIT('h0001)
	) name60 (
		\P2_reg3_reg[11]/NET0131 ,
		\P2_reg3_reg[12]/NET0131 ,
		\P2_reg3_reg[13]/NET0131 ,
		\P2_reg3_reg[14]/NET0131 ,
		_w523_
	);
	LUT2 #(
		.INIT('h8)
	) name61 (
		_w522_,
		_w523_,
		_w524_
	);
	LUT3 #(
		.INIT('h95)
	) name62 (
		\P2_reg3_reg[15]/NET0131 ,
		_w522_,
		_w523_,
		_w525_
	);
	LUT4 #(
		.INIT('h0084)
	) name63 (
		\P2_IR_reg[30]/NET0131 ,
		_w505_,
		_w516_,
		_w525_,
		_w526_
	);
	LUT4 #(
		.INIT('h0804)
	) name64 (
		\P2_IR_reg[30]/NET0131 ,
		\P2_reg2_reg[15]/NET0131 ,
		_w505_,
		_w516_,
		_w527_
	);
	LUT4 #(
		.INIT('h0001)
	) name65 (
		_w517_,
		_w518_,
		_w526_,
		_w527_,
		_w528_
	);
	LUT4 #(
		.INIT('hfffe)
	) name66 (
		_w517_,
		_w518_,
		_w526_,
		_w527_,
		_w529_
	);
	LUT3 #(
		.INIT('h80)
	) name67 (
		_w494_,
		_w499_,
		_w507_,
		_w530_
	);
	LUT4 #(
		.INIT('h0001)
	) name68 (
		\P2_IR_reg[19]/NET0131 ,
		\P2_IR_reg[20]/NET0131 ,
		\P2_IR_reg[21]/NET0131 ,
		\P2_IR_reg[22]/NET0131 ,
		_w531_
	);
	LUT4 #(
		.INIT('h0001)
	) name69 (
		\P2_IR_reg[16]/NET0131 ,
		\P2_IR_reg[17]/NET0131 ,
		\P2_IR_reg[18]/NET0131 ,
		\P2_IR_reg[23]/NET0131 ,
		_w532_
	);
	LUT2 #(
		.INIT('h8)
	) name70 (
		_w531_,
		_w532_,
		_w533_
	);
	LUT4 #(
		.INIT('h2aaa)
	) name71 (
		\P2_IR_reg[31]/NET0131 ,
		_w506_,
		_w530_,
		_w533_,
		_w534_
	);
	LUT4 #(
		.INIT('h0001)
	) name72 (
		\P2_IR_reg[24]/NET0131 ,
		\P2_IR_reg[25]/NET0131 ,
		\P2_IR_reg[26]/NET0131 ,
		\P2_IR_reg[27]/NET0131 ,
		_w535_
	);
	LUT2 #(
		.INIT('h2)
	) name73 (
		\P2_IR_reg[31]/NET0131 ,
		_w535_,
		_w536_
	);
	LUT3 #(
		.INIT('h56)
	) name74 (
		\P2_IR_reg[28]/NET0131 ,
		_w534_,
		_w536_,
		_w537_
	);
	LUT4 #(
		.INIT('h0001)
	) name75 (
		\P2_IR_reg[10]/NET0131 ,
		\P2_IR_reg[7]/NET0131 ,
		\P2_IR_reg[8]/NET0131 ,
		\P2_IR_reg[9]/NET0131 ,
		_w538_
	);
	LUT4 #(
		.INIT('h0001)
	) name76 (
		\P2_IR_reg[11]/NET0131 ,
		\P2_IR_reg[12]/NET0131 ,
		\P2_IR_reg[13]/NET0131 ,
		\P2_IR_reg[14]/NET0131 ,
		_w539_
	);
	LUT4 #(
		.INIT('h8000)
	) name77 (
		_w496_,
		_w497_,
		_w538_,
		_w539_,
		_w540_
	);
	LUT4 #(
		.INIT('h0001)
	) name78 (
		\P2_IR_reg[15]/NET0131 ,
		\P2_IR_reg[16]/NET0131 ,
		\P2_IR_reg[17]/NET0131 ,
		\P2_IR_reg[18]/NET0131 ,
		_w541_
	);
	LUT4 #(
		.INIT('h0001)
	) name79 (
		\P2_IR_reg[23]/NET0131 ,
		\P2_IR_reg[24]/NET0131 ,
		\P2_IR_reg[25]/NET0131 ,
		\P2_IR_reg[26]/NET0131 ,
		_w542_
	);
	LUT3 #(
		.INIT('h2a)
	) name80 (
		\P2_IR_reg[31]/NET0131 ,
		_w531_,
		_w542_,
		_w543_
	);
	LUT4 #(
		.INIT('h00d5)
	) name81 (
		\P2_IR_reg[31]/NET0131 ,
		_w540_,
		_w541_,
		_w543_,
		_w544_
	);
	LUT2 #(
		.INIT('h9)
	) name82 (
		\P2_IR_reg[27]/NET0131 ,
		_w544_,
		_w545_
	);
	LUT2 #(
		.INIT('h1)
	) name83 (
		_w537_,
		_w545_,
		_w546_
	);
	LUT4 #(
		.INIT('hfe5e)
	) name84 (
		\P1_addr_reg[19]/NET0131 ,
		\P1_rd_reg/NET0131 ,
		\P2_addr_reg[19]/NET0131 ,
		\P2_rd_reg/NET0131 ,
		_w547_
	);
	LUT2 #(
		.INIT('h2)
	) name85 (
		\P1_datao_reg[15]/NET0131 ,
		_w547_,
		_w548_
	);
	LUT2 #(
		.INIT('h1)
	) name86 (
		\P1_datao_reg[6]/NET0131 ,
		\si[6]_pad ,
		_w549_
	);
	LUT2 #(
		.INIT('h8)
	) name87 (
		\P1_datao_reg[6]/NET0131 ,
		\si[6]_pad ,
		_w550_
	);
	LUT4 #(
		.INIT('hec80)
	) name88 (
		\P1_datao_reg[5]/NET0131 ,
		\P1_datao_reg[6]/NET0131 ,
		\si[5]_pad ,
		\si[6]_pad ,
		_w551_
	);
	LUT2 #(
		.INIT('h1)
	) name89 (
		\P1_datao_reg[3]/NET0131 ,
		\si[3]_pad ,
		_w552_
	);
	LUT2 #(
		.INIT('h1)
	) name90 (
		\P1_datao_reg[2]/NET0131 ,
		\si[2]_pad ,
		_w553_
	);
	LUT2 #(
		.INIT('h8)
	) name91 (
		\P1_datao_reg[0]/NET0131 ,
		\si[0]_pad ,
		_w554_
	);
	LUT4 #(
		.INIT('ha080)
	) name92 (
		\P1_datao_reg[0]/NET0131 ,
		\P1_datao_reg[1]/NET0131 ,
		\si[0]_pad ,
		\si[1]_pad ,
		_w555_
	);
	LUT4 #(
		.INIT('h135f)
	) name93 (
		\P1_datao_reg[1]/NET0131 ,
		\P1_datao_reg[2]/NET0131 ,
		\si[1]_pad ,
		\si[2]_pad ,
		_w556_
	);
	LUT3 #(
		.INIT('h45)
	) name94 (
		_w553_,
		_w555_,
		_w556_,
		_w557_
	);
	LUT4 #(
		.INIT('h1011)
	) name95 (
		_w552_,
		_w553_,
		_w555_,
		_w556_,
		_w558_
	);
	LUT4 #(
		.INIT('h135f)
	) name96 (
		\P1_datao_reg[3]/NET0131 ,
		\P1_datao_reg[4]/NET0131 ,
		\si[3]_pad ,
		\si[4]_pad ,
		_w559_
	);
	LUT2 #(
		.INIT('h1)
	) name97 (
		\P1_datao_reg[4]/NET0131 ,
		\si[4]_pad ,
		_w560_
	);
	LUT4 #(
		.INIT('hfac8)
	) name98 (
		\P1_datao_reg[4]/NET0131 ,
		\P1_datao_reg[5]/NET0131 ,
		\si[4]_pad ,
		\si[5]_pad ,
		_w561_
	);
	LUT2 #(
		.INIT('h4)
	) name99 (
		_w549_,
		_w561_,
		_w562_
	);
	LUT4 #(
		.INIT('h1055)
	) name100 (
		_w551_,
		_w558_,
		_w559_,
		_w562_,
		_w563_
	);
	LUT2 #(
		.INIT('h1)
	) name101 (
		\P1_datao_reg[8]/NET0131 ,
		\si[8]_pad ,
		_w564_
	);
	LUT2 #(
		.INIT('h1)
	) name102 (
		\P1_datao_reg[9]/NET0131 ,
		\si[9]_pad ,
		_w565_
	);
	LUT4 #(
		.INIT('hfac8)
	) name103 (
		\P1_datao_reg[10]/NET0131 ,
		\P1_datao_reg[9]/NET0131 ,
		\si[10]_pad ,
		\si[9]_pad ,
		_w566_
	);
	LUT2 #(
		.INIT('h1)
	) name104 (
		\P1_datao_reg[7]/NET0131 ,
		\si[7]_pad ,
		_w567_
	);
	LUT3 #(
		.INIT('h04)
	) name105 (
		_w564_,
		_w566_,
		_w567_,
		_w568_
	);
	LUT2 #(
		.INIT('h8)
	) name106 (
		\P1_datao_reg[10]/NET0131 ,
		\si[10]_pad ,
		_w569_
	);
	LUT4 #(
		.INIT('he8a0)
	) name107 (
		\P1_datao_reg[10]/NET0131 ,
		\P1_datao_reg[9]/NET0131 ,
		\si[10]_pad ,
		\si[9]_pad ,
		_w570_
	);
	LUT2 #(
		.INIT('h8)
	) name108 (
		\P1_datao_reg[8]/NET0131 ,
		\si[8]_pad ,
		_w571_
	);
	LUT2 #(
		.INIT('h8)
	) name109 (
		\P1_datao_reg[7]/NET0131 ,
		\si[7]_pad ,
		_w572_
	);
	LUT4 #(
		.INIT('h135f)
	) name110 (
		\P1_datao_reg[7]/NET0131 ,
		\P1_datao_reg[8]/NET0131 ,
		\si[7]_pad ,
		\si[8]_pad ,
		_w573_
	);
	LUT4 #(
		.INIT('h5545)
	) name111 (
		_w570_,
		_w564_,
		_w566_,
		_w573_,
		_w574_
	);
	LUT3 #(
		.INIT('hb0)
	) name112 (
		_w563_,
		_w568_,
		_w574_,
		_w575_
	);
	LUT2 #(
		.INIT('h1)
	) name113 (
		\P1_datao_reg[12]/NET0131 ,
		\si[12]_pad ,
		_w576_
	);
	LUT2 #(
		.INIT('h1)
	) name114 (
		\P1_datao_reg[11]/NET0131 ,
		\si[11]_pad ,
		_w577_
	);
	LUT4 #(
		.INIT('hfac8)
	) name115 (
		\P1_datao_reg[11]/NET0131 ,
		\P1_datao_reg[12]/NET0131 ,
		\si[11]_pad ,
		\si[12]_pad ,
		_w578_
	);
	LUT2 #(
		.INIT('h1)
	) name116 (
		\P1_datao_reg[13]/NET0131 ,
		\si[13]_pad ,
		_w579_
	);
	LUT4 #(
		.INIT('hfac8)
	) name117 (
		\P1_datao_reg[13]/NET0131 ,
		\P1_datao_reg[14]/NET0131 ,
		\si[13]_pad ,
		\si[14]_pad ,
		_w580_
	);
	LUT2 #(
		.INIT('h8)
	) name118 (
		_w578_,
		_w580_,
		_w581_
	);
	LUT4 #(
		.INIT('h4f00)
	) name119 (
		_w563_,
		_w568_,
		_w574_,
		_w581_,
		_w582_
	);
	LUT4 #(
		.INIT('hec80)
	) name120 (
		\P1_datao_reg[13]/NET0131 ,
		\P1_datao_reg[14]/NET0131 ,
		\si[13]_pad ,
		\si[14]_pad ,
		_w583_
	);
	LUT2 #(
		.INIT('h8)
	) name121 (
		\P1_datao_reg[12]/NET0131 ,
		\si[12]_pad ,
		_w584_
	);
	LUT2 #(
		.INIT('h8)
	) name122 (
		\P1_datao_reg[11]/NET0131 ,
		\si[11]_pad ,
		_w585_
	);
	LUT4 #(
		.INIT('h135f)
	) name123 (
		\P1_datao_reg[11]/NET0131 ,
		\P1_datao_reg[12]/NET0131 ,
		\si[11]_pad ,
		\si[12]_pad ,
		_w586_
	);
	LUT4 #(
		.INIT('h0f0b)
	) name124 (
		_w576_,
		_w580_,
		_w583_,
		_w586_,
		_w587_
	);
	LUT2 #(
		.INIT('h1)
	) name125 (
		\P1_datao_reg[15]/NET0131 ,
		\si[15]_pad ,
		_w588_
	);
	LUT2 #(
		.INIT('h8)
	) name126 (
		\P1_datao_reg[15]/NET0131 ,
		\si[15]_pad ,
		_w589_
	);
	LUT2 #(
		.INIT('h6)
	) name127 (
		\P1_datao_reg[15]/NET0131 ,
		\si[15]_pad ,
		_w590_
	);
	LUT4 #(
		.INIT('h208a)
	) name128 (
		_w547_,
		_w582_,
		_w587_,
		_w590_,
		_w591_
	);
	LUT3 #(
		.INIT('ha6)
	) name129 (
		\P2_IR_reg[15]/NET0131 ,
		\P2_IR_reg[31]/NET0131 ,
		_w540_,
		_w592_
	);
	LUT3 #(
		.INIT('h10)
	) name130 (
		_w537_,
		_w545_,
		_w592_,
		_w593_
	);
	LUT4 #(
		.INIT('h00ab)
	) name131 (
		_w546_,
		_w548_,
		_w591_,
		_w593_,
		_w594_
	);
	LUT4 #(
		.INIT('h135f)
	) name132 (
		\P1_datao_reg[12]/NET0131 ,
		\P1_datao_reg[13]/NET0131 ,
		\si[12]_pad ,
		\si[13]_pad ,
		_w595_
	);
	LUT4 #(
		.INIT('h135f)
	) name133 (
		\P1_datao_reg[10]/NET0131 ,
		\P1_datao_reg[11]/NET0131 ,
		\si[10]_pad ,
		\si[11]_pad ,
		_w596_
	);
	LUT4 #(
		.INIT('h0323)
	) name134 (
		_w578_,
		_w579_,
		_w595_,
		_w596_,
		_w597_
	);
	LUT4 #(
		.INIT('h137f)
	) name135 (
		\P1_datao_reg[0]/NET0131 ,
		\P1_datao_reg[1]/NET0131 ,
		\si[0]_pad ,
		\si[1]_pad ,
		_w598_
	);
	LUT4 #(
		.INIT('h135f)
	) name136 (
		\P1_datao_reg[2]/NET0131 ,
		\P1_datao_reg[3]/NET0131 ,
		\si[2]_pad ,
		\si[3]_pad ,
		_w599_
	);
	LUT4 #(
		.INIT('h0155)
	) name137 (
		_w552_,
		_w553_,
		_w598_,
		_w599_,
		_w600_
	);
	LUT4 #(
		.INIT('hec80)
	) name138 (
		\P1_datao_reg[4]/NET0131 ,
		\P1_datao_reg[5]/NET0131 ,
		\si[4]_pad ,
		\si[5]_pad ,
		_w601_
	);
	LUT3 #(
		.INIT('h07)
	) name139 (
		_w561_,
		_w600_,
		_w601_,
		_w602_
	);
	LUT4 #(
		.INIT('hfac8)
	) name140 (
		\P1_datao_reg[7]/NET0131 ,
		\P1_datao_reg[8]/NET0131 ,
		\si[7]_pad ,
		\si[8]_pad ,
		_w603_
	);
	LUT3 #(
		.INIT('h10)
	) name141 (
		_w565_,
		_w549_,
		_w603_,
		_w604_
	);
	LUT4 #(
		.INIT('hf800)
	) name142 (
		_w561_,
		_w600_,
		_w601_,
		_w604_,
		_w605_
	);
	LUT4 #(
		.INIT('hec80)
	) name143 (
		\P1_datao_reg[8]/NET0131 ,
		\P1_datao_reg[9]/NET0131 ,
		\si[8]_pad ,
		\si[9]_pad ,
		_w606_
	);
	LUT4 #(
		.INIT('h135f)
	) name144 (
		\P1_datao_reg[6]/NET0131 ,
		\P1_datao_reg[7]/NET0131 ,
		\si[6]_pad ,
		\si[7]_pad ,
		_w607_
	);
	LUT4 #(
		.INIT('h0f0b)
	) name145 (
		_w565_,
		_w603_,
		_w606_,
		_w607_,
		_w608_
	);
	LUT4 #(
		.INIT('hfac8)
	) name146 (
		\P1_datao_reg[10]/NET0131 ,
		\P1_datao_reg[13]/NET0131 ,
		\si[10]_pad ,
		\si[13]_pad ,
		_w609_
	);
	LUT2 #(
		.INIT('h8)
	) name147 (
		_w578_,
		_w609_,
		_w610_
	);
	LUT4 #(
		.INIT('h1055)
	) name148 (
		_w597_,
		_w605_,
		_w608_,
		_w610_,
		_w611_
	);
	LUT4 #(
		.INIT('h9565)
	) name149 (
		\P1_datao_reg[14]/NET0131 ,
		\si[14]_pad ,
		_w547_,
		_w611_,
		_w612_
	);
	LUT4 #(
		.INIT('ha666)
	) name150 (
		\P2_IR_reg[14]/NET0131 ,
		\P2_IR_reg[31]/NET0131 ,
		_w506_,
		_w508_,
		_w613_
	);
	LUT3 #(
		.INIT('h10)
	) name151 (
		_w537_,
		_w545_,
		_w613_,
		_w614_
	);
	LUT3 #(
		.INIT('h0e)
	) name152 (
		_w546_,
		_w612_,
		_w614_,
		_w615_
	);
	LUT4 #(
		.INIT('h0804)
	) name153 (
		\P2_IR_reg[30]/NET0131 ,
		\P2_reg2_reg[14]/NET0131 ,
		_w505_,
		_w516_,
		_w616_
	);
	LUT4 #(
		.INIT('h0408)
	) name154 (
		\P2_IR_reg[30]/NET0131 ,
		\P2_reg0_reg[14]/NET0131 ,
		_w505_,
		_w516_,
		_w617_
	);
	LUT2 #(
		.INIT('h1)
	) name155 (
		_w616_,
		_w617_,
		_w618_
	);
	LUT4 #(
		.INIT('h0100)
	) name156 (
		\P2_reg3_reg[11]/NET0131 ,
		\P2_reg3_reg[12]/NET0131 ,
		\P2_reg3_reg[13]/NET0131 ,
		_w522_,
		_w619_
	);
	LUT3 #(
		.INIT('h31)
	) name157 (
		\P2_reg3_reg[14]/NET0131 ,
		_w524_,
		_w619_,
		_w620_
	);
	LUT4 #(
		.INIT('h4080)
	) name158 (
		\P2_IR_reg[30]/NET0131 ,
		\P2_reg1_reg[14]/NET0131 ,
		_w505_,
		_w516_,
		_w621_
	);
	LUT3 #(
		.INIT('h0d)
	) name159 (
		_w519_,
		_w620_,
		_w621_,
		_w622_
	);
	LUT2 #(
		.INIT('h8)
	) name160 (
		_w618_,
		_w622_,
		_w623_
	);
	LUT2 #(
		.INIT('h7)
	) name161 (
		_w618_,
		_w622_,
		_w624_
	);
	LUT4 #(
		.INIT('hd0dd)
	) name162 (
		_w528_,
		_w594_,
		_w615_,
		_w623_,
		_w625_
	);
	LUT4 #(
		.INIT('h4080)
	) name163 (
		\P2_IR_reg[30]/NET0131 ,
		\P2_reg1_reg[13]/NET0131 ,
		_w505_,
		_w516_,
		_w626_
	);
	LUT4 #(
		.INIT('h1e0f)
	) name164 (
		\P2_reg3_reg[11]/NET0131 ,
		\P2_reg3_reg[12]/NET0131 ,
		\P2_reg3_reg[13]/NET0131 ,
		_w522_,
		_w627_
	);
	LUT4 #(
		.INIT('h0084)
	) name165 (
		\P2_IR_reg[30]/NET0131 ,
		_w505_,
		_w516_,
		_w627_,
		_w628_
	);
	LUT4 #(
		.INIT('h0408)
	) name166 (
		\P2_IR_reg[30]/NET0131 ,
		\P2_reg0_reg[13]/NET0131 ,
		_w505_,
		_w516_,
		_w629_
	);
	LUT4 #(
		.INIT('h0804)
	) name167 (
		\P2_IR_reg[30]/NET0131 ,
		\P2_reg2_reg[13]/NET0131 ,
		_w505_,
		_w516_,
		_w630_
	);
	LUT4 #(
		.INIT('h0001)
	) name168 (
		_w626_,
		_w628_,
		_w629_,
		_w630_,
		_w631_
	);
	LUT4 #(
		.INIT('hfffe)
	) name169 (
		_w626_,
		_w628_,
		_w629_,
		_w630_,
		_w632_
	);
	LUT3 #(
		.INIT('h0b)
	) name170 (
		_w558_,
		_w559_,
		_w560_,
		_w633_
	);
	LUT4 #(
		.INIT('hfac8)
	) name171 (
		\P1_datao_reg[6]/NET0131 ,
		\P1_datao_reg[7]/NET0131 ,
		\si[6]_pad ,
		\si[7]_pad ,
		_w634_
	);
	LUT4 #(
		.INIT('hfac8)
	) name172 (
		\P1_datao_reg[5]/NET0131 ,
		\P1_datao_reg[8]/NET0131 ,
		\si[5]_pad ,
		\si[8]_pad ,
		_w635_
	);
	LUT2 #(
		.INIT('h8)
	) name173 (
		_w634_,
		_w635_,
		_w636_
	);
	LUT4 #(
		.INIT('h0b00)
	) name174 (
		_w558_,
		_w559_,
		_w560_,
		_w636_,
		_w637_
	);
	LUT4 #(
		.INIT('h0155)
	) name175 (
		_w571_,
		_w572_,
		_w551_,
		_w603_,
		_w638_
	);
	LUT2 #(
		.INIT('h8)
	) name176 (
		_w566_,
		_w578_,
		_w639_
	);
	LUT4 #(
		.INIT('h0307)
	) name177 (
		_w570_,
		_w578_,
		_w584_,
		_w585_,
		_w640_
	);
	LUT4 #(
		.INIT('h4f00)
	) name178 (
		_w637_,
		_w638_,
		_w639_,
		_w640_,
		_w641_
	);
	LUT4 #(
		.INIT('h9565)
	) name179 (
		\P1_datao_reg[13]/NET0131 ,
		\si[13]_pad ,
		_w547_,
		_w641_,
		_w642_
	);
	LUT3 #(
		.INIT('ha6)
	) name180 (
		\P2_IR_reg[13]/NET0131 ,
		\P2_IR_reg[31]/NET0131 ,
		_w498_,
		_w643_
	);
	LUT3 #(
		.INIT('h10)
	) name181 (
		_w537_,
		_w545_,
		_w643_,
		_w644_
	);
	LUT3 #(
		.INIT('h0e)
	) name182 (
		_w546_,
		_w642_,
		_w644_,
		_w645_
	);
	LUT4 #(
		.INIT('hcc04)
	) name183 (
		_w546_,
		_w631_,
		_w642_,
		_w644_,
		_w646_
	);
	LUT4 #(
		.INIT('h0032)
	) name184 (
		_w546_,
		_w631_,
		_w642_,
		_w644_,
		_w647_
	);
	LUT3 #(
		.INIT('h63)
	) name185 (
		\P2_reg3_reg[11]/NET0131 ,
		\P2_reg3_reg[12]/NET0131 ,
		_w522_,
		_w648_
	);
	LUT4 #(
		.INIT('h0084)
	) name186 (
		\P2_IR_reg[30]/NET0131 ,
		_w505_,
		_w516_,
		_w648_,
		_w649_
	);
	LUT4 #(
		.INIT('h0408)
	) name187 (
		\P2_IR_reg[30]/NET0131 ,
		\P2_reg0_reg[12]/NET0131 ,
		_w505_,
		_w516_,
		_w650_
	);
	LUT4 #(
		.INIT('h0804)
	) name188 (
		\P2_IR_reg[30]/NET0131 ,
		\P2_reg2_reg[12]/NET0131 ,
		_w505_,
		_w516_,
		_w651_
	);
	LUT4 #(
		.INIT('h4080)
	) name189 (
		\P2_IR_reg[30]/NET0131 ,
		\P2_reg1_reg[12]/NET0131 ,
		_w505_,
		_w516_,
		_w652_
	);
	LUT4 #(
		.INIT('h0001)
	) name190 (
		_w649_,
		_w650_,
		_w651_,
		_w652_,
		_w653_
	);
	LUT4 #(
		.INIT('hfffe)
	) name191 (
		_w649_,
		_w650_,
		_w651_,
		_w652_,
		_w654_
	);
	LUT4 #(
		.INIT('h0155)
	) name192 (
		_w572_,
		_w550_,
		_w601_,
		_w634_,
		_w655_
	);
	LUT4 #(
		.INIT('h7f00)
	) name193 (
		_w561_,
		_w600_,
		_w634_,
		_w655_,
		_w656_
	);
	LUT3 #(
		.INIT('h04)
	) name194 (
		_w564_,
		_w566_,
		_w577_,
		_w657_
	);
	LUT4 #(
		.INIT('hfac8)
	) name195 (
		\P1_datao_reg[10]/NET0131 ,
		\P1_datao_reg[11]/NET0131 ,
		\si[10]_pad ,
		\si[11]_pad ,
		_w658_
	);
	LUT4 #(
		.INIT('h0133)
	) name196 (
		_w569_,
		_w585_,
		_w606_,
		_w658_,
		_w659_
	);
	LUT3 #(
		.INIT('hb0)
	) name197 (
		_w656_,
		_w657_,
		_w659_,
		_w660_
	);
	LUT4 #(
		.INIT('h9565)
	) name198 (
		\P1_datao_reg[12]/NET0131 ,
		\si[12]_pad ,
		_w547_,
		_w660_,
		_w661_
	);
	LUT4 #(
		.INIT('h2aaa)
	) name199 (
		\P2_IR_reg[31]/NET0131 ,
		_w495_,
		_w496_,
		_w497_,
		_w662_
	);
	LUT4 #(
		.INIT('hf0e0)
	) name200 (
		\P2_IR_reg[10]/NET0131 ,
		\P2_IR_reg[11]/NET0131 ,
		\P2_IR_reg[31]/NET0131 ,
		\P2_IR_reg[9]/NET0131 ,
		_w663_
	);
	LUT3 #(
		.INIT('h56)
	) name201 (
		\P2_IR_reg[12]/NET0131 ,
		_w662_,
		_w663_,
		_w664_
	);
	LUT3 #(
		.INIT('h10)
	) name202 (
		_w537_,
		_w545_,
		_w664_,
		_w665_
	);
	LUT3 #(
		.INIT('h0e)
	) name203 (
		_w546_,
		_w661_,
		_w665_,
		_w666_
	);
	LUT4 #(
		.INIT('h0032)
	) name204 (
		_w546_,
		_w653_,
		_w661_,
		_w665_,
		_w667_
	);
	LUT2 #(
		.INIT('h1)
	) name205 (
		_w647_,
		_w667_,
		_w668_
	);
	LUT3 #(
		.INIT('h54)
	) name206 (
		_w646_,
		_w647_,
		_w667_,
		_w669_
	);
	LUT2 #(
		.INIT('h4)
	) name207 (
		_w528_,
		_w594_,
		_w670_
	);
	LUT4 #(
		.INIT('hbb0b)
	) name208 (
		_w528_,
		_w594_,
		_w615_,
		_w623_,
		_w671_
	);
	LUT4 #(
		.INIT('h44d4)
	) name209 (
		_w528_,
		_w594_,
		_w615_,
		_w623_,
		_w672_
	);
	LUT3 #(
		.INIT('h07)
	) name210 (
		_w625_,
		_w669_,
		_w672_,
		_w673_
	);
	LUT2 #(
		.INIT('h9)
	) name211 (
		\P2_reg3_reg[11]/NET0131 ,
		_w522_,
		_w674_
	);
	LUT4 #(
		.INIT('h0084)
	) name212 (
		\P2_IR_reg[30]/NET0131 ,
		_w505_,
		_w516_,
		_w674_,
		_w675_
	);
	LUT4 #(
		.INIT('h0408)
	) name213 (
		\P2_IR_reg[30]/NET0131 ,
		\P2_reg0_reg[11]/NET0131 ,
		_w505_,
		_w516_,
		_w676_
	);
	LUT4 #(
		.INIT('h0804)
	) name214 (
		\P2_IR_reg[30]/NET0131 ,
		\P2_reg2_reg[11]/NET0131 ,
		_w505_,
		_w516_,
		_w677_
	);
	LUT4 #(
		.INIT('h4080)
	) name215 (
		\P2_IR_reg[30]/NET0131 ,
		\P2_reg1_reg[11]/NET0131 ,
		_w505_,
		_w516_,
		_w678_
	);
	LUT4 #(
		.INIT('h0001)
	) name216 (
		_w675_,
		_w676_,
		_w677_,
		_w678_,
		_w679_
	);
	LUT4 #(
		.INIT('hfffe)
	) name217 (
		_w675_,
		_w676_,
		_w677_,
		_w678_,
		_w680_
	);
	LUT4 #(
		.INIT('h9565)
	) name218 (
		\P1_datao_reg[11]/NET0131 ,
		\si[11]_pad ,
		_w547_,
		_w575_,
		_w681_
	);
	LUT4 #(
		.INIT('h2aaa)
	) name219 (
		\P2_IR_reg[31]/NET0131 ,
		_w496_,
		_w497_,
		_w538_,
		_w682_
	);
	LUT2 #(
		.INIT('h6)
	) name220 (
		\P2_IR_reg[11]/NET0131 ,
		_w682_,
		_w683_
	);
	LUT3 #(
		.INIT('h10)
	) name221 (
		_w537_,
		_w545_,
		_w683_,
		_w684_
	);
	LUT3 #(
		.INIT('h0e)
	) name222 (
		_w546_,
		_w681_,
		_w684_,
		_w685_
	);
	LUT4 #(
		.INIT('h0032)
	) name223 (
		_w546_,
		_w679_,
		_w681_,
		_w684_,
		_w686_
	);
	LUT4 #(
		.INIT('hcc04)
	) name224 (
		_w546_,
		_w679_,
		_w681_,
		_w684_,
		_w687_
	);
	LUT4 #(
		.INIT('h4080)
	) name225 (
		\P2_IR_reg[30]/NET0131 ,
		\P2_reg1_reg[10]/NET0131 ,
		_w505_,
		_w516_,
		_w688_
	);
	LUT4 #(
		.INIT('h0804)
	) name226 (
		\P2_IR_reg[30]/NET0131 ,
		\P2_reg2_reg[10]/NET0131 ,
		_w505_,
		_w516_,
		_w689_
	);
	LUT4 #(
		.INIT('h6555)
	) name227 (
		\P2_reg3_reg[10]/NET0131 ,
		\P2_reg3_reg[7]/NET0131 ,
		_w520_,
		_w521_,
		_w690_
	);
	LUT4 #(
		.INIT('h0084)
	) name228 (
		\P2_IR_reg[30]/NET0131 ,
		_w505_,
		_w516_,
		_w690_,
		_w691_
	);
	LUT4 #(
		.INIT('h0408)
	) name229 (
		\P2_IR_reg[30]/NET0131 ,
		\P2_reg0_reg[10]/NET0131 ,
		_w505_,
		_w516_,
		_w692_
	);
	LUT4 #(
		.INIT('h0001)
	) name230 (
		_w688_,
		_w689_,
		_w691_,
		_w692_,
		_w693_
	);
	LUT4 #(
		.INIT('hfffe)
	) name231 (
		_w688_,
		_w689_,
		_w691_,
		_w692_,
		_w694_
	);
	LUT2 #(
		.INIT('h2)
	) name232 (
		\P1_datao_reg[10]/NET0131 ,
		_w547_,
		_w695_
	);
	LUT2 #(
		.INIT('h6)
	) name233 (
		\P1_datao_reg[10]/NET0131 ,
		\si[10]_pad ,
		_w696_
	);
	LUT4 #(
		.INIT('h208a)
	) name234 (
		_w547_,
		_w605_,
		_w608_,
		_w696_,
		_w697_
	);
	LUT4 #(
		.INIT('heee0)
	) name235 (
		_w537_,
		_w545_,
		_w695_,
		_w697_,
		_w698_
	);
	LUT4 #(
		.INIT('haaa8)
	) name236 (
		\P2_IR_reg[31]/NET0131 ,
		\P2_IR_reg[7]/NET0131 ,
		\P2_IR_reg[8]/NET0131 ,
		\P2_IR_reg[9]/NET0131 ,
		_w699_
	);
	LUT4 #(
		.INIT('h00d5)
	) name237 (
		\P2_IR_reg[31]/NET0131 ,
		_w496_,
		_w497_,
		_w699_,
		_w700_
	);
	LUT2 #(
		.INIT('h9)
	) name238 (
		\P2_IR_reg[10]/NET0131 ,
		_w700_,
		_w701_
	);
	LUT3 #(
		.INIT('h10)
	) name239 (
		_w537_,
		_w545_,
		_w701_,
		_w702_
	);
	LUT2 #(
		.INIT('h1)
	) name240 (
		_w698_,
		_w702_,
		_w703_
	);
	LUT3 #(
		.INIT('ha8)
	) name241 (
		_w693_,
		_w698_,
		_w702_,
		_w704_
	);
	LUT2 #(
		.INIT('h1)
	) name242 (
		_w687_,
		_w704_,
		_w705_
	);
	LUT4 #(
		.INIT('h0408)
	) name243 (
		\P2_IR_reg[30]/NET0131 ,
		\P2_reg0_reg[9]/NET0131 ,
		_w505_,
		_w516_,
		_w706_
	);
	LUT4 #(
		.INIT('h1e0f)
	) name244 (
		\P2_reg3_reg[7]/NET0131 ,
		\P2_reg3_reg[8]/NET0131 ,
		\P2_reg3_reg[9]/NET0131 ,
		_w520_,
		_w707_
	);
	LUT4 #(
		.INIT('h0084)
	) name245 (
		\P2_IR_reg[30]/NET0131 ,
		_w505_,
		_w516_,
		_w707_,
		_w708_
	);
	LUT4 #(
		.INIT('h4080)
	) name246 (
		\P2_IR_reg[30]/NET0131 ,
		\P2_reg1_reg[9]/NET0131 ,
		_w505_,
		_w516_,
		_w709_
	);
	LUT4 #(
		.INIT('h0804)
	) name247 (
		\P2_IR_reg[30]/NET0131 ,
		\P2_reg2_reg[9]/NET0131 ,
		_w505_,
		_w516_,
		_w710_
	);
	LUT4 #(
		.INIT('h0001)
	) name248 (
		_w706_,
		_w708_,
		_w709_,
		_w710_,
		_w711_
	);
	LUT4 #(
		.INIT('hfffe)
	) name249 (
		_w706_,
		_w708_,
		_w709_,
		_w710_,
		_w712_
	);
	LUT2 #(
		.INIT('h2)
	) name250 (
		\P1_datao_reg[9]/NET0131 ,
		_w547_,
		_w713_
	);
	LUT2 #(
		.INIT('h6)
	) name251 (
		\P1_datao_reg[9]/NET0131 ,
		\si[9]_pad ,
		_w714_
	);
	LUT4 #(
		.INIT('h208a)
	) name252 (
		_w547_,
		_w637_,
		_w638_,
		_w714_,
		_w715_
	);
	LUT4 #(
		.INIT('heee0)
	) name253 (
		_w537_,
		_w545_,
		_w713_,
		_w715_,
		_w716_
	);
	LUT2 #(
		.INIT('h9)
	) name254 (
		\P2_IR_reg[9]/NET0131 ,
		_w662_,
		_w717_
	);
	LUT3 #(
		.INIT('h01)
	) name255 (
		_w537_,
		_w545_,
		_w717_,
		_w718_
	);
	LUT2 #(
		.INIT('h1)
	) name256 (
		_w716_,
		_w718_,
		_w719_
	);
	LUT3 #(
		.INIT('ha8)
	) name257 (
		_w711_,
		_w716_,
		_w718_,
		_w720_
	);
	LUT4 #(
		.INIT('h0804)
	) name258 (
		\P2_IR_reg[30]/NET0131 ,
		\P2_reg2_reg[8]/NET0131 ,
		_w505_,
		_w516_,
		_w721_
	);
	LUT4 #(
		.INIT('h0408)
	) name259 (
		\P2_IR_reg[30]/NET0131 ,
		\P2_reg0_reg[8]/NET0131 ,
		_w505_,
		_w516_,
		_w722_
	);
	LUT3 #(
		.INIT('h63)
	) name260 (
		\P2_reg3_reg[7]/NET0131 ,
		\P2_reg3_reg[8]/NET0131 ,
		_w520_,
		_w723_
	);
	LUT4 #(
		.INIT('h0084)
	) name261 (
		\P2_IR_reg[30]/NET0131 ,
		_w505_,
		_w516_,
		_w723_,
		_w724_
	);
	LUT4 #(
		.INIT('h4080)
	) name262 (
		\P2_IR_reg[30]/NET0131 ,
		\P2_reg1_reg[8]/NET0131 ,
		_w505_,
		_w516_,
		_w725_
	);
	LUT4 #(
		.INIT('h0001)
	) name263 (
		_w721_,
		_w722_,
		_w724_,
		_w725_,
		_w726_
	);
	LUT4 #(
		.INIT('hfffe)
	) name264 (
		_w721_,
		_w722_,
		_w724_,
		_w725_,
		_w727_
	);
	LUT4 #(
		.INIT('h9565)
	) name265 (
		\P1_datao_reg[8]/NET0131 ,
		\si[8]_pad ,
		_w547_,
		_w656_,
		_w728_
	);
	LUT4 #(
		.INIT('h8aaa)
	) name266 (
		\P2_IR_reg[31]/NET0131 ,
		\P2_IR_reg[7]/NET0131 ,
		_w496_,
		_w497_,
		_w729_
	);
	LUT2 #(
		.INIT('h6)
	) name267 (
		\P2_IR_reg[8]/NET0131 ,
		_w729_,
		_w730_
	);
	LUT4 #(
		.INIT('he0f1)
	) name268 (
		_w537_,
		_w545_,
		_w728_,
		_w730_,
		_w731_
	);
	LUT2 #(
		.INIT('h2)
	) name269 (
		_w726_,
		_w731_,
		_w732_
	);
	LUT3 #(
		.INIT('h01)
	) name270 (
		_w711_,
		_w716_,
		_w718_,
		_w733_
	);
	LUT3 #(
		.INIT('h01)
	) name271 (
		_w693_,
		_w698_,
		_w702_,
		_w734_
	);
	LUT4 #(
		.INIT('h00b2)
	) name272 (
		_w711_,
		_w719_,
		_w732_,
		_w734_,
		_w735_
	);
	LUT3 #(
		.INIT('h51)
	) name273 (
		_w686_,
		_w705_,
		_w735_,
		_w736_
	);
	LUT4 #(
		.INIT('hcc04)
	) name274 (
		_w546_,
		_w653_,
		_w661_,
		_w665_,
		_w737_
	);
	LUT2 #(
		.INIT('h1)
	) name275 (
		_w646_,
		_w737_,
		_w738_
	);
	LUT3 #(
		.INIT('h0d)
	) name276 (
		_w615_,
		_w623_,
		_w647_,
		_w739_
	);
	LUT4 #(
		.INIT('h1311)
	) name277 (
		_w625_,
		_w670_,
		_w738_,
		_w739_,
		_w740_
	);
	LUT3 #(
		.INIT('ha8)
	) name278 (
		_w673_,
		_w736_,
		_w740_,
		_w741_
	);
	LUT4 #(
		.INIT('h0408)
	) name279 (
		\P2_IR_reg[30]/NET0131 ,
		\P2_reg0_reg[6]/NET0131 ,
		_w505_,
		_w516_,
		_w742_
	);
	LUT4 #(
		.INIT('h0804)
	) name280 (
		\P2_IR_reg[30]/NET0131 ,
		\P2_reg2_reg[6]/NET0131 ,
		_w505_,
		_w516_,
		_w743_
	);
	LUT4 #(
		.INIT('h01fe)
	) name281 (
		\P2_reg3_reg[3]/NET0131 ,
		\P2_reg3_reg[4]/NET0131 ,
		\P2_reg3_reg[5]/NET0131 ,
		\P2_reg3_reg[6]/NET0131 ,
		_w744_
	);
	LUT4 #(
		.INIT('h0084)
	) name282 (
		\P2_IR_reg[30]/NET0131 ,
		_w505_,
		_w516_,
		_w744_,
		_w745_
	);
	LUT4 #(
		.INIT('h4080)
	) name283 (
		\P2_IR_reg[30]/NET0131 ,
		\P2_reg1_reg[6]/NET0131 ,
		_w505_,
		_w516_,
		_w746_
	);
	LUT4 #(
		.INIT('h0001)
	) name284 (
		_w742_,
		_w743_,
		_w745_,
		_w746_,
		_w747_
	);
	LUT4 #(
		.INIT('hfffe)
	) name285 (
		_w742_,
		_w743_,
		_w745_,
		_w746_,
		_w748_
	);
	LUT4 #(
		.INIT('h9565)
	) name286 (
		\P1_datao_reg[6]/NET0131 ,
		\si[6]_pad ,
		_w547_,
		_w602_,
		_w749_
	);
	LUT4 #(
		.INIT('h5755)
	) name287 (
		\P2_IR_reg[31]/NET0131 ,
		\P2_IR_reg[4]/NET0131 ,
		\P2_IR_reg[5]/NET0131 ,
		_w496_,
		_w750_
	);
	LUT2 #(
		.INIT('h9)
	) name288 (
		\P2_IR_reg[6]/NET0131 ,
		_w750_,
		_w751_
	);
	LUT4 #(
		.INIT('he0f1)
	) name289 (
		_w537_,
		_w545_,
		_w749_,
		_w751_,
		_w752_
	);
	LUT2 #(
		.INIT('h2)
	) name290 (
		_w747_,
		_w752_,
		_w753_
	);
	LUT4 #(
		.INIT('h0408)
	) name291 (
		\P2_IR_reg[30]/NET0131 ,
		\P2_reg0_reg[7]/NET0131 ,
		_w505_,
		_w516_,
		_w754_
	);
	LUT2 #(
		.INIT('h9)
	) name292 (
		\P2_reg3_reg[7]/NET0131 ,
		_w520_,
		_w755_
	);
	LUT4 #(
		.INIT('h0084)
	) name293 (
		\P2_IR_reg[30]/NET0131 ,
		_w505_,
		_w516_,
		_w755_,
		_w756_
	);
	LUT4 #(
		.INIT('h0804)
	) name294 (
		\P2_IR_reg[30]/NET0131 ,
		\P2_reg2_reg[7]/NET0131 ,
		_w505_,
		_w516_,
		_w757_
	);
	LUT4 #(
		.INIT('h4080)
	) name295 (
		\P2_IR_reg[30]/NET0131 ,
		\P2_reg1_reg[7]/NET0131 ,
		_w505_,
		_w516_,
		_w758_
	);
	LUT4 #(
		.INIT('h0001)
	) name296 (
		_w754_,
		_w756_,
		_w757_,
		_w758_,
		_w759_
	);
	LUT4 #(
		.INIT('hfffe)
	) name297 (
		_w754_,
		_w756_,
		_w757_,
		_w758_,
		_w760_
	);
	LUT4 #(
		.INIT('h9565)
	) name298 (
		\P1_datao_reg[7]/NET0131 ,
		\si[7]_pad ,
		_w547_,
		_w563_,
		_w761_
	);
	LUT4 #(
		.INIT('hc666)
	) name299 (
		\P2_IR_reg[31]/NET0131 ,
		\P2_IR_reg[7]/NET0131 ,
		_w496_,
		_w497_,
		_w762_
	);
	LUT4 #(
		.INIT('he0f1)
	) name300 (
		_w537_,
		_w545_,
		_w761_,
		_w762_,
		_w763_
	);
	LUT4 #(
		.INIT('hdd0d)
	) name301 (
		_w747_,
		_w752_,
		_w759_,
		_w763_,
		_w764_
	);
	LUT3 #(
		.INIT('h1e)
	) name302 (
		\P2_reg3_reg[3]/NET0131 ,
		\P2_reg3_reg[4]/NET0131 ,
		\P2_reg3_reg[5]/NET0131 ,
		_w765_
	);
	LUT4 #(
		.INIT('h0084)
	) name303 (
		\P2_IR_reg[30]/NET0131 ,
		_w505_,
		_w516_,
		_w765_,
		_w766_
	);
	LUT4 #(
		.INIT('h0408)
	) name304 (
		\P2_IR_reg[30]/NET0131 ,
		\P2_reg0_reg[5]/NET0131 ,
		_w505_,
		_w516_,
		_w767_
	);
	LUT4 #(
		.INIT('h4080)
	) name305 (
		\P2_IR_reg[30]/NET0131 ,
		\P2_reg1_reg[5]/NET0131 ,
		_w505_,
		_w516_,
		_w768_
	);
	LUT4 #(
		.INIT('h0804)
	) name306 (
		\P2_IR_reg[30]/NET0131 ,
		\P2_reg2_reg[5]/NET0131 ,
		_w505_,
		_w516_,
		_w769_
	);
	LUT4 #(
		.INIT('h0001)
	) name307 (
		_w766_,
		_w767_,
		_w768_,
		_w769_,
		_w770_
	);
	LUT4 #(
		.INIT('hfffe)
	) name308 (
		_w766_,
		_w767_,
		_w768_,
		_w769_,
		_w771_
	);
	LUT4 #(
		.INIT('h6595)
	) name309 (
		\P1_datao_reg[5]/NET0131 ,
		\si[5]_pad ,
		_w547_,
		_w633_,
		_w772_
	);
	LUT4 #(
		.INIT('h87a5)
	) name310 (
		\P2_IR_reg[31]/NET0131 ,
		\P2_IR_reg[4]/NET0131 ,
		\P2_IR_reg[5]/NET0131 ,
		_w496_,
		_w773_
	);
	LUT4 #(
		.INIT('hf1e0)
	) name311 (
		_w537_,
		_w545_,
		_w772_,
		_w773_,
		_w774_
	);
	LUT4 #(
		.INIT('hb0bb)
	) name312 (
		_w747_,
		_w752_,
		_w770_,
		_w774_,
		_w775_
	);
	LUT2 #(
		.INIT('h6)
	) name313 (
		\P2_reg3_reg[3]/NET0131 ,
		\P2_reg3_reg[4]/NET0131 ,
		_w776_
	);
	LUT4 #(
		.INIT('h0084)
	) name314 (
		\P2_IR_reg[30]/NET0131 ,
		_w505_,
		_w516_,
		_w776_,
		_w777_
	);
	LUT4 #(
		.INIT('h0408)
	) name315 (
		\P2_IR_reg[30]/NET0131 ,
		\P2_reg0_reg[4]/NET0131 ,
		_w505_,
		_w516_,
		_w778_
	);
	LUT4 #(
		.INIT('h4080)
	) name316 (
		\P2_IR_reg[30]/NET0131 ,
		\P2_reg1_reg[4]/NET0131 ,
		_w505_,
		_w516_,
		_w779_
	);
	LUT4 #(
		.INIT('h0804)
	) name317 (
		\P2_IR_reg[30]/NET0131 ,
		\P2_reg2_reg[4]/NET0131 ,
		_w505_,
		_w516_,
		_w780_
	);
	LUT4 #(
		.INIT('h0001)
	) name318 (
		_w777_,
		_w778_,
		_w779_,
		_w780_,
		_w781_
	);
	LUT4 #(
		.INIT('hfffe)
	) name319 (
		_w777_,
		_w778_,
		_w779_,
		_w780_,
		_w782_
	);
	LUT4 #(
		.INIT('h6595)
	) name320 (
		\P1_datao_reg[4]/NET0131 ,
		\si[4]_pad ,
		_w547_,
		_w600_,
		_w783_
	);
	LUT3 #(
		.INIT('hc6)
	) name321 (
		\P2_IR_reg[31]/NET0131 ,
		\P2_IR_reg[4]/NET0131 ,
		_w496_,
		_w784_
	);
	LUT4 #(
		.INIT('he0f1)
	) name322 (
		_w537_,
		_w545_,
		_w783_,
		_w784_,
		_w785_
	);
	LUT2 #(
		.INIT('h2)
	) name323 (
		_w781_,
		_w785_,
		_w786_
	);
	LUT4 #(
		.INIT('hdd0d)
	) name324 (
		_w770_,
		_w774_,
		_w781_,
		_w785_,
		_w787_
	);
	LUT4 #(
		.INIT('h0408)
	) name325 (
		\P2_IR_reg[30]/NET0131 ,
		\P2_reg0_reg[3]/NET0131 ,
		_w505_,
		_w516_,
		_w788_
	);
	LUT4 #(
		.INIT('h0804)
	) name326 (
		\P2_IR_reg[30]/NET0131 ,
		\P2_reg2_reg[3]/NET0131 ,
		_w505_,
		_w516_,
		_w789_
	);
	LUT4 #(
		.INIT('h2010)
	) name327 (
		\P2_IR_reg[30]/NET0131 ,
		\P2_reg3_reg[3]/NET0131 ,
		_w505_,
		_w516_,
		_w790_
	);
	LUT4 #(
		.INIT('h4080)
	) name328 (
		\P2_IR_reg[30]/NET0131 ,
		\P2_reg1_reg[3]/NET0131 ,
		_w505_,
		_w516_,
		_w791_
	);
	LUT4 #(
		.INIT('h0001)
	) name329 (
		_w788_,
		_w789_,
		_w790_,
		_w791_,
		_w792_
	);
	LUT4 #(
		.INIT('hfffe)
	) name330 (
		_w788_,
		_w789_,
		_w790_,
		_w791_,
		_w793_
	);
	LUT4 #(
		.INIT('hfe00)
	) name331 (
		\P2_IR_reg[0]/NET0131 ,
		\P2_IR_reg[1]/NET0131 ,
		\P2_IR_reg[2]/NET0131 ,
		\P2_IR_reg[31]/NET0131 ,
		_w794_
	);
	LUT2 #(
		.INIT('h6)
	) name332 (
		\P2_IR_reg[3]/NET0131 ,
		_w794_,
		_w795_
	);
	LUT4 #(
		.INIT('h9a6a)
	) name333 (
		\P1_datao_reg[3]/NET0131 ,
		\si[3]_pad ,
		_w547_,
		_w557_,
		_w796_
	);
	LUT4 #(
		.INIT('h01ef)
	) name334 (
		_w537_,
		_w545_,
		_w795_,
		_w796_,
		_w797_
	);
	LUT4 #(
		.INIT('hb0bb)
	) name335 (
		_w781_,
		_w785_,
		_w792_,
		_w797_,
		_w798_
	);
	LUT4 #(
		.INIT('h0804)
	) name336 (
		\P2_IR_reg[30]/NET0131 ,
		\P2_reg2_reg[2]/NET0131 ,
		_w505_,
		_w516_,
		_w799_
	);
	LUT4 #(
		.INIT('h0408)
	) name337 (
		\P2_IR_reg[30]/NET0131 ,
		\P2_reg0_reg[2]/NET0131 ,
		_w505_,
		_w516_,
		_w800_
	);
	LUT4 #(
		.INIT('h8040)
	) name338 (
		\P2_IR_reg[30]/NET0131 ,
		\P2_reg3_reg[2]/NET0131 ,
		_w505_,
		_w516_,
		_w801_
	);
	LUT4 #(
		.INIT('h4080)
	) name339 (
		\P2_IR_reg[30]/NET0131 ,
		\P2_reg1_reg[2]/NET0131 ,
		_w505_,
		_w516_,
		_w802_
	);
	LUT4 #(
		.INIT('h0001)
	) name340 (
		_w799_,
		_w800_,
		_w801_,
		_w802_,
		_w803_
	);
	LUT4 #(
		.INIT('hfffe)
	) name341 (
		_w799_,
		_w800_,
		_w801_,
		_w802_,
		_w804_
	);
	LUT4 #(
		.INIT('h9565)
	) name342 (
		\P1_datao_reg[2]/NET0131 ,
		\si[2]_pad ,
		_w547_,
		_w598_,
		_w805_
	);
	LUT4 #(
		.INIT('he10f)
	) name343 (
		\P2_IR_reg[0]/NET0131 ,
		\P2_IR_reg[1]/NET0131 ,
		\P2_IR_reg[2]/NET0131 ,
		\P2_IR_reg[31]/NET0131 ,
		_w806_
	);
	LUT4 #(
		.INIT('hf1e0)
	) name344 (
		_w537_,
		_w545_,
		_w805_,
		_w806_,
		_w807_
	);
	LUT2 #(
		.INIT('h2)
	) name345 (
		_w803_,
		_w807_,
		_w808_
	);
	LUT4 #(
		.INIT('hdd0d)
	) name346 (
		_w792_,
		_w797_,
		_w803_,
		_w807_,
		_w809_
	);
	LUT4 #(
		.INIT('h4080)
	) name347 (
		\P2_IR_reg[30]/NET0131 ,
		\P2_reg1_reg[1]/NET0131 ,
		_w505_,
		_w516_,
		_w810_
	);
	LUT4 #(
		.INIT('h8040)
	) name348 (
		\P2_IR_reg[30]/NET0131 ,
		\P2_reg3_reg[1]/NET0131 ,
		_w505_,
		_w516_,
		_w811_
	);
	LUT4 #(
		.INIT('h0804)
	) name349 (
		\P2_IR_reg[30]/NET0131 ,
		\P2_reg2_reg[1]/NET0131 ,
		_w505_,
		_w516_,
		_w812_
	);
	LUT4 #(
		.INIT('h0408)
	) name350 (
		\P2_IR_reg[30]/NET0131 ,
		\P2_reg0_reg[1]/NET0131 ,
		_w505_,
		_w516_,
		_w813_
	);
	LUT4 #(
		.INIT('h0001)
	) name351 (
		_w810_,
		_w811_,
		_w812_,
		_w813_,
		_w814_
	);
	LUT4 #(
		.INIT('hfffe)
	) name352 (
		_w810_,
		_w811_,
		_w812_,
		_w813_,
		_w815_
	);
	LUT3 #(
		.INIT('h93)
	) name353 (
		\P2_IR_reg[0]/NET0131 ,
		\P2_IR_reg[1]/NET0131 ,
		\P2_IR_reg[31]/NET0131 ,
		_w816_
	);
	LUT4 #(
		.INIT('h9a6a)
	) name354 (
		\P1_datao_reg[1]/NET0131 ,
		\si[1]_pad ,
		_w547_,
		_w554_,
		_w817_
	);
	LUT4 #(
		.INIT('h10fe)
	) name355 (
		_w537_,
		_w545_,
		_w816_,
		_w817_,
		_w818_
	);
	LUT4 #(
		.INIT('h8040)
	) name356 (
		\P2_IR_reg[30]/NET0131 ,
		\P2_reg3_reg[0]/NET0131 ,
		_w505_,
		_w516_,
		_w819_
	);
	LUT4 #(
		.INIT('h0804)
	) name357 (
		\P2_IR_reg[30]/NET0131 ,
		\P2_reg2_reg[0]/NET0131 ,
		_w505_,
		_w516_,
		_w820_
	);
	LUT4 #(
		.INIT('h4080)
	) name358 (
		\P2_IR_reg[30]/NET0131 ,
		\P2_reg1_reg[0]/NET0131 ,
		_w505_,
		_w516_,
		_w821_
	);
	LUT4 #(
		.INIT('h0408)
	) name359 (
		\P2_IR_reg[30]/NET0131 ,
		\P2_reg0_reg[0]/NET0131 ,
		_w505_,
		_w516_,
		_w822_
	);
	LUT4 #(
		.INIT('h0001)
	) name360 (
		_w819_,
		_w820_,
		_w821_,
		_w822_,
		_w823_
	);
	LUT4 #(
		.INIT('hfffe)
	) name361 (
		_w819_,
		_w820_,
		_w821_,
		_w822_,
		_w824_
	);
	LUT3 #(
		.INIT('h6a)
	) name362 (
		\P1_datao_reg[0]/NET0131 ,
		\si[0]_pad ,
		_w547_,
		_w825_
	);
	LUT4 #(
		.INIT('h01fd)
	) name363 (
		\P2_IR_reg[0]/NET0131 ,
		_w537_,
		_w545_,
		_w825_,
		_w826_
	);
	LUT4 #(
		.INIT('h0d00)
	) name364 (
		_w814_,
		_w818_,
		_w823_,
		_w826_,
		_w827_
	);
	LUT2 #(
		.INIT('h4)
	) name365 (
		_w803_,
		_w807_,
		_w828_
	);
	LUT4 #(
		.INIT('hb0bb)
	) name366 (
		_w803_,
		_w807_,
		_w814_,
		_w818_,
		_w829_
	);
	LUT4 #(
		.INIT('h2a22)
	) name367 (
		_w798_,
		_w809_,
		_w827_,
		_w829_,
		_w830_
	);
	LUT4 #(
		.INIT('h22a2)
	) name368 (
		_w764_,
		_w775_,
		_w787_,
		_w830_,
		_w831_
	);
	LUT2 #(
		.INIT('h1)
	) name369 (
		_w686_,
		_w734_,
		_w832_
	);
	LUT2 #(
		.INIT('h4)
	) name370 (
		_w726_,
		_w731_,
		_w833_
	);
	LUT2 #(
		.INIT('h4)
	) name371 (
		_w759_,
		_w763_,
		_w834_
	);
	LUT3 #(
		.INIT('h01)
	) name372 (
		_w733_,
		_w833_,
		_w834_,
		_w835_
	);
	LUT4 #(
		.INIT('h8000)
	) name373 (
		_w668_,
		_w671_,
		_w832_,
		_w835_,
		_w836_
	);
	LUT2 #(
		.INIT('h4)
	) name374 (
		_w831_,
		_w836_,
		_w837_
	);
	LUT4 #(
		.INIT('h0804)
	) name375 (
		\P2_IR_reg[30]/NET0131 ,
		\P2_reg2_reg[17]/NET0131 ,
		_w505_,
		_w516_,
		_w838_
	);
	LUT4 #(
		.INIT('h0408)
	) name376 (
		\P2_IR_reg[30]/NET0131 ,
		\P2_reg0_reg[17]/NET0131 ,
		_w505_,
		_w516_,
		_w839_
	);
	LUT2 #(
		.INIT('h1)
	) name377 (
		\P2_reg3_reg[15]/NET0131 ,
		\P2_reg3_reg[16]/NET0131 ,
		_w840_
	);
	LUT3 #(
		.INIT('h80)
	) name378 (
		_w522_,
		_w523_,
		_w840_,
		_w841_
	);
	LUT4 #(
		.INIT('h9555)
	) name379 (
		\P2_reg3_reg[17]/NET0131 ,
		_w522_,
		_w523_,
		_w840_,
		_w842_
	);
	LUT4 #(
		.INIT('h0084)
	) name380 (
		\P2_IR_reg[30]/NET0131 ,
		_w505_,
		_w516_,
		_w842_,
		_w843_
	);
	LUT4 #(
		.INIT('h4080)
	) name381 (
		\P2_IR_reg[30]/NET0131 ,
		\P2_reg1_reg[17]/NET0131 ,
		_w505_,
		_w516_,
		_w844_
	);
	LUT4 #(
		.INIT('h0001)
	) name382 (
		_w838_,
		_w839_,
		_w843_,
		_w844_,
		_w845_
	);
	LUT4 #(
		.INIT('hfffe)
	) name383 (
		_w838_,
		_w839_,
		_w843_,
		_w844_,
		_w846_
	);
	LUT2 #(
		.INIT('h2)
	) name384 (
		\P1_datao_reg[17]/NET0131 ,
		_w547_,
		_w847_
	);
	LUT2 #(
		.INIT('h1)
	) name385 (
		\P1_datao_reg[17]/NET0131 ,
		\si[17]_pad ,
		_w848_
	);
	LUT2 #(
		.INIT('h8)
	) name386 (
		\P1_datao_reg[17]/NET0131 ,
		\si[17]_pad ,
		_w849_
	);
	LUT2 #(
		.INIT('h6)
	) name387 (
		\P1_datao_reg[17]/NET0131 ,
		\si[17]_pad ,
		_w850_
	);
	LUT4 #(
		.INIT('hfac8)
	) name388 (
		\P1_datao_reg[15]/NET0131 ,
		\P1_datao_reg[16]/NET0131 ,
		\si[15]_pad ,
		\si[16]_pad ,
		_w851_
	);
	LUT2 #(
		.INIT('h8)
	) name389 (
		_w580_,
		_w851_,
		_w852_
	);
	LUT4 #(
		.INIT('hb000)
	) name390 (
		_w637_,
		_w638_,
		_w639_,
		_w852_,
		_w853_
	);
	LUT2 #(
		.INIT('h8)
	) name391 (
		\P1_datao_reg[16]/NET0131 ,
		\si[16]_pad ,
		_w854_
	);
	LUT4 #(
		.INIT('h001f)
	) name392 (
		_w583_,
		_w589_,
		_w851_,
		_w854_,
		_w855_
	);
	LUT3 #(
		.INIT('hb0)
	) name393 (
		_w640_,
		_w852_,
		_w855_,
		_w856_
	);
	LUT4 #(
		.INIT('h2822)
	) name394 (
		_w547_,
		_w850_,
		_w853_,
		_w856_,
		_w857_
	);
	LUT4 #(
		.INIT('ha666)
	) name395 (
		\P2_IR_reg[17]/NET0131 ,
		\P2_IR_reg[31]/NET0131 ,
		_w498_,
		_w500_,
		_w858_
	);
	LUT3 #(
		.INIT('h10)
	) name396 (
		_w537_,
		_w545_,
		_w858_,
		_w859_
	);
	LUT4 #(
		.INIT('h00ab)
	) name397 (
		_w546_,
		_w847_,
		_w857_,
		_w859_,
		_w860_
	);
	LUT4 #(
		.INIT('h0804)
	) name398 (
		\P2_IR_reg[30]/NET0131 ,
		\P2_reg2_reg[16]/NET0131 ,
		_w505_,
		_w516_,
		_w861_
	);
	LUT4 #(
		.INIT('h4080)
	) name399 (
		\P2_IR_reg[30]/NET0131 ,
		\P2_reg1_reg[16]/NET0131 ,
		_w505_,
		_w516_,
		_w862_
	);
	LUT4 #(
		.INIT('h6333)
	) name400 (
		\P2_reg3_reg[15]/NET0131 ,
		\P2_reg3_reg[16]/NET0131 ,
		_w522_,
		_w523_,
		_w863_
	);
	LUT4 #(
		.INIT('h0084)
	) name401 (
		\P2_IR_reg[30]/NET0131 ,
		_w505_,
		_w516_,
		_w863_,
		_w864_
	);
	LUT4 #(
		.INIT('h0408)
	) name402 (
		\P2_IR_reg[30]/NET0131 ,
		\P2_reg0_reg[16]/NET0131 ,
		_w505_,
		_w516_,
		_w865_
	);
	LUT4 #(
		.INIT('h0001)
	) name403 (
		_w861_,
		_w862_,
		_w864_,
		_w865_,
		_w866_
	);
	LUT4 #(
		.INIT('hfffe)
	) name404 (
		_w861_,
		_w862_,
		_w864_,
		_w865_,
		_w867_
	);
	LUT2 #(
		.INIT('h2)
	) name405 (
		\P1_datao_reg[16]/NET0131 ,
		_w547_,
		_w868_
	);
	LUT2 #(
		.INIT('h2)
	) name406 (
		_w580_,
		_w588_,
		_w869_
	);
	LUT3 #(
		.INIT('h04)
	) name407 (
		_w576_,
		_w580_,
		_w588_,
		_w870_
	);
	LUT3 #(
		.INIT('h40)
	) name408 (
		_w656_,
		_w657_,
		_w870_,
		_w871_
	);
	LUT4 #(
		.INIT('hec80)
	) name409 (
		\P1_datao_reg[14]/NET0131 ,
		\P1_datao_reg[15]/NET0131 ,
		\si[14]_pad ,
		\si[15]_pad ,
		_w872_
	);
	LUT4 #(
		.INIT('h3700)
	) name410 (
		_w576_,
		_w595_,
		_w659_,
		_w869_,
		_w873_
	);
	LUT2 #(
		.INIT('h1)
	) name411 (
		_w872_,
		_w873_,
		_w874_
	);
	LUT2 #(
		.INIT('h6)
	) name412 (
		\P1_datao_reg[16]/NET0131 ,
		\si[16]_pad ,
		_w875_
	);
	LUT4 #(
		.INIT('h208a)
	) name413 (
		_w547_,
		_w871_,
		_w874_,
		_w875_,
		_w876_
	);
	LUT4 #(
		.INIT('ha666)
	) name414 (
		\P2_IR_reg[16]/NET0131 ,
		\P2_IR_reg[31]/NET0131 ,
		_w506_,
		_w530_,
		_w877_
	);
	LUT3 #(
		.INIT('h10)
	) name415 (
		_w537_,
		_w545_,
		_w877_,
		_w878_
	);
	LUT4 #(
		.INIT('h00ab)
	) name416 (
		_w546_,
		_w868_,
		_w876_,
		_w878_,
		_w879_
	);
	LUT4 #(
		.INIT('hb0bb)
	) name417 (
		_w845_,
		_w860_,
		_w866_,
		_w879_,
		_w880_
	);
	LUT4 #(
		.INIT('h4080)
	) name418 (
		\P2_IR_reg[30]/NET0131 ,
		\P2_reg1_reg[19]/NET0131 ,
		_w505_,
		_w516_,
		_w881_
	);
	LUT4 #(
		.INIT('h0804)
	) name419 (
		\P2_IR_reg[30]/NET0131 ,
		\P2_reg2_reg[19]/NET0131 ,
		_w505_,
		_w516_,
		_w882_
	);
	LUT2 #(
		.INIT('h1)
	) name420 (
		_w881_,
		_w882_,
		_w883_
	);
	LUT2 #(
		.INIT('h1)
	) name421 (
		\P2_reg3_reg[17]/NET0131 ,
		\P2_reg3_reg[18]/NET0131 ,
		_w884_
	);
	LUT4 #(
		.INIT('h8000)
	) name422 (
		_w522_,
		_w523_,
		_w840_,
		_w884_,
		_w885_
	);
	LUT2 #(
		.INIT('h9)
	) name423 (
		\P2_reg3_reg[19]/NET0131 ,
		_w885_,
		_w886_
	);
	LUT4 #(
		.INIT('h0408)
	) name424 (
		\P2_IR_reg[30]/NET0131 ,
		\P2_reg0_reg[19]/NET0131 ,
		_w505_,
		_w516_,
		_w887_
	);
	LUT3 #(
		.INIT('h0d)
	) name425 (
		_w519_,
		_w886_,
		_w887_,
		_w888_
	);
	LUT2 #(
		.INIT('h8)
	) name426 (
		_w883_,
		_w888_,
		_w889_
	);
	LUT2 #(
		.INIT('h7)
	) name427 (
		_w883_,
		_w888_,
		_w890_
	);
	LUT4 #(
		.INIT('hfac8)
	) name428 (
		\P1_datao_reg[17]/NET0131 ,
		\P1_datao_reg[18]/NET0131 ,
		\si[17]_pad ,
		\si[18]_pad ,
		_w891_
	);
	LUT2 #(
		.INIT('h8)
	) name429 (
		_w851_,
		_w891_,
		_w892_
	);
	LUT4 #(
		.INIT('h0137)
	) name430 (
		\P1_datao_reg[17]/NET0131 ,
		\P1_datao_reg[18]/NET0131 ,
		\si[17]_pad ,
		\si[18]_pad ,
		_w893_
	);
	LUT4 #(
		.INIT('hec80)
	) name431 (
		\P1_datao_reg[17]/NET0131 ,
		\P1_datao_reg[18]/NET0131 ,
		\si[17]_pad ,
		\si[18]_pad ,
		_w894_
	);
	LUT4 #(
		.INIT('h137f)
	) name432 (
		\P1_datao_reg[15]/NET0131 ,
		\P1_datao_reg[16]/NET0131 ,
		\si[15]_pad ,
		\si[16]_pad ,
		_w895_
	);
	LUT3 #(
		.INIT('h45)
	) name433 (
		_w893_,
		_w894_,
		_w895_,
		_w896_
	);
	LUT3 #(
		.INIT('h0b)
	) name434 (
		_w587_,
		_w892_,
		_w896_,
		_w897_
	);
	LUT3 #(
		.INIT('h70)
	) name435 (
		_w582_,
		_w892_,
		_w897_,
		_w898_
	);
	LUT4 #(
		.INIT('h9565)
	) name436 (
		\P1_datao_reg[19]/NET0131 ,
		\si[19]_pad ,
		_w547_,
		_w898_,
		_w899_
	);
	LUT4 #(
		.INIT('h5999)
	) name437 (
		\P2_IR_reg[19]/NET0131 ,
		\P2_IR_reg[31]/NET0131 ,
		_w540_,
		_w541_,
		_w900_
	);
	LUT3 #(
		.INIT('h01)
	) name438 (
		_w537_,
		_w545_,
		_w900_,
		_w901_
	);
	LUT3 #(
		.INIT('h0e)
	) name439 (
		_w546_,
		_w899_,
		_w901_,
		_w902_
	);
	LUT4 #(
		.INIT('h0032)
	) name440 (
		_w546_,
		_w889_,
		_w899_,
		_w901_,
		_w903_
	);
	LUT4 #(
		.INIT('h0804)
	) name441 (
		\P2_IR_reg[30]/NET0131 ,
		\P2_reg2_reg[18]/NET0131 ,
		_w505_,
		_w516_,
		_w904_
	);
	LUT4 #(
		.INIT('h0408)
	) name442 (
		\P2_IR_reg[30]/NET0131 ,
		\P2_reg0_reg[18]/NET0131 ,
		_w505_,
		_w516_,
		_w905_
	);
	LUT2 #(
		.INIT('h1)
	) name443 (
		_w904_,
		_w905_,
		_w906_
	);
	LUT3 #(
		.INIT('h63)
	) name444 (
		\P2_reg3_reg[17]/NET0131 ,
		\P2_reg3_reg[18]/NET0131 ,
		_w841_,
		_w907_
	);
	LUT4 #(
		.INIT('h4080)
	) name445 (
		\P2_IR_reg[30]/NET0131 ,
		\P2_reg1_reg[18]/NET0131 ,
		_w505_,
		_w516_,
		_w908_
	);
	LUT3 #(
		.INIT('h0d)
	) name446 (
		_w519_,
		_w907_,
		_w908_,
		_w909_
	);
	LUT2 #(
		.INIT('h8)
	) name447 (
		_w906_,
		_w909_,
		_w910_
	);
	LUT2 #(
		.INIT('h7)
	) name448 (
		_w906_,
		_w909_,
		_w911_
	);
	LUT2 #(
		.INIT('h2)
	) name449 (
		\P1_datao_reg[18]/NET0131 ,
		_w547_,
		_w912_
	);
	LUT2 #(
		.INIT('h6)
	) name450 (
		\P1_datao_reg[18]/NET0131 ,
		\si[18]_pad ,
		_w913_
	);
	LUT4 #(
		.INIT('hfac8)
	) name451 (
		\P1_datao_reg[14]/NET0131 ,
		\P1_datao_reg[17]/NET0131 ,
		\si[14]_pad ,
		\si[17]_pad ,
		_w914_
	);
	LUT2 #(
		.INIT('h8)
	) name452 (
		_w851_,
		_w914_,
		_w915_
	);
	LUT4 #(
		.INIT('hb000)
	) name453 (
		_w605_,
		_w608_,
		_w610_,
		_w915_,
		_w916_
	);
	LUT4 #(
		.INIT('hfac8)
	) name454 (
		\P1_datao_reg[16]/NET0131 ,
		\P1_datao_reg[17]/NET0131 ,
		\si[16]_pad ,
		\si[17]_pad ,
		_w917_
	);
	LUT4 #(
		.INIT('h0155)
	) name455 (
		_w849_,
		_w854_,
		_w872_,
		_w917_,
		_w918_
	);
	LUT3 #(
		.INIT('h70)
	) name456 (
		_w597_,
		_w915_,
		_w918_,
		_w919_
	);
	LUT4 #(
		.INIT('h2822)
	) name457 (
		_w547_,
		_w913_,
		_w916_,
		_w919_,
		_w920_
	);
	LUT2 #(
		.INIT('h2)
	) name458 (
		\P2_IR_reg[31]/NET0131 ,
		_w509_,
		_w921_
	);
	LUT4 #(
		.INIT('h00d5)
	) name459 (
		\P2_IR_reg[31]/NET0131 ,
		_w506_,
		_w508_,
		_w921_,
		_w922_
	);
	LUT2 #(
		.INIT('h9)
	) name460 (
		\P2_IR_reg[18]/NET0131 ,
		_w922_,
		_w923_
	);
	LUT3 #(
		.INIT('h10)
	) name461 (
		_w537_,
		_w545_,
		_w923_,
		_w924_
	);
	LUT4 #(
		.INIT('h00ab)
	) name462 (
		_w546_,
		_w912_,
		_w920_,
		_w924_,
		_w925_
	);
	LUT2 #(
		.INIT('h4)
	) name463 (
		_w910_,
		_w925_,
		_w926_
	);
	LUT3 #(
		.INIT('h02)
	) name464 (
		_w880_,
		_w903_,
		_w926_,
		_w927_
	);
	LUT2 #(
		.INIT('h2)
	) name465 (
		_w910_,
		_w925_,
		_w928_
	);
	LUT4 #(
		.INIT('hcc04)
	) name466 (
		_w546_,
		_w889_,
		_w899_,
		_w901_,
		_w929_
	);
	LUT4 #(
		.INIT('hdd0d)
	) name467 (
		_w845_,
		_w860_,
		_w866_,
		_w879_,
		_w930_
	);
	LUT4 #(
		.INIT('hb0bb)
	) name468 (
		_w845_,
		_w860_,
		_w910_,
		_w925_,
		_w931_
	);
	LUT4 #(
		.INIT('h1011)
	) name469 (
		_w928_,
		_w929_,
		_w930_,
		_w931_,
		_w932_
	);
	LUT2 #(
		.INIT('h1)
	) name470 (
		_w903_,
		_w932_,
		_w933_
	);
	LUT4 #(
		.INIT('h001f)
	) name471 (
		_w741_,
		_w837_,
		_w927_,
		_w933_,
		_w934_
	);
	LUT2 #(
		.INIT('h2)
	) name472 (
		\P1_datao_reg[21]/NET0131 ,
		_w547_,
		_w935_
	);
	LUT2 #(
		.INIT('h1)
	) name473 (
		\P1_datao_reg[21]/NET0131 ,
		\si[21]_pad ,
		_w936_
	);
	LUT2 #(
		.INIT('h8)
	) name474 (
		\P1_datao_reg[21]/NET0131 ,
		\si[21]_pad ,
		_w937_
	);
	LUT2 #(
		.INIT('h6)
	) name475 (
		\P1_datao_reg[21]/NET0131 ,
		\si[21]_pad ,
		_w938_
	);
	LUT4 #(
		.INIT('hec80)
	) name476 (
		\P1_datao_reg[19]/NET0131 ,
		\P1_datao_reg[20]/NET0131 ,
		\si[19]_pad ,
		\si[20]_pad ,
		_w939_
	);
	LUT4 #(
		.INIT('hfac8)
	) name477 (
		\P1_datao_reg[19]/NET0131 ,
		\P1_datao_reg[20]/NET0131 ,
		\si[19]_pad ,
		\si[20]_pad ,
		_w940_
	);
	LUT3 #(
		.INIT('h13)
	) name478 (
		_w894_,
		_w939_,
		_w940_,
		_w941_
	);
	LUT2 #(
		.INIT('h8)
	) name479 (
		_w891_,
		_w940_,
		_w942_
	);
	LUT4 #(
		.INIT('h4f00)
	) name480 (
		_w641_,
		_w852_,
		_w855_,
		_w942_,
		_w943_
	);
	LUT4 #(
		.INIT('h2282)
	) name481 (
		_w547_,
		_w938_,
		_w941_,
		_w943_,
		_w944_
	);
	LUT3 #(
		.INIT('h54)
	) name482 (
		_w546_,
		_w935_,
		_w944_,
		_w945_
	);
	LUT4 #(
		.INIT('h0100)
	) name483 (
		\P2_reg3_reg[19]/NET0131 ,
		\P2_reg3_reg[20]/NET0131 ,
		\P2_reg3_reg[21]/NET0131 ,
		_w885_,
		_w946_
	);
	LUT4 #(
		.INIT('h1e0f)
	) name484 (
		\P2_reg3_reg[19]/NET0131 ,
		\P2_reg3_reg[20]/NET0131 ,
		\P2_reg3_reg[21]/NET0131 ,
		_w885_,
		_w947_
	);
	LUT2 #(
		.INIT('h2)
	) name485 (
		_w519_,
		_w947_,
		_w948_
	);
	LUT4 #(
		.INIT('h0804)
	) name486 (
		\P2_IR_reg[30]/NET0131 ,
		\P2_reg2_reg[21]/NET0131 ,
		_w505_,
		_w516_,
		_w949_
	);
	LUT4 #(
		.INIT('h4080)
	) name487 (
		\P2_IR_reg[30]/NET0131 ,
		\P2_reg1_reg[21]/NET0131 ,
		_w505_,
		_w516_,
		_w950_
	);
	LUT4 #(
		.INIT('h0408)
	) name488 (
		\P2_IR_reg[30]/NET0131 ,
		\P2_reg0_reg[21]/NET0131 ,
		_w505_,
		_w516_,
		_w951_
	);
	LUT3 #(
		.INIT('h01)
	) name489 (
		_w950_,
		_w951_,
		_w949_,
		_w952_
	);
	LUT2 #(
		.INIT('h4)
	) name490 (
		_w948_,
		_w952_,
		_w953_
	);
	LUT2 #(
		.INIT('hb)
	) name491 (
		_w948_,
		_w952_,
		_w954_
	);
	LUT4 #(
		.INIT('h00ab)
	) name492 (
		_w546_,
		_w935_,
		_w944_,
		_w953_,
		_w955_
	);
	LUT4 #(
		.INIT('hfac8)
	) name493 (
		\P1_datao_reg[18]/NET0131 ,
		\P1_datao_reg[19]/NET0131 ,
		\si[18]_pad ,
		\si[19]_pad ,
		_w956_
	);
	LUT2 #(
		.INIT('h8)
	) name494 (
		_w917_,
		_w956_,
		_w957_
	);
	LUT4 #(
		.INIT('hec80)
	) name495 (
		\P1_datao_reg[18]/NET0131 ,
		\P1_datao_reg[19]/NET0131 ,
		\si[18]_pad ,
		\si[19]_pad ,
		_w958_
	);
	LUT4 #(
		.INIT('h135f)
	) name496 (
		\P1_datao_reg[16]/NET0131 ,
		\P1_datao_reg[17]/NET0131 ,
		\si[16]_pad ,
		\si[17]_pad ,
		_w959_
	);
	LUT4 #(
		.INIT('h0f0b)
	) name497 (
		_w848_,
		_w956_,
		_w958_,
		_w959_,
		_w960_
	);
	LUT4 #(
		.INIT('h4f00)
	) name498 (
		_w871_,
		_w874_,
		_w957_,
		_w960_,
		_w961_
	);
	LUT4 #(
		.INIT('h9565)
	) name499 (
		\P1_datao_reg[20]/NET0131 ,
		\si[20]_pad ,
		_w547_,
		_w961_,
		_w962_
	);
	LUT3 #(
		.INIT('h63)
	) name500 (
		\P2_reg3_reg[19]/NET0131 ,
		\P2_reg3_reg[20]/NET0131 ,
		_w885_,
		_w963_
	);
	LUT2 #(
		.INIT('h2)
	) name501 (
		_w519_,
		_w963_,
		_w964_
	);
	LUT4 #(
		.INIT('h0408)
	) name502 (
		\P2_IR_reg[30]/NET0131 ,
		\P2_reg0_reg[20]/NET0131 ,
		_w505_,
		_w516_,
		_w965_
	);
	LUT4 #(
		.INIT('h4080)
	) name503 (
		\P2_IR_reg[30]/NET0131 ,
		\P2_reg1_reg[20]/NET0131 ,
		_w505_,
		_w516_,
		_w966_
	);
	LUT4 #(
		.INIT('h0804)
	) name504 (
		\P2_IR_reg[30]/NET0131 ,
		\P2_reg2_reg[20]/NET0131 ,
		_w505_,
		_w516_,
		_w967_
	);
	LUT3 #(
		.INIT('h01)
	) name505 (
		_w966_,
		_w967_,
		_w965_,
		_w968_
	);
	LUT2 #(
		.INIT('h4)
	) name506 (
		_w964_,
		_w968_,
		_w969_
	);
	LUT2 #(
		.INIT('hb)
	) name507 (
		_w964_,
		_w968_,
		_w970_
	);
	LUT3 #(
		.INIT('h0e)
	) name508 (
		_w546_,
		_w962_,
		_w969_,
		_w971_
	);
	LUT2 #(
		.INIT('h1)
	) name509 (
		\P1_datao_reg[23]/NET0131 ,
		\si[23]_pad ,
		_w972_
	);
	LUT2 #(
		.INIT('h8)
	) name510 (
		\P1_datao_reg[23]/NET0131 ,
		\si[23]_pad ,
		_w973_
	);
	LUT2 #(
		.INIT('h8)
	) name511 (
		\P1_datao_reg[22]/NET0131 ,
		\si[22]_pad ,
		_w974_
	);
	LUT4 #(
		.INIT('hfac8)
	) name512 (
		\P1_datao_reg[21]/NET0131 ,
		\P1_datao_reg[22]/NET0131 ,
		\si[21]_pad ,
		\si[22]_pad ,
		_w975_
	);
	LUT4 #(
		.INIT('h010f)
	) name513 (
		_w937_,
		_w939_,
		_w974_,
		_w975_,
		_w976_
	);
	LUT2 #(
		.INIT('h8)
	) name514 (
		_w940_,
		_w975_,
		_w977_
	);
	LUT3 #(
		.INIT('h4c)
	) name515 (
		_w896_,
		_w976_,
		_w977_,
		_w978_
	);
	LUT4 #(
		.INIT('h8000)
	) name516 (
		_w851_,
		_w891_,
		_w940_,
		_w975_,
		_w979_
	);
	LUT4 #(
		.INIT('h40f0)
	) name517 (
		_w582_,
		_w587_,
		_w978_,
		_w979_,
		_w980_
	);
	LUT4 #(
		.INIT('h9565)
	) name518 (
		\P1_datao_reg[23]/NET0131 ,
		\si[23]_pad ,
		_w547_,
		_w980_,
		_w981_
	);
	LUT2 #(
		.INIT('h1)
	) name519 (
		_w546_,
		_w981_,
		_w982_
	);
	LUT3 #(
		.INIT('h63)
	) name520 (
		\P2_reg3_reg[22]/NET0131 ,
		\P2_reg3_reg[23]/NET0131 ,
		_w946_,
		_w983_
	);
	LUT4 #(
		.INIT('h90c0)
	) name521 (
		\P2_reg3_reg[22]/NET0131 ,
		\P2_reg3_reg[23]/NET0131 ,
		_w519_,
		_w946_,
		_w984_
	);
	LUT4 #(
		.INIT('h4080)
	) name522 (
		\P2_IR_reg[30]/NET0131 ,
		\P2_reg1_reg[23]/NET0131 ,
		_w505_,
		_w516_,
		_w985_
	);
	LUT4 #(
		.INIT('h0408)
	) name523 (
		\P2_IR_reg[30]/NET0131 ,
		\P2_reg0_reg[23]/NET0131 ,
		_w505_,
		_w516_,
		_w986_
	);
	LUT4 #(
		.INIT('h0804)
	) name524 (
		\P2_IR_reg[30]/NET0131 ,
		\P2_reg2_reg[23]/NET0131 ,
		_w505_,
		_w516_,
		_w987_
	);
	LUT3 #(
		.INIT('h01)
	) name525 (
		_w986_,
		_w987_,
		_w985_,
		_w988_
	);
	LUT2 #(
		.INIT('h4)
	) name526 (
		_w984_,
		_w988_,
		_w989_
	);
	LUT2 #(
		.INIT('hb)
	) name527 (
		_w984_,
		_w988_,
		_w990_
	);
	LUT3 #(
		.INIT('h0e)
	) name528 (
		_w546_,
		_w981_,
		_w989_,
		_w991_
	);
	LUT4 #(
		.INIT('hfac8)
	) name529 (
		\P1_datao_reg[20]/NET0131 ,
		\P1_datao_reg[21]/NET0131 ,
		\si[20]_pad ,
		\si[21]_pad ,
		_w992_
	);
	LUT4 #(
		.INIT('hec80)
	) name530 (
		\P1_datao_reg[20]/NET0131 ,
		\P1_datao_reg[21]/NET0131 ,
		\si[20]_pad ,
		\si[21]_pad ,
		_w993_
	);
	LUT3 #(
		.INIT('h07)
	) name531 (
		_w958_,
		_w992_,
		_w993_,
		_w994_
	);
	LUT2 #(
		.INIT('h8)
	) name532 (
		_w956_,
		_w992_,
		_w995_
	);
	LUT3 #(
		.INIT('h8c)
	) name533 (
		_w918_,
		_w994_,
		_w995_,
		_w996_
	);
	LUT4 #(
		.INIT('h8000)
	) name534 (
		_w851_,
		_w914_,
		_w956_,
		_w992_,
		_w997_
	);
	LUT3 #(
		.INIT('h8c)
	) name535 (
		_w611_,
		_w996_,
		_w997_,
		_w998_
	);
	LUT4 #(
		.INIT('h9565)
	) name536 (
		\P1_datao_reg[22]/NET0131 ,
		\si[22]_pad ,
		_w547_,
		_w998_,
		_w999_
	);
	LUT2 #(
		.INIT('h9)
	) name537 (
		\P2_reg3_reg[22]/NET0131 ,
		_w946_,
		_w1000_
	);
	LUT3 #(
		.INIT('h48)
	) name538 (
		\P2_reg3_reg[22]/NET0131 ,
		_w519_,
		_w946_,
		_w1001_
	);
	LUT4 #(
		.INIT('h0804)
	) name539 (
		\P2_IR_reg[30]/NET0131 ,
		\P2_reg2_reg[22]/NET0131 ,
		_w505_,
		_w516_,
		_w1002_
	);
	LUT4 #(
		.INIT('h0408)
	) name540 (
		\P2_IR_reg[30]/NET0131 ,
		\P2_reg0_reg[22]/NET0131 ,
		_w505_,
		_w516_,
		_w1003_
	);
	LUT4 #(
		.INIT('h4080)
	) name541 (
		\P2_IR_reg[30]/NET0131 ,
		\P2_reg1_reg[22]/NET0131 ,
		_w505_,
		_w516_,
		_w1004_
	);
	LUT3 #(
		.INIT('h01)
	) name542 (
		_w1003_,
		_w1004_,
		_w1002_,
		_w1005_
	);
	LUT2 #(
		.INIT('h4)
	) name543 (
		_w1001_,
		_w1005_,
		_w1006_
	);
	LUT2 #(
		.INIT('hb)
	) name544 (
		_w1001_,
		_w1005_,
		_w1007_
	);
	LUT3 #(
		.INIT('h0e)
	) name545 (
		_w546_,
		_w999_,
		_w1006_,
		_w1008_
	);
	LUT4 #(
		.INIT('h0001)
	) name546 (
		_w955_,
		_w971_,
		_w991_,
		_w1008_,
		_w1009_
	);
	LUT3 #(
		.INIT('h10)
	) name547 (
		_w546_,
		_w999_,
		_w1006_,
		_w1010_
	);
	LUT3 #(
		.INIT('h10)
	) name548 (
		_w546_,
		_w981_,
		_w989_,
		_w1011_
	);
	LUT2 #(
		.INIT('h1)
	) name549 (
		_w1010_,
		_w1011_,
		_w1012_
	);
	LUT4 #(
		.INIT('h5400)
	) name550 (
		_w546_,
		_w935_,
		_w944_,
		_w953_,
		_w1013_
	);
	LUT3 #(
		.INIT('h10)
	) name551 (
		_w546_,
		_w962_,
		_w969_,
		_w1014_
	);
	LUT2 #(
		.INIT('h1)
	) name552 (
		_w1013_,
		_w1014_,
		_w1015_
	);
	LUT4 #(
		.INIT('h0e08)
	) name553 (
		_w945_,
		_w953_,
		_w1008_,
		_w1014_,
		_w1016_
	);
	LUT3 #(
		.INIT('h51)
	) name554 (
		_w991_,
		_w1012_,
		_w1016_,
		_w1017_
	);
	LUT2 #(
		.INIT('h1)
	) name555 (
		\P1_datao_reg[24]/NET0131 ,
		\si[24]_pad ,
		_w1018_
	);
	LUT4 #(
		.INIT('hec80)
	) name556 (
		\P1_datao_reg[23]/NET0131 ,
		\P1_datao_reg[24]/NET0131 ,
		\si[23]_pad ,
		\si[24]_pad ,
		_w1019_
	);
	LUT4 #(
		.INIT('hfac8)
	) name557 (
		\P1_datao_reg[22]/NET0131 ,
		\P1_datao_reg[23]/NET0131 ,
		\si[22]_pad ,
		\si[23]_pad ,
		_w1020_
	);
	LUT4 #(
		.INIT('h135f)
	) name558 (
		\P1_datao_reg[21]/NET0131 ,
		\P1_datao_reg[22]/NET0131 ,
		\si[21]_pad ,
		\si[22]_pad ,
		_w1021_
	);
	LUT4 #(
		.INIT('h3323)
	) name559 (
		_w1018_,
		_w1019_,
		_w1020_,
		_w1021_,
		_w1022_
	);
	LUT3 #(
		.INIT('h10)
	) name560 (
		_w936_,
		_w1018_,
		_w1020_,
		_w1023_
	);
	LUT4 #(
		.INIT('h40f0)
	) name561 (
		_w853_,
		_w856_,
		_w941_,
		_w942_,
		_w1024_
	);
	LUT3 #(
		.INIT('ha2)
	) name562 (
		_w1022_,
		_w1023_,
		_w1024_,
		_w1025_
	);
	LUT4 #(
		.INIT('h9565)
	) name563 (
		\P1_datao_reg[25]/NET0131 ,
		\si[25]_pad ,
		_w547_,
		_w1025_,
		_w1026_
	);
	LUT2 #(
		.INIT('h1)
	) name564 (
		_w546_,
		_w1026_,
		_w1027_
	);
	LUT2 #(
		.INIT('h1)
	) name565 (
		\P2_reg3_reg[23]/NET0131 ,
		\P2_reg3_reg[24]/NET0131 ,
		_w1028_
	);
	LUT4 #(
		.INIT('h1000)
	) name566 (
		\P2_reg3_reg[22]/NET0131 ,
		\P2_reg3_reg[25]/NET0131 ,
		_w946_,
		_w1028_,
		_w1029_
	);
	LUT4 #(
		.INIT('h6333)
	) name567 (
		\P2_reg3_reg[22]/NET0131 ,
		\P2_reg3_reg[25]/NET0131 ,
		_w946_,
		_w1028_,
		_w1030_
	);
	LUT4 #(
		.INIT('h0804)
	) name568 (
		\P2_IR_reg[30]/NET0131 ,
		\P2_reg2_reg[25]/NET0131 ,
		_w505_,
		_w516_,
		_w1031_
	);
	LUT4 #(
		.INIT('h4080)
	) name569 (
		\P2_IR_reg[30]/NET0131 ,
		\P2_reg1_reg[25]/NET0131 ,
		_w505_,
		_w516_,
		_w1032_
	);
	LUT4 #(
		.INIT('h0408)
	) name570 (
		\P2_IR_reg[30]/NET0131 ,
		\P2_reg0_reg[25]/NET0131 ,
		_w505_,
		_w516_,
		_w1033_
	);
	LUT3 #(
		.INIT('h01)
	) name571 (
		_w1032_,
		_w1033_,
		_w1031_,
		_w1034_
	);
	LUT3 #(
		.INIT('hd0)
	) name572 (
		_w519_,
		_w1030_,
		_w1034_,
		_w1035_
	);
	LUT3 #(
		.INIT('h2f)
	) name573 (
		_w519_,
		_w1030_,
		_w1034_,
		_w1036_
	);
	LUT3 #(
		.INIT('h0e)
	) name574 (
		_w546_,
		_w1026_,
		_w1035_,
		_w1037_
	);
	LUT4 #(
		.INIT('h0155)
	) name575 (
		_w973_,
		_w974_,
		_w993_,
		_w1020_,
		_w1038_
	);
	LUT2 #(
		.INIT('h8)
	) name576 (
		_w992_,
		_w1020_,
		_w1039_
	);
	LUT3 #(
		.INIT('h8c)
	) name577 (
		_w961_,
		_w1038_,
		_w1039_,
		_w1040_
	);
	LUT4 #(
		.INIT('h9565)
	) name578 (
		\P1_datao_reg[24]/NET0131 ,
		\si[24]_pad ,
		_w547_,
		_w1040_,
		_w1041_
	);
	LUT4 #(
		.INIT('h1e0f)
	) name579 (
		\P2_reg3_reg[22]/NET0131 ,
		\P2_reg3_reg[23]/NET0131 ,
		\P2_reg3_reg[24]/NET0131 ,
		_w946_,
		_w1042_
	);
	LUT4 #(
		.INIT('h4080)
	) name580 (
		\P2_IR_reg[30]/NET0131 ,
		\P2_reg1_reg[24]/NET0131 ,
		_w505_,
		_w516_,
		_w1043_
	);
	LUT4 #(
		.INIT('h0804)
	) name581 (
		\P2_IR_reg[30]/NET0131 ,
		\P2_reg2_reg[24]/NET0131 ,
		_w505_,
		_w516_,
		_w1044_
	);
	LUT4 #(
		.INIT('h0408)
	) name582 (
		\P2_IR_reg[30]/NET0131 ,
		\P2_reg0_reg[24]/NET0131 ,
		_w505_,
		_w516_,
		_w1045_
	);
	LUT3 #(
		.INIT('h01)
	) name583 (
		_w1044_,
		_w1045_,
		_w1043_,
		_w1046_
	);
	LUT3 #(
		.INIT('hd0)
	) name584 (
		_w519_,
		_w1042_,
		_w1046_,
		_w1047_
	);
	LUT3 #(
		.INIT('h2f)
	) name585 (
		_w519_,
		_w1042_,
		_w1046_,
		_w1048_
	);
	LUT3 #(
		.INIT('h0e)
	) name586 (
		_w546_,
		_w1041_,
		_w1047_,
		_w1049_
	);
	LUT2 #(
		.INIT('h1)
	) name587 (
		\P1_datao_reg[26]/NET0131 ,
		\si[26]_pad ,
		_w1050_
	);
	LUT4 #(
		.INIT('hec80)
	) name588 (
		\P1_datao_reg[24]/NET0131 ,
		\P1_datao_reg[25]/NET0131 ,
		\si[24]_pad ,
		\si[25]_pad ,
		_w1051_
	);
	LUT4 #(
		.INIT('hfac8)
	) name589 (
		\P1_datao_reg[24]/NET0131 ,
		\P1_datao_reg[25]/NET0131 ,
		\si[24]_pad ,
		\si[25]_pad ,
		_w1052_
	);
	LUT4 #(
		.INIT('h135f)
	) name590 (
		\P1_datao_reg[22]/NET0131 ,
		\P1_datao_reg[23]/NET0131 ,
		\si[22]_pad ,
		\si[23]_pad ,
		_w1053_
	);
	LUT4 #(
		.INIT('h3323)
	) name591 (
		_w972_,
		_w1051_,
		_w1052_,
		_w1053_,
		_w1054_
	);
	LUT4 #(
		.INIT('h40f0)
	) name592 (
		_w916_,
		_w919_,
		_w994_,
		_w995_,
		_w1055_
	);
	LUT2 #(
		.INIT('h8)
	) name593 (
		_w1020_,
		_w1052_,
		_w1056_
	);
	LUT3 #(
		.INIT('h8a)
	) name594 (
		_w1054_,
		_w1055_,
		_w1056_,
		_w1057_
	);
	LUT4 #(
		.INIT('h9565)
	) name595 (
		\P1_datao_reg[26]/NET0131 ,
		\si[26]_pad ,
		_w547_,
		_w1057_,
		_w1058_
	);
	LUT2 #(
		.INIT('h1)
	) name596 (
		_w546_,
		_w1058_,
		_w1059_
	);
	LUT4 #(
		.INIT('h0001)
	) name597 (
		\P2_reg3_reg[21]/NET0131 ,
		\P2_reg3_reg[22]/NET0131 ,
		\P2_reg3_reg[25]/NET0131 ,
		\P2_reg3_reg[26]/NET0131 ,
		_w1060_
	);
	LUT2 #(
		.INIT('h8)
	) name598 (
		_w1028_,
		_w1060_,
		_w1061_
	);
	LUT4 #(
		.INIT('h1000)
	) name599 (
		\P2_reg3_reg[19]/NET0131 ,
		\P2_reg3_reg[20]/NET0131 ,
		_w885_,
		_w1061_,
		_w1062_
	);
	LUT3 #(
		.INIT('h0d)
	) name600 (
		\P2_reg3_reg[26]/NET0131 ,
		_w1029_,
		_w1062_,
		_w1063_
	);
	LUT4 #(
		.INIT('hcc08)
	) name601 (
		\P2_reg3_reg[26]/NET0131 ,
		_w519_,
		_w1029_,
		_w1062_,
		_w1064_
	);
	LUT4 #(
		.INIT('h0408)
	) name602 (
		\P2_IR_reg[30]/NET0131 ,
		\P2_reg0_reg[26]/NET0131 ,
		_w505_,
		_w516_,
		_w1065_
	);
	LUT4 #(
		.INIT('h0804)
	) name603 (
		\P2_IR_reg[30]/NET0131 ,
		\P2_reg2_reg[26]/NET0131 ,
		_w505_,
		_w516_,
		_w1066_
	);
	LUT4 #(
		.INIT('h4080)
	) name604 (
		\P2_IR_reg[30]/NET0131 ,
		\P2_reg1_reg[26]/NET0131 ,
		_w505_,
		_w516_,
		_w1067_
	);
	LUT3 #(
		.INIT('h01)
	) name605 (
		_w1066_,
		_w1067_,
		_w1065_,
		_w1068_
	);
	LUT2 #(
		.INIT('h4)
	) name606 (
		_w1064_,
		_w1068_,
		_w1069_
	);
	LUT2 #(
		.INIT('hb)
	) name607 (
		_w1064_,
		_w1068_,
		_w1070_
	);
	LUT3 #(
		.INIT('h0e)
	) name608 (
		_w546_,
		_w1058_,
		_w1069_,
		_w1071_
	);
	LUT4 #(
		.INIT('hec80)
	) name609 (
		\P1_datao_reg[25]/NET0131 ,
		\P1_datao_reg[26]/NET0131 ,
		\si[25]_pad ,
		\si[26]_pad ,
		_w1072_
	);
	LUT4 #(
		.INIT('hfac8)
	) name610 (
		\P1_datao_reg[25]/NET0131 ,
		\P1_datao_reg[26]/NET0131 ,
		\si[25]_pad ,
		\si[26]_pad ,
		_w1073_
	);
	LUT3 #(
		.INIT('h13)
	) name611 (
		_w1019_,
		_w1072_,
		_w1073_,
		_w1074_
	);
	LUT3 #(
		.INIT('h10)
	) name612 (
		_w972_,
		_w1050_,
		_w1052_,
		_w1075_
	);
	LUT4 #(
		.INIT('h8f00)
	) name613 (
		_w582_,
		_w892_,
		_w897_,
		_w977_,
		_w1076_
	);
	LUT4 #(
		.INIT('h0c8c)
	) name614 (
		_w976_,
		_w1074_,
		_w1075_,
		_w1076_,
		_w1077_
	);
	LUT4 #(
		.INIT('h9565)
	) name615 (
		\P1_datao_reg[27]/NET0131 ,
		\si[27]_pad ,
		_w547_,
		_w1077_,
		_w1078_
	);
	LUT2 #(
		.INIT('h9)
	) name616 (
		\P2_reg3_reg[27]/NET0131 ,
		_w1062_,
		_w1079_
	);
	LUT3 #(
		.INIT('h48)
	) name617 (
		\P2_reg3_reg[27]/NET0131 ,
		_w519_,
		_w1062_,
		_w1080_
	);
	LUT4 #(
		.INIT('h0408)
	) name618 (
		\P2_IR_reg[30]/NET0131 ,
		\P2_reg0_reg[27]/NET0131 ,
		_w505_,
		_w516_,
		_w1081_
	);
	LUT4 #(
		.INIT('h4080)
	) name619 (
		\P2_IR_reg[30]/NET0131 ,
		\P2_reg1_reg[27]/NET0131 ,
		_w505_,
		_w516_,
		_w1082_
	);
	LUT4 #(
		.INIT('h0804)
	) name620 (
		\P2_IR_reg[30]/NET0131 ,
		\P2_reg2_reg[27]/NET0131 ,
		_w505_,
		_w516_,
		_w1083_
	);
	LUT3 #(
		.INIT('h01)
	) name621 (
		_w1082_,
		_w1083_,
		_w1081_,
		_w1084_
	);
	LUT2 #(
		.INIT('h4)
	) name622 (
		_w1080_,
		_w1084_,
		_w1085_
	);
	LUT2 #(
		.INIT('hb)
	) name623 (
		_w1080_,
		_w1084_,
		_w1086_
	);
	LUT3 #(
		.INIT('h0e)
	) name624 (
		_w546_,
		_w1078_,
		_w1085_,
		_w1087_
	);
	LUT2 #(
		.INIT('h1)
	) name625 (
		_w1071_,
		_w1087_,
		_w1088_
	);
	LUT4 #(
		.INIT('h0001)
	) name626 (
		_w1037_,
		_w1049_,
		_w1071_,
		_w1087_,
		_w1089_
	);
	LUT4 #(
		.INIT('hf400)
	) name627 (
		_w934_,
		_w1009_,
		_w1017_,
		_w1089_,
		_w1090_
	);
	LUT3 #(
		.INIT('h10)
	) name628 (
		_w546_,
		_w1058_,
		_w1069_,
		_w1091_
	);
	LUT3 #(
		.INIT('h10)
	) name629 (
		_w546_,
		_w1078_,
		_w1085_,
		_w1092_
	);
	LUT2 #(
		.INIT('h1)
	) name630 (
		_w1091_,
		_w1092_,
		_w1093_
	);
	LUT3 #(
		.INIT('h10)
	) name631 (
		_w546_,
		_w1026_,
		_w1035_,
		_w1094_
	);
	LUT3 #(
		.INIT('h10)
	) name632 (
		_w546_,
		_w1041_,
		_w1047_,
		_w1095_
	);
	LUT4 #(
		.INIT('h0e08)
	) name633 (
		_w1027_,
		_w1035_,
		_w1071_,
		_w1095_,
		_w1096_
	);
	LUT3 #(
		.INIT('h51)
	) name634 (
		_w1087_,
		_w1093_,
		_w1096_,
		_w1097_
	);
	LUT2 #(
		.INIT('h8)
	) name635 (
		\P1_datao_reg[29]/NET0131 ,
		\si[29]_pad ,
		_w1098_
	);
	LUT4 #(
		.INIT('hfac8)
	) name636 (
		\P1_datao_reg[27]/NET0131 ,
		\P1_datao_reg[28]/NET0131 ,
		\si[27]_pad ,
		\si[28]_pad ,
		_w1099_
	);
	LUT2 #(
		.INIT('h8)
	) name637 (
		_w1073_,
		_w1099_,
		_w1100_
	);
	LUT2 #(
		.INIT('h8)
	) name638 (
		_w1023_,
		_w1100_,
		_w1101_
	);
	LUT2 #(
		.INIT('h8)
	) name639 (
		\P1_datao_reg[28]/NET0131 ,
		\si[28]_pad ,
		_w1102_
	);
	LUT4 #(
		.INIT('hec80)
	) name640 (
		\P1_datao_reg[27]/NET0131 ,
		\P1_datao_reg[28]/NET0131 ,
		\si[27]_pad ,
		\si[28]_pad ,
		_w1103_
	);
	LUT4 #(
		.INIT('hdc00)
	) name641 (
		_w1022_,
		_w1072_,
		_w1073_,
		_w1099_,
		_w1104_
	);
	LUT2 #(
		.INIT('h1)
	) name642 (
		_w1103_,
		_w1104_,
		_w1105_
	);
	LUT4 #(
		.INIT('h2f00)
	) name643 (
		_w941_,
		_w943_,
		_w1101_,
		_w1105_,
		_w1106_
	);
	LUT4 #(
		.INIT('h9565)
	) name644 (
		\P1_datao_reg[29]/NET0131 ,
		\si[29]_pad ,
		_w547_,
		_w1106_,
		_w1107_
	);
	LUT2 #(
		.INIT('h1)
	) name645 (
		_w546_,
		_w1107_,
		_w1108_
	);
	LUT2 #(
		.INIT('h1)
	) name646 (
		\P2_reg3_reg[27]/NET0131 ,
		\P2_reg3_reg[28]/NET0131 ,
		_w1109_
	);
	LUT3 #(
		.INIT('h80)
	) name647 (
		_w519_,
		_w1062_,
		_w1109_,
		_w1110_
	);
	LUT4 #(
		.INIT('h0408)
	) name648 (
		\P2_IR_reg[30]/NET0131 ,
		\P2_reg0_reg[29]/NET0131 ,
		_w505_,
		_w516_,
		_w1111_
	);
	LUT4 #(
		.INIT('h0804)
	) name649 (
		\P2_IR_reg[30]/NET0131 ,
		\P2_reg2_reg[29]/NET0131 ,
		_w505_,
		_w516_,
		_w1112_
	);
	LUT4 #(
		.INIT('h4080)
	) name650 (
		\P2_IR_reg[30]/NET0131 ,
		\P2_reg1_reg[29]/NET0131 ,
		_w505_,
		_w516_,
		_w1113_
	);
	LUT3 #(
		.INIT('h01)
	) name651 (
		_w1112_,
		_w1113_,
		_w1111_,
		_w1114_
	);
	LUT2 #(
		.INIT('h4)
	) name652 (
		_w1110_,
		_w1114_,
		_w1115_
	);
	LUT2 #(
		.INIT('hb)
	) name653 (
		_w1110_,
		_w1114_,
		_w1116_
	);
	LUT3 #(
		.INIT('h0e)
	) name654 (
		_w546_,
		_w1107_,
		_w1115_,
		_w1117_
	);
	LUT4 #(
		.INIT('hfac8)
	) name655 (
		\P1_datao_reg[26]/NET0131 ,
		\P1_datao_reg[27]/NET0131 ,
		\si[26]_pad ,
		\si[27]_pad ,
		_w1118_
	);
	LUT2 #(
		.INIT('h8)
	) name656 (
		_w1052_,
		_w1118_,
		_w1119_
	);
	LUT4 #(
		.INIT('hec80)
	) name657 (
		\P1_datao_reg[26]/NET0131 ,
		\P1_datao_reg[27]/NET0131 ,
		\si[26]_pad ,
		\si[27]_pad ,
		_w1120_
	);
	LUT4 #(
		.INIT('hdc00)
	) name658 (
		_w1038_,
		_w1051_,
		_w1052_,
		_w1118_,
		_w1121_
	);
	LUT2 #(
		.INIT('h1)
	) name659 (
		_w1120_,
		_w1121_,
		_w1122_
	);
	LUT4 #(
		.INIT('hbf00)
	) name660 (
		_w961_,
		_w1039_,
		_w1119_,
		_w1122_,
		_w1123_
	);
	LUT4 #(
		.INIT('h9565)
	) name661 (
		\P1_datao_reg[28]/NET0131 ,
		\si[28]_pad ,
		_w547_,
		_w1123_,
		_w1124_
	);
	LUT3 #(
		.INIT('h63)
	) name662 (
		\P2_reg3_reg[27]/NET0131 ,
		\P2_reg3_reg[28]/NET0131 ,
		_w1062_,
		_w1125_
	);
	LUT4 #(
		.INIT('h90c0)
	) name663 (
		\P2_reg3_reg[27]/NET0131 ,
		\P2_reg3_reg[28]/NET0131 ,
		_w519_,
		_w1062_,
		_w1126_
	);
	LUT4 #(
		.INIT('h4080)
	) name664 (
		\P2_IR_reg[30]/NET0131 ,
		\P2_reg1_reg[28]/NET0131 ,
		_w505_,
		_w516_,
		_w1127_
	);
	LUT4 #(
		.INIT('h0408)
	) name665 (
		\P2_IR_reg[30]/NET0131 ,
		\P2_reg0_reg[28]/NET0131 ,
		_w505_,
		_w516_,
		_w1128_
	);
	LUT4 #(
		.INIT('h0804)
	) name666 (
		\P2_IR_reg[30]/NET0131 ,
		\P2_reg2_reg[28]/NET0131 ,
		_w505_,
		_w516_,
		_w1129_
	);
	LUT3 #(
		.INIT('h01)
	) name667 (
		_w1128_,
		_w1129_,
		_w1127_,
		_w1130_
	);
	LUT2 #(
		.INIT('h4)
	) name668 (
		_w1126_,
		_w1130_,
		_w1131_
	);
	LUT2 #(
		.INIT('hb)
	) name669 (
		_w1126_,
		_w1130_,
		_w1132_
	);
	LUT3 #(
		.INIT('h0e)
	) name670 (
		_w546_,
		_w1124_,
		_w1131_,
		_w1133_
	);
	LUT4 #(
		.INIT('h4080)
	) name671 (
		\P2_IR_reg[30]/NET0131 ,
		\P2_reg1_reg[31]/NET0131 ,
		_w505_,
		_w516_,
		_w1134_
	);
	LUT4 #(
		.INIT('h0804)
	) name672 (
		\P2_IR_reg[30]/NET0131 ,
		\P2_reg2_reg[31]/NET0131 ,
		_w505_,
		_w516_,
		_w1135_
	);
	LUT4 #(
		.INIT('h0408)
	) name673 (
		\P2_IR_reg[30]/NET0131 ,
		\P2_reg0_reg[31]/NET0131 ,
		_w505_,
		_w516_,
		_w1136_
	);
	LUT3 #(
		.INIT('h01)
	) name674 (
		_w1135_,
		_w1136_,
		_w1134_,
		_w1137_
	);
	LUT2 #(
		.INIT('h4)
	) name675 (
		_w1110_,
		_w1137_,
		_w1138_
	);
	LUT2 #(
		.INIT('hb)
	) name676 (
		_w1110_,
		_w1137_,
		_w1139_
	);
	LUT4 #(
		.INIT('hfac8)
	) name677 (
		\P1_datao_reg[29]/NET0131 ,
		\P1_datao_reg[30]/NET0131 ,
		\si[29]_pad ,
		\si[30]_pad ,
		_w1140_
	);
	LUT2 #(
		.INIT('h8)
	) name678 (
		_w1099_,
		_w1140_,
		_w1141_
	);
	LUT2 #(
		.INIT('h8)
	) name679 (
		_w1075_,
		_w1141_,
		_w1142_
	);
	LUT4 #(
		.INIT('hb000)
	) name680 (
		_w582_,
		_w587_,
		_w979_,
		_w1142_,
		_w1143_
	);
	LUT4 #(
		.INIT('hb300)
	) name681 (
		_w896_,
		_w976_,
		_w977_,
		_w1075_,
		_w1144_
	);
	LUT2 #(
		.INIT('h8)
	) name682 (
		\P1_datao_reg[30]/NET0131 ,
		\si[30]_pad ,
		_w1145_
	);
	LUT4 #(
		.INIT('h001f)
	) name683 (
		_w1098_,
		_w1103_,
		_w1140_,
		_w1145_,
		_w1146_
	);
	LUT4 #(
		.INIT('h3b00)
	) name684 (
		_w1074_,
		_w1141_,
		_w1144_,
		_w1146_,
		_w1147_
	);
	LUT4 #(
		.INIT('h4844)
	) name685 (
		\si[31]_pad ,
		_w547_,
		_w1143_,
		_w1147_,
		_w1148_
	);
	LUT3 #(
		.INIT('h12)
	) name686 (
		\P1_datao_reg[31]/NET0131 ,
		_w546_,
		_w1148_,
		_w1149_
	);
	LUT4 #(
		.INIT('h1020)
	) name687 (
		\P1_datao_reg[31]/NET0131 ,
		_w546_,
		_w1138_,
		_w1148_,
		_w1150_
	);
	LUT4 #(
		.INIT('hfac8)
	) name688 (
		\P1_datao_reg[28]/NET0131 ,
		\P1_datao_reg[29]/NET0131 ,
		\si[28]_pad ,
		\si[29]_pad ,
		_w1151_
	);
	LUT2 #(
		.INIT('h8)
	) name689 (
		_w1118_,
		_w1151_,
		_w1152_
	);
	LUT4 #(
		.INIT('h8000)
	) name690 (
		_w1020_,
		_w1052_,
		_w1118_,
		_w1151_,
		_w1153_
	);
	LUT4 #(
		.INIT('h7300)
	) name691 (
		_w918_,
		_w994_,
		_w995_,
		_w1056_,
		_w1154_
	);
	LUT4 #(
		.INIT('h0155)
	) name692 (
		_w1098_,
		_w1102_,
		_w1120_,
		_w1151_,
		_w1155_
	);
	LUT4 #(
		.INIT('h3b00)
	) name693 (
		_w1054_,
		_w1152_,
		_w1154_,
		_w1155_,
		_w1156_
	);
	LUT4 #(
		.INIT('hbf00)
	) name694 (
		_w611_,
		_w997_,
		_w1153_,
		_w1156_,
		_w1157_
	);
	LUT4 #(
		.INIT('h9565)
	) name695 (
		\P1_datao_reg[30]/NET0131 ,
		\si[30]_pad ,
		_w547_,
		_w1157_,
		_w1158_
	);
	LUT4 #(
		.INIT('h4080)
	) name696 (
		\P2_IR_reg[30]/NET0131 ,
		\P2_reg1_reg[30]/NET0131 ,
		_w505_,
		_w516_,
		_w1159_
	);
	LUT4 #(
		.INIT('h0804)
	) name697 (
		\P2_IR_reg[30]/NET0131 ,
		\P2_reg2_reg[30]/NET0131 ,
		_w505_,
		_w516_,
		_w1160_
	);
	LUT4 #(
		.INIT('h0408)
	) name698 (
		\P2_IR_reg[30]/NET0131 ,
		\P2_reg0_reg[30]/NET0131 ,
		_w505_,
		_w516_,
		_w1161_
	);
	LUT3 #(
		.INIT('h01)
	) name699 (
		_w1160_,
		_w1161_,
		_w1159_,
		_w1162_
	);
	LUT2 #(
		.INIT('h4)
	) name700 (
		_w1110_,
		_w1162_,
		_w1163_
	);
	LUT2 #(
		.INIT('hb)
	) name701 (
		_w1110_,
		_w1162_,
		_w1164_
	);
	LUT3 #(
		.INIT('h0e)
	) name702 (
		_w546_,
		_w1158_,
		_w1163_,
		_w1165_
	);
	LUT2 #(
		.INIT('h1)
	) name703 (
		_w1150_,
		_w1165_,
		_w1166_
	);
	LUT3 #(
		.INIT('h10)
	) name704 (
		_w1117_,
		_w1133_,
		_w1166_,
		_w1167_
	);
	LUT4 #(
		.INIT('h0e0d)
	) name705 (
		\P1_datao_reg[31]/NET0131 ,
		_w546_,
		_w1138_,
		_w1148_,
		_w1168_
	);
	LUT3 #(
		.INIT('h10)
	) name706 (
		_w546_,
		_w1158_,
		_w1163_,
		_w1169_
	);
	LUT2 #(
		.INIT('h1)
	) name707 (
		_w1168_,
		_w1169_,
		_w1170_
	);
	LUT3 #(
		.INIT('h54)
	) name708 (
		_w1150_,
		_w1168_,
		_w1169_,
		_w1171_
	);
	LUT3 #(
		.INIT('h10)
	) name709 (
		_w546_,
		_w1107_,
		_w1115_,
		_w1172_
	);
	LUT3 #(
		.INIT('h10)
	) name710 (
		_w546_,
		_w1124_,
		_w1131_,
		_w1173_
	);
	LUT4 #(
		.INIT('he080)
	) name711 (
		_w1108_,
		_w1115_,
		_w1166_,
		_w1173_,
		_w1174_
	);
	LUT2 #(
		.INIT('h1)
	) name712 (
		_w1171_,
		_w1174_,
		_w1175_
	);
	LUT4 #(
		.INIT('h1f00)
	) name713 (
		_w1090_,
		_w1097_,
		_w1167_,
		_w1175_,
		_w1176_
	);
	LUT2 #(
		.INIT('h2)
	) name714 (
		\P2_IR_reg[31]/NET0131 ,
		_w501_,
		_w1177_
	);
	LUT4 #(
		.INIT('h00d5)
	) name715 (
		\P2_IR_reg[31]/NET0131 ,
		_w498_,
		_w500_,
		_w1177_,
		_w1178_
	);
	LUT2 #(
		.INIT('h9)
	) name716 (
		\P2_IR_reg[21]/NET0131 ,
		_w1178_,
		_w1179_
	);
	LUT4 #(
		.INIT('h0001)
	) name717 (
		\P2_IR_reg[16]/NET0131 ,
		\P2_IR_reg[17]/NET0131 ,
		\P2_IR_reg[18]/NET0131 ,
		\P2_IR_reg[19]/NET0131 ,
		_w1180_
	);
	LUT2 #(
		.INIT('h2)
	) name718 (
		\P2_IR_reg[31]/NET0131 ,
		_w1180_,
		_w1181_
	);
	LUT4 #(
		.INIT('h00d5)
	) name719 (
		\P2_IR_reg[31]/NET0131 ,
		_w506_,
		_w530_,
		_w1181_,
		_w1182_
	);
	LUT2 #(
		.INIT('h9)
	) name720 (
		\P2_IR_reg[20]/NET0131 ,
		_w1182_,
		_w1183_
	);
	LUT4 #(
		.INIT('h1428)
	) name721 (
		\P2_IR_reg[20]/NET0131 ,
		\P2_IR_reg[21]/NET0131 ,
		_w1178_,
		_w1182_,
		_w1184_
	);
	LUT4 #(
		.INIT('h2aaa)
	) name722 (
		\P2_IR_reg[31]/NET0131 ,
		_w506_,
		_w508_,
		_w511_,
		_w1185_
	);
	LUT2 #(
		.INIT('h6)
	) name723 (
		\P2_IR_reg[22]/NET0131 ,
		_w1185_,
		_w1186_
	);
	LUT2 #(
		.INIT('h2)
	) name724 (
		\P2_IR_reg[31]/NET0131 ,
		_w531_,
		_w1187_
	);
	LUT4 #(
		.INIT('h00d5)
	) name725 (
		\P2_IR_reg[31]/NET0131 ,
		_w540_,
		_w541_,
		_w1187_,
		_w1188_
	);
	LUT2 #(
		.INIT('h9)
	) name726 (
		\P2_IR_reg[23]/NET0131 ,
		_w1188_,
		_w1189_
	);
	LUT4 #(
		.INIT('h4812)
	) name727 (
		\P2_IR_reg[22]/NET0131 ,
		\P2_IR_reg[23]/NET0131 ,
		_w1185_,
		_w1188_,
		_w1190_
	);
	LUT2 #(
		.INIT('h8)
	) name728 (
		_w1184_,
		_w1190_,
		_w1191_
	);
	LUT3 #(
		.INIT('hb0)
	) name729 (
		\P2_B_reg/NET0131 ,
		_w1176_,
		_w1191_,
		_w1192_
	);
	LUT4 #(
		.INIT('h000e)
	) name730 (
		_w1117_,
		_w1133_,
		_w1169_,
		_w1172_,
		_w1193_
	);
	LUT3 #(
		.INIT('h31)
	) name731 (
		_w1166_,
		_w1168_,
		_w1193_,
		_w1194_
	);
	LUT4 #(
		.INIT('h0001)
	) name732 (
		_w1091_,
		_w1092_,
		_w1094_,
		_w1095_,
		_w1195_
	);
	LUT4 #(
		.INIT('h0001)
	) name733 (
		_w1010_,
		_w1011_,
		_w1013_,
		_w1014_,
		_w1196_
	);
	LUT4 #(
		.INIT('h4d44)
	) name734 (
		_w845_,
		_w860_,
		_w866_,
		_w879_,
		_w1197_
	);
	LUT3 #(
		.INIT('h10)
	) name735 (
		_w928_,
		_w929_,
		_w1197_,
		_w1198_
	);
	LUT3 #(
		.INIT('hd4)
	) name736 (
		_w889_,
		_w902_,
		_w926_,
		_w1199_
	);
	LUT2 #(
		.INIT('h1)
	) name737 (
		_w1198_,
		_w1199_,
		_w1200_
	);
	LUT3 #(
		.INIT('h10)
	) name738 (
		_w928_,
		_w929_,
		_w930_,
		_w1201_
	);
	LUT2 #(
		.INIT('h8)
	) name739 (
		_w625_,
		_w738_,
		_w1202_
	);
	LUT3 #(
		.INIT('h54)
	) name740 (
		_w720_,
		_w733_,
		_w833_,
		_w1203_
	);
	LUT3 #(
		.INIT('h32)
	) name741 (
		_w686_,
		_w687_,
		_w734_,
		_w1204_
	);
	LUT3 #(
		.INIT('h07)
	) name742 (
		_w705_,
		_w1203_,
		_w1204_,
		_w1205_
	);
	LUT3 #(
		.INIT('ha2)
	) name743 (
		_w673_,
		_w1202_,
		_w1205_,
		_w1206_
	);
	LUT4 #(
		.INIT('h44c4)
	) name744 (
		_w673_,
		_w1201_,
		_w1202_,
		_w1205_,
		_w1207_
	);
	LUT3 #(
		.INIT('ha2)
	) name745 (
		_w1196_,
		_w1200_,
		_w1207_,
		_w1208_
	);
	LUT2 #(
		.INIT('h8)
	) name746 (
		_w1196_,
		_w1201_,
		_w1209_
	);
	LUT4 #(
		.INIT('hdd4d)
	) name747 (
		_w814_,
		_w818_,
		_w823_,
		_w826_,
		_w1210_
	);
	LUT4 #(
		.INIT('h4d44)
	) name748 (
		_w792_,
		_w797_,
		_w803_,
		_w807_,
		_w1211_
	);
	LUT4 #(
		.INIT('haa80)
	) name749 (
		_w787_,
		_w809_,
		_w1210_,
		_w1211_,
		_w1212_
	);
	LUT4 #(
		.INIT('h4d44)
	) name750 (
		_w770_,
		_w774_,
		_w781_,
		_w785_,
		_w1213_
	);
	LUT4 #(
		.INIT('h4f04)
	) name751 (
		_w747_,
		_w752_,
		_w759_,
		_w763_,
		_w1214_
	);
	LUT4 #(
		.INIT('h0057)
	) name752 (
		_w764_,
		_w1212_,
		_w1213_,
		_w1214_,
		_w1215_
	);
	LUT4 #(
		.INIT('h0001)
	) name753 (
		_w687_,
		_w704_,
		_w720_,
		_w732_,
		_w1216_
	);
	LUT3 #(
		.INIT('h20)
	) name754 (
		_w1202_,
		_w1215_,
		_w1216_,
		_w1217_
	);
	LUT3 #(
		.INIT('h71)
	) name755 (
		_w945_,
		_w953_,
		_w971_,
		_w1218_
	);
	LUT3 #(
		.INIT('h71)
	) name756 (
		_w982_,
		_w989_,
		_w1008_,
		_w1219_
	);
	LUT3 #(
		.INIT('h07)
	) name757 (
		_w1012_,
		_w1218_,
		_w1219_,
		_w1220_
	);
	LUT3 #(
		.INIT('h70)
	) name758 (
		_w1209_,
		_w1217_,
		_w1220_,
		_w1221_
	);
	LUT3 #(
		.INIT('h71)
	) name759 (
		_w1027_,
		_w1035_,
		_w1049_,
		_w1222_
	);
	LUT4 #(
		.INIT('h000e)
	) name760 (
		_w1037_,
		_w1049_,
		_w1091_,
		_w1094_,
		_w1223_
	);
	LUT3 #(
		.INIT('h31)
	) name761 (
		_w1088_,
		_w1092_,
		_w1223_,
		_w1224_
	);
	LUT4 #(
		.INIT('h0075)
	) name762 (
		_w1195_,
		_w1208_,
		_w1221_,
		_w1224_,
		_w1225_
	);
	LUT3 #(
		.INIT('h02)
	) name763 (
		_w1170_,
		_w1172_,
		_w1173_,
		_w1226_
	);
	LUT4 #(
		.INIT('h1011)
	) name764 (
		\P2_B_reg/NET0131 ,
		_w1194_,
		_w1225_,
		_w1226_,
		_w1227_
	);
	LUT4 #(
		.INIT('h8421)
	) name765 (
		\P2_IR_reg[22]/NET0131 ,
		\P2_IR_reg[23]/NET0131 ,
		_w1185_,
		_w1188_,
		_w1228_
	);
	LUT4 #(
		.INIT('h2814)
	) name766 (
		\P2_IR_reg[20]/NET0131 ,
		\P2_IR_reg[21]/NET0131 ,
		_w1178_,
		_w1182_,
		_w1229_
	);
	LUT2 #(
		.INIT('h8)
	) name767 (
		_w1228_,
		_w1229_,
		_w1230_
	);
	LUT2 #(
		.INIT('h4)
	) name768 (
		_w1227_,
		_w1230_,
		_w1231_
	);
	LUT4 #(
		.INIT('h2184)
	) name769 (
		\P2_IR_reg[22]/NET0131 ,
		\P2_IR_reg[23]/NET0131 ,
		_w1185_,
		_w1188_,
		_w1232_
	);
	LUT2 #(
		.INIT('h8)
	) name770 (
		_w1229_,
		_w1232_,
		_w1233_
	);
	LUT4 #(
		.INIT('hba00)
	) name771 (
		_w1194_,
		_w1225_,
		_w1226_,
		_w1233_,
		_w1234_
	);
	LUT3 #(
		.INIT('h8a)
	) name772 (
		_w1209_,
		_w1217_,
		_w1206_,
		_w1235_
	);
	LUT3 #(
		.INIT('ha8)
	) name773 (
		_w1196_,
		_w1198_,
		_w1199_,
		_w1236_
	);
	LUT2 #(
		.INIT('h2)
	) name774 (
		_w1220_,
		_w1236_,
		_w1237_
	);
	LUT3 #(
		.INIT('hab)
	) name775 (
		_w1110_,
		_w1137_,
		_w1162_,
		_w1238_
	);
	LUT3 #(
		.INIT('h01)
	) name776 (
		_w546_,
		_w1158_,
		_w1238_,
		_w1239_
	);
	LUT2 #(
		.INIT('h1)
	) name777 (
		_w1168_,
		_w1239_,
		_w1240_
	);
	LUT3 #(
		.INIT('h10)
	) name778 (
		_w1172_,
		_w1173_,
		_w1240_,
		_w1241_
	);
	LUT2 #(
		.INIT('h8)
	) name779 (
		_w1195_,
		_w1241_,
		_w1242_
	);
	LUT3 #(
		.INIT('hb0)
	) name780 (
		_w1235_,
		_w1237_,
		_w1242_,
		_w1243_
	);
	LUT4 #(
		.INIT('h3100)
	) name781 (
		_w1088_,
		_w1092_,
		_w1223_,
		_w1241_,
		_w1244_
	);
	LUT4 #(
		.INIT('h0e00)
	) name782 (
		_w1117_,
		_w1133_,
		_w1172_,
		_w1240_,
		_w1245_
	);
	LUT4 #(
		.INIT('h3301)
	) name783 (
		_w546_,
		_w1138_,
		_w1158_,
		_w1163_,
		_w1246_
	);
	LUT2 #(
		.INIT('h2)
	) name784 (
		_w1149_,
		_w1246_,
		_w1247_
	);
	LUT2 #(
		.INIT('h1)
	) name785 (
		_w1245_,
		_w1247_,
		_w1248_
	);
	LUT2 #(
		.INIT('h4)
	) name786 (
		_w1244_,
		_w1248_,
		_w1249_
	);
	LUT3 #(
		.INIT('h20)
	) name787 (
		_w1179_,
		_w1183_,
		_w1190_,
		_w1250_
	);
	LUT4 #(
		.INIT('hba00)
	) name788 (
		\P2_B_reg/NET0131 ,
		_w1243_,
		_w1249_,
		_w1250_,
		_w1251_
	);
	LUT3 #(
		.INIT('h80)
	) name789 (
		_w1179_,
		_w1183_,
		_w1190_,
		_w1252_
	);
	LUT4 #(
		.INIT('h447f)
	) name790 (
		_w1179_,
		_w1183_,
		_w1190_,
		_w1228_,
		_w1253_
	);
	LUT2 #(
		.INIT('h2)
	) name791 (
		\P2_B_reg/NET0131 ,
		_w1253_,
		_w1254_
	);
	LUT3 #(
		.INIT('he0)
	) name792 (
		_w546_,
		_w1058_,
		_w1069_,
		_w1255_
	);
	LUT3 #(
		.INIT('h01)
	) name793 (
		_w546_,
		_w1058_,
		_w1069_,
		_w1256_
	);
	LUT3 #(
		.INIT('h1e)
	) name794 (
		_w546_,
		_w1058_,
		_w1069_,
		_w1257_
	);
	LUT3 #(
		.INIT('he0)
	) name795 (
		_w546_,
		_w1124_,
		_w1131_,
		_w1258_
	);
	LUT3 #(
		.INIT('h01)
	) name796 (
		_w546_,
		_w1124_,
		_w1131_,
		_w1259_
	);
	LUT3 #(
		.INIT('h1e)
	) name797 (
		_w546_,
		_w1124_,
		_w1131_,
		_w1260_
	);
	LUT3 #(
		.INIT('h01)
	) name798 (
		_w546_,
		_w1078_,
		_w1085_,
		_w1261_
	);
	LUT3 #(
		.INIT('he0)
	) name799 (
		_w546_,
		_w1078_,
		_w1085_,
		_w1262_
	);
	LUT3 #(
		.INIT('h1e)
	) name800 (
		_w546_,
		_w1078_,
		_w1085_,
		_w1263_
	);
	LUT3 #(
		.INIT('he1)
	) name801 (
		_w546_,
		_w1107_,
		_w1115_,
		_w1264_
	);
	LUT4 #(
		.INIT('h0100)
	) name802 (
		_w1257_,
		_w1260_,
		_w1263_,
		_w1264_,
		_w1265_
	);
	LUT3 #(
		.INIT('he0)
	) name803 (
		_w546_,
		_w1041_,
		_w1047_,
		_w1266_
	);
	LUT3 #(
		.INIT('h01)
	) name804 (
		_w546_,
		_w1041_,
		_w1047_,
		_w1267_
	);
	LUT3 #(
		.INIT('h1e)
	) name805 (
		_w546_,
		_w1041_,
		_w1047_,
		_w1268_
	);
	LUT3 #(
		.INIT('he0)
	) name806 (
		_w546_,
		_w1026_,
		_w1035_,
		_w1269_
	);
	LUT3 #(
		.INIT('h01)
	) name807 (
		_w546_,
		_w1026_,
		_w1035_,
		_w1270_
	);
	LUT3 #(
		.INIT('h1e)
	) name808 (
		_w546_,
		_w1026_,
		_w1035_,
		_w1271_
	);
	LUT4 #(
		.INIT('h33c9)
	) name809 (
		_w546_,
		_w889_,
		_w899_,
		_w901_,
		_w1272_
	);
	LUT3 #(
		.INIT('he0)
	) name810 (
		_w546_,
		_w999_,
		_w1006_,
		_w1273_
	);
	LUT3 #(
		.INIT('h01)
	) name811 (
		_w546_,
		_w999_,
		_w1006_,
		_w1274_
	);
	LUT3 #(
		.INIT('h1e)
	) name812 (
		_w546_,
		_w999_,
		_w1006_,
		_w1275_
	);
	LUT3 #(
		.INIT('h01)
	) name813 (
		_w546_,
		_w981_,
		_w989_,
		_w1276_
	);
	LUT3 #(
		.INIT('he0)
	) name814 (
		_w546_,
		_w981_,
		_w989_,
		_w1277_
	);
	LUT3 #(
		.INIT('h1e)
	) name815 (
		_w546_,
		_w981_,
		_w989_,
		_w1278_
	);
	LUT3 #(
		.INIT('h10)
	) name816 (
		_w1275_,
		_w1278_,
		_w1272_,
		_w1279_
	);
	LUT3 #(
		.INIT('h10)
	) name817 (
		_w1271_,
		_w1268_,
		_w1279_,
		_w1280_
	);
	LUT4 #(
		.INIT('h0054)
	) name818 (
		_w546_,
		_w935_,
		_w944_,
		_w953_,
		_w1281_
	);
	LUT4 #(
		.INIT('hab00)
	) name819 (
		_w546_,
		_w935_,
		_w944_,
		_w953_,
		_w1282_
	);
	LUT4 #(
		.INIT('h54ab)
	) name820 (
		_w546_,
		_w935_,
		_w944_,
		_w953_,
		_w1283_
	);
	LUT4 #(
		.INIT('he1d2)
	) name821 (
		\P1_datao_reg[31]/NET0131 ,
		_w546_,
		_w1138_,
		_w1148_,
		_w1284_
	);
	LUT2 #(
		.INIT('h4)
	) name822 (
		_w1283_,
		_w1284_,
		_w1285_
	);
	LUT3 #(
		.INIT('he1)
	) name823 (
		_w546_,
		_w1158_,
		_w1163_,
		_w1286_
	);
	LUT3 #(
		.INIT('he0)
	) name824 (
		_w546_,
		_w962_,
		_w969_,
		_w1287_
	);
	LUT3 #(
		.INIT('h01)
	) name825 (
		_w546_,
		_w962_,
		_w969_,
		_w1288_
	);
	LUT3 #(
		.INIT('h1e)
	) name826 (
		_w546_,
		_w962_,
		_w969_,
		_w1289_
	);
	LUT2 #(
		.INIT('h8)
	) name827 (
		_w910_,
		_w925_,
		_w1290_
	);
	LUT2 #(
		.INIT('h1)
	) name828 (
		_w910_,
		_w925_,
		_w1291_
	);
	LUT2 #(
		.INIT('h6)
	) name829 (
		_w910_,
		_w925_,
		_w1292_
	);
	LUT3 #(
		.INIT('h10)
	) name830 (
		_w1289_,
		_w1292_,
		_w1286_,
		_w1293_
	);
	LUT2 #(
		.INIT('h9)
	) name831 (
		_w866_,
		_w879_,
		_w1294_
	);
	LUT2 #(
		.INIT('h6)
	) name832 (
		_w528_,
		_w594_,
		_w1295_
	);
	LUT2 #(
		.INIT('h9)
	) name833 (
		_w615_,
		_w623_,
		_w1296_
	);
	LUT4 #(
		.INIT('h9009)
	) name834 (
		_w528_,
		_w594_,
		_w615_,
		_w623_,
		_w1297_
	);
	LUT2 #(
		.INIT('h8)
	) name835 (
		_w1294_,
		_w1297_,
		_w1298_
	);
	LUT4 #(
		.INIT('h33c9)
	) name836 (
		_w546_,
		_w631_,
		_w642_,
		_w644_,
		_w1299_
	);
	LUT4 #(
		.INIT('h00c8)
	) name837 (
		_w546_,
		_w653_,
		_w661_,
		_w665_,
		_w1300_
	);
	LUT4 #(
		.INIT('h3301)
	) name838 (
		_w546_,
		_w653_,
		_w661_,
		_w665_,
		_w1301_
	);
	LUT4 #(
		.INIT('hcc36)
	) name839 (
		_w546_,
		_w653_,
		_w661_,
		_w665_,
		_w1302_
	);
	LUT2 #(
		.INIT('h9)
	) name840 (
		_w759_,
		_w763_,
		_w1303_
	);
	LUT4 #(
		.INIT('h9009)
	) name841 (
		_w759_,
		_w763_,
		_w814_,
		_w818_,
		_w1304_
	);
	LUT2 #(
		.INIT('h9)
	) name842 (
		_w823_,
		_w826_,
		_w1305_
	);
	LUT2 #(
		.INIT('h9)
	) name843 (
		_w770_,
		_w774_,
		_w1306_
	);
	LUT4 #(
		.INIT('h9009)
	) name844 (
		_w770_,
		_w774_,
		_w823_,
		_w826_,
		_w1307_
	);
	LUT2 #(
		.INIT('h8)
	) name845 (
		_w726_,
		_w731_,
		_w1308_
	);
	LUT2 #(
		.INIT('h1)
	) name846 (
		_w726_,
		_w731_,
		_w1309_
	);
	LUT2 #(
		.INIT('h6)
	) name847 (
		_w726_,
		_w731_,
		_w1310_
	);
	LUT3 #(
		.INIT('h56)
	) name848 (
		_w711_,
		_w716_,
		_w718_,
		_w1311_
	);
	LUT4 #(
		.INIT('h4000)
	) name849 (
		_w1310_,
		_w1311_,
		_w1304_,
		_w1307_,
		_w1312_
	);
	LUT3 #(
		.INIT('h40)
	) name850 (
		_w1302_,
		_w1299_,
		_w1312_,
		_w1313_
	);
	LUT2 #(
		.INIT('h9)
	) name851 (
		_w845_,
		_w860_,
		_w1314_
	);
	LUT3 #(
		.INIT('h54)
	) name852 (
		_w693_,
		_w698_,
		_w702_,
		_w1315_
	);
	LUT3 #(
		.INIT('h02)
	) name853 (
		_w693_,
		_w698_,
		_w702_,
		_w1316_
	);
	LUT3 #(
		.INIT('ha9)
	) name854 (
		_w693_,
		_w698_,
		_w702_,
		_w1317_
	);
	LUT4 #(
		.INIT('h00c8)
	) name855 (
		_w546_,
		_w679_,
		_w681_,
		_w684_,
		_w1318_
	);
	LUT4 #(
		.INIT('h3301)
	) name856 (
		_w546_,
		_w679_,
		_w681_,
		_w684_,
		_w1319_
	);
	LUT4 #(
		.INIT('hcc36)
	) name857 (
		_w546_,
		_w679_,
		_w681_,
		_w684_,
		_w1320_
	);
	LUT2 #(
		.INIT('h9)
	) name858 (
		_w803_,
		_w807_,
		_w1321_
	);
	LUT2 #(
		.INIT('h6)
	) name859 (
		_w747_,
		_w752_,
		_w1322_
	);
	LUT4 #(
		.INIT('h9009)
	) name860 (
		_w747_,
		_w752_,
		_w803_,
		_w807_,
		_w1323_
	);
	LUT2 #(
		.INIT('h8)
	) name861 (
		_w781_,
		_w785_,
		_w1324_
	);
	LUT2 #(
		.INIT('h6)
	) name862 (
		_w781_,
		_w785_,
		_w1325_
	);
	LUT2 #(
		.INIT('h6)
	) name863 (
		_w792_,
		_w797_,
		_w1326_
	);
	LUT4 #(
		.INIT('h9009)
	) name864 (
		_w781_,
		_w785_,
		_w792_,
		_w797_,
		_w1327_
	);
	LUT4 #(
		.INIT('h1000)
	) name865 (
		_w1320_,
		_w1317_,
		_w1323_,
		_w1327_,
		_w1328_
	);
	LUT2 #(
		.INIT('h8)
	) name866 (
		_w1314_,
		_w1328_,
		_w1329_
	);
	LUT4 #(
		.INIT('h8000)
	) name867 (
		_w1313_,
		_w1329_,
		_w1298_,
		_w1293_,
		_w1330_
	);
	LUT4 #(
		.INIT('h8000)
	) name868 (
		_w1285_,
		_w1330_,
		_w1280_,
		_w1265_,
		_w1331_
	);
	LUT4 #(
		.INIT('h8421)
	) name869 (
		\P2_IR_reg[21]/NET0131 ,
		\P2_IR_reg[22]/NET0131 ,
		_w1178_,
		_w1185_,
		_w1332_
	);
	LUT4 #(
		.INIT('h2133)
	) name870 (
		_w1183_,
		_w1254_,
		_w1331_,
		_w1332_,
		_w1333_
	);
	LUT4 #(
		.INIT('h4f00)
	) name871 (
		_w1243_,
		_w1249_,
		_w1252_,
		_w1333_,
		_w1334_
	);
	LUT3 #(
		.INIT('h10)
	) name872 (
		_w1234_,
		_w1251_,
		_w1334_,
		_w1335_
	);
	LUT2 #(
		.INIT('h2)
	) name873 (
		_w1184_,
		_w1186_,
		_w1336_
	);
	LUT4 #(
		.INIT('h4500)
	) name874 (
		_w1194_,
		_w1225_,
		_w1226_,
		_w1336_,
		_w1337_
	);
	LUT4 #(
		.INIT('h1248)
	) name875 (
		\P2_IR_reg[22]/NET0131 ,
		\P2_IR_reg[23]/NET0131 ,
		_w1185_,
		_w1188_,
		_w1338_
	);
	LUT2 #(
		.INIT('h8)
	) name876 (
		_w1179_,
		_w1338_,
		_w1339_
	);
	LUT4 #(
		.INIT('h9a00)
	) name877 (
		_w1183_,
		_w1243_,
		_w1249_,
		_w1339_,
		_w1340_
	);
	LUT2 #(
		.INIT('h1)
	) name878 (
		_w1337_,
		_w1340_,
		_w1341_
	);
	LUT4 #(
		.INIT('h1000)
	) name879 (
		_w1192_,
		_w1231_,
		_w1335_,
		_w1341_,
		_w1342_
	);
	LUT2 #(
		.INIT('h8)
	) name880 (
		_w1190_,
		_w1229_,
		_w1343_
	);
	LUT3 #(
		.INIT('he0)
	) name881 (
		\P2_B_reg/NET0131 ,
		_w1176_,
		_w1343_,
		_w1344_
	);
	LUT3 #(
		.INIT('h40)
	) name882 (
		_w1179_,
		_w1183_,
		_w1338_,
		_w1345_
	);
	LUT3 #(
		.INIT('h10)
	) name883 (
		_w1179_,
		_w1183_,
		_w1338_,
		_w1346_
	);
	LUT3 #(
		.INIT('hd8)
	) name884 (
		_w1176_,
		_w1345_,
		_w1346_,
		_w1347_
	);
	LUT2 #(
		.INIT('h1)
	) name885 (
		_w1344_,
		_w1347_,
		_w1348_
	);
	LUT3 #(
		.INIT('h82)
	) name886 (
		\P1_state_reg[0]/NET0131 ,
		\P2_IR_reg[23]/NET0131 ,
		_w1188_,
		_w1349_
	);
	LUT4 #(
		.INIT('h3faa)
	) name887 (
		\P2_B_reg/NET0131 ,
		_w1342_,
		_w1348_,
		_w1349_,
		_w1350_
	);
	LUT2 #(
		.INIT('h2)
	) name888 (
		\P2_IR_reg[31]/NET0131 ,
		_w512_,
		_w1351_
	);
	LUT3 #(
		.INIT('h56)
	) name889 (
		\P2_IR_reg[26]/NET0131 ,
		_w1185_,
		_w1351_,
		_w1352_
	);
	LUT4 #(
		.INIT('h2aaa)
	) name890 (
		\P2_IR_reg[31]/NET0131 ,
		_w500_,
		_w501_,
		_w502_,
		_w1353_
	);
	LUT4 #(
		.INIT('h55a6)
	) name891 (
		\P2_IR_reg[25]/NET0131 ,
		\P2_IR_reg[31]/NET0131 ,
		_w498_,
		_w1353_,
		_w1354_
	);
	LUT2 #(
		.INIT('h6)
	) name892 (
		\P2_IR_reg[24]/NET0131 ,
		_w534_,
		_w1355_
	);
	LUT3 #(
		.INIT('h60)
	) name893 (
		\P2_IR_reg[24]/NET0131 ,
		_w534_,
		_w1354_,
		_w1356_
	);
	LUT3 #(
		.INIT('h40)
	) name894 (
		_w1189_,
		_w1352_,
		_w1356_,
		_w1357_
	);
	LUT2 #(
		.INIT('h4)
	) name895 (
		_w1079_,
		_w1357_,
		_w1358_
	);
	LUT3 #(
		.INIT('h15)
	) name896 (
		_w1189_,
		_w1352_,
		_w1356_,
		_w1359_
	);
	LUT2 #(
		.INIT('h1)
	) name897 (
		\P2_B_reg/NET0131 ,
		_w1354_,
		_w1360_
	);
	LUT3 #(
		.INIT('ha2)
	) name898 (
		_w1355_,
		_w1352_,
		_w1360_,
		_w1361_
	);
	LUT4 #(
		.INIT('h0082)
	) name899 (
		\P2_B_reg/NET0131 ,
		\P2_IR_reg[24]/NET0131 ,
		_w534_,
		_w1354_,
		_w1362_
	);
	LUT3 #(
		.INIT('hc8)
	) name900 (
		\P2_d_reg[0]/NET0131 ,
		_w1352_,
		_w1362_,
		_w1363_
	);
	LUT2 #(
		.INIT('he)
	) name901 (
		_w1361_,
		_w1363_,
		_w1364_
	);
	LUT4 #(
		.INIT('h0096)
	) name902 (
		\P2_B_reg/NET0131 ,
		\P2_IR_reg[24]/NET0131 ,
		_w534_,
		_w1354_,
		_w1365_
	);
	LUT4 #(
		.INIT('h1112)
	) name903 (
		\P2_IR_reg[26]/NET0131 ,
		\P2_d_reg[1]/NET0131 ,
		_w1185_,
		_w1351_,
		_w1366_
	);
	LUT4 #(
		.INIT('h0a09)
	) name904 (
		\P2_IR_reg[26]/NET0131 ,
		_w1185_,
		_w1354_,
		_w1351_,
		_w1367_
	);
	LUT3 #(
		.INIT('h0b)
	) name905 (
		_w1365_,
		_w1366_,
		_w1367_,
		_w1368_
	);
	LUT3 #(
		.INIT('he0)
	) name906 (
		_w1361_,
		_w1363_,
		_w1368_,
		_w1369_
	);
	LUT4 #(
		.INIT('h0155)
	) name907 (
		_w1079_,
		_w1361_,
		_w1363_,
		_w1368_,
		_w1370_
	);
	LUT4 #(
		.INIT('hdd0d)
	) name908 (
		_w528_,
		_w594_,
		_w866_,
		_w879_,
		_w1371_
	);
	LUT4 #(
		.INIT('hdd0d)
	) name909 (
		_w845_,
		_w860_,
		_w910_,
		_w925_,
		_w1372_
	);
	LUT2 #(
		.INIT('h8)
	) name910 (
		_w1371_,
		_w1372_,
		_w1373_
	);
	LUT4 #(
		.INIT('h4d44)
	) name911 (
		_w747_,
		_w752_,
		_w770_,
		_w774_,
		_w1374_
	);
	LUT4 #(
		.INIT('h222a)
	) name912 (
		_w798_,
		_w809_,
		_w828_,
		_w1210_,
		_w1375_
	);
	LUT2 #(
		.INIT('h4)
	) name913 (
		_w753_,
		_w787_,
		_w1376_
	);
	LUT4 #(
		.INIT('hdd0d)
	) name914 (
		_w726_,
		_w731_,
		_w759_,
		_w763_,
		_w1377_
	);
	LUT3 #(
		.INIT('h10)
	) name915 (
		_w704_,
		_w720_,
		_w1377_,
		_w1378_
	);
	LUT4 #(
		.INIT('hba00)
	) name916 (
		_w1374_,
		_w1375_,
		_w1376_,
		_w1378_,
		_w1379_
	);
	LUT4 #(
		.INIT('h4d44)
	) name917 (
		_w726_,
		_w731_,
		_w759_,
		_w763_,
		_w1380_
	);
	LUT3 #(
		.INIT('h10)
	) name918 (
		_w704_,
		_w720_,
		_w1380_,
		_w1381_
	);
	LUT3 #(
		.INIT('h54)
	) name919 (
		_w704_,
		_w733_,
		_w734_,
		_w1382_
	);
	LUT2 #(
		.INIT('h1)
	) name920 (
		_w1381_,
		_w1382_,
		_w1383_
	);
	LUT3 #(
		.INIT('h0b)
	) name921 (
		_w615_,
		_w623_,
		_w646_,
		_w1384_
	);
	LUT2 #(
		.INIT('h1)
	) name922 (
		_w687_,
		_w737_,
		_w1385_
	);
	LUT2 #(
		.INIT('h8)
	) name923 (
		_w1384_,
		_w1385_,
		_w1386_
	);
	LUT4 #(
		.INIT('h8a00)
	) name924 (
		_w1373_,
		_w1379_,
		_w1383_,
		_w1386_,
		_w1387_
	);
	LUT3 #(
		.INIT('h51)
	) name925 (
		_w667_,
		_w686_,
		_w737_,
		_w1388_
	);
	LUT3 #(
		.INIT('hb2)
	) name926 (
		_w615_,
		_w623_,
		_w647_,
		_w1389_
	);
	LUT3 #(
		.INIT('h0d)
	) name927 (
		_w1384_,
		_w1388_,
		_w1389_,
		_w1390_
	);
	LUT4 #(
		.INIT('h4f04)
	) name928 (
		_w528_,
		_w594_,
		_w866_,
		_w879_,
		_w1391_
	);
	LUT4 #(
		.INIT('h4f04)
	) name929 (
		_w845_,
		_w860_,
		_w910_,
		_w925_,
		_w1392_
	);
	LUT3 #(
		.INIT('h07)
	) name930 (
		_w1372_,
		_w1391_,
		_w1392_,
		_w1393_
	);
	LUT3 #(
		.INIT('hd0)
	) name931 (
		_w1373_,
		_w1390_,
		_w1393_,
		_w1394_
	);
	LUT2 #(
		.INIT('h1)
	) name932 (
		_w1010_,
		_w1013_,
		_w1395_
	);
	LUT4 #(
		.INIT('h0001)
	) name933 (
		_w929_,
		_w1010_,
		_w1013_,
		_w1014_,
		_w1396_
	);
	LUT4 #(
		.INIT('h3233)
	) name934 (
		_w546_,
		_w1011_,
		_w1041_,
		_w1047_,
		_w1397_
	);
	LUT3 #(
		.INIT('h10)
	) name935 (
		_w1091_,
		_w1094_,
		_w1397_,
		_w1398_
	);
	LUT4 #(
		.INIT('h1000)
	) name936 (
		_w1091_,
		_w1094_,
		_w1396_,
		_w1397_,
		_w1399_
	);
	LUT3 #(
		.INIT('hb0)
	) name937 (
		_w1387_,
		_w1394_,
		_w1399_,
		_w1400_
	);
	LUT3 #(
		.INIT('h31)
	) name938 (
		_w903_,
		_w971_,
		_w1014_,
		_w1401_
	);
	LUT3 #(
		.INIT('h0e)
	) name939 (
		_w955_,
		_w1008_,
		_w1010_,
		_w1402_
	);
	LUT3 #(
		.INIT('h0d)
	) name940 (
		_w1395_,
		_w1401_,
		_w1402_,
		_w1403_
	);
	LUT4 #(
		.INIT('h3701)
	) name941 (
		_w546_,
		_w991_,
		_w1041_,
		_w1047_,
		_w1404_
	);
	LUT3 #(
		.INIT('h01)
	) name942 (
		_w1091_,
		_w1094_,
		_w1404_,
		_w1405_
	);
	LUT3 #(
		.INIT('h0e)
	) name943 (
		_w1037_,
		_w1071_,
		_w1091_,
		_w1406_
	);
	LUT4 #(
		.INIT('h0031)
	) name944 (
		_w1398_,
		_w1405_,
		_w1403_,
		_w1406_,
		_w1407_
	);
	LUT4 #(
		.INIT('h8488)
	) name945 (
		_w1263_,
		_w1369_,
		_w1400_,
		_w1407_,
		_w1408_
	);
	LUT4 #(
		.INIT('hfcaf)
	) name946 (
		_w1179_,
		_w1183_,
		_w1186_,
		_w1189_,
		_w1409_
	);
	LUT3 #(
		.INIT('h0e)
	) name947 (
		_w1370_,
		_w1408_,
		_w1409_,
		_w1410_
	);
	LUT3 #(
		.INIT('h01)
	) name948 (
		_w1361_,
		_w1363_,
		_w1368_,
		_w1411_
	);
	LUT4 #(
		.INIT('h5554)
	) name949 (
		_w1079_,
		_w1361_,
		_w1363_,
		_w1368_,
		_w1412_
	);
	LUT3 #(
		.INIT('h45)
	) name950 (
		_w823_,
		_w1110_,
		_w1137_,
		_w1413_
	);
	LUT4 #(
		.INIT('h1011)
	) name951 (
		_w814_,
		_w823_,
		_w1110_,
		_w1137_,
		_w1414_
	);
	LUT4 #(
		.INIT('h0001)
	) name952 (
		_w747_,
		_w770_,
		_w781_,
		_w792_,
		_w1415_
	);
	LUT3 #(
		.INIT('h40)
	) name953 (
		_w803_,
		_w1414_,
		_w1415_,
		_w1416_
	);
	LUT2 #(
		.INIT('h1)
	) name954 (
		_w726_,
		_w759_,
		_w1417_
	);
	LUT4 #(
		.INIT('h4000)
	) name955 (
		_w803_,
		_w1414_,
		_w1415_,
		_w1417_,
		_w1418_
	);
	LUT4 #(
		.INIT('h0001)
	) name956 (
		_w653_,
		_w679_,
		_w693_,
		_w711_,
		_w1419_
	);
	LUT3 #(
		.INIT('h40)
	) name957 (
		_w631_,
		_w1418_,
		_w1419_,
		_w1420_
	);
	LUT3 #(
		.INIT('h15)
	) name958 (
		_w528_,
		_w618_,
		_w622_,
		_w1421_
	);
	LUT4 #(
		.INIT('h0015)
	) name959 (
		_w528_,
		_w618_,
		_w622_,
		_w866_,
		_w1422_
	);
	LUT4 #(
		.INIT('h4000)
	) name960 (
		_w631_,
		_w1418_,
		_w1419_,
		_w1422_,
		_w1423_
	);
	LUT4 #(
		.INIT('h7077)
	) name961 (
		_w883_,
		_w888_,
		_w964_,
		_w968_,
		_w1424_
	);
	LUT4 #(
		.INIT('h7077)
	) name962 (
		_w906_,
		_w909_,
		_w948_,
		_w952_,
		_w1425_
	);
	LUT2 #(
		.INIT('h8)
	) name963 (
		_w1424_,
		_w1425_,
		_w1426_
	);
	LUT3 #(
		.INIT('h45)
	) name964 (
		_w845_,
		_w1001_,
		_w1005_,
		_w1427_
	);
	LUT4 #(
		.INIT('h4000)
	) name965 (
		_w989_,
		_w1424_,
		_w1425_,
		_w1427_,
		_w1428_
	);
	LUT2 #(
		.INIT('h4)
	) name966 (
		_w1047_,
		_w1428_,
		_w1429_
	);
	LUT4 #(
		.INIT('h0045)
	) name967 (
		_w1035_,
		_w1064_,
		_w1068_,
		_w1085_,
		_w1430_
	);
	LUT3 #(
		.INIT('h80)
	) name968 (
		_w1423_,
		_w1429_,
		_w1430_,
		_w1431_
	);
	LUT4 #(
		.INIT('h4000)
	) name969 (
		_w1131_,
		_w1423_,
		_w1429_,
		_w1430_,
		_w1432_
	);
	LUT2 #(
		.INIT('h2)
	) name970 (
		_w537_,
		_w545_,
		_w1433_
	);
	LUT2 #(
		.INIT('h4)
	) name971 (
		_w537_,
		_w545_,
		_w1434_
	);
	LUT2 #(
		.INIT('h9)
	) name972 (
		_w537_,
		_w545_,
		_w1435_
	);
	LUT3 #(
		.INIT('h0b)
	) name973 (
		_w1064_,
		_w1068_,
		_w1435_,
		_w1436_
	);
	LUT4 #(
		.INIT('h006f)
	) name974 (
		_w1131_,
		_w1431_,
		_w1435_,
		_w1436_,
		_w1437_
	);
	LUT4 #(
		.INIT('h04c4)
	) name975 (
		_w1079_,
		_w1191_,
		_w1411_,
		_w1437_,
		_w1438_
	);
	LUT4 #(
		.INIT('h0155)
	) name976 (
		_w1229_,
		_w1361_,
		_w1363_,
		_w1368_,
		_w1439_
	);
	LUT2 #(
		.INIT('h2)
	) name977 (
		_w1232_,
		_w1439_,
		_w1440_
	);
	LUT2 #(
		.INIT('h4)
	) name978 (
		_w1184_,
		_w1190_,
		_w1441_
	);
	LUT2 #(
		.INIT('h4)
	) name979 (
		_w1229_,
		_w1232_,
		_w1442_
	);
	LUT4 #(
		.INIT('h1f00)
	) name980 (
		_w1361_,
		_w1363_,
		_w1368_,
		_w1442_,
		_w1443_
	);
	LUT3 #(
		.INIT('h54)
	) name981 (
		_w1079_,
		_w1441_,
		_w1443_,
		_w1444_
	);
	LUT4 #(
		.INIT('h00ef)
	) name982 (
		_w546_,
		_w1078_,
		_w1440_,
		_w1444_,
		_w1445_
	);
	LUT2 #(
		.INIT('h4)
	) name983 (
		_w1438_,
		_w1445_,
		_w1446_
	);
	LUT3 #(
		.INIT('h80)
	) name984 (
		_w1179_,
		_w1183_,
		_w1228_,
		_w1447_
	);
	LUT4 #(
		.INIT('h0777)
	) name985 (
		_w845_,
		_w860_,
		_w910_,
		_w925_,
		_w1448_
	);
	LUT4 #(
		.INIT('h0777)
	) name986 (
		_w528_,
		_w594_,
		_w866_,
		_w879_,
		_w1449_
	);
	LUT2 #(
		.INIT('h8)
	) name987 (
		_w1448_,
		_w1449_,
		_w1450_
	);
	LUT2 #(
		.INIT('h1)
	) name988 (
		_w803_,
		_w807_,
		_w1451_
	);
	LUT4 #(
		.INIT('heee8)
	) name989 (
		_w814_,
		_w818_,
		_w823_,
		_w826_,
		_w1452_
	);
	LUT4 #(
		.INIT('h0777)
	) name990 (
		_w792_,
		_w797_,
		_w803_,
		_w807_,
		_w1453_
	);
	LUT4 #(
		.INIT('h4500)
	) name991 (
		_w1324_,
		_w1451_,
		_w1452_,
		_w1453_,
		_w1454_
	);
	LUT4 #(
		.INIT('h1117)
	) name992 (
		_w781_,
		_w785_,
		_w792_,
		_w797_,
		_w1455_
	);
	LUT4 #(
		.INIT('h0777)
	) name993 (
		_w747_,
		_w752_,
		_w770_,
		_w774_,
		_w1456_
	);
	LUT4 #(
		.INIT('heee8)
	) name994 (
		_w747_,
		_w752_,
		_w770_,
		_w774_,
		_w1457_
	);
	LUT4 #(
		.INIT('h1f00)
	) name995 (
		_w1454_,
		_w1455_,
		_w1456_,
		_w1457_,
		_w1458_
	);
	LUT3 #(
		.INIT('h02)
	) name996 (
		_w711_,
		_w716_,
		_w718_,
		_w1459_
	);
	LUT4 #(
		.INIT('h0777)
	) name997 (
		_w726_,
		_w731_,
		_w759_,
		_w763_,
		_w1460_
	);
	LUT3 #(
		.INIT('h10)
	) name998 (
		_w1316_,
		_w1459_,
		_w1460_,
		_w1461_
	);
	LUT4 #(
		.INIT('h1117)
	) name999 (
		_w726_,
		_w731_,
		_w759_,
		_w763_,
		_w1462_
	);
	LUT3 #(
		.INIT('h10)
	) name1000 (
		_w1316_,
		_w1459_,
		_w1462_,
		_w1463_
	);
	LUT3 #(
		.INIT('h54)
	) name1001 (
		_w711_,
		_w716_,
		_w718_,
		_w1464_
	);
	LUT3 #(
		.INIT('h45)
	) name1002 (
		_w1315_,
		_w1316_,
		_w1464_,
		_w1465_
	);
	LUT2 #(
		.INIT('h4)
	) name1003 (
		_w1463_,
		_w1465_,
		_w1466_
	);
	LUT4 #(
		.INIT('h00c8)
	) name1004 (
		_w546_,
		_w631_,
		_w642_,
		_w644_,
		_w1467_
	);
	LUT3 #(
		.INIT('h07)
	) name1005 (
		_w615_,
		_w623_,
		_w1467_,
		_w1468_
	);
	LUT2 #(
		.INIT('h1)
	) name1006 (
		_w1318_,
		_w1300_,
		_w1469_
	);
	LUT2 #(
		.INIT('h8)
	) name1007 (
		_w1468_,
		_w1469_,
		_w1470_
	);
	LUT4 #(
		.INIT('h4f00)
	) name1008 (
		_w1458_,
		_w1461_,
		_w1466_,
		_w1470_,
		_w1471_
	);
	LUT3 #(
		.INIT('h0d)
	) name1009 (
		_w1319_,
		_w1300_,
		_w1301_,
		_w1472_
	);
	LUT4 #(
		.INIT('h3301)
	) name1010 (
		_w546_,
		_w631_,
		_w642_,
		_w644_,
		_w1473_
	);
	LUT3 #(
		.INIT('h8e)
	) name1011 (
		_w615_,
		_w623_,
		_w1473_,
		_w1474_
	);
	LUT3 #(
		.INIT('hd0)
	) name1012 (
		_w1468_,
		_w1472_,
		_w1474_,
		_w1475_
	);
	LUT4 #(
		.INIT('hfee0)
	) name1013 (
		_w528_,
		_w594_,
		_w866_,
		_w879_,
		_w1476_
	);
	LUT4 #(
		.INIT('hfee0)
	) name1014 (
		_w845_,
		_w860_,
		_w910_,
		_w925_,
		_w1477_
	);
	LUT3 #(
		.INIT('hd0)
	) name1015 (
		_w1448_,
		_w1476_,
		_w1477_,
		_w1478_
	);
	LUT3 #(
		.INIT('hd0)
	) name1016 (
		_w1450_,
		_w1475_,
		_w1478_,
		_w1479_
	);
	LUT4 #(
		.INIT('h001f)
	) name1017 (
		_w546_,
		_w1041_,
		_w1047_,
		_w1277_,
		_w1480_
	);
	LUT2 #(
		.INIT('h4)
	) name1018 (
		_w1269_,
		_w1480_,
		_w1481_
	);
	LUT2 #(
		.INIT('h1)
	) name1019 (
		_w1282_,
		_w1273_,
		_w1482_
	);
	LUT4 #(
		.INIT('h00c8)
	) name1020 (
		_w546_,
		_w889_,
		_w899_,
		_w901_,
		_w1483_
	);
	LUT4 #(
		.INIT('h0001)
	) name1021 (
		_w1287_,
		_w1282_,
		_w1273_,
		_w1483_,
		_w1484_
	);
	LUT4 #(
		.INIT('h1000)
	) name1022 (
		_w1255_,
		_w1269_,
		_w1480_,
		_w1484_,
		_w1485_
	);
	LUT4 #(
		.INIT('h8f00)
	) name1023 (
		_w1450_,
		_w1471_,
		_w1479_,
		_w1485_,
		_w1486_
	);
	LUT4 #(
		.INIT('h3301)
	) name1024 (
		_w546_,
		_w889_,
		_w899_,
		_w901_,
		_w1487_
	);
	LUT3 #(
		.INIT('h23)
	) name1025 (
		_w1287_,
		_w1288_,
		_w1487_,
		_w1488_
	);
	LUT3 #(
		.INIT('h0d)
	) name1026 (
		_w1281_,
		_w1273_,
		_w1274_,
		_w1489_
	);
	LUT3 #(
		.INIT('hd0)
	) name1027 (
		_w1482_,
		_w1488_,
		_w1489_,
		_w1490_
	);
	LUT4 #(
		.INIT('he0fe)
	) name1028 (
		_w546_,
		_w1041_,
		_w1047_,
		_w1276_,
		_w1491_
	);
	LUT4 #(
		.INIT('h0d04)
	) name1029 (
		_w1027_,
		_w1035_,
		_w1256_,
		_w1491_,
		_w1492_
	);
	LUT4 #(
		.INIT('h0455)
	) name1030 (
		_w1255_,
		_w1481_,
		_w1490_,
		_w1492_,
		_w1493_
	);
	LUT4 #(
		.INIT('h4448)
	) name1031 (
		_w1263_,
		_w1411_,
		_w1486_,
		_w1493_,
		_w1494_
	);
	LUT3 #(
		.INIT('ha8)
	) name1032 (
		_w1447_,
		_w1412_,
		_w1494_,
		_w1495_
	);
	LUT4 #(
		.INIT('hc7f7)
	) name1033 (
		_w1179_,
		_w1186_,
		_w1189_,
		_w1229_,
		_w1496_
	);
	LUT4 #(
		.INIT('h4448)
	) name1034 (
		_w1263_,
		_w1369_,
		_w1486_,
		_w1493_,
		_w1497_
	);
	LUT3 #(
		.INIT('h32)
	) name1035 (
		_w1370_,
		_w1496_,
		_w1497_,
		_w1498_
	);
	LUT4 #(
		.INIT('h0100)
	) name1036 (
		_w1410_,
		_w1495_,
		_w1498_,
		_w1446_,
		_w1499_
	);
	LUT4 #(
		.INIT('h88a8)
	) name1037 (
		\P1_state_reg[0]/NET0131 ,
		_w1358_,
		_w1359_,
		_w1499_,
		_w1500_
	);
	LUT4 #(
		.INIT('h93bb)
	) name1038 (
		\P1_state_reg[0]/NET0131 ,
		\P2_reg3_reg[27]/NET0131 ,
		_w1062_,
		_w1189_,
		_w1501_
	);
	LUT2 #(
		.INIT('hb)
	) name1039 (
		_w1500_,
		_w1501_,
		_w1502_
	);
	LUT3 #(
		.INIT('h28)
	) name1040 (
		\P1_state_reg[0]/NET0131 ,
		\P2_IR_reg[23]/NET0131 ,
		_w1188_,
		_w1503_
	);
	LUT4 #(
		.INIT('hd070)
	) name1041 (
		\P1_state_reg[0]/NET0131 ,
		\P2_IR_reg[23]/NET0131 ,
		\P2_reg2_reg[28]/NET0131 ,
		_w1188_,
		_w1504_
	);
	LUT4 #(
		.INIT('h2000)
	) name1042 (
		\P2_reg2_reg[28]/NET0131 ,
		_w1189_,
		_w1352_,
		_w1356_,
		_w1505_
	);
	LUT4 #(
		.INIT('hfeaf)
	) name1043 (
		_w1179_,
		_w1183_,
		_w1186_,
		_w1189_,
		_w1506_
	);
	LUT3 #(
		.INIT('h10)
	) name1044 (
		_w1361_,
		_w1363_,
		_w1368_,
		_w1507_
	);
	LUT3 #(
		.INIT('hb0)
	) name1045 (
		_w1215_,
		_w1216_,
		_w1205_,
		_w1508_
	);
	LUT2 #(
		.INIT('h8)
	) name1046 (
		_w1201_,
		_w1202_,
		_w1509_
	);
	LUT4 #(
		.INIT('h000b)
	) name1047 (
		_w673_,
		_w1201_,
		_w1198_,
		_w1199_,
		_w1510_
	);
	LUT3 #(
		.INIT('hb0)
	) name1048 (
		_w1508_,
		_w1509_,
		_w1510_,
		_w1511_
	);
	LUT2 #(
		.INIT('h8)
	) name1049 (
		_w1195_,
		_w1196_,
		_w1512_
	);
	LUT2 #(
		.INIT('h2)
	) name1050 (
		_w1195_,
		_w1220_,
		_w1513_
	);
	LUT4 #(
		.INIT('h0045)
	) name1051 (
		_w1224_,
		_w1511_,
		_w1512_,
		_w1513_,
		_w1514_
	);
	LUT4 #(
		.INIT('hc535)
	) name1052 (
		\P2_reg2_reg[28]/NET0131 ,
		_w1260_,
		_w1507_,
		_w1514_,
		_w1515_
	);
	LUT3 #(
		.INIT('h0e)
	) name1053 (
		_w1361_,
		_w1363_,
		_w1368_,
		_w1516_
	);
	LUT3 #(
		.INIT('h0b)
	) name1054 (
		_w1080_,
		_w1084_,
		_w1435_,
		_w1517_
	);
	LUT4 #(
		.INIT('hb0bb)
	) name1055 (
		_w1110_,
		_w1114_,
		_w1126_,
		_w1130_,
		_w1518_
	);
	LUT4 #(
		.INIT('h8000)
	) name1056 (
		_w1423_,
		_w1429_,
		_w1430_,
		_w1518_,
		_w1519_
	);
	LUT4 #(
		.INIT('h00d0)
	) name1057 (
		_w1115_,
		_w1432_,
		_w1435_,
		_w1519_,
		_w1520_
	);
	LUT4 #(
		.INIT('h111d)
	) name1058 (
		\P2_reg2_reg[28]/NET0131 ,
		_w1516_,
		_w1517_,
		_w1520_,
		_w1521_
	);
	LUT4 #(
		.INIT('h1000)
	) name1059 (
		_w1361_,
		_w1363_,
		_w1368_,
		_w1442_,
		_w1522_
	);
	LUT4 #(
		.INIT('hef00)
	) name1060 (
		_w1361_,
		_w1363_,
		_w1368_,
		_w1442_,
		_w1523_
	);
	LUT2 #(
		.INIT('h4)
	) name1061 (
		_w1125_,
		_w1233_,
		_w1524_
	);
	LUT4 #(
		.INIT('h0057)
	) name1062 (
		\P2_reg2_reg[28]/NET0131 ,
		_w1441_,
		_w1523_,
		_w1524_,
		_w1525_
	);
	LUT4 #(
		.INIT('hef00)
	) name1063 (
		_w546_,
		_w1124_,
		_w1522_,
		_w1525_,
		_w1526_
	);
	LUT3 #(
		.INIT('hd0)
	) name1064 (
		_w1191_,
		_w1521_,
		_w1526_,
		_w1527_
	);
	LUT3 #(
		.INIT('he0)
	) name1065 (
		_w1506_,
		_w1515_,
		_w1527_,
		_w1528_
	);
	LUT4 #(
		.INIT('hc355)
	) name1066 (
		\P2_reg2_reg[28]/NET0131 ,
		_w1260_,
		_w1514_,
		_w1516_,
		_w1529_
	);
	LUT3 #(
		.INIT('h20)
	) name1067 (
		_w1179_,
		_w1183_,
		_w1228_,
		_w1530_
	);
	LUT4 #(
		.INIT('h0777)
	) name1068 (
		_w747_,
		_w752_,
		_w759_,
		_w763_,
		_w1531_
	);
	LUT4 #(
		.INIT('h1117)
	) name1069 (
		_w792_,
		_w797_,
		_w803_,
		_w807_,
		_w1532_
	);
	LUT4 #(
		.INIT('h0777)
	) name1070 (
		_w770_,
		_w774_,
		_w781_,
		_w785_,
		_w1533_
	);
	LUT4 #(
		.INIT('hf400)
	) name1071 (
		_w1452_,
		_w1453_,
		_w1532_,
		_w1533_,
		_w1534_
	);
	LUT4 #(
		.INIT('heee8)
	) name1072 (
		_w770_,
		_w774_,
		_w781_,
		_w785_,
		_w1535_
	);
	LUT4 #(
		.INIT('hfee0)
	) name1073 (
		_w747_,
		_w752_,
		_w759_,
		_w763_,
		_w1536_
	);
	LUT4 #(
		.INIT('h7500)
	) name1074 (
		_w1531_,
		_w1534_,
		_w1535_,
		_w1536_,
		_w1537_
	);
	LUT2 #(
		.INIT('h1)
	) name1075 (
		_w1318_,
		_w1316_,
		_w1538_
	);
	LUT4 #(
		.INIT('h0001)
	) name1076 (
		_w1318_,
		_w1316_,
		_w1308_,
		_w1459_,
		_w1539_
	);
	LUT2 #(
		.INIT('h4)
	) name1077 (
		_w1537_,
		_w1539_,
		_w1540_
	);
	LUT3 #(
		.INIT('h32)
	) name1078 (
		_w1309_,
		_w1459_,
		_w1464_,
		_w1541_
	);
	LUT3 #(
		.INIT('h23)
	) name1079 (
		_w1318_,
		_w1319_,
		_w1315_,
		_w1542_
	);
	LUT3 #(
		.INIT('h70)
	) name1080 (
		_w1538_,
		_w1541_,
		_w1542_,
		_w1543_
	);
	LUT3 #(
		.INIT('hb0)
	) name1081 (
		_w1537_,
		_w1539_,
		_w1543_,
		_w1544_
	);
	LUT4 #(
		.INIT('h0777)
	) name1082 (
		_w528_,
		_w594_,
		_w615_,
		_w623_,
		_w1545_
	);
	LUT2 #(
		.INIT('h1)
	) name1083 (
		_w1300_,
		_w1467_,
		_w1546_
	);
	LUT2 #(
		.INIT('h8)
	) name1084 (
		_w1545_,
		_w1546_,
		_w1547_
	);
	LUT4 #(
		.INIT('h0777)
	) name1085 (
		_w845_,
		_w860_,
		_w866_,
		_w879_,
		_w1548_
	);
	LUT3 #(
		.INIT('h10)
	) name1086 (
		_w1290_,
		_w1483_,
		_w1548_,
		_w1549_
	);
	LUT2 #(
		.INIT('h8)
	) name1087 (
		_w1547_,
		_w1549_,
		_w1550_
	);
	LUT3 #(
		.INIT('h32)
	) name1088 (
		_w1301_,
		_w1467_,
		_w1473_,
		_w1551_
	);
	LUT4 #(
		.INIT('heee8)
	) name1089 (
		_w528_,
		_w594_,
		_w615_,
		_w623_,
		_w1552_
	);
	LUT3 #(
		.INIT('h70)
	) name1090 (
		_w1545_,
		_w1551_,
		_w1552_,
		_w1553_
	);
	LUT4 #(
		.INIT('heee8)
	) name1091 (
		_w845_,
		_w860_,
		_w866_,
		_w879_,
		_w1554_
	);
	LUT3 #(
		.INIT('h01)
	) name1092 (
		_w1290_,
		_w1483_,
		_w1554_,
		_w1555_
	);
	LUT3 #(
		.INIT('h32)
	) name1093 (
		_w1291_,
		_w1483_,
		_w1487_,
		_w1556_
	);
	LUT2 #(
		.INIT('h1)
	) name1094 (
		_w1555_,
		_w1556_,
		_w1557_
	);
	LUT4 #(
		.INIT('h000d)
	) name1095 (
		_w1549_,
		_w1553_,
		_w1555_,
		_w1556_,
		_w1558_
	);
	LUT3 #(
		.INIT('hb0)
	) name1096 (
		_w1544_,
		_w1550_,
		_w1558_,
		_w1559_
	);
	LUT2 #(
		.INIT('h1)
	) name1097 (
		_w1255_,
		_w1262_,
		_w1560_
	);
	LUT4 #(
		.INIT('h0001)
	) name1098 (
		_w1255_,
		_w1262_,
		_w1269_,
		_w1266_,
		_w1561_
	);
	LUT2 #(
		.INIT('h1)
	) name1099 (
		_w1287_,
		_w1282_,
		_w1562_
	);
	LUT2 #(
		.INIT('h1)
	) name1100 (
		_w1273_,
		_w1277_,
		_w1563_
	);
	LUT4 #(
		.INIT('h0001)
	) name1101 (
		_w1287_,
		_w1282_,
		_w1273_,
		_w1277_,
		_w1564_
	);
	LUT2 #(
		.INIT('h8)
	) name1102 (
		_w1561_,
		_w1564_,
		_w1565_
	);
	LUT3 #(
		.INIT('h31)
	) name1103 (
		_w1288_,
		_w1281_,
		_w1282_,
		_w1566_
	);
	LUT3 #(
		.INIT('h31)
	) name1104 (
		_w1274_,
		_w1276_,
		_w1277_,
		_w1567_
	);
	LUT3 #(
		.INIT('hd0)
	) name1105 (
		_w1563_,
		_w1566_,
		_w1567_,
		_w1568_
	);
	LUT2 #(
		.INIT('h2)
	) name1106 (
		_w1561_,
		_w1568_,
		_w1569_
	);
	LUT3 #(
		.INIT('h23)
	) name1107 (
		_w1269_,
		_w1270_,
		_w1267_,
		_w1570_
	);
	LUT3 #(
		.INIT('h31)
	) name1108 (
		_w1256_,
		_w1261_,
		_w1262_,
		_w1571_
	);
	LUT3 #(
		.INIT('hd0)
	) name1109 (
		_w1560_,
		_w1570_,
		_w1571_,
		_w1572_
	);
	LUT4 #(
		.INIT('h0b00)
	) name1110 (
		_w1559_,
		_w1565_,
		_w1569_,
		_w1572_,
		_w1573_
	);
	LUT4 #(
		.INIT('h35c5)
	) name1111 (
		\P2_reg2_reg[28]/NET0131 ,
		_w1260_,
		_w1507_,
		_w1573_,
		_w1574_
	);
	LUT4 #(
		.INIT('hf35f)
	) name1112 (
		_w1179_,
		_w1183_,
		_w1186_,
		_w1189_,
		_w1575_
	);
	LUT4 #(
		.INIT('hbbb0)
	) name1113 (
		_w1529_,
		_w1530_,
		_w1574_,
		_w1575_,
		_w1576_
	);
	LUT4 #(
		.INIT('h3111)
	) name1114 (
		_w1359_,
		_w1505_,
		_w1528_,
		_w1576_,
		_w1577_
	);
	LUT3 #(
		.INIT('hce)
	) name1115 (
		\P1_state_reg[0]/NET0131 ,
		_w1504_,
		_w1577_,
		_w1578_
	);
	LUT2 #(
		.INIT('h4)
	) name1116 (
		_w1125_,
		_w1357_,
		_w1579_
	);
	LUT4 #(
		.INIT('h0155)
	) name1117 (
		_w1125_,
		_w1361_,
		_w1363_,
		_w1368_,
		_w1580_
	);
	LUT4 #(
		.INIT('h00b7)
	) name1118 (
		_w1260_,
		_w1369_,
		_w1514_,
		_w1580_,
		_w1581_
	);
	LUT4 #(
		.INIT('h5554)
	) name1119 (
		_w1125_,
		_w1361_,
		_w1363_,
		_w1368_,
		_w1582_
	);
	LUT4 #(
		.INIT('h0057)
	) name1120 (
		_w1411_,
		_w1517_,
		_w1520_,
		_w1582_,
		_w1583_
	);
	LUT3 #(
		.INIT('h54)
	) name1121 (
		_w1125_,
		_w1441_,
		_w1443_,
		_w1584_
	);
	LUT4 #(
		.INIT('h00ef)
	) name1122 (
		_w546_,
		_w1124_,
		_w1440_,
		_w1584_,
		_w1585_
	);
	LUT3 #(
		.INIT('hd0)
	) name1123 (
		_w1191_,
		_w1583_,
		_w1585_,
		_w1586_
	);
	LUT3 #(
		.INIT('he0)
	) name1124 (
		_w1409_,
		_w1581_,
		_w1586_,
		_w1587_
	);
	LUT4 #(
		.INIT('h007b)
	) name1125 (
		_w1260_,
		_w1411_,
		_w1573_,
		_w1582_,
		_w1588_
	);
	LUT4 #(
		.INIT('h007b)
	) name1126 (
		_w1260_,
		_w1369_,
		_w1573_,
		_w1580_,
		_w1589_
	);
	LUT4 #(
		.INIT('hf5c4)
	) name1127 (
		_w1447_,
		_w1496_,
		_w1588_,
		_w1589_,
		_w1590_
	);
	LUT4 #(
		.INIT('h3111)
	) name1128 (
		_w1359_,
		_w1579_,
		_w1587_,
		_w1590_,
		_w1591_
	);
	LUT2 #(
		.INIT('h4)
	) name1129 (
		\P1_state_reg[0]/NET0131 ,
		\P2_reg3_reg[28]/NET0131 ,
		_w1592_
	);
	LUT4 #(
		.INIT('h9c00)
	) name1130 (
		\P2_reg3_reg[27]/NET0131 ,
		\P2_reg3_reg[28]/NET0131 ,
		_w1062_,
		_w1349_,
		_w1593_
	);
	LUT2 #(
		.INIT('h1)
	) name1131 (
		_w1592_,
		_w1593_,
		_w1594_
	);
	LUT3 #(
		.INIT('h2f)
	) name1132 (
		\P1_state_reg[0]/NET0131 ,
		_w1591_,
		_w1594_,
		_w1595_
	);
	LUT4 #(
		.INIT('hd070)
	) name1133 (
		\P1_state_reg[0]/NET0131 ,
		\P2_IR_reg[23]/NET0131 ,
		\P2_reg2_reg[27]/NET0131 ,
		_w1188_,
		_w1596_
	);
	LUT4 #(
		.INIT('h2000)
	) name1134 (
		\P2_reg2_reg[27]/NET0131 ,
		_w1189_,
		_w1352_,
		_w1356_,
		_w1597_
	);
	LUT4 #(
		.INIT('ha8aa)
	) name1135 (
		\P2_reg2_reg[27]/NET0131 ,
		_w1361_,
		_w1363_,
		_w1368_,
		_w1598_
	);
	LUT4 #(
		.INIT('h9a00)
	) name1136 (
		_w1263_,
		_w1400_,
		_w1407_,
		_w1507_,
		_w1599_
	);
	LUT3 #(
		.INIT('h54)
	) name1137 (
		_w1506_,
		_w1598_,
		_w1599_,
		_w1600_
	);
	LUT4 #(
		.INIT('haa02)
	) name1138 (
		\P2_reg2_reg[27]/NET0131 ,
		_w1361_,
		_w1363_,
		_w1368_,
		_w1601_
	);
	LUT4 #(
		.INIT('h0c88)
	) name1139 (
		\P2_reg2_reg[27]/NET0131 ,
		_w1191_,
		_w1437_,
		_w1516_,
		_w1602_
	);
	LUT4 #(
		.INIT('h6000)
	) name1140 (
		\P2_reg3_reg[27]/NET0131 ,
		_w1062_,
		_w1229_,
		_w1232_,
		_w1603_
	);
	LUT4 #(
		.INIT('h0057)
	) name1141 (
		\P2_reg2_reg[27]/NET0131 ,
		_w1441_,
		_w1523_,
		_w1603_,
		_w1604_
	);
	LUT4 #(
		.INIT('hef00)
	) name1142 (
		_w546_,
		_w1078_,
		_w1522_,
		_w1604_,
		_w1605_
	);
	LUT2 #(
		.INIT('h4)
	) name1143 (
		_w1602_,
		_w1605_,
		_w1606_
	);
	LUT4 #(
		.INIT('h5600)
	) name1144 (
		_w1263_,
		_w1486_,
		_w1493_,
		_w1507_,
		_w1607_
	);
	LUT3 #(
		.INIT('h54)
	) name1145 (
		_w1575_,
		_w1598_,
		_w1607_,
		_w1608_
	);
	LUT4 #(
		.INIT('h9a00)
	) name1146 (
		_w1263_,
		_w1400_,
		_w1407_,
		_w1516_,
		_w1609_
	);
	LUT3 #(
		.INIT('ha8)
	) name1147 (
		_w1530_,
		_w1601_,
		_w1609_,
		_w1610_
	);
	LUT4 #(
		.INIT('h0100)
	) name1148 (
		_w1600_,
		_w1608_,
		_w1610_,
		_w1606_,
		_w1611_
	);
	LUT4 #(
		.INIT('ha0a8)
	) name1149 (
		\P1_state_reg[0]/NET0131 ,
		_w1359_,
		_w1597_,
		_w1611_,
		_w1612_
	);
	LUT2 #(
		.INIT('he)
	) name1150 (
		_w1596_,
		_w1612_,
		_w1613_
	);
	LUT2 #(
		.INIT('h4)
	) name1151 (
		_w1042_,
		_w1357_,
		_w1614_
	);
	LUT4 #(
		.INIT('h0155)
	) name1152 (
		_w1042_,
		_w1361_,
		_w1363_,
		_w1368_,
		_w1615_
	);
	LUT4 #(
		.INIT('hb400)
	) name1153 (
		_w1208_,
		_w1221_,
		_w1268_,
		_w1369_,
		_w1616_
	);
	LUT3 #(
		.INIT('h54)
	) name1154 (
		_w1409_,
		_w1615_,
		_w1616_,
		_w1617_
	);
	LUT4 #(
		.INIT('h5554)
	) name1155 (
		_w1042_,
		_w1361_,
		_w1363_,
		_w1368_,
		_w1618_
	);
	LUT4 #(
		.INIT('h40f0)
	) name1156 (
		_w1543_,
		_w1547_,
		_w1549_,
		_w1553_,
		_w1619_
	);
	LUT3 #(
		.INIT('hc4)
	) name1157 (
		_w1557_,
		_w1564_,
		_w1619_,
		_w1620_
	);
	LUT3 #(
		.INIT('h80)
	) name1158 (
		_w1547_,
		_w1549_,
		_w1564_,
		_w1621_
	);
	LUT3 #(
		.INIT('h4c)
	) name1159 (
		_w1540_,
		_w1568_,
		_w1621_,
		_w1622_
	);
	LUT4 #(
		.INIT('h4844)
	) name1160 (
		_w1268_,
		_w1411_,
		_w1620_,
		_w1622_,
		_w1623_
	);
	LUT3 #(
		.INIT('ha8)
	) name1161 (
		_w1447_,
		_w1618_,
		_w1623_,
		_w1624_
	);
	LUT4 #(
		.INIT('h4844)
	) name1162 (
		_w1268_,
		_w1369_,
		_w1620_,
		_w1622_,
		_w1625_
	);
	LUT3 #(
		.INIT('h40)
	) name1163 (
		_w1035_,
		_w1423_,
		_w1429_,
		_w1626_
	);
	LUT4 #(
		.INIT('h9500)
	) name1164 (
		_w1035_,
		_w1423_,
		_w1429_,
		_w1435_,
		_w1627_
	);
	LUT3 #(
		.INIT('h0b)
	) name1165 (
		_w984_,
		_w988_,
		_w1435_,
		_w1628_
	);
	LUT4 #(
		.INIT('h1113)
	) name1166 (
		_w1411_,
		_w1618_,
		_w1627_,
		_w1628_,
		_w1629_
	);
	LUT3 #(
		.INIT('h54)
	) name1167 (
		_w1042_,
		_w1441_,
		_w1443_,
		_w1630_
	);
	LUT4 #(
		.INIT('h00ef)
	) name1168 (
		_w546_,
		_w1041_,
		_w1440_,
		_w1630_,
		_w1631_
	);
	LUT3 #(
		.INIT('hd0)
	) name1169 (
		_w1191_,
		_w1629_,
		_w1631_,
		_w1632_
	);
	LUT4 #(
		.INIT('hab00)
	) name1170 (
		_w1496_,
		_w1615_,
		_w1625_,
		_w1632_,
		_w1633_
	);
	LUT4 #(
		.INIT('ha8aa)
	) name1171 (
		_w1359_,
		_w1624_,
		_w1617_,
		_w1633_,
		_w1634_
	);
	LUT2 #(
		.INIT('h4)
	) name1172 (
		\P1_state_reg[0]/NET0131 ,
		\P2_reg3_reg[24]/NET0131 ,
		_w1635_
	);
	LUT3 #(
		.INIT('h0b)
	) name1173 (
		_w1042_,
		_w1349_,
		_w1635_,
		_w1636_
	);
	LUT4 #(
		.INIT('ha8ff)
	) name1174 (
		\P1_state_reg[0]/NET0131 ,
		_w1614_,
		_w1634_,
		_w1636_,
		_w1637_
	);
	LUT4 #(
		.INIT('hd070)
	) name1175 (
		\P1_state_reg[0]/NET0131 ,
		\P2_IR_reg[23]/NET0131 ,
		\P2_reg2_reg[24]/NET0131 ,
		_w1188_,
		_w1638_
	);
	LUT4 #(
		.INIT('h2000)
	) name1176 (
		\P2_reg2_reg[24]/NET0131 ,
		_w1189_,
		_w1352_,
		_w1356_,
		_w1639_
	);
	LUT4 #(
		.INIT('ha8aa)
	) name1177 (
		\P2_reg2_reg[24]/NET0131 ,
		_w1361_,
		_w1363_,
		_w1368_,
		_w1640_
	);
	LUT4 #(
		.INIT('hb400)
	) name1178 (
		_w1208_,
		_w1221_,
		_w1268_,
		_w1507_,
		_w1641_
	);
	LUT3 #(
		.INIT('h54)
	) name1179 (
		_w1506_,
		_w1640_,
		_w1641_,
		_w1642_
	);
	LUT4 #(
		.INIT('haa02)
	) name1180 (
		\P2_reg2_reg[24]/NET0131 ,
		_w1361_,
		_w1363_,
		_w1368_,
		_w1643_
	);
	LUT4 #(
		.INIT('hb400)
	) name1181 (
		_w1208_,
		_w1221_,
		_w1268_,
		_w1516_,
		_w1644_
	);
	LUT3 #(
		.INIT('ha8)
	) name1182 (
		_w1530_,
		_w1643_,
		_w1644_,
		_w1645_
	);
	LUT4 #(
		.INIT('h4844)
	) name1183 (
		_w1268_,
		_w1507_,
		_w1620_,
		_w1622_,
		_w1646_
	);
	LUT4 #(
		.INIT('h111d)
	) name1184 (
		\P2_reg2_reg[24]/NET0131 ,
		_w1516_,
		_w1627_,
		_w1628_,
		_w1647_
	);
	LUT2 #(
		.INIT('h4)
	) name1185 (
		_w1042_,
		_w1233_,
		_w1648_
	);
	LUT4 #(
		.INIT('h0057)
	) name1186 (
		\P2_reg2_reg[24]/NET0131 ,
		_w1441_,
		_w1523_,
		_w1648_,
		_w1649_
	);
	LUT4 #(
		.INIT('hef00)
	) name1187 (
		_w546_,
		_w1041_,
		_w1522_,
		_w1649_,
		_w1650_
	);
	LUT3 #(
		.INIT('hd0)
	) name1188 (
		_w1191_,
		_w1647_,
		_w1650_,
		_w1651_
	);
	LUT4 #(
		.INIT('hab00)
	) name1189 (
		_w1575_,
		_w1640_,
		_w1646_,
		_w1651_,
		_w1652_
	);
	LUT4 #(
		.INIT('ha8aa)
	) name1190 (
		_w1359_,
		_w1645_,
		_w1642_,
		_w1652_,
		_w1653_
	);
	LUT4 #(
		.INIT('heeec)
	) name1191 (
		\P1_state_reg[0]/NET0131 ,
		_w1638_,
		_w1639_,
		_w1653_,
		_w1654_
	);
	LUT4 #(
		.INIT('hd070)
	) name1192 (
		\P1_state_reg[0]/NET0131 ,
		\P2_IR_reg[23]/NET0131 ,
		\P2_reg0_reg[29]/NET0131 ,
		_w1188_,
		_w1655_
	);
	LUT4 #(
		.INIT('h2000)
	) name1193 (
		\P2_reg0_reg[29]/NET0131 ,
		_w1189_,
		_w1352_,
		_w1356_,
		_w1656_
	);
	LUT3 #(
		.INIT('h10)
	) name1194 (
		_w929_,
		_w1014_,
		_w1372_,
		_w1657_
	);
	LUT2 #(
		.INIT('h8)
	) name1195 (
		_w1371_,
		_w1384_,
		_w1658_
	);
	LUT2 #(
		.INIT('h8)
	) name1196 (
		_w1657_,
		_w1658_,
		_w1659_
	);
	LUT3 #(
		.INIT('h70)
	) name1197 (
		_w1382_,
		_w1385_,
		_w1388_,
		_w1660_
	);
	LUT3 #(
		.INIT('h07)
	) name1198 (
		_w1374_,
		_w1377_,
		_w1380_,
		_w1661_
	);
	LUT4 #(
		.INIT('hbf00)
	) name1199 (
		_w1375_,
		_w1376_,
		_w1377_,
		_w1661_,
		_w1662_
	);
	LUT4 #(
		.INIT('h0001)
	) name1200 (
		_w687_,
		_w704_,
		_w720_,
		_w737_,
		_w1663_
	);
	LUT3 #(
		.INIT('h8a)
	) name1201 (
		_w1660_,
		_w1662_,
		_w1663_,
		_w1664_
	);
	LUT3 #(
		.INIT('h07)
	) name1202 (
		_w1371_,
		_w1389_,
		_w1391_,
		_w1665_
	);
	LUT3 #(
		.INIT('h10)
	) name1203 (
		_w929_,
		_w1014_,
		_w1392_,
		_w1666_
	);
	LUT2 #(
		.INIT('h2)
	) name1204 (
		_w1401_,
		_w1666_,
		_w1667_
	);
	LUT4 #(
		.INIT('h00a2)
	) name1205 (
		_w1401_,
		_w1657_,
		_w1665_,
		_w1666_,
		_w1668_
	);
	LUT3 #(
		.INIT('hd0)
	) name1206 (
		_w1659_,
		_w1664_,
		_w1668_,
		_w1669_
	);
	LUT2 #(
		.INIT('h8)
	) name1207 (
		_w1395_,
		_w1397_,
		_w1670_
	);
	LUT2 #(
		.INIT('h1)
	) name1208 (
		_w1092_,
		_w1173_,
		_w1671_
	);
	LUT4 #(
		.INIT('h0001)
	) name1209 (
		_w1091_,
		_w1092_,
		_w1094_,
		_w1173_,
		_w1672_
	);
	LUT2 #(
		.INIT('h8)
	) name1210 (
		_w1670_,
		_w1672_,
		_w1673_
	);
	LUT3 #(
		.INIT('h4c)
	) name1211 (
		_w1397_,
		_w1404_,
		_w1402_,
		_w1674_
	);
	LUT2 #(
		.INIT('h2)
	) name1212 (
		_w1672_,
		_w1674_,
		_w1675_
	);
	LUT3 #(
		.INIT('h31)
	) name1213 (
		_w1087_,
		_w1133_,
		_w1173_,
		_w1676_
	);
	LUT3 #(
		.INIT('h70)
	) name1214 (
		_w1406_,
		_w1671_,
		_w1676_,
		_w1677_
	);
	LUT4 #(
		.INIT('h0b00)
	) name1215 (
		_w1669_,
		_w1673_,
		_w1675_,
		_w1677_,
		_w1678_
	);
	LUT4 #(
		.INIT('h35c5)
	) name1216 (
		\P2_reg0_reg[29]/NET0131 ,
		_w1264_,
		_w1411_,
		_w1678_,
		_w1679_
	);
	LUT3 #(
		.INIT('h0b)
	) name1217 (
		_w1126_,
		_w1130_,
		_w1435_,
		_w1680_
	);
	LUT3 #(
		.INIT('h43)
	) name1218 (
		\P2_B_reg/NET0131 ,
		_w537_,
		_w545_,
		_w1681_
	);
	LUT4 #(
		.INIT('h060f)
	) name1219 (
		_w1163_,
		_w1519_,
		_w1680_,
		_w1681_,
		_w1682_
	);
	LUT4 #(
		.INIT('h08c8)
	) name1220 (
		\P2_reg0_reg[29]/NET0131 ,
		_w1191_,
		_w1369_,
		_w1682_,
		_w1683_
	);
	LUT4 #(
		.INIT('h1b1f)
	) name1221 (
		_w1179_,
		_w1183_,
		_w1190_,
		_w1232_,
		_w1684_
	);
	LUT4 #(
		.INIT('hfe00)
	) name1222 (
		_w1361_,
		_w1363_,
		_w1368_,
		_w1442_,
		_w1685_
	);
	LUT3 #(
		.INIT('ha2)
	) name1223 (
		\P2_reg0_reg[29]/NET0131 ,
		_w1684_,
		_w1685_,
		_w1686_
	);
	LUT4 #(
		.INIT('h0100)
	) name1224 (
		_w1361_,
		_w1363_,
		_w1368_,
		_w1442_,
		_w1687_
	);
	LUT4 #(
		.INIT('h0e0f)
	) name1225 (
		_w546_,
		_w1107_,
		_w1686_,
		_w1687_,
		_w1688_
	);
	LUT2 #(
		.INIT('h4)
	) name1226 (
		_w1683_,
		_w1688_,
		_w1689_
	);
	LUT3 #(
		.INIT('he0)
	) name1227 (
		_w1409_,
		_w1679_,
		_w1689_,
		_w1690_
	);
	LUT3 #(
		.INIT('h04)
	) name1228 (
		_w1287_,
		_w1448_,
		_w1483_,
		_w1691_
	);
	LUT2 #(
		.INIT('h8)
	) name1229 (
		_w1449_,
		_w1468_,
		_w1692_
	);
	LUT2 #(
		.INIT('h8)
	) name1230 (
		_w1691_,
		_w1692_,
		_w1693_
	);
	LUT3 #(
		.INIT('hb0)
	) name1231 (
		_w1465_,
		_w1469_,
		_w1472_,
		_w1694_
	);
	LUT4 #(
		.INIT('he000)
	) name1232 (
		_w1454_,
		_w1455_,
		_w1456_,
		_w1460_,
		_w1695_
	);
	LUT3 #(
		.INIT('h0b)
	) name1233 (
		_w1457_,
		_w1460_,
		_w1462_,
		_w1696_
	);
	LUT4 #(
		.INIT('h0001)
	) name1234 (
		_w1318_,
		_w1316_,
		_w1300_,
		_w1459_,
		_w1697_
	);
	LUT3 #(
		.INIT('hb0)
	) name1235 (
		_w1695_,
		_w1696_,
		_w1697_,
		_w1698_
	);
	LUT4 #(
		.INIT('h20aa)
	) name1236 (
		_w1694_,
		_w1695_,
		_w1696_,
		_w1697_,
		_w1699_
	);
	LUT3 #(
		.INIT('hd0)
	) name1237 (
		_w1449_,
		_w1474_,
		_w1476_,
		_w1700_
	);
	LUT3 #(
		.INIT('h01)
	) name1238 (
		_w1287_,
		_w1477_,
		_w1483_,
		_w1701_
	);
	LUT2 #(
		.INIT('h2)
	) name1239 (
		_w1488_,
		_w1701_,
		_w1702_
	);
	LUT4 #(
		.INIT('h00a2)
	) name1240 (
		_w1488_,
		_w1691_,
		_w1700_,
		_w1701_,
		_w1703_
	);
	LUT3 #(
		.INIT('hd0)
	) name1241 (
		_w1693_,
		_w1699_,
		_w1703_,
		_w1704_
	);
	LUT2 #(
		.INIT('h8)
	) name1242 (
		_w1480_,
		_w1482_,
		_w1705_
	);
	LUT4 #(
		.INIT('h0001)
	) name1243 (
		_w1255_,
		_w1258_,
		_w1262_,
		_w1269_,
		_w1706_
	);
	LUT2 #(
		.INIT('h8)
	) name1244 (
		_w1705_,
		_w1706_,
		_w1707_
	);
	LUT4 #(
		.INIT('h0b02)
	) name1245 (
		_w1059_,
		_w1069_,
		_w1262_,
		_w1270_,
		_w1708_
	);
	LUT3 #(
		.INIT('h54)
	) name1246 (
		_w1258_,
		_w1261_,
		_w1708_,
		_w1709_
	);
	LUT3 #(
		.INIT('hc4)
	) name1247 (
		_w1480_,
		_w1491_,
		_w1489_,
		_w1710_
	);
	LUT3 #(
		.INIT('h51)
	) name1248 (
		_w1259_,
		_w1706_,
		_w1710_,
		_w1711_
	);
	LUT4 #(
		.INIT('h0b00)
	) name1249 (
		_w1704_,
		_w1707_,
		_w1709_,
		_w1711_,
		_w1712_
	);
	LUT4 #(
		.INIT('hc535)
	) name1250 (
		\P2_reg0_reg[29]/NET0131 ,
		_w1264_,
		_w1369_,
		_w1712_,
		_w1713_
	);
	LUT4 #(
		.INIT('hc535)
	) name1251 (
		\P2_reg0_reg[29]/NET0131 ,
		_w1264_,
		_w1411_,
		_w1712_,
		_w1714_
	);
	LUT4 #(
		.INIT('hf5c4)
	) name1252 (
		_w1447_,
		_w1496_,
		_w1713_,
		_w1714_,
		_w1715_
	);
	LUT4 #(
		.INIT('h3111)
	) name1253 (
		_w1359_,
		_w1656_,
		_w1690_,
		_w1715_,
		_w1716_
	);
	LUT3 #(
		.INIT('hce)
	) name1254 (
		\P1_state_reg[0]/NET0131 ,
		_w1655_,
		_w1716_,
		_w1717_
	);
	LUT4 #(
		.INIT('h4000)
	) name1255 (
		\P1_IR_reg[10]/NET0131 ,
		_w465_,
		_w466_,
		_w479_,
		_w1718_
	);
	LUT4 #(
		.INIT('h0001)
	) name1256 (
		\P1_IR_reg[11]/NET0131 ,
		\P1_IR_reg[12]/NET0131 ,
		\P1_IR_reg[13]/NET0131 ,
		\P1_IR_reg[14]/NET0131 ,
		_w1719_
	);
	LUT4 #(
		.INIT('h0001)
	) name1257 (
		\P1_IR_reg[15]/NET0131 ,
		\P1_IR_reg[16]/NET0131 ,
		\P1_IR_reg[17]/NET0131 ,
		\P1_IR_reg[18]/NET0131 ,
		_w1720_
	);
	LUT4 #(
		.INIT('h0001)
	) name1258 (
		\P1_IR_reg[19]/NET0131 ,
		\P1_IR_reg[20]/NET0131 ,
		\P1_IR_reg[21]/NET0131 ,
		\P1_IR_reg[22]/NET0131 ,
		_w1721_
	);
	LUT4 #(
		.INIT('h8000)
	) name1259 (
		_w1718_,
		_w1719_,
		_w1720_,
		_w1721_,
		_w1722_
	);
	LUT3 #(
		.INIT('ha6)
	) name1260 (
		\P1_IR_reg[23]/NET0131 ,
		\P1_IR_reg[31]/NET0131 ,
		_w1722_,
		_w1723_
	);
	LUT4 #(
		.INIT('h0001)
	) name1261 (
		\P1_IR_reg[16]/NET0131 ,
		\P1_IR_reg[17]/NET0131 ,
		\P1_IR_reg[18]/NET0131 ,
		\P1_IR_reg[19]/NET0131 ,
		_w1724_
	);
	LUT4 #(
		.INIT('h0001)
	) name1262 (
		\P1_IR_reg[20]/NET0131 ,
		\P1_IR_reg[21]/NET0131 ,
		\P1_IR_reg[22]/NET0131 ,
		\P1_IR_reg[23]/NET0131 ,
		_w1725_
	);
	LUT4 #(
		.INIT('h8000)
	) name1263 (
		_w468_,
		_w480_,
		_w1724_,
		_w1725_,
		_w1726_
	);
	LUT3 #(
		.INIT('ha6)
	) name1264 (
		\P1_IR_reg[24]/NET0131 ,
		\P1_IR_reg[31]/NET0131 ,
		_w1726_,
		_w1727_
	);
	LUT2 #(
		.INIT('h9)
	) name1265 (
		\P1_IR_reg[25]/NET0131 ,
		_w475_,
		_w1728_
	);
	LUT2 #(
		.INIT('h6)
	) name1266 (
		\P1_IR_reg[26]/NET0131 ,
		_w484_,
		_w1729_
	);
	LUT4 #(
		.INIT('h1248)
	) name1267 (
		\P1_IR_reg[25]/NET0131 ,
		\P1_IR_reg[26]/NET0131 ,
		_w475_,
		_w484_,
		_w1730_
	);
	LUT3 #(
		.INIT('h15)
	) name1268 (
		_w1723_,
		_w1727_,
		_w1730_,
		_w1731_
	);
	LUT4 #(
		.INIT('h2184)
	) name1269 (
		\P1_IR_reg[25]/NET0131 ,
		\P1_IR_reg[26]/NET0131 ,
		_w475_,
		_w484_,
		_w1732_
	);
	LUT4 #(
		.INIT('h4414)
	) name1270 (
		\P1_B_reg/NET0131 ,
		\P1_IR_reg[24]/NET0131 ,
		\P1_IR_reg[31]/NET0131 ,
		_w1726_,
		_w1733_
	);
	LUT2 #(
		.INIT('h8)
	) name1271 (
		_w1732_,
		_w1733_,
		_w1734_
	);
	LUT4 #(
		.INIT('he0a0)
	) name1272 (
		\P1_d_reg[0]/NET0131 ,
		_w1728_,
		_w1729_,
		_w1733_,
		_w1735_
	);
	LUT4 #(
		.INIT('h2282)
	) name1273 (
		\P1_B_reg/NET0131 ,
		\P1_IR_reg[24]/NET0131 ,
		\P1_IR_reg[31]/NET0131 ,
		_w1726_,
		_w1736_
	);
	LUT4 #(
		.INIT('hc5cf)
	) name1274 (
		\P1_B_reg/NET0131 ,
		_w1729_,
		_w1727_,
		_w1732_,
		_w1737_
	);
	LUT2 #(
		.INIT('hb)
	) name1275 (
		_w1735_,
		_w1737_,
		_w1738_
	);
	LUT4 #(
		.INIT('h1c5c)
	) name1276 (
		\P1_d_reg[1]/NET0131 ,
		_w1728_,
		_w1729_,
		_w1736_,
		_w1739_
	);
	LUT2 #(
		.INIT('hb)
	) name1277 (
		_w1734_,
		_w1739_,
		_w1740_
	);
	LUT4 #(
		.INIT('h2030)
	) name1278 (
		_w1734_,
		_w1735_,
		_w1737_,
		_w1739_,
		_w1741_
	);
	LUT4 #(
		.INIT('h0001)
	) name1279 (
		\P1_IR_reg[23]/NET0131 ,
		\P1_IR_reg[24]/NET0131 ,
		\P1_IR_reg[25]/NET0131 ,
		\P1_IR_reg[26]/NET0131 ,
		_w1742_
	);
	LUT2 #(
		.INIT('h2)
	) name1280 (
		\P1_IR_reg[31]/NET0131 ,
		_w1742_,
		_w1743_
	);
	LUT4 #(
		.INIT('h55a6)
	) name1281 (
		\P1_IR_reg[27]/NET0131 ,
		\P1_IR_reg[31]/NET0131 ,
		_w1722_,
		_w1743_,
		_w1744_
	);
	LUT4 #(
		.INIT('h0001)
	) name1282 (
		\P1_IR_reg[24]/NET0131 ,
		\P1_IR_reg[25]/NET0131 ,
		\P1_IR_reg[26]/NET0131 ,
		\P1_IR_reg[27]/NET0131 ,
		_w1745_
	);
	LUT2 #(
		.INIT('h2)
	) name1283 (
		\P1_IR_reg[31]/NET0131 ,
		_w1745_,
		_w1746_
	);
	LUT4 #(
		.INIT('h55a6)
	) name1284 (
		\P1_IR_reg[28]/NET0131 ,
		\P1_IR_reg[31]/NET0131 ,
		_w1726_,
		_w1746_,
		_w1747_
	);
	LUT2 #(
		.INIT('h1)
	) name1285 (
		_w1744_,
		_w1747_,
		_w1748_
	);
	LUT2 #(
		.INIT('h1)
	) name1286 (
		\P2_datao_reg[28]/NET0131 ,
		\si[28]_pad ,
		_w1749_
	);
	LUT4 #(
		.INIT('hfac8)
	) name1287 (
		\P2_datao_reg[18]/NET0131 ,
		\P2_datao_reg[19]/NET0131 ,
		\si[18]_pad ,
		\si[19]_pad ,
		_w1750_
	);
	LUT2 #(
		.INIT('h1)
	) name1288 (
		\P2_datao_reg[17]/NET0131 ,
		\si[17]_pad ,
		_w1751_
	);
	LUT4 #(
		.INIT('hec80)
	) name1289 (
		\P2_datao_reg[16]/NET0131 ,
		\P2_datao_reg[17]/NET0131 ,
		\si[16]_pad ,
		\si[17]_pad ,
		_w1752_
	);
	LUT4 #(
		.INIT('hec80)
	) name1290 (
		\P2_datao_reg[18]/NET0131 ,
		\P2_datao_reg[19]/NET0131 ,
		\si[18]_pad ,
		\si[19]_pad ,
		_w1753_
	);
	LUT3 #(
		.INIT('h07)
	) name1291 (
		_w1750_,
		_w1752_,
		_w1753_,
		_w1754_
	);
	LUT4 #(
		.INIT('hfac8)
	) name1292 (
		\P2_datao_reg[16]/NET0131 ,
		\P2_datao_reg[17]/NET0131 ,
		\si[16]_pad ,
		\si[17]_pad ,
		_w1755_
	);
	LUT2 #(
		.INIT('h8)
	) name1293 (
		_w1750_,
		_w1755_,
		_w1756_
	);
	LUT2 #(
		.INIT('h8)
	) name1294 (
		\P2_datao_reg[7]/NET0131 ,
		\si[7]_pad ,
		_w1757_
	);
	LUT4 #(
		.INIT('hfac8)
	) name1295 (
		\P2_datao_reg[4]/NET0131 ,
		\P2_datao_reg[5]/NET0131 ,
		\si[4]_pad ,
		\si[5]_pad ,
		_w1758_
	);
	LUT2 #(
		.INIT('h1)
	) name1296 (
		\P2_datao_reg[3]/NET0131 ,
		\si[3]_pad ,
		_w1759_
	);
	LUT2 #(
		.INIT('h1)
	) name1297 (
		\P2_datao_reg[2]/NET0131 ,
		\si[2]_pad ,
		_w1760_
	);
	LUT2 #(
		.INIT('h8)
	) name1298 (
		\P2_datao_reg[0]/NET0131 ,
		\si[0]_pad ,
		_w1761_
	);
	LUT4 #(
		.INIT('hec80)
	) name1299 (
		\P2_datao_reg[0]/NET0131 ,
		\P2_datao_reg[1]/NET0131 ,
		\si[0]_pad ,
		\si[1]_pad ,
		_w1762_
	);
	LUT4 #(
		.INIT('h135f)
	) name1300 (
		\P2_datao_reg[2]/NET0131 ,
		\P2_datao_reg[3]/NET0131 ,
		\si[2]_pad ,
		\si[3]_pad ,
		_w1763_
	);
	LUT4 #(
		.INIT('h1055)
	) name1301 (
		_w1759_,
		_w1760_,
		_w1762_,
		_w1763_,
		_w1764_
	);
	LUT2 #(
		.INIT('h8)
	) name1302 (
		\P2_datao_reg[6]/NET0131 ,
		\si[6]_pad ,
		_w1765_
	);
	LUT2 #(
		.INIT('h8)
	) name1303 (
		\P2_datao_reg[4]/NET0131 ,
		\si[4]_pad ,
		_w1766_
	);
	LUT4 #(
		.INIT('hec80)
	) name1304 (
		\P2_datao_reg[4]/NET0131 ,
		\P2_datao_reg[5]/NET0131 ,
		\si[4]_pad ,
		\si[5]_pad ,
		_w1767_
	);
	LUT2 #(
		.INIT('h1)
	) name1305 (
		_w1765_,
		_w1767_,
		_w1768_
	);
	LUT2 #(
		.INIT('h1)
	) name1306 (
		\P2_datao_reg[6]/NET0131 ,
		\si[6]_pad ,
		_w1769_
	);
	LUT4 #(
		.INIT('hfac8)
	) name1307 (
		\P2_datao_reg[6]/NET0131 ,
		\P2_datao_reg[7]/NET0131 ,
		\si[6]_pad ,
		\si[7]_pad ,
		_w1770_
	);
	LUT4 #(
		.INIT('h8f00)
	) name1308 (
		_w1758_,
		_w1764_,
		_w1768_,
		_w1770_,
		_w1771_
	);
	LUT2 #(
		.INIT('h1)
	) name1309 (
		\P2_datao_reg[9]/NET0131 ,
		\si[9]_pad ,
		_w1772_
	);
	LUT4 #(
		.INIT('hfac8)
	) name1310 (
		\P2_datao_reg[10]/NET0131 ,
		\P2_datao_reg[9]/NET0131 ,
		\si[10]_pad ,
		\si[9]_pad ,
		_w1773_
	);
	LUT2 #(
		.INIT('h1)
	) name1311 (
		\P2_datao_reg[8]/NET0131 ,
		\si[8]_pad ,
		_w1774_
	);
	LUT2 #(
		.INIT('h1)
	) name1312 (
		\P2_datao_reg[11]/NET0131 ,
		\si[11]_pad ,
		_w1775_
	);
	LUT3 #(
		.INIT('h02)
	) name1313 (
		_w1773_,
		_w1774_,
		_w1775_,
		_w1776_
	);
	LUT2 #(
		.INIT('h1)
	) name1314 (
		\P2_datao_reg[14]/NET0131 ,
		\si[14]_pad ,
		_w1777_
	);
	LUT4 #(
		.INIT('hfac8)
	) name1315 (
		\P2_datao_reg[14]/NET0131 ,
		\P2_datao_reg[15]/NET0131 ,
		\si[14]_pad ,
		\si[15]_pad ,
		_w1778_
	);
	LUT2 #(
		.INIT('h1)
	) name1316 (
		\P2_datao_reg[13]/NET0131 ,
		\si[13]_pad ,
		_w1779_
	);
	LUT4 #(
		.INIT('hfac8)
	) name1317 (
		\P2_datao_reg[12]/NET0131 ,
		\P2_datao_reg[13]/NET0131 ,
		\si[12]_pad ,
		\si[13]_pad ,
		_w1780_
	);
	LUT2 #(
		.INIT('h8)
	) name1318 (
		_w1778_,
		_w1780_,
		_w1781_
	);
	LUT4 #(
		.INIT('he000)
	) name1319 (
		_w1757_,
		_w1771_,
		_w1776_,
		_w1781_,
		_w1782_
	);
	LUT2 #(
		.INIT('h8)
	) name1320 (
		\P2_datao_reg[11]/NET0131 ,
		\si[11]_pad ,
		_w1783_
	);
	LUT2 #(
		.INIT('h8)
	) name1321 (
		\P2_datao_reg[10]/NET0131 ,
		\si[10]_pad ,
		_w1784_
	);
	LUT2 #(
		.INIT('h8)
	) name1322 (
		\P2_datao_reg[8]/NET0131 ,
		\si[8]_pad ,
		_w1785_
	);
	LUT4 #(
		.INIT('hec80)
	) name1323 (
		\P2_datao_reg[8]/NET0131 ,
		\P2_datao_reg[9]/NET0131 ,
		\si[8]_pad ,
		\si[9]_pad ,
		_w1786_
	);
	LUT4 #(
		.INIT('hfac8)
	) name1324 (
		\P2_datao_reg[10]/NET0131 ,
		\P2_datao_reg[11]/NET0131 ,
		\si[10]_pad ,
		\si[11]_pad ,
		_w1787_
	);
	LUT4 #(
		.INIT('h0155)
	) name1325 (
		_w1783_,
		_w1784_,
		_w1786_,
		_w1787_,
		_w1788_
	);
	LUT2 #(
		.INIT('h8)
	) name1326 (
		\P2_datao_reg[12]/NET0131 ,
		\si[12]_pad ,
		_w1789_
	);
	LUT4 #(
		.INIT('hec80)
	) name1327 (
		\P2_datao_reg[12]/NET0131 ,
		\P2_datao_reg[13]/NET0131 ,
		\si[12]_pad ,
		\si[13]_pad ,
		_w1790_
	);
	LUT4 #(
		.INIT('hec80)
	) name1328 (
		\P2_datao_reg[14]/NET0131 ,
		\P2_datao_reg[15]/NET0131 ,
		\si[14]_pad ,
		\si[15]_pad ,
		_w1791_
	);
	LUT3 #(
		.INIT('h07)
	) name1329 (
		_w1778_,
		_w1790_,
		_w1791_,
		_w1792_
	);
	LUT3 #(
		.INIT('hd0)
	) name1330 (
		_w1781_,
		_w1788_,
		_w1792_,
		_w1793_
	);
	LUT4 #(
		.INIT('h2a22)
	) name1331 (
		_w1754_,
		_w1756_,
		_w1782_,
		_w1793_,
		_w1794_
	);
	LUT2 #(
		.INIT('h1)
	) name1332 (
		\P2_datao_reg[20]/NET0131 ,
		\si[20]_pad ,
		_w1795_
	);
	LUT2 #(
		.INIT('h1)
	) name1333 (
		\P2_datao_reg[26]/NET0131 ,
		\si[26]_pad ,
		_w1796_
	);
	LUT2 #(
		.INIT('h1)
	) name1334 (
		\P2_datao_reg[24]/NET0131 ,
		\si[24]_pad ,
		_w1797_
	);
	LUT4 #(
		.INIT('hfac8)
	) name1335 (
		\P2_datao_reg[24]/NET0131 ,
		\P2_datao_reg[25]/NET0131 ,
		\si[24]_pad ,
		\si[25]_pad ,
		_w1798_
	);
	LUT2 #(
		.INIT('h4)
	) name1336 (
		_w1796_,
		_w1798_,
		_w1799_
	);
	LUT2 #(
		.INIT('h1)
	) name1337 (
		\P2_datao_reg[23]/NET0131 ,
		\si[23]_pad ,
		_w1800_
	);
	LUT2 #(
		.INIT('h1)
	) name1338 (
		\P2_datao_reg[21]/NET0131 ,
		\si[21]_pad ,
		_w1801_
	);
	LUT4 #(
		.INIT('hfac8)
	) name1339 (
		\P2_datao_reg[21]/NET0131 ,
		\P2_datao_reg[22]/NET0131 ,
		\si[21]_pad ,
		\si[22]_pad ,
		_w1802_
	);
	LUT2 #(
		.INIT('h1)
	) name1340 (
		\P2_datao_reg[27]/NET0131 ,
		\si[27]_pad ,
		_w1803_
	);
	LUT3 #(
		.INIT('h04)
	) name1341 (
		_w1800_,
		_w1802_,
		_w1803_,
		_w1804_
	);
	LUT2 #(
		.INIT('h8)
	) name1342 (
		_w1799_,
		_w1804_,
		_w1805_
	);
	LUT3 #(
		.INIT('h40)
	) name1343 (
		_w1795_,
		_w1799_,
		_w1804_,
		_w1806_
	);
	LUT4 #(
		.INIT('hec80)
	) name1344 (
		\P2_datao_reg[22]/NET0131 ,
		\P2_datao_reg[23]/NET0131 ,
		\si[22]_pad ,
		\si[23]_pad ,
		_w1807_
	);
	LUT4 #(
		.INIT('h135f)
	) name1345 (
		\P2_datao_reg[20]/NET0131 ,
		\P2_datao_reg[21]/NET0131 ,
		\si[20]_pad ,
		\si[21]_pad ,
		_w1808_
	);
	LUT4 #(
		.INIT('h0f0b)
	) name1346 (
		_w1800_,
		_w1802_,
		_w1807_,
		_w1808_,
		_w1809_
	);
	LUT4 #(
		.INIT('h135f)
	) name1347 (
		\P2_datao_reg[26]/NET0131 ,
		\P2_datao_reg[27]/NET0131 ,
		\si[26]_pad ,
		\si[27]_pad ,
		_w1810_
	);
	LUT4 #(
		.INIT('hec80)
	) name1348 (
		\P2_datao_reg[24]/NET0131 ,
		\P2_datao_reg[25]/NET0131 ,
		\si[24]_pad ,
		\si[25]_pad ,
		_w1811_
	);
	LUT3 #(
		.INIT('h8c)
	) name1349 (
		_w1796_,
		_w1810_,
		_w1811_,
		_w1812_
	);
	LUT4 #(
		.INIT('h0233)
	) name1350 (
		_w1799_,
		_w1803_,
		_w1809_,
		_w1812_,
		_w1813_
	);
	LUT3 #(
		.INIT('h0b)
	) name1351 (
		_w1794_,
		_w1806_,
		_w1813_,
		_w1814_
	);
	LUT4 #(
		.INIT('h5956)
	) name1352 (
		\P2_datao_reg[28]/NET0131 ,
		\si[28]_pad ,
		_w547_,
		_w1814_,
		_w1815_
	);
	LUT2 #(
		.INIT('h1)
	) name1353 (
		_w1748_,
		_w1815_,
		_w1816_
	);
	LUT4 #(
		.INIT('h8000)
	) name1354 (
		\P1_reg3_reg[3]/NET0131 ,
		\P1_reg3_reg[4]/NET0131 ,
		\P1_reg3_reg[5]/NET0131 ,
		\P1_reg3_reg[6]/NET0131 ,
		_w1817_
	);
	LUT4 #(
		.INIT('h8000)
	) name1355 (
		\P1_reg3_reg[10]/NET0131 ,
		\P1_reg3_reg[7]/NET0131 ,
		\P1_reg3_reg[8]/NET0131 ,
		\P1_reg3_reg[9]/NET0131 ,
		_w1818_
	);
	LUT2 #(
		.INIT('h8)
	) name1356 (
		_w1817_,
		_w1818_,
		_w1819_
	);
	LUT2 #(
		.INIT('h8)
	) name1357 (
		\P1_reg3_reg[11]/NET0131 ,
		\P1_reg3_reg[12]/NET0131 ,
		_w1820_
	);
	LUT4 #(
		.INIT('h8000)
	) name1358 (
		\P1_reg3_reg[13]/NET0131 ,
		_w1817_,
		_w1818_,
		_w1820_,
		_w1821_
	);
	LUT2 #(
		.INIT('h8)
	) name1359 (
		\P1_reg3_reg[16]/NET0131 ,
		\P1_reg3_reg[17]/NET0131 ,
		_w1822_
	);
	LUT4 #(
		.INIT('h8000)
	) name1360 (
		\P1_reg3_reg[15]/NET0131 ,
		\P1_reg3_reg[18]/NET0131 ,
		\P1_reg3_reg[19]/NET0131 ,
		\P1_reg3_reg[20]/NET0131 ,
		_w1823_
	);
	LUT2 #(
		.INIT('h8)
	) name1361 (
		_w1822_,
		_w1823_,
		_w1824_
	);
	LUT3 #(
		.INIT('h80)
	) name1362 (
		\P1_reg3_reg[14]/NET0131 ,
		_w1821_,
		_w1824_,
		_w1825_
	);
	LUT2 #(
		.INIT('h8)
	) name1363 (
		\P1_reg3_reg[21]/NET0131 ,
		\P1_reg3_reg[22]/NET0131 ,
		_w1826_
	);
	LUT4 #(
		.INIT('h8000)
	) name1364 (
		\P1_reg3_reg[14]/NET0131 ,
		_w1821_,
		_w1824_,
		_w1826_,
		_w1827_
	);
	LUT3 #(
		.INIT('h80)
	) name1365 (
		\P1_reg3_reg[23]/NET0131 ,
		\P1_reg3_reg[24]/NET0131 ,
		_w1827_,
		_w1828_
	);
	LUT2 #(
		.INIT('h8)
	) name1366 (
		\P1_reg3_reg[25]/NET0131 ,
		\P1_reg3_reg[26]/NET0131 ,
		_w1829_
	);
	LUT4 #(
		.INIT('h8000)
	) name1367 (
		\P1_reg3_reg[23]/NET0131 ,
		\P1_reg3_reg[24]/NET0131 ,
		_w1827_,
		_w1829_,
		_w1830_
	);
	LUT4 #(
		.INIT('h8000)
	) name1368 (
		\P1_reg3_reg[25]/NET0131 ,
		\P1_reg3_reg[26]/NET0131 ,
		\P1_reg3_reg[27]/NET0131 ,
		\P1_reg3_reg[28]/NET0131 ,
		_w1831_
	);
	LUT4 #(
		.INIT('h8000)
	) name1369 (
		\P1_reg3_reg[23]/NET0131 ,
		\P1_reg3_reg[24]/NET0131 ,
		_w1827_,
		_w1831_,
		_w1832_
	);
	LUT4 #(
		.INIT('h6ccc)
	) name1370 (
		\P1_reg3_reg[27]/NET0131 ,
		\P1_reg3_reg[28]/NET0131 ,
		_w1828_,
		_w1829_,
		_w1833_
	);
	LUT3 #(
		.INIT('h02)
	) name1371 (
		\P1_reg0_reg[28]/NET0131 ,
		_w478_,
		_w488_,
		_w1834_
	);
	LUT4 #(
		.INIT('hf35f)
	) name1372 (
		\P1_reg1_reg[28]/NET0131 ,
		\P1_reg2_reg[28]/NET0131 ,
		_w478_,
		_w488_,
		_w1835_
	);
	LUT4 #(
		.INIT('h1300)
	) name1373 (
		_w490_,
		_w1834_,
		_w1833_,
		_w1835_,
		_w1836_
	);
	LUT4 #(
		.INIT('hecff)
	) name1374 (
		_w490_,
		_w1834_,
		_w1833_,
		_w1835_,
		_w1837_
	);
	LUT3 #(
		.INIT('he0)
	) name1375 (
		_w1748_,
		_w1815_,
		_w1836_,
		_w1838_
	);
	LUT2 #(
		.INIT('h8)
	) name1376 (
		\P2_datao_reg[25]/NET0131 ,
		_w547_,
		_w1839_
	);
	LUT2 #(
		.INIT('h6)
	) name1377 (
		\P2_datao_reg[25]/NET0131 ,
		\si[25]_pad ,
		_w1840_
	);
	LUT4 #(
		.INIT('hec80)
	) name1378 (
		\P2_datao_reg[17]/NET0131 ,
		\P2_datao_reg[18]/NET0131 ,
		\si[17]_pad ,
		\si[18]_pad ,
		_w1841_
	);
	LUT4 #(
		.INIT('hfac8)
	) name1379 (
		\P2_datao_reg[19]/NET0131 ,
		\P2_datao_reg[20]/NET0131 ,
		\si[19]_pad ,
		\si[20]_pad ,
		_w1842_
	);
	LUT4 #(
		.INIT('hec80)
	) name1380 (
		\P2_datao_reg[19]/NET0131 ,
		\P2_datao_reg[20]/NET0131 ,
		\si[19]_pad ,
		\si[20]_pad ,
		_w1843_
	);
	LUT3 #(
		.INIT('h07)
	) name1381 (
		_w1841_,
		_w1842_,
		_w1843_,
		_w1844_
	);
	LUT4 #(
		.INIT('hfac8)
	) name1382 (
		\P2_datao_reg[17]/NET0131 ,
		\P2_datao_reg[18]/NET0131 ,
		\si[17]_pad ,
		\si[18]_pad ,
		_w1845_
	);
	LUT2 #(
		.INIT('h8)
	) name1383 (
		_w1842_,
		_w1845_,
		_w1846_
	);
	LUT2 #(
		.INIT('h2)
	) name1384 (
		_w1758_,
		_w1769_,
		_w1847_
	);
	LUT4 #(
		.INIT('hfac8)
	) name1385 (
		\P2_datao_reg[7]/NET0131 ,
		\P2_datao_reg[8]/NET0131 ,
		\si[7]_pad ,
		\si[8]_pad ,
		_w1848_
	);
	LUT3 #(
		.INIT('h20)
	) name1386 (
		_w1758_,
		_w1769_,
		_w1848_,
		_w1849_
	);
	LUT4 #(
		.INIT('hec80)
	) name1387 (
		\P2_datao_reg[5]/NET0131 ,
		\P2_datao_reg[6]/NET0131 ,
		\si[5]_pad ,
		\si[6]_pad ,
		_w1850_
	);
	LUT4 #(
		.INIT('h0313)
	) name1388 (
		_w1757_,
		_w1785_,
		_w1848_,
		_w1850_,
		_w1851_
	);
	LUT4 #(
		.INIT('h1f00)
	) name1389 (
		_w1764_,
		_w1766_,
		_w1849_,
		_w1851_,
		_w1852_
	);
	LUT4 #(
		.INIT('hfac8)
	) name1390 (
		\P2_datao_reg[11]/NET0131 ,
		\P2_datao_reg[12]/NET0131 ,
		\si[11]_pad ,
		\si[12]_pad ,
		_w1853_
	);
	LUT2 #(
		.INIT('h8)
	) name1391 (
		_w1773_,
		_w1853_,
		_w1854_
	);
	LUT4 #(
		.INIT('hfac8)
	) name1392 (
		\P2_datao_reg[15]/NET0131 ,
		\P2_datao_reg[16]/NET0131 ,
		\si[15]_pad ,
		\si[16]_pad ,
		_w1855_
	);
	LUT3 #(
		.INIT('h10)
	) name1393 (
		_w1777_,
		_w1779_,
		_w1855_,
		_w1856_
	);
	LUT4 #(
		.INIT('hec80)
	) name1394 (
		\P2_datao_reg[15]/NET0131 ,
		\P2_datao_reg[16]/NET0131 ,
		\si[15]_pad ,
		\si[16]_pad ,
		_w1857_
	);
	LUT4 #(
		.INIT('h135f)
	) name1395 (
		\P2_datao_reg[13]/NET0131 ,
		\P2_datao_reg[14]/NET0131 ,
		\si[13]_pad ,
		\si[14]_pad ,
		_w1858_
	);
	LUT4 #(
		.INIT('h0f0b)
	) name1396 (
		_w1777_,
		_w1855_,
		_w1857_,
		_w1858_,
		_w1859_
	);
	LUT4 #(
		.INIT('he8a0)
	) name1397 (
		\P2_datao_reg[10]/NET0131 ,
		\P2_datao_reg[9]/NET0131 ,
		\si[10]_pad ,
		\si[9]_pad ,
		_w1860_
	);
	LUT4 #(
		.INIT('h0515)
	) name1398 (
		_w1789_,
		_w1783_,
		_w1853_,
		_w1860_,
		_w1861_
	);
	LUT3 #(
		.INIT('hc4)
	) name1399 (
		_w1856_,
		_w1859_,
		_w1861_,
		_w1862_
	);
	LUT4 #(
		.INIT('hbf00)
	) name1400 (
		_w1852_,
		_w1854_,
		_w1856_,
		_w1862_,
		_w1863_
	);
	LUT3 #(
		.INIT('h04)
	) name1401 (
		_w1800_,
		_w1802_,
		_w1797_,
		_w1864_
	);
	LUT4 #(
		.INIT('h5d00)
	) name1402 (
		_w1844_,
		_w1846_,
		_w1863_,
		_w1864_,
		_w1865_
	);
	LUT4 #(
		.INIT('h135f)
	) name1403 (
		\P2_datao_reg[23]/NET0131 ,
		\P2_datao_reg[24]/NET0131 ,
		\si[23]_pad ,
		\si[24]_pad ,
		_w1866_
	);
	LUT4 #(
		.INIT('hec80)
	) name1404 (
		\P2_datao_reg[21]/NET0131 ,
		\P2_datao_reg[22]/NET0131 ,
		\si[21]_pad ,
		\si[22]_pad ,
		_w1867_
	);
	LUT3 #(
		.INIT('h8c)
	) name1405 (
		_w1800_,
		_w1866_,
		_w1867_,
		_w1868_
	);
	LUT4 #(
		.INIT('h1303)
	) name1406 (
		_w1800_,
		_w1797_,
		_w1866_,
		_w1867_,
		_w1869_
	);
	LUT4 #(
		.INIT('h1114)
	) name1407 (
		_w547_,
		_w1840_,
		_w1865_,
		_w1869_,
		_w1870_
	);
	LUT3 #(
		.INIT('h54)
	) name1408 (
		_w1748_,
		_w1839_,
		_w1870_,
		_w1871_
	);
	LUT4 #(
		.INIT('h78f0)
	) name1409 (
		\P1_reg3_reg[23]/NET0131 ,
		\P1_reg3_reg[24]/NET0131 ,
		\P1_reg3_reg[25]/NET0131 ,
		_w1827_,
		_w1872_
	);
	LUT3 #(
		.INIT('h80)
	) name1410 (
		_w478_,
		_w488_,
		_w1872_,
		_w1873_
	);
	LUT3 #(
		.INIT('h20)
	) name1411 (
		\P1_reg2_reg[25]/NET0131 ,
		_w478_,
		_w488_,
		_w1874_
	);
	LUT4 #(
		.INIT('hff35)
	) name1412 (
		\P1_reg0_reg[25]/NET0131 ,
		\P1_reg1_reg[25]/NET0131 ,
		_w478_,
		_w488_,
		_w1875_
	);
	LUT3 #(
		.INIT('h10)
	) name1413 (
		_w1874_,
		_w1873_,
		_w1875_,
		_w1876_
	);
	LUT3 #(
		.INIT('hef)
	) name1414 (
		_w1874_,
		_w1873_,
		_w1875_,
		_w1877_
	);
	LUT4 #(
		.INIT('hab00)
	) name1415 (
		_w1748_,
		_w1839_,
		_w1870_,
		_w1876_,
		_w1878_
	);
	LUT3 #(
		.INIT('h07)
	) name1416 (
		_w1758_,
		_w1764_,
		_w1767_,
		_w1879_
	);
	LUT3 #(
		.INIT('h10)
	) name1417 (
		_w1769_,
		_w1772_,
		_w1848_,
		_w1880_
	);
	LUT4 #(
		.INIT('hf800)
	) name1418 (
		_w1758_,
		_w1764_,
		_w1767_,
		_w1880_,
		_w1881_
	);
	LUT4 #(
		.INIT('h135f)
	) name1419 (
		\P2_datao_reg[6]/NET0131 ,
		\P2_datao_reg[7]/NET0131 ,
		\si[6]_pad ,
		\si[7]_pad ,
		_w1882_
	);
	LUT4 #(
		.INIT('h3323)
	) name1420 (
		_w1772_,
		_w1786_,
		_w1848_,
		_w1882_,
		_w1883_
	);
	LUT2 #(
		.INIT('h8)
	) name1421 (
		_w1780_,
		_w1787_,
		_w1884_
	);
	LUT3 #(
		.INIT('h10)
	) name1422 (
		_w1751_,
		_w1777_,
		_w1855_,
		_w1885_
	);
	LUT4 #(
		.INIT('hb000)
	) name1423 (
		_w1881_,
		_w1883_,
		_w1884_,
		_w1885_,
		_w1886_
	);
	LUT4 #(
		.INIT('h135f)
	) name1424 (
		\P2_datao_reg[10]/NET0131 ,
		\P2_datao_reg[11]/NET0131 ,
		\si[10]_pad ,
		\si[11]_pad ,
		_w1887_
	);
	LUT4 #(
		.INIT('h3323)
	) name1425 (
		_w1779_,
		_w1790_,
		_w1853_,
		_w1887_,
		_w1888_
	);
	LUT3 #(
		.INIT('h15)
	) name1426 (
		_w1752_,
		_w1755_,
		_w1791_,
		_w1889_
	);
	LUT3 #(
		.INIT('hd0)
	) name1427 (
		_w1885_,
		_w1888_,
		_w1889_,
		_w1890_
	);
	LUT4 #(
		.INIT('hfac8)
	) name1428 (
		\P2_datao_reg[20]/NET0131 ,
		\P2_datao_reg[21]/NET0131 ,
		\si[20]_pad ,
		\si[21]_pad ,
		_w1891_
	);
	LUT2 #(
		.INIT('h8)
	) name1429 (
		_w1750_,
		_w1891_,
		_w1892_
	);
	LUT4 #(
		.INIT('h020f)
	) name1430 (
		_w1753_,
		_w1795_,
		_w1801_,
		_w1808_,
		_w1893_
	);
	LUT4 #(
		.INIT('h004f)
	) name1431 (
		_w1886_,
		_w1890_,
		_w1892_,
		_w1893_,
		_w1894_
	);
	LUT4 #(
		.INIT('hfac8)
	) name1432 (
		\P2_datao_reg[22]/NET0131 ,
		\P2_datao_reg[23]/NET0131 ,
		\si[22]_pad ,
		\si[23]_pad ,
		_w1895_
	);
	LUT2 #(
		.INIT('h8)
	) name1433 (
		_w1798_,
		_w1895_,
		_w1896_
	);
	LUT3 #(
		.INIT('h07)
	) name1434 (
		_w1798_,
		_w1807_,
		_w1811_,
		_w1897_
	);
	LUT3 #(
		.INIT('hb0)
	) name1435 (
		_w1894_,
		_w1896_,
		_w1897_,
		_w1898_
	);
	LUT4 #(
		.INIT('h5956)
	) name1436 (
		\P2_datao_reg[26]/NET0131 ,
		\si[26]_pad ,
		_w547_,
		_w1898_,
		_w1899_
	);
	LUT2 #(
		.INIT('h1)
	) name1437 (
		_w1748_,
		_w1899_,
		_w1900_
	);
	LUT3 #(
		.INIT('h6c)
	) name1438 (
		\P1_reg3_reg[25]/NET0131 ,
		\P1_reg3_reg[26]/NET0131 ,
		_w1828_,
		_w1901_
	);
	LUT3 #(
		.INIT('h02)
	) name1439 (
		\P1_reg0_reg[26]/NET0131 ,
		_w478_,
		_w488_,
		_w1902_
	);
	LUT4 #(
		.INIT('hf35f)
	) name1440 (
		\P1_reg1_reg[26]/NET0131 ,
		\P1_reg2_reg[26]/NET0131 ,
		_w478_,
		_w488_,
		_w1903_
	);
	LUT4 #(
		.INIT('h1300)
	) name1441 (
		_w490_,
		_w1902_,
		_w1901_,
		_w1903_,
		_w1904_
	);
	LUT4 #(
		.INIT('hecff)
	) name1442 (
		_w490_,
		_w1902_,
		_w1901_,
		_w1903_,
		_w1905_
	);
	LUT3 #(
		.INIT('he0)
	) name1443 (
		_w1748_,
		_w1899_,
		_w1904_,
		_w1906_
	);
	LUT2 #(
		.INIT('h8)
	) name1444 (
		\P2_datao_reg[27]/NET0131 ,
		_w547_,
		_w1907_
	);
	LUT2 #(
		.INIT('h6)
	) name1445 (
		\P2_datao_reg[27]/NET0131 ,
		\si[27]_pad ,
		_w1908_
	);
	LUT4 #(
		.INIT('hec80)
	) name1446 (
		\P2_datao_reg[25]/NET0131 ,
		\P2_datao_reg[26]/NET0131 ,
		\si[25]_pad ,
		\si[26]_pad ,
		_w1909_
	);
	LUT4 #(
		.INIT('h00fb)
	) name1447 (
		_w1796_,
		_w1798_,
		_w1866_,
		_w1909_,
		_w1910_
	);
	LUT3 #(
		.INIT('h10)
	) name1448 (
		_w1800_,
		_w1796_,
		_w1798_,
		_w1911_
	);
	LUT4 #(
		.INIT('h001f)
	) name1449 (
		_w1764_,
		_w1766_,
		_w1847_,
		_w1850_,
		_w1912_
	);
	LUT2 #(
		.INIT('h8)
	) name1450 (
		_w1773_,
		_w1848_,
		_w1913_
	);
	LUT4 #(
		.INIT('h135f)
	) name1451 (
		\P2_datao_reg[7]/NET0131 ,
		\P2_datao_reg[8]/NET0131 ,
		\si[7]_pad ,
		\si[8]_pad ,
		_w1914_
	);
	LUT4 #(
		.INIT('h0f0d)
	) name1452 (
		_w1773_,
		_w1774_,
		_w1860_,
		_w1914_,
		_w1915_
	);
	LUT3 #(
		.INIT('hb0)
	) name1453 (
		_w1912_,
		_w1913_,
		_w1915_,
		_w1916_
	);
	LUT3 #(
		.INIT('h10)
	) name1454 (
		_w1777_,
		_w1779_,
		_w1853_,
		_w1917_
	);
	LUT4 #(
		.INIT('h4f00)
	) name1455 (
		_w1912_,
		_w1913_,
		_w1915_,
		_w1917_,
		_w1918_
	);
	LUT2 #(
		.INIT('h8)
	) name1456 (
		_w1802_,
		_w1842_,
		_w1919_
	);
	LUT2 #(
		.INIT('h8)
	) name1457 (
		_w1845_,
		_w1855_,
		_w1920_
	);
	LUT4 #(
		.INIT('h8000)
	) name1458 (
		_w1802_,
		_w1842_,
		_w1845_,
		_w1855_,
		_w1921_
	);
	LUT3 #(
		.INIT('h07)
	) name1459 (
		_w1802_,
		_w1843_,
		_w1867_,
		_w1922_
	);
	LUT4 #(
		.INIT('h135f)
	) name1460 (
		\P2_datao_reg[11]/NET0131 ,
		\P2_datao_reg[12]/NET0131 ,
		\si[11]_pad ,
		\si[12]_pad ,
		_w1923_
	);
	LUT4 #(
		.INIT('h0545)
	) name1461 (
		_w1777_,
		_w1780_,
		_w1858_,
		_w1923_,
		_w1924_
	);
	LUT3 #(
		.INIT('h15)
	) name1462 (
		_w1841_,
		_w1845_,
		_w1857_,
		_w1925_
	);
	LUT4 #(
		.INIT('h80aa)
	) name1463 (
		_w1919_,
		_w1920_,
		_w1924_,
		_w1925_,
		_w1926_
	);
	LUT2 #(
		.INIT('h2)
	) name1464 (
		_w1922_,
		_w1926_,
		_w1927_
	);
	LUT4 #(
		.INIT('h80aa)
	) name1465 (
		_w1911_,
		_w1918_,
		_w1921_,
		_w1927_,
		_w1928_
	);
	LUT4 #(
		.INIT('h1141)
	) name1466 (
		_w547_,
		_w1908_,
		_w1910_,
		_w1928_,
		_w1929_
	);
	LUT2 #(
		.INIT('h1)
	) name1467 (
		_w1907_,
		_w1929_,
		_w1930_
	);
	LUT3 #(
		.INIT('h54)
	) name1468 (
		_w1748_,
		_w1907_,
		_w1929_,
		_w1931_
	);
	LUT2 #(
		.INIT('h6)
	) name1469 (
		\P1_reg3_reg[27]/NET0131 ,
		_w1830_,
		_w1932_
	);
	LUT4 #(
		.INIT('h4080)
	) name1470 (
		\P1_reg3_reg[27]/NET0131 ,
		_w478_,
		_w488_,
		_w1830_,
		_w1933_
	);
	LUT3 #(
		.INIT('h08)
	) name1471 (
		\P1_reg1_reg[27]/NET0131 ,
		_w478_,
		_w488_,
		_w1934_
	);
	LUT4 #(
		.INIT('hf3f5)
	) name1472 (
		\P1_reg0_reg[27]/NET0131 ,
		\P1_reg2_reg[27]/NET0131 ,
		_w478_,
		_w488_,
		_w1935_
	);
	LUT3 #(
		.INIT('h10)
	) name1473 (
		_w1934_,
		_w1933_,
		_w1935_,
		_w1936_
	);
	LUT3 #(
		.INIT('hef)
	) name1474 (
		_w1934_,
		_w1933_,
		_w1935_,
		_w1937_
	);
	LUT4 #(
		.INIT('hab00)
	) name1475 (
		_w1748_,
		_w1907_,
		_w1929_,
		_w1936_,
		_w1938_
	);
	LUT4 #(
		.INIT('h001f)
	) name1476 (
		_w1748_,
		_w1899_,
		_w1904_,
		_w1938_,
		_w1939_
	);
	LUT2 #(
		.INIT('h4)
	) name1477 (
		_w1878_,
		_w1939_,
		_w1940_
	);
	LUT2 #(
		.INIT('h8)
	) name1478 (
		\P2_datao_reg[24]/NET0131 ,
		_w547_,
		_w1941_
	);
	LUT2 #(
		.INIT('h6)
	) name1479 (
		\P2_datao_reg[24]/NET0131 ,
		\si[24]_pad ,
		_w1942_
	);
	LUT4 #(
		.INIT('h08aa)
	) name1480 (
		_w1756_,
		_w1781_,
		_w1788_,
		_w1792_,
		_w1943_
	);
	LUT2 #(
		.INIT('h2)
	) name1481 (
		_w1754_,
		_w1943_,
		_w1944_
	);
	LUT3 #(
		.INIT('h10)
	) name1482 (
		_w1795_,
		_w1800_,
		_w1802_,
		_w1945_
	);
	LUT4 #(
		.INIT('h8f00)
	) name1483 (
		_w1756_,
		_w1782_,
		_w1944_,
		_w1945_,
		_w1946_
	);
	LUT4 #(
		.INIT('h0541)
	) name1484 (
		_w547_,
		_w1809_,
		_w1942_,
		_w1946_,
		_w1947_
	);
	LUT3 #(
		.INIT('h54)
	) name1485 (
		_w1748_,
		_w1941_,
		_w1947_,
		_w1948_
	);
	LUT4 #(
		.INIT('hff35)
	) name1486 (
		\P1_reg0_reg[24]/NET0131 ,
		\P1_reg1_reg[24]/NET0131 ,
		_w478_,
		_w488_,
		_w1949_
	);
	LUT3 #(
		.INIT('h6c)
	) name1487 (
		\P1_reg3_reg[23]/NET0131 ,
		\P1_reg3_reg[24]/NET0131 ,
		_w1827_,
		_w1950_
	);
	LUT4 #(
		.INIT('h1fdf)
	) name1488 (
		\P1_reg2_reg[24]/NET0131 ,
		_w478_,
		_w488_,
		_w1950_,
		_w1951_
	);
	LUT2 #(
		.INIT('h8)
	) name1489 (
		_w1949_,
		_w1951_,
		_w1952_
	);
	LUT2 #(
		.INIT('h7)
	) name1490 (
		_w1949_,
		_w1951_,
		_w1953_
	);
	LUT4 #(
		.INIT('hab00)
	) name1491 (
		_w1748_,
		_w1941_,
		_w1947_,
		_w1952_,
		_w1954_
	);
	LUT3 #(
		.INIT('ha2)
	) name1492 (
		_w1922_,
		_w1919_,
		_w1925_,
		_w1955_
	);
	LUT4 #(
		.INIT('h3700)
	) name1493 (
		_w1918_,
		_w1921_,
		_w1924_,
		_w1955_,
		_w1956_
	);
	LUT4 #(
		.INIT('h5956)
	) name1494 (
		\P2_datao_reg[23]/NET0131 ,
		\si[23]_pad ,
		_w547_,
		_w1956_,
		_w1957_
	);
	LUT2 #(
		.INIT('h1)
	) name1495 (
		_w1748_,
		_w1957_,
		_w1958_
	);
	LUT2 #(
		.INIT('h6)
	) name1496 (
		\P1_reg3_reg[23]/NET0131 ,
		_w1827_,
		_w1959_
	);
	LUT4 #(
		.INIT('h37f7)
	) name1497 (
		\P1_reg1_reg[23]/NET0131 ,
		_w478_,
		_w488_,
		_w1959_,
		_w1960_
	);
	LUT4 #(
		.INIT('hf3f5)
	) name1498 (
		\P1_reg0_reg[23]/NET0131 ,
		\P1_reg2_reg[23]/NET0131 ,
		_w478_,
		_w488_,
		_w1961_
	);
	LUT2 #(
		.INIT('h8)
	) name1499 (
		_w1960_,
		_w1961_,
		_w1962_
	);
	LUT2 #(
		.INIT('h7)
	) name1500 (
		_w1960_,
		_w1961_,
		_w1963_
	);
	LUT3 #(
		.INIT('he0)
	) name1501 (
		_w1748_,
		_w1957_,
		_w1962_,
		_w1964_
	);
	LUT2 #(
		.INIT('h1)
	) name1502 (
		_w1954_,
		_w1964_,
		_w1965_
	);
	LUT2 #(
		.INIT('h8)
	) name1503 (
		\P2_datao_reg[22]/NET0131 ,
		_w547_,
		_w1966_
	);
	LUT2 #(
		.INIT('h6)
	) name1504 (
		\P2_datao_reg[22]/NET0131 ,
		\si[22]_pad ,
		_w1967_
	);
	LUT4 #(
		.INIT('h4f00)
	) name1505 (
		_w1881_,
		_w1883_,
		_w1884_,
		_w1888_,
		_w1968_
	);
	LUT4 #(
		.INIT('h30b0)
	) name1506 (
		_w1885_,
		_w1889_,
		_w1892_,
		_w1968_,
		_w1969_
	);
	LUT4 #(
		.INIT('h0514)
	) name1507 (
		_w547_,
		_w1893_,
		_w1967_,
		_w1969_,
		_w1970_
	);
	LUT3 #(
		.INIT('h54)
	) name1508 (
		_w1748_,
		_w1966_,
		_w1970_,
		_w1971_
	);
	LUT4 #(
		.INIT('hff35)
	) name1509 (
		\P1_reg0_reg[22]/NET0131 ,
		\P1_reg1_reg[22]/NET0131 ,
		_w478_,
		_w488_,
		_w1972_
	);
	LUT3 #(
		.INIT('h6c)
	) name1510 (
		\P1_reg3_reg[21]/NET0131 ,
		\P1_reg3_reg[22]/NET0131 ,
		_w1825_,
		_w1973_
	);
	LUT4 #(
		.INIT('h1fdf)
	) name1511 (
		\P1_reg2_reg[22]/NET0131 ,
		_w478_,
		_w488_,
		_w1973_,
		_w1974_
	);
	LUT2 #(
		.INIT('h8)
	) name1512 (
		_w1972_,
		_w1974_,
		_w1975_
	);
	LUT2 #(
		.INIT('h7)
	) name1513 (
		_w1972_,
		_w1974_,
		_w1976_
	);
	LUT4 #(
		.INIT('h0054)
	) name1514 (
		_w1748_,
		_w1966_,
		_w1970_,
		_w1975_,
		_w1977_
	);
	LUT4 #(
		.INIT('hab00)
	) name1515 (
		_w1748_,
		_w1966_,
		_w1970_,
		_w1975_,
		_w1978_
	);
	LUT3 #(
		.INIT('hb0)
	) name1516 (
		_w1852_,
		_w1854_,
		_w1861_,
		_w1979_
	);
	LUT4 #(
		.INIT('h40f0)
	) name1517 (
		_w1852_,
		_w1854_,
		_w1856_,
		_w1861_,
		_w1980_
	);
	LUT4 #(
		.INIT('h22a2)
	) name1518 (
		_w1844_,
		_w1846_,
		_w1859_,
		_w1980_,
		_w1981_
	);
	LUT4 #(
		.INIT('h5956)
	) name1519 (
		\P2_datao_reg[21]/NET0131 ,
		\si[21]_pad ,
		_w547_,
		_w1981_,
		_w1982_
	);
	LUT2 #(
		.INIT('h1)
	) name1520 (
		_w1748_,
		_w1982_,
		_w1983_
	);
	LUT4 #(
		.INIT('hf35f)
	) name1521 (
		\P1_reg1_reg[21]/NET0131 ,
		\P1_reg2_reg[21]/NET0131 ,
		_w478_,
		_w488_,
		_w1984_
	);
	LUT4 #(
		.INIT('h6ccc)
	) name1522 (
		\P1_reg3_reg[14]/NET0131 ,
		\P1_reg3_reg[21]/NET0131 ,
		_w1821_,
		_w1824_,
		_w1985_
	);
	LUT4 #(
		.INIT('h3dfd)
	) name1523 (
		\P1_reg0_reg[21]/NET0131 ,
		_w478_,
		_w488_,
		_w1985_,
		_w1986_
	);
	LUT2 #(
		.INIT('h8)
	) name1524 (
		_w1984_,
		_w1986_,
		_w1987_
	);
	LUT2 #(
		.INIT('h7)
	) name1525 (
		_w1984_,
		_w1986_,
		_w1988_
	);
	LUT3 #(
		.INIT('h01)
	) name1526 (
		_w1748_,
		_w1982_,
		_w1987_,
		_w1989_
	);
	LUT3 #(
		.INIT('h45)
	) name1527 (
		_w1977_,
		_w1978_,
		_w1989_,
		_w1990_
	);
	LUT4 #(
		.INIT('h0054)
	) name1528 (
		_w1748_,
		_w1941_,
		_w1947_,
		_w1952_,
		_w1991_
	);
	LUT3 #(
		.INIT('h01)
	) name1529 (
		_w1748_,
		_w1957_,
		_w1962_,
		_w1992_
	);
	LUT3 #(
		.INIT('h23)
	) name1530 (
		_w1954_,
		_w1991_,
		_w1992_,
		_w1993_
	);
	LUT3 #(
		.INIT('hd0)
	) name1531 (
		_w1965_,
		_w1990_,
		_w1993_,
		_w1994_
	);
	LUT4 #(
		.INIT('h0054)
	) name1532 (
		_w1748_,
		_w1839_,
		_w1870_,
		_w1876_,
		_w1995_
	);
	LUT4 #(
		.INIT('h00fe)
	) name1533 (
		_w1748_,
		_w1899_,
		_w1904_,
		_w1995_,
		_w1996_
	);
	LUT4 #(
		.INIT('h0054)
	) name1534 (
		_w1748_,
		_w1907_,
		_w1929_,
		_w1936_,
		_w1997_
	);
	LUT4 #(
		.INIT('h00fe)
	) name1535 (
		_w1748_,
		_w1815_,
		_w1836_,
		_w1997_,
		_w1998_
	);
	LUT3 #(
		.INIT('hd0)
	) name1536 (
		_w1939_,
		_w1996_,
		_w1998_,
		_w1999_
	);
	LUT4 #(
		.INIT('h0455)
	) name1537 (
		_w1838_,
		_w1940_,
		_w1994_,
		_w1999_,
		_w2000_
	);
	LUT3 #(
		.INIT('h59)
	) name1538 (
		\P1_IR_reg[11]/NET0131 ,
		\P1_IR_reg[31]/NET0131 ,
		_w1718_,
		_w2001_
	);
	LUT3 #(
		.INIT('h10)
	) name1539 (
		_w1744_,
		_w1747_,
		_w2001_,
		_w2002_
	);
	LUT4 #(
		.INIT('h5956)
	) name1540 (
		\P2_datao_reg[11]/NET0131 ,
		\si[11]_pad ,
		_w547_,
		_w1916_,
		_w2003_
	);
	LUT3 #(
		.INIT('h23)
	) name1541 (
		_w1748_,
		_w2002_,
		_w2003_,
		_w2004_
	);
	LUT3 #(
		.INIT('h6a)
	) name1542 (
		\P1_reg3_reg[11]/NET0131 ,
		_w1817_,
		_w1818_,
		_w2005_
	);
	LUT4 #(
		.INIT('h37f7)
	) name1543 (
		\P1_reg1_reg[11]/NET0131 ,
		_w478_,
		_w488_,
		_w2005_,
		_w2006_
	);
	LUT4 #(
		.INIT('hf3f5)
	) name1544 (
		\P1_reg0_reg[11]/NET0131 ,
		\P1_reg2_reg[11]/NET0131 ,
		_w478_,
		_w488_,
		_w2007_
	);
	LUT2 #(
		.INIT('h8)
	) name1545 (
		_w2006_,
		_w2007_,
		_w2008_
	);
	LUT2 #(
		.INIT('h7)
	) name1546 (
		_w2006_,
		_w2007_,
		_w2009_
	);
	LUT4 #(
		.INIT('h2aaa)
	) name1547 (
		\P1_IR_reg[31]/NET0131 ,
		_w465_,
		_w466_,
		_w479_,
		_w2010_
	);
	LUT3 #(
		.INIT('he0)
	) name1548 (
		\P1_IR_reg[10]/NET0131 ,
		\P1_IR_reg[11]/NET0131 ,
		\P1_IR_reg[31]/NET0131 ,
		_w2011_
	);
	LUT3 #(
		.INIT('h56)
	) name1549 (
		\P1_IR_reg[12]/NET0131 ,
		_w2010_,
		_w2011_,
		_w2012_
	);
	LUT3 #(
		.INIT('h01)
	) name1550 (
		_w1744_,
		_w1747_,
		_w2012_,
		_w2013_
	);
	LUT4 #(
		.INIT('h1f00)
	) name1551 (
		_w1757_,
		_w1771_,
		_w1776_,
		_w1788_,
		_w2014_
	);
	LUT4 #(
		.INIT('h5956)
	) name1552 (
		\P2_datao_reg[12]/NET0131 ,
		\si[12]_pad ,
		_w547_,
		_w2014_,
		_w2015_
	);
	LUT3 #(
		.INIT('h23)
	) name1553 (
		_w1748_,
		_w2013_,
		_w2015_,
		_w2016_
	);
	LUT4 #(
		.INIT('hf35f)
	) name1554 (
		\P1_reg1_reg[12]/NET0131 ,
		\P1_reg2_reg[12]/NET0131 ,
		_w478_,
		_w488_,
		_w2017_
	);
	LUT4 #(
		.INIT('h6ccc)
	) name1555 (
		\P1_reg3_reg[11]/NET0131 ,
		\P1_reg3_reg[12]/NET0131 ,
		_w1817_,
		_w1818_,
		_w2018_
	);
	LUT4 #(
		.INIT('h3dfd)
	) name1556 (
		\P1_reg0_reg[12]/NET0131 ,
		_w478_,
		_w488_,
		_w2018_,
		_w2019_
	);
	LUT2 #(
		.INIT('h8)
	) name1557 (
		_w2017_,
		_w2019_,
		_w2020_
	);
	LUT2 #(
		.INIT('h7)
	) name1558 (
		_w2017_,
		_w2019_,
		_w2021_
	);
	LUT4 #(
		.INIT('hb0bb)
	) name1559 (
		_w2004_,
		_w2008_,
		_w2016_,
		_w2020_,
		_w2022_
	);
	LUT2 #(
		.INIT('h9)
	) name1560 (
		\P1_IR_reg[10]/NET0131 ,
		_w2010_,
		_w2023_
	);
	LUT3 #(
		.INIT('h10)
	) name1561 (
		_w1744_,
		_w1747_,
		_w2023_,
		_w2024_
	);
	LUT2 #(
		.INIT('h8)
	) name1562 (
		\P2_datao_reg[10]/NET0131 ,
		_w547_,
		_w2025_
	);
	LUT2 #(
		.INIT('h6)
	) name1563 (
		\P2_datao_reg[10]/NET0131 ,
		\si[10]_pad ,
		_w2026_
	);
	LUT4 #(
		.INIT('h1045)
	) name1564 (
		_w547_,
		_w1881_,
		_w1883_,
		_w2026_,
		_w2027_
	);
	LUT4 #(
		.INIT('h000e)
	) name1565 (
		_w1744_,
		_w1747_,
		_w2025_,
		_w2027_,
		_w2028_
	);
	LUT2 #(
		.INIT('h1)
	) name1566 (
		_w2024_,
		_w2028_,
		_w2029_
	);
	LUT4 #(
		.INIT('hf35f)
	) name1567 (
		\P1_reg1_reg[10]/NET0131 ,
		\P1_reg2_reg[10]/NET0131 ,
		_w478_,
		_w488_,
		_w2030_
	);
	LUT4 #(
		.INIT('h8000)
	) name1568 (
		\P1_reg3_reg[7]/NET0131 ,
		\P1_reg3_reg[8]/NET0131 ,
		\P1_reg3_reg[9]/NET0131 ,
		_w1817_,
		_w2031_
	);
	LUT3 #(
		.INIT('h32)
	) name1569 (
		\P1_reg3_reg[10]/NET0131 ,
		_w1819_,
		_w2031_,
		_w2032_
	);
	LUT4 #(
		.INIT('h3dfd)
	) name1570 (
		\P1_reg0_reg[10]/NET0131 ,
		_w478_,
		_w488_,
		_w2032_,
		_w2033_
	);
	LUT2 #(
		.INIT('h8)
	) name1571 (
		_w2030_,
		_w2033_,
		_w2034_
	);
	LUT2 #(
		.INIT('h7)
	) name1572 (
		_w2030_,
		_w2033_,
		_w2035_
	);
	LUT4 #(
		.INIT('he000)
	) name1573 (
		_w2024_,
		_w2028_,
		_w2030_,
		_w2033_,
		_w2036_
	);
	LUT4 #(
		.INIT('h0111)
	) name1574 (
		_w2024_,
		_w2028_,
		_w2030_,
		_w2033_,
		_w2037_
	);
	LUT3 #(
		.INIT('h39)
	) name1575 (
		\P1_IR_reg[31]/NET0131 ,
		\P1_IR_reg[9]/NET0131 ,
		_w467_,
		_w2038_
	);
	LUT4 #(
		.INIT('h5956)
	) name1576 (
		\P2_datao_reg[9]/NET0131 ,
		\si[9]_pad ,
		_w547_,
		_w1852_,
		_w2039_
	);
	LUT4 #(
		.INIT('h01ef)
	) name1577 (
		_w1744_,
		_w1747_,
		_w2038_,
		_w2039_,
		_w2040_
	);
	LUT4 #(
		.INIT('hf35f)
	) name1578 (
		\P1_reg1_reg[9]/NET0131 ,
		\P1_reg2_reg[9]/NET0131 ,
		_w478_,
		_w488_,
		_w2041_
	);
	LUT4 #(
		.INIT('h78f0)
	) name1579 (
		\P1_reg3_reg[7]/NET0131 ,
		\P1_reg3_reg[8]/NET0131 ,
		\P1_reg3_reg[9]/NET0131 ,
		_w1817_,
		_w2042_
	);
	LUT4 #(
		.INIT('h3dfd)
	) name1580 (
		\P1_reg0_reg[9]/NET0131 ,
		_w478_,
		_w488_,
		_w2042_,
		_w2043_
	);
	LUT2 #(
		.INIT('h8)
	) name1581 (
		_w2041_,
		_w2043_,
		_w2044_
	);
	LUT2 #(
		.INIT('h7)
	) name1582 (
		_w2041_,
		_w2043_,
		_w2045_
	);
	LUT3 #(
		.INIT('h2a)
	) name1583 (
		_w2040_,
		_w2041_,
		_w2043_,
		_w2046_
	);
	LUT3 #(
		.INIT('h54)
	) name1584 (
		_w2036_,
		_w2037_,
		_w2046_,
		_w2047_
	);
	LUT4 #(
		.INIT('h20f2)
	) name1585 (
		_w2004_,
		_w2008_,
		_w2016_,
		_w2020_,
		_w2048_
	);
	LUT3 #(
		.INIT('h07)
	) name1586 (
		_w2022_,
		_w2047_,
		_w2048_,
		_w2049_
	);
	LUT2 #(
		.INIT('h6)
	) name1587 (
		\P1_reg3_reg[3]/NET0131 ,
		\P1_reg3_reg[4]/NET0131 ,
		_w2050_
	);
	LUT4 #(
		.INIT('h3dfd)
	) name1588 (
		\P1_reg0_reg[4]/NET0131 ,
		_w478_,
		_w488_,
		_w2050_,
		_w2051_
	);
	LUT4 #(
		.INIT('hf35f)
	) name1589 (
		\P1_reg1_reg[4]/NET0131 ,
		\P1_reg2_reg[4]/NET0131 ,
		_w478_,
		_w488_,
		_w2052_
	);
	LUT2 #(
		.INIT('h8)
	) name1590 (
		_w2051_,
		_w2052_,
		_w2053_
	);
	LUT2 #(
		.INIT('h7)
	) name1591 (
		_w2051_,
		_w2052_,
		_w2054_
	);
	LUT4 #(
		.INIT('h5659)
	) name1592 (
		\P2_datao_reg[4]/NET0131 ,
		\si[4]_pad ,
		_w547_,
		_w1764_,
		_w2055_
	);
	LUT3 #(
		.INIT('h39)
	) name1593 (
		\P1_IR_reg[31]/NET0131 ,
		\P1_IR_reg[4]/NET0131 ,
		_w465_,
		_w2056_
	);
	LUT4 #(
		.INIT('hf1e0)
	) name1594 (
		_w1744_,
		_w1747_,
		_w2055_,
		_w2056_,
		_w2057_
	);
	LUT3 #(
		.INIT('h80)
	) name1595 (
		_w2051_,
		_w2052_,
		_w2057_,
		_w2058_
	);
	LUT4 #(
		.INIT('h3f5f)
	) name1596 (
		\P1_reg1_reg[2]/NET0131 ,
		\P1_reg3_reg[2]/NET0131 ,
		_w478_,
		_w488_,
		_w2059_
	);
	LUT4 #(
		.INIT('hf3f5)
	) name1597 (
		\P1_reg0_reg[2]/NET0131 ,
		\P1_reg2_reg[2]/NET0131 ,
		_w478_,
		_w488_,
		_w2060_
	);
	LUT2 #(
		.INIT('h8)
	) name1598 (
		_w2059_,
		_w2060_,
		_w2061_
	);
	LUT2 #(
		.INIT('h7)
	) name1599 (
		_w2059_,
		_w2060_,
		_w2062_
	);
	LUT4 #(
		.INIT('h5659)
	) name1600 (
		\P2_datao_reg[2]/NET0131 ,
		\si[2]_pad ,
		_w547_,
		_w1762_,
		_w2063_
	);
	LUT4 #(
		.INIT('h1ef0)
	) name1601 (
		\P1_IR_reg[0]/NET0131 ,
		\P1_IR_reg[1]/NET0131 ,
		\P1_IR_reg[2]/NET0131 ,
		\P1_IR_reg[31]/NET0131 ,
		_w2064_
	);
	LUT4 #(
		.INIT('he0f1)
	) name1602 (
		_w1744_,
		_w1747_,
		_w2063_,
		_w2064_,
		_w2065_
	);
	LUT3 #(
		.INIT('h80)
	) name1603 (
		_w2059_,
		_w2060_,
		_w2065_,
		_w2066_
	);
	LUT3 #(
		.INIT('h17)
	) name1604 (
		\P2_datao_reg[2]/NET0131 ,
		\si[2]_pad ,
		_w1762_,
		_w2067_
	);
	LUT4 #(
		.INIT('h5956)
	) name1605 (
		\P2_datao_reg[3]/NET0131 ,
		\si[3]_pad ,
		_w547_,
		_w2067_,
		_w2068_
	);
	LUT4 #(
		.INIT('h01ff)
	) name1606 (
		\P1_IR_reg[0]/NET0131 ,
		\P1_IR_reg[1]/NET0131 ,
		\P1_IR_reg[2]/NET0131 ,
		\P1_IR_reg[31]/NET0131 ,
		_w2069_
	);
	LUT2 #(
		.INIT('h9)
	) name1607 (
		\P1_IR_reg[3]/NET0131 ,
		_w2069_,
		_w2070_
	);
	LUT4 #(
		.INIT('he0f1)
	) name1608 (
		_w1744_,
		_w1747_,
		_w2068_,
		_w2070_,
		_w2071_
	);
	LUT3 #(
		.INIT('h80)
	) name1609 (
		_w489_,
		_w491_,
		_w2071_,
		_w2072_
	);
	LUT2 #(
		.INIT('h1)
	) name1610 (
		_w2066_,
		_w2072_,
		_w2073_
	);
	LUT3 #(
		.INIT('h07)
	) name1611 (
		_w2059_,
		_w2060_,
		_w2065_,
		_w2074_
	);
	LUT4 #(
		.INIT('h35ff)
	) name1612 (
		\P1_reg2_reg[1]/NET0131 ,
		\P1_reg3_reg[1]/NET0131 ,
		_w478_,
		_w488_,
		_w2075_
	);
	LUT4 #(
		.INIT('hff35)
	) name1613 (
		\P1_reg0_reg[1]/NET0131 ,
		\P1_reg1_reg[1]/NET0131 ,
		_w478_,
		_w488_,
		_w2076_
	);
	LUT2 #(
		.INIT('h8)
	) name1614 (
		_w2075_,
		_w2076_,
		_w2077_
	);
	LUT2 #(
		.INIT('h7)
	) name1615 (
		_w2075_,
		_w2076_,
		_w2078_
	);
	LUT3 #(
		.INIT('h6c)
	) name1616 (
		\P1_IR_reg[0]/NET0131 ,
		\P1_IR_reg[1]/NET0131 ,
		\P1_IR_reg[31]/NET0131 ,
		_w2079_
	);
	LUT4 #(
		.INIT('ha9a6)
	) name1617 (
		\P2_datao_reg[1]/NET0131 ,
		\si[1]_pad ,
		_w547_,
		_w1761_,
		_w2080_
	);
	LUT4 #(
		.INIT('h01ef)
	) name1618 (
		_w1744_,
		_w1747_,
		_w2079_,
		_w2080_,
		_w2081_
	);
	LUT3 #(
		.INIT('h07)
	) name1619 (
		_w2075_,
		_w2076_,
		_w2081_,
		_w2082_
	);
	LUT3 #(
		.INIT('h80)
	) name1620 (
		_w2075_,
		_w2076_,
		_w2081_,
		_w2083_
	);
	LUT4 #(
		.INIT('hff35)
	) name1621 (
		\P1_reg0_reg[0]/NET0131 ,
		\P1_reg1_reg[0]/NET0131 ,
		_w478_,
		_w488_,
		_w2084_
	);
	LUT4 #(
		.INIT('h35ff)
	) name1622 (
		\P1_reg2_reg[0]/NET0131 ,
		\P1_reg3_reg[0]/NET0131 ,
		_w478_,
		_w488_,
		_w2085_
	);
	LUT2 #(
		.INIT('h8)
	) name1623 (
		_w2084_,
		_w2085_,
		_w2086_
	);
	LUT2 #(
		.INIT('h7)
	) name1624 (
		_w2084_,
		_w2085_,
		_w2087_
	);
	LUT3 #(
		.INIT('ha6)
	) name1625 (
		\P2_datao_reg[0]/NET0131 ,
		\si[0]_pad ,
		_w547_,
		_w2088_
	);
	LUT4 #(
		.INIT('h01fd)
	) name1626 (
		\P1_IR_reg[0]/NET0131 ,
		_w1744_,
		_w1747_,
		_w2088_,
		_w2089_
	);
	LUT3 #(
		.INIT('h07)
	) name1627 (
		_w2084_,
		_w2085_,
		_w2089_,
		_w2090_
	);
	LUT3 #(
		.INIT('h45)
	) name1628 (
		_w2082_,
		_w2083_,
		_w2090_,
		_w2091_
	);
	LUT4 #(
		.INIT('h4054)
	) name1629 (
		_w2074_,
		_w2077_,
		_w2081_,
		_w2090_,
		_w2092_
	);
	LUT3 #(
		.INIT('h07)
	) name1630 (
		_w2051_,
		_w2052_,
		_w2057_,
		_w2093_
	);
	LUT3 #(
		.INIT('h07)
	) name1631 (
		_w489_,
		_w491_,
		_w2071_,
		_w2094_
	);
	LUT2 #(
		.INIT('h1)
	) name1632 (
		_w2093_,
		_w2094_,
		_w2095_
	);
	LUT4 #(
		.INIT('h0455)
	) name1633 (
		_w2058_,
		_w2073_,
		_w2092_,
		_w2095_,
		_w2096_
	);
	LUT4 #(
		.INIT('h2aaa)
	) name1634 (
		\P1_IR_reg[31]/NET0131 ,
		_w464_,
		_w465_,
		_w466_,
		_w2097_
	);
	LUT2 #(
		.INIT('h6)
	) name1635 (
		\P1_IR_reg[8]/NET0131 ,
		_w2097_,
		_w2098_
	);
	LUT3 #(
		.INIT('h01)
	) name1636 (
		_w1744_,
		_w1747_,
		_w2098_,
		_w2099_
	);
	LUT2 #(
		.INIT('h8)
	) name1637 (
		\P2_datao_reg[8]/NET0131 ,
		_w547_,
		_w2100_
	);
	LUT2 #(
		.INIT('h6)
	) name1638 (
		\P2_datao_reg[8]/NET0131 ,
		\si[8]_pad ,
		_w2101_
	);
	LUT4 #(
		.INIT('h0154)
	) name1639 (
		_w547_,
		_w1757_,
		_w1771_,
		_w2101_,
		_w2102_
	);
	LUT4 #(
		.INIT('h000e)
	) name1640 (
		_w1744_,
		_w1747_,
		_w2100_,
		_w2102_,
		_w2103_
	);
	LUT2 #(
		.INIT('h1)
	) name1641 (
		_w2099_,
		_w2103_,
		_w2104_
	);
	LUT4 #(
		.INIT('hf35f)
	) name1642 (
		\P1_reg1_reg[8]/NET0131 ,
		\P1_reg2_reg[8]/NET0131 ,
		_w478_,
		_w488_,
		_w2105_
	);
	LUT3 #(
		.INIT('h6c)
	) name1643 (
		\P1_reg3_reg[7]/NET0131 ,
		\P1_reg3_reg[8]/NET0131 ,
		_w1817_,
		_w2106_
	);
	LUT4 #(
		.INIT('h3dfd)
	) name1644 (
		\P1_reg0_reg[8]/NET0131 ,
		_w478_,
		_w488_,
		_w2106_,
		_w2107_
	);
	LUT2 #(
		.INIT('h8)
	) name1645 (
		_w2105_,
		_w2107_,
		_w2108_
	);
	LUT2 #(
		.INIT('h7)
	) name1646 (
		_w2105_,
		_w2107_,
		_w2109_
	);
	LUT4 #(
		.INIT('he000)
	) name1647 (
		_w2099_,
		_w2103_,
		_w2105_,
		_w2107_,
		_w2110_
	);
	LUT4 #(
		.INIT('h7555)
	) name1648 (
		\P1_IR_reg[31]/NET0131 ,
		\P1_IR_reg[6]/NET0131 ,
		_w465_,
		_w466_,
		_w2111_
	);
	LUT2 #(
		.INIT('h9)
	) name1649 (
		\P1_IR_reg[7]/NET0131 ,
		_w2111_,
		_w2112_
	);
	LUT4 #(
		.INIT('h5956)
	) name1650 (
		\P2_datao_reg[7]/NET0131 ,
		\si[7]_pad ,
		_w547_,
		_w1912_,
		_w2113_
	);
	LUT4 #(
		.INIT('h10fe)
	) name1651 (
		_w1744_,
		_w1747_,
		_w2112_,
		_w2113_,
		_w2114_
	);
	LUT2 #(
		.INIT('h6)
	) name1652 (
		\P1_reg3_reg[7]/NET0131 ,
		_w1817_,
		_w2115_
	);
	LUT4 #(
		.INIT('h3dfd)
	) name1653 (
		\P1_reg0_reg[7]/NET0131 ,
		_w478_,
		_w488_,
		_w2115_,
		_w2116_
	);
	LUT4 #(
		.INIT('hf35f)
	) name1654 (
		\P1_reg1_reg[7]/NET0131 ,
		\P1_reg2_reg[7]/NET0131 ,
		_w478_,
		_w488_,
		_w2117_
	);
	LUT2 #(
		.INIT('h8)
	) name1655 (
		_w2116_,
		_w2117_,
		_w2118_
	);
	LUT2 #(
		.INIT('h7)
	) name1656 (
		_w2116_,
		_w2117_,
		_w2119_
	);
	LUT3 #(
		.INIT('h40)
	) name1657 (
		_w2114_,
		_w2116_,
		_w2117_,
		_w2120_
	);
	LUT2 #(
		.INIT('h1)
	) name1658 (
		_w2110_,
		_w2120_,
		_w2121_
	);
	LUT4 #(
		.INIT('h5956)
	) name1659 (
		\P2_datao_reg[6]/NET0131 ,
		\si[6]_pad ,
		_w547_,
		_w1879_,
		_w2122_
	);
	LUT4 #(
		.INIT('hc666)
	) name1660 (
		\P1_IR_reg[31]/NET0131 ,
		\P1_IR_reg[6]/NET0131 ,
		_w465_,
		_w466_,
		_w2123_
	);
	LUT4 #(
		.INIT('he0f1)
	) name1661 (
		_w1744_,
		_w1747_,
		_w2122_,
		_w2123_,
		_w2124_
	);
	LUT4 #(
		.INIT('hf35f)
	) name1662 (
		\P1_reg1_reg[6]/NET0131 ,
		\P1_reg2_reg[6]/NET0131 ,
		_w478_,
		_w488_,
		_w2125_
	);
	LUT4 #(
		.INIT('h7f80)
	) name1663 (
		\P1_reg3_reg[3]/NET0131 ,
		\P1_reg3_reg[4]/NET0131 ,
		\P1_reg3_reg[5]/NET0131 ,
		\P1_reg3_reg[6]/NET0131 ,
		_w2126_
	);
	LUT4 #(
		.INIT('h3dfd)
	) name1664 (
		\P1_reg0_reg[6]/NET0131 ,
		_w478_,
		_w488_,
		_w2126_,
		_w2127_
	);
	LUT2 #(
		.INIT('h8)
	) name1665 (
		_w2125_,
		_w2127_,
		_w2128_
	);
	LUT2 #(
		.INIT('h7)
	) name1666 (
		_w2125_,
		_w2127_,
		_w2129_
	);
	LUT3 #(
		.INIT('h80)
	) name1667 (
		_w2124_,
		_w2125_,
		_w2127_,
		_w2130_
	);
	LUT3 #(
		.INIT('he8)
	) name1668 (
		\P2_datao_reg[4]/NET0131 ,
		\si[4]_pad ,
		_w1764_,
		_w2131_
	);
	LUT4 #(
		.INIT('h5659)
	) name1669 (
		\P2_datao_reg[5]/NET0131 ,
		\si[5]_pad ,
		_w547_,
		_w2131_,
		_w2132_
	);
	LUT4 #(
		.INIT('h785a)
	) name1670 (
		\P1_IR_reg[31]/NET0131 ,
		\P1_IR_reg[4]/NET0131 ,
		\P1_IR_reg[5]/NET0131 ,
		_w465_,
		_w2133_
	);
	LUT4 #(
		.INIT('he0f1)
	) name1671 (
		_w1744_,
		_w1747_,
		_w2132_,
		_w2133_,
		_w2134_
	);
	LUT4 #(
		.INIT('hf35f)
	) name1672 (
		\P1_reg1_reg[5]/NET0131 ,
		\P1_reg2_reg[5]/NET0131 ,
		_w478_,
		_w488_,
		_w2135_
	);
	LUT3 #(
		.INIT('h78)
	) name1673 (
		\P1_reg3_reg[3]/NET0131 ,
		\P1_reg3_reg[4]/NET0131 ,
		\P1_reg3_reg[5]/NET0131 ,
		_w2136_
	);
	LUT4 #(
		.INIT('h3dfd)
	) name1674 (
		\P1_reg0_reg[5]/NET0131 ,
		_w478_,
		_w488_,
		_w2136_,
		_w2137_
	);
	LUT2 #(
		.INIT('h8)
	) name1675 (
		_w2135_,
		_w2137_,
		_w2138_
	);
	LUT2 #(
		.INIT('h7)
	) name1676 (
		_w2135_,
		_w2137_,
		_w2139_
	);
	LUT3 #(
		.INIT('h80)
	) name1677 (
		_w2134_,
		_w2135_,
		_w2137_,
		_w2140_
	);
	LUT2 #(
		.INIT('h1)
	) name1678 (
		_w2130_,
		_w2140_,
		_w2141_
	);
	LUT4 #(
		.INIT('h0001)
	) name1679 (
		_w2110_,
		_w2120_,
		_w2130_,
		_w2140_,
		_w2142_
	);
	LUT3 #(
		.INIT('h15)
	) name1680 (
		_w2124_,
		_w2125_,
		_w2127_,
		_w2143_
	);
	LUT3 #(
		.INIT('h15)
	) name1681 (
		_w2134_,
		_w2135_,
		_w2137_,
		_w2144_
	);
	LUT3 #(
		.INIT('h54)
	) name1682 (
		_w2130_,
		_w2143_,
		_w2144_,
		_w2145_
	);
	LUT4 #(
		.INIT('h0111)
	) name1683 (
		_w2099_,
		_w2103_,
		_w2105_,
		_w2107_,
		_w2146_
	);
	LUT3 #(
		.INIT('h2a)
	) name1684 (
		_w2114_,
		_w2116_,
		_w2117_,
		_w2147_
	);
	LUT3 #(
		.INIT('h23)
	) name1685 (
		_w2110_,
		_w2146_,
		_w2147_,
		_w2148_
	);
	LUT3 #(
		.INIT('h70)
	) name1686 (
		_w2121_,
		_w2145_,
		_w2148_,
		_w2149_
	);
	LUT3 #(
		.INIT('h40)
	) name1687 (
		_w2040_,
		_w2041_,
		_w2043_,
		_w2150_
	);
	LUT2 #(
		.INIT('h1)
	) name1688 (
		_w2036_,
		_w2150_,
		_w2151_
	);
	LUT2 #(
		.INIT('h8)
	) name1689 (
		_w2022_,
		_w2151_,
		_w2152_
	);
	LUT4 #(
		.INIT('h8f00)
	) name1690 (
		_w2096_,
		_w2142_,
		_w2149_,
		_w2152_,
		_w2153_
	);
	LUT4 #(
		.INIT('h5956)
	) name1691 (
		\P2_datao_reg[20]/NET0131 ,
		\si[20]_pad ,
		_w547_,
		_w1794_,
		_w2154_
	);
	LUT2 #(
		.INIT('h1)
	) name1692 (
		_w1748_,
		_w2154_,
		_w2155_
	);
	LUT3 #(
		.INIT('h80)
	) name1693 (
		\P1_reg3_reg[14]/NET0131 ,
		\P1_reg3_reg[15]/NET0131 ,
		_w1821_,
		_w2156_
	);
	LUT4 #(
		.INIT('h8000)
	) name1694 (
		\P1_reg3_reg[14]/NET0131 ,
		\P1_reg3_reg[15]/NET0131 ,
		_w1821_,
		_w1822_,
		_w2157_
	);
	LUT4 #(
		.INIT('h070f)
	) name1695 (
		\P1_reg3_reg[18]/NET0131 ,
		\P1_reg3_reg[19]/NET0131 ,
		\P1_reg3_reg[20]/NET0131 ,
		_w2157_,
		_w2158_
	);
	LUT2 #(
		.INIT('h1)
	) name1696 (
		_w1825_,
		_w2158_,
		_w2159_
	);
	LUT4 #(
		.INIT('h0008)
	) name1697 (
		_w478_,
		_w488_,
		_w1825_,
		_w2158_,
		_w2160_
	);
	LUT3 #(
		.INIT('h08)
	) name1698 (
		\P1_reg1_reg[20]/NET0131 ,
		_w478_,
		_w488_,
		_w2161_
	);
	LUT4 #(
		.INIT('hf3f5)
	) name1699 (
		\P1_reg0_reg[20]/NET0131 ,
		\P1_reg2_reg[20]/NET0131 ,
		_w478_,
		_w488_,
		_w2162_
	);
	LUT3 #(
		.INIT('h10)
	) name1700 (
		_w2161_,
		_w2160_,
		_w2162_,
		_w2163_
	);
	LUT3 #(
		.INIT('hef)
	) name1701 (
		_w2161_,
		_w2160_,
		_w2162_,
		_w2164_
	);
	LUT3 #(
		.INIT('he0)
	) name1702 (
		_w1748_,
		_w2154_,
		_w2163_,
		_w2165_
	);
	LUT4 #(
		.INIT('h2aaa)
	) name1703 (
		\P1_IR_reg[31]/NET0131 ,
		_w1718_,
		_w1719_,
		_w1720_,
		_w2166_
	);
	LUT2 #(
		.INIT('h9)
	) name1704 (
		\P1_IR_reg[19]/NET0131 ,
		_w2166_,
		_w2167_
	);
	LUT3 #(
		.INIT('h10)
	) name1705 (
		_w1744_,
		_w1747_,
		_w2167_,
		_w2168_
	);
	LUT4 #(
		.INIT('h3700)
	) name1706 (
		_w1918_,
		_w1920_,
		_w1924_,
		_w1925_,
		_w2169_
	);
	LUT4 #(
		.INIT('h5956)
	) name1707 (
		\P2_datao_reg[19]/NET0131 ,
		\si[19]_pad ,
		_w547_,
		_w2169_,
		_w2170_
	);
	LUT3 #(
		.INIT('h23)
	) name1708 (
		_w1748_,
		_w2168_,
		_w2170_,
		_w2171_
	);
	LUT3 #(
		.INIT('h6c)
	) name1709 (
		\P1_reg3_reg[18]/NET0131 ,
		\P1_reg3_reg[19]/NET0131 ,
		_w2157_,
		_w2172_
	);
	LUT4 #(
		.INIT('h37f7)
	) name1710 (
		\P1_reg1_reg[19]/NET0131 ,
		_w478_,
		_w488_,
		_w2172_,
		_w2173_
	);
	LUT4 #(
		.INIT('hf3f5)
	) name1711 (
		\P1_reg0_reg[19]/NET0131 ,
		\P1_reg2_reg[19]/NET0131 ,
		_w478_,
		_w488_,
		_w2174_
	);
	LUT2 #(
		.INIT('h8)
	) name1712 (
		_w2173_,
		_w2174_,
		_w2175_
	);
	LUT2 #(
		.INIT('h7)
	) name1713 (
		_w2173_,
		_w2174_,
		_w2176_
	);
	LUT4 #(
		.INIT('hdc00)
	) name1714 (
		_w1748_,
		_w2168_,
		_w2170_,
		_w2175_,
		_w2177_
	);
	LUT4 #(
		.INIT('h5999)
	) name1715 (
		\P1_IR_reg[17]/NET0131 ,
		\P1_IR_reg[31]/NET0131 ,
		_w467_,
		_w471_,
		_w2178_
	);
	LUT3 #(
		.INIT('h10)
	) name1716 (
		_w1744_,
		_w1747_,
		_w2178_,
		_w2179_
	);
	LUT2 #(
		.INIT('h8)
	) name1717 (
		\P2_datao_reg[17]/NET0131 ,
		_w547_,
		_w2180_
	);
	LUT2 #(
		.INIT('h6)
	) name1718 (
		\P2_datao_reg[17]/NET0131 ,
		\si[17]_pad ,
		_w2181_
	);
	LUT4 #(
		.INIT('h0451)
	) name1719 (
		_w547_,
		_w1859_,
		_w1980_,
		_w2181_,
		_w2182_
	);
	LUT4 #(
		.INIT('h3332)
	) name1720 (
		_w1748_,
		_w2179_,
		_w2180_,
		_w2182_,
		_w2183_
	);
	LUT4 #(
		.INIT('hf35f)
	) name1721 (
		\P1_reg1_reg[17]/NET0131 ,
		\P1_reg2_reg[17]/NET0131 ,
		_w478_,
		_w488_,
		_w2184_
	);
	LUT3 #(
		.INIT('h6c)
	) name1722 (
		\P1_reg3_reg[16]/NET0131 ,
		\P1_reg3_reg[17]/NET0131 ,
		_w2156_,
		_w2185_
	);
	LUT4 #(
		.INIT('h3dfd)
	) name1723 (
		\P1_reg0_reg[17]/NET0131 ,
		_w478_,
		_w488_,
		_w2185_,
		_w2186_
	);
	LUT2 #(
		.INIT('h8)
	) name1724 (
		_w2184_,
		_w2186_,
		_w2187_
	);
	LUT2 #(
		.INIT('h7)
	) name1725 (
		_w2184_,
		_w2186_,
		_w2188_
	);
	LUT4 #(
		.INIT('h0001)
	) name1726 (
		\P1_IR_reg[14]/NET0131 ,
		\P1_IR_reg[15]/NET0131 ,
		\P1_IR_reg[16]/NET0131 ,
		\P1_IR_reg[17]/NET0131 ,
		_w2189_
	);
	LUT2 #(
		.INIT('h2)
	) name1727 (
		\P1_IR_reg[31]/NET0131 ,
		_w2189_,
		_w2190_
	);
	LUT4 #(
		.INIT('h55a6)
	) name1728 (
		\P1_IR_reg[18]/NET0131 ,
		\P1_IR_reg[31]/NET0131 ,
		_w480_,
		_w2190_,
		_w2191_
	);
	LUT3 #(
		.INIT('h01)
	) name1729 (
		_w1744_,
		_w1747_,
		_w2191_,
		_w2192_
	);
	LUT2 #(
		.INIT('h8)
	) name1730 (
		\P2_datao_reg[18]/NET0131 ,
		_w547_,
		_w2193_
	);
	LUT2 #(
		.INIT('h6)
	) name1731 (
		\P2_datao_reg[18]/NET0131 ,
		\si[18]_pad ,
		_w2194_
	);
	LUT4 #(
		.INIT('h1045)
	) name1732 (
		_w547_,
		_w1886_,
		_w1890_,
		_w2194_,
		_w2195_
	);
	LUT4 #(
		.INIT('h3332)
	) name1733 (
		_w1748_,
		_w2192_,
		_w2193_,
		_w2195_,
		_w2196_
	);
	LUT2 #(
		.INIT('h6)
	) name1734 (
		\P1_reg3_reg[18]/NET0131 ,
		_w2157_,
		_w2197_
	);
	LUT4 #(
		.INIT('h3dfd)
	) name1735 (
		\P1_reg0_reg[18]/NET0131 ,
		_w478_,
		_w488_,
		_w2197_,
		_w2198_
	);
	LUT4 #(
		.INIT('hf35f)
	) name1736 (
		\P1_reg1_reg[18]/NET0131 ,
		\P1_reg2_reg[18]/NET0131 ,
		_w478_,
		_w488_,
		_w2199_
	);
	LUT2 #(
		.INIT('h8)
	) name1737 (
		_w2198_,
		_w2199_,
		_w2200_
	);
	LUT2 #(
		.INIT('h7)
	) name1738 (
		_w2198_,
		_w2199_,
		_w2201_
	);
	LUT2 #(
		.INIT('h4)
	) name1739 (
		_w2196_,
		_w2200_,
		_w2202_
	);
	LUT4 #(
		.INIT('hb0bb)
	) name1740 (
		_w2183_,
		_w2187_,
		_w2196_,
		_w2200_,
		_w2203_
	);
	LUT3 #(
		.INIT('h10)
	) name1741 (
		_w2165_,
		_w2177_,
		_w2203_,
		_w2204_
	);
	LUT3 #(
		.INIT('ha6)
	) name1742 (
		\P1_IR_reg[14]/NET0131 ,
		\P1_IR_reg[31]/NET0131 ,
		_w480_,
		_w2205_
	);
	LUT3 #(
		.INIT('h01)
	) name1743 (
		_w1744_,
		_w1747_,
		_w2205_,
		_w2206_
	);
	LUT4 #(
		.INIT('h5956)
	) name1744 (
		\P2_datao_reg[14]/NET0131 ,
		\si[14]_pad ,
		_w547_,
		_w1968_,
		_w2207_
	);
	LUT3 #(
		.INIT('h23)
	) name1745 (
		_w1748_,
		_w2206_,
		_w2207_,
		_w2208_
	);
	LUT2 #(
		.INIT('h6)
	) name1746 (
		\P1_reg3_reg[14]/NET0131 ,
		_w1821_,
		_w2209_
	);
	LUT4 #(
		.INIT('h1fdf)
	) name1747 (
		\P1_reg2_reg[14]/NET0131 ,
		_w478_,
		_w488_,
		_w2209_,
		_w2210_
	);
	LUT4 #(
		.INIT('hff35)
	) name1748 (
		\P1_reg0_reg[14]/NET0131 ,
		\P1_reg1_reg[14]/NET0131 ,
		_w478_,
		_w488_,
		_w2211_
	);
	LUT2 #(
		.INIT('h8)
	) name1749 (
		_w2210_,
		_w2211_,
		_w2212_
	);
	LUT2 #(
		.INIT('h7)
	) name1750 (
		_w2210_,
		_w2211_,
		_w2213_
	);
	LUT2 #(
		.INIT('h1)
	) name1751 (
		\P1_IR_reg[12]/NET0131 ,
		\P1_IR_reg[9]/NET0131 ,
		_w2214_
	);
	LUT4 #(
		.INIT('h0d05)
	) name1752 (
		\P1_IR_reg[31]/NET0131 ,
		_w467_,
		_w2011_,
		_w2214_,
		_w2215_
	);
	LUT2 #(
		.INIT('h9)
	) name1753 (
		\P1_IR_reg[13]/NET0131 ,
		_w2215_,
		_w2216_
	);
	LUT3 #(
		.INIT('h01)
	) name1754 (
		_w1744_,
		_w1747_,
		_w2216_,
		_w2217_
	);
	LUT4 #(
		.INIT('h5956)
	) name1755 (
		\P2_datao_reg[13]/NET0131 ,
		\si[13]_pad ,
		_w547_,
		_w1979_,
		_w2218_
	);
	LUT3 #(
		.INIT('h23)
	) name1756 (
		_w1748_,
		_w2217_,
		_w2218_,
		_w2219_
	);
	LUT4 #(
		.INIT('h6aaa)
	) name1757 (
		\P1_reg3_reg[13]/NET0131 ,
		_w1817_,
		_w1818_,
		_w1820_,
		_w2220_
	);
	LUT4 #(
		.INIT('h3dfd)
	) name1758 (
		\P1_reg0_reg[13]/NET0131 ,
		_w478_,
		_w488_,
		_w2220_,
		_w2221_
	);
	LUT4 #(
		.INIT('hf35f)
	) name1759 (
		\P1_reg1_reg[13]/NET0131 ,
		\P1_reg2_reg[13]/NET0131 ,
		_w478_,
		_w488_,
		_w2222_
	);
	LUT2 #(
		.INIT('h8)
	) name1760 (
		_w2221_,
		_w2222_,
		_w2223_
	);
	LUT2 #(
		.INIT('h7)
	) name1761 (
		_w2221_,
		_w2222_,
		_w2224_
	);
	LUT4 #(
		.INIT('hb0bb)
	) name1762 (
		_w2208_,
		_w2212_,
		_w2219_,
		_w2223_,
		_w2225_
	);
	LUT4 #(
		.INIT('ha666)
	) name1763 (
		\P1_IR_reg[16]/NET0131 ,
		\P1_IR_reg[31]/NET0131 ,
		_w468_,
		_w480_,
		_w2226_
	);
	LUT3 #(
		.INIT('h01)
	) name1764 (
		_w1744_,
		_w1747_,
		_w2226_,
		_w2227_
	);
	LUT2 #(
		.INIT('h8)
	) name1765 (
		\P2_datao_reg[16]/NET0131 ,
		_w547_,
		_w2228_
	);
	LUT2 #(
		.INIT('h6)
	) name1766 (
		\P2_datao_reg[16]/NET0131 ,
		\si[16]_pad ,
		_w2229_
	);
	LUT4 #(
		.INIT('h1045)
	) name1767 (
		_w547_,
		_w1782_,
		_w1793_,
		_w2229_,
		_w2230_
	);
	LUT4 #(
		.INIT('h3332)
	) name1768 (
		_w1748_,
		_w2227_,
		_w2228_,
		_w2230_,
		_w2231_
	);
	LUT4 #(
		.INIT('hf35f)
	) name1769 (
		\P1_reg1_reg[16]/NET0131 ,
		\P1_reg2_reg[16]/NET0131 ,
		_w478_,
		_w488_,
		_w2232_
	);
	LUT4 #(
		.INIT('h78f0)
	) name1770 (
		\P1_reg3_reg[14]/NET0131 ,
		\P1_reg3_reg[15]/NET0131 ,
		\P1_reg3_reg[16]/NET0131 ,
		_w1821_,
		_w2233_
	);
	LUT4 #(
		.INIT('h3dfd)
	) name1771 (
		\P1_reg0_reg[16]/NET0131 ,
		_w478_,
		_w488_,
		_w2233_,
		_w2234_
	);
	LUT2 #(
		.INIT('h8)
	) name1772 (
		_w2232_,
		_w2234_,
		_w2235_
	);
	LUT2 #(
		.INIT('h7)
	) name1773 (
		_w2232_,
		_w2234_,
		_w2236_
	);
	LUT4 #(
		.INIT('ha666)
	) name1774 (
		\P1_IR_reg[15]/NET0131 ,
		\P1_IR_reg[31]/NET0131 ,
		_w1718_,
		_w1719_,
		_w2237_
	);
	LUT3 #(
		.INIT('h01)
	) name1775 (
		_w1744_,
		_w1747_,
		_w2237_,
		_w2238_
	);
	LUT2 #(
		.INIT('h8)
	) name1776 (
		\P2_datao_reg[15]/NET0131 ,
		_w547_,
		_w2239_
	);
	LUT2 #(
		.INIT('h6)
	) name1777 (
		\P2_datao_reg[15]/NET0131 ,
		\si[15]_pad ,
		_w2240_
	);
	LUT4 #(
		.INIT('h0154)
	) name1778 (
		_w547_,
		_w1918_,
		_w1924_,
		_w2240_,
		_w2241_
	);
	LUT4 #(
		.INIT('h3332)
	) name1779 (
		_w1748_,
		_w2238_,
		_w2239_,
		_w2241_,
		_w2242_
	);
	LUT3 #(
		.INIT('h6c)
	) name1780 (
		\P1_reg3_reg[14]/NET0131 ,
		\P1_reg3_reg[15]/NET0131 ,
		_w1821_,
		_w2243_
	);
	LUT4 #(
		.INIT('h1fdf)
	) name1781 (
		\P1_reg2_reg[15]/NET0131 ,
		_w478_,
		_w488_,
		_w2243_,
		_w2244_
	);
	LUT4 #(
		.INIT('hff35)
	) name1782 (
		\P1_reg0_reg[15]/NET0131 ,
		\P1_reg1_reg[15]/NET0131 ,
		_w478_,
		_w488_,
		_w2245_
	);
	LUT2 #(
		.INIT('h8)
	) name1783 (
		_w2244_,
		_w2245_,
		_w2246_
	);
	LUT2 #(
		.INIT('h7)
	) name1784 (
		_w2244_,
		_w2245_,
		_w2247_
	);
	LUT4 #(
		.INIT('hb0bb)
	) name1785 (
		_w2231_,
		_w2235_,
		_w2242_,
		_w2246_,
		_w2248_
	);
	LUT2 #(
		.INIT('h8)
	) name1786 (
		_w2225_,
		_w2248_,
		_w2249_
	);
	LUT2 #(
		.INIT('h8)
	) name1787 (
		_w2204_,
		_w2249_,
		_w2250_
	);
	LUT4 #(
		.INIT('h22b2)
	) name1788 (
		_w2208_,
		_w2212_,
		_w2219_,
		_w2223_,
		_w2251_
	);
	LUT4 #(
		.INIT('h22b2)
	) name1789 (
		_w2231_,
		_w2235_,
		_w2242_,
		_w2246_,
		_w2252_
	);
	LUT3 #(
		.INIT('h07)
	) name1790 (
		_w2248_,
		_w2251_,
		_w2252_,
		_w2253_
	);
	LUT2 #(
		.INIT('h2)
	) name1791 (
		_w2196_,
		_w2200_,
		_w2254_
	);
	LUT4 #(
		.INIT('h20f2)
	) name1792 (
		_w2183_,
		_w2187_,
		_w2196_,
		_w2200_,
		_w2255_
	);
	LUT3 #(
		.INIT('h10)
	) name1793 (
		_w2165_,
		_w2177_,
		_w2255_,
		_w2256_
	);
	LUT3 #(
		.INIT('h01)
	) name1794 (
		_w1748_,
		_w2154_,
		_w2163_,
		_w2257_
	);
	LUT4 #(
		.INIT('h0023)
	) name1795 (
		_w1748_,
		_w2168_,
		_w2170_,
		_w2175_,
		_w2258_
	);
	LUT3 #(
		.INIT('h23)
	) name1796 (
		_w2165_,
		_w2257_,
		_w2258_,
		_w2259_
	);
	LUT2 #(
		.INIT('h4)
	) name1797 (
		_w2256_,
		_w2259_,
		_w2260_
	);
	LUT4 #(
		.INIT('h0d00)
	) name1798 (
		_w2204_,
		_w2253_,
		_w2256_,
		_w2259_,
		_w2261_
	);
	LUT4 #(
		.INIT('h2f00)
	) name1799 (
		_w2049_,
		_w2153_,
		_w2250_,
		_w2261_,
		_w2262_
	);
	LUT3 #(
		.INIT('he0)
	) name1800 (
		_w1748_,
		_w1982_,
		_w1987_,
		_w2263_
	);
	LUT2 #(
		.INIT('h1)
	) name1801 (
		_w1978_,
		_w2263_,
		_w2264_
	);
	LUT4 #(
		.INIT('h0001)
	) name1802 (
		_w1954_,
		_w1964_,
		_w1978_,
		_w2263_,
		_w2265_
	);
	LUT4 #(
		.INIT('h1000)
	) name1803 (
		_w1838_,
		_w1878_,
		_w1939_,
		_w2265_,
		_w2266_
	);
	LUT2 #(
		.INIT('h8)
	) name1804 (
		\P2_datao_reg[29]/NET0131 ,
		\si[29]_pad ,
		_w2267_
	);
	LUT4 #(
		.INIT('h135f)
	) name1805 (
		\P2_datao_reg[27]/NET0131 ,
		\P2_datao_reg[28]/NET0131 ,
		\si[27]_pad ,
		\si[28]_pad ,
		_w2268_
	);
	LUT4 #(
		.INIT('h3302)
	) name1806 (
		_w1799_,
		_w1803_,
		_w1868_,
		_w1909_,
		_w2269_
	);
	LUT2 #(
		.INIT('h2)
	) name1807 (
		_w2268_,
		_w2269_,
		_w2270_
	);
	LUT4 #(
		.INIT('h0455)
	) name1808 (
		_w1749_,
		_w1805_,
		_w1981_,
		_w2270_,
		_w2271_
	);
	LUT4 #(
		.INIT('h5659)
	) name1809 (
		\P2_datao_reg[29]/NET0131 ,
		\si[29]_pad ,
		_w547_,
		_w2271_,
		_w2272_
	);
	LUT2 #(
		.INIT('h1)
	) name1810 (
		_w1748_,
		_w2272_,
		_w2273_
	);
	LUT4 #(
		.INIT('h37f7)
	) name1811 (
		\P1_reg1_reg[29]/NET0131 ,
		_w478_,
		_w488_,
		_w1832_,
		_w2274_
	);
	LUT4 #(
		.INIT('hf3f5)
	) name1812 (
		\P1_reg0_reg[29]/NET0131 ,
		\P1_reg2_reg[29]/NET0131 ,
		_w478_,
		_w488_,
		_w2275_
	);
	LUT2 #(
		.INIT('h8)
	) name1813 (
		_w2274_,
		_w2275_,
		_w2276_
	);
	LUT2 #(
		.INIT('h7)
	) name1814 (
		_w2274_,
		_w2275_,
		_w2277_
	);
	LUT3 #(
		.INIT('h10)
	) name1815 (
		_w1748_,
		_w2272_,
		_w2276_,
		_w2278_
	);
	LUT3 #(
		.INIT('h0e)
	) name1816 (
		_w1748_,
		_w2272_,
		_w2276_,
		_w2279_
	);
	LUT3 #(
		.INIT('he1)
	) name1817 (
		_w1748_,
		_w2272_,
		_w2276_,
		_w2280_
	);
	LUT4 #(
		.INIT('h45ba)
	) name1818 (
		_w2000_,
		_w2262_,
		_w2266_,
		_w2280_,
		_w2281_
	);
	LUT4 #(
		.INIT('ha666)
	) name1819 (
		\P1_IR_reg[22]/NET0131 ,
		\P1_IR_reg[31]/NET0131 ,
		_w480_,
		_w482_,
		_w2282_
	);
	LUT4 #(
		.INIT('ha600)
	) name1820 (
		\P1_IR_reg[23]/NET0131 ,
		\P1_IR_reg[31]/NET0131 ,
		_w1722_,
		_w2282_,
		_w2283_
	);
	LUT4 #(
		.INIT('h0059)
	) name1821 (
		\P1_IR_reg[23]/NET0131 ,
		\P1_IR_reg[31]/NET0131 ,
		_w1722_,
		_w2282_,
		_w2284_
	);
	LUT4 #(
		.INIT('h59a6)
	) name1822 (
		\P1_IR_reg[23]/NET0131 ,
		\P1_IR_reg[31]/NET0131 ,
		_w1722_,
		_w2282_,
		_w2285_
	);
	LUT2 #(
		.INIT('h2)
	) name1823 (
		\P1_IR_reg[31]/NET0131 ,
		_w472_,
		_w2286_
	);
	LUT4 #(
		.INIT('h00d5)
	) name1824 (
		\P1_IR_reg[31]/NET0131 ,
		_w467_,
		_w471_,
		_w2286_,
		_w2287_
	);
	LUT2 #(
		.INIT('h9)
	) name1825 (
		\P1_IR_reg[21]/NET0131 ,
		_w2287_,
		_w2288_
	);
	LUT3 #(
		.INIT('h84)
	) name1826 (
		\P1_IR_reg[21]/NET0131 ,
		_w2282_,
		_w2287_,
		_w2289_
	);
	LUT4 #(
		.INIT('h2aaa)
	) name1827 (
		\P1_IR_reg[31]/NET0131 ,
		_w468_,
		_w480_,
		_w1724_,
		_w2290_
	);
	LUT2 #(
		.INIT('h9)
	) name1828 (
		\P1_IR_reg[20]/NET0131 ,
		_w2290_,
		_w2291_
	);
	LUT4 #(
		.INIT('h0c04)
	) name1829 (
		_w1723_,
		_w2285_,
		_w2289_,
		_w2291_,
		_w2292_
	);
	LUT4 #(
		.INIT('h2e00)
	) name1830 (
		\P1_reg2_reg[29]/NET0131 ,
		_w1741_,
		_w2281_,
		_w2292_,
		_w2293_
	);
	LUT4 #(
		.INIT('h0777)
	) name1831 (
		_w2004_,
		_w2008_,
		_w2016_,
		_w2020_,
		_w2294_
	);
	LUT4 #(
		.INIT('h1000)
	) name1832 (
		_w2024_,
		_w2028_,
		_w2030_,
		_w2033_,
		_w2295_
	);
	LUT3 #(
		.INIT('h15)
	) name1833 (
		_w2040_,
		_w2041_,
		_w2043_,
		_w2296_
	);
	LUT4 #(
		.INIT('h0eee)
	) name1834 (
		_w2024_,
		_w2028_,
		_w2030_,
		_w2033_,
		_w2297_
	);
	LUT3 #(
		.INIT('h54)
	) name1835 (
		_w2295_,
		_w2296_,
		_w2297_,
		_w2298_
	);
	LUT2 #(
		.INIT('h1)
	) name1836 (
		_w2004_,
		_w2008_,
		_w2299_
	);
	LUT4 #(
		.INIT('hfee0)
	) name1837 (
		_w2004_,
		_w2008_,
		_w2016_,
		_w2020_,
		_w2300_
	);
	LUT3 #(
		.INIT('h70)
	) name1838 (
		_w2294_,
		_w2298_,
		_w2300_,
		_w2301_
	);
	LUT3 #(
		.INIT('h70)
	) name1839 (
		_w2051_,
		_w2052_,
		_w2057_,
		_w2302_
	);
	LUT3 #(
		.INIT('h70)
	) name1840 (
		_w489_,
		_w491_,
		_w2071_,
		_w2303_
	);
	LUT2 #(
		.INIT('h1)
	) name1841 (
		_w2302_,
		_w2303_,
		_w2304_
	);
	LUT3 #(
		.INIT('h08)
	) name1842 (
		_w2084_,
		_w2085_,
		_w2089_,
		_w2305_
	);
	LUT3 #(
		.INIT('h70)
	) name1843 (
		_w2059_,
		_w2060_,
		_w2065_,
		_w2306_
	);
	LUT4 #(
		.INIT('h00b2)
	) name1844 (
		_w2077_,
		_w2081_,
		_w2305_,
		_w2306_,
		_w2307_
	);
	LUT3 #(
		.INIT('h08)
	) name1845 (
		_w2059_,
		_w2060_,
		_w2065_,
		_w2308_
	);
	LUT3 #(
		.INIT('h08)
	) name1846 (
		_w489_,
		_w491_,
		_w2071_,
		_w2309_
	);
	LUT2 #(
		.INIT('h1)
	) name1847 (
		_w2308_,
		_w2309_,
		_w2310_
	);
	LUT3 #(
		.INIT('h40)
	) name1848 (
		_w2124_,
		_w2125_,
		_w2127_,
		_w2311_
	);
	LUT3 #(
		.INIT('h08)
	) name1849 (
		_w2051_,
		_w2052_,
		_w2057_,
		_w2312_
	);
	LUT3 #(
		.INIT('h40)
	) name1850 (
		_w2134_,
		_w2135_,
		_w2137_,
		_w2313_
	);
	LUT2 #(
		.INIT('h1)
	) name1851 (
		_w2312_,
		_w2313_,
		_w2314_
	);
	LUT3 #(
		.INIT('h01)
	) name1852 (
		_w2311_,
		_w2312_,
		_w2313_,
		_w2315_
	);
	LUT4 #(
		.INIT('h7500)
	) name1853 (
		_w2304_,
		_w2307_,
		_w2310_,
		_w2315_,
		_w2316_
	);
	LUT3 #(
		.INIT('h2a)
	) name1854 (
		_w2124_,
		_w2125_,
		_w2127_,
		_w2317_
	);
	LUT3 #(
		.INIT('h2a)
	) name1855 (
		_w2134_,
		_w2135_,
		_w2137_,
		_w2318_
	);
	LUT2 #(
		.INIT('h1)
	) name1856 (
		_w2317_,
		_w2318_,
		_w2319_
	);
	LUT3 #(
		.INIT('h54)
	) name1857 (
		_w2311_,
		_w2317_,
		_w2318_,
		_w2320_
	);
	LUT4 #(
		.INIT('h1000)
	) name1858 (
		_w2099_,
		_w2103_,
		_w2105_,
		_w2107_,
		_w2321_
	);
	LUT3 #(
		.INIT('h80)
	) name1859 (
		_w2114_,
		_w2116_,
		_w2117_,
		_w2322_
	);
	LUT2 #(
		.INIT('h1)
	) name1860 (
		_w2321_,
		_w2322_,
		_w2323_
	);
	LUT4 #(
		.INIT('h0eee)
	) name1861 (
		_w2099_,
		_w2103_,
		_w2105_,
		_w2107_,
		_w2324_
	);
	LUT3 #(
		.INIT('h15)
	) name1862 (
		_w2114_,
		_w2116_,
		_w2117_,
		_w2325_
	);
	LUT3 #(
		.INIT('h54)
	) name1863 (
		_w2321_,
		_w2324_,
		_w2325_,
		_w2326_
	);
	LUT4 #(
		.INIT('h001f)
	) name1864 (
		_w2316_,
		_w2320_,
		_w2323_,
		_w2326_,
		_w2327_
	);
	LUT3 #(
		.INIT('h80)
	) name1865 (
		_w2040_,
		_w2041_,
		_w2043_,
		_w2328_
	);
	LUT2 #(
		.INIT('h1)
	) name1866 (
		_w2295_,
		_w2328_,
		_w2329_
	);
	LUT2 #(
		.INIT('h8)
	) name1867 (
		_w2294_,
		_w2329_,
		_w2330_
	);
	LUT4 #(
		.INIT('h0777)
	) name1868 (
		_w2231_,
		_w2235_,
		_w2242_,
		_w2246_,
		_w2331_
	);
	LUT4 #(
		.INIT('heee0)
	) name1869 (
		_w2208_,
		_w2212_,
		_w2219_,
		_w2223_,
		_w2332_
	);
	LUT4 #(
		.INIT('h1117)
	) name1870 (
		_w2208_,
		_w2212_,
		_w2219_,
		_w2223_,
		_w2333_
	);
	LUT2 #(
		.INIT('h1)
	) name1871 (
		_w2242_,
		_w2246_,
		_w2334_
	);
	LUT4 #(
		.INIT('h1117)
	) name1872 (
		_w2231_,
		_w2235_,
		_w2242_,
		_w2246_,
		_w2335_
	);
	LUT3 #(
		.INIT('h07)
	) name1873 (
		_w2331_,
		_w2333_,
		_w2335_,
		_w2336_
	);
	LUT3 #(
		.INIT('h10)
	) name1874 (
		_w1748_,
		_w2154_,
		_w2163_,
		_w2337_
	);
	LUT4 #(
		.INIT('h2300)
	) name1875 (
		_w1748_,
		_w2168_,
		_w2170_,
		_w2175_,
		_w2338_
	);
	LUT2 #(
		.INIT('h8)
	) name1876 (
		_w2196_,
		_w2200_,
		_w2339_
	);
	LUT2 #(
		.INIT('h1)
	) name1877 (
		_w2196_,
		_w2200_,
		_w2340_
	);
	LUT4 #(
		.INIT('heee0)
	) name1878 (
		_w2183_,
		_w2187_,
		_w2196_,
		_w2200_,
		_w2341_
	);
	LUT4 #(
		.INIT('h011f)
	) name1879 (
		_w2183_,
		_w2187_,
		_w2196_,
		_w2200_,
		_w2342_
	);
	LUT3 #(
		.INIT('h10)
	) name1880 (
		_w2337_,
		_w2338_,
		_w2342_,
		_w2343_
	);
	LUT3 #(
		.INIT('h0e)
	) name1881 (
		_w1748_,
		_w2154_,
		_w2163_,
		_w2344_
	);
	LUT4 #(
		.INIT('h00dc)
	) name1882 (
		_w1748_,
		_w2168_,
		_w2170_,
		_w2175_,
		_w2345_
	);
	LUT3 #(
		.INIT('h54)
	) name1883 (
		_w2337_,
		_w2344_,
		_w2345_,
		_w2346_
	);
	LUT2 #(
		.INIT('h1)
	) name1884 (
		_w2343_,
		_w2346_,
		_w2347_
	);
	LUT3 #(
		.INIT('h02)
	) name1885 (
		_w2336_,
		_w2343_,
		_w2346_,
		_w2348_
	);
	LUT4 #(
		.INIT('h8a00)
	) name1886 (
		_w2301_,
		_w2327_,
		_w2330_,
		_w2348_,
		_w2349_
	);
	LUT4 #(
		.INIT('h0777)
	) name1887 (
		_w2183_,
		_w2187_,
		_w2196_,
		_w2200_,
		_w2350_
	);
	LUT3 #(
		.INIT('h10)
	) name1888 (
		_w2337_,
		_w2338_,
		_w2350_,
		_w2351_
	);
	LUT4 #(
		.INIT('h0777)
	) name1889 (
		_w2208_,
		_w2212_,
		_w2219_,
		_w2223_,
		_w2352_
	);
	LUT2 #(
		.INIT('h8)
	) name1890 (
		_w2331_,
		_w2352_,
		_w2353_
	);
	LUT4 #(
		.INIT('h0507)
	) name1891 (
		_w2331_,
		_w2333_,
		_w2335_,
		_w2352_,
		_w2354_
	);
	LUT4 #(
		.INIT('h1101)
	) name1892 (
		_w2343_,
		_w2346_,
		_w2351_,
		_w2354_,
		_w2355_
	);
	LUT4 #(
		.INIT('h5400)
	) name1893 (
		_w1748_,
		_w1907_,
		_w1929_,
		_w1936_,
		_w2356_
	);
	LUT3 #(
		.INIT('h10)
	) name1894 (
		_w1748_,
		_w1815_,
		_w1836_,
		_w2357_
	);
	LUT4 #(
		.INIT('h00ef)
	) name1895 (
		_w1748_,
		_w1815_,
		_w1836_,
		_w2356_,
		_w2358_
	);
	LUT4 #(
		.INIT('h5400)
	) name1896 (
		_w1748_,
		_w1839_,
		_w1870_,
		_w1876_,
		_w2359_
	);
	LUT3 #(
		.INIT('h10)
	) name1897 (
		_w1748_,
		_w1899_,
		_w1904_,
		_w2360_
	);
	LUT4 #(
		.INIT('h00ef)
	) name1898 (
		_w1748_,
		_w1899_,
		_w1904_,
		_w2359_,
		_w2361_
	);
	LUT2 #(
		.INIT('h8)
	) name1899 (
		_w2358_,
		_w2361_,
		_w2362_
	);
	LUT3 #(
		.INIT('h10)
	) name1900 (
		_w1748_,
		_w1982_,
		_w1987_,
		_w2363_
	);
	LUT4 #(
		.INIT('h5400)
	) name1901 (
		_w1748_,
		_w1966_,
		_w1970_,
		_w1975_,
		_w2364_
	);
	LUT2 #(
		.INIT('h1)
	) name1902 (
		_w2363_,
		_w2364_,
		_w2365_
	);
	LUT3 #(
		.INIT('h10)
	) name1903 (
		_w1748_,
		_w1957_,
		_w1962_,
		_w2366_
	);
	LUT4 #(
		.INIT('h5400)
	) name1904 (
		_w1748_,
		_w1941_,
		_w1947_,
		_w1952_,
		_w2367_
	);
	LUT2 #(
		.INIT('h1)
	) name1905 (
		_w2366_,
		_w2367_,
		_w2368_
	);
	LUT4 #(
		.INIT('h0001)
	) name1906 (
		_w2363_,
		_w2364_,
		_w2366_,
		_w2367_,
		_w2369_
	);
	LUT3 #(
		.INIT('h80)
	) name1907 (
		_w2358_,
		_w2361_,
		_w2369_,
		_w2370_
	);
	LUT2 #(
		.INIT('h4)
	) name1908 (
		_w2355_,
		_w2370_,
		_w2371_
	);
	LUT4 #(
		.INIT('h00ab)
	) name1909 (
		_w1748_,
		_w1966_,
		_w1970_,
		_w1975_,
		_w2372_
	);
	LUT3 #(
		.INIT('h0e)
	) name1910 (
		_w1748_,
		_w1982_,
		_w1987_,
		_w2373_
	);
	LUT3 #(
		.INIT('h54)
	) name1911 (
		_w2364_,
		_w2372_,
		_w2373_,
		_w2374_
	);
	LUT4 #(
		.INIT('h00ab)
	) name1912 (
		_w1748_,
		_w1941_,
		_w1947_,
		_w1952_,
		_w2375_
	);
	LUT3 #(
		.INIT('h0e)
	) name1913 (
		_w1748_,
		_w1957_,
		_w1962_,
		_w2376_
	);
	LUT3 #(
		.INIT('h23)
	) name1914 (
		_w2367_,
		_w2375_,
		_w2376_,
		_w2377_
	);
	LUT3 #(
		.INIT('h70)
	) name1915 (
		_w2368_,
		_w2374_,
		_w2377_,
		_w2378_
	);
	LUT4 #(
		.INIT('h00ab)
	) name1916 (
		_w1748_,
		_w1839_,
		_w1870_,
		_w1876_,
		_w2379_
	);
	LUT4 #(
		.INIT('h00f1)
	) name1917 (
		_w1748_,
		_w1899_,
		_w1904_,
		_w2379_,
		_w2380_
	);
	LUT4 #(
		.INIT('hef0e)
	) name1918 (
		_w1748_,
		_w1899_,
		_w1904_,
		_w2379_,
		_w2381_
	);
	LUT3 #(
		.INIT('h0e)
	) name1919 (
		_w1748_,
		_w1815_,
		_w1836_,
		_w2382_
	);
	LUT4 #(
		.INIT('h00ab)
	) name1920 (
		_w1748_,
		_w1907_,
		_w1929_,
		_w1936_,
		_w2383_
	);
	LUT4 #(
		.INIT('h10f1)
	) name1921 (
		_w1748_,
		_w1815_,
		_w1836_,
		_w2383_,
		_w2384_
	);
	LUT3 #(
		.INIT('h70)
	) name1922 (
		_w2358_,
		_w2381_,
		_w2384_,
		_w2385_
	);
	LUT3 #(
		.INIT('hd0)
	) name1923 (
		_w2362_,
		_w2378_,
		_w2385_,
		_w2386_
	);
	LUT4 #(
		.INIT('h9a55)
	) name1924 (
		_w2280_,
		_w2349_,
		_w2371_,
		_w2386_,
		_w2387_
	);
	LUT4 #(
		.INIT('h3032)
	) name1925 (
		_w1723_,
		_w2283_,
		_w2289_,
		_w2291_,
		_w2388_
	);
	LUT4 #(
		.INIT('he200)
	) name1926 (
		\P1_reg2_reg[29]/NET0131 ,
		_w1741_,
		_w2387_,
		_w2388_,
		_w2389_
	);
	LUT2 #(
		.INIT('h2)
	) name1927 (
		_w1747_,
		_w1836_,
		_w2390_
	);
	LUT4 #(
		.INIT('h0777)
	) name1928 (
		_w2173_,
		_w2174_,
		_w2198_,
		_w2199_,
		_w2391_
	);
	LUT2 #(
		.INIT('h4)
	) name1929 (
		_w2163_,
		_w2391_,
		_w2392_
	);
	LUT4 #(
		.INIT('h0777)
	) name1930 (
		_w1984_,
		_w1986_,
		_w2184_,
		_w2186_,
		_w2393_
	);
	LUT4 #(
		.INIT('h1000)
	) name1931 (
		_w2163_,
		_w2235_,
		_w2391_,
		_w2393_,
		_w2394_
	);
	LUT4 #(
		.INIT('h1fdf)
	) name1932 (
		\P1_reg2_reg[31]/NET0131 ,
		_w478_,
		_w488_,
		_w1832_,
		_w2395_
	);
	LUT4 #(
		.INIT('hff35)
	) name1933 (
		\P1_reg0_reg[31]/NET0131 ,
		\P1_reg1_reg[31]/NET0131 ,
		_w478_,
		_w488_,
		_w2396_
	);
	LUT2 #(
		.INIT('h8)
	) name1934 (
		_w2395_,
		_w2396_,
		_w2397_
	);
	LUT2 #(
		.INIT('h7)
	) name1935 (
		_w2395_,
		_w2396_,
		_w2398_
	);
	LUT4 #(
		.INIT('h0777)
	) name1936 (
		_w2084_,
		_w2085_,
		_w2395_,
		_w2396_,
		_w2399_
	);
	LUT4 #(
		.INIT('h0100)
	) name1937 (
		_w492_,
		_w2061_,
		_w2077_,
		_w2399_,
		_w2400_
	);
	LUT4 #(
		.INIT('h0777)
	) name1938 (
		_w2041_,
		_w2043_,
		_w2105_,
		_w2107_,
		_w2401_
	);
	LUT4 #(
		.INIT('h0777)
	) name1939 (
		_w2116_,
		_w2117_,
		_w2125_,
		_w2127_,
		_w2402_
	);
	LUT2 #(
		.INIT('h8)
	) name1940 (
		_w2401_,
		_w2402_,
		_w2403_
	);
	LUT4 #(
		.INIT('h1000)
	) name1941 (
		_w2053_,
		_w2138_,
		_w2400_,
		_w2403_,
		_w2404_
	);
	LUT4 #(
		.INIT('h0777)
	) name1942 (
		_w2006_,
		_w2007_,
		_w2030_,
		_w2033_,
		_w2405_
	);
	LUT2 #(
		.INIT('h4)
	) name1943 (
		_w2020_,
		_w2405_,
		_w2406_
	);
	LUT4 #(
		.INIT('h0777)
	) name1944 (
		_w2210_,
		_w2211_,
		_w2221_,
		_w2222_,
		_w2407_
	);
	LUT4 #(
		.INIT('h1000)
	) name1945 (
		_w2020_,
		_w2246_,
		_w2405_,
		_w2407_,
		_w2408_
	);
	LUT2 #(
		.INIT('h8)
	) name1946 (
		_w2404_,
		_w2408_,
		_w2409_
	);
	LUT3 #(
		.INIT('h80)
	) name1947 (
		_w2394_,
		_w2404_,
		_w2408_,
		_w2410_
	);
	LUT4 #(
		.INIT('h0777)
	) name1948 (
		_w1949_,
		_w1951_,
		_w1960_,
		_w1961_,
		_w2411_
	);
	LUT3 #(
		.INIT('h10)
	) name1949 (
		_w1876_,
		_w1904_,
		_w2411_,
		_w2412_
	);
	LUT2 #(
		.INIT('h1)
	) name1950 (
		_w1936_,
		_w1975_,
		_w2413_
	);
	LUT2 #(
		.INIT('h8)
	) name1951 (
		_w2412_,
		_w2413_,
		_w2414_
	);
	LUT3 #(
		.INIT('h40)
	) name1952 (
		_w1836_,
		_w2412_,
		_w2413_,
		_w2415_
	);
	LUT4 #(
		.INIT('h8000)
	) name1953 (
		_w2394_,
		_w2404_,
		_w2408_,
		_w2415_,
		_w2416_
	);
	LUT4 #(
		.INIT('h1fdf)
	) name1954 (
		\P1_reg2_reg[30]/NET0131 ,
		_w478_,
		_w488_,
		_w1832_,
		_w2417_
	);
	LUT4 #(
		.INIT('hff35)
	) name1955 (
		\P1_reg0_reg[30]/NET0131 ,
		\P1_reg1_reg[30]/NET0131 ,
		_w478_,
		_w488_,
		_w2418_
	);
	LUT2 #(
		.INIT('h8)
	) name1956 (
		_w2417_,
		_w2418_,
		_w2419_
	);
	LUT2 #(
		.INIT('h7)
	) name1957 (
		_w2417_,
		_w2418_,
		_w2420_
	);
	LUT3 #(
		.INIT('hf8)
	) name1958 (
		\P1_B_reg/NET0131 ,
		_w1744_,
		_w1747_,
		_w2421_
	);
	LUT4 #(
		.INIT('h1023)
	) name1959 (
		_w2276_,
		_w2421_,
		_w2416_,
		_w2419_,
		_w2422_
	);
	LUT4 #(
		.INIT('h111d)
	) name1960 (
		\P1_reg2_reg[29]/NET0131 ,
		_w1741_,
		_w2390_,
		_w2422_,
		_w2423_
	);
	LUT4 #(
		.INIT('h0800)
	) name1961 (
		_w1723_,
		_w2282_,
		_w2288_,
		_w2291_,
		_w2424_
	);
	LUT3 #(
		.INIT('h21)
	) name1962 (
		\P1_IR_reg[21]/NET0131 ,
		_w2282_,
		_w2287_,
		_w2425_
	);
	LUT2 #(
		.INIT('h4)
	) name1963 (
		_w1723_,
		_w2425_,
		_w2426_
	);
	LUT3 #(
		.INIT('h10)
	) name1964 (
		_w1748_,
		_w2272_,
		_w2426_,
		_w2427_
	);
	LUT3 #(
		.INIT('h80)
	) name1965 (
		_w2065_,
		_w2081_,
		_w2089_,
		_w2428_
	);
	LUT4 #(
		.INIT('h8000)
	) name1966 (
		_w2065_,
		_w2071_,
		_w2081_,
		_w2089_,
		_w2429_
	);
	LUT2 #(
		.INIT('h8)
	) name1967 (
		_w2124_,
		_w2134_,
		_w2430_
	);
	LUT4 #(
		.INIT('h2000)
	) name1968 (
		_w2057_,
		_w2114_,
		_w2429_,
		_w2430_,
		_w2431_
	);
	LUT2 #(
		.INIT('h1)
	) name1969 (
		_w2004_,
		_w2016_,
		_w2432_
	);
	LUT3 #(
		.INIT('h0e)
	) name1970 (
		_w2024_,
		_w2028_,
		_w2040_,
		_w2433_
	);
	LUT3 #(
		.INIT('h10)
	) name1971 (
		_w2104_,
		_w2219_,
		_w2433_,
		_w2434_
	);
	LUT4 #(
		.INIT('h0001)
	) name1972 (
		_w2183_,
		_w2208_,
		_w2231_,
		_w2242_,
		_w2435_
	);
	LUT4 #(
		.INIT('h8000)
	) name1973 (
		_w2431_,
		_w2432_,
		_w2434_,
		_w2435_,
		_w2436_
	);
	LUT3 #(
		.INIT('h0e)
	) name1974 (
		_w1748_,
		_w2154_,
		_w2196_,
		_w2437_
	);
	LUT2 #(
		.INIT('h4)
	) name1975 (
		_w2171_,
		_w2437_,
		_w2438_
	);
	LUT4 #(
		.INIT('habaa)
	) name1976 (
		_w1748_,
		_w1966_,
		_w1970_,
		_w1982_,
		_w2439_
	);
	LUT3 #(
		.INIT('h80)
	) name1977 (
		_w2436_,
		_w2438_,
		_w2439_,
		_w2440_
	);
	LUT4 #(
		.INIT('habaa)
	) name1978 (
		_w1748_,
		_w1839_,
		_w1870_,
		_w1957_,
		_w2441_
	);
	LUT2 #(
		.INIT('h4)
	) name1979 (
		_w1948_,
		_w2441_,
		_w2442_
	);
	LUT4 #(
		.INIT('h8000)
	) name1980 (
		_w2436_,
		_w2438_,
		_w2439_,
		_w2442_,
		_w2443_
	);
	LUT4 #(
		.INIT('heaaa)
	) name1981 (
		_w1748_,
		_w1815_,
		_w1899_,
		_w1930_,
		_w2444_
	);
	LUT2 #(
		.INIT('h8)
	) name1982 (
		_w2443_,
		_w2444_,
		_w2445_
	);
	LUT2 #(
		.INIT('h2)
	) name1983 (
		_w2284_,
		_w2288_,
		_w2446_
	);
	LUT3 #(
		.INIT('h20)
	) name1984 (
		_w2284_,
		_w2288_,
		_w2291_,
		_w2447_
	);
	LUT4 #(
		.INIT('h9500)
	) name1985 (
		_w2273_,
		_w2443_,
		_w2444_,
		_w2447_,
		_w2448_
	);
	LUT4 #(
		.INIT('h2814)
	) name1986 (
		\P1_IR_reg[20]/NET0131 ,
		\P1_IR_reg[21]/NET0131 ,
		_w2287_,
		_w2290_,
		_w2449_
	);
	LUT2 #(
		.INIT('h2)
	) name1987 (
		_w2283_,
		_w2449_,
		_w2450_
	);
	LUT4 #(
		.INIT('h1428)
	) name1988 (
		\P1_IR_reg[20]/NET0131 ,
		\P1_IR_reg[21]/NET0131 ,
		_w2287_,
		_w2290_,
		_w2451_
	);
	LUT2 #(
		.INIT('h2)
	) name1989 (
		_w2284_,
		_w2451_,
		_w2452_
	);
	LUT4 #(
		.INIT('ha2a0)
	) name1990 (
		\P1_reg2_reg[29]/NET0131 ,
		_w1741_,
		_w2450_,
		_w2452_,
		_w2453_
	);
	LUT3 #(
		.INIT('h02)
	) name1991 (
		_w2284_,
		_w2288_,
		_w2291_,
		_w2454_
	);
	LUT4 #(
		.INIT('h0008)
	) name1992 (
		_w1832_,
		_w2284_,
		_w2288_,
		_w2291_,
		_w2455_
	);
	LUT2 #(
		.INIT('h1)
	) name1993 (
		_w2453_,
		_w2455_,
		_w2456_
	);
	LUT4 #(
		.INIT('h5700)
	) name1994 (
		_w1741_,
		_w2427_,
		_w2448_,
		_w2456_,
		_w2457_
	);
	LUT3 #(
		.INIT('hb0)
	) name1995 (
		_w2423_,
		_w2424_,
		_w2457_,
		_w2458_
	);
	LUT4 #(
		.INIT('ha8aa)
	) name1996 (
		_w1731_,
		_w2293_,
		_w2389_,
		_w2458_,
		_w2459_
	);
	LUT3 #(
		.INIT('h40)
	) name1997 (
		_w1723_,
		_w1727_,
		_w1730_,
		_w2460_
	);
	LUT4 #(
		.INIT('h2000)
	) name1998 (
		\P1_reg2_reg[29]/NET0131 ,
		_w1723_,
		_w1727_,
		_w1730_,
		_w2461_
	);
	LUT4 #(
		.INIT('h5090)
	) name1999 (
		\P1_IR_reg[23]/NET0131 ,
		\P1_IR_reg[31]/NET0131 ,
		\P1_state_reg[0]/NET0131 ,
		_w1722_,
		_w2462_
	);
	LUT2 #(
		.INIT('h2)
	) name2000 (
		\P1_reg2_reg[29]/NET0131 ,
		_w2462_,
		_w2463_
	);
	LUT4 #(
		.INIT('hffa8)
	) name2001 (
		\P1_state_reg[0]/NET0131 ,
		_w2459_,
		_w2461_,
		_w2463_,
		_w2464_
	);
	LUT4 #(
		.INIT('hd070)
	) name2002 (
		\P1_state_reg[0]/NET0131 ,
		\P2_IR_reg[23]/NET0131 ,
		\P2_reg1_reg[29]/NET0131 ,
		_w1188_,
		_w2465_
	);
	LUT4 #(
		.INIT('h2000)
	) name2003 (
		\P2_reg1_reg[29]/NET0131 ,
		_w1189_,
		_w1352_,
		_w1356_,
		_w2466_
	);
	LUT4 #(
		.INIT('h35c5)
	) name2004 (
		\P2_reg1_reg[29]/NET0131 ,
		_w1264_,
		_w1516_,
		_w1678_,
		_w2467_
	);
	LUT4 #(
		.INIT('h08c8)
	) name2005 (
		\P2_reg1_reg[29]/NET0131 ,
		_w1191_,
		_w1507_,
		_w1682_,
		_w2468_
	);
	LUT4 #(
		.INIT('hf100)
	) name2006 (
		_w1361_,
		_w1363_,
		_w1368_,
		_w1442_,
		_w2469_
	);
	LUT3 #(
		.INIT('ha2)
	) name2007 (
		\P2_reg1_reg[29]/NET0131 ,
		_w1684_,
		_w2469_,
		_w2470_
	);
	LUT4 #(
		.INIT('h0e00)
	) name2008 (
		_w1361_,
		_w1363_,
		_w1368_,
		_w1442_,
		_w2471_
	);
	LUT4 #(
		.INIT('h0e0f)
	) name2009 (
		_w546_,
		_w1107_,
		_w2470_,
		_w2471_,
		_w2472_
	);
	LUT2 #(
		.INIT('h4)
	) name2010 (
		_w2468_,
		_w2472_,
		_w2473_
	);
	LUT3 #(
		.INIT('he0)
	) name2011 (
		_w1506_,
		_w2467_,
		_w2473_,
		_w2474_
	);
	LUT4 #(
		.INIT('hc535)
	) name2012 (
		\P2_reg1_reg[29]/NET0131 ,
		_w1264_,
		_w1516_,
		_w1712_,
		_w2475_
	);
	LUT4 #(
		.INIT('h35c5)
	) name2013 (
		\P2_reg1_reg[29]/NET0131 ,
		_w1264_,
		_w1507_,
		_w1678_,
		_w2476_
	);
	LUT4 #(
		.INIT('hfc54)
	) name2014 (
		_w1530_,
		_w1575_,
		_w2475_,
		_w2476_,
		_w2477_
	);
	LUT4 #(
		.INIT('h3111)
	) name2015 (
		_w1359_,
		_w2466_,
		_w2474_,
		_w2477_,
		_w2478_
	);
	LUT3 #(
		.INIT('hce)
	) name2016 (
		\P1_state_reg[0]/NET0131 ,
		_w2465_,
		_w2478_,
		_w2479_
	);
	LUT4 #(
		.INIT('hd070)
	) name2017 (
		\P1_state_reg[0]/NET0131 ,
		\P2_IR_reg[23]/NET0131 ,
		\P2_reg2_reg[25]/NET0131 ,
		_w1188_,
		_w2480_
	);
	LUT4 #(
		.INIT('h2000)
	) name2018 (
		\P2_reg2_reg[25]/NET0131 ,
		_w1189_,
		_w1352_,
		_w1356_,
		_w2481_
	);
	LUT4 #(
		.INIT('ha8aa)
	) name2019 (
		\P2_reg2_reg[25]/NET0131 ,
		_w1361_,
		_w1363_,
		_w1368_,
		_w2482_
	);
	LUT4 #(
		.INIT('h0800)
	) name2020 (
		_w1657_,
		_w1658_,
		_w1662_,
		_w1663_,
		_w2483_
	);
	LUT4 #(
		.INIT('h08aa)
	) name2021 (
		_w1657_,
		_w1658_,
		_w1660_,
		_w1665_,
		_w2484_
	);
	LUT4 #(
		.INIT('hccc4)
	) name2022 (
		_w1667_,
		_w1670_,
		_w2484_,
		_w2483_,
		_w2485_
	);
	LUT4 #(
		.INIT('h8848)
	) name2023 (
		_w1271_,
		_w1507_,
		_w1674_,
		_w2485_,
		_w2486_
	);
	LUT3 #(
		.INIT('h54)
	) name2024 (
		_w1506_,
		_w2482_,
		_w2486_,
		_w2487_
	);
	LUT4 #(
		.INIT('haa02)
	) name2025 (
		\P2_reg2_reg[25]/NET0131 ,
		_w1361_,
		_w1363_,
		_w1368_,
		_w2488_
	);
	LUT4 #(
		.INIT('h1000)
	) name2026 (
		_w1035_,
		_w1069_,
		_w1423_,
		_w1429_,
		_w2489_
	);
	LUT4 #(
		.INIT('h002f)
	) name2027 (
		_w519_,
		_w1042_,
		_w1046_,
		_w1435_,
		_w2490_
	);
	LUT4 #(
		.INIT('h007b)
	) name2028 (
		_w1069_,
		_w1435_,
		_w1626_,
		_w2490_,
		_w2491_
	);
	LUT4 #(
		.INIT('h08c8)
	) name2029 (
		\P2_reg2_reg[25]/NET0131 ,
		_w1191_,
		_w1516_,
		_w2491_,
		_w2492_
	);
	LUT2 #(
		.INIT('h4)
	) name2030 (
		_w1030_,
		_w1233_,
		_w2493_
	);
	LUT4 #(
		.INIT('h0057)
	) name2031 (
		\P2_reg2_reg[25]/NET0131 ,
		_w1441_,
		_w1523_,
		_w2493_,
		_w2494_
	);
	LUT4 #(
		.INIT('hef00)
	) name2032 (
		_w546_,
		_w1026_,
		_w1522_,
		_w2494_,
		_w2495_
	);
	LUT2 #(
		.INIT('h4)
	) name2033 (
		_w2492_,
		_w2495_,
		_w2496_
	);
	LUT4 #(
		.INIT('h08aa)
	) name2034 (
		_w1691_,
		_w1692_,
		_w1694_,
		_w1700_,
		_w2497_
	);
	LUT4 #(
		.INIT('h0070)
	) name2035 (
		_w1693_,
		_w1698_,
		_w1702_,
		_w2497_,
		_w2498_
	);
	LUT4 #(
		.INIT('h5a9a)
	) name2036 (
		_w1271_,
		_w1705_,
		_w1710_,
		_w2498_,
		_w2499_
	);
	LUT4 #(
		.INIT('h020e)
	) name2037 (
		\P2_reg2_reg[25]/NET0131 ,
		_w1507_,
		_w1575_,
		_w2499_,
		_w2500_
	);
	LUT4 #(
		.INIT('h8848)
	) name2038 (
		_w1271_,
		_w1516_,
		_w1674_,
		_w2485_,
		_w2501_
	);
	LUT3 #(
		.INIT('ha8)
	) name2039 (
		_w1530_,
		_w2488_,
		_w2501_,
		_w2502_
	);
	LUT4 #(
		.INIT('h0100)
	) name2040 (
		_w2487_,
		_w2500_,
		_w2502_,
		_w2496_,
		_w2503_
	);
	LUT4 #(
		.INIT('ha0a8)
	) name2041 (
		\P1_state_reg[0]/NET0131 ,
		_w1359_,
		_w2481_,
		_w2503_,
		_w2504_
	);
	LUT2 #(
		.INIT('he)
	) name2042 (
		_w2480_,
		_w2504_,
		_w2505_
	);
	LUT4 #(
		.INIT('hd070)
	) name2043 (
		\P1_state_reg[0]/NET0131 ,
		\P2_IR_reg[23]/NET0131 ,
		\P2_reg2_reg[29]/NET0131 ,
		_w1188_,
		_w2506_
	);
	LUT4 #(
		.INIT('h2000)
	) name2044 (
		\P2_reg2_reg[29]/NET0131 ,
		_w1189_,
		_w1352_,
		_w1356_,
		_w2507_
	);
	LUT4 #(
		.INIT('h35c5)
	) name2045 (
		\P2_reg2_reg[29]/NET0131 ,
		_w1264_,
		_w1507_,
		_w1678_,
		_w2508_
	);
	LUT4 #(
		.INIT('h08c8)
	) name2046 (
		\P2_reg2_reg[29]/NET0131 ,
		_w1191_,
		_w1516_,
		_w1682_,
		_w2509_
	);
	LUT4 #(
		.INIT('h8000)
	) name2047 (
		_w1062_,
		_w1109_,
		_w1229_,
		_w1232_,
		_w2510_
	);
	LUT4 #(
		.INIT('h0057)
	) name2048 (
		\P2_reg2_reg[29]/NET0131 ,
		_w1441_,
		_w1523_,
		_w2510_,
		_w2511_
	);
	LUT4 #(
		.INIT('hef00)
	) name2049 (
		_w546_,
		_w1107_,
		_w1522_,
		_w2511_,
		_w2512_
	);
	LUT2 #(
		.INIT('h4)
	) name2050 (
		_w2509_,
		_w2512_,
		_w2513_
	);
	LUT3 #(
		.INIT('he0)
	) name2051 (
		_w1506_,
		_w2508_,
		_w2513_,
		_w2514_
	);
	LUT4 #(
		.INIT('hc535)
	) name2052 (
		\P2_reg2_reg[29]/NET0131 ,
		_w1264_,
		_w1507_,
		_w1712_,
		_w2515_
	);
	LUT4 #(
		.INIT('h35c5)
	) name2053 (
		\P2_reg2_reg[29]/NET0131 ,
		_w1264_,
		_w1516_,
		_w1678_,
		_w2516_
	);
	LUT4 #(
		.INIT('hfc54)
	) name2054 (
		_w1530_,
		_w1575_,
		_w2515_,
		_w2516_,
		_w2517_
	);
	LUT4 #(
		.INIT('h3111)
	) name2055 (
		_w1359_,
		_w2507_,
		_w2514_,
		_w2517_,
		_w2518_
	);
	LUT3 #(
		.INIT('hce)
	) name2056 (
		\P1_state_reg[0]/NET0131 ,
		_w2506_,
		_w2518_,
		_w2519_
	);
	LUT4 #(
		.INIT('h4500)
	) name2057 (
		_w1734_,
		_w1735_,
		_w1737_,
		_w1739_,
		_w2520_
	);
	LUT4 #(
		.INIT('h30a0)
	) name2058 (
		\P1_reg1_reg[29]/NET0131 ,
		_w2281_,
		_w2292_,
		_w2520_,
		_w2521_
	);
	LUT4 #(
		.INIT('hc0a0)
	) name2059 (
		\P1_reg1_reg[29]/NET0131 ,
		_w2387_,
		_w2388_,
		_w2520_,
		_w2522_
	);
	LUT4 #(
		.INIT('h0355)
	) name2060 (
		\P1_reg1_reg[29]/NET0131 ,
		_w2390_,
		_w2422_,
		_w2520_,
		_w2523_
	);
	LUT4 #(
		.INIT('h5f51)
	) name2061 (
		_w2283_,
		_w2284_,
		_w2288_,
		_w2291_,
		_w2524_
	);
	LUT4 #(
		.INIT('hf100)
	) name2062 (
		_w2426_,
		_w2447_,
		_w2520_,
		_w2524_,
		_w2525_
	);
	LUT2 #(
		.INIT('h2)
	) name2063 (
		\P1_reg1_reg[29]/NET0131 ,
		_w2525_,
		_w2526_
	);
	LUT4 #(
		.INIT('h001f)
	) name2064 (
		_w2427_,
		_w2448_,
		_w2520_,
		_w2526_,
		_w2527_
	);
	LUT3 #(
		.INIT('hd0)
	) name2065 (
		_w2424_,
		_w2523_,
		_w2527_,
		_w2528_
	);
	LUT4 #(
		.INIT('ha8aa)
	) name2066 (
		_w1731_,
		_w2521_,
		_w2522_,
		_w2528_,
		_w2529_
	);
	LUT4 #(
		.INIT('h2000)
	) name2067 (
		\P1_reg1_reg[29]/NET0131 ,
		_w1723_,
		_w1727_,
		_w1730_,
		_w2530_
	);
	LUT2 #(
		.INIT('h2)
	) name2068 (
		\P1_reg1_reg[29]/NET0131 ,
		_w2462_,
		_w2531_
	);
	LUT4 #(
		.INIT('hffa8)
	) name2069 (
		\P1_state_reg[0]/NET0131 ,
		_w2529_,
		_w2530_,
		_w2531_,
		_w2532_
	);
	LUT4 #(
		.INIT('h1000)
	) name2070 (
		_w907_,
		_w1189_,
		_w1352_,
		_w1356_,
		_w2533_
	);
	LUT3 #(
		.INIT('h10)
	) name2071 (
		_w1308_,
		_w1459_,
		_w1531_,
		_w2534_
	);
	LUT3 #(
		.INIT('hb0)
	) name2072 (
		_w1534_,
		_w1535_,
		_w2534_,
		_w2535_
	);
	LUT3 #(
		.INIT('h01)
	) name2073 (
		_w1308_,
		_w1459_,
		_w1536_,
		_w2536_
	);
	LUT2 #(
		.INIT('h1)
	) name2074 (
		_w1541_,
		_w2536_,
		_w2537_
	);
	LUT4 #(
		.INIT('h0001)
	) name2075 (
		_w1318_,
		_w1316_,
		_w1300_,
		_w1467_,
		_w2538_
	);
	LUT3 #(
		.INIT('h0b)
	) name2076 (
		_w1542_,
		_w1546_,
		_w1551_,
		_w2539_
	);
	LUT4 #(
		.INIT('h4f00)
	) name2077 (
		_w2535_,
		_w2537_,
		_w2538_,
		_w2539_,
		_w2540_
	);
	LUT2 #(
		.INIT('h8)
	) name2078 (
		_w1545_,
		_w1548_,
		_w2541_
	);
	LUT3 #(
		.INIT('hd0)
	) name2079 (
		_w1548_,
		_w1552_,
		_w1554_,
		_w2542_
	);
	LUT4 #(
		.INIT('h9a55)
	) name2080 (
		_w1292_,
		_w2540_,
		_w2541_,
		_w2542_,
		_w2543_
	);
	LUT4 #(
		.INIT('h0d01)
	) name2081 (
		_w907_,
		_w1369_,
		_w1496_,
		_w2543_,
		_w2544_
	);
	LUT3 #(
		.INIT('h04)
	) name2082 (
		_w925_,
		_w1232_,
		_w1439_,
		_w2545_
	);
	LUT3 #(
		.INIT('h54)
	) name2083 (
		_w907_,
		_w1441_,
		_w1443_,
		_w2546_
	);
	LUT2 #(
		.INIT('h1)
	) name2084 (
		_w2545_,
		_w2546_,
		_w2547_
	);
	LUT2 #(
		.INIT('h4)
	) name2085 (
		_w2544_,
		_w2547_,
		_w2548_
	);
	LUT3 #(
		.INIT('h07)
	) name2086 (
		_w672_,
		_w930_,
		_w1197_,
		_w2549_
	);
	LUT2 #(
		.INIT('h8)
	) name2087 (
		_w625_,
		_w930_,
		_w2550_
	);
	LUT3 #(
		.INIT('h15)
	) name2088 (
		_w669_,
		_w738_,
		_w1204_,
		_w2551_
	);
	LUT3 #(
		.INIT('h10)
	) name2089 (
		_w720_,
		_w732_,
		_w1214_,
		_w2552_
	);
	LUT2 #(
		.INIT('h1)
	) name2090 (
		_w1203_,
		_w2552_,
		_w2553_
	);
	LUT3 #(
		.INIT('h10)
	) name2091 (
		_w720_,
		_w732_,
		_w764_,
		_w2554_
	);
	LUT3 #(
		.INIT('he0)
	) name2092 (
		_w1212_,
		_w1213_,
		_w2554_,
		_w2555_
	);
	LUT4 #(
		.INIT('h0001)
	) name2093 (
		_w646_,
		_w687_,
		_w704_,
		_w737_,
		_w2556_
	);
	LUT4 #(
		.INIT('h08aa)
	) name2094 (
		_w2551_,
		_w2553_,
		_w2555_,
		_w2556_,
		_w2557_
	);
	LUT4 #(
		.INIT('h9959)
	) name2095 (
		_w1292_,
		_w2549_,
		_w2550_,
		_w2557_,
		_w2558_
	);
	LUT4 #(
		.INIT('h010d)
	) name2096 (
		_w907_,
		_w1369_,
		_w1409_,
		_w2558_,
		_w2559_
	);
	LUT4 #(
		.INIT('hc404)
	) name2097 (
		_w907_,
		_w1447_,
		_w1411_,
		_w2543_,
		_w2560_
	);
	LUT3 #(
		.INIT('h10)
	) name2098 (
		_w845_,
		_w910_,
		_w1423_,
		_w2561_
	);
	LUT4 #(
		.INIT('h0100)
	) name2099 (
		_w845_,
		_w889_,
		_w910_,
		_w1423_,
		_w2562_
	);
	LUT2 #(
		.INIT('h1)
	) name2100 (
		_w845_,
		_w1435_,
		_w2563_
	);
	LUT4 #(
		.INIT('h007b)
	) name2101 (
		_w889_,
		_w1435_,
		_w2561_,
		_w2563_,
		_w2564_
	);
	LUT4 #(
		.INIT('h04c4)
	) name2102 (
		_w907_,
		_w1191_,
		_w1411_,
		_w2564_,
		_w2565_
	);
	LUT3 #(
		.INIT('h01)
	) name2103 (
		_w2560_,
		_w2565_,
		_w2559_,
		_w2566_
	);
	LUT4 #(
		.INIT('h3111)
	) name2104 (
		_w1359_,
		_w2533_,
		_w2548_,
		_w2566_,
		_w2567_
	);
	LUT2 #(
		.INIT('h4)
	) name2105 (
		\P1_state_reg[0]/NET0131 ,
		\P2_reg3_reg[18]/NET0131 ,
		_w2568_
	);
	LUT3 #(
		.INIT('h0b)
	) name2106 (
		_w907_,
		_w1349_,
		_w2568_,
		_w2569_
	);
	LUT3 #(
		.INIT('h2f)
	) name2107 (
		\P1_state_reg[0]/NET0131 ,
		_w2567_,
		_w2569_,
		_w2570_
	);
	LUT4 #(
		.INIT('h1000)
	) name2108 (
		_w886_,
		_w1189_,
		_w1352_,
		_w1356_,
		_w2571_
	);
	LUT4 #(
		.INIT('h0155)
	) name2109 (
		_w886_,
		_w1361_,
		_w1363_,
		_w1368_,
		_w2572_
	);
	LUT4 #(
		.INIT('h6a55)
	) name2110 (
		_w1272_,
		_w1450_,
		_w1471_,
		_w1479_,
		_w2573_
	);
	LUT4 #(
		.INIT('h010d)
	) name2111 (
		_w886_,
		_w1369_,
		_w1496_,
		_w2573_,
		_w2574_
	);
	LUT3 #(
		.INIT('h54)
	) name2112 (
		_w886_,
		_w1441_,
		_w1443_,
		_w2575_
	);
	LUT3 #(
		.INIT('h0b)
	) name2113 (
		_w902_,
		_w1440_,
		_w2575_,
		_w2576_
	);
	LUT2 #(
		.INIT('h4)
	) name2114 (
		_w2574_,
		_w2576_,
		_w2577_
	);
	LUT4 #(
		.INIT('h4844)
	) name2115 (
		_w1272_,
		_w1369_,
		_w1387_,
		_w1394_,
		_w2578_
	);
	LUT3 #(
		.INIT('h54)
	) name2116 (
		_w1409_,
		_w2572_,
		_w2578_,
		_w2579_
	);
	LUT4 #(
		.INIT('h5554)
	) name2117 (
		_w886_,
		_w1361_,
		_w1363_,
		_w1368_,
		_w2580_
	);
	LUT3 #(
		.INIT('h07)
	) name2118 (
		_w906_,
		_w909_,
		_w1435_,
		_w2581_
	);
	LUT4 #(
		.INIT('h1000)
	) name2119 (
		_w845_,
		_w910_,
		_w1423_,
		_w1424_,
		_w2582_
	);
	LUT4 #(
		.INIT('h00c4)
	) name2120 (
		_w969_,
		_w1435_,
		_w2562_,
		_w2582_,
		_w2583_
	);
	LUT4 #(
		.INIT('h1113)
	) name2121 (
		_w1411_,
		_w2580_,
		_w2581_,
		_w2583_,
		_w2584_
	);
	LUT4 #(
		.INIT('h04c4)
	) name2122 (
		_w886_,
		_w1447_,
		_w1411_,
		_w2573_,
		_w2585_
	);
	LUT4 #(
		.INIT('h000d)
	) name2123 (
		_w1191_,
		_w2584_,
		_w2585_,
		_w2579_,
		_w2586_
	);
	LUT4 #(
		.INIT('h3111)
	) name2124 (
		_w1359_,
		_w2571_,
		_w2577_,
		_w2586_,
		_w2587_
	);
	LUT2 #(
		.INIT('h4)
	) name2125 (
		\P1_state_reg[0]/NET0131 ,
		\P2_reg3_reg[19]/NET0131 ,
		_w2588_
	);
	LUT3 #(
		.INIT('h0b)
	) name2126 (
		_w886_,
		_w1349_,
		_w2588_,
		_w2589_
	);
	LUT3 #(
		.INIT('h2f)
	) name2127 (
		\P1_state_reg[0]/NET0131 ,
		_w2587_,
		_w2589_,
		_w2590_
	);
	LUT4 #(
		.INIT('h1000)
	) name2128 (
		_w842_,
		_w1189_,
		_w1352_,
		_w1356_,
		_w2591_
	);
	LUT4 #(
		.INIT('h0155)
	) name2129 (
		_w842_,
		_w1361_,
		_w1363_,
		_w1368_,
		_w2592_
	);
	LUT4 #(
		.INIT('h59aa)
	) name2130 (
		_w1314_,
		_w1692_,
		_w1699_,
		_w1700_,
		_w2593_
	);
	LUT4 #(
		.INIT('h0d01)
	) name2131 (
		_w842_,
		_w1369_,
		_w1496_,
		_w2593_,
		_w2594_
	);
	LUT4 #(
		.INIT('h5554)
	) name2132 (
		_w842_,
		_w1361_,
		_w1363_,
		_w1368_,
		_w2595_
	);
	LUT4 #(
		.INIT('h6300)
	) name2133 (
		_w845_,
		_w910_,
		_w1423_,
		_w1435_,
		_w2596_
	);
	LUT2 #(
		.INIT('h1)
	) name2134 (
		_w866_,
		_w1435_,
		_w2597_
	);
	LUT4 #(
		.INIT('h1113)
	) name2135 (
		_w1411_,
		_w2595_,
		_w2596_,
		_w2597_,
		_w2598_
	);
	LUT3 #(
		.INIT('h54)
	) name2136 (
		_w842_,
		_w1441_,
		_w1443_,
		_w2599_
	);
	LUT3 #(
		.INIT('h04)
	) name2137 (
		_w860_,
		_w1232_,
		_w1439_,
		_w2600_
	);
	LUT2 #(
		.INIT('h1)
	) name2138 (
		_w2599_,
		_w2600_,
		_w2601_
	);
	LUT3 #(
		.INIT('hd0)
	) name2139 (
		_w1191_,
		_w2598_,
		_w2601_,
		_w2602_
	);
	LUT4 #(
		.INIT('hc404)
	) name2140 (
		_w842_,
		_w1447_,
		_w1411_,
		_w2593_,
		_w2603_
	);
	LUT4 #(
		.INIT('h2a22)
	) name2141 (
		_w1658_,
		_w1660_,
		_w1662_,
		_w1663_,
		_w2604_
	);
	LUT4 #(
		.INIT('h4484)
	) name2142 (
		_w1314_,
		_w1369_,
		_w1665_,
		_w2604_,
		_w2605_
	);
	LUT3 #(
		.INIT('h54)
	) name2143 (
		_w1409_,
		_w2592_,
		_w2605_,
		_w2606_
	);
	LUT4 #(
		.INIT('h0100)
	) name2144 (
		_w2594_,
		_w2603_,
		_w2606_,
		_w2602_,
		_w2607_
	);
	LUT4 #(
		.INIT('ha0a8)
	) name2145 (
		\P1_state_reg[0]/NET0131 ,
		_w1359_,
		_w2591_,
		_w2607_,
		_w2608_
	);
	LUT2 #(
		.INIT('h4)
	) name2146 (
		\P1_state_reg[0]/NET0131 ,
		\P2_reg3_reg[17]/NET0131 ,
		_w2609_
	);
	LUT4 #(
		.INIT('h0802)
	) name2147 (
		\P1_state_reg[0]/NET0131 ,
		\P2_IR_reg[23]/NET0131 ,
		_w842_,
		_w1188_,
		_w2610_
	);
	LUT2 #(
		.INIT('h1)
	) name2148 (
		_w2609_,
		_w2610_,
		_w2611_
	);
	LUT2 #(
		.INIT('hb)
	) name2149 (
		_w2608_,
		_w2611_,
		_w2612_
	);
	LUT2 #(
		.INIT('h4)
	) name2150 (
		_w1000_,
		_w1357_,
		_w2613_
	);
	LUT4 #(
		.INIT('h5554)
	) name2151 (
		_w1000_,
		_w1361_,
		_w1363_,
		_w1368_,
		_w2614_
	);
	LUT3 #(
		.INIT('h70)
	) name2152 (
		_w1556_,
		_w1562_,
		_w1566_,
		_w2615_
	);
	LUT4 #(
		.INIT('h0001)
	) name2153 (
		_w1287_,
		_w1290_,
		_w1282_,
		_w1483_,
		_w2616_
	);
	LUT4 #(
		.INIT('h4f00)
	) name2154 (
		_w2540_,
		_w2541_,
		_w2542_,
		_w2616_,
		_w2617_
	);
	LUT4 #(
		.INIT('h4484)
	) name2155 (
		_w1275_,
		_w1411_,
		_w2615_,
		_w2617_,
		_w2618_
	);
	LUT3 #(
		.INIT('ha8)
	) name2156 (
		_w1447_,
		_w2614_,
		_w2618_,
		_w2619_
	);
	LUT4 #(
		.INIT('h0155)
	) name2157 (
		_w1000_,
		_w1361_,
		_w1363_,
		_w1368_,
		_w2620_
	);
	LUT4 #(
		.INIT('h4484)
	) name2158 (
		_w1275_,
		_w1369_,
		_w2615_,
		_w2617_,
		_w2621_
	);
	LUT3 #(
		.INIT('h54)
	) name2159 (
		_w1496_,
		_w2620_,
		_w2621_,
		_w2622_
	);
	LUT3 #(
		.INIT('h40)
	) name2160 (
		_w845_,
		_w1423_,
		_w1426_,
		_w2623_
	);
	LUT4 #(
		.INIT('h1000)
	) name2161 (
		_w845_,
		_w1006_,
		_w1423_,
		_w1426_,
		_w2624_
	);
	LUT3 #(
		.INIT('h0b)
	) name2162 (
		_w948_,
		_w952_,
		_w1435_,
		_w2625_
	);
	LUT4 #(
		.INIT('h007b)
	) name2163 (
		_w989_,
		_w1435_,
		_w2624_,
		_w2625_,
		_w2626_
	);
	LUT4 #(
		.INIT('h04c4)
	) name2164 (
		_w1000_,
		_w1191_,
		_w1411_,
		_w2626_,
		_w2627_
	);
	LUT3 #(
		.INIT('h07)
	) name2165 (
		_w1015_,
		_w1199_,
		_w1218_,
		_w2628_
	);
	LUT4 #(
		.INIT('h0001)
	) name2166 (
		_w928_,
		_w929_,
		_w1013_,
		_w1014_,
		_w2629_
	);
	LUT3 #(
		.INIT('h80)
	) name2167 (
		_w625_,
		_w930_,
		_w2556_,
		_w2630_
	);
	LUT2 #(
		.INIT('h8)
	) name2168 (
		_w2555_,
		_w2630_,
		_w2631_
	);
	LUT3 #(
		.INIT('he0)
	) name2169 (
		_w1203_,
		_w2552_,
		_w2556_,
		_w2632_
	);
	LUT4 #(
		.INIT('h22a2)
	) name2170 (
		_w2549_,
		_w2550_,
		_w2551_,
		_w2632_,
		_w2633_
	);
	LUT4 #(
		.INIT('h2a22)
	) name2171 (
		_w2628_,
		_w2629_,
		_w2631_,
		_w2633_,
		_w2634_
	);
	LUT4 #(
		.INIT('h0b07)
	) name2172 (
		_w1275_,
		_w1369_,
		_w2620_,
		_w2634_,
		_w2635_
	);
	LUT3 #(
		.INIT('h54)
	) name2173 (
		_w1000_,
		_w1441_,
		_w1443_,
		_w2636_
	);
	LUT4 #(
		.INIT('h0010)
	) name2174 (
		_w546_,
		_w999_,
		_w1232_,
		_w1439_,
		_w2637_
	);
	LUT2 #(
		.INIT('h1)
	) name2175 (
		_w2636_,
		_w2637_,
		_w2638_
	);
	LUT4 #(
		.INIT('h3200)
	) name2176 (
		_w1409_,
		_w2627_,
		_w2635_,
		_w2638_,
		_w2639_
	);
	LUT4 #(
		.INIT('ha8aa)
	) name2177 (
		_w1359_,
		_w2622_,
		_w2619_,
		_w2639_,
		_w2640_
	);
	LUT4 #(
		.INIT('h93bb)
	) name2178 (
		\P1_state_reg[0]/NET0131 ,
		\P2_reg3_reg[22]/NET0131 ,
		_w946_,
		_w1189_,
		_w2641_
	);
	LUT4 #(
		.INIT('ha8ff)
	) name2179 (
		\P1_state_reg[0]/NET0131 ,
		_w2613_,
		_w2640_,
		_w2641_,
		_w2642_
	);
	LUT2 #(
		.INIT('h8)
	) name2180 (
		_w1932_,
		_w2460_,
		_w2643_
	);
	LUT4 #(
		.INIT('h8acf)
	) name2181 (
		_w1734_,
		_w1735_,
		_w1737_,
		_w1739_,
		_w2644_
	);
	LUT2 #(
		.INIT('h2)
	) name2182 (
		_w1932_,
		_w2644_,
		_w2645_
	);
	LUT4 #(
		.INIT('h54ab)
	) name2183 (
		_w1748_,
		_w1907_,
		_w1929_,
		_w1936_,
		_w2646_
	);
	LUT3 #(
		.INIT('h8a)
	) name2184 (
		_w1990_,
		_w2259_,
		_w2264_,
		_w2647_
	);
	LUT3 #(
		.INIT('h01)
	) name2185 (
		_w1878_,
		_w1954_,
		_w1964_,
		_w2648_
	);
	LUT4 #(
		.INIT('h7500)
	) name2186 (
		_w1990_,
		_w2259_,
		_w2264_,
		_w2648_,
		_w2649_
	);
	LUT4 #(
		.INIT('h4504)
	) name2187 (
		_w1878_,
		_w1948_,
		_w1952_,
		_w1992_,
		_w2650_
	);
	LUT2 #(
		.INIT('h2)
	) name2188 (
		_w1996_,
		_w2650_,
		_w2651_
	);
	LUT3 #(
		.INIT('h45)
	) name2189 (
		_w1906_,
		_w2649_,
		_w2651_,
		_w2652_
	);
	LUT4 #(
		.INIT('h0001)
	) name2190 (
		_w2036_,
		_w2110_,
		_w2120_,
		_w2150_,
		_w2653_
	);
	LUT4 #(
		.INIT('hf800)
	) name2191 (
		_w2096_,
		_w2141_,
		_w2145_,
		_w2653_,
		_w2654_
	);
	LUT3 #(
		.INIT('h45)
	) name2192 (
		_w2047_,
		_w2148_,
		_w2151_,
		_w2655_
	);
	LUT2 #(
		.INIT('h8)
	) name2193 (
		_w2022_,
		_w2225_,
		_w2656_
	);
	LUT2 #(
		.INIT('h8)
	) name2194 (
		_w2203_,
		_w2248_,
		_w2657_
	);
	LUT4 #(
		.INIT('h8000)
	) name2195 (
		_w2022_,
		_w2203_,
		_w2225_,
		_w2248_,
		_w2658_
	);
	LUT3 #(
		.INIT('h07)
	) name2196 (
		_w2048_,
		_w2225_,
		_w2251_,
		_w2659_
	);
	LUT3 #(
		.INIT('h07)
	) name2197 (
		_w2203_,
		_w2252_,
		_w2255_,
		_w2660_
	);
	LUT3 #(
		.INIT('hd0)
	) name2198 (
		_w2657_,
		_w2659_,
		_w2660_,
		_w2661_
	);
	LUT4 #(
		.INIT('h4f00)
	) name2199 (
		_w2654_,
		_w2655_,
		_w2658_,
		_w2661_,
		_w2662_
	);
	LUT4 #(
		.INIT('h0001)
	) name2200 (
		_w1978_,
		_w2165_,
		_w2177_,
		_w2263_,
		_w2663_
	);
	LUT3 #(
		.INIT('h40)
	) name2201 (
		_w1906_,
		_w2648_,
		_w2663_,
		_w2664_
	);
	LUT4 #(
		.INIT('h9a99)
	) name2202 (
		_w2646_,
		_w2652_,
		_w2662_,
		_w2664_,
		_w2665_
	);
	LUT4 #(
		.INIT('h08c8)
	) name2203 (
		_w1932_,
		_w2292_,
		_w2644_,
		_w2665_,
		_w2666_
	);
	LUT4 #(
		.INIT('he000)
	) name2204 (
		_w2316_,
		_w2320_,
		_w2323_,
		_w2329_,
		_w2667_
	);
	LUT3 #(
		.INIT('h15)
	) name2205 (
		_w2298_,
		_w2326_,
		_w2329_,
		_w2668_
	);
	LUT2 #(
		.INIT('h8)
	) name2206 (
		_w2294_,
		_w2352_,
		_w2669_
	);
	LUT2 #(
		.INIT('h8)
	) name2207 (
		_w2331_,
		_w2350_,
		_w2670_
	);
	LUT4 #(
		.INIT('h8000)
	) name2208 (
		_w2294_,
		_w2331_,
		_w2350_,
		_w2352_,
		_w2671_
	);
	LUT3 #(
		.INIT('h23)
	) name2209 (
		_w2300_,
		_w2333_,
		_w2352_,
		_w2672_
	);
	LUT3 #(
		.INIT('h13)
	) name2210 (
		_w2335_,
		_w2342_,
		_w2350_,
		_w2673_
	);
	LUT3 #(
		.INIT('hd0)
	) name2211 (
		_w2670_,
		_w2672_,
		_w2673_,
		_w2674_
	);
	LUT4 #(
		.INIT('h4f00)
	) name2212 (
		_w2667_,
		_w2668_,
		_w2671_,
		_w2674_,
		_w2675_
	);
	LUT4 #(
		.INIT('h0001)
	) name2213 (
		_w2337_,
		_w2338_,
		_w2363_,
		_w2364_,
		_w2676_
	);
	LUT2 #(
		.INIT('h8)
	) name2214 (
		_w2361_,
		_w2368_,
		_w2677_
	);
	LUT3 #(
		.INIT('h80)
	) name2215 (
		_w2361_,
		_w2368_,
		_w2676_,
		_w2678_
	);
	LUT3 #(
		.INIT('h07)
	) name2216 (
		_w2346_,
		_w2365_,
		_w2374_,
		_w2679_
	);
	LUT3 #(
		.INIT('h0d)
	) name2217 (
		_w2361_,
		_w2377_,
		_w2381_,
		_w2680_
	);
	LUT3 #(
		.INIT('hd0)
	) name2218 (
		_w2677_,
		_w2679_,
		_w2680_,
		_w2681_
	);
	LUT4 #(
		.INIT('h9a55)
	) name2219 (
		_w2646_,
		_w2675_,
		_w2678_,
		_w2681_,
		_w2682_
	);
	LUT4 #(
		.INIT('h08c8)
	) name2220 (
		_w1932_,
		_w2388_,
		_w2644_,
		_w2682_,
		_w2683_
	);
	LUT2 #(
		.INIT('h2)
	) name2221 (
		_w1747_,
		_w1904_,
		_w2684_
	);
	LUT4 #(
		.INIT('h8000)
	) name2222 (
		_w2394_,
		_w2404_,
		_w2408_,
		_w2414_,
		_w2685_
	);
	LUT4 #(
		.INIT('h0501)
	) name2223 (
		_w1747_,
		_w1836_,
		_w2416_,
		_w2685_,
		_w2686_
	);
	LUT4 #(
		.INIT('h1113)
	) name2224 (
		_w2644_,
		_w2645_,
		_w2684_,
		_w2686_,
		_w2687_
	);
	LUT4 #(
		.INIT('h6300)
	) name2225 (
		_w1900_,
		_w1931_,
		_w2443_,
		_w2447_,
		_w2688_
	);
	LUT3 #(
		.INIT('h13)
	) name2226 (
		_w2426_,
		_w2454_,
		_w2644_,
		_w2689_
	);
	LUT4 #(
		.INIT('h0f01)
	) name2227 (
		_w2426_,
		_w2447_,
		_w2450_,
		_w2644_,
		_w2690_
	);
	LUT4 #(
		.INIT('hf531)
	) name2228 (
		_w1931_,
		_w1932_,
		_w2689_,
		_w2690_,
		_w2691_
	);
	LUT3 #(
		.INIT('h70)
	) name2229 (
		_w2644_,
		_w2688_,
		_w2691_,
		_w2692_
	);
	LUT3 #(
		.INIT('hd0)
	) name2230 (
		_w2424_,
		_w2687_,
		_w2692_,
		_w2693_
	);
	LUT4 #(
		.INIT('ha8aa)
	) name2231 (
		_w1731_,
		_w2666_,
		_w2683_,
		_w2693_,
		_w2694_
	);
	LUT4 #(
		.INIT('ha060)
	) name2232 (
		\P1_IR_reg[23]/NET0131 ,
		\P1_IR_reg[31]/NET0131 ,
		\P1_state_reg[0]/NET0131 ,
		_w1722_,
		_w2695_
	);
	LUT4 #(
		.INIT('h9d5d)
	) name2233 (
		\P1_reg3_reg[27]/NET0131 ,
		\P1_state_reg[0]/NET0131 ,
		_w1723_,
		_w1830_,
		_w2696_
	);
	LUT4 #(
		.INIT('ha8ff)
	) name2234 (
		\P1_state_reg[0]/NET0131 ,
		_w2643_,
		_w2694_,
		_w2696_,
		_w2697_
	);
	LUT4 #(
		.INIT('hd070)
	) name2235 (
		\P1_state_reg[0]/NET0131 ,
		\P2_IR_reg[23]/NET0131 ,
		\P2_reg2_reg[22]/NET0131 ,
		_w1188_,
		_w2698_
	);
	LUT4 #(
		.INIT('h2000)
	) name2236 (
		\P2_reg2_reg[22]/NET0131 ,
		_w1189_,
		_w1352_,
		_w1356_,
		_w2699_
	);
	LUT4 #(
		.INIT('ha8aa)
	) name2237 (
		\P2_reg2_reg[22]/NET0131 ,
		_w1361_,
		_w1363_,
		_w1368_,
		_w2700_
	);
	LUT4 #(
		.INIT('h4484)
	) name2238 (
		_w1275_,
		_w1507_,
		_w2615_,
		_w2617_,
		_w2701_
	);
	LUT3 #(
		.INIT('h54)
	) name2239 (
		_w1575_,
		_w2700_,
		_w2701_,
		_w2702_
	);
	LUT4 #(
		.INIT('h08c8)
	) name2240 (
		\P2_reg2_reg[22]/NET0131 ,
		_w1191_,
		_w1516_,
		_w2626_,
		_w2703_
	);
	LUT4 #(
		.INIT('hc535)
	) name2241 (
		\P2_reg2_reg[22]/NET0131 ,
		_w1275_,
		_w1516_,
		_w2634_,
		_w2704_
	);
	LUT2 #(
		.INIT('h2)
	) name2242 (
		_w1530_,
		_w2704_,
		_w2705_
	);
	LUT4 #(
		.INIT('hc535)
	) name2243 (
		\P2_reg2_reg[22]/NET0131 ,
		_w1275_,
		_w1507_,
		_w2634_,
		_w2706_
	);
	LUT4 #(
		.INIT('h1000)
	) name2244 (
		_w546_,
		_w999_,
		_w1442_,
		_w1507_,
		_w2707_
	);
	LUT4 #(
		.INIT('h6000)
	) name2245 (
		\P2_reg3_reg[22]/NET0131 ,
		_w946_,
		_w1229_,
		_w1232_,
		_w2708_
	);
	LUT4 #(
		.INIT('h0057)
	) name2246 (
		\P2_reg2_reg[22]/NET0131 ,
		_w1441_,
		_w1523_,
		_w2708_,
		_w2709_
	);
	LUT2 #(
		.INIT('h4)
	) name2247 (
		_w2707_,
		_w2709_,
		_w2710_
	);
	LUT3 #(
		.INIT('he0)
	) name2248 (
		_w1506_,
		_w2706_,
		_w2710_,
		_w2711_
	);
	LUT4 #(
		.INIT('h0100)
	) name2249 (
		_w2702_,
		_w2703_,
		_w2705_,
		_w2711_,
		_w2712_
	);
	LUT4 #(
		.INIT('ha0a8)
	) name2250 (
		\P1_state_reg[0]/NET0131 ,
		_w1359_,
		_w2699_,
		_w2712_,
		_w2713_
	);
	LUT2 #(
		.INIT('he)
	) name2251 (
		_w2698_,
		_w2713_,
		_w2714_
	);
	LUT4 #(
		.INIT('hd070)
	) name2252 (
		\P1_state_reg[0]/NET0131 ,
		\P2_IR_reg[23]/NET0131 ,
		\P2_reg0_reg[27]/NET0131 ,
		_w1188_,
		_w2715_
	);
	LUT4 #(
		.INIT('h2000)
	) name2253 (
		\P2_reg0_reg[27]/NET0131 ,
		_w1189_,
		_w1352_,
		_w1356_,
		_w2716_
	);
	LUT4 #(
		.INIT('haaa8)
	) name2254 (
		\P2_reg0_reg[27]/NET0131 ,
		_w1361_,
		_w1363_,
		_w1368_,
		_w2717_
	);
	LUT4 #(
		.INIT('h9a00)
	) name2255 (
		_w1263_,
		_w1400_,
		_w1407_,
		_w1411_,
		_w2718_
	);
	LUT3 #(
		.INIT('h54)
	) name2256 (
		_w1409_,
		_w2717_,
		_w2718_,
		_w2719_
	);
	LUT4 #(
		.INIT('h02aa)
	) name2257 (
		\P2_reg0_reg[27]/NET0131 ,
		_w1361_,
		_w1363_,
		_w1368_,
		_w2720_
	);
	LUT4 #(
		.INIT('h08c8)
	) name2258 (
		\P2_reg0_reg[27]/NET0131 ,
		_w1191_,
		_w1369_,
		_w1437_,
		_w2721_
	);
	LUT3 #(
		.INIT('ha2)
	) name2259 (
		\P2_reg0_reg[27]/NET0131 ,
		_w1684_,
		_w1685_,
		_w2722_
	);
	LUT4 #(
		.INIT('h00ef)
	) name2260 (
		_w546_,
		_w1078_,
		_w1687_,
		_w2722_,
		_w2723_
	);
	LUT2 #(
		.INIT('h4)
	) name2261 (
		_w2721_,
		_w2723_,
		_w2724_
	);
	LUT3 #(
		.INIT('ha8)
	) name2262 (
		_w1447_,
		_w1497_,
		_w2720_,
		_w2725_
	);
	LUT3 #(
		.INIT('h32)
	) name2263 (
		_w1494_,
		_w1496_,
		_w2717_,
		_w2726_
	);
	LUT4 #(
		.INIT('h0100)
	) name2264 (
		_w2719_,
		_w2725_,
		_w2726_,
		_w2724_,
		_w2727_
	);
	LUT4 #(
		.INIT('ha0a8)
	) name2265 (
		\P1_state_reg[0]/NET0131 ,
		_w1359_,
		_w2716_,
		_w2727_,
		_w2728_
	);
	LUT2 #(
		.INIT('he)
	) name2266 (
		_w2715_,
		_w2728_,
		_w2729_
	);
	LUT4 #(
		.INIT('hd070)
	) name2267 (
		\P1_state_reg[0]/NET0131 ,
		\P2_IR_reg[23]/NET0131 ,
		\P2_reg0_reg[28]/NET0131 ,
		_w1188_,
		_w2730_
	);
	LUT4 #(
		.INIT('h2000)
	) name2268 (
		\P2_reg0_reg[28]/NET0131 ,
		_w1189_,
		_w1352_,
		_w1356_,
		_w2731_
	);
	LUT4 #(
		.INIT('hc535)
	) name2269 (
		\P2_reg0_reg[28]/NET0131 ,
		_w1260_,
		_w1411_,
		_w1514_,
		_w2732_
	);
	LUT4 #(
		.INIT('h111d)
	) name2270 (
		\P2_reg0_reg[28]/NET0131 ,
		_w1369_,
		_w1517_,
		_w1520_,
		_w2733_
	);
	LUT4 #(
		.INIT('h1000)
	) name2271 (
		_w546_,
		_w1124_,
		_w1411_,
		_w1442_,
		_w2734_
	);
	LUT3 #(
		.INIT('ha2)
	) name2272 (
		\P2_reg0_reg[28]/NET0131 ,
		_w1684_,
		_w1685_,
		_w2735_
	);
	LUT2 #(
		.INIT('h1)
	) name2273 (
		_w2734_,
		_w2735_,
		_w2736_
	);
	LUT3 #(
		.INIT('hd0)
	) name2274 (
		_w1191_,
		_w2733_,
		_w2736_,
		_w2737_
	);
	LUT3 #(
		.INIT('he0)
	) name2275 (
		_w1409_,
		_w2732_,
		_w2737_,
		_w2738_
	);
	LUT4 #(
		.INIT('h35c5)
	) name2276 (
		\P2_reg0_reg[28]/NET0131 ,
		_w1260_,
		_w1411_,
		_w1573_,
		_w2739_
	);
	LUT4 #(
		.INIT('h35c5)
	) name2277 (
		\P2_reg0_reg[28]/NET0131 ,
		_w1260_,
		_w1369_,
		_w1573_,
		_w2740_
	);
	LUT4 #(
		.INIT('hfc54)
	) name2278 (
		_w1447_,
		_w1496_,
		_w2739_,
		_w2740_,
		_w2741_
	);
	LUT4 #(
		.INIT('h3111)
	) name2279 (
		_w1359_,
		_w2731_,
		_w2738_,
		_w2741_,
		_w2742_
	);
	LUT3 #(
		.INIT('hce)
	) name2280 (
		\P1_state_reg[0]/NET0131 ,
		_w2730_,
		_w2742_,
		_w2743_
	);
	LUT2 #(
		.INIT('h2)
	) name2281 (
		\P1_reg2_reg[28]/NET0131 ,
		_w2462_,
		_w2744_
	);
	LUT4 #(
		.INIT('h2000)
	) name2282 (
		\P1_reg2_reg[28]/NET0131 ,
		_w1723_,
		_w1727_,
		_w1730_,
		_w2745_
	);
	LUT2 #(
		.INIT('h1)
	) name2283 (
		_w2120_,
		_w2130_,
		_w2746_
	);
	LUT3 #(
		.INIT('h0b)
	) name2284 (
		_w2072_,
		_w2074_,
		_w2094_,
		_w2747_
	);
	LUT2 #(
		.INIT('h1)
	) name2285 (
		_w2058_,
		_w2140_,
		_w2748_
	);
	LUT4 #(
		.INIT('h2f00)
	) name2286 (
		_w2073_,
		_w2091_,
		_w2747_,
		_w2748_,
		_w2749_
	);
	LUT3 #(
		.INIT('h32)
	) name2287 (
		_w2093_,
		_w2140_,
		_w2144_,
		_w2750_
	);
	LUT3 #(
		.INIT('h54)
	) name2288 (
		_w2120_,
		_w2143_,
		_w2147_,
		_w2751_
	);
	LUT4 #(
		.INIT('h0057)
	) name2289 (
		_w2746_,
		_w2749_,
		_w2750_,
		_w2751_,
		_w2752_
	);
	LUT2 #(
		.INIT('h1)
	) name2290 (
		_w2110_,
		_w2150_,
		_w2753_
	);
	LUT3 #(
		.INIT('h0b)
	) name2291 (
		_w2004_,
		_w2008_,
		_w2036_,
		_w2754_
	);
	LUT2 #(
		.INIT('h8)
	) name2292 (
		_w2753_,
		_w2754_,
		_w2755_
	);
	LUT3 #(
		.INIT('h51)
	) name2293 (
		_w2046_,
		_w2146_,
		_w2150_,
		_w2756_
	);
	LUT3 #(
		.INIT('h4d)
	) name2294 (
		_w2004_,
		_w2008_,
		_w2037_,
		_w2757_
	);
	LUT3 #(
		.INIT('hd0)
	) name2295 (
		_w2754_,
		_w2756_,
		_w2757_,
		_w2758_
	);
	LUT4 #(
		.INIT('hb0bb)
	) name2296 (
		_w2208_,
		_w2212_,
		_w2242_,
		_w2246_,
		_w2759_
	);
	LUT4 #(
		.INIT('hb0bb)
	) name2297 (
		_w2016_,
		_w2020_,
		_w2219_,
		_w2223_,
		_w2760_
	);
	LUT2 #(
		.INIT('h8)
	) name2298 (
		_w2759_,
		_w2760_,
		_w2761_
	);
	LUT4 #(
		.INIT('hb0bb)
	) name2299 (
		_w2183_,
		_w2187_,
		_w2231_,
		_w2235_,
		_w2762_
	);
	LUT3 #(
		.INIT('h10)
	) name2300 (
		_w2177_,
		_w2202_,
		_w2762_,
		_w2763_
	);
	LUT2 #(
		.INIT('h8)
	) name2301 (
		_w2761_,
		_w2763_,
		_w2764_
	);
	LUT4 #(
		.INIT('h4f00)
	) name2302 (
		_w2752_,
		_w2755_,
		_w2758_,
		_w2764_,
		_w2765_
	);
	LUT4 #(
		.INIT('h20f2)
	) name2303 (
		_w2016_,
		_w2020_,
		_w2219_,
		_w2223_,
		_w2766_
	);
	LUT4 #(
		.INIT('h20f2)
	) name2304 (
		_w2208_,
		_w2212_,
		_w2242_,
		_w2246_,
		_w2767_
	);
	LUT3 #(
		.INIT('h07)
	) name2305 (
		_w2759_,
		_w2766_,
		_w2767_,
		_w2768_
	);
	LUT4 #(
		.INIT('hdd4d)
	) name2306 (
		_w2183_,
		_w2187_,
		_w2231_,
		_w2235_,
		_w2769_
	);
	LUT3 #(
		.INIT('h01)
	) name2307 (
		_w2177_,
		_w2202_,
		_w2769_,
		_w2770_
	);
	LUT3 #(
		.INIT('h54)
	) name2308 (
		_w2177_,
		_w2254_,
		_w2258_,
		_w2771_
	);
	LUT2 #(
		.INIT('h1)
	) name2309 (
		_w2770_,
		_w2771_,
		_w2772_
	);
	LUT4 #(
		.INIT('h000d)
	) name2310 (
		_w2763_,
		_w2768_,
		_w2770_,
		_w2771_,
		_w2773_
	);
	LUT2 #(
		.INIT('h1)
	) name2311 (
		_w2165_,
		_w2263_,
		_w2774_
	);
	LUT2 #(
		.INIT('h1)
	) name2312 (
		_w1964_,
		_w1978_,
		_w2775_
	);
	LUT4 #(
		.INIT('h0001)
	) name2313 (
		_w1964_,
		_w1978_,
		_w2165_,
		_w2263_,
		_w2776_
	);
	LUT3 #(
		.INIT('h04)
	) name2314 (
		_w1878_,
		_w1939_,
		_w1954_,
		_w2777_
	);
	LUT4 #(
		.INIT('h0400)
	) name2315 (
		_w1878_,
		_w1939_,
		_w1954_,
		_w2776_,
		_w2778_
	);
	LUT3 #(
		.INIT('h51)
	) name2316 (
		_w1989_,
		_w2257_,
		_w2263_,
		_w2779_
	);
	LUT3 #(
		.INIT('h0b)
	) name2317 (
		_w1964_,
		_w1977_,
		_w1992_,
		_w2780_
	);
	LUT3 #(
		.INIT('hd0)
	) name2318 (
		_w2775_,
		_w2779_,
		_w2780_,
		_w2781_
	);
	LUT2 #(
		.INIT('h1)
	) name2319 (
		_w1991_,
		_w1995_,
		_w2782_
	);
	LUT3 #(
		.INIT('h04)
	) name2320 (
		_w1878_,
		_w1939_,
		_w2782_,
		_w2783_
	);
	LUT4 #(
		.INIT('h0001)
	) name2321 (
		_w1748_,
		_w1899_,
		_w1904_,
		_w1938_,
		_w2784_
	);
	LUT2 #(
		.INIT('h1)
	) name2322 (
		_w1997_,
		_w2784_,
		_w2785_
	);
	LUT4 #(
		.INIT('h0d00)
	) name2323 (
		_w2777_,
		_w2781_,
		_w2783_,
		_w2785_,
		_w2786_
	);
	LUT4 #(
		.INIT('h4f00)
	) name2324 (
		_w2765_,
		_w2773_,
		_w2778_,
		_w2786_,
		_w2787_
	);
	LUT3 #(
		.INIT('h1e)
	) name2325 (
		_w1748_,
		_w1815_,
		_w1836_,
		_w2788_
	);
	LUT4 #(
		.INIT('h1dd1)
	) name2326 (
		\P1_reg2_reg[28]/NET0131 ,
		_w1741_,
		_w2787_,
		_w2788_,
		_w2789_
	);
	LUT4 #(
		.INIT('h0777)
	) name2327 (
		_w2183_,
		_w2187_,
		_w2231_,
		_w2235_,
		_w2790_
	);
	LUT3 #(
		.INIT('h10)
	) name2328 (
		_w2338_,
		_w2339_,
		_w2790_,
		_w2791_
	);
	LUT3 #(
		.INIT('hb2)
	) name2329 (
		_w2077_,
		_w2081_,
		_w2305_,
		_w2792_
	);
	LUT3 #(
		.INIT('h0e)
	) name2330 (
		_w2303_,
		_w2306_,
		_w2309_,
		_w2793_
	);
	LUT2 #(
		.INIT('h1)
	) name2331 (
		_w2311_,
		_w2322_,
		_w2794_
	);
	LUT4 #(
		.INIT('h0001)
	) name2332 (
		_w2311_,
		_w2312_,
		_w2313_,
		_w2322_,
		_w2795_
	);
	LUT4 #(
		.INIT('hf200)
	) name2333 (
		_w2310_,
		_w2792_,
		_w2793_,
		_w2795_,
		_w2796_
	);
	LUT3 #(
		.INIT('h32)
	) name2334 (
		_w2302_,
		_w2313_,
		_w2318_,
		_w2797_
	);
	LUT3 #(
		.INIT('h0d)
	) name2335 (
		_w2317_,
		_w2322_,
		_w2325_,
		_w2798_
	);
	LUT3 #(
		.INIT('h70)
	) name2336 (
		_w2794_,
		_w2797_,
		_w2798_,
		_w2799_
	);
	LUT2 #(
		.INIT('h1)
	) name2337 (
		_w2321_,
		_w2328_,
		_w2800_
	);
	LUT3 #(
		.INIT('h07)
	) name2338 (
		_w2004_,
		_w2008_,
		_w2295_,
		_w2801_
	);
	LUT2 #(
		.INIT('h8)
	) name2339 (
		_w2800_,
		_w2801_,
		_w2802_
	);
	LUT3 #(
		.INIT('h0e)
	) name2340 (
		_w2296_,
		_w2324_,
		_w2328_,
		_w2803_
	);
	LUT3 #(
		.INIT('h0e)
	) name2341 (
		_w2004_,
		_w2008_,
		_w2297_,
		_w2804_
	);
	LUT3 #(
		.INIT('h71)
	) name2342 (
		_w2004_,
		_w2008_,
		_w2297_,
		_w2805_
	);
	LUT3 #(
		.INIT('h07)
	) name2343 (
		_w2801_,
		_w2803_,
		_w2805_,
		_w2806_
	);
	LUT4 #(
		.INIT('h4f00)
	) name2344 (
		_w2796_,
		_w2799_,
		_w2802_,
		_w2806_,
		_w2807_
	);
	LUT4 #(
		.INIT('h0777)
	) name2345 (
		_w2208_,
		_w2212_,
		_w2242_,
		_w2246_,
		_w2808_
	);
	LUT4 #(
		.INIT('h0777)
	) name2346 (
		_w2016_,
		_w2020_,
		_w2219_,
		_w2223_,
		_w2809_
	);
	LUT2 #(
		.INIT('h8)
	) name2347 (
		_w2808_,
		_w2809_,
		_w2810_
	);
	LUT4 #(
		.INIT('heee0)
	) name2348 (
		_w2016_,
		_w2020_,
		_w2219_,
		_w2223_,
		_w2811_
	);
	LUT4 #(
		.INIT('h011f)
	) name2349 (
		_w2016_,
		_w2020_,
		_w2219_,
		_w2223_,
		_w2812_
	);
	LUT4 #(
		.INIT('heee0)
	) name2350 (
		_w2208_,
		_w2212_,
		_w2242_,
		_w2246_,
		_w2813_
	);
	LUT4 #(
		.INIT('h011f)
	) name2351 (
		_w2208_,
		_w2212_,
		_w2242_,
		_w2246_,
		_w2814_
	);
	LUT3 #(
		.INIT('h07)
	) name2352 (
		_w2808_,
		_w2812_,
		_w2814_,
		_w2815_
	);
	LUT4 #(
		.INIT('heee0)
	) name2353 (
		_w2183_,
		_w2187_,
		_w2231_,
		_w2235_,
		_w2816_
	);
	LUT4 #(
		.INIT('h1117)
	) name2354 (
		_w2183_,
		_w2187_,
		_w2231_,
		_w2235_,
		_w2817_
	);
	LUT3 #(
		.INIT('h10)
	) name2355 (
		_w2338_,
		_w2339_,
		_w2817_,
		_w2818_
	);
	LUT3 #(
		.INIT('h54)
	) name2356 (
		_w2338_,
		_w2340_,
		_w2345_,
		_w2819_
	);
	LUT2 #(
		.INIT('h1)
	) name2357 (
		_w2818_,
		_w2819_,
		_w2820_
	);
	LUT4 #(
		.INIT('h000d)
	) name2358 (
		_w2791_,
		_w2815_,
		_w2818_,
		_w2819_,
		_w2821_
	);
	LUT4 #(
		.INIT('hdf00)
	) name2359 (
		_w2791_,
		_w2807_,
		_w2810_,
		_w2821_,
		_w2822_
	);
	LUT2 #(
		.INIT('h1)
	) name2360 (
		_w2337_,
		_w2363_,
		_w2823_
	);
	LUT2 #(
		.INIT('h1)
	) name2361 (
		_w2364_,
		_w2366_,
		_w2824_
	);
	LUT4 #(
		.INIT('h0001)
	) name2362 (
		_w2337_,
		_w2363_,
		_w2364_,
		_w2366_,
		_w2825_
	);
	LUT2 #(
		.INIT('h1)
	) name2363 (
		_w2359_,
		_w2367_,
		_w2826_
	);
	LUT4 #(
		.INIT('h00ef)
	) name2364 (
		_w1748_,
		_w1899_,
		_w1904_,
		_w2356_,
		_w2827_
	);
	LUT2 #(
		.INIT('h8)
	) name2365 (
		_w2826_,
		_w2827_,
		_w2828_
	);
	LUT3 #(
		.INIT('h80)
	) name2366 (
		_w2825_,
		_w2826_,
		_w2827_,
		_w2829_
	);
	LUT3 #(
		.INIT('h0d)
	) name2367 (
		_w2344_,
		_w2363_,
		_w2373_,
		_w2830_
	);
	LUT2 #(
		.INIT('h1)
	) name2368 (
		_w2372_,
		_w2376_,
		_w2831_
	);
	LUT3 #(
		.INIT('h54)
	) name2369 (
		_w2366_,
		_w2372_,
		_w2376_,
		_w2832_
	);
	LUT3 #(
		.INIT('h0d)
	) name2370 (
		_w2824_,
		_w2830_,
		_w2832_,
		_w2833_
	);
	LUT4 #(
		.INIT('h00f1)
	) name2371 (
		_w1748_,
		_w1899_,
		_w1904_,
		_w2383_,
		_w2834_
	);
	LUT2 #(
		.INIT('h1)
	) name2372 (
		_w2375_,
		_w2379_,
		_w2835_
	);
	LUT3 #(
		.INIT('h54)
	) name2373 (
		_w2359_,
		_w2375_,
		_w2379_,
		_w2836_
	);
	LUT4 #(
		.INIT('h1505)
	) name2374 (
		_w2356_,
		_w2360_,
		_w2834_,
		_w2836_,
		_w2837_
	);
	LUT3 #(
		.INIT('h0d)
	) name2375 (
		_w2828_,
		_w2833_,
		_w2837_,
		_w2838_
	);
	LUT4 #(
		.INIT('h9a55)
	) name2376 (
		_w2788_,
		_w2822_,
		_w2829_,
		_w2838_,
		_w2839_
	);
	LUT4 #(
		.INIT('h20e0)
	) name2377 (
		\P1_reg2_reg[28]/NET0131 ,
		_w1741_,
		_w2388_,
		_w2839_,
		_w2840_
	);
	LUT3 #(
		.INIT('h10)
	) name2378 (
		_w1748_,
		_w1815_,
		_w2426_,
		_w2841_
	);
	LUT4 #(
		.INIT('ha8aa)
	) name2379 (
		_w1816_,
		_w1900_,
		_w1931_,
		_w2443_,
		_w2842_
	);
	LUT4 #(
		.INIT('h0f0b)
	) name2380 (
		_w2445_,
		_w2447_,
		_w2841_,
		_w2842_,
		_w2843_
	);
	LUT4 #(
		.INIT('h0200)
	) name2381 (
		_w1747_,
		_w1934_,
		_w1933_,
		_w1935_,
		_w2844_
	);
	LUT4 #(
		.INIT('h00eb)
	) name2382 (
		_w1747_,
		_w2276_,
		_w2416_,
		_w2844_,
		_w2845_
	);
	LUT4 #(
		.INIT('he020)
	) name2383 (
		\P1_reg2_reg[28]/NET0131 ,
		_w1741_,
		_w2424_,
		_w2845_,
		_w2846_
	);
	LUT4 #(
		.INIT('ha2a0)
	) name2384 (
		\P1_reg2_reg[28]/NET0131 ,
		_w1741_,
		_w2450_,
		_w2452_,
		_w2847_
	);
	LUT2 #(
		.INIT('h8)
	) name2385 (
		_w1833_,
		_w2454_,
		_w2848_
	);
	LUT2 #(
		.INIT('h1)
	) name2386 (
		_w2847_,
		_w2848_,
		_w2849_
	);
	LUT4 #(
		.INIT('h0d00)
	) name2387 (
		_w1741_,
		_w2843_,
		_w2846_,
		_w2849_,
		_w2850_
	);
	LUT4 #(
		.INIT('h0d00)
	) name2388 (
		_w2292_,
		_w2789_,
		_w2840_,
		_w2850_,
		_w2851_
	);
	LUT4 #(
		.INIT('ha0a8)
	) name2389 (
		\P1_state_reg[0]/NET0131 ,
		_w1731_,
		_w2745_,
		_w2851_,
		_w2852_
	);
	LUT2 #(
		.INIT('he)
	) name2390 (
		_w2744_,
		_w2852_,
		_w2853_
	);
	LUT4 #(
		.INIT('hd070)
	) name2391 (
		\P1_state_reg[0]/NET0131 ,
		\P2_IR_reg[23]/NET0131 ,
		\P2_reg1_reg[27]/NET0131 ,
		_w1188_,
		_w2854_
	);
	LUT4 #(
		.INIT('h2000)
	) name2392 (
		\P2_reg1_reg[27]/NET0131 ,
		_w1189_,
		_w1352_,
		_w1356_,
		_w2855_
	);
	LUT4 #(
		.INIT('haa02)
	) name2393 (
		\P2_reg1_reg[27]/NET0131 ,
		_w1361_,
		_w1363_,
		_w1368_,
		_w2856_
	);
	LUT3 #(
		.INIT('h54)
	) name2394 (
		_w1506_,
		_w1609_,
		_w2856_,
		_w2857_
	);
	LUT4 #(
		.INIT('ha8aa)
	) name2395 (
		\P2_reg1_reg[27]/NET0131 ,
		_w1361_,
		_w1363_,
		_w1368_,
		_w2858_
	);
	LUT4 #(
		.INIT('h0c88)
	) name2396 (
		\P2_reg1_reg[27]/NET0131 ,
		_w1191_,
		_w1437_,
		_w1507_,
		_w2859_
	);
	LUT3 #(
		.INIT('ha2)
	) name2397 (
		\P2_reg1_reg[27]/NET0131 ,
		_w1684_,
		_w2469_,
		_w2860_
	);
	LUT4 #(
		.INIT('h00ef)
	) name2398 (
		_w546_,
		_w1078_,
		_w2471_,
		_w2860_,
		_w2861_
	);
	LUT2 #(
		.INIT('h4)
	) name2399 (
		_w2859_,
		_w2861_,
		_w2862_
	);
	LUT4 #(
		.INIT('h5600)
	) name2400 (
		_w1263_,
		_w1486_,
		_w1493_,
		_w1516_,
		_w2863_
	);
	LUT3 #(
		.INIT('h54)
	) name2401 (
		_w1575_,
		_w2856_,
		_w2863_,
		_w2864_
	);
	LUT3 #(
		.INIT('ha8)
	) name2402 (
		_w1530_,
		_w1599_,
		_w2858_,
		_w2865_
	);
	LUT4 #(
		.INIT('h0100)
	) name2403 (
		_w2857_,
		_w2864_,
		_w2865_,
		_w2862_,
		_w2866_
	);
	LUT4 #(
		.INIT('ha0a8)
	) name2404 (
		\P1_state_reg[0]/NET0131 ,
		_w1359_,
		_w2855_,
		_w2866_,
		_w2867_
	);
	LUT2 #(
		.INIT('he)
	) name2405 (
		_w2854_,
		_w2867_,
		_w2868_
	);
	LUT4 #(
		.INIT('hd070)
	) name2406 (
		\P1_state_reg[0]/NET0131 ,
		\P2_IR_reg[23]/NET0131 ,
		\P2_reg1_reg[28]/NET0131 ,
		_w1188_,
		_w2869_
	);
	LUT4 #(
		.INIT('h2000)
	) name2407 (
		\P2_reg1_reg[28]/NET0131 ,
		_w1189_,
		_w1352_,
		_w1356_,
		_w2870_
	);
	LUT4 #(
		.INIT('hc355)
	) name2408 (
		\P2_reg1_reg[28]/NET0131 ,
		_w1260_,
		_w1514_,
		_w1516_,
		_w2871_
	);
	LUT4 #(
		.INIT('h111d)
	) name2409 (
		\P2_reg1_reg[28]/NET0131 ,
		_w1507_,
		_w1517_,
		_w1520_,
		_w2872_
	);
	LUT4 #(
		.INIT('h1000)
	) name2410 (
		_w546_,
		_w1124_,
		_w1442_,
		_w1516_,
		_w2873_
	);
	LUT3 #(
		.INIT('ha2)
	) name2411 (
		\P2_reg1_reg[28]/NET0131 ,
		_w1684_,
		_w2469_,
		_w2874_
	);
	LUT2 #(
		.INIT('h1)
	) name2412 (
		_w2873_,
		_w2874_,
		_w2875_
	);
	LUT3 #(
		.INIT('hd0)
	) name2413 (
		_w1191_,
		_w2872_,
		_w2875_,
		_w2876_
	);
	LUT3 #(
		.INIT('he0)
	) name2414 (
		_w1506_,
		_w2871_,
		_w2876_,
		_w2877_
	);
	LUT4 #(
		.INIT('h35c5)
	) name2415 (
		\P2_reg1_reg[28]/NET0131 ,
		_w1260_,
		_w1516_,
		_w1573_,
		_w2878_
	);
	LUT4 #(
		.INIT('hc535)
	) name2416 (
		\P2_reg1_reg[28]/NET0131 ,
		_w1260_,
		_w1507_,
		_w1514_,
		_w2879_
	);
	LUT4 #(
		.INIT('hfc54)
	) name2417 (
		_w1530_,
		_w1575_,
		_w2878_,
		_w2879_,
		_w2880_
	);
	LUT4 #(
		.INIT('h3111)
	) name2418 (
		_w1359_,
		_w2870_,
		_w2877_,
		_w2880_,
		_w2881_
	);
	LUT3 #(
		.INIT('hce)
	) name2419 (
		\P1_state_reg[0]/NET0131 ,
		_w2869_,
		_w2881_,
		_w2882_
	);
	LUT4 #(
		.INIT('h1000)
	) name2420 (
		_w1734_,
		_w1735_,
		_w1737_,
		_w1739_,
		_w2883_
	);
	LUT2 #(
		.INIT('h2)
	) name2421 (
		\P1_reg0_reg[29]/NET0131 ,
		_w2883_,
		_w2884_
	);
	LUT4 #(
		.INIT('h30a0)
	) name2422 (
		\P1_reg0_reg[29]/NET0131 ,
		_w2281_,
		_w2292_,
		_w2883_,
		_w2885_
	);
	LUT4 #(
		.INIT('hc0a0)
	) name2423 (
		\P1_reg0_reg[29]/NET0131 ,
		_w2387_,
		_w2388_,
		_w2883_,
		_w2886_
	);
	LUT4 #(
		.INIT('h0355)
	) name2424 (
		\P1_reg0_reg[29]/NET0131 ,
		_w2390_,
		_w2422_,
		_w2883_,
		_w2887_
	);
	LUT4 #(
		.INIT('h9500)
	) name2425 (
		_w2273_,
		_w2443_,
		_w2444_,
		_w2883_,
		_w2888_
	);
	LUT2 #(
		.INIT('h2)
	) name2426 (
		\P1_reg0_reg[29]/NET0131 ,
		_w2524_,
		_w2889_
	);
	LUT4 #(
		.INIT('hfc55)
	) name2427 (
		\P1_reg0_reg[29]/NET0131 ,
		_w1748_,
		_w2272_,
		_w2883_,
		_w2890_
	);
	LUT3 #(
		.INIT('h31)
	) name2428 (
		_w2426_,
		_w2889_,
		_w2890_,
		_w2891_
	);
	LUT4 #(
		.INIT('h5700)
	) name2429 (
		_w2447_,
		_w2884_,
		_w2888_,
		_w2891_,
		_w2892_
	);
	LUT3 #(
		.INIT('hd0)
	) name2430 (
		_w2424_,
		_w2887_,
		_w2892_,
		_w2893_
	);
	LUT4 #(
		.INIT('ha8aa)
	) name2431 (
		_w1731_,
		_w2885_,
		_w2886_,
		_w2893_,
		_w2894_
	);
	LUT4 #(
		.INIT('h2000)
	) name2432 (
		\P1_reg0_reg[29]/NET0131 ,
		_w1723_,
		_w1727_,
		_w1730_,
		_w2895_
	);
	LUT2 #(
		.INIT('h2)
	) name2433 (
		\P1_reg0_reg[29]/NET0131 ,
		_w2462_,
		_w2896_
	);
	LUT4 #(
		.INIT('hffa8)
	) name2434 (
		\P1_state_reg[0]/NET0131 ,
		_w2894_,
		_w2895_,
		_w2896_,
		_w2897_
	);
	LUT4 #(
		.INIT('hd070)
	) name2435 (
		\P1_state_reg[0]/NET0131 ,
		\P2_IR_reg[23]/NET0131 ,
		\P2_reg2_reg[20]/NET0131 ,
		_w1188_,
		_w2898_
	);
	LUT4 #(
		.INIT('h2000)
	) name2436 (
		\P2_reg2_reg[20]/NET0131 ,
		_w1189_,
		_w1352_,
		_w1356_,
		_w2899_
	);
	LUT3 #(
		.INIT('h07)
	) name2437 (
		_w883_,
		_w888_,
		_w1435_,
		_w2900_
	);
	LUT4 #(
		.INIT('hbf00)
	) name2438 (
		_w845_,
		_w1423_,
		_w1426_,
		_w1435_,
		_w2901_
	);
	LUT4 #(
		.INIT('h020f)
	) name2439 (
		_w953_,
		_w2582_,
		_w2900_,
		_w2901_,
		_w2902_
	);
	LUT4 #(
		.INIT('h08c8)
	) name2440 (
		\P2_reg2_reg[20]/NET0131 ,
		_w1191_,
		_w1516_,
		_w2902_,
		_w2903_
	);
	LUT3 #(
		.INIT('h10)
	) name2441 (
		_w546_,
		_w962_,
		_w1522_,
		_w2904_
	);
	LUT3 #(
		.INIT('h40)
	) name2442 (
		_w963_,
		_w1229_,
		_w1232_,
		_w2905_
	);
	LUT4 #(
		.INIT('h0057)
	) name2443 (
		\P2_reg2_reg[20]/NET0131 ,
		_w1441_,
		_w1523_,
		_w2905_,
		_w2906_
	);
	LUT2 #(
		.INIT('h4)
	) name2444 (
		_w2904_,
		_w2906_,
		_w2907_
	);
	LUT2 #(
		.INIT('h4)
	) name2445 (
		_w2903_,
		_w2907_,
		_w2908_
	);
	LUT4 #(
		.INIT('h9a55)
	) name2446 (
		_w1289_,
		_w1508_,
		_w1509_,
		_w1510_,
		_w2909_
	);
	LUT4 #(
		.INIT('h0232)
	) name2447 (
		\P2_reg2_reg[20]/NET0131 ,
		_w1506_,
		_w1507_,
		_w2909_,
		_w2910_
	);
	LUT4 #(
		.INIT('h65aa)
	) name2448 (
		_w1289_,
		_w1544_,
		_w1550_,
		_w1558_,
		_w2911_
	);
	LUT4 #(
		.INIT('h020e)
	) name2449 (
		\P2_reg2_reg[20]/NET0131 ,
		_w1507_,
		_w1575_,
		_w2911_,
		_w2912_
	);
	LUT4 #(
		.INIT('h20e0)
	) name2450 (
		\P2_reg2_reg[20]/NET0131 ,
		_w1516_,
		_w1530_,
		_w2909_,
		_w2913_
	);
	LUT3 #(
		.INIT('h01)
	) name2451 (
		_w2912_,
		_w2913_,
		_w2910_,
		_w2914_
	);
	LUT4 #(
		.INIT('h3111)
	) name2452 (
		_w1359_,
		_w2899_,
		_w2908_,
		_w2914_,
		_w2915_
	);
	LUT3 #(
		.INIT('hce)
	) name2453 (
		\P1_state_reg[0]/NET0131 ,
		_w2898_,
		_w2915_,
		_w2916_
	);
	LUT2 #(
		.INIT('h8)
	) name2454 (
		_w1901_,
		_w2460_,
		_w2917_
	);
	LUT2 #(
		.INIT('h2)
	) name2455 (
		_w1901_,
		_w2644_,
		_w2918_
	);
	LUT4 #(
		.INIT('h1000)
	) name2456 (
		_w2212_,
		_w2223_,
		_w2404_,
		_w2406_,
		_w2919_
	);
	LUT4 #(
		.INIT('h0777)
	) name2457 (
		_w1972_,
		_w1974_,
		_w2244_,
		_w2245_,
		_w2920_
	);
	LUT2 #(
		.INIT('h8)
	) name2458 (
		_w2394_,
		_w2920_,
		_w2921_
	);
	LUT4 #(
		.INIT('h4000)
	) name2459 (
		_w1936_,
		_w2412_,
		_w2919_,
		_w2921_,
		_w2922_
	);
	LUT4 #(
		.INIT('h9555)
	) name2460 (
		_w1936_,
		_w2412_,
		_w2919_,
		_w2921_,
		_w2923_
	);
	LUT4 #(
		.INIT('h7020)
	) name2461 (
		_w1747_,
		_w1876_,
		_w2644_,
		_w2923_,
		_w2924_
	);
	LUT4 #(
		.INIT('h006f)
	) name2462 (
		_w1900_,
		_w2443_,
		_w2644_,
		_w2918_,
		_w2925_
	);
	LUT4 #(
		.INIT('ha0a8)
	) name2463 (
		_w1901_,
		_w2426_,
		_w2450_,
		_w2644_,
		_w2926_
	);
	LUT4 #(
		.INIT('h00fe)
	) name2464 (
		_w1748_,
		_w1899_,
		_w2689_,
		_w2926_,
		_w2927_
	);
	LUT3 #(
		.INIT('hd0)
	) name2465 (
		_w2447_,
		_w2925_,
		_w2927_,
		_w2928_
	);
	LUT4 #(
		.INIT('h5700)
	) name2466 (
		_w2424_,
		_w2918_,
		_w2924_,
		_w2928_,
		_w2929_
	);
	LUT3 #(
		.INIT('h1e)
	) name2467 (
		_w1748_,
		_w1899_,
		_w1904_,
		_w2930_
	);
	LUT2 #(
		.INIT('h8)
	) name2468 (
		_w2790_,
		_w2808_,
		_w2931_
	);
	LUT4 #(
		.INIT('hcc08)
	) name2469 (
		_w2310_,
		_w2314_,
		_w2792_,
		_w2793_,
		_w2932_
	);
	LUT4 #(
		.INIT('h0001)
	) name2470 (
		_w2311_,
		_w2321_,
		_w2322_,
		_w2328_,
		_w2933_
	);
	LUT3 #(
		.INIT('h0b)
	) name2471 (
		_w2798_,
		_w2800_,
		_w2803_,
		_w2934_
	);
	LUT4 #(
		.INIT('h1f00)
	) name2472 (
		_w2797_,
		_w2932_,
		_w2933_,
		_w2934_,
		_w2935_
	);
	LUT2 #(
		.INIT('h8)
	) name2473 (
		_w2801_,
		_w2809_,
		_w2936_
	);
	LUT3 #(
		.INIT('h07)
	) name2474 (
		_w2805_,
		_w2809_,
		_w2812_,
		_w2937_
	);
	LUT3 #(
		.INIT('h07)
	) name2475 (
		_w2790_,
		_w2814_,
		_w2817_,
		_w2938_
	);
	LUT3 #(
		.INIT('hd0)
	) name2476 (
		_w2931_,
		_w2937_,
		_w2938_,
		_w2939_
	);
	LUT4 #(
		.INIT('hdf00)
	) name2477 (
		_w2931_,
		_w2935_,
		_w2936_,
		_w2939_,
		_w2940_
	);
	LUT4 #(
		.INIT('h0001)
	) name2478 (
		_w2359_,
		_w2364_,
		_w2366_,
		_w2367_,
		_w2941_
	);
	LUT4 #(
		.INIT('h0001)
	) name2479 (
		_w2337_,
		_w2338_,
		_w2339_,
		_w2363_,
		_w2942_
	);
	LUT2 #(
		.INIT('h8)
	) name2480 (
		_w2941_,
		_w2942_,
		_w2943_
	);
	LUT3 #(
		.INIT('h70)
	) name2481 (
		_w2819_,
		_w2823_,
		_w2830_,
		_w2944_
	);
	LUT4 #(
		.INIT('h8f00)
	) name2482 (
		_w2819_,
		_w2823_,
		_w2830_,
		_w2941_,
		_w2945_
	);
	LUT3 #(
		.INIT('h07)
	) name2483 (
		_w2826_,
		_w2832_,
		_w2836_,
		_w2946_
	);
	LUT2 #(
		.INIT('h4)
	) name2484 (
		_w2945_,
		_w2946_,
		_w2947_
	);
	LUT4 #(
		.INIT('h9a55)
	) name2485 (
		_w2930_,
		_w2940_,
		_w2943_,
		_w2947_,
		_w2948_
	);
	LUT4 #(
		.INIT('h08c8)
	) name2486 (
		_w1901_,
		_w2388_,
		_w2644_,
		_w2948_,
		_w2949_
	);
	LUT2 #(
		.INIT('h8)
	) name2487 (
		_w2759_,
		_w2762_,
		_w2950_
	);
	LUT4 #(
		.INIT('h0001)
	) name2488 (
		_w2110_,
		_w2120_,
		_w2130_,
		_w2150_,
		_w2951_
	);
	LUT3 #(
		.INIT('h70)
	) name2489 (
		_w2751_,
		_w2753_,
		_w2756_,
		_w2952_
	);
	LUT4 #(
		.INIT('h1f00)
	) name2490 (
		_w2749_,
		_w2750_,
		_w2951_,
		_w2952_,
		_w2953_
	);
	LUT2 #(
		.INIT('h8)
	) name2491 (
		_w2754_,
		_w2760_,
		_w2954_
	);
	LUT3 #(
		.INIT('h0b)
	) name2492 (
		_w2757_,
		_w2760_,
		_w2766_,
		_w2955_
	);
	LUT3 #(
		.INIT('h70)
	) name2493 (
		_w2762_,
		_w2767_,
		_w2769_,
		_w2956_
	);
	LUT3 #(
		.INIT('hd0)
	) name2494 (
		_w2950_,
		_w2955_,
		_w2956_,
		_w2957_
	);
	LUT4 #(
		.INIT('hdf00)
	) name2495 (
		_w2950_,
		_w2953_,
		_w2954_,
		_w2957_,
		_w2958_
	);
	LUT4 #(
		.INIT('h0001)
	) name2496 (
		_w2165_,
		_w2177_,
		_w2202_,
		_w2263_,
		_w2959_
	);
	LUT4 #(
		.INIT('h0001)
	) name2497 (
		_w1878_,
		_w1954_,
		_w1964_,
		_w1978_,
		_w2960_
	);
	LUT2 #(
		.INIT('h8)
	) name2498 (
		_w2959_,
		_w2960_,
		_w2961_
	);
	LUT3 #(
		.INIT('h70)
	) name2499 (
		_w2771_,
		_w2774_,
		_w2779_,
		_w2962_
	);
	LUT4 #(
		.INIT('h8f00)
	) name2500 (
		_w2771_,
		_w2774_,
		_w2779_,
		_w2960_,
		_w2963_
	);
	LUT4 #(
		.INIT('h4504)
	) name2501 (
		_w1954_,
		_w1958_,
		_w1962_,
		_w1977_,
		_w2964_
	);
	LUT3 #(
		.INIT('h51)
	) name2502 (
		_w1878_,
		_w2782_,
		_w2964_,
		_w2965_
	);
	LUT2 #(
		.INIT('h1)
	) name2503 (
		_w2963_,
		_w2965_,
		_w2966_
	);
	LUT4 #(
		.INIT('h65aa)
	) name2504 (
		_w2930_,
		_w2958_,
		_w2961_,
		_w2966_,
		_w2967_
	);
	LUT4 #(
		.INIT('h08c8)
	) name2505 (
		_w1901_,
		_w2292_,
		_w2644_,
		_w2967_,
		_w2968_
	);
	LUT4 #(
		.INIT('ha8aa)
	) name2506 (
		_w1731_,
		_w2949_,
		_w2968_,
		_w2929_,
		_w2969_
	);
	LUT2 #(
		.INIT('h2)
	) name2507 (
		\P1_reg3_reg[26]/NET0131 ,
		\P1_state_reg[0]/NET0131 ,
		_w2970_
	);
	LUT4 #(
		.INIT('h6c00)
	) name2508 (
		\P1_reg3_reg[25]/NET0131 ,
		\P1_reg3_reg[26]/NET0131 ,
		_w1828_,
		_w2695_,
		_w2971_
	);
	LUT2 #(
		.INIT('h1)
	) name2509 (
		_w2970_,
		_w2971_,
		_w2972_
	);
	LUT4 #(
		.INIT('ha8ff)
	) name2510 (
		\P1_state_reg[0]/NET0131 ,
		_w2917_,
		_w2969_,
		_w2972_,
		_w2973_
	);
	LUT4 #(
		.INIT('h54ab)
	) name2511 (
		_w1748_,
		_w1941_,
		_w1947_,
		_w1952_,
		_w2974_
	);
	LUT4 #(
		.INIT('h20aa)
	) name2512 (
		_w2791_,
		_w2807_,
		_w2810_,
		_w2815_,
		_w2975_
	);
	LUT4 #(
		.INIT('h30b0)
	) name2513 (
		_w2820_,
		_w2825_,
		_w2833_,
		_w2975_,
		_w2976_
	);
	LUT4 #(
		.INIT('hd11d)
	) name2514 (
		\P1_reg2_reg[24]/NET0131 ,
		_w1741_,
		_w2974_,
		_w2976_,
		_w2977_
	);
	LUT2 #(
		.INIT('h2)
	) name2515 (
		_w2388_,
		_w2977_,
		_w2978_
	);
	LUT3 #(
		.INIT('h40)
	) name2516 (
		_w2752_,
		_w2755_,
		_w2764_,
		_w2979_
	);
	LUT4 #(
		.INIT('h40f0)
	) name2517 (
		_w2758_,
		_w2761_,
		_w2763_,
		_w2768_,
		_w2980_
	);
	LUT2 #(
		.INIT('h2)
	) name2518 (
		_w2772_,
		_w2980_,
		_w2981_
	);
	LUT4 #(
		.INIT('h4c44)
	) name2519 (
		_w2776_,
		_w2781_,
		_w2979_,
		_w2981_,
		_w2982_
	);
	LUT4 #(
		.INIT('h1dd1)
	) name2520 (
		\P1_reg2_reg[24]/NET0131 ,
		_w1741_,
		_w2974_,
		_w2982_,
		_w2983_
	);
	LUT4 #(
		.INIT('h0777)
	) name2521 (
		_w1960_,
		_w1961_,
		_w1972_,
		_w1974_,
		_w2984_
	);
	LUT4 #(
		.INIT('h8000)
	) name2522 (
		_w2394_,
		_w2404_,
		_w2408_,
		_w2984_,
		_w2985_
	);
	LUT4 #(
		.INIT('h4144)
	) name2523 (
		_w1747_,
		_w1876_,
		_w1952_,
		_w2985_,
		_w2986_
	);
	LUT3 #(
		.INIT('h80)
	) name2524 (
		_w1747_,
		_w1960_,
		_w1961_,
		_w2987_
	);
	LUT4 #(
		.INIT('hddd1)
	) name2525 (
		\P1_reg2_reg[24]/NET0131 ,
		_w1741_,
		_w2986_,
		_w2987_,
		_w2988_
	);
	LUT4 #(
		.INIT('h5400)
	) name2526 (
		_w1748_,
		_w1941_,
		_w1947_,
		_w2426_,
		_w2989_
	);
	LUT4 #(
		.INIT('h4000)
	) name2527 (
		_w1958_,
		_w2436_,
		_w2438_,
		_w2439_,
		_w2990_
	);
	LUT4 #(
		.INIT('h070b)
	) name2528 (
		_w1948_,
		_w2447_,
		_w2989_,
		_w2990_,
		_w2991_
	);
	LUT4 #(
		.INIT('ha2a0)
	) name2529 (
		\P1_reg2_reg[24]/NET0131 ,
		_w1741_,
		_w2450_,
		_w2452_,
		_w2992_
	);
	LUT4 #(
		.INIT('h0008)
	) name2530 (
		_w1950_,
		_w2284_,
		_w2288_,
		_w2291_,
		_w2993_
	);
	LUT2 #(
		.INIT('h1)
	) name2531 (
		_w2992_,
		_w2993_,
		_w2994_
	);
	LUT3 #(
		.INIT('hd0)
	) name2532 (
		_w1741_,
		_w2991_,
		_w2994_,
		_w2995_
	);
	LUT3 #(
		.INIT('hd0)
	) name2533 (
		_w2424_,
		_w2988_,
		_w2995_,
		_w2996_
	);
	LUT3 #(
		.INIT('hd0)
	) name2534 (
		_w2292_,
		_w2983_,
		_w2996_,
		_w2997_
	);
	LUT4 #(
		.INIT('h2000)
	) name2535 (
		\P1_reg2_reg[24]/NET0131 ,
		_w1723_,
		_w1727_,
		_w1730_,
		_w2998_
	);
	LUT4 #(
		.INIT('h0075)
	) name2536 (
		_w1731_,
		_w2978_,
		_w2997_,
		_w2998_,
		_w2999_
	);
	LUT2 #(
		.INIT('h2)
	) name2537 (
		\P1_reg2_reg[24]/NET0131 ,
		_w2462_,
		_w3000_
	);
	LUT3 #(
		.INIT('hf2)
	) name2538 (
		\P1_state_reg[0]/NET0131 ,
		_w2999_,
		_w3000_,
		_w3001_
	);
	LUT2 #(
		.INIT('h2)
	) name2539 (
		\P1_reg2_reg[25]/NET0131 ,
		_w2462_,
		_w3002_
	);
	LUT4 #(
		.INIT('h2000)
	) name2540 (
		\P1_reg2_reg[25]/NET0131 ,
		_w1723_,
		_w1727_,
		_w1730_,
		_w3003_
	);
	LUT2 #(
		.INIT('h2)
	) name2541 (
		\P1_reg2_reg[25]/NET0131 ,
		_w1741_,
		_w3004_
	);
	LUT4 #(
		.INIT('hc9cc)
	) name2542 (
		_w1876_,
		_w1904_,
		_w1952_,
		_w2985_,
		_w3005_
	);
	LUT4 #(
		.INIT('h082a)
	) name2543 (
		_w1741_,
		_w1747_,
		_w1952_,
		_w3005_,
		_w3006_
	);
	LUT3 #(
		.INIT('ha8)
	) name2544 (
		_w2424_,
		_w3004_,
		_w3006_,
		_w3007_
	);
	LUT4 #(
		.INIT('h0705)
	) name2545 (
		_w1871_,
		_w1948_,
		_w2443_,
		_w2990_,
		_w3008_
	);
	LUT4 #(
		.INIT('he020)
	) name2546 (
		\P1_reg2_reg[25]/NET0131 ,
		_w1741_,
		_w2447_,
		_w3008_,
		_w3009_
	);
	LUT4 #(
		.INIT('h5400)
	) name2547 (
		_w1748_,
		_w1839_,
		_w1870_,
		_w2426_,
		_w3010_
	);
	LUT4 #(
		.INIT('haa20)
	) name2548 (
		\P1_reg2_reg[25]/NET0131 ,
		_w1741_,
		_w2426_,
		_w2450_,
		_w3011_
	);
	LUT4 #(
		.INIT('h0008)
	) name2549 (
		_w1872_,
		_w2284_,
		_w2288_,
		_w2291_,
		_w3012_
	);
	LUT4 #(
		.INIT('h0103)
	) name2550 (
		_w1741_,
		_w3011_,
		_w3012_,
		_w3010_,
		_w3013_
	);
	LUT2 #(
		.INIT('h4)
	) name2551 (
		_w3009_,
		_w3013_,
		_w3014_
	);
	LUT2 #(
		.INIT('h4)
	) name2552 (
		_w3007_,
		_w3014_,
		_w3015_
	);
	LUT4 #(
		.INIT('h54ab)
	) name2553 (
		_w1748_,
		_w1839_,
		_w1870_,
		_w1876_,
		_w3016_
	);
	LUT4 #(
		.INIT('h40cc)
	) name2554 (
		_w2049_,
		_w2204_,
		_w2249_,
		_w2253_,
		_w3017_
	);
	LUT4 #(
		.INIT('h0070)
	) name2555 (
		_w2153_,
		_w2250_,
		_w2260_,
		_w3017_,
		_w3018_
	);
	LUT4 #(
		.INIT('h5ad2)
	) name2556 (
		_w1994_,
		_w2265_,
		_w3016_,
		_w3018_,
		_w3019_
	);
	LUT4 #(
		.INIT('h20e0)
	) name2557 (
		\P1_reg2_reg[25]/NET0131 ,
		_w1741_,
		_w2292_,
		_w3019_,
		_w3020_
	);
	LUT2 #(
		.INIT('h8)
	) name2558 (
		_w2351_,
		_w2353_,
		_w3021_
	);
	LUT3 #(
		.INIT('h40)
	) name2559 (
		_w2327_,
		_w2330_,
		_w3021_,
		_w3022_
	);
	LUT4 #(
		.INIT('h7030)
	) name2560 (
		_w2301_,
		_w2336_,
		_w2351_,
		_w2353_,
		_w3023_
	);
	LUT2 #(
		.INIT('h2)
	) name2561 (
		_w2347_,
		_w3023_,
		_w3024_
	);
	LUT4 #(
		.INIT('h4c44)
	) name2562 (
		_w2369_,
		_w2378_,
		_w3022_,
		_w3024_,
		_w3025_
	);
	LUT4 #(
		.INIT('hd11d)
	) name2563 (
		\P1_reg2_reg[25]/NET0131 ,
		_w1741_,
		_w3016_,
		_w3025_,
		_w3026_
	);
	LUT3 #(
		.INIT('h31)
	) name2564 (
		_w2388_,
		_w3020_,
		_w3026_,
		_w3027_
	);
	LUT4 #(
		.INIT('h3111)
	) name2565 (
		_w1731_,
		_w3003_,
		_w3015_,
		_w3027_,
		_w3028_
	);
	LUT3 #(
		.INIT('hce)
	) name2566 (
		\P1_state_reg[0]/NET0131 ,
		_w3002_,
		_w3028_,
		_w3029_
	);
	LUT4 #(
		.INIT('hd070)
	) name2567 (
		\P1_state_reg[0]/NET0131 ,
		\P2_IR_reg[23]/NET0131 ,
		\P2_reg2_reg[17]/NET0131 ,
		_w1188_,
		_w3030_
	);
	LUT4 #(
		.INIT('h2000)
	) name2568 (
		\P2_reg2_reg[17]/NET0131 ,
		_w1189_,
		_w1352_,
		_w1356_,
		_w3031_
	);
	LUT4 #(
		.INIT('ha8aa)
	) name2569 (
		\P2_reg2_reg[17]/NET0131 ,
		_w1361_,
		_w1363_,
		_w1368_,
		_w3032_
	);
	LUT4 #(
		.INIT('h0e02)
	) name2570 (
		\P2_reg2_reg[17]/NET0131 ,
		_w1507_,
		_w1575_,
		_w2593_,
		_w3033_
	);
	LUT4 #(
		.INIT('haa02)
	) name2571 (
		\P2_reg2_reg[17]/NET0131 ,
		_w1361_,
		_w1363_,
		_w1368_,
		_w3034_
	);
	LUT4 #(
		.INIT('h111d)
	) name2572 (
		\P2_reg2_reg[17]/NET0131 ,
		_w1516_,
		_w2596_,
		_w2597_,
		_w3035_
	);
	LUT3 #(
		.INIT('h40)
	) name2573 (
		_w860_,
		_w1442_,
		_w1507_,
		_w3036_
	);
	LUT3 #(
		.INIT('h40)
	) name2574 (
		_w842_,
		_w1229_,
		_w1232_,
		_w3037_
	);
	LUT4 #(
		.INIT('h0057)
	) name2575 (
		\P2_reg2_reg[17]/NET0131 ,
		_w1441_,
		_w1523_,
		_w3037_,
		_w3038_
	);
	LUT2 #(
		.INIT('h4)
	) name2576 (
		_w3036_,
		_w3038_,
		_w3039_
	);
	LUT3 #(
		.INIT('hd0)
	) name2577 (
		_w1191_,
		_w3035_,
		_w3039_,
		_w3040_
	);
	LUT4 #(
		.INIT('h4484)
	) name2578 (
		_w1314_,
		_w1516_,
		_w1665_,
		_w2604_,
		_w3041_
	);
	LUT3 #(
		.INIT('ha8)
	) name2579 (
		_w1530_,
		_w3034_,
		_w3041_,
		_w3042_
	);
	LUT4 #(
		.INIT('h4484)
	) name2580 (
		_w1314_,
		_w1507_,
		_w1665_,
		_w2604_,
		_w3043_
	);
	LUT3 #(
		.INIT('h54)
	) name2581 (
		_w1506_,
		_w3032_,
		_w3043_,
		_w3044_
	);
	LUT4 #(
		.INIT('h0100)
	) name2582 (
		_w3033_,
		_w3042_,
		_w3044_,
		_w3040_,
		_w3045_
	);
	LUT4 #(
		.INIT('ha0a8)
	) name2583 (
		\P1_state_reg[0]/NET0131 ,
		_w1359_,
		_w3031_,
		_w3045_,
		_w3046_
	);
	LUT2 #(
		.INIT('he)
	) name2584 (
		_w3030_,
		_w3046_,
		_w3047_
	);
	LUT4 #(
		.INIT('hd070)
	) name2585 (
		\P1_state_reg[0]/NET0131 ,
		\P2_IR_reg[23]/NET0131 ,
		\P2_reg2_reg[18]/NET0131 ,
		_w1188_,
		_w3048_
	);
	LUT4 #(
		.INIT('h2000)
	) name2586 (
		\P2_reg2_reg[18]/NET0131 ,
		_w1189_,
		_w1352_,
		_w1356_,
		_w3049_
	);
	LUT4 #(
		.INIT('h08c8)
	) name2587 (
		\P2_reg2_reg[18]/NET0131 ,
		_w1191_,
		_w1516_,
		_w2564_,
		_w3050_
	);
	LUT3 #(
		.INIT('h40)
	) name2588 (
		_w925_,
		_w1442_,
		_w1507_,
		_w3051_
	);
	LUT3 #(
		.INIT('h40)
	) name2589 (
		_w907_,
		_w1229_,
		_w1232_,
		_w3052_
	);
	LUT4 #(
		.INIT('h0057)
	) name2590 (
		\P2_reg2_reg[18]/NET0131 ,
		_w1441_,
		_w1523_,
		_w3052_,
		_w3053_
	);
	LUT2 #(
		.INIT('h4)
	) name2591 (
		_w3051_,
		_w3053_,
		_w3054_
	);
	LUT2 #(
		.INIT('h4)
	) name2592 (
		_w3050_,
		_w3054_,
		_w3055_
	);
	LUT4 #(
		.INIT('h20e0)
	) name2593 (
		\P2_reg2_reg[18]/NET0131 ,
		_w1516_,
		_w1530_,
		_w2558_,
		_w3056_
	);
	LUT4 #(
		.INIT('h0e02)
	) name2594 (
		\P2_reg2_reg[18]/NET0131 ,
		_w1507_,
		_w1575_,
		_w2543_,
		_w3057_
	);
	LUT4 #(
		.INIT('h0232)
	) name2595 (
		\P2_reg2_reg[18]/NET0131 ,
		_w1506_,
		_w1507_,
		_w2558_,
		_w3058_
	);
	LUT3 #(
		.INIT('h01)
	) name2596 (
		_w3057_,
		_w3058_,
		_w3056_,
		_w3059_
	);
	LUT4 #(
		.INIT('h3111)
	) name2597 (
		_w1359_,
		_w3049_,
		_w3055_,
		_w3059_,
		_w3060_
	);
	LUT3 #(
		.INIT('hce)
	) name2598 (
		\P1_state_reg[0]/NET0131 ,
		_w3048_,
		_w3060_,
		_w3061_
	);
	LUT4 #(
		.INIT('hd070)
	) name2599 (
		\P1_state_reg[0]/NET0131 ,
		\P2_IR_reg[23]/NET0131 ,
		\P2_reg2_reg[19]/NET0131 ,
		_w1188_,
		_w3062_
	);
	LUT4 #(
		.INIT('h2000)
	) name2600 (
		\P2_reg2_reg[19]/NET0131 ,
		_w1189_,
		_w1352_,
		_w1356_,
		_w3063_
	);
	LUT4 #(
		.INIT('haa02)
	) name2601 (
		\P2_reg2_reg[19]/NET0131 ,
		_w1361_,
		_w1363_,
		_w1368_,
		_w3064_
	);
	LUT4 #(
		.INIT('h111d)
	) name2602 (
		\P2_reg2_reg[19]/NET0131 ,
		_w1516_,
		_w2581_,
		_w2583_,
		_w3065_
	);
	LUT4 #(
		.INIT('hf100)
	) name2603 (
		_w546_,
		_w899_,
		_w901_,
		_w1442_,
		_w3066_
	);
	LUT3 #(
		.INIT('h40)
	) name2604 (
		_w886_,
		_w1229_,
		_w1232_,
		_w3067_
	);
	LUT4 #(
		.INIT('h0057)
	) name2605 (
		\P2_reg2_reg[19]/NET0131 ,
		_w1441_,
		_w1523_,
		_w3067_,
		_w3068_
	);
	LUT3 #(
		.INIT('h70)
	) name2606 (
		_w1507_,
		_w3066_,
		_w3068_,
		_w3069_
	);
	LUT3 #(
		.INIT('hd0)
	) name2607 (
		_w1191_,
		_w3065_,
		_w3069_,
		_w3070_
	);
	LUT4 #(
		.INIT('ha8aa)
	) name2608 (
		\P2_reg2_reg[19]/NET0131 ,
		_w1361_,
		_w1363_,
		_w1368_,
		_w3071_
	);
	LUT4 #(
		.INIT('h020e)
	) name2609 (
		\P2_reg2_reg[19]/NET0131 ,
		_w1507_,
		_w1575_,
		_w2573_,
		_w3072_
	);
	LUT4 #(
		.INIT('h6500)
	) name2610 (
		_w1272_,
		_w1387_,
		_w1394_,
		_w1516_,
		_w3073_
	);
	LUT3 #(
		.INIT('ha8)
	) name2611 (
		_w1530_,
		_w3064_,
		_w3073_,
		_w3074_
	);
	LUT4 #(
		.INIT('h6500)
	) name2612 (
		_w1272_,
		_w1387_,
		_w1394_,
		_w1507_,
		_w3075_
	);
	LUT3 #(
		.INIT('h54)
	) name2613 (
		_w1506_,
		_w3071_,
		_w3075_,
		_w3076_
	);
	LUT3 #(
		.INIT('h01)
	) name2614 (
		_w3074_,
		_w3076_,
		_w3072_,
		_w3077_
	);
	LUT4 #(
		.INIT('h3111)
	) name2615 (
		_w1359_,
		_w3063_,
		_w3070_,
		_w3077_,
		_w3078_
	);
	LUT3 #(
		.INIT('hce)
	) name2616 (
		\P1_state_reg[0]/NET0131 ,
		_w3062_,
		_w3078_,
		_w3079_
	);
	LUT4 #(
		.INIT('h1000)
	) name2617 (
		_w963_,
		_w1189_,
		_w1352_,
		_w1356_,
		_w3080_
	);
	LUT4 #(
		.INIT('h04c4)
	) name2618 (
		_w963_,
		_w1447_,
		_w1411_,
		_w2911_,
		_w3081_
	);
	LUT4 #(
		.INIT('h0010)
	) name2619 (
		_w546_,
		_w962_,
		_w1232_,
		_w1439_,
		_w3082_
	);
	LUT3 #(
		.INIT('h54)
	) name2620 (
		_w963_,
		_w1441_,
		_w1443_,
		_w3083_
	);
	LUT2 #(
		.INIT('h1)
	) name2621 (
		_w3082_,
		_w3083_,
		_w3084_
	);
	LUT2 #(
		.INIT('h4)
	) name2622 (
		_w3081_,
		_w3084_,
		_w3085_
	);
	LUT4 #(
		.INIT('h04c4)
	) name2623 (
		_w963_,
		_w1191_,
		_w1411_,
		_w2902_,
		_w3086_
	);
	LUT4 #(
		.INIT('h010d)
	) name2624 (
		_w963_,
		_w1369_,
		_w1496_,
		_w2911_,
		_w3087_
	);
	LUT4 #(
		.INIT('h010d)
	) name2625 (
		_w963_,
		_w1369_,
		_w1409_,
		_w2909_,
		_w3088_
	);
	LUT3 #(
		.INIT('h01)
	) name2626 (
		_w3087_,
		_w3088_,
		_w3086_,
		_w3089_
	);
	LUT4 #(
		.INIT('h3111)
	) name2627 (
		_w1359_,
		_w3080_,
		_w3085_,
		_w3089_,
		_w3090_
	);
	LUT2 #(
		.INIT('h4)
	) name2628 (
		\P1_state_reg[0]/NET0131 ,
		\P2_reg3_reg[20]/NET0131 ,
		_w3091_
	);
	LUT3 #(
		.INIT('h0b)
	) name2629 (
		_w963_,
		_w1349_,
		_w3091_,
		_w3092_
	);
	LUT3 #(
		.INIT('h2f)
	) name2630 (
		\P1_state_reg[0]/NET0131 ,
		_w3090_,
		_w3092_,
		_w3093_
	);
	LUT4 #(
		.INIT('h8828)
	) name2631 (
		\P1_B_reg/NET0131 ,
		\P1_IR_reg[23]/NET0131 ,
		\P1_IR_reg[31]/NET0131 ,
		_w1722_,
		_w3094_
	);
	LUT4 #(
		.INIT('h0323)
	) name2632 (
		_w2332_,
		_w2334_,
		_w2808_,
		_w2809_,
		_w3095_
	);
	LUT4 #(
		.INIT('h0e08)
	) name2633 (
		_w2040_,
		_w2044_,
		_w2297_,
		_w2321_,
		_w3096_
	);
	LUT3 #(
		.INIT('h51)
	) name2634 (
		_w2299_,
		_w2801_,
		_w3096_,
		_w3097_
	);
	LUT3 #(
		.INIT('ha8)
	) name2635 (
		_w2815_,
		_w3095_,
		_w3097_,
		_w3098_
	);
	LUT3 #(
		.INIT('h70)
	) name2636 (
		_w2084_,
		_w2085_,
		_w2089_,
		_w3099_
	);
	LUT4 #(
		.INIT('h020b)
	) name2637 (
		_w2077_,
		_w2081_,
		_w2306_,
		_w3099_,
		_w3100_
	);
	LUT4 #(
		.INIT('h50d0)
	) name2638 (
		_w2304_,
		_w2310_,
		_w2314_,
		_w3100_,
		_w3101_
	);
	LUT3 #(
		.INIT('h01)
	) name2639 (
		_w2296_,
		_w2324_,
		_w2325_,
		_w3102_
	);
	LUT4 #(
		.INIT('h8000)
	) name2640 (
		_w2804_,
		_w2811_,
		_w2813_,
		_w3102_,
		_w3103_
	);
	LUT4 #(
		.INIT('h3b00)
	) name2641 (
		_w2319_,
		_w2794_,
		_w3101_,
		_w3103_,
		_w3104_
	);
	LUT3 #(
		.INIT('h01)
	) name2642 (
		_w2344_,
		_w2345_,
		_w2373_,
		_w3105_
	);
	LUT2 #(
		.INIT('h4)
	) name2643 (
		_w2340_,
		_w2816_,
		_w3106_
	);
	LUT3 #(
		.INIT('h80)
	) name2644 (
		_w2831_,
		_w3105_,
		_w3106_,
		_w3107_
	);
	LUT3 #(
		.INIT('he0)
	) name2645 (
		_w3098_,
		_w3104_,
		_w3107_,
		_w3108_
	);
	LUT4 #(
		.INIT('h00e8)
	) name2646 (
		_w1983_,
		_w1987_,
		_w2337_,
		_w2372_,
		_w3109_
	);
	LUT3 #(
		.INIT('h51)
	) name2647 (
		_w2376_,
		_w2824_,
		_w3109_,
		_w3110_
	);
	LUT4 #(
		.INIT('h1101)
	) name2648 (
		_w2338_,
		_w2339_,
		_w2341_,
		_w2790_,
		_w3111_
	);
	LUT3 #(
		.INIT('h20)
	) name2649 (
		_w2831_,
		_w3111_,
		_w3105_,
		_w3112_
	);
	LUT2 #(
		.INIT('h1)
	) name2650 (
		_w3110_,
		_w3112_,
		_w3113_
	);
	LUT2 #(
		.INIT('h8)
	) name2651 (
		_w2834_,
		_w2835_,
		_w3114_
	);
	LUT4 #(
		.INIT('h0233)
	) name2652 (
		_w2380_,
		_w2383_,
		_w2826_,
		_w2827_,
		_w3115_
	);
	LUT4 #(
		.INIT('h004f)
	) name2653 (
		_w3108_,
		_w3113_,
		_w3114_,
		_w3115_,
		_w3116_
	);
	LUT2 #(
		.INIT('h1)
	) name2654 (
		\P2_datao_reg[30]/NET0131 ,
		\si[30]_pad ,
		_w3117_
	);
	LUT4 #(
		.INIT('hfac8)
	) name2655 (
		\P2_datao_reg[28]/NET0131 ,
		\P2_datao_reg[29]/NET0131 ,
		\si[28]_pad ,
		\si[29]_pad ,
		_w3118_
	);
	LUT3 #(
		.INIT('h10)
	) name2656 (
		_w1803_,
		_w3117_,
		_w3118_,
		_w3119_
	);
	LUT2 #(
		.INIT('h8)
	) name2657 (
		_w1911_,
		_w3119_,
		_w3120_
	);
	LUT2 #(
		.INIT('h8)
	) name2658 (
		\P2_datao_reg[30]/NET0131 ,
		\si[30]_pad ,
		_w3121_
	);
	LUT4 #(
		.INIT('h0b0a)
	) name2659 (
		_w2267_,
		_w2268_,
		_w3117_,
		_w3118_,
		_w3122_
	);
	LUT4 #(
		.INIT('h0023)
	) name2660 (
		_w1910_,
		_w3121_,
		_w3119_,
		_w3122_,
		_w3123_
	);
	LUT3 #(
		.INIT('hb0)
	) name2661 (
		_w1956_,
		_w3120_,
		_w3123_,
		_w3124_
	);
	LUT4 #(
		.INIT('ha6a9)
	) name2662 (
		\P2_datao_reg[31]/NET0131 ,
		\si[31]_pad ,
		_w547_,
		_w3124_,
		_w3125_
	);
	LUT2 #(
		.INIT('h4)
	) name2663 (
		_w1748_,
		_w3125_,
		_w3126_
	);
	LUT3 #(
		.INIT('h40)
	) name2664 (
		_w1748_,
		_w2397_,
		_w3125_,
		_w3127_
	);
	LUT3 #(
		.INIT('h10)
	) name2665 (
		_w1796_,
		_w1803_,
		_w3118_,
		_w3128_
	);
	LUT2 #(
		.INIT('h8)
	) name2666 (
		_w1896_,
		_w3128_,
		_w3129_
	);
	LUT4 #(
		.INIT('h137f)
	) name2667 (
		\P2_datao_reg[28]/NET0131 ,
		\P2_datao_reg[29]/NET0131 ,
		\si[28]_pad ,
		\si[29]_pad ,
		_w3130_
	);
	LUT4 #(
		.INIT('hef00)
	) name2668 (
		_w1803_,
		_w1810_,
		_w3118_,
		_w3130_,
		_w3131_
	);
	LUT3 #(
		.INIT('hb0)
	) name2669 (
		_w1897_,
		_w3128_,
		_w3131_,
		_w3132_
	);
	LUT4 #(
		.INIT('h1f00)
	) name2670 (
		_w1893_,
		_w1969_,
		_w3129_,
		_w3132_,
		_w3133_
	);
	LUT4 #(
		.INIT('h5956)
	) name2671 (
		\P2_datao_reg[30]/NET0131 ,
		\si[30]_pad ,
		_w547_,
		_w3133_,
		_w3134_
	);
	LUT2 #(
		.INIT('h1)
	) name2672 (
		_w1748_,
		_w3134_,
		_w3135_
	);
	LUT3 #(
		.INIT('h32)
	) name2673 (
		_w1748_,
		_w2419_,
		_w3134_,
		_w3136_
	);
	LUT2 #(
		.INIT('h1)
	) name2674 (
		_w3127_,
		_w3136_,
		_w3137_
	);
	LUT4 #(
		.INIT('h0001)
	) name2675 (
		_w2279_,
		_w2382_,
		_w3127_,
		_w3136_,
		_w3138_
	);
	LUT3 #(
		.INIT('h23)
	) name2676 (
		_w1748_,
		_w2397_,
		_w3125_,
		_w3139_
	);
	LUT3 #(
		.INIT('h04)
	) name2677 (
		_w1748_,
		_w2419_,
		_w3134_,
		_w3140_
	);
	LUT2 #(
		.INIT('h1)
	) name2678 (
		_w3139_,
		_w3140_,
		_w3141_
	);
	LUT4 #(
		.INIT('h00e8)
	) name2679 (
		_w2273_,
		_w2276_,
		_w2357_,
		_w3136_,
		_w3142_
	);
	LUT3 #(
		.INIT('h51)
	) name2680 (
		_w3127_,
		_w3141_,
		_w3142_,
		_w3143_
	);
	LUT4 #(
		.INIT('h5510)
	) name2681 (
		_w3094_,
		_w3116_,
		_w3138_,
		_w3143_,
		_w3144_
	);
	LUT4 #(
		.INIT('h0045)
	) name2682 (
		_w3094_,
		_w3116_,
		_w3138_,
		_w3143_,
		_w3145_
	);
	LUT4 #(
		.INIT('hfeba)
	) name2683 (
		_w2288_,
		_w2291_,
		_w3144_,
		_w3145_,
		_w3146_
	);
	LUT4 #(
		.INIT('h0001)
	) name2684 (
		_w2278_,
		_w2357_,
		_w3139_,
		_w3140_,
		_w3147_
	);
	LUT3 #(
		.INIT('he0)
	) name2685 (
		_w2818_,
		_w2819_,
		_w2825_,
		_w3148_
	);
	LUT4 #(
		.INIT('h050d)
	) name2686 (
		_w2828_,
		_w2833_,
		_w2837_,
		_w3148_,
		_w3149_
	);
	LUT2 #(
		.INIT('h2)
	) name2687 (
		_w3147_,
		_w3149_,
		_w3150_
	);
	LUT3 #(
		.INIT('h54)
	) name2688 (
		_w2278_,
		_w2279_,
		_w2382_,
		_w3151_
	);
	LUT4 #(
		.INIT('h0071)
	) name2689 (
		_w2273_,
		_w2276_,
		_w2382_,
		_w3140_,
		_w3152_
	);
	LUT3 #(
		.INIT('h31)
	) name2690 (
		_w3137_,
		_w3139_,
		_w3152_,
		_w3153_
	);
	LUT2 #(
		.INIT('h8)
	) name2691 (
		_w2829_,
		_w3147_,
		_w3154_
	);
	LUT3 #(
		.INIT('h13)
	) name2692 (
		_w2975_,
		_w3153_,
		_w3154_,
		_w3155_
	);
	LUT4 #(
		.INIT('h1311)
	) name2693 (
		_w2451_,
		_w3094_,
		_w3150_,
		_w3155_,
		_w3156_
	);
	LUT2 #(
		.INIT('h4)
	) name2694 (
		_w2282_,
		_w2449_,
		_w3157_
	);
	LUT3 #(
		.INIT('h02)
	) name2695 (
		_w2280_,
		_w3127_,
		_w3136_,
		_w3158_
	);
	LUT2 #(
		.INIT('h8)
	) name2696 (
		_w3141_,
		_w3158_,
		_w3159_
	);
	LUT3 #(
		.INIT('h1e)
	) name2697 (
		_w1748_,
		_w1982_,
		_w1987_,
		_w3160_
	);
	LUT3 #(
		.INIT('h1e)
	) name2698 (
		_w1748_,
		_w1957_,
		_w1962_,
		_w3161_
	);
	LUT3 #(
		.INIT('h1e)
	) name2699 (
		_w1748_,
		_w2154_,
		_w2163_,
		_w3162_
	);
	LUT3 #(
		.INIT('h01)
	) name2700 (
		_w3161_,
		_w3162_,
		_w3160_,
		_w3163_
	);
	LUT3 #(
		.INIT('h10)
	) name2701 (
		_w2788_,
		_w2930_,
		_w3163_,
		_w3164_
	);
	LUT4 #(
		.INIT('hdc23)
	) name2702 (
		_w1748_,
		_w2168_,
		_w2170_,
		_w2175_,
		_w3165_
	);
	LUT4 #(
		.INIT('h54ab)
	) name2703 (
		_w1748_,
		_w1966_,
		_w1970_,
		_w1975_,
		_w3166_
	);
	LUT3 #(
		.INIT('h10)
	) name2704 (
		_w3016_,
		_w3166_,
		_w3165_,
		_w3167_
	);
	LUT2 #(
		.INIT('h9)
	) name2705 (
		_w2231_,
		_w2235_,
		_w3168_
	);
	LUT2 #(
		.INIT('h9)
	) name2706 (
		_w2242_,
		_w2246_,
		_w3169_
	);
	LUT2 #(
		.INIT('h9)
	) name2707 (
		_w2183_,
		_w2187_,
		_w3170_
	);
	LUT4 #(
		.INIT('h0660)
	) name2708 (
		_w2183_,
		_w2187_,
		_w2242_,
		_w2246_,
		_w3171_
	);
	LUT2 #(
		.INIT('h4)
	) name2709 (
		_w3168_,
		_w3171_,
		_w3172_
	);
	LUT2 #(
		.INIT('h9)
	) name2710 (
		_w2016_,
		_w2020_,
		_w3173_
	);
	LUT2 #(
		.INIT('h9)
	) name2711 (
		_w2208_,
		_w2212_,
		_w3174_
	);
	LUT4 #(
		.INIT('h1eee)
	) name2712 (
		_w2099_,
		_w2103_,
		_w2105_,
		_w2107_,
		_w3175_
	);
	LUT4 #(
		.INIT('h1eee)
	) name2713 (
		_w2024_,
		_w2028_,
		_w2030_,
		_w2033_,
		_w3176_
	);
	LUT3 #(
		.INIT('h87)
	) name2714 (
		_w2084_,
		_w2085_,
		_w2089_,
		_w3177_
	);
	LUT3 #(
		.INIT('h87)
	) name2715 (
		_w2051_,
		_w2052_,
		_w2057_,
		_w3178_
	);
	LUT4 #(
		.INIT('h0040)
	) name2716 (
		_w3176_,
		_w3177_,
		_w3178_,
		_w3175_,
		_w3179_
	);
	LUT3 #(
		.INIT('h10)
	) name2717 (
		_w3174_,
		_w3173_,
		_w3179_,
		_w3180_
	);
	LUT2 #(
		.INIT('h9)
	) name2718 (
		_w2196_,
		_w2200_,
		_w3181_
	);
	LUT3 #(
		.INIT('h6a)
	) name2719 (
		_w2124_,
		_w2125_,
		_w2127_,
		_w3182_
	);
	LUT3 #(
		.INIT('h95)
	) name2720 (
		_w2114_,
		_w2116_,
		_w2117_,
		_w3183_
	);
	LUT3 #(
		.INIT('h87)
	) name2721 (
		_w2059_,
		_w2060_,
		_w2065_,
		_w3184_
	);
	LUT3 #(
		.INIT('h04)
	) name2722 (
		_w3183_,
		_w3184_,
		_w3182_,
		_w3185_
	);
	LUT3 #(
		.INIT('h6a)
	) name2723 (
		_w2040_,
		_w2041_,
		_w2043_,
		_w3186_
	);
	LUT3 #(
		.INIT('h6a)
	) name2724 (
		_w2134_,
		_w2135_,
		_w2137_,
		_w3187_
	);
	LUT3 #(
		.INIT('h78)
	) name2725 (
		_w489_,
		_w491_,
		_w2071_,
		_w3188_
	);
	LUT3 #(
		.INIT('h87)
	) name2726 (
		_w2075_,
		_w2076_,
		_w2081_,
		_w3189_
	);
	LUT4 #(
		.INIT('h0200)
	) name2727 (
		_w3186_,
		_w3187_,
		_w3188_,
		_w3189_,
		_w3190_
	);
	LUT2 #(
		.INIT('h6)
	) name2728 (
		_w2004_,
		_w2008_,
		_w3191_
	);
	LUT2 #(
		.INIT('h9)
	) name2729 (
		_w2219_,
		_w2223_,
		_w3192_
	);
	LUT4 #(
		.INIT('h0660)
	) name2730 (
		_w2004_,
		_w2008_,
		_w2219_,
		_w2223_,
		_w3193_
	);
	LUT4 #(
		.INIT('h4000)
	) name2731 (
		_w3181_,
		_w3185_,
		_w3190_,
		_w3193_,
		_w3194_
	);
	LUT2 #(
		.INIT('h1)
	) name2732 (
		_w2646_,
		_w2974_,
		_w3195_
	);
	LUT4 #(
		.INIT('h8000)
	) name2733 (
		_w3180_,
		_w3194_,
		_w3172_,
		_w3195_,
		_w3196_
	);
	LUT3 #(
		.INIT('h80)
	) name2734 (
		_w3167_,
		_w3196_,
		_w3164_,
		_w3197_
	);
	LUT4 #(
		.INIT('h8444)
	) name2735 (
		_w2291_,
		_w2425_,
		_w3159_,
		_w3197_,
		_w3198_
	);
	LUT4 #(
		.INIT('h00bf)
	) name2736 (
		_w3150_,
		_w3155_,
		_w3157_,
		_w3198_,
		_w3199_
	);
	LUT3 #(
		.INIT('he0)
	) name2737 (
		_w2282_,
		_w3156_,
		_w3199_,
		_w3200_
	);
	LUT4 #(
		.INIT('h0777)
	) name2738 (
		_w2395_,
		_w2396_,
		_w2417_,
		_w2418_,
		_w3201_
	);
	LUT3 #(
		.INIT('h01)
	) name2739 (
		_w1748_,
		_w3134_,
		_w3201_,
		_w3202_
	);
	LUT2 #(
		.INIT('h1)
	) name2740 (
		_w3139_,
		_w3202_,
		_w3203_
	);
	LUT4 #(
		.INIT('h0001)
	) name2741 (
		_w2278_,
		_w2357_,
		_w3139_,
		_w3202_,
		_w3204_
	);
	LUT2 #(
		.INIT('h8)
	) name2742 (
		_w2828_,
		_w3204_,
		_w3205_
	);
	LUT2 #(
		.INIT('h8)
	) name2743 (
		_w2837_,
		_w3204_,
		_w3206_
	);
	LUT4 #(
		.INIT('h3031)
	) name2744 (
		_w1748_,
		_w2397_,
		_w2419_,
		_w3134_,
		_w3207_
	);
	LUT2 #(
		.INIT('h2)
	) name2745 (
		_w3126_,
		_w3207_,
		_w3208_
	);
	LUT3 #(
		.INIT('h07)
	) name2746 (
		_w3151_,
		_w3203_,
		_w3208_,
		_w3209_
	);
	LUT2 #(
		.INIT('h4)
	) name2747 (
		_w3206_,
		_w3209_,
		_w3210_
	);
	LUT3 #(
		.INIT('hb0)
	) name2748 (
		_w2976_,
		_w3205_,
		_w3210_,
		_w3211_
	);
	LUT3 #(
		.INIT('h08)
	) name2749 (
		_w1723_,
		_w2289_,
		_w2291_,
		_w3212_
	);
	LUT3 #(
		.INIT('h80)
	) name2750 (
		_w1723_,
		_w2289_,
		_w2291_,
		_w3213_
	);
	LUT4 #(
		.INIT('h014f)
	) name2751 (
		\P1_B_reg/NET0131 ,
		_w3211_,
		_w3212_,
		_w3213_,
		_w3214_
	);
	LUT4 #(
		.INIT('hd000)
	) name2752 (
		_w2282_,
		_w3146_,
		_w3200_,
		_w3214_,
		_w3215_
	);
	LUT3 #(
		.INIT('h2e)
	) name2753 (
		\P1_B_reg/NET0131 ,
		_w2695_,
		_w3215_,
		_w3216_
	);
	LUT2 #(
		.INIT('h8)
	) name2754 (
		_w1833_,
		_w2460_,
		_w3217_
	);
	LUT2 #(
		.INIT('h2)
	) name2755 (
		_w1833_,
		_w2644_,
		_w3218_
	);
	LUT4 #(
		.INIT('h007d)
	) name2756 (
		_w2644_,
		_w2787_,
		_w2788_,
		_w3218_,
		_w3219_
	);
	LUT4 #(
		.INIT('h08c8)
	) name2757 (
		_w1833_,
		_w2388_,
		_w2644_,
		_w2839_,
		_w3220_
	);
	LUT4 #(
		.INIT('h0040)
	) name2758 (
		_w2445_,
		_w2447_,
		_w2644_,
		_w2842_,
		_w3221_
	);
	LUT4 #(
		.INIT('hc808)
	) name2759 (
		_w1833_,
		_w2424_,
		_w2644_,
		_w2845_,
		_w3222_
	);
	LUT3 #(
		.INIT('h01)
	) name2760 (
		_w1748_,
		_w1815_,
		_w2689_,
		_w3223_
	);
	LUT2 #(
		.INIT('h2)
	) name2761 (
		_w1833_,
		_w2690_,
		_w3224_
	);
	LUT2 #(
		.INIT('h1)
	) name2762 (
		_w3223_,
		_w3224_,
		_w3225_
	);
	LUT3 #(
		.INIT('h10)
	) name2763 (
		_w3222_,
		_w3221_,
		_w3225_,
		_w3226_
	);
	LUT4 #(
		.INIT('h0d00)
	) name2764 (
		_w2292_,
		_w3219_,
		_w3220_,
		_w3226_,
		_w3227_
	);
	LUT4 #(
		.INIT('ha0a8)
	) name2765 (
		\P1_state_reg[0]/NET0131 ,
		_w1731_,
		_w3217_,
		_w3227_,
		_w3228_
	);
	LUT2 #(
		.INIT('h2)
	) name2766 (
		\P1_reg3_reg[28]/NET0131 ,
		\P1_state_reg[0]/NET0131 ,
		_w3229_
	);
	LUT3 #(
		.INIT('h07)
	) name2767 (
		_w1833_,
		_w2695_,
		_w3229_,
		_w3230_
	);
	LUT2 #(
		.INIT('hb)
	) name2768 (
		_w3228_,
		_w3230_,
		_w3231_
	);
	LUT2 #(
		.INIT('h4)
	) name2769 (
		_w1030_,
		_w1357_,
		_w3232_
	);
	LUT4 #(
		.INIT('h0155)
	) name2770 (
		_w1030_,
		_w1361_,
		_w1363_,
		_w1368_,
		_w3233_
	);
	LUT4 #(
		.INIT('h8848)
	) name2771 (
		_w1271_,
		_w1369_,
		_w1674_,
		_w2485_,
		_w3234_
	);
	LUT3 #(
		.INIT('h54)
	) name2772 (
		_w1409_,
		_w3233_,
		_w3234_,
		_w3235_
	);
	LUT4 #(
		.INIT('h04c4)
	) name2773 (
		_w1030_,
		_w1191_,
		_w1411_,
		_w2491_,
		_w3236_
	);
	LUT3 #(
		.INIT('h54)
	) name2774 (
		_w1030_,
		_w1441_,
		_w1443_,
		_w3237_
	);
	LUT4 #(
		.INIT('h00ef)
	) name2775 (
		_w546_,
		_w1026_,
		_w1440_,
		_w3237_,
		_w3238_
	);
	LUT2 #(
		.INIT('h4)
	) name2776 (
		_w3236_,
		_w3238_,
		_w3239_
	);
	LUT4 #(
		.INIT('h010d)
	) name2777 (
		_w1030_,
		_w1369_,
		_w1496_,
		_w2499_,
		_w3240_
	);
	LUT4 #(
		.INIT('h04c4)
	) name2778 (
		_w1030_,
		_w1447_,
		_w1411_,
		_w2499_,
		_w3241_
	);
	LUT4 #(
		.INIT('h0100)
	) name2779 (
		_w3235_,
		_w3240_,
		_w3241_,
		_w3239_,
		_w3242_
	);
	LUT4 #(
		.INIT('ha0a8)
	) name2780 (
		\P1_state_reg[0]/NET0131 ,
		_w1359_,
		_w3232_,
		_w3242_,
		_w3243_
	);
	LUT2 #(
		.INIT('h4)
	) name2781 (
		\P1_state_reg[0]/NET0131 ,
		\P2_reg3_reg[25]/NET0131 ,
		_w3244_
	);
	LUT3 #(
		.INIT('h0b)
	) name2782 (
		_w1030_,
		_w1349_,
		_w3244_,
		_w3245_
	);
	LUT2 #(
		.INIT('hb)
	) name2783 (
		_w3243_,
		_w3245_,
		_w3246_
	);
	LUT4 #(
		.INIT('hf200)
	) name2784 (
		\P2_reg3_reg[26]/NET0131 ,
		_w1029_,
		_w1062_,
		_w1357_,
		_w3247_
	);
	LUT2 #(
		.INIT('h1)
	) name2785 (
		_w1063_,
		_w1411_,
		_w3248_
	);
	LUT3 #(
		.INIT('h10)
	) name2786 (
		_w1269_,
		_w1273_,
		_w1480_,
		_w3249_
	);
	LUT4 #(
		.INIT('h1000)
	) name2787 (
		_w1269_,
		_w1273_,
		_w1480_,
		_w2616_,
		_w3250_
	);
	LUT4 #(
		.INIT('h4f00)
	) name2788 (
		_w2540_,
		_w2541_,
		_w2542_,
		_w3250_,
		_w3251_
	);
	LUT3 #(
		.INIT('h01)
	) name2789 (
		_w1269_,
		_w1266_,
		_w1567_,
		_w3252_
	);
	LUT4 #(
		.INIT('h008a)
	) name2790 (
		_w1570_,
		_w2615_,
		_w3249_,
		_w3252_,
		_w3253_
	);
	LUT4 #(
		.INIT('h4844)
	) name2791 (
		_w1257_,
		_w1411_,
		_w3251_,
		_w3253_,
		_w3254_
	);
	LUT3 #(
		.INIT('ha8)
	) name2792 (
		_w1447_,
		_w3248_,
		_w3254_,
		_w3255_
	);
	LUT4 #(
		.INIT('h002f)
	) name2793 (
		_w519_,
		_w1030_,
		_w1034_,
		_w1435_,
		_w3256_
	);
	LUT4 #(
		.INIT('h7f00)
	) name2794 (
		_w1423_,
		_w1429_,
		_w1430_,
		_w1435_,
		_w3257_
	);
	LUT4 #(
		.INIT('h020f)
	) name2795 (
		_w1085_,
		_w2489_,
		_w3256_,
		_w3257_,
		_w3258_
	);
	LUT4 #(
		.INIT('h04c4)
	) name2796 (
		_w1063_,
		_w1191_,
		_w1411_,
		_w3258_,
		_w3259_
	);
	LUT3 #(
		.INIT('h54)
	) name2797 (
		_w1063_,
		_w1441_,
		_w1443_,
		_w3260_
	);
	LUT4 #(
		.INIT('h00ef)
	) name2798 (
		_w546_,
		_w1058_,
		_w1440_,
		_w3260_,
		_w3261_
	);
	LUT2 #(
		.INIT('h4)
	) name2799 (
		_w3259_,
		_w3261_,
		_w3262_
	);
	LUT2 #(
		.INIT('h1)
	) name2800 (
		_w1063_,
		_w1369_,
		_w3263_
	);
	LUT4 #(
		.INIT('h4844)
	) name2801 (
		_w1257_,
		_w1369_,
		_w3251_,
		_w3253_,
		_w3264_
	);
	LUT3 #(
		.INIT('h54)
	) name2802 (
		_w1496_,
		_w3263_,
		_w3264_,
		_w3265_
	);
	LUT3 #(
		.INIT('h02)
	) name2803 (
		_w1012_,
		_w1094_,
		_w1095_,
		_w3266_
	);
	LUT4 #(
		.INIT('h0200)
	) name2804 (
		_w1012_,
		_w1094_,
		_w1095_,
		_w2629_,
		_w3267_
	);
	LUT4 #(
		.INIT('h5d00)
	) name2805 (
		_w2549_,
		_w2550_,
		_w2557_,
		_w3267_,
		_w3268_
	);
	LUT3 #(
		.INIT('h10)
	) name2806 (
		_w1094_,
		_w1095_,
		_w1219_,
		_w3269_
	);
	LUT4 #(
		.INIT('h0045)
	) name2807 (
		_w1222_,
		_w2628_,
		_w3266_,
		_w3269_,
		_w3270_
	);
	LUT4 #(
		.INIT('h8488)
	) name2808 (
		_w1257_,
		_w1369_,
		_w3268_,
		_w3270_,
		_w3271_
	);
	LUT3 #(
		.INIT('h54)
	) name2809 (
		_w1409_,
		_w3263_,
		_w3271_,
		_w3272_
	);
	LUT4 #(
		.INIT('h0100)
	) name2810 (
		_w3255_,
		_w3265_,
		_w3272_,
		_w3262_,
		_w3273_
	);
	LUT4 #(
		.INIT('ha0a8)
	) name2811 (
		\P1_state_reg[0]/NET0131 ,
		_w1359_,
		_w3247_,
		_w3273_,
		_w3274_
	);
	LUT2 #(
		.INIT('h4)
	) name2812 (
		\P1_state_reg[0]/NET0131 ,
		\P2_reg3_reg[26]/NET0131 ,
		_w3275_
	);
	LUT4 #(
		.INIT('hf200)
	) name2813 (
		\P2_reg3_reg[26]/NET0131 ,
		_w1029_,
		_w1062_,
		_w1349_,
		_w3276_
	);
	LUT2 #(
		.INIT('h1)
	) name2814 (
		_w3275_,
		_w3276_,
		_w3277_
	);
	LUT2 #(
		.INIT('hb)
	) name2815 (
		_w3274_,
		_w3277_,
		_w3278_
	);
	LUT4 #(
		.INIT('hd070)
	) name2816 (
		\P1_state_reg[0]/NET0131 ,
		\P2_IR_reg[23]/NET0131 ,
		\P2_reg2_reg[21]/NET0131 ,
		_w1188_,
		_w3279_
	);
	LUT4 #(
		.INIT('h2000)
	) name2817 (
		\P2_reg2_reg[21]/NET0131 ,
		_w1189_,
		_w1352_,
		_w1356_,
		_w3280_
	);
	LUT4 #(
		.INIT('h59aa)
	) name2818 (
		_w1283_,
		_w1693_,
		_w1699_,
		_w1703_,
		_w3281_
	);
	LUT4 #(
		.INIT('h020e)
	) name2819 (
		\P2_reg2_reg[21]/NET0131 ,
		_w1507_,
		_w1575_,
		_w3281_,
		_w3282_
	);
	LUT4 #(
		.INIT('h5400)
	) name2820 (
		_w546_,
		_w935_,
		_w944_,
		_w1442_,
		_w3283_
	);
	LUT3 #(
		.INIT('h40)
	) name2821 (
		_w947_,
		_w1229_,
		_w1232_,
		_w3284_
	);
	LUT4 #(
		.INIT('h0057)
	) name2822 (
		\P2_reg2_reg[21]/NET0131 ,
		_w1441_,
		_w1523_,
		_w3284_,
		_w3285_
	);
	LUT3 #(
		.INIT('h70)
	) name2823 (
		_w1507_,
		_w3283_,
		_w3285_,
		_w3286_
	);
	LUT2 #(
		.INIT('h4)
	) name2824 (
		_w3282_,
		_w3286_,
		_w3287_
	);
	LUT3 #(
		.INIT('h0b)
	) name2825 (
		_w964_,
		_w968_,
		_w1435_,
		_w3288_
	);
	LUT4 #(
		.INIT('h007b)
	) name2826 (
		_w1006_,
		_w1435_,
		_w2623_,
		_w3288_,
		_w3289_
	);
	LUT4 #(
		.INIT('h08c8)
	) name2827 (
		\P2_reg2_reg[21]/NET0131 ,
		_w1191_,
		_w1516_,
		_w3289_,
		_w3290_
	);
	LUT4 #(
		.INIT('ha655)
	) name2828 (
		_w1283_,
		_w1659_,
		_w1664_,
		_w1668_,
		_w3291_
	);
	LUT4 #(
		.INIT('h0232)
	) name2829 (
		\P2_reg2_reg[21]/NET0131 ,
		_w1506_,
		_w1507_,
		_w3291_,
		_w3292_
	);
	LUT4 #(
		.INIT('h20e0)
	) name2830 (
		\P2_reg2_reg[21]/NET0131 ,
		_w1516_,
		_w1530_,
		_w3291_,
		_w3293_
	);
	LUT3 #(
		.INIT('h01)
	) name2831 (
		_w3292_,
		_w3293_,
		_w3290_,
		_w3294_
	);
	LUT4 #(
		.INIT('h3111)
	) name2832 (
		_w1359_,
		_w3280_,
		_w3287_,
		_w3294_,
		_w3295_
	);
	LUT3 #(
		.INIT('hce)
	) name2833 (
		\P1_state_reg[0]/NET0131 ,
		_w3279_,
		_w3295_,
		_w3296_
	);
	LUT4 #(
		.INIT('hd070)
	) name2834 (
		\P1_state_reg[0]/NET0131 ,
		\P2_IR_reg[23]/NET0131 ,
		\P2_reg0_reg[24]/NET0131 ,
		_w1188_,
		_w3297_
	);
	LUT4 #(
		.INIT('h2000)
	) name2835 (
		\P2_reg0_reg[24]/NET0131 ,
		_w1189_,
		_w1352_,
		_w1356_,
		_w3298_
	);
	LUT4 #(
		.INIT('haaa8)
	) name2836 (
		\P2_reg0_reg[24]/NET0131 ,
		_w1361_,
		_w1363_,
		_w1368_,
		_w3299_
	);
	LUT4 #(
		.INIT('hb400)
	) name2837 (
		_w1208_,
		_w1221_,
		_w1268_,
		_w1411_,
		_w3300_
	);
	LUT3 #(
		.INIT('h54)
	) name2838 (
		_w1409_,
		_w3299_,
		_w3300_,
		_w3301_
	);
	LUT4 #(
		.INIT('h02aa)
	) name2839 (
		\P2_reg0_reg[24]/NET0131 ,
		_w1361_,
		_w1363_,
		_w1368_,
		_w3302_
	);
	LUT3 #(
		.INIT('ha8)
	) name2840 (
		_w1447_,
		_w1625_,
		_w3302_,
		_w3303_
	);
	LUT4 #(
		.INIT('h111d)
	) name2841 (
		\P2_reg0_reg[24]/NET0131 ,
		_w1369_,
		_w1627_,
		_w1628_,
		_w3304_
	);
	LUT3 #(
		.INIT('ha2)
	) name2842 (
		\P2_reg0_reg[24]/NET0131 ,
		_w1684_,
		_w1685_,
		_w3305_
	);
	LUT4 #(
		.INIT('h1000)
	) name2843 (
		_w546_,
		_w1041_,
		_w1411_,
		_w1442_,
		_w3306_
	);
	LUT2 #(
		.INIT('h1)
	) name2844 (
		_w3305_,
		_w3306_,
		_w3307_
	);
	LUT3 #(
		.INIT('hd0)
	) name2845 (
		_w1191_,
		_w3304_,
		_w3307_,
		_w3308_
	);
	LUT4 #(
		.INIT('hab00)
	) name2846 (
		_w1496_,
		_w1623_,
		_w3299_,
		_w3308_,
		_w3309_
	);
	LUT4 #(
		.INIT('ha8aa)
	) name2847 (
		_w1359_,
		_w3303_,
		_w3301_,
		_w3309_,
		_w3310_
	);
	LUT4 #(
		.INIT('heeec)
	) name2848 (
		\P1_state_reg[0]/NET0131 ,
		_w3297_,
		_w3298_,
		_w3310_,
		_w3311_
	);
	LUT4 #(
		.INIT('hd070)
	) name2849 (
		\P1_state_reg[0]/NET0131 ,
		\P2_IR_reg[23]/NET0131 ,
		\P2_reg0_reg[25]/NET0131 ,
		_w1188_,
		_w3312_
	);
	LUT4 #(
		.INIT('h2000)
	) name2850 (
		\P2_reg0_reg[25]/NET0131 ,
		_w1189_,
		_w1352_,
		_w1356_,
		_w3313_
	);
	LUT4 #(
		.INIT('haaa8)
	) name2851 (
		\P2_reg0_reg[25]/NET0131 ,
		_w1361_,
		_w1363_,
		_w1368_,
		_w3314_
	);
	LUT4 #(
		.INIT('h8848)
	) name2852 (
		_w1271_,
		_w1411_,
		_w1674_,
		_w2485_,
		_w3315_
	);
	LUT3 #(
		.INIT('h54)
	) name2853 (
		_w1409_,
		_w3314_,
		_w3315_,
		_w3316_
	);
	LUT4 #(
		.INIT('h08c8)
	) name2854 (
		\P2_reg0_reg[25]/NET0131 ,
		_w1191_,
		_w1369_,
		_w2491_,
		_w3317_
	);
	LUT4 #(
		.INIT('h1000)
	) name2855 (
		_w546_,
		_w1026_,
		_w1411_,
		_w1442_,
		_w3318_
	);
	LUT3 #(
		.INIT('ha2)
	) name2856 (
		\P2_reg0_reg[25]/NET0131 ,
		_w1684_,
		_w1685_,
		_w3319_
	);
	LUT2 #(
		.INIT('h1)
	) name2857 (
		_w3318_,
		_w3319_,
		_w3320_
	);
	LUT2 #(
		.INIT('h4)
	) name2858 (
		_w3317_,
		_w3320_,
		_w3321_
	);
	LUT4 #(
		.INIT('h020e)
	) name2859 (
		\P2_reg0_reg[25]/NET0131 ,
		_w1411_,
		_w1496_,
		_w2499_,
		_w3322_
	);
	LUT4 #(
		.INIT('h20e0)
	) name2860 (
		\P2_reg0_reg[25]/NET0131 ,
		_w1369_,
		_w1447_,
		_w2499_,
		_w3323_
	);
	LUT4 #(
		.INIT('h0100)
	) name2861 (
		_w3316_,
		_w3322_,
		_w3323_,
		_w3321_,
		_w3324_
	);
	LUT4 #(
		.INIT('ha0a8)
	) name2862 (
		\P1_state_reg[0]/NET0131 ,
		_w1359_,
		_w3313_,
		_w3324_,
		_w3325_
	);
	LUT2 #(
		.INIT('he)
	) name2863 (
		_w3312_,
		_w3325_,
		_w3326_
	);
	LUT4 #(
		.INIT('hd070)
	) name2864 (
		\P1_state_reg[0]/NET0131 ,
		\P2_IR_reg[23]/NET0131 ,
		\P2_reg0_reg[26]/NET0131 ,
		_w1188_,
		_w3327_
	);
	LUT4 #(
		.INIT('h2000)
	) name2865 (
		\P2_reg0_reg[26]/NET0131 ,
		_w1189_,
		_w1352_,
		_w1356_,
		_w3328_
	);
	LUT4 #(
		.INIT('haaa8)
	) name2866 (
		\P2_reg0_reg[26]/NET0131 ,
		_w1361_,
		_w1363_,
		_w1368_,
		_w3329_
	);
	LUT4 #(
		.INIT('h8488)
	) name2867 (
		_w1257_,
		_w1411_,
		_w3268_,
		_w3270_,
		_w3330_
	);
	LUT3 #(
		.INIT('h54)
	) name2868 (
		_w1409_,
		_w3329_,
		_w3330_,
		_w3331_
	);
	LUT4 #(
		.INIT('h02aa)
	) name2869 (
		\P2_reg0_reg[26]/NET0131 ,
		_w1361_,
		_w1363_,
		_w1368_,
		_w3332_
	);
	LUT4 #(
		.INIT('h08c8)
	) name2870 (
		\P2_reg0_reg[26]/NET0131 ,
		_w1191_,
		_w1369_,
		_w3258_,
		_w3333_
	);
	LUT3 #(
		.INIT('ha2)
	) name2871 (
		\P2_reg0_reg[26]/NET0131 ,
		_w1684_,
		_w1685_,
		_w3334_
	);
	LUT4 #(
		.INIT('h00ef)
	) name2872 (
		_w546_,
		_w1058_,
		_w1687_,
		_w3334_,
		_w3335_
	);
	LUT2 #(
		.INIT('h4)
	) name2873 (
		_w3333_,
		_w3335_,
		_w3336_
	);
	LUT3 #(
		.INIT('ha8)
	) name2874 (
		_w1447_,
		_w3264_,
		_w3332_,
		_w3337_
	);
	LUT3 #(
		.INIT('h54)
	) name2875 (
		_w1496_,
		_w3254_,
		_w3329_,
		_w3338_
	);
	LUT4 #(
		.INIT('h0100)
	) name2876 (
		_w3331_,
		_w3337_,
		_w3338_,
		_w3336_,
		_w3339_
	);
	LUT4 #(
		.INIT('ha0a8)
	) name2877 (
		\P1_state_reg[0]/NET0131 ,
		_w1359_,
		_w3328_,
		_w3339_,
		_w3340_
	);
	LUT2 #(
		.INIT('he)
	) name2878 (
		_w3327_,
		_w3340_,
		_w3341_
	);
	LUT4 #(
		.INIT('h2000)
	) name2879 (
		\P1_reg2_reg[27]/NET0131 ,
		_w1723_,
		_w1727_,
		_w1730_,
		_w3342_
	);
	LUT4 #(
		.INIT('h20e0)
	) name2880 (
		\P1_reg2_reg[27]/NET0131 ,
		_w1741_,
		_w2292_,
		_w2665_,
		_w3343_
	);
	LUT4 #(
		.INIT('h20e0)
	) name2881 (
		\P1_reg2_reg[27]/NET0131 ,
		_w1741_,
		_w2388_,
		_w2682_,
		_w3344_
	);
	LUT4 #(
		.INIT('h5400)
	) name2882 (
		_w1748_,
		_w1907_,
		_w1929_,
		_w2426_,
		_w3345_
	);
	LUT3 #(
		.INIT('ha8)
	) name2883 (
		_w1741_,
		_w2688_,
		_w3345_,
		_w3346_
	);
	LUT4 #(
		.INIT('h111d)
	) name2884 (
		\P1_reg2_reg[27]/NET0131 ,
		_w1741_,
		_w2684_,
		_w2686_,
		_w3347_
	);
	LUT4 #(
		.INIT('ha2a0)
	) name2885 (
		\P1_reg2_reg[27]/NET0131 ,
		_w1741_,
		_w2450_,
		_w2452_,
		_w3348_
	);
	LUT2 #(
		.INIT('h8)
	) name2886 (
		_w1932_,
		_w2454_,
		_w3349_
	);
	LUT2 #(
		.INIT('h1)
	) name2887 (
		_w3348_,
		_w3349_,
		_w3350_
	);
	LUT4 #(
		.INIT('h3100)
	) name2888 (
		_w2424_,
		_w3346_,
		_w3347_,
		_w3350_,
		_w3351_
	);
	LUT4 #(
		.INIT('ha8aa)
	) name2889 (
		_w1731_,
		_w3343_,
		_w3344_,
		_w3351_,
		_w3352_
	);
	LUT2 #(
		.INIT('h2)
	) name2890 (
		\P1_reg2_reg[27]/NET0131 ,
		_w2462_,
		_w3353_
	);
	LUT4 #(
		.INIT('hffa8)
	) name2891 (
		\P1_state_reg[0]/NET0131 ,
		_w3342_,
		_w3352_,
		_w3353_,
		_w3354_
	);
	LUT4 #(
		.INIT('hd070)
	) name2892 (
		\P1_state_reg[0]/NET0131 ,
		\P2_IR_reg[23]/NET0131 ,
		\P2_reg1_reg[24]/NET0131 ,
		_w1188_,
		_w3355_
	);
	LUT4 #(
		.INIT('h2000)
	) name2893 (
		\P2_reg1_reg[24]/NET0131 ,
		_w1189_,
		_w1352_,
		_w1356_,
		_w3356_
	);
	LUT4 #(
		.INIT('ha8aa)
	) name2894 (
		\P2_reg1_reg[24]/NET0131 ,
		_w1361_,
		_w1363_,
		_w1368_,
		_w3357_
	);
	LUT3 #(
		.INIT('ha8)
	) name2895 (
		_w1530_,
		_w1641_,
		_w3357_,
		_w3358_
	);
	LUT4 #(
		.INIT('haa02)
	) name2896 (
		\P2_reg1_reg[24]/NET0131 ,
		_w1361_,
		_w1363_,
		_w1368_,
		_w3359_
	);
	LUT3 #(
		.INIT('h54)
	) name2897 (
		_w1506_,
		_w1644_,
		_w3359_,
		_w3360_
	);
	LUT4 #(
		.INIT('h4844)
	) name2898 (
		_w1268_,
		_w1516_,
		_w1620_,
		_w1622_,
		_w3361_
	);
	LUT4 #(
		.INIT('h111d)
	) name2899 (
		\P2_reg1_reg[24]/NET0131 ,
		_w1507_,
		_w1627_,
		_w1628_,
		_w3362_
	);
	LUT4 #(
		.INIT('h1000)
	) name2900 (
		_w546_,
		_w1041_,
		_w1442_,
		_w1516_,
		_w3363_
	);
	LUT3 #(
		.INIT('ha2)
	) name2901 (
		\P2_reg1_reg[24]/NET0131 ,
		_w1684_,
		_w2469_,
		_w3364_
	);
	LUT2 #(
		.INIT('h1)
	) name2902 (
		_w3363_,
		_w3364_,
		_w3365_
	);
	LUT3 #(
		.INIT('hd0)
	) name2903 (
		_w1191_,
		_w3362_,
		_w3365_,
		_w3366_
	);
	LUT4 #(
		.INIT('hab00)
	) name2904 (
		_w1575_,
		_w3359_,
		_w3361_,
		_w3366_,
		_w3367_
	);
	LUT4 #(
		.INIT('ha8aa)
	) name2905 (
		_w1359_,
		_w3360_,
		_w3358_,
		_w3367_,
		_w3368_
	);
	LUT4 #(
		.INIT('heeec)
	) name2906 (
		\P1_state_reg[0]/NET0131 ,
		_w3355_,
		_w3356_,
		_w3368_,
		_w3369_
	);
	LUT4 #(
		.INIT('hd070)
	) name2907 (
		\P1_state_reg[0]/NET0131 ,
		\P2_IR_reg[23]/NET0131 ,
		\P2_reg1_reg[26]/NET0131 ,
		_w1188_,
		_w3370_
	);
	LUT4 #(
		.INIT('h2000)
	) name2908 (
		\P2_reg1_reg[26]/NET0131 ,
		_w1189_,
		_w1352_,
		_w1356_,
		_w3371_
	);
	LUT4 #(
		.INIT('haa02)
	) name2909 (
		\P2_reg1_reg[26]/NET0131 ,
		_w1361_,
		_w1363_,
		_w1368_,
		_w3372_
	);
	LUT4 #(
		.INIT('h8488)
	) name2910 (
		_w1257_,
		_w1516_,
		_w3268_,
		_w3270_,
		_w3373_
	);
	LUT3 #(
		.INIT('h54)
	) name2911 (
		_w1506_,
		_w3372_,
		_w3373_,
		_w3374_
	);
	LUT4 #(
		.INIT('ha8aa)
	) name2912 (
		\P2_reg1_reg[26]/NET0131 ,
		_w1361_,
		_w1363_,
		_w1368_,
		_w3375_
	);
	LUT4 #(
		.INIT('h08c8)
	) name2913 (
		\P2_reg1_reg[26]/NET0131 ,
		_w1191_,
		_w1507_,
		_w3258_,
		_w3376_
	);
	LUT3 #(
		.INIT('ha2)
	) name2914 (
		\P2_reg1_reg[26]/NET0131 ,
		_w1684_,
		_w2469_,
		_w3377_
	);
	LUT4 #(
		.INIT('h00ef)
	) name2915 (
		_w546_,
		_w1058_,
		_w2471_,
		_w3377_,
		_w3378_
	);
	LUT2 #(
		.INIT('h4)
	) name2916 (
		_w3376_,
		_w3378_,
		_w3379_
	);
	LUT4 #(
		.INIT('h8488)
	) name2917 (
		_w1257_,
		_w1507_,
		_w3268_,
		_w3270_,
		_w3380_
	);
	LUT3 #(
		.INIT('ha8)
	) name2918 (
		_w1530_,
		_w3375_,
		_w3380_,
		_w3381_
	);
	LUT4 #(
		.INIT('h4844)
	) name2919 (
		_w1257_,
		_w1516_,
		_w3251_,
		_w3253_,
		_w3382_
	);
	LUT3 #(
		.INIT('h54)
	) name2920 (
		_w1575_,
		_w3372_,
		_w3382_,
		_w3383_
	);
	LUT4 #(
		.INIT('h0100)
	) name2921 (
		_w3374_,
		_w3381_,
		_w3383_,
		_w3379_,
		_w3384_
	);
	LUT4 #(
		.INIT('ha0a8)
	) name2922 (
		\P1_state_reg[0]/NET0131 ,
		_w1359_,
		_w3371_,
		_w3384_,
		_w3385_
	);
	LUT2 #(
		.INIT('he)
	) name2923 (
		_w3370_,
		_w3385_,
		_w3386_
	);
	LUT4 #(
		.INIT('hd070)
	) name2924 (
		\P1_state_reg[0]/NET0131 ,
		\P2_IR_reg[23]/NET0131 ,
		\P2_reg1_reg[25]/NET0131 ,
		_w1188_,
		_w3387_
	);
	LUT4 #(
		.INIT('h2000)
	) name2925 (
		\P2_reg1_reg[25]/NET0131 ,
		_w1189_,
		_w1352_,
		_w1356_,
		_w3388_
	);
	LUT4 #(
		.INIT('haa02)
	) name2926 (
		\P2_reg1_reg[25]/NET0131 ,
		_w1361_,
		_w1363_,
		_w1368_,
		_w3389_
	);
	LUT3 #(
		.INIT('h54)
	) name2927 (
		_w1506_,
		_w2501_,
		_w3389_,
		_w3390_
	);
	LUT4 #(
		.INIT('ha8aa)
	) name2928 (
		\P2_reg1_reg[25]/NET0131 ,
		_w1361_,
		_w1363_,
		_w1368_,
		_w3391_
	);
	LUT4 #(
		.INIT('h08c8)
	) name2929 (
		\P2_reg1_reg[25]/NET0131 ,
		_w1191_,
		_w1507_,
		_w2491_,
		_w3392_
	);
	LUT4 #(
		.INIT('h1000)
	) name2930 (
		_w546_,
		_w1026_,
		_w1442_,
		_w1516_,
		_w3393_
	);
	LUT3 #(
		.INIT('ha2)
	) name2931 (
		\P2_reg1_reg[25]/NET0131 ,
		_w1684_,
		_w2469_,
		_w3394_
	);
	LUT2 #(
		.INIT('h1)
	) name2932 (
		_w3393_,
		_w3394_,
		_w3395_
	);
	LUT2 #(
		.INIT('h4)
	) name2933 (
		_w3392_,
		_w3395_,
		_w3396_
	);
	LUT4 #(
		.INIT('h020e)
	) name2934 (
		\P2_reg1_reg[25]/NET0131 ,
		_w1516_,
		_w1575_,
		_w2499_,
		_w3397_
	);
	LUT3 #(
		.INIT('ha8)
	) name2935 (
		_w1530_,
		_w2486_,
		_w3391_,
		_w3398_
	);
	LUT4 #(
		.INIT('h0100)
	) name2936 (
		_w3390_,
		_w3397_,
		_w3398_,
		_w3396_,
		_w3399_
	);
	LUT4 #(
		.INIT('ha0a8)
	) name2937 (
		\P1_state_reg[0]/NET0131 ,
		_w1359_,
		_w3388_,
		_w3399_,
		_w3400_
	);
	LUT2 #(
		.INIT('he)
	) name2938 (
		_w3387_,
		_w3400_,
		_w3401_
	);
	LUT2 #(
		.INIT('h2)
	) name2939 (
		\P1_reg0_reg[26]/NET0131 ,
		_w2462_,
		_w3402_
	);
	LUT4 #(
		.INIT('h2000)
	) name2940 (
		\P1_reg0_reg[26]/NET0131 ,
		_w1723_,
		_w1727_,
		_w1730_,
		_w3403_
	);
	LUT2 #(
		.INIT('h2)
	) name2941 (
		\P1_reg0_reg[26]/NET0131 ,
		_w2883_,
		_w3404_
	);
	LUT4 #(
		.INIT('h7020)
	) name2942 (
		_w1747_,
		_w1876_,
		_w2883_,
		_w2923_,
		_w3405_
	);
	LUT3 #(
		.INIT('h10)
	) name2943 (
		_w1748_,
		_w1899_,
		_w2426_,
		_w3406_
	);
	LUT4 #(
		.INIT('h006f)
	) name2944 (
		_w1900_,
		_w2443_,
		_w2447_,
		_w3406_,
		_w3407_
	);
	LUT3 #(
		.INIT('hc4)
	) name2945 (
		_w2452_,
		_w2524_,
		_w2883_,
		_w3408_
	);
	LUT4 #(
		.INIT('h0a8a)
	) name2946 (
		\P1_reg0_reg[26]/NET0131 ,
		_w2452_,
		_w2524_,
		_w2883_,
		_w3409_
	);
	LUT3 #(
		.INIT('h0d)
	) name2947 (
		_w2883_,
		_w3407_,
		_w3409_,
		_w3410_
	);
	LUT4 #(
		.INIT('h5700)
	) name2948 (
		_w2424_,
		_w3404_,
		_w3405_,
		_w3410_,
		_w3411_
	);
	LUT4 #(
		.INIT('h08c8)
	) name2949 (
		\P1_reg0_reg[26]/NET0131 ,
		_w2292_,
		_w2883_,
		_w2967_,
		_w3412_
	);
	LUT4 #(
		.INIT('h08c8)
	) name2950 (
		\P1_reg0_reg[26]/NET0131 ,
		_w2388_,
		_w2883_,
		_w2948_,
		_w3413_
	);
	LUT4 #(
		.INIT('ha8aa)
	) name2951 (
		_w1731_,
		_w3412_,
		_w3413_,
		_w3411_,
		_w3414_
	);
	LUT4 #(
		.INIT('heeec)
	) name2952 (
		\P1_state_reg[0]/NET0131 ,
		_w3402_,
		_w3403_,
		_w3414_,
		_w3415_
	);
	LUT4 #(
		.INIT('h2000)
	) name2953 (
		\P1_reg0_reg[27]/NET0131 ,
		_w1723_,
		_w1727_,
		_w1730_,
		_w3416_
	);
	LUT4 #(
		.INIT('h0c88)
	) name2954 (
		\P1_reg0_reg[27]/NET0131 ,
		_w2292_,
		_w2665_,
		_w2883_,
		_w3417_
	);
	LUT4 #(
		.INIT('h0c88)
	) name2955 (
		\P1_reg0_reg[27]/NET0131 ,
		_w2388_,
		_w2682_,
		_w2883_,
		_w3418_
	);
	LUT3 #(
		.INIT('hc8)
	) name2956 (
		_w2688_,
		_w2883_,
		_w3345_,
		_w3419_
	);
	LUT4 #(
		.INIT('hf010)
	) name2957 (
		_w2426_,
		_w2447_,
		_w2524_,
		_w2883_,
		_w3420_
	);
	LUT2 #(
		.INIT('h2)
	) name2958 (
		\P1_reg0_reg[27]/NET0131 ,
		_w3420_,
		_w3421_
	);
	LUT4 #(
		.INIT('h0355)
	) name2959 (
		\P1_reg0_reg[27]/NET0131 ,
		_w2684_,
		_w2686_,
		_w2883_,
		_w3422_
	);
	LUT4 #(
		.INIT('h0301)
	) name2960 (
		_w2424_,
		_w3419_,
		_w3421_,
		_w3422_,
		_w3423_
	);
	LUT4 #(
		.INIT('ha8aa)
	) name2961 (
		_w1731_,
		_w3417_,
		_w3418_,
		_w3423_,
		_w3424_
	);
	LUT2 #(
		.INIT('h2)
	) name2962 (
		\P1_reg0_reg[27]/NET0131 ,
		_w2462_,
		_w3425_
	);
	LUT4 #(
		.INIT('hffa8)
	) name2963 (
		\P1_state_reg[0]/NET0131 ,
		_w3416_,
		_w3424_,
		_w3425_,
		_w3426_
	);
	LUT2 #(
		.INIT('h2)
	) name2964 (
		\P1_reg0_reg[28]/NET0131 ,
		_w2462_,
		_w3427_
	);
	LUT4 #(
		.INIT('h2000)
	) name2965 (
		\P1_reg0_reg[28]/NET0131 ,
		_w1723_,
		_w1727_,
		_w1730_,
		_w3428_
	);
	LUT4 #(
		.INIT('h3c55)
	) name2966 (
		\P1_reg0_reg[28]/NET0131 ,
		_w2787_,
		_w2788_,
		_w2883_,
		_w3429_
	);
	LUT4 #(
		.INIT('h0c88)
	) name2967 (
		\P1_reg0_reg[28]/NET0131 ,
		_w2388_,
		_w2839_,
		_w2883_,
		_w3430_
	);
	LUT2 #(
		.INIT('h2)
	) name2968 (
		\P1_reg0_reg[28]/NET0131 ,
		_w3420_,
		_w3431_
	);
	LUT4 #(
		.INIT('hc088)
	) name2969 (
		\P1_reg0_reg[28]/NET0131 ,
		_w2424_,
		_w2845_,
		_w2883_,
		_w3432_
	);
	LUT4 #(
		.INIT('h000b)
	) name2970 (
		_w2843_,
		_w2883_,
		_w3431_,
		_w3432_,
		_w3433_
	);
	LUT4 #(
		.INIT('h0d00)
	) name2971 (
		_w2292_,
		_w3429_,
		_w3430_,
		_w3433_,
		_w3434_
	);
	LUT4 #(
		.INIT('ha0a8)
	) name2972 (
		\P1_state_reg[0]/NET0131 ,
		_w1731_,
		_w3428_,
		_w3434_,
		_w3435_
	);
	LUT2 #(
		.INIT('he)
	) name2973 (
		_w3427_,
		_w3435_,
		_w3436_
	);
	LUT2 #(
		.INIT('h2)
	) name2974 (
		\P1_reg1_reg[27]/NET0131 ,
		_w2462_,
		_w3437_
	);
	LUT2 #(
		.INIT('h2)
	) name2975 (
		\P1_reg1_reg[27]/NET0131 ,
		_w2520_,
		_w3438_
	);
	LUT4 #(
		.INIT('h08c8)
	) name2976 (
		\P1_reg1_reg[27]/NET0131 ,
		_w2292_,
		_w2520_,
		_w2665_,
		_w3439_
	);
	LUT4 #(
		.INIT('h08c8)
	) name2977 (
		\P1_reg1_reg[27]/NET0131 ,
		_w2388_,
		_w2520_,
		_w2682_,
		_w3440_
	);
	LUT4 #(
		.INIT('h6300)
	) name2978 (
		_w1900_,
		_w1931_,
		_w2443_,
		_w2520_,
		_w3441_
	);
	LUT3 #(
		.INIT('ha8)
	) name2979 (
		_w2447_,
		_w3438_,
		_w3441_,
		_w3442_
	);
	LUT4 #(
		.INIT('h111d)
	) name2980 (
		\P1_reg1_reg[27]/NET0131 ,
		_w2520_,
		_w2684_,
		_w2686_,
		_w3443_
	);
	LUT4 #(
		.INIT('h08aa)
	) name2981 (
		\P1_reg1_reg[27]/NET0131 ,
		_w2426_,
		_w2520_,
		_w2524_,
		_w3444_
	);
	LUT3 #(
		.INIT('h07)
	) name2982 (
		_w2520_,
		_w3345_,
		_w3444_,
		_w3445_
	);
	LUT4 #(
		.INIT('h3100)
	) name2983 (
		_w2424_,
		_w3442_,
		_w3443_,
		_w3445_,
		_w3446_
	);
	LUT4 #(
		.INIT('ha8aa)
	) name2984 (
		_w1731_,
		_w3439_,
		_w3440_,
		_w3446_,
		_w3447_
	);
	LUT4 #(
		.INIT('h2000)
	) name2985 (
		\P1_reg1_reg[27]/NET0131 ,
		_w1723_,
		_w1727_,
		_w1730_,
		_w3448_
	);
	LUT4 #(
		.INIT('heeec)
	) name2986 (
		\P1_state_reg[0]/NET0131 ,
		_w3437_,
		_w3447_,
		_w3448_,
		_w3449_
	);
	LUT2 #(
		.INIT('h2)
	) name2987 (
		\P1_reg1_reg[28]/NET0131 ,
		_w2462_,
		_w3450_
	);
	LUT4 #(
		.INIT('h2000)
	) name2988 (
		\P1_reg1_reg[28]/NET0131 ,
		_w1723_,
		_w1727_,
		_w1730_,
		_w3451_
	);
	LUT4 #(
		.INIT('h1dd1)
	) name2989 (
		\P1_reg1_reg[28]/NET0131 ,
		_w2520_,
		_w2787_,
		_w2788_,
		_w3452_
	);
	LUT4 #(
		.INIT('h08c8)
	) name2990 (
		\P1_reg1_reg[28]/NET0131 ,
		_w2388_,
		_w2520_,
		_w2839_,
		_w3453_
	);
	LUT4 #(
		.INIT('hf5c5)
	) name2991 (
		\P1_reg1_reg[28]/NET0131 ,
		_w2445_,
		_w2520_,
		_w2842_,
		_w3454_
	);
	LUT4 #(
		.INIT('hc808)
	) name2992 (
		\P1_reg1_reg[28]/NET0131 ,
		_w2424_,
		_w2520_,
		_w2845_,
		_w3455_
	);
	LUT4 #(
		.INIT('h08aa)
	) name2993 (
		\P1_reg1_reg[28]/NET0131 ,
		_w2426_,
		_w2520_,
		_w2524_,
		_w3456_
	);
	LUT4 #(
		.INIT('h1000)
	) name2994 (
		_w1748_,
		_w1815_,
		_w2426_,
		_w2520_,
		_w3457_
	);
	LUT2 #(
		.INIT('h1)
	) name2995 (
		_w3456_,
		_w3457_,
		_w3458_
	);
	LUT4 #(
		.INIT('h0d00)
	) name2996 (
		_w2447_,
		_w3454_,
		_w3455_,
		_w3458_,
		_w3459_
	);
	LUT4 #(
		.INIT('h0d00)
	) name2997 (
		_w2292_,
		_w3452_,
		_w3453_,
		_w3459_,
		_w3460_
	);
	LUT4 #(
		.INIT('ha0a8)
	) name2998 (
		\P1_state_reg[0]/NET0131 ,
		_w1731_,
		_w3451_,
		_w3460_,
		_w3461_
	);
	LUT2 #(
		.INIT('he)
	) name2999 (
		_w3450_,
		_w3461_,
		_w3462_
	);
	LUT4 #(
		.INIT('h4000)
	) name3000 (
		_w1723_,
		_w1727_,
		_w1730_,
		_w2197_,
		_w3463_
	);
	LUT2 #(
		.INIT('h2)
	) name3001 (
		_w2197_,
		_w2644_,
		_w3464_
	);
	LUT4 #(
		.INIT('h1000)
	) name3002 (
		_w2187_,
		_w2235_,
		_w2404_,
		_w2408_,
		_w3465_
	);
	LUT4 #(
		.INIT('h4144)
	) name3003 (
		_w1747_,
		_w2175_,
		_w2200_,
		_w3465_,
		_w3466_
	);
	LUT3 #(
		.INIT('h80)
	) name3004 (
		_w1747_,
		_w2184_,
		_w2186_,
		_w3467_
	);
	LUT4 #(
		.INIT('h3331)
	) name3005 (
		_w2644_,
		_w3464_,
		_w3466_,
		_w3467_,
		_w3468_
	);
	LUT2 #(
		.INIT('h2)
	) name3006 (
		_w2424_,
		_w3468_,
		_w3469_
	);
	LUT4 #(
		.INIT('h007d)
	) name3007 (
		_w2644_,
		_w2958_,
		_w3181_,
		_w3464_,
		_w3470_
	);
	LUT2 #(
		.INIT('h2)
	) name3008 (
		_w2292_,
		_w3470_,
		_w3471_
	);
	LUT4 #(
		.INIT('h00d7)
	) name3009 (
		_w2644_,
		_w2940_,
		_w3181_,
		_w3464_,
		_w3472_
	);
	LUT4 #(
		.INIT('had88)
	) name3010 (
		_w2196_,
		_w2426_,
		_w2436_,
		_w2447_,
		_w3473_
	);
	LUT2 #(
		.INIT('h8)
	) name3011 (
		_w2196_,
		_w2454_,
		_w3474_
	);
	LUT3 #(
		.INIT('h51)
	) name3012 (
		_w2450_,
		_w2452_,
		_w2644_,
		_w3475_
	);
	LUT4 #(
		.INIT('h88a8)
	) name3013 (
		_w2197_,
		_w2450_,
		_w2452_,
		_w2644_,
		_w3476_
	);
	LUT2 #(
		.INIT('h1)
	) name3014 (
		_w3474_,
		_w3476_,
		_w3477_
	);
	LUT3 #(
		.INIT('h70)
	) name3015 (
		_w2644_,
		_w3473_,
		_w3477_,
		_w3478_
	);
	LUT3 #(
		.INIT('hd0)
	) name3016 (
		_w2388_,
		_w3472_,
		_w3478_,
		_w3479_
	);
	LUT4 #(
		.INIT('ha8aa)
	) name3017 (
		_w1731_,
		_w3469_,
		_w3471_,
		_w3479_,
		_w3480_
	);
	LUT2 #(
		.INIT('h2)
	) name3018 (
		\P1_reg3_reg[18]/NET0131 ,
		\P1_state_reg[0]/NET0131 ,
		_w3481_
	);
	LUT3 #(
		.INIT('h07)
	) name3019 (
		_w2197_,
		_w2695_,
		_w3481_,
		_w3482_
	);
	LUT4 #(
		.INIT('ha8ff)
	) name3020 (
		\P1_state_reg[0]/NET0131 ,
		_w3463_,
		_w3480_,
		_w3482_,
		_w3483_
	);
	LUT4 #(
		.INIT('h4000)
	) name3021 (
		_w1723_,
		_w1727_,
		_w1730_,
		_w2185_,
		_w3484_
	);
	LUT2 #(
		.INIT('h2)
	) name3022 (
		_w2185_,
		_w2644_,
		_w3485_
	);
	LUT4 #(
		.INIT('h7500)
	) name3023 (
		_w2301_,
		_w2327_,
		_w2330_,
		_w2353_,
		_w3486_
	);
	LUT4 #(
		.INIT('hc048)
	) name3024 (
		_w2336_,
		_w2644_,
		_w3170_,
		_w3486_,
		_w3487_
	);
	LUT3 #(
		.INIT('ha8)
	) name3025 (
		_w2388_,
		_w3485_,
		_w3487_,
		_w3488_
	);
	LUT4 #(
		.INIT('h2f00)
	) name3026 (
		_w2049_,
		_w2153_,
		_w2249_,
		_w2253_,
		_w3489_
	);
	LUT4 #(
		.INIT('h070d)
	) name3027 (
		_w2644_,
		_w3170_,
		_w3485_,
		_w3489_,
		_w3490_
	);
	LUT3 #(
		.INIT('h80)
	) name3028 (
		_w1747_,
		_w2232_,
		_w2234_,
		_w3491_
	);
	LUT4 #(
		.INIT('h00eb)
	) name3029 (
		_w1747_,
		_w2200_,
		_w3465_,
		_w3491_,
		_w3492_
	);
	LUT4 #(
		.INIT('hc808)
	) name3030 (
		_w2185_,
		_w2424_,
		_w2644_,
		_w3492_,
		_w3493_
	);
	LUT4 #(
		.INIT('h4000)
	) name3031 (
		_w2208_,
		_w2431_,
		_w2432_,
		_w2434_,
		_w3494_
	);
	LUT4 #(
		.INIT('ha8aa)
	) name3032 (
		_w2183_,
		_w2231_,
		_w2242_,
		_w3494_,
		_w3495_
	);
	LUT4 #(
		.INIT('h0040)
	) name3033 (
		_w2436_,
		_w2447_,
		_w2644_,
		_w3495_,
		_w3496_
	);
	LUT4 #(
		.INIT('ha8a0)
	) name3034 (
		_w2183_,
		_w2426_,
		_w2454_,
		_w2644_,
		_w3497_
	);
	LUT3 #(
		.INIT('h0d)
	) name3035 (
		_w2185_,
		_w2690_,
		_w3497_,
		_w3498_
	);
	LUT2 #(
		.INIT('h4)
	) name3036 (
		_w3496_,
		_w3498_,
		_w3499_
	);
	LUT4 #(
		.INIT('h0d00)
	) name3037 (
		_w2292_,
		_w3490_,
		_w3493_,
		_w3499_,
		_w3500_
	);
	LUT4 #(
		.INIT('h1311)
	) name3038 (
		_w1731_,
		_w3484_,
		_w3488_,
		_w3500_,
		_w3501_
	);
	LUT2 #(
		.INIT('h2)
	) name3039 (
		\P1_reg3_reg[17]/NET0131 ,
		\P1_state_reg[0]/NET0131 ,
		_w3502_
	);
	LUT3 #(
		.INIT('h07)
	) name3040 (
		_w2185_,
		_w2695_,
		_w3502_,
		_w3503_
	);
	LUT3 #(
		.INIT('h2f)
	) name3041 (
		\P1_state_reg[0]/NET0131 ,
		_w3501_,
		_w3503_,
		_w3504_
	);
	LUT4 #(
		.INIT('h4000)
	) name3042 (
		_w1723_,
		_w1727_,
		_w1730_,
		_w2172_,
		_w3505_
	);
	LUT2 #(
		.INIT('h2)
	) name3043 (
		_w2172_,
		_w2644_,
		_w3506_
	);
	LUT4 #(
		.INIT('ha8aa)
	) name3044 (
		_w2163_,
		_w2175_,
		_w2200_,
		_w3465_,
		_w3507_
	);
	LUT2 #(
		.INIT('h8)
	) name3045 (
		_w2392_,
		_w3465_,
		_w3508_
	);
	LUT3 #(
		.INIT('h80)
	) name3046 (
		_w1747_,
		_w2198_,
		_w2199_,
		_w3509_
	);
	LUT4 #(
		.INIT('h00ab)
	) name3047 (
		_w1747_,
		_w3507_,
		_w3508_,
		_w3509_,
		_w3510_
	);
	LUT4 #(
		.INIT('hc808)
	) name3048 (
		_w2172_,
		_w2424_,
		_w2644_,
		_w3510_,
		_w3511_
	);
	LUT4 #(
		.INIT('h00d7)
	) name3049 (
		_w2644_,
		_w2662_,
		_w3165_,
		_w3506_,
		_w3512_
	);
	LUT2 #(
		.INIT('h2)
	) name3050 (
		_w2292_,
		_w3512_,
		_w3513_
	);
	LUT4 #(
		.INIT('h007d)
	) name3051 (
		_w2644_,
		_w2675_,
		_w3165_,
		_w3506_,
		_w3514_
	);
	LUT4 #(
		.INIT('h2300)
	) name3052 (
		_w1748_,
		_w2168_,
		_w2170_,
		_w2426_,
		_w3515_
	);
	LUT4 #(
		.INIT('h6500)
	) name3053 (
		_w2171_,
		_w2196_,
		_w2436_,
		_w2447_,
		_w3516_
	);
	LUT4 #(
		.INIT('h2300)
	) name3054 (
		_w1748_,
		_w2168_,
		_w2170_,
		_w2454_,
		_w3517_
	);
	LUT4 #(
		.INIT('h88a8)
	) name3055 (
		_w2172_,
		_w2450_,
		_w2452_,
		_w2644_,
		_w3518_
	);
	LUT2 #(
		.INIT('h1)
	) name3056 (
		_w3517_,
		_w3518_,
		_w3519_
	);
	LUT4 #(
		.INIT('h5700)
	) name3057 (
		_w2644_,
		_w3515_,
		_w3516_,
		_w3519_,
		_w3520_
	);
	LUT3 #(
		.INIT('hd0)
	) name3058 (
		_w2388_,
		_w3514_,
		_w3520_,
		_w3521_
	);
	LUT4 #(
		.INIT('ha8aa)
	) name3059 (
		_w1731_,
		_w3511_,
		_w3513_,
		_w3521_,
		_w3522_
	);
	LUT2 #(
		.INIT('h2)
	) name3060 (
		\P1_reg3_reg[19]/NET0131 ,
		\P1_state_reg[0]/NET0131 ,
		_w3523_
	);
	LUT3 #(
		.INIT('h07)
	) name3061 (
		_w2172_,
		_w2695_,
		_w3523_,
		_w3524_
	);
	LUT4 #(
		.INIT('ha8ff)
	) name3062 (
		\P1_state_reg[0]/NET0131 ,
		_w3505_,
		_w3522_,
		_w3524_,
		_w3525_
	);
	LUT4 #(
		.INIT('h1000)
	) name3063 (
		_w863_,
		_w1189_,
		_w1352_,
		_w1356_,
		_w3526_
	);
	LUT4 #(
		.INIT('h0155)
	) name3064 (
		_w863_,
		_w1361_,
		_w1363_,
		_w1368_,
		_w3527_
	);
	LUT4 #(
		.INIT('h4f00)
	) name3065 (
		_w1537_,
		_w1539_,
		_w1543_,
		_w1547_,
		_w3528_
	);
	LUT4 #(
		.INIT('h8848)
	) name3066 (
		_w1294_,
		_w1369_,
		_w1553_,
		_w3528_,
		_w3529_
	);
	LUT3 #(
		.INIT('h54)
	) name3067 (
		_w1496_,
		_w3527_,
		_w3529_,
		_w3530_
	);
	LUT4 #(
		.INIT('h5554)
	) name3068 (
		_w863_,
		_w1361_,
		_w1363_,
		_w1368_,
		_w3531_
	);
	LUT4 #(
		.INIT('h8848)
	) name3069 (
		_w1294_,
		_w1411_,
		_w1553_,
		_w3528_,
		_w3532_
	);
	LUT3 #(
		.INIT('ha8)
	) name3070 (
		_w1447_,
		_w3531_,
		_w3532_,
		_w3533_
	);
	LUT4 #(
		.INIT('h4b00)
	) name3071 (
		_w1217_,
		_w1206_,
		_w1294_,
		_w1369_,
		_w3534_
	);
	LUT3 #(
		.INIT('h54)
	) name3072 (
		_w1409_,
		_w3527_,
		_w3534_,
		_w3535_
	);
	LUT2 #(
		.INIT('h1)
	) name3073 (
		_w528_,
		_w1435_,
		_w3536_
	);
	LUT4 #(
		.INIT('h006f)
	) name3074 (
		_w845_,
		_w1423_,
		_w1435_,
		_w3536_,
		_w3537_
	);
	LUT4 #(
		.INIT('h04c4)
	) name3075 (
		_w863_,
		_w1191_,
		_w1411_,
		_w3537_,
		_w3538_
	);
	LUT3 #(
		.INIT('h04)
	) name3076 (
		_w879_,
		_w1232_,
		_w1439_,
		_w3539_
	);
	LUT3 #(
		.INIT('h54)
	) name3077 (
		_w863_,
		_w1441_,
		_w1443_,
		_w3540_
	);
	LUT2 #(
		.INIT('h1)
	) name3078 (
		_w3539_,
		_w3540_,
		_w3541_
	);
	LUT2 #(
		.INIT('h4)
	) name3079 (
		_w3538_,
		_w3541_,
		_w3542_
	);
	LUT4 #(
		.INIT('h0100)
	) name3080 (
		_w3533_,
		_w3530_,
		_w3535_,
		_w3542_,
		_w3543_
	);
	LUT4 #(
		.INIT('ha0a8)
	) name3081 (
		\P1_state_reg[0]/NET0131 ,
		_w1359_,
		_w3526_,
		_w3543_,
		_w3544_
	);
	LUT4 #(
		.INIT('h0802)
	) name3082 (
		\P1_state_reg[0]/NET0131 ,
		\P2_IR_reg[23]/NET0131 ,
		_w863_,
		_w1188_,
		_w3545_
	);
	LUT2 #(
		.INIT('h4)
	) name3083 (
		\P1_state_reg[0]/NET0131 ,
		\P2_reg3_reg[16]/NET0131 ,
		_w3546_
	);
	LUT2 #(
		.INIT('h1)
	) name3084 (
		_w3545_,
		_w3546_,
		_w3547_
	);
	LUT2 #(
		.INIT('hb)
	) name3085 (
		_w3544_,
		_w3547_,
		_w3548_
	);
	LUT2 #(
		.INIT('h2)
	) name3086 (
		_w1950_,
		_w2644_,
		_w3549_
	);
	LUT4 #(
		.INIT('h00d7)
	) name3087 (
		_w2644_,
		_w2974_,
		_w2976_,
		_w3549_,
		_w3550_
	);
	LUT2 #(
		.INIT('h2)
	) name3088 (
		_w2388_,
		_w3550_,
		_w3551_
	);
	LUT4 #(
		.INIT('h007d)
	) name3089 (
		_w2644_,
		_w2974_,
		_w2982_,
		_w3549_,
		_w3552_
	);
	LUT4 #(
		.INIT('h00fd)
	) name3090 (
		_w2644_,
		_w2986_,
		_w2987_,
		_w3549_,
		_w3553_
	);
	LUT4 #(
		.INIT('h8040)
	) name3091 (
		_w1948_,
		_w2447_,
		_w2644_,
		_w2990_,
		_w3554_
	);
	LUT4 #(
		.INIT('hf531)
	) name3092 (
		_w1948_,
		_w1950_,
		_w2689_,
		_w2690_,
		_w3555_
	);
	LUT2 #(
		.INIT('h4)
	) name3093 (
		_w3554_,
		_w3555_,
		_w3556_
	);
	LUT3 #(
		.INIT('hd0)
	) name3094 (
		_w2424_,
		_w3553_,
		_w3556_,
		_w3557_
	);
	LUT3 #(
		.INIT('hd0)
	) name3095 (
		_w2292_,
		_w3552_,
		_w3557_,
		_w3558_
	);
	LUT4 #(
		.INIT('h4000)
	) name3096 (
		_w1723_,
		_w1727_,
		_w1730_,
		_w1950_,
		_w3559_
	);
	LUT4 #(
		.INIT('h0075)
	) name3097 (
		_w1731_,
		_w3551_,
		_w3558_,
		_w3559_,
		_w3560_
	);
	LUT2 #(
		.INIT('h2)
	) name3098 (
		\P1_reg3_reg[24]/NET0131 ,
		\P1_state_reg[0]/NET0131 ,
		_w3561_
	);
	LUT3 #(
		.INIT('h07)
	) name3099 (
		_w1950_,
		_w2695_,
		_w3561_,
		_w3562_
	);
	LUT3 #(
		.INIT('h2f)
	) name3100 (
		\P1_state_reg[0]/NET0131 ,
		_w3560_,
		_w3562_,
		_w3563_
	);
	LUT2 #(
		.INIT('h2)
	) name3101 (
		\P1_reg2_reg[31]/NET0131 ,
		_w2462_,
		_w3564_
	);
	LUT4 #(
		.INIT('h2000)
	) name3102 (
		\P1_reg2_reg[31]/NET0131 ,
		_w1723_,
		_w1727_,
		_w1730_,
		_w3565_
	);
	LUT4 #(
		.INIT('h0040)
	) name3103 (
		_w2273_,
		_w2443_,
		_w2444_,
		_w3135_,
		_w3566_
	);
	LUT4 #(
		.INIT('h1dd1)
	) name3104 (
		\P1_reg2_reg[31]/NET0131 ,
		_w1741_,
		_w3126_,
		_w3566_,
		_w3567_
	);
	LUT4 #(
		.INIT('h0777)
	) name3105 (
		_w2274_,
		_w2275_,
		_w2417_,
		_w2418_,
		_w3568_
	);
	LUT2 #(
		.INIT('h4)
	) name3106 (
		_w1836_,
		_w3568_,
		_w3569_
	);
	LUT3 #(
		.INIT('h15)
	) name3107 (
		_w2421_,
		_w2395_,
		_w2396_,
		_w3570_
	);
	LUT2 #(
		.INIT('h8)
	) name3108 (
		_w1741_,
		_w2424_,
		_w3571_
	);
	LUT4 #(
		.INIT('h7000)
	) name3109 (
		_w2922_,
		_w3569_,
		_w3570_,
		_w3571_,
		_w3572_
	);
	LUT4 #(
		.INIT('hd1dd)
	) name3110 (
		\P1_reg2_reg[31]/NET0131 ,
		_w1741_,
		_w1748_,
		_w3125_,
		_w3573_
	);
	LUT4 #(
		.INIT('h3133)
	) name3111 (
		_w1723_,
		_w2285_,
		_w2288_,
		_w2291_,
		_w3574_
	);
	LUT4 #(
		.INIT('ha0a2)
	) name3112 (
		\P1_reg2_reg[31]/NET0131 ,
		_w1741_,
		_w2450_,
		_w3574_,
		_w3575_
	);
	LUT2 #(
		.INIT('h1)
	) name3113 (
		_w2455_,
		_w3575_,
		_w3576_
	);
	LUT3 #(
		.INIT('hd0)
	) name3114 (
		_w2426_,
		_w3573_,
		_w3576_,
		_w3577_
	);
	LUT4 #(
		.INIT('h0d00)
	) name3115 (
		_w2447_,
		_w3567_,
		_w3572_,
		_w3577_,
		_w3578_
	);
	LUT4 #(
		.INIT('ha0a8)
	) name3116 (
		\P1_state_reg[0]/NET0131 ,
		_w1731_,
		_w3565_,
		_w3578_,
		_w3579_
	);
	LUT2 #(
		.INIT('he)
	) name3117 (
		_w3564_,
		_w3579_,
		_w3580_
	);
	LUT4 #(
		.INIT('hd070)
	) name3118 (
		\P1_state_reg[0]/NET0131 ,
		\P2_IR_reg[23]/NET0131 ,
		\P2_reg2_reg[23]/NET0131 ,
		_w1188_,
		_w3581_
	);
	LUT4 #(
		.INIT('h2000)
	) name3119 (
		\P2_reg2_reg[23]/NET0131 ,
		_w1189_,
		_w1352_,
		_w1356_,
		_w3582_
	);
	LUT4 #(
		.INIT('h6030)
	) name3120 (
		_w989_,
		_w1047_,
		_w1435_,
		_w2624_,
		_w3583_
	);
	LUT3 #(
		.INIT('h0b)
	) name3121 (
		_w1001_,
		_w1005_,
		_w1435_,
		_w3584_
	);
	LUT4 #(
		.INIT('h111d)
	) name3122 (
		\P2_reg2_reg[23]/NET0131 ,
		_w1516_,
		_w3583_,
		_w3584_,
		_w3585_
	);
	LUT2 #(
		.INIT('h2)
	) name3123 (
		_w1191_,
		_w3585_,
		_w3586_
	);
	LUT4 #(
		.INIT('ha8aa)
	) name3124 (
		\P2_reg2_reg[23]/NET0131 ,
		_w1361_,
		_w1363_,
		_w1368_,
		_w3587_
	);
	LUT2 #(
		.INIT('h8)
	) name3125 (
		_w1450_,
		_w1484_,
		_w3588_
	);
	LUT3 #(
		.INIT('hb0)
	) name3126 (
		_w1471_,
		_w1475_,
		_w3588_,
		_w3589_
	);
	LUT2 #(
		.INIT('h4)
	) name3127 (
		_w1478_,
		_w1484_,
		_w3590_
	);
	LUT2 #(
		.INIT('h2)
	) name3128 (
		_w1490_,
		_w3590_,
		_w3591_
	);
	LUT4 #(
		.INIT('h4844)
	) name3129 (
		_w1278_,
		_w1507_,
		_w3589_,
		_w3591_,
		_w3592_
	);
	LUT4 #(
		.INIT('h1000)
	) name3130 (
		_w546_,
		_w981_,
		_w1442_,
		_w1507_,
		_w3593_
	);
	LUT2 #(
		.INIT('h4)
	) name3131 (
		_w983_,
		_w1233_,
		_w3594_
	);
	LUT4 #(
		.INIT('h0057)
	) name3132 (
		\P2_reg2_reg[23]/NET0131 ,
		_w1441_,
		_w1523_,
		_w3594_,
		_w3595_
	);
	LUT2 #(
		.INIT('h4)
	) name3133 (
		_w3593_,
		_w3595_,
		_w3596_
	);
	LUT4 #(
		.INIT('hab00)
	) name3134 (
		_w1575_,
		_w3587_,
		_w3592_,
		_w3596_,
		_w3597_
	);
	LUT4 #(
		.INIT('h4f00)
	) name3135 (
		_w1379_,
		_w1383_,
		_w1386_,
		_w1390_,
		_w3598_
	);
	LUT2 #(
		.INIT('h8)
	) name3136 (
		_w1373_,
		_w1396_,
		_w3599_
	);
	LUT2 #(
		.INIT('h4)
	) name3137 (
		_w1393_,
		_w1396_,
		_w3600_
	);
	LUT4 #(
		.INIT('h008a)
	) name3138 (
		_w1403_,
		_w3598_,
		_w3599_,
		_w3600_,
		_w3601_
	);
	LUT4 #(
		.INIT('hc535)
	) name3139 (
		\P2_reg2_reg[23]/NET0131 ,
		_w1278_,
		_w1507_,
		_w3601_,
		_w3602_
	);
	LUT4 #(
		.INIT('hc535)
	) name3140 (
		\P2_reg2_reg[23]/NET0131 ,
		_w1278_,
		_w1516_,
		_w3601_,
		_w3603_
	);
	LUT4 #(
		.INIT('hfa32)
	) name3141 (
		_w1506_,
		_w1530_,
		_w3602_,
		_w3603_,
		_w3604_
	);
	LUT4 #(
		.INIT('h8aaa)
	) name3142 (
		_w1359_,
		_w3586_,
		_w3597_,
		_w3604_,
		_w3605_
	);
	LUT4 #(
		.INIT('heeec)
	) name3143 (
		\P1_state_reg[0]/NET0131 ,
		_w3581_,
		_w3582_,
		_w3605_,
		_w3606_
	);
	LUT2 #(
		.INIT('h4)
	) name3144 (
		_w983_,
		_w1357_,
		_w3607_
	);
	LUT4 #(
		.INIT('h5554)
	) name3145 (
		_w983_,
		_w1361_,
		_w1363_,
		_w1368_,
		_w3608_
	);
	LUT4 #(
		.INIT('h0057)
	) name3146 (
		_w1411_,
		_w3583_,
		_w3584_,
		_w3608_,
		_w3609_
	);
	LUT2 #(
		.INIT('h2)
	) name3147 (
		_w1191_,
		_w3609_,
		_w3610_
	);
	LUT4 #(
		.INIT('h4844)
	) name3148 (
		_w1278_,
		_w1411_,
		_w3589_,
		_w3591_,
		_w3611_
	);
	LUT3 #(
		.INIT('h54)
	) name3149 (
		_w983_,
		_w1441_,
		_w1443_,
		_w3612_
	);
	LUT4 #(
		.INIT('h0010)
	) name3150 (
		_w546_,
		_w981_,
		_w1232_,
		_w1439_,
		_w3613_
	);
	LUT2 #(
		.INIT('h1)
	) name3151 (
		_w3612_,
		_w3613_,
		_w3614_
	);
	LUT4 #(
		.INIT('h5700)
	) name3152 (
		_w1447_,
		_w3608_,
		_w3611_,
		_w3614_,
		_w3615_
	);
	LUT4 #(
		.INIT('h0155)
	) name3153 (
		_w983_,
		_w1361_,
		_w1363_,
		_w1368_,
		_w3616_
	);
	LUT4 #(
		.INIT('h00b7)
	) name3154 (
		_w1278_,
		_w1369_,
		_w3601_,
		_w3616_,
		_w3617_
	);
	LUT2 #(
		.INIT('h1)
	) name3155 (
		_w1409_,
		_w3617_,
		_w3618_
	);
	LUT4 #(
		.INIT('h4844)
	) name3156 (
		_w1278_,
		_w1369_,
		_w3589_,
		_w3591_,
		_w3619_
	);
	LUT3 #(
		.INIT('h54)
	) name3157 (
		_w1496_,
		_w3616_,
		_w3619_,
		_w3620_
	);
	LUT4 #(
		.INIT('h0100)
	) name3158 (
		_w3610_,
		_w3618_,
		_w3620_,
		_w3615_,
		_w3621_
	);
	LUT4 #(
		.INIT('ha0a8)
	) name3159 (
		\P1_state_reg[0]/NET0131 ,
		_w1359_,
		_w3607_,
		_w3621_,
		_w3622_
	);
	LUT2 #(
		.INIT('h4)
	) name3160 (
		\P1_state_reg[0]/NET0131 ,
		\P2_reg3_reg[23]/NET0131 ,
		_w3623_
	);
	LUT4 #(
		.INIT('h9c00)
	) name3161 (
		\P2_reg3_reg[22]/NET0131 ,
		\P2_reg3_reg[23]/NET0131 ,
		_w946_,
		_w1349_,
		_w3624_
	);
	LUT2 #(
		.INIT('h1)
	) name3162 (
		_w3623_,
		_w3624_,
		_w3625_
	);
	LUT2 #(
		.INIT('hb)
	) name3163 (
		_w3622_,
		_w3625_,
		_w3626_
	);
	LUT4 #(
		.INIT('h4000)
	) name3164 (
		_w1723_,
		_w1727_,
		_w1730_,
		_w1872_,
		_w3627_
	);
	LUT2 #(
		.INIT('h2)
	) name3165 (
		_w1872_,
		_w2644_,
		_w3628_
	);
	LUT4 #(
		.INIT('h2070)
	) name3166 (
		_w1747_,
		_w1952_,
		_w2644_,
		_w3005_,
		_w3629_
	);
	LUT3 #(
		.INIT('ha8)
	) name3167 (
		_w2424_,
		_w3628_,
		_w3629_,
		_w3630_
	);
	LUT4 #(
		.INIT('hc808)
	) name3168 (
		_w1872_,
		_w2447_,
		_w2644_,
		_w3008_,
		_w3631_
	);
	LUT4 #(
		.INIT('ha0a8)
	) name3169 (
		_w1872_,
		_w2426_,
		_w2450_,
		_w2644_,
		_w3632_
	);
	LUT3 #(
		.INIT('h0d)
	) name3170 (
		_w1871_,
		_w2689_,
		_w3632_,
		_w3633_
	);
	LUT2 #(
		.INIT('h4)
	) name3171 (
		_w3631_,
		_w3633_,
		_w3634_
	);
	LUT2 #(
		.INIT('h4)
	) name3172 (
		_w3630_,
		_w3634_,
		_w3635_
	);
	LUT4 #(
		.INIT('h08c8)
	) name3173 (
		_w1872_,
		_w2292_,
		_w2644_,
		_w3019_,
		_w3636_
	);
	LUT4 #(
		.INIT('h00d7)
	) name3174 (
		_w2644_,
		_w3016_,
		_w3025_,
		_w3628_,
		_w3637_
	);
	LUT3 #(
		.INIT('h31)
	) name3175 (
		_w2388_,
		_w3636_,
		_w3637_,
		_w3638_
	);
	LUT4 #(
		.INIT('h3111)
	) name3176 (
		_w1731_,
		_w3627_,
		_w3635_,
		_w3638_,
		_w3639_
	);
	LUT2 #(
		.INIT('h2)
	) name3177 (
		\P1_reg3_reg[25]/NET0131 ,
		\P1_state_reg[0]/NET0131 ,
		_w3640_
	);
	LUT3 #(
		.INIT('h07)
	) name3178 (
		_w1872_,
		_w2695_,
		_w3640_,
		_w3641_
	);
	LUT3 #(
		.INIT('h2f)
	) name3179 (
		\P1_state_reg[0]/NET0131 ,
		_w3639_,
		_w3641_,
		_w3642_
	);
	LUT4 #(
		.INIT('hd070)
	) name3180 (
		\P1_state_reg[0]/NET0131 ,
		\P2_IR_reg[23]/NET0131 ,
		\P2_reg0_reg[22]/NET0131 ,
		_w1188_,
		_w3643_
	);
	LUT4 #(
		.INIT('h2000)
	) name3181 (
		\P2_reg0_reg[22]/NET0131 ,
		_w1189_,
		_w1352_,
		_w1356_,
		_w3644_
	);
	LUT4 #(
		.INIT('h02aa)
	) name3182 (
		\P2_reg0_reg[22]/NET0131 ,
		_w1361_,
		_w1363_,
		_w1368_,
		_w3645_
	);
	LUT3 #(
		.INIT('ha8)
	) name3183 (
		_w1447_,
		_w2621_,
		_w3645_,
		_w3646_
	);
	LUT4 #(
		.INIT('haaa8)
	) name3184 (
		\P2_reg0_reg[22]/NET0131 ,
		_w1361_,
		_w1363_,
		_w1368_,
		_w3647_
	);
	LUT3 #(
		.INIT('h54)
	) name3185 (
		_w1496_,
		_w2618_,
		_w3647_,
		_w3648_
	);
	LUT4 #(
		.INIT('h08c8)
	) name3186 (
		\P2_reg0_reg[22]/NET0131 ,
		_w1191_,
		_w1369_,
		_w2626_,
		_w3649_
	);
	LUT4 #(
		.INIT('hc535)
	) name3187 (
		\P2_reg0_reg[22]/NET0131 ,
		_w1275_,
		_w1411_,
		_w2634_,
		_w3650_
	);
	LUT4 #(
		.INIT('h1000)
	) name3188 (
		_w546_,
		_w999_,
		_w1411_,
		_w1442_,
		_w3651_
	);
	LUT3 #(
		.INIT('ha2)
	) name3189 (
		\P2_reg0_reg[22]/NET0131 ,
		_w1684_,
		_w1685_,
		_w3652_
	);
	LUT2 #(
		.INIT('h1)
	) name3190 (
		_w3651_,
		_w3652_,
		_w3653_
	);
	LUT4 #(
		.INIT('h3200)
	) name3191 (
		_w1409_,
		_w3649_,
		_w3650_,
		_w3653_,
		_w3654_
	);
	LUT4 #(
		.INIT('ha8aa)
	) name3192 (
		_w1359_,
		_w3648_,
		_w3646_,
		_w3654_,
		_w3655_
	);
	LUT4 #(
		.INIT('heeec)
	) name3193 (
		\P1_state_reg[0]/NET0131 ,
		_w3643_,
		_w3644_,
		_w3655_,
		_w3656_
	);
	LUT2 #(
		.INIT('h2)
	) name3194 (
		\P1_reg2_reg[26]/NET0131 ,
		_w2462_,
		_w3657_
	);
	LUT4 #(
		.INIT('h2000)
	) name3195 (
		\P1_reg2_reg[26]/NET0131 ,
		_w1723_,
		_w1727_,
		_w1730_,
		_w3658_
	);
	LUT2 #(
		.INIT('h2)
	) name3196 (
		\P1_reg2_reg[26]/NET0131 ,
		_w1741_,
		_w3659_
	);
	LUT4 #(
		.INIT('h2a08)
	) name3197 (
		_w1741_,
		_w1747_,
		_w1876_,
		_w2923_,
		_w3660_
	);
	LUT4 #(
		.INIT('ha2a0)
	) name3198 (
		\P1_reg2_reg[26]/NET0131 ,
		_w1741_,
		_w2450_,
		_w2452_,
		_w3661_
	);
	LUT2 #(
		.INIT('h8)
	) name3199 (
		_w1901_,
		_w2454_,
		_w3662_
	);
	LUT2 #(
		.INIT('h1)
	) name3200 (
		_w3661_,
		_w3662_,
		_w3663_
	);
	LUT3 #(
		.INIT('hd0)
	) name3201 (
		_w1741_,
		_w3407_,
		_w3663_,
		_w3664_
	);
	LUT4 #(
		.INIT('h5700)
	) name3202 (
		_w2424_,
		_w3659_,
		_w3660_,
		_w3664_,
		_w3665_
	);
	LUT4 #(
		.INIT('h20e0)
	) name3203 (
		\P1_reg2_reg[26]/NET0131 ,
		_w1741_,
		_w2388_,
		_w2948_,
		_w3666_
	);
	LUT4 #(
		.INIT('h20e0)
	) name3204 (
		\P1_reg2_reg[26]/NET0131 ,
		_w1741_,
		_w2292_,
		_w2967_,
		_w3667_
	);
	LUT4 #(
		.INIT('ha8aa)
	) name3205 (
		_w1731_,
		_w3666_,
		_w3667_,
		_w3665_,
		_w3668_
	);
	LUT4 #(
		.INIT('heeec)
	) name3206 (
		\P1_state_reg[0]/NET0131 ,
		_w3657_,
		_w3658_,
		_w3668_,
		_w3669_
	);
	LUT4 #(
		.INIT('hd070)
	) name3207 (
		\P1_state_reg[0]/NET0131 ,
		\P2_IR_reg[23]/NET0131 ,
		\P2_reg1_reg[22]/NET0131 ,
		_w1188_,
		_w3670_
	);
	LUT4 #(
		.INIT('h2000)
	) name3208 (
		\P2_reg1_reg[22]/NET0131 ,
		_w1189_,
		_w1352_,
		_w1356_,
		_w3671_
	);
	LUT4 #(
		.INIT('h4484)
	) name3209 (
		_w1275_,
		_w1516_,
		_w2615_,
		_w2617_,
		_w3672_
	);
	LUT4 #(
		.INIT('haa02)
	) name3210 (
		\P2_reg1_reg[22]/NET0131 ,
		_w1361_,
		_w1363_,
		_w1368_,
		_w3673_
	);
	LUT3 #(
		.INIT('h54)
	) name3211 (
		_w1575_,
		_w3672_,
		_w3673_,
		_w3674_
	);
	LUT4 #(
		.INIT('h08c8)
	) name3212 (
		\P2_reg1_reg[22]/NET0131 ,
		_w1191_,
		_w1507_,
		_w2626_,
		_w3675_
	);
	LUT4 #(
		.INIT('hc535)
	) name3213 (
		\P2_reg1_reg[22]/NET0131 ,
		_w1275_,
		_w1507_,
		_w2634_,
		_w3676_
	);
	LUT2 #(
		.INIT('h2)
	) name3214 (
		_w1530_,
		_w3676_,
		_w3677_
	);
	LUT4 #(
		.INIT('hc535)
	) name3215 (
		\P2_reg1_reg[22]/NET0131 ,
		_w1275_,
		_w1516_,
		_w2634_,
		_w3678_
	);
	LUT4 #(
		.INIT('h1000)
	) name3216 (
		_w546_,
		_w999_,
		_w1442_,
		_w1516_,
		_w3679_
	);
	LUT3 #(
		.INIT('ha2)
	) name3217 (
		\P2_reg1_reg[22]/NET0131 ,
		_w1684_,
		_w2469_,
		_w3680_
	);
	LUT2 #(
		.INIT('h1)
	) name3218 (
		_w3679_,
		_w3680_,
		_w3681_
	);
	LUT3 #(
		.INIT('he0)
	) name3219 (
		_w1506_,
		_w3678_,
		_w3681_,
		_w3682_
	);
	LUT4 #(
		.INIT('h0100)
	) name3220 (
		_w3674_,
		_w3675_,
		_w3677_,
		_w3682_,
		_w3683_
	);
	LUT4 #(
		.INIT('ha0a8)
	) name3221 (
		\P1_state_reg[0]/NET0131 ,
		_w1359_,
		_w3671_,
		_w3683_,
		_w3684_
	);
	LUT2 #(
		.INIT('he)
	) name3222 (
		_w3670_,
		_w3684_,
		_w3685_
	);
	LUT2 #(
		.INIT('h2)
	) name3223 (
		\P1_reg0_reg[22]/NET0131 ,
		_w2462_,
		_w3686_
	);
	LUT4 #(
		.INIT('h2000)
	) name3224 (
		\P1_reg0_reg[22]/NET0131 ,
		_w1723_,
		_w1727_,
		_w1730_,
		_w3687_
	);
	LUT2 #(
		.INIT('h2)
	) name3225 (
		\P1_reg0_reg[22]/NET0131 ,
		_w2883_,
		_w3688_
	);
	LUT4 #(
		.INIT('h1444)
	) name3226 (
		_w1747_,
		_w1962_,
		_w2919_,
		_w2921_,
		_w3689_
	);
	LUT3 #(
		.INIT('h80)
	) name3227 (
		_w1747_,
		_w1984_,
		_w1986_,
		_w3690_
	);
	LUT4 #(
		.INIT('hddd1)
	) name3228 (
		\P1_reg0_reg[22]/NET0131 ,
		_w2883_,
		_w3689_,
		_w3690_,
		_w3691_
	);
	LUT4 #(
		.INIT('h5400)
	) name3229 (
		_w1748_,
		_w1966_,
		_w1970_,
		_w2426_,
		_w3692_
	);
	LUT4 #(
		.INIT('h6555)
	) name3230 (
		_w1971_,
		_w1983_,
		_w2436_,
		_w2438_,
		_w3693_
	);
	LUT4 #(
		.INIT('hc8c0)
	) name3231 (
		_w2447_,
		_w2883_,
		_w3692_,
		_w3693_,
		_w3694_
	);
	LUT4 #(
		.INIT('h0a8a)
	) name3232 (
		\P1_reg0_reg[22]/NET0131 ,
		_w2452_,
		_w2524_,
		_w2883_,
		_w3695_
	);
	LUT2 #(
		.INIT('h1)
	) name3233 (
		_w3694_,
		_w3695_,
		_w3696_
	);
	LUT3 #(
		.INIT('hd0)
	) name3234 (
		_w2424_,
		_w3691_,
		_w3696_,
		_w3697_
	);
	LUT2 #(
		.INIT('h8)
	) name3235 (
		_w2950_,
		_w2959_,
		_w3698_
	);
	LUT4 #(
		.INIT('h4f00)
	) name3236 (
		_w2953_,
		_w2954_,
		_w2955_,
		_w3698_,
		_w3699_
	);
	LUT2 #(
		.INIT('h4)
	) name3237 (
		_w2956_,
		_w2959_,
		_w3700_
	);
	LUT2 #(
		.INIT('h2)
	) name3238 (
		_w2962_,
		_w3700_,
		_w3701_
	);
	LUT4 #(
		.INIT('h2822)
	) name3239 (
		_w2883_,
		_w3166_,
		_w3699_,
		_w3701_,
		_w3702_
	);
	LUT3 #(
		.INIT('ha8)
	) name3240 (
		_w2292_,
		_w3688_,
		_w3702_,
		_w3703_
	);
	LUT2 #(
		.INIT('h8)
	) name3241 (
		_w2931_,
		_w2942_,
		_w3704_
	);
	LUT4 #(
		.INIT('h4f00)
	) name3242 (
		_w2935_,
		_w2936_,
		_w2937_,
		_w3704_,
		_w3705_
	);
	LUT2 #(
		.INIT('h4)
	) name3243 (
		_w2938_,
		_w2942_,
		_w3706_
	);
	LUT2 #(
		.INIT('h2)
	) name3244 (
		_w2944_,
		_w3706_,
		_w3707_
	);
	LUT4 #(
		.INIT('h8288)
	) name3245 (
		_w2883_,
		_w3166_,
		_w3705_,
		_w3707_,
		_w3708_
	);
	LUT3 #(
		.INIT('ha8)
	) name3246 (
		_w2388_,
		_w3688_,
		_w3708_,
		_w3709_
	);
	LUT4 #(
		.INIT('ha8aa)
	) name3247 (
		_w1731_,
		_w3703_,
		_w3709_,
		_w3697_,
		_w3710_
	);
	LUT4 #(
		.INIT('heeec)
	) name3248 (
		\P1_state_reg[0]/NET0131 ,
		_w3686_,
		_w3687_,
		_w3710_,
		_w3711_
	);
	LUT2 #(
		.INIT('h2)
	) name3249 (
		\P1_reg0_reg[25]/NET0131 ,
		_w2462_,
		_w3712_
	);
	LUT4 #(
		.INIT('h2000)
	) name3250 (
		\P1_reg0_reg[25]/NET0131 ,
		_w1723_,
		_w1727_,
		_w1730_,
		_w3713_
	);
	LUT2 #(
		.INIT('h2)
	) name3251 (
		\P1_reg0_reg[25]/NET0131 ,
		_w2883_,
		_w3714_
	);
	LUT4 #(
		.INIT('h2070)
	) name3252 (
		_w1747_,
		_w1952_,
		_w2883_,
		_w3005_,
		_w3715_
	);
	LUT3 #(
		.INIT('ha8)
	) name3253 (
		_w2424_,
		_w3714_,
		_w3715_,
		_w3716_
	);
	LUT4 #(
		.INIT('hc808)
	) name3254 (
		\P1_reg0_reg[25]/NET0131 ,
		_w2447_,
		_w2883_,
		_w3008_,
		_w3717_
	);
	LUT4 #(
		.INIT('h0a8a)
	) name3255 (
		\P1_reg0_reg[25]/NET0131 ,
		_w2426_,
		_w2524_,
		_w2883_,
		_w3718_
	);
	LUT3 #(
		.INIT('h07)
	) name3256 (
		_w2883_,
		_w3010_,
		_w3718_,
		_w3719_
	);
	LUT2 #(
		.INIT('h4)
	) name3257 (
		_w3717_,
		_w3719_,
		_w3720_
	);
	LUT2 #(
		.INIT('h4)
	) name3258 (
		_w3716_,
		_w3720_,
		_w3721_
	);
	LUT4 #(
		.INIT('h08c8)
	) name3259 (
		\P1_reg0_reg[25]/NET0131 ,
		_w2292_,
		_w2883_,
		_w3019_,
		_w3722_
	);
	LUT4 #(
		.INIT('hd11d)
	) name3260 (
		\P1_reg0_reg[25]/NET0131 ,
		_w2883_,
		_w3016_,
		_w3025_,
		_w3723_
	);
	LUT3 #(
		.INIT('h31)
	) name3261 (
		_w2388_,
		_w3722_,
		_w3723_,
		_w3724_
	);
	LUT4 #(
		.INIT('h3111)
	) name3262 (
		_w1731_,
		_w3713_,
		_w3721_,
		_w3724_,
		_w3725_
	);
	LUT3 #(
		.INIT('hce)
	) name3263 (
		\P1_state_reg[0]/NET0131 ,
		_w3712_,
		_w3725_,
		_w3726_
	);
	LUT4 #(
		.INIT('hd11d)
	) name3264 (
		\P1_reg0_reg[24]/NET0131 ,
		_w2883_,
		_w2974_,
		_w2976_,
		_w3727_
	);
	LUT2 #(
		.INIT('h2)
	) name3265 (
		_w2388_,
		_w3727_,
		_w3728_
	);
	LUT4 #(
		.INIT('h1dd1)
	) name3266 (
		\P1_reg0_reg[24]/NET0131 ,
		_w2883_,
		_w2974_,
		_w2982_,
		_w3729_
	);
	LUT4 #(
		.INIT('hddd1)
	) name3267 (
		\P1_reg0_reg[24]/NET0131 ,
		_w2883_,
		_w2986_,
		_w2987_,
		_w3730_
	);
	LUT2 #(
		.INIT('h2)
	) name3268 (
		\P1_reg0_reg[24]/NET0131 ,
		_w3420_,
		_w3731_
	);
	LUT3 #(
		.INIT('h0d)
	) name3269 (
		_w2883_,
		_w2991_,
		_w3731_,
		_w3732_
	);
	LUT3 #(
		.INIT('hd0)
	) name3270 (
		_w2424_,
		_w3730_,
		_w3732_,
		_w3733_
	);
	LUT3 #(
		.INIT('hd0)
	) name3271 (
		_w2292_,
		_w3729_,
		_w3733_,
		_w3734_
	);
	LUT4 #(
		.INIT('h2000)
	) name3272 (
		\P1_reg0_reg[24]/NET0131 ,
		_w1723_,
		_w1727_,
		_w1730_,
		_w3735_
	);
	LUT4 #(
		.INIT('h0075)
	) name3273 (
		_w1731_,
		_w3728_,
		_w3734_,
		_w3735_,
		_w3736_
	);
	LUT2 #(
		.INIT('h2)
	) name3274 (
		\P1_reg0_reg[24]/NET0131 ,
		_w2462_,
		_w3737_
	);
	LUT3 #(
		.INIT('hf2)
	) name3275 (
		\P1_state_reg[0]/NET0131 ,
		_w3736_,
		_w3737_,
		_w3738_
	);
	LUT2 #(
		.INIT('h2)
	) name3276 (
		\P1_reg1_reg[22]/NET0131 ,
		_w2462_,
		_w3739_
	);
	LUT4 #(
		.INIT('h2000)
	) name3277 (
		\P1_reg1_reg[22]/NET0131 ,
		_w1723_,
		_w1727_,
		_w1730_,
		_w3740_
	);
	LUT2 #(
		.INIT('h2)
	) name3278 (
		\P1_reg1_reg[22]/NET0131 ,
		_w2520_,
		_w3741_
	);
	LUT4 #(
		.INIT('hddd1)
	) name3279 (
		\P1_reg1_reg[22]/NET0131 ,
		_w2520_,
		_w3689_,
		_w3690_,
		_w3742_
	);
	LUT4 #(
		.INIT('hc8c0)
	) name3280 (
		_w2447_,
		_w2520_,
		_w3692_,
		_w3693_,
		_w3743_
	);
	LUT3 #(
		.INIT('hd0)
	) name3281 (
		_w2452_,
		_w2520_,
		_w2524_,
		_w3744_
	);
	LUT4 #(
		.INIT('h08aa)
	) name3282 (
		\P1_reg1_reg[22]/NET0131 ,
		_w2452_,
		_w2520_,
		_w2524_,
		_w3745_
	);
	LUT2 #(
		.INIT('h1)
	) name3283 (
		_w3743_,
		_w3745_,
		_w3746_
	);
	LUT3 #(
		.INIT('hd0)
	) name3284 (
		_w2424_,
		_w3742_,
		_w3746_,
		_w3747_
	);
	LUT4 #(
		.INIT('h8288)
	) name3285 (
		_w2520_,
		_w3166_,
		_w3705_,
		_w3707_,
		_w3748_
	);
	LUT3 #(
		.INIT('ha8)
	) name3286 (
		_w2388_,
		_w3741_,
		_w3748_,
		_w3749_
	);
	LUT4 #(
		.INIT('h2822)
	) name3287 (
		_w2520_,
		_w3166_,
		_w3699_,
		_w3701_,
		_w3750_
	);
	LUT3 #(
		.INIT('ha8)
	) name3288 (
		_w2292_,
		_w3741_,
		_w3750_,
		_w3751_
	);
	LUT4 #(
		.INIT('ha8aa)
	) name3289 (
		_w1731_,
		_w3749_,
		_w3751_,
		_w3747_,
		_w3752_
	);
	LUT4 #(
		.INIT('heeec)
	) name3290 (
		\P1_state_reg[0]/NET0131 ,
		_w3739_,
		_w3740_,
		_w3752_,
		_w3753_
	);
	LUT2 #(
		.INIT('h2)
	) name3291 (
		\P1_reg1_reg[24]/NET0131 ,
		_w2520_,
		_w3754_
	);
	LUT4 #(
		.INIT('hd11d)
	) name3292 (
		\P1_reg1_reg[24]/NET0131 ,
		_w2520_,
		_w2974_,
		_w2976_,
		_w3755_
	);
	LUT2 #(
		.INIT('h2)
	) name3293 (
		_w2388_,
		_w3755_,
		_w3756_
	);
	LUT4 #(
		.INIT('h1dd1)
	) name3294 (
		\P1_reg1_reg[24]/NET0131 ,
		_w2520_,
		_w2974_,
		_w2982_,
		_w3757_
	);
	LUT4 #(
		.INIT('hddd1)
	) name3295 (
		\P1_reg1_reg[24]/NET0131 ,
		_w2520_,
		_w2986_,
		_w2987_,
		_w3758_
	);
	LUT4 #(
		.INIT('h35c5)
	) name3296 (
		\P1_reg1_reg[24]/NET0131 ,
		_w1948_,
		_w2520_,
		_w2990_,
		_w3759_
	);
	LUT2 #(
		.INIT('h2)
	) name3297 (
		\P1_reg1_reg[24]/NET0131 ,
		_w2524_,
		_w3760_
	);
	LUT4 #(
		.INIT('h5400)
	) name3298 (
		_w1748_,
		_w1941_,
		_w1947_,
		_w2520_,
		_w3761_
	);
	LUT4 #(
		.INIT('h0507)
	) name3299 (
		_w2426_,
		_w3754_,
		_w3760_,
		_w3761_,
		_w3762_
	);
	LUT3 #(
		.INIT('hd0)
	) name3300 (
		_w2447_,
		_w3759_,
		_w3762_,
		_w3763_
	);
	LUT3 #(
		.INIT('hd0)
	) name3301 (
		_w2424_,
		_w3758_,
		_w3763_,
		_w3764_
	);
	LUT3 #(
		.INIT('hd0)
	) name3302 (
		_w2292_,
		_w3757_,
		_w3764_,
		_w3765_
	);
	LUT4 #(
		.INIT('h2000)
	) name3303 (
		\P1_reg1_reg[24]/NET0131 ,
		_w1723_,
		_w1727_,
		_w1730_,
		_w3766_
	);
	LUT4 #(
		.INIT('h0075)
	) name3304 (
		_w1731_,
		_w3756_,
		_w3765_,
		_w3766_,
		_w3767_
	);
	LUT2 #(
		.INIT('h2)
	) name3305 (
		\P1_reg1_reg[24]/NET0131 ,
		_w2462_,
		_w3768_
	);
	LUT3 #(
		.INIT('hf2)
	) name3306 (
		\P1_state_reg[0]/NET0131 ,
		_w3767_,
		_w3768_,
		_w3769_
	);
	LUT2 #(
		.INIT('h2)
	) name3307 (
		\P1_reg1_reg[25]/NET0131 ,
		_w2462_,
		_w3770_
	);
	LUT4 #(
		.INIT('h2000)
	) name3308 (
		\P1_reg1_reg[25]/NET0131 ,
		_w1723_,
		_w1727_,
		_w1730_,
		_w3771_
	);
	LUT2 #(
		.INIT('h2)
	) name3309 (
		\P1_reg1_reg[25]/NET0131 ,
		_w2520_,
		_w3772_
	);
	LUT4 #(
		.INIT('h2070)
	) name3310 (
		_w1747_,
		_w1952_,
		_w2520_,
		_w3005_,
		_w3773_
	);
	LUT3 #(
		.INIT('ha8)
	) name3311 (
		_w2424_,
		_w3772_,
		_w3773_,
		_w3774_
	);
	LUT4 #(
		.INIT('hc808)
	) name3312 (
		\P1_reg1_reg[25]/NET0131 ,
		_w2447_,
		_w2520_,
		_w3008_,
		_w3775_
	);
	LUT4 #(
		.INIT('h08aa)
	) name3313 (
		\P1_reg1_reg[25]/NET0131 ,
		_w2426_,
		_w2520_,
		_w2524_,
		_w3776_
	);
	LUT3 #(
		.INIT('h07)
	) name3314 (
		_w2520_,
		_w3010_,
		_w3776_,
		_w3777_
	);
	LUT2 #(
		.INIT('h4)
	) name3315 (
		_w3775_,
		_w3777_,
		_w3778_
	);
	LUT2 #(
		.INIT('h4)
	) name3316 (
		_w3774_,
		_w3778_,
		_w3779_
	);
	LUT4 #(
		.INIT('h08c8)
	) name3317 (
		\P1_reg1_reg[25]/NET0131 ,
		_w2292_,
		_w2520_,
		_w3019_,
		_w3780_
	);
	LUT4 #(
		.INIT('hd11d)
	) name3318 (
		\P1_reg1_reg[25]/NET0131 ,
		_w2520_,
		_w3016_,
		_w3025_,
		_w3781_
	);
	LUT3 #(
		.INIT('h31)
	) name3319 (
		_w2388_,
		_w3780_,
		_w3781_,
		_w3782_
	);
	LUT4 #(
		.INIT('h3111)
	) name3320 (
		_w1731_,
		_w3771_,
		_w3779_,
		_w3782_,
		_w3783_
	);
	LUT3 #(
		.INIT('hce)
	) name3321 (
		\P1_state_reg[0]/NET0131 ,
		_w3770_,
		_w3783_,
		_w3784_
	);
	LUT2 #(
		.INIT('h2)
	) name3322 (
		\P1_reg1_reg[26]/NET0131 ,
		_w2462_,
		_w3785_
	);
	LUT4 #(
		.INIT('h2000)
	) name3323 (
		\P1_reg1_reg[26]/NET0131 ,
		_w1723_,
		_w1727_,
		_w1730_,
		_w3786_
	);
	LUT2 #(
		.INIT('h2)
	) name3324 (
		\P1_reg1_reg[26]/NET0131 ,
		_w2520_,
		_w3787_
	);
	LUT4 #(
		.INIT('h7020)
	) name3325 (
		_w1747_,
		_w1876_,
		_w2520_,
		_w2923_,
		_w3788_
	);
	LUT4 #(
		.INIT('h08aa)
	) name3326 (
		\P1_reg1_reg[26]/NET0131 ,
		_w2452_,
		_w2520_,
		_w2524_,
		_w3789_
	);
	LUT3 #(
		.INIT('h0d)
	) name3327 (
		_w2520_,
		_w3407_,
		_w3789_,
		_w3790_
	);
	LUT4 #(
		.INIT('h5700)
	) name3328 (
		_w2424_,
		_w3787_,
		_w3788_,
		_w3790_,
		_w3791_
	);
	LUT4 #(
		.INIT('h08c8)
	) name3329 (
		\P1_reg1_reg[26]/NET0131 ,
		_w2292_,
		_w2520_,
		_w2967_,
		_w3792_
	);
	LUT4 #(
		.INIT('h08c8)
	) name3330 (
		\P1_reg1_reg[26]/NET0131 ,
		_w2388_,
		_w2520_,
		_w2948_,
		_w3793_
	);
	LUT4 #(
		.INIT('ha8aa)
	) name3331 (
		_w1731_,
		_w3792_,
		_w3793_,
		_w3791_,
		_w3794_
	);
	LUT4 #(
		.INIT('heeec)
	) name3332 (
		\P1_state_reg[0]/NET0131 ,
		_w3785_,
		_w3786_,
		_w3794_,
		_w3795_
	);
	LUT4 #(
		.INIT('h4000)
	) name3333 (
		_w1723_,
		_w1727_,
		_w1730_,
		_w2018_,
		_w3796_
	);
	LUT2 #(
		.INIT('h2)
	) name3334 (
		_w2018_,
		_w2644_,
		_w3797_
	);
	LUT4 #(
		.INIT('hb04f)
	) name3335 (
		_w2752_,
		_w2755_,
		_w2758_,
		_w3173_,
		_w3798_
	);
	LUT4 #(
		.INIT('hc808)
	) name3336 (
		_w2018_,
		_w2292_,
		_w2644_,
		_w3798_,
		_w3799_
	);
	LUT4 #(
		.INIT('h1444)
	) name3337 (
		_w1747_,
		_w2223_,
		_w2404_,
		_w2406_,
		_w3800_
	);
	LUT3 #(
		.INIT('h80)
	) name3338 (
		_w1747_,
		_w2006_,
		_w2007_,
		_w3801_
	);
	LUT4 #(
		.INIT('h3331)
	) name3339 (
		_w2644_,
		_w3797_,
		_w3800_,
		_w3801_,
		_w3802_
	);
	LUT2 #(
		.INIT('h2)
	) name3340 (
		_w2424_,
		_w3802_,
		_w3803_
	);
	LUT4 #(
		.INIT('h0100)
	) name3341 (
		_w2029_,
		_w2040_,
		_w2104_,
		_w2431_,
		_w3804_
	);
	LUT4 #(
		.INIT('h6030)
	) name3342 (
		_w2004_,
		_w2016_,
		_w2447_,
		_w3804_,
		_w3805_
	);
	LUT2 #(
		.INIT('h8)
	) name3343 (
		_w2644_,
		_w3805_,
		_w3806_
	);
	LUT4 #(
		.INIT('h00d7)
	) name3344 (
		_w2644_,
		_w2807_,
		_w3173_,
		_w3797_,
		_w3807_
	);
	LUT4 #(
		.INIT('ha8a0)
	) name3345 (
		_w2016_,
		_w2426_,
		_w2454_,
		_w2644_,
		_w3808_
	);
	LUT3 #(
		.INIT('h0d)
	) name3346 (
		_w2018_,
		_w2690_,
		_w3808_,
		_w3809_
	);
	LUT4 #(
		.INIT('h0d00)
	) name3347 (
		_w2388_,
		_w3807_,
		_w3806_,
		_w3809_,
		_w3810_
	);
	LUT4 #(
		.INIT('ha8aa)
	) name3348 (
		_w1731_,
		_w3799_,
		_w3803_,
		_w3810_,
		_w3811_
	);
	LUT2 #(
		.INIT('h2)
	) name3349 (
		\P1_reg3_reg[12]/NET0131 ,
		\P1_state_reg[0]/NET0131 ,
		_w3812_
	);
	LUT3 #(
		.INIT('h07)
	) name3350 (
		_w2018_,
		_w2695_,
		_w3812_,
		_w3813_
	);
	LUT4 #(
		.INIT('ha8ff)
	) name3351 (
		\P1_state_reg[0]/NET0131 ,
		_w3796_,
		_w3811_,
		_w3813_,
		_w3814_
	);
	LUT4 #(
		.INIT('h4000)
	) name3352 (
		_w1723_,
		_w1727_,
		_w1730_,
		_w2233_,
		_w3815_
	);
	LUT2 #(
		.INIT('h2)
	) name3353 (
		_w2233_,
		_w2644_,
		_w3816_
	);
	LUT4 #(
		.INIT('h4f00)
	) name3354 (
		_w2752_,
		_w2755_,
		_w2758_,
		_w2761_,
		_w3817_
	);
	LUT4 #(
		.INIT('h0a82)
	) name3355 (
		_w2644_,
		_w2768_,
		_w3168_,
		_w3817_,
		_w3818_
	);
	LUT3 #(
		.INIT('ha8)
	) name3356 (
		_w2292_,
		_w3816_,
		_w3818_,
		_w3819_
	);
	LUT4 #(
		.INIT('hb04f)
	) name3357 (
		_w2807_,
		_w2810_,
		_w2815_,
		_w3168_,
		_w3820_
	);
	LUT4 #(
		.INIT('h08c8)
	) name3358 (
		_w2233_,
		_w2388_,
		_w2644_,
		_w3820_,
		_w3821_
	);
	LUT4 #(
		.INIT('h6555)
	) name3359 (
		_w2187_,
		_w2235_,
		_w2404_,
		_w2408_,
		_w3822_
	);
	LUT4 #(
		.INIT('h7020)
	) name3360 (
		_w1747_,
		_w2246_,
		_w2644_,
		_w3822_,
		_w3823_
	);
	LUT4 #(
		.INIT('h6050)
	) name3361 (
		_w2231_,
		_w2242_,
		_w2447_,
		_w3494_,
		_w3824_
	);
	LUT4 #(
		.INIT('ha8a0)
	) name3362 (
		_w2231_,
		_w2426_,
		_w2454_,
		_w2644_,
		_w3825_
	);
	LUT3 #(
		.INIT('h0d)
	) name3363 (
		_w2233_,
		_w2690_,
		_w3825_,
		_w3826_
	);
	LUT3 #(
		.INIT('h70)
	) name3364 (
		_w2644_,
		_w3824_,
		_w3826_,
		_w3827_
	);
	LUT4 #(
		.INIT('h5700)
	) name3365 (
		_w2424_,
		_w3816_,
		_w3823_,
		_w3827_,
		_w3828_
	);
	LUT2 #(
		.INIT('h4)
	) name3366 (
		_w3821_,
		_w3828_,
		_w3829_
	);
	LUT4 #(
		.INIT('h1311)
	) name3367 (
		_w1731_,
		_w3815_,
		_w3819_,
		_w3829_,
		_w3830_
	);
	LUT2 #(
		.INIT('h2)
	) name3368 (
		\P1_reg3_reg[16]/NET0131 ,
		\P1_state_reg[0]/NET0131 ,
		_w3831_
	);
	LUT3 #(
		.INIT('h07)
	) name3369 (
		_w2233_,
		_w2695_,
		_w3831_,
		_w3832_
	);
	LUT3 #(
		.INIT('h2f)
	) name3370 (
		\P1_state_reg[0]/NET0131 ,
		_w3830_,
		_w3832_,
		_w3833_
	);
	LUT2 #(
		.INIT('h2)
	) name3371 (
		_w1985_,
		_w2644_,
		_w3834_
	);
	LUT4 #(
		.INIT('h0c8c)
	) name3372 (
		_w2336_,
		_w2347_,
		_w2351_,
		_w3486_,
		_w3835_
	);
	LUT4 #(
		.INIT('h0d07)
	) name3373 (
		_w2644_,
		_w3160_,
		_w3834_,
		_w3835_,
		_w3836_
	);
	LUT4 #(
		.INIT('h007b)
	) name3374 (
		_w2262_,
		_w2644_,
		_w3160_,
		_w3834_,
		_w3837_
	);
	LUT4 #(
		.INIT('h9555)
	) name3375 (
		_w1975_,
		_w2394_,
		_w2404_,
		_w2408_,
		_w3838_
	);
	LUT4 #(
		.INIT('h0200)
	) name3376 (
		_w1747_,
		_w2161_,
		_w2160_,
		_w2162_,
		_w3839_
	);
	LUT2 #(
		.INIT('h2)
	) name3377 (
		_w2424_,
		_w3839_,
		_w3840_
	);
	LUT4 #(
		.INIT('h9500)
	) name3378 (
		_w1983_,
		_w2436_,
		_w2438_,
		_w2447_,
		_w3841_
	);
	LUT4 #(
		.INIT('h001f)
	) name3379 (
		_w1747_,
		_w3838_,
		_w3840_,
		_w3841_,
		_w3842_
	);
	LUT4 #(
		.INIT('h66ef)
	) name3380 (
		_w1723_,
		_w2282_,
		_w2288_,
		_w2449_,
		_w3843_
	);
	LUT4 #(
		.INIT('h888a)
	) name3381 (
		_w1985_,
		_w2450_,
		_w2644_,
		_w3843_,
		_w3844_
	);
	LUT3 #(
		.INIT('h0d)
	) name3382 (
		_w1983_,
		_w2689_,
		_w3844_,
		_w3845_
	);
	LUT3 #(
		.INIT('hd0)
	) name3383 (
		_w2644_,
		_w3842_,
		_w3845_,
		_w3846_
	);
	LUT3 #(
		.INIT('hd0)
	) name3384 (
		_w2292_,
		_w3837_,
		_w3846_,
		_w3847_
	);
	LUT4 #(
		.INIT('h08aa)
	) name3385 (
		_w1731_,
		_w2388_,
		_w3836_,
		_w3847_,
		_w3848_
	);
	LUT4 #(
		.INIT('h4000)
	) name3386 (
		_w1723_,
		_w1727_,
		_w1730_,
		_w1985_,
		_w3849_
	);
	LUT2 #(
		.INIT('h2)
	) name3387 (
		\P1_reg3_reg[21]/NET0131 ,
		\P1_state_reg[0]/NET0131 ,
		_w3850_
	);
	LUT3 #(
		.INIT('h07)
	) name3388 (
		_w1985_,
		_w2695_,
		_w3850_,
		_w3851_
	);
	LUT4 #(
		.INIT('ha8ff)
	) name3389 (
		\P1_state_reg[0]/NET0131 ,
		_w3848_,
		_w3849_,
		_w3851_,
		_w3852_
	);
	LUT2 #(
		.INIT('h8)
	) name3390 (
		_w2159_,
		_w2460_,
		_w3853_
	);
	LUT2 #(
		.INIT('h2)
	) name3391 (
		_w2159_,
		_w2644_,
		_w3854_
	);
	LUT4 #(
		.INIT('h208a)
	) name3392 (
		_w2644_,
		_w2765_,
		_w2773_,
		_w3162_,
		_w3855_
	);
	LUT3 #(
		.INIT('ha8)
	) name3393 (
		_w2292_,
		_w3854_,
		_w3855_,
		_w3856_
	);
	LUT4 #(
		.INIT('h0d05)
	) name3394 (
		_w1987_,
		_w2392_,
		_w2410_,
		_w3465_,
		_w3857_
	);
	LUT4 #(
		.INIT('h7020)
	) name3395 (
		_w1747_,
		_w2175_,
		_w2644_,
		_w3857_,
		_w3858_
	);
	LUT3 #(
		.INIT('ha8)
	) name3396 (
		_w2424_,
		_w3854_,
		_w3858_,
		_w3859_
	);
	LUT4 #(
		.INIT('h00d7)
	) name3397 (
		_w2644_,
		_w2822_,
		_w3162_,
		_w3854_,
		_w3860_
	);
	LUT4 #(
		.INIT('h5655)
	) name3398 (
		_w2155_,
		_w2171_,
		_w2196_,
		_w2436_,
		_w3861_
	);
	LUT4 #(
		.INIT('hf531)
	) name3399 (
		_w2155_,
		_w2159_,
		_w2689_,
		_w2690_,
		_w3862_
	);
	LUT4 #(
		.INIT('h7f00)
	) name3400 (
		_w2447_,
		_w2644_,
		_w3861_,
		_w3862_,
		_w3863_
	);
	LUT3 #(
		.INIT('hd0)
	) name3401 (
		_w2388_,
		_w3860_,
		_w3863_,
		_w3864_
	);
	LUT4 #(
		.INIT('ha8aa)
	) name3402 (
		_w1731_,
		_w3859_,
		_w3856_,
		_w3864_,
		_w3865_
	);
	LUT2 #(
		.INIT('h2)
	) name3403 (
		\P1_reg3_reg[20]/NET0131 ,
		\P1_state_reg[0]/NET0131 ,
		_w3866_
	);
	LUT4 #(
		.INIT('h00ef)
	) name3404 (
		_w1825_,
		_w2158_,
		_w2695_,
		_w3866_,
		_w3867_
	);
	LUT4 #(
		.INIT('ha8ff)
	) name3405 (
		\P1_state_reg[0]/NET0131 ,
		_w3853_,
		_w3865_,
		_w3867_,
		_w3868_
	);
	LUT2 #(
		.INIT('h2)
	) name3406 (
		\P1_reg2_reg[21]/NET0131 ,
		_w2462_,
		_w3869_
	);
	LUT4 #(
		.INIT('hd11d)
	) name3407 (
		\P1_reg2_reg[21]/NET0131 ,
		_w1741_,
		_w3160_,
		_w3835_,
		_w3870_
	);
	LUT4 #(
		.INIT('h1dd1)
	) name3408 (
		\P1_reg2_reg[21]/NET0131 ,
		_w1741_,
		_w2262_,
		_w3160_,
		_w3871_
	);
	LUT3 #(
		.INIT('h10)
	) name3409 (
		_w1748_,
		_w1982_,
		_w2426_,
		_w3872_
	);
	LUT4 #(
		.INIT('ha0a2)
	) name3410 (
		\P1_reg2_reg[21]/NET0131 ,
		_w1741_,
		_w2450_,
		_w3843_,
		_w3873_
	);
	LUT4 #(
		.INIT('h0008)
	) name3411 (
		_w1985_,
		_w2284_,
		_w2288_,
		_w2291_,
		_w3874_
	);
	LUT2 #(
		.INIT('h1)
	) name3412 (
		_w3873_,
		_w3874_,
		_w3875_
	);
	LUT4 #(
		.INIT('h5d00)
	) name3413 (
		_w1741_,
		_w3842_,
		_w3872_,
		_w3875_,
		_w3876_
	);
	LUT3 #(
		.INIT('hd0)
	) name3414 (
		_w2292_,
		_w3871_,
		_w3876_,
		_w3877_
	);
	LUT4 #(
		.INIT('h08aa)
	) name3415 (
		_w1731_,
		_w2388_,
		_w3870_,
		_w3877_,
		_w3878_
	);
	LUT4 #(
		.INIT('h2000)
	) name3416 (
		\P1_reg2_reg[21]/NET0131 ,
		_w1723_,
		_w1727_,
		_w1730_,
		_w3879_
	);
	LUT4 #(
		.INIT('heeec)
	) name3417 (
		\P1_state_reg[0]/NET0131 ,
		_w3869_,
		_w3878_,
		_w3879_,
		_w3880_
	);
	LUT2 #(
		.INIT('h2)
	) name3418 (
		\P1_reg2_reg[18]/NET0131 ,
		_w2462_,
		_w3881_
	);
	LUT4 #(
		.INIT('h2000)
	) name3419 (
		\P1_reg2_reg[18]/NET0131 ,
		_w1723_,
		_w1727_,
		_w1730_,
		_w3882_
	);
	LUT4 #(
		.INIT('hddd1)
	) name3420 (
		\P1_reg2_reg[18]/NET0131 ,
		_w1741_,
		_w3466_,
		_w3467_,
		_w3883_
	);
	LUT2 #(
		.INIT('h2)
	) name3421 (
		_w2424_,
		_w3883_,
		_w3884_
	);
	LUT4 #(
		.INIT('hd11d)
	) name3422 (
		\P1_reg2_reg[18]/NET0131 ,
		_w1741_,
		_w2940_,
		_w3181_,
		_w3885_
	);
	LUT2 #(
		.INIT('h2)
	) name3423 (
		_w2388_,
		_w3885_,
		_w3886_
	);
	LUT4 #(
		.INIT('h1dd1)
	) name3424 (
		\P1_reg2_reg[18]/NET0131 ,
		_w1741_,
		_w2958_,
		_w3181_,
		_w3887_
	);
	LUT4 #(
		.INIT('h0008)
	) name3425 (
		_w2197_,
		_w2284_,
		_w2288_,
		_w2291_,
		_w3888_
	);
	LUT4 #(
		.INIT('ha2a0)
	) name3426 (
		\P1_reg2_reg[18]/NET0131 ,
		_w1741_,
		_w2450_,
		_w2452_,
		_w3889_
	);
	LUT2 #(
		.INIT('h1)
	) name3427 (
		_w3888_,
		_w3889_,
		_w3890_
	);
	LUT3 #(
		.INIT('h70)
	) name3428 (
		_w1741_,
		_w3473_,
		_w3890_,
		_w3891_
	);
	LUT3 #(
		.INIT('hd0)
	) name3429 (
		_w2292_,
		_w3887_,
		_w3891_,
		_w3892_
	);
	LUT4 #(
		.INIT('ha8aa)
	) name3430 (
		_w1731_,
		_w3884_,
		_w3886_,
		_w3892_,
		_w3893_
	);
	LUT4 #(
		.INIT('heeec)
	) name3431 (
		\P1_state_reg[0]/NET0131 ,
		_w3881_,
		_w3882_,
		_w3893_,
		_w3894_
	);
	LUT2 #(
		.INIT('h2)
	) name3432 (
		\P1_reg2_reg[17]/NET0131 ,
		_w2462_,
		_w3895_
	);
	LUT4 #(
		.INIT('h2000)
	) name3433 (
		\P1_reg2_reg[17]/NET0131 ,
		_w1723_,
		_w1727_,
		_w1730_,
		_w3896_
	);
	LUT2 #(
		.INIT('h2)
	) name3434 (
		\P1_reg2_reg[17]/NET0131 ,
		_w1741_,
		_w3897_
	);
	LUT4 #(
		.INIT('ha028)
	) name3435 (
		_w1741_,
		_w2336_,
		_w3170_,
		_w3486_,
		_w3898_
	);
	LUT3 #(
		.INIT('ha8)
	) name3436 (
		_w2388_,
		_w3897_,
		_w3898_,
		_w3899_
	);
	LUT4 #(
		.INIT('h1dd1)
	) name3437 (
		\P1_reg2_reg[17]/NET0131 ,
		_w1741_,
		_w3170_,
		_w3489_,
		_w3900_
	);
	LUT4 #(
		.INIT('he020)
	) name3438 (
		\P1_reg2_reg[17]/NET0131 ,
		_w1741_,
		_w2424_,
		_w3492_,
		_w3901_
	);
	LUT4 #(
		.INIT('hddd1)
	) name3439 (
		\P1_reg2_reg[17]/NET0131 ,
		_w1741_,
		_w2436_,
		_w3495_,
		_w3902_
	);
	LUT2 #(
		.INIT('h8)
	) name3440 (
		_w2183_,
		_w2426_,
		_w3903_
	);
	LUT3 #(
		.INIT('h80)
	) name3441 (
		_w1741_,
		_w2183_,
		_w2426_,
		_w3904_
	);
	LUT4 #(
		.INIT('haa20)
	) name3442 (
		\P1_reg2_reg[17]/NET0131 ,
		_w1741_,
		_w2426_,
		_w2450_,
		_w3905_
	);
	LUT4 #(
		.INIT('h0008)
	) name3443 (
		_w2185_,
		_w2284_,
		_w2288_,
		_w2291_,
		_w3906_
	);
	LUT3 #(
		.INIT('h01)
	) name3444 (
		_w3905_,
		_w3906_,
		_w3904_,
		_w3907_
	);
	LUT3 #(
		.INIT('hd0)
	) name3445 (
		_w2447_,
		_w3902_,
		_w3907_,
		_w3908_
	);
	LUT4 #(
		.INIT('h0d00)
	) name3446 (
		_w2292_,
		_w3900_,
		_w3901_,
		_w3908_,
		_w3909_
	);
	LUT4 #(
		.INIT('h1311)
	) name3447 (
		_w1731_,
		_w3896_,
		_w3899_,
		_w3909_,
		_w3910_
	);
	LUT3 #(
		.INIT('hce)
	) name3448 (
		\P1_state_reg[0]/NET0131 ,
		_w3895_,
		_w3910_,
		_w3911_
	);
	LUT2 #(
		.INIT('h2)
	) name3449 (
		\P1_reg2_reg[19]/NET0131 ,
		_w2462_,
		_w3912_
	);
	LUT4 #(
		.INIT('h2000)
	) name3450 (
		\P1_reg2_reg[19]/NET0131 ,
		_w1723_,
		_w1727_,
		_w1730_,
		_w3913_
	);
	LUT4 #(
		.INIT('he020)
	) name3451 (
		\P1_reg2_reg[19]/NET0131 ,
		_w1741_,
		_w2424_,
		_w3510_,
		_w3914_
	);
	LUT4 #(
		.INIT('hd11d)
	) name3452 (
		\P1_reg2_reg[19]/NET0131 ,
		_w1741_,
		_w2662_,
		_w3165_,
		_w3915_
	);
	LUT2 #(
		.INIT('h2)
	) name3453 (
		_w2292_,
		_w3915_,
		_w3916_
	);
	LUT4 #(
		.INIT('h1dd1)
	) name3454 (
		\P1_reg2_reg[19]/NET0131 ,
		_w1741_,
		_w2675_,
		_w3165_,
		_w3917_
	);
	LUT4 #(
		.INIT('h0008)
	) name3455 (
		_w2172_,
		_w2284_,
		_w2288_,
		_w2291_,
		_w3918_
	);
	LUT4 #(
		.INIT('ha2a0)
	) name3456 (
		\P1_reg2_reg[19]/NET0131 ,
		_w1741_,
		_w2450_,
		_w2452_,
		_w3919_
	);
	LUT2 #(
		.INIT('h1)
	) name3457 (
		_w3918_,
		_w3919_,
		_w3920_
	);
	LUT4 #(
		.INIT('h5700)
	) name3458 (
		_w1741_,
		_w3515_,
		_w3516_,
		_w3920_,
		_w3921_
	);
	LUT3 #(
		.INIT('hd0)
	) name3459 (
		_w2388_,
		_w3917_,
		_w3921_,
		_w3922_
	);
	LUT4 #(
		.INIT('ha8aa)
	) name3460 (
		_w1731_,
		_w3914_,
		_w3916_,
		_w3922_,
		_w3923_
	);
	LUT4 #(
		.INIT('heeec)
	) name3461 (
		\P1_state_reg[0]/NET0131 ,
		_w3912_,
		_w3913_,
		_w3923_,
		_w3924_
	);
	LUT4 #(
		.INIT('h1000)
	) name3462 (
		_w947_,
		_w1189_,
		_w1352_,
		_w1356_,
		_w3925_
	);
	LUT4 #(
		.INIT('h04c4)
	) name3463 (
		_w947_,
		_w1191_,
		_w1411_,
		_w3289_,
		_w3926_
	);
	LUT3 #(
		.INIT('h54)
	) name3464 (
		_w947_,
		_w1441_,
		_w1443_,
		_w3927_
	);
	LUT3 #(
		.INIT('h07)
	) name3465 (
		_w945_,
		_w1440_,
		_w3927_,
		_w3928_
	);
	LUT2 #(
		.INIT('h4)
	) name3466 (
		_w3926_,
		_w3928_,
		_w3929_
	);
	LUT4 #(
		.INIT('h010d)
	) name3467 (
		_w947_,
		_w1369_,
		_w1409_,
		_w3291_,
		_w3930_
	);
	LUT4 #(
		.INIT('h04c4)
	) name3468 (
		_w947_,
		_w1447_,
		_w1411_,
		_w3281_,
		_w3931_
	);
	LUT4 #(
		.INIT('h010d)
	) name3469 (
		_w947_,
		_w1369_,
		_w1496_,
		_w3281_,
		_w3932_
	);
	LUT3 #(
		.INIT('h01)
	) name3470 (
		_w3931_,
		_w3932_,
		_w3930_,
		_w3933_
	);
	LUT4 #(
		.INIT('h3111)
	) name3471 (
		_w1359_,
		_w3925_,
		_w3929_,
		_w3933_,
		_w3934_
	);
	LUT2 #(
		.INIT('h4)
	) name3472 (
		\P1_state_reg[0]/NET0131 ,
		\P2_reg3_reg[21]/NET0131 ,
		_w3935_
	);
	LUT3 #(
		.INIT('h0b)
	) name3473 (
		_w947_,
		_w1349_,
		_w3935_,
		_w3936_
	);
	LUT3 #(
		.INIT('h2f)
	) name3474 (
		\P1_state_reg[0]/NET0131 ,
		_w3934_,
		_w3936_,
		_w3937_
	);
	LUT4 #(
		.INIT('h4000)
	) name3475 (
		_w1723_,
		_w1727_,
		_w1730_,
		_w1973_,
		_w3938_
	);
	LUT2 #(
		.INIT('h2)
	) name3476 (
		_w1973_,
		_w2644_,
		_w3939_
	);
	LUT4 #(
		.INIT('h00fd)
	) name3477 (
		_w2644_,
		_w3689_,
		_w3690_,
		_w3939_,
		_w3940_
	);
	LUT4 #(
		.INIT('hf531)
	) name3478 (
		_w1971_,
		_w1973_,
		_w2689_,
		_w2690_,
		_w3941_
	);
	LUT4 #(
		.INIT('h7f00)
	) name3479 (
		_w2447_,
		_w2644_,
		_w3693_,
		_w3941_,
		_w3942_
	);
	LUT3 #(
		.INIT('hd0)
	) name3480 (
		_w2424_,
		_w3940_,
		_w3942_,
		_w3943_
	);
	LUT4 #(
		.INIT('h2822)
	) name3481 (
		_w2644_,
		_w3166_,
		_w3699_,
		_w3701_,
		_w3944_
	);
	LUT3 #(
		.INIT('ha8)
	) name3482 (
		_w2292_,
		_w3939_,
		_w3944_,
		_w3945_
	);
	LUT4 #(
		.INIT('h8288)
	) name3483 (
		_w2644_,
		_w3166_,
		_w3705_,
		_w3707_,
		_w3946_
	);
	LUT3 #(
		.INIT('ha8)
	) name3484 (
		_w2388_,
		_w3939_,
		_w3946_,
		_w3947_
	);
	LUT4 #(
		.INIT('ha8aa)
	) name3485 (
		_w1731_,
		_w3945_,
		_w3947_,
		_w3943_,
		_w3948_
	);
	LUT2 #(
		.INIT('h2)
	) name3486 (
		\P1_reg3_reg[22]/NET0131 ,
		\P1_state_reg[0]/NET0131 ,
		_w3949_
	);
	LUT3 #(
		.INIT('h07)
	) name3487 (
		_w1973_,
		_w2695_,
		_w3949_,
		_w3950_
	);
	LUT4 #(
		.INIT('ha8ff)
	) name3488 (
		\P1_state_reg[0]/NET0131 ,
		_w3938_,
		_w3948_,
		_w3950_,
		_w3951_
	);
	LUT4 #(
		.INIT('hd070)
	) name3489 (
		\P1_state_reg[0]/NET0131 ,
		\P2_IR_reg[23]/NET0131 ,
		\P2_reg0_reg[18]/NET0131 ,
		_w1188_,
		_w3952_
	);
	LUT4 #(
		.INIT('h2000)
	) name3490 (
		\P2_reg0_reg[18]/NET0131 ,
		_w1189_,
		_w1352_,
		_w1356_,
		_w3953_
	);
	LUT4 #(
		.INIT('h0e02)
	) name3491 (
		\P2_reg0_reg[18]/NET0131 ,
		_w1411_,
		_w1496_,
		_w2543_,
		_w3954_
	);
	LUT3 #(
		.INIT('ha2)
	) name3492 (
		\P2_reg0_reg[18]/NET0131 ,
		_w1684_,
		_w1685_,
		_w3955_
	);
	LUT3 #(
		.INIT('h40)
	) name3493 (
		_w925_,
		_w1411_,
		_w1442_,
		_w3956_
	);
	LUT2 #(
		.INIT('h1)
	) name3494 (
		_w3955_,
		_w3956_,
		_w3957_
	);
	LUT2 #(
		.INIT('h4)
	) name3495 (
		_w3954_,
		_w3957_,
		_w3958_
	);
	LUT4 #(
		.INIT('h0232)
	) name3496 (
		\P2_reg0_reg[18]/NET0131 ,
		_w1409_,
		_w1411_,
		_w2558_,
		_w3959_
	);
	LUT4 #(
		.INIT('he020)
	) name3497 (
		\P2_reg0_reg[18]/NET0131 ,
		_w1369_,
		_w1447_,
		_w2543_,
		_w3960_
	);
	LUT4 #(
		.INIT('h08c8)
	) name3498 (
		\P2_reg0_reg[18]/NET0131 ,
		_w1191_,
		_w1369_,
		_w2564_,
		_w3961_
	);
	LUT3 #(
		.INIT('h01)
	) name3499 (
		_w3960_,
		_w3961_,
		_w3959_,
		_w3962_
	);
	LUT4 #(
		.INIT('h3111)
	) name3500 (
		_w1359_,
		_w3953_,
		_w3958_,
		_w3962_,
		_w3963_
	);
	LUT3 #(
		.INIT('hce)
	) name3501 (
		\P1_state_reg[0]/NET0131 ,
		_w3952_,
		_w3963_,
		_w3964_
	);
	LUT2 #(
		.INIT('h2)
	) name3502 (
		\P1_reg1_reg[31]/NET0131 ,
		_w2462_,
		_w3965_
	);
	LUT4 #(
		.INIT('h2000)
	) name3503 (
		\P1_reg1_reg[31]/NET0131 ,
		_w1723_,
		_w1727_,
		_w1730_,
		_w3966_
	);
	LUT4 #(
		.INIT('h1dd1)
	) name3504 (
		\P1_reg1_reg[31]/NET0131 ,
		_w2520_,
		_w3126_,
		_w3566_,
		_w3967_
	);
	LUT2 #(
		.INIT('h8)
	) name3505 (
		_w2424_,
		_w2520_,
		_w3968_
	);
	LUT4 #(
		.INIT('h7000)
	) name3506 (
		_w2922_,
		_w3569_,
		_w3570_,
		_w3968_,
		_w3969_
	);
	LUT4 #(
		.INIT('hc5f5)
	) name3507 (
		\P1_reg1_reg[31]/NET0131 ,
		_w1748_,
		_w2520_,
		_w3125_,
		_w3970_
	);
	LUT4 #(
		.INIT('h0a2a)
	) name3508 (
		\P1_reg1_reg[31]/NET0131 ,
		_w2520_,
		_w2524_,
		_w3574_,
		_w3971_
	);
	LUT3 #(
		.INIT('h0d)
	) name3509 (
		_w2426_,
		_w3970_,
		_w3971_,
		_w3972_
	);
	LUT4 #(
		.INIT('h0d00)
	) name3510 (
		_w2447_,
		_w3967_,
		_w3969_,
		_w3972_,
		_w3973_
	);
	LUT4 #(
		.INIT('ha0a8)
	) name3511 (
		\P1_state_reg[0]/NET0131 ,
		_w1731_,
		_w3966_,
		_w3973_,
		_w3974_
	);
	LUT2 #(
		.INIT('he)
	) name3512 (
		_w3965_,
		_w3974_,
		_w3975_
	);
	LUT4 #(
		.INIT('hd070)
	) name3513 (
		\P1_state_reg[0]/NET0131 ,
		\P2_IR_reg[23]/NET0131 ,
		\P2_reg0_reg[19]/NET0131 ,
		_w1188_,
		_w3976_
	);
	LUT4 #(
		.INIT('h2000)
	) name3514 (
		\P2_reg0_reg[19]/NET0131 ,
		_w1189_,
		_w1352_,
		_w1356_,
		_w3977_
	);
	LUT4 #(
		.INIT('haaa8)
	) name3515 (
		\P2_reg0_reg[19]/NET0131 ,
		_w1361_,
		_w1363_,
		_w1368_,
		_w3978_
	);
	LUT4 #(
		.INIT('h020e)
	) name3516 (
		\P2_reg0_reg[19]/NET0131 ,
		_w1411_,
		_w1496_,
		_w2573_,
		_w3979_
	);
	LUT3 #(
		.INIT('ha2)
	) name3517 (
		\P2_reg0_reg[19]/NET0131 ,
		_w1684_,
		_w1685_,
		_w3980_
	);
	LUT3 #(
		.INIT('h07)
	) name3518 (
		_w1411_,
		_w3066_,
		_w3980_,
		_w3981_
	);
	LUT2 #(
		.INIT('h4)
	) name3519 (
		_w3979_,
		_w3981_,
		_w3982_
	);
	LUT4 #(
		.INIT('h6500)
	) name3520 (
		_w1272_,
		_w1387_,
		_w1394_,
		_w1411_,
		_w3983_
	);
	LUT3 #(
		.INIT('h54)
	) name3521 (
		_w1409_,
		_w3978_,
		_w3983_,
		_w3984_
	);
	LUT4 #(
		.INIT('h111d)
	) name3522 (
		\P2_reg0_reg[19]/NET0131 ,
		_w1369_,
		_w2581_,
		_w2583_,
		_w3985_
	);
	LUT4 #(
		.INIT('h20e0)
	) name3523 (
		\P2_reg0_reg[19]/NET0131 ,
		_w1369_,
		_w1447_,
		_w2573_,
		_w3986_
	);
	LUT4 #(
		.INIT('h000d)
	) name3524 (
		_w1191_,
		_w3985_,
		_w3986_,
		_w3984_,
		_w3987_
	);
	LUT4 #(
		.INIT('h3111)
	) name3525 (
		_w1359_,
		_w3977_,
		_w3982_,
		_w3987_,
		_w3988_
	);
	LUT3 #(
		.INIT('hce)
	) name3526 (
		\P1_state_reg[0]/NET0131 ,
		_w3976_,
		_w3988_,
		_w3989_
	);
	LUT4 #(
		.INIT('hd070)
	) name3527 (
		\P1_state_reg[0]/NET0131 ,
		\P2_IR_reg[23]/NET0131 ,
		\P2_reg0_reg[17]/NET0131 ,
		_w1188_,
		_w3990_
	);
	LUT4 #(
		.INIT('h2000)
	) name3528 (
		\P2_reg0_reg[17]/NET0131 ,
		_w1189_,
		_w1352_,
		_w1356_,
		_w3991_
	);
	LUT4 #(
		.INIT('haaa8)
	) name3529 (
		\P2_reg0_reg[17]/NET0131 ,
		_w1361_,
		_w1363_,
		_w1368_,
		_w3992_
	);
	LUT4 #(
		.INIT('h0e02)
	) name3530 (
		\P2_reg0_reg[17]/NET0131 ,
		_w1411_,
		_w1496_,
		_w2593_,
		_w3993_
	);
	LUT4 #(
		.INIT('h111d)
	) name3531 (
		\P2_reg0_reg[17]/NET0131 ,
		_w1369_,
		_w2596_,
		_w2597_,
		_w3994_
	);
	LUT3 #(
		.INIT('h40)
	) name3532 (
		_w860_,
		_w1411_,
		_w1442_,
		_w3995_
	);
	LUT3 #(
		.INIT('ha2)
	) name3533 (
		\P2_reg0_reg[17]/NET0131 ,
		_w1684_,
		_w1685_,
		_w3996_
	);
	LUT2 #(
		.INIT('h1)
	) name3534 (
		_w3995_,
		_w3996_,
		_w3997_
	);
	LUT3 #(
		.INIT('hd0)
	) name3535 (
		_w1191_,
		_w3994_,
		_w3997_,
		_w3998_
	);
	LUT4 #(
		.INIT('he020)
	) name3536 (
		\P2_reg0_reg[17]/NET0131 ,
		_w1369_,
		_w1447_,
		_w2593_,
		_w3999_
	);
	LUT4 #(
		.INIT('h4484)
	) name3537 (
		_w1314_,
		_w1411_,
		_w1665_,
		_w2604_,
		_w4000_
	);
	LUT3 #(
		.INIT('h54)
	) name3538 (
		_w1409_,
		_w3992_,
		_w4000_,
		_w4001_
	);
	LUT4 #(
		.INIT('h0100)
	) name3539 (
		_w3993_,
		_w3999_,
		_w4001_,
		_w3998_,
		_w4002_
	);
	LUT4 #(
		.INIT('ha0a8)
	) name3540 (
		\P1_state_reg[0]/NET0131 ,
		_w1359_,
		_w3991_,
		_w4002_,
		_w4003_
	);
	LUT2 #(
		.INIT('he)
	) name3541 (
		_w3990_,
		_w4003_,
		_w4004_
	);
	LUT4 #(
		.INIT('hd070)
	) name3542 (
		\P1_state_reg[0]/NET0131 ,
		\P2_IR_reg[23]/NET0131 ,
		\P2_reg0_reg[21]/NET0131 ,
		_w1188_,
		_w4005_
	);
	LUT4 #(
		.INIT('h2000)
	) name3543 (
		\P2_reg0_reg[21]/NET0131 ,
		_w1189_,
		_w1352_,
		_w1356_,
		_w4006_
	);
	LUT4 #(
		.INIT('h08c8)
	) name3544 (
		\P2_reg0_reg[21]/NET0131 ,
		_w1191_,
		_w1369_,
		_w3289_,
		_w4007_
	);
	LUT3 #(
		.INIT('ha2)
	) name3545 (
		\P2_reg0_reg[21]/NET0131 ,
		_w1684_,
		_w1685_,
		_w4008_
	);
	LUT3 #(
		.INIT('h07)
	) name3546 (
		_w1411_,
		_w3283_,
		_w4008_,
		_w4009_
	);
	LUT2 #(
		.INIT('h4)
	) name3547 (
		_w4007_,
		_w4009_,
		_w4010_
	);
	LUT4 #(
		.INIT('h0232)
	) name3548 (
		\P2_reg0_reg[21]/NET0131 ,
		_w1409_,
		_w1411_,
		_w3291_,
		_w4011_
	);
	LUT4 #(
		.INIT('h20e0)
	) name3549 (
		\P2_reg0_reg[21]/NET0131 ,
		_w1369_,
		_w1447_,
		_w3281_,
		_w4012_
	);
	LUT4 #(
		.INIT('h020e)
	) name3550 (
		\P2_reg0_reg[21]/NET0131 ,
		_w1411_,
		_w1496_,
		_w3281_,
		_w4013_
	);
	LUT3 #(
		.INIT('h01)
	) name3551 (
		_w4012_,
		_w4013_,
		_w4011_,
		_w4014_
	);
	LUT4 #(
		.INIT('h3111)
	) name3552 (
		_w1359_,
		_w4006_,
		_w4010_,
		_w4014_,
		_w4015_
	);
	LUT3 #(
		.INIT('hce)
	) name3553 (
		\P1_state_reg[0]/NET0131 ,
		_w4005_,
		_w4015_,
		_w4016_
	);
	LUT4 #(
		.INIT('hd070)
	) name3554 (
		\P1_state_reg[0]/NET0131 ,
		\P2_IR_reg[23]/NET0131 ,
		\P2_reg0_reg[20]/NET0131 ,
		_w1188_,
		_w4017_
	);
	LUT4 #(
		.INIT('h2000)
	) name3555 (
		\P2_reg0_reg[20]/NET0131 ,
		_w1189_,
		_w1352_,
		_w1356_,
		_w4018_
	);
	LUT4 #(
		.INIT('h020e)
	) name3556 (
		\P2_reg0_reg[20]/NET0131 ,
		_w1411_,
		_w1496_,
		_w2911_,
		_w4019_
	);
	LUT3 #(
		.INIT('ha2)
	) name3557 (
		\P2_reg0_reg[20]/NET0131 ,
		_w1684_,
		_w1685_,
		_w4020_
	);
	LUT3 #(
		.INIT('h10)
	) name3558 (
		_w546_,
		_w962_,
		_w1687_,
		_w4021_
	);
	LUT2 #(
		.INIT('h1)
	) name3559 (
		_w4020_,
		_w4021_,
		_w4022_
	);
	LUT2 #(
		.INIT('h4)
	) name3560 (
		_w4019_,
		_w4022_,
		_w4023_
	);
	LUT4 #(
		.INIT('h08c8)
	) name3561 (
		\P2_reg0_reg[20]/NET0131 ,
		_w1191_,
		_w1369_,
		_w2902_,
		_w4024_
	);
	LUT4 #(
		.INIT('h20e0)
	) name3562 (
		\P2_reg0_reg[20]/NET0131 ,
		_w1369_,
		_w1447_,
		_w2911_,
		_w4025_
	);
	LUT4 #(
		.INIT('h0232)
	) name3563 (
		\P2_reg0_reg[20]/NET0131 ,
		_w1409_,
		_w1411_,
		_w2909_,
		_w4026_
	);
	LUT3 #(
		.INIT('h01)
	) name3564 (
		_w4025_,
		_w4026_,
		_w4024_,
		_w4027_
	);
	LUT4 #(
		.INIT('h3111)
	) name3565 (
		_w1359_,
		_w4018_,
		_w4023_,
		_w4027_,
		_w4028_
	);
	LUT3 #(
		.INIT('hce)
	) name3566 (
		\P1_state_reg[0]/NET0131 ,
		_w4017_,
		_w4028_,
		_w4029_
	);
	LUT2 #(
		.INIT('h2)
	) name3567 (
		\P1_reg2_reg[20]/NET0131 ,
		_w2462_,
		_w4030_
	);
	LUT4 #(
		.INIT('h2000)
	) name3568 (
		\P1_reg2_reg[20]/NET0131 ,
		_w1723_,
		_w1727_,
		_w1730_,
		_w4031_
	);
	LUT2 #(
		.INIT('h2)
	) name3569 (
		\P1_reg2_reg[20]/NET0131 ,
		_w1741_,
		_w4032_
	);
	LUT4 #(
		.INIT('h208a)
	) name3570 (
		_w1741_,
		_w2765_,
		_w2773_,
		_w3162_,
		_w4033_
	);
	LUT3 #(
		.INIT('ha8)
	) name3571 (
		_w2292_,
		_w4032_,
		_w4033_,
		_w4034_
	);
	LUT4 #(
		.INIT('h2a08)
	) name3572 (
		_w1741_,
		_w1747_,
		_w2175_,
		_w3857_,
		_w4035_
	);
	LUT3 #(
		.INIT('ha8)
	) name3573 (
		_w2424_,
		_w4032_,
		_w4035_,
		_w4036_
	);
	LUT4 #(
		.INIT('hd11d)
	) name3574 (
		\P1_reg2_reg[20]/NET0131 ,
		_w1741_,
		_w2822_,
		_w3162_,
		_w4037_
	);
	LUT3 #(
		.INIT('h10)
	) name3575 (
		_w1748_,
		_w2154_,
		_w2426_,
		_w4038_
	);
	LUT4 #(
		.INIT('haa80)
	) name3576 (
		_w1741_,
		_w2447_,
		_w3861_,
		_w4038_,
		_w4039_
	);
	LUT4 #(
		.INIT('h00ab)
	) name3577 (
		_w1741_,
		_w2426_,
		_w2447_,
		_w2450_,
		_w4040_
	);
	LUT2 #(
		.INIT('h8)
	) name3578 (
		_w2159_,
		_w2454_,
		_w4041_
	);
	LUT3 #(
		.INIT('h0d)
	) name3579 (
		\P1_reg2_reg[20]/NET0131 ,
		_w4040_,
		_w4041_,
		_w4042_
	);
	LUT2 #(
		.INIT('h4)
	) name3580 (
		_w4039_,
		_w4042_,
		_w4043_
	);
	LUT3 #(
		.INIT('hd0)
	) name3581 (
		_w2388_,
		_w4037_,
		_w4043_,
		_w4044_
	);
	LUT4 #(
		.INIT('ha8aa)
	) name3582 (
		_w1731_,
		_w4036_,
		_w4034_,
		_w4044_,
		_w4045_
	);
	LUT4 #(
		.INIT('heeec)
	) name3583 (
		\P1_state_reg[0]/NET0131 ,
		_w4030_,
		_w4031_,
		_w4045_,
		_w4046_
	);
	LUT4 #(
		.INIT('hd070)
	) name3584 (
		\P1_state_reg[0]/NET0131 ,
		\P2_IR_reg[23]/NET0131 ,
		\P2_reg1_reg[17]/NET0131 ,
		_w1188_,
		_w4047_
	);
	LUT4 #(
		.INIT('h2000)
	) name3585 (
		\P2_reg1_reg[17]/NET0131 ,
		_w1189_,
		_w1352_,
		_w1356_,
		_w4048_
	);
	LUT4 #(
		.INIT('haa02)
	) name3586 (
		\P2_reg1_reg[17]/NET0131 ,
		_w1361_,
		_w1363_,
		_w1368_,
		_w4049_
	);
	LUT4 #(
		.INIT('h0e02)
	) name3587 (
		\P2_reg1_reg[17]/NET0131 ,
		_w1516_,
		_w1575_,
		_w2593_,
		_w4050_
	);
	LUT4 #(
		.INIT('ha8aa)
	) name3588 (
		\P2_reg1_reg[17]/NET0131 ,
		_w1361_,
		_w1363_,
		_w1368_,
		_w4051_
	);
	LUT4 #(
		.INIT('h111d)
	) name3589 (
		\P2_reg1_reg[17]/NET0131 ,
		_w1507_,
		_w2596_,
		_w2597_,
		_w4052_
	);
	LUT3 #(
		.INIT('h40)
	) name3590 (
		_w860_,
		_w1442_,
		_w1516_,
		_w4053_
	);
	LUT3 #(
		.INIT('ha2)
	) name3591 (
		\P2_reg1_reg[17]/NET0131 ,
		_w1684_,
		_w2469_,
		_w4054_
	);
	LUT2 #(
		.INIT('h1)
	) name3592 (
		_w4053_,
		_w4054_,
		_w4055_
	);
	LUT3 #(
		.INIT('hd0)
	) name3593 (
		_w1191_,
		_w4052_,
		_w4055_,
		_w4056_
	);
	LUT3 #(
		.INIT('ha8)
	) name3594 (
		_w1530_,
		_w3043_,
		_w4051_,
		_w4057_
	);
	LUT3 #(
		.INIT('h54)
	) name3595 (
		_w1506_,
		_w3041_,
		_w4049_,
		_w4058_
	);
	LUT4 #(
		.INIT('h0100)
	) name3596 (
		_w4050_,
		_w4057_,
		_w4058_,
		_w4056_,
		_w4059_
	);
	LUT4 #(
		.INIT('ha0a8)
	) name3597 (
		\P1_state_reg[0]/NET0131 ,
		_w1359_,
		_w4048_,
		_w4059_,
		_w4060_
	);
	LUT2 #(
		.INIT('he)
	) name3598 (
		_w4047_,
		_w4060_,
		_w4061_
	);
	LUT4 #(
		.INIT('hd070)
	) name3599 (
		\P1_state_reg[0]/NET0131 ,
		\P2_IR_reg[23]/NET0131 ,
		\P2_reg1_reg[18]/NET0131 ,
		_w1188_,
		_w4062_
	);
	LUT4 #(
		.INIT('h2000)
	) name3600 (
		\P2_reg1_reg[18]/NET0131 ,
		_w1189_,
		_w1352_,
		_w1356_,
		_w4063_
	);
	LUT4 #(
		.INIT('h0e02)
	) name3601 (
		\P2_reg1_reg[18]/NET0131 ,
		_w1516_,
		_w1575_,
		_w2543_,
		_w4064_
	);
	LUT3 #(
		.INIT('ha2)
	) name3602 (
		\P2_reg1_reg[18]/NET0131 ,
		_w1684_,
		_w2469_,
		_w4065_
	);
	LUT3 #(
		.INIT('h40)
	) name3603 (
		_w925_,
		_w1442_,
		_w1516_,
		_w4066_
	);
	LUT2 #(
		.INIT('h1)
	) name3604 (
		_w4065_,
		_w4066_,
		_w4067_
	);
	LUT2 #(
		.INIT('h4)
	) name3605 (
		_w4064_,
		_w4067_,
		_w4068_
	);
	LUT4 #(
		.INIT('h0232)
	) name3606 (
		\P2_reg1_reg[18]/NET0131 ,
		_w1506_,
		_w1516_,
		_w2558_,
		_w4069_
	);
	LUT4 #(
		.INIT('h20e0)
	) name3607 (
		\P2_reg1_reg[18]/NET0131 ,
		_w1507_,
		_w1530_,
		_w2558_,
		_w4070_
	);
	LUT4 #(
		.INIT('h08c8)
	) name3608 (
		\P2_reg1_reg[18]/NET0131 ,
		_w1191_,
		_w1507_,
		_w2564_,
		_w4071_
	);
	LUT3 #(
		.INIT('h01)
	) name3609 (
		_w4070_,
		_w4071_,
		_w4069_,
		_w4072_
	);
	LUT4 #(
		.INIT('h3111)
	) name3610 (
		_w1359_,
		_w4063_,
		_w4068_,
		_w4072_,
		_w4073_
	);
	LUT3 #(
		.INIT('hce)
	) name3611 (
		\P1_state_reg[0]/NET0131 ,
		_w4062_,
		_w4073_,
		_w4074_
	);
	LUT4 #(
		.INIT('hd070)
	) name3612 (
		\P1_state_reg[0]/NET0131 ,
		\P2_IR_reg[23]/NET0131 ,
		\P2_reg1_reg[19]/NET0131 ,
		_w1188_,
		_w4075_
	);
	LUT4 #(
		.INIT('h2000)
	) name3613 (
		\P2_reg1_reg[19]/NET0131 ,
		_w1189_,
		_w1352_,
		_w1356_,
		_w4076_
	);
	LUT4 #(
		.INIT('ha8aa)
	) name3614 (
		\P2_reg1_reg[19]/NET0131 ,
		_w1361_,
		_w1363_,
		_w1368_,
		_w4077_
	);
	LUT4 #(
		.INIT('h111d)
	) name3615 (
		\P2_reg1_reg[19]/NET0131 ,
		_w1507_,
		_w2581_,
		_w2583_,
		_w4078_
	);
	LUT3 #(
		.INIT('ha2)
	) name3616 (
		\P2_reg1_reg[19]/NET0131 ,
		_w1684_,
		_w2469_,
		_w4079_
	);
	LUT3 #(
		.INIT('h07)
	) name3617 (
		_w1516_,
		_w3066_,
		_w4079_,
		_w4080_
	);
	LUT3 #(
		.INIT('hd0)
	) name3618 (
		_w1191_,
		_w4078_,
		_w4080_,
		_w4081_
	);
	LUT4 #(
		.INIT('haa02)
	) name3619 (
		\P2_reg1_reg[19]/NET0131 ,
		_w1361_,
		_w1363_,
		_w1368_,
		_w4082_
	);
	LUT4 #(
		.INIT('h020e)
	) name3620 (
		\P2_reg1_reg[19]/NET0131 ,
		_w1516_,
		_w1575_,
		_w2573_,
		_w4083_
	);
	LUT3 #(
		.INIT('ha8)
	) name3621 (
		_w1530_,
		_w3075_,
		_w4077_,
		_w4084_
	);
	LUT3 #(
		.INIT('h54)
	) name3622 (
		_w1506_,
		_w3073_,
		_w4082_,
		_w4085_
	);
	LUT3 #(
		.INIT('h01)
	) name3623 (
		_w4084_,
		_w4085_,
		_w4083_,
		_w4086_
	);
	LUT4 #(
		.INIT('h3111)
	) name3624 (
		_w1359_,
		_w4076_,
		_w4081_,
		_w4086_,
		_w4087_
	);
	LUT3 #(
		.INIT('hce)
	) name3625 (
		\P1_state_reg[0]/NET0131 ,
		_w4075_,
		_w4087_,
		_w4088_
	);
	LUT4 #(
		.INIT('hd070)
	) name3626 (
		\P1_state_reg[0]/NET0131 ,
		\P2_IR_reg[23]/NET0131 ,
		\P2_reg1_reg[20]/NET0131 ,
		_w1188_,
		_w4089_
	);
	LUT4 #(
		.INIT('h2000)
	) name3627 (
		\P2_reg1_reg[20]/NET0131 ,
		_w1189_,
		_w1352_,
		_w1356_,
		_w4090_
	);
	LUT4 #(
		.INIT('h020e)
	) name3628 (
		\P2_reg1_reg[20]/NET0131 ,
		_w1516_,
		_w1575_,
		_w2911_,
		_w4091_
	);
	LUT3 #(
		.INIT('ha2)
	) name3629 (
		\P2_reg1_reg[20]/NET0131 ,
		_w1684_,
		_w2469_,
		_w4092_
	);
	LUT3 #(
		.INIT('h10)
	) name3630 (
		_w546_,
		_w962_,
		_w2471_,
		_w4093_
	);
	LUT2 #(
		.INIT('h1)
	) name3631 (
		_w4092_,
		_w4093_,
		_w4094_
	);
	LUT2 #(
		.INIT('h4)
	) name3632 (
		_w4091_,
		_w4094_,
		_w4095_
	);
	LUT4 #(
		.INIT('h08c8)
	) name3633 (
		\P2_reg1_reg[20]/NET0131 ,
		_w1191_,
		_w1507_,
		_w2902_,
		_w4096_
	);
	LUT4 #(
		.INIT('h0232)
	) name3634 (
		\P2_reg1_reg[20]/NET0131 ,
		_w1506_,
		_w1516_,
		_w2909_,
		_w4097_
	);
	LUT4 #(
		.INIT('h20e0)
	) name3635 (
		\P2_reg1_reg[20]/NET0131 ,
		_w1507_,
		_w1530_,
		_w2909_,
		_w4098_
	);
	LUT3 #(
		.INIT('h01)
	) name3636 (
		_w4097_,
		_w4098_,
		_w4096_,
		_w4099_
	);
	LUT4 #(
		.INIT('h3111)
	) name3637 (
		_w1359_,
		_w4090_,
		_w4095_,
		_w4099_,
		_w4100_
	);
	LUT3 #(
		.INIT('hce)
	) name3638 (
		\P1_state_reg[0]/NET0131 ,
		_w4089_,
		_w4100_,
		_w4101_
	);
	LUT4 #(
		.INIT('hd070)
	) name3639 (
		\P1_state_reg[0]/NET0131 ,
		\P2_IR_reg[23]/NET0131 ,
		\P2_reg1_reg[21]/NET0131 ,
		_w1188_,
		_w4102_
	);
	LUT4 #(
		.INIT('h2000)
	) name3640 (
		\P2_reg1_reg[21]/NET0131 ,
		_w1189_,
		_w1352_,
		_w1356_,
		_w4103_
	);
	LUT4 #(
		.INIT('h020e)
	) name3641 (
		\P2_reg1_reg[21]/NET0131 ,
		_w1516_,
		_w1575_,
		_w3281_,
		_w4104_
	);
	LUT3 #(
		.INIT('ha2)
	) name3642 (
		\P2_reg1_reg[21]/NET0131 ,
		_w1684_,
		_w2469_,
		_w4105_
	);
	LUT3 #(
		.INIT('h07)
	) name3643 (
		_w1516_,
		_w3283_,
		_w4105_,
		_w4106_
	);
	LUT2 #(
		.INIT('h4)
	) name3644 (
		_w4104_,
		_w4106_,
		_w4107_
	);
	LUT4 #(
		.INIT('h08c8)
	) name3645 (
		\P2_reg1_reg[21]/NET0131 ,
		_w1191_,
		_w1507_,
		_w3289_,
		_w4108_
	);
	LUT4 #(
		.INIT('h0232)
	) name3646 (
		\P2_reg1_reg[21]/NET0131 ,
		_w1506_,
		_w1516_,
		_w3291_,
		_w4109_
	);
	LUT4 #(
		.INIT('h20e0)
	) name3647 (
		\P2_reg1_reg[21]/NET0131 ,
		_w1507_,
		_w1530_,
		_w3291_,
		_w4110_
	);
	LUT3 #(
		.INIT('h01)
	) name3648 (
		_w4109_,
		_w4110_,
		_w4108_,
		_w4111_
	);
	LUT4 #(
		.INIT('h3111)
	) name3649 (
		_w1359_,
		_w4103_,
		_w4107_,
		_w4111_,
		_w4112_
	);
	LUT3 #(
		.INIT('hce)
	) name3650 (
		\P1_state_reg[0]/NET0131 ,
		_w4102_,
		_w4112_,
		_w4113_
	);
	LUT2 #(
		.INIT('h2)
	) name3651 (
		\P1_reg0_reg[17]/NET0131 ,
		_w2462_,
		_w4114_
	);
	LUT4 #(
		.INIT('h2000)
	) name3652 (
		\P1_reg0_reg[17]/NET0131 ,
		_w1723_,
		_w1727_,
		_w1730_,
		_w4115_
	);
	LUT2 #(
		.INIT('h2)
	) name3653 (
		\P1_reg0_reg[17]/NET0131 ,
		_w2883_,
		_w4116_
	);
	LUT4 #(
		.INIT('hc048)
	) name3654 (
		_w2336_,
		_w2883_,
		_w3170_,
		_w3486_,
		_w4117_
	);
	LUT3 #(
		.INIT('ha8)
	) name3655 (
		_w2388_,
		_w4116_,
		_w4117_,
		_w4118_
	);
	LUT4 #(
		.INIT('h1dd1)
	) name3656 (
		\P1_reg0_reg[17]/NET0131 ,
		_w2883_,
		_w3170_,
		_w3489_,
		_w4119_
	);
	LUT4 #(
		.INIT('hc808)
	) name3657 (
		\P1_reg0_reg[17]/NET0131 ,
		_w2424_,
		_w2883_,
		_w3492_,
		_w4120_
	);
	LUT2 #(
		.INIT('h2)
	) name3658 (
		\P1_reg0_reg[17]/NET0131 ,
		_w3420_,
		_w4121_
	);
	LUT4 #(
		.INIT('h00fb)
	) name3659 (
		_w2436_,
		_w2447_,
		_w3495_,
		_w3903_,
		_w4122_
	);
	LUT3 #(
		.INIT('h31)
	) name3660 (
		_w2883_,
		_w4121_,
		_w4122_,
		_w4123_
	);
	LUT4 #(
		.INIT('h0d00)
	) name3661 (
		_w2292_,
		_w4119_,
		_w4120_,
		_w4123_,
		_w4124_
	);
	LUT4 #(
		.INIT('h1311)
	) name3662 (
		_w1731_,
		_w4115_,
		_w4118_,
		_w4124_,
		_w4125_
	);
	LUT3 #(
		.INIT('hce)
	) name3663 (
		\P1_state_reg[0]/NET0131 ,
		_w4114_,
		_w4125_,
		_w4126_
	);
	LUT2 #(
		.INIT('h2)
	) name3664 (
		\P1_reg0_reg[18]/NET0131 ,
		_w2462_,
		_w4127_
	);
	LUT4 #(
		.INIT('h2000)
	) name3665 (
		\P1_reg0_reg[18]/NET0131 ,
		_w1723_,
		_w1727_,
		_w1730_,
		_w4128_
	);
	LUT4 #(
		.INIT('hddd1)
	) name3666 (
		\P1_reg0_reg[18]/NET0131 ,
		_w2883_,
		_w3466_,
		_w3467_,
		_w4129_
	);
	LUT2 #(
		.INIT('h2)
	) name3667 (
		_w2424_,
		_w4129_,
		_w4130_
	);
	LUT4 #(
		.INIT('hd11d)
	) name3668 (
		\P1_reg0_reg[18]/NET0131 ,
		_w2883_,
		_w2940_,
		_w3181_,
		_w4131_
	);
	LUT2 #(
		.INIT('h2)
	) name3669 (
		_w2388_,
		_w4131_,
		_w4132_
	);
	LUT4 #(
		.INIT('h1dd1)
	) name3670 (
		\P1_reg0_reg[18]/NET0131 ,
		_w2883_,
		_w2958_,
		_w3181_,
		_w4133_
	);
	LUT4 #(
		.INIT('h0a8a)
	) name3671 (
		\P1_reg0_reg[18]/NET0131 ,
		_w2452_,
		_w2524_,
		_w2883_,
		_w4134_
	);
	LUT3 #(
		.INIT('h07)
	) name3672 (
		_w2883_,
		_w3473_,
		_w4134_,
		_w4135_
	);
	LUT3 #(
		.INIT('hd0)
	) name3673 (
		_w2292_,
		_w4133_,
		_w4135_,
		_w4136_
	);
	LUT4 #(
		.INIT('ha8aa)
	) name3674 (
		_w1731_,
		_w4130_,
		_w4132_,
		_w4136_,
		_w4137_
	);
	LUT4 #(
		.INIT('heeec)
	) name3675 (
		\P1_state_reg[0]/NET0131 ,
		_w4127_,
		_w4128_,
		_w4137_,
		_w4138_
	);
	LUT2 #(
		.INIT('h2)
	) name3676 (
		\P1_reg0_reg[19]/NET0131 ,
		_w2462_,
		_w4139_
	);
	LUT4 #(
		.INIT('h2000)
	) name3677 (
		\P1_reg0_reg[19]/NET0131 ,
		_w1723_,
		_w1727_,
		_w1730_,
		_w4140_
	);
	LUT4 #(
		.INIT('hc808)
	) name3678 (
		\P1_reg0_reg[19]/NET0131 ,
		_w2424_,
		_w2883_,
		_w3510_,
		_w4141_
	);
	LUT4 #(
		.INIT('hc535)
	) name3679 (
		\P1_reg0_reg[19]/NET0131 ,
		_w2662_,
		_w2883_,
		_w3165_,
		_w4142_
	);
	LUT2 #(
		.INIT('h2)
	) name3680 (
		_w2292_,
		_w4142_,
		_w4143_
	);
	LUT4 #(
		.INIT('h35c5)
	) name3681 (
		\P1_reg0_reg[19]/NET0131 ,
		_w2675_,
		_w2883_,
		_w3165_,
		_w4144_
	);
	LUT4 #(
		.INIT('h0a8a)
	) name3682 (
		\P1_reg0_reg[19]/NET0131 ,
		_w2452_,
		_w2524_,
		_w2883_,
		_w4145_
	);
	LUT4 #(
		.INIT('h0057)
	) name3683 (
		_w2883_,
		_w3515_,
		_w3516_,
		_w4145_,
		_w4146_
	);
	LUT3 #(
		.INIT('hd0)
	) name3684 (
		_w2388_,
		_w4144_,
		_w4146_,
		_w4147_
	);
	LUT4 #(
		.INIT('ha8aa)
	) name3685 (
		_w1731_,
		_w4141_,
		_w4143_,
		_w4147_,
		_w4148_
	);
	LUT4 #(
		.INIT('heeec)
	) name3686 (
		\P1_state_reg[0]/NET0131 ,
		_w4139_,
		_w4140_,
		_w4148_,
		_w4149_
	);
	LUT2 #(
		.INIT('h2)
	) name3687 (
		\P1_reg0_reg[21]/NET0131 ,
		_w2462_,
		_w4150_
	);
	LUT4 #(
		.INIT('h2000)
	) name3688 (
		\P1_reg0_reg[21]/NET0131 ,
		_w1723_,
		_w1727_,
		_w1730_,
		_w4151_
	);
	LUT4 #(
		.INIT('hd11d)
	) name3689 (
		\P1_reg0_reg[21]/NET0131 ,
		_w2883_,
		_w3160_,
		_w3835_,
		_w4152_
	);
	LUT4 #(
		.INIT('h35c5)
	) name3690 (
		\P1_reg0_reg[21]/NET0131 ,
		_w2262_,
		_w2883_,
		_w3160_,
		_w4153_
	);
	LUT4 #(
		.INIT('h222a)
	) name3691 (
		\P1_reg0_reg[21]/NET0131 ,
		_w2524_,
		_w2883_,
		_w3843_,
		_w4154_
	);
	LUT4 #(
		.INIT('h005d)
	) name3692 (
		_w2883_,
		_w3842_,
		_w3872_,
		_w4154_,
		_w4155_
	);
	LUT3 #(
		.INIT('hd0)
	) name3693 (
		_w2292_,
		_w4153_,
		_w4155_,
		_w4156_
	);
	LUT4 #(
		.INIT('h08aa)
	) name3694 (
		_w1731_,
		_w2388_,
		_w4152_,
		_w4156_,
		_w4157_
	);
	LUT4 #(
		.INIT('heeec)
	) name3695 (
		\P1_state_reg[0]/NET0131 ,
		_w4150_,
		_w4151_,
		_w4157_,
		_w4158_
	);
	LUT2 #(
		.INIT('h2)
	) name3696 (
		\P1_reg0_reg[31]/NET0131 ,
		_w2462_,
		_w4159_
	);
	LUT4 #(
		.INIT('h2000)
	) name3697 (
		\P1_reg0_reg[31]/NET0131 ,
		_w1723_,
		_w1727_,
		_w1730_,
		_w4160_
	);
	LUT4 #(
		.INIT('h1dd1)
	) name3698 (
		\P1_reg0_reg[31]/NET0131 ,
		_w2883_,
		_w3126_,
		_w3566_,
		_w4161_
	);
	LUT2 #(
		.INIT('h8)
	) name3699 (
		_w2424_,
		_w2883_,
		_w4162_
	);
	LUT4 #(
		.INIT('h7000)
	) name3700 (
		_w2922_,
		_w3569_,
		_w3570_,
		_w4162_,
		_w4163_
	);
	LUT4 #(
		.INIT('hc5f5)
	) name3701 (
		\P1_reg0_reg[31]/NET0131 ,
		_w1748_,
		_w2883_,
		_w3125_,
		_w4164_
	);
	LUT2 #(
		.INIT('h1)
	) name3702 (
		_w2883_,
		_w3574_,
		_w4165_
	);
	LUT4 #(
		.INIT('h222a)
	) name3703 (
		\P1_reg0_reg[31]/NET0131 ,
		_w2524_,
		_w2883_,
		_w3574_,
		_w4166_
	);
	LUT3 #(
		.INIT('h0d)
	) name3704 (
		_w2426_,
		_w4164_,
		_w4166_,
		_w4167_
	);
	LUT4 #(
		.INIT('h0d00)
	) name3705 (
		_w2447_,
		_w4161_,
		_w4163_,
		_w4167_,
		_w4168_
	);
	LUT4 #(
		.INIT('ha0a8)
	) name3706 (
		\P1_state_reg[0]/NET0131 ,
		_w1731_,
		_w4160_,
		_w4168_,
		_w4169_
	);
	LUT2 #(
		.INIT('he)
	) name3707 (
		_w4159_,
		_w4169_,
		_w4170_
	);
	LUT2 #(
		.INIT('h2)
	) name3708 (
		\P1_reg1_reg[17]/NET0131 ,
		_w2462_,
		_w4171_
	);
	LUT4 #(
		.INIT('h2000)
	) name3709 (
		\P1_reg1_reg[17]/NET0131 ,
		_w1723_,
		_w1727_,
		_w1730_,
		_w4172_
	);
	LUT2 #(
		.INIT('h2)
	) name3710 (
		\P1_reg1_reg[17]/NET0131 ,
		_w2520_,
		_w4173_
	);
	LUT4 #(
		.INIT('hc048)
	) name3711 (
		_w2336_,
		_w2520_,
		_w3170_,
		_w3486_,
		_w4174_
	);
	LUT3 #(
		.INIT('ha8)
	) name3712 (
		_w2388_,
		_w4173_,
		_w4174_,
		_w4175_
	);
	LUT4 #(
		.INIT('h1dd1)
	) name3713 (
		\P1_reg1_reg[17]/NET0131 ,
		_w2520_,
		_w3170_,
		_w3489_,
		_w4176_
	);
	LUT4 #(
		.INIT('hc808)
	) name3714 (
		\P1_reg1_reg[17]/NET0131 ,
		_w2424_,
		_w2520_,
		_w3492_,
		_w4177_
	);
	LUT2 #(
		.INIT('h2)
	) name3715 (
		\P1_reg1_reg[17]/NET0131 ,
		_w2525_,
		_w4178_
	);
	LUT3 #(
		.INIT('h0d)
	) name3716 (
		_w2520_,
		_w4122_,
		_w4178_,
		_w4179_
	);
	LUT4 #(
		.INIT('h0d00)
	) name3717 (
		_w2292_,
		_w4176_,
		_w4177_,
		_w4179_,
		_w4180_
	);
	LUT4 #(
		.INIT('h1311)
	) name3718 (
		_w1731_,
		_w4172_,
		_w4175_,
		_w4180_,
		_w4181_
	);
	LUT3 #(
		.INIT('hce)
	) name3719 (
		\P1_state_reg[0]/NET0131 ,
		_w4171_,
		_w4181_,
		_w4182_
	);
	LUT2 #(
		.INIT('h2)
	) name3720 (
		\P1_reg1_reg[18]/NET0131 ,
		_w2462_,
		_w4183_
	);
	LUT4 #(
		.INIT('h2000)
	) name3721 (
		\P1_reg1_reg[18]/NET0131 ,
		_w1723_,
		_w1727_,
		_w1730_,
		_w4184_
	);
	LUT4 #(
		.INIT('hddd1)
	) name3722 (
		\P1_reg1_reg[18]/NET0131 ,
		_w2520_,
		_w3466_,
		_w3467_,
		_w4185_
	);
	LUT2 #(
		.INIT('h2)
	) name3723 (
		_w2424_,
		_w4185_,
		_w4186_
	);
	LUT4 #(
		.INIT('hd11d)
	) name3724 (
		\P1_reg1_reg[18]/NET0131 ,
		_w2520_,
		_w2940_,
		_w3181_,
		_w4187_
	);
	LUT2 #(
		.INIT('h2)
	) name3725 (
		_w2388_,
		_w4187_,
		_w4188_
	);
	LUT4 #(
		.INIT('h1dd1)
	) name3726 (
		\P1_reg1_reg[18]/NET0131 ,
		_w2520_,
		_w2958_,
		_w3181_,
		_w4189_
	);
	LUT4 #(
		.INIT('h08aa)
	) name3727 (
		\P1_reg1_reg[18]/NET0131 ,
		_w2452_,
		_w2520_,
		_w2524_,
		_w4190_
	);
	LUT3 #(
		.INIT('h07)
	) name3728 (
		_w2520_,
		_w3473_,
		_w4190_,
		_w4191_
	);
	LUT3 #(
		.INIT('hd0)
	) name3729 (
		_w2292_,
		_w4189_,
		_w4191_,
		_w4192_
	);
	LUT4 #(
		.INIT('ha8aa)
	) name3730 (
		_w1731_,
		_w4186_,
		_w4188_,
		_w4192_,
		_w4193_
	);
	LUT4 #(
		.INIT('heeec)
	) name3731 (
		\P1_state_reg[0]/NET0131 ,
		_w4183_,
		_w4184_,
		_w4193_,
		_w4194_
	);
	LUT2 #(
		.INIT('h2)
	) name3732 (
		\P1_reg1_reg[19]/NET0131 ,
		_w2462_,
		_w4195_
	);
	LUT4 #(
		.INIT('h2000)
	) name3733 (
		\P1_reg1_reg[19]/NET0131 ,
		_w1723_,
		_w1727_,
		_w1730_,
		_w4196_
	);
	LUT4 #(
		.INIT('hc808)
	) name3734 (
		\P1_reg1_reg[19]/NET0131 ,
		_w2424_,
		_w2520_,
		_w3510_,
		_w4197_
	);
	LUT4 #(
		.INIT('hd11d)
	) name3735 (
		\P1_reg1_reg[19]/NET0131 ,
		_w2520_,
		_w2662_,
		_w3165_,
		_w4198_
	);
	LUT2 #(
		.INIT('h2)
	) name3736 (
		_w2292_,
		_w4198_,
		_w4199_
	);
	LUT4 #(
		.INIT('h1dd1)
	) name3737 (
		\P1_reg1_reg[19]/NET0131 ,
		_w2520_,
		_w2675_,
		_w3165_,
		_w4200_
	);
	LUT4 #(
		.INIT('h08aa)
	) name3738 (
		\P1_reg1_reg[19]/NET0131 ,
		_w2452_,
		_w2520_,
		_w2524_,
		_w4201_
	);
	LUT4 #(
		.INIT('h0057)
	) name3739 (
		_w2520_,
		_w3515_,
		_w3516_,
		_w4201_,
		_w4202_
	);
	LUT3 #(
		.INIT('hd0)
	) name3740 (
		_w2388_,
		_w4200_,
		_w4202_,
		_w4203_
	);
	LUT4 #(
		.INIT('ha8aa)
	) name3741 (
		_w1731_,
		_w4197_,
		_w4199_,
		_w4203_,
		_w4204_
	);
	LUT4 #(
		.INIT('heeec)
	) name3742 (
		\P1_state_reg[0]/NET0131 ,
		_w4195_,
		_w4196_,
		_w4204_,
		_w4205_
	);
	LUT2 #(
		.INIT('h2)
	) name3743 (
		\P1_reg1_reg[21]/NET0131 ,
		_w2462_,
		_w4206_
	);
	LUT4 #(
		.INIT('h2000)
	) name3744 (
		\P1_reg1_reg[21]/NET0131 ,
		_w1723_,
		_w1727_,
		_w1730_,
		_w4207_
	);
	LUT4 #(
		.INIT('hd11d)
	) name3745 (
		\P1_reg1_reg[21]/NET0131 ,
		_w2520_,
		_w3160_,
		_w3835_,
		_w4208_
	);
	LUT4 #(
		.INIT('h35c5)
	) name3746 (
		\P1_reg1_reg[21]/NET0131 ,
		_w2262_,
		_w2520_,
		_w3160_,
		_w4209_
	);
	LUT4 #(
		.INIT('h0a2a)
	) name3747 (
		\P1_reg1_reg[21]/NET0131 ,
		_w2520_,
		_w2524_,
		_w3843_,
		_w4210_
	);
	LUT4 #(
		.INIT('h005d)
	) name3748 (
		_w2520_,
		_w3842_,
		_w3872_,
		_w4210_,
		_w4211_
	);
	LUT3 #(
		.INIT('hd0)
	) name3749 (
		_w2292_,
		_w4209_,
		_w4211_,
		_w4212_
	);
	LUT4 #(
		.INIT('h08aa)
	) name3750 (
		_w1731_,
		_w2388_,
		_w4208_,
		_w4212_,
		_w4213_
	);
	LUT4 #(
		.INIT('heeec)
	) name3751 (
		\P1_state_reg[0]/NET0131 ,
		_w4206_,
		_w4207_,
		_w4213_,
		_w4214_
	);
	LUT4 #(
		.INIT('h4000)
	) name3752 (
		_w1723_,
		_w1727_,
		_w1730_,
		_w2032_,
		_w4215_
	);
	LUT2 #(
		.INIT('h2)
	) name3753 (
		_w2032_,
		_w2644_,
		_w4216_
	);
	LUT4 #(
		.INIT('h4144)
	) name3754 (
		_w1747_,
		_w2008_,
		_w2034_,
		_w2404_,
		_w4217_
	);
	LUT3 #(
		.INIT('h80)
	) name3755 (
		_w1747_,
		_w2041_,
		_w2043_,
		_w4218_
	);
	LUT4 #(
		.INIT('h3331)
	) name3756 (
		_w2644_,
		_w4216_,
		_w4217_,
		_w4218_,
		_w4219_
	);
	LUT2 #(
		.INIT('h2)
	) name3757 (
		_w2424_,
		_w4219_,
		_w4220_
	);
	LUT4 #(
		.INIT('h00d7)
	) name3758 (
		_w2644_,
		_w2935_,
		_w3176_,
		_w4216_,
		_w4221_
	);
	LUT2 #(
		.INIT('h2)
	) name3759 (
		_w2388_,
		_w4221_,
		_w4222_
	);
	LUT4 #(
		.INIT('h007d)
	) name3760 (
		_w2644_,
		_w2953_,
		_w3176_,
		_w4216_,
		_w4223_
	);
	LUT4 #(
		.INIT('h5655)
	) name3761 (
		_w2029_,
		_w2040_,
		_w2104_,
		_w2431_,
		_w4224_
	);
	LUT4 #(
		.INIT('hc808)
	) name3762 (
		_w2032_,
		_w2447_,
		_w2644_,
		_w4224_,
		_w4225_
	);
	LUT4 #(
		.INIT('ha8a0)
	) name3763 (
		_w2029_,
		_w2426_,
		_w2454_,
		_w2644_,
		_w4226_
	);
	LUT4 #(
		.INIT('ha0a8)
	) name3764 (
		_w2032_,
		_w2426_,
		_w2450_,
		_w2644_,
		_w4227_
	);
	LUT2 #(
		.INIT('h1)
	) name3765 (
		_w4226_,
		_w4227_,
		_w4228_
	);
	LUT2 #(
		.INIT('h4)
	) name3766 (
		_w4225_,
		_w4228_,
		_w4229_
	);
	LUT3 #(
		.INIT('hd0)
	) name3767 (
		_w2292_,
		_w4223_,
		_w4229_,
		_w4230_
	);
	LUT4 #(
		.INIT('ha8aa)
	) name3768 (
		_w1731_,
		_w4220_,
		_w4222_,
		_w4230_,
		_w4231_
	);
	LUT2 #(
		.INIT('h2)
	) name3769 (
		\P1_reg3_reg[10]/NET0131 ,
		\P1_state_reg[0]/NET0131 ,
		_w4232_
	);
	LUT3 #(
		.INIT('h07)
	) name3770 (
		_w2032_,
		_w2695_,
		_w4232_,
		_w4233_
	);
	LUT4 #(
		.INIT('ha8ff)
	) name3771 (
		\P1_state_reg[0]/NET0131 ,
		_w4215_,
		_w4231_,
		_w4233_,
		_w4234_
	);
	LUT4 #(
		.INIT('h4000)
	) name3772 (
		_w1723_,
		_w1727_,
		_w1730_,
		_w2220_,
		_w4235_
	);
	LUT2 #(
		.INIT('h2)
	) name3773 (
		_w2220_,
		_w2644_,
		_w4236_
	);
	LUT4 #(
		.INIT('h6555)
	) name3774 (
		_w2212_,
		_w2223_,
		_w2404_,
		_w2406_,
		_w4237_
	);
	LUT4 #(
		.INIT('h7020)
	) name3775 (
		_w1747_,
		_w2020_,
		_w2644_,
		_w4237_,
		_w4238_
	);
	LUT4 #(
		.INIT('h7f00)
	) name3776 (
		_w2431_,
		_w2432_,
		_w2434_,
		_w2447_,
		_w4239_
	);
	LUT4 #(
		.INIT('hd500)
	) name3777 (
		_w2219_,
		_w2432_,
		_w3804_,
		_w4239_,
		_w4240_
	);
	LUT4 #(
		.INIT('ha8a0)
	) name3778 (
		_w2219_,
		_w2426_,
		_w2454_,
		_w2644_,
		_w4241_
	);
	LUT3 #(
		.INIT('h0d)
	) name3779 (
		_w2220_,
		_w2690_,
		_w4241_,
		_w4242_
	);
	LUT3 #(
		.INIT('h70)
	) name3780 (
		_w2644_,
		_w4240_,
		_w4242_,
		_w4243_
	);
	LUT4 #(
		.INIT('h5700)
	) name3781 (
		_w2424_,
		_w4236_,
		_w4238_,
		_w4243_,
		_w4244_
	);
	LUT4 #(
		.INIT('h8a75)
	) name3782 (
		_w2301_,
		_w2327_,
		_w2330_,
		_w3192_,
		_w4245_
	);
	LUT4 #(
		.INIT('h08c8)
	) name3783 (
		_w2220_,
		_w2388_,
		_w2644_,
		_w4245_,
		_w4246_
	);
	LUT4 #(
		.INIT('h20d0)
	) name3784 (
		_w2049_,
		_w2153_,
		_w2644_,
		_w3192_,
		_w4247_
	);
	LUT3 #(
		.INIT('ha8)
	) name3785 (
		_w2292_,
		_w4236_,
		_w4247_,
		_w4248_
	);
	LUT4 #(
		.INIT('ha8aa)
	) name3786 (
		_w1731_,
		_w4246_,
		_w4248_,
		_w4244_,
		_w4249_
	);
	LUT2 #(
		.INIT('h2)
	) name3787 (
		\P1_reg3_reg[13]/NET0131 ,
		\P1_state_reg[0]/NET0131 ,
		_w4250_
	);
	LUT3 #(
		.INIT('h07)
	) name3788 (
		_w2220_,
		_w2695_,
		_w4250_,
		_w4251_
	);
	LUT4 #(
		.INIT('ha8ff)
	) name3789 (
		\P1_state_reg[0]/NET0131 ,
		_w4235_,
		_w4249_,
		_w4251_,
		_w4252_
	);
	LUT4 #(
		.INIT('h1000)
	) name3790 (
		_w690_,
		_w1189_,
		_w1352_,
		_w1356_,
		_w4253_
	);
	LUT4 #(
		.INIT('h5554)
	) name3791 (
		_w690_,
		_w1361_,
		_w1363_,
		_w1368_,
		_w4254_
	);
	LUT3 #(
		.INIT('h10)
	) name3792 (
		_w693_,
		_w711_,
		_w1418_,
		_w4255_
	);
	LUT4 #(
		.INIT('h0100)
	) name3793 (
		_w679_,
		_w693_,
		_w711_,
		_w1418_,
		_w4256_
	);
	LUT2 #(
		.INIT('h1)
	) name3794 (
		_w711_,
		_w1435_,
		_w4257_
	);
	LUT4 #(
		.INIT('h007b)
	) name3795 (
		_w679_,
		_w1435_,
		_w4255_,
		_w4257_,
		_w4258_
	);
	LUT4 #(
		.INIT('h04c4)
	) name3796 (
		_w690_,
		_w1191_,
		_w1411_,
		_w4258_,
		_w4259_
	);
	LUT4 #(
		.INIT('h0155)
	) name3797 (
		_w690_,
		_w1361_,
		_w1363_,
		_w1368_,
		_w4260_
	);
	LUT4 #(
		.INIT('h8848)
	) name3798 (
		_w1317_,
		_w1369_,
		_w2553_,
		_w2555_,
		_w4261_
	);
	LUT3 #(
		.INIT('h04)
	) name3799 (
		_w703_,
		_w1232_,
		_w1439_,
		_w4262_
	);
	LUT3 #(
		.INIT('h54)
	) name3800 (
		_w690_,
		_w1441_,
		_w1443_,
		_w4263_
	);
	LUT2 #(
		.INIT('h1)
	) name3801 (
		_w4262_,
		_w4263_,
		_w4264_
	);
	LUT4 #(
		.INIT('hab00)
	) name3802 (
		_w1409_,
		_w4260_,
		_w4261_,
		_w4264_,
		_w4265_
	);
	LUT4 #(
		.INIT('h4844)
	) name3803 (
		_w1317_,
		_w1369_,
		_w2535_,
		_w2537_,
		_w4266_
	);
	LUT3 #(
		.INIT('h54)
	) name3804 (
		_w1496_,
		_w4260_,
		_w4266_,
		_w4267_
	);
	LUT4 #(
		.INIT('h4844)
	) name3805 (
		_w1317_,
		_w1411_,
		_w2535_,
		_w2537_,
		_w4268_
	);
	LUT3 #(
		.INIT('ha8)
	) name3806 (
		_w1447_,
		_w4254_,
		_w4268_,
		_w4269_
	);
	LUT4 #(
		.INIT('h0100)
	) name3807 (
		_w4267_,
		_w4269_,
		_w4259_,
		_w4265_,
		_w4270_
	);
	LUT4 #(
		.INIT('ha0a8)
	) name3808 (
		\P1_state_reg[0]/NET0131 ,
		_w1359_,
		_w4253_,
		_w4270_,
		_w4271_
	);
	LUT2 #(
		.INIT('h4)
	) name3809 (
		\P1_state_reg[0]/NET0131 ,
		\P2_reg3_reg[10]/NET0131 ,
		_w4272_
	);
	LUT4 #(
		.INIT('h0802)
	) name3810 (
		\P1_state_reg[0]/NET0131 ,
		\P2_IR_reg[23]/NET0131 ,
		_w690_,
		_w1188_,
		_w4273_
	);
	LUT2 #(
		.INIT('h1)
	) name3811 (
		_w4272_,
		_w4273_,
		_w4274_
	);
	LUT2 #(
		.INIT('hb)
	) name3812 (
		_w4271_,
		_w4274_,
		_w4275_
	);
	LUT4 #(
		.INIT('h1000)
	) name3813 (
		_w648_,
		_w1189_,
		_w1352_,
		_w1356_,
		_w4276_
	);
	LUT4 #(
		.INIT('hb04f)
	) name3814 (
		_w1215_,
		_w1216_,
		_w1205_,
		_w1302_,
		_w4277_
	);
	LUT4 #(
		.INIT('h010d)
	) name3815 (
		_w648_,
		_w1369_,
		_w1409_,
		_w4277_,
		_w4278_
	);
	LUT4 #(
		.INIT('h5554)
	) name3816 (
		_w648_,
		_w1361_,
		_w1363_,
		_w1368_,
		_w4279_
	);
	LUT4 #(
		.INIT('h9500)
	) name3817 (
		_w631_,
		_w1418_,
		_w1419_,
		_w1435_,
		_w4280_
	);
	LUT2 #(
		.INIT('h1)
	) name3818 (
		_w679_,
		_w1435_,
		_w4281_
	);
	LUT4 #(
		.INIT('h1113)
	) name3819 (
		_w1411_,
		_w4279_,
		_w4280_,
		_w4281_,
		_w4282_
	);
	LUT3 #(
		.INIT('h04)
	) name3820 (
		_w666_,
		_w1232_,
		_w1439_,
		_w4283_
	);
	LUT3 #(
		.INIT('h54)
	) name3821 (
		_w648_,
		_w1441_,
		_w1443_,
		_w4284_
	);
	LUT2 #(
		.INIT('h1)
	) name3822 (
		_w4283_,
		_w4284_,
		_w4285_
	);
	LUT3 #(
		.INIT('hd0)
	) name3823 (
		_w1191_,
		_w4282_,
		_w4285_,
		_w4286_
	);
	LUT4 #(
		.INIT('h9a55)
	) name3824 (
		_w1302_,
		_w1537_,
		_w1539_,
		_w1543_,
		_w4287_
	);
	LUT4 #(
		.INIT('h0d01)
	) name3825 (
		_w648_,
		_w1369_,
		_w1496_,
		_w4287_,
		_w4288_
	);
	LUT4 #(
		.INIT('hc404)
	) name3826 (
		_w648_,
		_w1447_,
		_w1411_,
		_w4287_,
		_w4289_
	);
	LUT4 #(
		.INIT('h0100)
	) name3827 (
		_w4278_,
		_w4288_,
		_w4289_,
		_w4286_,
		_w4290_
	);
	LUT4 #(
		.INIT('ha0a8)
	) name3828 (
		\P1_state_reg[0]/NET0131 ,
		_w1359_,
		_w4276_,
		_w4290_,
		_w4291_
	);
	LUT2 #(
		.INIT('h4)
	) name3829 (
		\P1_state_reg[0]/NET0131 ,
		\P2_reg3_reg[12]/NET0131 ,
		_w4292_
	);
	LUT4 #(
		.INIT('h0802)
	) name3830 (
		\P1_state_reg[0]/NET0131 ,
		\P2_IR_reg[23]/NET0131 ,
		_w648_,
		_w1188_,
		_w4293_
	);
	LUT2 #(
		.INIT('h1)
	) name3831 (
		_w4292_,
		_w4293_,
		_w4294_
	);
	LUT2 #(
		.INIT('hb)
	) name3832 (
		_w4291_,
		_w4294_,
		_w4295_
	);
	LUT4 #(
		.INIT('h1000)
	) name3833 (
		_w627_,
		_w1189_,
		_w1352_,
		_w1356_,
		_w4296_
	);
	LUT4 #(
		.INIT('h5554)
	) name3834 (
		_w627_,
		_w1361_,
		_w1363_,
		_w1368_,
		_w4297_
	);
	LUT4 #(
		.INIT('h00b7)
	) name3835 (
		_w1299_,
		_w1411_,
		_w1699_,
		_w4297_,
		_w4298_
	);
	LUT4 #(
		.INIT('h1000)
	) name3836 (
		_w623_,
		_w631_,
		_w1418_,
		_w1419_,
		_w4299_
	);
	LUT2 #(
		.INIT('h1)
	) name3837 (
		_w653_,
		_w1435_,
		_w4300_
	);
	LUT4 #(
		.INIT('h006f)
	) name3838 (
		_w623_,
		_w1420_,
		_w1435_,
		_w4300_,
		_w4301_
	);
	LUT4 #(
		.INIT('h04c4)
	) name3839 (
		_w627_,
		_w1191_,
		_w1411_,
		_w4301_,
		_w4302_
	);
	LUT3 #(
		.INIT('h04)
	) name3840 (
		_w645_,
		_w1232_,
		_w1439_,
		_w4303_
	);
	LUT3 #(
		.INIT('h54)
	) name3841 (
		_w627_,
		_w1441_,
		_w1443_,
		_w4304_
	);
	LUT2 #(
		.INIT('h1)
	) name3842 (
		_w4303_,
		_w4304_,
		_w4305_
	);
	LUT4 #(
		.INIT('h0d00)
	) name3843 (
		_w1447_,
		_w4298_,
		_w4302_,
		_w4305_,
		_w4306_
	);
	LUT4 #(
		.INIT('h0155)
	) name3844 (
		_w627_,
		_w1361_,
		_w1363_,
		_w1368_,
		_w4307_
	);
	LUT4 #(
		.INIT('h00b7)
	) name3845 (
		_w1299_,
		_w1369_,
		_w1699_,
		_w4307_,
		_w4308_
	);
	LUT4 #(
		.INIT('h9599)
	) name3846 (
		_w1299_,
		_w1660_,
		_w1662_,
		_w1663_,
		_w4309_
	);
	LUT4 #(
		.INIT('h0d01)
	) name3847 (
		_w627_,
		_w1369_,
		_w1409_,
		_w4309_,
		_w4310_
	);
	LUT3 #(
		.INIT('h0e)
	) name3848 (
		_w1496_,
		_w4308_,
		_w4310_,
		_w4311_
	);
	LUT4 #(
		.INIT('h3111)
	) name3849 (
		_w1359_,
		_w4296_,
		_w4306_,
		_w4311_,
		_w4312_
	);
	LUT2 #(
		.INIT('h4)
	) name3850 (
		\P1_state_reg[0]/NET0131 ,
		\P2_reg3_reg[13]/NET0131 ,
		_w4313_
	);
	LUT4 #(
		.INIT('h0802)
	) name3851 (
		\P1_state_reg[0]/NET0131 ,
		\P2_IR_reg[23]/NET0131 ,
		_w627_,
		_w1188_,
		_w4314_
	);
	LUT2 #(
		.INIT('h1)
	) name3852 (
		_w4313_,
		_w4314_,
		_w4315_
	);
	LUT3 #(
		.INIT('h2f)
	) name3853 (
		\P1_state_reg[0]/NET0131 ,
		_w4312_,
		_w4315_,
		_w4316_
	);
	LUT4 #(
		.INIT('h4000)
	) name3854 (
		_w1723_,
		_w1727_,
		_w1730_,
		_w2042_,
		_w4317_
	);
	LUT2 #(
		.INIT('h2)
	) name3855 (
		_w2042_,
		_w2644_,
		_w4318_
	);
	LUT4 #(
		.INIT('h007b)
	) name3856 (
		_w2327_,
		_w2644_,
		_w3186_,
		_w4318_,
		_w4319_
	);
	LUT4 #(
		.INIT('h6500)
	) name3857 (
		_w2040_,
		_w2104_,
		_w2431_,
		_w2644_,
		_w4320_
	);
	LUT4 #(
		.INIT('ha8a0)
	) name3858 (
		_w2040_,
		_w2426_,
		_w2454_,
		_w2644_,
		_w4321_
	);
	LUT4 #(
		.INIT('ha0a8)
	) name3859 (
		_w2042_,
		_w2426_,
		_w2450_,
		_w2644_,
		_w4322_
	);
	LUT2 #(
		.INIT('h1)
	) name3860 (
		_w4321_,
		_w4322_,
		_w4323_
	);
	LUT4 #(
		.INIT('h5700)
	) name3861 (
		_w2447_,
		_w4318_,
		_w4320_,
		_w4323_,
		_w4324_
	);
	LUT3 #(
		.INIT('hd0)
	) name3862 (
		_w2388_,
		_w4319_,
		_w4324_,
		_w4325_
	);
	LUT4 #(
		.INIT('h708f)
	) name3863 (
		_w2096_,
		_w2142_,
		_w2149_,
		_w3186_,
		_w4326_
	);
	LUT4 #(
		.INIT('h08c8)
	) name3864 (
		_w2042_,
		_w2292_,
		_w2644_,
		_w4326_,
		_w4327_
	);
	LUT3 #(
		.INIT('h80)
	) name3865 (
		_w1747_,
		_w2105_,
		_w2107_,
		_w4328_
	);
	LUT4 #(
		.INIT('h00eb)
	) name3866 (
		_w1747_,
		_w2034_,
		_w2404_,
		_w4328_,
		_w4329_
	);
	LUT4 #(
		.INIT('hc808)
	) name3867 (
		_w2042_,
		_w2424_,
		_w2644_,
		_w4329_,
		_w4330_
	);
	LUT2 #(
		.INIT('h1)
	) name3868 (
		_w4327_,
		_w4330_,
		_w4331_
	);
	LUT4 #(
		.INIT('h3111)
	) name3869 (
		_w1731_,
		_w4317_,
		_w4325_,
		_w4331_,
		_w4332_
	);
	LUT2 #(
		.INIT('h2)
	) name3870 (
		\P1_reg3_reg[9]/NET0131 ,
		\P1_state_reg[0]/NET0131 ,
		_w4333_
	);
	LUT3 #(
		.INIT('h07)
	) name3871 (
		_w2042_,
		_w2695_,
		_w4333_,
		_w4334_
	);
	LUT3 #(
		.INIT('h2f)
	) name3872 (
		\P1_state_reg[0]/NET0131 ,
		_w4332_,
		_w4334_,
		_w4335_
	);
	LUT4 #(
		.INIT('h1000)
	) name3873 (
		_w707_,
		_w1189_,
		_w1352_,
		_w1356_,
		_w4336_
	);
	LUT4 #(
		.INIT('h5554)
	) name3874 (
		_w707_,
		_w1361_,
		_w1363_,
		_w1368_,
		_w4337_
	);
	LUT4 #(
		.INIT('h8488)
	) name3875 (
		_w1311_,
		_w1411_,
		_w1695_,
		_w1696_,
		_w4338_
	);
	LUT3 #(
		.INIT('h04)
	) name3876 (
		_w719_,
		_w1232_,
		_w1439_,
		_w4339_
	);
	LUT3 #(
		.INIT('h54)
	) name3877 (
		_w707_,
		_w1441_,
		_w1443_,
		_w4340_
	);
	LUT2 #(
		.INIT('h1)
	) name3878 (
		_w4339_,
		_w4340_,
		_w4341_
	);
	LUT4 #(
		.INIT('h5700)
	) name3879 (
		_w1447_,
		_w4337_,
		_w4338_,
		_w4341_,
		_w4342_
	);
	LUT4 #(
		.INIT('h0155)
	) name3880 (
		_w707_,
		_w1361_,
		_w1363_,
		_w1368_,
		_w4343_
	);
	LUT4 #(
		.INIT('h007b)
	) name3881 (
		_w1311_,
		_w1369_,
		_w1662_,
		_w4343_,
		_w4344_
	);
	LUT2 #(
		.INIT('h1)
	) name3882 (
		_w1409_,
		_w4344_,
		_w4345_
	);
	LUT4 #(
		.INIT('h6500)
	) name3883 (
		_w693_,
		_w711_,
		_w1418_,
		_w1435_,
		_w4346_
	);
	LUT2 #(
		.INIT('h1)
	) name3884 (
		_w726_,
		_w1435_,
		_w4347_
	);
	LUT4 #(
		.INIT('h1113)
	) name3885 (
		_w1411_,
		_w4337_,
		_w4346_,
		_w4347_,
		_w4348_
	);
	LUT2 #(
		.INIT('h2)
	) name3886 (
		_w1191_,
		_w4348_,
		_w4349_
	);
	LUT4 #(
		.INIT('h8488)
	) name3887 (
		_w1311_,
		_w1369_,
		_w1695_,
		_w1696_,
		_w4350_
	);
	LUT3 #(
		.INIT('h54)
	) name3888 (
		_w1496_,
		_w4343_,
		_w4350_,
		_w4351_
	);
	LUT4 #(
		.INIT('h0100)
	) name3889 (
		_w4349_,
		_w4351_,
		_w4345_,
		_w4342_,
		_w4352_
	);
	LUT4 #(
		.INIT('ha0a8)
	) name3890 (
		\P1_state_reg[0]/NET0131 ,
		_w1359_,
		_w4336_,
		_w4352_,
		_w4353_
	);
	LUT2 #(
		.INIT('h4)
	) name3891 (
		\P1_state_reg[0]/NET0131 ,
		\P2_reg3_reg[9]/NET0131 ,
		_w4354_
	);
	LUT4 #(
		.INIT('h0802)
	) name3892 (
		\P1_state_reg[0]/NET0131 ,
		\P2_IR_reg[23]/NET0131 ,
		_w707_,
		_w1188_,
		_w4355_
	);
	LUT2 #(
		.INIT('h1)
	) name3893 (
		_w4354_,
		_w4355_,
		_w4356_
	);
	LUT2 #(
		.INIT('hb)
	) name3894 (
		_w4353_,
		_w4356_,
		_w4357_
	);
	LUT4 #(
		.INIT('h4f00)
	) name3895 (
		_w2654_,
		_w2655_,
		_w2656_,
		_w2659_,
		_w4358_
	);
	LUT2 #(
		.INIT('h8)
	) name3896 (
		_w2657_,
		_w2663_,
		_w4359_
	);
	LUT2 #(
		.INIT('h4)
	) name3897 (
		_w2660_,
		_w2663_,
		_w4360_
	);
	LUT2 #(
		.INIT('h2)
	) name3898 (
		_w2647_,
		_w4360_,
		_w4361_
	);
	LUT4 #(
		.INIT('h65aa)
	) name3899 (
		_w3161_,
		_w4358_,
		_w4359_,
		_w4361_,
		_w4362_
	);
	LUT4 #(
		.INIT('h08c8)
	) name3900 (
		_w1959_,
		_w2292_,
		_w2644_,
		_w4362_,
		_w4363_
	);
	LUT4 #(
		.INIT('h4f00)
	) name3901 (
		_w2667_,
		_w2668_,
		_w2669_,
		_w2672_,
		_w4364_
	);
	LUT2 #(
		.INIT('h8)
	) name3902 (
		_w2670_,
		_w2676_,
		_w4365_
	);
	LUT2 #(
		.INIT('h4)
	) name3903 (
		_w2673_,
		_w2676_,
		_w4366_
	);
	LUT2 #(
		.INIT('h2)
	) name3904 (
		_w2679_,
		_w4366_,
		_w4367_
	);
	LUT4 #(
		.INIT('h9a55)
	) name3905 (
		_w3161_,
		_w4364_,
		_w4365_,
		_w4367_,
		_w4368_
	);
	LUT4 #(
		.INIT('h08c8)
	) name3906 (
		_w1959_,
		_w2388_,
		_w2644_,
		_w4368_,
		_w4369_
	);
	LUT3 #(
		.INIT('h80)
	) name3907 (
		_w1747_,
		_w1972_,
		_w1974_,
		_w4370_
	);
	LUT4 #(
		.INIT('h00eb)
	) name3908 (
		_w1747_,
		_w1952_,
		_w2985_,
		_w4370_,
		_w4371_
	);
	LUT4 #(
		.INIT('hc808)
	) name3909 (
		_w1959_,
		_w2424_,
		_w2644_,
		_w4371_,
		_w4372_
	);
	LUT3 #(
		.INIT('h10)
	) name3910 (
		_w1748_,
		_w1957_,
		_w2426_,
		_w4373_
	);
	LUT4 #(
		.INIT('h006f)
	) name3911 (
		_w1958_,
		_w2440_,
		_w2447_,
		_w4373_,
		_w4374_
	);
	LUT3 #(
		.INIT('h10)
	) name3912 (
		_w1748_,
		_w1957_,
		_w2454_,
		_w4375_
	);
	LUT4 #(
		.INIT('h88a8)
	) name3913 (
		_w1959_,
		_w2450_,
		_w2452_,
		_w2644_,
		_w4376_
	);
	LUT2 #(
		.INIT('h1)
	) name3914 (
		_w4375_,
		_w4376_,
		_w4377_
	);
	LUT3 #(
		.INIT('hd0)
	) name3915 (
		_w2644_,
		_w4374_,
		_w4377_,
		_w4378_
	);
	LUT2 #(
		.INIT('h4)
	) name3916 (
		_w4372_,
		_w4378_,
		_w4379_
	);
	LUT4 #(
		.INIT('ha8aa)
	) name3917 (
		_w1731_,
		_w4363_,
		_w4369_,
		_w4379_,
		_w4380_
	);
	LUT4 #(
		.INIT('h4000)
	) name3918 (
		_w1723_,
		_w1727_,
		_w1730_,
		_w1959_,
		_w4381_
	);
	LUT2 #(
		.INIT('h2)
	) name3919 (
		\P1_reg3_reg[23]/NET0131 ,
		\P1_state_reg[0]/NET0131 ,
		_w4382_
	);
	LUT3 #(
		.INIT('h07)
	) name3920 (
		_w1959_,
		_w2695_,
		_w4382_,
		_w4383_
	);
	LUT4 #(
		.INIT('ha8ff)
	) name3921 (
		\P1_state_reg[0]/NET0131 ,
		_w4380_,
		_w4381_,
		_w4383_,
		_w4384_
	);
	LUT2 #(
		.INIT('h2)
	) name3922 (
		\P1_reg2_reg[16]/NET0131 ,
		_w2462_,
		_w4385_
	);
	LUT4 #(
		.INIT('h2000)
	) name3923 (
		\P1_reg2_reg[16]/NET0131 ,
		_w1723_,
		_w1727_,
		_w1730_,
		_w4386_
	);
	LUT2 #(
		.INIT('h2)
	) name3924 (
		\P1_reg2_reg[16]/NET0131 ,
		_w1741_,
		_w4387_
	);
	LUT4 #(
		.INIT('h0a82)
	) name3925 (
		_w1741_,
		_w2768_,
		_w3168_,
		_w3817_,
		_w4388_
	);
	LUT3 #(
		.INIT('ha8)
	) name3926 (
		_w2292_,
		_w4387_,
		_w4388_,
		_w4389_
	);
	LUT4 #(
		.INIT('h20e0)
	) name3927 (
		\P1_reg2_reg[16]/NET0131 ,
		_w1741_,
		_w2388_,
		_w3820_,
		_w4390_
	);
	LUT4 #(
		.INIT('h2a08)
	) name3928 (
		_w1741_,
		_w1747_,
		_w2246_,
		_w3822_,
		_w4391_
	);
	LUT4 #(
		.INIT('h2822)
	) name3929 (
		_w1741_,
		_w2231_,
		_w2242_,
		_w3494_,
		_w4392_
	);
	LUT2 #(
		.INIT('h8)
	) name3930 (
		_w2231_,
		_w2426_,
		_w4393_
	);
	LUT3 #(
		.INIT('h80)
	) name3931 (
		_w1741_,
		_w2231_,
		_w2426_,
		_w4394_
	);
	LUT4 #(
		.INIT('haa20)
	) name3932 (
		\P1_reg2_reg[16]/NET0131 ,
		_w1741_,
		_w2426_,
		_w2450_,
		_w4395_
	);
	LUT4 #(
		.INIT('h0008)
	) name3933 (
		_w2233_,
		_w2284_,
		_w2288_,
		_w2291_,
		_w4396_
	);
	LUT3 #(
		.INIT('h01)
	) name3934 (
		_w4395_,
		_w4396_,
		_w4394_,
		_w4397_
	);
	LUT4 #(
		.INIT('h5700)
	) name3935 (
		_w2447_,
		_w4387_,
		_w4392_,
		_w4397_,
		_w4398_
	);
	LUT4 #(
		.INIT('h5700)
	) name3936 (
		_w2424_,
		_w4387_,
		_w4391_,
		_w4398_,
		_w4399_
	);
	LUT2 #(
		.INIT('h4)
	) name3937 (
		_w4390_,
		_w4399_,
		_w4400_
	);
	LUT4 #(
		.INIT('h1311)
	) name3938 (
		_w1731_,
		_w4386_,
		_w4389_,
		_w4400_,
		_w4401_
	);
	LUT3 #(
		.INIT('hce)
	) name3939 (
		\P1_state_reg[0]/NET0131 ,
		_w4385_,
		_w4401_,
		_w4402_
	);
	LUT2 #(
		.INIT('h2)
	) name3940 (
		\P1_reg2_reg[12]/NET0131 ,
		_w2462_,
		_w4403_
	);
	LUT4 #(
		.INIT('h2000)
	) name3941 (
		\P1_reg2_reg[12]/NET0131 ,
		_w1723_,
		_w1727_,
		_w1730_,
		_w4404_
	);
	LUT2 #(
		.INIT('h2)
	) name3942 (
		\P1_reg2_reg[12]/NET0131 ,
		_w1741_,
		_w4405_
	);
	LUT4 #(
		.INIT('he020)
	) name3943 (
		\P1_reg2_reg[12]/NET0131 ,
		_w1741_,
		_w2292_,
		_w3798_,
		_w4406_
	);
	LUT4 #(
		.INIT('h280a)
	) name3944 (
		_w1741_,
		_w2004_,
		_w2016_,
		_w3804_,
		_w4407_
	);
	LUT3 #(
		.INIT('ha8)
	) name3945 (
		_w2447_,
		_w4405_,
		_w4407_,
		_w4408_
	);
	LUT4 #(
		.INIT('hddd1)
	) name3946 (
		\P1_reg2_reg[12]/NET0131 ,
		_w1741_,
		_w3800_,
		_w3801_,
		_w4409_
	);
	LUT2 #(
		.INIT('h2)
	) name3947 (
		_w2424_,
		_w4409_,
		_w4410_
	);
	LUT4 #(
		.INIT('hd11d)
	) name3948 (
		\P1_reg2_reg[12]/NET0131 ,
		_w1741_,
		_w2807_,
		_w3173_,
		_w4411_
	);
	LUT4 #(
		.INIT('h2300)
	) name3949 (
		_w1748_,
		_w2013_,
		_w2015_,
		_w2426_,
		_w4412_
	);
	LUT2 #(
		.INIT('h8)
	) name3950 (
		_w1741_,
		_w4412_,
		_w4413_
	);
	LUT4 #(
		.INIT('haa20)
	) name3951 (
		\P1_reg2_reg[12]/NET0131 ,
		_w1741_,
		_w2426_,
		_w2450_,
		_w4414_
	);
	LUT4 #(
		.INIT('h0008)
	) name3952 (
		_w2018_,
		_w2284_,
		_w2288_,
		_w2291_,
		_w4415_
	);
	LUT3 #(
		.INIT('h01)
	) name3953 (
		_w4414_,
		_w4415_,
		_w4413_,
		_w4416_
	);
	LUT3 #(
		.INIT('hd0)
	) name3954 (
		_w2388_,
		_w4411_,
		_w4416_,
		_w4417_
	);
	LUT4 #(
		.INIT('h0100)
	) name3955 (
		_w4406_,
		_w4410_,
		_w4408_,
		_w4417_,
		_w4418_
	);
	LUT4 #(
		.INIT('ha0a8)
	) name3956 (
		\P1_state_reg[0]/NET0131 ,
		_w1731_,
		_w4404_,
		_w4418_,
		_w4419_
	);
	LUT2 #(
		.INIT('he)
	) name3957 (
		_w4403_,
		_w4419_,
		_w4420_
	);
	LUT4 #(
		.INIT('hd070)
	) name3958 (
		\P1_state_reg[0]/NET0131 ,
		\P2_IR_reg[23]/NET0131 ,
		\P2_reg0_reg[23]/NET0131 ,
		_w1188_,
		_w4421_
	);
	LUT4 #(
		.INIT('h2000)
	) name3959 (
		\P2_reg0_reg[23]/NET0131 ,
		_w1189_,
		_w1352_,
		_w1356_,
		_w4422_
	);
	LUT4 #(
		.INIT('h02aa)
	) name3960 (
		\P2_reg0_reg[23]/NET0131 ,
		_w1361_,
		_w1363_,
		_w1368_,
		_w4423_
	);
	LUT4 #(
		.INIT('h111d)
	) name3961 (
		\P2_reg0_reg[23]/NET0131 ,
		_w1369_,
		_w3583_,
		_w3584_,
		_w4424_
	);
	LUT2 #(
		.INIT('h2)
	) name3962 (
		_w1191_,
		_w4424_,
		_w4425_
	);
	LUT3 #(
		.INIT('ha2)
	) name3963 (
		\P2_reg0_reg[23]/NET0131 ,
		_w1684_,
		_w1685_,
		_w4426_
	);
	LUT4 #(
		.INIT('h1000)
	) name3964 (
		_w546_,
		_w981_,
		_w1411_,
		_w1442_,
		_w4427_
	);
	LUT2 #(
		.INIT('h1)
	) name3965 (
		_w4426_,
		_w4427_,
		_w4428_
	);
	LUT4 #(
		.INIT('h5700)
	) name3966 (
		_w1447_,
		_w3619_,
		_w4423_,
		_w4428_,
		_w4429_
	);
	LUT4 #(
		.INIT('haaa8)
	) name3967 (
		\P2_reg0_reg[23]/NET0131 ,
		_w1361_,
		_w1363_,
		_w1368_,
		_w4430_
	);
	LUT4 #(
		.INIT('hc535)
	) name3968 (
		\P2_reg0_reg[23]/NET0131 ,
		_w1278_,
		_w1411_,
		_w3601_,
		_w4431_
	);
	LUT2 #(
		.INIT('h1)
	) name3969 (
		_w1409_,
		_w4431_,
		_w4432_
	);
	LUT3 #(
		.INIT('h54)
	) name3970 (
		_w1496_,
		_w3611_,
		_w4430_,
		_w4433_
	);
	LUT4 #(
		.INIT('h0100)
	) name3971 (
		_w4425_,
		_w4432_,
		_w4433_,
		_w4429_,
		_w4434_
	);
	LUT4 #(
		.INIT('ha0a8)
	) name3972 (
		\P1_state_reg[0]/NET0131 ,
		_w1359_,
		_w4422_,
		_w4434_,
		_w4435_
	);
	LUT2 #(
		.INIT('he)
	) name3973 (
		_w4421_,
		_w4435_,
		_w4436_
	);
	LUT2 #(
		.INIT('h2)
	) name3974 (
		\P1_reg0_reg[12]/NET0131 ,
		_w2462_,
		_w4437_
	);
	LUT4 #(
		.INIT('h2000)
	) name3975 (
		\P1_reg0_reg[12]/NET0131 ,
		_w1723_,
		_w1727_,
		_w1730_,
		_w4438_
	);
	LUT4 #(
		.INIT('hc808)
	) name3976 (
		\P1_reg0_reg[12]/NET0131 ,
		_w2292_,
		_w2883_,
		_w3798_,
		_w4439_
	);
	LUT4 #(
		.INIT('hddd1)
	) name3977 (
		\P1_reg0_reg[12]/NET0131 ,
		_w2883_,
		_w3800_,
		_w3801_,
		_w4440_
	);
	LUT2 #(
		.INIT('h2)
	) name3978 (
		_w2424_,
		_w4440_,
		_w4441_
	);
	LUT3 #(
		.INIT('ha8)
	) name3979 (
		_w2883_,
		_w3805_,
		_w4412_,
		_w4442_
	);
	LUT4 #(
		.INIT('hc535)
	) name3980 (
		\P1_reg0_reg[12]/NET0131 ,
		_w2807_,
		_w2883_,
		_w3173_,
		_w4443_
	);
	LUT2 #(
		.INIT('h2)
	) name3981 (
		\P1_reg0_reg[12]/NET0131 ,
		_w3420_,
		_w4444_
	);
	LUT4 #(
		.INIT('h0031)
	) name3982 (
		_w2388_,
		_w4442_,
		_w4443_,
		_w4444_,
		_w4445_
	);
	LUT4 #(
		.INIT('ha8aa)
	) name3983 (
		_w1731_,
		_w4439_,
		_w4441_,
		_w4445_,
		_w4446_
	);
	LUT4 #(
		.INIT('heeec)
	) name3984 (
		\P1_state_reg[0]/NET0131 ,
		_w4437_,
		_w4438_,
		_w4446_,
		_w4447_
	);
	LUT4 #(
		.INIT('hd070)
	) name3985 (
		\P1_state_reg[0]/NET0131 ,
		\P2_IR_reg[23]/NET0131 ,
		\P2_reg1_reg[23]/NET0131 ,
		_w1188_,
		_w4448_
	);
	LUT4 #(
		.INIT('h2000)
	) name3986 (
		\P2_reg1_reg[23]/NET0131 ,
		_w1189_,
		_w1352_,
		_w1356_,
		_w4449_
	);
	LUT4 #(
		.INIT('h111d)
	) name3987 (
		\P2_reg1_reg[23]/NET0131 ,
		_w1507_,
		_w3583_,
		_w3584_,
		_w4450_
	);
	LUT2 #(
		.INIT('h2)
	) name3988 (
		_w1191_,
		_w4450_,
		_w4451_
	);
	LUT4 #(
		.INIT('haa02)
	) name3989 (
		\P2_reg1_reg[23]/NET0131 ,
		_w1361_,
		_w1363_,
		_w1368_,
		_w4452_
	);
	LUT4 #(
		.INIT('h4844)
	) name3990 (
		_w1278_,
		_w1516_,
		_w3589_,
		_w3591_,
		_w4453_
	);
	LUT3 #(
		.INIT('ha2)
	) name3991 (
		\P2_reg1_reg[23]/NET0131 ,
		_w1684_,
		_w2469_,
		_w4454_
	);
	LUT4 #(
		.INIT('h1000)
	) name3992 (
		_w546_,
		_w981_,
		_w1442_,
		_w1516_,
		_w4455_
	);
	LUT2 #(
		.INIT('h1)
	) name3993 (
		_w4454_,
		_w4455_,
		_w4456_
	);
	LUT4 #(
		.INIT('hab00)
	) name3994 (
		_w1575_,
		_w4452_,
		_w4453_,
		_w4456_,
		_w4457_
	);
	LUT4 #(
		.INIT('hc535)
	) name3995 (
		\P2_reg1_reg[23]/NET0131 ,
		_w1278_,
		_w1516_,
		_w3601_,
		_w4458_
	);
	LUT4 #(
		.INIT('hc535)
	) name3996 (
		\P2_reg1_reg[23]/NET0131 ,
		_w1278_,
		_w1507_,
		_w3601_,
		_w4459_
	);
	LUT4 #(
		.INIT('hfa32)
	) name3997 (
		_w1506_,
		_w1530_,
		_w4458_,
		_w4459_,
		_w4460_
	);
	LUT4 #(
		.INIT('h8aaa)
	) name3998 (
		_w1359_,
		_w4451_,
		_w4457_,
		_w4460_,
		_w4461_
	);
	LUT4 #(
		.INIT('heeec)
	) name3999 (
		\P1_state_reg[0]/NET0131 ,
		_w4448_,
		_w4449_,
		_w4461_,
		_w4462_
	);
	LUT2 #(
		.INIT('h2)
	) name4000 (
		\P1_reg0_reg[16]/NET0131 ,
		_w2462_,
		_w4463_
	);
	LUT4 #(
		.INIT('h2000)
	) name4001 (
		\P1_reg0_reg[16]/NET0131 ,
		_w1723_,
		_w1727_,
		_w1730_,
		_w4464_
	);
	LUT2 #(
		.INIT('h2)
	) name4002 (
		\P1_reg0_reg[16]/NET0131 ,
		_w2883_,
		_w4465_
	);
	LUT4 #(
		.INIT('h0c84)
	) name4003 (
		_w2768_,
		_w2883_,
		_w3168_,
		_w3817_,
		_w4466_
	);
	LUT3 #(
		.INIT('ha8)
	) name4004 (
		_w2292_,
		_w4465_,
		_w4466_,
		_w4467_
	);
	LUT4 #(
		.INIT('h08c8)
	) name4005 (
		\P1_reg0_reg[16]/NET0131 ,
		_w2388_,
		_w2883_,
		_w3820_,
		_w4468_
	);
	LUT4 #(
		.INIT('h7020)
	) name4006 (
		_w1747_,
		_w2246_,
		_w2883_,
		_w3822_,
		_w4469_
	);
	LUT2 #(
		.INIT('h2)
	) name4007 (
		\P1_reg0_reg[16]/NET0131 ,
		_w3420_,
		_w4470_
	);
	LUT4 #(
		.INIT('h0057)
	) name4008 (
		_w2883_,
		_w3824_,
		_w4393_,
		_w4470_,
		_w4471_
	);
	LUT4 #(
		.INIT('h5700)
	) name4009 (
		_w2424_,
		_w4465_,
		_w4469_,
		_w4471_,
		_w4472_
	);
	LUT2 #(
		.INIT('h4)
	) name4010 (
		_w4468_,
		_w4472_,
		_w4473_
	);
	LUT4 #(
		.INIT('h1311)
	) name4011 (
		_w1731_,
		_w4464_,
		_w4467_,
		_w4473_,
		_w4474_
	);
	LUT3 #(
		.INIT('hce)
	) name4012 (
		\P1_state_reg[0]/NET0131 ,
		_w4463_,
		_w4474_,
		_w4475_
	);
	LUT2 #(
		.INIT('h2)
	) name4013 (
		\P1_reg0_reg[20]/NET0131 ,
		_w2462_,
		_w4476_
	);
	LUT4 #(
		.INIT('h2000)
	) name4014 (
		\P1_reg0_reg[20]/NET0131 ,
		_w1723_,
		_w1727_,
		_w1730_,
		_w4477_
	);
	LUT2 #(
		.INIT('h2)
	) name4015 (
		\P1_reg0_reg[20]/NET0131 ,
		_w2883_,
		_w4478_
	);
	LUT4 #(
		.INIT('h40b0)
	) name4016 (
		_w2765_,
		_w2773_,
		_w2883_,
		_w3162_,
		_w4479_
	);
	LUT3 #(
		.INIT('ha8)
	) name4017 (
		_w2292_,
		_w4478_,
		_w4479_,
		_w4480_
	);
	LUT4 #(
		.INIT('h7020)
	) name4018 (
		_w1747_,
		_w2175_,
		_w2883_,
		_w3857_,
		_w4481_
	);
	LUT3 #(
		.INIT('ha8)
	) name4019 (
		_w2424_,
		_w4478_,
		_w4481_,
		_w4482_
	);
	LUT4 #(
		.INIT('hc535)
	) name4020 (
		\P1_reg0_reg[20]/NET0131 ,
		_w2822_,
		_w2883_,
		_w3162_,
		_w4483_
	);
	LUT4 #(
		.INIT('hcc80)
	) name4021 (
		_w2447_,
		_w2883_,
		_w3861_,
		_w4038_,
		_w4484_
	);
	LUT2 #(
		.INIT('h2)
	) name4022 (
		\P1_reg0_reg[20]/NET0131 ,
		_w3420_,
		_w4485_
	);
	LUT2 #(
		.INIT('h1)
	) name4023 (
		_w4484_,
		_w4485_,
		_w4486_
	);
	LUT3 #(
		.INIT('hd0)
	) name4024 (
		_w2388_,
		_w4483_,
		_w4486_,
		_w4487_
	);
	LUT4 #(
		.INIT('ha8aa)
	) name4025 (
		_w1731_,
		_w4482_,
		_w4480_,
		_w4487_,
		_w4488_
	);
	LUT4 #(
		.INIT('heeec)
	) name4026 (
		\P1_state_reg[0]/NET0131 ,
		_w4476_,
		_w4477_,
		_w4488_,
		_w4489_
	);
	LUT2 #(
		.INIT('h2)
	) name4027 (
		\P1_reg1_reg[12]/NET0131 ,
		_w2462_,
		_w4490_
	);
	LUT4 #(
		.INIT('h2000)
	) name4028 (
		\P1_reg1_reg[12]/NET0131 ,
		_w1723_,
		_w1727_,
		_w1730_,
		_w4491_
	);
	LUT4 #(
		.INIT('hc808)
	) name4029 (
		\P1_reg1_reg[12]/NET0131 ,
		_w2292_,
		_w2520_,
		_w3798_,
		_w4492_
	);
	LUT4 #(
		.INIT('hddd1)
	) name4030 (
		\P1_reg1_reg[12]/NET0131 ,
		_w2520_,
		_w3800_,
		_w3801_,
		_w4493_
	);
	LUT2 #(
		.INIT('h2)
	) name4031 (
		_w2424_,
		_w4493_,
		_w4494_
	);
	LUT3 #(
		.INIT('ha8)
	) name4032 (
		_w2520_,
		_w3805_,
		_w4412_,
		_w4495_
	);
	LUT4 #(
		.INIT('hd11d)
	) name4033 (
		\P1_reg1_reg[12]/NET0131 ,
		_w2520_,
		_w2807_,
		_w3173_,
		_w4496_
	);
	LUT2 #(
		.INIT('h2)
	) name4034 (
		\P1_reg1_reg[12]/NET0131 ,
		_w2525_,
		_w4497_
	);
	LUT4 #(
		.INIT('h0031)
	) name4035 (
		_w2388_,
		_w4495_,
		_w4496_,
		_w4497_,
		_w4498_
	);
	LUT4 #(
		.INIT('ha8aa)
	) name4036 (
		_w1731_,
		_w4492_,
		_w4494_,
		_w4498_,
		_w4499_
	);
	LUT4 #(
		.INIT('heeec)
	) name4037 (
		\P1_state_reg[0]/NET0131 ,
		_w4490_,
		_w4491_,
		_w4499_,
		_w4500_
	);
	LUT2 #(
		.INIT('h2)
	) name4038 (
		\P1_reg1_reg[16]/NET0131 ,
		_w2462_,
		_w4501_
	);
	LUT4 #(
		.INIT('h2000)
	) name4039 (
		\P1_reg1_reg[16]/NET0131 ,
		_w1723_,
		_w1727_,
		_w1730_,
		_w4502_
	);
	LUT2 #(
		.INIT('h2)
	) name4040 (
		\P1_reg1_reg[16]/NET0131 ,
		_w2520_,
		_w4503_
	);
	LUT4 #(
		.INIT('h0a82)
	) name4041 (
		_w2520_,
		_w2768_,
		_w3168_,
		_w3817_,
		_w4504_
	);
	LUT3 #(
		.INIT('ha8)
	) name4042 (
		_w2292_,
		_w4503_,
		_w4504_,
		_w4505_
	);
	LUT4 #(
		.INIT('h08c8)
	) name4043 (
		\P1_reg1_reg[16]/NET0131 ,
		_w2388_,
		_w2520_,
		_w3820_,
		_w4506_
	);
	LUT4 #(
		.INIT('h7020)
	) name4044 (
		_w1747_,
		_w2246_,
		_w2520_,
		_w3822_,
		_w4507_
	);
	LUT2 #(
		.INIT('h2)
	) name4045 (
		\P1_reg1_reg[16]/NET0131 ,
		_w2525_,
		_w4508_
	);
	LUT4 #(
		.INIT('h0057)
	) name4046 (
		_w2520_,
		_w3824_,
		_w4393_,
		_w4508_,
		_w4509_
	);
	LUT4 #(
		.INIT('h5700)
	) name4047 (
		_w2424_,
		_w4503_,
		_w4507_,
		_w4509_,
		_w4510_
	);
	LUT2 #(
		.INIT('h4)
	) name4048 (
		_w4506_,
		_w4510_,
		_w4511_
	);
	LUT4 #(
		.INIT('h1311)
	) name4049 (
		_w1731_,
		_w4502_,
		_w4505_,
		_w4511_,
		_w4512_
	);
	LUT3 #(
		.INIT('hce)
	) name4050 (
		\P1_state_reg[0]/NET0131 ,
		_w4501_,
		_w4512_,
		_w4513_
	);
	LUT2 #(
		.INIT('h2)
	) name4051 (
		\P1_reg1_reg[20]/NET0131 ,
		_w2462_,
		_w4514_
	);
	LUT4 #(
		.INIT('h2000)
	) name4052 (
		\P1_reg1_reg[20]/NET0131 ,
		_w1723_,
		_w1727_,
		_w1730_,
		_w4515_
	);
	LUT2 #(
		.INIT('h2)
	) name4053 (
		\P1_reg1_reg[20]/NET0131 ,
		_w2520_,
		_w4516_
	);
	LUT4 #(
		.INIT('h208a)
	) name4054 (
		_w2520_,
		_w2765_,
		_w2773_,
		_w3162_,
		_w4517_
	);
	LUT3 #(
		.INIT('ha8)
	) name4055 (
		_w2292_,
		_w4516_,
		_w4517_,
		_w4518_
	);
	LUT4 #(
		.INIT('h7020)
	) name4056 (
		_w1747_,
		_w2175_,
		_w2520_,
		_w3857_,
		_w4519_
	);
	LUT3 #(
		.INIT('ha8)
	) name4057 (
		_w2424_,
		_w4516_,
		_w4519_,
		_w4520_
	);
	LUT4 #(
		.INIT('hd11d)
	) name4058 (
		\P1_reg1_reg[20]/NET0131 ,
		_w2520_,
		_w2822_,
		_w3162_,
		_w4521_
	);
	LUT4 #(
		.INIT('hc808)
	) name4059 (
		\P1_reg1_reg[20]/NET0131 ,
		_w2447_,
		_w2520_,
		_w3861_,
		_w4522_
	);
	LUT4 #(
		.INIT('h1000)
	) name4060 (
		_w1748_,
		_w2154_,
		_w2426_,
		_w2520_,
		_w4523_
	);
	LUT4 #(
		.INIT('h08aa)
	) name4061 (
		\P1_reg1_reg[20]/NET0131 ,
		_w2426_,
		_w2520_,
		_w2524_,
		_w4524_
	);
	LUT2 #(
		.INIT('h1)
	) name4062 (
		_w4523_,
		_w4524_,
		_w4525_
	);
	LUT2 #(
		.INIT('h4)
	) name4063 (
		_w4522_,
		_w4525_,
		_w4526_
	);
	LUT3 #(
		.INIT('hd0)
	) name4064 (
		_w2388_,
		_w4521_,
		_w4526_,
		_w4527_
	);
	LUT4 #(
		.INIT('ha8aa)
	) name4065 (
		_w1731_,
		_w4520_,
		_w4518_,
		_w4527_,
		_w4528_
	);
	LUT4 #(
		.INIT('heeec)
	) name4066 (
		\P1_state_reg[0]/NET0131 ,
		_w4514_,
		_w4515_,
		_w4528_,
		_w4529_
	);
	LUT4 #(
		.INIT('h4000)
	) name4067 (
		_w1723_,
		_w1727_,
		_w1730_,
		_w2005_,
		_w4530_
	);
	LUT2 #(
		.INIT('h2)
	) name4068 (
		_w2005_,
		_w2644_,
		_w4531_
	);
	LUT4 #(
		.INIT('h8a20)
	) name4069 (
		_w2644_,
		_w2654_,
		_w2655_,
		_w3191_,
		_w4532_
	);
	LUT3 #(
		.INIT('ha8)
	) name4070 (
		_w2292_,
		_w4531_,
		_w4532_,
		_w4533_
	);
	LUT4 #(
		.INIT('h208a)
	) name4071 (
		_w2644_,
		_w2667_,
		_w2668_,
		_w3191_,
		_w4534_
	);
	LUT3 #(
		.INIT('ha8)
	) name4072 (
		_w2388_,
		_w4531_,
		_w4534_,
		_w4535_
	);
	LUT4 #(
		.INIT('h1444)
	) name4073 (
		_w1747_,
		_w2020_,
		_w2404_,
		_w2405_,
		_w4536_
	);
	LUT3 #(
		.INIT('h80)
	) name4074 (
		_w1747_,
		_w2030_,
		_w2033_,
		_w4537_
	);
	LUT4 #(
		.INIT('h3331)
	) name4075 (
		_w2644_,
		_w4531_,
		_w4536_,
		_w4537_,
		_w4538_
	);
	LUT4 #(
		.INIT('h8040)
	) name4076 (
		_w2004_,
		_w2447_,
		_w2644_,
		_w3804_,
		_w4539_
	);
	LUT4 #(
		.INIT('ha8a0)
	) name4077 (
		_w2004_,
		_w2426_,
		_w2454_,
		_w2644_,
		_w4540_
	);
	LUT3 #(
		.INIT('h0d)
	) name4078 (
		_w2005_,
		_w2690_,
		_w4540_,
		_w4541_
	);
	LUT2 #(
		.INIT('h4)
	) name4079 (
		_w4539_,
		_w4541_,
		_w4542_
	);
	LUT3 #(
		.INIT('hd0)
	) name4080 (
		_w2424_,
		_w4538_,
		_w4542_,
		_w4543_
	);
	LUT4 #(
		.INIT('ha8aa)
	) name4081 (
		_w1731_,
		_w4533_,
		_w4535_,
		_w4543_,
		_w4544_
	);
	LUT2 #(
		.INIT('h2)
	) name4082 (
		\P1_reg3_reg[11]/NET0131 ,
		\P1_state_reg[0]/NET0131 ,
		_w4545_
	);
	LUT3 #(
		.INIT('h07)
	) name4083 (
		_w2005_,
		_w2695_,
		_w4545_,
		_w4546_
	);
	LUT4 #(
		.INIT('ha8ff)
	) name4084 (
		\P1_state_reg[0]/NET0131 ,
		_w4530_,
		_w4544_,
		_w4546_,
		_w4547_
	);
	LUT2 #(
		.INIT('h2)
	) name4085 (
		_w2243_,
		_w2644_,
		_w4548_
	);
	LUT4 #(
		.INIT('h007d)
	) name4086 (
		_w2644_,
		_w3169_,
		_w4358_,
		_w4548_,
		_w4549_
	);
	LUT2 #(
		.INIT('h2)
	) name4087 (
		_w2292_,
		_w4549_,
		_w4550_
	);
	LUT4 #(
		.INIT('h00d7)
	) name4088 (
		_w2644_,
		_w3169_,
		_w4364_,
		_w4548_,
		_w4551_
	);
	LUT4 #(
		.INIT('h1444)
	) name4089 (
		_w1747_,
		_w2235_,
		_w2404_,
		_w2408_,
		_w4552_
	);
	LUT3 #(
		.INIT('h80)
	) name4090 (
		_w1747_,
		_w2210_,
		_w2211_,
		_w4553_
	);
	LUT4 #(
		.INIT('h3331)
	) name4091 (
		_w2644_,
		_w4548_,
		_w4552_,
		_w4553_,
		_w4554_
	);
	LUT4 #(
		.INIT('ha8d8)
	) name4092 (
		_w2242_,
		_w2426_,
		_w2447_,
		_w3494_,
		_w4555_
	);
	LUT2 #(
		.INIT('h8)
	) name4093 (
		_w2242_,
		_w2454_,
		_w4556_
	);
	LUT4 #(
		.INIT('h88a8)
	) name4094 (
		_w2243_,
		_w2450_,
		_w2452_,
		_w2644_,
		_w4557_
	);
	LUT2 #(
		.INIT('h1)
	) name4095 (
		_w4556_,
		_w4557_,
		_w4558_
	);
	LUT3 #(
		.INIT('h70)
	) name4096 (
		_w2644_,
		_w4555_,
		_w4558_,
		_w4559_
	);
	LUT3 #(
		.INIT('hd0)
	) name4097 (
		_w2424_,
		_w4554_,
		_w4559_,
		_w4560_
	);
	LUT3 #(
		.INIT('hd0)
	) name4098 (
		_w2388_,
		_w4551_,
		_w4560_,
		_w4561_
	);
	LUT4 #(
		.INIT('h4000)
	) name4099 (
		_w1723_,
		_w1727_,
		_w1730_,
		_w2243_,
		_w4562_
	);
	LUT4 #(
		.INIT('h0075)
	) name4100 (
		_w1731_,
		_w4550_,
		_w4561_,
		_w4562_,
		_w4563_
	);
	LUT2 #(
		.INIT('h2)
	) name4101 (
		\P1_reg3_reg[15]/NET0131 ,
		\P1_state_reg[0]/NET0131 ,
		_w4564_
	);
	LUT3 #(
		.INIT('h07)
	) name4102 (
		_w2243_,
		_w2695_,
		_w4564_,
		_w4565_
	);
	LUT3 #(
		.INIT('h2f)
	) name4103 (
		\P1_state_reg[0]/NET0131 ,
		_w4563_,
		_w4565_,
		_w4566_
	);
	LUT4 #(
		.INIT('h4000)
	) name4104 (
		_w1723_,
		_w1727_,
		_w1730_,
		_w2209_,
		_w4567_
	);
	LUT2 #(
		.INIT('h2)
	) name4105 (
		_w2209_,
		_w2644_,
		_w4568_
	);
	LUT4 #(
		.INIT('h5054)
	) name4106 (
		_w1747_,
		_w2246_,
		_w2409_,
		_w2919_,
		_w4569_
	);
	LUT3 #(
		.INIT('h80)
	) name4107 (
		_w1747_,
		_w2221_,
		_w2222_,
		_w4570_
	);
	LUT4 #(
		.INIT('h3331)
	) name4108 (
		_w2644_,
		_w4568_,
		_w4569_,
		_w4570_,
		_w4571_
	);
	LUT2 #(
		.INIT('h2)
	) name4109 (
		_w2424_,
		_w4571_,
		_w4572_
	);
	LUT4 #(
		.INIT('hb04f)
	) name4110 (
		_w2935_,
		_w2936_,
		_w2937_,
		_w3174_,
		_w4573_
	);
	LUT4 #(
		.INIT('h08c8)
	) name4111 (
		_w2209_,
		_w2388_,
		_w2644_,
		_w4573_,
		_w4574_
	);
	LUT4 #(
		.INIT('hb04f)
	) name4112 (
		_w2953_,
		_w2954_,
		_w2955_,
		_w3174_,
		_w4575_
	);
	LUT4 #(
		.INIT('hc808)
	) name4113 (
		_w2209_,
		_w2292_,
		_w2644_,
		_w4575_,
		_w4576_
	);
	LUT4 #(
		.INIT('h2300)
	) name4114 (
		_w1748_,
		_w2206_,
		_w2207_,
		_w2426_,
		_w4577_
	);
	LUT4 #(
		.INIT('h2aaa)
	) name4115 (
		_w2208_,
		_w2431_,
		_w2432_,
		_w2434_,
		_w4578_
	);
	LUT4 #(
		.INIT('h0f0d)
	) name4116 (
		_w2447_,
		_w3494_,
		_w4577_,
		_w4578_,
		_w4579_
	);
	LUT4 #(
		.INIT('h2300)
	) name4117 (
		_w1748_,
		_w2206_,
		_w2207_,
		_w2454_,
		_w4580_
	);
	LUT4 #(
		.INIT('h88a8)
	) name4118 (
		_w2209_,
		_w2450_,
		_w2452_,
		_w2644_,
		_w4581_
	);
	LUT2 #(
		.INIT('h1)
	) name4119 (
		_w4580_,
		_w4581_,
		_w4582_
	);
	LUT3 #(
		.INIT('hd0)
	) name4120 (
		_w2644_,
		_w4579_,
		_w4582_,
		_w4583_
	);
	LUT3 #(
		.INIT('h10)
	) name4121 (
		_w4576_,
		_w4574_,
		_w4583_,
		_w4584_
	);
	LUT4 #(
		.INIT('h1311)
	) name4122 (
		_w1731_,
		_w4567_,
		_w4572_,
		_w4584_,
		_w4585_
	);
	LUT2 #(
		.INIT('h2)
	) name4123 (
		\P1_reg3_reg[14]/NET0131 ,
		\P1_state_reg[0]/NET0131 ,
		_w4586_
	);
	LUT3 #(
		.INIT('h07)
	) name4124 (
		_w2209_,
		_w2695_,
		_w4586_,
		_w4587_
	);
	LUT3 #(
		.INIT('h2f)
	) name4125 (
		\P1_state_reg[0]/NET0131 ,
		_w4585_,
		_w4587_,
		_w4588_
	);
	LUT4 #(
		.INIT('h1000)
	) name4126 (
		_w674_,
		_w1189_,
		_w1352_,
		_w1356_,
		_w4589_
	);
	LUT4 #(
		.INIT('h0155)
	) name4127 (
		_w674_,
		_w1361_,
		_w1363_,
		_w1368_,
		_w4590_
	);
	LUT4 #(
		.INIT('h8488)
	) name4128 (
		_w1320_,
		_w1369_,
		_w1379_,
		_w1383_,
		_w4591_
	);
	LUT3 #(
		.INIT('h04)
	) name4129 (
		_w685_,
		_w1232_,
		_w1439_,
		_w4592_
	);
	LUT3 #(
		.INIT('h54)
	) name4130 (
		_w674_,
		_w1441_,
		_w1443_,
		_w4593_
	);
	LUT2 #(
		.INIT('h1)
	) name4131 (
		_w4592_,
		_w4593_,
		_w4594_
	);
	LUT4 #(
		.INIT('hab00)
	) name4132 (
		_w1409_,
		_w4590_,
		_w4591_,
		_w4594_,
		_w4595_
	);
	LUT2 #(
		.INIT('h1)
	) name4133 (
		_w693_,
		_w1435_,
		_w4596_
	);
	LUT3 #(
		.INIT('h70)
	) name4134 (
		_w1418_,
		_w1419_,
		_w1435_,
		_w4597_
	);
	LUT4 #(
		.INIT('h020f)
	) name4135 (
		_w653_,
		_w4256_,
		_w4596_,
		_w4597_,
		_w4598_
	);
	LUT4 #(
		.INIT('h04c4)
	) name4136 (
		_w674_,
		_w1191_,
		_w1411_,
		_w4598_,
		_w4599_
	);
	LUT4 #(
		.INIT('h9a55)
	) name4137 (
		_w1320_,
		_w1458_,
		_w1461_,
		_w1466_,
		_w4600_
	);
	LUT4 #(
		.INIT('h0d01)
	) name4138 (
		_w674_,
		_w1369_,
		_w1496_,
		_w4600_,
		_w4601_
	);
	LUT4 #(
		.INIT('hc404)
	) name4139 (
		_w674_,
		_w1447_,
		_w1411_,
		_w4600_,
		_w4602_
	);
	LUT4 #(
		.INIT('h0100)
	) name4140 (
		_w4601_,
		_w4602_,
		_w4599_,
		_w4595_,
		_w4603_
	);
	LUT4 #(
		.INIT('ha0a8)
	) name4141 (
		\P1_state_reg[0]/NET0131 ,
		_w1359_,
		_w4589_,
		_w4603_,
		_w4604_
	);
	LUT2 #(
		.INIT('h4)
	) name4142 (
		\P1_state_reg[0]/NET0131 ,
		\P2_reg3_reg[11]/NET0131 ,
		_w4605_
	);
	LUT4 #(
		.INIT('h0802)
	) name4143 (
		\P1_state_reg[0]/NET0131 ,
		\P2_IR_reg[23]/NET0131 ,
		_w674_,
		_w1188_,
		_w4606_
	);
	LUT2 #(
		.INIT('h1)
	) name4144 (
		_w4605_,
		_w4606_,
		_w4607_
	);
	LUT2 #(
		.INIT('hb)
	) name4145 (
		_w4604_,
		_w4607_,
		_w4608_
	);
	LUT4 #(
		.INIT('h1000)
	) name4146 (
		_w620_,
		_w1189_,
		_w1352_,
		_w1356_,
		_w4609_
	);
	LUT4 #(
		.INIT('h5554)
	) name4147 (
		_w620_,
		_w1361_,
		_w1363_,
		_w1368_,
		_w4610_
	);
	LUT4 #(
		.INIT('h00b7)
	) name4148 (
		_w1296_,
		_w1411_,
		_w2540_,
		_w4610_,
		_w4611_
	);
	LUT2 #(
		.INIT('h2)
	) name4149 (
		_w1447_,
		_w4611_,
		_w4612_
	);
	LUT4 #(
		.INIT('h4000)
	) name4150 (
		_w631_,
		_w1418_,
		_w1419_,
		_w1421_,
		_w4613_
	);
	LUT4 #(
		.INIT('h00c4)
	) name4151 (
		_w528_,
		_w1435_,
		_w4299_,
		_w4613_,
		_w4614_
	);
	LUT2 #(
		.INIT('h1)
	) name4152 (
		_w631_,
		_w1435_,
		_w4615_
	);
	LUT4 #(
		.INIT('h1113)
	) name4153 (
		_w1411_,
		_w4610_,
		_w4614_,
		_w4615_,
		_w4616_
	);
	LUT3 #(
		.INIT('h04)
	) name4154 (
		_w615_,
		_w1232_,
		_w1439_,
		_w4617_
	);
	LUT3 #(
		.INIT('h54)
	) name4155 (
		_w620_,
		_w1441_,
		_w1443_,
		_w4618_
	);
	LUT2 #(
		.INIT('h1)
	) name4156 (
		_w4617_,
		_w4618_,
		_w4619_
	);
	LUT3 #(
		.INIT('hd0)
	) name4157 (
		_w1191_,
		_w4616_,
		_w4619_,
		_w4620_
	);
	LUT4 #(
		.INIT('h0155)
	) name4158 (
		_w620_,
		_w1361_,
		_w1363_,
		_w1368_,
		_w4621_
	);
	LUT4 #(
		.INIT('h00b7)
	) name4159 (
		_w1296_,
		_w1369_,
		_w2540_,
		_w4621_,
		_w4622_
	);
	LUT4 #(
		.INIT('h007b)
	) name4160 (
		_w1296_,
		_w1369_,
		_w2557_,
		_w4621_,
		_w4623_
	);
	LUT4 #(
		.INIT('hfca8)
	) name4161 (
		_w1409_,
		_w1496_,
		_w4622_,
		_w4623_,
		_w4624_
	);
	LUT4 #(
		.INIT('h8aaa)
	) name4162 (
		_w1359_,
		_w4612_,
		_w4620_,
		_w4624_,
		_w4625_
	);
	LUT2 #(
		.INIT('h4)
	) name4163 (
		\P1_state_reg[0]/NET0131 ,
		\P2_reg3_reg[14]/NET0131 ,
		_w4626_
	);
	LUT3 #(
		.INIT('h0b)
	) name4164 (
		_w620_,
		_w1349_,
		_w4626_,
		_w4627_
	);
	LUT4 #(
		.INIT('ha8ff)
	) name4165 (
		\P1_state_reg[0]/NET0131 ,
		_w4609_,
		_w4625_,
		_w4627_,
		_w4628_
	);
	LUT4 #(
		.INIT('h1000)
	) name4166 (
		_w525_,
		_w1189_,
		_w1352_,
		_w1356_,
		_w4629_
	);
	LUT4 #(
		.INIT('h5554)
	) name4167 (
		_w525_,
		_w1361_,
		_w1363_,
		_w1368_,
		_w4630_
	);
	LUT4 #(
		.INIT('h4844)
	) name4168 (
		_w1295_,
		_w1411_,
		_w1471_,
		_w1475_,
		_w4631_
	);
	LUT3 #(
		.INIT('ha8)
	) name4169 (
		_w1447_,
		_w4630_,
		_w4631_,
		_w4632_
	);
	LUT3 #(
		.INIT('h07)
	) name4170 (
		_w618_,
		_w622_,
		_w1435_,
		_w4633_
	);
	LUT4 #(
		.INIT('h3010)
	) name4171 (
		_w866_,
		_w1423_,
		_w1435_,
		_w4613_,
		_w4634_
	);
	LUT4 #(
		.INIT('h1113)
	) name4172 (
		_w1411_,
		_w4630_,
		_w4633_,
		_w4634_,
		_w4635_
	);
	LUT3 #(
		.INIT('h04)
	) name4173 (
		_w594_,
		_w1232_,
		_w1439_,
		_w4636_
	);
	LUT3 #(
		.INIT('h54)
	) name4174 (
		_w525_,
		_w1441_,
		_w1443_,
		_w4637_
	);
	LUT2 #(
		.INIT('h1)
	) name4175 (
		_w4636_,
		_w4637_,
		_w4638_
	);
	LUT3 #(
		.INIT('hd0)
	) name4176 (
		_w1191_,
		_w4635_,
		_w4638_,
		_w4639_
	);
	LUT4 #(
		.INIT('h0155)
	) name4177 (
		_w525_,
		_w1361_,
		_w1363_,
		_w1368_,
		_w4640_
	);
	LUT4 #(
		.INIT('h4844)
	) name4178 (
		_w1295_,
		_w1369_,
		_w1471_,
		_w1475_,
		_w4641_
	);
	LUT3 #(
		.INIT('h54)
	) name4179 (
		_w1496_,
		_w4640_,
		_w4641_,
		_w4642_
	);
	LUT4 #(
		.INIT('h00b7)
	) name4180 (
		_w1295_,
		_w1369_,
		_w3598_,
		_w4640_,
		_w4643_
	);
	LUT2 #(
		.INIT('h1)
	) name4181 (
		_w1409_,
		_w4643_,
		_w4644_
	);
	LUT4 #(
		.INIT('h0100)
	) name4182 (
		_w4632_,
		_w4642_,
		_w4644_,
		_w4639_,
		_w4645_
	);
	LUT4 #(
		.INIT('ha0a8)
	) name4183 (
		\P1_state_reg[0]/NET0131 ,
		_w1359_,
		_w4629_,
		_w4645_,
		_w4646_
	);
	LUT4 #(
		.INIT('h0802)
	) name4184 (
		\P1_state_reg[0]/NET0131 ,
		\P2_IR_reg[23]/NET0131 ,
		_w525_,
		_w1188_,
		_w4647_
	);
	LUT2 #(
		.INIT('h4)
	) name4185 (
		\P1_state_reg[0]/NET0131 ,
		\P2_reg3_reg[15]/NET0131 ,
		_w4648_
	);
	LUT2 #(
		.INIT('h1)
	) name4186 (
		_w4647_,
		_w4648_,
		_w4649_
	);
	LUT2 #(
		.INIT('hb)
	) name4187 (
		_w4646_,
		_w4649_,
		_w4650_
	);
	LUT4 #(
		.INIT('h4000)
	) name4188 (
		_w1723_,
		_w1727_,
		_w1730_,
		_w2106_,
		_w4651_
	);
	LUT3 #(
		.INIT('h2a)
	) name4189 (
		_w1747_,
		_w2116_,
		_w2117_,
		_w4652_
	);
	LUT4 #(
		.INIT('h0100)
	) name4190 (
		_w2053_,
		_w2128_,
		_w2138_,
		_w2400_,
		_w4653_
	);
	LUT4 #(
		.INIT('ha8aa)
	) name4191 (
		_w2044_,
		_w2108_,
		_w2118_,
		_w4653_,
		_w4654_
	);
	LUT2 #(
		.INIT('h1)
	) name4192 (
		_w1747_,
		_w2404_,
		_w4655_
	);
	LUT4 #(
		.INIT('h8a88)
	) name4193 (
		_w2424_,
		_w4652_,
		_w4654_,
		_w4655_,
		_w4656_
	);
	LUT4 #(
		.INIT('h8a20)
	) name4194 (
		_w2388_,
		_w2796_,
		_w2799_,
		_w3175_,
		_w4657_
	);
	LUT4 #(
		.INIT('h007d)
	) name4195 (
		_w2292_,
		_w2752_,
		_w3175_,
		_w4657_,
		_w4658_
	);
	LUT3 #(
		.INIT('h90)
	) name4196 (
		_w2104_,
		_w2431_,
		_w2447_,
		_w4659_
	);
	LUT4 #(
		.INIT('haaa2)
	) name4197 (
		_w2644_,
		_w4658_,
		_w4656_,
		_w4659_,
		_w4660_
	);
	LUT4 #(
		.INIT('ha8a0)
	) name4198 (
		_w2104_,
		_w2426_,
		_w2454_,
		_w2644_,
		_w4661_
	);
	LUT2 #(
		.INIT('h1)
	) name4199 (
		_w2644_,
		_w3574_,
		_w4662_
	);
	LUT4 #(
		.INIT('h050d)
	) name4200 (
		_w2106_,
		_w2690_,
		_w4661_,
		_w4662_,
		_w4663_
	);
	LUT4 #(
		.INIT('h1311)
	) name4201 (
		_w1731_,
		_w4651_,
		_w4660_,
		_w4663_,
		_w4664_
	);
	LUT2 #(
		.INIT('h2)
	) name4202 (
		\P1_reg3_reg[8]/NET0131 ,
		\P1_state_reg[0]/NET0131 ,
		_w4665_
	);
	LUT3 #(
		.INIT('h07)
	) name4203 (
		_w2106_,
		_w2695_,
		_w4665_,
		_w4666_
	);
	LUT3 #(
		.INIT('h2f)
	) name4204 (
		\P1_state_reg[0]/NET0131 ,
		_w4664_,
		_w4666_,
		_w4667_
	);
	LUT4 #(
		.INIT('h1000)
	) name4205 (
		_w723_,
		_w1189_,
		_w1352_,
		_w1356_,
		_w4668_
	);
	LUT4 #(
		.INIT('h5554)
	) name4206 (
		_w723_,
		_w1361_,
		_w1363_,
		_w1368_,
		_w4669_
	);
	LUT4 #(
		.INIT('h007b)
	) name4207 (
		_w1310_,
		_w1411_,
		_w1537_,
		_w4669_,
		_w4670_
	);
	LUT2 #(
		.INIT('h1)
	) name4208 (
		_w759_,
		_w1435_,
		_w4671_
	);
	LUT4 #(
		.INIT('h006f)
	) name4209 (
		_w711_,
		_w1418_,
		_w1435_,
		_w4671_,
		_w4672_
	);
	LUT4 #(
		.INIT('h04c4)
	) name4210 (
		_w723_,
		_w1191_,
		_w1411_,
		_w4672_,
		_w4673_
	);
	LUT3 #(
		.INIT('h04)
	) name4211 (
		_w731_,
		_w1232_,
		_w1439_,
		_w4674_
	);
	LUT3 #(
		.INIT('h54)
	) name4212 (
		_w723_,
		_w1441_,
		_w1443_,
		_w4675_
	);
	LUT2 #(
		.INIT('h1)
	) name4213 (
		_w4674_,
		_w4675_,
		_w4676_
	);
	LUT4 #(
		.INIT('h0d00)
	) name4214 (
		_w1447_,
		_w4670_,
		_w4673_,
		_w4676_,
		_w4677_
	);
	LUT4 #(
		.INIT('h0155)
	) name4215 (
		_w723_,
		_w1361_,
		_w1363_,
		_w1368_,
		_w4678_
	);
	LUT4 #(
		.INIT('h007b)
	) name4216 (
		_w1310_,
		_w1369_,
		_w1537_,
		_w4678_,
		_w4679_
	);
	LUT4 #(
		.INIT('h009f)
	) name4217 (
		_w1215_,
		_w1310_,
		_w1369_,
		_w4678_,
		_w4680_
	);
	LUT4 #(
		.INIT('hfca8)
	) name4218 (
		_w1409_,
		_w1496_,
		_w4679_,
		_w4680_,
		_w4681_
	);
	LUT4 #(
		.INIT('h3111)
	) name4219 (
		_w1359_,
		_w4668_,
		_w4677_,
		_w4681_,
		_w4682_
	);
	LUT2 #(
		.INIT('h4)
	) name4220 (
		\P1_state_reg[0]/NET0131 ,
		\P2_reg3_reg[8]/NET0131 ,
		_w4683_
	);
	LUT4 #(
		.INIT('h0802)
	) name4221 (
		\P1_state_reg[0]/NET0131 ,
		\P2_IR_reg[23]/NET0131 ,
		_w723_,
		_w1188_,
		_w4684_
	);
	LUT2 #(
		.INIT('h1)
	) name4222 (
		_w4683_,
		_w4684_,
		_w4685_
	);
	LUT3 #(
		.INIT('h2f)
	) name4223 (
		\P1_state_reg[0]/NET0131 ,
		_w4682_,
		_w4685_,
		_w4686_
	);
	LUT2 #(
		.INIT('h2)
	) name4224 (
		\P1_reg2_reg[10]/NET0131 ,
		_w2462_,
		_w4687_
	);
	LUT4 #(
		.INIT('h2000)
	) name4225 (
		\P1_reg2_reg[10]/NET0131 ,
		_w1723_,
		_w1727_,
		_w1730_,
		_w4688_
	);
	LUT4 #(
		.INIT('hddd1)
	) name4226 (
		\P1_reg2_reg[10]/NET0131 ,
		_w1741_,
		_w4217_,
		_w4218_,
		_w4689_
	);
	LUT2 #(
		.INIT('h2)
	) name4227 (
		_w2424_,
		_w4689_,
		_w4690_
	);
	LUT4 #(
		.INIT('hd11d)
	) name4228 (
		\P1_reg2_reg[10]/NET0131 ,
		_w1741_,
		_w2935_,
		_w3176_,
		_w4691_
	);
	LUT2 #(
		.INIT('h2)
	) name4229 (
		_w2388_,
		_w4691_,
		_w4692_
	);
	LUT4 #(
		.INIT('h1dd1)
	) name4230 (
		\P1_reg2_reg[10]/NET0131 ,
		_w1741_,
		_w2953_,
		_w3176_,
		_w4693_
	);
	LUT4 #(
		.INIT('he020)
	) name4231 (
		\P1_reg2_reg[10]/NET0131 ,
		_w1741_,
		_w2447_,
		_w4224_,
		_w4694_
	);
	LUT4 #(
		.INIT('haa20)
	) name4232 (
		\P1_reg2_reg[10]/NET0131 ,
		_w1741_,
		_w2426_,
		_w2450_,
		_w4695_
	);
	LUT4 #(
		.INIT('h0008)
	) name4233 (
		_w2032_,
		_w2284_,
		_w2288_,
		_w2291_,
		_w4696_
	);
	LUT3 #(
		.INIT('h10)
	) name4234 (
		_w2024_,
		_w2028_,
		_w2426_,
		_w4697_
	);
	LUT3 #(
		.INIT('h13)
	) name4235 (
		_w1741_,
		_w4696_,
		_w4697_,
		_w4698_
	);
	LUT2 #(
		.INIT('h4)
	) name4236 (
		_w4695_,
		_w4698_,
		_w4699_
	);
	LUT2 #(
		.INIT('h4)
	) name4237 (
		_w4694_,
		_w4699_,
		_w4700_
	);
	LUT3 #(
		.INIT('hd0)
	) name4238 (
		_w2292_,
		_w4693_,
		_w4700_,
		_w4701_
	);
	LUT4 #(
		.INIT('ha8aa)
	) name4239 (
		_w1731_,
		_w4690_,
		_w4692_,
		_w4701_,
		_w4702_
	);
	LUT4 #(
		.INIT('heeec)
	) name4240 (
		\P1_state_reg[0]/NET0131 ,
		_w4687_,
		_w4688_,
		_w4702_,
		_w4703_
	);
	LUT2 #(
		.INIT('h2)
	) name4241 (
		\P1_reg2_reg[13]/NET0131 ,
		_w2462_,
		_w4704_
	);
	LUT4 #(
		.INIT('h2000)
	) name4242 (
		\P1_reg2_reg[13]/NET0131 ,
		_w1723_,
		_w1727_,
		_w1730_,
		_w4705_
	);
	LUT2 #(
		.INIT('h2)
	) name4243 (
		\P1_reg2_reg[13]/NET0131 ,
		_w1741_,
		_w4706_
	);
	LUT4 #(
		.INIT('h20e0)
	) name4244 (
		\P1_reg2_reg[13]/NET0131 ,
		_w1741_,
		_w2388_,
		_w4245_,
		_w4707_
	);
	LUT4 #(
		.INIT('h2300)
	) name4245 (
		_w1748_,
		_w2217_,
		_w2218_,
		_w2426_,
		_w4708_
	);
	LUT4 #(
		.INIT('h0008)
	) name4246 (
		_w2220_,
		_w2284_,
		_w2288_,
		_w2291_,
		_w4709_
	);
	LUT3 #(
		.INIT('h0d)
	) name4247 (
		\P1_reg2_reg[13]/NET0131 ,
		_w4040_,
		_w4709_,
		_w4710_
	);
	LUT4 #(
		.INIT('h5700)
	) name4248 (
		_w1741_,
		_w4240_,
		_w4708_,
		_w4710_,
		_w4711_
	);
	LUT4 #(
		.INIT('h08a2)
	) name4249 (
		_w1741_,
		_w2049_,
		_w2153_,
		_w3192_,
		_w4712_
	);
	LUT3 #(
		.INIT('ha8)
	) name4250 (
		_w2292_,
		_w4706_,
		_w4712_,
		_w4713_
	);
	LUT4 #(
		.INIT('h2a08)
	) name4251 (
		_w1741_,
		_w1747_,
		_w2020_,
		_w4237_,
		_w4714_
	);
	LUT3 #(
		.INIT('ha8)
	) name4252 (
		_w2424_,
		_w4706_,
		_w4714_,
		_w4715_
	);
	LUT4 #(
		.INIT('h0100)
	) name4253 (
		_w4707_,
		_w4713_,
		_w4715_,
		_w4711_,
		_w4716_
	);
	LUT4 #(
		.INIT('ha0a8)
	) name4254 (
		\P1_state_reg[0]/NET0131 ,
		_w1731_,
		_w4705_,
		_w4716_,
		_w4717_
	);
	LUT2 #(
		.INIT('he)
	) name4255 (
		_w4704_,
		_w4717_,
		_w4718_
	);
	LUT2 #(
		.INIT('h2)
	) name4256 (
		\P1_reg2_reg[9]/NET0131 ,
		_w2462_,
		_w4719_
	);
	LUT4 #(
		.INIT('h2000)
	) name4257 (
		\P1_reg2_reg[9]/NET0131 ,
		_w1723_,
		_w1727_,
		_w1730_,
		_w4720_
	);
	LUT2 #(
		.INIT('h2)
	) name4258 (
		\P1_reg2_reg[9]/NET0131 ,
		_w1741_,
		_w4721_
	);
	LUT4 #(
		.INIT('h20e0)
	) name4259 (
		\P1_reg2_reg[9]/NET0131 ,
		_w1741_,
		_w2292_,
		_w4326_,
		_w4722_
	);
	LUT4 #(
		.INIT('h2822)
	) name4260 (
		_w1741_,
		_w2040_,
		_w2104_,
		_w2431_,
		_w4723_
	);
	LUT4 #(
		.INIT('haa20)
	) name4261 (
		\P1_reg2_reg[9]/NET0131 ,
		_w1741_,
		_w2426_,
		_w2450_,
		_w4724_
	);
	LUT4 #(
		.INIT('h0008)
	) name4262 (
		_w2042_,
		_w2284_,
		_w2288_,
		_w2291_,
		_w4725_
	);
	LUT2 #(
		.INIT('h8)
	) name4263 (
		_w2040_,
		_w2426_,
		_w4726_
	);
	LUT3 #(
		.INIT('h13)
	) name4264 (
		_w1741_,
		_w4725_,
		_w4726_,
		_w4727_
	);
	LUT2 #(
		.INIT('h4)
	) name4265 (
		_w4724_,
		_w4727_,
		_w4728_
	);
	LUT4 #(
		.INIT('h5700)
	) name4266 (
		_w2447_,
		_w4721_,
		_w4723_,
		_w4728_,
		_w4729_
	);
	LUT2 #(
		.INIT('h4)
	) name4267 (
		_w4722_,
		_w4729_,
		_w4730_
	);
	LUT4 #(
		.INIT('he020)
	) name4268 (
		\P1_reg2_reg[9]/NET0131 ,
		_w1741_,
		_w2424_,
		_w4329_,
		_w4731_
	);
	LUT4 #(
		.INIT('h1dd1)
	) name4269 (
		\P1_reg2_reg[9]/NET0131 ,
		_w1741_,
		_w2327_,
		_w3186_,
		_w4732_
	);
	LUT3 #(
		.INIT('h31)
	) name4270 (
		_w2388_,
		_w4731_,
		_w4732_,
		_w4733_
	);
	LUT4 #(
		.INIT('h3111)
	) name4271 (
		_w1731_,
		_w4720_,
		_w4730_,
		_w4733_,
		_w4734_
	);
	LUT3 #(
		.INIT('hce)
	) name4272 (
		\P1_state_reg[0]/NET0131 ,
		_w4719_,
		_w4734_,
		_w4735_
	);
	LUT4 #(
		.INIT('hd070)
	) name4273 (
		\P1_state_reg[0]/NET0131 ,
		\P2_IR_reg[23]/NET0131 ,
		\P2_reg0_reg[16]/NET0131 ,
		_w1188_,
		_w4736_
	);
	LUT4 #(
		.INIT('h2000)
	) name4274 (
		\P2_reg0_reg[16]/NET0131 ,
		_w1189_,
		_w1352_,
		_w1356_,
		_w4737_
	);
	LUT4 #(
		.INIT('haaa8)
	) name4275 (
		\P2_reg0_reg[16]/NET0131 ,
		_w1361_,
		_w1363_,
		_w1368_,
		_w4738_
	);
	LUT3 #(
		.INIT('h54)
	) name4276 (
		_w1496_,
		_w3532_,
		_w4738_,
		_w4739_
	);
	LUT4 #(
		.INIT('h02aa)
	) name4277 (
		\P2_reg0_reg[16]/NET0131 ,
		_w1361_,
		_w1363_,
		_w1368_,
		_w4740_
	);
	LUT3 #(
		.INIT('ha8)
	) name4278 (
		_w1447_,
		_w3529_,
		_w4740_,
		_w4741_
	);
	LUT4 #(
		.INIT('h4b00)
	) name4279 (
		_w1217_,
		_w1206_,
		_w1294_,
		_w1411_,
		_w4742_
	);
	LUT3 #(
		.INIT('h54)
	) name4280 (
		_w1409_,
		_w4738_,
		_w4742_,
		_w4743_
	);
	LUT4 #(
		.INIT('h08c8)
	) name4281 (
		\P2_reg0_reg[16]/NET0131 ,
		_w1191_,
		_w1369_,
		_w3537_,
		_w4744_
	);
	LUT2 #(
		.INIT('h4)
	) name4282 (
		_w879_,
		_w1687_,
		_w4745_
	);
	LUT3 #(
		.INIT('ha2)
	) name4283 (
		\P2_reg0_reg[16]/NET0131 ,
		_w1684_,
		_w1685_,
		_w4746_
	);
	LUT2 #(
		.INIT('h1)
	) name4284 (
		_w4745_,
		_w4746_,
		_w4747_
	);
	LUT2 #(
		.INIT('h4)
	) name4285 (
		_w4744_,
		_w4747_,
		_w4748_
	);
	LUT4 #(
		.INIT('h0100)
	) name4286 (
		_w4741_,
		_w4739_,
		_w4743_,
		_w4748_,
		_w4749_
	);
	LUT4 #(
		.INIT('ha0a8)
	) name4287 (
		\P1_state_reg[0]/NET0131 ,
		_w1359_,
		_w4737_,
		_w4749_,
		_w4750_
	);
	LUT2 #(
		.INIT('he)
	) name4288 (
		_w4736_,
		_w4750_,
		_w4751_
	);
	LUT2 #(
		.INIT('h2)
	) name4289 (
		\P1_reg1_reg[9]/NET0131 ,
		_w2462_,
		_w4752_
	);
	LUT4 #(
		.INIT('h2000)
	) name4290 (
		\P1_reg1_reg[9]/NET0131 ,
		_w1723_,
		_w1727_,
		_w1730_,
		_w4753_
	);
	LUT2 #(
		.INIT('h2)
	) name4291 (
		\P1_reg1_reg[9]/NET0131 ,
		_w2520_,
		_w4754_
	);
	LUT4 #(
		.INIT('h35c5)
	) name4292 (
		\P1_reg1_reg[9]/NET0131 ,
		_w2327_,
		_w2520_,
		_w3186_,
		_w4755_
	);
	LUT4 #(
		.INIT('h6500)
	) name4293 (
		_w2040_,
		_w2104_,
		_w2431_,
		_w2520_,
		_w4756_
	);
	LUT2 #(
		.INIT('h8)
	) name4294 (
		_w2520_,
		_w4726_,
		_w4757_
	);
	LUT4 #(
		.INIT('h08aa)
	) name4295 (
		\P1_reg1_reg[9]/NET0131 ,
		_w2426_,
		_w2520_,
		_w2524_,
		_w4758_
	);
	LUT2 #(
		.INIT('h1)
	) name4296 (
		_w4757_,
		_w4758_,
		_w4759_
	);
	LUT4 #(
		.INIT('h5700)
	) name4297 (
		_w2447_,
		_w4754_,
		_w4756_,
		_w4759_,
		_w4760_
	);
	LUT3 #(
		.INIT('hd0)
	) name4298 (
		_w2388_,
		_w4755_,
		_w4760_,
		_w4761_
	);
	LUT4 #(
		.INIT('hc808)
	) name4299 (
		\P1_reg1_reg[9]/NET0131 ,
		_w2424_,
		_w2520_,
		_w4329_,
		_w4762_
	);
	LUT4 #(
		.INIT('h08c8)
	) name4300 (
		\P1_reg1_reg[9]/NET0131 ,
		_w2292_,
		_w2520_,
		_w4326_,
		_w4763_
	);
	LUT2 #(
		.INIT('h1)
	) name4301 (
		_w4762_,
		_w4763_,
		_w4764_
	);
	LUT4 #(
		.INIT('h3111)
	) name4302 (
		_w1731_,
		_w4753_,
		_w4761_,
		_w4764_,
		_w4765_
	);
	LUT3 #(
		.INIT('hce)
	) name4303 (
		\P1_state_reg[0]/NET0131 ,
		_w4752_,
		_w4765_,
		_w4766_
	);
	LUT4 #(
		.INIT('hd070)
	) name4304 (
		\P1_state_reg[0]/NET0131 ,
		\P2_IR_reg[23]/NET0131 ,
		\P2_reg0_reg[9]/NET0131 ,
		_w1188_,
		_w4767_
	);
	LUT4 #(
		.INIT('h2000)
	) name4305 (
		\P2_reg0_reg[9]/NET0131 ,
		_w1189_,
		_w1352_,
		_w1356_,
		_w4768_
	);
	LUT4 #(
		.INIT('h02aa)
	) name4306 (
		\P2_reg0_reg[9]/NET0131 ,
		_w1361_,
		_w1363_,
		_w1368_,
		_w4769_
	);
	LUT3 #(
		.INIT('he0)
	) name4307 (
		_w716_,
		_w718_,
		_w1442_,
		_w4770_
	);
	LUT2 #(
		.INIT('h8)
	) name4308 (
		_w1411_,
		_w4770_,
		_w4771_
	);
	LUT3 #(
		.INIT('ha2)
	) name4309 (
		\P2_reg0_reg[9]/NET0131 ,
		_w1684_,
		_w1685_,
		_w4772_
	);
	LUT2 #(
		.INIT('h1)
	) name4310 (
		_w4771_,
		_w4772_,
		_w4773_
	);
	LUT4 #(
		.INIT('h5700)
	) name4311 (
		_w1447_,
		_w4350_,
		_w4769_,
		_w4773_,
		_w4774_
	);
	LUT4 #(
		.INIT('haaa8)
	) name4312 (
		\P2_reg0_reg[9]/NET0131 ,
		_w1361_,
		_w1363_,
		_w1368_,
		_w4775_
	);
	LUT4 #(
		.INIT('h35c5)
	) name4313 (
		\P2_reg0_reg[9]/NET0131 ,
		_w1311_,
		_w1411_,
		_w1662_,
		_w4776_
	);
	LUT2 #(
		.INIT('h1)
	) name4314 (
		_w1409_,
		_w4776_,
		_w4777_
	);
	LUT4 #(
		.INIT('h111d)
	) name4315 (
		\P2_reg0_reg[9]/NET0131 ,
		_w1369_,
		_w4346_,
		_w4347_,
		_w4778_
	);
	LUT2 #(
		.INIT('h2)
	) name4316 (
		_w1191_,
		_w4778_,
		_w4779_
	);
	LUT3 #(
		.INIT('h54)
	) name4317 (
		_w1496_,
		_w4338_,
		_w4775_,
		_w4780_
	);
	LUT4 #(
		.INIT('h0100)
	) name4318 (
		_w4779_,
		_w4780_,
		_w4777_,
		_w4774_,
		_w4781_
	);
	LUT4 #(
		.INIT('ha0a8)
	) name4319 (
		\P1_state_reg[0]/NET0131 ,
		_w1359_,
		_w4768_,
		_w4781_,
		_w4782_
	);
	LUT2 #(
		.INIT('he)
	) name4320 (
		_w4767_,
		_w4782_,
		_w4783_
	);
	LUT4 #(
		.INIT('h20e0)
	) name4321 (
		\P1_reg2_reg[23]/NET0131 ,
		_w1741_,
		_w2292_,
		_w4362_,
		_w4784_
	);
	LUT4 #(
		.INIT('h20e0)
	) name4322 (
		\P1_reg2_reg[23]/NET0131 ,
		_w1741_,
		_w2388_,
		_w4368_,
		_w4785_
	);
	LUT4 #(
		.INIT('he020)
	) name4323 (
		\P1_reg2_reg[23]/NET0131 ,
		_w1741_,
		_w2424_,
		_w4371_,
		_w4786_
	);
	LUT4 #(
		.INIT('h0008)
	) name4324 (
		_w1959_,
		_w2284_,
		_w2288_,
		_w2291_,
		_w4787_
	);
	LUT4 #(
		.INIT('ha2a0)
	) name4325 (
		\P1_reg2_reg[23]/NET0131 ,
		_w1741_,
		_w2450_,
		_w2452_,
		_w4788_
	);
	LUT2 #(
		.INIT('h1)
	) name4326 (
		_w4787_,
		_w4788_,
		_w4789_
	);
	LUT3 #(
		.INIT('hd0)
	) name4327 (
		_w1741_,
		_w4374_,
		_w4789_,
		_w4790_
	);
	LUT2 #(
		.INIT('h4)
	) name4328 (
		_w4786_,
		_w4790_,
		_w4791_
	);
	LUT4 #(
		.INIT('ha8aa)
	) name4329 (
		_w1731_,
		_w4784_,
		_w4785_,
		_w4791_,
		_w4792_
	);
	LUT4 #(
		.INIT('h2000)
	) name4330 (
		\P1_reg2_reg[23]/NET0131 ,
		_w1723_,
		_w1727_,
		_w1730_,
		_w4793_
	);
	LUT2 #(
		.INIT('h2)
	) name4331 (
		\P1_reg2_reg[23]/NET0131 ,
		_w2462_,
		_w4794_
	);
	LUT4 #(
		.INIT('hffa8)
	) name4332 (
		\P1_state_reg[0]/NET0131 ,
		_w4792_,
		_w4793_,
		_w4794_,
		_w4795_
	);
	LUT4 #(
		.INIT('hd070)
	) name4333 (
		\P1_state_reg[0]/NET0131 ,
		\P2_IR_reg[23]/NET0131 ,
		\P2_reg1_reg[10]/NET0131 ,
		_w1188_,
		_w4796_
	);
	LUT4 #(
		.INIT('h2000)
	) name4334 (
		\P2_reg1_reg[10]/NET0131 ,
		_w1189_,
		_w1352_,
		_w1356_,
		_w4797_
	);
	LUT4 #(
		.INIT('ha8aa)
	) name4335 (
		\P2_reg1_reg[10]/NET0131 ,
		_w1361_,
		_w1363_,
		_w1368_,
		_w4798_
	);
	LUT4 #(
		.INIT('h08c8)
	) name4336 (
		\P2_reg1_reg[10]/NET0131 ,
		_w1191_,
		_w1507_,
		_w4258_,
		_w4799_
	);
	LUT4 #(
		.INIT('haa02)
	) name4337 (
		\P2_reg1_reg[10]/NET0131 ,
		_w1361_,
		_w1363_,
		_w1368_,
		_w4800_
	);
	LUT4 #(
		.INIT('h4844)
	) name4338 (
		_w1317_,
		_w1516_,
		_w2535_,
		_w2537_,
		_w4801_
	);
	LUT3 #(
		.INIT('he0)
	) name4339 (
		_w698_,
		_w702_,
		_w1442_,
		_w4802_
	);
	LUT2 #(
		.INIT('h8)
	) name4340 (
		_w1516_,
		_w4802_,
		_w4803_
	);
	LUT3 #(
		.INIT('ha2)
	) name4341 (
		\P2_reg1_reg[10]/NET0131 ,
		_w1684_,
		_w2469_,
		_w4804_
	);
	LUT2 #(
		.INIT('h1)
	) name4342 (
		_w4803_,
		_w4804_,
		_w4805_
	);
	LUT4 #(
		.INIT('hab00)
	) name4343 (
		_w1575_,
		_w4800_,
		_w4801_,
		_w4805_,
		_w4806_
	);
	LUT4 #(
		.INIT('h8848)
	) name4344 (
		_w1317_,
		_w1507_,
		_w2553_,
		_w2555_,
		_w4807_
	);
	LUT3 #(
		.INIT('ha8)
	) name4345 (
		_w1530_,
		_w4798_,
		_w4807_,
		_w4808_
	);
	LUT4 #(
		.INIT('h8848)
	) name4346 (
		_w1317_,
		_w1516_,
		_w2553_,
		_w2555_,
		_w4809_
	);
	LUT3 #(
		.INIT('h54)
	) name4347 (
		_w1506_,
		_w4800_,
		_w4809_,
		_w4810_
	);
	LUT4 #(
		.INIT('h0100)
	) name4348 (
		_w4808_,
		_w4810_,
		_w4799_,
		_w4806_,
		_w4811_
	);
	LUT4 #(
		.INIT('ha0a8)
	) name4349 (
		\P1_state_reg[0]/NET0131 ,
		_w1359_,
		_w4797_,
		_w4811_,
		_w4812_
	);
	LUT2 #(
		.INIT('he)
	) name4350 (
		_w4796_,
		_w4812_,
		_w4813_
	);
	LUT4 #(
		.INIT('hd070)
	) name4351 (
		\P1_state_reg[0]/NET0131 ,
		\P2_IR_reg[23]/NET0131 ,
		\P2_reg1_reg[12]/NET0131 ,
		_w1188_,
		_w4814_
	);
	LUT4 #(
		.INIT('h2000)
	) name4352 (
		\P2_reg1_reg[12]/NET0131 ,
		_w1189_,
		_w1352_,
		_w1356_,
		_w4815_
	);
	LUT4 #(
		.INIT('h0232)
	) name4353 (
		\P2_reg1_reg[12]/NET0131 ,
		_w1506_,
		_w1516_,
		_w4277_,
		_w4816_
	);
	LUT4 #(
		.INIT('h111d)
	) name4354 (
		\P2_reg1_reg[12]/NET0131 ,
		_w1507_,
		_w4280_,
		_w4281_,
		_w4817_
	);
	LUT4 #(
		.INIT('hf100)
	) name4355 (
		_w546_,
		_w661_,
		_w665_,
		_w1442_,
		_w4818_
	);
	LUT2 #(
		.INIT('h8)
	) name4356 (
		_w1516_,
		_w4818_,
		_w4819_
	);
	LUT3 #(
		.INIT('ha2)
	) name4357 (
		\P2_reg1_reg[12]/NET0131 ,
		_w1684_,
		_w2469_,
		_w4820_
	);
	LUT2 #(
		.INIT('h1)
	) name4358 (
		_w4819_,
		_w4820_,
		_w4821_
	);
	LUT3 #(
		.INIT('hd0)
	) name4359 (
		_w1191_,
		_w4817_,
		_w4821_,
		_w4822_
	);
	LUT4 #(
		.INIT('h20e0)
	) name4360 (
		\P2_reg1_reg[12]/NET0131 ,
		_w1507_,
		_w1530_,
		_w4277_,
		_w4823_
	);
	LUT4 #(
		.INIT('h0e02)
	) name4361 (
		\P2_reg1_reg[12]/NET0131 ,
		_w1516_,
		_w1575_,
		_w4287_,
		_w4824_
	);
	LUT4 #(
		.INIT('h0100)
	) name4362 (
		_w4816_,
		_w4823_,
		_w4824_,
		_w4822_,
		_w4825_
	);
	LUT4 #(
		.INIT('ha0a8)
	) name4363 (
		\P1_state_reg[0]/NET0131 ,
		_w1359_,
		_w4815_,
		_w4825_,
		_w4826_
	);
	LUT2 #(
		.INIT('he)
	) name4364 (
		_w4814_,
		_w4826_,
		_w4827_
	);
	LUT4 #(
		.INIT('hd070)
	) name4365 (
		\P1_state_reg[0]/NET0131 ,
		\P2_IR_reg[23]/NET0131 ,
		\P2_reg1_reg[13]/NET0131 ,
		_w1188_,
		_w4828_
	);
	LUT4 #(
		.INIT('h2000)
	) name4366 (
		\P2_reg1_reg[13]/NET0131 ,
		_w1189_,
		_w1352_,
		_w1356_,
		_w4829_
	);
	LUT4 #(
		.INIT('hc535)
	) name4367 (
		\P2_reg1_reg[13]/NET0131 ,
		_w1299_,
		_w1516_,
		_w1699_,
		_w4830_
	);
	LUT4 #(
		.INIT('h08c8)
	) name4368 (
		\P2_reg1_reg[13]/NET0131 ,
		_w1191_,
		_w1507_,
		_w4301_,
		_w4831_
	);
	LUT4 #(
		.INIT('hf100)
	) name4369 (
		_w546_,
		_w642_,
		_w644_,
		_w1442_,
		_w4832_
	);
	LUT2 #(
		.INIT('h8)
	) name4370 (
		_w1516_,
		_w4832_,
		_w4833_
	);
	LUT3 #(
		.INIT('ha2)
	) name4371 (
		\P2_reg1_reg[13]/NET0131 ,
		_w1684_,
		_w2469_,
		_w4834_
	);
	LUT2 #(
		.INIT('h1)
	) name4372 (
		_w4833_,
		_w4834_,
		_w4835_
	);
	LUT4 #(
		.INIT('h0e00)
	) name4373 (
		_w1575_,
		_w4830_,
		_w4831_,
		_w4835_,
		_w4836_
	);
	LUT4 #(
		.INIT('he020)
	) name4374 (
		\P2_reg1_reg[13]/NET0131 ,
		_w1507_,
		_w1530_,
		_w4309_,
		_w4837_
	);
	LUT4 #(
		.INIT('h3202)
	) name4375 (
		\P2_reg1_reg[13]/NET0131 ,
		_w1506_,
		_w1516_,
		_w4309_,
		_w4838_
	);
	LUT2 #(
		.INIT('h1)
	) name4376 (
		_w4837_,
		_w4838_,
		_w4839_
	);
	LUT4 #(
		.INIT('h3111)
	) name4377 (
		_w1359_,
		_w4829_,
		_w4836_,
		_w4839_,
		_w4840_
	);
	LUT3 #(
		.INIT('hce)
	) name4378 (
		\P1_state_reg[0]/NET0131 ,
		_w4828_,
		_w4840_,
		_w4841_
	);
	LUT4 #(
		.INIT('hd070)
	) name4379 (
		\P1_state_reg[0]/NET0131 ,
		\P2_IR_reg[23]/NET0131 ,
		\P2_reg1_reg[16]/NET0131 ,
		_w1188_,
		_w4842_
	);
	LUT4 #(
		.INIT('h2000)
	) name4380 (
		\P2_reg1_reg[16]/NET0131 ,
		_w1189_,
		_w1352_,
		_w1356_,
		_w4843_
	);
	LUT4 #(
		.INIT('haa02)
	) name4381 (
		\P2_reg1_reg[16]/NET0131 ,
		_w1361_,
		_w1363_,
		_w1368_,
		_w4844_
	);
	LUT4 #(
		.INIT('h8848)
	) name4382 (
		_w1294_,
		_w1516_,
		_w1553_,
		_w3528_,
		_w4845_
	);
	LUT3 #(
		.INIT('h54)
	) name4383 (
		_w1575_,
		_w4844_,
		_w4845_,
		_w4846_
	);
	LUT4 #(
		.INIT('h4b00)
	) name4384 (
		_w1217_,
		_w1206_,
		_w1294_,
		_w1516_,
		_w4847_
	);
	LUT3 #(
		.INIT('h54)
	) name4385 (
		_w1506_,
		_w4844_,
		_w4847_,
		_w4848_
	);
	LUT4 #(
		.INIT('ha8aa)
	) name4386 (
		\P2_reg1_reg[16]/NET0131 ,
		_w1361_,
		_w1363_,
		_w1368_,
		_w4849_
	);
	LUT4 #(
		.INIT('h4b00)
	) name4387 (
		_w1217_,
		_w1206_,
		_w1294_,
		_w1507_,
		_w4850_
	);
	LUT3 #(
		.INIT('ha8)
	) name4388 (
		_w1530_,
		_w4849_,
		_w4850_,
		_w4851_
	);
	LUT4 #(
		.INIT('h08c8)
	) name4389 (
		\P2_reg1_reg[16]/NET0131 ,
		_w1191_,
		_w1507_,
		_w3537_,
		_w4852_
	);
	LUT3 #(
		.INIT('ha2)
	) name4390 (
		\P2_reg1_reg[16]/NET0131 ,
		_w1684_,
		_w2469_,
		_w4853_
	);
	LUT2 #(
		.INIT('h4)
	) name4391 (
		_w879_,
		_w2471_,
		_w4854_
	);
	LUT2 #(
		.INIT('h1)
	) name4392 (
		_w4853_,
		_w4854_,
		_w4855_
	);
	LUT2 #(
		.INIT('h4)
	) name4393 (
		_w4852_,
		_w4855_,
		_w4856_
	);
	LUT4 #(
		.INIT('h0100)
	) name4394 (
		_w4851_,
		_w4848_,
		_w4846_,
		_w4856_,
		_w4857_
	);
	LUT4 #(
		.INIT('ha0a8)
	) name4395 (
		\P1_state_reg[0]/NET0131 ,
		_w1359_,
		_w4843_,
		_w4857_,
		_w4858_
	);
	LUT2 #(
		.INIT('he)
	) name4396 (
		_w4842_,
		_w4858_,
		_w4859_
	);
	LUT2 #(
		.INIT('h2)
	) name4397 (
		\P1_reg2_reg[30]/NET0131 ,
		_w2462_,
		_w4860_
	);
	LUT4 #(
		.INIT('h2000)
	) name4398 (
		\P1_reg2_reg[30]/NET0131 ,
		_w1723_,
		_w1727_,
		_w1730_,
		_w4861_
	);
	LUT4 #(
		.INIT('h40bf)
	) name4399 (
		_w2273_,
		_w2443_,
		_w2444_,
		_w3135_,
		_w4862_
	);
	LUT3 #(
		.INIT('he0)
	) name4400 (
		\P1_reg2_reg[30]/NET0131 ,
		_w1741_,
		_w2447_,
		_w4863_
	);
	LUT3 #(
		.INIT('hd0)
	) name4401 (
		_w1741_,
		_w4862_,
		_w4863_,
		_w4864_
	);
	LUT2 #(
		.INIT('h8)
	) name4402 (
		_w1741_,
		_w2426_,
		_w4865_
	);
	LUT3 #(
		.INIT('h10)
	) name4403 (
		_w1748_,
		_w3134_,
		_w4865_,
		_w4866_
	);
	LUT4 #(
		.INIT('haa02)
	) name4404 (
		\P1_reg2_reg[30]/NET0131 ,
		_w1741_,
		_w2446_,
		_w2450_,
		_w4867_
	);
	LUT2 #(
		.INIT('h1)
	) name4405 (
		_w2455_,
		_w4867_,
		_w4868_
	);
	LUT2 #(
		.INIT('h4)
	) name4406 (
		_w4866_,
		_w4868_,
		_w4869_
	);
	LUT4 #(
		.INIT('ha8aa)
	) name4407 (
		_w1731_,
		_w3572_,
		_w4864_,
		_w4869_,
		_w4870_
	);
	LUT4 #(
		.INIT('heeec)
	) name4408 (
		\P1_state_reg[0]/NET0131 ,
		_w4860_,
		_w4861_,
		_w4870_,
		_w4871_
	);
	LUT4 #(
		.INIT('hd070)
	) name4409 (
		\P1_state_reg[0]/NET0131 ,
		\P2_IR_reg[23]/NET0131 ,
		\P2_reg1_reg[9]/NET0131 ,
		_w1188_,
		_w4872_
	);
	LUT4 #(
		.INIT('h2000)
	) name4410 (
		\P2_reg1_reg[9]/NET0131 ,
		_w1189_,
		_w1352_,
		_w1356_,
		_w4873_
	);
	LUT4 #(
		.INIT('h111d)
	) name4411 (
		\P2_reg1_reg[9]/NET0131 ,
		_w1507_,
		_w4346_,
		_w4347_,
		_w4874_
	);
	LUT2 #(
		.INIT('h8)
	) name4412 (
		_w1516_,
		_w4770_,
		_w4875_
	);
	LUT3 #(
		.INIT('ha2)
	) name4413 (
		\P2_reg1_reg[9]/NET0131 ,
		_w1684_,
		_w2469_,
		_w4876_
	);
	LUT2 #(
		.INIT('h1)
	) name4414 (
		_w4875_,
		_w4876_,
		_w4877_
	);
	LUT3 #(
		.INIT('hd0)
	) name4415 (
		_w1191_,
		_w4874_,
		_w4877_,
		_w4878_
	);
	LUT4 #(
		.INIT('haa02)
	) name4416 (
		\P2_reg1_reg[9]/NET0131 ,
		_w1361_,
		_w1363_,
		_w1368_,
		_w4879_
	);
	LUT4 #(
		.INIT('h8488)
	) name4417 (
		_w1311_,
		_w1516_,
		_w1695_,
		_w1696_,
		_w4880_
	);
	LUT3 #(
		.INIT('h54)
	) name4418 (
		_w1575_,
		_w4879_,
		_w4880_,
		_w4881_
	);
	LUT4 #(
		.INIT('h35c5)
	) name4419 (
		\P2_reg1_reg[9]/NET0131 ,
		_w1311_,
		_w1507_,
		_w1662_,
		_w4882_
	);
	LUT4 #(
		.INIT('h35c5)
	) name4420 (
		\P2_reg1_reg[9]/NET0131 ,
		_w1311_,
		_w1516_,
		_w1662_,
		_w4883_
	);
	LUT4 #(
		.INIT('hf3a2)
	) name4421 (
		_w1506_,
		_w1530_,
		_w4882_,
		_w4883_,
		_w4884_
	);
	LUT4 #(
		.INIT('h8aaa)
	) name4422 (
		_w1359_,
		_w4881_,
		_w4878_,
		_w4884_,
		_w4885_
	);
	LUT4 #(
		.INIT('heeec)
	) name4423 (
		\P1_state_reg[0]/NET0131 ,
		_w4872_,
		_w4873_,
		_w4885_,
		_w4886_
	);
	LUT4 #(
		.INIT('hd070)
	) name4424 (
		\P1_state_reg[0]/NET0131 ,
		\P2_IR_reg[23]/NET0131 ,
		\P2_reg2_reg[10]/NET0131 ,
		_w1188_,
		_w4887_
	);
	LUT4 #(
		.INIT('h2000)
	) name4425 (
		\P2_reg2_reg[10]/NET0131 ,
		_w1189_,
		_w1352_,
		_w1356_,
		_w4888_
	);
	LUT4 #(
		.INIT('haa02)
	) name4426 (
		\P2_reg2_reg[10]/NET0131 ,
		_w1361_,
		_w1363_,
		_w1368_,
		_w4889_
	);
	LUT4 #(
		.INIT('h08c8)
	) name4427 (
		\P2_reg2_reg[10]/NET0131 ,
		_w1191_,
		_w1516_,
		_w4258_,
		_w4890_
	);
	LUT4 #(
		.INIT('ha8aa)
	) name4428 (
		\P2_reg2_reg[10]/NET0131 ,
		_w1361_,
		_w1363_,
		_w1368_,
		_w4891_
	);
	LUT4 #(
		.INIT('h4844)
	) name4429 (
		_w1317_,
		_w1507_,
		_w2535_,
		_w2537_,
		_w4892_
	);
	LUT3 #(
		.INIT('ha8)
	) name4430 (
		\P2_reg2_reg[10]/NET0131 ,
		_w1441_,
		_w1523_,
		_w4893_
	);
	LUT3 #(
		.INIT('h40)
	) name4431 (
		_w690_,
		_w1229_,
		_w1232_,
		_w4894_
	);
	LUT3 #(
		.INIT('h07)
	) name4432 (
		_w1507_,
		_w4802_,
		_w4894_,
		_w4895_
	);
	LUT2 #(
		.INIT('h4)
	) name4433 (
		_w4893_,
		_w4895_,
		_w4896_
	);
	LUT4 #(
		.INIT('hab00)
	) name4434 (
		_w1575_,
		_w4891_,
		_w4892_,
		_w4896_,
		_w4897_
	);
	LUT3 #(
		.INIT('ha8)
	) name4435 (
		_w1530_,
		_w4809_,
		_w4889_,
		_w4898_
	);
	LUT3 #(
		.INIT('h54)
	) name4436 (
		_w1506_,
		_w4807_,
		_w4891_,
		_w4899_
	);
	LUT4 #(
		.INIT('h0100)
	) name4437 (
		_w4898_,
		_w4899_,
		_w4890_,
		_w4897_,
		_w4900_
	);
	LUT4 #(
		.INIT('ha0a8)
	) name4438 (
		\P1_state_reg[0]/NET0131 ,
		_w1359_,
		_w4888_,
		_w4900_,
		_w4901_
	);
	LUT2 #(
		.INIT('he)
	) name4439 (
		_w4887_,
		_w4901_,
		_w4902_
	);
	LUT4 #(
		.INIT('hd070)
	) name4440 (
		\P1_state_reg[0]/NET0131 ,
		\P2_IR_reg[23]/NET0131 ,
		\P2_reg2_reg[12]/NET0131 ,
		_w1188_,
		_w4903_
	);
	LUT4 #(
		.INIT('h2000)
	) name4441 (
		\P2_reg2_reg[12]/NET0131 ,
		_w1189_,
		_w1352_,
		_w1356_,
		_w4904_
	);
	LUT4 #(
		.INIT('h0e02)
	) name4442 (
		\P2_reg2_reg[12]/NET0131 ,
		_w1507_,
		_w1575_,
		_w4287_,
		_w4905_
	);
	LUT4 #(
		.INIT('h111d)
	) name4443 (
		\P2_reg2_reg[12]/NET0131 ,
		_w1516_,
		_w4280_,
		_w4281_,
		_w4906_
	);
	LUT3 #(
		.INIT('ha8)
	) name4444 (
		\P2_reg2_reg[12]/NET0131 ,
		_w1441_,
		_w1523_,
		_w4907_
	);
	LUT3 #(
		.INIT('h40)
	) name4445 (
		_w648_,
		_w1229_,
		_w1232_,
		_w4908_
	);
	LUT3 #(
		.INIT('h07)
	) name4446 (
		_w1507_,
		_w4818_,
		_w4908_,
		_w4909_
	);
	LUT2 #(
		.INIT('h4)
	) name4447 (
		_w4907_,
		_w4909_,
		_w4910_
	);
	LUT3 #(
		.INIT('hd0)
	) name4448 (
		_w1191_,
		_w4906_,
		_w4910_,
		_w4911_
	);
	LUT4 #(
		.INIT('h20e0)
	) name4449 (
		\P2_reg2_reg[12]/NET0131 ,
		_w1516_,
		_w1530_,
		_w4277_,
		_w4912_
	);
	LUT4 #(
		.INIT('h0232)
	) name4450 (
		\P2_reg2_reg[12]/NET0131 ,
		_w1506_,
		_w1507_,
		_w4277_,
		_w4913_
	);
	LUT4 #(
		.INIT('h0100)
	) name4451 (
		_w4905_,
		_w4912_,
		_w4913_,
		_w4911_,
		_w4914_
	);
	LUT4 #(
		.INIT('ha0a8)
	) name4452 (
		\P1_state_reg[0]/NET0131 ,
		_w1359_,
		_w4904_,
		_w4914_,
		_w4915_
	);
	LUT2 #(
		.INIT('he)
	) name4453 (
		_w4903_,
		_w4915_,
		_w4916_
	);
	LUT4 #(
		.INIT('hd070)
	) name4454 (
		\P1_state_reg[0]/NET0131 ,
		\P2_IR_reg[23]/NET0131 ,
		\P2_reg2_reg[13]/NET0131 ,
		_w1188_,
		_w4917_
	);
	LUT4 #(
		.INIT('h2000)
	) name4455 (
		\P2_reg2_reg[13]/NET0131 ,
		_w1189_,
		_w1352_,
		_w1356_,
		_w4918_
	);
	LUT4 #(
		.INIT('hc535)
	) name4456 (
		\P2_reg2_reg[13]/NET0131 ,
		_w1299_,
		_w1507_,
		_w1699_,
		_w4919_
	);
	LUT4 #(
		.INIT('h08c8)
	) name4457 (
		\P2_reg2_reg[13]/NET0131 ,
		_w1191_,
		_w1516_,
		_w4301_,
		_w4920_
	);
	LUT3 #(
		.INIT('ha8)
	) name4458 (
		\P2_reg2_reg[13]/NET0131 ,
		_w1441_,
		_w1523_,
		_w4921_
	);
	LUT3 #(
		.INIT('h40)
	) name4459 (
		_w627_,
		_w1229_,
		_w1232_,
		_w4922_
	);
	LUT3 #(
		.INIT('h07)
	) name4460 (
		_w1507_,
		_w4832_,
		_w4922_,
		_w4923_
	);
	LUT2 #(
		.INIT('h4)
	) name4461 (
		_w4921_,
		_w4923_,
		_w4924_
	);
	LUT4 #(
		.INIT('h3200)
	) name4462 (
		_w1575_,
		_w4920_,
		_w4919_,
		_w4924_,
		_w4925_
	);
	LUT4 #(
		.INIT('he020)
	) name4463 (
		\P2_reg2_reg[13]/NET0131 ,
		_w1516_,
		_w1530_,
		_w4309_,
		_w4926_
	);
	LUT4 #(
		.INIT('h3202)
	) name4464 (
		\P2_reg2_reg[13]/NET0131 ,
		_w1506_,
		_w1507_,
		_w4309_,
		_w4927_
	);
	LUT2 #(
		.INIT('h1)
	) name4465 (
		_w4926_,
		_w4927_,
		_w4928_
	);
	LUT4 #(
		.INIT('h3111)
	) name4466 (
		_w1359_,
		_w4918_,
		_w4925_,
		_w4928_,
		_w4929_
	);
	LUT3 #(
		.INIT('hce)
	) name4467 (
		\P1_state_reg[0]/NET0131 ,
		_w4917_,
		_w4929_,
		_w4930_
	);
	LUT4 #(
		.INIT('hd070)
	) name4468 (
		\P1_state_reg[0]/NET0131 ,
		\P2_IR_reg[23]/NET0131 ,
		\P2_reg2_reg[16]/NET0131 ,
		_w1188_,
		_w4931_
	);
	LUT4 #(
		.INIT('h2000)
	) name4469 (
		\P2_reg2_reg[16]/NET0131 ,
		_w1189_,
		_w1352_,
		_w1356_,
		_w4932_
	);
	LUT4 #(
		.INIT('ha8aa)
	) name4470 (
		\P2_reg2_reg[16]/NET0131 ,
		_w1361_,
		_w1363_,
		_w1368_,
		_w4933_
	);
	LUT4 #(
		.INIT('h8848)
	) name4471 (
		_w1294_,
		_w1507_,
		_w1553_,
		_w3528_,
		_w4934_
	);
	LUT3 #(
		.INIT('h54)
	) name4472 (
		_w1575_,
		_w4933_,
		_w4934_,
		_w4935_
	);
	LUT3 #(
		.INIT('h54)
	) name4473 (
		_w1506_,
		_w4850_,
		_w4933_,
		_w4936_
	);
	LUT4 #(
		.INIT('haa02)
	) name4474 (
		\P2_reg2_reg[16]/NET0131 ,
		_w1361_,
		_w1363_,
		_w1368_,
		_w4937_
	);
	LUT3 #(
		.INIT('ha8)
	) name4475 (
		_w1530_,
		_w4847_,
		_w4937_,
		_w4938_
	);
	LUT4 #(
		.INIT('h08c8)
	) name4476 (
		\P2_reg2_reg[16]/NET0131 ,
		_w1191_,
		_w1516_,
		_w3537_,
		_w4939_
	);
	LUT3 #(
		.INIT('ha8)
	) name4477 (
		\P2_reg2_reg[16]/NET0131 ,
		_w1441_,
		_w1523_,
		_w4940_
	);
	LUT3 #(
		.INIT('h40)
	) name4478 (
		_w863_,
		_w1229_,
		_w1232_,
		_w4941_
	);
	LUT3 #(
		.INIT('h0b)
	) name4479 (
		_w879_,
		_w1522_,
		_w4941_,
		_w4942_
	);
	LUT2 #(
		.INIT('h4)
	) name4480 (
		_w4940_,
		_w4942_,
		_w4943_
	);
	LUT2 #(
		.INIT('h4)
	) name4481 (
		_w4939_,
		_w4943_,
		_w4944_
	);
	LUT4 #(
		.INIT('h0100)
	) name4482 (
		_w4938_,
		_w4936_,
		_w4935_,
		_w4944_,
		_w4945_
	);
	LUT4 #(
		.INIT('ha0a8)
	) name4483 (
		\P1_state_reg[0]/NET0131 ,
		_w1359_,
		_w4932_,
		_w4945_,
		_w4946_
	);
	LUT2 #(
		.INIT('he)
	) name4484 (
		_w4931_,
		_w4946_,
		_w4947_
	);
	LUT2 #(
		.INIT('h2)
	) name4485 (
		\P1_reg0_reg[10]/NET0131 ,
		_w2462_,
		_w4948_
	);
	LUT4 #(
		.INIT('h2000)
	) name4486 (
		\P1_reg0_reg[10]/NET0131 ,
		_w1723_,
		_w1727_,
		_w1730_,
		_w4949_
	);
	LUT4 #(
		.INIT('hddd1)
	) name4487 (
		\P1_reg0_reg[10]/NET0131 ,
		_w2883_,
		_w4217_,
		_w4218_,
		_w4950_
	);
	LUT2 #(
		.INIT('h2)
	) name4488 (
		_w2424_,
		_w4950_,
		_w4951_
	);
	LUT4 #(
		.INIT('h1dd1)
	) name4489 (
		\P1_reg0_reg[10]/NET0131 ,
		_w2883_,
		_w2953_,
		_w3176_,
		_w4952_
	);
	LUT2 #(
		.INIT('h2)
	) name4490 (
		_w2292_,
		_w4952_,
		_w4953_
	);
	LUT4 #(
		.INIT('hd11d)
	) name4491 (
		\P1_reg0_reg[10]/NET0131 ,
		_w2883_,
		_w2935_,
		_w3176_,
		_w4954_
	);
	LUT4 #(
		.INIT('hc808)
	) name4492 (
		\P1_reg0_reg[10]/NET0131 ,
		_w2447_,
		_w2883_,
		_w4224_,
		_w4955_
	);
	LUT2 #(
		.INIT('h8)
	) name4493 (
		_w2883_,
		_w4697_,
		_w4956_
	);
	LUT4 #(
		.INIT('h0a8a)
	) name4494 (
		\P1_reg0_reg[10]/NET0131 ,
		_w2426_,
		_w2524_,
		_w2883_,
		_w4957_
	);
	LUT2 #(
		.INIT('h1)
	) name4495 (
		_w4956_,
		_w4957_,
		_w4958_
	);
	LUT2 #(
		.INIT('h4)
	) name4496 (
		_w4955_,
		_w4958_,
		_w4959_
	);
	LUT3 #(
		.INIT('hd0)
	) name4497 (
		_w2388_,
		_w4954_,
		_w4959_,
		_w4960_
	);
	LUT4 #(
		.INIT('ha8aa)
	) name4498 (
		_w1731_,
		_w4951_,
		_w4953_,
		_w4960_,
		_w4961_
	);
	LUT4 #(
		.INIT('heeec)
	) name4499 (
		\P1_state_reg[0]/NET0131 ,
		_w4948_,
		_w4949_,
		_w4961_,
		_w4962_
	);
	LUT4 #(
		.INIT('hd070)
	) name4500 (
		\P1_state_reg[0]/NET0131 ,
		\P2_IR_reg[23]/NET0131 ,
		\P2_reg2_reg[9]/NET0131 ,
		_w1188_,
		_w4963_
	);
	LUT4 #(
		.INIT('h2000)
	) name4501 (
		\P2_reg2_reg[9]/NET0131 ,
		_w1189_,
		_w1352_,
		_w1356_,
		_w4964_
	);
	LUT4 #(
		.INIT('h111d)
	) name4502 (
		\P2_reg2_reg[9]/NET0131 ,
		_w1516_,
		_w4346_,
		_w4347_,
		_w4965_
	);
	LUT3 #(
		.INIT('ha8)
	) name4503 (
		\P2_reg2_reg[9]/NET0131 ,
		_w1441_,
		_w1523_,
		_w4966_
	);
	LUT3 #(
		.INIT('h40)
	) name4504 (
		_w707_,
		_w1229_,
		_w1232_,
		_w4967_
	);
	LUT3 #(
		.INIT('h07)
	) name4505 (
		_w1507_,
		_w4770_,
		_w4967_,
		_w4968_
	);
	LUT2 #(
		.INIT('h4)
	) name4506 (
		_w4966_,
		_w4968_,
		_w4969_
	);
	LUT3 #(
		.INIT('hd0)
	) name4507 (
		_w1191_,
		_w4965_,
		_w4969_,
		_w4970_
	);
	LUT4 #(
		.INIT('ha8aa)
	) name4508 (
		\P2_reg2_reg[9]/NET0131 ,
		_w1361_,
		_w1363_,
		_w1368_,
		_w4971_
	);
	LUT4 #(
		.INIT('h8488)
	) name4509 (
		_w1311_,
		_w1507_,
		_w1695_,
		_w1696_,
		_w4972_
	);
	LUT3 #(
		.INIT('h54)
	) name4510 (
		_w1575_,
		_w4971_,
		_w4972_,
		_w4973_
	);
	LUT4 #(
		.INIT('h35c5)
	) name4511 (
		\P2_reg2_reg[9]/NET0131 ,
		_w1311_,
		_w1516_,
		_w1662_,
		_w4974_
	);
	LUT4 #(
		.INIT('h35c5)
	) name4512 (
		\P2_reg2_reg[9]/NET0131 ,
		_w1311_,
		_w1507_,
		_w1662_,
		_w4975_
	);
	LUT4 #(
		.INIT('hf3a2)
	) name4513 (
		_w1506_,
		_w1530_,
		_w4974_,
		_w4975_,
		_w4976_
	);
	LUT4 #(
		.INIT('h8aaa)
	) name4514 (
		_w1359_,
		_w4973_,
		_w4970_,
		_w4976_,
		_w4977_
	);
	LUT4 #(
		.INIT('heeec)
	) name4515 (
		\P1_state_reg[0]/NET0131 ,
		_w4963_,
		_w4964_,
		_w4977_,
		_w4978_
	);
	LUT2 #(
		.INIT('h2)
	) name4516 (
		\P1_reg0_reg[13]/NET0131 ,
		_w2462_,
		_w4979_
	);
	LUT4 #(
		.INIT('h2000)
	) name4517 (
		\P1_reg0_reg[13]/NET0131 ,
		_w1723_,
		_w1727_,
		_w1730_,
		_w4980_
	);
	LUT2 #(
		.INIT('h2)
	) name4518 (
		\P1_reg0_reg[13]/NET0131 ,
		_w2883_,
		_w4981_
	);
	LUT4 #(
		.INIT('h7020)
	) name4519 (
		_w1747_,
		_w2020_,
		_w2883_,
		_w4237_,
		_w4982_
	);
	LUT2 #(
		.INIT('h2)
	) name4520 (
		\P1_reg0_reg[13]/NET0131 ,
		_w3420_,
		_w4983_
	);
	LUT4 #(
		.INIT('h0057)
	) name4521 (
		_w2883_,
		_w4240_,
		_w4708_,
		_w4983_,
		_w4984_
	);
	LUT4 #(
		.INIT('h5700)
	) name4522 (
		_w2424_,
		_w4981_,
		_w4982_,
		_w4984_,
		_w4985_
	);
	LUT4 #(
		.INIT('h20d0)
	) name4523 (
		_w2049_,
		_w2153_,
		_w2883_,
		_w3192_,
		_w4986_
	);
	LUT3 #(
		.INIT('ha8)
	) name4524 (
		_w2292_,
		_w4981_,
		_w4986_,
		_w4987_
	);
	LUT4 #(
		.INIT('h08c8)
	) name4525 (
		\P1_reg0_reg[13]/NET0131 ,
		_w2388_,
		_w2883_,
		_w4245_,
		_w4988_
	);
	LUT4 #(
		.INIT('ha8aa)
	) name4526 (
		_w1731_,
		_w4987_,
		_w4988_,
		_w4985_,
		_w4989_
	);
	LUT4 #(
		.INIT('heeec)
	) name4527 (
		\P1_state_reg[0]/NET0131 ,
		_w4979_,
		_w4980_,
		_w4989_,
		_w4990_
	);
	LUT2 #(
		.INIT('h2)
	) name4528 (
		\P1_reg0_reg[23]/NET0131 ,
		_w2462_,
		_w4991_
	);
	LUT4 #(
		.INIT('h08c8)
	) name4529 (
		\P1_reg0_reg[23]/NET0131 ,
		_w2292_,
		_w2883_,
		_w4362_,
		_w4992_
	);
	LUT4 #(
		.INIT('h08c8)
	) name4530 (
		\P1_reg0_reg[23]/NET0131 ,
		_w2388_,
		_w2883_,
		_w4368_,
		_w4993_
	);
	LUT4 #(
		.INIT('hc808)
	) name4531 (
		\P1_reg0_reg[23]/NET0131 ,
		_w2424_,
		_w2883_,
		_w4371_,
		_w4994_
	);
	LUT4 #(
		.INIT('h0a8a)
	) name4532 (
		\P1_reg0_reg[23]/NET0131 ,
		_w2452_,
		_w2524_,
		_w2883_,
		_w4995_
	);
	LUT3 #(
		.INIT('h0d)
	) name4533 (
		_w2883_,
		_w4374_,
		_w4995_,
		_w4996_
	);
	LUT2 #(
		.INIT('h4)
	) name4534 (
		_w4994_,
		_w4996_,
		_w4997_
	);
	LUT4 #(
		.INIT('ha8aa)
	) name4535 (
		_w1731_,
		_w4992_,
		_w4993_,
		_w4997_,
		_w4998_
	);
	LUT4 #(
		.INIT('h2000)
	) name4536 (
		\P1_reg0_reg[23]/NET0131 ,
		_w1723_,
		_w1727_,
		_w1730_,
		_w4999_
	);
	LUT4 #(
		.INIT('heeec)
	) name4537 (
		\P1_state_reg[0]/NET0131 ,
		_w4991_,
		_w4998_,
		_w4999_,
		_w5000_
	);
	LUT2 #(
		.INIT('h2)
	) name4538 (
		\P1_reg0_reg[30]/NET0131 ,
		_w2462_,
		_w5001_
	);
	LUT4 #(
		.INIT('h2000)
	) name4539 (
		\P1_reg0_reg[30]/NET0131 ,
		_w1723_,
		_w1727_,
		_w1730_,
		_w5002_
	);
	LUT4 #(
		.INIT('hc808)
	) name4540 (
		\P1_reg0_reg[30]/NET0131 ,
		_w2447_,
		_w2883_,
		_w4862_,
		_w5003_
	);
	LUT4 #(
		.INIT('hf5c5)
	) name4541 (
		\P1_reg0_reg[30]/NET0131 ,
		_w1748_,
		_w2883_,
		_w3134_,
		_w5004_
	);
	LUT4 #(
		.INIT('h222a)
	) name4542 (
		\P1_reg0_reg[30]/NET0131 ,
		_w2524_,
		_w2883_,
		_w3574_,
		_w5005_
	);
	LUT3 #(
		.INIT('h0d)
	) name4543 (
		_w2426_,
		_w5004_,
		_w5005_,
		_w5006_
	);
	LUT4 #(
		.INIT('ha8aa)
	) name4544 (
		_w1731_,
		_w4163_,
		_w5003_,
		_w5006_,
		_w5007_
	);
	LUT4 #(
		.INIT('heeec)
	) name4545 (
		\P1_state_reg[0]/NET0131 ,
		_w5001_,
		_w5002_,
		_w5007_,
		_w5008_
	);
	LUT2 #(
		.INIT('h2)
	) name4546 (
		\P1_reg0_reg[9]/NET0131 ,
		_w2462_,
		_w5009_
	);
	LUT4 #(
		.INIT('h2000)
	) name4547 (
		\P1_reg0_reg[9]/NET0131 ,
		_w1723_,
		_w1727_,
		_w1730_,
		_w5010_
	);
	LUT2 #(
		.INIT('h2)
	) name4548 (
		\P1_reg0_reg[9]/NET0131 ,
		_w2883_,
		_w5011_
	);
	LUT4 #(
		.INIT('h35c5)
	) name4549 (
		\P1_reg0_reg[9]/NET0131 ,
		_w2327_,
		_w2883_,
		_w3186_,
		_w5012_
	);
	LUT4 #(
		.INIT('h6500)
	) name4550 (
		_w2040_,
		_w2104_,
		_w2431_,
		_w2883_,
		_w5013_
	);
	LUT2 #(
		.INIT('h8)
	) name4551 (
		_w2883_,
		_w4726_,
		_w5014_
	);
	LUT4 #(
		.INIT('h0a8a)
	) name4552 (
		\P1_reg0_reg[9]/NET0131 ,
		_w2426_,
		_w2524_,
		_w2883_,
		_w5015_
	);
	LUT2 #(
		.INIT('h1)
	) name4553 (
		_w5014_,
		_w5015_,
		_w5016_
	);
	LUT4 #(
		.INIT('h5700)
	) name4554 (
		_w2447_,
		_w5011_,
		_w5013_,
		_w5016_,
		_w5017_
	);
	LUT3 #(
		.INIT('hd0)
	) name4555 (
		_w2388_,
		_w5012_,
		_w5017_,
		_w5018_
	);
	LUT4 #(
		.INIT('hc808)
	) name4556 (
		\P1_reg0_reg[9]/NET0131 ,
		_w2424_,
		_w2883_,
		_w4329_,
		_w5019_
	);
	LUT4 #(
		.INIT('h08c8)
	) name4557 (
		\P1_reg0_reg[9]/NET0131 ,
		_w2292_,
		_w2883_,
		_w4326_,
		_w5020_
	);
	LUT2 #(
		.INIT('h1)
	) name4558 (
		_w5019_,
		_w5020_,
		_w5021_
	);
	LUT4 #(
		.INIT('h3111)
	) name4559 (
		_w1731_,
		_w5010_,
		_w5018_,
		_w5021_,
		_w5022_
	);
	LUT3 #(
		.INIT('hce)
	) name4560 (
		\P1_state_reg[0]/NET0131 ,
		_w5009_,
		_w5022_,
		_w5023_
	);
	LUT2 #(
		.INIT('h2)
	) name4561 (
		\P1_reg1_reg[10]/NET0131 ,
		_w2462_,
		_w5024_
	);
	LUT4 #(
		.INIT('h2000)
	) name4562 (
		\P1_reg1_reg[10]/NET0131 ,
		_w1723_,
		_w1727_,
		_w1730_,
		_w5025_
	);
	LUT4 #(
		.INIT('hddd1)
	) name4563 (
		\P1_reg1_reg[10]/NET0131 ,
		_w2520_,
		_w4217_,
		_w4218_,
		_w5026_
	);
	LUT2 #(
		.INIT('h2)
	) name4564 (
		_w2424_,
		_w5026_,
		_w5027_
	);
	LUT4 #(
		.INIT('h1dd1)
	) name4565 (
		\P1_reg1_reg[10]/NET0131 ,
		_w2520_,
		_w2953_,
		_w3176_,
		_w5028_
	);
	LUT2 #(
		.INIT('h2)
	) name4566 (
		_w2292_,
		_w5028_,
		_w5029_
	);
	LUT4 #(
		.INIT('hd11d)
	) name4567 (
		\P1_reg1_reg[10]/NET0131 ,
		_w2520_,
		_w2935_,
		_w3176_,
		_w5030_
	);
	LUT4 #(
		.INIT('hc808)
	) name4568 (
		\P1_reg1_reg[10]/NET0131 ,
		_w2447_,
		_w2520_,
		_w4224_,
		_w5031_
	);
	LUT2 #(
		.INIT('h8)
	) name4569 (
		_w2520_,
		_w4697_,
		_w5032_
	);
	LUT4 #(
		.INIT('h08aa)
	) name4570 (
		\P1_reg1_reg[10]/NET0131 ,
		_w2426_,
		_w2520_,
		_w2524_,
		_w5033_
	);
	LUT2 #(
		.INIT('h1)
	) name4571 (
		_w5032_,
		_w5033_,
		_w5034_
	);
	LUT2 #(
		.INIT('h4)
	) name4572 (
		_w5031_,
		_w5034_,
		_w5035_
	);
	LUT3 #(
		.INIT('hd0)
	) name4573 (
		_w2388_,
		_w5030_,
		_w5035_,
		_w5036_
	);
	LUT4 #(
		.INIT('ha8aa)
	) name4574 (
		_w1731_,
		_w5027_,
		_w5029_,
		_w5036_,
		_w5037_
	);
	LUT4 #(
		.INIT('heeec)
	) name4575 (
		\P1_state_reg[0]/NET0131 ,
		_w5024_,
		_w5025_,
		_w5037_,
		_w5038_
	);
	LUT2 #(
		.INIT('h2)
	) name4576 (
		\P1_reg1_reg[13]/NET0131 ,
		_w2462_,
		_w5039_
	);
	LUT4 #(
		.INIT('h2000)
	) name4577 (
		\P1_reg1_reg[13]/NET0131 ,
		_w1723_,
		_w1727_,
		_w1730_,
		_w5040_
	);
	LUT2 #(
		.INIT('h2)
	) name4578 (
		\P1_reg1_reg[13]/NET0131 ,
		_w2520_,
		_w5041_
	);
	LUT4 #(
		.INIT('h20d0)
	) name4579 (
		_w2049_,
		_w2153_,
		_w2520_,
		_w3192_,
		_w5042_
	);
	LUT2 #(
		.INIT('h2)
	) name4580 (
		\P1_reg1_reg[13]/NET0131 ,
		_w2525_,
		_w5043_
	);
	LUT4 #(
		.INIT('h0057)
	) name4581 (
		_w2520_,
		_w4240_,
		_w4708_,
		_w5043_,
		_w5044_
	);
	LUT4 #(
		.INIT('h5700)
	) name4582 (
		_w2292_,
		_w5041_,
		_w5042_,
		_w5044_,
		_w5045_
	);
	LUT4 #(
		.INIT('h7020)
	) name4583 (
		_w1747_,
		_w2020_,
		_w2520_,
		_w4237_,
		_w5046_
	);
	LUT3 #(
		.INIT('ha8)
	) name4584 (
		_w2424_,
		_w5041_,
		_w5046_,
		_w5047_
	);
	LUT4 #(
		.INIT('h08c8)
	) name4585 (
		\P1_reg1_reg[13]/NET0131 ,
		_w2388_,
		_w2520_,
		_w4245_,
		_w5048_
	);
	LUT4 #(
		.INIT('ha8aa)
	) name4586 (
		_w1731_,
		_w5047_,
		_w5048_,
		_w5045_,
		_w5049_
	);
	LUT4 #(
		.INIT('heeec)
	) name4587 (
		\P1_state_reg[0]/NET0131 ,
		_w5039_,
		_w5040_,
		_w5049_,
		_w5050_
	);
	LUT4 #(
		.INIT('h08c8)
	) name4588 (
		\P1_reg1_reg[23]/NET0131 ,
		_w2292_,
		_w2520_,
		_w4362_,
		_w5051_
	);
	LUT4 #(
		.INIT('h08c8)
	) name4589 (
		\P1_reg1_reg[23]/NET0131 ,
		_w2388_,
		_w2520_,
		_w4368_,
		_w5052_
	);
	LUT4 #(
		.INIT('hc808)
	) name4590 (
		\P1_reg1_reg[23]/NET0131 ,
		_w2424_,
		_w2520_,
		_w4371_,
		_w5053_
	);
	LUT4 #(
		.INIT('h08aa)
	) name4591 (
		\P1_reg1_reg[23]/NET0131 ,
		_w2452_,
		_w2520_,
		_w2524_,
		_w5054_
	);
	LUT3 #(
		.INIT('h0d)
	) name4592 (
		_w2520_,
		_w4374_,
		_w5054_,
		_w5055_
	);
	LUT2 #(
		.INIT('h4)
	) name4593 (
		_w5053_,
		_w5055_,
		_w5056_
	);
	LUT4 #(
		.INIT('ha8aa)
	) name4594 (
		_w1731_,
		_w5051_,
		_w5052_,
		_w5056_,
		_w5057_
	);
	LUT4 #(
		.INIT('h2000)
	) name4595 (
		\P1_reg1_reg[23]/NET0131 ,
		_w1723_,
		_w1727_,
		_w1730_,
		_w5058_
	);
	LUT2 #(
		.INIT('h2)
	) name4596 (
		\P1_reg1_reg[23]/NET0131 ,
		_w2462_,
		_w5059_
	);
	LUT4 #(
		.INIT('hffa8)
	) name4597 (
		\P1_state_reg[0]/NET0131 ,
		_w5057_,
		_w5058_,
		_w5059_,
		_w5060_
	);
	LUT4 #(
		.INIT('hd070)
	) name4598 (
		\P1_state_reg[0]/NET0131 ,
		\P2_IR_reg[23]/NET0131 ,
		\P2_reg0_reg[10]/NET0131 ,
		_w1188_,
		_w5061_
	);
	LUT4 #(
		.INIT('h2000)
	) name4599 (
		\P2_reg0_reg[10]/NET0131 ,
		_w1189_,
		_w1352_,
		_w1356_,
		_w5062_
	);
	LUT4 #(
		.INIT('h02aa)
	) name4600 (
		\P2_reg0_reg[10]/NET0131 ,
		_w1361_,
		_w1363_,
		_w1368_,
		_w5063_
	);
	LUT4 #(
		.INIT('h08c8)
	) name4601 (
		\P2_reg0_reg[10]/NET0131 ,
		_w1191_,
		_w1369_,
		_w4258_,
		_w5064_
	);
	LUT4 #(
		.INIT('haaa8)
	) name4602 (
		\P2_reg0_reg[10]/NET0131 ,
		_w1361_,
		_w1363_,
		_w1368_,
		_w5065_
	);
	LUT2 #(
		.INIT('h8)
	) name4603 (
		_w1411_,
		_w4802_,
		_w5066_
	);
	LUT3 #(
		.INIT('ha2)
	) name4604 (
		\P2_reg0_reg[10]/NET0131 ,
		_w1684_,
		_w1685_,
		_w5067_
	);
	LUT2 #(
		.INIT('h1)
	) name4605 (
		_w5066_,
		_w5067_,
		_w5068_
	);
	LUT4 #(
		.INIT('hab00)
	) name4606 (
		_w1496_,
		_w4268_,
		_w5065_,
		_w5068_,
		_w5069_
	);
	LUT4 #(
		.INIT('h8848)
	) name4607 (
		_w1317_,
		_w1411_,
		_w2553_,
		_w2555_,
		_w5070_
	);
	LUT3 #(
		.INIT('h54)
	) name4608 (
		_w1409_,
		_w5065_,
		_w5070_,
		_w5071_
	);
	LUT3 #(
		.INIT('ha8)
	) name4609 (
		_w1447_,
		_w4266_,
		_w5063_,
		_w5072_
	);
	LUT4 #(
		.INIT('h0100)
	) name4610 (
		_w5071_,
		_w5072_,
		_w5064_,
		_w5069_,
		_w5073_
	);
	LUT4 #(
		.INIT('ha0a8)
	) name4611 (
		\P1_state_reg[0]/NET0131 ,
		_w1359_,
		_w5062_,
		_w5073_,
		_w5074_
	);
	LUT2 #(
		.INIT('he)
	) name4612 (
		_w5061_,
		_w5074_,
		_w5075_
	);
	LUT4 #(
		.INIT('hd070)
	) name4613 (
		\P1_state_reg[0]/NET0131 ,
		\P2_IR_reg[23]/NET0131 ,
		\P2_reg0_reg[12]/NET0131 ,
		_w1188_,
		_w5076_
	);
	LUT4 #(
		.INIT('h2000)
	) name4614 (
		\P2_reg0_reg[12]/NET0131 ,
		_w1189_,
		_w1352_,
		_w1356_,
		_w5077_
	);
	LUT4 #(
		.INIT('h0232)
	) name4615 (
		\P2_reg0_reg[12]/NET0131 ,
		_w1409_,
		_w1411_,
		_w4277_,
		_w5078_
	);
	LUT4 #(
		.INIT('h111d)
	) name4616 (
		\P2_reg0_reg[12]/NET0131 ,
		_w1369_,
		_w4280_,
		_w4281_,
		_w5079_
	);
	LUT2 #(
		.INIT('h8)
	) name4617 (
		_w1411_,
		_w4818_,
		_w5080_
	);
	LUT3 #(
		.INIT('ha2)
	) name4618 (
		\P2_reg0_reg[12]/NET0131 ,
		_w1684_,
		_w1685_,
		_w5081_
	);
	LUT2 #(
		.INIT('h1)
	) name4619 (
		_w5080_,
		_w5081_,
		_w5082_
	);
	LUT3 #(
		.INIT('hd0)
	) name4620 (
		_w1191_,
		_w5079_,
		_w5082_,
		_w5083_
	);
	LUT4 #(
		.INIT('h0e02)
	) name4621 (
		\P2_reg0_reg[12]/NET0131 ,
		_w1411_,
		_w1496_,
		_w4287_,
		_w5084_
	);
	LUT4 #(
		.INIT('he020)
	) name4622 (
		\P2_reg0_reg[12]/NET0131 ,
		_w1369_,
		_w1447_,
		_w4287_,
		_w5085_
	);
	LUT4 #(
		.INIT('h0100)
	) name4623 (
		_w5078_,
		_w5084_,
		_w5085_,
		_w5083_,
		_w5086_
	);
	LUT4 #(
		.INIT('ha0a8)
	) name4624 (
		\P1_state_reg[0]/NET0131 ,
		_w1359_,
		_w5077_,
		_w5086_,
		_w5087_
	);
	LUT2 #(
		.INIT('he)
	) name4625 (
		_w5076_,
		_w5087_,
		_w5088_
	);
	LUT4 #(
		.INIT('hd070)
	) name4626 (
		\P1_state_reg[0]/NET0131 ,
		\P2_IR_reg[23]/NET0131 ,
		\P2_reg0_reg[13]/NET0131 ,
		_w1188_,
		_w5089_
	);
	LUT4 #(
		.INIT('h2000)
	) name4627 (
		\P2_reg0_reg[13]/NET0131 ,
		_w1189_,
		_w1352_,
		_w1356_,
		_w5090_
	);
	LUT4 #(
		.INIT('hc535)
	) name4628 (
		\P2_reg0_reg[13]/NET0131 ,
		_w1299_,
		_w1411_,
		_w1699_,
		_w5091_
	);
	LUT4 #(
		.INIT('h08c8)
	) name4629 (
		\P2_reg0_reg[13]/NET0131 ,
		_w1191_,
		_w1369_,
		_w4301_,
		_w5092_
	);
	LUT2 #(
		.INIT('h8)
	) name4630 (
		_w1411_,
		_w4832_,
		_w5093_
	);
	LUT3 #(
		.INIT('ha2)
	) name4631 (
		\P2_reg0_reg[13]/NET0131 ,
		_w1684_,
		_w1685_,
		_w5094_
	);
	LUT2 #(
		.INIT('h1)
	) name4632 (
		_w5093_,
		_w5094_,
		_w5095_
	);
	LUT4 #(
		.INIT('h0e00)
	) name4633 (
		_w1496_,
		_w5091_,
		_w5092_,
		_w5095_,
		_w5096_
	);
	LUT4 #(
		.INIT('hc535)
	) name4634 (
		\P2_reg0_reg[13]/NET0131 ,
		_w1299_,
		_w1369_,
		_w1699_,
		_w5097_
	);
	LUT4 #(
		.INIT('h3202)
	) name4635 (
		\P2_reg0_reg[13]/NET0131 ,
		_w1409_,
		_w1411_,
		_w4309_,
		_w5098_
	);
	LUT3 #(
		.INIT('h0d)
	) name4636 (
		_w1447_,
		_w5097_,
		_w5098_,
		_w5099_
	);
	LUT4 #(
		.INIT('h3111)
	) name4637 (
		_w1359_,
		_w5090_,
		_w5096_,
		_w5099_,
		_w5100_
	);
	LUT3 #(
		.INIT('hce)
	) name4638 (
		\P1_state_reg[0]/NET0131 ,
		_w5089_,
		_w5100_,
		_w5101_
	);
	LUT2 #(
		.INIT('h2)
	) name4639 (
		\P1_reg1_reg[30]/NET0131 ,
		_w2462_,
		_w5102_
	);
	LUT4 #(
		.INIT('h2000)
	) name4640 (
		\P1_reg1_reg[30]/NET0131 ,
		_w1723_,
		_w1727_,
		_w1730_,
		_w5103_
	);
	LUT4 #(
		.INIT('hc808)
	) name4641 (
		\P1_reg1_reg[30]/NET0131 ,
		_w2447_,
		_w2520_,
		_w4862_,
		_w5104_
	);
	LUT4 #(
		.INIT('hf5c5)
	) name4642 (
		\P1_reg1_reg[30]/NET0131 ,
		_w1748_,
		_w2520_,
		_w3134_,
		_w5105_
	);
	LUT4 #(
		.INIT('h0a2a)
	) name4643 (
		\P1_reg1_reg[30]/NET0131 ,
		_w2520_,
		_w2524_,
		_w3574_,
		_w5106_
	);
	LUT3 #(
		.INIT('h0d)
	) name4644 (
		_w2426_,
		_w5105_,
		_w5106_,
		_w5107_
	);
	LUT4 #(
		.INIT('ha8aa)
	) name4645 (
		_w1731_,
		_w3969_,
		_w5104_,
		_w5107_,
		_w5108_
	);
	LUT4 #(
		.INIT('heeec)
	) name4646 (
		\P1_state_reg[0]/NET0131 ,
		_w5102_,
		_w5103_,
		_w5108_,
		_w5109_
	);
	LUT4 #(
		.INIT('h4000)
	) name4647 (
		_w1723_,
		_w1727_,
		_w1730_,
		_w2050_,
		_w5110_
	);
	LUT2 #(
		.INIT('h2)
	) name4648 (
		_w2050_,
		_w2644_,
		_w5111_
	);
	LUT4 #(
		.INIT('h4150)
	) name4649 (
		_w1747_,
		_w2053_,
		_w2138_,
		_w2400_,
		_w5112_
	);
	LUT3 #(
		.INIT('h80)
	) name4650 (
		_w489_,
		_w491_,
		_w1747_,
		_w5113_
	);
	LUT4 #(
		.INIT('h3331)
	) name4651 (
		_w2644_,
		_w5111_,
		_w5112_,
		_w5113_,
		_w5114_
	);
	LUT2 #(
		.INIT('h2)
	) name4652 (
		_w2424_,
		_w5114_,
		_w5115_
	);
	LUT4 #(
		.INIT('h0df2)
	) name4653 (
		_w2310_,
		_w2792_,
		_w2793_,
		_w3178_,
		_w5116_
	);
	LUT4 #(
		.INIT('hc808)
	) name4654 (
		_w2050_,
		_w2388_,
		_w2644_,
		_w5116_,
		_w5117_
	);
	LUT4 #(
		.INIT('hd02f)
	) name4655 (
		_w2073_,
		_w2091_,
		_w2747_,
		_w3178_,
		_w5118_
	);
	LUT4 #(
		.INIT('h08c8)
	) name4656 (
		_w2050_,
		_w2292_,
		_w2644_,
		_w5118_,
		_w5119_
	);
	LUT4 #(
		.INIT('hc355)
	) name4657 (
		_w2050_,
		_w2057_,
		_w2429_,
		_w2644_,
		_w5120_
	);
	LUT4 #(
		.INIT('h5450)
	) name4658 (
		_w2057_,
		_w2426_,
		_w2454_,
		_w2644_,
		_w5121_
	);
	LUT4 #(
		.INIT('ha0a8)
	) name4659 (
		_w2050_,
		_w2426_,
		_w2450_,
		_w2644_,
		_w5122_
	);
	LUT4 #(
		.INIT('h0031)
	) name4660 (
		_w2447_,
		_w5121_,
		_w5120_,
		_w5122_,
		_w5123_
	);
	LUT3 #(
		.INIT('h10)
	) name4661 (
		_w5119_,
		_w5117_,
		_w5123_,
		_w5124_
	);
	LUT4 #(
		.INIT('h1311)
	) name4662 (
		_w1731_,
		_w5110_,
		_w5115_,
		_w5124_,
		_w5125_
	);
	LUT2 #(
		.INIT('h2)
	) name4663 (
		\P1_reg3_reg[4]/NET0131 ,
		\P1_state_reg[0]/NET0131 ,
		_w5126_
	);
	LUT3 #(
		.INIT('h07)
	) name4664 (
		_w2050_,
		_w2695_,
		_w5126_,
		_w5127_
	);
	LUT3 #(
		.INIT('h2f)
	) name4665 (
		\P1_state_reg[0]/NET0131 ,
		_w5125_,
		_w5127_,
		_w5128_
	);
	LUT2 #(
		.INIT('h2)
	) name4666 (
		_w2136_,
		_w2644_,
		_w5129_
	);
	LUT4 #(
		.INIT('h3633)
	) name4667 (
		_w2053_,
		_w2128_,
		_w2138_,
		_w2400_,
		_w5130_
	);
	LUT4 #(
		.INIT('h7020)
	) name4668 (
		_w1747_,
		_w2053_,
		_w2644_,
		_w5130_,
		_w5131_
	);
	LUT3 #(
		.INIT('ha8)
	) name4669 (
		_w2424_,
		_w5129_,
		_w5131_,
		_w5132_
	);
	LUT4 #(
		.INIT('h00b7)
	) name4670 (
		_w2096_,
		_w2644_,
		_w3187_,
		_w5129_,
		_w5133_
	);
	LUT2 #(
		.INIT('h2)
	) name4671 (
		_w2292_,
		_w5133_,
		_w5134_
	);
	LUT4 #(
		.INIT('h0075)
	) name4672 (
		_w2304_,
		_w2307_,
		_w2310_,
		_w2312_,
		_w5135_
	);
	LUT4 #(
		.INIT('h070d)
	) name4673 (
		_w2644_,
		_w3187_,
		_w5129_,
		_w5135_,
		_w5136_
	);
	LUT4 #(
		.INIT('h6c00)
	) name4674 (
		_w2057_,
		_w2134_,
		_w2429_,
		_w2447_,
		_w5137_
	);
	LUT2 #(
		.INIT('h8)
	) name4675 (
		_w2644_,
		_w5137_,
		_w5138_
	);
	LUT4 #(
		.INIT('h5450)
	) name4676 (
		_w2134_,
		_w2426_,
		_w2454_,
		_w2644_,
		_w5139_
	);
	LUT3 #(
		.INIT('h0d)
	) name4677 (
		_w2136_,
		_w2690_,
		_w5139_,
		_w5140_
	);
	LUT2 #(
		.INIT('h4)
	) name4678 (
		_w5138_,
		_w5140_,
		_w5141_
	);
	LUT3 #(
		.INIT('hd0)
	) name4679 (
		_w2388_,
		_w5136_,
		_w5141_,
		_w5142_
	);
	LUT4 #(
		.INIT('ha8aa)
	) name4680 (
		_w1731_,
		_w5132_,
		_w5134_,
		_w5142_,
		_w5143_
	);
	LUT4 #(
		.INIT('h4000)
	) name4681 (
		_w1723_,
		_w1727_,
		_w1730_,
		_w2136_,
		_w5144_
	);
	LUT2 #(
		.INIT('h2)
	) name4682 (
		\P1_reg3_reg[5]/NET0131 ,
		\P1_state_reg[0]/NET0131 ,
		_w5145_
	);
	LUT3 #(
		.INIT('h07)
	) name4683 (
		_w2136_,
		_w2695_,
		_w5145_,
		_w5146_
	);
	LUT4 #(
		.INIT('ha8ff)
	) name4684 (
		\P1_state_reg[0]/NET0131 ,
		_w5143_,
		_w5144_,
		_w5146_,
		_w5147_
	);
	LUT4 #(
		.INIT('h1000)
	) name4685 (
		_w765_,
		_w1189_,
		_w1352_,
		_w1356_,
		_w5148_
	);
	LUT4 #(
		.INIT('h5554)
	) name4686 (
		_w765_,
		_w1361_,
		_w1363_,
		_w1368_,
		_w5149_
	);
	LUT2 #(
		.INIT('h1)
	) name4687 (
		_w781_,
		_w1435_,
		_w5150_
	);
	LUT3 #(
		.INIT('h10)
	) name4688 (
		_w792_,
		_w803_,
		_w1414_,
		_w5151_
	);
	LUT4 #(
		.INIT('h0100)
	) name4689 (
		_w781_,
		_w792_,
		_w803_,
		_w1414_,
		_w5152_
	);
	LUT4 #(
		.INIT('hbf00)
	) name4690 (
		_w803_,
		_w1414_,
		_w1415_,
		_w1435_,
		_w5153_
	);
	LUT4 #(
		.INIT('h7500)
	) name4691 (
		_w747_,
		_w770_,
		_w5152_,
		_w5153_,
		_w5154_
	);
	LUT4 #(
		.INIT('h1113)
	) name4692 (
		_w1411_,
		_w5149_,
		_w5150_,
		_w5154_,
		_w5155_
	);
	LUT2 #(
		.INIT('h2)
	) name4693 (
		_w1191_,
		_w5155_,
		_w5156_
	);
	LUT4 #(
		.INIT('h0155)
	) name4694 (
		_w765_,
		_w1361_,
		_w1363_,
		_w1368_,
		_w5157_
	);
	LUT4 #(
		.INIT('hc090)
	) name4695 (
		_w786_,
		_w1306_,
		_w1369_,
		_w1375_,
		_w5158_
	);
	LUT3 #(
		.INIT('h54)
	) name4696 (
		_w1409_,
		_w5157_,
		_w5158_,
		_w5159_
	);
	LUT4 #(
		.INIT('h8884)
	) name4697 (
		_w1306_,
		_w1369_,
		_w1454_,
		_w1455_,
		_w5160_
	);
	LUT3 #(
		.INIT('h54)
	) name4698 (
		_w1496_,
		_w5157_,
		_w5160_,
		_w5161_
	);
	LUT4 #(
		.INIT('h8884)
	) name4699 (
		_w1306_,
		_w1411_,
		_w1454_,
		_w1455_,
		_w5162_
	);
	LUT3 #(
		.INIT('h04)
	) name4700 (
		_w774_,
		_w1232_,
		_w1439_,
		_w5163_
	);
	LUT3 #(
		.INIT('h54)
	) name4701 (
		_w765_,
		_w1441_,
		_w1443_,
		_w5164_
	);
	LUT2 #(
		.INIT('h1)
	) name4702 (
		_w5163_,
		_w5164_,
		_w5165_
	);
	LUT4 #(
		.INIT('h5700)
	) name4703 (
		_w1447_,
		_w5149_,
		_w5162_,
		_w5165_,
		_w5166_
	);
	LUT3 #(
		.INIT('h10)
	) name4704 (
		_w5159_,
		_w5161_,
		_w5166_,
		_w5167_
	);
	LUT4 #(
		.INIT('h1311)
	) name4705 (
		_w1359_,
		_w5148_,
		_w5156_,
		_w5167_,
		_w5168_
	);
	LUT2 #(
		.INIT('h4)
	) name4706 (
		\P1_state_reg[0]/NET0131 ,
		\P2_reg3_reg[5]/NET0131 ,
		_w5169_
	);
	LUT4 #(
		.INIT('h0802)
	) name4707 (
		\P1_state_reg[0]/NET0131 ,
		\P2_IR_reg[23]/NET0131 ,
		_w765_,
		_w1188_,
		_w5170_
	);
	LUT2 #(
		.INIT('h1)
	) name4708 (
		_w5169_,
		_w5170_,
		_w5171_
	);
	LUT3 #(
		.INIT('h2f)
	) name4709 (
		\P1_state_reg[0]/NET0131 ,
		_w5168_,
		_w5171_,
		_w5172_
	);
	LUT4 #(
		.INIT('h1000)
	) name4710 (
		_w744_,
		_w1189_,
		_w1352_,
		_w1356_,
		_w5173_
	);
	LUT4 #(
		.INIT('h0155)
	) name4711 (
		_w744_,
		_w1361_,
		_w1363_,
		_w1368_,
		_w5174_
	);
	LUT4 #(
		.INIT('h4844)
	) name4712 (
		_w1322_,
		_w1369_,
		_w1534_,
		_w1535_,
		_w5175_
	);
	LUT3 #(
		.INIT('h04)
	) name4713 (
		_w752_,
		_w1232_,
		_w1439_,
		_w5176_
	);
	LUT3 #(
		.INIT('h54)
	) name4714 (
		_w744_,
		_w1441_,
		_w1443_,
		_w5177_
	);
	LUT2 #(
		.INIT('h1)
	) name4715 (
		_w5176_,
		_w5177_,
		_w5178_
	);
	LUT4 #(
		.INIT('hab00)
	) name4716 (
		_w1496_,
		_w5174_,
		_w5175_,
		_w5178_,
		_w5179_
	);
	LUT4 #(
		.INIT('he100)
	) name4717 (
		_w1212_,
		_w1213_,
		_w1322_,
		_w1369_,
		_w5180_
	);
	LUT3 #(
		.INIT('h54)
	) name4718 (
		_w1409_,
		_w5174_,
		_w5180_,
		_w5181_
	);
	LUT4 #(
		.INIT('h5554)
	) name4719 (
		_w744_,
		_w1361_,
		_w1363_,
		_w1368_,
		_w5182_
	);
	LUT4 #(
		.INIT('h4844)
	) name4720 (
		_w1322_,
		_w1411_,
		_w1534_,
		_w1535_,
		_w5183_
	);
	LUT3 #(
		.INIT('ha8)
	) name4721 (
		_w1447_,
		_w5182_,
		_w5183_,
		_w5184_
	);
	LUT4 #(
		.INIT('h1000)
	) name4722 (
		_w759_,
		_w803_,
		_w1414_,
		_w1415_,
		_w5185_
	);
	LUT2 #(
		.INIT('h1)
	) name4723 (
		_w770_,
		_w1435_,
		_w5186_
	);
	LUT4 #(
		.INIT('h006f)
	) name4724 (
		_w759_,
		_w1416_,
		_w1435_,
		_w5186_,
		_w5187_
	);
	LUT4 #(
		.INIT('h04c4)
	) name4725 (
		_w744_,
		_w1191_,
		_w1411_,
		_w5187_,
		_w5188_
	);
	LUT4 #(
		.INIT('h0100)
	) name4726 (
		_w5184_,
		_w5188_,
		_w5181_,
		_w5179_,
		_w5189_
	);
	LUT4 #(
		.INIT('ha0a8)
	) name4727 (
		\P1_state_reg[0]/NET0131 ,
		_w1359_,
		_w5173_,
		_w5189_,
		_w5190_
	);
	LUT2 #(
		.INIT('h4)
	) name4728 (
		\P1_state_reg[0]/NET0131 ,
		\P2_reg3_reg[6]/NET0131 ,
		_w5191_
	);
	LUT4 #(
		.INIT('h0802)
	) name4729 (
		\P1_state_reg[0]/NET0131 ,
		\P2_IR_reg[23]/NET0131 ,
		_w744_,
		_w1188_,
		_w5192_
	);
	LUT2 #(
		.INIT('h1)
	) name4730 (
		_w5191_,
		_w5192_,
		_w5193_
	);
	LUT2 #(
		.INIT('hb)
	) name4731 (
		_w5190_,
		_w5193_,
		_w5194_
	);
	LUT4 #(
		.INIT('h1000)
	) name4732 (
		_w755_,
		_w1189_,
		_w1352_,
		_w1356_,
		_w5195_
	);
	LUT4 #(
		.INIT('h0155)
	) name4733 (
		_w755_,
		_w1361_,
		_w1363_,
		_w1368_,
		_w5196_
	);
	LUT4 #(
		.INIT('h00b7)
	) name4734 (
		_w1303_,
		_w1369_,
		_w1458_,
		_w5196_,
		_w5197_
	);
	LUT2 #(
		.INIT('h1)
	) name4735 (
		_w1496_,
		_w5197_,
		_w5198_
	);
	LUT4 #(
		.INIT('h5554)
	) name4736 (
		_w755_,
		_w1361_,
		_w1363_,
		_w1368_,
		_w5199_
	);
	LUT2 #(
		.INIT('h1)
	) name4737 (
		_w747_,
		_w1435_,
		_w5200_
	);
	LUT4 #(
		.INIT('h3010)
	) name4738 (
		_w726_,
		_w1418_,
		_w1435_,
		_w5185_,
		_w5201_
	);
	LUT4 #(
		.INIT('h1113)
	) name4739 (
		_w1411_,
		_w5199_,
		_w5200_,
		_w5201_,
		_w5202_
	);
	LUT3 #(
		.INIT('h04)
	) name4740 (
		_w763_,
		_w1232_,
		_w1439_,
		_w5203_
	);
	LUT3 #(
		.INIT('h54)
	) name4741 (
		_w755_,
		_w1441_,
		_w1443_,
		_w5204_
	);
	LUT2 #(
		.INIT('h1)
	) name4742 (
		_w5203_,
		_w5204_,
		_w5205_
	);
	LUT3 #(
		.INIT('hd0)
	) name4743 (
		_w1191_,
		_w5202_,
		_w5205_,
		_w5206_
	);
	LUT4 #(
		.INIT('h00b7)
	) name4744 (
		_w1303_,
		_w1411_,
		_w1458_,
		_w5199_,
		_w5207_
	);
	LUT4 #(
		.INIT('h6566)
	) name4745 (
		_w1303_,
		_w1374_,
		_w1375_,
		_w1376_,
		_w5208_
	);
	LUT4 #(
		.INIT('h0d01)
	) name4746 (
		_w755_,
		_w1369_,
		_w1409_,
		_w5208_,
		_w5209_
	);
	LUT3 #(
		.INIT('h0d)
	) name4747 (
		_w1447_,
		_w5207_,
		_w5209_,
		_w5210_
	);
	LUT4 #(
		.INIT('h8aaa)
	) name4748 (
		_w1359_,
		_w5198_,
		_w5206_,
		_w5210_,
		_w5211_
	);
	LUT2 #(
		.INIT('h4)
	) name4749 (
		\P1_state_reg[0]/NET0131 ,
		\P2_reg3_reg[7]/NET0131 ,
		_w5212_
	);
	LUT4 #(
		.INIT('h0802)
	) name4750 (
		\P1_state_reg[0]/NET0131 ,
		\P2_IR_reg[23]/NET0131 ,
		_w755_,
		_w1188_,
		_w5213_
	);
	LUT2 #(
		.INIT('h1)
	) name4751 (
		_w5212_,
		_w5213_,
		_w5214_
	);
	LUT4 #(
		.INIT('ha8ff)
	) name4752 (
		\P1_state_reg[0]/NET0131 ,
		_w5195_,
		_w5211_,
		_w5214_,
		_w5215_
	);
	LUT2 #(
		.INIT('h2)
	) name4753 (
		\P1_reg1_reg[4]/NET0131 ,
		_w2462_,
		_w5216_
	);
	LUT4 #(
		.INIT('h2000)
	) name4754 (
		\P1_reg1_reg[4]/NET0131 ,
		_w1723_,
		_w1727_,
		_w1730_,
		_w5217_
	);
	LUT4 #(
		.INIT('hddd1)
	) name4755 (
		\P1_reg1_reg[4]/NET0131 ,
		_w2520_,
		_w5112_,
		_w5113_,
		_w5218_
	);
	LUT2 #(
		.INIT('h2)
	) name4756 (
		_w2424_,
		_w5218_,
		_w5219_
	);
	LUT4 #(
		.INIT('hc808)
	) name4757 (
		\P1_reg1_reg[4]/NET0131 ,
		_w2388_,
		_w2520_,
		_w5116_,
		_w5220_
	);
	LUT4 #(
		.INIT('h08c8)
	) name4758 (
		\P1_reg1_reg[4]/NET0131 ,
		_w2292_,
		_w2520_,
		_w5118_,
		_w5221_
	);
	LUT4 #(
		.INIT('hc355)
	) name4759 (
		\P1_reg1_reg[4]/NET0131 ,
		_w2057_,
		_w2429_,
		_w2520_,
		_w5222_
	);
	LUT2 #(
		.INIT('h4)
	) name4760 (
		_w2057_,
		_w2426_,
		_w5223_
	);
	LUT2 #(
		.INIT('h8)
	) name4761 (
		_w2520_,
		_w5223_,
		_w5224_
	);
	LUT4 #(
		.INIT('h08aa)
	) name4762 (
		\P1_reg1_reg[4]/NET0131 ,
		_w2426_,
		_w2520_,
		_w2524_,
		_w5225_
	);
	LUT4 #(
		.INIT('h0031)
	) name4763 (
		_w2447_,
		_w5224_,
		_w5222_,
		_w5225_,
		_w5226_
	);
	LUT3 #(
		.INIT('h10)
	) name4764 (
		_w5221_,
		_w5220_,
		_w5226_,
		_w5227_
	);
	LUT4 #(
		.INIT('h1311)
	) name4765 (
		_w1731_,
		_w5217_,
		_w5219_,
		_w5227_,
		_w5228_
	);
	LUT3 #(
		.INIT('hce)
	) name4766 (
		\P1_state_reg[0]/NET0131 ,
		_w5216_,
		_w5228_,
		_w5229_
	);
	LUT2 #(
		.INIT('h2)
	) name4767 (
		\P1_reg0_reg[4]/NET0131 ,
		_w2462_,
		_w5230_
	);
	LUT4 #(
		.INIT('h2000)
	) name4768 (
		\P1_reg0_reg[4]/NET0131 ,
		_w1723_,
		_w1727_,
		_w1730_,
		_w5231_
	);
	LUT4 #(
		.INIT('hddd1)
	) name4769 (
		\P1_reg0_reg[4]/NET0131 ,
		_w2883_,
		_w5112_,
		_w5113_,
		_w5232_
	);
	LUT2 #(
		.INIT('h2)
	) name4770 (
		_w2424_,
		_w5232_,
		_w5233_
	);
	LUT4 #(
		.INIT('hc808)
	) name4771 (
		\P1_reg0_reg[4]/NET0131 ,
		_w2388_,
		_w2883_,
		_w5116_,
		_w5234_
	);
	LUT4 #(
		.INIT('h08c8)
	) name4772 (
		\P1_reg0_reg[4]/NET0131 ,
		_w2292_,
		_w2883_,
		_w5118_,
		_w5235_
	);
	LUT4 #(
		.INIT('hc355)
	) name4773 (
		\P1_reg0_reg[4]/NET0131 ,
		_w2057_,
		_w2429_,
		_w2883_,
		_w5236_
	);
	LUT2 #(
		.INIT('h8)
	) name4774 (
		_w2883_,
		_w5223_,
		_w5237_
	);
	LUT4 #(
		.INIT('h0a8a)
	) name4775 (
		\P1_reg0_reg[4]/NET0131 ,
		_w2426_,
		_w2524_,
		_w2883_,
		_w5238_
	);
	LUT4 #(
		.INIT('h0031)
	) name4776 (
		_w2447_,
		_w5237_,
		_w5236_,
		_w5238_,
		_w5239_
	);
	LUT3 #(
		.INIT('h10)
	) name4777 (
		_w5235_,
		_w5234_,
		_w5239_,
		_w5240_
	);
	LUT4 #(
		.INIT('h1311)
	) name4778 (
		_w1731_,
		_w5231_,
		_w5233_,
		_w5240_,
		_w5241_
	);
	LUT3 #(
		.INIT('hce)
	) name4779 (
		\P1_state_reg[0]/NET0131 ,
		_w5230_,
		_w5241_,
		_w5242_
	);
	LUT2 #(
		.INIT('h1)
	) name4780 (
		\P1_reg2_reg[8]/NET0131 ,
		_w1741_,
		_w5243_
	);
	LUT4 #(
		.INIT('h0222)
	) name4781 (
		\P1_state_reg[0]/NET0131 ,
		_w1723_,
		_w1727_,
		_w1730_,
		_w5244_
	);
	LUT4 #(
		.INIT('h0d0f)
	) name4782 (
		_w4658_,
		_w4656_,
		_w5243_,
		_w5244_,
		_w5245_
	);
	LUT4 #(
		.INIT('had88)
	) name4783 (
		_w2104_,
		_w2426_,
		_w2431_,
		_w2447_,
		_w5246_
	);
	LUT4 #(
		.INIT('h0008)
	) name4784 (
		_w2106_,
		_w2284_,
		_w2288_,
		_w2291_,
		_w5247_
	);
	LUT4 #(
		.INIT('h2322)
	) name4785 (
		_w1741_,
		_w2450_,
		_w2452_,
		_w3574_,
		_w5248_
	);
	LUT3 #(
		.INIT('h31)
	) name4786 (
		\P1_reg2_reg[8]/NET0131 ,
		_w5247_,
		_w5248_,
		_w5249_
	);
	LUT3 #(
		.INIT('h70)
	) name4787 (
		_w1741_,
		_w5246_,
		_w5249_,
		_w5250_
	);
	LUT2 #(
		.INIT('h1)
	) name4788 (
		\P1_reg2_reg[8]/NET0131 ,
		_w5244_,
		_w5251_
	);
	LUT3 #(
		.INIT('h0b)
	) name4789 (
		_w5245_,
		_w5250_,
		_w5251_,
		_w5252_
	);
	LUT4 #(
		.INIT('hd070)
	) name4790 (
		\P1_state_reg[0]/NET0131 ,
		\P2_IR_reg[23]/NET0131 ,
		\P2_reg0_reg[15]/NET0131 ,
		_w1188_,
		_w5253_
	);
	LUT4 #(
		.INIT('h2000)
	) name4791 (
		\P2_reg0_reg[15]/NET0131 ,
		_w1189_,
		_w1352_,
		_w1356_,
		_w5254_
	);
	LUT4 #(
		.INIT('h02aa)
	) name4792 (
		\P2_reg0_reg[15]/NET0131 ,
		_w1361_,
		_w1363_,
		_w1368_,
		_w5255_
	);
	LUT3 #(
		.INIT('ha8)
	) name4793 (
		_w1447_,
		_w4641_,
		_w5255_,
		_w5256_
	);
	LUT4 #(
		.INIT('h111d)
	) name4794 (
		\P2_reg0_reg[15]/NET0131 ,
		_w1369_,
		_w4633_,
		_w4634_,
		_w5257_
	);
	LUT3 #(
		.INIT('h40)
	) name4795 (
		_w594_,
		_w1411_,
		_w1442_,
		_w5258_
	);
	LUT3 #(
		.INIT('ha2)
	) name4796 (
		\P2_reg0_reg[15]/NET0131 ,
		_w1684_,
		_w1685_,
		_w5259_
	);
	LUT2 #(
		.INIT('h1)
	) name4797 (
		_w5258_,
		_w5259_,
		_w5260_
	);
	LUT3 #(
		.INIT('hd0)
	) name4798 (
		_w1191_,
		_w5257_,
		_w5260_,
		_w5261_
	);
	LUT4 #(
		.INIT('haaa8)
	) name4799 (
		\P2_reg0_reg[15]/NET0131 ,
		_w1361_,
		_w1363_,
		_w1368_,
		_w5262_
	);
	LUT3 #(
		.INIT('h54)
	) name4800 (
		_w1496_,
		_w4631_,
		_w5262_,
		_w5263_
	);
	LUT4 #(
		.INIT('hc535)
	) name4801 (
		\P2_reg0_reg[15]/NET0131 ,
		_w1295_,
		_w1411_,
		_w3598_,
		_w5264_
	);
	LUT2 #(
		.INIT('h1)
	) name4802 (
		_w1409_,
		_w5264_,
		_w5265_
	);
	LUT4 #(
		.INIT('h0100)
	) name4803 (
		_w5256_,
		_w5263_,
		_w5265_,
		_w5261_,
		_w5266_
	);
	LUT4 #(
		.INIT('ha0a8)
	) name4804 (
		\P1_state_reg[0]/NET0131 ,
		_w1359_,
		_w5254_,
		_w5266_,
		_w5267_
	);
	LUT2 #(
		.INIT('he)
	) name4805 (
		_w5253_,
		_w5267_,
		_w5268_
	);
	LUT4 #(
		.INIT('h2022)
	) name4806 (
		_w2520_,
		_w4652_,
		_w4654_,
		_w4655_,
		_w5269_
	);
	LUT2 #(
		.INIT('h2)
	) name4807 (
		_w2424_,
		_w5269_,
		_w5270_
	);
	LUT2 #(
		.INIT('h2)
	) name4808 (
		_w2285_,
		_w2520_,
		_w5271_
	);
	LUT3 #(
		.INIT('h07)
	) name4809 (
		_w2520_,
		_w5246_,
		_w5271_,
		_w5272_
	);
	LUT3 #(
		.INIT('h80)
	) name4810 (
		_w4658_,
		_w5244_,
		_w5272_,
		_w5273_
	);
	LUT3 #(
		.INIT('h20)
	) name4811 (
		_w3744_,
		_w5270_,
		_w5273_,
		_w5274_
	);
	LUT2 #(
		.INIT('h8)
	) name4812 (
		_w2520_,
		_w5244_,
		_w5275_
	);
	LUT4 #(
		.INIT('h1055)
	) name4813 (
		\P1_reg1_reg[8]/NET0131 ,
		_w5270_,
		_w5273_,
		_w5275_,
		_w5276_
	);
	LUT2 #(
		.INIT('h1)
	) name4814 (
		_w5274_,
		_w5276_,
		_w5277_
	);
	LUT2 #(
		.INIT('h2)
	) name4815 (
		\P1_reg2_reg[11]/NET0131 ,
		_w2462_,
		_w5278_
	);
	LUT4 #(
		.INIT('h2000)
	) name4816 (
		\P1_reg2_reg[11]/NET0131 ,
		_w1723_,
		_w1727_,
		_w1730_,
		_w5279_
	);
	LUT2 #(
		.INIT('h2)
	) name4817 (
		\P1_reg2_reg[11]/NET0131 ,
		_w1741_,
		_w5280_
	);
	LUT4 #(
		.INIT('h8a20)
	) name4818 (
		_w1741_,
		_w2654_,
		_w2655_,
		_w3191_,
		_w5281_
	);
	LUT3 #(
		.INIT('ha8)
	) name4819 (
		_w2292_,
		_w5280_,
		_w5281_,
		_w5282_
	);
	LUT4 #(
		.INIT('h208a)
	) name4820 (
		_w1741_,
		_w2667_,
		_w2668_,
		_w3191_,
		_w5283_
	);
	LUT3 #(
		.INIT('ha8)
	) name4821 (
		_w2388_,
		_w5280_,
		_w5283_,
		_w5284_
	);
	LUT4 #(
		.INIT('hddd1)
	) name4822 (
		\P1_reg2_reg[11]/NET0131 ,
		_w1741_,
		_w4536_,
		_w4537_,
		_w5285_
	);
	LUT4 #(
		.INIT('h2300)
	) name4823 (
		_w1748_,
		_w2002_,
		_w2003_,
		_w2426_,
		_w5286_
	);
	LUT4 #(
		.INIT('h007b)
	) name4824 (
		_w2004_,
		_w2447_,
		_w3804_,
		_w5286_,
		_w5287_
	);
	LUT4 #(
		.INIT('h0008)
	) name4825 (
		_w2005_,
		_w2284_,
		_w2288_,
		_w2291_,
		_w5288_
	);
	LUT4 #(
		.INIT('ha2a0)
	) name4826 (
		\P1_reg2_reg[11]/NET0131 ,
		_w1741_,
		_w2450_,
		_w2452_,
		_w5289_
	);
	LUT2 #(
		.INIT('h1)
	) name4827 (
		_w5288_,
		_w5289_,
		_w5290_
	);
	LUT3 #(
		.INIT('hd0)
	) name4828 (
		_w1741_,
		_w5287_,
		_w5290_,
		_w5291_
	);
	LUT3 #(
		.INIT('hd0)
	) name4829 (
		_w2424_,
		_w5285_,
		_w5291_,
		_w5292_
	);
	LUT4 #(
		.INIT('ha8aa)
	) name4830 (
		_w1731_,
		_w5282_,
		_w5284_,
		_w5292_,
		_w5293_
	);
	LUT4 #(
		.INIT('heeec)
	) name4831 (
		\P1_state_reg[0]/NET0131 ,
		_w5278_,
		_w5279_,
		_w5293_,
		_w5294_
	);
	LUT4 #(
		.INIT('h1dd1)
	) name4832 (
		\P1_reg2_reg[15]/NET0131 ,
		_w1741_,
		_w3169_,
		_w4358_,
		_w5295_
	);
	LUT2 #(
		.INIT('h2)
	) name4833 (
		_w2292_,
		_w5295_,
		_w5296_
	);
	LUT4 #(
		.INIT('hd11d)
	) name4834 (
		\P1_reg2_reg[15]/NET0131 ,
		_w1741_,
		_w3169_,
		_w4364_,
		_w5297_
	);
	LUT4 #(
		.INIT('hddd1)
	) name4835 (
		\P1_reg2_reg[15]/NET0131 ,
		_w1741_,
		_w4552_,
		_w4553_,
		_w5298_
	);
	LUT4 #(
		.INIT('h0008)
	) name4836 (
		_w2243_,
		_w2284_,
		_w2288_,
		_w2291_,
		_w5299_
	);
	LUT4 #(
		.INIT('ha2a0)
	) name4837 (
		\P1_reg2_reg[15]/NET0131 ,
		_w1741_,
		_w2450_,
		_w2452_,
		_w5300_
	);
	LUT2 #(
		.INIT('h1)
	) name4838 (
		_w5299_,
		_w5300_,
		_w5301_
	);
	LUT3 #(
		.INIT('h70)
	) name4839 (
		_w1741_,
		_w4555_,
		_w5301_,
		_w5302_
	);
	LUT3 #(
		.INIT('hd0)
	) name4840 (
		_w2424_,
		_w5298_,
		_w5302_,
		_w5303_
	);
	LUT3 #(
		.INIT('hd0)
	) name4841 (
		_w2388_,
		_w5297_,
		_w5303_,
		_w5304_
	);
	LUT4 #(
		.INIT('h2000)
	) name4842 (
		\P1_reg2_reg[15]/NET0131 ,
		_w1723_,
		_w1727_,
		_w1730_,
		_w5305_
	);
	LUT4 #(
		.INIT('h0075)
	) name4843 (
		_w1731_,
		_w5296_,
		_w5304_,
		_w5305_,
		_w5306_
	);
	LUT2 #(
		.INIT('h2)
	) name4844 (
		\P1_reg2_reg[15]/NET0131 ,
		_w2462_,
		_w5307_
	);
	LUT3 #(
		.INIT('hf2)
	) name4845 (
		\P1_state_reg[0]/NET0131 ,
		_w5306_,
		_w5307_,
		_w5308_
	);
	LUT2 #(
		.INIT('h2)
	) name4846 (
		\P1_reg2_reg[14]/NET0131 ,
		_w2462_,
		_w5309_
	);
	LUT4 #(
		.INIT('h2000)
	) name4847 (
		\P1_reg2_reg[14]/NET0131 ,
		_w1723_,
		_w1727_,
		_w1730_,
		_w5310_
	);
	LUT4 #(
		.INIT('hddd1)
	) name4848 (
		\P1_reg2_reg[14]/NET0131 ,
		_w1741_,
		_w4569_,
		_w4570_,
		_w5311_
	);
	LUT2 #(
		.INIT('h2)
	) name4849 (
		_w2424_,
		_w5311_,
		_w5312_
	);
	LUT4 #(
		.INIT('he020)
	) name4850 (
		\P1_reg2_reg[14]/NET0131 ,
		_w1741_,
		_w2292_,
		_w4575_,
		_w5313_
	);
	LUT4 #(
		.INIT('h20e0)
	) name4851 (
		\P1_reg2_reg[14]/NET0131 ,
		_w1741_,
		_w2388_,
		_w4573_,
		_w5314_
	);
	LUT4 #(
		.INIT('h0008)
	) name4852 (
		_w2209_,
		_w2284_,
		_w2288_,
		_w2291_,
		_w5315_
	);
	LUT4 #(
		.INIT('ha2a0)
	) name4853 (
		\P1_reg2_reg[14]/NET0131 ,
		_w1741_,
		_w2450_,
		_w2452_,
		_w5316_
	);
	LUT2 #(
		.INIT('h1)
	) name4854 (
		_w5315_,
		_w5316_,
		_w5317_
	);
	LUT3 #(
		.INIT('hd0)
	) name4855 (
		_w1741_,
		_w4579_,
		_w5317_,
		_w5318_
	);
	LUT3 #(
		.INIT('h10)
	) name4856 (
		_w5314_,
		_w5313_,
		_w5318_,
		_w5319_
	);
	LUT4 #(
		.INIT('h1311)
	) name4857 (
		_w1731_,
		_w5310_,
		_w5312_,
		_w5319_,
		_w5320_
	);
	LUT3 #(
		.INIT('hce)
	) name4858 (
		\P1_state_reg[0]/NET0131 ,
		_w5309_,
		_w5320_,
		_w5321_
	);
	LUT4 #(
		.INIT('hd070)
	) name4859 (
		\P1_state_reg[0]/NET0131 ,
		\P2_IR_reg[23]/NET0131 ,
		\P2_reg1_reg[11]/NET0131 ,
		_w1188_,
		_w5322_
	);
	LUT4 #(
		.INIT('h2000)
	) name4860 (
		\P2_reg1_reg[11]/NET0131 ,
		_w1189_,
		_w1352_,
		_w1356_,
		_w5323_
	);
	LUT4 #(
		.INIT('haa02)
	) name4861 (
		\P2_reg1_reg[11]/NET0131 ,
		_w1361_,
		_w1363_,
		_w1368_,
		_w5324_
	);
	LUT4 #(
		.INIT('h0e02)
	) name4862 (
		\P2_reg1_reg[11]/NET0131 ,
		_w1516_,
		_w1575_,
		_w4600_,
		_w5325_
	);
	LUT2 #(
		.INIT('h4)
	) name4863 (
		_w685_,
		_w2471_,
		_w5326_
	);
	LUT3 #(
		.INIT('ha2)
	) name4864 (
		\P2_reg1_reg[11]/NET0131 ,
		_w1684_,
		_w2469_,
		_w5327_
	);
	LUT2 #(
		.INIT('h1)
	) name4865 (
		_w5326_,
		_w5327_,
		_w5328_
	);
	LUT2 #(
		.INIT('h4)
	) name4866 (
		_w5325_,
		_w5328_,
		_w5329_
	);
	LUT4 #(
		.INIT('ha8aa)
	) name4867 (
		\P2_reg1_reg[11]/NET0131 ,
		_w1361_,
		_w1363_,
		_w1368_,
		_w5330_
	);
	LUT4 #(
		.INIT('h08c8)
	) name4868 (
		\P2_reg1_reg[11]/NET0131 ,
		_w1191_,
		_w1507_,
		_w4598_,
		_w5331_
	);
	LUT4 #(
		.INIT('h9a00)
	) name4869 (
		_w1320_,
		_w1379_,
		_w1383_,
		_w1507_,
		_w5332_
	);
	LUT3 #(
		.INIT('ha8)
	) name4870 (
		_w1530_,
		_w5330_,
		_w5332_,
		_w5333_
	);
	LUT4 #(
		.INIT('h9a00)
	) name4871 (
		_w1320_,
		_w1379_,
		_w1383_,
		_w1516_,
		_w5334_
	);
	LUT3 #(
		.INIT('h54)
	) name4872 (
		_w1506_,
		_w5324_,
		_w5334_,
		_w5335_
	);
	LUT3 #(
		.INIT('h01)
	) name4873 (
		_w5333_,
		_w5335_,
		_w5331_,
		_w5336_
	);
	LUT4 #(
		.INIT('h3111)
	) name4874 (
		_w1359_,
		_w5323_,
		_w5329_,
		_w5336_,
		_w5337_
	);
	LUT3 #(
		.INIT('hce)
	) name4875 (
		\P1_state_reg[0]/NET0131 ,
		_w5322_,
		_w5337_,
		_w5338_
	);
	LUT4 #(
		.INIT('hd070)
	) name4876 (
		\P1_state_reg[0]/NET0131 ,
		\P2_IR_reg[23]/NET0131 ,
		\P2_reg1_reg[14]/NET0131 ,
		_w1188_,
		_w5339_
	);
	LUT4 #(
		.INIT('h2000)
	) name4877 (
		\P2_reg1_reg[14]/NET0131 ,
		_w1189_,
		_w1352_,
		_w1356_,
		_w5340_
	);
	LUT4 #(
		.INIT('h35c5)
	) name4878 (
		\P2_reg1_reg[14]/NET0131 ,
		_w1296_,
		_w1507_,
		_w2557_,
		_w5341_
	);
	LUT2 #(
		.INIT('h2)
	) name4879 (
		_w1530_,
		_w5341_,
		_w5342_
	);
	LUT4 #(
		.INIT('h111d)
	) name4880 (
		\P2_reg1_reg[14]/NET0131 ,
		_w1507_,
		_w4614_,
		_w4615_,
		_w5343_
	);
	LUT4 #(
		.INIT('hf100)
	) name4881 (
		_w546_,
		_w612_,
		_w614_,
		_w1442_,
		_w5344_
	);
	LUT2 #(
		.INIT('h8)
	) name4882 (
		_w1516_,
		_w5344_,
		_w5345_
	);
	LUT3 #(
		.INIT('ha2)
	) name4883 (
		\P2_reg1_reg[14]/NET0131 ,
		_w1684_,
		_w2469_,
		_w5346_
	);
	LUT2 #(
		.INIT('h1)
	) name4884 (
		_w5345_,
		_w5346_,
		_w5347_
	);
	LUT3 #(
		.INIT('hd0)
	) name4885 (
		_w1191_,
		_w5343_,
		_w5347_,
		_w5348_
	);
	LUT4 #(
		.INIT('h35c5)
	) name4886 (
		\P2_reg1_reg[14]/NET0131 ,
		_w1296_,
		_w1516_,
		_w2557_,
		_w5349_
	);
	LUT4 #(
		.INIT('hc535)
	) name4887 (
		\P2_reg1_reg[14]/NET0131 ,
		_w1296_,
		_w1516_,
		_w2540_,
		_w5350_
	);
	LUT4 #(
		.INIT('hfac8)
	) name4888 (
		_w1506_,
		_w1575_,
		_w5349_,
		_w5350_,
		_w5351_
	);
	LUT4 #(
		.INIT('h8aaa)
	) name4889 (
		_w1359_,
		_w5342_,
		_w5348_,
		_w5351_,
		_w5352_
	);
	LUT4 #(
		.INIT('heeec)
	) name4890 (
		\P1_state_reg[0]/NET0131 ,
		_w5339_,
		_w5340_,
		_w5352_,
		_w5353_
	);
	LUT4 #(
		.INIT('hd070)
	) name4891 (
		\P1_state_reg[0]/NET0131 ,
		\P2_IR_reg[23]/NET0131 ,
		\P2_reg1_reg[15]/NET0131 ,
		_w1188_,
		_w5354_
	);
	LUT4 #(
		.INIT('h2000)
	) name4892 (
		\P2_reg1_reg[15]/NET0131 ,
		_w1189_,
		_w1352_,
		_w1356_,
		_w5355_
	);
	LUT4 #(
		.INIT('hc535)
	) name4893 (
		\P2_reg1_reg[15]/NET0131 ,
		_w1295_,
		_w1507_,
		_w3598_,
		_w5356_
	);
	LUT2 #(
		.INIT('h2)
	) name4894 (
		_w1530_,
		_w5356_,
		_w5357_
	);
	LUT4 #(
		.INIT('h111d)
	) name4895 (
		\P2_reg1_reg[15]/NET0131 ,
		_w1507_,
		_w4633_,
		_w4634_,
		_w5358_
	);
	LUT3 #(
		.INIT('h40)
	) name4896 (
		_w594_,
		_w1442_,
		_w1516_,
		_w5359_
	);
	LUT3 #(
		.INIT('ha2)
	) name4897 (
		\P2_reg1_reg[15]/NET0131 ,
		_w1684_,
		_w2469_,
		_w5360_
	);
	LUT2 #(
		.INIT('h1)
	) name4898 (
		_w5359_,
		_w5360_,
		_w5361_
	);
	LUT3 #(
		.INIT('hd0)
	) name4899 (
		_w1191_,
		_w5358_,
		_w5361_,
		_w5362_
	);
	LUT4 #(
		.INIT('haa02)
	) name4900 (
		\P2_reg1_reg[15]/NET0131 ,
		_w1361_,
		_w1363_,
		_w1368_,
		_w5363_
	);
	LUT4 #(
		.INIT('h6500)
	) name4901 (
		_w1295_,
		_w1471_,
		_w1475_,
		_w1516_,
		_w5364_
	);
	LUT3 #(
		.INIT('h54)
	) name4902 (
		_w1575_,
		_w5363_,
		_w5364_,
		_w5365_
	);
	LUT4 #(
		.INIT('hc535)
	) name4903 (
		\P2_reg1_reg[15]/NET0131 ,
		_w1295_,
		_w1516_,
		_w3598_,
		_w5366_
	);
	LUT2 #(
		.INIT('h1)
	) name4904 (
		_w1506_,
		_w5366_,
		_w5367_
	);
	LUT4 #(
		.INIT('h0100)
	) name4905 (
		_w5357_,
		_w5365_,
		_w5367_,
		_w5362_,
		_w5368_
	);
	LUT4 #(
		.INIT('ha0a8)
	) name4906 (
		\P1_state_reg[0]/NET0131 ,
		_w1359_,
		_w5355_,
		_w5368_,
		_w5369_
	);
	LUT2 #(
		.INIT('he)
	) name4907 (
		_w5354_,
		_w5369_,
		_w5370_
	);
	LUT4 #(
		.INIT('hd070)
	) name4908 (
		\P1_state_reg[0]/NET0131 ,
		\P2_IR_reg[23]/NET0131 ,
		\P2_reg2_reg[11]/NET0131 ,
		_w1188_,
		_w5371_
	);
	LUT4 #(
		.INIT('h2000)
	) name4909 (
		\P2_reg2_reg[11]/NET0131 ,
		_w1189_,
		_w1352_,
		_w1356_,
		_w5372_
	);
	LUT4 #(
		.INIT('ha8aa)
	) name4910 (
		\P2_reg2_reg[11]/NET0131 ,
		_w1361_,
		_w1363_,
		_w1368_,
		_w5373_
	);
	LUT4 #(
		.INIT('h0e02)
	) name4911 (
		\P2_reg2_reg[11]/NET0131 ,
		_w1507_,
		_w1575_,
		_w4600_,
		_w5374_
	);
	LUT3 #(
		.INIT('ha8)
	) name4912 (
		\P2_reg2_reg[11]/NET0131 ,
		_w1441_,
		_w1523_,
		_w5375_
	);
	LUT3 #(
		.INIT('h40)
	) name4913 (
		_w674_,
		_w1229_,
		_w1232_,
		_w5376_
	);
	LUT3 #(
		.INIT('h0b)
	) name4914 (
		_w685_,
		_w1522_,
		_w5376_,
		_w5377_
	);
	LUT2 #(
		.INIT('h4)
	) name4915 (
		_w5375_,
		_w5377_,
		_w5378_
	);
	LUT2 #(
		.INIT('h4)
	) name4916 (
		_w5374_,
		_w5378_,
		_w5379_
	);
	LUT4 #(
		.INIT('haa02)
	) name4917 (
		\P2_reg2_reg[11]/NET0131 ,
		_w1361_,
		_w1363_,
		_w1368_,
		_w5380_
	);
	LUT4 #(
		.INIT('h08c8)
	) name4918 (
		\P2_reg2_reg[11]/NET0131 ,
		_w1191_,
		_w1516_,
		_w4598_,
		_w5381_
	);
	LUT3 #(
		.INIT('ha8)
	) name4919 (
		_w1530_,
		_w5334_,
		_w5380_,
		_w5382_
	);
	LUT3 #(
		.INIT('h54)
	) name4920 (
		_w1506_,
		_w5332_,
		_w5373_,
		_w5383_
	);
	LUT3 #(
		.INIT('h01)
	) name4921 (
		_w5382_,
		_w5383_,
		_w5381_,
		_w5384_
	);
	LUT4 #(
		.INIT('h3111)
	) name4922 (
		_w1359_,
		_w5372_,
		_w5379_,
		_w5384_,
		_w5385_
	);
	LUT3 #(
		.INIT('hce)
	) name4923 (
		\P1_state_reg[0]/NET0131 ,
		_w5371_,
		_w5385_,
		_w5386_
	);
	LUT4 #(
		.INIT('hd070)
	) name4924 (
		\P1_state_reg[0]/NET0131 ,
		\P2_IR_reg[23]/NET0131 ,
		\P2_reg2_reg[14]/NET0131 ,
		_w1188_,
		_w5387_
	);
	LUT4 #(
		.INIT('h2000)
	) name4925 (
		\P2_reg2_reg[14]/NET0131 ,
		_w1189_,
		_w1352_,
		_w1356_,
		_w5388_
	);
	LUT4 #(
		.INIT('h35c5)
	) name4926 (
		\P2_reg2_reg[14]/NET0131 ,
		_w1296_,
		_w1516_,
		_w2557_,
		_w5389_
	);
	LUT2 #(
		.INIT('h2)
	) name4927 (
		_w1530_,
		_w5389_,
		_w5390_
	);
	LUT4 #(
		.INIT('h111d)
	) name4928 (
		\P2_reg2_reg[14]/NET0131 ,
		_w1516_,
		_w4614_,
		_w4615_,
		_w5391_
	);
	LUT2 #(
		.INIT('h8)
	) name4929 (
		_w1507_,
		_w5344_,
		_w5392_
	);
	LUT3 #(
		.INIT('h40)
	) name4930 (
		_w620_,
		_w1229_,
		_w1232_,
		_w5393_
	);
	LUT4 #(
		.INIT('h0057)
	) name4931 (
		\P2_reg2_reg[14]/NET0131 ,
		_w1441_,
		_w1523_,
		_w5393_,
		_w5394_
	);
	LUT2 #(
		.INIT('h4)
	) name4932 (
		_w5392_,
		_w5394_,
		_w5395_
	);
	LUT3 #(
		.INIT('hd0)
	) name4933 (
		_w1191_,
		_w5391_,
		_w5395_,
		_w5396_
	);
	LUT4 #(
		.INIT('h35c5)
	) name4934 (
		\P2_reg2_reg[14]/NET0131 ,
		_w1296_,
		_w1507_,
		_w2557_,
		_w5397_
	);
	LUT4 #(
		.INIT('hc535)
	) name4935 (
		\P2_reg2_reg[14]/NET0131 ,
		_w1296_,
		_w1507_,
		_w2540_,
		_w5398_
	);
	LUT4 #(
		.INIT('hfac8)
	) name4936 (
		_w1506_,
		_w1575_,
		_w5397_,
		_w5398_,
		_w5399_
	);
	LUT4 #(
		.INIT('h8aaa)
	) name4937 (
		_w1359_,
		_w5390_,
		_w5396_,
		_w5399_,
		_w5400_
	);
	LUT4 #(
		.INIT('heeec)
	) name4938 (
		\P1_state_reg[0]/NET0131 ,
		_w5387_,
		_w5388_,
		_w5400_,
		_w5401_
	);
	LUT4 #(
		.INIT('hd070)
	) name4939 (
		\P1_state_reg[0]/NET0131 ,
		\P2_IR_reg[23]/NET0131 ,
		\P2_reg2_reg[15]/NET0131 ,
		_w1188_,
		_w5402_
	);
	LUT4 #(
		.INIT('h2000)
	) name4940 (
		\P2_reg2_reg[15]/NET0131 ,
		_w1189_,
		_w1352_,
		_w1356_,
		_w5403_
	);
	LUT4 #(
		.INIT('hc535)
	) name4941 (
		\P2_reg2_reg[15]/NET0131 ,
		_w1295_,
		_w1516_,
		_w3598_,
		_w5404_
	);
	LUT2 #(
		.INIT('h2)
	) name4942 (
		_w1530_,
		_w5404_,
		_w5405_
	);
	LUT4 #(
		.INIT('h111d)
	) name4943 (
		\P2_reg2_reg[15]/NET0131 ,
		_w1516_,
		_w4633_,
		_w4634_,
		_w5406_
	);
	LUT3 #(
		.INIT('h40)
	) name4944 (
		_w594_,
		_w1442_,
		_w1507_,
		_w5407_
	);
	LUT3 #(
		.INIT('h40)
	) name4945 (
		_w525_,
		_w1229_,
		_w1232_,
		_w5408_
	);
	LUT4 #(
		.INIT('h0057)
	) name4946 (
		\P2_reg2_reg[15]/NET0131 ,
		_w1441_,
		_w1523_,
		_w5408_,
		_w5409_
	);
	LUT2 #(
		.INIT('h4)
	) name4947 (
		_w5407_,
		_w5409_,
		_w5410_
	);
	LUT3 #(
		.INIT('hd0)
	) name4948 (
		_w1191_,
		_w5406_,
		_w5410_,
		_w5411_
	);
	LUT4 #(
		.INIT('ha8aa)
	) name4949 (
		\P2_reg2_reg[15]/NET0131 ,
		_w1361_,
		_w1363_,
		_w1368_,
		_w5412_
	);
	LUT4 #(
		.INIT('h6500)
	) name4950 (
		_w1295_,
		_w1471_,
		_w1475_,
		_w1507_,
		_w5413_
	);
	LUT3 #(
		.INIT('h54)
	) name4951 (
		_w1575_,
		_w5412_,
		_w5413_,
		_w5414_
	);
	LUT4 #(
		.INIT('hc535)
	) name4952 (
		\P2_reg2_reg[15]/NET0131 ,
		_w1295_,
		_w1507_,
		_w3598_,
		_w5415_
	);
	LUT2 #(
		.INIT('h1)
	) name4953 (
		_w1506_,
		_w5415_,
		_w5416_
	);
	LUT4 #(
		.INIT('h0100)
	) name4954 (
		_w5405_,
		_w5414_,
		_w5416_,
		_w5411_,
		_w5417_
	);
	LUT4 #(
		.INIT('ha0a8)
	) name4955 (
		\P1_state_reg[0]/NET0131 ,
		_w1359_,
		_w5403_,
		_w5417_,
		_w5418_
	);
	LUT2 #(
		.INIT('he)
	) name4956 (
		_w5402_,
		_w5418_,
		_w5419_
	);
	LUT2 #(
		.INIT('h2)
	) name4957 (
		\P1_reg0_reg[15]/NET0131 ,
		_w2462_,
		_w5420_
	);
	LUT4 #(
		.INIT('h1dd1)
	) name4958 (
		\P1_reg0_reg[15]/NET0131 ,
		_w2883_,
		_w3169_,
		_w4358_,
		_w5421_
	);
	LUT2 #(
		.INIT('h2)
	) name4959 (
		_w2292_,
		_w5421_,
		_w5422_
	);
	LUT4 #(
		.INIT('hd11d)
	) name4960 (
		\P1_reg0_reg[15]/NET0131 ,
		_w2883_,
		_w3169_,
		_w4364_,
		_w5423_
	);
	LUT4 #(
		.INIT('hddd1)
	) name4961 (
		\P1_reg0_reg[15]/NET0131 ,
		_w2883_,
		_w4552_,
		_w4553_,
		_w5424_
	);
	LUT4 #(
		.INIT('h0a8a)
	) name4962 (
		\P1_reg0_reg[15]/NET0131 ,
		_w2452_,
		_w2524_,
		_w2883_,
		_w5425_
	);
	LUT3 #(
		.INIT('h07)
	) name4963 (
		_w2883_,
		_w4555_,
		_w5425_,
		_w5426_
	);
	LUT3 #(
		.INIT('hd0)
	) name4964 (
		_w2424_,
		_w5424_,
		_w5426_,
		_w5427_
	);
	LUT3 #(
		.INIT('hd0)
	) name4965 (
		_w2388_,
		_w5423_,
		_w5427_,
		_w5428_
	);
	LUT4 #(
		.INIT('h2000)
	) name4966 (
		\P1_reg0_reg[15]/NET0131 ,
		_w1723_,
		_w1727_,
		_w1730_,
		_w5429_
	);
	LUT4 #(
		.INIT('h0075)
	) name4967 (
		_w1731_,
		_w5422_,
		_w5428_,
		_w5429_,
		_w5430_
	);
	LUT3 #(
		.INIT('hce)
	) name4968 (
		\P1_state_reg[0]/NET0131 ,
		_w5420_,
		_w5430_,
		_w5431_
	);
	LUT4 #(
		.INIT('h0020)
	) name4969 (
		_w4658_,
		_w4656_,
		_w5244_,
		_w5246_,
		_w5432_
	);
	LUT4 #(
		.INIT('h5515)
	) name4970 (
		\P1_reg0_reg[8]/NET0131 ,
		_w2883_,
		_w5244_,
		_w5432_,
		_w5433_
	);
	LUT4 #(
		.INIT('h0400)
	) name4971 (
		_w4165_,
		_w4658_,
		_w4656_,
		_w5244_,
		_w5434_
	);
	LUT2 #(
		.INIT('h2)
	) name4972 (
		\P1_reg0_reg[8]/NET0131 ,
		_w5434_,
		_w5435_
	);
	LUT3 #(
		.INIT('hc4)
	) name4973 (
		_w2883_,
		_w3408_,
		_w5432_,
		_w5436_
	);
	LUT3 #(
		.INIT('h45)
	) name4974 (
		_w5433_,
		_w5435_,
		_w5436_,
		_w5437_
	);
	LUT4 #(
		.INIT('h1dd1)
	) name4975 (
		\P1_reg1_reg[15]/NET0131 ,
		_w2520_,
		_w3169_,
		_w4358_,
		_w5438_
	);
	LUT2 #(
		.INIT('h2)
	) name4976 (
		_w2292_,
		_w5438_,
		_w5439_
	);
	LUT4 #(
		.INIT('hd11d)
	) name4977 (
		\P1_reg1_reg[15]/NET0131 ,
		_w2520_,
		_w3169_,
		_w4364_,
		_w5440_
	);
	LUT4 #(
		.INIT('hddd1)
	) name4978 (
		\P1_reg1_reg[15]/NET0131 ,
		_w2520_,
		_w4552_,
		_w4553_,
		_w5441_
	);
	LUT4 #(
		.INIT('h08aa)
	) name4979 (
		\P1_reg1_reg[15]/NET0131 ,
		_w2452_,
		_w2520_,
		_w2524_,
		_w5442_
	);
	LUT3 #(
		.INIT('h07)
	) name4980 (
		_w2520_,
		_w4555_,
		_w5442_,
		_w5443_
	);
	LUT3 #(
		.INIT('hd0)
	) name4981 (
		_w2424_,
		_w5441_,
		_w5443_,
		_w5444_
	);
	LUT3 #(
		.INIT('hd0)
	) name4982 (
		_w2388_,
		_w5440_,
		_w5444_,
		_w5445_
	);
	LUT4 #(
		.INIT('h2000)
	) name4983 (
		\P1_reg1_reg[15]/NET0131 ,
		_w1723_,
		_w1727_,
		_w1730_,
		_w5446_
	);
	LUT4 #(
		.INIT('h0075)
	) name4984 (
		_w1731_,
		_w5439_,
		_w5445_,
		_w5446_,
		_w5447_
	);
	LUT2 #(
		.INIT('h2)
	) name4985 (
		\P1_reg1_reg[15]/NET0131 ,
		_w2462_,
		_w5448_
	);
	LUT3 #(
		.INIT('hf2)
	) name4986 (
		\P1_state_reg[0]/NET0131 ,
		_w5447_,
		_w5448_,
		_w5449_
	);
	LUT4 #(
		.INIT('hd070)
	) name4987 (
		\P1_state_reg[0]/NET0131 ,
		\P2_IR_reg[23]/NET0131 ,
		\P2_reg0_reg[11]/NET0131 ,
		_w1188_,
		_w5450_
	);
	LUT4 #(
		.INIT('h2000)
	) name4988 (
		\P2_reg0_reg[11]/NET0131 ,
		_w1189_,
		_w1352_,
		_w1356_,
		_w5451_
	);
	LUT4 #(
		.INIT('haaa8)
	) name4989 (
		\P2_reg0_reg[11]/NET0131 ,
		_w1361_,
		_w1363_,
		_w1368_,
		_w5452_
	);
	LUT4 #(
		.INIT('h9a00)
	) name4990 (
		_w1320_,
		_w1379_,
		_w1383_,
		_w1411_,
		_w5453_
	);
	LUT2 #(
		.INIT('h4)
	) name4991 (
		_w685_,
		_w1687_,
		_w5454_
	);
	LUT3 #(
		.INIT('ha2)
	) name4992 (
		\P2_reg0_reg[11]/NET0131 ,
		_w1684_,
		_w1685_,
		_w5455_
	);
	LUT2 #(
		.INIT('h1)
	) name4993 (
		_w5454_,
		_w5455_,
		_w5456_
	);
	LUT4 #(
		.INIT('hab00)
	) name4994 (
		_w1409_,
		_w5452_,
		_w5453_,
		_w5456_,
		_w5457_
	);
	LUT4 #(
		.INIT('h08c8)
	) name4995 (
		\P2_reg0_reg[11]/NET0131 ,
		_w1191_,
		_w1369_,
		_w4598_,
		_w5458_
	);
	LUT4 #(
		.INIT('h0e02)
	) name4996 (
		\P2_reg0_reg[11]/NET0131 ,
		_w1411_,
		_w1496_,
		_w4600_,
		_w5459_
	);
	LUT4 #(
		.INIT('he020)
	) name4997 (
		\P2_reg0_reg[11]/NET0131 ,
		_w1369_,
		_w1447_,
		_w4600_,
		_w5460_
	);
	LUT4 #(
		.INIT('h0100)
	) name4998 (
		_w5459_,
		_w5460_,
		_w5458_,
		_w5457_,
		_w5461_
	);
	LUT4 #(
		.INIT('ha0a8)
	) name4999 (
		\P1_state_reg[0]/NET0131 ,
		_w1359_,
		_w5451_,
		_w5461_,
		_w5462_
	);
	LUT2 #(
		.INIT('he)
	) name5000 (
		_w5450_,
		_w5462_,
		_w5463_
	);
	LUT4 #(
		.INIT('hd070)
	) name5001 (
		\P1_state_reg[0]/NET0131 ,
		\P2_IR_reg[23]/NET0131 ,
		\P2_reg0_reg[14]/NET0131 ,
		_w1188_,
		_w5464_
	);
	LUT4 #(
		.INIT('h2000)
	) name5002 (
		\P2_reg0_reg[14]/NET0131 ,
		_w1189_,
		_w1352_,
		_w1356_,
		_w5465_
	);
	LUT4 #(
		.INIT('hc535)
	) name5003 (
		\P2_reg0_reg[14]/NET0131 ,
		_w1296_,
		_w1369_,
		_w2540_,
		_w5466_
	);
	LUT2 #(
		.INIT('h2)
	) name5004 (
		_w1447_,
		_w5466_,
		_w5467_
	);
	LUT4 #(
		.INIT('h111d)
	) name5005 (
		\P2_reg0_reg[14]/NET0131 ,
		_w1369_,
		_w4614_,
		_w4615_,
		_w5468_
	);
	LUT2 #(
		.INIT('h8)
	) name5006 (
		_w1411_,
		_w5344_,
		_w5469_
	);
	LUT3 #(
		.INIT('ha2)
	) name5007 (
		\P2_reg0_reg[14]/NET0131 ,
		_w1684_,
		_w1685_,
		_w5470_
	);
	LUT2 #(
		.INIT('h1)
	) name5008 (
		_w5469_,
		_w5470_,
		_w5471_
	);
	LUT3 #(
		.INIT('hd0)
	) name5009 (
		_w1191_,
		_w5468_,
		_w5471_,
		_w5472_
	);
	LUT4 #(
		.INIT('hc535)
	) name5010 (
		\P2_reg0_reg[14]/NET0131 ,
		_w1296_,
		_w1411_,
		_w2540_,
		_w5473_
	);
	LUT4 #(
		.INIT('h35c5)
	) name5011 (
		\P2_reg0_reg[14]/NET0131 ,
		_w1296_,
		_w1411_,
		_w2557_,
		_w5474_
	);
	LUT4 #(
		.INIT('hfca8)
	) name5012 (
		_w1409_,
		_w1496_,
		_w5473_,
		_w5474_,
		_w5475_
	);
	LUT4 #(
		.INIT('h8aaa)
	) name5013 (
		_w1359_,
		_w5467_,
		_w5472_,
		_w5475_,
		_w5476_
	);
	LUT4 #(
		.INIT('heeec)
	) name5014 (
		\P1_state_reg[0]/NET0131 ,
		_w5464_,
		_w5465_,
		_w5476_,
		_w5477_
	);
	LUT2 #(
		.INIT('h1)
	) name5015 (
		\P1_reg3_reg[3]/NET0131 ,
		_w2644_,
		_w5478_
	);
	LUT3 #(
		.INIT('h80)
	) name5016 (
		_w1747_,
		_w2059_,
		_w2060_,
		_w5479_
	);
	LUT4 #(
		.INIT('h00eb)
	) name5017 (
		_w1747_,
		_w2053_,
		_w2400_,
		_w5479_,
		_w5480_
	);
	LUT4 #(
		.INIT('hc404)
	) name5018 (
		\P1_reg3_reg[3]/NET0131 ,
		_w2424_,
		_w2644_,
		_w5480_,
		_w5481_
	);
	LUT4 #(
		.INIT('he010)
	) name5019 (
		_w2066_,
		_w2092_,
		_w2644_,
		_w3188_,
		_w5482_
	);
	LUT3 #(
		.INIT('ha8)
	) name5020 (
		_w2292_,
		_w5478_,
		_w5482_,
		_w5483_
	);
	LUT4 #(
		.INIT('h10e0)
	) name5021 (
		_w2307_,
		_w2308_,
		_w2644_,
		_w3188_,
		_w5484_
	);
	LUT4 #(
		.INIT('h6000)
	) name5022 (
		_w2071_,
		_w2428_,
		_w2447_,
		_w2644_,
		_w5485_
	);
	LUT4 #(
		.INIT('h5450)
	) name5023 (
		_w2071_,
		_w2426_,
		_w2454_,
		_w2644_,
		_w5486_
	);
	LUT4 #(
		.INIT('h000e)
	) name5024 (
		\P1_reg3_reg[3]/NET0131 ,
		_w2690_,
		_w5486_,
		_w5485_,
		_w5487_
	);
	LUT4 #(
		.INIT('h5700)
	) name5025 (
		_w2388_,
		_w5478_,
		_w5484_,
		_w5487_,
		_w5488_
	);
	LUT4 #(
		.INIT('ha8aa)
	) name5026 (
		_w1731_,
		_w5481_,
		_w5483_,
		_w5488_,
		_w5489_
	);
	LUT4 #(
		.INIT('h1000)
	) name5027 (
		\P1_reg3_reg[3]/NET0131 ,
		_w1723_,
		_w1727_,
		_w1730_,
		_w5490_
	);
	LUT3 #(
		.INIT('h9d)
	) name5028 (
		\P1_reg3_reg[3]/NET0131 ,
		\P1_state_reg[0]/NET0131 ,
		_w1723_,
		_w5491_
	);
	LUT4 #(
		.INIT('ha8ff)
	) name5029 (
		\P1_state_reg[0]/NET0131 ,
		_w5489_,
		_w5490_,
		_w5491_,
		_w5492_
	);
	LUT4 #(
		.INIT('h4000)
	) name5030 (
		_w1723_,
		_w1727_,
		_w1730_,
		_w2126_,
		_w5493_
	);
	LUT2 #(
		.INIT('h2)
	) name5031 (
		_w2126_,
		_w2644_,
		_w5494_
	);
	LUT3 #(
		.INIT('h80)
	) name5032 (
		_w1747_,
		_w2135_,
		_w2137_,
		_w5495_
	);
	LUT4 #(
		.INIT('h00eb)
	) name5033 (
		_w1747_,
		_w2118_,
		_w4653_,
		_w5495_,
		_w5496_
	);
	LUT4 #(
		.INIT('hc808)
	) name5034 (
		_w2126_,
		_w2424_,
		_w2644_,
		_w5496_,
		_w5497_
	);
	LUT4 #(
		.INIT('h02a8)
	) name5035 (
		_w2644_,
		_w2749_,
		_w2750_,
		_w3182_,
		_w5498_
	);
	LUT3 #(
		.INIT('ha8)
	) name5036 (
		_w2292_,
		_w5494_,
		_w5498_,
		_w5499_
	);
	LUT4 #(
		.INIT('ha802)
	) name5037 (
		_w2644_,
		_w2797_,
		_w2932_,
		_w3182_,
		_w5500_
	);
	LUT4 #(
		.INIT('h6ccc)
	) name5038 (
		_w2057_,
		_w2124_,
		_w2134_,
		_w2429_,
		_w5501_
	);
	LUT4 #(
		.INIT('hc808)
	) name5039 (
		_w2126_,
		_w2447_,
		_w2644_,
		_w5501_,
		_w5502_
	);
	LUT4 #(
		.INIT('h5450)
	) name5040 (
		_w2124_,
		_w2426_,
		_w2454_,
		_w2644_,
		_w5503_
	);
	LUT4 #(
		.INIT('ha0a8)
	) name5041 (
		_w2126_,
		_w2426_,
		_w2450_,
		_w2644_,
		_w5504_
	);
	LUT2 #(
		.INIT('h1)
	) name5042 (
		_w5503_,
		_w5504_,
		_w5505_
	);
	LUT2 #(
		.INIT('h4)
	) name5043 (
		_w5502_,
		_w5505_,
		_w5506_
	);
	LUT4 #(
		.INIT('h5700)
	) name5044 (
		_w2388_,
		_w5494_,
		_w5500_,
		_w5506_,
		_w5507_
	);
	LUT4 #(
		.INIT('ha8aa)
	) name5045 (
		_w1731_,
		_w5499_,
		_w5497_,
		_w5507_,
		_w5508_
	);
	LUT2 #(
		.INIT('h2)
	) name5046 (
		\P1_reg3_reg[6]/NET0131 ,
		\P1_state_reg[0]/NET0131 ,
		_w5509_
	);
	LUT3 #(
		.INIT('h07)
	) name5047 (
		_w2126_,
		_w2695_,
		_w5509_,
		_w5510_
	);
	LUT4 #(
		.INIT('ha8ff)
	) name5048 (
		\P1_state_reg[0]/NET0131 ,
		_w5493_,
		_w5508_,
		_w5510_,
		_w5511_
	);
	LUT2 #(
		.INIT('h2)
	) name5049 (
		_w2115_,
		_w2644_,
		_w5512_
	);
	LUT4 #(
		.INIT('h4144)
	) name5050 (
		_w1747_,
		_w2108_,
		_w2118_,
		_w4653_,
		_w5513_
	);
	LUT3 #(
		.INIT('h80)
	) name5051 (
		_w1747_,
		_w2125_,
		_w2127_,
		_w5514_
	);
	LUT4 #(
		.INIT('h3331)
	) name5052 (
		_w2644_,
		_w5512_,
		_w5513_,
		_w5514_,
		_w5515_
	);
	LUT4 #(
		.INIT('h07f8)
	) name5053 (
		_w2096_,
		_w2141_,
		_w2145_,
		_w3183_,
		_w5516_
	);
	LUT4 #(
		.INIT('hc808)
	) name5054 (
		_w2115_,
		_w2292_,
		_w2644_,
		_w5516_,
		_w5517_
	);
	LUT4 #(
		.INIT('he010)
	) name5055 (
		_w2316_,
		_w2320_,
		_w2644_,
		_w3183_,
		_w5518_
	);
	LUT4 #(
		.INIT('h4ccc)
	) name5056 (
		_w2057_,
		_w2114_,
		_w2429_,
		_w2430_,
		_w5519_
	);
	LUT4 #(
		.INIT('h0040)
	) name5057 (
		_w2431_,
		_w2447_,
		_w2644_,
		_w5519_,
		_w5520_
	);
	LUT4 #(
		.INIT('ha8a0)
	) name5058 (
		_w2114_,
		_w2426_,
		_w2454_,
		_w2644_,
		_w5521_
	);
	LUT3 #(
		.INIT('h0d)
	) name5059 (
		_w2115_,
		_w2690_,
		_w5521_,
		_w5522_
	);
	LUT2 #(
		.INIT('h4)
	) name5060 (
		_w5520_,
		_w5522_,
		_w5523_
	);
	LUT4 #(
		.INIT('h5700)
	) name5061 (
		_w2388_,
		_w5512_,
		_w5518_,
		_w5523_,
		_w5524_
	);
	LUT4 #(
		.INIT('h0d00)
	) name5062 (
		_w2424_,
		_w5515_,
		_w5517_,
		_w5524_,
		_w5525_
	);
	LUT4 #(
		.INIT('h4000)
	) name5063 (
		_w1723_,
		_w1727_,
		_w1730_,
		_w2115_,
		_w5526_
	);
	LUT4 #(
		.INIT('haa08)
	) name5064 (
		\P1_state_reg[0]/NET0131 ,
		_w1731_,
		_w5525_,
		_w5526_,
		_w5527_
	);
	LUT2 #(
		.INIT('h2)
	) name5065 (
		\P1_reg3_reg[7]/NET0131 ,
		\P1_state_reg[0]/NET0131 ,
		_w5528_
	);
	LUT3 #(
		.INIT('h07)
	) name5066 (
		_w2115_,
		_w2695_,
		_w5528_,
		_w5529_
	);
	LUT2 #(
		.INIT('hb)
	) name5067 (
		_w5527_,
		_w5529_,
		_w5530_
	);
	LUT4 #(
		.INIT('h1000)
	) name5068 (
		_w776_,
		_w1189_,
		_w1352_,
		_w1356_,
		_w5531_
	);
	LUT2 #(
		.INIT('h1)
	) name5069 (
		_w792_,
		_w1435_,
		_w5532_
	);
	LUT4 #(
		.INIT('h007b)
	) name5070 (
		_w770_,
		_w1435_,
		_w5152_,
		_w5532_,
		_w5533_
	);
	LUT4 #(
		.INIT('h04c4)
	) name5071 (
		_w776_,
		_w1191_,
		_w1411_,
		_w5533_,
		_w5534_
	);
	LUT4 #(
		.INIT('h07f8)
	) name5072 (
		_w809_,
		_w1210_,
		_w1211_,
		_w1325_,
		_w5535_
	);
	LUT4 #(
		.INIT('h010d)
	) name5073 (
		_w776_,
		_w1369_,
		_w1409_,
		_w5535_,
		_w5536_
	);
	LUT3 #(
		.INIT('h04)
	) name5074 (
		_w785_,
		_w1232_,
		_w1439_,
		_w5537_
	);
	LUT3 #(
		.INIT('h54)
	) name5075 (
		_w776_,
		_w1441_,
		_w1443_,
		_w5538_
	);
	LUT2 #(
		.INIT('h1)
	) name5076 (
		_w5537_,
		_w5538_,
		_w5539_
	);
	LUT4 #(
		.INIT('h559a)
	) name5077 (
		_w1325_,
		_w1452_,
		_w1453_,
		_w1532_,
		_w5540_
	);
	LUT4 #(
		.INIT('h0d01)
	) name5078 (
		_w776_,
		_w1369_,
		_w1496_,
		_w5540_,
		_w5541_
	);
	LUT4 #(
		.INIT('hc404)
	) name5079 (
		_w776_,
		_w1447_,
		_w1411_,
		_w5540_,
		_w5542_
	);
	LUT4 #(
		.INIT('h0100)
	) name5080 (
		_w5536_,
		_w5541_,
		_w5542_,
		_w5539_,
		_w5543_
	);
	LUT4 #(
		.INIT('h1311)
	) name5081 (
		_w1359_,
		_w5531_,
		_w5534_,
		_w5543_,
		_w5544_
	);
	LUT2 #(
		.INIT('h4)
	) name5082 (
		\P1_state_reg[0]/NET0131 ,
		\P2_reg3_reg[4]/NET0131 ,
		_w5545_
	);
	LUT4 #(
		.INIT('h0802)
	) name5083 (
		\P1_state_reg[0]/NET0131 ,
		\P2_IR_reg[23]/NET0131 ,
		_w776_,
		_w1188_,
		_w5546_
	);
	LUT2 #(
		.INIT('h1)
	) name5084 (
		_w5545_,
		_w5546_,
		_w5547_
	);
	LUT3 #(
		.INIT('h2f)
	) name5085 (
		\P1_state_reg[0]/NET0131 ,
		_w5544_,
		_w5547_,
		_w5548_
	);
	LUT2 #(
		.INIT('h2)
	) name5086 (
		\P1_reg2_reg[5]/NET0131 ,
		_w2462_,
		_w5549_
	);
	LUT2 #(
		.INIT('h2)
	) name5087 (
		\P1_reg2_reg[5]/NET0131 ,
		_w1741_,
		_w5550_
	);
	LUT4 #(
		.INIT('h2a08)
	) name5088 (
		_w1741_,
		_w1747_,
		_w2053_,
		_w5130_,
		_w5551_
	);
	LUT3 #(
		.INIT('ha8)
	) name5089 (
		_w2424_,
		_w5550_,
		_w5551_,
		_w5552_
	);
	LUT4 #(
		.INIT('hd11d)
	) name5090 (
		\P1_reg2_reg[5]/NET0131 ,
		_w1741_,
		_w2096_,
		_w3187_,
		_w5553_
	);
	LUT2 #(
		.INIT('h2)
	) name5091 (
		_w2292_,
		_w5553_,
		_w5554_
	);
	LUT4 #(
		.INIT('h1dd1)
	) name5092 (
		\P1_reg2_reg[5]/NET0131 ,
		_w1741_,
		_w3187_,
		_w5135_,
		_w5555_
	);
	LUT2 #(
		.INIT('h4)
	) name5093 (
		_w2134_,
		_w2426_,
		_w5556_
	);
	LUT3 #(
		.INIT('ha8)
	) name5094 (
		_w1741_,
		_w5137_,
		_w5556_,
		_w5557_
	);
	LUT4 #(
		.INIT('h0008)
	) name5095 (
		_w2136_,
		_w2284_,
		_w2288_,
		_w2291_,
		_w5558_
	);
	LUT4 #(
		.INIT('ha2a0)
	) name5096 (
		\P1_reg2_reg[5]/NET0131 ,
		_w1741_,
		_w2450_,
		_w2452_,
		_w5559_
	);
	LUT2 #(
		.INIT('h1)
	) name5097 (
		_w5558_,
		_w5559_,
		_w5560_
	);
	LUT2 #(
		.INIT('h4)
	) name5098 (
		_w5557_,
		_w5560_,
		_w5561_
	);
	LUT3 #(
		.INIT('hd0)
	) name5099 (
		_w2388_,
		_w5555_,
		_w5561_,
		_w5562_
	);
	LUT4 #(
		.INIT('ha8aa)
	) name5100 (
		_w1731_,
		_w5552_,
		_w5554_,
		_w5562_,
		_w5563_
	);
	LUT4 #(
		.INIT('h2000)
	) name5101 (
		\P1_reg2_reg[5]/NET0131 ,
		_w1723_,
		_w1727_,
		_w1730_,
		_w5564_
	);
	LUT4 #(
		.INIT('heeec)
	) name5102 (
		\P1_state_reg[0]/NET0131 ,
		_w5549_,
		_w5563_,
		_w5564_,
		_w5565_
	);
	LUT2 #(
		.INIT('h2)
	) name5103 (
		\P1_reg1_reg[5]/NET0131 ,
		_w2520_,
		_w5566_
	);
	LUT4 #(
		.INIT('h7020)
	) name5104 (
		_w1747_,
		_w2053_,
		_w2520_,
		_w5130_,
		_w5567_
	);
	LUT3 #(
		.INIT('ha8)
	) name5105 (
		_w2424_,
		_w5566_,
		_w5567_,
		_w5568_
	);
	LUT4 #(
		.INIT('hc535)
	) name5106 (
		\P1_reg1_reg[5]/NET0131 ,
		_w2096_,
		_w2520_,
		_w3187_,
		_w5569_
	);
	LUT2 #(
		.INIT('h2)
	) name5107 (
		_w2292_,
		_w5569_,
		_w5570_
	);
	LUT4 #(
		.INIT('h1dd1)
	) name5108 (
		\P1_reg1_reg[5]/NET0131 ,
		_w2520_,
		_w3187_,
		_w5135_,
		_w5571_
	);
	LUT2 #(
		.INIT('h2)
	) name5109 (
		\P1_reg1_reg[5]/NET0131 ,
		_w2525_,
		_w5572_
	);
	LUT3 #(
		.INIT('ha8)
	) name5110 (
		_w2520_,
		_w5137_,
		_w5556_,
		_w5573_
	);
	LUT2 #(
		.INIT('h1)
	) name5111 (
		_w5572_,
		_w5573_,
		_w5574_
	);
	LUT3 #(
		.INIT('hd0)
	) name5112 (
		_w2388_,
		_w5571_,
		_w5574_,
		_w5575_
	);
	LUT4 #(
		.INIT('ha8aa)
	) name5113 (
		_w1731_,
		_w5568_,
		_w5570_,
		_w5575_,
		_w5576_
	);
	LUT4 #(
		.INIT('h2000)
	) name5114 (
		\P1_reg1_reg[5]/NET0131 ,
		_w1723_,
		_w1727_,
		_w1730_,
		_w5577_
	);
	LUT2 #(
		.INIT('h2)
	) name5115 (
		\P1_reg1_reg[5]/NET0131 ,
		_w2462_,
		_w5578_
	);
	LUT4 #(
		.INIT('hffa8)
	) name5116 (
		\P1_state_reg[0]/NET0131 ,
		_w5576_,
		_w5577_,
		_w5578_,
		_w5579_
	);
	LUT4 #(
		.INIT('hd070)
	) name5117 (
		\P1_state_reg[0]/NET0131 ,
		\P2_IR_reg[23]/NET0131 ,
		\P2_reg0_reg[5]/NET0131 ,
		_w1188_,
		_w5580_
	);
	LUT4 #(
		.INIT('h2000)
	) name5118 (
		\P2_reg0_reg[5]/NET0131 ,
		_w1189_,
		_w1352_,
		_w1356_,
		_w5581_
	);
	LUT4 #(
		.INIT('h02aa)
	) name5119 (
		\P2_reg0_reg[5]/NET0131 ,
		_w1361_,
		_w1363_,
		_w1368_,
		_w5582_
	);
	LUT4 #(
		.INIT('h111d)
	) name5120 (
		\P2_reg0_reg[5]/NET0131 ,
		_w1369_,
		_w5150_,
		_w5154_,
		_w5583_
	);
	LUT2 #(
		.INIT('h2)
	) name5121 (
		_w1191_,
		_w5583_,
		_w5584_
	);
	LUT4 #(
		.INIT('haaa8)
	) name5122 (
		\P2_reg0_reg[5]/NET0131 ,
		_w1361_,
		_w1363_,
		_w1368_,
		_w5585_
	);
	LUT4 #(
		.INIT('hc900)
	) name5123 (
		_w786_,
		_w1306_,
		_w1375_,
		_w1411_,
		_w5586_
	);
	LUT3 #(
		.INIT('h54)
	) name5124 (
		_w1409_,
		_w5585_,
		_w5586_,
		_w5587_
	);
	LUT3 #(
		.INIT('h54)
	) name5125 (
		_w1496_,
		_w5162_,
		_w5585_,
		_w5588_
	);
	LUT2 #(
		.INIT('h4)
	) name5126 (
		_w774_,
		_w1442_,
		_w5589_
	);
	LUT2 #(
		.INIT('h8)
	) name5127 (
		_w1411_,
		_w5589_,
		_w5590_
	);
	LUT3 #(
		.INIT('ha2)
	) name5128 (
		\P2_reg0_reg[5]/NET0131 ,
		_w1684_,
		_w1685_,
		_w5591_
	);
	LUT2 #(
		.INIT('h1)
	) name5129 (
		_w5590_,
		_w5591_,
		_w5592_
	);
	LUT4 #(
		.INIT('h5700)
	) name5130 (
		_w1447_,
		_w5160_,
		_w5582_,
		_w5592_,
		_w5593_
	);
	LUT3 #(
		.INIT('h10)
	) name5131 (
		_w5587_,
		_w5588_,
		_w5593_,
		_w5594_
	);
	LUT4 #(
		.INIT('h1311)
	) name5132 (
		_w1359_,
		_w5581_,
		_w5584_,
		_w5594_,
		_w5595_
	);
	LUT3 #(
		.INIT('hce)
	) name5133 (
		\P1_state_reg[0]/NET0131 ,
		_w5580_,
		_w5595_,
		_w5596_
	);
	LUT4 #(
		.INIT('hd070)
	) name5134 (
		\P1_state_reg[0]/NET0131 ,
		\P2_IR_reg[23]/NET0131 ,
		\P2_reg0_reg[6]/NET0131 ,
		_w1188_,
		_w5597_
	);
	LUT4 #(
		.INIT('h2000)
	) name5135 (
		\P2_reg0_reg[6]/NET0131 ,
		_w1189_,
		_w1352_,
		_w1356_,
		_w5598_
	);
	LUT4 #(
		.INIT('haaa8)
	) name5136 (
		\P2_reg0_reg[6]/NET0131 ,
		_w1361_,
		_w1363_,
		_w1368_,
		_w5599_
	);
	LUT4 #(
		.INIT('he100)
	) name5137 (
		_w1212_,
		_w1213_,
		_w1322_,
		_w1411_,
		_w5600_
	);
	LUT2 #(
		.INIT('h4)
	) name5138 (
		_w752_,
		_w1442_,
		_w5601_
	);
	LUT2 #(
		.INIT('h8)
	) name5139 (
		_w1411_,
		_w5601_,
		_w5602_
	);
	LUT3 #(
		.INIT('ha2)
	) name5140 (
		\P2_reg0_reg[6]/NET0131 ,
		_w1684_,
		_w1685_,
		_w5603_
	);
	LUT2 #(
		.INIT('h1)
	) name5141 (
		_w5602_,
		_w5603_,
		_w5604_
	);
	LUT4 #(
		.INIT('hab00)
	) name5142 (
		_w1409_,
		_w5599_,
		_w5600_,
		_w5604_,
		_w5605_
	);
	LUT3 #(
		.INIT('h54)
	) name5143 (
		_w1496_,
		_w5183_,
		_w5599_,
		_w5606_
	);
	LUT4 #(
		.INIT('h02aa)
	) name5144 (
		\P2_reg0_reg[6]/NET0131 ,
		_w1361_,
		_w1363_,
		_w1368_,
		_w5607_
	);
	LUT3 #(
		.INIT('ha8)
	) name5145 (
		_w1447_,
		_w5175_,
		_w5607_,
		_w5608_
	);
	LUT4 #(
		.INIT('h08c8)
	) name5146 (
		\P2_reg0_reg[6]/NET0131 ,
		_w1191_,
		_w1369_,
		_w5187_,
		_w5609_
	);
	LUT4 #(
		.INIT('h0100)
	) name5147 (
		_w5608_,
		_w5609_,
		_w5606_,
		_w5605_,
		_w5610_
	);
	LUT4 #(
		.INIT('ha0a8)
	) name5148 (
		\P1_state_reg[0]/NET0131 ,
		_w1359_,
		_w5598_,
		_w5610_,
		_w5611_
	);
	LUT2 #(
		.INIT('he)
	) name5149 (
		_w5597_,
		_w5611_,
		_w5612_
	);
	LUT4 #(
		.INIT('hd070)
	) name5150 (
		\P1_state_reg[0]/NET0131 ,
		\P2_IR_reg[23]/NET0131 ,
		\P2_reg0_reg[7]/NET0131 ,
		_w1188_,
		_w5613_
	);
	LUT4 #(
		.INIT('h2000)
	) name5151 (
		\P2_reg0_reg[7]/NET0131 ,
		_w1189_,
		_w1352_,
		_w1356_,
		_w5614_
	);
	LUT4 #(
		.INIT('h3202)
	) name5152 (
		\P2_reg0_reg[7]/NET0131 ,
		_w1409_,
		_w1411_,
		_w5208_,
		_w5615_
	);
	LUT4 #(
		.INIT('h111d)
	) name5153 (
		\P2_reg0_reg[7]/NET0131 ,
		_w1369_,
		_w5200_,
		_w5201_,
		_w5616_
	);
	LUT2 #(
		.INIT('h4)
	) name5154 (
		_w763_,
		_w1442_,
		_w5617_
	);
	LUT2 #(
		.INIT('h8)
	) name5155 (
		_w1411_,
		_w5617_,
		_w5618_
	);
	LUT3 #(
		.INIT('ha2)
	) name5156 (
		\P2_reg0_reg[7]/NET0131 ,
		_w1684_,
		_w1685_,
		_w5619_
	);
	LUT2 #(
		.INIT('h1)
	) name5157 (
		_w5618_,
		_w5619_,
		_w5620_
	);
	LUT4 #(
		.INIT('h3100)
	) name5158 (
		_w1191_,
		_w5615_,
		_w5616_,
		_w5620_,
		_w5621_
	);
	LUT4 #(
		.INIT('hc535)
	) name5159 (
		\P2_reg0_reg[7]/NET0131 ,
		_w1303_,
		_w1369_,
		_w1458_,
		_w5622_
	);
	LUT4 #(
		.INIT('hc535)
	) name5160 (
		\P2_reg0_reg[7]/NET0131 ,
		_w1303_,
		_w1411_,
		_w1458_,
		_w5623_
	);
	LUT4 #(
		.INIT('hf5c4)
	) name5161 (
		_w1447_,
		_w1496_,
		_w5622_,
		_w5623_,
		_w5624_
	);
	LUT4 #(
		.INIT('h3111)
	) name5162 (
		_w1359_,
		_w5614_,
		_w5621_,
		_w5624_,
		_w5625_
	);
	LUT3 #(
		.INIT('hce)
	) name5163 (
		\P1_state_reg[0]/NET0131 ,
		_w5613_,
		_w5625_,
		_w5626_
	);
	LUT4 #(
		.INIT('hd070)
	) name5164 (
		\P1_state_reg[0]/NET0131 ,
		\P2_IR_reg[23]/NET0131 ,
		\P2_reg0_reg[8]/NET0131 ,
		_w1188_,
		_w5627_
	);
	LUT4 #(
		.INIT('h2000)
	) name5165 (
		\P2_reg0_reg[8]/NET0131 ,
		_w1189_,
		_w1352_,
		_w1356_,
		_w5628_
	);
	LUT4 #(
		.INIT('h35c5)
	) name5166 (
		\P2_reg0_reg[8]/NET0131 ,
		_w1310_,
		_w1369_,
		_w1537_,
		_w5629_
	);
	LUT4 #(
		.INIT('h08c8)
	) name5167 (
		\P2_reg0_reg[8]/NET0131 ,
		_w1191_,
		_w1369_,
		_w4672_,
		_w5630_
	);
	LUT2 #(
		.INIT('h4)
	) name5168 (
		_w731_,
		_w1442_,
		_w5631_
	);
	LUT2 #(
		.INIT('h8)
	) name5169 (
		_w1411_,
		_w5631_,
		_w5632_
	);
	LUT3 #(
		.INIT('ha2)
	) name5170 (
		\P2_reg0_reg[8]/NET0131 ,
		_w1684_,
		_w1685_,
		_w5633_
	);
	LUT2 #(
		.INIT('h1)
	) name5171 (
		_w5632_,
		_w5633_,
		_w5634_
	);
	LUT4 #(
		.INIT('h0d00)
	) name5172 (
		_w1447_,
		_w5629_,
		_w5630_,
		_w5634_,
		_w5635_
	);
	LUT4 #(
		.INIT('h35c5)
	) name5173 (
		\P2_reg0_reg[8]/NET0131 ,
		_w1310_,
		_w1411_,
		_w1537_,
		_w5636_
	);
	LUT4 #(
		.INIT('hc355)
	) name5174 (
		\P2_reg0_reg[8]/NET0131 ,
		_w1215_,
		_w1310_,
		_w1411_,
		_w5637_
	);
	LUT4 #(
		.INIT('hfca8)
	) name5175 (
		_w1409_,
		_w1496_,
		_w5636_,
		_w5637_,
		_w5638_
	);
	LUT4 #(
		.INIT('h3111)
	) name5176 (
		_w1359_,
		_w5628_,
		_w5635_,
		_w5638_,
		_w5639_
	);
	LUT3 #(
		.INIT('hce)
	) name5177 (
		\P1_state_reg[0]/NET0131 ,
		_w5627_,
		_w5639_,
		_w5640_
	);
	LUT2 #(
		.INIT('h2)
	) name5178 (
		\P1_reg2_reg[4]/NET0131 ,
		_w2462_,
		_w5641_
	);
	LUT4 #(
		.INIT('h2000)
	) name5179 (
		\P1_reg2_reg[4]/NET0131 ,
		_w1723_,
		_w1727_,
		_w1730_,
		_w5642_
	);
	LUT4 #(
		.INIT('hddd1)
	) name5180 (
		\P1_reg2_reg[4]/NET0131 ,
		_w1741_,
		_w5112_,
		_w5113_,
		_w5643_
	);
	LUT2 #(
		.INIT('h2)
	) name5181 (
		_w2424_,
		_w5643_,
		_w5644_
	);
	LUT4 #(
		.INIT('he020)
	) name5182 (
		\P1_reg2_reg[4]/NET0131 ,
		_w1741_,
		_w2388_,
		_w5116_,
		_w5645_
	);
	LUT4 #(
		.INIT('h20e0)
	) name5183 (
		\P1_reg2_reg[4]/NET0131 ,
		_w1741_,
		_w2292_,
		_w5118_,
		_w5646_
	);
	LUT4 #(
		.INIT('hd11d)
	) name5184 (
		\P1_reg2_reg[4]/NET0131 ,
		_w1741_,
		_w2057_,
		_w2429_,
		_w5647_
	);
	LUT4 #(
		.INIT('haa20)
	) name5185 (
		\P1_reg2_reg[4]/NET0131 ,
		_w1741_,
		_w2426_,
		_w2450_,
		_w5648_
	);
	LUT4 #(
		.INIT('h0008)
	) name5186 (
		_w2050_,
		_w2284_,
		_w2288_,
		_w2291_,
		_w5649_
	);
	LUT3 #(
		.INIT('h07)
	) name5187 (
		_w1741_,
		_w5223_,
		_w5649_,
		_w5650_
	);
	LUT4 #(
		.INIT('h3100)
	) name5188 (
		_w2447_,
		_w5648_,
		_w5647_,
		_w5650_,
		_w5651_
	);
	LUT3 #(
		.INIT('h10)
	) name5189 (
		_w5646_,
		_w5645_,
		_w5651_,
		_w5652_
	);
	LUT4 #(
		.INIT('h1311)
	) name5190 (
		_w1731_,
		_w5642_,
		_w5644_,
		_w5652_,
		_w5653_
	);
	LUT3 #(
		.INIT('hce)
	) name5191 (
		\P1_state_reg[0]/NET0131 ,
		_w5641_,
		_w5653_,
		_w5654_
	);
	LUT4 #(
		.INIT('hd070)
	) name5192 (
		\P1_state_reg[0]/NET0131 ,
		\P2_IR_reg[23]/NET0131 ,
		\P2_reg1_reg[5]/NET0131 ,
		_w1188_,
		_w5655_
	);
	LUT4 #(
		.INIT('h2000)
	) name5193 (
		\P2_reg1_reg[5]/NET0131 ,
		_w1189_,
		_w1352_,
		_w1356_,
		_w5656_
	);
	LUT4 #(
		.INIT('ha8aa)
	) name5194 (
		\P2_reg1_reg[5]/NET0131 ,
		_w1361_,
		_w1363_,
		_w1368_,
		_w5657_
	);
	LUT4 #(
		.INIT('h111d)
	) name5195 (
		\P2_reg1_reg[5]/NET0131 ,
		_w1507_,
		_w5150_,
		_w5154_,
		_w5658_
	);
	LUT2 #(
		.INIT('h2)
	) name5196 (
		_w1191_,
		_w5658_,
		_w5659_
	);
	LUT4 #(
		.INIT('hc900)
	) name5197 (
		_w786_,
		_w1306_,
		_w1375_,
		_w1507_,
		_w5660_
	);
	LUT3 #(
		.INIT('ha8)
	) name5198 (
		_w1530_,
		_w5657_,
		_w5660_,
		_w5661_
	);
	LUT4 #(
		.INIT('haa02)
	) name5199 (
		\P2_reg1_reg[5]/NET0131 ,
		_w1361_,
		_w1363_,
		_w1368_,
		_w5662_
	);
	LUT4 #(
		.INIT('hc900)
	) name5200 (
		_w786_,
		_w1306_,
		_w1375_,
		_w1516_,
		_w5663_
	);
	LUT3 #(
		.INIT('h54)
	) name5201 (
		_w1506_,
		_w5662_,
		_w5663_,
		_w5664_
	);
	LUT4 #(
		.INIT('ha900)
	) name5202 (
		_w1306_,
		_w1454_,
		_w1455_,
		_w1516_,
		_w5665_
	);
	LUT2 #(
		.INIT('h8)
	) name5203 (
		_w1516_,
		_w5589_,
		_w5666_
	);
	LUT3 #(
		.INIT('ha2)
	) name5204 (
		\P2_reg1_reg[5]/NET0131 ,
		_w1684_,
		_w2469_,
		_w5667_
	);
	LUT2 #(
		.INIT('h1)
	) name5205 (
		_w5666_,
		_w5667_,
		_w5668_
	);
	LUT4 #(
		.INIT('hab00)
	) name5206 (
		_w1575_,
		_w5662_,
		_w5665_,
		_w5668_,
		_w5669_
	);
	LUT3 #(
		.INIT('h10)
	) name5207 (
		_w5664_,
		_w5661_,
		_w5669_,
		_w5670_
	);
	LUT4 #(
		.INIT('h1311)
	) name5208 (
		_w1359_,
		_w5656_,
		_w5659_,
		_w5670_,
		_w5671_
	);
	LUT3 #(
		.INIT('hce)
	) name5209 (
		\P1_state_reg[0]/NET0131 ,
		_w5655_,
		_w5671_,
		_w5672_
	);
	LUT4 #(
		.INIT('hd070)
	) name5210 (
		\P1_state_reg[0]/NET0131 ,
		\P2_IR_reg[23]/NET0131 ,
		\P2_reg1_reg[6]/NET0131 ,
		_w1188_,
		_w5673_
	);
	LUT4 #(
		.INIT('h2000)
	) name5211 (
		\P2_reg1_reg[6]/NET0131 ,
		_w1189_,
		_w1352_,
		_w1356_,
		_w5674_
	);
	LUT4 #(
		.INIT('haa02)
	) name5212 (
		\P2_reg1_reg[6]/NET0131 ,
		_w1361_,
		_w1363_,
		_w1368_,
		_w5675_
	);
	LUT4 #(
		.INIT('h4844)
	) name5213 (
		_w1322_,
		_w1516_,
		_w1534_,
		_w1535_,
		_w5676_
	);
	LUT2 #(
		.INIT('h8)
	) name5214 (
		_w1516_,
		_w5601_,
		_w5677_
	);
	LUT3 #(
		.INIT('ha2)
	) name5215 (
		\P2_reg1_reg[6]/NET0131 ,
		_w1684_,
		_w2469_,
		_w5678_
	);
	LUT2 #(
		.INIT('h1)
	) name5216 (
		_w5677_,
		_w5678_,
		_w5679_
	);
	LUT4 #(
		.INIT('hab00)
	) name5217 (
		_w1575_,
		_w5675_,
		_w5676_,
		_w5679_,
		_w5680_
	);
	LUT4 #(
		.INIT('he100)
	) name5218 (
		_w1212_,
		_w1213_,
		_w1322_,
		_w1516_,
		_w5681_
	);
	LUT3 #(
		.INIT('h54)
	) name5219 (
		_w1506_,
		_w5675_,
		_w5681_,
		_w5682_
	);
	LUT4 #(
		.INIT('ha8aa)
	) name5220 (
		\P2_reg1_reg[6]/NET0131 ,
		_w1361_,
		_w1363_,
		_w1368_,
		_w5683_
	);
	LUT4 #(
		.INIT('he100)
	) name5221 (
		_w1212_,
		_w1213_,
		_w1322_,
		_w1507_,
		_w5684_
	);
	LUT3 #(
		.INIT('ha8)
	) name5222 (
		_w1530_,
		_w5683_,
		_w5684_,
		_w5685_
	);
	LUT4 #(
		.INIT('h08c8)
	) name5223 (
		\P2_reg1_reg[6]/NET0131 ,
		_w1191_,
		_w1507_,
		_w5187_,
		_w5686_
	);
	LUT4 #(
		.INIT('h0100)
	) name5224 (
		_w5685_,
		_w5686_,
		_w5682_,
		_w5680_,
		_w5687_
	);
	LUT4 #(
		.INIT('ha0a8)
	) name5225 (
		\P1_state_reg[0]/NET0131 ,
		_w1359_,
		_w5674_,
		_w5687_,
		_w5688_
	);
	LUT2 #(
		.INIT('he)
	) name5226 (
		_w5673_,
		_w5688_,
		_w5689_
	);
	LUT4 #(
		.INIT('hd070)
	) name5227 (
		\P1_state_reg[0]/NET0131 ,
		\P2_IR_reg[23]/NET0131 ,
		\P2_reg1_reg[7]/NET0131 ,
		_w1188_,
		_w5690_
	);
	LUT4 #(
		.INIT('h2000)
	) name5228 (
		\P2_reg1_reg[7]/NET0131 ,
		_w1189_,
		_w1352_,
		_w1356_,
		_w5691_
	);
	LUT4 #(
		.INIT('hc355)
	) name5229 (
		\P2_reg1_reg[7]/NET0131 ,
		_w1303_,
		_w1458_,
		_w1516_,
		_w5692_
	);
	LUT2 #(
		.INIT('h1)
	) name5230 (
		_w1575_,
		_w5692_,
		_w5693_
	);
	LUT4 #(
		.INIT('h111d)
	) name5231 (
		\P2_reg1_reg[7]/NET0131 ,
		_w1507_,
		_w5200_,
		_w5201_,
		_w5694_
	);
	LUT2 #(
		.INIT('h8)
	) name5232 (
		_w1516_,
		_w5617_,
		_w5695_
	);
	LUT3 #(
		.INIT('ha2)
	) name5233 (
		\P2_reg1_reg[7]/NET0131 ,
		_w1684_,
		_w2469_,
		_w5696_
	);
	LUT2 #(
		.INIT('h1)
	) name5234 (
		_w5695_,
		_w5696_,
		_w5697_
	);
	LUT3 #(
		.INIT('hd0)
	) name5235 (
		_w1191_,
		_w5694_,
		_w5697_,
		_w5698_
	);
	LUT4 #(
		.INIT('he020)
	) name5236 (
		\P2_reg1_reg[7]/NET0131 ,
		_w1507_,
		_w1530_,
		_w5208_,
		_w5699_
	);
	LUT4 #(
		.INIT('h3202)
	) name5237 (
		\P2_reg1_reg[7]/NET0131 ,
		_w1506_,
		_w1516_,
		_w5208_,
		_w5700_
	);
	LUT2 #(
		.INIT('h1)
	) name5238 (
		_w5699_,
		_w5700_,
		_w5701_
	);
	LUT4 #(
		.INIT('h8aaa)
	) name5239 (
		_w1359_,
		_w5693_,
		_w5698_,
		_w5701_,
		_w5702_
	);
	LUT4 #(
		.INIT('heeec)
	) name5240 (
		\P1_state_reg[0]/NET0131 ,
		_w5690_,
		_w5691_,
		_w5702_,
		_w5703_
	);
	LUT4 #(
		.INIT('hd070)
	) name5241 (
		\P1_state_reg[0]/NET0131 ,
		\P2_IR_reg[23]/NET0131 ,
		\P2_reg1_reg[8]/NET0131 ,
		_w1188_,
		_w5704_
	);
	LUT4 #(
		.INIT('h2000)
	) name5242 (
		\P2_reg1_reg[8]/NET0131 ,
		_w1189_,
		_w1352_,
		_w1356_,
		_w5705_
	);
	LUT4 #(
		.INIT('h35c5)
	) name5243 (
		\P2_reg1_reg[8]/NET0131 ,
		_w1310_,
		_w1516_,
		_w1537_,
		_w5706_
	);
	LUT4 #(
		.INIT('h08c8)
	) name5244 (
		\P2_reg1_reg[8]/NET0131 ,
		_w1191_,
		_w1507_,
		_w4672_,
		_w5707_
	);
	LUT2 #(
		.INIT('h8)
	) name5245 (
		_w1516_,
		_w5631_,
		_w5708_
	);
	LUT3 #(
		.INIT('ha2)
	) name5246 (
		\P2_reg1_reg[8]/NET0131 ,
		_w1684_,
		_w2469_,
		_w5709_
	);
	LUT2 #(
		.INIT('h1)
	) name5247 (
		_w5708_,
		_w5709_,
		_w5710_
	);
	LUT4 #(
		.INIT('h0e00)
	) name5248 (
		_w1575_,
		_w5706_,
		_w5707_,
		_w5710_,
		_w5711_
	);
	LUT4 #(
		.INIT('hc355)
	) name5249 (
		\P2_reg1_reg[8]/NET0131 ,
		_w1215_,
		_w1310_,
		_w1516_,
		_w5712_
	);
	LUT4 #(
		.INIT('hc355)
	) name5250 (
		\P2_reg1_reg[8]/NET0131 ,
		_w1215_,
		_w1310_,
		_w1507_,
		_w5713_
	);
	LUT4 #(
		.INIT('hfa32)
	) name5251 (
		_w1506_,
		_w1530_,
		_w5712_,
		_w5713_,
		_w5714_
	);
	LUT4 #(
		.INIT('h3111)
	) name5252 (
		_w1359_,
		_w5705_,
		_w5711_,
		_w5714_,
		_w5715_
	);
	LUT3 #(
		.INIT('hce)
	) name5253 (
		\P1_state_reg[0]/NET0131 ,
		_w5704_,
		_w5715_,
		_w5716_
	);
	LUT2 #(
		.INIT('h2)
	) name5254 (
		\P1_reg0_reg[11]/NET0131 ,
		_w2462_,
		_w5717_
	);
	LUT4 #(
		.INIT('h2000)
	) name5255 (
		\P1_reg0_reg[11]/NET0131 ,
		_w1723_,
		_w1727_,
		_w1730_,
		_w5718_
	);
	LUT2 #(
		.INIT('h2)
	) name5256 (
		\P1_reg0_reg[11]/NET0131 ,
		_w2883_,
		_w5719_
	);
	LUT4 #(
		.INIT('hb040)
	) name5257 (
		_w2654_,
		_w2655_,
		_w2883_,
		_w3191_,
		_w5720_
	);
	LUT3 #(
		.INIT('ha8)
	) name5258 (
		_w2292_,
		_w5719_,
		_w5720_,
		_w5721_
	);
	LUT4 #(
		.INIT('h40b0)
	) name5259 (
		_w2667_,
		_w2668_,
		_w2883_,
		_w3191_,
		_w5722_
	);
	LUT3 #(
		.INIT('ha8)
	) name5260 (
		_w2388_,
		_w5719_,
		_w5722_,
		_w5723_
	);
	LUT4 #(
		.INIT('hddd1)
	) name5261 (
		\P1_reg0_reg[11]/NET0131 ,
		_w2883_,
		_w4536_,
		_w4537_,
		_w5724_
	);
	LUT2 #(
		.INIT('h2)
	) name5262 (
		\P1_reg0_reg[11]/NET0131 ,
		_w3420_,
		_w5725_
	);
	LUT3 #(
		.INIT('h0d)
	) name5263 (
		_w2883_,
		_w5287_,
		_w5725_,
		_w5726_
	);
	LUT3 #(
		.INIT('hd0)
	) name5264 (
		_w2424_,
		_w5724_,
		_w5726_,
		_w5727_
	);
	LUT4 #(
		.INIT('ha8aa)
	) name5265 (
		_w1731_,
		_w5721_,
		_w5723_,
		_w5727_,
		_w5728_
	);
	LUT4 #(
		.INIT('heeec)
	) name5266 (
		\P1_state_reg[0]/NET0131 ,
		_w5717_,
		_w5718_,
		_w5728_,
		_w5729_
	);
	LUT4 #(
		.INIT('hd070)
	) name5267 (
		\P1_state_reg[0]/NET0131 ,
		\P2_IR_reg[23]/NET0131 ,
		\P2_reg2_reg[5]/NET0131 ,
		_w1188_,
		_w5730_
	);
	LUT4 #(
		.INIT('h2000)
	) name5268 (
		\P2_reg2_reg[5]/NET0131 ,
		_w1189_,
		_w1352_,
		_w1356_,
		_w5731_
	);
	LUT4 #(
		.INIT('haa02)
	) name5269 (
		\P2_reg2_reg[5]/NET0131 ,
		_w1361_,
		_w1363_,
		_w1368_,
		_w5732_
	);
	LUT4 #(
		.INIT('h111d)
	) name5270 (
		\P2_reg2_reg[5]/NET0131 ,
		_w1516_,
		_w5150_,
		_w5154_,
		_w5733_
	);
	LUT2 #(
		.INIT('h2)
	) name5271 (
		_w1191_,
		_w5733_,
		_w5734_
	);
	LUT3 #(
		.INIT('ha8)
	) name5272 (
		_w1530_,
		_w5663_,
		_w5732_,
		_w5735_
	);
	LUT4 #(
		.INIT('ha8aa)
	) name5273 (
		\P2_reg2_reg[5]/NET0131 ,
		_w1361_,
		_w1363_,
		_w1368_,
		_w5736_
	);
	LUT3 #(
		.INIT('h54)
	) name5274 (
		_w1506_,
		_w5660_,
		_w5736_,
		_w5737_
	);
	LUT4 #(
		.INIT('ha900)
	) name5275 (
		_w1306_,
		_w1454_,
		_w1455_,
		_w1507_,
		_w5738_
	);
	LUT3 #(
		.INIT('ha8)
	) name5276 (
		\P2_reg2_reg[5]/NET0131 ,
		_w1441_,
		_w1523_,
		_w5739_
	);
	LUT3 #(
		.INIT('h40)
	) name5277 (
		_w765_,
		_w1229_,
		_w1232_,
		_w5740_
	);
	LUT3 #(
		.INIT('h07)
	) name5278 (
		_w1507_,
		_w5589_,
		_w5740_,
		_w5741_
	);
	LUT2 #(
		.INIT('h4)
	) name5279 (
		_w5739_,
		_w5741_,
		_w5742_
	);
	LUT4 #(
		.INIT('hab00)
	) name5280 (
		_w1575_,
		_w5736_,
		_w5738_,
		_w5742_,
		_w5743_
	);
	LUT3 #(
		.INIT('h10)
	) name5281 (
		_w5737_,
		_w5735_,
		_w5743_,
		_w5744_
	);
	LUT4 #(
		.INIT('h1311)
	) name5282 (
		_w1359_,
		_w5731_,
		_w5734_,
		_w5744_,
		_w5745_
	);
	LUT3 #(
		.INIT('hce)
	) name5283 (
		\P1_state_reg[0]/NET0131 ,
		_w5730_,
		_w5745_,
		_w5746_
	);
	LUT4 #(
		.INIT('hd070)
	) name5284 (
		\P1_state_reg[0]/NET0131 ,
		\P2_IR_reg[23]/NET0131 ,
		\P2_reg2_reg[6]/NET0131 ,
		_w1188_,
		_w5747_
	);
	LUT4 #(
		.INIT('h2000)
	) name5285 (
		\P2_reg2_reg[6]/NET0131 ,
		_w1189_,
		_w1352_,
		_w1356_,
		_w5748_
	);
	LUT4 #(
		.INIT('ha8aa)
	) name5286 (
		\P2_reg2_reg[6]/NET0131 ,
		_w1361_,
		_w1363_,
		_w1368_,
		_w5749_
	);
	LUT3 #(
		.INIT('ha8)
	) name5287 (
		\P2_reg2_reg[6]/NET0131 ,
		_w1441_,
		_w1523_,
		_w5750_
	);
	LUT3 #(
		.INIT('h40)
	) name5288 (
		_w744_,
		_w1229_,
		_w1232_,
		_w5751_
	);
	LUT3 #(
		.INIT('h07)
	) name5289 (
		_w1507_,
		_w5601_,
		_w5751_,
		_w5752_
	);
	LUT2 #(
		.INIT('h4)
	) name5290 (
		_w5750_,
		_w5752_,
		_w5753_
	);
	LUT4 #(
		.INIT('hab00)
	) name5291 (
		_w1506_,
		_w5684_,
		_w5749_,
		_w5753_,
		_w5754_
	);
	LUT4 #(
		.INIT('h4844)
	) name5292 (
		_w1322_,
		_w1507_,
		_w1534_,
		_w1535_,
		_w5755_
	);
	LUT3 #(
		.INIT('h54)
	) name5293 (
		_w1575_,
		_w5749_,
		_w5755_,
		_w5756_
	);
	LUT4 #(
		.INIT('haa02)
	) name5294 (
		\P2_reg2_reg[6]/NET0131 ,
		_w1361_,
		_w1363_,
		_w1368_,
		_w5757_
	);
	LUT3 #(
		.INIT('ha8)
	) name5295 (
		_w1530_,
		_w5681_,
		_w5757_,
		_w5758_
	);
	LUT4 #(
		.INIT('h08c8)
	) name5296 (
		\P2_reg2_reg[6]/NET0131 ,
		_w1191_,
		_w1516_,
		_w5187_,
		_w5759_
	);
	LUT4 #(
		.INIT('h0100)
	) name5297 (
		_w5758_,
		_w5759_,
		_w5756_,
		_w5754_,
		_w5760_
	);
	LUT4 #(
		.INIT('ha0a8)
	) name5298 (
		\P1_state_reg[0]/NET0131 ,
		_w1359_,
		_w5748_,
		_w5760_,
		_w5761_
	);
	LUT2 #(
		.INIT('he)
	) name5299 (
		_w5747_,
		_w5761_,
		_w5762_
	);
	LUT4 #(
		.INIT('hd070)
	) name5300 (
		\P1_state_reg[0]/NET0131 ,
		\P2_IR_reg[23]/NET0131 ,
		\P2_reg2_reg[7]/NET0131 ,
		_w1188_,
		_w5763_
	);
	LUT4 #(
		.INIT('h2000)
	) name5301 (
		\P2_reg2_reg[7]/NET0131 ,
		_w1189_,
		_w1352_,
		_w1356_,
		_w5764_
	);
	LUT4 #(
		.INIT('hc355)
	) name5302 (
		\P2_reg2_reg[7]/NET0131 ,
		_w1303_,
		_w1458_,
		_w1507_,
		_w5765_
	);
	LUT2 #(
		.INIT('h1)
	) name5303 (
		_w1575_,
		_w5765_,
		_w5766_
	);
	LUT4 #(
		.INIT('h111d)
	) name5304 (
		\P2_reg2_reg[7]/NET0131 ,
		_w1516_,
		_w5200_,
		_w5201_,
		_w5767_
	);
	LUT3 #(
		.INIT('ha8)
	) name5305 (
		\P2_reg2_reg[7]/NET0131 ,
		_w1441_,
		_w1523_,
		_w5768_
	);
	LUT3 #(
		.INIT('h40)
	) name5306 (
		_w755_,
		_w1229_,
		_w1232_,
		_w5769_
	);
	LUT3 #(
		.INIT('h07)
	) name5307 (
		_w1507_,
		_w5617_,
		_w5769_,
		_w5770_
	);
	LUT2 #(
		.INIT('h4)
	) name5308 (
		_w5768_,
		_w5770_,
		_w5771_
	);
	LUT3 #(
		.INIT('hd0)
	) name5309 (
		_w1191_,
		_w5767_,
		_w5771_,
		_w5772_
	);
	LUT4 #(
		.INIT('he020)
	) name5310 (
		\P2_reg2_reg[7]/NET0131 ,
		_w1516_,
		_w1530_,
		_w5208_,
		_w5773_
	);
	LUT4 #(
		.INIT('h3202)
	) name5311 (
		\P2_reg2_reg[7]/NET0131 ,
		_w1506_,
		_w1507_,
		_w5208_,
		_w5774_
	);
	LUT2 #(
		.INIT('h1)
	) name5312 (
		_w5773_,
		_w5774_,
		_w5775_
	);
	LUT4 #(
		.INIT('h8aaa)
	) name5313 (
		_w1359_,
		_w5766_,
		_w5772_,
		_w5775_,
		_w5776_
	);
	LUT4 #(
		.INIT('heeec)
	) name5314 (
		\P1_state_reg[0]/NET0131 ,
		_w5763_,
		_w5764_,
		_w5776_,
		_w5777_
	);
	LUT4 #(
		.INIT('hd070)
	) name5315 (
		\P1_state_reg[0]/NET0131 ,
		\P2_IR_reg[23]/NET0131 ,
		\P2_reg2_reg[8]/NET0131 ,
		_w1188_,
		_w5778_
	);
	LUT4 #(
		.INIT('h2000)
	) name5316 (
		\P2_reg2_reg[8]/NET0131 ,
		_w1189_,
		_w1352_,
		_w1356_,
		_w5779_
	);
	LUT4 #(
		.INIT('h35c5)
	) name5317 (
		\P2_reg2_reg[8]/NET0131 ,
		_w1310_,
		_w1507_,
		_w1537_,
		_w5780_
	);
	LUT4 #(
		.INIT('h08c8)
	) name5318 (
		\P2_reg2_reg[8]/NET0131 ,
		_w1191_,
		_w1516_,
		_w4672_,
		_w5781_
	);
	LUT3 #(
		.INIT('ha8)
	) name5319 (
		\P2_reg2_reg[8]/NET0131 ,
		_w1441_,
		_w1523_,
		_w5782_
	);
	LUT3 #(
		.INIT('h40)
	) name5320 (
		_w723_,
		_w1229_,
		_w1232_,
		_w5783_
	);
	LUT3 #(
		.INIT('h07)
	) name5321 (
		_w1507_,
		_w5631_,
		_w5783_,
		_w5784_
	);
	LUT2 #(
		.INIT('h4)
	) name5322 (
		_w5782_,
		_w5784_,
		_w5785_
	);
	LUT4 #(
		.INIT('h3200)
	) name5323 (
		_w1575_,
		_w5781_,
		_w5780_,
		_w5785_,
		_w5786_
	);
	LUT4 #(
		.INIT('hc355)
	) name5324 (
		\P2_reg2_reg[8]/NET0131 ,
		_w1215_,
		_w1310_,
		_w1516_,
		_w5787_
	);
	LUT4 #(
		.INIT('hc355)
	) name5325 (
		\P2_reg2_reg[8]/NET0131 ,
		_w1215_,
		_w1310_,
		_w1507_,
		_w5788_
	);
	LUT4 #(
		.INIT('hf3a2)
	) name5326 (
		_w1506_,
		_w1530_,
		_w5787_,
		_w5788_,
		_w5789_
	);
	LUT4 #(
		.INIT('h3111)
	) name5327 (
		_w1359_,
		_w5779_,
		_w5786_,
		_w5789_,
		_w5790_
	);
	LUT3 #(
		.INIT('hce)
	) name5328 (
		\P1_state_reg[0]/NET0131 ,
		_w5778_,
		_w5790_,
		_w5791_
	);
	LUT2 #(
		.INIT('h2)
	) name5329 (
		\P1_reg0_reg[14]/NET0131 ,
		_w2462_,
		_w5792_
	);
	LUT4 #(
		.INIT('h2000)
	) name5330 (
		\P1_reg0_reg[14]/NET0131 ,
		_w1723_,
		_w1727_,
		_w1730_,
		_w5793_
	);
	LUT4 #(
		.INIT('hddd1)
	) name5331 (
		\P1_reg0_reg[14]/NET0131 ,
		_w2883_,
		_w4569_,
		_w4570_,
		_w5794_
	);
	LUT2 #(
		.INIT('h2)
	) name5332 (
		_w2424_,
		_w5794_,
		_w5795_
	);
	LUT4 #(
		.INIT('hc808)
	) name5333 (
		\P1_reg0_reg[14]/NET0131 ,
		_w2292_,
		_w2883_,
		_w4575_,
		_w5796_
	);
	LUT4 #(
		.INIT('h08c8)
	) name5334 (
		\P1_reg0_reg[14]/NET0131 ,
		_w2388_,
		_w2883_,
		_w4573_,
		_w5797_
	);
	LUT4 #(
		.INIT('h0a8a)
	) name5335 (
		\P1_reg0_reg[14]/NET0131 ,
		_w2452_,
		_w2524_,
		_w2883_,
		_w5798_
	);
	LUT3 #(
		.INIT('h0d)
	) name5336 (
		_w2883_,
		_w4579_,
		_w5798_,
		_w5799_
	);
	LUT3 #(
		.INIT('h10)
	) name5337 (
		_w5797_,
		_w5796_,
		_w5799_,
		_w5800_
	);
	LUT4 #(
		.INIT('h1311)
	) name5338 (
		_w1731_,
		_w5793_,
		_w5795_,
		_w5800_,
		_w5801_
	);
	LUT3 #(
		.INIT('hce)
	) name5339 (
		\P1_state_reg[0]/NET0131 ,
		_w5792_,
		_w5801_,
		_w5802_
	);
	LUT2 #(
		.INIT('h2)
	) name5340 (
		\P1_reg0_reg[5]/NET0131 ,
		_w2462_,
		_w5803_
	);
	LUT2 #(
		.INIT('h2)
	) name5341 (
		\P1_reg0_reg[5]/NET0131 ,
		_w2883_,
		_w5804_
	);
	LUT4 #(
		.INIT('h7020)
	) name5342 (
		_w1747_,
		_w2053_,
		_w2883_,
		_w5130_,
		_w5805_
	);
	LUT3 #(
		.INIT('ha8)
	) name5343 (
		_w2424_,
		_w5804_,
		_w5805_,
		_w5806_
	);
	LUT4 #(
		.INIT('hc535)
	) name5344 (
		\P1_reg0_reg[5]/NET0131 ,
		_w2096_,
		_w2883_,
		_w3187_,
		_w5807_
	);
	LUT2 #(
		.INIT('h2)
	) name5345 (
		_w2292_,
		_w5807_,
		_w5808_
	);
	LUT4 #(
		.INIT('h1dd1)
	) name5346 (
		\P1_reg0_reg[5]/NET0131 ,
		_w2883_,
		_w3187_,
		_w5135_,
		_w5809_
	);
	LUT4 #(
		.INIT('h0a8a)
	) name5347 (
		\P1_reg0_reg[5]/NET0131 ,
		_w2452_,
		_w2524_,
		_w2883_,
		_w5810_
	);
	LUT4 #(
		.INIT('h0057)
	) name5348 (
		_w2883_,
		_w5137_,
		_w5556_,
		_w5810_,
		_w5811_
	);
	LUT3 #(
		.INIT('hd0)
	) name5349 (
		_w2388_,
		_w5809_,
		_w5811_,
		_w5812_
	);
	LUT4 #(
		.INIT('ha8aa)
	) name5350 (
		_w1731_,
		_w5806_,
		_w5808_,
		_w5812_,
		_w5813_
	);
	LUT4 #(
		.INIT('h2000)
	) name5351 (
		\P1_reg0_reg[5]/NET0131 ,
		_w1723_,
		_w1727_,
		_w1730_,
		_w5814_
	);
	LUT4 #(
		.INIT('heeec)
	) name5352 (
		\P1_state_reg[0]/NET0131 ,
		_w5803_,
		_w5813_,
		_w5814_,
		_w5815_
	);
	LUT2 #(
		.INIT('h2)
	) name5353 (
		\P1_reg1_reg[11]/NET0131 ,
		_w2462_,
		_w5816_
	);
	LUT4 #(
		.INIT('h2000)
	) name5354 (
		\P1_reg1_reg[11]/NET0131 ,
		_w1723_,
		_w1727_,
		_w1730_,
		_w5817_
	);
	LUT2 #(
		.INIT('h2)
	) name5355 (
		\P1_reg1_reg[11]/NET0131 ,
		_w2520_,
		_w5818_
	);
	LUT4 #(
		.INIT('h8a20)
	) name5356 (
		_w2520_,
		_w2654_,
		_w2655_,
		_w3191_,
		_w5819_
	);
	LUT3 #(
		.INIT('ha8)
	) name5357 (
		_w2292_,
		_w5818_,
		_w5819_,
		_w5820_
	);
	LUT4 #(
		.INIT('h208a)
	) name5358 (
		_w2520_,
		_w2667_,
		_w2668_,
		_w3191_,
		_w5821_
	);
	LUT3 #(
		.INIT('ha8)
	) name5359 (
		_w2388_,
		_w5818_,
		_w5821_,
		_w5822_
	);
	LUT4 #(
		.INIT('hddd1)
	) name5360 (
		\P1_reg1_reg[11]/NET0131 ,
		_w2520_,
		_w4536_,
		_w4537_,
		_w5823_
	);
	LUT4 #(
		.INIT('h08aa)
	) name5361 (
		\P1_reg1_reg[11]/NET0131 ,
		_w2452_,
		_w2520_,
		_w2524_,
		_w5824_
	);
	LUT3 #(
		.INIT('h0d)
	) name5362 (
		_w2520_,
		_w5287_,
		_w5824_,
		_w5825_
	);
	LUT3 #(
		.INIT('hd0)
	) name5363 (
		_w2424_,
		_w5823_,
		_w5825_,
		_w5826_
	);
	LUT4 #(
		.INIT('ha8aa)
	) name5364 (
		_w1731_,
		_w5820_,
		_w5822_,
		_w5826_,
		_w5827_
	);
	LUT4 #(
		.INIT('heeec)
	) name5365 (
		\P1_state_reg[0]/NET0131 ,
		_w5816_,
		_w5817_,
		_w5827_,
		_w5828_
	);
	LUT2 #(
		.INIT('h2)
	) name5366 (
		\P1_reg1_reg[14]/NET0131 ,
		_w2462_,
		_w5829_
	);
	LUT4 #(
		.INIT('h2000)
	) name5367 (
		\P1_reg1_reg[14]/NET0131 ,
		_w1723_,
		_w1727_,
		_w1730_,
		_w5830_
	);
	LUT4 #(
		.INIT('hddd1)
	) name5368 (
		\P1_reg1_reg[14]/NET0131 ,
		_w2520_,
		_w4569_,
		_w4570_,
		_w5831_
	);
	LUT2 #(
		.INIT('h2)
	) name5369 (
		_w2424_,
		_w5831_,
		_w5832_
	);
	LUT4 #(
		.INIT('h08c8)
	) name5370 (
		\P1_reg1_reg[14]/NET0131 ,
		_w2388_,
		_w2520_,
		_w4573_,
		_w5833_
	);
	LUT4 #(
		.INIT('hc808)
	) name5371 (
		\P1_reg1_reg[14]/NET0131 ,
		_w2292_,
		_w2520_,
		_w4575_,
		_w5834_
	);
	LUT4 #(
		.INIT('h08aa)
	) name5372 (
		\P1_reg1_reg[14]/NET0131 ,
		_w2452_,
		_w2520_,
		_w2524_,
		_w5835_
	);
	LUT3 #(
		.INIT('h0d)
	) name5373 (
		_w2520_,
		_w4579_,
		_w5835_,
		_w5836_
	);
	LUT3 #(
		.INIT('h10)
	) name5374 (
		_w5834_,
		_w5833_,
		_w5836_,
		_w5837_
	);
	LUT4 #(
		.INIT('h1311)
	) name5375 (
		_w1731_,
		_w5830_,
		_w5832_,
		_w5837_,
		_w5838_
	);
	LUT3 #(
		.INIT('hce)
	) name5376 (
		\P1_state_reg[0]/NET0131 ,
		_w5829_,
		_w5838_,
		_w5839_
	);
	LUT4 #(
		.INIT('h1000)
	) name5377 (
		\P2_reg3_reg[3]/NET0131 ,
		_w1189_,
		_w1352_,
		_w1356_,
		_w5840_
	);
	LUT2 #(
		.INIT('h1)
	) name5378 (
		_w803_,
		_w1435_,
		_w5841_
	);
	LUT4 #(
		.INIT('h007b)
	) name5379 (
		_w781_,
		_w1435_,
		_w5151_,
		_w5841_,
		_w5842_
	);
	LUT4 #(
		.INIT('h04c4)
	) name5380 (
		\P2_reg3_reg[3]/NET0131 ,
		_w1191_,
		_w1411_,
		_w5842_,
		_w5843_
	);
	LUT4 #(
		.INIT('h54ab)
	) name5381 (
		_w808_,
		_w828_,
		_w1210_,
		_w1326_,
		_w5844_
	);
	LUT4 #(
		.INIT('h1e78)
	) name5382 (
		_w803_,
		_w807_,
		_w1326_,
		_w1452_,
		_w5845_
	);
	LUT4 #(
		.INIT('ha8fc)
	) name5383 (
		_w1409_,
		_w1496_,
		_w5845_,
		_w5844_,
		_w5846_
	);
	LUT4 #(
		.INIT('h04c4)
	) name5384 (
		\P2_reg3_reg[3]/NET0131 ,
		_w1447_,
		_w1411_,
		_w5845_,
		_w5847_
	);
	LUT3 #(
		.INIT('h04)
	) name5385 (
		_w797_,
		_w1232_,
		_w1439_,
		_w5848_
	);
	LUT4 #(
		.INIT('h008f)
	) name5386 (
		_w1179_,
		_w1183_,
		_w1228_,
		_w1338_,
		_w5849_
	);
	LUT4 #(
		.INIT('h001f)
	) name5387 (
		_w1361_,
		_w1363_,
		_w1368_,
		_w5849_,
		_w5850_
	);
	LUT4 #(
		.INIT('h5554)
	) name5388 (
		\P2_reg3_reg[3]/NET0131 ,
		_w1441_,
		_w1443_,
		_w5850_,
		_w5851_
	);
	LUT2 #(
		.INIT('h1)
	) name5389 (
		_w5848_,
		_w5851_,
		_w5852_
	);
	LUT4 #(
		.INIT('h3100)
	) name5390 (
		_w1369_,
		_w5847_,
		_w5846_,
		_w5852_,
		_w5853_
	);
	LUT4 #(
		.INIT('h1311)
	) name5391 (
		_w1359_,
		_w5840_,
		_w5843_,
		_w5853_,
		_w5854_
	);
	LUT2 #(
		.INIT('h4)
	) name5392 (
		\P1_state_reg[0]/NET0131 ,
		\P2_reg3_reg[3]/NET0131 ,
		_w5855_
	);
	LUT4 #(
		.INIT('ha7ad)
	) name5393 (
		\P1_state_reg[0]/NET0131 ,
		\P2_IR_reg[23]/NET0131 ,
		\P2_reg3_reg[3]/NET0131 ,
		_w1188_,
		_w5856_
	);
	LUT3 #(
		.INIT('h2f)
	) name5394 (
		\P1_state_reg[0]/NET0131 ,
		_w5854_,
		_w5856_,
		_w5857_
	);
	LUT2 #(
		.INIT('h2)
	) name5395 (
		\P1_reg1_reg[3]/NET0131 ,
		_w2520_,
		_w5858_
	);
	LUT4 #(
		.INIT('hc808)
	) name5396 (
		\P1_reg1_reg[3]/NET0131 ,
		_w2424_,
		_w2520_,
		_w5480_,
		_w5859_
	);
	LUT4 #(
		.INIT('he010)
	) name5397 (
		_w2066_,
		_w2092_,
		_w2520_,
		_w3188_,
		_w5860_
	);
	LUT3 #(
		.INIT('ha8)
	) name5398 (
		_w2292_,
		_w5858_,
		_w5860_,
		_w5861_
	);
	LUT4 #(
		.INIT('h10e0)
	) name5399 (
		_w2307_,
		_w2308_,
		_w2520_,
		_w3188_,
		_w5862_
	);
	LUT2 #(
		.INIT('h4)
	) name5400 (
		_w2071_,
		_w2426_,
		_w5863_
	);
	LUT4 #(
		.INIT('h009f)
	) name5401 (
		_w2071_,
		_w2428_,
		_w2447_,
		_w5863_,
		_w5864_
	);
	LUT4 #(
		.INIT('hf531)
	) name5402 (
		\P1_reg1_reg[3]/NET0131 ,
		_w2520_,
		_w2525_,
		_w5864_,
		_w5865_
	);
	LUT4 #(
		.INIT('h5700)
	) name5403 (
		_w2388_,
		_w5858_,
		_w5862_,
		_w5865_,
		_w5866_
	);
	LUT4 #(
		.INIT('ha8aa)
	) name5404 (
		_w1731_,
		_w5859_,
		_w5861_,
		_w5866_,
		_w5867_
	);
	LUT4 #(
		.INIT('h2000)
	) name5405 (
		\P1_reg1_reg[3]/NET0131 ,
		_w1723_,
		_w1727_,
		_w1730_,
		_w5868_
	);
	LUT2 #(
		.INIT('h2)
	) name5406 (
		\P1_reg1_reg[3]/NET0131 ,
		_w2462_,
		_w5869_
	);
	LUT4 #(
		.INIT('hffa8)
	) name5407 (
		\P1_state_reg[0]/NET0131 ,
		_w5867_,
		_w5868_,
		_w5869_,
		_w5870_
	);
	LUT2 #(
		.INIT('h2)
	) name5408 (
		\P1_reg1_reg[7]/NET0131 ,
		_w2520_,
		_w5871_
	);
	LUT4 #(
		.INIT('hddd1)
	) name5409 (
		\P1_reg1_reg[7]/NET0131 ,
		_w2520_,
		_w5513_,
		_w5514_,
		_w5872_
	);
	LUT4 #(
		.INIT('hc808)
	) name5410 (
		\P1_reg1_reg[7]/NET0131 ,
		_w2292_,
		_w2520_,
		_w5516_,
		_w5873_
	);
	LUT4 #(
		.INIT('he010)
	) name5411 (
		_w2316_,
		_w2320_,
		_w2520_,
		_w3183_,
		_w5874_
	);
	LUT2 #(
		.INIT('h2)
	) name5412 (
		\P1_reg1_reg[7]/NET0131 ,
		_w2525_,
		_w5875_
	);
	LUT2 #(
		.INIT('h8)
	) name5413 (
		_w2114_,
		_w2426_,
		_w5876_
	);
	LUT4 #(
		.INIT('h00fb)
	) name5414 (
		_w2431_,
		_w2447_,
		_w5519_,
		_w5876_,
		_w5877_
	);
	LUT3 #(
		.INIT('h31)
	) name5415 (
		_w2520_,
		_w5875_,
		_w5877_,
		_w5878_
	);
	LUT4 #(
		.INIT('h5700)
	) name5416 (
		_w2388_,
		_w5871_,
		_w5874_,
		_w5878_,
		_w5879_
	);
	LUT4 #(
		.INIT('h0d00)
	) name5417 (
		_w2424_,
		_w5872_,
		_w5873_,
		_w5879_,
		_w5880_
	);
	LUT4 #(
		.INIT('h2000)
	) name5418 (
		\P1_reg1_reg[7]/NET0131 ,
		_w1723_,
		_w1727_,
		_w1730_,
		_w5881_
	);
	LUT4 #(
		.INIT('haa08)
	) name5419 (
		\P1_state_reg[0]/NET0131 ,
		_w1731_,
		_w5880_,
		_w5881_,
		_w5882_
	);
	LUT2 #(
		.INIT('h2)
	) name5420 (
		\P1_reg1_reg[7]/NET0131 ,
		_w2462_,
		_w5883_
	);
	LUT2 #(
		.INIT('he)
	) name5421 (
		_w5882_,
		_w5883_,
		_w5884_
	);
	LUT2 #(
		.INIT('h2)
	) name5422 (
		\P1_reg2_reg[3]/NET0131 ,
		_w1741_,
		_w5885_
	);
	LUT4 #(
		.INIT('he020)
	) name5423 (
		\P1_reg2_reg[3]/NET0131 ,
		_w1741_,
		_w2424_,
		_w5480_,
		_w5886_
	);
	LUT4 #(
		.INIT('ha802)
	) name5424 (
		_w1741_,
		_w2066_,
		_w2092_,
		_w3188_,
		_w5887_
	);
	LUT3 #(
		.INIT('ha8)
	) name5425 (
		_w2292_,
		_w5885_,
		_w5887_,
		_w5888_
	);
	LUT4 #(
		.INIT('h02a8)
	) name5426 (
		_w1741_,
		_w2307_,
		_w2308_,
		_w3188_,
		_w5889_
	);
	LUT4 #(
		.INIT('ha2a0)
	) name5427 (
		\P1_reg2_reg[3]/NET0131 ,
		_w1741_,
		_w2450_,
		_w2452_,
		_w5890_
	);
	LUT4 #(
		.INIT('h0004)
	) name5428 (
		\P1_reg3_reg[3]/NET0131 ,
		_w2284_,
		_w2288_,
		_w2291_,
		_w5891_
	);
	LUT4 #(
		.INIT('h000d)
	) name5429 (
		_w1741_,
		_w5864_,
		_w5890_,
		_w5891_,
		_w5892_
	);
	LUT4 #(
		.INIT('h5700)
	) name5430 (
		_w2388_,
		_w5885_,
		_w5889_,
		_w5892_,
		_w5893_
	);
	LUT4 #(
		.INIT('ha8aa)
	) name5431 (
		_w1731_,
		_w5886_,
		_w5888_,
		_w5893_,
		_w5894_
	);
	LUT4 #(
		.INIT('h2000)
	) name5432 (
		\P1_reg2_reg[3]/NET0131 ,
		_w1723_,
		_w1727_,
		_w1730_,
		_w5895_
	);
	LUT2 #(
		.INIT('h2)
	) name5433 (
		\P1_reg2_reg[3]/NET0131 ,
		_w2462_,
		_w5896_
	);
	LUT4 #(
		.INIT('hffa8)
	) name5434 (
		\P1_state_reg[0]/NET0131 ,
		_w5894_,
		_w5895_,
		_w5896_,
		_w5897_
	);
	LUT2 #(
		.INIT('h2)
	) name5435 (
		\P1_reg2_reg[6]/NET0131 ,
		_w2462_,
		_w5898_
	);
	LUT4 #(
		.INIT('h2000)
	) name5436 (
		\P1_reg2_reg[6]/NET0131 ,
		_w1723_,
		_w1727_,
		_w1730_,
		_w5899_
	);
	LUT2 #(
		.INIT('h2)
	) name5437 (
		\P1_reg2_reg[6]/NET0131 ,
		_w1741_,
		_w5900_
	);
	LUT4 #(
		.INIT('he020)
	) name5438 (
		\P1_reg2_reg[6]/NET0131 ,
		_w1741_,
		_w2424_,
		_w5496_,
		_w5901_
	);
	LUT4 #(
		.INIT('h02a8)
	) name5439 (
		_w1741_,
		_w2749_,
		_w2750_,
		_w3182_,
		_w5902_
	);
	LUT3 #(
		.INIT('ha8)
	) name5440 (
		_w2292_,
		_w5900_,
		_w5902_,
		_w5903_
	);
	LUT4 #(
		.INIT('ha802)
	) name5441 (
		_w1741_,
		_w2797_,
		_w2932_,
		_w3182_,
		_w5904_
	);
	LUT4 #(
		.INIT('he020)
	) name5442 (
		\P1_reg2_reg[6]/NET0131 ,
		_w1741_,
		_w2447_,
		_w5501_,
		_w5905_
	);
	LUT4 #(
		.INIT('haa20)
	) name5443 (
		\P1_reg2_reg[6]/NET0131 ,
		_w1741_,
		_w2426_,
		_w2450_,
		_w5906_
	);
	LUT4 #(
		.INIT('h0008)
	) name5444 (
		_w2126_,
		_w2284_,
		_w2288_,
		_w2291_,
		_w5907_
	);
	LUT2 #(
		.INIT('h4)
	) name5445 (
		_w2124_,
		_w2426_,
		_w5908_
	);
	LUT3 #(
		.INIT('h13)
	) name5446 (
		_w1741_,
		_w5907_,
		_w5908_,
		_w5909_
	);
	LUT2 #(
		.INIT('h4)
	) name5447 (
		_w5906_,
		_w5909_,
		_w5910_
	);
	LUT2 #(
		.INIT('h4)
	) name5448 (
		_w5905_,
		_w5910_,
		_w5911_
	);
	LUT4 #(
		.INIT('h5700)
	) name5449 (
		_w2388_,
		_w5900_,
		_w5904_,
		_w5911_,
		_w5912_
	);
	LUT4 #(
		.INIT('ha8aa)
	) name5450 (
		_w1731_,
		_w5903_,
		_w5901_,
		_w5912_,
		_w5913_
	);
	LUT4 #(
		.INIT('heeec)
	) name5451 (
		\P1_state_reg[0]/NET0131 ,
		_w5898_,
		_w5899_,
		_w5913_,
		_w5914_
	);
	LUT2 #(
		.INIT('h2)
	) name5452 (
		\P1_reg2_reg[7]/NET0131 ,
		_w1741_,
		_w5915_
	);
	LUT4 #(
		.INIT('hddd1)
	) name5453 (
		\P1_reg2_reg[7]/NET0131 ,
		_w1741_,
		_w5513_,
		_w5514_,
		_w5916_
	);
	LUT4 #(
		.INIT('he020)
	) name5454 (
		\P1_reg2_reg[7]/NET0131 ,
		_w1741_,
		_w2292_,
		_w5516_,
		_w5917_
	);
	LUT4 #(
		.INIT('ha802)
	) name5455 (
		_w1741_,
		_w2316_,
		_w2320_,
		_w3183_,
		_w5918_
	);
	LUT4 #(
		.INIT('h0008)
	) name5456 (
		_w2115_,
		_w2284_,
		_w2288_,
		_w2291_,
		_w5919_
	);
	LUT4 #(
		.INIT('ha2a0)
	) name5457 (
		\P1_reg2_reg[7]/NET0131 ,
		_w1741_,
		_w2450_,
		_w2452_,
		_w5920_
	);
	LUT2 #(
		.INIT('h1)
	) name5458 (
		_w5919_,
		_w5920_,
		_w5921_
	);
	LUT3 #(
		.INIT('hd0)
	) name5459 (
		_w1741_,
		_w5877_,
		_w5921_,
		_w5922_
	);
	LUT4 #(
		.INIT('h5700)
	) name5460 (
		_w2388_,
		_w5915_,
		_w5918_,
		_w5922_,
		_w5923_
	);
	LUT4 #(
		.INIT('h0d00)
	) name5461 (
		_w2424_,
		_w5916_,
		_w5917_,
		_w5923_,
		_w5924_
	);
	LUT4 #(
		.INIT('h2000)
	) name5462 (
		\P1_reg2_reg[7]/NET0131 ,
		_w1723_,
		_w1727_,
		_w1730_,
		_w5925_
	);
	LUT4 #(
		.INIT('haa08)
	) name5463 (
		\P1_state_reg[0]/NET0131 ,
		_w1731_,
		_w5924_,
		_w5925_,
		_w5926_
	);
	LUT2 #(
		.INIT('h2)
	) name5464 (
		\P1_reg2_reg[7]/NET0131 ,
		_w2462_,
		_w5927_
	);
	LUT2 #(
		.INIT('he)
	) name5465 (
		_w5926_,
		_w5927_,
		_w5928_
	);
	LUT2 #(
		.INIT('h2)
	) name5466 (
		\P1_reg0_reg[3]/NET0131 ,
		_w2462_,
		_w5929_
	);
	LUT2 #(
		.INIT('h2)
	) name5467 (
		\P1_reg0_reg[3]/NET0131 ,
		_w2883_,
		_w5930_
	);
	LUT4 #(
		.INIT('hc808)
	) name5468 (
		\P1_reg0_reg[3]/NET0131 ,
		_w2424_,
		_w2883_,
		_w5480_,
		_w5931_
	);
	LUT4 #(
		.INIT('he010)
	) name5469 (
		_w2066_,
		_w2092_,
		_w2883_,
		_w3188_,
		_w5932_
	);
	LUT3 #(
		.INIT('ha8)
	) name5470 (
		_w2292_,
		_w5930_,
		_w5932_,
		_w5933_
	);
	LUT4 #(
		.INIT('h10e0)
	) name5471 (
		_w2307_,
		_w2308_,
		_w2883_,
		_w3188_,
		_w5934_
	);
	LUT4 #(
		.INIT('h0a8a)
	) name5472 (
		\P1_reg0_reg[3]/NET0131 ,
		_w2452_,
		_w2524_,
		_w2883_,
		_w5935_
	);
	LUT3 #(
		.INIT('h0d)
	) name5473 (
		_w2883_,
		_w5864_,
		_w5935_,
		_w5936_
	);
	LUT4 #(
		.INIT('h5700)
	) name5474 (
		_w2388_,
		_w5930_,
		_w5934_,
		_w5936_,
		_w5937_
	);
	LUT4 #(
		.INIT('ha8aa)
	) name5475 (
		_w1731_,
		_w5931_,
		_w5933_,
		_w5937_,
		_w5938_
	);
	LUT4 #(
		.INIT('h2000)
	) name5476 (
		\P1_reg0_reg[3]/NET0131 ,
		_w1723_,
		_w1727_,
		_w1730_,
		_w5939_
	);
	LUT4 #(
		.INIT('heeec)
	) name5477 (
		\P1_state_reg[0]/NET0131 ,
		_w5929_,
		_w5938_,
		_w5939_,
		_w5940_
	);
	LUT2 #(
		.INIT('h2)
	) name5478 (
		\P1_reg0_reg[7]/NET0131 ,
		_w2462_,
		_w5941_
	);
	LUT2 #(
		.INIT('h2)
	) name5479 (
		\P1_reg0_reg[7]/NET0131 ,
		_w2883_,
		_w5942_
	);
	LUT4 #(
		.INIT('hddd1)
	) name5480 (
		\P1_reg0_reg[7]/NET0131 ,
		_w2883_,
		_w5513_,
		_w5514_,
		_w5943_
	);
	LUT4 #(
		.INIT('hc808)
	) name5481 (
		\P1_reg0_reg[7]/NET0131 ,
		_w2292_,
		_w2883_,
		_w5516_,
		_w5944_
	);
	LUT4 #(
		.INIT('he010)
	) name5482 (
		_w2316_,
		_w2320_,
		_w2883_,
		_w3183_,
		_w5945_
	);
	LUT4 #(
		.INIT('h0a8a)
	) name5483 (
		\P1_reg0_reg[7]/NET0131 ,
		_w2452_,
		_w2524_,
		_w2883_,
		_w5946_
	);
	LUT3 #(
		.INIT('h0d)
	) name5484 (
		_w2883_,
		_w5877_,
		_w5946_,
		_w5947_
	);
	LUT4 #(
		.INIT('h5700)
	) name5485 (
		_w2388_,
		_w5942_,
		_w5945_,
		_w5947_,
		_w5948_
	);
	LUT4 #(
		.INIT('h0d00)
	) name5486 (
		_w2424_,
		_w5943_,
		_w5944_,
		_w5948_,
		_w5949_
	);
	LUT4 #(
		.INIT('h2000)
	) name5487 (
		\P1_reg0_reg[7]/NET0131 ,
		_w1723_,
		_w1727_,
		_w1730_,
		_w5950_
	);
	LUT4 #(
		.INIT('haa08)
	) name5488 (
		\P1_state_reg[0]/NET0131 ,
		_w1731_,
		_w5949_,
		_w5950_,
		_w5951_
	);
	LUT2 #(
		.INIT('he)
	) name5489 (
		_w5941_,
		_w5951_,
		_w5952_
	);
	LUT4 #(
		.INIT('hd070)
	) name5490 (
		\P1_state_reg[0]/NET0131 ,
		\P2_IR_reg[23]/NET0131 ,
		\P2_reg3_reg[2]/NET0131 ,
		_w1188_,
		_w5953_
	);
	LUT4 #(
		.INIT('h2000)
	) name5491 (
		\P2_reg3_reg[2]/NET0131 ,
		_w1189_,
		_w1352_,
		_w1356_,
		_w5954_
	);
	LUT4 #(
		.INIT('h6500)
	) name5492 (
		_w792_,
		_w803_,
		_w1414_,
		_w1435_,
		_w5955_
	);
	LUT2 #(
		.INIT('h1)
	) name5493 (
		_w814_,
		_w1435_,
		_w5956_
	);
	LUT4 #(
		.INIT('h111d)
	) name5494 (
		\P2_reg3_reg[2]/NET0131 ,
		_w1411_,
		_w5955_,
		_w5956_,
		_w5957_
	);
	LUT4 #(
		.INIT('hc355)
	) name5495 (
		\P2_reg3_reg[2]/NET0131 ,
		_w1210_,
		_w1321_,
		_w1369_,
		_w5958_
	);
	LUT3 #(
		.INIT('ha8)
	) name5496 (
		\P2_reg3_reg[2]/NET0131 ,
		_w1441_,
		_w1443_,
		_w5959_
	);
	LUT3 #(
		.INIT('h04)
	) name5497 (
		_w807_,
		_w1232_,
		_w1439_,
		_w5960_
	);
	LUT4 #(
		.INIT('h0032)
	) name5498 (
		_w1409_,
		_w5959_,
		_w5958_,
		_w5960_,
		_w5961_
	);
	LUT4 #(
		.INIT('hc535)
	) name5499 (
		\P2_reg3_reg[2]/NET0131 ,
		_w1321_,
		_w1411_,
		_w1452_,
		_w5962_
	);
	LUT4 #(
		.INIT('hc535)
	) name5500 (
		\P2_reg3_reg[2]/NET0131 ,
		_w1321_,
		_w1369_,
		_w1452_,
		_w5963_
	);
	LUT4 #(
		.INIT('hf5c4)
	) name5501 (
		_w1447_,
		_w1496_,
		_w5962_,
		_w5963_,
		_w5964_
	);
	LUT4 #(
		.INIT('hd000)
	) name5502 (
		_w1191_,
		_w5957_,
		_w5961_,
		_w5964_,
		_w5965_
	);
	LUT4 #(
		.INIT('ha0a8)
	) name5503 (
		\P1_state_reg[0]/NET0131 ,
		_w1359_,
		_w5954_,
		_w5965_,
		_w5966_
	);
	LUT2 #(
		.INIT('he)
	) name5504 (
		_w5953_,
		_w5966_,
		_w5967_
	);
	LUT2 #(
		.INIT('h2)
	) name5505 (
		\P1_reg1_reg[6]/NET0131 ,
		_w2462_,
		_w5968_
	);
	LUT4 #(
		.INIT('h2000)
	) name5506 (
		\P1_reg1_reg[6]/NET0131 ,
		_w1723_,
		_w1727_,
		_w1730_,
		_w5969_
	);
	LUT2 #(
		.INIT('h2)
	) name5507 (
		\P1_reg1_reg[6]/NET0131 ,
		_w2520_,
		_w5970_
	);
	LUT4 #(
		.INIT('hc808)
	) name5508 (
		\P1_reg1_reg[6]/NET0131 ,
		_w2424_,
		_w2520_,
		_w5496_,
		_w5971_
	);
	LUT4 #(
		.INIT('ha802)
	) name5509 (
		_w2520_,
		_w2797_,
		_w2932_,
		_w3182_,
		_w5972_
	);
	LUT3 #(
		.INIT('ha8)
	) name5510 (
		_w2388_,
		_w5970_,
		_w5972_,
		_w5973_
	);
	LUT4 #(
		.INIT('h02a8)
	) name5511 (
		_w2520_,
		_w2749_,
		_w2750_,
		_w3182_,
		_w5974_
	);
	LUT4 #(
		.INIT('hc808)
	) name5512 (
		\P1_reg1_reg[6]/NET0131 ,
		_w2447_,
		_w2520_,
		_w5501_,
		_w5975_
	);
	LUT2 #(
		.INIT('h8)
	) name5513 (
		_w2520_,
		_w5908_,
		_w5976_
	);
	LUT4 #(
		.INIT('h08aa)
	) name5514 (
		\P1_reg1_reg[6]/NET0131 ,
		_w2426_,
		_w2520_,
		_w2524_,
		_w5977_
	);
	LUT2 #(
		.INIT('h1)
	) name5515 (
		_w5976_,
		_w5977_,
		_w5978_
	);
	LUT2 #(
		.INIT('h4)
	) name5516 (
		_w5975_,
		_w5978_,
		_w5979_
	);
	LUT4 #(
		.INIT('h5700)
	) name5517 (
		_w2292_,
		_w5970_,
		_w5974_,
		_w5979_,
		_w5980_
	);
	LUT4 #(
		.INIT('ha8aa)
	) name5518 (
		_w1731_,
		_w5973_,
		_w5971_,
		_w5980_,
		_w5981_
	);
	LUT4 #(
		.INIT('heeec)
	) name5519 (
		\P1_state_reg[0]/NET0131 ,
		_w5968_,
		_w5969_,
		_w5981_,
		_w5982_
	);
	LUT4 #(
		.INIT('hd070)
	) name5520 (
		\P1_state_reg[0]/NET0131 ,
		\P2_IR_reg[23]/NET0131 ,
		\P2_reg0_reg[3]/NET0131 ,
		_w1188_,
		_w5983_
	);
	LUT4 #(
		.INIT('h2000)
	) name5521 (
		\P2_reg0_reg[3]/NET0131 ,
		_w1189_,
		_w1352_,
		_w1356_,
		_w5984_
	);
	LUT4 #(
		.INIT('h0155)
	) name5522 (
		\P2_reg0_reg[3]/NET0131 ,
		_w1361_,
		_w1363_,
		_w1368_,
		_w5985_
	);
	LUT2 #(
		.INIT('h2)
	) name5523 (
		_w1191_,
		_w5985_,
		_w5986_
	);
	LUT3 #(
		.INIT('h70)
	) name5524 (
		_w1369_,
		_w5842_,
		_w5986_,
		_w5987_
	);
	LUT4 #(
		.INIT('h3202)
	) name5525 (
		\P2_reg0_reg[3]/NET0131 ,
		_w1409_,
		_w1411_,
		_w5844_,
		_w5988_
	);
	LUT4 #(
		.INIT('h020e)
	) name5526 (
		\P2_reg0_reg[3]/NET0131 ,
		_w1411_,
		_w1496_,
		_w5845_,
		_w5989_
	);
	LUT2 #(
		.INIT('h2)
	) name5527 (
		_w1447_,
		_w5985_,
		_w5990_
	);
	LUT3 #(
		.INIT('h70)
	) name5528 (
		_w1369_,
		_w5845_,
		_w5990_,
		_w5991_
	);
	LUT2 #(
		.INIT('h4)
	) name5529 (
		_w797_,
		_w1442_,
		_w5992_
	);
	LUT2 #(
		.INIT('h8)
	) name5530 (
		_w1411_,
		_w5992_,
		_w5993_
	);
	LUT3 #(
		.INIT('ha2)
	) name5531 (
		\P2_reg0_reg[3]/NET0131 ,
		_w1684_,
		_w1685_,
		_w5994_
	);
	LUT2 #(
		.INIT('h1)
	) name5532 (
		_w5993_,
		_w5994_,
		_w5995_
	);
	LUT4 #(
		.INIT('h0100)
	) name5533 (
		_w5989_,
		_w5988_,
		_w5991_,
		_w5995_,
		_w5996_
	);
	LUT4 #(
		.INIT('h1311)
	) name5534 (
		_w1359_,
		_w5984_,
		_w5987_,
		_w5996_,
		_w5997_
	);
	LUT3 #(
		.INIT('hce)
	) name5535 (
		\P1_state_reg[0]/NET0131 ,
		_w5983_,
		_w5997_,
		_w5998_
	);
	LUT4 #(
		.INIT('hd070)
	) name5536 (
		\P1_state_reg[0]/NET0131 ,
		\P2_IR_reg[23]/NET0131 ,
		\P2_reg0_reg[4]/NET0131 ,
		_w1188_,
		_w5999_
	);
	LUT4 #(
		.INIT('h2000)
	) name5537 (
		\P2_reg0_reg[4]/NET0131 ,
		_w1189_,
		_w1352_,
		_w1356_,
		_w6000_
	);
	LUT4 #(
		.INIT('h08c8)
	) name5538 (
		\P2_reg0_reg[4]/NET0131 ,
		_w1191_,
		_w1369_,
		_w5533_,
		_w6001_
	);
	LUT4 #(
		.INIT('h0232)
	) name5539 (
		\P2_reg0_reg[4]/NET0131 ,
		_w1409_,
		_w1411_,
		_w5535_,
		_w6002_
	);
	LUT2 #(
		.INIT('h4)
	) name5540 (
		_w785_,
		_w1442_,
		_w6003_
	);
	LUT2 #(
		.INIT('h8)
	) name5541 (
		_w1411_,
		_w6003_,
		_w6004_
	);
	LUT3 #(
		.INIT('ha2)
	) name5542 (
		\P2_reg0_reg[4]/NET0131 ,
		_w1684_,
		_w1685_,
		_w6005_
	);
	LUT2 #(
		.INIT('h1)
	) name5543 (
		_w6004_,
		_w6005_,
		_w6006_
	);
	LUT4 #(
		.INIT('h0e02)
	) name5544 (
		\P2_reg0_reg[4]/NET0131 ,
		_w1411_,
		_w1496_,
		_w5540_,
		_w6007_
	);
	LUT4 #(
		.INIT('he020)
	) name5545 (
		\P2_reg0_reg[4]/NET0131 ,
		_w1369_,
		_w1447_,
		_w5540_,
		_w6008_
	);
	LUT4 #(
		.INIT('h0100)
	) name5546 (
		_w6002_,
		_w6007_,
		_w6008_,
		_w6006_,
		_w6009_
	);
	LUT4 #(
		.INIT('h1311)
	) name5547 (
		_w1359_,
		_w6000_,
		_w6001_,
		_w6009_,
		_w6010_
	);
	LUT3 #(
		.INIT('hce)
	) name5548 (
		\P1_state_reg[0]/NET0131 ,
		_w5999_,
		_w6010_,
		_w6011_
	);
	LUT4 #(
		.INIT('hd070)
	) name5549 (
		\P1_state_reg[0]/NET0131 ,
		\P2_IR_reg[23]/NET0131 ,
		\P2_reg1_reg[3]/NET0131 ,
		_w1188_,
		_w6012_
	);
	LUT4 #(
		.INIT('h2000)
	) name5550 (
		\P2_reg1_reg[3]/NET0131 ,
		_w1189_,
		_w1352_,
		_w1356_,
		_w6013_
	);
	LUT4 #(
		.INIT('h08c8)
	) name5551 (
		\P2_reg1_reg[3]/NET0131 ,
		_w1191_,
		_w1507_,
		_w5842_,
		_w6014_
	);
	LUT4 #(
		.INIT('h020e)
	) name5552 (
		\P2_reg1_reg[3]/NET0131 ,
		_w1516_,
		_w1575_,
		_w5845_,
		_w6015_
	);
	LUT2 #(
		.INIT('h8)
	) name5553 (
		_w1516_,
		_w5992_,
		_w6016_
	);
	LUT3 #(
		.INIT('ha2)
	) name5554 (
		\P2_reg1_reg[3]/NET0131 ,
		_w1684_,
		_w2469_,
		_w6017_
	);
	LUT2 #(
		.INIT('h1)
	) name5555 (
		_w6016_,
		_w6017_,
		_w6018_
	);
	LUT4 #(
		.INIT('h3202)
	) name5556 (
		\P2_reg1_reg[3]/NET0131 ,
		_w1506_,
		_w1516_,
		_w5844_,
		_w6019_
	);
	LUT4 #(
		.INIT('he020)
	) name5557 (
		\P2_reg1_reg[3]/NET0131 ,
		_w1507_,
		_w1530_,
		_w5844_,
		_w6020_
	);
	LUT4 #(
		.INIT('h0100)
	) name5558 (
		_w6015_,
		_w6019_,
		_w6020_,
		_w6018_,
		_w6021_
	);
	LUT4 #(
		.INIT('h1311)
	) name5559 (
		_w1359_,
		_w6013_,
		_w6014_,
		_w6021_,
		_w6022_
	);
	LUT3 #(
		.INIT('hce)
	) name5560 (
		\P1_state_reg[0]/NET0131 ,
		_w6012_,
		_w6022_,
		_w6023_
	);
	LUT4 #(
		.INIT('hd070)
	) name5561 (
		\P1_state_reg[0]/NET0131 ,
		\P2_IR_reg[23]/NET0131 ,
		\P2_reg1_reg[4]/NET0131 ,
		_w1188_,
		_w6024_
	);
	LUT4 #(
		.INIT('h2000)
	) name5562 (
		\P2_reg1_reg[4]/NET0131 ,
		_w1189_,
		_w1352_,
		_w1356_,
		_w6025_
	);
	LUT4 #(
		.INIT('h08c8)
	) name5563 (
		\P2_reg1_reg[4]/NET0131 ,
		_w1191_,
		_w1507_,
		_w5533_,
		_w6026_
	);
	LUT4 #(
		.INIT('h20e0)
	) name5564 (
		\P2_reg1_reg[4]/NET0131 ,
		_w1507_,
		_w1530_,
		_w5535_,
		_w6027_
	);
	LUT2 #(
		.INIT('h8)
	) name5565 (
		_w1516_,
		_w6003_,
		_w6028_
	);
	LUT3 #(
		.INIT('ha2)
	) name5566 (
		\P2_reg1_reg[4]/NET0131 ,
		_w1684_,
		_w2469_,
		_w6029_
	);
	LUT2 #(
		.INIT('h1)
	) name5567 (
		_w6028_,
		_w6029_,
		_w6030_
	);
	LUT4 #(
		.INIT('h0232)
	) name5568 (
		\P2_reg1_reg[4]/NET0131 ,
		_w1506_,
		_w1516_,
		_w5535_,
		_w6031_
	);
	LUT4 #(
		.INIT('h0e02)
	) name5569 (
		\P2_reg1_reg[4]/NET0131 ,
		_w1516_,
		_w1575_,
		_w5540_,
		_w6032_
	);
	LUT4 #(
		.INIT('h0100)
	) name5570 (
		_w6027_,
		_w6031_,
		_w6032_,
		_w6030_,
		_w6033_
	);
	LUT4 #(
		.INIT('h1311)
	) name5571 (
		_w1359_,
		_w6025_,
		_w6026_,
		_w6033_,
		_w6034_
	);
	LUT3 #(
		.INIT('hce)
	) name5572 (
		\P1_state_reg[0]/NET0131 ,
		_w6024_,
		_w6034_,
		_w6035_
	);
	LUT4 #(
		.INIT('hd070)
	) name5573 (
		\P1_state_reg[0]/NET0131 ,
		\P2_IR_reg[23]/NET0131 ,
		\P2_reg2_reg[3]/NET0131 ,
		_w1188_,
		_w6036_
	);
	LUT4 #(
		.INIT('h2000)
	) name5574 (
		\P2_reg2_reg[3]/NET0131 ,
		_w1189_,
		_w1352_,
		_w1356_,
		_w6037_
	);
	LUT4 #(
		.INIT('h08c8)
	) name5575 (
		\P2_reg2_reg[3]/NET0131 ,
		_w1191_,
		_w1516_,
		_w5842_,
		_w6038_
	);
	LUT4 #(
		.INIT('he020)
	) name5576 (
		\P2_reg2_reg[3]/NET0131 ,
		_w1516_,
		_w1530_,
		_w5844_,
		_w6039_
	);
	LUT3 #(
		.INIT('ha8)
	) name5577 (
		\P2_reg2_reg[3]/NET0131 ,
		_w1441_,
		_w1523_,
		_w6040_
	);
	LUT3 #(
		.INIT('h40)
	) name5578 (
		\P2_reg3_reg[3]/NET0131 ,
		_w1229_,
		_w1232_,
		_w6041_
	);
	LUT3 #(
		.INIT('h07)
	) name5579 (
		_w1507_,
		_w5992_,
		_w6041_,
		_w6042_
	);
	LUT2 #(
		.INIT('h4)
	) name5580 (
		_w6040_,
		_w6042_,
		_w6043_
	);
	LUT4 #(
		.INIT('h020e)
	) name5581 (
		\P2_reg2_reg[3]/NET0131 ,
		_w1507_,
		_w1575_,
		_w5845_,
		_w6044_
	);
	LUT4 #(
		.INIT('h3202)
	) name5582 (
		\P2_reg2_reg[3]/NET0131 ,
		_w1506_,
		_w1507_,
		_w5844_,
		_w6045_
	);
	LUT4 #(
		.INIT('h0100)
	) name5583 (
		_w6039_,
		_w6044_,
		_w6045_,
		_w6043_,
		_w6046_
	);
	LUT4 #(
		.INIT('h1311)
	) name5584 (
		_w1359_,
		_w6037_,
		_w6038_,
		_w6046_,
		_w6047_
	);
	LUT3 #(
		.INIT('hce)
	) name5585 (
		\P1_state_reg[0]/NET0131 ,
		_w6036_,
		_w6047_,
		_w6048_
	);
	LUT4 #(
		.INIT('hd070)
	) name5586 (
		\P1_state_reg[0]/NET0131 ,
		\P2_IR_reg[23]/NET0131 ,
		\P2_reg2_reg[4]/NET0131 ,
		_w1188_,
		_w6049_
	);
	LUT4 #(
		.INIT('h2000)
	) name5587 (
		\P2_reg2_reg[4]/NET0131 ,
		_w1189_,
		_w1352_,
		_w1356_,
		_w6050_
	);
	LUT4 #(
		.INIT('h08c8)
	) name5588 (
		\P2_reg2_reg[4]/NET0131 ,
		_w1191_,
		_w1516_,
		_w5533_,
		_w6051_
	);
	LUT4 #(
		.INIT('h0232)
	) name5589 (
		\P2_reg2_reg[4]/NET0131 ,
		_w1506_,
		_w1507_,
		_w5535_,
		_w6052_
	);
	LUT3 #(
		.INIT('ha8)
	) name5590 (
		\P2_reg2_reg[4]/NET0131 ,
		_w1441_,
		_w1523_,
		_w6053_
	);
	LUT3 #(
		.INIT('h40)
	) name5591 (
		_w776_,
		_w1229_,
		_w1232_,
		_w6054_
	);
	LUT3 #(
		.INIT('h07)
	) name5592 (
		_w1507_,
		_w6003_,
		_w6054_,
		_w6055_
	);
	LUT2 #(
		.INIT('h4)
	) name5593 (
		_w6053_,
		_w6055_,
		_w6056_
	);
	LUT4 #(
		.INIT('h20e0)
	) name5594 (
		\P2_reg2_reg[4]/NET0131 ,
		_w1516_,
		_w1530_,
		_w5535_,
		_w6057_
	);
	LUT4 #(
		.INIT('h0e02)
	) name5595 (
		\P2_reg2_reg[4]/NET0131 ,
		_w1507_,
		_w1575_,
		_w5540_,
		_w6058_
	);
	LUT4 #(
		.INIT('h0100)
	) name5596 (
		_w6052_,
		_w6057_,
		_w6058_,
		_w6056_,
		_w6059_
	);
	LUT4 #(
		.INIT('h1311)
	) name5597 (
		_w1359_,
		_w6050_,
		_w6051_,
		_w6059_,
		_w6060_
	);
	LUT3 #(
		.INIT('hce)
	) name5598 (
		\P1_state_reg[0]/NET0131 ,
		_w6049_,
		_w6060_,
		_w6061_
	);
	LUT2 #(
		.INIT('h2)
	) name5599 (
		\P1_reg0_reg[6]/NET0131 ,
		_w2462_,
		_w6062_
	);
	LUT4 #(
		.INIT('h2000)
	) name5600 (
		\P1_reg0_reg[6]/NET0131 ,
		_w1723_,
		_w1727_,
		_w1730_,
		_w6063_
	);
	LUT2 #(
		.INIT('h2)
	) name5601 (
		\P1_reg0_reg[6]/NET0131 ,
		_w2883_,
		_w6064_
	);
	LUT4 #(
		.INIT('hc808)
	) name5602 (
		\P1_reg0_reg[6]/NET0131 ,
		_w2424_,
		_w2883_,
		_w5496_,
		_w6065_
	);
	LUT4 #(
		.INIT('hc804)
	) name5603 (
		_w2797_,
		_w2883_,
		_w2932_,
		_w3182_,
		_w6066_
	);
	LUT3 #(
		.INIT('ha8)
	) name5604 (
		_w2388_,
		_w6064_,
		_w6066_,
		_w6067_
	);
	LUT4 #(
		.INIT('h10e0)
	) name5605 (
		_w2749_,
		_w2750_,
		_w2883_,
		_w3182_,
		_w6068_
	);
	LUT4 #(
		.INIT('hc808)
	) name5606 (
		\P1_reg0_reg[6]/NET0131 ,
		_w2447_,
		_w2883_,
		_w5501_,
		_w6069_
	);
	LUT2 #(
		.INIT('h8)
	) name5607 (
		_w2883_,
		_w5908_,
		_w6070_
	);
	LUT4 #(
		.INIT('h0a8a)
	) name5608 (
		\P1_reg0_reg[6]/NET0131 ,
		_w2426_,
		_w2524_,
		_w2883_,
		_w6071_
	);
	LUT2 #(
		.INIT('h1)
	) name5609 (
		_w6070_,
		_w6071_,
		_w6072_
	);
	LUT2 #(
		.INIT('h4)
	) name5610 (
		_w6069_,
		_w6072_,
		_w6073_
	);
	LUT4 #(
		.INIT('h5700)
	) name5611 (
		_w2292_,
		_w6064_,
		_w6068_,
		_w6073_,
		_w6074_
	);
	LUT4 #(
		.INIT('ha8aa)
	) name5612 (
		_w1731_,
		_w6067_,
		_w6065_,
		_w6074_,
		_w6075_
	);
	LUT4 #(
		.INIT('heeec)
	) name5613 (
		\P1_state_reg[0]/NET0131 ,
		_w6062_,
		_w6063_,
		_w6075_,
		_w6076_
	);
	LUT2 #(
		.INIT('h2)
	) name5614 (
		\P1_reg3_reg[1]/NET0131 ,
		_w2462_,
		_w6077_
	);
	LUT4 #(
		.INIT('h2000)
	) name5615 (
		\P1_reg3_reg[1]/NET0131 ,
		_w1723_,
		_w1727_,
		_w1730_,
		_w6078_
	);
	LUT4 #(
		.INIT('h20d0)
	) name5616 (
		_w2086_,
		_w2089_,
		_w2388_,
		_w3189_,
		_w6079_
	);
	LUT3 #(
		.INIT('h60)
	) name5617 (
		_w2081_,
		_w2089_,
		_w2447_,
		_w6080_
	);
	LUT4 #(
		.INIT('h007b)
	) name5618 (
		_w2090_,
		_w2292_,
		_w3189_,
		_w6080_,
		_w6081_
	);
	LUT3 #(
		.INIT('h8a)
	) name5619 (
		_w2644_,
		_w6079_,
		_w6081_,
		_w6082_
	);
	LUT4 #(
		.INIT('h4144)
	) name5620 (
		_w1747_,
		_w2061_,
		_w2077_,
		_w2399_,
		_w6083_
	);
	LUT3 #(
		.INIT('h80)
	) name5621 (
		_w1747_,
		_w2084_,
		_w2085_,
		_w6084_
	);
	LUT4 #(
		.INIT('hddd1)
	) name5622 (
		\P1_reg3_reg[1]/NET0131 ,
		_w2644_,
		_w6083_,
		_w6084_,
		_w6085_
	);
	LUT4 #(
		.INIT('h30a0)
	) name5623 (
		\P1_reg3_reg[1]/NET0131 ,
		_w2081_,
		_w2426_,
		_w2644_,
		_w6086_
	);
	LUT2 #(
		.INIT('h4)
	) name5624 (
		_w2081_,
		_w2454_,
		_w6087_
	);
	LUT3 #(
		.INIT('h23)
	) name5625 (
		_w2282_,
		_w2285_,
		_w2449_,
		_w6088_
	);
	LUT4 #(
		.INIT('h888a)
	) name5626 (
		\P1_reg3_reg[1]/NET0131 ,
		_w2450_,
		_w2644_,
		_w6088_,
		_w6089_
	);
	LUT3 #(
		.INIT('h01)
	) name5627 (
		_w6087_,
		_w6089_,
		_w6086_,
		_w6090_
	);
	LUT4 #(
		.INIT('h0d00)
	) name5628 (
		_w2424_,
		_w6085_,
		_w6082_,
		_w6090_,
		_w6091_
	);
	LUT4 #(
		.INIT('ha0a8)
	) name5629 (
		\P1_state_reg[0]/NET0131 ,
		_w1731_,
		_w6078_,
		_w6091_,
		_w6092_
	);
	LUT2 #(
		.INIT('he)
	) name5630 (
		_w6077_,
		_w6092_,
		_w6093_
	);
	LUT4 #(
		.INIT('hd070)
	) name5631 (
		\P1_state_reg[0]/NET0131 ,
		\P2_IR_reg[23]/NET0131 ,
		\P2_reg3_reg[1]/NET0131 ,
		_w1188_,
		_w6094_
	);
	LUT4 #(
		.INIT('h2000)
	) name5632 (
		\P2_reg3_reg[1]/NET0131 ,
		_w1189_,
		_w1352_,
		_w1356_,
		_w6095_
	);
	LUT2 #(
		.INIT('h1)
	) name5633 (
		_w823_,
		_w1435_,
		_w6096_
	);
	LUT4 #(
		.INIT('h006f)
	) name5634 (
		_w803_,
		_w1414_,
		_w1435_,
		_w6096_,
		_w6097_
	);
	LUT4 #(
		.INIT('h08c8)
	) name5635 (
		\P2_reg3_reg[1]/NET0131 ,
		_w1191_,
		_w1411_,
		_w6097_,
		_w6098_
	);
	LUT4 #(
		.INIT('h02aa)
	) name5636 (
		\P2_reg3_reg[1]/NET0131 ,
		_w1361_,
		_w1363_,
		_w1368_,
		_w6099_
	);
	LUT4 #(
		.INIT('h9969)
	) name5637 (
		_w814_,
		_w818_,
		_w823_,
		_w826_,
		_w6100_
	);
	LUT4 #(
		.INIT('h020e)
	) name5638 (
		\P2_reg3_reg[1]/NET0131 ,
		_w1369_,
		_w1409_,
		_w6100_,
		_w6101_
	);
	LUT4 #(
		.INIT('h5400)
	) name5639 (
		_w818_,
		_w1361_,
		_w1363_,
		_w1368_,
		_w6102_
	);
	LUT3 #(
		.INIT('h20)
	) name5640 (
		\P2_reg3_reg[1]/NET0131 ,
		_w1184_,
		_w1190_,
		_w6103_
	);
	LUT3 #(
		.INIT('h0b)
	) name5641 (
		_w818_,
		_w1233_,
		_w6103_,
		_w6104_
	);
	LUT4 #(
		.INIT('h5700)
	) name5642 (
		_w1442_,
		_w6099_,
		_w6102_,
		_w6104_,
		_w6105_
	);
	LUT4 #(
		.INIT('h6669)
	) name5643 (
		_w814_,
		_w818_,
		_w823_,
		_w826_,
		_w6106_
	);
	LUT4 #(
		.INIT('h0e02)
	) name5644 (
		\P2_reg3_reg[1]/NET0131 ,
		_w1369_,
		_w1496_,
		_w6106_,
		_w6107_
	);
	LUT4 #(
		.INIT('hc808)
	) name5645 (
		\P2_reg3_reg[1]/NET0131 ,
		_w1447_,
		_w1411_,
		_w6106_,
		_w6108_
	);
	LUT4 #(
		.INIT('h0100)
	) name5646 (
		_w6101_,
		_w6107_,
		_w6108_,
		_w6105_,
		_w6109_
	);
	LUT4 #(
		.INIT('h1311)
	) name5647 (
		_w1359_,
		_w6095_,
		_w6098_,
		_w6109_,
		_w6110_
	);
	LUT3 #(
		.INIT('hce)
	) name5648 (
		\P1_state_reg[0]/NET0131 ,
		_w6094_,
		_w6110_,
		_w6111_
	);
	LUT2 #(
		.INIT('h2)
	) name5649 (
		\P1_reg3_reg[2]/NET0131 ,
		_w2462_,
		_w6112_
	);
	LUT4 #(
		.INIT('h2000)
	) name5650 (
		\P1_reg3_reg[2]/NET0131 ,
		_w1723_,
		_w1727_,
		_w1730_,
		_w6113_
	);
	LUT2 #(
		.INIT('h2)
	) name5651 (
		\P1_reg3_reg[2]/NET0131 ,
		_w2644_,
		_w6114_
	);
	LUT4 #(
		.INIT('h5655)
	) name5652 (
		_w492_,
		_w2061_,
		_w2077_,
		_w2399_,
		_w6115_
	);
	LUT4 #(
		.INIT('h7020)
	) name5653 (
		_w1747_,
		_w2077_,
		_w2644_,
		_w6115_,
		_w6116_
	);
	LUT3 #(
		.INIT('ha8)
	) name5654 (
		_w2424_,
		_w6114_,
		_w6116_,
		_w6117_
	);
	LUT4 #(
		.INIT('hb24d)
	) name5655 (
		_w2077_,
		_w2081_,
		_w2305_,
		_w3184_,
		_w6118_
	);
	LUT4 #(
		.INIT('hc808)
	) name5656 (
		\P1_reg3_reg[2]/NET0131 ,
		_w2388_,
		_w2644_,
		_w6118_,
		_w6119_
	);
	LUT4 #(
		.INIT('h45ba)
	) name5657 (
		_w2082_,
		_w2083_,
		_w2090_,
		_w3184_,
		_w6120_
	);
	LUT4 #(
		.INIT('h08c8)
	) name5658 (
		\P1_reg3_reg[2]/NET0131 ,
		_w2292_,
		_w2644_,
		_w6120_,
		_w6121_
	);
	LUT3 #(
		.INIT('h6a)
	) name5659 (
		_w2065_,
		_w2081_,
		_w2089_,
		_w6122_
	);
	LUT4 #(
		.INIT('hc808)
	) name5660 (
		\P1_reg3_reg[2]/NET0131 ,
		_w2447_,
		_w2644_,
		_w6122_,
		_w6123_
	);
	LUT4 #(
		.INIT('h5450)
	) name5661 (
		_w2065_,
		_w2426_,
		_w2454_,
		_w2644_,
		_w6124_
	);
	LUT4 #(
		.INIT('ha0a8)
	) name5662 (
		\P1_reg3_reg[2]/NET0131 ,
		_w2426_,
		_w2450_,
		_w2644_,
		_w6125_
	);
	LUT3 #(
		.INIT('h01)
	) name5663 (
		_w6124_,
		_w6123_,
		_w6125_,
		_w6126_
	);
	LUT3 #(
		.INIT('h10)
	) name5664 (
		_w6121_,
		_w6119_,
		_w6126_,
		_w6127_
	);
	LUT4 #(
		.INIT('h1311)
	) name5665 (
		_w1731_,
		_w6113_,
		_w6117_,
		_w6127_,
		_w6128_
	);
	LUT3 #(
		.INIT('hce)
	) name5666 (
		\P1_state_reg[0]/NET0131 ,
		_w6112_,
		_w6128_,
		_w6129_
	);
	LUT4 #(
		.INIT('hd070)
	) name5667 (
		\P1_state_reg[0]/NET0131 ,
		\P2_IR_reg[23]/NET0131 ,
		\P2_reg0_reg[2]/NET0131 ,
		_w1188_,
		_w6130_
	);
	LUT4 #(
		.INIT('h2000)
	) name5668 (
		\P2_reg0_reg[2]/NET0131 ,
		_w1189_,
		_w1352_,
		_w1356_,
		_w6131_
	);
	LUT4 #(
		.INIT('h111d)
	) name5669 (
		\P2_reg0_reg[2]/NET0131 ,
		_w1369_,
		_w5955_,
		_w5956_,
		_w6132_
	);
	LUT4 #(
		.INIT('hc535)
	) name5670 (
		\P2_reg0_reg[2]/NET0131 ,
		_w1321_,
		_w1411_,
		_w1452_,
		_w6133_
	);
	LUT2 #(
		.INIT('h4)
	) name5671 (
		_w807_,
		_w1442_,
		_w6134_
	);
	LUT2 #(
		.INIT('h8)
	) name5672 (
		_w1411_,
		_w6134_,
		_w6135_
	);
	LUT3 #(
		.INIT('ha2)
	) name5673 (
		\P2_reg0_reg[2]/NET0131 ,
		_w1684_,
		_w1685_,
		_w6136_
	);
	LUT4 #(
		.INIT('h0032)
	) name5674 (
		_w1496_,
		_w6135_,
		_w6133_,
		_w6136_,
		_w6137_
	);
	LUT4 #(
		.INIT('hc535)
	) name5675 (
		\P2_reg0_reg[2]/NET0131 ,
		_w1321_,
		_w1369_,
		_w1452_,
		_w6138_
	);
	LUT4 #(
		.INIT('hc355)
	) name5676 (
		\P2_reg0_reg[2]/NET0131 ,
		_w1210_,
		_w1321_,
		_w1411_,
		_w6139_
	);
	LUT4 #(
		.INIT('hf3a2)
	) name5677 (
		_w1409_,
		_w1447_,
		_w6138_,
		_w6139_,
		_w6140_
	);
	LUT4 #(
		.INIT('hd000)
	) name5678 (
		_w1191_,
		_w6132_,
		_w6137_,
		_w6140_,
		_w6141_
	);
	LUT4 #(
		.INIT('ha0a8)
	) name5679 (
		\P1_state_reg[0]/NET0131 ,
		_w1359_,
		_w6131_,
		_w6141_,
		_w6142_
	);
	LUT2 #(
		.INIT('he)
	) name5680 (
		_w6130_,
		_w6142_,
		_w6143_
	);
	LUT4 #(
		.INIT('hd070)
	) name5681 (
		\P1_state_reg[0]/NET0131 ,
		\P2_IR_reg[23]/NET0131 ,
		\P2_reg1_reg[2]/NET0131 ,
		_w1188_,
		_w6144_
	);
	LUT4 #(
		.INIT('h2000)
	) name5682 (
		\P2_reg1_reg[2]/NET0131 ,
		_w1189_,
		_w1352_,
		_w1356_,
		_w6145_
	);
	LUT4 #(
		.INIT('h111d)
	) name5683 (
		\P2_reg1_reg[2]/NET0131 ,
		_w1507_,
		_w5955_,
		_w5956_,
		_w6146_
	);
	LUT3 #(
		.INIT('h06)
	) name5684 (
		_w1210_,
		_w1321_,
		_w1506_,
		_w6147_
	);
	LUT4 #(
		.INIT('h00f9)
	) name5685 (
		_w1321_,
		_w1452_,
		_w1575_,
		_w6134_,
		_w6148_
	);
	LUT3 #(
		.INIT('h8a)
	) name5686 (
		_w1516_,
		_w6147_,
		_w6148_,
		_w6149_
	);
	LUT4 #(
		.INIT('hc355)
	) name5687 (
		\P2_reg1_reg[2]/NET0131 ,
		_w1210_,
		_w1321_,
		_w1507_,
		_w6150_
	);
	LUT4 #(
		.INIT('hf20f)
	) name5688 (
		_w1179_,
		_w1183_,
		_w1186_,
		_w1189_,
		_w6151_
	);
	LUT4 #(
		.INIT('h00f1)
	) name5689 (
		_w1361_,
		_w1363_,
		_w1368_,
		_w6151_,
		_w6152_
	);
	LUT3 #(
		.INIT('h02)
	) name5690 (
		_w1684_,
		_w2469_,
		_w6152_,
		_w6153_
	);
	LUT4 #(
		.INIT('haaa2)
	) name5691 (
		\P2_reg1_reg[2]/NET0131 ,
		_w1684_,
		_w2469_,
		_w6152_,
		_w6154_
	);
	LUT3 #(
		.INIT('h0d)
	) name5692 (
		_w1530_,
		_w6150_,
		_w6154_,
		_w6155_
	);
	LUT4 #(
		.INIT('h3100)
	) name5693 (
		_w1191_,
		_w6149_,
		_w6146_,
		_w6155_,
		_w6156_
	);
	LUT4 #(
		.INIT('ha0a8)
	) name5694 (
		\P1_state_reg[0]/NET0131 ,
		_w1359_,
		_w6145_,
		_w6156_,
		_w6157_
	);
	LUT2 #(
		.INIT('he)
	) name5695 (
		_w6144_,
		_w6157_,
		_w6158_
	);
	LUT4 #(
		.INIT('hd070)
	) name5696 (
		\P1_state_reg[0]/NET0131 ,
		\P2_IR_reg[23]/NET0131 ,
		\P2_reg2_reg[2]/NET0131 ,
		_w1188_,
		_w6159_
	);
	LUT4 #(
		.INIT('h2000)
	) name5697 (
		\P2_reg2_reg[2]/NET0131 ,
		_w1189_,
		_w1352_,
		_w1356_,
		_w6160_
	);
	LUT4 #(
		.INIT('h111d)
	) name5698 (
		\P2_reg2_reg[2]/NET0131 ,
		_w1516_,
		_w5955_,
		_w5956_,
		_w6161_
	);
	LUT4 #(
		.INIT('hc355)
	) name5699 (
		\P2_reg2_reg[2]/NET0131 ,
		_w1210_,
		_w1321_,
		_w1507_,
		_w6162_
	);
	LUT3 #(
		.INIT('ha8)
	) name5700 (
		\P2_reg2_reg[2]/NET0131 ,
		_w1441_,
		_w1523_,
		_w6163_
	);
	LUT3 #(
		.INIT('h80)
	) name5701 (
		\P2_reg3_reg[2]/NET0131 ,
		_w1229_,
		_w1232_,
		_w6164_
	);
	LUT3 #(
		.INIT('h07)
	) name5702 (
		_w1507_,
		_w6134_,
		_w6164_,
		_w6165_
	);
	LUT4 #(
		.INIT('h0e00)
	) name5703 (
		_w1506_,
		_w6162_,
		_w6163_,
		_w6165_,
		_w6166_
	);
	LUT4 #(
		.INIT('hc355)
	) name5704 (
		\P2_reg2_reg[2]/NET0131 ,
		_w1321_,
		_w1452_,
		_w1507_,
		_w6167_
	);
	LUT4 #(
		.INIT('hc355)
	) name5705 (
		\P2_reg2_reg[2]/NET0131 ,
		_w1210_,
		_w1321_,
		_w1516_,
		_w6168_
	);
	LUT4 #(
		.INIT('hfc54)
	) name5706 (
		_w1530_,
		_w1575_,
		_w6167_,
		_w6168_,
		_w6169_
	);
	LUT4 #(
		.INIT('hd000)
	) name5707 (
		_w1191_,
		_w6161_,
		_w6166_,
		_w6169_,
		_w6170_
	);
	LUT4 #(
		.INIT('ha0a8)
	) name5708 (
		\P1_state_reg[0]/NET0131 ,
		_w1359_,
		_w6160_,
		_w6170_,
		_w6171_
	);
	LUT2 #(
		.INIT('he)
	) name5709 (
		_w6159_,
		_w6171_,
		_w6172_
	);
	LUT2 #(
		.INIT('h2)
	) name5710 (
		\P1_reg0_reg[2]/NET0131 ,
		_w2462_,
		_w6173_
	);
	LUT4 #(
		.INIT('h2000)
	) name5711 (
		\P1_reg0_reg[2]/NET0131 ,
		_w1723_,
		_w1727_,
		_w1730_,
		_w6174_
	);
	LUT2 #(
		.INIT('h2)
	) name5712 (
		\P1_reg0_reg[2]/NET0131 ,
		_w2883_,
		_w6175_
	);
	LUT4 #(
		.INIT('h7020)
	) name5713 (
		_w1747_,
		_w2077_,
		_w2883_,
		_w6115_,
		_w6176_
	);
	LUT3 #(
		.INIT('ha8)
	) name5714 (
		_w2424_,
		_w6175_,
		_w6176_,
		_w6177_
	);
	LUT4 #(
		.INIT('h08c8)
	) name5715 (
		\P1_reg0_reg[2]/NET0131 ,
		_w2292_,
		_w2883_,
		_w6120_,
		_w6178_
	);
	LUT4 #(
		.INIT('hc808)
	) name5716 (
		\P1_reg0_reg[2]/NET0131 ,
		_w2388_,
		_w2883_,
		_w6118_,
		_w6179_
	);
	LUT4 #(
		.INIT('hc808)
	) name5717 (
		\P1_reg0_reg[2]/NET0131 ,
		_w2447_,
		_w2883_,
		_w6122_,
		_w6180_
	);
	LUT2 #(
		.INIT('h4)
	) name5718 (
		_w2065_,
		_w2426_,
		_w6181_
	);
	LUT2 #(
		.INIT('h8)
	) name5719 (
		_w2883_,
		_w6181_,
		_w6182_
	);
	LUT4 #(
		.INIT('h0a8a)
	) name5720 (
		\P1_reg0_reg[2]/NET0131 ,
		_w2426_,
		_w2524_,
		_w2883_,
		_w6183_
	);
	LUT3 #(
		.INIT('h01)
	) name5721 (
		_w6182_,
		_w6180_,
		_w6183_,
		_w6184_
	);
	LUT3 #(
		.INIT('h10)
	) name5722 (
		_w6179_,
		_w6178_,
		_w6184_,
		_w6185_
	);
	LUT4 #(
		.INIT('h1311)
	) name5723 (
		_w1731_,
		_w6174_,
		_w6177_,
		_w6185_,
		_w6186_
	);
	LUT3 #(
		.INIT('hce)
	) name5724 (
		\P1_state_reg[0]/NET0131 ,
		_w6173_,
		_w6186_,
		_w6187_
	);
	LUT2 #(
		.INIT('h2)
	) name5725 (
		\P1_reg1_reg[2]/NET0131 ,
		_w2462_,
		_w6188_
	);
	LUT4 #(
		.INIT('h2000)
	) name5726 (
		\P1_reg1_reg[2]/NET0131 ,
		_w1723_,
		_w1727_,
		_w1730_,
		_w6189_
	);
	LUT2 #(
		.INIT('h2)
	) name5727 (
		\P1_reg1_reg[2]/NET0131 ,
		_w2520_,
		_w6190_
	);
	LUT4 #(
		.INIT('h7020)
	) name5728 (
		_w1747_,
		_w2077_,
		_w2520_,
		_w6115_,
		_w6191_
	);
	LUT3 #(
		.INIT('ha8)
	) name5729 (
		_w2424_,
		_w6190_,
		_w6191_,
		_w6192_
	);
	LUT4 #(
		.INIT('h08c8)
	) name5730 (
		\P1_reg1_reg[2]/NET0131 ,
		_w2292_,
		_w2520_,
		_w6120_,
		_w6193_
	);
	LUT4 #(
		.INIT('hc808)
	) name5731 (
		\P1_reg1_reg[2]/NET0131 ,
		_w2388_,
		_w2520_,
		_w6118_,
		_w6194_
	);
	LUT4 #(
		.INIT('hc808)
	) name5732 (
		\P1_reg1_reg[2]/NET0131 ,
		_w2447_,
		_w2520_,
		_w6122_,
		_w6195_
	);
	LUT2 #(
		.INIT('h8)
	) name5733 (
		_w2520_,
		_w6181_,
		_w6196_
	);
	LUT4 #(
		.INIT('h08aa)
	) name5734 (
		\P1_reg1_reg[2]/NET0131 ,
		_w2426_,
		_w2520_,
		_w2524_,
		_w6197_
	);
	LUT3 #(
		.INIT('h01)
	) name5735 (
		_w6196_,
		_w6195_,
		_w6197_,
		_w6198_
	);
	LUT3 #(
		.INIT('h10)
	) name5736 (
		_w6194_,
		_w6193_,
		_w6198_,
		_w6199_
	);
	LUT4 #(
		.INIT('h1311)
	) name5737 (
		_w1731_,
		_w6189_,
		_w6192_,
		_w6199_,
		_w6200_
	);
	LUT3 #(
		.INIT('hce)
	) name5738 (
		\P1_state_reg[0]/NET0131 ,
		_w6188_,
		_w6200_,
		_w6201_
	);
	LUT4 #(
		.INIT('hd070)
	) name5739 (
		\P1_state_reg[0]/NET0131 ,
		\P2_IR_reg[23]/NET0131 ,
		\P2_reg0_reg[1]/NET0131 ,
		_w1188_,
		_w6202_
	);
	LUT4 #(
		.INIT('h2000)
	) name5740 (
		\P2_reg0_reg[1]/NET0131 ,
		_w1189_,
		_w1352_,
		_w1356_,
		_w6203_
	);
	LUT4 #(
		.INIT('h08c8)
	) name5741 (
		\P2_reg0_reg[1]/NET0131 ,
		_w1191_,
		_w1369_,
		_w6097_,
		_w6204_
	);
	LUT4 #(
		.INIT('he020)
	) name5742 (
		\P2_reg0_reg[1]/NET0131 ,
		_w1369_,
		_w1447_,
		_w6106_,
		_w6205_
	);
	LUT2 #(
		.INIT('h2)
	) name5743 (
		\P2_reg0_reg[1]/NET0131 ,
		_w1684_,
		_w6206_
	);
	LUT4 #(
		.INIT('haaa8)
	) name5744 (
		\P2_reg0_reg[1]/NET0131 ,
		_w1361_,
		_w1363_,
		_w1368_,
		_w6207_
	);
	LUT4 #(
		.INIT('h0001)
	) name5745 (
		_w818_,
		_w1361_,
		_w1363_,
		_w1368_,
		_w6208_
	);
	LUT4 #(
		.INIT('h1113)
	) name5746 (
		_w1442_,
		_w6206_,
		_w6207_,
		_w6208_,
		_w6209_
	);
	LUT4 #(
		.INIT('h0e02)
	) name5747 (
		\P2_reg0_reg[1]/NET0131 ,
		_w1411_,
		_w1496_,
		_w6106_,
		_w6210_
	);
	LUT4 #(
		.INIT('h0232)
	) name5748 (
		\P2_reg0_reg[1]/NET0131 ,
		_w1409_,
		_w1411_,
		_w6100_,
		_w6211_
	);
	LUT4 #(
		.INIT('h0100)
	) name5749 (
		_w6205_,
		_w6210_,
		_w6211_,
		_w6209_,
		_w6212_
	);
	LUT4 #(
		.INIT('h1311)
	) name5750 (
		_w1359_,
		_w6203_,
		_w6204_,
		_w6212_,
		_w6213_
	);
	LUT3 #(
		.INIT('hce)
	) name5751 (
		\P1_state_reg[0]/NET0131 ,
		_w6202_,
		_w6213_,
		_w6214_
	);
	LUT4 #(
		.INIT('hd070)
	) name5752 (
		\P1_state_reg[0]/NET0131 ,
		\P2_IR_reg[23]/NET0131 ,
		\P2_reg1_reg[1]/NET0131 ,
		_w1188_,
		_w6215_
	);
	LUT4 #(
		.INIT('h2000)
	) name5753 (
		\P2_reg1_reg[1]/NET0131 ,
		_w1189_,
		_w1352_,
		_w1356_,
		_w6216_
	);
	LUT4 #(
		.INIT('h08c8)
	) name5754 (
		\P2_reg1_reg[1]/NET0131 ,
		_w1191_,
		_w1507_,
		_w6097_,
		_w6217_
	);
	LUT4 #(
		.INIT('h20e0)
	) name5755 (
		\P2_reg1_reg[1]/NET0131 ,
		_w1507_,
		_w1530_,
		_w6100_,
		_w6218_
	);
	LUT2 #(
		.INIT('h2)
	) name5756 (
		\P2_reg1_reg[1]/NET0131 ,
		_w1684_,
		_w6219_
	);
	LUT4 #(
		.INIT('haa02)
	) name5757 (
		\P2_reg1_reg[1]/NET0131 ,
		_w1361_,
		_w1363_,
		_w1368_,
		_w6220_
	);
	LUT4 #(
		.INIT('h0054)
	) name5758 (
		_w818_,
		_w1361_,
		_w1363_,
		_w1368_,
		_w6221_
	);
	LUT4 #(
		.INIT('h1113)
	) name5759 (
		_w1442_,
		_w6219_,
		_w6220_,
		_w6221_,
		_w6222_
	);
	LUT4 #(
		.INIT('h0232)
	) name5760 (
		\P2_reg1_reg[1]/NET0131 ,
		_w1506_,
		_w1516_,
		_w6100_,
		_w6223_
	);
	LUT4 #(
		.INIT('h0e02)
	) name5761 (
		\P2_reg1_reg[1]/NET0131 ,
		_w1516_,
		_w1575_,
		_w6106_,
		_w6224_
	);
	LUT4 #(
		.INIT('h0100)
	) name5762 (
		_w6218_,
		_w6223_,
		_w6224_,
		_w6222_,
		_w6225_
	);
	LUT4 #(
		.INIT('h1311)
	) name5763 (
		_w1359_,
		_w6216_,
		_w6217_,
		_w6225_,
		_w6226_
	);
	LUT3 #(
		.INIT('hce)
	) name5764 (
		\P1_state_reg[0]/NET0131 ,
		_w6215_,
		_w6226_,
		_w6227_
	);
	LUT2 #(
		.INIT('h2)
	) name5765 (
		\P1_reg2_reg[2]/NET0131 ,
		_w2462_,
		_w6228_
	);
	LUT4 #(
		.INIT('h2000)
	) name5766 (
		\P1_reg2_reg[2]/NET0131 ,
		_w1723_,
		_w1727_,
		_w1730_,
		_w6229_
	);
	LUT2 #(
		.INIT('h2)
	) name5767 (
		\P1_reg2_reg[2]/NET0131 ,
		_w1741_,
		_w6230_
	);
	LUT4 #(
		.INIT('h2a08)
	) name5768 (
		_w1741_,
		_w1747_,
		_w2077_,
		_w6115_,
		_w6231_
	);
	LUT3 #(
		.INIT('ha8)
	) name5769 (
		_w2424_,
		_w6230_,
		_w6231_,
		_w6232_
	);
	LUT2 #(
		.INIT('h2)
	) name5770 (
		_w2292_,
		_w6120_,
		_w6233_
	);
	LUT4 #(
		.INIT('h6a00)
	) name5771 (
		_w2065_,
		_w2081_,
		_w2089_,
		_w2447_,
		_w6234_
	);
	LUT3 #(
		.INIT('h07)
	) name5772 (
		_w2388_,
		_w6118_,
		_w6234_,
		_w6235_
	);
	LUT4 #(
		.INIT('h00ab)
	) name5773 (
		_w1741_,
		_w2285_,
		_w2447_,
		_w2450_,
		_w6236_
	);
	LUT4 #(
		.INIT('h0008)
	) name5774 (
		\P1_reg3_reg[2]/NET0131 ,
		_w2284_,
		_w2288_,
		_w2291_,
		_w6237_
	);
	LUT4 #(
		.INIT('h2e00)
	) name5775 (
		\P1_reg2_reg[2]/NET0131 ,
		_w1741_,
		_w2065_,
		_w2426_,
		_w6238_
	);
	LUT4 #(
		.INIT('h0301)
	) name5776 (
		\P1_reg2_reg[2]/NET0131 ,
		_w6237_,
		_w6238_,
		_w6236_,
		_w6239_
	);
	LUT4 #(
		.INIT('h7500)
	) name5777 (
		_w1741_,
		_w6233_,
		_w6235_,
		_w6239_,
		_w6240_
	);
	LUT4 #(
		.INIT('h1311)
	) name5778 (
		_w1731_,
		_w6229_,
		_w6232_,
		_w6240_,
		_w6241_
	);
	LUT3 #(
		.INIT('hce)
	) name5779 (
		\P1_state_reg[0]/NET0131 ,
		_w6228_,
		_w6241_,
		_w6242_
	);
	LUT4 #(
		.INIT('hd070)
	) name5780 (
		\P1_state_reg[0]/NET0131 ,
		\P2_IR_reg[23]/NET0131 ,
		\P2_reg2_reg[1]/NET0131 ,
		_w1188_,
		_w6243_
	);
	LUT4 #(
		.INIT('h2000)
	) name5781 (
		\P2_reg2_reg[1]/NET0131 ,
		_w1189_,
		_w1352_,
		_w1356_,
		_w6244_
	);
	LUT4 #(
		.INIT('h08c8)
	) name5782 (
		\P2_reg2_reg[1]/NET0131 ,
		_w1191_,
		_w1516_,
		_w6097_,
		_w6245_
	);
	LUT4 #(
		.INIT('h20e0)
	) name5783 (
		\P2_reg2_reg[1]/NET0131 ,
		_w1516_,
		_w1530_,
		_w6100_,
		_w6246_
	);
	LUT4 #(
		.INIT('ha8aa)
	) name5784 (
		\P2_reg2_reg[1]/NET0131 ,
		_w1361_,
		_w1363_,
		_w1368_,
		_w6247_
	);
	LUT4 #(
		.INIT('h0100)
	) name5785 (
		_w818_,
		_w1361_,
		_w1363_,
		_w1368_,
		_w6248_
	);
	LUT3 #(
		.INIT('h80)
	) name5786 (
		\P2_reg3_reg[1]/NET0131 ,
		_w1229_,
		_w1232_,
		_w6249_
	);
	LUT3 #(
		.INIT('h20)
	) name5787 (
		\P2_reg2_reg[1]/NET0131 ,
		_w1184_,
		_w1190_,
		_w6250_
	);
	LUT2 #(
		.INIT('h1)
	) name5788 (
		_w6249_,
		_w6250_,
		_w6251_
	);
	LUT4 #(
		.INIT('h5700)
	) name5789 (
		_w1442_,
		_w6247_,
		_w6248_,
		_w6251_,
		_w6252_
	);
	LUT4 #(
		.INIT('h0232)
	) name5790 (
		\P2_reg2_reg[1]/NET0131 ,
		_w1506_,
		_w1507_,
		_w6100_,
		_w6253_
	);
	LUT4 #(
		.INIT('h0e02)
	) name5791 (
		\P2_reg2_reg[1]/NET0131 ,
		_w1507_,
		_w1575_,
		_w6106_,
		_w6254_
	);
	LUT4 #(
		.INIT('h0100)
	) name5792 (
		_w6246_,
		_w6253_,
		_w6254_,
		_w6252_,
		_w6255_
	);
	LUT4 #(
		.INIT('h1311)
	) name5793 (
		_w1359_,
		_w6244_,
		_w6245_,
		_w6255_,
		_w6256_
	);
	LUT3 #(
		.INIT('hce)
	) name5794 (
		\P1_state_reg[0]/NET0131 ,
		_w6243_,
		_w6256_,
		_w6257_
	);
	LUT2 #(
		.INIT('h2)
	) name5795 (
		\P1_reg0_reg[1]/NET0131 ,
		_w2462_,
		_w6258_
	);
	LUT4 #(
		.INIT('h2000)
	) name5796 (
		\P1_reg0_reg[1]/NET0131 ,
		_w1723_,
		_w1727_,
		_w1730_,
		_w6259_
	);
	LUT3 #(
		.INIT('h8a)
	) name5797 (
		_w2883_,
		_w6079_,
		_w6081_,
		_w6260_
	);
	LUT4 #(
		.INIT('hddd1)
	) name5798 (
		\P1_reg0_reg[1]/NET0131 ,
		_w2883_,
		_w6083_,
		_w6084_,
		_w6261_
	);
	LUT4 #(
		.INIT('h30a0)
	) name5799 (
		\P1_reg0_reg[1]/NET0131 ,
		_w2081_,
		_w2426_,
		_w2883_,
		_w6262_
	);
	LUT4 #(
		.INIT('h222a)
	) name5800 (
		\P1_reg0_reg[1]/NET0131 ,
		_w2524_,
		_w2883_,
		_w6088_,
		_w6263_
	);
	LUT2 #(
		.INIT('h1)
	) name5801 (
		_w6262_,
		_w6263_,
		_w6264_
	);
	LUT4 #(
		.INIT('h0d00)
	) name5802 (
		_w2424_,
		_w6261_,
		_w6260_,
		_w6264_,
		_w6265_
	);
	LUT4 #(
		.INIT('ha0a8)
	) name5803 (
		\P1_state_reg[0]/NET0131 ,
		_w1731_,
		_w6259_,
		_w6265_,
		_w6266_
	);
	LUT2 #(
		.INIT('he)
	) name5804 (
		_w6258_,
		_w6266_,
		_w6267_
	);
	LUT2 #(
		.INIT('h2)
	) name5805 (
		\P1_reg1_reg[1]/NET0131 ,
		_w2462_,
		_w6268_
	);
	LUT4 #(
		.INIT('h2000)
	) name5806 (
		\P1_reg1_reg[1]/NET0131 ,
		_w1723_,
		_w1727_,
		_w1730_,
		_w6269_
	);
	LUT2 #(
		.INIT('h2)
	) name5807 (
		\P1_reg1_reg[1]/NET0131 ,
		_w2520_,
		_w6270_
	);
	LUT4 #(
		.INIT('hddd1)
	) name5808 (
		\P1_reg1_reg[1]/NET0131 ,
		_w2520_,
		_w6083_,
		_w6084_,
		_w6271_
	);
	LUT2 #(
		.INIT('h2)
	) name5809 (
		_w2424_,
		_w6271_,
		_w6272_
	);
	LUT4 #(
		.INIT('h20d0)
	) name5810 (
		_w2086_,
		_w2089_,
		_w2520_,
		_w3189_,
		_w6273_
	);
	LUT3 #(
		.INIT('ha8)
	) name5811 (
		_w2388_,
		_w6270_,
		_w6273_,
		_w6274_
	);
	LUT4 #(
		.INIT('h35c5)
	) name5812 (
		\P1_reg1_reg[1]/NET0131 ,
		_w2090_,
		_w2520_,
		_w3189_,
		_w6275_
	);
	LUT2 #(
		.INIT('h2)
	) name5813 (
		_w2292_,
		_w6275_,
		_w6276_
	);
	LUT4 #(
		.INIT('h89af)
	) name5814 (
		_w2081_,
		_w2089_,
		_w2426_,
		_w2447_,
		_w6277_
	);
	LUT2 #(
		.INIT('h2)
	) name5815 (
		_w2520_,
		_w6277_,
		_w6278_
	);
	LUT3 #(
		.INIT('h0d)
	) name5816 (
		\P1_reg1_reg[1]/NET0131 ,
		_w2525_,
		_w6278_,
		_w6279_
	);
	LUT3 #(
		.INIT('h10)
	) name5817 (
		_w6274_,
		_w6276_,
		_w6279_,
		_w6280_
	);
	LUT4 #(
		.INIT('h1311)
	) name5818 (
		_w1731_,
		_w6269_,
		_w6272_,
		_w6280_,
		_w6281_
	);
	LUT3 #(
		.INIT('hce)
	) name5819 (
		\P1_state_reg[0]/NET0131 ,
		_w6268_,
		_w6281_,
		_w6282_
	);
	LUT4 #(
		.INIT('hd070)
	) name5820 (
		\P1_state_reg[0]/NET0131 ,
		\P2_IR_reg[23]/NET0131 ,
		\P2_reg3_reg[0]/NET0131 ,
		_w1188_,
		_w6283_
	);
	LUT4 #(
		.INIT('h2000)
	) name5821 (
		\P2_reg3_reg[0]/NET0131 ,
		_w1189_,
		_w1352_,
		_w1356_,
		_w6284_
	);
	LUT4 #(
		.INIT('haaa8)
	) name5822 (
		\P2_reg3_reg[0]/NET0131 ,
		_w1361_,
		_w1363_,
		_w1368_,
		_w6285_
	);
	LUT4 #(
		.INIT('h8400)
	) name5823 (
		_w814_,
		_w1411_,
		_w1413_,
		_w1435_,
		_w6286_
	);
	LUT3 #(
		.INIT('ha8)
	) name5824 (
		_w1191_,
		_w6285_,
		_w6286_,
		_w6287_
	);
	LUT4 #(
		.INIT('h30a0)
	) name5825 (
		\P2_reg3_reg[0]/NET0131 ,
		_w1305_,
		_w1447_,
		_w1411_,
		_w6288_
	);
	LUT3 #(
		.INIT('h20)
	) name5826 (
		\P2_reg3_reg[0]/NET0131 ,
		_w1184_,
		_w1190_,
		_w6289_
	);
	LUT3 #(
		.INIT('h0b)
	) name5827 (
		_w826_,
		_w1233_,
		_w6289_,
		_w6290_
	);
	LUT4 #(
		.INIT('h02aa)
	) name5828 (
		\P2_reg3_reg[0]/NET0131 ,
		_w1361_,
		_w1363_,
		_w1368_,
		_w6291_
	);
	LUT4 #(
		.INIT('h5400)
	) name5829 (
		_w826_,
		_w1361_,
		_w1363_,
		_w1368_,
		_w6292_
	);
	LUT3 #(
		.INIT('ha8)
	) name5830 (
		_w1442_,
		_w6291_,
		_w6292_,
		_w6293_
	);
	LUT4 #(
		.INIT('h003a)
	) name5831 (
		\P2_reg3_reg[0]/NET0131 ,
		_w1305_,
		_w1369_,
		_w5849_,
		_w6294_
	);
	LUT4 #(
		.INIT('h0100)
	) name5832 (
		_w6288_,
		_w6293_,
		_w6294_,
		_w6290_,
		_w6295_
	);
	LUT4 #(
		.INIT('h1311)
	) name5833 (
		_w1359_,
		_w6284_,
		_w6287_,
		_w6295_,
		_w6296_
	);
	LUT3 #(
		.INIT('hce)
	) name5834 (
		\P1_state_reg[0]/NET0131 ,
		_w6283_,
		_w6296_,
		_w6297_
	);
	LUT2 #(
		.INIT('h2)
	) name5835 (
		\P1_reg2_reg[1]/NET0131 ,
		_w2462_,
		_w6298_
	);
	LUT4 #(
		.INIT('h2000)
	) name5836 (
		\P1_reg2_reg[1]/NET0131 ,
		_w1723_,
		_w1727_,
		_w1730_,
		_w6299_
	);
	LUT2 #(
		.INIT('h2)
	) name5837 (
		\P1_reg2_reg[1]/NET0131 ,
		_w1741_,
		_w6300_
	);
	LUT4 #(
		.INIT('hddd1)
	) name5838 (
		\P1_reg2_reg[1]/NET0131 ,
		_w1741_,
		_w6083_,
		_w6084_,
		_w6301_
	);
	LUT2 #(
		.INIT('h2)
	) name5839 (
		_w2424_,
		_w6301_,
		_w6302_
	);
	LUT4 #(
		.INIT('h08a2)
	) name5840 (
		_w1741_,
		_w2086_,
		_w2089_,
		_w3189_,
		_w6303_
	);
	LUT3 #(
		.INIT('ha8)
	) name5841 (
		_w2388_,
		_w6300_,
		_w6303_,
		_w6304_
	);
	LUT4 #(
		.INIT('h1dd1)
	) name5842 (
		\P1_reg2_reg[1]/NET0131 ,
		_w1741_,
		_w2090_,
		_w3189_,
		_w6305_
	);
	LUT2 #(
		.INIT('h2)
	) name5843 (
		_w2292_,
		_w6305_,
		_w6306_
	);
	LUT2 #(
		.INIT('h2)
	) name5844 (
		_w1741_,
		_w6277_,
		_w6307_
	);
	LUT4 #(
		.INIT('ha2a0)
	) name5845 (
		\P1_reg2_reg[1]/NET0131 ,
		_w1741_,
		_w2450_,
		_w2452_,
		_w6308_
	);
	LUT4 #(
		.INIT('h0008)
	) name5846 (
		\P1_reg3_reg[1]/NET0131 ,
		_w2284_,
		_w2288_,
		_w2291_,
		_w6309_
	);
	LUT3 #(
		.INIT('h01)
	) name5847 (
		_w6308_,
		_w6307_,
		_w6309_,
		_w6310_
	);
	LUT3 #(
		.INIT('h10)
	) name5848 (
		_w6304_,
		_w6306_,
		_w6310_,
		_w6311_
	);
	LUT4 #(
		.INIT('h1311)
	) name5849 (
		_w1731_,
		_w6299_,
		_w6302_,
		_w6311_,
		_w6312_
	);
	LUT3 #(
		.INIT('hce)
	) name5850 (
		\P1_state_reg[0]/NET0131 ,
		_w6298_,
		_w6312_,
		_w6313_
	);
	LUT4 #(
		.INIT('hd070)
	) name5851 (
		\P1_state_reg[0]/NET0131 ,
		\P2_IR_reg[23]/NET0131 ,
		\P2_reg1_reg[0]/NET0131 ,
		_w1188_,
		_w6314_
	);
	LUT4 #(
		.INIT('h2000)
	) name5852 (
		\P2_reg1_reg[0]/NET0131 ,
		_w1189_,
		_w1352_,
		_w1356_,
		_w6315_
	);
	LUT4 #(
		.INIT('h6f00)
	) name5853 (
		_w814_,
		_w1413_,
		_w1435_,
		_w1507_,
		_w6316_
	);
	LUT4 #(
		.INIT('h5455)
	) name5854 (
		\P2_reg1_reg[0]/NET0131 ,
		_w1361_,
		_w1363_,
		_w1368_,
		_w6317_
	);
	LUT2 #(
		.INIT('h2)
	) name5855 (
		_w1191_,
		_w6317_,
		_w6318_
	);
	LUT2 #(
		.INIT('h4)
	) name5856 (
		_w6316_,
		_w6318_,
		_w6319_
	);
	LUT4 #(
		.INIT('haa02)
	) name5857 (
		\P2_reg1_reg[0]/NET0131 ,
		_w1361_,
		_w1363_,
		_w1368_,
		_w6320_
	);
	LUT4 #(
		.INIT('h003a)
	) name5858 (
		\P2_reg1_reg[0]/NET0131 ,
		_w1305_,
		_w1516_,
		_w6151_,
		_w6321_
	);
	LUT2 #(
		.INIT('h2)
	) name5859 (
		\P2_reg1_reg[0]/NET0131 ,
		_w1684_,
		_w6322_
	);
	LUT4 #(
		.INIT('h0054)
	) name5860 (
		_w826_,
		_w1361_,
		_w1363_,
		_w1368_,
		_w6323_
	);
	LUT3 #(
		.INIT('ha8)
	) name5861 (
		_w1442_,
		_w6320_,
		_w6323_,
		_w6324_
	);
	LUT4 #(
		.INIT('h3a00)
	) name5862 (
		\P2_reg1_reg[0]/NET0131 ,
		_w1305_,
		_w1507_,
		_w1530_,
		_w6325_
	);
	LUT4 #(
		.INIT('h0001)
	) name5863 (
		_w6321_,
		_w6322_,
		_w6324_,
		_w6325_,
		_w6326_
	);
	LUT4 #(
		.INIT('h1311)
	) name5864 (
		_w1359_,
		_w6315_,
		_w6319_,
		_w6326_,
		_w6327_
	);
	LUT3 #(
		.INIT('hce)
	) name5865 (
		\P1_state_reg[0]/NET0131 ,
		_w6314_,
		_w6327_,
		_w6328_
	);
	LUT4 #(
		.INIT('hd070)
	) name5866 (
		\P1_state_reg[0]/NET0131 ,
		\P2_IR_reg[23]/NET0131 ,
		\P2_reg2_reg[0]/NET0131 ,
		_w1188_,
		_w6329_
	);
	LUT4 #(
		.INIT('h2000)
	) name5867 (
		\P2_reg2_reg[0]/NET0131 ,
		_w1189_,
		_w1352_,
		_w1356_,
		_w6330_
	);
	LUT4 #(
		.INIT('haa02)
	) name5868 (
		\P2_reg2_reg[0]/NET0131 ,
		_w1361_,
		_w1363_,
		_w1368_,
		_w6331_
	);
	LUT4 #(
		.INIT('h9000)
	) name5869 (
		_w814_,
		_w1413_,
		_w1435_,
		_w1516_,
		_w6332_
	);
	LUT3 #(
		.INIT('ha8)
	) name5870 (
		_w1191_,
		_w6331_,
		_w6332_,
		_w6333_
	);
	LUT4 #(
		.INIT('h5455)
	) name5871 (
		\P2_reg2_reg[0]/NET0131 ,
		_w1361_,
		_w1363_,
		_w1368_,
		_w6334_
	);
	LUT4 #(
		.INIT('h0200)
	) name5872 (
		_w826_,
		_w1361_,
		_w1363_,
		_w1368_,
		_w6335_
	);
	LUT2 #(
		.INIT('h2)
	) name5873 (
		_w1442_,
		_w6335_,
		_w6336_
	);
	LUT3 #(
		.INIT('h07)
	) name5874 (
		_w1305_,
		_w1507_,
		_w6151_,
		_w6337_
	);
	LUT3 #(
		.INIT('h54)
	) name5875 (
		_w6334_,
		_w6336_,
		_w6337_,
		_w6338_
	);
	LUT4 #(
		.INIT('h3a00)
	) name5876 (
		\P2_reg2_reg[0]/NET0131 ,
		_w1305_,
		_w1516_,
		_w1530_,
		_w6339_
	);
	LUT3 #(
		.INIT('h80)
	) name5877 (
		\P2_reg3_reg[0]/NET0131 ,
		_w1229_,
		_w1232_,
		_w6340_
	);
	LUT3 #(
		.INIT('h20)
	) name5878 (
		\P2_reg2_reg[0]/NET0131 ,
		_w1184_,
		_w1190_,
		_w6341_
	);
	LUT2 #(
		.INIT('h1)
	) name5879 (
		_w6340_,
		_w6341_,
		_w6342_
	);
	LUT2 #(
		.INIT('h4)
	) name5880 (
		_w6339_,
		_w6342_,
		_w6343_
	);
	LUT4 #(
		.INIT('ha8aa)
	) name5881 (
		_w1359_,
		_w6338_,
		_w6333_,
		_w6343_,
		_w6344_
	);
	LUT4 #(
		.INIT('heeec)
	) name5882 (
		\P1_state_reg[0]/NET0131 ,
		_w6329_,
		_w6330_,
		_w6344_,
		_w6345_
	);
	LUT4 #(
		.INIT('hd070)
	) name5883 (
		\P1_state_reg[0]/NET0131 ,
		\P2_IR_reg[23]/NET0131 ,
		\P2_reg0_reg[0]/NET0131 ,
		_w1188_,
		_w6346_
	);
	LUT4 #(
		.INIT('h2000)
	) name5884 (
		\P2_reg0_reg[0]/NET0131 ,
		_w1189_,
		_w1352_,
		_w1356_,
		_w6347_
	);
	LUT4 #(
		.INIT('h02aa)
	) name5885 (
		\P2_reg0_reg[0]/NET0131 ,
		_w1361_,
		_w1363_,
		_w1368_,
		_w6348_
	);
	LUT4 #(
		.INIT('h8400)
	) name5886 (
		_w814_,
		_w1369_,
		_w1413_,
		_w1435_,
		_w6349_
	);
	LUT3 #(
		.INIT('ha8)
	) name5887 (
		_w1191_,
		_w6348_,
		_w6349_,
		_w6350_
	);
	LUT4 #(
		.INIT('haaa8)
	) name5888 (
		\P2_reg0_reg[0]/NET0131 ,
		_w1361_,
		_w1363_,
		_w1368_,
		_w6351_
	);
	LUT4 #(
		.INIT('h0001)
	) name5889 (
		_w826_,
		_w1361_,
		_w1363_,
		_w1368_,
		_w6352_
	);
	LUT2 #(
		.INIT('h2)
	) name5890 (
		\P2_reg0_reg[0]/NET0131 ,
		_w1684_,
		_w6353_
	);
	LUT4 #(
		.INIT('h0057)
	) name5891 (
		_w1442_,
		_w6351_,
		_w6352_,
		_w6353_,
		_w6354_
	);
	LUT4 #(
		.INIT('h3a00)
	) name5892 (
		\P2_reg0_reg[0]/NET0131 ,
		_w1305_,
		_w1369_,
		_w1447_,
		_w6355_
	);
	LUT4 #(
		.INIT('h003a)
	) name5893 (
		\P2_reg0_reg[0]/NET0131 ,
		_w1305_,
		_w1411_,
		_w5849_,
		_w6356_
	);
	LUT3 #(
		.INIT('h10)
	) name5894 (
		_w6355_,
		_w6356_,
		_w6354_,
		_w6357_
	);
	LUT4 #(
		.INIT('h1311)
	) name5895 (
		_w1359_,
		_w6347_,
		_w6350_,
		_w6357_,
		_w6358_
	);
	LUT3 #(
		.INIT('hce)
	) name5896 (
		\P1_state_reg[0]/NET0131 ,
		_w6346_,
		_w6358_,
		_w6359_
	);
	LUT4 #(
		.INIT('h7800)
	) name5897 (
		_w2084_,
		_w2085_,
		_w2089_,
		_w2285_,
		_w6360_
	);
	LUT2 #(
		.INIT('h4)
	) name5898 (
		_w1747_,
		_w2424_,
		_w6361_
	);
	LUT4 #(
		.INIT('h060f)
	) name5899 (
		_w2077_,
		_w2399_,
		_w6360_,
		_w6361_,
		_w6362_
	);
	LUT2 #(
		.INIT('h4)
	) name5900 (
		_w2089_,
		_w2284_,
		_w6363_
	);
	LUT3 #(
		.INIT('he0)
	) name5901 (
		_w2451_,
		_w2644_,
		_w6363_,
		_w6364_
	);
	LUT4 #(
		.INIT('hcc08)
	) name5902 (
		_w2644_,
		_w5244_,
		_w6362_,
		_w6364_,
		_w6365_
	);
	LUT3 #(
		.INIT('he0)
	) name5903 (
		_w2644_,
		_w3574_,
		_w5244_,
		_w6366_
	);
	LUT3 #(
		.INIT('h2a)
	) name5904 (
		\P1_reg3_reg[0]/NET0131 ,
		_w3475_,
		_w6366_,
		_w6367_
	);
	LUT2 #(
		.INIT('he)
	) name5905 (
		_w6365_,
		_w6367_,
		_w6368_
	);
	LUT4 #(
		.INIT('h0008)
	) name5906 (
		\P1_reg3_reg[0]/NET0131 ,
		_w2284_,
		_w2288_,
		_w2291_,
		_w6369_
	);
	LUT2 #(
		.INIT('h4)
	) name5907 (
		_w2089_,
		_w2452_,
		_w6370_
	);
	LUT4 #(
		.INIT('h050d)
	) name5908 (
		_w1741_,
		_w6362_,
		_w6369_,
		_w6370_,
		_w6371_
	);
	LUT3 #(
		.INIT('h2a)
	) name5909 (
		\P1_reg2_reg[0]/NET0131 ,
		_w5244_,
		_w5248_,
		_w6372_
	);
	LUT3 #(
		.INIT('hf2)
	) name5910 (
		_w5244_,
		_w6371_,
		_w6372_,
		_w6373_
	);
	LUT4 #(
		.INIT('h8808)
	) name5911 (
		_w2883_,
		_w5244_,
		_w6362_,
		_w6370_,
		_w6374_
	);
	LUT3 #(
		.INIT('he0)
	) name5912 (
		_w2883_,
		_w3574_,
		_w5244_,
		_w6375_
	);
	LUT3 #(
		.INIT('h2a)
	) name5913 (
		\P1_reg0_reg[0]/NET0131 ,
		_w3408_,
		_w6375_,
		_w6376_
	);
	LUT2 #(
		.INIT('he)
	) name5914 (
		_w6374_,
		_w6376_,
		_w6377_
	);
	LUT4 #(
		.INIT('h8808)
	) name5915 (
		_w2520_,
		_w5244_,
		_w6362_,
		_w6370_,
		_w6378_
	);
	LUT3 #(
		.INIT('he0)
	) name5916 (
		_w2520_,
		_w3574_,
		_w5244_,
		_w6379_
	);
	LUT3 #(
		.INIT('h2a)
	) name5917 (
		\P1_reg1_reg[0]/NET0131 ,
		_w3744_,
		_w6379_,
		_w6380_
	);
	LUT2 #(
		.INIT('he)
	) name5918 (
		_w6378_,
		_w6380_,
		_w6381_
	);
	LUT4 #(
		.INIT('h1f00)
	) name5919 (
		_w546_,
		_w1158_,
		_w1411_,
		_w1442_,
		_w6382_
	);
	LUT4 #(
		.INIT('h67ef)
	) name5920 (
		_w1179_,
		_w1183_,
		_w1190_,
		_w1228_,
		_w6383_
	);
	LUT4 #(
		.INIT('h001f)
	) name5921 (
		_w1361_,
		_w1363_,
		_w1368_,
		_w6383_,
		_w6384_
	);
	LUT4 #(
		.INIT('h00fe)
	) name5922 (
		_w1361_,
		_w1363_,
		_w1368_,
		_w5849_,
		_w6385_
	);
	LUT3 #(
		.INIT('h70)
	) name5923 (
		_w1352_,
		_w1356_,
		_w1503_,
		_w6386_
	);
	LUT2 #(
		.INIT('h4)
	) name5924 (
		_w1233_,
		_w6386_,
		_w6387_
	);
	LUT3 #(
		.INIT('h10)
	) name5925 (
		_w6385_,
		_w6384_,
		_w6387_,
		_w6388_
	);
	LUT3 #(
		.INIT('h8a)
	) name5926 (
		\P2_reg0_reg[30]/NET0131 ,
		_w6382_,
		_w6388_,
		_w6389_
	);
	LUT3 #(
		.INIT('hb0)
	) name5927 (
		_w1110_,
		_w1137_,
		_w1191_,
		_w6390_
	);
	LUT4 #(
		.INIT('hb000)
	) name5928 (
		_w1163_,
		_w1519_,
		_w1681_,
		_w6390_,
		_w6391_
	);
	LUT4 #(
		.INIT('h1000)
	) name5929 (
		_w546_,
		_w1158_,
		_w1411_,
		_w1442_,
		_w6392_
	);
	LUT4 #(
		.INIT('hcc80)
	) name5930 (
		_w1369_,
		_w6386_,
		_w6391_,
		_w6392_,
		_w6393_
	);
	LUT2 #(
		.INIT('he)
	) name5931 (
		_w6389_,
		_w6393_,
		_w6394_
	);
	LUT4 #(
		.INIT('hed00)
	) name5932 (
		\P1_datao_reg[31]/NET0131 ,
		_w546_,
		_w1148_,
		_w1411_,
		_w6395_
	);
	LUT4 #(
		.INIT('h0a8a)
	) name5933 (
		\P2_reg0_reg[31]/NET0131 ,
		_w1442_,
		_w6388_,
		_w6395_,
		_w6396_
	);
	LUT3 #(
		.INIT('h80)
	) name5934 (
		_w1149_,
		_w1411_,
		_w1442_,
		_w6397_
	);
	LUT4 #(
		.INIT('hcc80)
	) name5935 (
		_w1369_,
		_w6386_,
		_w6391_,
		_w6397_,
		_w6398_
	);
	LUT2 #(
		.INIT('he)
	) name5936 (
		_w6396_,
		_w6398_,
		_w6399_
	);
	LUT3 #(
		.INIT('h10)
	) name5937 (
		_w546_,
		_w1158_,
		_w2471_,
		_w6400_
	);
	LUT4 #(
		.INIT('hcc80)
	) name5938 (
		_w1507_,
		_w6386_,
		_w6391_,
		_w6400_,
		_w6401_
	);
	LUT4 #(
		.INIT('hcdef)
	) name5939 (
		_w1179_,
		_w1183_,
		_w1190_,
		_w1228_,
		_w6402_
	);
	LUT4 #(
		.INIT('h00ef)
	) name5940 (
		_w1361_,
		_w1363_,
		_w1368_,
		_w6402_,
		_w6403_
	);
	LUT2 #(
		.INIT('h2)
	) name5941 (
		_w6386_,
		_w6403_,
		_w6404_
	);
	LUT3 #(
		.INIT('h2a)
	) name5942 (
		\P2_reg1_reg[30]/NET0131 ,
		_w6153_,
		_w6404_,
		_w6405_
	);
	LUT2 #(
		.INIT('he)
	) name5943 (
		_w6401_,
		_w6405_,
		_w6406_
	);
	LUT4 #(
		.INIT('he0c0)
	) name5944 (
		_w1516_,
		_w2510_,
		_w6386_,
		_w6391_,
		_w6407_
	);
	LUT4 #(
		.INIT('h00ef)
	) name5945 (
		_w1361_,
		_w1363_,
		_w1368_,
		_w6151_,
		_w6408_
	);
	LUT4 #(
		.INIT('h00f1)
	) name5946 (
		_w1361_,
		_w1363_,
		_w1368_,
		_w6402_,
		_w6409_
	);
	LUT4 #(
		.INIT('haaa2)
	) name5947 (
		\P2_reg2_reg[30]/NET0131 ,
		_w6386_,
		_w6409_,
		_w6408_,
		_w6410_
	);
	LUT4 #(
		.INIT('ha8aa)
	) name5948 (
		\P2_reg2_reg[30]/NET0131 ,
		_w1361_,
		_w1363_,
		_w1368_,
		_w6411_
	);
	LUT4 #(
		.INIT('h1000)
	) name5949 (
		_w1361_,
		_w1363_,
		_w1368_,
		_w6386_,
		_w6412_
	);
	LUT4 #(
		.INIT('h0e0f)
	) name5950 (
		_w546_,
		_w1158_,
		_w6411_,
		_w6412_,
		_w6413_
	);
	LUT3 #(
		.INIT('h31)
	) name5951 (
		_w1442_,
		_w6410_,
		_w6413_,
		_w6414_
	);
	LUT2 #(
		.INIT('hb)
	) name5952 (
		_w6407_,
		_w6414_,
		_w6415_
	);
	LUT4 #(
		.INIT('h1200)
	) name5953 (
		\P1_datao_reg[31]/NET0131 ,
		_w546_,
		_w1148_,
		_w2471_,
		_w6416_
	);
	LUT4 #(
		.INIT('hcc80)
	) name5954 (
		_w1507_,
		_w6386_,
		_w6391_,
		_w6416_,
		_w6417_
	);
	LUT3 #(
		.INIT('h2a)
	) name5955 (
		\P2_reg1_reg[31]/NET0131 ,
		_w6153_,
		_w6404_,
		_w6418_
	);
	LUT2 #(
		.INIT('he)
	) name5956 (
		_w6417_,
		_w6418_,
		_w6419_
	);
	LUT4 #(
		.INIT('haaa2)
	) name5957 (
		\P2_reg2_reg[31]/NET0131 ,
		_w6386_,
		_w6409_,
		_w6408_,
		_w6420_
	);
	LUT4 #(
		.INIT('ha8aa)
	) name5958 (
		\P2_reg2_reg[31]/NET0131 ,
		_w1361_,
		_w1363_,
		_w1368_,
		_w6421_
	);
	LUT4 #(
		.INIT('h1200)
	) name5959 (
		\P1_datao_reg[31]/NET0131 ,
		_w546_,
		_w1148_,
		_w6412_,
		_w6422_
	);
	LUT4 #(
		.INIT('h1113)
	) name5960 (
		_w1442_,
		_w6420_,
		_w6421_,
		_w6422_,
		_w6423_
	);
	LUT2 #(
		.INIT('hb)
	) name5961 (
		_w6407_,
		_w6423_,
		_w6424_
	);
	LUT2 #(
		.INIT('h8)
	) name5962 (
		\P1_state_reg[0]/NET0131 ,
		_w1744_,
		_w6425_
	);
	LUT4 #(
		.INIT('hff54)
	) name5963 (
		\P1_state_reg[0]/NET0131 ,
		_w1907_,
		_w1929_,
		_w6425_,
		_w6426_
	);
	LUT2 #(
		.INIT('h2)
	) name5964 (
		\P1_state_reg[0]/NET0131 ,
		_w1354_,
		_w6427_
	);
	LUT3 #(
		.INIT('h0b)
	) name5965 (
		\P1_state_reg[0]/NET0131 ,
		_w1026_,
		_w6427_,
		_w6428_
	);
	LUT4 #(
		.INIT('h8882)
	) name5966 (
		\P1_state_reg[0]/NET0131 ,
		\P2_IR_reg[26]/NET0131 ,
		_w1185_,
		_w1351_,
		_w6429_
	);
	LUT3 #(
		.INIT('h0b)
	) name5967 (
		\P1_state_reg[0]/NET0131 ,
		_w1058_,
		_w6429_,
		_w6430_
	);
	LUT3 #(
		.INIT('h82)
	) name5968 (
		\P1_state_reg[0]/NET0131 ,
		\P2_IR_reg[27]/NET0131 ,
		_w544_,
		_w6431_
	);
	LUT3 #(
		.INIT('hf1)
	) name5969 (
		\P1_state_reg[0]/NET0131 ,
		_w1078_,
		_w6431_,
		_w6432_
	);
	LUT3 #(
		.INIT('h48)
	) name5970 (
		\P1_IR_reg[25]/NET0131 ,
		\P1_state_reg[0]/NET0131 ,
		_w475_,
		_w6433_
	);
	LUT4 #(
		.INIT('hff54)
	) name5971 (
		\P1_state_reg[0]/NET0131 ,
		_w1839_,
		_w1870_,
		_w6433_,
		_w6434_
	);
	LUT3 #(
		.INIT('h48)
	) name5972 (
		\P1_IR_reg[26]/NET0131 ,
		\P1_state_reg[0]/NET0131 ,
		_w484_,
		_w6435_
	);
	LUT3 #(
		.INIT('hf1)
	) name5973 (
		\P1_state_reg[0]/NET0131 ,
		_w1899_,
		_w6435_,
		_w6436_
	);
	LUT4 #(
		.INIT('h0200)
	) name5974 (
		\P1_state_reg[0]/NET0131 ,
		\P2_IR_reg[27]/NET0131 ,
		\P2_IR_reg[30]/NET0131 ,
		\P2_IR_reg[31]/NET0131 ,
		_w6437_
	);
	LUT4 #(
		.INIT('h8000)
	) name5975 (
		_w513_,
		_w531_,
		_w542_,
		_w6437_,
		_w6438_
	);
	LUT3 #(
		.INIT('h80)
	) name5976 (
		_w540_,
		_w541_,
		_w6438_,
		_w6439_
	);
	LUT4 #(
		.INIT('hff12)
	) name5977 (
		\P1_datao_reg[31]/NET0131 ,
		\P1_state_reg[0]/NET0131 ,
		_w1148_,
		_w6439_,
		_w6440_
	);
	LUT2 #(
		.INIT('h8)
	) name5978 (
		\P1_state_reg[0]/NET0131 ,
		_w877_,
		_w6441_
	);
	LUT4 #(
		.INIT('hff54)
	) name5979 (
		\P1_state_reg[0]/NET0131 ,
		_w868_,
		_w876_,
		_w6441_,
		_w6442_
	);
	LUT3 #(
		.INIT('h0b)
	) name5980 (
		\P1_state_reg[0]/NET0131 ,
		_w981_,
		_w1503_,
		_w6443_
	);
	LUT3 #(
		.INIT('h82)
	) name5981 (
		\P1_state_reg[0]/NET0131 ,
		\P2_IR_reg[10]/NET0131 ,
		_w700_,
		_w6444_
	);
	LUT4 #(
		.INIT('hff54)
	) name5982 (
		\P1_state_reg[0]/NET0131 ,
		_w695_,
		_w697_,
		_w6444_,
		_w6445_
	);
	LUT3 #(
		.INIT('h28)
	) name5983 (
		\P1_state_reg[0]/NET0131 ,
		\P2_IR_reg[11]/NET0131 ,
		_w682_,
		_w6446_
	);
	LUT3 #(
		.INIT('hf1)
	) name5984 (
		\P1_state_reg[0]/NET0131 ,
		_w681_,
		_w6446_,
		_w6447_
	);
	LUT4 #(
		.INIT('h2228)
	) name5985 (
		\P1_state_reg[0]/NET0131 ,
		\P2_IR_reg[12]/NET0131 ,
		_w662_,
		_w663_,
		_w6448_
	);
	LUT3 #(
		.INIT('hf1)
	) name5986 (
		\P1_state_reg[0]/NET0131 ,
		_w661_,
		_w6448_,
		_w6449_
	);
	LUT4 #(
		.INIT('h8828)
	) name5987 (
		\P1_state_reg[0]/NET0131 ,
		\P2_IR_reg[13]/NET0131 ,
		\P2_IR_reg[31]/NET0131 ,
		_w498_,
		_w6450_
	);
	LUT3 #(
		.INIT('hf1)
	) name5988 (
		\P1_state_reg[0]/NET0131 ,
		_w642_,
		_w6450_,
		_w6451_
	);
	LUT2 #(
		.INIT('h8)
	) name5989 (
		\P1_state_reg[0]/NET0131 ,
		_w613_,
		_w6452_
	);
	LUT3 #(
		.INIT('hf1)
	) name5990 (
		\P1_state_reg[0]/NET0131 ,
		_w612_,
		_w6452_,
		_w6453_
	);
	LUT4 #(
		.INIT('h8828)
	) name5991 (
		\P1_state_reg[0]/NET0131 ,
		\P2_IR_reg[15]/NET0131 ,
		\P2_IR_reg[31]/NET0131 ,
		_w540_,
		_w6454_
	);
	LUT4 #(
		.INIT('hff54)
	) name5992 (
		\P1_state_reg[0]/NET0131 ,
		_w548_,
		_w591_,
		_w6454_,
		_w6455_
	);
	LUT2 #(
		.INIT('h8)
	) name5993 (
		\P1_state_reg[0]/NET0131 ,
		_w858_,
		_w6456_
	);
	LUT4 #(
		.INIT('hff54)
	) name5994 (
		\P1_state_reg[0]/NET0131 ,
		_w847_,
		_w857_,
		_w6456_,
		_w6457_
	);
	LUT3 #(
		.INIT('h82)
	) name5995 (
		\P1_state_reg[0]/NET0131 ,
		\P2_IR_reg[18]/NET0131 ,
		_w922_,
		_w6458_
	);
	LUT4 #(
		.INIT('hff54)
	) name5996 (
		\P1_state_reg[0]/NET0131 ,
		_w912_,
		_w920_,
		_w6458_,
		_w6459_
	);
	LUT2 #(
		.INIT('h2)
	) name5997 (
		\P1_state_reg[0]/NET0131 ,
		_w900_,
		_w6460_
	);
	LUT3 #(
		.INIT('hf1)
	) name5998 (
		\P1_state_reg[0]/NET0131 ,
		_w899_,
		_w6460_,
		_w6461_
	);
	LUT4 #(
		.INIT('h28a0)
	) name5999 (
		\P1_state_reg[0]/NET0131 ,
		\P2_IR_reg[0]/NET0131 ,
		\P2_IR_reg[1]/NET0131 ,
		\P2_IR_reg[31]/NET0131 ,
		_w6462_
	);
	LUT3 #(
		.INIT('hf4)
	) name6000 (
		\P1_state_reg[0]/NET0131 ,
		_w817_,
		_w6462_,
		_w6463_
	);
	LUT3 #(
		.INIT('h28)
	) name6001 (
		\P1_state_reg[0]/NET0131 ,
		\P2_IR_reg[20]/NET0131 ,
		_w1182_,
		_w6464_
	);
	LUT3 #(
		.INIT('h0b)
	) name6002 (
		\P1_state_reg[0]/NET0131 ,
		_w962_,
		_w6464_,
		_w6465_
	);
	LUT3 #(
		.INIT('h28)
	) name6003 (
		\P1_state_reg[0]/NET0131 ,
		\P2_IR_reg[21]/NET0131 ,
		_w1178_,
		_w6466_
	);
	LUT4 #(
		.INIT('h00fe)
	) name6004 (
		\P1_state_reg[0]/NET0131 ,
		_w935_,
		_w944_,
		_w6466_,
		_w6467_
	);
	LUT3 #(
		.INIT('h28)
	) name6005 (
		\P1_state_reg[0]/NET0131 ,
		\P2_IR_reg[22]/NET0131 ,
		_w1185_,
		_w6468_
	);
	LUT3 #(
		.INIT('hf1)
	) name6006 (
		\P1_state_reg[0]/NET0131 ,
		_w999_,
		_w6468_,
		_w6469_
	);
	LUT3 #(
		.INIT('h28)
	) name6007 (
		\P1_state_reg[0]/NET0131 ,
		\P2_IR_reg[24]/NET0131 ,
		_w534_,
		_w6470_
	);
	LUT3 #(
		.INIT('hf1)
	) name6008 (
		\P1_state_reg[0]/NET0131 ,
		_w1041_,
		_w6470_,
		_w6471_
	);
	LUT4 #(
		.INIT('h2228)
	) name6009 (
		\P1_state_reg[0]/NET0131 ,
		\P2_IR_reg[28]/NET0131 ,
		_w534_,
		_w536_,
		_w6472_
	);
	LUT3 #(
		.INIT('hf1)
	) name6010 (
		\P1_state_reg[0]/NET0131 ,
		_w1124_,
		_w6472_,
		_w6473_
	);
	LUT2 #(
		.INIT('h8)
	) name6011 (
		\P1_state_reg[0]/NET0131 ,
		_w505_,
		_w6474_
	);
	LUT3 #(
		.INIT('hf1)
	) name6012 (
		\P1_state_reg[0]/NET0131 ,
		_w1107_,
		_w6474_,
		_w6475_
	);
	LUT2 #(
		.INIT('h2)
	) name6013 (
		\P1_state_reg[0]/NET0131 ,
		_w806_,
		_w6476_
	);
	LUT3 #(
		.INIT('hf1)
	) name6014 (
		\P1_state_reg[0]/NET0131 ,
		_w805_,
		_w6476_,
		_w6477_
	);
	LUT3 #(
		.INIT('h82)
	) name6015 (
		\P1_state_reg[0]/NET0131 ,
		\P2_IR_reg[30]/NET0131 ,
		_w516_,
		_w6478_
	);
	LUT3 #(
		.INIT('hf1)
	) name6016 (
		\P1_state_reg[0]/NET0131 ,
		_w1158_,
		_w6478_,
		_w6479_
	);
	LUT3 #(
		.INIT('h28)
	) name6017 (
		\P1_state_reg[0]/NET0131 ,
		\P2_IR_reg[3]/NET0131 ,
		_w794_,
		_w6480_
	);
	LUT3 #(
		.INIT('hf4)
	) name6018 (
		\P1_state_reg[0]/NET0131 ,
		_w796_,
		_w6480_,
		_w6481_
	);
	LUT4 #(
		.INIT('ha028)
	) name6019 (
		\P1_state_reg[0]/NET0131 ,
		\P2_IR_reg[31]/NET0131 ,
		\P2_IR_reg[4]/NET0131 ,
		_w496_,
		_w6482_
	);
	LUT3 #(
		.INIT('hf1)
	) name6020 (
		\P1_state_reg[0]/NET0131 ,
		_w783_,
		_w6482_,
		_w6483_
	);
	LUT2 #(
		.INIT('h2)
	) name6021 (
		\P1_state_reg[0]/NET0131 ,
		_w773_,
		_w6484_
	);
	LUT3 #(
		.INIT('hf1)
	) name6022 (
		\P1_state_reg[0]/NET0131 ,
		_w772_,
		_w6484_,
		_w6485_
	);
	LUT3 #(
		.INIT('h82)
	) name6023 (
		\P1_state_reg[0]/NET0131 ,
		\P2_IR_reg[6]/NET0131 ,
		_w750_,
		_w6486_
	);
	LUT3 #(
		.INIT('hf1)
	) name6024 (
		\P1_state_reg[0]/NET0131 ,
		_w749_,
		_w6486_,
		_w6487_
	);
	LUT2 #(
		.INIT('h8)
	) name6025 (
		\P1_state_reg[0]/NET0131 ,
		_w762_,
		_w6488_
	);
	LUT3 #(
		.INIT('hf1)
	) name6026 (
		\P1_state_reg[0]/NET0131 ,
		_w761_,
		_w6488_,
		_w6489_
	);
	LUT3 #(
		.INIT('h28)
	) name6027 (
		\P1_state_reg[0]/NET0131 ,
		\P2_IR_reg[8]/NET0131 ,
		_w729_,
		_w6490_
	);
	LUT3 #(
		.INIT('hf1)
	) name6028 (
		\P1_state_reg[0]/NET0131 ,
		_w728_,
		_w6490_,
		_w6491_
	);
	LUT3 #(
		.INIT('h28)
	) name6029 (
		\P1_state_reg[0]/NET0131 ,
		\P2_IR_reg[9]/NET0131 ,
		_w662_,
		_w6492_
	);
	LUT4 #(
		.INIT('hff54)
	) name6030 (
		\P1_state_reg[0]/NET0131 ,
		_w713_,
		_w715_,
		_w6492_,
		_w6493_
	);
	LUT3 #(
		.INIT('h48)
	) name6031 (
		\P1_IR_reg[10]/NET0131 ,
		\P1_state_reg[0]/NET0131 ,
		_w2010_,
		_w6494_
	);
	LUT4 #(
		.INIT('hff54)
	) name6032 (
		\P1_state_reg[0]/NET0131 ,
		_w2025_,
		_w2027_,
		_w6494_,
		_w6495_
	);
	LUT4 #(
		.INIT('ha060)
	) name6033 (
		\P1_IR_reg[11]/NET0131 ,
		\P1_IR_reg[31]/NET0131 ,
		\P1_state_reg[0]/NET0131 ,
		_w1718_,
		_w6496_
	);
	LUT3 #(
		.INIT('hf1)
	) name6034 (
		\P1_state_reg[0]/NET0131 ,
		_w2003_,
		_w6496_,
		_w6497_
	);
	LUT4 #(
		.INIT('h8884)
	) name6035 (
		\P1_IR_reg[12]/NET0131 ,
		\P1_state_reg[0]/NET0131 ,
		_w2010_,
		_w2011_,
		_w6498_
	);
	LUT3 #(
		.INIT('h0b)
	) name6036 (
		\P1_state_reg[0]/NET0131 ,
		_w2015_,
		_w6498_,
		_w6499_
	);
	LUT3 #(
		.INIT('h48)
	) name6037 (
		\P1_IR_reg[13]/NET0131 ,
		\P1_state_reg[0]/NET0131 ,
		_w2215_,
		_w6500_
	);
	LUT3 #(
		.INIT('h0b)
	) name6038 (
		\P1_state_reg[0]/NET0131 ,
		_w2218_,
		_w6500_,
		_w6501_
	);
	LUT4 #(
		.INIT('ha060)
	) name6039 (
		\P1_IR_reg[14]/NET0131 ,
		\P1_IR_reg[31]/NET0131 ,
		\P1_state_reg[0]/NET0131 ,
		_w480_,
		_w6502_
	);
	LUT3 #(
		.INIT('hf1)
	) name6040 (
		\P1_state_reg[0]/NET0131 ,
		_w2207_,
		_w6502_,
		_w6503_
	);
	LUT2 #(
		.INIT('h8)
	) name6041 (
		\P1_state_reg[0]/NET0131 ,
		_w2237_,
		_w6504_
	);
	LUT4 #(
		.INIT('hff54)
	) name6042 (
		\P1_state_reg[0]/NET0131 ,
		_w2239_,
		_w2241_,
		_w6504_,
		_w6505_
	);
	LUT2 #(
		.INIT('h8)
	) name6043 (
		\P1_state_reg[0]/NET0131 ,
		_w2226_,
		_w6506_
	);
	LUT4 #(
		.INIT('hff54)
	) name6044 (
		\P1_state_reg[0]/NET0131 ,
		_w2228_,
		_w2230_,
		_w6506_,
		_w6507_
	);
	LUT2 #(
		.INIT('h8)
	) name6045 (
		\P1_state_reg[0]/NET0131 ,
		_w2178_,
		_w6508_
	);
	LUT4 #(
		.INIT('h00fe)
	) name6046 (
		\P1_state_reg[0]/NET0131 ,
		_w2180_,
		_w2182_,
		_w6508_,
		_w6509_
	);
	LUT2 #(
		.INIT('h2)
	) name6047 (
		\P1_state_reg[0]/NET0131 ,
		_w2191_,
		_w6510_
	);
	LUT4 #(
		.INIT('h00fe)
	) name6048 (
		\P1_state_reg[0]/NET0131 ,
		_w2193_,
		_w2195_,
		_w6510_,
		_w6511_
	);
	LUT3 #(
		.INIT('h48)
	) name6049 (
		\P1_IR_reg[19]/NET0131 ,
		\P1_state_reg[0]/NET0131 ,
		_w2166_,
		_w6512_
	);
	LUT3 #(
		.INIT('hf1)
	) name6050 (
		\P1_state_reg[0]/NET0131 ,
		_w2170_,
		_w6512_,
		_w6513_
	);
	LUT4 #(
		.INIT('h6c00)
	) name6051 (
		\P1_IR_reg[0]/NET0131 ,
		\P1_IR_reg[1]/NET0131 ,
		\P1_IR_reg[31]/NET0131 ,
		\P1_state_reg[0]/NET0131 ,
		_w6514_
	);
	LUT3 #(
		.INIT('hf4)
	) name6052 (
		\P1_state_reg[0]/NET0131 ,
		_w2080_,
		_w6514_,
		_w6515_
	);
	LUT3 #(
		.INIT('h48)
	) name6053 (
		\P1_IR_reg[20]/NET0131 ,
		\P1_state_reg[0]/NET0131 ,
		_w2290_,
		_w6516_
	);
	LUT3 #(
		.INIT('hf1)
	) name6054 (
		\P1_state_reg[0]/NET0131 ,
		_w2154_,
		_w6516_,
		_w6517_
	);
	LUT3 #(
		.INIT('h48)
	) name6055 (
		\P1_IR_reg[21]/NET0131 ,
		\P1_state_reg[0]/NET0131 ,
		_w2287_,
		_w6518_
	);
	LUT3 #(
		.INIT('h0b)
	) name6056 (
		\P1_state_reg[0]/NET0131 ,
		_w1982_,
		_w6518_,
		_w6519_
	);
	LUT2 #(
		.INIT('h8)
	) name6057 (
		\P1_state_reg[0]/NET0131 ,
		_w2282_,
		_w6520_
	);
	LUT4 #(
		.INIT('hff54)
	) name6058 (
		\P1_state_reg[0]/NET0131 ,
		_w1966_,
		_w1970_,
		_w6520_,
		_w6521_
	);
	LUT3 #(
		.INIT('hf1)
	) name6059 (
		\P1_state_reg[0]/NET0131 ,
		_w1957_,
		_w2695_,
		_w6522_
	);
	LUT4 #(
		.INIT('ha060)
	) name6060 (
		\P1_IR_reg[24]/NET0131 ,
		\P1_IR_reg[31]/NET0131 ,
		\P1_state_reg[0]/NET0131 ,
		_w1726_,
		_w6523_
	);
	LUT4 #(
		.INIT('hff54)
	) name6061 (
		\P1_state_reg[0]/NET0131 ,
		_w1941_,
		_w1947_,
		_w6523_,
		_w6524_
	);
	LUT2 #(
		.INIT('h8)
	) name6062 (
		\P1_state_reg[0]/NET0131 ,
		_w1747_,
		_w6525_
	);
	LUT3 #(
		.INIT('hf1)
	) name6063 (
		\P1_state_reg[0]/NET0131 ,
		_w1815_,
		_w6525_,
		_w6526_
	);
	LUT4 #(
		.INIT('h4448)
	) name6064 (
		\P1_IR_reg[29]/NET0131 ,
		\P1_state_reg[0]/NET0131 ,
		_w475_,
		_w477_,
		_w6527_
	);
	LUT3 #(
		.INIT('hf1)
	) name6065 (
		\P1_state_reg[0]/NET0131 ,
		_w2272_,
		_w6527_,
		_w6528_
	);
	LUT2 #(
		.INIT('h8)
	) name6066 (
		\P1_state_reg[0]/NET0131 ,
		_w2064_,
		_w6529_
	);
	LUT3 #(
		.INIT('hf1)
	) name6067 (
		\P1_state_reg[0]/NET0131 ,
		_w2063_,
		_w6529_,
		_w6530_
	);
	LUT4 #(
		.INIT('h4448)
	) name6068 (
		\P1_IR_reg[30]/NET0131 ,
		\P1_state_reg[0]/NET0131 ,
		_w484_,
		_w487_,
		_w6531_
	);
	LUT3 #(
		.INIT('hf1)
	) name6069 (
		\P1_state_reg[0]/NET0131 ,
		_w3134_,
		_w6531_,
		_w6532_
	);
	LUT3 #(
		.INIT('h40)
	) name6070 (
		\P1_IR_reg[30]/NET0131 ,
		\P1_IR_reg[31]/NET0131 ,
		\P1_state_reg[0]/NET0131 ,
		_w6533_
	);
	LUT3 #(
		.INIT('h80)
	) name6071 (
		_w485_,
		_w1742_,
		_w6533_,
		_w6534_
	);
	LUT2 #(
		.INIT('h8)
	) name6072 (
		_w1722_,
		_w6534_,
		_w6535_
	);
	LUT3 #(
		.INIT('hf4)
	) name6073 (
		\P1_state_reg[0]/NET0131 ,
		_w3125_,
		_w6535_,
		_w6536_
	);
	LUT3 #(
		.INIT('h84)
	) name6074 (
		\P1_IR_reg[3]/NET0131 ,
		\P1_state_reg[0]/NET0131 ,
		_w2069_,
		_w6537_
	);
	LUT3 #(
		.INIT('hf1)
	) name6075 (
		\P1_state_reg[0]/NET0131 ,
		_w2068_,
		_w6537_,
		_w6538_
	);
	LUT4 #(
		.INIT('hc060)
	) name6076 (
		\P1_IR_reg[31]/NET0131 ,
		\P1_IR_reg[4]/NET0131 ,
		\P1_state_reg[0]/NET0131 ,
		_w465_,
		_w6539_
	);
	LUT3 #(
		.INIT('hf1)
	) name6077 (
		\P1_state_reg[0]/NET0131 ,
		_w2055_,
		_w6539_,
		_w6540_
	);
	LUT2 #(
		.INIT('h8)
	) name6078 (
		\P1_state_reg[0]/NET0131 ,
		_w2133_,
		_w6541_
	);
	LUT3 #(
		.INIT('hf1)
	) name6079 (
		\P1_state_reg[0]/NET0131 ,
		_w2132_,
		_w6541_,
		_w6542_
	);
	LUT3 #(
		.INIT('h48)
	) name6080 (
		\P1_IR_reg[7]/NET0131 ,
		\P1_state_reg[0]/NET0131 ,
		_w2111_,
		_w6543_
	);
	LUT3 #(
		.INIT('h0b)
	) name6081 (
		\P1_state_reg[0]/NET0131 ,
		_w2113_,
		_w6543_,
		_w6544_
	);
	LUT2 #(
		.INIT('h8)
	) name6082 (
		\P1_state_reg[0]/NET0131 ,
		_w2123_,
		_w6545_
	);
	LUT3 #(
		.INIT('hf1)
	) name6083 (
		\P1_state_reg[0]/NET0131 ,
		_w2122_,
		_w6545_,
		_w6546_
	);
	LUT3 #(
		.INIT('h84)
	) name6084 (
		\P1_IR_reg[8]/NET0131 ,
		\P1_state_reg[0]/NET0131 ,
		_w2097_,
		_w6547_
	);
	LUT4 #(
		.INIT('h00fe)
	) name6085 (
		\P1_state_reg[0]/NET0131 ,
		_w2100_,
		_w2102_,
		_w6547_,
		_w6548_
	);
	LUT4 #(
		.INIT('hc060)
	) name6086 (
		\P1_IR_reg[31]/NET0131 ,
		\P1_IR_reg[9]/NET0131 ,
		\P1_state_reg[0]/NET0131 ,
		_w467_,
		_w6549_
	);
	LUT3 #(
		.INIT('hf1)
	) name6087 (
		\P1_state_reg[0]/NET0131 ,
		_w2039_,
		_w6549_,
		_w6550_
	);
	LUT3 #(
		.INIT('h96)
	) name6088 (
		\P1_IR_reg[8]/NET0131 ,
		\P1_reg1_reg[8]/NET0131 ,
		_w2097_,
		_w6551_
	);
	LUT2 #(
		.INIT('h8)
	) name6089 (
		\P1_reg1_reg[6]/NET0131 ,
		_w2123_,
		_w6552_
	);
	LUT2 #(
		.INIT('h1)
	) name6090 (
		\P1_reg1_reg[6]/NET0131 ,
		_w2123_,
		_w6553_
	);
	LUT3 #(
		.INIT('h12)
	) name6091 (
		\P1_IR_reg[3]/NET0131 ,
		\P1_reg1_reg[3]/NET0131 ,
		_w2069_,
		_w6554_
	);
	LUT3 #(
		.INIT('h84)
	) name6092 (
		\P1_IR_reg[3]/NET0131 ,
		\P1_reg1_reg[3]/NET0131 ,
		_w2069_,
		_w6555_
	);
	LUT2 #(
		.INIT('h8)
	) name6093 (
		\P1_IR_reg[0]/NET0131 ,
		\P1_reg1_reg[0]/NET0131 ,
		_w6556_
	);
	LUT3 #(
		.INIT('he8)
	) name6094 (
		\P1_reg1_reg[1]/NET0131 ,
		_w2079_,
		_w6556_,
		_w6557_
	);
	LUT4 #(
		.INIT('h0107)
	) name6095 (
		\P1_reg1_reg[2]/NET0131 ,
		_w2064_,
		_w6555_,
		_w6557_,
		_w6558_
	);
	LUT4 #(
		.INIT('hddd4)
	) name6096 (
		\P1_reg1_reg[4]/NET0131 ,
		_w2056_,
		_w6554_,
		_w6558_,
		_w6559_
	);
	LUT4 #(
		.INIT('h080e)
	) name6097 (
		\P1_reg1_reg[5]/NET0131 ,
		_w2133_,
		_w6553_,
		_w6559_,
		_w6560_
	);
	LUT4 #(
		.INIT('h1117)
	) name6098 (
		\P1_reg1_reg[7]/NET0131 ,
		_w2112_,
		_w6552_,
		_w6560_,
		_w6561_
	);
	LUT2 #(
		.INIT('h4)
	) name6099 (
		_w1744_,
		_w1747_,
		_w6562_
	);
	LUT3 #(
		.INIT('h82)
	) name6100 (
		_w6562_,
		_w6551_,
		_w6561_,
		_w6563_
	);
	LUT3 #(
		.INIT('h48)
	) name6101 (
		\P1_IR_reg[8]/NET0131 ,
		\P1_reg2_reg[8]/NET0131 ,
		_w2097_,
		_w6564_
	);
	LUT3 #(
		.INIT('h21)
	) name6102 (
		\P1_IR_reg[8]/NET0131 ,
		\P1_reg2_reg[8]/NET0131 ,
		_w2097_,
		_w6565_
	);
	LUT3 #(
		.INIT('h96)
	) name6103 (
		\P1_IR_reg[8]/NET0131 ,
		\P1_reg2_reg[8]/NET0131 ,
		_w2097_,
		_w6566_
	);
	LUT2 #(
		.INIT('h8)
	) name6104 (
		\P1_reg2_reg[6]/NET0131 ,
		_w2123_,
		_w6567_
	);
	LUT2 #(
		.INIT('h1)
	) name6105 (
		\P1_reg2_reg[6]/NET0131 ,
		_w2123_,
		_w6568_
	);
	LUT3 #(
		.INIT('h12)
	) name6106 (
		\P1_IR_reg[3]/NET0131 ,
		\P1_reg2_reg[3]/NET0131 ,
		_w2069_,
		_w6569_
	);
	LUT3 #(
		.INIT('h84)
	) name6107 (
		\P1_IR_reg[3]/NET0131 ,
		\P1_reg2_reg[3]/NET0131 ,
		_w2069_,
		_w6570_
	);
	LUT2 #(
		.INIT('h8)
	) name6108 (
		\P1_IR_reg[0]/NET0131 ,
		\P1_reg2_reg[0]/NET0131 ,
		_w6571_
	);
	LUT3 #(
		.INIT('he8)
	) name6109 (
		\P1_reg2_reg[1]/NET0131 ,
		_w2079_,
		_w6571_,
		_w6572_
	);
	LUT4 #(
		.INIT('h0107)
	) name6110 (
		\P1_reg2_reg[2]/NET0131 ,
		_w2064_,
		_w6570_,
		_w6572_,
		_w6573_
	);
	LUT4 #(
		.INIT('hddd4)
	) name6111 (
		\P1_reg2_reg[4]/NET0131 ,
		_w2056_,
		_w6569_,
		_w6573_,
		_w6574_
	);
	LUT4 #(
		.INIT('h080e)
	) name6112 (
		\P1_reg2_reg[5]/NET0131 ,
		_w2133_,
		_w6568_,
		_w6574_,
		_w6575_
	);
	LUT4 #(
		.INIT('h1117)
	) name6113 (
		\P1_reg2_reg[7]/NET0131 ,
		_w2112_,
		_w6567_,
		_w6575_,
		_w6576_
	);
	LUT2 #(
		.INIT('h8)
	) name6114 (
		_w1744_,
		_w1747_,
		_w6577_
	);
	LUT4 #(
		.INIT('h00bf)
	) name6115 (
		_w1723_,
		_w1727_,
		_w1730_,
		_w1744_,
		_w6578_
	);
	LUT4 #(
		.INIT('h2230)
	) name6116 (
		\P1_addr_reg[8]/NET0131 ,
		_w1747_,
		_w2098_,
		_w6578_,
		_w6579_
	);
	LUT4 #(
		.INIT('h007d)
	) name6117 (
		_w6577_,
		_w6566_,
		_w6576_,
		_w6579_,
		_w6580_
	);
	LUT4 #(
		.INIT('he2ee)
	) name6118 (
		\P1_reg3_reg[8]/NET0131 ,
		\P1_state_reg[0]/NET0131 ,
		_w6563_,
		_w6580_,
		_w6581_
	);
	LUT4 #(
		.INIT('h4448)
	) name6119 (
		\P1_IR_reg[12]/NET0131 ,
		\P1_reg1_reg[12]/NET0131 ,
		_w2010_,
		_w2011_,
		_w6582_
	);
	LUT4 #(
		.INIT('h2221)
	) name6120 (
		\P1_IR_reg[12]/NET0131 ,
		\P1_reg1_reg[12]/NET0131 ,
		_w2010_,
		_w2011_,
		_w6583_
	);
	LUT4 #(
		.INIT('h9996)
	) name6121 (
		\P1_IR_reg[12]/NET0131 ,
		\P1_reg1_reg[12]/NET0131 ,
		_w2010_,
		_w2011_,
		_w6584_
	);
	LUT4 #(
		.INIT('ha060)
	) name6122 (
		\P1_IR_reg[11]/NET0131 ,
		\P1_IR_reg[31]/NET0131 ,
		\P1_reg1_reg[11]/NET0131 ,
		_w1718_,
		_w6585_
	);
	LUT3 #(
		.INIT('h48)
	) name6123 (
		\P1_IR_reg[10]/NET0131 ,
		\P1_reg1_reg[10]/NET0131 ,
		_w2010_,
		_w6586_
	);
	LUT4 #(
		.INIT('hc060)
	) name6124 (
		\P1_IR_reg[31]/NET0131 ,
		\P1_IR_reg[9]/NET0131 ,
		\P1_reg1_reg[9]/NET0131 ,
		_w467_,
		_w6587_
	);
	LUT3 #(
		.INIT('h71)
	) name6125 (
		\P1_reg1_reg[8]/NET0131 ,
		_w2098_,
		_w6561_,
		_w6588_
	);
	LUT4 #(
		.INIT('h0071)
	) name6126 (
		\P1_reg1_reg[8]/NET0131 ,
		_w2098_,
		_w6561_,
		_w6587_,
		_w6589_
	);
	LUT3 #(
		.INIT('h21)
	) name6127 (
		\P1_IR_reg[10]/NET0131 ,
		\P1_reg1_reg[10]/NET0131 ,
		_w2010_,
		_w6590_
	);
	LUT4 #(
		.INIT('h0309)
	) name6128 (
		\P1_IR_reg[31]/NET0131 ,
		\P1_IR_reg[9]/NET0131 ,
		\P1_reg1_reg[9]/NET0131 ,
		_w467_,
		_w6591_
	);
	LUT2 #(
		.INIT('h1)
	) name6129 (
		_w6590_,
		_w6591_,
		_w6592_
	);
	LUT3 #(
		.INIT('h45)
	) name6130 (
		_w6586_,
		_w6589_,
		_w6592_,
		_w6593_
	);
	LUT4 #(
		.INIT('h1011)
	) name6131 (
		_w6585_,
		_w6586_,
		_w6589_,
		_w6592_,
		_w6594_
	);
	LUT4 #(
		.INIT('h0509)
	) name6132 (
		\P1_IR_reg[11]/NET0131 ,
		\P1_IR_reg[31]/NET0131 ,
		\P1_reg1_reg[11]/NET0131 ,
		_w1718_,
		_w6595_
	);
	LUT4 #(
		.INIT('h8882)
	) name6133 (
		_w6562_,
		_w6584_,
		_w6594_,
		_w6595_,
		_w6596_
	);
	LUT4 #(
		.INIT('h2230)
	) name6134 (
		\P1_addr_reg[12]/NET0131 ,
		_w1747_,
		_w2012_,
		_w6578_,
		_w6597_
	);
	LUT4 #(
		.INIT('h4448)
	) name6135 (
		\P1_IR_reg[12]/NET0131 ,
		\P1_reg2_reg[12]/NET0131 ,
		_w2010_,
		_w2011_,
		_w6598_
	);
	LUT4 #(
		.INIT('h2221)
	) name6136 (
		\P1_IR_reg[12]/NET0131 ,
		\P1_reg2_reg[12]/NET0131 ,
		_w2010_,
		_w2011_,
		_w6599_
	);
	LUT4 #(
		.INIT('h9996)
	) name6137 (
		\P1_IR_reg[12]/NET0131 ,
		\P1_reg2_reg[12]/NET0131 ,
		_w2010_,
		_w2011_,
		_w6600_
	);
	LUT4 #(
		.INIT('h0509)
	) name6138 (
		\P1_IR_reg[11]/NET0131 ,
		\P1_IR_reg[31]/NET0131 ,
		\P1_reg2_reg[11]/NET0131 ,
		_w1718_,
		_w6601_
	);
	LUT3 #(
		.INIT('h21)
	) name6139 (
		\P1_IR_reg[10]/NET0131 ,
		\P1_reg2_reg[10]/NET0131 ,
		_w2010_,
		_w6602_
	);
	LUT4 #(
		.INIT('h0309)
	) name6140 (
		\P1_IR_reg[31]/NET0131 ,
		\P1_IR_reg[9]/NET0131 ,
		\P1_reg2_reg[9]/NET0131 ,
		_w467_,
		_w6603_
	);
	LUT2 #(
		.INIT('h1)
	) name6141 (
		_w6565_,
		_w6603_,
		_w6604_
	);
	LUT4 #(
		.INIT('hc060)
	) name6142 (
		\P1_IR_reg[31]/NET0131 ,
		\P1_IR_reg[9]/NET0131 ,
		\P1_reg2_reg[9]/NET0131 ,
		_w467_,
		_w6605_
	);
	LUT3 #(
		.INIT('h4d)
	) name6143 (
		\P1_reg2_reg[9]/NET0131 ,
		_w2038_,
		_w6564_,
		_w6606_
	);
	LUT3 #(
		.INIT('hb0)
	) name6144 (
		_w6576_,
		_w6604_,
		_w6606_,
		_w6607_
	);
	LUT4 #(
		.INIT('h1033)
	) name6145 (
		_w6576_,
		_w6602_,
		_w6604_,
		_w6606_,
		_w6608_
	);
	LUT4 #(
		.INIT('ha060)
	) name6146 (
		\P1_IR_reg[11]/NET0131 ,
		\P1_IR_reg[31]/NET0131 ,
		\P1_reg2_reg[11]/NET0131 ,
		_w1718_,
		_w6609_
	);
	LUT3 #(
		.INIT('h48)
	) name6147 (
		\P1_IR_reg[10]/NET0131 ,
		\P1_reg2_reg[10]/NET0131 ,
		_w2010_,
		_w6610_
	);
	LUT2 #(
		.INIT('h1)
	) name6148 (
		_w6609_,
		_w6610_,
		_w6611_
	);
	LUT3 #(
		.INIT('h45)
	) name6149 (
		_w6601_,
		_w6608_,
		_w6611_,
		_w6612_
	);
	LUT4 #(
		.INIT('h3113)
	) name6150 (
		_w6577_,
		_w6597_,
		_w6600_,
		_w6612_,
		_w6613_
	);
	LUT4 #(
		.INIT('he2ee)
	) name6151 (
		\P1_reg3_reg[12]/NET0131 ,
		\P1_state_reg[0]/NET0131 ,
		_w6596_,
		_w6613_,
		_w6614_
	);
	LUT4 #(
		.INIT('h3c96)
	) name6152 (
		\P1_IR_reg[31]/NET0131 ,
		\P1_IR_reg[9]/NET0131 ,
		\P1_reg2_reg[9]/NET0131 ,
		_w467_,
		_w6615_
	);
	LUT4 #(
		.INIT('h8e00)
	) name6153 (
		\P1_reg2_reg[8]/NET0131 ,
		_w2098_,
		_w6576_,
		_w6615_,
		_w6616_
	);
	LUT4 #(
		.INIT('h0071)
	) name6154 (
		\P1_reg2_reg[8]/NET0131 ,
		_w2098_,
		_w6576_,
		_w6615_,
		_w6617_
	);
	LUT3 #(
		.INIT('h02)
	) name6155 (
		_w6577_,
		_w6617_,
		_w6616_,
		_w6618_
	);
	LUT4 #(
		.INIT('h3c96)
	) name6156 (
		\P1_IR_reg[31]/NET0131 ,
		\P1_IR_reg[9]/NET0131 ,
		\P1_reg1_reg[9]/NET0131 ,
		_w467_,
		_w6619_
	);
	LUT4 #(
		.INIT('h2203)
	) name6157 (
		\P1_addr_reg[9]/NET0131 ,
		_w1747_,
		_w2038_,
		_w6578_,
		_w6620_
	);
	LUT4 #(
		.INIT('h007d)
	) name6158 (
		_w6562_,
		_w6588_,
		_w6619_,
		_w6620_,
		_w6621_
	);
	LUT4 #(
		.INIT('he2ee)
	) name6159 (
		\P1_reg3_reg[9]/NET0131 ,
		\P1_state_reg[0]/NET0131 ,
		_w6618_,
		_w6621_,
		_w6622_
	);
	LUT3 #(
		.INIT('h69)
	) name6160 (
		\P1_IR_reg[7]/NET0131 ,
		\P1_reg1_reg[7]/NET0131 ,
		_w2111_,
		_w6623_
	);
	LUT4 #(
		.INIT('h02a8)
	) name6161 (
		_w6562_,
		_w6552_,
		_w6560_,
		_w6623_,
		_w6624_
	);
	LUT4 #(
		.INIT('h2230)
	) name6162 (
		\P1_addr_reg[7]/NET0131 ,
		_w1747_,
		_w2112_,
		_w6578_,
		_w6625_
	);
	LUT3 #(
		.INIT('h69)
	) name6163 (
		\P1_IR_reg[7]/NET0131 ,
		\P1_reg2_reg[7]/NET0131 ,
		_w2111_,
		_w6626_
	);
	LUT4 #(
		.INIT('h02a8)
	) name6164 (
		_w6577_,
		_w6567_,
		_w6575_,
		_w6626_,
		_w6627_
	);
	LUT4 #(
		.INIT('haaa8)
	) name6165 (
		\P1_state_reg[0]/NET0131 ,
		_w6625_,
		_w6627_,
		_w6624_,
		_w6628_
	);
	LUT2 #(
		.INIT('he)
	) name6166 (
		_w5528_,
		_w6628_,
		_w6629_
	);
	LUT4 #(
		.INIT('ha060)
	) name6167 (
		\P1_IR_reg[14]/NET0131 ,
		\P1_IR_reg[31]/NET0131 ,
		\P1_reg1_reg[14]/NET0131 ,
		_w480_,
		_w6630_
	);
	LUT4 #(
		.INIT('h0509)
	) name6168 (
		\P1_IR_reg[14]/NET0131 ,
		\P1_IR_reg[31]/NET0131 ,
		\P1_reg1_reg[14]/NET0131 ,
		_w480_,
		_w6631_
	);
	LUT4 #(
		.INIT('h5a96)
	) name6169 (
		\P1_IR_reg[14]/NET0131 ,
		\P1_IR_reg[31]/NET0131 ,
		\P1_reg1_reg[14]/NET0131 ,
		_w480_,
		_w6632_
	);
	LUT3 #(
		.INIT('h84)
	) name6170 (
		\P1_IR_reg[13]/NET0131 ,
		\P1_reg1_reg[13]/NET0131 ,
		_w2215_,
		_w6633_
	);
	LUT3 #(
		.INIT('h12)
	) name6171 (
		\P1_IR_reg[13]/NET0131 ,
		\P1_reg1_reg[13]/NET0131 ,
		_w2215_,
		_w6634_
	);
	LUT2 #(
		.INIT('h1)
	) name6172 (
		_w6583_,
		_w6595_,
		_w6635_
	);
	LUT3 #(
		.INIT('h45)
	) name6173 (
		_w6582_,
		_w6594_,
		_w6635_,
		_w6636_
	);
	LUT4 #(
		.INIT('h0b0a)
	) name6174 (
		_w6582_,
		_w6594_,
		_w6634_,
		_w6635_,
		_w6637_
	);
	LUT4 #(
		.INIT('h2228)
	) name6175 (
		_w6562_,
		_w6632_,
		_w6633_,
		_w6637_,
		_w6638_
	);
	LUT4 #(
		.INIT('h2230)
	) name6176 (
		\P1_addr_reg[14]/NET0131 ,
		_w1747_,
		_w2205_,
		_w6578_,
		_w6639_
	);
	LUT4 #(
		.INIT('ha060)
	) name6177 (
		\P1_IR_reg[14]/NET0131 ,
		\P1_IR_reg[31]/NET0131 ,
		\P1_reg2_reg[14]/NET0131 ,
		_w480_,
		_w6640_
	);
	LUT4 #(
		.INIT('h0509)
	) name6178 (
		\P1_IR_reg[14]/NET0131 ,
		\P1_IR_reg[31]/NET0131 ,
		\P1_reg2_reg[14]/NET0131 ,
		_w480_,
		_w6641_
	);
	LUT4 #(
		.INIT('h5a96)
	) name6179 (
		\P1_IR_reg[14]/NET0131 ,
		\P1_IR_reg[31]/NET0131 ,
		\P1_reg2_reg[14]/NET0131 ,
		_w480_,
		_w6642_
	);
	LUT3 #(
		.INIT('h12)
	) name6180 (
		\P1_IR_reg[13]/NET0131 ,
		\P1_reg2_reg[13]/NET0131 ,
		_w2215_,
		_w6643_
	);
	LUT4 #(
		.INIT('h1011)
	) name6181 (
		_w6599_,
		_w6601_,
		_w6608_,
		_w6611_,
		_w6644_
	);
	LUT4 #(
		.INIT('h007b)
	) name6182 (
		\P1_IR_reg[13]/NET0131 ,
		\P1_reg2_reg[13]/NET0131 ,
		_w2215_,
		_w6598_,
		_w6645_
	);
	LUT3 #(
		.INIT('h45)
	) name6183 (
		_w6643_,
		_w6644_,
		_w6645_,
		_w6646_
	);
	LUT4 #(
		.INIT('h3113)
	) name6184 (
		_w6577_,
		_w6639_,
		_w6642_,
		_w6646_,
		_w6647_
	);
	LUT4 #(
		.INIT('he2ee)
	) name6185 (
		\P1_reg3_reg[14]/NET0131 ,
		\P1_state_reg[0]/NET0131 ,
		_w6638_,
		_w6647_,
		_w6648_
	);
	LUT3 #(
		.INIT('h12)
	) name6186 (
		\P2_IR_reg[9]/NET0131 ,
		\P2_reg1_reg[9]/NET0131 ,
		_w662_,
		_w6649_
	);
	LUT3 #(
		.INIT('h84)
	) name6187 (
		\P2_IR_reg[9]/NET0131 ,
		\P2_reg1_reg[9]/NET0131 ,
		_w662_,
		_w6650_
	);
	LUT3 #(
		.INIT('h69)
	) name6188 (
		\P2_IR_reg[9]/NET0131 ,
		\P2_reg1_reg[9]/NET0131 ,
		_w662_,
		_w6651_
	);
	LUT3 #(
		.INIT('h84)
	) name6189 (
		\P2_IR_reg[8]/NET0131 ,
		\P2_reg1_reg[8]/NET0131 ,
		_w729_,
		_w6652_
	);
	LUT3 #(
		.INIT('h12)
	) name6190 (
		\P2_IR_reg[8]/NET0131 ,
		\P2_reg1_reg[8]/NET0131 ,
		_w729_,
		_w6653_
	);
	LUT3 #(
		.INIT('h48)
	) name6191 (
		\P2_IR_reg[6]/NET0131 ,
		\P2_reg1_reg[6]/NET0131 ,
		_w750_,
		_w6654_
	);
	LUT3 #(
		.INIT('h21)
	) name6192 (
		\P2_IR_reg[6]/NET0131 ,
		\P2_reg1_reg[6]/NET0131 ,
		_w750_,
		_w6655_
	);
	LUT2 #(
		.INIT('h1)
	) name6193 (
		\P2_reg1_reg[5]/NET0131 ,
		_w773_,
		_w6656_
	);
	LUT4 #(
		.INIT('h3090)
	) name6194 (
		\P2_IR_reg[31]/NET0131 ,
		\P2_IR_reg[4]/NET0131 ,
		\P2_reg1_reg[4]/NET0131 ,
		_w496_,
		_w6657_
	);
	LUT4 #(
		.INIT('h0c06)
	) name6195 (
		\P2_IR_reg[31]/NET0131 ,
		\P2_IR_reg[4]/NET0131 ,
		\P2_reg1_reg[4]/NET0131 ,
		_w496_,
		_w6658_
	);
	LUT3 #(
		.INIT('h84)
	) name6196 (
		\P2_IR_reg[3]/NET0131 ,
		\P2_reg1_reg[3]/NET0131 ,
		_w794_,
		_w6659_
	);
	LUT3 #(
		.INIT('h12)
	) name6197 (
		\P2_IR_reg[3]/NET0131 ,
		\P2_reg1_reg[3]/NET0131 ,
		_w794_,
		_w6660_
	);
	LUT2 #(
		.INIT('h2)
	) name6198 (
		\P2_IR_reg[0]/NET0131 ,
		\P2_reg1_reg[0]/NET0131 ,
		_w6661_
	);
	LUT3 #(
		.INIT('h71)
	) name6199 (
		\P2_reg1_reg[1]/NET0131 ,
		_w816_,
		_w6661_,
		_w6662_
	);
	LUT4 #(
		.INIT('h080e)
	) name6200 (
		\P2_reg1_reg[2]/NET0131 ,
		_w806_,
		_w6660_,
		_w6662_,
		_w6663_
	);
	LUT4 #(
		.INIT('h444d)
	) name6201 (
		\P2_reg1_reg[4]/NET0131 ,
		_w784_,
		_w6659_,
		_w6663_,
		_w6664_
	);
	LUT4 #(
		.INIT('h080e)
	) name6202 (
		\P2_reg1_reg[5]/NET0131 ,
		_w773_,
		_w6655_,
		_w6664_,
		_w6665_
	);
	LUT4 #(
		.INIT('h444d)
	) name6203 (
		\P2_reg1_reg[7]/NET0131 ,
		_w762_,
		_w6654_,
		_w6665_,
		_w6666_
	);
	LUT4 #(
		.INIT('h0d04)
	) name6204 (
		\P2_reg1_reg[8]/NET0131 ,
		_w730_,
		_w6651_,
		_w6666_,
		_w6667_
	);
	LUT4 #(
		.INIT('h20b0)
	) name6205 (
		\P2_reg1_reg[8]/NET0131 ,
		_w730_,
		_w6651_,
		_w6666_,
		_w6668_
	);
	LUT3 #(
		.INIT('h02)
	) name6206 (
		_w546_,
		_w6668_,
		_w6667_,
		_w6669_
	);
	LUT3 #(
		.INIT('h84)
	) name6207 (
		\P2_IR_reg[9]/NET0131 ,
		\P2_reg2_reg[9]/NET0131 ,
		_w662_,
		_w6670_
	);
	LUT3 #(
		.INIT('h12)
	) name6208 (
		\P2_IR_reg[9]/NET0131 ,
		\P2_reg2_reg[9]/NET0131 ,
		_w662_,
		_w6671_
	);
	LUT3 #(
		.INIT('h69)
	) name6209 (
		\P2_IR_reg[9]/NET0131 ,
		\P2_reg2_reg[9]/NET0131 ,
		_w662_,
		_w6672_
	);
	LUT3 #(
		.INIT('h84)
	) name6210 (
		\P2_IR_reg[8]/NET0131 ,
		\P2_reg2_reg[8]/NET0131 ,
		_w729_,
		_w6673_
	);
	LUT3 #(
		.INIT('h12)
	) name6211 (
		\P2_IR_reg[8]/NET0131 ,
		\P2_reg2_reg[8]/NET0131 ,
		_w729_,
		_w6674_
	);
	LUT2 #(
		.INIT('h2)
	) name6212 (
		\P2_reg2_reg[7]/NET0131 ,
		_w762_,
		_w6675_
	);
	LUT2 #(
		.INIT('h4)
	) name6213 (
		\P2_reg2_reg[7]/NET0131 ,
		_w762_,
		_w6676_
	);
	LUT3 #(
		.INIT('h48)
	) name6214 (
		\P2_IR_reg[6]/NET0131 ,
		\P2_reg2_reg[6]/NET0131 ,
		_w750_,
		_w6677_
	);
	LUT3 #(
		.INIT('h21)
	) name6215 (
		\P2_IR_reg[6]/NET0131 ,
		\P2_reg2_reg[6]/NET0131 ,
		_w750_,
		_w6678_
	);
	LUT2 #(
		.INIT('h8)
	) name6216 (
		\P2_reg2_reg[5]/NET0131 ,
		_w773_,
		_w6679_
	);
	LUT2 #(
		.INIT('h1)
	) name6217 (
		\P2_reg2_reg[5]/NET0131 ,
		_w773_,
		_w6680_
	);
	LUT3 #(
		.INIT('h84)
	) name6218 (
		\P2_IR_reg[3]/NET0131 ,
		\P2_reg2_reg[3]/NET0131 ,
		_w794_,
		_w6681_
	);
	LUT3 #(
		.INIT('h12)
	) name6219 (
		\P2_IR_reg[3]/NET0131 ,
		\P2_reg2_reg[3]/NET0131 ,
		_w794_,
		_w6682_
	);
	LUT2 #(
		.INIT('h2)
	) name6220 (
		\P2_IR_reg[0]/NET0131 ,
		\P2_reg2_reg[0]/NET0131 ,
		_w6683_
	);
	LUT3 #(
		.INIT('h71)
	) name6221 (
		\P2_reg2_reg[1]/NET0131 ,
		_w816_,
		_w6683_,
		_w6684_
	);
	LUT4 #(
		.INIT('h080e)
	) name6222 (
		\P2_reg2_reg[2]/NET0131 ,
		_w806_,
		_w6682_,
		_w6684_,
		_w6685_
	);
	LUT4 #(
		.INIT('h444d)
	) name6223 (
		\P2_reg2_reg[4]/NET0131 ,
		_w784_,
		_w6681_,
		_w6685_,
		_w6686_
	);
	LUT3 #(
		.INIT('h71)
	) name6224 (
		\P2_reg2_reg[5]/NET0131 ,
		_w773_,
		_w6686_,
		_w6687_
	);
	LUT4 #(
		.INIT('h080e)
	) name6225 (
		\P2_reg2_reg[5]/NET0131 ,
		_w773_,
		_w6678_,
		_w6686_,
		_w6688_
	);
	LUT4 #(
		.INIT('h444d)
	) name6226 (
		\P2_reg2_reg[7]/NET0131 ,
		_w762_,
		_w6677_,
		_w6688_,
		_w6689_
	);
	LUT3 #(
		.INIT('hd4)
	) name6227 (
		\P2_reg2_reg[8]/NET0131 ,
		_w730_,
		_w6689_,
		_w6690_
	);
	LUT4 #(
		.INIT('h0056)
	) name6228 (
		\P2_IR_reg[28]/NET0131 ,
		_w534_,
		_w536_,
		_w717_,
		_w6691_
	);
	LUT4 #(
		.INIT('h0040)
	) name6229 (
		_w1189_,
		_w1352_,
		_w1356_,
		_w6691_,
		_w6692_
	);
	LUT4 #(
		.INIT('h7d00)
	) name6230 (
		_w1434_,
		_w6672_,
		_w6690_,
		_w6692_,
		_w6693_
	);
	LUT2 #(
		.INIT('h4)
	) name6231 (
		\P2_IR_reg[0]/NET0131 ,
		\P2_reg1_reg[0]/NET0131 ,
		_w6694_
	);
	LUT3 #(
		.INIT('he8)
	) name6232 (
		\P2_reg1_reg[1]/NET0131 ,
		_w816_,
		_w6694_,
		_w6695_
	);
	LUT4 #(
		.INIT('h0107)
	) name6233 (
		\P2_reg1_reg[2]/NET0131 ,
		_w806_,
		_w6659_,
		_w6695_,
		_w6696_
	);
	LUT3 #(
		.INIT('h07)
	) name6234 (
		\P2_reg1_reg[5]/NET0131 ,
		_w773_,
		_w6657_,
		_w6697_
	);
	LUT4 #(
		.INIT('hfe00)
	) name6235 (
		_w6658_,
		_w6660_,
		_w6696_,
		_w6697_,
		_w6698_
	);
	LUT4 #(
		.INIT('h222b)
	) name6236 (
		\P2_reg1_reg[6]/NET0131 ,
		_w751_,
		_w6656_,
		_w6698_,
		_w6699_
	);
	LUT4 #(
		.INIT('h0b02)
	) name6237 (
		\P2_reg1_reg[7]/NET0131 ,
		_w762_,
		_w6653_,
		_w6699_,
		_w6700_
	);
	LUT4 #(
		.INIT('h8882)
	) name6238 (
		_w1433_,
		_w6651_,
		_w6700_,
		_w6652_,
		_w6701_
	);
	LUT2 #(
		.INIT('h4)
	) name6239 (
		\P2_IR_reg[0]/NET0131 ,
		\P2_reg2_reg[0]/NET0131 ,
		_w6702_
	);
	LUT3 #(
		.INIT('he8)
	) name6240 (
		\P2_reg2_reg[1]/NET0131 ,
		_w816_,
		_w6702_,
		_w6703_
	);
	LUT4 #(
		.INIT('h0e08)
	) name6241 (
		\P2_reg2_reg[2]/NET0131 ,
		_w806_,
		_w6682_,
		_w6703_,
		_w6704_
	);
	LUT4 #(
		.INIT('h444d)
	) name6242 (
		\P2_reg2_reg[4]/NET0131 ,
		_w784_,
		_w6681_,
		_w6704_,
		_w6705_
	);
	LUT2 #(
		.INIT('h1)
	) name6243 (
		_w6678_,
		_w6680_,
		_w6706_
	);
	LUT4 #(
		.INIT('h1055)
	) name6244 (
		_w6677_,
		_w6679_,
		_w6705_,
		_w6706_,
		_w6707_
	);
	LUT2 #(
		.INIT('h1)
	) name6245 (
		_w6674_,
		_w6676_,
		_w6708_
	);
	LUT4 #(
		.INIT('h1055)
	) name6246 (
		_w6673_,
		_w6675_,
		_w6707_,
		_w6708_,
		_w6709_
	);
	LUT2 #(
		.INIT('h8)
	) name6247 (
		_w537_,
		_w545_,
		_w6710_
	);
	LUT3 #(
		.INIT('h02)
	) name6248 (
		\P2_addr_reg[9]/NET0131 ,
		_w537_,
		_w545_,
		_w6711_
	);
	LUT3 #(
		.INIT('h04)
	) name6249 (
		_w537_,
		_w545_,
		_w717_,
		_w6712_
	);
	LUT3 #(
		.INIT('h01)
	) name6250 (
		_w1357_,
		_w6712_,
		_w6711_,
		_w6713_
	);
	LUT4 #(
		.INIT('h9f00)
	) name6251 (
		_w6672_,
		_w6709_,
		_w6710_,
		_w6713_,
		_w6714_
	);
	LUT3 #(
		.INIT('h8a)
	) name6252 (
		\P1_state_reg[0]/NET0131 ,
		_w6701_,
		_w6714_,
		_w6715_
	);
	LUT4 #(
		.INIT('hefaa)
	) name6253 (
		_w4354_,
		_w6669_,
		_w6693_,
		_w6715_,
		_w6716_
	);
	LUT2 #(
		.INIT('h2)
	) name6254 (
		\P1_reg3_reg[0]/NET0131 ,
		\P1_state_reg[0]/NET0131 ,
		_w6717_
	);
	LUT3 #(
		.INIT('hb0)
	) name6255 (
		\P1_reg2_reg[0]/NET0131 ,
		_w1744_,
		_w1747_,
		_w6718_
	);
	LUT3 #(
		.INIT('h01)
	) name6256 (
		\P1_IR_reg[0]/NET0131 ,
		_w6578_,
		_w6718_,
		_w6719_
	);
	LUT2 #(
		.INIT('h6)
	) name6257 (
		\P1_IR_reg[0]/NET0131 ,
		\P1_reg1_reg[0]/NET0131 ,
		_w6720_
	);
	LUT4 #(
		.INIT('h80c4)
	) name6258 (
		_w1744_,
		_w1747_,
		_w6571_,
		_w6720_,
		_w6721_
	);
	LUT2 #(
		.INIT('h1)
	) name6259 (
		\P1_addr_reg[0]/NET0131 ,
		_w1747_,
		_w6722_
	);
	LUT4 #(
		.INIT('h002a)
	) name6260 (
		\P1_state_reg[0]/NET0131 ,
		_w6578_,
		_w6722_,
		_w6721_,
		_w6723_
	);
	LUT3 #(
		.INIT('hba)
	) name6261 (
		_w6717_,
		_w6719_,
		_w6723_,
		_w6724_
	);
	LUT3 #(
		.INIT('h96)
	) name6262 (
		\P1_IR_reg[10]/NET0131 ,
		\P1_reg1_reg[10]/NET0131 ,
		_w2010_,
		_w6725_
	);
	LUT4 #(
		.INIT('ha802)
	) name6263 (
		_w6562_,
		_w6589_,
		_w6591_,
		_w6725_,
		_w6726_
	);
	LUT4 #(
		.INIT('h2203)
	) name6264 (
		\P1_addr_reg[10]/NET0131 ,
		_w1747_,
		_w2023_,
		_w6578_,
		_w6727_
	);
	LUT3 #(
		.INIT('h96)
	) name6265 (
		\P1_IR_reg[10]/NET0131 ,
		\P1_reg2_reg[10]/NET0131 ,
		_w2010_,
		_w6728_
	);
	LUT4 #(
		.INIT('h070d)
	) name6266 (
		_w6577_,
		_w6607_,
		_w6727_,
		_w6728_,
		_w6729_
	);
	LUT4 #(
		.INIT('he2ee)
	) name6267 (
		\P1_reg3_reg[10]/NET0131 ,
		\P1_state_reg[0]/NET0131 ,
		_w6726_,
		_w6729_,
		_w6730_
	);
	LUT4 #(
		.INIT('h5a96)
	) name6268 (
		\P1_IR_reg[11]/NET0131 ,
		\P1_IR_reg[31]/NET0131 ,
		\P1_reg1_reg[11]/NET0131 ,
		_w1718_,
		_w6731_
	);
	LUT4 #(
		.INIT('h5a96)
	) name6269 (
		\P1_IR_reg[11]/NET0131 ,
		\P1_IR_reg[31]/NET0131 ,
		\P1_reg2_reg[11]/NET0131 ,
		_w1718_,
		_w6732_
	);
	LUT3 #(
		.INIT('h01)
	) name6270 (
		_w6565_,
		_w6602_,
		_w6603_,
		_w6733_
	);
	LUT3 #(
		.INIT('h4d)
	) name6271 (
		\P1_reg2_reg[10]/NET0131 ,
		_w2023_,
		_w6605_,
		_w6734_
	);
	LUT4 #(
		.INIT('h4f00)
	) name6272 (
		_w6564_,
		_w6576_,
		_w6733_,
		_w6734_,
		_w6735_
	);
	LUT4 #(
		.INIT('h2203)
	) name6273 (
		\P1_addr_reg[11]/NET0131 ,
		_w1747_,
		_w2001_,
		_w6578_,
		_w6736_
	);
	LUT4 #(
		.INIT('h007d)
	) name6274 (
		_w6577_,
		_w6732_,
		_w6735_,
		_w6736_,
		_w6737_
	);
	LUT4 #(
		.INIT('h7d00)
	) name6275 (
		_w6562_,
		_w6593_,
		_w6731_,
		_w6737_,
		_w6738_
	);
	LUT3 #(
		.INIT('h2e)
	) name6276 (
		\P1_reg3_reg[11]/NET0131 ,
		\P1_state_reg[0]/NET0131 ,
		_w6738_,
		_w6739_
	);
	LUT3 #(
		.INIT('h69)
	) name6277 (
		\P1_IR_reg[13]/NET0131 ,
		\P1_reg1_reg[13]/NET0131 ,
		_w2215_,
		_w6740_
	);
	LUT4 #(
		.INIT('h2230)
	) name6278 (
		\P1_addr_reg[13]/NET0131 ,
		_w1747_,
		_w2216_,
		_w6578_,
		_w6741_
	);
	LUT3 #(
		.INIT('h69)
	) name6279 (
		\P1_IR_reg[13]/NET0131 ,
		\P1_reg2_reg[13]/NET0131 ,
		_w2215_,
		_w6742_
	);
	LUT2 #(
		.INIT('h1)
	) name6280 (
		_w6599_,
		_w6601_,
		_w6743_
	);
	LUT4 #(
		.INIT('h1055)
	) name6281 (
		_w6598_,
		_w6609_,
		_w6735_,
		_w6743_,
		_w6744_
	);
	LUT4 #(
		.INIT('h1331)
	) name6282 (
		_w6577_,
		_w6741_,
		_w6742_,
		_w6744_,
		_w6745_
	);
	LUT4 #(
		.INIT('h7d00)
	) name6283 (
		_w6562_,
		_w6636_,
		_w6740_,
		_w6745_,
		_w6746_
	);
	LUT3 #(
		.INIT('h2e)
	) name6284 (
		\P1_reg3_reg[13]/NET0131 ,
		\P1_state_reg[0]/NET0131 ,
		_w6746_,
		_w6747_
	);
	LUT4 #(
		.INIT('h2228)
	) name6285 (
		\P2_IR_reg[0]/NET0131 ,
		\P2_IR_reg[28]/NET0131 ,
		_w534_,
		_w536_,
		_w6748_
	);
	LUT4 #(
		.INIT('h0040)
	) name6286 (
		_w1189_,
		_w1352_,
		_w1356_,
		_w6748_,
		_w6749_
	);
	LUT2 #(
		.INIT('h9)
	) name6287 (
		\P2_IR_reg[0]/NET0131 ,
		\P2_reg2_reg[0]/NET0131 ,
		_w6750_
	);
	LUT2 #(
		.INIT('h9)
	) name6288 (
		\P2_IR_reg[0]/NET0131 ,
		\P2_reg1_reg[0]/NET0131 ,
		_w6751_
	);
	LUT4 #(
		.INIT('hfbea)
	) name6289 (
		_w537_,
		_w545_,
		_w6750_,
		_w6751_,
		_w6752_
	);
	LUT2 #(
		.INIT('h8)
	) name6290 (
		_w6749_,
		_w6752_,
		_w6753_
	);
	LUT3 #(
		.INIT('h02)
	) name6291 (
		\P2_addr_reg[0]/NET0131 ,
		_w537_,
		_w545_,
		_w6754_
	);
	LUT3 #(
		.INIT('h02)
	) name6292 (
		_w537_,
		_w545_,
		_w6751_,
		_w6755_
	);
	LUT4 #(
		.INIT('h95ff)
	) name6293 (
		\P2_IR_reg[0]/NET0131 ,
		\P2_reg2_reg[0]/NET0131 ,
		_w537_,
		_w545_,
		_w6756_
	);
	LUT4 #(
		.INIT('h0100)
	) name6294 (
		_w1357_,
		_w6754_,
		_w6755_,
		_w6756_,
		_w6757_
	);
	LUT4 #(
		.INIT('h444e)
	) name6295 (
		\P1_state_reg[0]/NET0131 ,
		\P2_reg3_reg[0]/NET0131 ,
		_w6753_,
		_w6757_,
		_w6758_
	);
	LUT2 #(
		.INIT('h1)
	) name6296 (
		\P1_reg1_reg[15]/NET0131 ,
		_w2237_,
		_w6759_
	);
	LUT2 #(
		.INIT('h6)
	) name6297 (
		\P1_reg1_reg[15]/NET0131 ,
		_w2237_,
		_w6760_
	);
	LUT4 #(
		.INIT('h1117)
	) name6298 (
		\P1_reg1_reg[14]/NET0131 ,
		_w2205_,
		_w6633_,
		_w6637_,
		_w6761_
	);
	LUT3 #(
		.INIT('h82)
	) name6299 (
		_w6562_,
		_w6760_,
		_w6761_,
		_w6762_
	);
	LUT4 #(
		.INIT('h007b)
	) name6300 (
		\P1_IR_reg[13]/NET0131 ,
		\P1_reg2_reg[13]/NET0131 ,
		_w2215_,
		_w6640_,
		_w6763_
	);
	LUT4 #(
		.INIT('h0155)
	) name6301 (
		_w6641_,
		_w6643_,
		_w6744_,
		_w6763_,
		_w6764_
	);
	LUT2 #(
		.INIT('h1)
	) name6302 (
		\P1_reg2_reg[15]/NET0131 ,
		_w2237_,
		_w6765_
	);
	LUT4 #(
		.INIT('h9060)
	) name6303 (
		\P1_reg2_reg[15]/NET0131 ,
		_w2237_,
		_w6577_,
		_w6764_,
		_w6766_
	);
	LUT4 #(
		.INIT('h2230)
	) name6304 (
		\P1_addr_reg[15]/NET0131 ,
		_w1747_,
		_w2237_,
		_w6578_,
		_w6767_
	);
	LUT2 #(
		.INIT('h1)
	) name6305 (
		_w6766_,
		_w6767_,
		_w6768_
	);
	LUT4 #(
		.INIT('he2ee)
	) name6306 (
		\P1_reg3_reg[15]/NET0131 ,
		\P1_state_reg[0]/NET0131 ,
		_w6762_,
		_w6768_,
		_w6769_
	);
	LUT4 #(
		.INIT('h1112)
	) name6307 (
		\P2_IR_reg[12]/NET0131 ,
		\P2_reg2_reg[12]/NET0131 ,
		_w662_,
		_w663_,
		_w6770_
	);
	LUT4 #(
		.INIT('h8884)
	) name6308 (
		\P2_IR_reg[12]/NET0131 ,
		\P2_reg2_reg[12]/NET0131 ,
		_w662_,
		_w663_,
		_w6771_
	);
	LUT4 #(
		.INIT('h6669)
	) name6309 (
		\P2_IR_reg[12]/NET0131 ,
		\P2_reg2_reg[12]/NET0131 ,
		_w662_,
		_w663_,
		_w6772_
	);
	LUT3 #(
		.INIT('h84)
	) name6310 (
		\P2_IR_reg[11]/NET0131 ,
		\P2_reg2_reg[11]/NET0131 ,
		_w682_,
		_w6773_
	);
	LUT3 #(
		.INIT('h12)
	) name6311 (
		\P2_IR_reg[11]/NET0131 ,
		\P2_reg2_reg[11]/NET0131 ,
		_w682_,
		_w6774_
	);
	LUT3 #(
		.INIT('h48)
	) name6312 (
		\P2_IR_reg[10]/NET0131 ,
		\P2_reg2_reg[10]/NET0131 ,
		_w700_,
		_w6775_
	);
	LUT3 #(
		.INIT('h21)
	) name6313 (
		\P2_IR_reg[10]/NET0131 ,
		\P2_reg2_reg[10]/NET0131 ,
		_w700_,
		_w6776_
	);
	LUT4 #(
		.INIT('h0d04)
	) name6314 (
		\P2_reg2_reg[8]/NET0131 ,
		_w730_,
		_w6670_,
		_w6689_,
		_w6777_
	);
	LUT4 #(
		.INIT('hddd4)
	) name6315 (
		\P2_reg2_reg[10]/NET0131 ,
		_w701_,
		_w6671_,
		_w6777_,
		_w6778_
	);
	LUT4 #(
		.INIT('h0d04)
	) name6316 (
		\P2_reg2_reg[11]/NET0131 ,
		_w683_,
		_w6772_,
		_w6778_,
		_w6779_
	);
	LUT4 #(
		.INIT('h20b0)
	) name6317 (
		\P2_reg2_reg[11]/NET0131 ,
		_w683_,
		_w6772_,
		_w6778_,
		_w6780_
	);
	LUT3 #(
		.INIT('h02)
	) name6318 (
		_w1434_,
		_w6780_,
		_w6779_,
		_w6781_
	);
	LUT4 #(
		.INIT('h1112)
	) name6319 (
		\P2_IR_reg[12]/NET0131 ,
		\P2_reg1_reg[12]/NET0131 ,
		_w662_,
		_w663_,
		_w6782_
	);
	LUT4 #(
		.INIT('h8884)
	) name6320 (
		\P2_IR_reg[12]/NET0131 ,
		\P2_reg1_reg[12]/NET0131 ,
		_w662_,
		_w663_,
		_w6783_
	);
	LUT4 #(
		.INIT('h6669)
	) name6321 (
		\P2_IR_reg[12]/NET0131 ,
		\P2_reg1_reg[12]/NET0131 ,
		_w662_,
		_w663_,
		_w6784_
	);
	LUT3 #(
		.INIT('h84)
	) name6322 (
		\P2_IR_reg[11]/NET0131 ,
		\P2_reg1_reg[11]/NET0131 ,
		_w682_,
		_w6785_
	);
	LUT3 #(
		.INIT('h12)
	) name6323 (
		\P2_IR_reg[11]/NET0131 ,
		\P2_reg1_reg[11]/NET0131 ,
		_w682_,
		_w6786_
	);
	LUT3 #(
		.INIT('h48)
	) name6324 (
		\P2_IR_reg[10]/NET0131 ,
		\P2_reg1_reg[10]/NET0131 ,
		_w700_,
		_w6787_
	);
	LUT3 #(
		.INIT('h21)
	) name6325 (
		\P2_IR_reg[10]/NET0131 ,
		\P2_reg1_reg[10]/NET0131 ,
		_w700_,
		_w6788_
	);
	LUT4 #(
		.INIT('h0d04)
	) name6326 (
		\P2_reg1_reg[8]/NET0131 ,
		_w730_,
		_w6650_,
		_w6666_,
		_w6789_
	);
	LUT4 #(
		.INIT('hddd4)
	) name6327 (
		\P2_reg1_reg[10]/NET0131 ,
		_w701_,
		_w6649_,
		_w6789_,
		_w6790_
	);
	LUT3 #(
		.INIT('hd4)
	) name6328 (
		\P2_reg1_reg[11]/NET0131 ,
		_w683_,
		_w6790_,
		_w6791_
	);
	LUT4 #(
		.INIT('h5600)
	) name6329 (
		\P2_IR_reg[28]/NET0131 ,
		_w534_,
		_w536_,
		_w664_,
		_w6792_
	);
	LUT4 #(
		.INIT('h0040)
	) name6330 (
		_w1189_,
		_w1352_,
		_w1356_,
		_w6792_,
		_w6793_
	);
	LUT4 #(
		.INIT('h7d00)
	) name6331 (
		_w546_,
		_w6784_,
		_w6791_,
		_w6793_,
		_w6794_
	);
	LUT2 #(
		.INIT('h1)
	) name6332 (
		_w6650_,
		_w6652_,
		_w6795_
	);
	LUT3 #(
		.INIT('h45)
	) name6333 (
		_w6649_,
		_w6700_,
		_w6795_,
		_w6796_
	);
	LUT4 #(
		.INIT('h0b0a)
	) name6334 (
		_w6649_,
		_w6700_,
		_w6787_,
		_w6795_,
		_w6797_
	);
	LUT4 #(
		.INIT('h222b)
	) name6335 (
		\P2_reg1_reg[11]/NET0131 ,
		_w683_,
		_w6788_,
		_w6797_,
		_w6798_
	);
	LUT3 #(
		.INIT('h82)
	) name6336 (
		_w1433_,
		_w6784_,
		_w6798_,
		_w6799_
	);
	LUT4 #(
		.INIT('h0701)
	) name6337 (
		\P2_reg2_reg[5]/NET0131 ,
		_w773_,
		_w6677_,
		_w6705_,
		_w6800_
	);
	LUT2 #(
		.INIT('h1)
	) name6338 (
		_w6678_,
		_w6676_,
		_w6801_
	);
	LUT3 #(
		.INIT('h45)
	) name6339 (
		_w6675_,
		_w6800_,
		_w6801_,
		_w6802_
	);
	LUT4 #(
		.INIT('h1011)
	) name6340 (
		_w6673_,
		_w6675_,
		_w6800_,
		_w6801_,
		_w6803_
	);
	LUT2 #(
		.INIT('h1)
	) name6341 (
		_w6671_,
		_w6674_,
		_w6804_
	);
	LUT4 #(
		.INIT('h1011)
	) name6342 (
		_w6670_,
		_w6775_,
		_w6803_,
		_w6804_,
		_w6805_
	);
	LUT2 #(
		.INIT('h1)
	) name6343 (
		_w6774_,
		_w6776_,
		_w6806_
	);
	LUT3 #(
		.INIT('h45)
	) name6344 (
		_w6773_,
		_w6805_,
		_w6806_,
		_w6807_
	);
	LUT3 #(
		.INIT('h02)
	) name6345 (
		\P2_addr_reg[12]/NET0131 ,
		_w537_,
		_w545_,
		_w6808_
	);
	LUT3 #(
		.INIT('h40)
	) name6346 (
		_w537_,
		_w545_,
		_w664_,
		_w6809_
	);
	LUT3 #(
		.INIT('h01)
	) name6347 (
		_w1357_,
		_w6809_,
		_w6808_,
		_w6810_
	);
	LUT4 #(
		.INIT('hd700)
	) name6348 (
		_w6710_,
		_w6772_,
		_w6807_,
		_w6810_,
		_w6811_
	);
	LUT3 #(
		.INIT('h8a)
	) name6349 (
		\P1_state_reg[0]/NET0131 ,
		_w6799_,
		_w6811_,
		_w6812_
	);
	LUT4 #(
		.INIT('hefaa)
	) name6350 (
		_w4292_,
		_w6781_,
		_w6794_,
		_w6812_,
		_w6813_
	);
	LUT2 #(
		.INIT('h1)
	) name6351 (
		\P1_reg1_reg[16]/NET0131 ,
		_w2226_,
		_w6814_
	);
	LUT2 #(
		.INIT('h6)
	) name6352 (
		\P1_reg1_reg[16]/NET0131 ,
		_w2226_,
		_w6815_
	);
	LUT3 #(
		.INIT('h07)
	) name6353 (
		\P1_reg1_reg[15]/NET0131 ,
		_w2237_,
		_w6630_,
		_w6816_
	);
	LUT4 #(
		.INIT('hab00)
	) name6354 (
		_w6631_,
		_w6633_,
		_w6637_,
		_w6816_,
		_w6817_
	);
	LUT4 #(
		.INIT('ha082)
	) name6355 (
		_w6562_,
		_w6759_,
		_w6815_,
		_w6817_,
		_w6818_
	);
	LUT4 #(
		.INIT('h2230)
	) name6356 (
		\P1_addr_reg[16]/NET0131 ,
		_w1747_,
		_w2226_,
		_w6578_,
		_w6819_
	);
	LUT2 #(
		.INIT('h1)
	) name6357 (
		\P1_reg2_reg[16]/NET0131 ,
		_w2226_,
		_w6820_
	);
	LUT2 #(
		.INIT('h6)
	) name6358 (
		\P1_reg2_reg[16]/NET0131 ,
		_w2226_,
		_w6821_
	);
	LUT4 #(
		.INIT('h1011)
	) name6359 (
		_w6641_,
		_w6643_,
		_w6644_,
		_w6645_,
		_w6822_
	);
	LUT3 #(
		.INIT('h07)
	) name6360 (
		\P1_reg2_reg[15]/NET0131 ,
		_w2237_,
		_w6640_,
		_w6823_
	);
	LUT3 #(
		.INIT('h45)
	) name6361 (
		_w6765_,
		_w6822_,
		_w6823_,
		_w6824_
	);
	LUT4 #(
		.INIT('h3113)
	) name6362 (
		_w6577_,
		_w6819_,
		_w6821_,
		_w6824_,
		_w6825_
	);
	LUT4 #(
		.INIT('he2ee)
	) name6363 (
		\P1_reg3_reg[16]/NET0131 ,
		\P1_state_reg[0]/NET0131 ,
		_w6818_,
		_w6825_,
		_w6826_
	);
	LUT4 #(
		.INIT('h0a06)
	) name6364 (
		\P2_IR_reg[13]/NET0131 ,
		\P2_IR_reg[31]/NET0131 ,
		\P2_reg1_reg[13]/NET0131 ,
		_w498_,
		_w6827_
	);
	LUT4 #(
		.INIT('h5090)
	) name6365 (
		\P2_IR_reg[13]/NET0131 ,
		\P2_IR_reg[31]/NET0131 ,
		\P2_reg1_reg[13]/NET0131 ,
		_w498_,
		_w6828_
	);
	LUT4 #(
		.INIT('ha569)
	) name6366 (
		\P2_IR_reg[13]/NET0131 ,
		\P2_IR_reg[31]/NET0131 ,
		\P2_reg1_reg[13]/NET0131 ,
		_w498_,
		_w6829_
	);
	LUT2 #(
		.INIT('h1)
	) name6367 (
		_w6783_,
		_w6785_,
		_w6830_
	);
	LUT4 #(
		.INIT('h0155)
	) name6368 (
		_w6782_,
		_w6786_,
		_w6790_,
		_w6830_,
		_w6831_
	);
	LUT3 #(
		.INIT('h28)
	) name6369 (
		_w546_,
		_w6829_,
		_w6831_,
		_w6832_
	);
	LUT4 #(
		.INIT('h0a06)
	) name6370 (
		\P2_IR_reg[13]/NET0131 ,
		\P2_IR_reg[31]/NET0131 ,
		\P2_reg2_reg[13]/NET0131 ,
		_w498_,
		_w6833_
	);
	LUT4 #(
		.INIT('h5090)
	) name6371 (
		\P2_IR_reg[13]/NET0131 ,
		\P2_IR_reg[31]/NET0131 ,
		\P2_reg2_reg[13]/NET0131 ,
		_w498_,
		_w6834_
	);
	LUT4 #(
		.INIT('ha569)
	) name6372 (
		\P2_IR_reg[13]/NET0131 ,
		\P2_IR_reg[31]/NET0131 ,
		\P2_reg2_reg[13]/NET0131 ,
		_w498_,
		_w6835_
	);
	LUT2 #(
		.INIT('h1)
	) name6373 (
		_w6770_,
		_w6774_,
		_w6836_
	);
	LUT3 #(
		.INIT('h4d)
	) name6374 (
		\P2_reg2_reg[12]/NET0131 ,
		_w664_,
		_w6773_,
		_w6837_
	);
	LUT3 #(
		.INIT('hb0)
	) name6375 (
		_w6778_,
		_w6836_,
		_w6837_,
		_w6838_
	);
	LUT4 #(
		.INIT('h5600)
	) name6376 (
		\P2_IR_reg[28]/NET0131 ,
		_w534_,
		_w536_,
		_w643_,
		_w6839_
	);
	LUT4 #(
		.INIT('h0040)
	) name6377 (
		_w1189_,
		_w1352_,
		_w1356_,
		_w6839_,
		_w6840_
	);
	LUT4 #(
		.INIT('h7d00)
	) name6378 (
		_w1434_,
		_w6835_,
		_w6838_,
		_w6840_,
		_w6841_
	);
	LUT2 #(
		.INIT('h1)
	) name6379 (
		_w6782_,
		_w6786_,
		_w6842_
	);
	LUT4 #(
		.INIT('hab00)
	) name6380 (
		_w6785_,
		_w6788_,
		_w6797_,
		_w6842_,
		_w6843_
	);
	LUT4 #(
		.INIT('ha082)
	) name6381 (
		_w1433_,
		_w6783_,
		_w6829_,
		_w6843_,
		_w6844_
	);
	LUT2 #(
		.INIT('h1)
	) name6382 (
		_w6671_,
		_w6776_,
		_w6845_
	);
	LUT4 #(
		.INIT('h040f)
	) name6383 (
		_w6670_,
		_w6709_,
		_w6775_,
		_w6845_,
		_w6846_
	);
	LUT4 #(
		.INIT('h1505)
	) name6384 (
		_w6771_,
		_w6773_,
		_w6836_,
		_w6846_,
		_w6847_
	);
	LUT3 #(
		.INIT('h40)
	) name6385 (
		_w537_,
		_w545_,
		_w643_,
		_w6848_
	);
	LUT3 #(
		.INIT('h02)
	) name6386 (
		\P2_addr_reg[13]/NET0131 ,
		_w537_,
		_w545_,
		_w6849_
	);
	LUT3 #(
		.INIT('h01)
	) name6387 (
		_w1357_,
		_w6849_,
		_w6848_,
		_w6850_
	);
	LUT4 #(
		.INIT('hd700)
	) name6388 (
		_w6710_,
		_w6835_,
		_w6847_,
		_w6850_,
		_w6851_
	);
	LUT3 #(
		.INIT('h8a)
	) name6389 (
		\P1_state_reg[0]/NET0131 ,
		_w6844_,
		_w6851_,
		_w6852_
	);
	LUT4 #(
		.INIT('hefaa)
	) name6390 (
		_w4313_,
		_w6832_,
		_w6841_,
		_w6852_,
		_w6853_
	);
	LUT2 #(
		.INIT('h4)
	) name6391 (
		\P1_reg1_reg[17]/NET0131 ,
		_w2178_,
		_w6854_
	);
	LUT2 #(
		.INIT('h2)
	) name6392 (
		\P1_reg1_reg[17]/NET0131 ,
		_w2178_,
		_w6855_
	);
	LUT2 #(
		.INIT('h9)
	) name6393 (
		\P1_reg1_reg[17]/NET0131 ,
		_w2178_,
		_w6856_
	);
	LUT4 #(
		.INIT('h007b)
	) name6394 (
		\P1_IR_reg[13]/NET0131 ,
		\P1_reg1_reg[13]/NET0131 ,
		_w2215_,
		_w6630_,
		_w6857_
	);
	LUT3 #(
		.INIT('h0e)
	) name6395 (
		\P1_reg1_reg[15]/NET0131 ,
		_w2237_,
		_w6631_,
		_w6858_
	);
	LUT4 #(
		.INIT('h153f)
	) name6396 (
		\P1_reg1_reg[15]/NET0131 ,
		\P1_reg1_reg[16]/NET0131 ,
		_w2226_,
		_w2237_,
		_w6859_
	);
	LUT4 #(
		.INIT('h4f00)
	) name6397 (
		_w6637_,
		_w6857_,
		_w6858_,
		_w6859_,
		_w6860_
	);
	LUT4 #(
		.INIT('ha082)
	) name6398 (
		_w6562_,
		_w6814_,
		_w6856_,
		_w6860_,
		_w6861_
	);
	LUT2 #(
		.INIT('h4)
	) name6399 (
		\P1_reg2_reg[17]/NET0131 ,
		_w2178_,
		_w6862_
	);
	LUT2 #(
		.INIT('h2)
	) name6400 (
		\P1_reg2_reg[17]/NET0131 ,
		_w2178_,
		_w6863_
	);
	LUT2 #(
		.INIT('h9)
	) name6401 (
		\P1_reg2_reg[17]/NET0131 ,
		_w2178_,
		_w6864_
	);
	LUT4 #(
		.INIT('h153f)
	) name6402 (
		\P1_reg2_reg[15]/NET0131 ,
		\P1_reg2_reg[16]/NET0131 ,
		_w2226_,
		_w2237_,
		_w6865_
	);
	LUT4 #(
		.INIT('h020f)
	) name6403 (
		_w6764_,
		_w6765_,
		_w6820_,
		_w6865_,
		_w6866_
	);
	LUT4 #(
		.INIT('h2203)
	) name6404 (
		\P1_addr_reg[17]/NET0131 ,
		_w1747_,
		_w2178_,
		_w6578_,
		_w6867_
	);
	LUT4 #(
		.INIT('h00d7)
	) name6405 (
		_w6577_,
		_w6864_,
		_w6866_,
		_w6867_,
		_w6868_
	);
	LUT4 #(
		.INIT('he2ee)
	) name6406 (
		\P1_reg3_reg[17]/NET0131 ,
		\P1_state_reg[0]/NET0131 ,
		_w6861_,
		_w6868_,
		_w6869_
	);
	LUT4 #(
		.INIT('h0a06)
	) name6407 (
		\P2_IR_reg[15]/NET0131 ,
		\P2_IR_reg[31]/NET0131 ,
		\P2_reg1_reg[15]/NET0131 ,
		_w540_,
		_w6870_
	);
	LUT4 #(
		.INIT('h5090)
	) name6408 (
		\P2_IR_reg[15]/NET0131 ,
		\P2_IR_reg[31]/NET0131 ,
		\P2_reg1_reg[15]/NET0131 ,
		_w540_,
		_w6871_
	);
	LUT4 #(
		.INIT('ha569)
	) name6409 (
		\P2_IR_reg[15]/NET0131 ,
		\P2_IR_reg[31]/NET0131 ,
		\P2_reg1_reg[15]/NET0131 ,
		_w540_,
		_w6872_
	);
	LUT2 #(
		.INIT('h4)
	) name6410 (
		\P2_reg1_reg[14]/NET0131 ,
		_w613_,
		_w6873_
	);
	LUT3 #(
		.INIT('h0b)
	) name6411 (
		\P2_reg1_reg[14]/NET0131 ,
		_w613_,
		_w6827_,
		_w6874_
	);
	LUT2 #(
		.INIT('h2)
	) name6412 (
		\P2_reg1_reg[14]/NET0131 ,
		_w613_,
		_w6875_
	);
	LUT3 #(
		.INIT('h4d)
	) name6413 (
		\P2_reg1_reg[14]/NET0131 ,
		_w613_,
		_w6828_,
		_w6876_
	);
	LUT4 #(
		.INIT('h80cc)
	) name6414 (
		_w6831_,
		_w6872_,
		_w6874_,
		_w6876_,
		_w6877_
	);
	LUT4 #(
		.INIT('h1300)
	) name6415 (
		_w6831_,
		_w6872_,
		_w6874_,
		_w6876_,
		_w6878_
	);
	LUT3 #(
		.INIT('h02)
	) name6416 (
		_w546_,
		_w6878_,
		_w6877_,
		_w6879_
	);
	LUT4 #(
		.INIT('h0a06)
	) name6417 (
		\P2_IR_reg[15]/NET0131 ,
		\P2_IR_reg[31]/NET0131 ,
		\P2_reg2_reg[15]/NET0131 ,
		_w540_,
		_w6880_
	);
	LUT4 #(
		.INIT('h5090)
	) name6418 (
		\P2_IR_reg[15]/NET0131 ,
		\P2_IR_reg[31]/NET0131 ,
		\P2_reg2_reg[15]/NET0131 ,
		_w540_,
		_w6881_
	);
	LUT4 #(
		.INIT('ha569)
	) name6419 (
		\P2_IR_reg[15]/NET0131 ,
		\P2_IR_reg[31]/NET0131 ,
		\P2_reg2_reg[15]/NET0131 ,
		_w540_,
		_w6882_
	);
	LUT2 #(
		.INIT('h4)
	) name6420 (
		\P2_reg2_reg[14]/NET0131 ,
		_w613_,
		_w6883_
	);
	LUT3 #(
		.INIT('h0b)
	) name6421 (
		\P2_reg2_reg[14]/NET0131 ,
		_w613_,
		_w6833_,
		_w6884_
	);
	LUT4 #(
		.INIT('h4f00)
	) name6422 (
		_w6778_,
		_w6836_,
		_w6837_,
		_w6884_,
		_w6885_
	);
	LUT2 #(
		.INIT('h2)
	) name6423 (
		\P2_reg2_reg[14]/NET0131 ,
		_w613_,
		_w6886_
	);
	LUT3 #(
		.INIT('h4d)
	) name6424 (
		\P2_reg2_reg[14]/NET0131 ,
		_w613_,
		_w6834_,
		_w6887_
	);
	LUT4 #(
		.INIT('h2822)
	) name6425 (
		_w1434_,
		_w6882_,
		_w6885_,
		_w6887_,
		_w6888_
	);
	LUT4 #(
		.INIT('h5600)
	) name6426 (
		\P2_IR_reg[28]/NET0131 ,
		_w534_,
		_w536_,
		_w592_,
		_w6889_
	);
	LUT4 #(
		.INIT('h0040)
	) name6427 (
		_w1189_,
		_w1352_,
		_w1356_,
		_w6889_,
		_w6890_
	);
	LUT2 #(
		.INIT('h4)
	) name6428 (
		_w6888_,
		_w6890_,
		_w6891_
	);
	LUT4 #(
		.INIT('hfe00)
	) name6429 (
		_w6783_,
		_w6828_,
		_w6843_,
		_w6874_,
		_w6892_
	);
	LUT4 #(
		.INIT('h8882)
	) name6430 (
		_w1433_,
		_w6872_,
		_w6875_,
		_w6892_,
		_w6893_
	);
	LUT4 #(
		.INIT('h040f)
	) name6431 (
		_w6834_,
		_w6847_,
		_w6886_,
		_w6884_,
		_w6894_
	);
	LUT3 #(
		.INIT('h40)
	) name6432 (
		_w537_,
		_w545_,
		_w592_,
		_w6895_
	);
	LUT3 #(
		.INIT('h02)
	) name6433 (
		\P2_addr_reg[15]/NET0131 ,
		_w537_,
		_w545_,
		_w6896_
	);
	LUT3 #(
		.INIT('h01)
	) name6434 (
		_w1357_,
		_w6896_,
		_w6895_,
		_w6897_
	);
	LUT4 #(
		.INIT('hd700)
	) name6435 (
		_w6710_,
		_w6882_,
		_w6894_,
		_w6897_,
		_w6898_
	);
	LUT3 #(
		.INIT('h8a)
	) name6436 (
		\P1_state_reg[0]/NET0131 ,
		_w6893_,
		_w6898_,
		_w6899_
	);
	LUT4 #(
		.INIT('hefaa)
	) name6437 (
		_w4648_,
		_w6879_,
		_w6891_,
		_w6899_,
		_w6900_
	);
	LUT2 #(
		.INIT('h2)
	) name6438 (
		\P2_reg2_reg[16]/NET0131 ,
		_w877_,
		_w6901_
	);
	LUT2 #(
		.INIT('h9)
	) name6439 (
		\P2_reg2_reg[16]/NET0131 ,
		_w877_,
		_w6902_
	);
	LUT3 #(
		.INIT('h0d)
	) name6440 (
		\P2_reg2_reg[14]/NET0131 ,
		_w613_,
		_w6881_,
		_w6903_
	);
	LUT4 #(
		.INIT('h020b)
	) name6441 (
		\P2_reg2_reg[11]/NET0131 ,
		_w683_,
		_w6770_,
		_w6778_,
		_w6904_
	);
	LUT2 #(
		.INIT('h1)
	) name6442 (
		_w6771_,
		_w6834_,
		_w6905_
	);
	LUT4 #(
		.INIT('h1011)
	) name6443 (
		_w6833_,
		_w6883_,
		_w6904_,
		_w6905_,
		_w6906_
	);
	LUT4 #(
		.INIT('h4404)
	) name6444 (
		_w6880_,
		_w6902_,
		_w6903_,
		_w6906_,
		_w6907_
	);
	LUT4 #(
		.INIT('h2232)
	) name6445 (
		_w6880_,
		_w6902_,
		_w6903_,
		_w6906_,
		_w6908_
	);
	LUT3 #(
		.INIT('h02)
	) name6446 (
		_w1434_,
		_w6908_,
		_w6907_,
		_w6909_
	);
	LUT2 #(
		.INIT('h2)
	) name6447 (
		\P2_reg1_reg[16]/NET0131 ,
		_w877_,
		_w6910_
	);
	LUT2 #(
		.INIT('h9)
	) name6448 (
		\P2_reg1_reg[16]/NET0131 ,
		_w877_,
		_w6911_
	);
	LUT3 #(
		.INIT('h0d)
	) name6449 (
		\P2_reg1_reg[14]/NET0131 ,
		_w613_,
		_w6871_,
		_w6912_
	);
	LUT4 #(
		.INIT('h020b)
	) name6450 (
		\P2_reg1_reg[11]/NET0131 ,
		_w683_,
		_w6782_,
		_w6790_,
		_w6913_
	);
	LUT2 #(
		.INIT('h1)
	) name6451 (
		_w6783_,
		_w6828_,
		_w6914_
	);
	LUT3 #(
		.INIT('h45)
	) name6452 (
		_w6827_,
		_w6913_,
		_w6914_,
		_w6915_
	);
	LUT4 #(
		.INIT('h1011)
	) name6453 (
		_w6827_,
		_w6873_,
		_w6913_,
		_w6914_,
		_w6916_
	);
	LUT3 #(
		.INIT('h51)
	) name6454 (
		_w6870_,
		_w6912_,
		_w6916_,
		_w6917_
	);
	LUT4 #(
		.INIT('h5600)
	) name6455 (
		\P2_IR_reg[28]/NET0131 ,
		_w534_,
		_w536_,
		_w877_,
		_w6918_
	);
	LUT4 #(
		.INIT('h0040)
	) name6456 (
		_w1189_,
		_w1352_,
		_w1356_,
		_w6918_,
		_w6919_
	);
	LUT4 #(
		.INIT('hd700)
	) name6457 (
		_w546_,
		_w6911_,
		_w6917_,
		_w6919_,
		_w6920_
	);
	LUT3 #(
		.INIT('h0b)
	) name6458 (
		\P2_reg1_reg[14]/NET0131 ,
		_w613_,
		_w6870_,
		_w6921_
	);
	LUT2 #(
		.INIT('h1)
	) name6459 (
		_w6782_,
		_w6827_,
		_w6922_
	);
	LUT4 #(
		.INIT('h010f)
	) name6460 (
		_w6783_,
		_w6798_,
		_w6828_,
		_w6922_,
		_w6923_
	);
	LUT4 #(
		.INIT('h1505)
	) name6461 (
		_w6871_,
		_w6875_,
		_w6921_,
		_w6923_,
		_w6924_
	);
	LUT3 #(
		.INIT('h28)
	) name6462 (
		_w1433_,
		_w6911_,
		_w6924_,
		_w6925_
	);
	LUT3 #(
		.INIT('h0b)
	) name6463 (
		\P2_reg2_reg[14]/NET0131 ,
		_w613_,
		_w6880_,
		_w6926_
	);
	LUT4 #(
		.INIT('h1011)
	) name6464 (
		_w6771_,
		_w6773_,
		_w6805_,
		_w6806_,
		_w6927_
	);
	LUT2 #(
		.INIT('h1)
	) name6465 (
		_w6770_,
		_w6833_,
		_w6928_
	);
	LUT3 #(
		.INIT('h45)
	) name6466 (
		_w6834_,
		_w6927_,
		_w6928_,
		_w6929_
	);
	LUT4 #(
		.INIT('h1011)
	) name6467 (
		_w6834_,
		_w6886_,
		_w6927_,
		_w6928_,
		_w6930_
	);
	LUT3 #(
		.INIT('h51)
	) name6468 (
		_w6881_,
		_w6926_,
		_w6930_,
		_w6931_
	);
	LUT3 #(
		.INIT('h40)
	) name6469 (
		_w537_,
		_w545_,
		_w877_,
		_w6932_
	);
	LUT3 #(
		.INIT('h02)
	) name6470 (
		\P2_addr_reg[16]/NET0131 ,
		_w537_,
		_w545_,
		_w6933_
	);
	LUT3 #(
		.INIT('h01)
	) name6471 (
		_w1357_,
		_w6933_,
		_w6932_,
		_w6934_
	);
	LUT4 #(
		.INIT('hd700)
	) name6472 (
		_w6710_,
		_w6902_,
		_w6931_,
		_w6934_,
		_w6935_
	);
	LUT3 #(
		.INIT('h8a)
	) name6473 (
		\P1_state_reg[0]/NET0131 ,
		_w6925_,
		_w6935_,
		_w6936_
	);
	LUT4 #(
		.INIT('hefaa)
	) name6474 (
		_w3546_,
		_w6909_,
		_w6920_,
		_w6936_,
		_w6937_
	);
	LUT2 #(
		.INIT('h4)
	) name6475 (
		\P2_reg1_reg[17]/NET0131 ,
		_w858_,
		_w6938_
	);
	LUT2 #(
		.INIT('h2)
	) name6476 (
		\P2_reg1_reg[17]/NET0131 ,
		_w858_,
		_w6939_
	);
	LUT2 #(
		.INIT('h9)
	) name6477 (
		\P2_reg1_reg[17]/NET0131 ,
		_w858_,
		_w6940_
	);
	LUT3 #(
		.INIT('h0b)
	) name6478 (
		\P2_reg1_reg[16]/NET0131 ,
		_w877_,
		_w6870_,
		_w6941_
	);
	LUT4 #(
		.INIT('h010f)
	) name6479 (
		_w6828_,
		_w6831_,
		_w6875_,
		_w6874_,
		_w6942_
	);
	LUT3 #(
		.INIT('h4d)
	) name6480 (
		\P2_reg1_reg[16]/NET0131 ,
		_w877_,
		_w6871_,
		_w6943_
	);
	LUT4 #(
		.INIT('h08aa)
	) name6481 (
		_w6940_,
		_w6941_,
		_w6942_,
		_w6943_,
		_w6944_
	);
	LUT4 #(
		.INIT('h5100)
	) name6482 (
		_w6940_,
		_w6941_,
		_w6942_,
		_w6943_,
		_w6945_
	);
	LUT3 #(
		.INIT('h02)
	) name6483 (
		_w546_,
		_w6945_,
		_w6944_,
		_w6946_
	);
	LUT2 #(
		.INIT('h4)
	) name6484 (
		\P2_reg2_reg[17]/NET0131 ,
		_w858_,
		_w6947_
	);
	LUT2 #(
		.INIT('h2)
	) name6485 (
		\P2_reg2_reg[17]/NET0131 ,
		_w858_,
		_w6948_
	);
	LUT2 #(
		.INIT('h9)
	) name6486 (
		\P2_reg2_reg[17]/NET0131 ,
		_w858_,
		_w6949_
	);
	LUT3 #(
		.INIT('h0b)
	) name6487 (
		\P2_reg2_reg[16]/NET0131 ,
		_w877_,
		_w6880_,
		_w6950_
	);
	LUT4 #(
		.INIT('h2300)
	) name6488 (
		_w6778_,
		_w6834_,
		_w6836_,
		_w6837_,
		_w6951_
	);
	LUT4 #(
		.INIT('ha0e0)
	) name6489 (
		_w6886_,
		_w6884_,
		_w6950_,
		_w6951_,
		_w6952_
	);
	LUT3 #(
		.INIT('h4d)
	) name6490 (
		\P2_reg2_reg[16]/NET0131 ,
		_w877_,
		_w6881_,
		_w6953_
	);
	LUT4 #(
		.INIT('h2822)
	) name6491 (
		_w1434_,
		_w6949_,
		_w6952_,
		_w6953_,
		_w6954_
	);
	LUT4 #(
		.INIT('h5600)
	) name6492 (
		\P2_IR_reg[28]/NET0131 ,
		_w534_,
		_w536_,
		_w858_,
		_w6955_
	);
	LUT4 #(
		.INIT('h0040)
	) name6493 (
		_w1189_,
		_w1352_,
		_w1356_,
		_w6955_,
		_w6956_
	);
	LUT2 #(
		.INIT('h4)
	) name6494 (
		_w6954_,
		_w6956_,
		_w6957_
	);
	LUT4 #(
		.INIT('hfe00)
	) name6495 (
		_w6871_,
		_w6875_,
		_w6892_,
		_w6941_,
		_w6958_
	);
	LUT4 #(
		.INIT('ha082)
	) name6496 (
		_w1433_,
		_w6910_,
		_w6940_,
		_w6958_,
		_w6959_
	);
	LUT4 #(
		.INIT('h040f)
	) name6497 (
		_w6881_,
		_w6894_,
		_w6901_,
		_w6950_,
		_w6960_
	);
	LUT3 #(
		.INIT('h40)
	) name6498 (
		_w537_,
		_w545_,
		_w858_,
		_w6961_
	);
	LUT3 #(
		.INIT('h02)
	) name6499 (
		\P2_addr_reg[17]/NET0131 ,
		_w537_,
		_w545_,
		_w6962_
	);
	LUT3 #(
		.INIT('h01)
	) name6500 (
		_w1357_,
		_w6962_,
		_w6961_,
		_w6963_
	);
	LUT4 #(
		.INIT('hd700)
	) name6501 (
		_w6710_,
		_w6949_,
		_w6960_,
		_w6963_,
		_w6964_
	);
	LUT3 #(
		.INIT('h8a)
	) name6502 (
		\P1_state_reg[0]/NET0131 ,
		_w6959_,
		_w6964_,
		_w6965_
	);
	LUT4 #(
		.INIT('hefaa)
	) name6503 (
		_w2609_,
		_w6946_,
		_w6957_,
		_w6965_,
		_w6966_
	);
	LUT3 #(
		.INIT('h21)
	) name6504 (
		\P2_IR_reg[18]/NET0131 ,
		\P2_reg1_reg[18]/NET0131 ,
		_w922_,
		_w6967_
	);
	LUT3 #(
		.INIT('h48)
	) name6505 (
		\P2_IR_reg[18]/NET0131 ,
		\P2_reg1_reg[18]/NET0131 ,
		_w922_,
		_w6968_
	);
	LUT3 #(
		.INIT('h96)
	) name6506 (
		\P2_IR_reg[18]/NET0131 ,
		\P2_reg1_reg[18]/NET0131 ,
		_w922_,
		_w6969_
	);
	LUT4 #(
		.INIT('h8acf)
	) name6507 (
		\P2_reg1_reg[16]/NET0131 ,
		\P2_reg1_reg[17]/NET0131 ,
		_w858_,
		_w877_,
		_w6970_
	);
	LUT4 #(
		.INIT('h040f)
	) name6508 (
		_w6910_,
		_w6924_,
		_w6939_,
		_w6970_,
		_w6971_
	);
	LUT3 #(
		.INIT('h28)
	) name6509 (
		_w1433_,
		_w6969_,
		_w6971_,
		_w6972_
	);
	LUT3 #(
		.INIT('h21)
	) name6510 (
		\P2_IR_reg[18]/NET0131 ,
		\P2_reg2_reg[18]/NET0131 ,
		_w922_,
		_w6973_
	);
	LUT3 #(
		.INIT('h48)
	) name6511 (
		\P2_IR_reg[18]/NET0131 ,
		\P2_reg2_reg[18]/NET0131 ,
		_w922_,
		_w6974_
	);
	LUT3 #(
		.INIT('h96)
	) name6512 (
		\P2_IR_reg[18]/NET0131 ,
		\P2_reg2_reg[18]/NET0131 ,
		_w922_,
		_w6975_
	);
	LUT4 #(
		.INIT('h8acf)
	) name6513 (
		\P2_reg2_reg[16]/NET0131 ,
		\P2_reg2_reg[17]/NET0131 ,
		_w858_,
		_w877_,
		_w6976_
	);
	LUT4 #(
		.INIT('h1101)
	) name6514 (
		_w6881_,
		_w6901_,
		_w6926_,
		_w6930_,
		_w6977_
	);
	LUT3 #(
		.INIT('h51)
	) name6515 (
		_w6948_,
		_w6976_,
		_w6977_,
		_w6978_
	);
	LUT3 #(
		.INIT('h02)
	) name6516 (
		\P2_addr_reg[18]/NET0131 ,
		_w537_,
		_w545_,
		_w6979_
	);
	LUT3 #(
		.INIT('h40)
	) name6517 (
		_w537_,
		_w545_,
		_w923_,
		_w6980_
	);
	LUT3 #(
		.INIT('h01)
	) name6518 (
		_w1357_,
		_w6980_,
		_w6979_,
		_w6981_
	);
	LUT4 #(
		.INIT('hd700)
	) name6519 (
		_w6710_,
		_w6975_,
		_w6978_,
		_w6981_,
		_w6982_
	);
	LUT4 #(
		.INIT('hf351)
	) name6520 (
		\P2_reg2_reg[16]/NET0131 ,
		\P2_reg2_reg[17]/NET0131 ,
		_w858_,
		_w877_,
		_w6983_
	);
	LUT4 #(
		.INIT('h1033)
	) name6521 (
		_w6903_,
		_w6947_,
		_w6950_,
		_w6983_,
		_w6984_
	);
	LUT2 #(
		.INIT('h8)
	) name6522 (
		_w6926_,
		_w6976_,
		_w6985_
	);
	LUT4 #(
		.INIT('h4500)
	) name6523 (
		_w6833_,
		_w6904_,
		_w6905_,
		_w6985_,
		_w6986_
	);
	LUT4 #(
		.INIT('h2228)
	) name6524 (
		_w1434_,
		_w6975_,
		_w6984_,
		_w6986_,
		_w6987_
	);
	LUT4 #(
		.INIT('hf351)
	) name6525 (
		\P2_reg1_reg[16]/NET0131 ,
		\P2_reg1_reg[17]/NET0131 ,
		_w858_,
		_w877_,
		_w6988_
	);
	LUT4 #(
		.INIT('h1033)
	) name6526 (
		_w6912_,
		_w6938_,
		_w6941_,
		_w6988_,
		_w6989_
	);
	LUT2 #(
		.INIT('h8)
	) name6527 (
		_w6921_,
		_w6970_,
		_w6990_
	);
	LUT4 #(
		.INIT('h4500)
	) name6528 (
		_w6827_,
		_w6913_,
		_w6914_,
		_w6990_,
		_w6991_
	);
	LUT4 #(
		.INIT('h2228)
	) name6529 (
		_w546_,
		_w6969_,
		_w6989_,
		_w6991_,
		_w6992_
	);
	LUT2 #(
		.INIT('h8)
	) name6530 (
		_w537_,
		_w923_,
		_w6993_
	);
	LUT2 #(
		.INIT('h2)
	) name6531 (
		_w1357_,
		_w6993_,
		_w6994_
	);
	LUT4 #(
		.INIT('ha8aa)
	) name6532 (
		\P1_state_reg[0]/NET0131 ,
		_w6992_,
		_w6987_,
		_w6994_,
		_w6995_
	);
	LUT4 #(
		.INIT('hefaa)
	) name6533 (
		_w2568_,
		_w6972_,
		_w6982_,
		_w6995_,
		_w6996_
	);
	LUT3 #(
		.INIT('h96)
	) name6534 (
		\P2_IR_reg[6]/NET0131 ,
		\P2_reg1_reg[6]/NET0131 ,
		_w750_,
		_w6997_
	);
	LUT4 #(
		.INIT('h0071)
	) name6535 (
		\P2_reg1_reg[5]/NET0131 ,
		_w773_,
		_w6664_,
		_w6997_,
		_w6998_
	);
	LUT4 #(
		.INIT('h8e00)
	) name6536 (
		\P2_reg1_reg[5]/NET0131 ,
		_w773_,
		_w6664_,
		_w6997_,
		_w6999_
	);
	LUT3 #(
		.INIT('h02)
	) name6537 (
		_w546_,
		_w6999_,
		_w6998_,
		_w7000_
	);
	LUT3 #(
		.INIT('h96)
	) name6538 (
		\P2_IR_reg[6]/NET0131 ,
		\P2_reg2_reg[6]/NET0131 ,
		_w750_,
		_w7001_
	);
	LUT4 #(
		.INIT('h5600)
	) name6539 (
		\P2_IR_reg[28]/NET0131 ,
		_w534_,
		_w536_,
		_w751_,
		_w7002_
	);
	LUT4 #(
		.INIT('h0040)
	) name6540 (
		_w1189_,
		_w1352_,
		_w1356_,
		_w7002_,
		_w7003_
	);
	LUT4 #(
		.INIT('h7d00)
	) name6541 (
		_w1434_,
		_w6687_,
		_w7001_,
		_w7003_,
		_w7004_
	);
	LUT2 #(
		.INIT('h4)
	) name6542 (
		_w7000_,
		_w7004_,
		_w7005_
	);
	LUT4 #(
		.INIT('h7100)
	) name6543 (
		\P2_reg2_reg[5]/NET0131 ,
		_w773_,
		_w6705_,
		_w7001_,
		_w7006_
	);
	LUT4 #(
		.INIT('h008e)
	) name6544 (
		\P2_reg2_reg[5]/NET0131 ,
		_w773_,
		_w6705_,
		_w7001_,
		_w7007_
	);
	LUT3 #(
		.INIT('h02)
	) name6545 (
		_w6710_,
		_w7007_,
		_w7006_,
		_w7008_
	);
	LUT3 #(
		.INIT('he0)
	) name6546 (
		_w6656_,
		_w6698_,
		_w6997_,
		_w7009_
	);
	LUT3 #(
		.INIT('h01)
	) name6547 (
		_w6656_,
		_w6698_,
		_w6997_,
		_w7010_
	);
	LUT3 #(
		.INIT('h02)
	) name6548 (
		_w1433_,
		_w7010_,
		_w7009_,
		_w7011_
	);
	LUT3 #(
		.INIT('h02)
	) name6549 (
		\P2_addr_reg[6]/NET0131 ,
		_w537_,
		_w545_,
		_w7012_
	);
	LUT3 #(
		.INIT('h40)
	) name6550 (
		_w537_,
		_w545_,
		_w751_,
		_w7013_
	);
	LUT3 #(
		.INIT('h01)
	) name6551 (
		_w1357_,
		_w7013_,
		_w7012_,
		_w7014_
	);
	LUT4 #(
		.INIT('ha8aa)
	) name6552 (
		\P1_state_reg[0]/NET0131 ,
		_w7011_,
		_w7008_,
		_w7014_,
		_w7015_
	);
	LUT3 #(
		.INIT('hba)
	) name6553 (
		_w5191_,
		_w7005_,
		_w7015_,
		_w7016_
	);
	LUT4 #(
		.INIT('h936c)
	) name6554 (
		\P1_IR_reg[0]/NET0131 ,
		\P1_IR_reg[1]/NET0131 ,
		\P1_IR_reg[31]/NET0131 ,
		\P1_reg2_reg[1]/NET0131 ,
		_w7017_
	);
	LUT2 #(
		.INIT('h6)
	) name6555 (
		_w6571_,
		_w7017_,
		_w7018_
	);
	LUT4 #(
		.INIT('h936c)
	) name6556 (
		\P1_IR_reg[0]/NET0131 ,
		\P1_IR_reg[1]/NET0131 ,
		\P1_IR_reg[31]/NET0131 ,
		\P1_reg1_reg[1]/NET0131 ,
		_w7019_
	);
	LUT2 #(
		.INIT('h9)
	) name6557 (
		_w6556_,
		_w7019_,
		_w7020_
	);
	LUT4 #(
		.INIT('h40c8)
	) name6558 (
		_w1744_,
		_w1747_,
		_w7020_,
		_w7018_,
		_w7021_
	);
	LUT4 #(
		.INIT('h1103)
	) name6559 (
		\P1_addr_reg[1]/NET0131 ,
		_w1747_,
		_w2079_,
		_w6578_,
		_w7022_
	);
	LUT4 #(
		.INIT('h222e)
	) name6560 (
		\P1_reg3_reg[1]/NET0131 ,
		\P1_state_reg[0]/NET0131 ,
		_w7021_,
		_w7022_,
		_w7023_
	);
	LUT2 #(
		.INIT('h6)
	) name6561 (
		\P1_reg2_reg[2]/NET0131 ,
		_w2064_,
		_w7024_
	);
	LUT2 #(
		.INIT('h6)
	) name6562 (
		_w6572_,
		_w7024_,
		_w7025_
	);
	LUT2 #(
		.INIT('h6)
	) name6563 (
		\P1_reg1_reg[2]/NET0131 ,
		_w2064_,
		_w7026_
	);
	LUT2 #(
		.INIT('h9)
	) name6564 (
		_w6557_,
		_w7026_,
		_w7027_
	);
	LUT4 #(
		.INIT('h40c8)
	) name6565 (
		_w1744_,
		_w1747_,
		_w7027_,
		_w7025_,
		_w7028_
	);
	LUT4 #(
		.INIT('h1103)
	) name6566 (
		\P1_addr_reg[2]/NET0131 ,
		_w1747_,
		_w2064_,
		_w6578_,
		_w7029_
	);
	LUT4 #(
		.INIT('h222e)
	) name6567 (
		\P1_reg3_reg[2]/NET0131 ,
		\P1_state_reg[0]/NET0131 ,
		_w7028_,
		_w7029_,
		_w7030_
	);
	LUT4 #(
		.INIT('h2230)
	) name6568 (
		\P1_addr_reg[3]/NET0131 ,
		_w1747_,
		_w2070_,
		_w6578_,
		_w7031_
	);
	LUT3 #(
		.INIT('h69)
	) name6569 (
		\P1_IR_reg[3]/NET0131 ,
		\P1_reg1_reg[3]/NET0131 ,
		_w2069_,
		_w7032_
	);
	LUT4 #(
		.INIT('h17e8)
	) name6570 (
		\P1_reg1_reg[2]/NET0131 ,
		_w2064_,
		_w6557_,
		_w7032_,
		_w7033_
	);
	LUT3 #(
		.INIT('h69)
	) name6571 (
		\P1_IR_reg[3]/NET0131 ,
		\P1_reg2_reg[3]/NET0131 ,
		_w2069_,
		_w7034_
	);
	LUT4 #(
		.INIT('h17e8)
	) name6572 (
		\P1_reg2_reg[2]/NET0131 ,
		_w2064_,
		_w6572_,
		_w7034_,
		_w7035_
	);
	LUT4 #(
		.INIT('h37bf)
	) name6573 (
		_w1744_,
		_w1747_,
		_w7033_,
		_w7035_,
		_w7036_
	);
	LUT4 #(
		.INIT('he2ee)
	) name6574 (
		\P1_reg3_reg[3]/NET0131 ,
		\P1_state_reg[0]/NET0131 ,
		_w7031_,
		_w7036_,
		_w7037_
	);
	LUT4 #(
		.INIT('h2203)
	) name6575 (
		\P1_addr_reg[4]/NET0131 ,
		_w1747_,
		_w2056_,
		_w6578_,
		_w7038_
	);
	LUT4 #(
		.INIT('h3c96)
	) name6576 (
		\P1_IR_reg[31]/NET0131 ,
		\P1_IR_reg[4]/NET0131 ,
		\P1_reg1_reg[4]/NET0131 ,
		_w465_,
		_w7039_
	);
	LUT3 #(
		.INIT('he1)
	) name6577 (
		_w6554_,
		_w6558_,
		_w7039_,
		_w7040_
	);
	LUT4 #(
		.INIT('h3c96)
	) name6578 (
		\P1_IR_reg[31]/NET0131 ,
		\P1_IR_reg[4]/NET0131 ,
		\P1_reg2_reg[4]/NET0131 ,
		_w465_,
		_w7041_
	);
	LUT3 #(
		.INIT('he1)
	) name6579 (
		_w6569_,
		_w6573_,
		_w7041_,
		_w7042_
	);
	LUT4 #(
		.INIT('h37bf)
	) name6580 (
		_w1744_,
		_w1747_,
		_w7040_,
		_w7042_,
		_w7043_
	);
	LUT4 #(
		.INIT('he2ee)
	) name6581 (
		\P1_reg3_reg[4]/NET0131 ,
		\P1_state_reg[0]/NET0131 ,
		_w7038_,
		_w7043_,
		_w7044_
	);
	LUT4 #(
		.INIT('h2230)
	) name6582 (
		\P1_addr_reg[5]/NET0131 ,
		_w1747_,
		_w2133_,
		_w6578_,
		_w7045_
	);
	LUT2 #(
		.INIT('h6)
	) name6583 (
		\P1_reg2_reg[5]/NET0131 ,
		_w2133_,
		_w7046_
	);
	LUT4 #(
		.INIT('h8008)
	) name6584 (
		_w1744_,
		_w1747_,
		_w6574_,
		_w7046_,
		_w7047_
	);
	LUT2 #(
		.INIT('h6)
	) name6585 (
		\P1_reg1_reg[5]/NET0131 ,
		_w2133_,
		_w7048_
	);
	LUT4 #(
		.INIT('h4004)
	) name6586 (
		_w1744_,
		_w1747_,
		_w6559_,
		_w7048_,
		_w7049_
	);
	LUT2 #(
		.INIT('h1)
	) name6587 (
		_w7047_,
		_w7049_,
		_w7050_
	);
	LUT4 #(
		.INIT('he2ee)
	) name6588 (
		\P1_reg3_reg[5]/NET0131 ,
		\P1_state_reg[0]/NET0131 ,
		_w7045_,
		_w7050_,
		_w7051_
	);
	LUT2 #(
		.INIT('h6)
	) name6589 (
		\P1_reg2_reg[6]/NET0131 ,
		_w2123_,
		_w7052_
	);
	LUT4 #(
		.INIT('h8e00)
	) name6590 (
		\P1_reg2_reg[5]/NET0131 ,
		_w2133_,
		_w6574_,
		_w7052_,
		_w7053_
	);
	LUT4 #(
		.INIT('h0071)
	) name6591 (
		\P1_reg2_reg[5]/NET0131 ,
		_w2133_,
		_w6574_,
		_w7052_,
		_w7054_
	);
	LUT3 #(
		.INIT('h02)
	) name6592 (
		_w6577_,
		_w7054_,
		_w7053_,
		_w7055_
	);
	LUT4 #(
		.INIT('h2230)
	) name6593 (
		\P1_addr_reg[6]/NET0131 ,
		_w1747_,
		_w2123_,
		_w6578_,
		_w7056_
	);
	LUT2 #(
		.INIT('h6)
	) name6594 (
		\P1_reg1_reg[6]/NET0131 ,
		_w2123_,
		_w7057_
	);
	LUT4 #(
		.INIT('h8e00)
	) name6595 (
		\P1_reg1_reg[5]/NET0131 ,
		_w2133_,
		_w6559_,
		_w7057_,
		_w7058_
	);
	LUT4 #(
		.INIT('h0071)
	) name6596 (
		\P1_reg1_reg[5]/NET0131 ,
		_w2133_,
		_w6559_,
		_w7057_,
		_w7059_
	);
	LUT3 #(
		.INIT('h02)
	) name6597 (
		_w6562_,
		_w7059_,
		_w7058_,
		_w7060_
	);
	LUT4 #(
		.INIT('haaa8)
	) name6598 (
		\P1_state_reg[0]/NET0131 ,
		_w7056_,
		_w7060_,
		_w7055_,
		_w7061_
	);
	LUT2 #(
		.INIT('he)
	) name6599 (
		_w5509_,
		_w7061_,
		_w7062_
	);
	LUT3 #(
		.INIT('h96)
	) name6600 (
		\P2_IR_reg[10]/NET0131 ,
		\P2_reg1_reg[10]/NET0131 ,
		_w700_,
		_w7063_
	);
	LUT4 #(
		.INIT('ha802)
	) name6601 (
		_w546_,
		_w6649_,
		_w6789_,
		_w7063_,
		_w7064_
	);
	LUT3 #(
		.INIT('h96)
	) name6602 (
		\P2_IR_reg[10]/NET0131 ,
		\P2_reg2_reg[10]/NET0131 ,
		_w700_,
		_w7065_
	);
	LUT4 #(
		.INIT('ha802)
	) name6603 (
		_w1434_,
		_w6671_,
		_w6777_,
		_w7065_,
		_w7066_
	);
	LUT4 #(
		.INIT('h5600)
	) name6604 (
		\P2_IR_reg[28]/NET0131 ,
		_w534_,
		_w536_,
		_w701_,
		_w7067_
	);
	LUT4 #(
		.INIT('h0040)
	) name6605 (
		_w1189_,
		_w1352_,
		_w1356_,
		_w7067_,
		_w7068_
	);
	LUT3 #(
		.INIT('h10)
	) name6606 (
		_w7066_,
		_w7064_,
		_w7068_,
		_w7069_
	);
	LUT4 #(
		.INIT('h4500)
	) name6607 (
		_w6670_,
		_w6803_,
		_w6804_,
		_w7065_,
		_w7070_
	);
	LUT4 #(
		.INIT('h00ba)
	) name6608 (
		_w6670_,
		_w6803_,
		_w6804_,
		_w7065_,
		_w7071_
	);
	LUT3 #(
		.INIT('h02)
	) name6609 (
		_w6710_,
		_w7071_,
		_w7070_,
		_w7072_
	);
	LUT3 #(
		.INIT('h02)
	) name6610 (
		\P2_addr_reg[10]/NET0131 ,
		_w537_,
		_w545_,
		_w7073_
	);
	LUT3 #(
		.INIT('h40)
	) name6611 (
		_w537_,
		_w545_,
		_w701_,
		_w7074_
	);
	LUT3 #(
		.INIT('h01)
	) name6612 (
		_w1357_,
		_w7074_,
		_w7073_,
		_w7075_
	);
	LUT4 #(
		.INIT('h7d00)
	) name6613 (
		_w1433_,
		_w6796_,
		_w7063_,
		_w7075_,
		_w7076_
	);
	LUT3 #(
		.INIT('h8a)
	) name6614 (
		\P1_state_reg[0]/NET0131 ,
		_w7072_,
		_w7076_,
		_w7077_
	);
	LUT3 #(
		.INIT('hba)
	) name6615 (
		_w4272_,
		_w7069_,
		_w7077_,
		_w7078_
	);
	LUT3 #(
		.INIT('h69)
	) name6616 (
		\P2_IR_reg[11]/NET0131 ,
		\P2_reg2_reg[11]/NET0131 ,
		_w682_,
		_w7079_
	);
	LUT3 #(
		.INIT('h82)
	) name6617 (
		_w1434_,
		_w6778_,
		_w7079_,
		_w7080_
	);
	LUT3 #(
		.INIT('h69)
	) name6618 (
		\P2_IR_reg[11]/NET0131 ,
		\P2_reg1_reg[11]/NET0131 ,
		_w682_,
		_w7081_
	);
	LUT4 #(
		.INIT('h5600)
	) name6619 (
		\P2_IR_reg[28]/NET0131 ,
		_w534_,
		_w536_,
		_w683_,
		_w7082_
	);
	LUT4 #(
		.INIT('h0040)
	) name6620 (
		_w1189_,
		_w1352_,
		_w1356_,
		_w7082_,
		_w7083_
	);
	LUT4 #(
		.INIT('h7d00)
	) name6621 (
		_w546_,
		_w6790_,
		_w7081_,
		_w7083_,
		_w7084_
	);
	LUT4 #(
		.INIT('h02a8)
	) name6622 (
		_w1433_,
		_w6788_,
		_w6797_,
		_w7081_,
		_w7085_
	);
	LUT3 #(
		.INIT('h02)
	) name6623 (
		\P2_addr_reg[11]/NET0131 ,
		_w537_,
		_w545_,
		_w7086_
	);
	LUT3 #(
		.INIT('h40)
	) name6624 (
		_w537_,
		_w545_,
		_w683_,
		_w7087_
	);
	LUT3 #(
		.INIT('h01)
	) name6625 (
		_w1357_,
		_w7087_,
		_w7086_,
		_w7088_
	);
	LUT4 #(
		.INIT('hd700)
	) name6626 (
		_w6710_,
		_w6846_,
		_w7079_,
		_w7088_,
		_w7089_
	);
	LUT3 #(
		.INIT('h8a)
	) name6627 (
		\P1_state_reg[0]/NET0131 ,
		_w7085_,
		_w7089_,
		_w7090_
	);
	LUT4 #(
		.INIT('hefaa)
	) name6628 (
		_w4605_,
		_w7080_,
		_w7084_,
		_w7090_,
		_w7091_
	);
	LUT2 #(
		.INIT('h9)
	) name6629 (
		\P2_reg2_reg[14]/NET0131 ,
		_w613_,
		_w7092_
	);
	LUT4 #(
		.INIT('h00ba)
	) name6630 (
		_w6833_,
		_w6904_,
		_w6905_,
		_w7092_,
		_w7093_
	);
	LUT4 #(
		.INIT('h4500)
	) name6631 (
		_w6833_,
		_w6904_,
		_w6905_,
		_w7092_,
		_w7094_
	);
	LUT3 #(
		.INIT('h02)
	) name6632 (
		_w1434_,
		_w7094_,
		_w7093_,
		_w7095_
	);
	LUT2 #(
		.INIT('h9)
	) name6633 (
		\P2_reg1_reg[14]/NET0131 ,
		_w613_,
		_w7096_
	);
	LUT4 #(
		.INIT('h5600)
	) name6634 (
		\P2_IR_reg[28]/NET0131 ,
		_w534_,
		_w536_,
		_w613_,
		_w7097_
	);
	LUT4 #(
		.INIT('h0040)
	) name6635 (
		_w1189_,
		_w1352_,
		_w1356_,
		_w7097_,
		_w7098_
	);
	LUT4 #(
		.INIT('hd700)
	) name6636 (
		_w546_,
		_w6915_,
		_w7096_,
		_w7098_,
		_w7099_
	);
	LUT3 #(
		.INIT('h28)
	) name6637 (
		_w1433_,
		_w6923_,
		_w7096_,
		_w7100_
	);
	LUT3 #(
		.INIT('h40)
	) name6638 (
		_w537_,
		_w545_,
		_w613_,
		_w7101_
	);
	LUT3 #(
		.INIT('h02)
	) name6639 (
		\P2_addr_reg[14]/NET0131 ,
		_w537_,
		_w545_,
		_w7102_
	);
	LUT3 #(
		.INIT('h01)
	) name6640 (
		_w1357_,
		_w7102_,
		_w7101_,
		_w7103_
	);
	LUT4 #(
		.INIT('hd700)
	) name6641 (
		_w6710_,
		_w6929_,
		_w7092_,
		_w7103_,
		_w7104_
	);
	LUT3 #(
		.INIT('h8a)
	) name6642 (
		\P1_state_reg[0]/NET0131 ,
		_w7100_,
		_w7104_,
		_w7105_
	);
	LUT4 #(
		.INIT('hefaa)
	) name6643 (
		_w4626_,
		_w7095_,
		_w7099_,
		_w7105_,
		_w7106_
	);
	LUT2 #(
		.INIT('h6)
	) name6644 (
		\P2_reg2_reg[5]/NET0131 ,
		_w773_,
		_w7107_
	);
	LUT4 #(
		.INIT('h0880)
	) name6645 (
		_w537_,
		_w545_,
		_w6705_,
		_w7107_,
		_w7108_
	);
	LUT2 #(
		.INIT('h6)
	) name6646 (
		\P2_reg1_reg[5]/NET0131 ,
		_w773_,
		_w7109_
	);
	LUT4 #(
		.INIT('hddd4)
	) name6647 (
		\P2_reg1_reg[4]/NET0131 ,
		_w784_,
		_w6660_,
		_w6696_,
		_w7110_
	);
	LUT4 #(
		.INIT('h0220)
	) name6648 (
		_w537_,
		_w545_,
		_w7109_,
		_w7110_,
		_w7111_
	);
	LUT3 #(
		.INIT('h04)
	) name6649 (
		_w537_,
		_w545_,
		_w773_,
		_w7112_
	);
	LUT3 #(
		.INIT('h02)
	) name6650 (
		\P2_addr_reg[5]/NET0131 ,
		_w537_,
		_w545_,
		_w7113_
	);
	LUT4 #(
		.INIT('h0001)
	) name6651 (
		_w1357_,
		_w7113_,
		_w7112_,
		_w7111_,
		_w7114_
	);
	LUT4 #(
		.INIT('h1001)
	) name6652 (
		_w537_,
		_w545_,
		_w6664_,
		_w7109_,
		_w7115_
	);
	LUT4 #(
		.INIT('h4004)
	) name6653 (
		_w537_,
		_w545_,
		_w6686_,
		_w7107_,
		_w7116_
	);
	LUT4 #(
		.INIT('h0056)
	) name6654 (
		\P2_IR_reg[28]/NET0131 ,
		_w534_,
		_w536_,
		_w773_,
		_w7117_
	);
	LUT4 #(
		.INIT('h0040)
	) name6655 (
		_w1189_,
		_w1352_,
		_w1356_,
		_w7117_,
		_w7118_
	);
	LUT4 #(
		.INIT('ha8aa)
	) name6656 (
		\P1_state_reg[0]/NET0131 ,
		_w7116_,
		_w7115_,
		_w7118_,
		_w7119_
	);
	LUT4 #(
		.INIT('hefaa)
	) name6657 (
		_w5169_,
		_w7108_,
		_w7114_,
		_w7119_,
		_w7120_
	);
	LUT2 #(
		.INIT('h9)
	) name6658 (
		\P2_reg1_reg[7]/NET0131 ,
		_w762_,
		_w7121_
	);
	LUT4 #(
		.INIT('h02a8)
	) name6659 (
		_w546_,
		_w6654_,
		_w6665_,
		_w7121_,
		_w7122_
	);
	LUT2 #(
		.INIT('h9)
	) name6660 (
		\P2_reg2_reg[7]/NET0131 ,
		_w762_,
		_w7123_
	);
	LUT4 #(
		.INIT('h02a8)
	) name6661 (
		_w1434_,
		_w6677_,
		_w6688_,
		_w7123_,
		_w7124_
	);
	LUT4 #(
		.INIT('h5600)
	) name6662 (
		\P2_IR_reg[28]/NET0131 ,
		_w534_,
		_w536_,
		_w762_,
		_w7125_
	);
	LUT4 #(
		.INIT('h0040)
	) name6663 (
		_w1189_,
		_w1352_,
		_w1356_,
		_w7125_,
		_w7126_
	);
	LUT3 #(
		.INIT('h10)
	) name6664 (
		_w7124_,
		_w7122_,
		_w7126_,
		_w7127_
	);
	LUT3 #(
		.INIT('h48)
	) name6665 (
		_w6707_,
		_w6710_,
		_w7123_,
		_w7128_
	);
	LUT3 #(
		.INIT('h82)
	) name6666 (
		_w1433_,
		_w6699_,
		_w7121_,
		_w7129_
	);
	LUT3 #(
		.INIT('h40)
	) name6667 (
		_w537_,
		_w545_,
		_w762_,
		_w7130_
	);
	LUT3 #(
		.INIT('h02)
	) name6668 (
		\P2_addr_reg[7]/NET0131 ,
		_w537_,
		_w545_,
		_w7131_
	);
	LUT3 #(
		.INIT('h01)
	) name6669 (
		_w1357_,
		_w7131_,
		_w7130_,
		_w7132_
	);
	LUT4 #(
		.INIT('ha8aa)
	) name6670 (
		\P1_state_reg[0]/NET0131 ,
		_w7129_,
		_w7128_,
		_w7132_,
		_w7133_
	);
	LUT3 #(
		.INIT('hba)
	) name6671 (
		_w5212_,
		_w7127_,
		_w7133_,
		_w7134_
	);
	LUT3 #(
		.INIT('h69)
	) name6672 (
		\P2_IR_reg[8]/NET0131 ,
		\P2_reg2_reg[8]/NET0131 ,
		_w729_,
		_w7135_
	);
	LUT3 #(
		.INIT('h82)
	) name6673 (
		_w1434_,
		_w6689_,
		_w7135_,
		_w7136_
	);
	LUT3 #(
		.INIT('h69)
	) name6674 (
		\P2_IR_reg[8]/NET0131 ,
		\P2_reg1_reg[8]/NET0131 ,
		_w729_,
		_w7137_
	);
	LUT4 #(
		.INIT('h8448)
	) name6675 (
		\P2_reg1_reg[8]/NET0131 ,
		_w546_,
		_w730_,
		_w6666_,
		_w7138_
	);
	LUT4 #(
		.INIT('h5600)
	) name6676 (
		\P2_IR_reg[28]/NET0131 ,
		_w534_,
		_w536_,
		_w730_,
		_w7139_
	);
	LUT4 #(
		.INIT('h0040)
	) name6677 (
		_w1189_,
		_w1352_,
		_w1356_,
		_w7139_,
		_w7140_
	);
	LUT3 #(
		.INIT('h10)
	) name6678 (
		_w7138_,
		_w7136_,
		_w7140_,
		_w7141_
	);
	LUT4 #(
		.INIT('h4d00)
	) name6679 (
		\P2_reg1_reg[7]/NET0131 ,
		_w762_,
		_w6699_,
		_w7137_,
		_w7142_
	);
	LUT4 #(
		.INIT('h00b2)
	) name6680 (
		\P2_reg1_reg[7]/NET0131 ,
		_w762_,
		_w6699_,
		_w7137_,
		_w7143_
	);
	LUT3 #(
		.INIT('h02)
	) name6681 (
		_w1433_,
		_w7143_,
		_w7142_,
		_w7144_
	);
	LUT3 #(
		.INIT('h02)
	) name6682 (
		\P2_addr_reg[8]/NET0131 ,
		_w537_,
		_w545_,
		_w7145_
	);
	LUT3 #(
		.INIT('h40)
	) name6683 (
		_w537_,
		_w545_,
		_w730_,
		_w7146_
	);
	LUT3 #(
		.INIT('h01)
	) name6684 (
		_w1357_,
		_w7146_,
		_w7145_,
		_w7147_
	);
	LUT4 #(
		.INIT('hd700)
	) name6685 (
		_w6710_,
		_w6802_,
		_w7135_,
		_w7147_,
		_w7148_
	);
	LUT3 #(
		.INIT('h8a)
	) name6686 (
		\P1_state_reg[0]/NET0131 ,
		_w7144_,
		_w7148_,
		_w7149_
	);
	LUT3 #(
		.INIT('hba)
	) name6687 (
		_w4683_,
		_w7141_,
		_w7149_,
		_w7150_
	);
	LUT2 #(
		.INIT('h1)
	) name6688 (
		_w6938_,
		_w6967_,
		_w7151_
	);
	LUT4 #(
		.INIT('hfe00)
	) name6689 (
		_w6910_,
		_w6939_,
		_w6958_,
		_w7151_,
		_w7152_
	);
	LUT2 #(
		.INIT('h6)
	) name6690 (
		\P2_reg1_reg[19]/NET0131 ,
		_w900_,
		_w7153_
	);
	LUT4 #(
		.INIT('ha802)
	) name6691 (
		_w1433_,
		_w6968_,
		_w7152_,
		_w7153_,
		_w7154_
	);
	LUT2 #(
		.INIT('h1)
	) name6692 (
		_w6947_,
		_w6973_,
		_w7155_
	);
	LUT4 #(
		.INIT('h040f)
	) name6693 (
		_w6948_,
		_w6960_,
		_w6974_,
		_w7155_,
		_w7156_
	);
	LUT2 #(
		.INIT('h6)
	) name6694 (
		\P2_reg2_reg[19]/NET0131 ,
		_w900_,
		_w7157_
	);
	LUT3 #(
		.INIT('h02)
	) name6695 (
		\P2_addr_reg[19]/NET0131 ,
		_w537_,
		_w545_,
		_w7158_
	);
	LUT3 #(
		.INIT('h04)
	) name6696 (
		_w537_,
		_w545_,
		_w900_,
		_w7159_
	);
	LUT3 #(
		.INIT('h01)
	) name6697 (
		_w1357_,
		_w7159_,
		_w7158_,
		_w7160_
	);
	LUT4 #(
		.INIT('hd700)
	) name6698 (
		_w6710_,
		_w7156_,
		_w7157_,
		_w7160_,
		_w7161_
	);
	LUT2 #(
		.INIT('h4)
	) name6699 (
		_w7154_,
		_w7161_,
		_w7162_
	);
	LUT4 #(
		.INIT('h8f00)
	) name6700 (
		_w6831_,
		_w6874_,
		_w6876_,
		_w6941_,
		_w7163_
	);
	LUT2 #(
		.INIT('h4)
	) name6701 (
		_w6939_,
		_w6943_,
		_w7164_
	);
	LUT4 #(
		.INIT('h1511)
	) name6702 (
		_w6968_,
		_w7151_,
		_w7163_,
		_w7164_,
		_w7165_
	);
	LUT3 #(
		.INIT('h82)
	) name6703 (
		_w546_,
		_w7153_,
		_w7165_,
		_w7166_
	);
	LUT2 #(
		.INIT('h4)
	) name6704 (
		_w6948_,
		_w6953_,
		_w7167_
	);
	LUT4 #(
		.INIT('h4f00)
	) name6705 (
		_w6885_,
		_w6887_,
		_w6950_,
		_w7167_,
		_w7168_
	);
	LUT3 #(
		.INIT('h51)
	) name6706 (
		_w6974_,
		_w7155_,
		_w7168_,
		_w7169_
	);
	LUT4 #(
		.INIT('h0056)
	) name6707 (
		\P2_IR_reg[28]/NET0131 ,
		_w534_,
		_w536_,
		_w900_,
		_w7170_
	);
	LUT4 #(
		.INIT('h0040)
	) name6708 (
		_w1189_,
		_w1352_,
		_w1356_,
		_w7170_,
		_w7171_
	);
	LUT4 #(
		.INIT('h7d00)
	) name6709 (
		_w1434_,
		_w7157_,
		_w7169_,
		_w7171_,
		_w7172_
	);
	LUT3 #(
		.INIT('h8a)
	) name6710 (
		\P1_state_reg[0]/NET0131 ,
		_w7166_,
		_w7172_,
		_w7173_
	);
	LUT3 #(
		.INIT('hba)
	) name6711 (
		_w2588_,
		_w7162_,
		_w7173_,
		_w7174_
	);
	LUT4 #(
		.INIT('h0056)
	) name6712 (
		\P2_IR_reg[28]/NET0131 ,
		_w534_,
		_w536_,
		_w816_,
		_w7175_
	);
	LUT4 #(
		.INIT('h0040)
	) name6713 (
		_w1189_,
		_w1352_,
		_w1356_,
		_w7175_,
		_w7176_
	);
	LUT4 #(
		.INIT('h6c93)
	) name6714 (
		\P2_IR_reg[0]/NET0131 ,
		\P2_IR_reg[1]/NET0131 ,
		\P2_IR_reg[31]/NET0131 ,
		\P2_reg2_reg[1]/NET0131 ,
		_w7177_
	);
	LUT2 #(
		.INIT('h9)
	) name6715 (
		_w6683_,
		_w7177_,
		_w7178_
	);
	LUT4 #(
		.INIT('h6c93)
	) name6716 (
		\P2_IR_reg[0]/NET0131 ,
		\P2_IR_reg[1]/NET0131 ,
		\P2_IR_reg[31]/NET0131 ,
		\P2_reg1_reg[1]/NET0131 ,
		_w7179_
	);
	LUT2 #(
		.INIT('h9)
	) name6717 (
		_w6661_,
		_w7179_,
		_w7180_
	);
	LUT4 #(
		.INIT('haebf)
	) name6718 (
		_w537_,
		_w545_,
		_w7178_,
		_w7180_,
		_w7181_
	);
	LUT2 #(
		.INIT('h8)
	) name6719 (
		_w7176_,
		_w7181_,
		_w7182_
	);
	LUT3 #(
		.INIT('h02)
	) name6720 (
		\P2_addr_reg[1]/NET0131 ,
		_w537_,
		_w545_,
		_w7183_
	);
	LUT2 #(
		.INIT('h9)
	) name6721 (
		_w6702_,
		_w7177_,
		_w7184_
	);
	LUT3 #(
		.INIT('h80)
	) name6722 (
		_w537_,
		_w545_,
		_w7184_,
		_w7185_
	);
	LUT2 #(
		.INIT('h9)
	) name6723 (
		_w6694_,
		_w7179_,
		_w7186_
	);
	LUT4 #(
		.INIT('hd9fb)
	) name6724 (
		_w537_,
		_w545_,
		_w816_,
		_w7186_,
		_w7187_
	);
	LUT4 #(
		.INIT('h0100)
	) name6725 (
		_w1357_,
		_w7183_,
		_w7185_,
		_w7187_,
		_w7188_
	);
	LUT4 #(
		.INIT('h444e)
	) name6726 (
		\P1_state_reg[0]/NET0131 ,
		\P2_reg3_reg[1]/NET0131 ,
		_w7182_,
		_w7188_,
		_w7189_
	);
	LUT3 #(
		.INIT('h69)
	) name6727 (
		\P2_IR_reg[3]/NET0131 ,
		\P2_reg1_reg[3]/NET0131 ,
		_w794_,
		_w7190_
	);
	LUT4 #(
		.INIT('he817)
	) name6728 (
		\P2_reg1_reg[2]/NET0131 ,
		_w806_,
		_w6695_,
		_w7190_,
		_w7191_
	);
	LUT3 #(
		.INIT('h20)
	) name6729 (
		_w537_,
		_w545_,
		_w7191_,
		_w7192_
	);
	LUT3 #(
		.INIT('h69)
	) name6730 (
		\P2_IR_reg[3]/NET0131 ,
		\P2_reg2_reg[3]/NET0131 ,
		_w794_,
		_w7193_
	);
	LUT4 #(
		.INIT('he817)
	) name6731 (
		\P2_reg2_reg[2]/NET0131 ,
		_w806_,
		_w6703_,
		_w7193_,
		_w7194_
	);
	LUT3 #(
		.INIT('h80)
	) name6732 (
		_w537_,
		_w545_,
		_w7194_,
		_w7195_
	);
	LUT4 #(
		.INIT('hcdfd)
	) name6733 (
		\P2_addr_reg[3]/NET0131 ,
		_w537_,
		_w545_,
		_w795_,
		_w7196_
	);
	LUT4 #(
		.INIT('h0100)
	) name6734 (
		_w1357_,
		_w7192_,
		_w7195_,
		_w7196_,
		_w7197_
	);
	LUT4 #(
		.INIT('h5600)
	) name6735 (
		\P2_IR_reg[28]/NET0131 ,
		_w534_,
		_w536_,
		_w795_,
		_w7198_
	);
	LUT4 #(
		.INIT('h0040)
	) name6736 (
		_w1189_,
		_w1352_,
		_w1356_,
		_w7198_,
		_w7199_
	);
	LUT4 #(
		.INIT('h718e)
	) name6737 (
		\P2_reg1_reg[2]/NET0131 ,
		_w806_,
		_w6662_,
		_w7190_,
		_w7200_
	);
	LUT4 #(
		.INIT('h718e)
	) name6738 (
		\P2_reg2_reg[2]/NET0131 ,
		_w806_,
		_w6684_,
		_w7193_,
		_w7201_
	);
	LUT4 #(
		.INIT('habef)
	) name6739 (
		_w537_,
		_w545_,
		_w7200_,
		_w7201_,
		_w7202_
	);
	LUT3 #(
		.INIT('h2a)
	) name6740 (
		\P1_state_reg[0]/NET0131 ,
		_w7199_,
		_w7202_,
		_w7203_
	);
	LUT3 #(
		.INIT('hba)
	) name6741 (
		_w5855_,
		_w7197_,
		_w7203_,
		_w7204_
	);
	LUT2 #(
		.INIT('h8)
	) name6742 (
		\P1_reg1_reg[18]/NET0131 ,
		_w2191_,
		_w7205_
	);
	LUT4 #(
		.INIT('haf8c)
	) name6743 (
		\P1_reg1_reg[17]/NET0131 ,
		\P1_reg1_reg[18]/NET0131 ,
		_w2178_,
		_w2191_,
		_w7206_
	);
	LUT4 #(
		.INIT('hcd00)
	) name6744 (
		_w6814_,
		_w6855_,
		_w6860_,
		_w7206_,
		_w7207_
	);
	LUT3 #(
		.INIT('h69)
	) name6745 (
		\P1_IR_reg[19]/NET0131 ,
		\P1_reg1_reg[19]/NET0131 ,
		_w2166_,
		_w7208_
	);
	LUT4 #(
		.INIT('ha802)
	) name6746 (
		_w6562_,
		_w7205_,
		_w7207_,
		_w7208_,
		_w7209_
	);
	LUT2 #(
		.INIT('h8)
	) name6747 (
		\P1_reg2_reg[18]/NET0131 ,
		_w2191_,
		_w7210_
	);
	LUT4 #(
		.INIT('haf8c)
	) name6748 (
		\P1_reg2_reg[17]/NET0131 ,
		\P1_reg2_reg[18]/NET0131 ,
		_w2178_,
		_w2191_,
		_w7211_
	);
	LUT4 #(
		.INIT('h010f)
	) name6749 (
		_w6863_,
		_w6866_,
		_w7210_,
		_w7211_,
		_w7212_
	);
	LUT3 #(
		.INIT('h69)
	) name6750 (
		\P1_IR_reg[19]/NET0131 ,
		\P1_reg2_reg[19]/NET0131 ,
		_w2166_,
		_w7213_
	);
	LUT4 #(
		.INIT('h2203)
	) name6751 (
		\P1_addr_reg[19]/NET0131 ,
		_w1747_,
		_w2167_,
		_w6578_,
		_w7214_
	);
	LUT4 #(
		.INIT('h00d7)
	) name6752 (
		_w6577_,
		_w7212_,
		_w7213_,
		_w7214_,
		_w7215_
	);
	LUT4 #(
		.INIT('he2ee)
	) name6753 (
		\P1_reg3_reg[19]/NET0131 ,
		\P1_state_reg[0]/NET0131 ,
		_w7209_,
		_w7215_,
		_w7216_
	);
	LUT2 #(
		.INIT('h6)
	) name6754 (
		\P1_reg1_reg[18]/NET0131 ,
		_w2191_,
		_w7217_
	);
	LUT4 #(
		.INIT('h51f3)
	) name6755 (
		\P1_reg1_reg[16]/NET0131 ,
		\P1_reg1_reg[17]/NET0131 ,
		_w2178_,
		_w2226_,
		_w7218_
	);
	LUT4 #(
		.INIT('hfe00)
	) name6756 (
		_w6759_,
		_w6814_,
		_w6817_,
		_w7218_,
		_w7219_
	);
	LUT4 #(
		.INIT('ha082)
	) name6757 (
		_w6562_,
		_w6854_,
		_w7217_,
		_w7219_,
		_w7220_
	);
	LUT2 #(
		.INIT('h6)
	) name6758 (
		\P1_reg2_reg[18]/NET0131 ,
		_w2191_,
		_w7221_
	);
	LUT4 #(
		.INIT('h1011)
	) name6759 (
		_w6765_,
		_w6820_,
		_w6822_,
		_w6823_,
		_w7222_
	);
	LUT4 #(
		.INIT('h51f3)
	) name6760 (
		\P1_reg2_reg[16]/NET0131 ,
		\P1_reg2_reg[17]/NET0131 ,
		_w2178_,
		_w2226_,
		_w7223_
	);
	LUT3 #(
		.INIT('h45)
	) name6761 (
		_w6862_,
		_w7222_,
		_w7223_,
		_w7224_
	);
	LUT4 #(
		.INIT('h2230)
	) name6762 (
		\P1_addr_reg[18]/NET0131 ,
		_w1747_,
		_w2191_,
		_w6578_,
		_w7225_
	);
	LUT4 #(
		.INIT('h00d7)
	) name6763 (
		_w6577_,
		_w7221_,
		_w7224_,
		_w7225_,
		_w7226_
	);
	LUT4 #(
		.INIT('he2ee)
	) name6764 (
		\P1_reg3_reg[18]/NET0131 ,
		\P1_state_reg[0]/NET0131 ,
		_w7220_,
		_w7226_,
		_w7227_
	);
	LUT4 #(
		.INIT('h0056)
	) name6765 (
		\P2_IR_reg[28]/NET0131 ,
		_w534_,
		_w536_,
		_w806_,
		_w7228_
	);
	LUT4 #(
		.INIT('h0040)
	) name6766 (
		_w1189_,
		_w1352_,
		_w1356_,
		_w7228_,
		_w7229_
	);
	LUT2 #(
		.INIT('h6)
	) name6767 (
		\P2_reg2_reg[2]/NET0131 ,
		_w806_,
		_w7230_
	);
	LUT2 #(
		.INIT('h9)
	) name6768 (
		_w6684_,
		_w7230_,
		_w7231_
	);
	LUT2 #(
		.INIT('h6)
	) name6769 (
		\P2_reg1_reg[2]/NET0131 ,
		_w806_,
		_w7232_
	);
	LUT2 #(
		.INIT('h9)
	) name6770 (
		_w6662_,
		_w7232_,
		_w7233_
	);
	LUT4 #(
		.INIT('haebf)
	) name6771 (
		_w537_,
		_w545_,
		_w7231_,
		_w7233_,
		_w7234_
	);
	LUT2 #(
		.INIT('h8)
	) name6772 (
		_w7229_,
		_w7234_,
		_w7235_
	);
	LUT3 #(
		.INIT('h02)
	) name6773 (
		\P2_addr_reg[2]/NET0131 ,
		_w537_,
		_w545_,
		_w7236_
	);
	LUT2 #(
		.INIT('h9)
	) name6774 (
		_w6695_,
		_w7232_,
		_w7237_
	);
	LUT3 #(
		.INIT('h20)
	) name6775 (
		_w537_,
		_w545_,
		_w7237_,
		_w7238_
	);
	LUT2 #(
		.INIT('h9)
	) name6776 (
		_w6703_,
		_w7230_,
		_w7239_
	);
	LUT4 #(
		.INIT('h73fb)
	) name6777 (
		_w537_,
		_w545_,
		_w806_,
		_w7239_,
		_w7240_
	);
	LUT4 #(
		.INIT('h0100)
	) name6778 (
		_w1357_,
		_w7236_,
		_w7238_,
		_w7240_,
		_w7241_
	);
	LUT4 #(
		.INIT('h444e)
	) name6779 (
		\P1_state_reg[0]/NET0131 ,
		\P2_reg3_reg[2]/NET0131 ,
		_w7235_,
		_w7241_,
		_w7242_
	);
	LUT3 #(
		.INIT('h02)
	) name6780 (
		\P2_addr_reg[4]/NET0131 ,
		_w537_,
		_w545_,
		_w7243_
	);
	LUT4 #(
		.INIT('hc369)
	) name6781 (
		\P2_IR_reg[31]/NET0131 ,
		\P2_IR_reg[4]/NET0131 ,
		\P2_reg1_reg[4]/NET0131 ,
		_w496_,
		_w7244_
	);
	LUT3 #(
		.INIT('h1e)
	) name6782 (
		_w6660_,
		_w6696_,
		_w7244_,
		_w7245_
	);
	LUT3 #(
		.INIT('h20)
	) name6783 (
		_w537_,
		_w545_,
		_w7245_,
		_w7246_
	);
	LUT4 #(
		.INIT('hc369)
	) name6784 (
		\P2_IR_reg[31]/NET0131 ,
		\P2_IR_reg[4]/NET0131 ,
		\P2_reg2_reg[4]/NET0131 ,
		_w496_,
		_w7247_
	);
	LUT3 #(
		.INIT('he1)
	) name6785 (
		_w6681_,
		_w6704_,
		_w7247_,
		_w7248_
	);
	LUT4 #(
		.INIT('h37bf)
	) name6786 (
		_w537_,
		_w545_,
		_w784_,
		_w7248_,
		_w7249_
	);
	LUT4 #(
		.INIT('h0100)
	) name6787 (
		_w1357_,
		_w7243_,
		_w7246_,
		_w7249_,
		_w7250_
	);
	LUT4 #(
		.INIT('h5600)
	) name6788 (
		\P2_IR_reg[28]/NET0131 ,
		_w534_,
		_w536_,
		_w784_,
		_w7251_
	);
	LUT4 #(
		.INIT('h0040)
	) name6789 (
		_w1189_,
		_w1352_,
		_w1356_,
		_w7251_,
		_w7252_
	);
	LUT3 #(
		.INIT('h1e)
	) name6790 (
		_w6681_,
		_w6685_,
		_w7247_,
		_w7253_
	);
	LUT3 #(
		.INIT('h1e)
	) name6791 (
		_w6659_,
		_w6663_,
		_w7244_,
		_w7254_
	);
	LUT4 #(
		.INIT('haebf)
	) name6792 (
		_w537_,
		_w545_,
		_w7253_,
		_w7254_,
		_w7255_
	);
	LUT3 #(
		.INIT('h2a)
	) name6793 (
		\P1_state_reg[0]/NET0131 ,
		_w7252_,
		_w7255_,
		_w7256_
	);
	LUT3 #(
		.INIT('hba)
	) name6794 (
		_w5545_,
		_w7250_,
		_w7256_,
		_w7257_
	);
	LUT3 #(
		.INIT('h57)
	) name6795 (
		\P1_state_reg[0]/NET0131 ,
		_w1748_,
		_w2460_,
		_w7258_
	);
	LUT3 #(
		.INIT('h57)
	) name6796 (
		\P1_state_reg[0]/NET0131 ,
		_w546_,
		_w1357_,
		_w7259_
	);
	LUT4 #(
		.INIT('h2000)
	) name6797 (
		\P1_state_reg[0]/NET0131 ,
		_w1723_,
		_w1727_,
		_w1730_,
		_w7260_
	);
	LUT4 #(
		.INIT('h2000)
	) name6798 (
		\P1_state_reg[0]/NET0131 ,
		_w1189_,
		_w1352_,
		_w1356_,
		_w7261_
	);
	LUT2 #(
		.INIT('h2)
	) name6799 (
		\P1_reg2_reg[22]/NET0131 ,
		_w5244_,
		_w7262_
	);
	LUT2 #(
		.INIT('h2)
	) name6800 (
		\P1_reg2_reg[22]/NET0131 ,
		_w1741_,
		_w7263_
	);
	LUT4 #(
		.INIT('h8288)
	) name6801 (
		_w1741_,
		_w3166_,
		_w3705_,
		_w3707_,
		_w7264_
	);
	LUT4 #(
		.INIT('he020)
	) name6802 (
		\P1_reg2_reg[22]/NET0131 ,
		_w1741_,
		_w2447_,
		_w3693_,
		_w7265_
	);
	LUT4 #(
		.INIT('h0008)
	) name6803 (
		_w1973_,
		_w2284_,
		_w2288_,
		_w2291_,
		_w7266_
	);
	LUT4 #(
		.INIT('h2220)
	) name6804 (
		_w1741_,
		_w1748_,
		_w1966_,
		_w1970_,
		_w7267_
	);
	LUT4 #(
		.INIT('h1113)
	) name6805 (
		_w2426_,
		_w7266_,
		_w7263_,
		_w7267_,
		_w7268_
	);
	LUT2 #(
		.INIT('h4)
	) name6806 (
		_w7265_,
		_w7268_,
		_w7269_
	);
	LUT4 #(
		.INIT('h5700)
	) name6807 (
		_w2388_,
		_w7263_,
		_w7264_,
		_w7269_,
		_w7270_
	);
	LUT4 #(
		.INIT('h2822)
	) name6808 (
		_w1741_,
		_w3166_,
		_w3699_,
		_w3701_,
		_w7271_
	);
	LUT3 #(
		.INIT('ha8)
	) name6809 (
		_w2292_,
		_w7263_,
		_w7271_,
		_w7272_
	);
	LUT4 #(
		.INIT('hddd1)
	) name6810 (
		\P1_reg2_reg[22]/NET0131 ,
		_w1741_,
		_w3689_,
		_w3690_,
		_w7273_
	);
	LUT2 #(
		.INIT('h2)
	) name6811 (
		_w2424_,
		_w7273_,
		_w7274_
	);
	LUT4 #(
		.INIT('ha8aa)
	) name6812 (
		_w5244_,
		_w7272_,
		_w7274_,
		_w7270_,
		_w7275_
	);
	LUT2 #(
		.INIT('he)
	) name6813 (
		_w7262_,
		_w7275_,
		_w7276_
	);
	LUT4 #(
		.INIT('hd070)
	) name6814 (
		\P1_state_reg[0]/NET0131 ,
		\P2_IR_reg[23]/NET0131 ,
		\P2_reg2_reg[26]/NET0131 ,
		_w1188_,
		_w7277_
	);
	LUT4 #(
		.INIT('h2000)
	) name6815 (
		\P2_reg2_reg[26]/NET0131 ,
		_w1189_,
		_w1352_,
		_w1356_,
		_w7278_
	);
	LUT4 #(
		.INIT('haa02)
	) name6816 (
		\P2_reg2_reg[26]/NET0131 ,
		_w1361_,
		_w1363_,
		_w1368_,
		_w7279_
	);
	LUT3 #(
		.INIT('ha8)
	) name6817 (
		_w1530_,
		_w3373_,
		_w7279_,
		_w7280_
	);
	LUT4 #(
		.INIT('h08c8)
	) name6818 (
		\P2_reg2_reg[26]/NET0131 ,
		_w1191_,
		_w1516_,
		_w3258_,
		_w7281_
	);
	LUT4 #(
		.INIT('hf200)
	) name6819 (
		\P2_reg3_reg[26]/NET0131 ,
		_w1029_,
		_w1062_,
		_w1233_,
		_w7282_
	);
	LUT4 #(
		.INIT('h0057)
	) name6820 (
		\P2_reg2_reg[26]/NET0131 ,
		_w1441_,
		_w1523_,
		_w7282_,
		_w7283_
	);
	LUT4 #(
		.INIT('hef00)
	) name6821 (
		_w546_,
		_w1058_,
		_w1522_,
		_w7283_,
		_w7284_
	);
	LUT2 #(
		.INIT('h4)
	) name6822 (
		_w7281_,
		_w7284_,
		_w7285_
	);
	LUT4 #(
		.INIT('ha8aa)
	) name6823 (
		\P2_reg2_reg[26]/NET0131 ,
		_w1361_,
		_w1363_,
		_w1368_,
		_w7286_
	);
	LUT3 #(
		.INIT('h54)
	) name6824 (
		_w1506_,
		_w3380_,
		_w7286_,
		_w7287_
	);
	LUT4 #(
		.INIT('h4844)
	) name6825 (
		_w1257_,
		_w1507_,
		_w3251_,
		_w3253_,
		_w7288_
	);
	LUT3 #(
		.INIT('h54)
	) name6826 (
		_w1575_,
		_w7286_,
		_w7288_,
		_w7289_
	);
	LUT4 #(
		.INIT('h0100)
	) name6827 (
		_w7280_,
		_w7287_,
		_w7289_,
		_w7285_,
		_w7290_
	);
	LUT4 #(
		.INIT('ha0a8)
	) name6828 (
		\P1_state_reg[0]/NET0131 ,
		_w1359_,
		_w7278_,
		_w7290_,
		_w7291_
	);
	LUT2 #(
		.INIT('he)
	) name6829 (
		_w7277_,
		_w7291_,
		_w7292_
	);
	LUT2 #(
		.INIT('h9)
	) name6830 (
		\P1_rd_reg/NET0131 ,
		\P2_rd_reg/NET0131 ,
		_w7293_
	);
	LUT2 #(
		.INIT('h6)
	) name6831 (
		\P1_addr_reg[0]/NET0131 ,
		\P2_addr_reg[0]/NET0131 ,
		_w7294_
	);
	LUT2 #(
		.INIT('h6)
	) name6832 (
		\P1_addr_reg[10]/NET0131 ,
		\P2_addr_reg[10]/NET0131 ,
		_w7295_
	);
	LUT2 #(
		.INIT('h1)
	) name6833 (
		\P1_addr_reg[9]/NET0131 ,
		\P2_addr_reg[9]/NET0131 ,
		_w7296_
	);
	LUT2 #(
		.INIT('h8)
	) name6834 (
		\P1_addr_reg[9]/NET0131 ,
		\P2_addr_reg[9]/NET0131 ,
		_w7297_
	);
	LUT2 #(
		.INIT('h1)
	) name6835 (
		\P1_addr_reg[6]/NET0131 ,
		\P2_addr_reg[6]/NET0131 ,
		_w7298_
	);
	LUT2 #(
		.INIT('h8)
	) name6836 (
		\P1_addr_reg[6]/NET0131 ,
		\P2_addr_reg[6]/NET0131 ,
		_w7299_
	);
	LUT2 #(
		.INIT('h1)
	) name6837 (
		\P1_addr_reg[3]/NET0131 ,
		\P2_addr_reg[3]/NET0131 ,
		_w7300_
	);
	LUT2 #(
		.INIT('h8)
	) name6838 (
		\P1_addr_reg[3]/NET0131 ,
		\P2_addr_reg[3]/NET0131 ,
		_w7301_
	);
	LUT4 #(
		.INIT('hec80)
	) name6839 (
		\P1_addr_reg[0]/NET0131 ,
		\P1_addr_reg[1]/NET0131 ,
		\P2_addr_reg[0]/NET0131 ,
		\P2_addr_reg[1]/NET0131 ,
		_w7302_
	);
	LUT4 #(
		.INIT('h0107)
	) name6840 (
		\P1_addr_reg[2]/NET0131 ,
		\P2_addr_reg[2]/NET0131 ,
		_w7301_,
		_w7302_,
		_w7303_
	);
	LUT4 #(
		.INIT('h888e)
	) name6841 (
		\P1_addr_reg[4]/NET0131 ,
		\P2_addr_reg[4]/NET0131 ,
		_w7300_,
		_w7303_,
		_w7304_
	);
	LUT4 #(
		.INIT('h0107)
	) name6842 (
		\P1_addr_reg[5]/NET0131 ,
		\P2_addr_reg[5]/NET0131 ,
		_w7299_,
		_w7304_,
		_w7305_
	);
	LUT4 #(
		.INIT('h888e)
	) name6843 (
		\P1_addr_reg[7]/NET0131 ,
		\P2_addr_reg[7]/NET0131 ,
		_w7298_,
		_w7305_,
		_w7306_
	);
	LUT4 #(
		.INIT('h0107)
	) name6844 (
		\P1_addr_reg[8]/NET0131 ,
		\P2_addr_reg[8]/NET0131 ,
		_w7297_,
		_w7306_,
		_w7307_
	);
	LUT3 #(
		.INIT('ha9)
	) name6845 (
		_w7295_,
		_w7296_,
		_w7307_,
		_w7308_
	);
	LUT2 #(
		.INIT('h6)
	) name6846 (
		\P1_addr_reg[11]/NET0131 ,
		\P2_addr_reg[11]/NET0131 ,
		_w7309_
	);
	LUT4 #(
		.INIT('h888e)
	) name6847 (
		\P1_addr_reg[10]/NET0131 ,
		\P2_addr_reg[10]/NET0131 ,
		_w7296_,
		_w7307_,
		_w7310_
	);
	LUT2 #(
		.INIT('h6)
	) name6848 (
		_w7309_,
		_w7310_,
		_w7311_
	);
	LUT2 #(
		.INIT('h8)
	) name6849 (
		\P1_addr_reg[12]/NET0131 ,
		\P2_addr_reg[12]/NET0131 ,
		_w7312_
	);
	LUT2 #(
		.INIT('h1)
	) name6850 (
		\P1_addr_reg[12]/NET0131 ,
		\P2_addr_reg[12]/NET0131 ,
		_w7313_
	);
	LUT2 #(
		.INIT('h6)
	) name6851 (
		\P1_addr_reg[12]/NET0131 ,
		\P2_addr_reg[12]/NET0131 ,
		_w7314_
	);
	LUT4 #(
		.INIT('h17e8)
	) name6852 (
		\P1_addr_reg[11]/NET0131 ,
		\P2_addr_reg[11]/NET0131 ,
		_w7310_,
		_w7314_,
		_w7315_
	);
	LUT2 #(
		.INIT('h6)
	) name6853 (
		\P1_addr_reg[13]/NET0131 ,
		\P2_addr_reg[13]/NET0131 ,
		_w7316_
	);
	LUT4 #(
		.INIT('h0017)
	) name6854 (
		\P1_addr_reg[11]/NET0131 ,
		\P2_addr_reg[11]/NET0131 ,
		_w7310_,
		_w7312_,
		_w7317_
	);
	LUT3 #(
		.INIT('hc9)
	) name6855 (
		_w7313_,
		_w7316_,
		_w7317_,
		_w7318_
	);
	LUT2 #(
		.INIT('h6)
	) name6856 (
		\P1_addr_reg[14]/NET0131 ,
		\P2_addr_reg[14]/NET0131 ,
		_w7319_
	);
	LUT4 #(
		.INIT('h888e)
	) name6857 (
		\P1_addr_reg[13]/NET0131 ,
		\P2_addr_reg[13]/NET0131 ,
		_w7313_,
		_w7317_,
		_w7320_
	);
	LUT2 #(
		.INIT('h6)
	) name6858 (
		_w7319_,
		_w7320_,
		_w7321_
	);
	LUT2 #(
		.INIT('h8)
	) name6859 (
		\P1_addr_reg[15]/NET0131 ,
		\P2_addr_reg[15]/NET0131 ,
		_w7322_
	);
	LUT2 #(
		.INIT('h1)
	) name6860 (
		\P1_addr_reg[15]/NET0131 ,
		\P2_addr_reg[15]/NET0131 ,
		_w7323_
	);
	LUT2 #(
		.INIT('h6)
	) name6861 (
		\P1_addr_reg[15]/NET0131 ,
		\P2_addr_reg[15]/NET0131 ,
		_w7324_
	);
	LUT4 #(
		.INIT('h17e8)
	) name6862 (
		\P1_addr_reg[14]/NET0131 ,
		\P2_addr_reg[14]/NET0131 ,
		_w7320_,
		_w7324_,
		_w7325_
	);
	LUT2 #(
		.INIT('h6)
	) name6863 (
		\P1_addr_reg[16]/NET0131 ,
		\P2_addr_reg[16]/NET0131 ,
		_w7326_
	);
	LUT4 #(
		.INIT('h0017)
	) name6864 (
		\P1_addr_reg[14]/NET0131 ,
		\P2_addr_reg[14]/NET0131 ,
		_w7320_,
		_w7322_,
		_w7327_
	);
	LUT3 #(
		.INIT('hc9)
	) name6865 (
		_w7323_,
		_w7326_,
		_w7327_,
		_w7328_
	);
	LUT2 #(
		.INIT('h6)
	) name6866 (
		\P1_addr_reg[17]/NET0131 ,
		\P2_addr_reg[17]/NET0131 ,
		_w7329_
	);
	LUT4 #(
		.INIT('h888e)
	) name6867 (
		\P1_addr_reg[16]/NET0131 ,
		\P2_addr_reg[16]/NET0131 ,
		_w7323_,
		_w7327_,
		_w7330_
	);
	LUT2 #(
		.INIT('h6)
	) name6868 (
		_w7329_,
		_w7330_,
		_w7331_
	);
	LUT2 #(
		.INIT('h8)
	) name6869 (
		\P1_addr_reg[18]/NET0131 ,
		\P2_addr_reg[18]/NET0131 ,
		_w7332_
	);
	LUT2 #(
		.INIT('h1)
	) name6870 (
		\P1_addr_reg[18]/NET0131 ,
		\P2_addr_reg[18]/NET0131 ,
		_w7333_
	);
	LUT2 #(
		.INIT('h6)
	) name6871 (
		\P1_addr_reg[18]/NET0131 ,
		\P2_addr_reg[18]/NET0131 ,
		_w7334_
	);
	LUT4 #(
		.INIT('h17e8)
	) name6872 (
		\P1_addr_reg[17]/NET0131 ,
		\P2_addr_reg[17]/NET0131 ,
		_w7330_,
		_w7334_,
		_w7335_
	);
	LUT2 #(
		.INIT('h6)
	) name6873 (
		\P1_addr_reg[19]/NET0131 ,
		\P2_addr_reg[19]/NET0131 ,
		_w7336_
	);
	LUT4 #(
		.INIT('h0017)
	) name6874 (
		\P1_addr_reg[17]/NET0131 ,
		\P2_addr_reg[17]/NET0131 ,
		_w7330_,
		_w7332_,
		_w7337_
	);
	LUT3 #(
		.INIT('hc9)
	) name6875 (
		_w7333_,
		_w7336_,
		_w7337_,
		_w7338_
	);
	LUT4 #(
		.INIT('h936c)
	) name6876 (
		\P1_addr_reg[0]/NET0131 ,
		\P1_addr_reg[1]/NET0131 ,
		\P2_addr_reg[0]/NET0131 ,
		\P2_addr_reg[1]/NET0131 ,
		_w7339_
	);
	LUT2 #(
		.INIT('h6)
	) name6877 (
		\P1_addr_reg[2]/NET0131 ,
		\P2_addr_reg[2]/NET0131 ,
		_w7340_
	);
	LUT2 #(
		.INIT('h6)
	) name6878 (
		_w7302_,
		_w7340_,
		_w7341_
	);
	LUT2 #(
		.INIT('h6)
	) name6879 (
		\P1_addr_reg[3]/NET0131 ,
		\P2_addr_reg[3]/NET0131 ,
		_w7342_
	);
	LUT4 #(
		.INIT('h17e8)
	) name6880 (
		\P1_addr_reg[2]/NET0131 ,
		\P2_addr_reg[2]/NET0131 ,
		_w7302_,
		_w7342_,
		_w7343_
	);
	LUT2 #(
		.INIT('h6)
	) name6881 (
		\P1_addr_reg[4]/NET0131 ,
		\P2_addr_reg[4]/NET0131 ,
		_w7344_
	);
	LUT3 #(
		.INIT('he1)
	) name6882 (
		_w7300_,
		_w7303_,
		_w7344_,
		_w7345_
	);
	LUT2 #(
		.INIT('h6)
	) name6883 (
		\P1_addr_reg[5]/NET0131 ,
		\P2_addr_reg[5]/NET0131 ,
		_w7346_
	);
	LUT2 #(
		.INIT('h6)
	) name6884 (
		_w7304_,
		_w7346_,
		_w7347_
	);
	LUT2 #(
		.INIT('h6)
	) name6885 (
		\P1_addr_reg[6]/NET0131 ,
		\P2_addr_reg[6]/NET0131 ,
		_w7348_
	);
	LUT4 #(
		.INIT('h17e8)
	) name6886 (
		\P1_addr_reg[5]/NET0131 ,
		\P2_addr_reg[5]/NET0131 ,
		_w7304_,
		_w7348_,
		_w7349_
	);
	LUT2 #(
		.INIT('h6)
	) name6887 (
		\P1_addr_reg[7]/NET0131 ,
		\P2_addr_reg[7]/NET0131 ,
		_w7350_
	);
	LUT3 #(
		.INIT('he1)
	) name6888 (
		_w7298_,
		_w7305_,
		_w7350_,
		_w7351_
	);
	LUT2 #(
		.INIT('h6)
	) name6889 (
		\P1_addr_reg[8]/NET0131 ,
		\P2_addr_reg[8]/NET0131 ,
		_w7352_
	);
	LUT2 #(
		.INIT('h6)
	) name6890 (
		_w7306_,
		_w7352_,
		_w7353_
	);
	LUT2 #(
		.INIT('h6)
	) name6891 (
		\P1_addr_reg[9]/NET0131 ,
		\P2_addr_reg[9]/NET0131 ,
		_w7354_
	);
	LUT4 #(
		.INIT('h17e8)
	) name6892 (
		\P1_addr_reg[8]/NET0131 ,
		\P2_addr_reg[8]/NET0131 ,
		_w7306_,
		_w7354_,
		_w7355_
	);
	LUT2 #(
		.INIT('h9)
	) name6893 (
		\P1_wr_reg/NET0131 ,
		\P2_wr_reg/NET0131 ,
		_w7356_
	);
	assign \P1_state_reg[0]/NET0131_syn_2  = _w216_ ;
	assign \_al_n0  = 1'b0;
	assign \_al_n1  = 1'b1;
	assign \g35/_0_  = _w493_ ;
	assign \g73637/_0_  = _w1350_ ;
	assign \g73647/_0_  = _w1502_ ;
	assign \g73648/_0_  = _w1578_ ;
	assign \g73649/_0_  = _w1595_ ;
	assign \g73650/_0_  = _w1613_ ;
	assign \g73667/_0_  = _w1637_ ;
	assign \g73668/_0_  = _w1654_ ;
	assign \g73669/_0_  = _w1717_ ;
	assign \g73670/_0_  = _w2464_ ;
	assign \g73671/_0_  = _w2479_ ;
	assign \g73672/_0_  = _w2505_ ;
	assign \g73674/_0_  = _w2519_ ;
	assign \g73675/_0_  = _w2532_ ;
	assign \g73709/_0_  = _w2570_ ;
	assign \g73710/_0_  = _w2590_ ;
	assign \g73711/_0_  = _w2612_ ;
	assign \g73716/_0_  = _w2642_ ;
	assign \g73717/_0_  = _w2697_ ;
	assign \g73718/_0_  = _w2714_ ;
	assign \g73719/_0_  = _w2729_ ;
	assign \g73720/_0_  = _w2743_ ;
	assign \g73721/_0_  = _w2853_ ;
	assign \g73722/_0_  = _w2868_ ;
	assign \g73723/_0_  = _w2882_ ;
	assign \g73724/_0_  = _w2897_ ;
	assign \g73765/_0_  = _w2916_ ;
	assign \g73769/_0_  = _w2973_ ;
	assign \g73770/_0_  = _w3001_ ;
	assign \g73771/_0_  = _w3029_ ;
	assign \g73772/_0_  = _w3047_ ;
	assign \g73773/_0_  = _w3061_ ;
	assign \g73774/_0_  = _w3079_ ;
	assign \g73775/_0_  = _w3093_ ;
	assign \g73776/_0_  = _w3216_ ;
	assign \g73777/_0_  = _w3231_ ;
	assign \g73778/_0_  = _w3246_ ;
	assign \g73779/_0_  = _w3278_ ;
	assign \g73780/_0_  = _w3296_ ;
	assign \g73781/_0_  = _w3311_ ;
	assign \g73782/_0_  = _w3326_ ;
	assign \g73783/_0_  = _w3341_ ;
	assign \g73784/_0_  = _w3354_ ;
	assign \g73785/_0_  = _w3369_ ;
	assign \g73786/_0_  = _w3386_ ;
	assign \g73787/_0_  = _w3401_ ;
	assign \g73788/_0_  = _w3415_ ;
	assign \g73789/_0_  = _w3426_ ;
	assign \g73790/_0_  = _w3436_ ;
	assign \g73791/_0_  = _w3449_ ;
	assign \g73792/_0_  = _w3462_ ;
	assign \g73845/_0_  = _w3483_ ;
	assign \g73846/_0_  = _w3504_ ;
	assign \g73847/_0_  = _w3525_ ;
	assign \g73848/_0_  = _w3548_ ;
	assign \g73860/_0_  = _w3563_ ;
	assign \g73863/_0_  = _w3580_ ;
	assign \g73864/_0_  = _w3606_ ;
	assign \g73867/_0_  = _w3626_ ;
	assign \g73870/_0_  = _w3642_ ;
	assign \g73871/_0_  = _w3656_ ;
	assign \g73872/_0_  = _w3669_ ;
	assign \g73873/_0_  = _w3685_ ;
	assign \g73874/_0_  = _w3711_ ;
	assign \g73875/_0_  = _w3726_ ;
	assign \g73876/_0_  = _w3738_ ;
	assign \g73877/_0_  = _w3753_ ;
	assign \g73878/_0_  = _w3769_ ;
	assign \g73879/_0_  = _w3784_ ;
	assign \g73880/_0_  = _w3795_ ;
	assign \g73924/_0_  = _w3814_ ;
	assign \g73925/_0_  = _w3833_ ;
	assign \g73949/_0_  = _w3852_ ;
	assign \g73950/_0_  = _w3868_ ;
	assign \g73953/_0_  = _w3880_ ;
	assign \g73954/_0_  = _w3894_ ;
	assign \g73955/_0_  = _w3911_ ;
	assign \g73956/_0_  = _w3924_ ;
	assign \g73957/_0_  = _w3937_ ;
	assign \g73958/_0_  = _w3951_ ;
	assign \g73960/_0_  = _w3964_ ;
	assign \g73961/_0_  = _w3975_ ;
	assign \g73962/_0_  = _w3989_ ;
	assign \g73963/_0_  = _w4004_ ;
	assign \g73964/_0_  = _w4016_ ;
	assign \g73965/_0_  = _w4029_ ;
	assign \g73966/_0_  = _w4046_ ;
	assign \g73967/_0_  = _w4061_ ;
	assign \g73968/_0_  = _w4074_ ;
	assign \g73969/_0_  = _w4088_ ;
	assign \g73970/_0_  = _w4101_ ;
	assign \g73971/_0_  = _w4113_ ;
	assign \g73972/_0_  = _w4126_ ;
	assign \g73973/_0_  = _w4138_ ;
	assign \g73974/_0_  = _w4149_ ;
	assign \g73975/_0_  = _w4158_ ;
	assign \g73976/_0_  = _w4170_ ;
	assign \g73977/_0_  = _w4182_ ;
	assign \g73978/_0_  = _w4194_ ;
	assign \g73979/_0_  = _w4205_ ;
	assign \g73980/_0_  = _w4214_ ;
	assign \g74062/_0_  = _w4234_ ;
	assign \g74063/_0_  = _w4252_ ;
	assign \g74064/_0_  = _w4275_ ;
	assign \g74065/_0_  = _w4295_ ;
	assign \g74066/_0_  = _w4316_ ;
	assign \g74071/_0_  = _w4335_ ;
	assign \g74072/_0_  = _w4357_ ;
	assign \g74105/_0_  = _w4384_ ;
	assign \g74106/_0_  = _w4402_ ;
	assign \g74107/_0_  = _w4420_ ;
	assign \g74108/_0_  = _w4436_ ;
	assign \g74109/_0_  = _w4447_ ;
	assign \g74110/_0_  = _w4462_ ;
	assign \g74111/_0_  = _w4475_ ;
	assign \g74112/_0_  = _w4489_ ;
	assign \g74113/_0_  = _w4500_ ;
	assign \g74114/_0_  = _w4513_ ;
	assign \g74115/_0_  = _w4529_ ;
	assign \g74167/_0_  = _w4547_ ;
	assign \g74168/_0_  = _w4566_ ;
	assign \g74169/_0_  = _w4588_ ;
	assign \g74170/_0_  = _w4608_ ;
	assign \g74172/_0_  = _w4628_ ;
	assign \g74173/_0_  = _w4650_ ;
	assign \g74174/_0_  = _w4667_ ;
	assign \g74175/_0_  = _w4686_ ;
	assign \g74225/_0_  = _w4703_ ;
	assign \g74226/_0_  = _w4718_ ;
	assign \g74227/_0_  = _w4735_ ;
	assign \g74229/_0_  = _w4751_ ;
	assign \g74230/_0_  = _w4766_ ;
	assign \g74231/_0_  = _w4783_ ;
	assign \g74232/_0_  = _w4795_ ;
	assign \g74233/_0_  = _w4813_ ;
	assign \g74234/_0_  = _w4827_ ;
	assign \g74235/_0_  = _w4841_ ;
	assign \g74236/_0_  = _w4859_ ;
	assign \g74237/_0_  = _w4871_ ;
	assign \g74238/_0_  = _w4886_ ;
	assign \g74239/_0_  = _w4902_ ;
	assign \g74240/_0_  = _w4916_ ;
	assign \g74241/_0_  = _w4930_ ;
	assign \g74242/_0_  = _w4947_ ;
	assign \g74243/_0_  = _w4962_ ;
	assign \g74244/_0_  = _w4978_ ;
	assign \g74245/_0_  = _w4990_ ;
	assign \g74246/_0_  = _w5000_ ;
	assign \g74247/_0_  = _w5008_ ;
	assign \g74248/_0_  = _w5023_ ;
	assign \g74249/_0_  = _w5038_ ;
	assign \g74250/_0_  = _w5050_ ;
	assign \g74251/_0_  = _w5060_ ;
	assign \g74252/_0_  = _w5075_ ;
	assign \g74253/_0_  = _w5088_ ;
	assign \g74254/_0_  = _w5101_ ;
	assign \g74255/_0_  = _w5109_ ;
	assign \g74330/_0_  = _w5128_ ;
	assign \g74331/_0_  = _w5147_ ;
	assign \g74333/_0_  = _w5172_ ;
	assign \g74334/_0_  = _w5194_ ;
	assign \g74335/_0_  = _w5215_ ;
	assign \g74390/_0_  = _w5229_ ;
	assign \g74391/_0_  = _w5242_ ;
	assign \g74405/_0_  = _w5252_ ;
	assign \g74407/_0_  = _w5268_ ;
	assign \g74408/_0_  = _w5277_ ;
	assign \g74409/_0_  = _w5294_ ;
	assign \g74410/_0_  = _w5308_ ;
	assign \g74411/_0_  = _w5321_ ;
	assign \g74412/_0_  = _w5338_ ;
	assign \g74413/_0_  = _w5353_ ;
	assign \g74414/_0_  = _w5370_ ;
	assign \g74415/_0_  = _w5386_ ;
	assign \g74416/_0_  = _w5401_ ;
	assign \g74417/_0_  = _w5419_ ;
	assign \g74418/_0_  = _w5431_ ;
	assign \g74419/_0_  = _w5437_ ;
	assign \g74420/_0_  = _w5449_ ;
	assign \g74421/_0_  = _w5463_ ;
	assign \g74422/_0_  = _w5477_ ;
	assign \g74483/_0_  = _w5492_ ;
	assign \g74485/_0_  = _w5511_ ;
	assign \g74486/_0_  = _w5530_ ;
	assign \g74487/_0_  = _w5548_ ;
	assign \g74576/_0_  = _w5565_ ;
	assign \g74578/_0_  = _w5579_ ;
	assign \g74581/_0_  = _w5596_ ;
	assign \g74582/_0_  = _w5612_ ;
	assign \g74583/_0_  = _w5626_ ;
	assign \g74584/_0_  = _w5640_ ;
	assign \g74585/_0_  = _w5654_ ;
	assign \g74588/_0_  = _w5672_ ;
	assign \g74589/_0_  = _w5689_ ;
	assign \g74590/_0_  = _w5703_ ;
	assign \g74591/_0_  = _w5716_ ;
	assign \g74592/_0_  = _w5729_ ;
	assign \g74595/_0_  = _w5746_ ;
	assign \g74596/_0_  = _w5762_ ;
	assign \g74597/_0_  = _w5777_ ;
	assign \g74598/_0_  = _w5791_ ;
	assign \g74599/_0_  = _w5802_ ;
	assign \g74600/_0_  = _w5815_ ;
	assign \g74601/_0_  = _w5828_ ;
	assign \g74602/_0_  = _w5839_ ;
	assign \g74711/_0_  = _w5857_ ;
	assign \g74835/_0_  = _w5870_ ;
	assign \g74836/_0_  = _w5884_ ;
	assign \g74838/_0_  = _w5897_ ;
	assign \g74840/_0_  = _w5914_ ;
	assign \g74841/_0_  = _w5928_ ;
	assign \g74843/_0_  = _w5940_ ;
	assign \g74844/_0_  = _w5952_ ;
	assign \g74963/_0_  = _w5967_ ;
	assign \g75075/_0_  = _w5982_ ;
	assign \g75078/_0_  = _w5998_ ;
	assign \g75079/_0_  = _w6011_ ;
	assign \g75083/_0_  = _w6023_ ;
	assign \g75084/_0_  = _w6035_ ;
	assign \g75089/_0_  = _w6048_ ;
	assign \g75090/_0_  = _w6061_ ;
	assign \g75091/_0_  = _w6076_ ;
	assign \g75224/_0_  = _w6093_ ;
	assign \g75233/_0_  = _w6111_ ;
	assign \g75234/_0_  = _w6129_ ;
	assign \g75427/_0_  = _w6143_ ;
	assign \g75430/_0_  = _w6158_ ;
	assign \g75434/_0_  = _w6172_ ;
	assign \g75436/_0_  = _w6187_ ;
	assign \g75438/_0_  = _w6201_ ;
	assign \g75844/_0_  = _w6214_ ;
	assign \g75850/_0_  = _w6227_ ;
	assign \g75851/_0_  = _w6242_ ;
	assign \g75860/_0_  = _w6257_ ;
	assign \g75865/_0_  = _w6267_ ;
	assign \g75867/_0_  = _w6282_ ;
	assign \g76076/_0_  = _w6297_ ;
	assign \g76375/_0_  = _w6313_ ;
	assign \g76896/_0_  = _w6328_ ;
	assign \g76901/_0_  = _w6345_ ;
	assign \g76905/_0_  = _w6359_ ;
	assign \g77085/_0_  = _w6368_ ;
	assign \g77892/_0_  = _w6373_ ;
	assign \g77897/_0_  = _w6377_ ;
	assign \g77902/_0_  = _w6381_ ;
	assign \g78635/_0_  = _w6394_ ;
	assign \g78636/_0_  = _w6399_ ;
	assign \g78640/_0_  = _w6406_ ;
	assign \g78642/_0_  = _w6415_ ;
	assign \g78645/_0_  = _w6419_ ;
	assign \g78964/_0_  = _w6424_ ;
	assign \g83163/_3_  = _w6426_ ;
	assign \g83164/_3_  = _w6428_ ;
	assign \g83165/_3_  = _w6430_ ;
	assign \g83166/_3_  = _w6432_ ;
	assign \g83167/_3_  = _w6434_ ;
	assign \g83168/_3_  = _w6436_ ;
	assign \g83644/_0_  = _w6440_ ;
	assign \g83645/_0_  = _w6442_ ;
	assign \g83646/_0_  = _w6443_ ;
	assign \g83647/_0_  = _w6445_ ;
	assign \g83648/_0_  = _w6447_ ;
	assign \g83649/_0_  = _w6449_ ;
	assign \g83650/_0_  = _w6451_ ;
	assign \g83651/_0_  = _w6453_ ;
	assign \g83652/_0_  = _w6455_ ;
	assign \g83653/_0_  = _w6457_ ;
	assign \g83654/_0_  = _w6459_ ;
	assign \g83655/_0_  = _w6461_ ;
	assign \g83656/_0_  = _w6463_ ;
	assign \g83657/_0_  = _w6465_ ;
	assign \g83658/_0_  = _w6467_ ;
	assign \g83659/_0_  = _w6469_ ;
	assign \g83660/_0_  = _w6471_ ;
	assign \g83661/_0_  = _w6473_ ;
	assign \g83662/_0_  = _w6475_ ;
	assign \g83663/_0_  = _w6477_ ;
	assign \g83664/_0_  = _w6479_ ;
	assign \g83665/_0_  = _w6481_ ;
	assign \g83666/_0_  = _w6483_ ;
	assign \g83667/_3_  = _w6485_ ;
	assign \g83668/_0_  = _w6487_ ;
	assign \g83669/_0_  = _w6489_ ;
	assign \g83670/_0_  = _w6491_ ;
	assign \g83671/_0_  = _w6493_ ;
	assign \g83715/_3_  = _w6495_ ;
	assign \g83716/_3_  = _w6497_ ;
	assign \g83717/_3_  = _w6499_ ;
	assign \g83718/_3_  = _w6501_ ;
	assign \g83719/_3_  = _w6503_ ;
	assign \g83720/_3_  = _w6505_ ;
	assign \g83721/_3_  = _w6507_ ;
	assign \g83722/_3_  = _w6509_ ;
	assign \g83723/_3_  = _w6511_ ;
	assign \g83724/_3_  = _w6513_ ;
	assign \g83725/_0_  = _w6515_ ;
	assign \g83726/_3_  = _w6517_ ;
	assign \g83727/_3_  = _w6519_ ;
	assign \g83728/_3_  = _w6521_ ;
	assign \g83729/_3_  = _w6522_ ;
	assign \g83730/_3_  = _w6524_ ;
	assign \g83731/_3_  = _w6526_ ;
	assign \g83732/_3_  = _w6528_ ;
	assign \g83733/_3_  = _w6530_ ;
	assign \g83734/_3_  = _w6532_ ;
	assign \g83735/_0_  = _w6536_ ;
	assign \g83736/_0_  = _w6538_ ;
	assign \g83737/_0_  = _w6540_ ;
	assign \g83738/_3_  = _w6542_ ;
	assign \g83739/_3_  = _w6544_ ;
	assign \g83740/_0_  = _w6546_ ;
	assign \g83741/_3_  = _w6548_ ;
	assign \g83742/_3_  = _w6550_ ;
	assign \g84164/_0_  = _w2088_ ;
	assign \g84181/_0_  = _w825_ ;
	assign \g85146/_0_  = _w6581_ ;
	assign \g85147/_0_  = _w6614_ ;
	assign \g85148/_0_  = _w6622_ ;
	assign \g85149/_0_  = _w6629_ ;
	assign \g85151/_0_  = _w6648_ ;
	assign \g85152/_0_  = _w6716_ ;
	assign \g85154/_0_  = _w6724_ ;
	assign \g85155/_0_  = _w6730_ ;
	assign \g85156/_0_  = _w6739_ ;
	assign \g85157/_0_  = _w6747_ ;
	assign \g85158/_0_  = _w6758_ ;
	assign \g85159/_0_  = _w6769_ ;
	assign \g85160/_0_  = _w6813_ ;
	assign \g85161/_0_  = _w6826_ ;
	assign \g85162/_0_  = _w6853_ ;
	assign \g85163/_0_  = _w6869_ ;
	assign \g85164/_0_  = _w6900_ ;
	assign \g85165/_0_  = _w6937_ ;
	assign \g85166/_0_  = _w6966_ ;
	assign \g85167/_0_  = _w6996_ ;
	assign \g85168/_0_  = _w7016_ ;
	assign \g85169/_0_  = _w7023_ ;
	assign \g85171/_0_  = _w7030_ ;
	assign \g85173/_0_  = _w7037_ ;
	assign \g85174/_0_  = _w7044_ ;
	assign \g85175/_0_  = _w7051_ ;
	assign \g85176/_0_  = _w7062_ ;
	assign \g85178/_0_  = _w7078_ ;
	assign \g85179/_0_  = _w7091_ ;
	assign \g85180/_0_  = _w7106_ ;
	assign \g85181/_0_  = _w7120_ ;
	assign \g85182/_0_  = _w7134_ ;
	assign \g85183/_0_  = _w7150_ ;
	assign \g85184/_0_  = _w7174_ ;
	assign \g85185/_0_  = _w7189_ ;
	assign \g85186/_0_  = _w7204_ ;
	assign \g85187/_0_  = _w7216_ ;
	assign \g85188/_0_  = _w7227_ ;
	assign \g85189/_0_  = _w7242_ ;
	assign \g85190/_0_  = _w7257_ ;
	assign \g85510/_0_  = _w7258_ ;
	assign \g85711/u3_syn_4  = _w6386_ ;
	assign \g85972/_0_  = _w7259_ ;
	assign \g86107/_0_  = _w1738_ ;
	assign \g86200/u3_syn_4  = _w5244_ ;
	assign \g86477/_0_  = _w1740_ ;
	assign \g86548/_0_  = _w1368_ ;
	assign \g86652/u3_syn_4  = _w7260_ ;
	assign \g86807/u3_syn_4  = _w7261_ ;
	assign \g87581/_0_  = _w2277_ ;
	assign \g88104/_0_  = _w1116_ ;
	assign \g88112/_0_  = _w2021_ ;
	assign \g88136/_0_  = _w2087_ ;
	assign \g88148/_0_  = _w2139_ ;
	assign \g88157/_0_  = _w1988_ ;
	assign \g88171/_0_  = _w2062_ ;
	assign \g88179/_0_  = _w2109_ ;
	assign \g88208/_0_  = _w2164_ ;
	assign \g88217/_0_  = _w2201_ ;
	assign \g88222/_0_  = _w2176_ ;
	assign \g88228/_0_  = _w1976_ ;
	assign \g88236/_0_  = _w2236_ ;
	assign \g88242/_0_  = _w2188_ ;
	assign \g88252_dup/_0_  = _w1139_ ;
	assign \g88253/_2_  = _w1086_ ;
	assign \g88259/_0_  = _w1164_ ;
	assign \g88274/_0_  = _w1937_ ;
	assign \g88286/_0_  = _w1963_ ;
	assign \g88296/_0_  = _w1953_ ;
	assign \g88306/_0_  = _w1877_ ;
	assign \g88319/_0_  = _w1837_ ;
	assign \g88330/_0_  = _w2054_ ;
	assign \g88370/_0_  = _w2035_ ;
	assign \g88375/_0_  = _w2009_ ;
	assign \g88388/_0_  = _w2129_ ;
	assign \g88397/_0_  = _w2045_ ;
	assign \g88404/_0_  = _w2213_ ;
	assign \g88793/_0_  = _w890_ ;
	assign \g88834/_0_  = _w727_ ;
	assign \g88905/_0_  = _w712_ ;
	assign \g88910/_0_  = _w824_ ;
	assign \g88936_dup/_0_  = _w624_ ;
	assign \g88953/_0_  = _w782_ ;
	assign \g88962/_0_  = _w1132_ ;
	assign \g89007/_0_  = _w970_ ;
	assign \g89018/_0_  = _w954_ ;
	assign \g89024/_0_  = _w1007_ ;
	assign \g89031/_0_  = _w990_ ;
	assign \g89066/_0_  = _w748_ ;
	assign \g89082/_0_  = _w771_ ;
	assign \g89097/_0_  = _w815_ ;
	assign \g90677/_1__syn_2  = _w2462_ ;
	assign \g96226/_0_  = _w2247_ ;
	assign \g96236/_0_  = _w2119_ ;
	assign \g96261/_0_  = _w7276_ ;
	assign \g96339/_0_  = _w2078_ ;
	assign \g96380/_1_  = _w1905_ ;
	assign \g96418/_0_  = _w2224_ ;
	assign \g96566/_1_  = _w2420_ ;
	assign \g96574/_0_  = _w2398_ ;
	assign \g96620/_0_  = _w654_ ;
	assign \g96629/_0_  = _w911_ ;
	assign \g96735/_0_  = _w1364_ ;
	assign \g96866/_0_  = _w694_ ;
	assign \g96875/_0_  = _w760_ ;
	assign \g96910/_0_  = _w846_ ;
	assign \g96946/_0_  = _w867_ ;
	assign \g96965/_0_  = _w680_ ;
	assign \g97098/_0_  = _w632_ ;
	assign \g97228/_0_  = _w1070_ ;
	assign \g97231/_0_  = _w1036_ ;
	assign \g97242/_0_  = _w804_ ;
	assign \g97384/_0_  = _w793_ ;
	assign \g97409/_0_  = _w529_ ;
	assign \g97506/_0_  = _w1048_ ;
	assign \g97626/_0_  = _w7292_ ;
	assign rd_pad = _w7293_ ;
	assign \so[0]_pad  = _w7294_ ;
	assign \so[10]_pad  = _w7308_ ;
	assign \so[11]_pad  = _w7311_ ;
	assign \so[12]_pad  = _w7315_ ;
	assign \so[13]_pad  = _w7318_ ;
	assign \so[14]_pad  = _w7321_ ;
	assign \so[15]_pad  = _w7325_ ;
	assign \so[16]_pad  = _w7328_ ;
	assign \so[17]_pad  = _w7331_ ;
	assign \so[18]_pad  = _w7335_ ;
	assign \so[19]_pad  = _w7338_ ;
	assign \so[1]_pad  = _w7339_ ;
	assign \so[2]_pad  = _w7341_ ;
	assign \so[3]_pad  = _w7343_ ;
	assign \so[4]_pad  = _w7345_ ;
	assign \so[5]_pad  = _w7347_ ;
	assign \so[6]_pad  = _w7349_ ;
	assign \so[7]_pad  = _w7351_ ;
	assign \so[8]_pad  = _w7353_ ;
	assign \so[9]_pad  = _w7355_ ;
	assign wr_pad = _w7356_ ;
endmodule;