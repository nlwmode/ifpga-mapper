module top( \B_reg/NET0131  , \IR_reg[0]/NET0131  , \IR_reg[10]/NET0131  , \IR_reg[11]/NET0131  , \IR_reg[12]/NET0131  , \IR_reg[13]/NET0131  , \IR_reg[14]/NET0131  , \IR_reg[15]/NET0131  , \IR_reg[16]/NET0131  , \IR_reg[17]/NET0131  , \IR_reg[18]/NET0131  , \IR_reg[19]/NET0131  , \IR_reg[1]/NET0131  , \IR_reg[20]/NET0131  , \IR_reg[21]/NET0131  , \IR_reg[22]/NET0131  , \IR_reg[23]/NET0131  , \IR_reg[24]/NET0131  , \IR_reg[25]/NET0131  , \IR_reg[26]/NET0131  , \IR_reg[27]/NET0131  , \IR_reg[28]/NET0131  , \IR_reg[29]/NET0131  , \IR_reg[2]/NET0131  , \IR_reg[30]/NET0131  , \IR_reg[31]/NET0131  , \IR_reg[3]/NET0131  , \IR_reg[4]/NET0131  , \IR_reg[5]/NET0131  , \IR_reg[6]/NET0131  , \IR_reg[7]/NET0131  , \IR_reg[8]/NET0131  , \IR_reg[9]/NET0131  , \addr[0]_pad  , \addr[10]_pad  , \addr[11]_pad  , \addr[12]_pad  , \addr[13]_pad  , \addr[14]_pad  , \addr[15]_pad  , \addr[16]_pad  , \addr[17]_pad  , \addr[18]_pad  , \addr[19]_pad  , \addr[1]_pad  , \addr[2]_pad  , \addr[3]_pad  , \addr[4]_pad  , \addr[5]_pad  , \addr[6]_pad  , \addr[7]_pad  , \addr[8]_pad  , \addr[9]_pad  , \d_reg[0]/NET0131  , \d_reg[1]/NET0131  , \datai[0]_pad  , \datai[10]_pad  , \datai[11]_pad  , \datai[12]_pad  , \datai[13]_pad  , \datai[14]_pad  , \datai[15]_pad  , \datai[16]_pad  , \datai[17]_pad  , \datai[18]_pad  , \datai[19]_pad  , \datai[1]_pad  , \datai[20]_pad  , \datai[21]_pad  , \datai[22]_pad  , \datai[23]_pad  , \datai[24]_pad  , \datai[25]_pad  , \datai[26]_pad  , \datai[27]_pad  , \datai[28]_pad  , \datai[29]_pad  , \datai[2]_pad  , \datai[30]_pad  , \datai[31]_pad  , \datai[3]_pad  , \datai[4]_pad  , \datai[5]_pad  , \datai[6]_pad  , \datai[7]_pad  , \datai[8]_pad  , \datai[9]_pad  , \reg0_reg[0]/NET0131  , \reg0_reg[10]/NET0131  , \reg0_reg[11]/NET0131  , \reg0_reg[12]/NET0131  , \reg0_reg[13]/NET0131  , \reg0_reg[14]/NET0131  , \reg0_reg[15]/NET0131  , \reg0_reg[16]/NET0131  , \reg0_reg[17]/NET0131  , \reg0_reg[18]/NET0131  , \reg0_reg[19]/NET0131  , \reg0_reg[1]/NET0131  , \reg0_reg[20]/NET0131  , \reg0_reg[21]/NET0131  , \reg0_reg[22]/NET0131  , \reg0_reg[23]/NET0131  , \reg0_reg[24]/NET0131  , \reg0_reg[25]/NET0131  , \reg0_reg[26]/NET0131  , \reg0_reg[27]/NET0131  , \reg0_reg[28]/NET0131  , \reg0_reg[29]/NET0131  , \reg0_reg[2]/NET0131  , \reg0_reg[30]/NET0131  , \reg0_reg[31]/NET0131  , \reg0_reg[3]/NET0131  , \reg0_reg[4]/NET0131  , \reg0_reg[5]/NET0131  , \reg0_reg[6]/NET0131  , \reg0_reg[7]/NET0131  , \reg0_reg[8]/NET0131  , \reg0_reg[9]/NET0131  , \reg1_reg[0]/NET0131  , \reg1_reg[10]/NET0131  , \reg1_reg[11]/NET0131  , \reg1_reg[12]/NET0131  , \reg1_reg[13]/NET0131  , \reg1_reg[14]/NET0131  , \reg1_reg[15]/NET0131  , \reg1_reg[16]/NET0131  , \reg1_reg[17]/NET0131  , \reg1_reg[18]/NET0131  , \reg1_reg[19]/NET0131  , \reg1_reg[1]/NET0131  , \reg1_reg[20]/NET0131  , \reg1_reg[21]/NET0131  , \reg1_reg[22]/NET0131  , \reg1_reg[23]/NET0131  , \reg1_reg[24]/NET0131  , \reg1_reg[25]/NET0131  , \reg1_reg[26]/NET0131  , \reg1_reg[27]/NET0131  , \reg1_reg[28]/NET0131  , \reg1_reg[29]/NET0131  , \reg1_reg[2]/NET0131  , \reg1_reg[30]/NET0131  , \reg1_reg[31]/NET0131  , \reg1_reg[3]/NET0131  , \reg1_reg[4]/NET0131  , \reg1_reg[5]/NET0131  , \reg1_reg[6]/NET0131  , \reg1_reg[7]/NET0131  , \reg1_reg[8]/NET0131  , \reg1_reg[9]/NET0131  , \reg2_reg[0]/NET0131  , \reg2_reg[10]/NET0131  , \reg2_reg[11]/NET0131  , \reg2_reg[12]/NET0131  , \reg2_reg[13]/NET0131  , \reg2_reg[14]/NET0131  , \reg2_reg[15]/NET0131  , \reg2_reg[16]/NET0131  , \reg2_reg[17]/NET0131  , \reg2_reg[18]/NET0131  , \reg2_reg[19]/NET0131  , \reg2_reg[1]/NET0131  , \reg2_reg[20]/NET0131  , \reg2_reg[21]/NET0131  , \reg2_reg[22]/NET0131  , \reg2_reg[23]/NET0131  , \reg2_reg[24]/NET0131  , \reg2_reg[25]/NET0131  , \reg2_reg[26]/NET0131  , \reg2_reg[27]/NET0131  , \reg2_reg[28]/NET0131  , \reg2_reg[29]/NET0131  , \reg2_reg[2]/NET0131  , \reg2_reg[30]/NET0131  , \reg2_reg[31]/NET0131  , \reg2_reg[3]/NET0131  , \reg2_reg[4]/NET0131  , \reg2_reg[5]/NET0131  , \reg2_reg[6]/NET0131  , \reg2_reg[7]/NET0131  , \reg2_reg[8]/NET0131  , \reg2_reg[9]/NET0131  , \reg3_reg[0]/NET0131  , \reg3_reg[10]/NET0131  , \reg3_reg[11]/NET0131  , \reg3_reg[12]/NET0131  , \reg3_reg[13]/NET0131  , \reg3_reg[14]/NET0131  , \reg3_reg[15]/NET0131  , \reg3_reg[16]/NET0131  , \reg3_reg[17]/NET0131  , \reg3_reg[18]/NET0131  , \reg3_reg[19]/NET0131  , \reg3_reg[1]/NET0131  , \reg3_reg[20]/NET0131  , \reg3_reg[21]/NET0131  , \reg3_reg[22]/NET0131  , \reg3_reg[23]/NET0131  , \reg3_reg[24]/NET0131  , \reg3_reg[25]/NET0131  , \reg3_reg[26]/NET0131  , \reg3_reg[27]/NET0131  , \reg3_reg[28]/NET0131  , \reg3_reg[2]/NET0131  , \reg3_reg[3]/NET0131  , \reg3_reg[4]/NET0131  , \reg3_reg[5]/NET0131  , \reg3_reg[6]/NET0131  , \reg3_reg[7]/NET0131  , \reg3_reg[8]/NET0131  , \reg3_reg[9]/NET0131  , \state_reg[0]/NET0131  , \_al_n0  , \_al_n1  , \g29_dup/_0_  , \g33_dup47063/_0_  , \g36117/_0_  , \g36132/_0_  , \g36133/_0_  , \g36134/_0_  , \g36135/_0_  , \g36136/_0_  , \g36153/_0_  , \g36154/_0_  , \g36155/_0_  , \g36156/_0_  , \g36157/_0_  , \g36158/_0_  , \g36186/_0_  , \g36187/_0_  , \g36193/_0_  , \g36197/_0_  , \g36198/_0_  , \g36199/_0_  , \g36200/_0_  , \g36201/_0_  , \g36202/_0_  , \g36203/_0_  , \g36204/_0_  , \g36239/_0_  , \g36240/_0_  , \g36242/_0_  , \g36246/_0_  , \g36255/_0_  , \g36259/_0_  , \g36260/_0_  , \g36261/_0_  , \g36262/_0_  , \g36263/_0_  , \g36264/_0_  , \g36265/_0_  , \g36266/_0_  , \g36267/_0_  , \g36268/_0_  , \g36269/_0_  , \g36270/_0_  , \g36271/_0_  , \g36272/_0_  , \g36273/_0_  , \g36274/_0_  , \g36321/_0_  , \g36322/_0_  , \g36323/_0_  , \g36324/_0_  , \g36325/_0_  , \g36341/_0_  , \g36343/_0_  , \g36344/_0_  , \g36345/_0_  , \g36346/_0_  , \g36347/_0_  , \g36348/_0_  , \g36349/_0_  , \g36350/_0_  , \g36351/_0_  , \g36352/_0_  , \g36353/_0_  , \g36354/_0_  , \g36355/_0_  , \g36356/_0_  , \g36357/_0_  , \g36358/_0_  , \g36359/_0_  , \g36360/_0_  , \g36361/_0_  , \g36362/_0_  , \g36363/_0_  , \g36410/_0_  , \g36413/_0_  , \g36414/_0_  , \g36415/_0_  , \g36416/_0_  , \g36424/_0_  , \g36425/_0_  , \g36452/_0_  , \g36455/_0_  , \g36456/_0_  , \g36457/_0_  , \g36458/_0_  , \g36459/_0_  , \g36460/_0_  , \g36461/_0_  , \g36462/_0_  , \g36463/_0_  , \g36464/_0_  , \g36465/_0_  , \g36466/_0_  , \g36467/_0_  , \g36468/_0_  , \g36469/_0_  , \g36470/_0_  , \g36471/_0_  , \g36472/_0_  , \g36473/_0_  , \g36557/_0_  , \g36558/_0_  , \g36559/_0_  , \g36560/_0_  , \g36561/_0_  , \g36562/_0_  , \g36563/_0_  , \g36564/_0_  , \g36565/_0_  , \g36566/_0_  , \g36567/_0_  , \g36568/_0_  , \g36569/_0_  , \g36570/_0_  , \g36571/_0_  , \g36572/_0_  , \g36573/_0_  , \g36574/_0_  , \g36575/_0_  , \g36576/_0_  , \g36577/_0_  , \g36672/_0_  , \g36673/_0_  , \g36674/_0_  , \g38/_0_  , \g38_dup47616/_1_  , \g39789/u3_syn_4  , \g40089/_0_  , \g40090/_0_  , \g40092/_0_  , \g40093/_0_  , \g40095/_0_  , \g40096/_0_  , \g40097/_0_  , \g40098/_0_  , \g40099/_0_  , \g40100/_0_  , \g40105/_0_  , \g40106/_0_  , \g40108/_0_  , \g40109/_0_  , \g40219/_0_  , \g40220/_0_  , \g40221/_0_  , \g40222/_0_  , \g40223/_0_  , \g40228/_0_  , \g40434/_0_  , \g40495/_0_  , \g40760/_0_  , \g41149/u3_syn_4  , \g42397/_0_  , \g42487/_0_  , \g42553/_0_  , \g43089/_0_  , \g43163/_0_  , \g43169/_0_  , \g43180/_0_  , \g43189_dup/_0_  , \g43196/_0_  , \g43217/_0_  , \g43236/_0_  , \g43251/_0_  , \g43256/_0_  , \g43272/_0_  , \g43277/_0_  , \g43324/_0_  , \g43341/_0_  , \g43350/_0_  , \g43360/_0_  , \g44419/_3_  , \g44452/_3_  , \g44514/_3_  , \g44515/_3_  , \g44516/_3_  , \g44583/_3_  , \g44586/_3_  , \g44587/_3_  , \g44588/_3_  , \g44589/_3_  , \g44590/_3_  , \g44591/_3_  , \g44679/_0_  , \g44680/_3_  , \g44681/_3_  , \g44682/_3_  , \g44686/_3_  , \g44687/_3_  , \g44688/_3_  , \g44689/_3_  , \g44771/_3_  , \g44785/_3_  , \g44795/_3_  , \g44796/_3_  , \g44906/_3_  , \g44968/_3_  , \g44984/_3_  , \g45042/_3_  , \g45044/_3_  , \g45115/_3_  , \g45116/_3_  , \g46478/_1_  , \g46505/_0_  , \g46519/_0_  , \g46696/_0_  , \g47017/_2_  , \g47072_dup/_0_  , \g47395/_0_  , \g47397/_0_  , \g47401/_0_  , \g47404/_0_  , \g47458/_0_  , \g47540/_0_  , \g47791/_0_  , \state_reg[0]/NET0131_syn_2  );
  input \B_reg/NET0131  ;
  input \IR_reg[0]/NET0131  ;
  input \IR_reg[10]/NET0131  ;
  input \IR_reg[11]/NET0131  ;
  input \IR_reg[12]/NET0131  ;
  input \IR_reg[13]/NET0131  ;
  input \IR_reg[14]/NET0131  ;
  input \IR_reg[15]/NET0131  ;
  input \IR_reg[16]/NET0131  ;
  input \IR_reg[17]/NET0131  ;
  input \IR_reg[18]/NET0131  ;
  input \IR_reg[19]/NET0131  ;
  input \IR_reg[1]/NET0131  ;
  input \IR_reg[20]/NET0131  ;
  input \IR_reg[21]/NET0131  ;
  input \IR_reg[22]/NET0131  ;
  input \IR_reg[23]/NET0131  ;
  input \IR_reg[24]/NET0131  ;
  input \IR_reg[25]/NET0131  ;
  input \IR_reg[26]/NET0131  ;
  input \IR_reg[27]/NET0131  ;
  input \IR_reg[28]/NET0131  ;
  input \IR_reg[29]/NET0131  ;
  input \IR_reg[2]/NET0131  ;
  input \IR_reg[30]/NET0131  ;
  input \IR_reg[31]/NET0131  ;
  input \IR_reg[3]/NET0131  ;
  input \IR_reg[4]/NET0131  ;
  input \IR_reg[5]/NET0131  ;
  input \IR_reg[6]/NET0131  ;
  input \IR_reg[7]/NET0131  ;
  input \IR_reg[8]/NET0131  ;
  input \IR_reg[9]/NET0131  ;
  input \addr[0]_pad  ;
  input \addr[10]_pad  ;
  input \addr[11]_pad  ;
  input \addr[12]_pad  ;
  input \addr[13]_pad  ;
  input \addr[14]_pad  ;
  input \addr[15]_pad  ;
  input \addr[16]_pad  ;
  input \addr[17]_pad  ;
  input \addr[18]_pad  ;
  input \addr[19]_pad  ;
  input \addr[1]_pad  ;
  input \addr[2]_pad  ;
  input \addr[3]_pad  ;
  input \addr[4]_pad  ;
  input \addr[5]_pad  ;
  input \addr[6]_pad  ;
  input \addr[7]_pad  ;
  input \addr[8]_pad  ;
  input \addr[9]_pad  ;
  input \d_reg[0]/NET0131  ;
  input \d_reg[1]/NET0131  ;
  input \datai[0]_pad  ;
  input \datai[10]_pad  ;
  input \datai[11]_pad  ;
  input \datai[12]_pad  ;
  input \datai[13]_pad  ;
  input \datai[14]_pad  ;
  input \datai[15]_pad  ;
  input \datai[16]_pad  ;
  input \datai[17]_pad  ;
  input \datai[18]_pad  ;
  input \datai[19]_pad  ;
  input \datai[1]_pad  ;
  input \datai[20]_pad  ;
  input \datai[21]_pad  ;
  input \datai[22]_pad  ;
  input \datai[23]_pad  ;
  input \datai[24]_pad  ;
  input \datai[25]_pad  ;
  input \datai[26]_pad  ;
  input \datai[27]_pad  ;
  input \datai[28]_pad  ;
  input \datai[29]_pad  ;
  input \datai[2]_pad  ;
  input \datai[30]_pad  ;
  input \datai[31]_pad  ;
  input \datai[3]_pad  ;
  input \datai[4]_pad  ;
  input \datai[5]_pad  ;
  input \datai[6]_pad  ;
  input \datai[7]_pad  ;
  input \datai[8]_pad  ;
  input \datai[9]_pad  ;
  input \reg0_reg[0]/NET0131  ;
  input \reg0_reg[10]/NET0131  ;
  input \reg0_reg[11]/NET0131  ;
  input \reg0_reg[12]/NET0131  ;
  input \reg0_reg[13]/NET0131  ;
  input \reg0_reg[14]/NET0131  ;
  input \reg0_reg[15]/NET0131  ;
  input \reg0_reg[16]/NET0131  ;
  input \reg0_reg[17]/NET0131  ;
  input \reg0_reg[18]/NET0131  ;
  input \reg0_reg[19]/NET0131  ;
  input \reg0_reg[1]/NET0131  ;
  input \reg0_reg[20]/NET0131  ;
  input \reg0_reg[21]/NET0131  ;
  input \reg0_reg[22]/NET0131  ;
  input \reg0_reg[23]/NET0131  ;
  input \reg0_reg[24]/NET0131  ;
  input \reg0_reg[25]/NET0131  ;
  input \reg0_reg[26]/NET0131  ;
  input \reg0_reg[27]/NET0131  ;
  input \reg0_reg[28]/NET0131  ;
  input \reg0_reg[29]/NET0131  ;
  input \reg0_reg[2]/NET0131  ;
  input \reg0_reg[30]/NET0131  ;
  input \reg0_reg[31]/NET0131  ;
  input \reg0_reg[3]/NET0131  ;
  input \reg0_reg[4]/NET0131  ;
  input \reg0_reg[5]/NET0131  ;
  input \reg0_reg[6]/NET0131  ;
  input \reg0_reg[7]/NET0131  ;
  input \reg0_reg[8]/NET0131  ;
  input \reg0_reg[9]/NET0131  ;
  input \reg1_reg[0]/NET0131  ;
  input \reg1_reg[10]/NET0131  ;
  input \reg1_reg[11]/NET0131  ;
  input \reg1_reg[12]/NET0131  ;
  input \reg1_reg[13]/NET0131  ;
  input \reg1_reg[14]/NET0131  ;
  input \reg1_reg[15]/NET0131  ;
  input \reg1_reg[16]/NET0131  ;
  input \reg1_reg[17]/NET0131  ;
  input \reg1_reg[18]/NET0131  ;
  input \reg1_reg[19]/NET0131  ;
  input \reg1_reg[1]/NET0131  ;
  input \reg1_reg[20]/NET0131  ;
  input \reg1_reg[21]/NET0131  ;
  input \reg1_reg[22]/NET0131  ;
  input \reg1_reg[23]/NET0131  ;
  input \reg1_reg[24]/NET0131  ;
  input \reg1_reg[25]/NET0131  ;
  input \reg1_reg[26]/NET0131  ;
  input \reg1_reg[27]/NET0131  ;
  input \reg1_reg[28]/NET0131  ;
  input \reg1_reg[29]/NET0131  ;
  input \reg1_reg[2]/NET0131  ;
  input \reg1_reg[30]/NET0131  ;
  input \reg1_reg[31]/NET0131  ;
  input \reg1_reg[3]/NET0131  ;
  input \reg1_reg[4]/NET0131  ;
  input \reg1_reg[5]/NET0131  ;
  input \reg1_reg[6]/NET0131  ;
  input \reg1_reg[7]/NET0131  ;
  input \reg1_reg[8]/NET0131  ;
  input \reg1_reg[9]/NET0131  ;
  input \reg2_reg[0]/NET0131  ;
  input \reg2_reg[10]/NET0131  ;
  input \reg2_reg[11]/NET0131  ;
  input \reg2_reg[12]/NET0131  ;
  input \reg2_reg[13]/NET0131  ;
  input \reg2_reg[14]/NET0131  ;
  input \reg2_reg[15]/NET0131  ;
  input \reg2_reg[16]/NET0131  ;
  input \reg2_reg[17]/NET0131  ;
  input \reg2_reg[18]/NET0131  ;
  input \reg2_reg[19]/NET0131  ;
  input \reg2_reg[1]/NET0131  ;
  input \reg2_reg[20]/NET0131  ;
  input \reg2_reg[21]/NET0131  ;
  input \reg2_reg[22]/NET0131  ;
  input \reg2_reg[23]/NET0131  ;
  input \reg2_reg[24]/NET0131  ;
  input \reg2_reg[25]/NET0131  ;
  input \reg2_reg[26]/NET0131  ;
  input \reg2_reg[27]/NET0131  ;
  input \reg2_reg[28]/NET0131  ;
  input \reg2_reg[29]/NET0131  ;
  input \reg2_reg[2]/NET0131  ;
  input \reg2_reg[30]/NET0131  ;
  input \reg2_reg[31]/NET0131  ;
  input \reg2_reg[3]/NET0131  ;
  input \reg2_reg[4]/NET0131  ;
  input \reg2_reg[5]/NET0131  ;
  input \reg2_reg[6]/NET0131  ;
  input \reg2_reg[7]/NET0131  ;
  input \reg2_reg[8]/NET0131  ;
  input \reg2_reg[9]/NET0131  ;
  input \reg3_reg[0]/NET0131  ;
  input \reg3_reg[10]/NET0131  ;
  input \reg3_reg[11]/NET0131  ;
  input \reg3_reg[12]/NET0131  ;
  input \reg3_reg[13]/NET0131  ;
  input \reg3_reg[14]/NET0131  ;
  input \reg3_reg[15]/NET0131  ;
  input \reg3_reg[16]/NET0131  ;
  input \reg3_reg[17]/NET0131  ;
  input \reg3_reg[18]/NET0131  ;
  input \reg3_reg[19]/NET0131  ;
  input \reg3_reg[1]/NET0131  ;
  input \reg3_reg[20]/NET0131  ;
  input \reg3_reg[21]/NET0131  ;
  input \reg3_reg[22]/NET0131  ;
  input \reg3_reg[23]/NET0131  ;
  input \reg3_reg[24]/NET0131  ;
  input \reg3_reg[25]/NET0131  ;
  input \reg3_reg[26]/NET0131  ;
  input \reg3_reg[27]/NET0131  ;
  input \reg3_reg[28]/NET0131  ;
  input \reg3_reg[2]/NET0131  ;
  input \reg3_reg[3]/NET0131  ;
  input \reg3_reg[4]/NET0131  ;
  input \reg3_reg[5]/NET0131  ;
  input \reg3_reg[6]/NET0131  ;
  input \reg3_reg[7]/NET0131  ;
  input \reg3_reg[8]/NET0131  ;
  input \reg3_reg[9]/NET0131  ;
  input \state_reg[0]/NET0131  ;
  output \_al_n0  ;
  output \_al_n1  ;
  output \g29_dup/_0_  ;
  output \g33_dup47063/_0_  ;
  output \g36117/_0_  ;
  output \g36132/_0_  ;
  output \g36133/_0_  ;
  output \g36134/_0_  ;
  output \g36135/_0_  ;
  output \g36136/_0_  ;
  output \g36153/_0_  ;
  output \g36154/_0_  ;
  output \g36155/_0_  ;
  output \g36156/_0_  ;
  output \g36157/_0_  ;
  output \g36158/_0_  ;
  output \g36186/_0_  ;
  output \g36187/_0_  ;
  output \g36193/_0_  ;
  output \g36197/_0_  ;
  output \g36198/_0_  ;
  output \g36199/_0_  ;
  output \g36200/_0_  ;
  output \g36201/_0_  ;
  output \g36202/_0_  ;
  output \g36203/_0_  ;
  output \g36204/_0_  ;
  output \g36239/_0_  ;
  output \g36240/_0_  ;
  output \g36242/_0_  ;
  output \g36246/_0_  ;
  output \g36255/_0_  ;
  output \g36259/_0_  ;
  output \g36260/_0_  ;
  output \g36261/_0_  ;
  output \g36262/_0_  ;
  output \g36263/_0_  ;
  output \g36264/_0_  ;
  output \g36265/_0_  ;
  output \g36266/_0_  ;
  output \g36267/_0_  ;
  output \g36268/_0_  ;
  output \g36269/_0_  ;
  output \g36270/_0_  ;
  output \g36271/_0_  ;
  output \g36272/_0_  ;
  output \g36273/_0_  ;
  output \g36274/_0_  ;
  output \g36321/_0_  ;
  output \g36322/_0_  ;
  output \g36323/_0_  ;
  output \g36324/_0_  ;
  output \g36325/_0_  ;
  output \g36341/_0_  ;
  output \g36343/_0_  ;
  output \g36344/_0_  ;
  output \g36345/_0_  ;
  output \g36346/_0_  ;
  output \g36347/_0_  ;
  output \g36348/_0_  ;
  output \g36349/_0_  ;
  output \g36350/_0_  ;
  output \g36351/_0_  ;
  output \g36352/_0_  ;
  output \g36353/_0_  ;
  output \g36354/_0_  ;
  output \g36355/_0_  ;
  output \g36356/_0_  ;
  output \g36357/_0_  ;
  output \g36358/_0_  ;
  output \g36359/_0_  ;
  output \g36360/_0_  ;
  output \g36361/_0_  ;
  output \g36362/_0_  ;
  output \g36363/_0_  ;
  output \g36410/_0_  ;
  output \g36413/_0_  ;
  output \g36414/_0_  ;
  output \g36415/_0_  ;
  output \g36416/_0_  ;
  output \g36424/_0_  ;
  output \g36425/_0_  ;
  output \g36452/_0_  ;
  output \g36455/_0_  ;
  output \g36456/_0_  ;
  output \g36457/_0_  ;
  output \g36458/_0_  ;
  output \g36459/_0_  ;
  output \g36460/_0_  ;
  output \g36461/_0_  ;
  output \g36462/_0_  ;
  output \g36463/_0_  ;
  output \g36464/_0_  ;
  output \g36465/_0_  ;
  output \g36466/_0_  ;
  output \g36467/_0_  ;
  output \g36468/_0_  ;
  output \g36469/_0_  ;
  output \g36470/_0_  ;
  output \g36471/_0_  ;
  output \g36472/_0_  ;
  output \g36473/_0_  ;
  output \g36557/_0_  ;
  output \g36558/_0_  ;
  output \g36559/_0_  ;
  output \g36560/_0_  ;
  output \g36561/_0_  ;
  output \g36562/_0_  ;
  output \g36563/_0_  ;
  output \g36564/_0_  ;
  output \g36565/_0_  ;
  output \g36566/_0_  ;
  output \g36567/_0_  ;
  output \g36568/_0_  ;
  output \g36569/_0_  ;
  output \g36570/_0_  ;
  output \g36571/_0_  ;
  output \g36572/_0_  ;
  output \g36573/_0_  ;
  output \g36574/_0_  ;
  output \g36575/_0_  ;
  output \g36576/_0_  ;
  output \g36577/_0_  ;
  output \g36672/_0_  ;
  output \g36673/_0_  ;
  output \g36674/_0_  ;
  output \g38/_0_  ;
  output \g38_dup47616/_1_  ;
  output \g39789/u3_syn_4  ;
  output \g40089/_0_  ;
  output \g40090/_0_  ;
  output \g40092/_0_  ;
  output \g40093/_0_  ;
  output \g40095/_0_  ;
  output \g40096/_0_  ;
  output \g40097/_0_  ;
  output \g40098/_0_  ;
  output \g40099/_0_  ;
  output \g40100/_0_  ;
  output \g40105/_0_  ;
  output \g40106/_0_  ;
  output \g40108/_0_  ;
  output \g40109/_0_  ;
  output \g40219/_0_  ;
  output \g40220/_0_  ;
  output \g40221/_0_  ;
  output \g40222/_0_  ;
  output \g40223/_0_  ;
  output \g40228/_0_  ;
  output \g40434/_0_  ;
  output \g40495/_0_  ;
  output \g40760/_0_  ;
  output \g41149/u3_syn_4  ;
  output \g42397/_0_  ;
  output \g42487/_0_  ;
  output \g42553/_0_  ;
  output \g43089/_0_  ;
  output \g43163/_0_  ;
  output \g43169/_0_  ;
  output \g43180/_0_  ;
  output \g43189_dup/_0_  ;
  output \g43196/_0_  ;
  output \g43217/_0_  ;
  output \g43236/_0_  ;
  output \g43251/_0_  ;
  output \g43256/_0_  ;
  output \g43272/_0_  ;
  output \g43277/_0_  ;
  output \g43324/_0_  ;
  output \g43341/_0_  ;
  output \g43350/_0_  ;
  output \g43360/_0_  ;
  output \g44419/_3_  ;
  output \g44452/_3_  ;
  output \g44514/_3_  ;
  output \g44515/_3_  ;
  output \g44516/_3_  ;
  output \g44583/_3_  ;
  output \g44586/_3_  ;
  output \g44587/_3_  ;
  output \g44588/_3_  ;
  output \g44589/_3_  ;
  output \g44590/_3_  ;
  output \g44591/_3_  ;
  output \g44679/_0_  ;
  output \g44680/_3_  ;
  output \g44681/_3_  ;
  output \g44682/_3_  ;
  output \g44686/_3_  ;
  output \g44687/_3_  ;
  output \g44688/_3_  ;
  output \g44689/_3_  ;
  output \g44771/_3_  ;
  output \g44785/_3_  ;
  output \g44795/_3_  ;
  output \g44796/_3_  ;
  output \g44906/_3_  ;
  output \g44968/_3_  ;
  output \g44984/_3_  ;
  output \g45042/_3_  ;
  output \g45044/_3_  ;
  output \g45115/_3_  ;
  output \g45116/_3_  ;
  output \g46478/_1_  ;
  output \g46505/_0_  ;
  output \g46519/_0_  ;
  output \g46696/_0_  ;
  output \g47017/_2_  ;
  output \g47072_dup/_0_  ;
  output \g47395/_0_  ;
  output \g47397/_0_  ;
  output \g47401/_0_  ;
  output \g47404/_0_  ;
  output \g47458/_0_  ;
  output \g47540/_0_  ;
  output \g47791/_0_  ;
  output \state_reg[0]/NET0131_syn_2  ;
  wire n214 , n215 , n216 , n217 , n218 , n219 , n220 , n221 , n222 , n223 , n224 , n225 , n226 , n227 , n228 , n229 , n230 , n231 , n232 , n233 , n234 , n235 , n236 , n237 , n238 , n239 , n240 , n241 , n242 , n243 , n244 , n245 , n246 , n247 , n248 , n249 , n250 , n251 , n252 , n253 , n254 , n255 , n256 , n257 , n258 , n259 , n260 , n261 , n262 , n263 , n264 , n265 , n266 , n267 , n268 , n269 , n270 , n271 , n272 , n273 , n274 , n275 , n276 , n277 , n278 , n279 , n280 , n281 , n282 , n283 , n284 , n285 , n286 , n287 , n288 , n289 , n290 , n291 , n292 , n293 , n294 , n295 , n296 , n297 , n298 , n299 , n300 , n301 , n302 , n303 , n304 , n305 , n306 , n307 , n308 , n309 , n310 , n311 , n312 , n313 , n314 , n315 , n316 , n317 , n318 , n319 , n320 , n321 , n322 , n323 , n324 , n325 , n326 , n327 , n328 , n329 , n330 , n331 , n332 , n333 , n334 , n335 , n336 , n337 , n338 , n339 , n340 , n341 , n342 , n343 , n344 , n345 , n346 , n347 , n348 , n349 , n350 , n351 , n352 , n353 , n354 , n355 , n356 , n357 , n358 , n359 , n360 , n361 , n362 , n363 , n364 , n365 , n366 , n367 , n368 , n369 , n370 , n371 , n372 , n373 , n374 , n375 , n376 , n377 , n378 , n379 , n380 , n381 , n382 , n383 , n384 , n385 , n386 , n387 , n388 , n389 , n390 , n391 , n392 , n393 , n394 , n395 , n396 , n397 , n398 , n399 , n400 , n401 , n402 , n403 , n404 , n405 , n406 , n407 , n408 , n409 , n410 , n411 , n412 , n413 , n414 , n415 , n416 , n417 , n418 , n419 , n420 , n421 , n422 , n423 , n424 , n425 , n426 , n427 , n428 , n429 , n430 , n431 , n432 , n433 , n434 , n435 , n436 , n437 , n438 , n439 , n440 , n441 , n442 , n443 , n444 , n445 , n446 , n447 , n448 , n449 , n450 , n451 , n452 , n453 , n454 , n455 , n456 , n457 , n458 , n459 , n460 , n461 , n462 , n463 , n464 , n465 , n466 , n467 , n468 , n469 , n470 , n471 , n472 , n473 , n474 , n475 , n476 , n477 , n478 , n479 , n480 , n481 , n482 , n483 , n484 , n485 , n486 , n487 , n488 , n489 , n490 , n491 , n492 , n493 , n494 , n495 , n496 , n497 , n498 , n499 , n500 , n501 , n502 , n503 , n504 , n505 , n506 , n507 , n508 , n509 , n510 , n511 , n512 , n513 , n514 , n515 , n516 , n517 , n518 , n519 , n520 , n521 , n522 , n523 , n524 , n525 , n526 , n527 , n528 , n529 , n530 , n531 , n532 , n533 , n534 , n535 , n536 , n537 , n538 , n539 , n540 , n541 , n542 , n543 , n544 , n545 , n546 , n547 , n548 , n549 , n550 , n551 , n552 , n553 , n554 , n555 , n556 , n557 , n558 , n559 , n560 , n561 , n562 , n563 , n564 , n565 , n566 , n567 , n568 , n569 , n570 , n571 , n572 , n573 , n574 , n575 , n576 , n577 , n578 , n579 , n580 , n581 , n582 , n583 , n584 , n585 , n586 , n587 , n588 , n589 , n590 , n591 , n592 , n593 , n594 , n595 , n596 , n597 , n598 , n599 , n600 , n601 , n602 , n603 , n604 , n605 , n606 , n607 , n608 , n609 , n610 , n611 , n612 , n613 , n614 , n615 , n616 , n617 , n618 , n619 , n620 , n621 , n622 , n623 , n624 , n625 , n626 , n627 , n628 , n629 , n630 , n631 , n632 , n633 , n634 , n635 , n636 , n637 , n638 , n639 , n640 , n641 , n642 , n643 , n644 , n645 , n646 , n647 , n648 , n649 , n650 , n651 , n652 , n653 , n654 , n655 , n656 , n657 , n658 , n659 , n660 , n661 , n662 , n663 , n664 , n665 , n666 , n667 , n668 , n669 , n670 , n671 , n672 , n673 , n674 , n675 , n676 , n677 , n678 , n679 , n680 , n681 , n682 , n683 , n684 , n685 , n686 , n687 , n688 , n689 , n690 , n691 , n692 , n693 , n694 , n695 , n696 , n697 , n698 , n699 , n700 , n701 , n702 , n703 , n704 , n705 , n706 , n707 , n708 , n709 , n710 , n711 , n712 , n713 , n714 , n715 , n716 , n717 , n718 , n719 , n720 , n721 , n722 , n723 , n724 , n725 , n726 , n727 , n728 , n729 , n730 , n731 , n732 , n733 , n734 , n735 , n736 , n737 , n738 , n739 , n740 , n741 , n742 , n743 , n744 , n745 , n746 , n747 , n748 , n749 , n750 , n751 , n752 , n753 , n754 , n755 , n756 , n757 , n758 , n759 , n760 , n761 , n762 , n763 , n764 , n765 , n766 , n767 , n768 , n769 , n770 , n771 , n772 , n773 , n774 , n775 , n776 , n777 , n778 , n779 , n780 , n781 , n782 , n783 , n784 , n785 , n786 , n787 , n788 , n789 , n790 , n791 , n792 , n793 , n794 , n795 , n796 , n797 , n798 , n799 , n800 , n801 , n802 , n803 , n804 , n805 , n806 , n807 , n808 , n809 , n810 , n811 , n812 , n813 , n814 , n815 , n816 , n817 , n818 , n819 , n820 , n821 , n822 , n823 , n824 , n825 , n826 , n827 , n828 , n829 , n830 , n831 , n832 , n833 , n834 , n835 , n836 , n837 , n838 , n839 , n840 , n841 , n842 , n843 , n844 , n845 , n846 , n847 , n848 , n849 , n850 , n851 , n852 , n853 , n854 , n855 , n856 , n857 , n858 , n859 , n860 , n861 , n862 , n863 , n864 , n865 , n866 , n867 , n868 , n869 , n870 , n871 , n872 , n873 , n874 , n875 , n876 , n877 , n878 , n879 , n880 , n881 , n882 , n883 , n884 , n885 , n886 , n887 , n888 , n889 , n890 , n891 , n892 , n893 , n894 , n895 , n896 , n897 , n898 , n899 , n900 , n901 , n902 , n903 , n904 , n905 , n906 , n907 , n908 , n909 , n910 , n911 , n912 , n913 , n914 , n915 , n916 , n917 , n918 , n919 , n920 , n921 , n922 , n923 , n924 , n925 , n926 , n927 , n928 , n929 , n930 , n931 , n932 , n933 , n934 , n935 , n936 , n937 , n938 , n939 , n940 , n941 , n942 , n943 , n944 , n945 , n946 , n947 , n948 , n949 , n950 , n951 , n952 , n953 , n954 , n955 , n956 , n957 , n958 , n959 , n960 , n961 , n962 , n963 , n964 , n965 , n966 , n967 , n968 , n969 , n970 , n971 , n972 , n973 , n974 , n975 , n976 , n977 , n978 , n979 , n980 , n981 , n982 , n983 , n984 , n985 , n986 , n987 , n988 , n989 , n990 , n991 , n992 , n993 , n994 , n995 , n996 , n997 , n998 , n999 , n1000 , n1001 , n1002 , n1003 , n1004 , n1005 , n1006 , n1007 , n1008 , n1009 , n1010 , n1011 , n1012 , n1013 , n1014 , n1015 , n1016 , n1017 , n1018 , n1019 , n1020 , n1021 , n1022 , n1023 , n1024 , n1025 , n1026 , n1027 , n1028 , n1029 , n1030 , n1031 , n1032 , n1033 , n1034 , n1035 , n1036 , n1037 , n1038 , n1039 , n1040 , n1041 , n1042 , n1043 , n1044 , n1045 , n1046 , n1047 , n1048 , n1049 , n1050 , n1051 , n1052 , n1053 , n1054 , n1055 , n1056 , n1057 , n1058 , n1059 , n1060 , n1061 , n1062 , n1063 , n1064 , n1065 , n1066 , n1067 , n1068 , n1069 , n1070 , n1071 , n1072 , n1073 , n1074 , n1075 , n1076 , n1077 , n1078 , n1079 , n1080 , n1081 , n1082 , n1083 , n1084 , n1085 , n1086 , n1087 , n1088 , n1089 , n1090 , n1091 , n1092 , n1093 , n1094 , n1095 , n1096 , n1097 , n1098 , n1099 , n1100 , n1101 , n1102 , n1103 , n1104 , n1105 , n1106 , n1107 , n1108 , n1109 , n1110 , n1111 , n1112 , n1113 , n1114 , n1115 , n1116 , n1117 , n1118 , n1119 , n1120 , n1121 , n1122 , n1123 , n1124 , n1125 , n1126 , n1127 , n1128 , n1129 , n1130 , n1131 , n1132 , n1133 , n1134 , n1135 , n1136 , n1137 , n1138 , n1139 , n1140 , n1141 , n1142 , n1143 , n1144 , n1145 , n1146 , n1147 , n1148 , n1149 , n1150 , n1151 , n1152 , n1153 , n1154 , n1155 , n1156 , n1157 , n1158 , n1159 , n1160 , n1161 , n1162 , n1163 , n1164 , n1165 , n1166 , n1167 , n1168 , n1169 , n1170 , n1171 , n1172 , n1173 , n1174 , n1175 , n1176 , n1177 , n1178 , n1179 , n1180 , n1181 , n1182 , n1183 , n1184 , n1185 , n1186 , n1187 , n1188 , n1189 , n1190 , n1191 , n1192 , n1193 , n1194 , n1195 , n1196 , n1197 , n1198 , n1199 , n1200 , n1201 , n1202 , n1203 , n1204 , n1205 , n1206 , n1207 , n1208 , n1209 , n1210 , n1211 , n1212 , n1213 , n1214 , n1215 , n1216 , n1217 , n1218 , n1219 , n1220 , n1221 , n1222 , n1223 , n1224 , n1225 , n1226 , n1227 , n1228 , n1229 , n1230 , n1231 , n1232 , n1233 , n1234 , n1235 , n1236 , n1237 , n1238 , n1239 , n1240 , n1241 , n1242 , n1243 , n1244 , n1245 , n1246 , n1247 , n1248 , n1249 , n1250 , n1251 , n1252 , n1253 , n1254 , n1255 , n1256 , n1257 , n1258 , n1259 , n1260 , n1261 , n1262 , n1263 , n1264 , n1265 , n1266 , n1267 , n1268 , n1269 , n1270 , n1271 , n1272 , n1273 , n1274 , n1275 , n1276 , n1277 , n1278 , n1279 , n1280 , n1281 , n1282 , n1283 , n1284 , n1285 , n1286 , n1287 , n1288 , n1289 , n1290 , n1291 , n1292 , n1293 , n1294 , n1295 , n1296 , n1297 , n1298 , n1299 , n1300 , n1301 , n1302 , n1303 , n1304 , n1305 , n1306 , n1307 , n1308 , n1309 , n1310 , n1311 , n1312 , n1313 , n1314 , n1315 , n1316 , n1317 , n1318 , n1319 , n1320 , n1321 , n1322 , n1323 , n1324 , n1325 , n1326 , n1327 , n1328 , n1329 , n1330 , n1331 , n1332 , n1333 , n1334 , n1335 , n1336 , n1337 , n1338 , n1339 , n1340 , n1341 , n1342 , n1343 , n1344 , n1345 , n1346 , n1347 , n1348 , n1349 , n1350 , n1351 , n1352 , n1353 , n1354 , n1355 , n1356 , n1357 , n1358 , n1359 , n1360 , n1361 , n1362 , n1363 , n1364 , n1365 , n1366 , n1367 , n1368 , n1369 , n1370 , n1371 , n1372 , n1373 , n1374 , n1375 , n1376 , n1377 , n1378 , n1379 , n1380 , n1381 , n1382 , n1383 , n1384 , n1385 , n1386 , n1387 , n1388 , n1389 , n1390 , n1391 , n1392 , n1393 , n1394 , n1395 , n1396 , n1397 , n1398 , n1399 , n1400 , n1401 , n1402 , n1403 , n1404 , n1405 , n1406 , n1407 , n1408 , n1409 , n1410 , n1411 , n1412 , n1413 , n1414 , n1415 , n1416 , n1417 , n1418 , n1419 , n1420 , n1421 , n1422 , n1423 , n1424 , n1425 , n1426 , n1427 , n1428 , n1429 , n1430 , n1431 , n1432 , n1433 , n1434 , n1435 , n1436 , n1437 , n1438 , n1439 , n1440 , n1441 , n1442 , n1443 , n1444 , n1445 , n1446 , n1447 , n1448 , n1449 , n1450 , n1451 , n1452 , n1453 , n1454 , n1455 , n1456 , n1457 , n1458 , n1459 , n1460 , n1461 , n1462 , n1463 , n1464 , n1465 , n1466 , n1467 , n1468 , n1469 , n1470 , n1471 , n1472 , n1473 , n1474 , n1475 , n1476 , n1477 , n1478 , n1479 , n1480 , n1481 , n1482 , n1483 , n1484 , n1485 , n1486 , n1487 , n1488 , n1489 , n1490 , n1491 , n1492 , n1493 , n1494 , n1495 , n1496 , n1497 , n1498 , n1499 , n1500 , n1501 , n1502 , n1503 , n1504 , n1505 , n1506 , n1507 , n1508 , n1509 , n1510 , n1511 , n1512 , n1513 , n1514 , n1515 , n1516 , n1517 , n1518 , n1519 , n1520 , n1521 , n1522 , n1523 , n1524 , n1525 , n1526 , n1527 , n1528 , n1529 , n1530 , n1531 , n1532 , n1533 , n1534 , n1535 , n1536 , n1537 , n1538 , n1539 , n1540 , n1541 , n1542 , n1543 , n1544 , n1545 , n1546 , n1547 , n1548 , n1549 , n1550 , n1551 , n1552 , n1553 , n1554 , n1555 , n1556 , n1557 , n1558 , n1559 , n1560 , n1561 , n1562 , n1563 , n1564 , n1565 , n1566 , n1567 , n1568 , n1569 , n1570 , n1571 , n1572 , n1573 , n1574 , n1575 , n1576 , n1577 , n1578 , n1579 , n1580 , n1581 , n1582 , n1583 , n1584 , n1585 , n1586 , n1587 , n1588 , n1589 , n1590 , n1591 , n1592 , n1593 , n1594 , n1595 , n1596 , n1597 , n1598 , n1599 , n1600 , n1601 , n1602 , n1603 , n1604 , n1605 , n1606 , n1607 , n1608 , n1609 , n1610 , n1611 , n1612 , n1613 , n1614 , n1615 , n1616 , n1617 , n1618 , n1619 , n1620 , n1621 , n1622 , n1623 , n1624 , n1625 , n1626 , n1627 , n1628 , n1629 , n1630 , n1631 , n1632 , n1633 , n1634 , n1635 , n1636 , n1637 , n1638 , n1639 , n1640 , n1641 , n1642 , n1643 , n1644 , n1645 , n1646 , n1647 , n1648 , n1649 , n1650 , n1651 , n1652 , n1653 , n1654 , n1655 , n1656 , n1657 , n1658 , n1659 , n1660 , n1661 , n1662 , n1663 , n1664 , n1665 , n1666 , n1667 , n1668 , n1669 , n1670 , n1671 , n1672 , n1673 , n1674 , n1675 , n1676 , n1677 , n1678 , n1679 , n1680 , n1681 , n1682 , n1683 , n1684 , n1685 , n1686 , n1687 , n1688 , n1689 , n1690 , n1691 , n1692 , n1693 , n1694 , n1695 , n1696 , n1697 , n1698 , n1699 , n1700 , n1701 , n1702 , n1703 , n1704 , n1705 , n1706 , n1707 , n1708 , n1709 , n1710 , n1711 , n1712 , n1713 , n1714 , n1715 , n1716 , n1717 , n1718 , n1719 , n1720 , n1721 , n1722 , n1723 , n1724 , n1725 , n1726 , n1727 , n1728 , n1729 , n1730 , n1731 , n1732 , n1733 , n1734 , n1735 , n1736 , n1737 , n1738 , n1739 , n1740 , n1741 , n1742 , n1743 , n1744 , n1745 , n1746 , n1747 , n1748 , n1749 , n1750 , n1751 , n1752 , n1753 , n1754 , n1755 , n1756 , n1757 , n1758 , n1759 , n1760 , n1761 , n1762 , n1763 , n1764 , n1765 , n1766 , n1767 , n1768 , n1769 , n1770 , n1771 , n1772 , n1773 , n1774 , n1775 , n1776 , n1777 , n1778 , n1779 , n1780 , n1781 , n1782 , n1783 , n1784 , n1785 , n1786 , n1787 , n1788 , n1789 , n1790 , n1791 , n1792 , n1793 , n1794 , n1795 , n1796 , n1797 , n1798 , n1799 , n1800 , n1801 , n1802 , n1803 , n1804 , n1805 , n1806 , n1807 , n1808 , n1809 , n1810 , n1811 , n1812 , n1813 , n1814 , n1815 , n1816 , n1817 , n1818 , n1819 , n1820 , n1821 , n1822 , n1823 , n1824 , n1825 , n1826 , n1827 , n1828 , n1829 , n1830 , n1831 , n1832 , n1833 , n1834 , n1835 , n1836 , n1837 , n1838 , n1839 , n1840 , n1841 , n1842 , n1843 , n1844 , n1845 , n1846 , n1847 , n1848 , n1849 , n1850 , n1851 , n1852 , n1853 , n1854 , n1855 , n1856 , n1857 , n1858 , n1859 , n1860 , n1861 , n1862 , n1863 , n1864 , n1865 , n1866 , n1867 , n1868 , n1869 , n1870 , n1871 , n1872 , n1873 , n1874 , n1875 , n1876 , n1877 , n1878 , n1879 , n1880 , n1881 , n1882 , n1883 , n1884 , n1885 , n1886 , n1887 , n1888 , n1889 , n1890 , n1891 , n1892 , n1893 , n1894 , n1895 , n1896 , n1897 , n1898 , n1899 , n1900 , n1901 , n1902 , n1903 , n1904 , n1905 , n1906 , n1907 , n1908 , n1909 , n1910 , n1911 , n1912 , n1913 , n1914 , n1915 , n1916 , n1917 , n1918 , n1919 , n1920 , n1921 , n1922 , n1923 , n1924 , n1925 , n1926 , n1927 , n1928 , n1929 , n1930 , n1931 , n1932 , n1933 , n1934 , n1935 , n1936 , n1937 , n1938 , n1939 , n1940 , n1941 , n1942 , n1943 , n1944 , n1945 , n1946 , n1947 , n1948 , n1949 , n1950 , n1951 , n1952 , n1953 , n1954 , n1955 , n1956 , n1957 , n1958 , n1959 , n1960 , n1961 , n1962 , n1963 , n1964 , n1965 , n1966 , n1967 , n1968 , n1969 , n1970 , n1971 , n1972 , n1973 , n1974 , n1975 , n1976 , n1977 , n1978 , n1979 , n1980 , n1981 , n1982 , n1983 , n1984 , n1985 , n1986 , n1987 , n1988 , n1989 , n1990 , n1991 , n1992 , n1993 , n1994 , n1995 , n1996 , n1997 , n1998 , n1999 , n2000 , n2001 , n2002 , n2003 , n2004 , n2005 , n2006 , n2007 , n2008 , n2009 , n2010 , n2011 , n2012 , n2013 , n2014 , n2015 , n2016 , n2017 , n2018 , n2019 , n2020 , n2021 , n2022 , n2023 , n2024 , n2025 , n2026 , n2027 , n2028 , n2029 , n2030 , n2031 , n2032 , n2033 , n2034 , n2035 , n2036 , n2037 , n2038 , n2039 , n2040 , n2041 , n2042 , n2043 , n2044 , n2045 , n2046 , n2047 , n2048 , n2049 , n2050 , n2051 , n2052 , n2053 , n2054 , n2055 , n2056 , n2057 , n2058 , n2059 , n2060 , n2061 , n2062 , n2063 , n2064 , n2065 , n2066 , n2067 , n2068 , n2069 , n2070 , n2071 , n2072 , n2073 , n2074 , n2075 , n2076 , n2077 , n2078 , n2079 , n2080 , n2081 , n2082 , n2083 , n2084 , n2085 , n2086 , n2087 , n2088 , n2089 , n2090 , n2091 , n2092 , n2093 , n2094 , n2095 , n2096 , n2097 , n2098 , n2099 , n2100 , n2101 , n2102 , n2103 , n2104 , n2105 , n2106 , n2107 , n2108 , n2109 , n2110 , n2111 , n2112 , n2113 , n2114 , n2115 , n2116 , n2117 , n2118 , n2119 , n2120 , n2121 , n2122 , n2123 , n2124 , n2125 , n2126 , n2127 , n2128 , n2129 , n2130 , n2131 , n2132 , n2133 , n2134 , n2135 , n2136 , n2137 , n2138 , n2139 , n2140 , n2141 , n2142 , n2143 , n2144 , n2145 , n2146 , n2147 , n2148 , n2149 , n2150 , n2151 , n2152 , n2153 , n2154 , n2155 , n2156 , n2157 , n2158 , n2159 , n2160 , n2161 , n2162 , n2163 , n2164 , n2165 , n2166 , n2167 , n2168 , n2169 , n2170 , n2171 , n2172 , n2173 , n2174 , n2175 , n2176 , n2177 , n2178 , n2179 , n2180 , n2181 , n2182 , n2183 , n2184 , n2185 , n2186 , n2187 , n2188 , n2189 , n2190 , n2191 , n2192 , n2193 , n2194 , n2195 , n2196 , n2197 , n2198 , n2199 , n2200 , n2201 , n2202 , n2203 , n2204 , n2205 , n2206 , n2207 , n2208 , n2209 , n2210 , n2211 , n2212 , n2213 , n2214 , n2215 , n2216 , n2217 , n2218 , n2219 , n2220 , n2221 , n2222 , n2223 , n2224 , n2225 , n2226 , n2227 , n2228 , n2229 , n2230 , n2231 , n2232 , n2233 , n2234 , n2235 , n2236 , n2237 , n2238 , n2239 , n2240 , n2241 , n2242 , n2243 , n2244 , n2245 , n2246 , n2247 , n2248 , n2249 , n2250 , n2251 , n2252 , n2253 , n2254 , n2255 , n2256 , n2257 , n2258 , n2259 , n2260 , n2261 , n2262 , n2263 , n2264 , n2265 , n2266 , n2267 , n2268 , n2269 , n2270 , n2271 , n2272 , n2273 , n2274 , n2275 , n2276 , n2277 , n2278 , n2279 , n2280 , n2281 , n2282 , n2283 , n2284 , n2285 , n2286 , n2287 , n2288 , n2289 , n2290 , n2291 , n2292 , n2293 , n2294 , n2295 , n2296 , n2297 , n2298 , n2299 , n2300 , n2301 , n2302 , n2303 , n2304 , n2305 , n2306 , n2307 , n2308 , n2309 , n2310 , n2311 , n2312 , n2313 , n2314 , n2315 , n2316 , n2317 , n2318 , n2319 , n2320 , n2321 , n2322 , n2323 , n2324 , n2325 , n2326 , n2327 , n2328 , n2329 , n2330 , n2331 , n2332 , n2333 , n2334 , n2335 , n2336 , n2337 , n2338 , n2339 , n2340 , n2341 , n2342 , n2343 , n2344 , n2345 , n2346 , n2347 , n2348 , n2349 , n2350 , n2351 , n2352 , n2353 , n2354 , n2355 , n2356 , n2357 , n2358 , n2359 , n2360 , n2361 , n2362 , n2363 , n2364 , n2365 , n2366 , n2367 , n2368 , n2369 , n2370 , n2371 , n2372 , n2373 , n2374 , n2375 , n2376 , n2377 , n2378 , n2379 , n2380 , n2381 , n2382 , n2383 , n2384 , n2385 , n2386 , n2387 , n2388 , n2389 , n2390 , n2391 , n2392 , n2393 , n2394 , n2395 , n2396 , n2397 , n2398 , n2399 , n2400 , n2401 , n2402 , n2403 , n2404 , n2405 , n2406 , n2407 , n2408 , n2409 , n2410 , n2411 , n2412 , n2413 , n2414 , n2415 , n2416 , n2417 , n2418 , n2419 , n2420 , n2421 , n2422 , n2423 , n2424 , n2425 , n2426 , n2427 , n2428 , n2429 , n2430 , n2431 , n2432 , n2433 , n2434 , n2435 , n2436 , n2437 , n2438 , n2439 , n2440 , n2441 , n2442 , n2443 , n2444 , n2445 , n2446 , n2447 , n2448 , n2449 , n2450 , n2451 , n2452 , n2453 , n2454 , n2455 , n2456 , n2457 , n2458 , n2459 , n2460 , n2461 , n2462 , n2463 , n2464 , n2465 , n2466 , n2467 , n2468 , n2469 , n2470 , n2471 , n2472 , n2473 , n2474 , n2475 , n2476 , n2477 , n2478 , n2479 , n2480 , n2481 , n2482 , n2483 , n2484 , n2485 , n2486 , n2487 , n2488 , n2489 , n2490 , n2491 , n2492 , n2493 , n2494 , n2495 , n2496 , n2497 , n2498 , n2499 , n2500 , n2501 , n2502 , n2503 , n2504 , n2505 , n2506 , n2507 , n2508 , n2509 , n2510 , n2511 , n2512 , n2513 , n2514 , n2515 , n2516 , n2517 , n2518 , n2519 , n2520 , n2521 , n2522 , n2523 , n2524 , n2525 , n2526 , n2527 , n2528 , n2529 , n2530 , n2531 , n2532 , n2533 , n2534 , n2535 , n2536 , n2537 , n2538 , n2539 , n2540 , n2541 , n2542 , n2543 , n2544 , n2545 , n2546 , n2547 , n2548 , n2549 , n2550 , n2551 , n2552 , n2553 , n2554 , n2555 , n2556 , n2557 , n2558 , n2559 , n2560 , n2561 , n2562 , n2563 , n2564 , n2565 , n2566 , n2567 , n2568 , n2569 , n2570 , n2571 , n2572 , n2573 , n2574 , n2575 , n2576 , n2577 , n2578 , n2579 , n2580 , n2581 , n2582 , n2583 , n2584 , n2585 , n2586 , n2587 , n2588 , n2589 , n2590 , n2591 , n2592 , n2593 , n2594 , n2595 , n2596 , n2597 , n2598 , n2599 , n2600 , n2601 , n2602 , n2603 , n2604 , n2605 , n2606 , n2607 , n2608 , n2609 , n2610 , n2611 , n2612 , n2613 , n2614 , n2615 , n2616 , n2617 , n2618 , n2619 , n2620 , n2621 , n2622 , n2623 , n2624 , n2625 , n2626 , n2627 , n2628 , n2629 , n2630 , n2631 , n2632 , n2633 , n2634 , n2635 , n2636 , n2637 , n2638 , n2639 , n2640 , n2641 , n2642 , n2643 , n2644 , n2645 , n2646 , n2647 , n2648 , n2649 , n2650 , n2651 , n2652 , n2653 , n2654 , n2655 , n2656 , n2657 , n2658 , n2659 , n2660 , n2661 , n2662 , n2663 , n2664 , n2665 , n2666 , n2667 , n2668 , n2669 , n2670 , n2671 , n2672 , n2673 , n2674 , n2675 , n2676 , n2677 , n2678 , n2679 , n2680 , n2681 , n2682 , n2683 , n2684 , n2685 , n2686 , n2687 , n2688 , n2689 , n2690 , n2691 , n2692 , n2693 , n2694 , n2695 , n2696 , n2697 , n2698 , n2699 , n2700 , n2701 , n2702 , n2703 , n2704 , n2705 , n2706 , n2707 , n2708 , n2709 , n2710 , n2711 , n2712 , n2713 , n2714 , n2715 , n2716 , n2717 , n2718 , n2719 , n2720 , n2721 , n2722 , n2723 , n2724 , n2725 , n2726 , n2727 , n2728 , n2729 , n2730 , n2731 , n2732 , n2733 , n2734 , n2735 , n2736 , n2737 , n2738 , n2739 , n2740 , n2741 , n2742 , n2743 , n2744 , n2745 , n2746 , n2747 , n2748 , n2749 , n2750 , n2751 , n2752 , n2753 , n2754 , n2755 , n2756 , n2757 , n2758 , n2759 , n2760 , n2761 , n2762 , n2763 , n2764 , n2765 , n2766 , n2767 , n2768 , n2769 , n2770 , n2771 , n2772 , n2773 , n2774 , n2775 , n2776 , n2777 , n2778 , n2779 , n2780 , n2781 , n2782 , n2783 , n2784 , n2785 , n2786 , n2787 , n2788 , n2789 , n2790 , n2791 , n2792 , n2793 , n2794 , n2795 , n2796 , n2797 , n2798 , n2799 , n2800 , n2801 , n2802 , n2803 , n2804 , n2805 , n2806 , n2807 , n2808 , n2809 , n2810 , n2811 , n2812 , n2813 , n2814 , n2815 , n2816 , n2817 , n2818 , n2819 , n2820 , n2821 , n2822 , n2823 , n2824 , n2825 , n2826 , n2827 , n2828 , n2829 , n2830 , n2831 , n2832 , n2833 , n2834 , n2835 , n2836 , n2837 , n2838 , n2839 , n2840 , n2841 , n2842 , n2843 , n2844 , n2845 , n2846 , n2847 , n2848 , n2849 , n2850 , n2851 , n2852 , n2853 , n2854 , n2855 , n2856 , n2857 , n2858 , n2859 , n2860 , n2861 , n2862 , n2863 , n2864 , n2865 , n2866 , n2867 , n2868 , n2869 , n2870 , n2871 , n2872 , n2873 , n2874 , n2875 , n2876 , n2877 , n2878 , n2879 , n2880 , n2881 , n2882 , n2883 , n2884 , n2885 , n2886 , n2887 , n2888 , n2889 , n2890 , n2891 , n2892 , n2893 , n2894 , n2895 , n2896 , n2897 , n2898 , n2899 , n2900 , n2901 , n2902 , n2903 , n2904 , n2905 , n2906 , n2907 , n2908 , n2909 , n2910 , n2911 , n2912 , n2913 , n2914 , n2915 , n2916 , n2917 , n2918 , n2919 , n2920 , n2921 , n2922 , n2923 , n2924 , n2925 , n2926 , n2927 , n2928 , n2929 , n2930 , n2931 , n2932 , n2933 , n2934 , n2935 , n2936 , n2937 , n2938 , n2939 , n2940 , n2941 , n2942 , n2943 , n2944 , n2945 , n2946 , n2947 , n2948 , n2949 , n2950 , n2951 , n2952 , n2953 , n2954 , n2955 , n2956 , n2957 , n2958 , n2959 , n2960 , n2961 , n2962 , n2963 , n2964 , n2965 , n2966 , n2967 , n2968 , n2969 , n2970 , n2971 , n2972 , n2973 , n2974 , n2975 , n2976 , n2977 , n2978 , n2979 , n2980 , n2981 , n2982 , n2983 , n2984 , n2985 , n2986 , n2987 , n2988 , n2989 , n2990 , n2991 , n2992 , n2993 , n2994 , n2995 , n2996 , n2997 , n2998 , n2999 , n3000 , n3001 , n3002 , n3003 , n3004 , n3005 , n3006 , n3007 , n3008 , n3009 , n3010 , n3011 , n3012 , n3013 , n3014 , n3015 , n3016 , n3017 , n3018 , n3019 , n3020 , n3021 , n3022 , n3023 , n3024 , n3025 , n3026 , n3027 , n3028 , n3029 , n3030 , n3031 , n3032 , n3033 , n3034 , n3035 , n3036 , n3037 , n3038 , n3039 , n3040 , n3041 , n3042 , n3043 , n3044 , n3045 , n3046 , n3047 , n3048 , n3049 , n3050 , n3051 , n3052 , n3053 , n3054 , n3055 , n3056 , n3057 , n3058 , n3059 , n3060 , n3061 , n3062 , n3063 , n3064 , n3065 , n3066 , n3067 , n3068 , n3069 , n3070 , n3071 , n3072 , n3073 , n3074 , n3075 , n3076 , n3077 , n3078 , n3079 , n3080 , n3081 , n3082 , n3083 , n3084 , n3085 , n3086 , n3087 , n3088 , n3089 , n3090 , n3091 , n3092 , n3093 , n3094 , n3095 , n3096 , n3097 , n3098 , n3099 , n3100 , n3101 , n3102 , n3103 , n3104 , n3105 , n3106 , n3107 , n3108 , n3109 , n3110 , n3111 , n3112 , n3113 , n3114 , n3115 , n3116 , n3117 , n3118 , n3119 , n3120 , n3121 , n3122 , n3123 , n3124 , n3125 , n3126 , n3127 , n3128 , n3129 , n3130 , n3131 , n3132 , n3133 , n3134 , n3135 , n3136 , n3137 , n3138 , n3139 , n3140 , n3141 , n3142 , n3143 , n3144 , n3145 , n3146 , n3147 , n3148 , n3149 , n3150 , n3151 , n3152 , n3153 , n3154 , n3155 , n3156 , n3157 , n3158 , n3159 , n3160 , n3161 , n3162 , n3163 , n3164 , n3165 , n3166 , n3167 , n3168 , n3169 , n3170 , n3171 , n3172 , n3173 , n3174 , n3175 , n3176 , n3177 , n3178 , n3179 , n3180 , n3181 , n3182 , n3183 , n3184 , n3185 , n3186 , n3187 , n3188 , n3189 , n3190 , n3191 , n3192 , n3193 , n3194 , n3195 , n3196 , n3197 , n3198 , n3199 , n3200 , n3201 , n3202 , n3203 , n3204 , n3205 , n3206 , n3207 , n3208 , n3209 , n3210 , n3211 , n3212 , n3213 , n3214 , n3215 , n3216 , n3217 , n3218 , n3219 , n3220 , n3221 , n3222 , n3223 , n3224 , n3225 , n3226 , n3227 , n3228 , n3229 , n3230 , n3231 , n3232 , n3233 , n3234 , n3235 , n3236 , n3237 , n3238 , n3239 , n3240 , n3241 , n3242 , n3243 , n3244 , n3245 , n3246 , n3247 , n3248 , n3249 , n3250 , n3251 , n3252 , n3253 , n3254 , n3255 , n3256 , n3257 , n3258 , n3259 , n3260 , n3261 , n3262 , n3263 , n3264 , n3265 , n3266 , n3267 , n3268 , n3269 , n3270 , n3271 , n3272 , n3273 , n3274 , n3275 , n3276 , n3277 , n3278 , n3279 , n3280 , n3281 , n3282 , n3283 , n3284 , n3285 , n3286 , n3287 , n3288 , n3289 , n3290 , n3291 , n3292 , n3293 , n3294 , n3295 , n3296 , n3297 , n3298 , n3299 , n3300 , n3301 , n3302 , n3303 , n3304 , n3305 , n3306 , n3307 , n3308 , n3309 , n3310 , n3311 , n3312 , n3313 , n3314 , n3315 , n3316 , n3317 , n3318 , n3319 , n3320 , n3321 , n3322 , n3323 , n3324 , n3325 , n3326 , n3327 , n3328 , n3329 , n3330 , n3331 , n3332 , n3333 , n3334 , n3335 , n3336 , n3337 , n3338 , n3339 , n3340 , n3341 , n3342 , n3343 , n3344 , n3345 , n3346 , n3347 , n3348 , n3349 , n3350 , n3351 , n3352 , n3353 , n3354 , n3355 , n3356 , n3357 , n3358 , n3359 , n3360 , n3361 , n3362 , n3363 , n3364 , n3365 , n3366 , n3367 , n3368 , n3369 , n3370 , n3371 , n3372 , n3373 , n3374 , n3375 , n3376 , n3377 , n3378 , n3379 , n3380 , n3381 , n3382 , n3383 , n3384 , n3385 , n3386 , n3387 , n3388 , n3389 , n3390 , n3391 , n3392 , n3393 , n3394 , n3395 , n3396 , n3397 , n3398 , n3399 , n3400 , n3401 , n3402 , n3403 , n3404 , n3405 , n3406 , n3407 , n3408 , n3409 , n3410 , n3411 , n3412 , n3413 , n3414 , n3415 , n3416 , n3417 , n3418 , n3419 , n3420 , n3421 , n3422 , n3423 , n3424 , n3425 , n3426 , n3427 , n3428 , n3429 , n3430 , n3431 , n3432 , n3433 , n3434 , n3435 , n3436 , n3437 , n3438 , n3439 , n3440 , n3441 , n3442 , n3443 , n3444 , n3445 , n3446 , n3447 , n3448 , n3449 , n3450 , n3451 , n3452 , n3453 , n3454 , n3455 , n3456 , n3457 , n3458 , n3459 , n3460 , n3461 , n3462 , n3463 , n3464 , n3465 , n3466 , n3467 , n3468 , n3469 , n3470 , n3471 , n3472 , n3473 , n3474 , n3475 , n3476 , n3477 , n3478 , n3479 , n3480 , n3481 , n3482 , n3483 , n3484 , n3485 , n3486 , n3487 , n3488 , n3489 , n3490 , n3491 , n3492 , n3493 , n3494 , n3495 , n3496 , n3497 , n3498 , n3499 , n3500 , n3501 , n3502 , n3503 , n3504 , n3505 , n3506 , n3507 , n3508 , n3509 , n3510 , n3511 , n3512 , n3513 , n3514 , n3515 , n3516 , n3517 , n3518 , n3519 , n3520 , n3521 , n3522 , n3523 , n3524 , n3525 , n3526 , n3527 , n3528 , n3529 , n3530 , n3531 , n3532 , n3533 , n3534 , n3535 , n3536 , n3537 , n3538 , n3539 , n3540 , n3541 , n3542 , n3543 , n3544 , n3545 , n3546 , n3547 , n3548 , n3549 , n3550 , n3551 , n3552 , n3553 , n3554 , n3555 , n3556 , n3557 , n3558 , n3559 , n3560 , n3561 , n3562 , n3563 , n3564 , n3565 , n3566 , n3567 , n3568 , n3569 , n3570 , n3571 , n3572 , n3573 , n3574 , n3575 , n3576 , n3577 , n3578 , n3579 , n3580 , n3581 , n3582 , n3583 , n3584 , n3585 , n3586 , n3587 , n3588 , n3589 , n3590 , n3591 , n3592 , n3593 , n3594 , n3595 , n3596 , n3597 , n3598 , n3599 , n3600 , n3601 , n3602 , n3603 , n3604 , n3605 , n3606 , n3607 , n3608 , n3609 , n3610 , n3611 , n3612 , n3613 , n3614 , n3615 , n3616 , n3617 , n3618 , n3619 , n3620 , n3621 , n3622 , n3623 , n3624 , n3625 , n3626 , n3627 , n3628 , n3629 , n3630 , n3631 , n3632 , n3633 , n3634 , n3635 , n3636 , n3637 , n3638 , n3639 , n3640 , n3641 , n3642 , n3643 , n3644 , n3645 , n3646 , n3647 , n3648 , n3649 , n3650 , n3651 , n3652 , n3653 , n3654 , n3655 , n3656 , n3657 , n3658 , n3659 , n3660 , n3661 , n3662 , n3663 , n3664 , n3665 , n3666 , n3667 , n3668 , n3669 , n3670 , n3671 , n3672 , n3673 , n3674 , n3675 , n3676 , n3677 , n3678 , n3679 , n3680 , n3681 , n3682 , n3683 , n3684 , n3685 , n3686 , n3687 , n3688 , n3689 , n3690 , n3691 , n3692 , n3693 , n3694 , n3695 , n3696 , n3697 , n3698 , n3699 , n3700 , n3701 , n3702 , n3703 , n3704 , n3705 , n3706 , n3707 , n3708 , n3709 , n3710 , n3711 , n3712 , n3713 , n3714 , n3715 , n3716 , n3717 , n3718 , n3719 , n3720 , n3721 , n3722 , n3723 , n3724 , n3725 , n3726 , n3727 , n3728 , n3729 , n3730 , n3731 , n3732 , n3733 , n3734 , n3735 , n3736 , n3737 , n3738 , n3739 , n3740 , n3741 , n3742 , n3743 , n3744 , n3745 , n3746 , n3747 , n3748 , n3749 , n3750 , n3751 , n3752 , n3753 , n3754 , n3755 , n3756 , n3757 , n3758 , n3759 , n3760 , n3761 , n3762 , n3763 , n3764 , n3765 , n3766 , n3767 , n3768 , n3769 , n3770 , n3771 , n3772 , n3773 , n3774 , n3775 , n3776 , n3777 , n3778 , n3779 , n3780 , n3781 , n3782 , n3783 , n3784 , n3785 , n3786 , n3787 , n3788 , n3789 , n3790 , n3791 , n3792 , n3793 , n3794 , n3795 , n3796 , n3797 , n3798 , n3799 , n3800 , n3801 , n3802 , n3803 , n3804 , n3805 , n3806 , n3807 , n3808 , n3809 , n3810 , n3811 , n3812 , n3813 , n3814 , n3815 , n3816 , n3817 , n3818 , n3819 , n3820 , n3821 , n3822 , n3823 , n3824 , n3825 , n3826 , n3827 , n3828 , n3829 , n3830 , n3831 , n3832 , n3833 , n3834 , n3835 , n3836 , n3837 , n3838 , n3839 , n3840 , n3841 , n3842 , n3843 , n3844 , n3845 , n3846 , n3847 , n3848 , n3849 , n3850 , n3851 , n3852 , n3853 , n3854 , n3855 , n3856 , n3857 , n3858 , n3859 , n3860 , n3861 , n3862 , n3863 , n3864 , n3865 , n3866 , n3867 , n3868 , n3869 , n3870 , n3871 , n3872 , n3873 , n3874 , n3875 , n3876 , n3877 , n3878 , n3879 , n3880 , n3881 , n3882 , n3883 , n3884 , n3885 , n3886 , n3887 , n3888 , n3889 , n3890 , n3891 , n3892 , n3893 , n3894 , n3895 , n3896 , n3897 , n3898 , n3899 , n3900 , n3901 , n3902 , n3903 , n3904 , n3905 , n3906 , n3907 , n3908 , n3909 , n3910 , n3911 , n3912 , n3913 , n3914 , n3915 , n3916 , n3917 , n3918 , n3919 , n3920 , n3921 , n3922 , n3923 , n3924 , n3925 , n3926 , n3927 , n3928 , n3929 , n3930 , n3931 , n3932 , n3933 , n3934 , n3935 , n3936 , n3937 , n3938 , n3939 , n3940 , n3941 , n3942 , n3943 , n3944 , n3945 , n3946 , n3947 , n3948 , n3949 , n3950 , n3951 , n3952 , n3953 , n3954 , n3955 , n3956 , n3957 , n3958 , n3959 , n3960 , n3961 , n3962 , n3963 , n3964 , n3965 , n3966 , n3967 , n3968 , n3969 , n3970 , n3971 , n3972 , n3973 , n3974 , n3975 , n3976 , n3977 , n3978 , n3979 , n3980 , n3981 , n3982 , n3983 , n3984 , n3985 , n3986 , n3987 , n3988 , n3989 , n3990 , n3991 , n3992 , n3993 , n3994 , n3995 , n3996 , n3997 , n3998 , n3999 , n4000 , n4001 , n4002 , n4003 , n4004 , n4005 , n4006 , n4007 , n4008 , n4009 , n4010 , n4011 , n4012 , n4013 , n4014 , n4015 , n4016 , n4017 , n4018 , n4019 , n4020 , n4021 , n4022 , n4023 , n4024 , n4025 , n4026 , n4027 , n4028 , n4029 , n4030 , n4031 , n4032 , n4033 , n4034 , n4035 , n4036 , n4037 , n4038 , n4039 , n4040 , n4041 , n4042 , n4043 , n4044 , n4045 , n4046 , n4047 , n4048 , n4049 , n4050 , n4051 , n4052 , n4053 , n4054 , n4055 , n4056 , n4057 , n4058 , n4059 , n4060 , n4061 , n4062 , n4063 , n4064 , n4065 , n4066 , n4067 , n4068 , n4069 , n4070 , n4071 , n4072 , n4073 , n4074 , n4075 , n4076 , n4077 , n4078 , n4079 , n4080 , n4081 , n4082 , n4083 , n4084 , n4085 , n4086 , n4087 , n4088 , n4089 , n4090 , n4091 , n4092 , n4093 , n4094 , n4095 , n4096 , n4097 , n4098 , n4099 , n4100 , n4101 , n4102 , n4103 , n4104 , n4105 , n4106 , n4107 , n4108 , n4109 , n4110 , n4111 , n4112 , n4113 , n4114 , n4115 , n4116 , n4117 , n4118 , n4119 , n4120 , n4121 , n4122 , n4123 , n4124 , n4125 , n4126 , n4127 , n4128 , n4129 , n4130 , n4131 , n4132 , n4133 , n4134 , n4135 , n4136 , n4137 , n4138 , n4139 , n4140 , n4141 , n4142 , n4143 , n4144 , n4145 , n4146 , n4147 , n4148 , n4149 , n4150 , n4151 , n4152 , n4153 , n4154 , n4155 , n4156 , n4157 , n4158 , n4159 , n4160 , n4161 , n4162 , n4163 , n4164 , n4165 , n4166 , n4167 , n4168 , n4169 , n4170 , n4171 , n4172 , n4173 , n4174 , n4175 , n4176 , n4177 , n4178 , n4179 , n4180 , n4181 , n4182 , n4183 , n4184 , n4185 , n4186 , n4187 , n4188 , n4189 , n4190 , n4191 , n4192 , n4193 , n4194 , n4195 , n4196 , n4197 , n4198 , n4199 , n4200 , n4201 , n4202 , n4203 , n4204 , n4205 , n4206 , n4207 , n4208 , n4209 , n4210 , n4211 , n4212 , n4213 , n4214 , n4215 , n4216 , n4217 , n4218 , n4219 , n4220 , n4221 , n4222 , n4223 , n4224 , n4225 , n4226 , n4227 , n4228 , n4229 , n4230 , n4231 , n4232 , n4233 , n4234 , n4235 , n4236 , n4237 , n4238 , n4239 , n4240 , n4241 , n4242 , n4243 , n4244 , n4245 , n4246 , n4247 , n4248 , n4249 , n4250 , n4251 , n4252 , n4253 , n4254 , n4255 , n4256 , n4257 , n4258 , n4259 , n4260 , n4261 , n4262 , n4263 , n4264 , n4265 , n4266 , n4267 , n4268 , n4269 , n4270 , n4271 , n4272 , n4273 , n4274 , n4275 , n4276 , n4277 , n4278 , n4279 , n4280 , n4281 , n4282 , n4283 , n4284 , n4285 , n4286 , n4287 , n4288 , n4289 , n4290 , n4291 , n4292 , n4293 , n4294 , n4295 , n4296 , n4297 , n4298 , n4299 , n4300 , n4301 , n4302 , n4303 , n4304 , n4305 , n4306 , n4307 , n4308 , n4309 , n4310 , n4311 , n4312 , n4313 , n4314 , n4315 , n4316 , n4317 , n4318 , n4319 , n4320 , n4321 , n4322 , n4323 , n4324 , n4325 , n4326 , n4327 , n4328 , n4329 , n4330 , n4331 , n4332 , n4333 , n4334 , n4335 , n4336 , n4337 , n4338 , n4339 , n4340 , n4341 , n4342 , n4343 , n4344 , n4345 , n4346 , n4347 , n4348 , n4349 , n4350 , n4351 , n4352 , n4353 , n4354 , n4355 , n4356 , n4357 , n4358 , n4359 , n4360 , n4361 , n4362 , n4363 , n4364 , n4365 , n4366 , n4367 , n4368 , n4369 , n4370 , n4371 , n4372 , n4373 , n4374 , n4375 , n4376 , n4377 , n4378 , n4379 , n4380 , n4381 , n4382 , n4383 , n4384 , n4385 , n4386 , n4387 , n4388 , n4389 , n4390 , n4391 , n4392 , n4393 , n4394 , n4395 , n4396 , n4397 , n4398 , n4399 , n4400 , n4401 , n4402 , n4403 , n4404 , n4405 , n4406 , n4407 , n4408 , n4409 , n4410 , n4411 , n4412 , n4413 , n4414 , n4415 , n4416 , n4417 , n4418 , n4419 , n4420 , n4421 , n4422 , n4423 , n4424 , n4425 , n4426 , n4427 , n4428 , n4429 , n4430 , n4431 , n4432 , n4433 , n4434 , n4435 , n4436 , n4437 , n4438 , n4439 , n4440 , n4441 , n4442 , n4443 , n4444 , n4445 , n4446 , n4447 , n4448 , n4449 , n4450 , n4451 , n4452 , n4453 , n4454 , n4455 , n4456 , n4457 , n4458 , n4459 , n4460 , n4461 , n4462 , n4463 , n4464 , n4465 , n4466 , n4467 , n4468 , n4469 , n4470 , n4471 , n4472 , n4473 , n4474 , n4475 , n4476 , n4477 , n4478 , n4479 , n4480 , n4481 , n4482 , n4483 , n4484 , n4485 , n4486 , n4487 , n4488 , n4489 , n4490 , n4491 , n4492 , n4493 , n4494 , n4495 , n4496 , n4497 , n4498 , n4499 , n4500 , n4501 , n4502 , n4503 , n4504 , n4505 , n4506 , n4507 , n4508 , n4509 , n4510 , n4511 , n4512 , n4513 , n4514 , n4515 , n4516 , n4517 , n4518 , n4519 , n4520 , n4521 , n4522 , n4523 , n4524 , n4525 , n4526 , n4527 , n4528 , n4529 , n4530 , n4531 , n4532 , n4533 , n4534 , n4535 , n4536 , n4537 , n4538 , n4539 , n4540 , n4541 , n4542 , n4543 , n4544 , n4545 , n4546 , n4547 , n4548 , n4549 , n4550 , n4551 , n4552 , n4553 , n4554 , n4555 , n4556 , n4557 , n4558 , n4559 , n4560 , n4561 , n4562 , n4563 , n4564 , n4565 , n4566 , n4567 , n4568 , n4569 , n4570 , n4571 , n4572 , n4573 , n4574 , n4575 , n4576 , n4577 , n4578 , n4579 , n4580 , n4581 , n4582 , n4583 , n4584 , n4585 , n4586 , n4587 , n4588 , n4589 , n4590 , n4591 , n4592 , n4593 , n4594 , n4595 , n4596 , n4597 , n4598 , n4599 , n4600 , n4601 , n4602 , n4603 , n4604 , n4605 , n4606 , n4607 , n4608 , n4609 , n4610 , n4611 , n4612 , n4613 , n4614 , n4615 , n4616 , n4617 , n4618 , n4619 , n4620 , n4621 , n4622 , n4623 , n4624 , n4625 , n4626 , n4627 , n4628 , n4629 , n4630 , n4631 , n4632 , n4633 , n4634 , n4635 , n4636 , n4637 , n4638 , n4639 , n4640 , n4641 , n4642 , n4643 , n4644 , n4645 , n4646 , n4647 , n4648 , n4649 , n4650 , n4651 , n4652 , n4653 , n4654 , n4655 , n4656 , n4657 , n4658 , n4659 , n4660 , n4661 , n4662 , n4663 , n4664 , n4665 , n4666 , n4667 , n4668 , n4669 , n4670 , n4671 , n4672 , n4673 , n4674 , n4675 , n4676 , n4677 , n4678 , n4679 , n4680 , n4681 , n4682 , n4683 , n4684 , n4685 , n4686 , n4687 , n4688 , n4689 , n4690 , n4691 , n4692 , n4693 , n4694 , n4695 , n4696 , n4697 , n4698 , n4699 , n4700 , n4701 , n4702 , n4703 , n4704 , n4705 , n4706 , n4707 , n4708 , n4709 , n4710 , n4711 , n4712 , n4713 , n4714 , n4715 , n4716 , n4717 , n4718 , n4719 , n4720 , n4721 , n4722 , n4723 , n4724 , n4725 , n4726 , n4727 , n4728 , n4729 , n4730 , n4731 , n4732 , n4733 , n4734 , n4735 , n4736 , n4737 , n4738 , n4739 , n4740 , n4741 , n4742 , n4743 , n4744 , n4745 , n4746 , n4747 , n4748 , n4749 , n4750 , n4751 , n4752 , n4753 , n4754 , n4755 , n4756 , n4757 , n4758 , n4759 , n4760 , n4761 , n4762 , n4763 , n4764 , n4765 , n4766 , n4767 , n4768 , n4769 , n4770 , n4771 , n4772 , n4773 , n4774 , n4775 , n4776 , n4777 , n4778 , n4779 , n4780 , n4781 , n4782 , n4783 , n4784 , n4785 , n4786 , n4787 , n4788 , n4789 , n4790 , n4791 , n4792 , n4793 , n4794 , n4795 , n4796 , n4797 , n4798 , n4799 , n4800 , n4801 , n4802 , n4803 , n4804 , n4805 , n4806 , n4807 , n4808 , n4809 , n4810 , n4811 , n4812 , n4813 , n4814 , n4815 , n4816 , n4817 , n4818 , n4819 , n4820 , n4821 , n4822 , n4823 , n4824 , n4825 , n4826 , n4827 , n4828 , n4829 , n4830 , n4831 , n4832 , n4833 , n4834 , n4835 , n4836 , n4837 , n4838 , n4839 , n4840 , n4841 , n4842 , n4843 , n4844 , n4845 , n4846 , n4847 , n4848 , n4849 , n4850 , n4851 , n4852 , n4853 , n4854 , n4855 , n4856 , n4857 , n4858 , n4859 , n4860 , n4861 , n4862 , n4863 , n4864 , n4865 , n4866 , n4867 , n4868 , n4869 , n4870 , n4871 , n4872 , n4873 , n4874 , n4875 , n4876 , n4877 , n4878 , n4879 , n4880 , n4881 , n4882 , n4883 , n4884 , n4885 , n4886 , n4887 , n4888 , n4889 , n4890 , n4891 , n4892 , n4893 , n4894 , n4895 , n4896 , n4897 , n4898 , n4899 , n4900 , n4901 , n4902 , n4903 , n4904 , n4905 , n4906 , n4907 , n4908 , n4909 , n4910 , n4911 , n4912 , n4913 , n4914 , n4915 , n4916 , n4917 , n4918 , n4919 , n4920 , n4921 , n4922 , n4923 , n4924 , n4925 , n4926 , n4927 , n4928 , n4929 , n4930 , n4931 , n4932 , n4933 , n4934 , n4935 , n4936 , n4937 , n4938 , n4939 , n4940 , n4941 , n4942 , n4943 , n4944 , n4945 , n4946 , n4947 , n4948 , n4949 , n4950 , n4951 , n4952 , n4953 , n4954 , n4955 , n4956 , n4957 , n4958 , n4959 , n4960 , n4961 , n4962 , n4963 , n4964 , n4965 , n4966 , n4967 , n4968 , n4969 , n4970 , n4971 , n4972 , n4973 , n4974 , n4975 , n4976 , n4977 , n4978 , n4979 , n4980 , n4981 , n4982 , n4983 , n4984 , n4985 , n4986 , n4987 , n4988 , n4989 , n4990 , n4991 , n4992 , n4993 , n4994 , n4995 , n4996 , n4997 , n4998 , n4999 , n5000 , n5001 , n5002 , n5003 , n5004 , n5005 , n5006 , n5007 , n5008 , n5009 , n5010 , n5011 , n5012 , n5013 , n5014 , n5015 , n5016 , n5017 , n5018 , n5019 , n5020 , n5021 , n5022 , n5023 , n5024 , n5025 , n5026 , n5027 , n5028 , n5029 , n5030 , n5031 , n5032 , n5033 , n5034 , n5035 , n5036 , n5037 , n5038 , n5039 , n5040 , n5041 , n5042 , n5043 , n5044 , n5045 , n5046 , n5047 , n5048 , n5049 , n5050 , n5051 , n5052 , n5053 , n5054 , n5055 , n5056 , n5057 , n5058 , n5059 , n5060 , n5061 , n5062 , n5063 , n5064 , n5065 , n5066 , n5067 , n5068 , n5069 , n5070 , n5071 , n5072 , n5073 , n5074 , n5075 , n5076 , n5077 , n5078 , n5079 , n5080 , n5081 , n5082 , n5083 , n5084 , n5085 , n5086 , n5087 , n5088 , n5089 , n5090 , n5091 , n5092 , n5093 , n5094 , n5095 , n5096 , n5097 , n5098 , n5099 , n5100 , n5101 , n5102 , n5103 , n5104 , n5105 , n5106 , n5107 , n5108 , n5109 , n5110 , n5111 , n5112 , n5113 , n5114 , n5115 , n5116 , n5117 , n5118 , n5119 , n5120 , n5121 , n5122 , n5123 , n5124 , n5125 , n5126 , n5127 , n5128 , n5129 , n5130 , n5131 , n5132 , n5133 , n5134 , n5135 , n5136 , n5137 , n5138 , n5139 , n5140 , n5141 , n5142 , n5143 , n5144 , n5145 , n5146 , n5147 , n5148 , n5149 , n5150 , n5151 , n5152 , n5153 , n5154 , n5155 , n5156 , n5157 , n5158 , n5159 , n5160 , n5161 , n5162 , n5163 , n5164 , n5165 , n5166 , n5167 , n5168 , n5169 , n5170 , n5171 , n5172 , n5173 , n5174 , n5175 , n5176 , n5177 , n5178 , n5179 , n5180 , n5181 , n5182 , n5183 , n5184 , n5185 , n5186 , n5187 , n5188 , n5189 , n5190 , n5191 , n5192 , n5193 , n5194 , n5195 , n5196 , n5197 , n5198 , n5199 , n5200 , n5201 , n5202 , n5203 , n5204 , n5205 , n5206 , n5207 , n5208 , n5209 , n5210 , n5211 , n5212 , n5213 , n5214 , n5215 , n5216 , n5217 , n5218 , n5219 , n5220 , n5221 , n5222 , n5223 , n5224 , n5225 , n5226 , n5227 , n5228 , n5229 , n5230 , n5231 , n5232 , n5233 , n5234 , n5235 , n5236 , n5237 , n5238 , n5239 , n5240 , n5241 , n5242 , n5243 , n5244 , n5245 , n5246 , n5247 , n5248 , n5249 , n5250 , n5251 , n5252 , n5253 , n5254 , n5255 , n5256 , n5257 , n5258 , n5259 , n5260 , n5261 , n5262 , n5263 , n5264 , n5265 , n5266 , n5267 , n5268 , n5269 , n5270 , n5271 , n5272 , n5273 , n5274 , n5275 , n5276 , n5277 , n5278 , n5279 , n5280 , n5281 , n5282 , n5283 , n5284 , n5285 , n5286 , n5287 , n5288 , n5289 , n5290 , n5291 , n5292 , n5293 , n5294 , n5295 , n5296 , n5297 , n5298 , n5299 , n5300 , n5301 , n5302 , n5303 , n5304 , n5305 , n5306 , n5307 , n5308 , n5309 , n5310 , n5311 , n5312 , n5313 , n5314 , n5315 , n5316 , n5317 , n5318 , n5319 , n5320 , n5321 , n5322 , n5323 , n5324 , n5325 , n5326 , n5327 , n5328 , n5329 , n5330 , n5331 , n5332 , n5333 , n5334 , n5335 , n5336 , n5337 , n5338 , n5339 , n5340 , n5341 , n5342 , n5343 , n5344 , n5345 , n5346 , n5347 , n5348 , n5349 , n5350 , n5351 , n5352 , n5353 , n5354 , n5355 , n5356 , n5357 , n5358 , n5359 , n5360 , n5361 , n5362 , n5363 , n5364 , n5365 , n5366 , n5367 , n5368 , n5369 , n5370 , n5371 ;
  assign n214 = ~\IR_reg[6]/NET0131  & ~\IR_reg[7]/NET0131  ;
  assign n215 = ~\IR_reg[0]/NET0131  & ~\IR_reg[1]/NET0131  ;
  assign n216 = ~\IR_reg[2]/NET0131  & n215 ;
  assign n217 = ~\IR_reg[3]/NET0131  & n216 ;
  assign n218 = ~\IR_reg[4]/NET0131  & ~\IR_reg[5]/NET0131  ;
  assign n219 = n217 & n218 ;
  assign n220 = n214 & n219 ;
  assign n222 = ~\IR_reg[10]/NET0131  & ~\IR_reg[8]/NET0131  ;
  assign n223 = ~\IR_reg[9]/NET0131  & n222 ;
  assign n221 = ~\IR_reg[11]/NET0131  & ~\IR_reg[12]/NET0131  ;
  assign n224 = ~\IR_reg[13]/NET0131  & n221 ;
  assign n225 = n223 & n224 ;
  assign n226 = n220 & n225 ;
  assign n227 = \IR_reg[31]/NET0131  & ~n226 ;
  assign n228 = ~\IR_reg[14]/NET0131  & ~\IR_reg[15]/NET0131  ;
  assign n229 = ~\IR_reg[16]/NET0131  & ~\IR_reg[17]/NET0131  ;
  assign n230 = ~\IR_reg[18]/NET0131  & n229 ;
  assign n231 = ~\IR_reg[19]/NET0131  & n230 ;
  assign n232 = n228 & n231 ;
  assign n233 = ~\IR_reg[21]/NET0131  & ~\IR_reg[22]/NET0131  ;
  assign n234 = ~\IR_reg[23]/NET0131  & n233 ;
  assign n235 = ~\IR_reg[20]/NET0131  & n234 ;
  assign n236 = ~\IR_reg[24]/NET0131  & ~\IR_reg[25]/NET0131  ;
  assign n237 = n235 & n236 ;
  assign n238 = n232 & n237 ;
  assign n239 = ~\IR_reg[27]/NET0131  & ~\IR_reg[28]/NET0131  ;
  assign n240 = ~\IR_reg[29]/NET0131  & n239 ;
  assign n241 = ~\IR_reg[26]/NET0131  & n240 ;
  assign n242 = n238 & n241 ;
  assign n243 = \IR_reg[31]/NET0131  & ~n242 ;
  assign n244 = ~n227 & ~n243 ;
  assign n245 = \IR_reg[30]/NET0131  & ~n244 ;
  assign n246 = ~\IR_reg[30]/NET0131  & n244 ;
  assign n247 = ~n245 & ~n246 ;
  assign n248 = ~\IR_reg[8]/NET0131  & n214 ;
  assign n249 = n219 & n248 ;
  assign n250 = ~\IR_reg[10]/NET0131  & ~\IR_reg[9]/NET0131  ;
  assign n251 = n221 & n250 ;
  assign n252 = n249 & n251 ;
  assign n253 = \IR_reg[31]/NET0131  & ~n252 ;
  assign n254 = ~\IR_reg[13]/NET0131  & n228 ;
  assign n255 = ~\IR_reg[20]/NET0131  & n254 ;
  assign n256 = n231 & n255 ;
  assign n257 = ~\IR_reg[26]/NET0131  & n236 ;
  assign n258 = ~\IR_reg[27]/NET0131  & n257 ;
  assign n259 = ~\IR_reg[28]/NET0131  & n234 ;
  assign n260 = n258 & n259 ;
  assign n261 = n256 & n260 ;
  assign n262 = \IR_reg[31]/NET0131  & ~n261 ;
  assign n263 = ~n253 & ~n262 ;
  assign n264 = \IR_reg[29]/NET0131  & ~n263 ;
  assign n265 = ~\IR_reg[29]/NET0131  & n263 ;
  assign n266 = ~n264 & ~n265 ;
  assign n267 = n247 & ~n266 ;
  assign n268 = \reg2_reg[5]/NET0131  & n267 ;
  assign n269 = ~n247 & n266 ;
  assign n270 = \reg1_reg[5]/NET0131  & n269 ;
  assign n279 = ~n268 & ~n270 ;
  assign n271 = n247 & n266 ;
  assign n272 = \reg3_reg[3]/NET0131  & \reg3_reg[4]/NET0131  ;
  assign n273 = \reg3_reg[5]/NET0131  & n272 ;
  assign n274 = ~\reg3_reg[5]/NET0131  & ~n272 ;
  assign n275 = ~n273 & ~n274 ;
  assign n276 = n271 & n275 ;
  assign n277 = ~n247 & ~n266 ;
  assign n278 = \reg0_reg[5]/NET0131  & n277 ;
  assign n280 = ~n276 & ~n278 ;
  assign n281 = n279 & n280 ;
  assign n282 = \reg3_reg[6]/NET0131  & n273 ;
  assign n283 = \reg3_reg[7]/NET0131  & n282 ;
  assign n284 = \reg3_reg[8]/NET0131  & n283 ;
  assign n285 = \reg3_reg[9]/NET0131  & n284 ;
  assign n286 = \reg3_reg[10]/NET0131  & n285 ;
  assign n287 = \reg3_reg[11]/NET0131  & n286 ;
  assign n288 = \reg3_reg[12]/NET0131  & n287 ;
  assign n289 = ~\reg3_reg[13]/NET0131  & ~n288 ;
  assign n290 = \reg3_reg[13]/NET0131  & n288 ;
  assign n291 = ~n289 & ~n290 ;
  assign n292 = n271 & n291 ;
  assign n293 = \reg0_reg[13]/NET0131  & n277 ;
  assign n296 = ~n292 & ~n293 ;
  assign n294 = \reg1_reg[13]/NET0131  & n269 ;
  assign n295 = \reg2_reg[13]/NET0131  & n267 ;
  assign n297 = ~n294 & ~n295 ;
  assign n298 = n296 & n297 ;
  assign n299 = ~\IR_reg[14]/NET0131  & n225 ;
  assign n300 = n220 & n299 ;
  assign n301 = ~\IR_reg[15]/NET0131  & n230 ;
  assign n302 = n300 & n301 ;
  assign n303 = \IR_reg[31]/NET0131  & ~n302 ;
  assign n304 = ~\IR_reg[19]/NET0131  & ~\IR_reg[20]/NET0131  ;
  assign n305 = n233 & n304 ;
  assign n306 = \IR_reg[31]/NET0131  & ~n305 ;
  assign n307 = ~n303 & ~n306 ;
  assign n308 = \IR_reg[23]/NET0131  & ~n307 ;
  assign n309 = ~\IR_reg[23]/NET0131  & n307 ;
  assign n310 = ~n308 & ~n309 ;
  assign n311 = \state_reg[0]/NET0131  & n310 ;
  assign n312 = \B_reg/NET0131  & ~n311 ;
  assign n318 = n226 & n232 ;
  assign n319 = \IR_reg[31]/NET0131  & ~n318 ;
  assign n930 = \IR_reg[20]/NET0131  & ~n319 ;
  assign n931 = ~\IR_reg[20]/NET0131  & n319 ;
  assign n932 = ~n930 & ~n931 ;
  assign n326 = n234 & n304 ;
  assign n327 = n257 & n326 ;
  assign n328 = n302 & n327 ;
  assign n329 = \IR_reg[31]/NET0131  & ~n328 ;
  assign n330 = ~\IR_reg[27]/NET0131  & ~n329 ;
  assign n331 = \IR_reg[27]/NET0131  & n329 ;
  assign n332 = ~n330 & ~n331 ;
  assign n333 = n235 & n258 ;
  assign n334 = \IR_reg[31]/NET0131  & ~n333 ;
  assign n335 = ~n319 & ~n334 ;
  assign n336 = \IR_reg[28]/NET0131  & ~n335 ;
  assign n337 = ~\IR_reg[28]/NET0131  & n335 ;
  assign n338 = ~n336 & ~n337 ;
  assign n339 = ~n332 & ~n338 ;
  assign n340 = \datai[31]_pad  & ~n339 ;
  assign n341 = \reg3_reg[12]/NET0131  & \reg3_reg[13]/NET0131  ;
  assign n342 = \reg3_reg[14]/NET0131  & n341 ;
  assign n343 = \reg3_reg[15]/NET0131  & n342 ;
  assign n344 = \reg3_reg[16]/NET0131  & n343 ;
  assign n345 = n287 & n344 ;
  assign n346 = \reg3_reg[20]/NET0131  & \reg3_reg[21]/NET0131  ;
  assign n347 = \reg3_reg[22]/NET0131  & n346 ;
  assign n348 = \reg3_reg[17]/NET0131  & \reg3_reg[18]/NET0131  ;
  assign n349 = \reg3_reg[19]/NET0131  & \reg3_reg[23]/NET0131  ;
  assign n350 = \reg3_reg[24]/NET0131  & n349 ;
  assign n351 = n348 & n350 ;
  assign n352 = n347 & n351 ;
  assign n353 = n345 & n352 ;
  assign n354 = \reg3_reg[25]/NET0131  & \reg3_reg[26]/NET0131  ;
  assign n355 = \reg3_reg[27]/NET0131  & \reg3_reg[28]/NET0131  ;
  assign n356 = n354 & n355 ;
  assign n357 = n353 & n356 ;
  assign n358 = n271 & n357 ;
  assign n359 = \reg0_reg[31]/NET0131  & n277 ;
  assign n362 = ~n358 & ~n359 ;
  assign n360 = \reg1_reg[31]/NET0131  & n269 ;
  assign n361 = \reg2_reg[31]/NET0131  & n267 ;
  assign n363 = ~n360 & ~n361 ;
  assign n364 = n362 & n363 ;
  assign n367 = \datai[30]_pad  & ~n339 ;
  assign n368 = \reg0_reg[30]/NET0131  & n277 ;
  assign n371 = ~n358 & ~n368 ;
  assign n369 = \reg1_reg[30]/NET0131  & n269 ;
  assign n370 = \reg2_reg[30]/NET0131  & n267 ;
  assign n372 = ~n369 & ~n370 ;
  assign n373 = n371 & n372 ;
  assign n385 = ~n367 & ~n373 ;
  assign n1004 = ~n364 & ~n385 ;
  assign n1005 = n340 & ~n1004 ;
  assign n377 = \datai[29]_pad  & ~n339 ;
  assign n378 = \reg1_reg[29]/NET0131  & n269 ;
  assign n381 = ~n358 & ~n378 ;
  assign n379 = \reg2_reg[29]/NET0131  & n267 ;
  assign n380 = \reg0_reg[29]/NET0131  & n277 ;
  assign n382 = ~n379 & ~n380 ;
  assign n383 = n381 & n382 ;
  assign n384 = ~n377 & ~n383 ;
  assign n388 = n377 & n383 ;
  assign n389 = \datai[28]_pad  & ~n339 ;
  assign n393 = \reg3_reg[25]/NET0131  & n353 ;
  assign n394 = \reg3_reg[26]/NET0131  & n393 ;
  assign n395 = \reg3_reg[27]/NET0131  & n394 ;
  assign n396 = ~\reg3_reg[28]/NET0131  & ~n395 ;
  assign n397 = ~n357 & ~n396 ;
  assign n398 = n271 & n397 ;
  assign n392 = \reg2_reg[28]/NET0131  & n267 ;
  assign n390 = \reg1_reg[28]/NET0131  & n269 ;
  assign n391 = \reg0_reg[28]/NET0131  & n277 ;
  assign n399 = ~n390 & ~n391 ;
  assign n400 = ~n392 & n399 ;
  assign n401 = ~n398 & n400 ;
  assign n404 = ~n389 & ~n401 ;
  assign n941 = ~n388 & n404 ;
  assign n942 = ~n384 & ~n941 ;
  assign n402 = n389 & n401 ;
  assign n403 = ~n388 & ~n402 ;
  assign n405 = \datai[27]_pad  & ~n339 ;
  assign n409 = ~\reg3_reg[27]/NET0131  & ~n394 ;
  assign n410 = ~n395 & ~n409 ;
  assign n411 = n271 & n410 ;
  assign n408 = \reg0_reg[27]/NET0131  & n277 ;
  assign n406 = \reg1_reg[27]/NET0131  & n269 ;
  assign n407 = \reg2_reg[27]/NET0131  & n267 ;
  assign n412 = ~n406 & ~n407 ;
  assign n413 = ~n408 & n412 ;
  assign n414 = ~n411 & n413 ;
  assign n458 = n405 & n414 ;
  assign n445 = \datai[26]_pad  & ~n339 ;
  assign n449 = ~\reg3_reg[26]/NET0131  & ~n393 ;
  assign n450 = ~n394 & ~n449 ;
  assign n451 = n271 & n450 ;
  assign n448 = \reg1_reg[26]/NET0131  & n269 ;
  assign n446 = \reg2_reg[26]/NET0131  & n267 ;
  assign n447 = \reg0_reg[26]/NET0131  & n277 ;
  assign n452 = ~n446 & ~n447 ;
  assign n453 = ~n448 & n452 ;
  assign n454 = ~n451 & n453 ;
  assign n459 = n445 & n454 ;
  assign n417 = \datai[25]_pad  & ~n339 ;
  assign n421 = ~\reg3_reg[25]/NET0131  & ~n353 ;
  assign n422 = ~n393 & ~n421 ;
  assign n423 = n271 & n422 ;
  assign n420 = \reg2_reg[25]/NET0131  & n267 ;
  assign n418 = \reg1_reg[25]/NET0131  & n269 ;
  assign n419 = \reg0_reg[25]/NET0131  & n277 ;
  assign n424 = ~n418 & ~n419 ;
  assign n425 = ~n420 & n424 ;
  assign n426 = ~n423 & n425 ;
  assign n427 = n417 & n426 ;
  assign n444 = ~n417 & ~n426 ;
  assign n428 = \datai[24]_pad  & ~n339 ;
  assign n432 = n345 & n348 ;
  assign n433 = \reg3_reg[19]/NET0131  & n432 ;
  assign n434 = n347 & n433 ;
  assign n435 = \reg3_reg[23]/NET0131  & n434 ;
  assign n436 = ~\reg3_reg[24]/NET0131  & ~n435 ;
  assign n437 = ~n353 & ~n436 ;
  assign n438 = n271 & n437 ;
  assign n431 = \reg2_reg[24]/NET0131  & n267 ;
  assign n429 = \reg1_reg[24]/NET0131  & n269 ;
  assign n430 = \reg0_reg[24]/NET0131  & n277 ;
  assign n439 = ~n429 & ~n430 ;
  assign n440 = ~n431 & n439 ;
  assign n441 = ~n438 & n440 ;
  assign n922 = ~n428 & ~n441 ;
  assign n923 = ~n444 & ~n922 ;
  assign n990 = ~n427 & ~n923 ;
  assign n991 = ~n459 & n990 ;
  assign n415 = ~n405 & ~n414 ;
  assign n455 = ~n445 & ~n454 ;
  assign n992 = ~n415 & ~n455 ;
  assign n993 = ~n991 & n992 ;
  assign n994 = ~n458 & ~n993 ;
  assign n442 = n428 & n441 ;
  assign n986 = ~n427 & ~n459 ;
  assign n987 = ~n458 & n986 ;
  assign n988 = ~n442 & n987 ;
  assign n476 = \datai[22]_pad  & ~n339 ;
  assign n480 = n346 & n433 ;
  assign n481 = ~\reg3_reg[22]/NET0131  & ~n480 ;
  assign n482 = ~n434 & ~n481 ;
  assign n483 = n271 & n482 ;
  assign n479 = \reg0_reg[22]/NET0131  & n277 ;
  assign n477 = \reg1_reg[22]/NET0131  & n269 ;
  assign n478 = \reg2_reg[22]/NET0131  & n267 ;
  assign n484 = ~n477 & ~n478 ;
  assign n485 = ~n479 & n484 ;
  assign n486 = ~n483 & n485 ;
  assign n894 = n476 & n486 ;
  assign n465 = \datai[23]_pad  & ~n339 ;
  assign n469 = ~\reg3_reg[23]/NET0131  & ~n434 ;
  assign n470 = ~n435 & ~n469 ;
  assign n471 = n271 & n470 ;
  assign n468 = \reg1_reg[23]/NET0131  & n269 ;
  assign n466 = \reg2_reg[23]/NET0131  & n267 ;
  assign n467 = \reg0_reg[23]/NET0131  & n277 ;
  assign n472 = ~n466 & ~n467 ;
  assign n473 = ~n468 & n472 ;
  assign n474 = ~n471 & n473 ;
  assign n895 = n465 & n474 ;
  assign n896 = ~n894 & ~n895 ;
  assign n830 = \datai[21]_pad  & ~n339 ;
  assign n834 = \reg3_reg[20]/NET0131  & n433 ;
  assign n835 = ~\reg3_reg[21]/NET0131  & ~n834 ;
  assign n836 = ~n480 & ~n835 ;
  assign n837 = n271 & n836 ;
  assign n833 = \reg2_reg[21]/NET0131  & n267 ;
  assign n831 = \reg0_reg[21]/NET0131  & n277 ;
  assign n832 = \reg1_reg[21]/NET0131  & n269 ;
  assign n838 = ~n831 & ~n832 ;
  assign n839 = ~n833 & n838 ;
  assign n840 = ~n837 & n839 ;
  assign n841 = ~n830 & ~n840 ;
  assign n842 = \datai[20]_pad  & ~n339 ;
  assign n846 = ~\reg3_reg[20]/NET0131  & ~n433 ;
  assign n847 = ~n834 & ~n846 ;
  assign n848 = n271 & n847 ;
  assign n845 = \reg2_reg[20]/NET0131  & n267 ;
  assign n843 = \reg0_reg[20]/NET0131  & n277 ;
  assign n844 = \reg1_reg[20]/NET0131  & n269 ;
  assign n849 = ~n843 & ~n844 ;
  assign n850 = ~n845 & n849 ;
  assign n851 = ~n848 & n850 ;
  assign n852 = ~n842 & ~n851 ;
  assign n853 = ~n841 & ~n852 ;
  assign n897 = n830 & n840 ;
  assign n898 = ~n853 & ~n897 ;
  assign n899 = n896 & n898 ;
  assign n475 = ~n465 & ~n474 ;
  assign n487 = ~n476 & ~n486 ;
  assign n488 = ~n475 & ~n487 ;
  assign n900 = ~n488 & ~n895 ;
  assign n901 = ~n899 & ~n900 ;
  assign n792 = ~\IR_reg[19]/NET0131  & ~n303 ;
  assign n793 = \IR_reg[19]/NET0131  & n303 ;
  assign n794 = ~n792 & ~n793 ;
  assign n795 = n339 & n794 ;
  assign n796 = \datai[19]_pad  & ~n339 ;
  assign n797 = ~n795 & ~n796 ;
  assign n801 = ~\reg3_reg[19]/NET0131  & ~n432 ;
  assign n802 = ~n433 & ~n801 ;
  assign n803 = n271 & n802 ;
  assign n800 = \reg1_reg[19]/NET0131  & n269 ;
  assign n798 = \reg0_reg[19]/NET0131  & n277 ;
  assign n799 = \reg2_reg[19]/NET0131  & n267 ;
  assign n804 = ~n798 & ~n799 ;
  assign n805 = ~n800 & n804 ;
  assign n806 = ~n803 & n805 ;
  assign n902 = ~n797 & n806 ;
  assign n808 = ~\IR_reg[15]/NET0131  & n300 ;
  assign n809 = \IR_reg[31]/NET0131  & ~n808 ;
  assign n810 = \IR_reg[31]/NET0131  & ~n229 ;
  assign n811 = ~n809 & ~n810 ;
  assign n812 = \IR_reg[18]/NET0131  & ~n811 ;
  assign n813 = ~\IR_reg[18]/NET0131  & n811 ;
  assign n814 = ~n812 & ~n813 ;
  assign n815 = n339 & ~n814 ;
  assign n816 = ~\datai[18]_pad  & ~n339 ;
  assign n817 = ~n815 & ~n816 ;
  assign n821 = \reg3_reg[17]/NET0131  & n345 ;
  assign n822 = ~\reg3_reg[18]/NET0131  & ~n821 ;
  assign n823 = ~n432 & ~n822 ;
  assign n824 = n271 & n823 ;
  assign n820 = \reg2_reg[18]/NET0131  & n267 ;
  assign n818 = \reg0_reg[18]/NET0131  & n277 ;
  assign n819 = \reg1_reg[18]/NET0131  & n269 ;
  assign n825 = ~n818 & ~n819 ;
  assign n826 = ~n820 & n825 ;
  assign n827 = ~n824 & n826 ;
  assign n903 = n817 & n827 ;
  assign n904 = ~n902 & ~n903 ;
  assign n854 = \reg2_reg[17]/NET0131  & n267 ;
  assign n855 = \reg1_reg[17]/NET0131  & n269 ;
  assign n860 = ~n854 & ~n855 ;
  assign n856 = ~\reg3_reg[17]/NET0131  & ~n345 ;
  assign n857 = ~n821 & ~n856 ;
  assign n858 = n271 & n857 ;
  assign n859 = \reg0_reg[17]/NET0131  & n277 ;
  assign n861 = ~n858 & ~n859 ;
  assign n862 = n860 & n861 ;
  assign n863 = ~\IR_reg[16]/NET0131  & n254 ;
  assign n864 = n252 & n863 ;
  assign n865 = \IR_reg[31]/NET0131  & ~n864 ;
  assign n866 = \IR_reg[17]/NET0131  & n865 ;
  assign n867 = ~\IR_reg[17]/NET0131  & ~n865 ;
  assign n868 = ~n866 & ~n867 ;
  assign n869 = n339 & ~n868 ;
  assign n870 = ~\datai[17]_pad  & ~n339 ;
  assign n871 = ~n869 & ~n870 ;
  assign n872 = ~n862 & ~n871 ;
  assign n873 = ~\IR_reg[16]/NET0131  & ~n809 ;
  assign n874 = \IR_reg[16]/NET0131  & n809 ;
  assign n875 = ~n873 & ~n874 ;
  assign n876 = n339 & ~n875 ;
  assign n877 = ~\datai[16]_pad  & ~n339 ;
  assign n878 = ~n876 & ~n877 ;
  assign n507 = n287 & n343 ;
  assign n879 = ~\reg3_reg[16]/NET0131  & ~n507 ;
  assign n880 = ~n345 & ~n879 ;
  assign n881 = n271 & n880 ;
  assign n882 = \reg0_reg[16]/NET0131  & n277 ;
  assign n885 = ~n881 & ~n882 ;
  assign n883 = \reg1_reg[16]/NET0131  & n269 ;
  assign n884 = \reg2_reg[16]/NET0131  & n267 ;
  assign n886 = ~n883 & ~n884 ;
  assign n887 = n885 & n886 ;
  assign n888 = ~n878 & ~n887 ;
  assign n889 = ~n872 & ~n888 ;
  assign n905 = n862 & n871 ;
  assign n946 = ~n889 & ~n905 ;
  assign n947 = n904 & n946 ;
  assign n807 = n797 & ~n806 ;
  assign n828 = ~n817 & ~n827 ;
  assign n829 = ~n807 & ~n828 ;
  assign n948 = ~n829 & ~n902 ;
  assign n949 = ~n947 & ~n948 ;
  assign n912 = n842 & n851 ;
  assign n950 = ~n897 & ~n912 ;
  assign n951 = n896 & n950 ;
  assign n952 = ~n949 & n951 ;
  assign n953 = n901 & ~n952 ;
  assign n491 = ~\reg3_reg[14]/NET0131  & ~n290 ;
  assign n492 = n287 & n342 ;
  assign n493 = ~n491 & ~n492 ;
  assign n494 = n271 & n493 ;
  assign n495 = \reg1_reg[14]/NET0131  & n269 ;
  assign n489 = \reg0_reg[14]/NET0131  & n277 ;
  assign n490 = \reg2_reg[14]/NET0131  & n267 ;
  assign n496 = ~n489 & ~n490 ;
  assign n497 = ~n495 & n496 ;
  assign n498 = ~n494 & n497 ;
  assign n499 = ~\IR_reg[14]/NET0131  & ~n227 ;
  assign n500 = \IR_reg[14]/NET0131  & n227 ;
  assign n501 = ~n499 & ~n500 ;
  assign n502 = n339 & n501 ;
  assign n503 = \datai[14]_pad  & ~n339 ;
  assign n504 = ~n502 & ~n503 ;
  assign n505 = n498 & ~n504 ;
  assign n506 = ~\reg3_reg[15]/NET0131  & ~n492 ;
  assign n508 = ~n506 & ~n507 ;
  assign n509 = n271 & n508 ;
  assign n510 = \reg0_reg[15]/NET0131  & n277 ;
  assign n513 = ~n509 & ~n510 ;
  assign n511 = \reg2_reg[15]/NET0131  & n267 ;
  assign n512 = \reg1_reg[15]/NET0131  & n269 ;
  assign n514 = ~n511 & ~n512 ;
  assign n515 = n513 & n514 ;
  assign n516 = \IR_reg[31]/NET0131  & ~n300 ;
  assign n517 = \IR_reg[15]/NET0131  & n516 ;
  assign n518 = ~\IR_reg[15]/NET0131  & ~n516 ;
  assign n519 = ~n517 & ~n518 ;
  assign n520 = n339 & ~n519 ;
  assign n521 = ~\datai[15]_pad  & ~n339 ;
  assign n522 = ~n520 & ~n521 ;
  assign n523 = n515 & n522 ;
  assign n524 = ~n505 & ~n523 ;
  assign n525 = ~\IR_reg[13]/NET0131  & ~n253 ;
  assign n526 = \IR_reg[13]/NET0131  & n253 ;
  assign n527 = ~n525 & ~n526 ;
  assign n528 = n339 & n527 ;
  assign n529 = \datai[13]_pad  & ~n339 ;
  assign n530 = ~n528 & ~n529 ;
  assign n531 = n298 & ~n530 ;
  assign n532 = ~n298 & n530 ;
  assign n533 = \reg2_reg[12]/NET0131  & n267 ;
  assign n534 = \reg0_reg[12]/NET0131  & n277 ;
  assign n539 = ~n533 & ~n534 ;
  assign n535 = \reg1_reg[12]/NET0131  & n269 ;
  assign n536 = ~\reg3_reg[12]/NET0131  & ~n287 ;
  assign n537 = ~n288 & ~n536 ;
  assign n538 = n271 & n537 ;
  assign n540 = ~n535 & ~n538 ;
  assign n541 = n539 & n540 ;
  assign n542 = n220 & n223 ;
  assign n543 = \IR_reg[31]/NET0131  & ~n542 ;
  assign n544 = \IR_reg[11]/NET0131  & \IR_reg[31]/NET0131  ;
  assign n545 = ~n543 & ~n544 ;
  assign n546 = \IR_reg[12]/NET0131  & ~n545 ;
  assign n547 = ~\IR_reg[12]/NET0131  & n545 ;
  assign n548 = ~n546 & ~n547 ;
  assign n549 = n339 & ~n548 ;
  assign n550 = ~\datai[12]_pad  & ~n339 ;
  assign n551 = ~n549 & ~n550 ;
  assign n552 = ~n541 & ~n551 ;
  assign n553 = ~n532 & ~n552 ;
  assign n554 = ~n531 & ~n553 ;
  assign n555 = n524 & n554 ;
  assign n556 = ~n498 & n504 ;
  assign n557 = ~n515 & ~n522 ;
  assign n558 = ~n556 & ~n557 ;
  assign n559 = ~n523 & ~n558 ;
  assign n560 = ~n555 & ~n559 ;
  assign n567 = \datai[11]_pad  & ~n339 ;
  assign n568 = \IR_reg[11]/NET0131  & ~n543 ;
  assign n569 = ~\IR_reg[11]/NET0131  & n543 ;
  assign n570 = ~n568 & ~n569 ;
  assign n571 = n339 & ~n570 ;
  assign n572 = ~n567 & ~n571 ;
  assign n573 = \reg1_reg[11]/NET0131  & n269 ;
  assign n574 = ~\reg3_reg[11]/NET0131  & ~n286 ;
  assign n575 = ~n287 & ~n574 ;
  assign n576 = n271 & n575 ;
  assign n579 = ~n573 & ~n576 ;
  assign n577 = \reg2_reg[11]/NET0131  & n267 ;
  assign n578 = \reg0_reg[11]/NET0131  & n277 ;
  assign n580 = ~n577 & ~n578 ;
  assign n581 = n579 & n580 ;
  assign n583 = ~n572 & n581 ;
  assign n584 = ~\reg3_reg[10]/NET0131  & ~n285 ;
  assign n585 = ~n286 & ~n584 ;
  assign n586 = n271 & n585 ;
  assign n587 = \reg2_reg[10]/NET0131  & n267 ;
  assign n590 = ~n586 & ~n587 ;
  assign n588 = \reg0_reg[10]/NET0131  & n277 ;
  assign n589 = \reg1_reg[10]/NET0131  & n269 ;
  assign n591 = ~n588 & ~n589 ;
  assign n592 = n590 & n591 ;
  assign n593 = \IR_reg[31]/NET0131  & ~n249 ;
  assign n594 = \IR_reg[31]/NET0131  & \IR_reg[9]/NET0131  ;
  assign n595 = ~n593 & ~n594 ;
  assign n596 = \IR_reg[10]/NET0131  & ~n595 ;
  assign n597 = ~\IR_reg[10]/NET0131  & n595 ;
  assign n598 = ~n596 & ~n597 ;
  assign n599 = n339 & ~n598 ;
  assign n600 = ~\datai[10]_pad  & ~n339 ;
  assign n601 = ~n599 & ~n600 ;
  assign n602 = n592 & n601 ;
  assign n603 = ~n583 & ~n602 ;
  assign n604 = \datai[9]_pad  & ~n339 ;
  assign n605 = \IR_reg[9]/NET0131  & ~n593 ;
  assign n606 = ~\IR_reg[9]/NET0131  & n593 ;
  assign n607 = ~n605 & ~n606 ;
  assign n608 = n339 & ~n607 ;
  assign n609 = ~n604 & ~n608 ;
  assign n610 = ~\reg3_reg[9]/NET0131  & ~n284 ;
  assign n611 = ~n285 & ~n610 ;
  assign n612 = n271 & n611 ;
  assign n613 = \reg1_reg[9]/NET0131  & n269 ;
  assign n616 = ~n612 & ~n613 ;
  assign n614 = \reg2_reg[9]/NET0131  & n267 ;
  assign n615 = \reg0_reg[9]/NET0131  & n277 ;
  assign n617 = ~n614 & ~n615 ;
  assign n618 = n616 & n617 ;
  assign n638 = n609 & ~n618 ;
  assign n619 = ~n609 & n618 ;
  assign n620 = ~\reg3_reg[8]/NET0131  & ~n283 ;
  assign n621 = ~n284 & ~n620 ;
  assign n622 = n271 & n621 ;
  assign n623 = \reg1_reg[8]/NET0131  & n269 ;
  assign n626 = ~n622 & ~n623 ;
  assign n624 = \reg2_reg[8]/NET0131  & n267 ;
  assign n625 = \reg0_reg[8]/NET0131  & n277 ;
  assign n627 = ~n624 & ~n625 ;
  assign n628 = n626 & n627 ;
  assign n629 = \IR_reg[31]/NET0131  & ~n220 ;
  assign n630 = \IR_reg[8]/NET0131  & n629 ;
  assign n631 = ~\IR_reg[8]/NET0131  & ~n629 ;
  assign n632 = ~n630 & ~n631 ;
  assign n633 = n339 & ~n632 ;
  assign n634 = ~\datai[8]_pad  & ~n339 ;
  assign n635 = ~n633 & ~n634 ;
  assign n782 = ~n628 & ~n635 ;
  assign n956 = ~n619 & n782 ;
  assign n957 = ~n638 & ~n956 ;
  assign n958 = n603 & ~n957 ;
  assign n582 = n572 & ~n581 ;
  assign n639 = ~n592 & ~n601 ;
  assign n959 = ~n582 & ~n639 ;
  assign n960 = ~n583 & ~n959 ;
  assign n961 = ~n958 & ~n960 ;
  assign n561 = n541 & n551 ;
  assign n562 = ~n531 & ~n561 ;
  assign n962 = n524 & n562 ;
  assign n963 = ~n961 & n962 ;
  assign n964 = n560 & ~n963 ;
  assign n646 = \datai[6]_pad  & ~n339 ;
  assign n647 = \IR_reg[31]/NET0131  & ~n219 ;
  assign n648 = \IR_reg[6]/NET0131  & ~n647 ;
  assign n649 = ~\IR_reg[6]/NET0131  & n647 ;
  assign n650 = ~n648 & ~n649 ;
  assign n651 = n339 & ~n650 ;
  assign n652 = ~n646 & ~n651 ;
  assign n653 = \reg2_reg[6]/NET0131  & n267 ;
  assign n654 = \reg1_reg[6]/NET0131  & n269 ;
  assign n659 = ~n653 & ~n654 ;
  assign n655 = ~\reg3_reg[6]/NET0131  & ~n273 ;
  assign n656 = ~n282 & ~n655 ;
  assign n657 = n271 & n656 ;
  assign n658 = \reg0_reg[6]/NET0131  & n277 ;
  assign n660 = ~n657 & ~n658 ;
  assign n661 = n659 & n660 ;
  assign n662 = ~n652 & n661 ;
  assign n663 = \reg1_reg[7]/NET0131  & n269 ;
  assign n664 = \reg0_reg[7]/NET0131  & n277 ;
  assign n669 = ~n663 & ~n664 ;
  assign n665 = ~\reg3_reg[7]/NET0131  & ~n282 ;
  assign n666 = ~n283 & ~n665 ;
  assign n667 = n271 & n666 ;
  assign n668 = \reg2_reg[7]/NET0131  & n267 ;
  assign n670 = ~n667 & ~n668 ;
  assign n671 = n669 & n670 ;
  assign n672 = \IR_reg[31]/NET0131  & \IR_reg[6]/NET0131  ;
  assign n673 = ~n647 & ~n672 ;
  assign n674 = \IR_reg[7]/NET0131  & ~n673 ;
  assign n675 = ~\IR_reg[7]/NET0131  & n673 ;
  assign n676 = ~n674 & ~n675 ;
  assign n677 = n339 & ~n676 ;
  assign n678 = ~\datai[7]_pad  & ~n339 ;
  assign n679 = ~n677 & ~n678 ;
  assign n680 = n671 & n679 ;
  assign n681 = ~n662 & ~n680 ;
  assign n694 = \datai[4]_pad  & ~n339 ;
  assign n682 = \IR_reg[31]/NET0131  & ~n217 ;
  assign n695 = \IR_reg[4]/NET0131  & ~n682 ;
  assign n696 = ~\IR_reg[4]/NET0131  & n682 ;
  assign n697 = ~n695 & ~n696 ;
  assign n698 = n339 & ~n697 ;
  assign n699 = ~n694 & ~n698 ;
  assign n700 = ~\reg3_reg[3]/NET0131  & ~\reg3_reg[4]/NET0131  ;
  assign n701 = ~n272 & ~n700 ;
  assign n702 = n271 & n701 ;
  assign n703 = \reg1_reg[4]/NET0131  & n269 ;
  assign n706 = ~n702 & ~n703 ;
  assign n704 = \reg2_reg[4]/NET0131  & n267 ;
  assign n705 = \reg0_reg[4]/NET0131  & n277 ;
  assign n707 = ~n704 & ~n705 ;
  assign n708 = n706 & n707 ;
  assign n709 = ~n699 & n708 ;
  assign n683 = \IR_reg[31]/NET0131  & \IR_reg[4]/NET0131  ;
  assign n684 = ~n682 & ~n683 ;
  assign n685 = \IR_reg[5]/NET0131  & ~n684 ;
  assign n686 = ~\IR_reg[5]/NET0131  & n684 ;
  assign n687 = ~n685 & ~n686 ;
  assign n688 = n339 & ~n687 ;
  assign n689 = ~\datai[5]_pad  & ~n339 ;
  assign n690 = ~n688 & ~n689 ;
  assign n710 = n281 & n690 ;
  assign n711 = ~n709 & ~n710 ;
  assign n729 = \reg1_reg[2]/NET0131  & n269 ;
  assign n730 = \reg0_reg[2]/NET0131  & n277 ;
  assign n733 = ~n729 & ~n730 ;
  assign n731 = \reg2_reg[2]/NET0131  & n267 ;
  assign n732 = \reg3_reg[2]/NET0131  & n271 ;
  assign n734 = ~n731 & ~n732 ;
  assign n735 = n733 & n734 ;
  assign n736 = \datai[2]_pad  & ~n339 ;
  assign n737 = \IR_reg[31]/NET0131  & ~n215 ;
  assign n738 = \IR_reg[2]/NET0131  & ~n737 ;
  assign n739 = ~\IR_reg[2]/NET0131  & n737 ;
  assign n740 = ~n738 & ~n739 ;
  assign n741 = n339 & ~n740 ;
  assign n742 = ~n736 & ~n741 ;
  assign n743 = n735 & ~n742 ;
  assign n712 = ~\reg3_reg[3]/NET0131  & n271 ;
  assign n713 = \reg1_reg[3]/NET0131  & n269 ;
  assign n716 = ~n712 & ~n713 ;
  assign n714 = \reg2_reg[3]/NET0131  & n267 ;
  assign n715 = \reg0_reg[3]/NET0131  & n277 ;
  assign n717 = ~n714 & ~n715 ;
  assign n718 = n716 & n717 ;
  assign n719 = \IR_reg[31]/NET0131  & ~n216 ;
  assign n720 = \IR_reg[3]/NET0131  & n719 ;
  assign n721 = ~\IR_reg[3]/NET0131  & ~n719 ;
  assign n722 = ~n720 & ~n721 ;
  assign n723 = n339 & n722 ;
  assign n724 = \datai[3]_pad  & ~n339 ;
  assign n725 = ~n723 & ~n724 ;
  assign n744 = n718 & ~n725 ;
  assign n745 = ~n743 & ~n744 ;
  assign n746 = \reg3_reg[1]/NET0131  & n271 ;
  assign n747 = \reg1_reg[1]/NET0131  & n269 ;
  assign n750 = ~n746 & ~n747 ;
  assign n748 = \reg0_reg[1]/NET0131  & n277 ;
  assign n749 = \reg2_reg[1]/NET0131  & n267 ;
  assign n751 = ~n748 & ~n749 ;
  assign n752 = n750 & n751 ;
  assign n753 = \IR_reg[1]/NET0131  & ~\IR_reg[31]/NET0131  ;
  assign n754 = \IR_reg[0]/NET0131  & \IR_reg[1]/NET0131  ;
  assign n755 = n737 & ~n754 ;
  assign n756 = ~n753 & ~n755 ;
  assign n757 = n339 & ~n756 ;
  assign n758 = \datai[1]_pad  & ~n339 ;
  assign n759 = ~n757 & ~n758 ;
  assign n761 = n752 & ~n759 ;
  assign n760 = ~n752 & n759 ;
  assign n762 = \reg0_reg[0]/NET0131  & n277 ;
  assign n763 = \reg1_reg[0]/NET0131  & n269 ;
  assign n766 = ~n762 & ~n763 ;
  assign n764 = \reg2_reg[0]/NET0131  & n267 ;
  assign n765 = \reg3_reg[0]/NET0131  & n271 ;
  assign n767 = ~n764 & ~n765 ;
  assign n768 = n766 & n767 ;
  assign n769 = \datai[0]_pad  & ~n339 ;
  assign n770 = \IR_reg[0]/NET0131  & n339 ;
  assign n771 = ~n769 & ~n770 ;
  assign n965 = n768 & ~n771 ;
  assign n966 = ~n760 & n965 ;
  assign n967 = ~n761 & ~n966 ;
  assign n968 = n745 & n967 ;
  assign n726 = ~n718 & n725 ;
  assign n774 = ~n735 & n742 ;
  assign n969 = ~n726 & ~n774 ;
  assign n970 = ~n744 & ~n969 ;
  assign n971 = ~n968 & ~n970 ;
  assign n972 = n711 & ~n971 ;
  assign n691 = ~n281 & ~n690 ;
  assign n727 = n699 & ~n708 ;
  assign n973 = ~n710 & n727 ;
  assign n974 = ~n691 & ~n973 ;
  assign n975 = ~n972 & n974 ;
  assign n976 = n681 & ~n975 ;
  assign n692 = n652 & ~n661 ;
  assign n783 = ~n671 & ~n679 ;
  assign n977 = ~n692 & ~n783 ;
  assign n978 = ~n680 & ~n977 ;
  assign n979 = ~n976 & ~n978 ;
  assign n1006 = n964 & n979 ;
  assign n563 = ~n532 & ~n556 ;
  assign n564 = ~n562 & n563 ;
  assign n565 = n524 & ~n564 ;
  assign n566 = ~n557 & ~n565 ;
  assign n636 = n628 & n635 ;
  assign n637 = ~n619 & ~n636 ;
  assign n640 = ~n638 & ~n639 ;
  assign n641 = ~n637 & n640 ;
  assign n642 = n603 & ~n641 ;
  assign n643 = ~n582 & ~n642 ;
  assign n644 = ~n566 & ~n643 ;
  assign n645 = n560 & ~n644 ;
  assign n906 = n878 & n887 ;
  assign n907 = ~n905 & ~n906 ;
  assign n954 = n904 & n907 ;
  assign n955 = n951 & n954 ;
  assign n1007 = ~n645 & n955 ;
  assign n1008 = ~n1006 & n1007 ;
  assign n1009 = n953 & ~n1008 ;
  assign n1010 = n988 & ~n1009 ;
  assign n1011 = ~n994 & ~n1010 ;
  assign n1012 = n403 & ~n1011 ;
  assign n1013 = n942 & ~n1012 ;
  assign n366 = ~n340 & ~n364 ;
  assign n1014 = ~n364 & ~n373 ;
  assign n1015 = n367 & ~n1014 ;
  assign n1016 = ~n366 & ~n1015 ;
  assign n1017 = ~n1013 & n1016 ;
  assign n1018 = ~n1005 & ~n1017 ;
  assign n1020 = n932 & ~n1018 ;
  assign n313 = \IR_reg[31]/NET0131  & ~n256 ;
  assign n314 = ~n253 & ~n313 ;
  assign n315 = \IR_reg[21]/NET0131  & ~n314 ;
  assign n316 = ~\IR_reg[21]/NET0131  & n314 ;
  assign n317 = ~n315 & ~n316 ;
  assign n320 = ~\IR_reg[20]/NET0131  & ~\IR_reg[21]/NET0131  ;
  assign n321 = \IR_reg[31]/NET0131  & ~n320 ;
  assign n322 = ~n319 & ~n321 ;
  assign n323 = \IR_reg[22]/NET0131  & ~n322 ;
  assign n324 = ~\IR_reg[22]/NET0131  & n322 ;
  assign n325 = ~n323 & ~n324 ;
  assign n1003 = n317 & n325 ;
  assign n1019 = ~n932 & n1018 ;
  assign n1021 = n1003 & ~n1019 ;
  assign n1022 = ~n1020 & n1021 ;
  assign n365 = n340 & n364 ;
  assign n386 = ~n365 & ~n385 ;
  assign n374 = n367 & n373 ;
  assign n943 = ~n374 & ~n942 ;
  assign n944 = n386 & ~n943 ;
  assign n945 = ~n366 & ~n944 ;
  assign n980 = n603 & n637 ;
  assign n981 = ~n979 & n980 ;
  assign n982 = n962 & n981 ;
  assign n983 = n964 & ~n982 ;
  assign n984 = n955 & ~n983 ;
  assign n985 = n953 & ~n984 ;
  assign n989 = ~n985 & n988 ;
  assign n995 = ~n989 & ~n994 ;
  assign n375 = ~n366 & ~n374 ;
  assign n996 = n375 & n403 ;
  assign n997 = ~n995 & n996 ;
  assign n998 = ~n945 & ~n997 ;
  assign n1000 = ~n932 & n998 ;
  assign n940 = ~n317 & ~n325 ;
  assign n999 = n932 & ~n998 ;
  assign n1001 = n940 & ~n999 ;
  assign n1002 = ~n1000 & n1001 ;
  assign n693 = ~n691 & ~n692 ;
  assign n728 = ~n726 & ~n727 ;
  assign n772 = ~n768 & n771 ;
  assign n773 = ~n761 & n772 ;
  assign n775 = ~n760 & ~n774 ;
  assign n776 = ~n773 & n775 ;
  assign n777 = n745 & ~n776 ;
  assign n778 = n728 & ~n777 ;
  assign n779 = n711 & ~n778 ;
  assign n780 = n693 & ~n779 ;
  assign n781 = n681 & ~n780 ;
  assign n786 = ~n532 & n640 ;
  assign n784 = ~n782 & ~n783 ;
  assign n785 = ~n552 & ~n582 ;
  assign n787 = n784 & n785 ;
  assign n788 = n786 & n787 ;
  assign n789 = n558 & n788 ;
  assign n790 = ~n781 & n789 ;
  assign n791 = ~n645 & ~n790 ;
  assign n890 = n829 & n889 ;
  assign n891 = n488 & n890 ;
  assign n892 = n853 & n891 ;
  assign n893 = ~n791 & n892 ;
  assign n913 = ~n894 & ~n897 ;
  assign n914 = ~n912 & n913 ;
  assign n915 = n841 & ~n894 ;
  assign n916 = n488 & ~n915 ;
  assign n917 = ~n914 & n916 ;
  assign n908 = ~n828 & ~n872 ;
  assign n909 = ~n907 & n908 ;
  assign n910 = n904 & ~n909 ;
  assign n911 = ~n807 & ~n910 ;
  assign n918 = ~n895 & ~n911 ;
  assign n919 = ~n917 & n918 ;
  assign n920 = n901 & ~n919 ;
  assign n921 = ~n893 & ~n920 ;
  assign n416 = ~n404 & ~n415 ;
  assign n387 = ~n384 & n386 ;
  assign n924 = n387 & ~n455 ;
  assign n925 = n416 & n924 ;
  assign n926 = n923 & n925 ;
  assign n927 = ~n921 & n926 ;
  assign n376 = ~n365 & ~n375 ;
  assign n443 = ~n427 & ~n442 ;
  assign n456 = ~n444 & ~n455 ;
  assign n457 = ~n443 & n456 ;
  assign n460 = ~n458 & ~n459 ;
  assign n461 = ~n457 & n460 ;
  assign n462 = n416 & ~n461 ;
  assign n463 = n403 & ~n462 ;
  assign n464 = n387 & ~n463 ;
  assign n928 = ~n376 & ~n464 ;
  assign n929 = ~n927 & n928 ;
  assign n934 = ~n929 & n932 ;
  assign n933 = n929 & ~n932 ;
  assign n935 = \B_reg/NET0131  & n310 ;
  assign n936 = ~n933 & ~n935 ;
  assign n937 = ~n934 & n936 ;
  assign n938 = ~n317 & n325 ;
  assign n939 = ~n937 & n938 ;
  assign n1023 = n932 & n935 ;
  assign n1078 = ~n417 & n426 ;
  assign n1079 = n417 & ~n426 ;
  assign n1080 = ~n1078 & ~n1079 ;
  assign n1081 = ~n807 & ~n902 ;
  assign n1108 = ~n1080 & n1081 ;
  assign n1082 = n842 & ~n851 ;
  assign n1083 = ~n842 & n851 ;
  assign n1084 = ~n1082 & ~n1083 ;
  assign n1088 = n817 & ~n827 ;
  assign n1089 = ~n817 & n827 ;
  assign n1090 = ~n1088 & ~n1089 ;
  assign n1109 = ~n1084 & ~n1090 ;
  assign n1110 = n1108 & n1109 ;
  assign n1092 = n375 & n386 ;
  assign n1024 = n541 & ~n551 ;
  assign n1025 = ~n541 & n551 ;
  assign n1026 = ~n1024 & ~n1025 ;
  assign n1027 = ~n662 & ~n692 ;
  assign n1093 = ~n1026 & n1027 ;
  assign n1106 = n1092 & n1093 ;
  assign n1040 = ~n505 & ~n556 ;
  assign n1058 = n445 & ~n454 ;
  assign n1059 = ~n445 & n454 ;
  assign n1060 = ~n1058 & ~n1059 ;
  assign n1107 = n1040 & ~n1060 ;
  assign n1111 = n1106 & n1107 ;
  assign n1118 = n1110 & n1111 ;
  assign n1048 = n428 & ~n441 ;
  assign n1049 = ~n428 & n441 ;
  assign n1050 = ~n1048 & ~n1049 ;
  assign n1071 = ~n389 & n401 ;
  assign n1072 = n389 & ~n401 ;
  assign n1073 = ~n1071 & ~n1072 ;
  assign n1119 = ~n1050 & ~n1073 ;
  assign n1120 = n1118 & n1119 ;
  assign n1045 = n830 & ~n840 ;
  assign n1046 = ~n830 & n840 ;
  assign n1047 = ~n1045 & ~n1046 ;
  assign n1061 = n465 & ~n474 ;
  assign n1062 = ~n465 & n474 ;
  assign n1063 = ~n1061 & ~n1062 ;
  assign n1114 = ~n1047 & ~n1063 ;
  assign n1068 = n476 & ~n486 ;
  assign n1069 = ~n476 & n486 ;
  assign n1070 = ~n1068 & ~n1069 ;
  assign n1074 = ~n405 & n414 ;
  assign n1075 = n405 & ~n414 ;
  assign n1076 = ~n1074 & ~n1075 ;
  assign n1115 = ~n1070 & ~n1076 ;
  assign n1116 = n1114 & n1115 ;
  assign n1036 = ~n582 & ~n583 ;
  assign n1037 = n281 & ~n690 ;
  assign n1038 = ~n281 & n690 ;
  assign n1039 = ~n1037 & ~n1038 ;
  assign n1096 = n1036 & ~n1039 ;
  assign n1041 = n862 & ~n871 ;
  assign n1042 = ~n862 & n871 ;
  assign n1043 = ~n1041 & ~n1042 ;
  assign n1044 = ~n384 & ~n388 ;
  assign n1097 = ~n1043 & n1044 ;
  assign n1104 = n1096 & n1097 ;
  assign n1028 = n671 & ~n679 ;
  assign n1029 = ~n671 & n679 ;
  assign n1030 = ~n1028 & ~n1029 ;
  assign n1031 = ~n709 & ~n727 ;
  assign n1094 = ~n1030 & n1031 ;
  assign n1032 = ~n772 & ~n965 ;
  assign n1033 = ~n628 & n635 ;
  assign n1034 = n628 & ~n635 ;
  assign n1035 = ~n1033 & ~n1034 ;
  assign n1095 = n1032 & ~n1035 ;
  assign n1105 = n1094 & n1095 ;
  assign n1112 = n1104 & n1105 ;
  assign n1065 = n718 & n725 ;
  assign n1066 = ~n718 & ~n725 ;
  assign n1067 = ~n1065 & ~n1066 ;
  assign n1077 = ~n531 & ~n532 ;
  assign n1100 = ~n1067 & n1077 ;
  assign n1085 = n515 & ~n522 ;
  assign n1086 = ~n515 & n522 ;
  assign n1087 = ~n1085 & ~n1086 ;
  assign n1091 = ~n743 & ~n774 ;
  assign n1101 = ~n1087 & n1091 ;
  assign n1102 = n1100 & n1101 ;
  assign n1051 = ~n878 & n887 ;
  assign n1052 = n878 & ~n887 ;
  assign n1053 = ~n1051 & ~n1052 ;
  assign n1054 = ~n592 & n601 ;
  assign n1055 = n592 & ~n601 ;
  assign n1056 = ~n1054 & ~n1055 ;
  assign n1098 = ~n1053 & ~n1056 ;
  assign n1057 = ~n619 & ~n638 ;
  assign n1064 = ~n760 & ~n761 ;
  assign n1099 = n1057 & n1064 ;
  assign n1103 = n1098 & n1099 ;
  assign n1113 = n1102 & n1103 ;
  assign n1117 = n1112 & n1113 ;
  assign n1121 = n1116 & n1117 ;
  assign n1122 = n1120 & n1121 ;
  assign n1124 = ~n932 & ~n1122 ;
  assign n1123 = n932 & n1122 ;
  assign n1125 = ~n935 & ~n1123 ;
  assign n1126 = ~n1124 & n1125 ;
  assign n1127 = n317 & ~n1126 ;
  assign n1128 = ~n1023 & ~n1127 ;
  assign n1129 = ~n325 & ~n1128 ;
  assign n1130 = ~n940 & ~n1003 ;
  assign n1131 = ~n317 & n932 ;
  assign n1132 = n935 & ~n1131 ;
  assign n1133 = ~n1130 & n1132 ;
  assign n1134 = ~n1129 & ~n1133 ;
  assign n1135 = ~n939 & n1134 ;
  assign n1136 = ~n1002 & n1135 ;
  assign n1137 = ~n1022 & n1136 ;
  assign n1138 = n311 & ~n1137 ;
  assign n1139 = ~n312 & ~n1138 ;
  assign n1140 = \IR_reg[31]/NET0131  & ~n235 ;
  assign n1141 = ~n319 & ~n1140 ;
  assign n1142 = \IR_reg[24]/NET0131  & ~n1141 ;
  assign n1143 = ~\IR_reg[24]/NET0131  & n1141 ;
  assign n1144 = ~n1142 & ~n1143 ;
  assign n1145 = \IR_reg[31]/NET0131  & ~n238 ;
  assign n1146 = ~n227 & ~n1145 ;
  assign n1147 = \IR_reg[26]/NET0131  & ~n1146 ;
  assign n1148 = ~\IR_reg[26]/NET0131  & n1146 ;
  assign n1149 = ~n1147 & ~n1148 ;
  assign n1150 = ~n1144 & ~n1149 ;
  assign n1151 = ~\IR_reg[24]/NET0131  & n234 ;
  assign n1152 = n252 & n1151 ;
  assign n1153 = \IR_reg[31]/NET0131  & ~n1152 ;
  assign n1154 = ~n313 & ~n1153 ;
  assign n1155 = \IR_reg[25]/NET0131  & ~n1154 ;
  assign n1156 = ~\IR_reg[25]/NET0131  & n1154 ;
  assign n1157 = ~n1155 & ~n1156 ;
  assign n1158 = \B_reg/NET0131  & ~n1144 ;
  assign n1159 = ~\B_reg/NET0131  & n1144 ;
  assign n1160 = ~n1158 & ~n1159 ;
  assign n1161 = ~n1157 & ~n1160 ;
  assign n1162 = ~\d_reg[0]/NET0131  & n1149 ;
  assign n1163 = ~n1161 & n1162 ;
  assign n1164 = ~n1150 & ~n1163 ;
  assign n1165 = ~\d_reg[1]/NET0131  & n1149 ;
  assign n1166 = ~n1161 & n1165 ;
  assign n1167 = ~n1149 & ~n1157 ;
  assign n1168 = ~n1166 & ~n1167 ;
  assign n1169 = n1164 & n1168 ;
  assign n1170 = n397 & ~n1169 ;
  assign n1171 = n961 & ~n981 ;
  assign n1172 = n954 & n962 ;
  assign n1173 = ~n1171 & n1172 ;
  assign n1174 = ~n560 & n954 ;
  assign n1175 = n949 & ~n1174 ;
  assign n1176 = ~n1173 & n1175 ;
  assign n1177 = n951 & n988 ;
  assign n1178 = ~n1176 & n1177 ;
  assign n1179 = ~n901 & n988 ;
  assign n1180 = ~n994 & ~n1179 ;
  assign n1181 = ~n1178 & n1180 ;
  assign n1182 = n1073 & ~n1181 ;
  assign n1183 = ~n1073 & n1181 ;
  assign n1184 = ~n1182 & ~n1183 ;
  assign n1185 = n1169 & ~n1184 ;
  assign n1186 = ~n1170 & ~n1185 ;
  assign n1187 = n310 & n325 ;
  assign n1188 = n310 & ~n932 ;
  assign n1189 = ~n1003 & ~n1188 ;
  assign n1190 = ~n1187 & ~n1189 ;
  assign n1191 = ~n1186 & n1190 ;
  assign n1192 = n298 & n530 ;
  assign n1193 = ~n1024 & ~n1192 ;
  assign n1194 = n498 & n504 ;
  assign n1195 = ~n1085 & ~n1194 ;
  assign n1196 = n1193 & n1195 ;
  assign n1197 = ~n1041 & ~n1051 ;
  assign n1198 = n797 & n806 ;
  assign n1199 = ~n1089 & ~n1198 ;
  assign n1200 = n1197 & n1199 ;
  assign n1201 = n1196 & n1200 ;
  assign n1202 = n572 & n581 ;
  assign n1203 = ~n1055 & ~n1202 ;
  assign n1204 = ~n609 & ~n618 ;
  assign n1205 = n609 & n618 ;
  assign n1206 = n1033 & ~n1205 ;
  assign n1207 = ~n1204 & ~n1206 ;
  assign n1208 = n1203 & ~n1207 ;
  assign n1209 = ~n572 & ~n581 ;
  assign n1210 = ~n1054 & ~n1209 ;
  assign n1211 = ~n1202 & ~n1210 ;
  assign n1212 = ~n1208 & ~n1211 ;
  assign n1213 = n652 & n661 ;
  assign n1214 = ~n1028 & ~n1213 ;
  assign n1215 = n699 & n708 ;
  assign n1216 = ~n1037 & ~n1215 ;
  assign n1217 = ~n752 & ~n759 ;
  assign n1218 = ~n768 & ~n771 ;
  assign n1219 = n752 & n759 ;
  assign n1220 = n1218 & ~n1219 ;
  assign n1221 = ~n1217 & ~n1220 ;
  assign n1222 = n735 & n742 ;
  assign n1223 = ~n1065 & ~n1222 ;
  assign n1224 = ~n1221 & n1223 ;
  assign n1225 = ~n735 & ~n742 ;
  assign n1226 = ~n1066 & ~n1225 ;
  assign n1227 = ~n1065 & ~n1226 ;
  assign n1228 = ~n1224 & ~n1227 ;
  assign n1229 = n1216 & ~n1228 ;
  assign n1230 = n1214 & n1229 ;
  assign n1231 = ~n699 & ~n708 ;
  assign n1232 = ~n1037 & n1231 ;
  assign n1233 = ~n1038 & ~n1232 ;
  assign n1234 = n1214 & ~n1233 ;
  assign n1235 = ~n652 & ~n661 ;
  assign n1236 = ~n1028 & n1235 ;
  assign n1237 = ~n1029 & ~n1236 ;
  assign n1238 = ~n1234 & n1237 ;
  assign n1239 = ~n1230 & n1238 ;
  assign n1240 = ~n1034 & ~n1205 ;
  assign n1241 = n1203 & n1240 ;
  assign n1242 = ~n1239 & n1241 ;
  assign n1243 = n1212 & ~n1242 ;
  assign n1244 = n1201 & ~n1243 ;
  assign n1245 = ~n298 & ~n530 ;
  assign n1246 = n1025 & ~n1192 ;
  assign n1247 = ~n1245 & ~n1246 ;
  assign n1248 = n1195 & ~n1247 ;
  assign n1249 = ~n498 & ~n504 ;
  assign n1250 = ~n1085 & n1249 ;
  assign n1251 = ~n1086 & ~n1250 ;
  assign n1252 = ~n1248 & n1251 ;
  assign n1253 = n1200 & ~n1252 ;
  assign n1254 = ~n1042 & ~n1052 ;
  assign n1255 = ~n1041 & ~n1254 ;
  assign n1256 = n1199 & n1255 ;
  assign n1257 = ~n797 & ~n806 ;
  assign n1258 = n1088 & ~n1198 ;
  assign n1259 = ~n1257 & ~n1258 ;
  assign n1260 = ~n1256 & n1259 ;
  assign n1261 = ~n1253 & n1260 ;
  assign n1262 = ~n1244 & n1261 ;
  assign n1263 = ~n1059 & ~n1074 ;
  assign n1264 = ~n1078 & n1263 ;
  assign n1265 = ~n1049 & n1264 ;
  assign n1266 = ~n1046 & ~n1069 ;
  assign n1267 = ~n1083 & n1266 ;
  assign n1268 = ~n1062 & n1267 ;
  assign n1269 = n1265 & n1268 ;
  assign n1270 = ~n1262 & n1269 ;
  assign n1275 = ~n1061 & ~n1068 ;
  assign n1276 = ~n1046 & n1082 ;
  assign n1277 = ~n1045 & ~n1276 ;
  assign n1278 = ~n1069 & ~n1277 ;
  assign n1279 = n1275 & ~n1278 ;
  assign n1280 = ~n1062 & ~n1279 ;
  assign n1281 = n1265 & n1280 ;
  assign n1271 = n1048 & ~n1078 ;
  assign n1272 = ~n1079 & ~n1271 ;
  assign n1273 = ~n1058 & n1272 ;
  assign n1274 = n1263 & ~n1273 ;
  assign n1282 = ~n1075 & ~n1274 ;
  assign n1283 = ~n1281 & n1282 ;
  assign n1284 = ~n1270 & n1283 ;
  assign n1285 = n1073 & n1284 ;
  assign n1286 = ~n1073 & ~n1284 ;
  assign n1287 = ~n1285 & ~n1286 ;
  assign n1288 = n1169 & ~n1287 ;
  assign n1289 = ~n1170 & ~n1288 ;
  assign n1290 = ~n310 & ~n325 ;
  assign n1291 = ~n1187 & ~n1290 ;
  assign n1292 = n1189 & n1291 ;
  assign n1293 = ~n1289 & n1292 ;
  assign n1294 = n759 & n771 ;
  assign n1295 = n742 & n1294 ;
  assign n1296 = n725 & n1295 ;
  assign n1297 = n699 & n1296 ;
  assign n1298 = ~n690 & n1297 ;
  assign n1299 = n652 & ~n679 ;
  assign n1300 = n1298 & n1299 ;
  assign n1301 = n609 & ~n635 ;
  assign n1302 = n1300 & n1301 ;
  assign n1303 = n530 & ~n551 ;
  assign n1304 = n572 & ~n601 ;
  assign n1305 = n1303 & n1304 ;
  assign n1306 = n1302 & n1305 ;
  assign n1307 = n504 & ~n522 ;
  assign n1308 = ~n878 & n1307 ;
  assign n1309 = ~n871 & n1308 ;
  assign n1310 = n1306 & n1309 ;
  assign n1311 = n797 & ~n842 ;
  assign n1312 = ~n817 & n1311 ;
  assign n1313 = n1310 & n1312 ;
  assign n1314 = ~n428 & ~n465 ;
  assign n1315 = ~n476 & ~n830 ;
  assign n1316 = n1314 & n1315 ;
  assign n1317 = n1313 & n1316 ;
  assign n1318 = ~n417 & ~n445 ;
  assign n1319 = n1317 & n1318 ;
  assign n1320 = ~n405 & n1319 ;
  assign n1321 = n389 & ~n1320 ;
  assign n1322 = ~n389 & n1320 ;
  assign n1323 = ~n1321 & ~n1322 ;
  assign n1324 = n1169 & n1323 ;
  assign n1325 = ~n1170 & ~n1324 ;
  assign n1326 = n1131 & n1290 ;
  assign n1327 = ~n1325 & n1326 ;
  assign n1334 = ~n364 & ~n768 ;
  assign n1335 = ~n752 & n1334 ;
  assign n1336 = ~n735 & n1335 ;
  assign n1337 = ~n718 & n1336 ;
  assign n1338 = ~n281 & ~n708 ;
  assign n1339 = n1337 & n1338 ;
  assign n1340 = ~n661 & ~n671 ;
  assign n1341 = n1339 & n1340 ;
  assign n1342 = ~n581 & ~n592 ;
  assign n1343 = ~n618 & ~n628 ;
  assign n1344 = n1342 & n1343 ;
  assign n1345 = n1341 & n1344 ;
  assign n1346 = ~n298 & ~n515 ;
  assign n1347 = ~n541 & n1346 ;
  assign n1348 = ~n498 & n1347 ;
  assign n1349 = n1345 & n1348 ;
  assign n1350 = ~n862 & ~n887 ;
  assign n1351 = ~n806 & n1350 ;
  assign n1352 = ~n827 & n1351 ;
  assign n1353 = n1349 & n1352 ;
  assign n1354 = ~n486 & ~n840 ;
  assign n1355 = ~n474 & ~n851 ;
  assign n1356 = n1354 & n1355 ;
  assign n1357 = ~n426 & ~n441 ;
  assign n1358 = n1356 & n1357 ;
  assign n1359 = ~n414 & ~n454 ;
  assign n1360 = ~n401 & n1359 ;
  assign n1361 = n1358 & n1360 ;
  assign n1362 = n1353 & n1361 ;
  assign n1363 = n383 & ~n1362 ;
  assign n1364 = ~n383 & n1362 ;
  assign n1365 = ~n1363 & ~n1364 ;
  assign n1366 = ~n338 & ~n1365 ;
  assign n1367 = n338 & n414 ;
  assign n1368 = ~n1366 & ~n1367 ;
  assign n1369 = n325 & n1131 ;
  assign n1370 = n310 & n1369 ;
  assign n1371 = n1368 & n1370 ;
  assign n1372 = n1169 & n1371 ;
  assign n1328 = n317 & n1290 ;
  assign n1329 = n1169 & n1328 ;
  assign n1330 = ~n310 & ~n932 ;
  assign n1331 = n940 & n1330 ;
  assign n1332 = ~n1329 & ~n1331 ;
  assign n1333 = n389 & ~n1332 ;
  assign n1373 = ~n1131 & n1187 ;
  assign n1374 = ~n1169 & n1328 ;
  assign n1375 = ~n1373 & ~n1374 ;
  assign n1376 = ~n1169 & n1370 ;
  assign n1377 = n1375 & ~n1376 ;
  assign n1378 = n397 & ~n1377 ;
  assign n1379 = ~n1333 & ~n1378 ;
  assign n1380 = ~n1372 & n1379 ;
  assign n1381 = ~n1327 & n1380 ;
  assign n1382 = ~n1293 & n1381 ;
  assign n1383 = ~n1191 & n1382 ;
  assign n1384 = n1144 & n1149 ;
  assign n1385 = n1157 & n1384 ;
  assign n1386 = ~n310 & ~n1385 ;
  assign n1387 = ~n1383 & n1386 ;
  assign n1388 = ~n310 & n1385 ;
  assign n1389 = n397 & n1388 ;
  assign n1390 = ~n1387 & ~n1389 ;
  assign n1391 = \state_reg[0]/NET0131  & ~n1390 ;
  assign n1392 = \reg3_reg[28]/NET0131  & ~\state_reg[0]/NET0131  ;
  assign n1393 = n311 & n397 ;
  assign n1394 = ~n1392 & ~n1393 ;
  assign n1395 = ~n1391 & n1394 ;
  assign n1396 = ~n1164 & n1168 ;
  assign n1397 = \reg2_reg[28]/NET0131  & ~n1396 ;
  assign n1398 = ~n1184 & n1396 ;
  assign n1399 = ~n1397 & ~n1398 ;
  assign n1400 = n1190 & ~n1399 ;
  assign n1401 = ~n1287 & n1396 ;
  assign n1402 = ~n1397 & ~n1401 ;
  assign n1403 = n1292 & ~n1402 ;
  assign n1404 = n1323 & n1396 ;
  assign n1405 = ~n1397 & ~n1404 ;
  assign n1406 = n1326 & ~n1405 ;
  assign n1407 = n1368 & n1396 ;
  assign n1408 = ~n1397 & ~n1407 ;
  assign n1409 = n1370 & ~n1408 ;
  assign n1413 = n1328 & ~n1396 ;
  assign n1414 = ~n1373 & ~n1413 ;
  assign n1415 = \reg2_reg[28]/NET0131  & ~n1414 ;
  assign n1410 = n397 & n1331 ;
  assign n1411 = n389 & n1328 ;
  assign n1412 = n1396 & n1411 ;
  assign n1416 = ~n1410 & ~n1412 ;
  assign n1417 = ~n1415 & n1416 ;
  assign n1418 = ~n1409 & n1417 ;
  assign n1419 = ~n1406 & n1418 ;
  assign n1420 = ~n1403 & n1419 ;
  assign n1421 = ~n1400 & n1420 ;
  assign n1422 = n1386 & ~n1421 ;
  assign n1423 = \reg2_reg[28]/NET0131  & n1388 ;
  assign n1424 = ~n1422 & ~n1423 ;
  assign n1425 = \state_reg[0]/NET0131  & ~n1424 ;
  assign n1426 = \state_reg[0]/NET0131  & ~n310 ;
  assign n1427 = \reg2_reg[28]/NET0131  & ~n1426 ;
  assign n1428 = ~n1425 & ~n1427 ;
  assign n1429 = \reg2_reg[29]/NET0131  & ~n1426 ;
  assign n1430 = \reg2_reg[29]/NET0131  & n1388 ;
  assign n1431 = \reg2_reg[29]/NET0131  & ~n1396 ;
  assign n1432 = n377 & ~n1322 ;
  assign n1433 = ~n377 & n1322 ;
  assign n1434 = ~n1432 & ~n1433 ;
  assign n1435 = n1396 & n1434 ;
  assign n1436 = ~n1431 & ~n1435 ;
  assign n1437 = n1326 & ~n1436 ;
  assign n1438 = n338 & ~n401 ;
  assign n1439 = n373 & ~n1364 ;
  assign n1440 = ~n373 & n1364 ;
  assign n1441 = \B_reg/NET0131  & n332 ;
  assign n1442 = ~n338 & ~n1441 ;
  assign n1443 = ~n1440 & n1442 ;
  assign n1444 = ~n1439 & n1443 ;
  assign n1445 = ~n1438 & ~n1444 ;
  assign n1446 = n1396 & ~n1445 ;
  assign n1447 = ~n1431 & ~n1446 ;
  assign n1448 = n1370 & ~n1447 ;
  assign n1452 = \reg2_reg[29]/NET0131  & ~n1414 ;
  assign n1449 = n357 & n1331 ;
  assign n1450 = n377 & n1328 ;
  assign n1451 = n1396 & n1450 ;
  assign n1596 = ~n1449 & ~n1451 ;
  assign n1597 = ~n1452 & n1596 ;
  assign n1598 = ~n1448 & n1597 ;
  assign n1599 = ~n1437 & n1598 ;
  assign n1453 = ~n1192 & ~n1194 ;
  assign n1454 = ~n1051 & ~n1085 ;
  assign n1455 = n1453 & n1454 ;
  assign n1456 = ~n1041 & ~n1089 ;
  assign n1457 = ~n1083 & ~n1198 ;
  assign n1458 = n1456 & n1457 ;
  assign n1459 = n1455 & n1458 ;
  assign n1460 = ~n1024 & ~n1202 ;
  assign n1461 = ~n1055 & n1204 ;
  assign n1462 = ~n1054 & ~n1461 ;
  assign n1463 = n1460 & ~n1462 ;
  assign n1464 = ~n1024 & n1209 ;
  assign n1465 = ~n1025 & ~n1464 ;
  assign n1466 = ~n1463 & n1465 ;
  assign n1467 = ~n1028 & ~n1034 ;
  assign n1468 = ~n1217 & ~n1225 ;
  assign n1469 = ~n1220 & n1468 ;
  assign n1470 = n1223 & ~n1469 ;
  assign n1471 = ~n1066 & ~n1231 ;
  assign n1472 = ~n1470 & n1471 ;
  assign n1473 = ~n1213 & n1216 ;
  assign n1474 = ~n1472 & n1473 ;
  assign n1475 = n1467 & n1474 ;
  assign n1476 = n1038 & ~n1213 ;
  assign n1477 = ~n1235 & ~n1476 ;
  assign n1478 = n1467 & ~n1477 ;
  assign n1479 = n1029 & ~n1034 ;
  assign n1480 = ~n1033 & ~n1479 ;
  assign n1481 = ~n1478 & n1480 ;
  assign n1482 = ~n1475 & n1481 ;
  assign n1483 = ~n1055 & ~n1205 ;
  assign n1484 = n1460 & n1483 ;
  assign n1485 = ~n1482 & n1484 ;
  assign n1486 = n1466 & ~n1485 ;
  assign n1487 = n1459 & ~n1486 ;
  assign n1488 = ~n1194 & n1245 ;
  assign n1489 = ~n1249 & ~n1488 ;
  assign n1490 = n1454 & ~n1489 ;
  assign n1491 = ~n1052 & ~n1086 ;
  assign n1492 = ~n1051 & ~n1491 ;
  assign n1493 = ~n1490 & ~n1492 ;
  assign n1494 = n1458 & ~n1493 ;
  assign n1495 = ~n1082 & ~n1257 ;
  assign n1496 = n1042 & ~n1089 ;
  assign n1497 = ~n1088 & ~n1496 ;
  assign n1498 = ~n1198 & ~n1497 ;
  assign n1499 = n1495 & ~n1498 ;
  assign n1500 = ~n1083 & ~n1499 ;
  assign n1501 = ~n1494 & ~n1500 ;
  assign n1502 = ~n1487 & n1501 ;
  assign n1503 = ~n1071 & n1264 ;
  assign n1504 = ~n1049 & ~n1062 ;
  assign n1505 = n1266 & n1504 ;
  assign n1506 = n1503 & n1505 ;
  assign n1507 = ~n1502 & n1506 ;
  assign n1512 = n1045 & ~n1069 ;
  assign n1513 = ~n1068 & ~n1512 ;
  assign n1514 = n1504 & ~n1513 ;
  assign n1515 = ~n1049 & n1061 ;
  assign n1516 = ~n1048 & ~n1515 ;
  assign n1517 = ~n1514 & n1516 ;
  assign n1518 = n1503 & ~n1517 ;
  assign n1508 = ~n1058 & ~n1079 ;
  assign n1509 = n1263 & ~n1508 ;
  assign n1510 = ~n1075 & ~n1509 ;
  assign n1511 = ~n1071 & ~n1510 ;
  assign n1519 = ~n1072 & ~n1511 ;
  assign n1520 = ~n1518 & n1519 ;
  assign n1521 = ~n1507 & n1520 ;
  assign n1522 = ~n1044 & n1521 ;
  assign n1523 = n1044 & ~n1521 ;
  assign n1524 = ~n1522 & ~n1523 ;
  assign n1525 = n1396 & ~n1524 ;
  assign n1526 = ~n1431 & ~n1525 ;
  assign n1527 = n1292 & ~n1526 ;
  assign n1528 = ~n602 & ~n619 ;
  assign n1529 = ~n561 & ~n583 ;
  assign n1530 = n1528 & n1529 ;
  assign n1531 = ~n636 & ~n680 ;
  assign n1532 = ~n774 & ~n967 ;
  assign n1533 = ~n709 & n745 ;
  assign n1534 = ~n1532 & n1533 ;
  assign n1535 = ~n709 & ~n728 ;
  assign n1536 = ~n1534 & ~n1535 ;
  assign n1537 = ~n662 & ~n710 ;
  assign n1538 = ~n1536 & n1537 ;
  assign n1539 = n1531 & n1538 ;
  assign n1540 = n1530 & n1539 ;
  assign n1541 = ~n662 & ~n693 ;
  assign n1542 = n1531 & n1541 ;
  assign n1543 = ~n636 & ~n784 ;
  assign n1544 = ~n1542 & ~n1543 ;
  assign n1545 = n1530 & ~n1544 ;
  assign n1546 = ~n602 & ~n640 ;
  assign n1547 = n1529 & n1546 ;
  assign n1548 = ~n561 & ~n785 ;
  assign n1549 = ~n1547 & ~n1548 ;
  assign n1550 = ~n1545 & n1549 ;
  assign n1551 = ~n1540 & n1550 ;
  assign n1552 = ~n902 & ~n912 ;
  assign n1553 = ~n903 & ~n905 ;
  assign n1554 = n1552 & n1553 ;
  assign n1555 = ~n505 & ~n531 ;
  assign n1556 = ~n523 & ~n906 ;
  assign n1557 = n1555 & n1556 ;
  assign n1558 = n1554 & n1557 ;
  assign n1559 = ~n1551 & n1558 ;
  assign n1560 = ~n505 & ~n563 ;
  assign n1561 = n1556 & n1560 ;
  assign n1562 = n557 & ~n906 ;
  assign n1563 = ~n888 & ~n1562 ;
  assign n1564 = ~n1561 & n1563 ;
  assign n1565 = n1554 & ~n1564 ;
  assign n1566 = ~n807 & ~n852 ;
  assign n1567 = ~n903 & ~n908 ;
  assign n1568 = ~n902 & n1567 ;
  assign n1569 = n1566 & ~n1568 ;
  assign n1570 = ~n912 & ~n1569 ;
  assign n1571 = ~n1565 & ~n1570 ;
  assign n1572 = ~n1559 & n1571 ;
  assign n1573 = ~n442 & ~n895 ;
  assign n1574 = n913 & n1573 ;
  assign n1575 = ~n402 & n987 ;
  assign n1576 = n1574 & n1575 ;
  assign n1577 = ~n1572 & n1576 ;
  assign n1578 = ~n487 & ~n915 ;
  assign n1579 = n1573 & ~n1578 ;
  assign n1580 = ~n442 & n475 ;
  assign n1581 = ~n922 & ~n1580 ;
  assign n1582 = ~n1579 & n1581 ;
  assign n1583 = n987 & ~n1582 ;
  assign n1584 = ~n456 & ~n459 ;
  assign n1585 = ~n458 & n1584 ;
  assign n1586 = n416 & ~n1585 ;
  assign n1587 = ~n1583 & n1586 ;
  assign n1588 = ~n402 & ~n1587 ;
  assign n1589 = ~n1577 & ~n1588 ;
  assign n1590 = ~n1044 & n1589 ;
  assign n1591 = n1044 & ~n1589 ;
  assign n1592 = ~n1590 & ~n1591 ;
  assign n1593 = n1396 & n1592 ;
  assign n1594 = ~n1431 & ~n1593 ;
  assign n1595 = n1190 & ~n1594 ;
  assign n1600 = ~n1527 & ~n1595 ;
  assign n1601 = n1599 & n1600 ;
  assign n1602 = n1386 & ~n1601 ;
  assign n1603 = ~n1430 & ~n1602 ;
  assign n1604 = \state_reg[0]/NET0131  & ~n1603 ;
  assign n1605 = ~n1429 & ~n1604 ;
  assign n1606 = \reg0_reg[28]/NET0131  & ~n1426 ;
  assign n1607 = ~n1164 & ~n1168 ;
  assign n1608 = \reg0_reg[28]/NET0131  & ~n1607 ;
  assign n1609 = ~n1184 & n1607 ;
  assign n1610 = ~n1608 & ~n1609 ;
  assign n1611 = n1190 & ~n1610 ;
  assign n1612 = ~n1287 & n1607 ;
  assign n1613 = ~n1608 & ~n1612 ;
  assign n1614 = n1292 & ~n1613 ;
  assign n1615 = n1323 & n1326 ;
  assign n1616 = ~n1371 & ~n1411 ;
  assign n1617 = ~n1615 & n1616 ;
  assign n1618 = n1607 & ~n1617 ;
  assign n1619 = n1370 & ~n1607 ;
  assign n1620 = ~n1331 & ~n1373 ;
  assign n1621 = ~n1326 & ~n1328 ;
  assign n1622 = ~n1607 & ~n1621 ;
  assign n1623 = n1620 & ~n1622 ;
  assign n1624 = ~n1619 & n1623 ;
  assign n1625 = \reg0_reg[28]/NET0131  & ~n1624 ;
  assign n1626 = ~n1618 & ~n1625 ;
  assign n1627 = ~n1614 & n1626 ;
  assign n1628 = ~n1611 & n1627 ;
  assign n1629 = n1386 & ~n1628 ;
  assign n1630 = \reg0_reg[28]/NET0131  & n1388 ;
  assign n1631 = ~n1629 & ~n1630 ;
  assign n1632 = \state_reg[0]/NET0131  & ~n1631 ;
  assign n1633 = ~n1606 & ~n1632 ;
  assign n1634 = \reg1_reg[28]/NET0131  & ~n1426 ;
  assign n1635 = n1164 & ~n1168 ;
  assign n1636 = \reg1_reg[28]/NET0131  & ~n1635 ;
  assign n1637 = ~n1184 & n1635 ;
  assign n1638 = ~n1636 & ~n1637 ;
  assign n1639 = n1190 & ~n1638 ;
  assign n1640 = ~n1287 & n1635 ;
  assign n1641 = ~n1636 & ~n1640 ;
  assign n1642 = n1292 & ~n1641 ;
  assign n1643 = ~n1617 & n1635 ;
  assign n1644 = n1370 & ~n1635 ;
  assign n1645 = ~n1621 & ~n1635 ;
  assign n1646 = n1620 & ~n1645 ;
  assign n1647 = ~n1644 & n1646 ;
  assign n1648 = \reg1_reg[28]/NET0131  & ~n1647 ;
  assign n1649 = ~n1643 & ~n1648 ;
  assign n1650 = ~n1642 & n1649 ;
  assign n1651 = ~n1639 & n1650 ;
  assign n1652 = n1386 & ~n1651 ;
  assign n1653 = \reg1_reg[28]/NET0131  & n1388 ;
  assign n1654 = ~n1652 & ~n1653 ;
  assign n1655 = \state_reg[0]/NET0131  & ~n1654 ;
  assign n1656 = ~n1634 & ~n1655 ;
  assign n1660 = n508 & ~n1169 ;
  assign n1661 = n1548 & n1555 ;
  assign n1662 = ~n1560 & ~n1661 ;
  assign n1663 = n1529 & n1555 ;
  assign n1664 = ~n1538 & ~n1541 ;
  assign n1665 = n1528 & n1531 ;
  assign n1666 = ~n1664 & n1665 ;
  assign n1667 = n1528 & n1543 ;
  assign n1668 = ~n1546 & ~n1667 ;
  assign n1669 = ~n1666 & n1668 ;
  assign n1670 = n1663 & ~n1669 ;
  assign n1671 = n1662 & ~n1670 ;
  assign n1672 = n1087 & n1671 ;
  assign n1673 = ~n1087 & ~n1671 ;
  assign n1674 = ~n1672 & ~n1673 ;
  assign n1675 = n1169 & n1674 ;
  assign n1676 = ~n1660 & ~n1675 ;
  assign n1677 = n1190 & ~n1676 ;
  assign n1678 = ~n1474 & n1477 ;
  assign n1679 = n1467 & n1483 ;
  assign n1680 = ~n1678 & n1679 ;
  assign n1681 = ~n1480 & n1483 ;
  assign n1682 = n1462 & ~n1681 ;
  assign n1683 = ~n1680 & n1682 ;
  assign n1684 = n1453 & n1460 ;
  assign n1685 = ~n1683 & n1684 ;
  assign n1686 = n1453 & ~n1465 ;
  assign n1687 = n1489 & ~n1686 ;
  assign n1688 = ~n1685 & n1687 ;
  assign n1689 = n1087 & n1688 ;
  assign n1690 = ~n1087 & ~n1688 ;
  assign n1691 = ~n1689 & ~n1690 ;
  assign n1692 = n1169 & ~n1691 ;
  assign n1693 = ~n1660 & ~n1692 ;
  assign n1694 = n1292 & ~n1693 ;
  assign n1695 = ~n887 & n1349 ;
  assign n1696 = n887 & ~n1349 ;
  assign n1697 = ~n1695 & ~n1696 ;
  assign n1698 = ~n338 & ~n1697 ;
  assign n1699 = n338 & n498 ;
  assign n1700 = ~n1698 & ~n1699 ;
  assign n1701 = n1169 & n1700 ;
  assign n1702 = ~n1660 & ~n1701 ;
  assign n1703 = n1370 & ~n1702 ;
  assign n1704 = n504 & n1306 ;
  assign n1705 = n522 & ~n1704 ;
  assign n1706 = ~n522 & n1704 ;
  assign n1707 = ~n1705 & ~n1706 ;
  assign n1708 = n1169 & n1707 ;
  assign n1709 = ~n1660 & ~n1708 ;
  assign n1710 = n1326 & ~n1709 ;
  assign n1659 = n522 & ~n1332 ;
  assign n1711 = n508 & ~n1375 ;
  assign n1712 = ~n1659 & ~n1711 ;
  assign n1713 = ~n1710 & n1712 ;
  assign n1714 = ~n1703 & n1713 ;
  assign n1715 = ~n1694 & n1714 ;
  assign n1716 = ~n1677 & n1715 ;
  assign n1717 = \state_reg[0]/NET0131  & n1386 ;
  assign n1718 = ~n1716 & n1717 ;
  assign n1657 = \state_reg[0]/NET0131  & ~n1386 ;
  assign n1658 = n508 & n1657 ;
  assign n1719 = \reg3_reg[15]/NET0131  & ~\state_reg[0]/NET0131  ;
  assign n1720 = ~n1658 & ~n1719 ;
  assign n1721 = ~n1718 & n1720 ;
  assign n1722 = \reg2_reg[27]/NET0131  & ~n1396 ;
  assign n1723 = n1267 & ~n1495 ;
  assign n1724 = n1513 & ~n1723 ;
  assign n1725 = n1504 & ~n1724 ;
  assign n1726 = n1516 & ~n1725 ;
  assign n1727 = ~n1078 & ~n1726 ;
  assign n1728 = n1508 & ~n1727 ;
  assign n1729 = ~n1059 & ~n1728 ;
  assign n1730 = n1454 & n1456 ;
  assign n1731 = ~n1688 & n1730 ;
  assign n1732 = n1456 & n1492 ;
  assign n1733 = n1497 & ~n1732 ;
  assign n1734 = ~n1731 & n1733 ;
  assign n1736 = ~n1078 & n1504 ;
  assign n1735 = ~n1198 & n1267 ;
  assign n1737 = ~n1059 & n1735 ;
  assign n1738 = n1736 & n1737 ;
  assign n1739 = ~n1734 & n1738 ;
  assign n1740 = ~n1729 & ~n1739 ;
  assign n1741 = n1076 & n1740 ;
  assign n1742 = ~n1076 & ~n1740 ;
  assign n1743 = ~n1741 & ~n1742 ;
  assign n1744 = n1396 & ~n1743 ;
  assign n1745 = ~n1722 & ~n1744 ;
  assign n1746 = n1292 & ~n1745 ;
  assign n1752 = n1553 & n1556 ;
  assign n1753 = n1663 & n1752 ;
  assign n1754 = ~n1669 & n1753 ;
  assign n1755 = ~n1662 & n1752 ;
  assign n1756 = n1553 & ~n1563 ;
  assign n1757 = ~n1567 & ~n1756 ;
  assign n1758 = ~n1755 & n1757 ;
  assign n1759 = ~n1754 & n1758 ;
  assign n1760 = n986 & n1552 ;
  assign n1761 = n1574 & n1760 ;
  assign n1762 = ~n1759 & n1761 ;
  assign n1747 = n914 & ~n1566 ;
  assign n1748 = n1578 & ~n1747 ;
  assign n1749 = n1573 & ~n1748 ;
  assign n1750 = n1581 & ~n1749 ;
  assign n1751 = n986 & ~n1750 ;
  assign n1763 = ~n1584 & ~n1751 ;
  assign n1764 = ~n1762 & n1763 ;
  assign n1765 = n1076 & ~n1764 ;
  assign n1766 = ~n1076 & n1764 ;
  assign n1767 = ~n1765 & ~n1766 ;
  assign n1768 = n1396 & ~n1767 ;
  assign n1769 = ~n1722 & ~n1768 ;
  assign n1770 = n1190 & ~n1769 ;
  assign n1771 = n1353 & n1358 ;
  assign n1772 = n1359 & n1771 ;
  assign n1773 = n401 & ~n1772 ;
  assign n1774 = ~n1362 & ~n1773 ;
  assign n1775 = ~n338 & ~n1774 ;
  assign n1776 = n338 & n454 ;
  assign n1777 = ~n1775 & ~n1776 ;
  assign n1778 = n1396 & n1777 ;
  assign n1779 = ~n1722 & ~n1778 ;
  assign n1780 = n1370 & ~n1779 ;
  assign n1781 = n405 & ~n1319 ;
  assign n1782 = ~n1320 & ~n1781 ;
  assign n1783 = n1396 & n1782 ;
  assign n1784 = ~n1722 & ~n1783 ;
  assign n1785 = n1326 & ~n1784 ;
  assign n1789 = \reg2_reg[27]/NET0131  & ~n1414 ;
  assign n1786 = n410 & n1331 ;
  assign n1787 = n405 & n1328 ;
  assign n1788 = n1396 & n1787 ;
  assign n1790 = ~n1786 & ~n1788 ;
  assign n1791 = ~n1789 & n1790 ;
  assign n1792 = ~n1785 & n1791 ;
  assign n1793 = ~n1780 & n1792 ;
  assign n1794 = ~n1770 & n1793 ;
  assign n1795 = ~n1746 & n1794 ;
  assign n1796 = n1386 & ~n1795 ;
  assign n1797 = \reg2_reg[27]/NET0131  & n1388 ;
  assign n1798 = ~n1796 & ~n1797 ;
  assign n1799 = \state_reg[0]/NET0131  & ~n1798 ;
  assign n1800 = \reg2_reg[27]/NET0131  & ~n1426 ;
  assign n1801 = ~n1799 & ~n1800 ;
  assign n1802 = \reg0_reg[27]/NET0131  & ~n1426 ;
  assign n1803 = \reg0_reg[27]/NET0131  & ~n1607 ;
  assign n1804 = n1607 & ~n1743 ;
  assign n1805 = ~n1803 & ~n1804 ;
  assign n1806 = n1292 & ~n1805 ;
  assign n1807 = n1607 & ~n1767 ;
  assign n1808 = ~n1803 & ~n1807 ;
  assign n1809 = n1190 & ~n1808 ;
  assign n1810 = n1370 & n1777 ;
  assign n1811 = n1326 & n1782 ;
  assign n1812 = ~n1787 & ~n1811 ;
  assign n1813 = ~n1810 & n1812 ;
  assign n1814 = n1607 & ~n1813 ;
  assign n1815 = \reg0_reg[27]/NET0131  & ~n1624 ;
  assign n1816 = ~n1814 & ~n1815 ;
  assign n1817 = ~n1809 & n1816 ;
  assign n1818 = ~n1806 & n1817 ;
  assign n1819 = n1386 & ~n1818 ;
  assign n1820 = \reg0_reg[27]/NET0131  & n1388 ;
  assign n1821 = ~n1819 & ~n1820 ;
  assign n1822 = \state_reg[0]/NET0131  & ~n1821 ;
  assign n1823 = ~n1802 & ~n1822 ;
  assign n1824 = \reg0_reg[29]/NET0131  & ~n1426 ;
  assign n1825 = \reg0_reg[29]/NET0131  & n1388 ;
  assign n1826 = n1326 & n1434 ;
  assign n1827 = ~n1450 & ~n1826 ;
  assign n1828 = n1607 & ~n1827 ;
  assign n1829 = \reg0_reg[29]/NET0131  & ~n1607 ;
  assign n1830 = ~n1445 & n1607 ;
  assign n1831 = ~n1829 & ~n1830 ;
  assign n1832 = n1370 & ~n1831 ;
  assign n1833 = \reg0_reg[29]/NET0131  & ~n1623 ;
  assign n1840 = ~n1832 & ~n1833 ;
  assign n1841 = ~n1828 & n1840 ;
  assign n1834 = ~n1524 & n1607 ;
  assign n1835 = ~n1829 & ~n1834 ;
  assign n1836 = n1292 & ~n1835 ;
  assign n1837 = n1592 & n1607 ;
  assign n1838 = ~n1829 & ~n1837 ;
  assign n1839 = n1190 & ~n1838 ;
  assign n1842 = ~n1836 & ~n1839 ;
  assign n1843 = n1841 & n1842 ;
  assign n1844 = n1386 & ~n1843 ;
  assign n1845 = ~n1825 & ~n1844 ;
  assign n1846 = \state_reg[0]/NET0131  & ~n1845 ;
  assign n1847 = ~n1824 & ~n1846 ;
  assign n1848 = \reg1_reg[27]/NET0131  & ~n1426 ;
  assign n1849 = \reg1_reg[27]/NET0131  & ~n1635 ;
  assign n1850 = n1635 & ~n1743 ;
  assign n1851 = ~n1849 & ~n1850 ;
  assign n1852 = n1292 & ~n1851 ;
  assign n1853 = n1635 & ~n1767 ;
  assign n1854 = ~n1849 & ~n1853 ;
  assign n1855 = n1190 & ~n1854 ;
  assign n1856 = n1635 & ~n1813 ;
  assign n1857 = \reg1_reg[27]/NET0131  & ~n1647 ;
  assign n1858 = ~n1856 & ~n1857 ;
  assign n1859 = ~n1855 & n1858 ;
  assign n1860 = ~n1852 & n1859 ;
  assign n1861 = n1386 & ~n1860 ;
  assign n1862 = \reg1_reg[27]/NET0131  & n1388 ;
  assign n1863 = ~n1861 & ~n1862 ;
  assign n1864 = \state_reg[0]/NET0131  & ~n1863 ;
  assign n1865 = ~n1848 & ~n1864 ;
  assign n1866 = \reg1_reg[29]/NET0131  & ~n1426 ;
  assign n1867 = \reg1_reg[29]/NET0131  & n1388 ;
  assign n1868 = n1635 & ~n1827 ;
  assign n1869 = \reg1_reg[29]/NET0131  & ~n1635 ;
  assign n1870 = ~n1445 & n1635 ;
  assign n1871 = ~n1869 & ~n1870 ;
  assign n1872 = n1370 & ~n1871 ;
  assign n1873 = \reg1_reg[29]/NET0131  & ~n1646 ;
  assign n1880 = ~n1872 & ~n1873 ;
  assign n1881 = ~n1868 & n1880 ;
  assign n1874 = ~n1524 & n1635 ;
  assign n1875 = ~n1869 & ~n1874 ;
  assign n1876 = n1292 & ~n1875 ;
  assign n1877 = n1592 & n1635 ;
  assign n1878 = ~n1869 & ~n1877 ;
  assign n1879 = n1190 & ~n1878 ;
  assign n1882 = ~n1876 & ~n1879 ;
  assign n1883 = n1881 & n1882 ;
  assign n1884 = n1386 & ~n1883 ;
  assign n1885 = ~n1867 & ~n1884 ;
  assign n1886 = \state_reg[0]/NET0131  & ~n1885 ;
  assign n1887 = ~n1866 & ~n1886 ;
  assign n1890 = n575 & n1388 ;
  assign n1892 = n575 & ~n1169 ;
  assign n1893 = n1036 & ~n1669 ;
  assign n1894 = ~n1036 & n1669 ;
  assign n1895 = ~n1893 & ~n1894 ;
  assign n1896 = n1169 & n1895 ;
  assign n1897 = ~n1892 & ~n1896 ;
  assign n1898 = n1190 & ~n1897 ;
  assign n1905 = ~n541 & n1345 ;
  assign n1906 = n541 & ~n1345 ;
  assign n1907 = ~n1905 & ~n1906 ;
  assign n1908 = ~n338 & ~n1907 ;
  assign n1909 = n338 & n592 ;
  assign n1910 = ~n1908 & ~n1909 ;
  assign n1911 = n1169 & n1910 ;
  assign n1912 = ~n1892 & ~n1911 ;
  assign n1913 = n1370 & ~n1912 ;
  assign n1899 = n1036 & ~n1683 ;
  assign n1900 = ~n1036 & n1683 ;
  assign n1901 = ~n1899 & ~n1900 ;
  assign n1902 = n1169 & ~n1901 ;
  assign n1903 = ~n1892 & ~n1902 ;
  assign n1904 = n1292 & ~n1903 ;
  assign n1914 = ~n601 & n1302 ;
  assign n1915 = n572 & n1914 ;
  assign n1916 = ~n572 & ~n1914 ;
  assign n1917 = ~n1915 & ~n1916 ;
  assign n1918 = n1169 & n1917 ;
  assign n1919 = ~n1892 & ~n1918 ;
  assign n1920 = n1326 & ~n1919 ;
  assign n1891 = ~n572 & ~n1332 ;
  assign n1921 = n575 & ~n1375 ;
  assign n1922 = ~n1891 & ~n1921 ;
  assign n1923 = ~n1920 & n1922 ;
  assign n1924 = ~n1904 & n1923 ;
  assign n1925 = ~n1913 & n1924 ;
  assign n1926 = ~n1898 & n1925 ;
  assign n1927 = n1386 & ~n1926 ;
  assign n1928 = ~n1890 & ~n1927 ;
  assign n1929 = \state_reg[0]/NET0131  & ~n1928 ;
  assign n1888 = \reg3_reg[11]/NET0131  & ~\state_reg[0]/NET0131  ;
  assign n1889 = n311 & n575 ;
  assign n1930 = ~n1888 & ~n1889 ;
  assign n1931 = ~n1929 & n1930 ;
  assign n1934 = n537 & n1388 ;
  assign n1936 = n537 & ~n1169 ;
  assign n1937 = n1026 & n1171 ;
  assign n1938 = ~n1026 & ~n1171 ;
  assign n1939 = ~n1937 & ~n1938 ;
  assign n1940 = n1169 & n1939 ;
  assign n1941 = ~n1936 & ~n1940 ;
  assign n1942 = n1190 & ~n1941 ;
  assign n1952 = n1026 & n1243 ;
  assign n1953 = ~n1026 & ~n1243 ;
  assign n1954 = ~n1952 & ~n1953 ;
  assign n1955 = n1169 & ~n1954 ;
  assign n1956 = ~n1936 & ~n1955 ;
  assign n1957 = n1292 & ~n1956 ;
  assign n1943 = n298 & ~n1905 ;
  assign n1944 = ~n298 & n1905 ;
  assign n1945 = ~n1943 & ~n1944 ;
  assign n1946 = ~n338 & ~n1945 ;
  assign n1947 = n338 & n581 ;
  assign n1948 = ~n1946 & ~n1947 ;
  assign n1949 = n1169 & n1948 ;
  assign n1950 = ~n1936 & ~n1949 ;
  assign n1951 = n1370 & ~n1950 ;
  assign n1958 = n551 & ~n1915 ;
  assign n1959 = ~n551 & n1915 ;
  assign n1960 = ~n1958 & ~n1959 ;
  assign n1961 = n1169 & n1960 ;
  assign n1962 = ~n1936 & ~n1961 ;
  assign n1963 = n1326 & ~n1962 ;
  assign n1935 = n551 & ~n1332 ;
  assign n1964 = n537 & ~n1375 ;
  assign n1965 = ~n1935 & ~n1964 ;
  assign n1966 = ~n1963 & n1965 ;
  assign n1967 = ~n1951 & n1966 ;
  assign n1968 = ~n1957 & n1967 ;
  assign n1969 = ~n1942 & n1968 ;
  assign n1970 = n1386 & ~n1969 ;
  assign n1971 = ~n1934 & ~n1970 ;
  assign n1972 = \state_reg[0]/NET0131  & ~n1971 ;
  assign n1932 = \reg3_reg[12]/NET0131  & ~\state_reg[0]/NET0131  ;
  assign n1933 = n311 & n537 ;
  assign n1973 = ~n1932 & ~n1933 ;
  assign n1974 = ~n1972 & n1973 ;
  assign n1977 = n437 & n1388 ;
  assign n1978 = n437 & ~n1169 ;
  assign n1982 = n955 & n982 ;
  assign n1979 = n954 & ~n964 ;
  assign n1980 = n949 & ~n1979 ;
  assign n1981 = n951 & ~n1980 ;
  assign n1983 = n901 & ~n1981 ;
  assign n1984 = ~n1982 & n1983 ;
  assign n1985 = n1050 & ~n1984 ;
  assign n1986 = ~n1050 & n1984 ;
  assign n1987 = ~n1985 & ~n1986 ;
  assign n1988 = n1169 & ~n1987 ;
  assign n1989 = ~n1978 & ~n1988 ;
  assign n1990 = n1190 & ~n1989 ;
  assign n1991 = n338 & ~n474 ;
  assign n1992 = n1353 & n1356 ;
  assign n1993 = ~n441 & n1992 ;
  assign n1994 = n426 & ~n1993 ;
  assign n1995 = ~n338 & ~n1771 ;
  assign n1996 = ~n1994 & n1995 ;
  assign n1997 = ~n1991 & ~n1996 ;
  assign n1998 = n1169 & ~n1997 ;
  assign n1999 = ~n1978 & ~n1998 ;
  assign n2000 = n1370 & ~n1999 ;
  assign n2001 = n428 & ~n1332 ;
  assign n2002 = n437 & ~n1375 ;
  assign n2025 = ~n2001 & ~n2002 ;
  assign n2026 = ~n2000 & n2025 ;
  assign n2027 = ~n1990 & n2026 ;
  assign n2003 = ~n830 & n1313 ;
  assign n2004 = ~n476 & n2003 ;
  assign n2005 = ~n465 & n2004 ;
  assign n2006 = n428 & ~n2005 ;
  assign n2007 = ~n1317 & ~n2006 ;
  assign n2008 = n1169 & n2007 ;
  assign n2009 = ~n1978 & ~n2008 ;
  assign n2010 = n1326 & ~n2009 ;
  assign n2011 = n1201 & n1242 ;
  assign n2012 = n1196 & ~n1212 ;
  assign n2013 = n1252 & ~n2012 ;
  assign n2014 = n1200 & ~n2013 ;
  assign n2015 = n1260 & ~n2014 ;
  assign n2016 = ~n2011 & n2015 ;
  assign n2017 = n1268 & ~n2016 ;
  assign n2018 = ~n1280 & ~n2017 ;
  assign n2019 = n1050 & n2018 ;
  assign n2020 = ~n1050 & ~n2018 ;
  assign n2021 = ~n2019 & ~n2020 ;
  assign n2022 = n1169 & ~n2021 ;
  assign n2023 = ~n1978 & ~n2022 ;
  assign n2024 = n1292 & ~n2023 ;
  assign n2028 = ~n2010 & ~n2024 ;
  assign n2029 = n2027 & n2028 ;
  assign n2030 = n1386 & ~n2029 ;
  assign n2031 = ~n1977 & ~n2030 ;
  assign n2032 = \state_reg[0]/NET0131  & ~n2031 ;
  assign n1975 = \reg3_reg[24]/NET0131  & ~\state_reg[0]/NET0131  ;
  assign n1976 = n311 & n437 ;
  assign n2033 = ~n1975 & ~n1976 ;
  assign n2034 = ~n2032 & n2033 ;
  assign n2035 = n470 & n1388 ;
  assign n2036 = n470 & ~n1169 ;
  assign n2037 = ~n1734 & n1735 ;
  assign n2038 = n1724 & ~n2037 ;
  assign n2039 = n1063 & n2038 ;
  assign n2040 = ~n1063 & ~n2038 ;
  assign n2041 = ~n2039 & ~n2040 ;
  assign n2042 = n1169 & ~n2041 ;
  assign n2043 = ~n2036 & ~n2042 ;
  assign n2044 = n1292 & ~n2043 ;
  assign n2045 = n913 & n1552 ;
  assign n2046 = n1752 & n2045 ;
  assign n2047 = ~n1671 & n2046 ;
  assign n2048 = ~n1757 & n2045 ;
  assign n2049 = n1748 & ~n2048 ;
  assign n2050 = ~n2047 & n2049 ;
  assign n2051 = n1063 & ~n2050 ;
  assign n2052 = ~n1063 & n2050 ;
  assign n2053 = ~n2051 & ~n2052 ;
  assign n2054 = n1169 & ~n2053 ;
  assign n2055 = ~n2036 & ~n2054 ;
  assign n2056 = n1190 & ~n2055 ;
  assign n2065 = n465 & ~n2004 ;
  assign n2066 = ~n2005 & ~n2065 ;
  assign n2067 = n1169 & n2066 ;
  assign n2068 = ~n2036 & ~n2067 ;
  assign n2069 = n1326 & ~n2068 ;
  assign n2057 = n441 & ~n1992 ;
  assign n2058 = ~n1993 & ~n2057 ;
  assign n2059 = ~n338 & ~n2058 ;
  assign n2060 = n338 & n486 ;
  assign n2061 = ~n2059 & ~n2060 ;
  assign n2062 = n1169 & n2061 ;
  assign n2063 = ~n2036 & ~n2062 ;
  assign n2064 = n1370 & ~n2063 ;
  assign n2070 = n470 & ~n1375 ;
  assign n2071 = n465 & ~n1332 ;
  assign n2072 = ~n2070 & ~n2071 ;
  assign n2073 = ~n2064 & n2072 ;
  assign n2074 = ~n2069 & n2073 ;
  assign n2075 = ~n2056 & n2074 ;
  assign n2076 = ~n2044 & n2075 ;
  assign n2077 = n1386 & ~n2076 ;
  assign n2078 = ~n2035 & ~n2077 ;
  assign n2079 = \state_reg[0]/NET0131  & ~n2078 ;
  assign n2080 = \reg3_reg[23]/NET0131  & ~\state_reg[0]/NET0131  ;
  assign n2081 = n311 & n470 ;
  assign n2082 = ~n2080 & ~n2081 ;
  assign n2083 = ~n2079 & n2082 ;
  assign n2084 = \reg0_reg[15]/NET0131  & ~n1426 ;
  assign n2085 = \reg0_reg[15]/NET0131  & n1388 ;
  assign n2092 = \reg0_reg[15]/NET0131  & ~n1607 ;
  assign n2093 = n1607 & n1674 ;
  assign n2094 = ~n2092 & ~n2093 ;
  assign n2095 = n1190 & ~n2094 ;
  assign n2096 = n1607 & ~n1691 ;
  assign n2097 = ~n2092 & ~n2096 ;
  assign n2098 = n1292 & ~n2097 ;
  assign n2087 = n1370 & n1700 ;
  assign n2086 = n1326 & n1707 ;
  assign n2088 = n522 & n1328 ;
  assign n2089 = ~n2086 & ~n2088 ;
  assign n2090 = ~n2087 & n2089 ;
  assign n2091 = n1607 & ~n2090 ;
  assign n2099 = \reg0_reg[15]/NET0131  & ~n1624 ;
  assign n2100 = ~n2091 & ~n2099 ;
  assign n2101 = ~n2098 & n2100 ;
  assign n2102 = ~n2095 & n2101 ;
  assign n2103 = n1386 & ~n2102 ;
  assign n2104 = ~n2085 & ~n2103 ;
  assign n2105 = \state_reg[0]/NET0131  & ~n2104 ;
  assign n2106 = ~n2084 & ~n2105 ;
  assign n2107 = \reg0_reg[23]/NET0131  & ~n1426 ;
  assign n2108 = \reg0_reg[23]/NET0131  & n1388 ;
  assign n2109 = \reg0_reg[23]/NET0131  & ~n1607 ;
  assign n2110 = n1607 & ~n2041 ;
  assign n2111 = ~n2109 & ~n2110 ;
  assign n2112 = n1292 & ~n2111 ;
  assign n2113 = n1607 & ~n2053 ;
  assign n2114 = ~n2109 & ~n2113 ;
  assign n2115 = n1190 & ~n2114 ;
  assign n2118 = n1326 & n2066 ;
  assign n2116 = n465 & n1328 ;
  assign n2117 = n1370 & n2061 ;
  assign n2119 = ~n2116 & ~n2117 ;
  assign n2120 = ~n2118 & n2119 ;
  assign n2121 = n1607 & ~n2120 ;
  assign n2122 = \reg0_reg[23]/NET0131  & ~n1624 ;
  assign n2123 = ~n2121 & ~n2122 ;
  assign n2124 = ~n2115 & n2123 ;
  assign n2125 = ~n2112 & n2124 ;
  assign n2126 = n1386 & ~n2125 ;
  assign n2127 = ~n2108 & ~n2126 ;
  assign n2128 = \state_reg[0]/NET0131  & ~n2127 ;
  assign n2129 = ~n2107 & ~n2128 ;
  assign n2130 = \reg0_reg[24]/NET0131  & ~n1426 ;
  assign n2131 = \reg0_reg[24]/NET0131  & n1388 ;
  assign n2132 = \reg0_reg[24]/NET0131  & ~n1607 ;
  assign n2133 = n1607 & ~n1987 ;
  assign n2134 = ~n2132 & ~n2133 ;
  assign n2135 = n1190 & ~n2134 ;
  assign n2136 = n1607 & ~n1997 ;
  assign n2137 = ~n2132 & ~n2136 ;
  assign n2138 = n1370 & ~n2137 ;
  assign n2139 = n428 & n1328 ;
  assign n2140 = n1607 & n2139 ;
  assign n2141 = n1328 & ~n1607 ;
  assign n2142 = n1620 & ~n2141 ;
  assign n2143 = \reg0_reg[24]/NET0131  & ~n2142 ;
  assign n2150 = ~n2140 & ~n2143 ;
  assign n2151 = ~n2138 & n2150 ;
  assign n2152 = ~n2135 & n2151 ;
  assign n2144 = n1607 & n2007 ;
  assign n2145 = ~n2132 & ~n2144 ;
  assign n2146 = n1326 & ~n2145 ;
  assign n2147 = n1607 & ~n2021 ;
  assign n2148 = ~n2132 & ~n2147 ;
  assign n2149 = n1292 & ~n2148 ;
  assign n2153 = ~n2146 & ~n2149 ;
  assign n2154 = n2152 & n2153 ;
  assign n2155 = n1386 & ~n2154 ;
  assign n2156 = ~n2131 & ~n2155 ;
  assign n2157 = \state_reg[0]/NET0131  & ~n2156 ;
  assign n2158 = ~n2130 & ~n2157 ;
  assign n2159 = \reg1_reg[15]/NET0131  & ~n1426 ;
  assign n2160 = \reg1_reg[15]/NET0131  & n1388 ;
  assign n2162 = \reg1_reg[15]/NET0131  & ~n1635 ;
  assign n2163 = n1635 & n1674 ;
  assign n2164 = ~n2162 & ~n2163 ;
  assign n2165 = n1190 & ~n2164 ;
  assign n2166 = n1635 & ~n1691 ;
  assign n2167 = ~n2162 & ~n2166 ;
  assign n2168 = n1292 & ~n2167 ;
  assign n2161 = n1635 & ~n2090 ;
  assign n2169 = \reg1_reg[15]/NET0131  & ~n1647 ;
  assign n2170 = ~n2161 & ~n2169 ;
  assign n2171 = ~n2168 & n2170 ;
  assign n2172 = ~n2165 & n2171 ;
  assign n2173 = n1386 & ~n2172 ;
  assign n2174 = ~n2160 & ~n2173 ;
  assign n2175 = \state_reg[0]/NET0131  & ~n2174 ;
  assign n2176 = ~n2159 & ~n2175 ;
  assign n2177 = \reg1_reg[23]/NET0131  & ~n1426 ;
  assign n2178 = \reg1_reg[23]/NET0131  & n1388 ;
  assign n2179 = \reg1_reg[23]/NET0131  & ~n1635 ;
  assign n2180 = n1635 & ~n2041 ;
  assign n2181 = ~n2179 & ~n2180 ;
  assign n2182 = n1292 & ~n2181 ;
  assign n2183 = n1635 & ~n2053 ;
  assign n2184 = ~n2179 & ~n2183 ;
  assign n2185 = n1190 & ~n2184 ;
  assign n2186 = n1635 & ~n2120 ;
  assign n2187 = \reg1_reg[23]/NET0131  & ~n1647 ;
  assign n2188 = ~n2186 & ~n2187 ;
  assign n2189 = ~n2185 & n2188 ;
  assign n2190 = ~n2182 & n2189 ;
  assign n2191 = n1386 & ~n2190 ;
  assign n2192 = ~n2178 & ~n2191 ;
  assign n2193 = \state_reg[0]/NET0131  & ~n2192 ;
  assign n2194 = ~n2177 & ~n2193 ;
  assign n2195 = \reg2_reg[15]/NET0131  & ~n1426 ;
  assign n2196 = \reg2_reg[15]/NET0131  & n1388 ;
  assign n2198 = \reg2_reg[15]/NET0131  & ~n1396 ;
  assign n2199 = n1396 & n1674 ;
  assign n2200 = ~n2198 & ~n2199 ;
  assign n2201 = n1190 & ~n2200 ;
  assign n2203 = n1396 & ~n1691 ;
  assign n2204 = ~n2198 & ~n2203 ;
  assign n2205 = n1292 & ~n2204 ;
  assign n2197 = n1396 & ~n2090 ;
  assign n2202 = n508 & n1331 ;
  assign n2206 = n1370 & ~n1396 ;
  assign n2207 = ~n1396 & ~n1621 ;
  assign n2208 = ~n1373 & ~n2207 ;
  assign n2209 = ~n2206 & n2208 ;
  assign n2210 = \reg2_reg[15]/NET0131  & ~n2209 ;
  assign n2211 = ~n2202 & ~n2210 ;
  assign n2212 = ~n2197 & n2211 ;
  assign n2213 = ~n2205 & n2212 ;
  assign n2214 = ~n2201 & n2213 ;
  assign n2215 = n1386 & ~n2214 ;
  assign n2216 = ~n2196 & ~n2215 ;
  assign n2217 = \state_reg[0]/NET0131  & ~n2216 ;
  assign n2218 = ~n2195 & ~n2217 ;
  assign n2219 = \reg2_reg[23]/NET0131  & ~n1426 ;
  assign n2220 = \reg2_reg[23]/NET0131  & n1388 ;
  assign n2221 = \reg2_reg[23]/NET0131  & ~n1396 ;
  assign n2222 = n1396 & ~n2041 ;
  assign n2223 = ~n2221 & ~n2222 ;
  assign n2224 = n1292 & ~n2223 ;
  assign n2225 = n1396 & ~n2053 ;
  assign n2226 = ~n2221 & ~n2225 ;
  assign n2227 = n1190 & ~n2226 ;
  assign n2228 = n1396 & ~n2120 ;
  assign n2229 = n470 & n1331 ;
  assign n2230 = \reg2_reg[23]/NET0131  & ~n2209 ;
  assign n2231 = ~n2229 & ~n2230 ;
  assign n2232 = ~n2228 & n2231 ;
  assign n2233 = ~n2227 & n2232 ;
  assign n2234 = ~n2224 & n2233 ;
  assign n2235 = n1386 & ~n2234 ;
  assign n2236 = ~n2220 & ~n2235 ;
  assign n2237 = \state_reg[0]/NET0131  & ~n2236 ;
  assign n2238 = ~n2219 & ~n2237 ;
  assign n2240 = n493 & n1388 ;
  assign n2267 = n637 & n976 ;
  assign n2268 = n637 & n978 ;
  assign n2269 = n957 & ~n2268 ;
  assign n2270 = ~n2267 & n2269 ;
  assign n2271 = n562 & n603 ;
  assign n2272 = ~n2270 & n2271 ;
  assign n2273 = n562 & n960 ;
  assign n2274 = ~n554 & ~n2273 ;
  assign n2275 = ~n2272 & n2274 ;
  assign n2277 = ~n1040 & n2275 ;
  assign n2276 = n1040 & ~n2275 ;
  assign n2278 = n1190 & ~n2276 ;
  assign n2279 = ~n2277 & n2278 ;
  assign n2252 = n1193 & n1211 ;
  assign n2253 = n1247 & ~n2252 ;
  assign n2254 = ~n1229 & n1233 ;
  assign n2255 = n1214 & n1240 ;
  assign n2256 = ~n2254 & n2255 ;
  assign n2257 = ~n1237 & n1240 ;
  assign n2258 = n1207 & ~n2257 ;
  assign n2259 = ~n2256 & n2258 ;
  assign n2260 = n1193 & n1203 ;
  assign n2261 = ~n2259 & n2260 ;
  assign n2262 = n2253 & ~n2261 ;
  assign n2264 = ~n1040 & ~n2262 ;
  assign n2263 = n1040 & n2262 ;
  assign n2265 = n1292 & ~n2263 ;
  assign n2266 = ~n2264 & n2265 ;
  assign n2242 = ~n338 & ~n515 ;
  assign n2243 = ~n498 & n1944 ;
  assign n2244 = ~n2242 & ~n2243 ;
  assign n2245 = ~n1349 & ~n2244 ;
  assign n2246 = ~n298 & n338 ;
  assign n2247 = ~n2245 & ~n2246 ;
  assign n2248 = n1370 & ~n2247 ;
  assign n2249 = ~n504 & ~n1306 ;
  assign n2250 = n1326 & ~n1704 ;
  assign n2251 = ~n2249 & n2250 ;
  assign n2280 = ~n2248 & ~n2251 ;
  assign n2281 = ~n2266 & n2280 ;
  assign n2282 = ~n2279 & n2281 ;
  assign n2283 = n1169 & ~n2282 ;
  assign n2241 = ~n504 & ~n1332 ;
  assign n2284 = ~n1131 & ~n1291 ;
  assign n2285 = ~n1169 & ~n2284 ;
  assign n2286 = n1375 & ~n2285 ;
  assign n2287 = n493 & ~n2286 ;
  assign n2288 = ~n2241 & ~n2287 ;
  assign n2289 = ~n2283 & n2288 ;
  assign n2290 = n1386 & ~n2289 ;
  assign n2291 = ~n2240 & ~n2290 ;
  assign n2292 = \state_reg[0]/NET0131  & ~n2291 ;
  assign n2239 = n311 & n493 ;
  assign n2293 = \reg3_reg[14]/NET0131  & ~\state_reg[0]/NET0131  ;
  assign n2294 = ~n2239 & ~n2293 ;
  assign n2295 = ~n2292 & n2294 ;
  assign n2298 = n880 & n1388 ;
  assign n2300 = n880 & ~n1169 ;
  assign n2309 = n983 & n1053 ;
  assign n2310 = ~n983 & ~n1053 ;
  assign n2311 = ~n2309 & ~n2310 ;
  assign n2312 = n1169 & n2311 ;
  assign n2313 = ~n2300 & ~n2312 ;
  assign n2314 = n1190 & ~n2313 ;
  assign n2301 = n1196 & ~n1243 ;
  assign n2302 = n1252 & ~n2301 ;
  assign n2303 = n1053 & ~n2302 ;
  assign n2304 = ~n1053 & n2302 ;
  assign n2305 = ~n2303 & ~n2304 ;
  assign n2306 = n1169 & n2305 ;
  assign n2307 = ~n2300 & ~n2306 ;
  assign n2308 = n1292 & ~n2307 ;
  assign n2315 = n862 & ~n1695 ;
  assign n2316 = ~n862 & n1695 ;
  assign n2317 = ~n2315 & ~n2316 ;
  assign n2318 = ~n338 & ~n2317 ;
  assign n2319 = n338 & n515 ;
  assign n2320 = ~n2318 & ~n2319 ;
  assign n2321 = n1169 & n2320 ;
  assign n2322 = ~n2300 & ~n2321 ;
  assign n2323 = n1370 & ~n2322 ;
  assign n2324 = n878 & ~n1706 ;
  assign n2325 = n1306 & n1308 ;
  assign n2326 = ~n2324 & ~n2325 ;
  assign n2327 = n1169 & n2326 ;
  assign n2328 = ~n2300 & ~n2327 ;
  assign n2329 = n1326 & ~n2328 ;
  assign n2299 = n878 & ~n1332 ;
  assign n2330 = n880 & ~n1375 ;
  assign n2331 = ~n2299 & ~n2330 ;
  assign n2332 = ~n2329 & n2331 ;
  assign n2333 = ~n2323 & n2332 ;
  assign n2334 = ~n2308 & n2333 ;
  assign n2335 = ~n2314 & n2334 ;
  assign n2336 = n1386 & ~n2335 ;
  assign n2337 = ~n2298 & ~n2336 ;
  assign n2338 = \state_reg[0]/NET0131  & ~n2337 ;
  assign n2296 = n311 & n880 ;
  assign n2297 = \reg3_reg[16]/NET0131  & ~\state_reg[0]/NET0131  ;
  assign n2339 = ~n2296 & ~n2297 ;
  assign n2340 = ~n2338 & n2339 ;
  assign n2343 = n666 & n1388 ;
  assign n2347 = n666 & ~n1169 ;
  assign n2354 = n628 & ~n1341 ;
  assign n2355 = ~n628 & n1341 ;
  assign n2356 = ~n2354 & ~n2355 ;
  assign n2357 = ~n338 & ~n2356 ;
  assign n2358 = n338 & n661 ;
  assign n2359 = ~n2357 & ~n2358 ;
  assign n2360 = n1169 & n2359 ;
  assign n2361 = ~n2347 & ~n2360 ;
  assign n2362 = n1370 & ~n2361 ;
  assign n2348 = n1030 & n1664 ;
  assign n2349 = ~n1030 & ~n1664 ;
  assign n2350 = ~n2348 & ~n2349 ;
  assign n2351 = n1169 & n2350 ;
  assign n2352 = ~n2347 & ~n2351 ;
  assign n2353 = n1190 & ~n2352 ;
  assign n2363 = n1030 & n1678 ;
  assign n2364 = ~n1030 & ~n1678 ;
  assign n2365 = ~n2363 & ~n2364 ;
  assign n2366 = n1169 & ~n2365 ;
  assign n2367 = ~n2347 & ~n2366 ;
  assign n2368 = n1292 & ~n2367 ;
  assign n2369 = n652 & n1298 ;
  assign n2370 = n679 & ~n2369 ;
  assign n2371 = ~n1300 & n1326 ;
  assign n2372 = ~n2370 & n2371 ;
  assign n2373 = n1169 & n2372 ;
  assign n2344 = ~n1169 & ~n1621 ;
  assign n2345 = ~n1373 & ~n2344 ;
  assign n2346 = n666 & ~n2345 ;
  assign n2374 = n679 & ~n1332 ;
  assign n2375 = ~n2346 & ~n2374 ;
  assign n2376 = ~n2373 & n2375 ;
  assign n2377 = ~n2368 & n2376 ;
  assign n2378 = ~n2353 & n2377 ;
  assign n2379 = ~n2362 & n2378 ;
  assign n2380 = n1386 & ~n2379 ;
  assign n2381 = ~n2343 & ~n2380 ;
  assign n2382 = \state_reg[0]/NET0131  & ~n2381 ;
  assign n2341 = \reg3_reg[7]/NET0131  & ~\state_reg[0]/NET0131  ;
  assign n2342 = n311 & n666 ;
  assign n2383 = ~n2341 & ~n2342 ;
  assign n2384 = ~n2382 & n2383 ;
  assign n2385 = \reg3_reg[19]/NET0131  & ~\state_reg[0]/NET0131  ;
  assign n2388 = n802 & ~n1169 ;
  assign n2389 = n1081 & n1734 ;
  assign n2390 = ~n1081 & ~n1734 ;
  assign n2391 = ~n2389 & ~n2390 ;
  assign n2392 = n1169 & n2391 ;
  assign n2393 = ~n2388 & ~n2392 ;
  assign n2394 = n1292 & ~n2393 ;
  assign n2395 = n1081 & n1759 ;
  assign n2396 = ~n1081 & ~n1759 ;
  assign n2397 = ~n2395 & ~n2396 ;
  assign n2398 = n1169 & ~n2397 ;
  assign n2399 = ~n2388 & ~n2398 ;
  assign n2400 = n1190 & ~n2399 ;
  assign n2401 = ~n851 & n1353 ;
  assign n2402 = n851 & ~n1353 ;
  assign n2403 = ~n2401 & ~n2402 ;
  assign n2404 = ~n338 & ~n2403 ;
  assign n2405 = n338 & n827 ;
  assign n2406 = ~n2404 & ~n2405 ;
  assign n2407 = n1169 & n2406 ;
  assign n2408 = ~n2388 & ~n2407 ;
  assign n2409 = n1370 & ~n2408 ;
  assign n2410 = ~n817 & n1310 ;
  assign n2411 = ~n797 & ~n2410 ;
  assign n2412 = n797 & n2410 ;
  assign n2413 = ~n2411 & ~n2412 ;
  assign n2414 = n1169 & n2413 ;
  assign n2415 = ~n2388 & ~n2414 ;
  assign n2416 = n1326 & ~n2415 ;
  assign n2417 = ~n797 & ~n1332 ;
  assign n2387 = n802 & ~n1375 ;
  assign n2418 = n1386 & ~n2387 ;
  assign n2419 = ~n2417 & n2418 ;
  assign n2420 = ~n2416 & n2419 ;
  assign n2421 = ~n2409 & n2420 ;
  assign n2422 = ~n2400 & n2421 ;
  assign n2423 = ~n2394 & n2422 ;
  assign n2386 = ~n802 & ~n1386 ;
  assign n2424 = \state_reg[0]/NET0131  & ~n2386 ;
  assign n2425 = ~n2423 & n2424 ;
  assign n2426 = ~n2385 & ~n2425 ;
  assign n2429 = n847 & n1388 ;
  assign n2431 = n847 & ~n1169 ;
  assign n2432 = n1084 & ~n1176 ;
  assign n2433 = ~n1084 & n1176 ;
  assign n2434 = ~n2432 & ~n2433 ;
  assign n2435 = n1169 & ~n2434 ;
  assign n2436 = ~n2431 & ~n2435 ;
  assign n2437 = n1190 & ~n2436 ;
  assign n2447 = n1084 & n1262 ;
  assign n2448 = ~n1084 & ~n1262 ;
  assign n2449 = ~n2447 & ~n2448 ;
  assign n2450 = n1169 & ~n2449 ;
  assign n2451 = ~n2431 & ~n2450 ;
  assign n2452 = n1292 & ~n2451 ;
  assign n2438 = n840 & ~n2401 ;
  assign n2439 = ~n840 & n2401 ;
  assign n2440 = ~n2438 & ~n2439 ;
  assign n2441 = ~n338 & ~n2440 ;
  assign n2442 = n338 & n806 ;
  assign n2443 = ~n2441 & ~n2442 ;
  assign n2444 = n1169 & n2443 ;
  assign n2445 = ~n2431 & ~n2444 ;
  assign n2446 = n1370 & ~n2445 ;
  assign n2453 = n842 & ~n2412 ;
  assign n2454 = ~n1313 & ~n2453 ;
  assign n2455 = n1169 & n2454 ;
  assign n2456 = ~n2431 & ~n2455 ;
  assign n2457 = n1326 & ~n2456 ;
  assign n2430 = n842 & ~n1332 ;
  assign n2458 = n847 & ~n1375 ;
  assign n2459 = ~n2430 & ~n2458 ;
  assign n2460 = ~n2457 & n2459 ;
  assign n2461 = ~n2446 & n2460 ;
  assign n2462 = ~n2452 & n2461 ;
  assign n2463 = ~n2437 & n2462 ;
  assign n2464 = n1386 & ~n2463 ;
  assign n2465 = ~n2429 & ~n2464 ;
  assign n2466 = \state_reg[0]/NET0131  & ~n2465 ;
  assign n2427 = n311 & n847 ;
  assign n2428 = \reg3_reg[20]/NET0131  & ~\state_reg[0]/NET0131  ;
  assign n2467 = ~n2427 & ~n2428 ;
  assign n2468 = ~n2466 & n2467 ;
  assign n2469 = n559 & n907 ;
  assign n2470 = ~n946 & ~n2469 ;
  assign n2471 = n524 & n907 ;
  assign n2472 = ~n2275 & n2471 ;
  assign n2473 = n2470 & ~n2472 ;
  assign n2474 = n904 & n950 ;
  assign n2475 = n443 & n896 ;
  assign n2476 = n2474 & n2475 ;
  assign n2477 = ~n2473 & n2476 ;
  assign n2479 = n948 & n950 ;
  assign n2480 = ~n898 & ~n2479 ;
  assign n2481 = n2475 & ~n2480 ;
  assign n2478 = n443 & n900 ;
  assign n2482 = ~n990 & ~n2478 ;
  assign n2483 = ~n2481 & n2482 ;
  assign n2484 = ~n2477 & n2483 ;
  assign n2485 = n1060 & ~n2484 ;
  assign n2486 = ~n1060 & n2484 ;
  assign n2487 = ~n2485 & ~n2486 ;
  assign n2488 = n1169 & n2487 ;
  assign n2489 = ~n450 & ~n1169 ;
  assign n2490 = n1190 & ~n2489 ;
  assign n2491 = ~n2488 & n2490 ;
  assign n2500 = ~n1046 & ~n1083 ;
  assign n2501 = n1199 & n2500 ;
  assign n2502 = ~n1069 & n1736 ;
  assign n2503 = n2501 & n2502 ;
  assign n2504 = n1195 & n1197 ;
  assign n2505 = n2503 & n2504 ;
  assign n2506 = n2261 & n2505 ;
  assign n2507 = ~n2253 & n2504 ;
  assign n2508 = n1197 & ~n1251 ;
  assign n2509 = ~n1255 & ~n2508 ;
  assign n2510 = ~n2507 & n2509 ;
  assign n2511 = n2503 & ~n2510 ;
  assign n2512 = ~n1259 & n2500 ;
  assign n2513 = n1277 & ~n2512 ;
  assign n2514 = n2502 & ~n2513 ;
  assign n2515 = ~n1275 & n1736 ;
  assign n2516 = n1272 & ~n2515 ;
  assign n2517 = ~n2514 & n2516 ;
  assign n2518 = ~n2511 & n2517 ;
  assign n2519 = ~n2506 & n2518 ;
  assign n2521 = n1060 & ~n2519 ;
  assign n2520 = ~n1060 & n2519 ;
  assign n2522 = n1292 & ~n2520 ;
  assign n2523 = ~n2521 & n2522 ;
  assign n2493 = n338 & ~n426 ;
  assign n2494 = ~n338 & ~n414 ;
  assign n2495 = ~n454 & n1771 ;
  assign n2496 = ~n2494 & ~n2495 ;
  assign n2497 = ~n1772 & ~n2496 ;
  assign n2498 = ~n2493 & ~n2497 ;
  assign n2499 = n1370 & ~n2498 ;
  assign n2524 = ~n417 & n1317 ;
  assign n2525 = n445 & ~n2524 ;
  assign n2526 = ~n1319 & n1326 ;
  assign n2527 = ~n2525 & n2526 ;
  assign n2528 = ~n2499 & ~n2527 ;
  assign n2529 = ~n2523 & n2528 ;
  assign n2530 = n1169 & ~n2529 ;
  assign n2492 = n445 & ~n1332 ;
  assign n2531 = ~n1292 & ~n1326 ;
  assign n2532 = ~n1169 & ~n2531 ;
  assign n2533 = n1377 & ~n2532 ;
  assign n2534 = n450 & ~n2533 ;
  assign n2535 = ~n2492 & ~n2534 ;
  assign n2536 = ~n2530 & n2535 ;
  assign n2537 = ~n2491 & n2536 ;
  assign n2538 = n1386 & ~n2537 ;
  assign n2539 = n450 & n1388 ;
  assign n2540 = ~n2538 & ~n2539 ;
  assign n2541 = \state_reg[0]/NET0131  & ~n2540 ;
  assign n2542 = \reg3_reg[26]/NET0131  & ~\state_reg[0]/NET0131  ;
  assign n2543 = n311 & n450 ;
  assign n2544 = ~n2542 & ~n2543 ;
  assign n2545 = ~n2541 & n2544 ;
  assign n2549 = ~n367 & n1433 ;
  assign n2551 = ~n340 & n2549 ;
  assign n2550 = n340 & ~n2549 ;
  assign n2552 = n1326 & ~n2550 ;
  assign n2553 = ~n2551 & n2552 ;
  assign n2546 = n340 & n1328 ;
  assign n2547 = ~n364 & n1370 ;
  assign n2548 = n1443 & n2547 ;
  assign n2554 = ~n2546 & ~n2548 ;
  assign n2555 = ~n2553 & n2554 ;
  assign n2556 = n1396 & ~n2555 ;
  assign n2557 = ~n1449 & ~n2556 ;
  assign n2558 = n1717 & ~n2557 ;
  assign n2559 = ~n1331 & ~n1396 ;
  assign n2560 = ~n1373 & n1717 ;
  assign n2561 = ~n2559 & n2560 ;
  assign n2562 = \reg2_reg[31]/NET0131  & ~n2561 ;
  assign n2563 = ~n2558 & ~n2562 ;
  assign n2564 = \reg2_reg[26]/NET0131  & ~n1426 ;
  assign n2565 = n1396 & n2487 ;
  assign n2566 = ~\reg2_reg[26]/NET0131  & ~n1396 ;
  assign n2567 = n1190 & ~n2566 ;
  assign n2568 = ~n2565 & n2567 ;
  assign n2569 = n445 & n1328 ;
  assign n2570 = n2529 & ~n2569 ;
  assign n2571 = n1396 & ~n2570 ;
  assign n2572 = n450 & n1331 ;
  assign n2573 = n1292 & ~n1396 ;
  assign n2574 = n2208 & ~n2573 ;
  assign n2575 = ~n2206 & n2574 ;
  assign n2576 = \reg2_reg[26]/NET0131  & ~n2575 ;
  assign n2577 = ~n2572 & ~n2576 ;
  assign n2578 = ~n2571 & n2577 ;
  assign n2579 = ~n2568 & n2578 ;
  assign n2580 = n1386 & ~n2579 ;
  assign n2581 = \reg2_reg[26]/NET0131  & n1388 ;
  assign n2582 = ~n2580 & ~n2581 ;
  assign n2583 = \state_reg[0]/NET0131  & ~n2582 ;
  assign n2584 = ~n2564 & ~n2583 ;
  assign n2585 = \reg0_reg[20]/NET0131  & ~n1426 ;
  assign n2586 = \reg0_reg[20]/NET0131  & n1388 ;
  assign n2589 = \reg0_reg[20]/NET0131  & ~n1607 ;
  assign n2590 = n1607 & ~n2434 ;
  assign n2591 = ~n2589 & ~n2590 ;
  assign n2592 = n1190 & ~n2591 ;
  assign n2596 = n1607 & ~n2449 ;
  assign n2597 = ~n2589 & ~n2596 ;
  assign n2598 = n1292 & ~n2597 ;
  assign n2593 = n1607 & n2443 ;
  assign n2594 = ~n2589 & ~n2593 ;
  assign n2595 = n1370 & ~n2594 ;
  assign n2599 = n1607 & n2454 ;
  assign n2600 = ~n2589 & ~n2599 ;
  assign n2601 = n1326 & ~n2600 ;
  assign n2587 = n842 & n1328 ;
  assign n2588 = n1607 & n2587 ;
  assign n2602 = \reg0_reg[20]/NET0131  & ~n2142 ;
  assign n2603 = ~n2588 & ~n2602 ;
  assign n2604 = ~n2601 & n2603 ;
  assign n2605 = ~n2595 & n2604 ;
  assign n2606 = ~n2598 & n2605 ;
  assign n2607 = ~n2592 & n2606 ;
  assign n2608 = n1386 & ~n2607 ;
  assign n2609 = ~n2586 & ~n2608 ;
  assign n2610 = \state_reg[0]/NET0131  & ~n2609 ;
  assign n2611 = ~n2585 & ~n2610 ;
  assign n2612 = ~n1607 & ~n2531 ;
  assign n2613 = n2142 & ~n2612 ;
  assign n2614 = n1190 & ~n1607 ;
  assign n2615 = n1717 & ~n2614 ;
  assign n2616 = n2613 & n2615 ;
  assign n2617 = ~n1619 & n2616 ;
  assign n2618 = \reg0_reg[26]/NET0131  & ~n2617 ;
  assign n2619 = n1190 & ~n2487 ;
  assign n2620 = n2570 & ~n2619 ;
  assign n2621 = n1607 & n1717 ;
  assign n2622 = ~n2620 & n2621 ;
  assign n2623 = ~n2618 & ~n2622 ;
  assign n2624 = \reg1_reg[11]/NET0131  & ~n1426 ;
  assign n2625 = \reg1_reg[11]/NET0131  & n1388 ;
  assign n2627 = \reg1_reg[11]/NET0131  & ~n1635 ;
  assign n2628 = n1635 & n1895 ;
  assign n2629 = ~n2627 & ~n2628 ;
  assign n2630 = n1190 & ~n2629 ;
  assign n2634 = n1635 & n1910 ;
  assign n2635 = ~n2627 & ~n2634 ;
  assign n2636 = n1370 & ~n2635 ;
  assign n2631 = n1635 & ~n1901 ;
  assign n2632 = ~n2627 & ~n2631 ;
  assign n2633 = n1292 & ~n2632 ;
  assign n2626 = \reg1_reg[11]/NET0131  & ~n1646 ;
  assign n2637 = ~n572 & n1328 ;
  assign n2638 = n1326 & n1917 ;
  assign n2639 = ~n2637 & ~n2638 ;
  assign n2640 = n1635 & ~n2639 ;
  assign n2641 = ~n2626 & ~n2640 ;
  assign n2642 = ~n2633 & n2641 ;
  assign n2643 = ~n2636 & n2642 ;
  assign n2644 = ~n2630 & n2643 ;
  assign n2645 = n1386 & ~n2644 ;
  assign n2646 = ~n2625 & ~n2645 ;
  assign n2647 = \state_reg[0]/NET0131  & ~n2646 ;
  assign n2648 = ~n2624 & ~n2647 ;
  assign n2649 = \reg1_reg[12]/NET0131  & ~n1426 ;
  assign n2650 = \reg1_reg[12]/NET0131  & n1388 ;
  assign n2653 = \reg1_reg[12]/NET0131  & ~n1635 ;
  assign n2654 = n1635 & n1939 ;
  assign n2655 = ~n2653 & ~n2654 ;
  assign n2656 = n1190 & ~n2655 ;
  assign n2660 = n1635 & ~n1954 ;
  assign n2661 = ~n2653 & ~n2660 ;
  assign n2662 = n1292 & ~n2661 ;
  assign n2657 = n1635 & n1948 ;
  assign n2658 = ~n2653 & ~n2657 ;
  assign n2659 = n1370 & ~n2658 ;
  assign n2663 = n1635 & n1960 ;
  assign n2664 = ~n2653 & ~n2663 ;
  assign n2665 = n1326 & ~n2664 ;
  assign n2651 = n551 & n1328 ;
  assign n2652 = n1635 & n2651 ;
  assign n2666 = n1328 & ~n1635 ;
  assign n2667 = n1620 & ~n2666 ;
  assign n2668 = \reg1_reg[12]/NET0131  & ~n2667 ;
  assign n2669 = ~n2652 & ~n2668 ;
  assign n2670 = ~n2665 & n2669 ;
  assign n2671 = ~n2659 & n2670 ;
  assign n2672 = ~n2662 & n2671 ;
  assign n2673 = ~n2656 & n2672 ;
  assign n2674 = n1386 & ~n2673 ;
  assign n2675 = ~n2650 & ~n2674 ;
  assign n2676 = \state_reg[0]/NET0131  & ~n2675 ;
  assign n2677 = ~n2649 & ~n2676 ;
  assign n2678 = \reg1_reg[20]/NET0131  & ~n1426 ;
  assign n2679 = \reg1_reg[20]/NET0131  & n1388 ;
  assign n2681 = \reg1_reg[20]/NET0131  & ~n1635 ;
  assign n2682 = n1635 & ~n2434 ;
  assign n2683 = ~n2681 & ~n2682 ;
  assign n2684 = n1190 & ~n2683 ;
  assign n2688 = n1635 & ~n2449 ;
  assign n2689 = ~n2681 & ~n2688 ;
  assign n2690 = n1292 & ~n2689 ;
  assign n2685 = n1635 & n2443 ;
  assign n2686 = ~n2681 & ~n2685 ;
  assign n2687 = n1370 & ~n2686 ;
  assign n2691 = n1635 & n2454 ;
  assign n2692 = ~n2681 & ~n2691 ;
  assign n2693 = n1326 & ~n2692 ;
  assign n2680 = n1635 & n2587 ;
  assign n2694 = \reg1_reg[20]/NET0131  & ~n2667 ;
  assign n2695 = ~n2680 & ~n2694 ;
  assign n2696 = ~n2693 & n2695 ;
  assign n2697 = ~n2687 & n2696 ;
  assign n2698 = ~n2690 & n2697 ;
  assign n2699 = ~n2684 & n2698 ;
  assign n2700 = n1386 & ~n2699 ;
  assign n2701 = ~n2679 & ~n2700 ;
  assign n2702 = \state_reg[0]/NET0131  & ~n2701 ;
  assign n2703 = ~n2678 & ~n2702 ;
  assign n2704 = \reg1_reg[24]/NET0131  & ~n1426 ;
  assign n2705 = \reg1_reg[24]/NET0131  & n1388 ;
  assign n2706 = \reg1_reg[24]/NET0131  & ~n1635 ;
  assign n2707 = n1635 & ~n1987 ;
  assign n2708 = ~n2706 & ~n2707 ;
  assign n2709 = n1190 & ~n2708 ;
  assign n2710 = n1635 & ~n1997 ;
  assign n2711 = ~n2706 & ~n2710 ;
  assign n2712 = n1370 & ~n2711 ;
  assign n2713 = n1635 & n2139 ;
  assign n2714 = \reg1_reg[24]/NET0131  & ~n2667 ;
  assign n2721 = ~n2713 & ~n2714 ;
  assign n2722 = ~n2712 & n2721 ;
  assign n2723 = ~n2709 & n2722 ;
  assign n2715 = n1635 & n2007 ;
  assign n2716 = ~n2706 & ~n2715 ;
  assign n2717 = n1326 & ~n2716 ;
  assign n2718 = n1635 & ~n2021 ;
  assign n2719 = ~n2706 & ~n2718 ;
  assign n2720 = n1292 & ~n2719 ;
  assign n2724 = ~n2717 & ~n2720 ;
  assign n2725 = n2723 & n2724 ;
  assign n2726 = n1386 & ~n2725 ;
  assign n2727 = ~n2705 & ~n2726 ;
  assign n2728 = \state_reg[0]/NET0131  & ~n2727 ;
  assign n2729 = ~n2704 & ~n2728 ;
  assign n2730 = \reg1_reg[25]/NET0131  & ~n1426 ;
  assign n2731 = \reg1_reg[25]/NET0131  & n1388 ;
  assign n2732 = ~n1190 & ~n1292 ;
  assign n2733 = ~n1635 & ~n2732 ;
  assign n2734 = n1647 & ~n2733 ;
  assign n2735 = \reg1_reg[25]/NET0131  & ~n2734 ;
  assign n2739 = ~n1539 & n1544 ;
  assign n2740 = n1530 & ~n2739 ;
  assign n2741 = n1558 & n2740 ;
  assign n2736 = ~n1549 & n1557 ;
  assign n2737 = n1564 & ~n2736 ;
  assign n2738 = n1554 & ~n2737 ;
  assign n2742 = ~n1570 & ~n2738 ;
  assign n2743 = ~n2741 & n2742 ;
  assign n2744 = n1574 & ~n2743 ;
  assign n2745 = n1582 & ~n2744 ;
  assign n2746 = n1080 & ~n2745 ;
  assign n2747 = ~n1080 & n2745 ;
  assign n2748 = ~n2746 & ~n2747 ;
  assign n2749 = n1190 & ~n2748 ;
  assign n2757 = n1459 & n1485 ;
  assign n2758 = n1455 & ~n1466 ;
  assign n2759 = n1493 & ~n2758 ;
  assign n2760 = n1458 & ~n2759 ;
  assign n2761 = ~n1500 & ~n2760 ;
  assign n2762 = ~n2757 & n2761 ;
  assign n2763 = n1505 & ~n2762 ;
  assign n2764 = n1517 & ~n2763 ;
  assign n2765 = n1080 & n2764 ;
  assign n2766 = ~n1080 & ~n2764 ;
  assign n2767 = ~n2765 & ~n2766 ;
  assign n2768 = n1292 & ~n2767 ;
  assign n2750 = n454 & ~n1771 ;
  assign n2751 = ~n2495 & ~n2750 ;
  assign n2752 = ~n338 & ~n2751 ;
  assign n2753 = n338 & n441 ;
  assign n2754 = ~n2752 & ~n2753 ;
  assign n2755 = n1370 & n2754 ;
  assign n2756 = n417 & n1328 ;
  assign n2769 = n417 & ~n1317 ;
  assign n2770 = ~n2524 & ~n2769 ;
  assign n2771 = n1326 & n2770 ;
  assign n2772 = ~n2756 & ~n2771 ;
  assign n2773 = ~n2755 & n2772 ;
  assign n2774 = ~n2768 & n2773 ;
  assign n2775 = ~n2749 & n2774 ;
  assign n2776 = n1635 & ~n2775 ;
  assign n2777 = ~n2735 & ~n2776 ;
  assign n2778 = n1386 & ~n2777 ;
  assign n2779 = ~n2731 & ~n2778 ;
  assign n2780 = \state_reg[0]/NET0131  & ~n2779 ;
  assign n2781 = ~n2730 & ~n2780 ;
  assign n2782 = \reg2_reg[12]/NET0131  & ~n1426 ;
  assign n2783 = \reg2_reg[12]/NET0131  & n1388 ;
  assign n2785 = \reg2_reg[12]/NET0131  & ~n1396 ;
  assign n2786 = n1396 & n1939 ;
  assign n2787 = ~n2785 & ~n2786 ;
  assign n2788 = n1190 & ~n2787 ;
  assign n2792 = n1396 & ~n1954 ;
  assign n2793 = ~n2785 & ~n2792 ;
  assign n2794 = n1292 & ~n2793 ;
  assign n2789 = n1396 & n1948 ;
  assign n2790 = ~n2785 & ~n2789 ;
  assign n2791 = n1370 & ~n2790 ;
  assign n2795 = n1396 & n1960 ;
  assign n2796 = ~n2785 & ~n2795 ;
  assign n2797 = n1326 & ~n2796 ;
  assign n2799 = \reg2_reg[12]/NET0131  & ~n1414 ;
  assign n2784 = n1396 & n2651 ;
  assign n2798 = n537 & n1331 ;
  assign n2800 = ~n2784 & ~n2798 ;
  assign n2801 = ~n2799 & n2800 ;
  assign n2802 = ~n2797 & n2801 ;
  assign n2803 = ~n2791 & n2802 ;
  assign n2804 = ~n2794 & n2803 ;
  assign n2805 = ~n2788 & n2804 ;
  assign n2806 = n1386 & ~n2805 ;
  assign n2807 = ~n2783 & ~n2806 ;
  assign n2808 = \state_reg[0]/NET0131  & ~n2807 ;
  assign n2809 = ~n2782 & ~n2808 ;
  assign n2810 = \reg2_reg[11]/NET0131  & ~n1426 ;
  assign n2811 = \reg2_reg[11]/NET0131  & n1388 ;
  assign n2813 = \reg2_reg[11]/NET0131  & ~n1396 ;
  assign n2814 = n1396 & n1895 ;
  assign n2815 = ~n2813 & ~n2814 ;
  assign n2816 = n1190 & ~n2815 ;
  assign n2820 = n1396 & n1910 ;
  assign n2821 = ~n2813 & ~n2820 ;
  assign n2822 = n1370 & ~n2821 ;
  assign n2817 = n1396 & ~n1901 ;
  assign n2818 = ~n2813 & ~n2817 ;
  assign n2819 = n1292 & ~n2818 ;
  assign n2823 = n1396 & n1917 ;
  assign n2824 = ~n2813 & ~n2823 ;
  assign n2825 = n1326 & ~n2824 ;
  assign n2812 = \reg2_reg[11]/NET0131  & ~n1414 ;
  assign n2826 = n1396 & n2637 ;
  assign n2827 = n575 & n1331 ;
  assign n2828 = ~n2826 & ~n2827 ;
  assign n2829 = ~n2812 & n2828 ;
  assign n2830 = ~n2825 & n2829 ;
  assign n2831 = ~n2819 & n2830 ;
  assign n2832 = ~n2822 & n2831 ;
  assign n2833 = ~n2816 & n2832 ;
  assign n2834 = n1386 & ~n2833 ;
  assign n2835 = ~n2811 & ~n2834 ;
  assign n2836 = \state_reg[0]/NET0131  & ~n2835 ;
  assign n2837 = ~n2810 & ~n2836 ;
  assign n2838 = \reg0_reg[11]/NET0131  & ~n1426 ;
  assign n2839 = \reg0_reg[11]/NET0131  & n1388 ;
  assign n2841 = \reg0_reg[11]/NET0131  & ~n1607 ;
  assign n2842 = n1607 & n1895 ;
  assign n2843 = ~n2841 & ~n2842 ;
  assign n2844 = n1190 & ~n2843 ;
  assign n2848 = n1607 & n1910 ;
  assign n2849 = ~n2841 & ~n2848 ;
  assign n2850 = n1370 & ~n2849 ;
  assign n2845 = n1607 & ~n1901 ;
  assign n2846 = ~n2841 & ~n2845 ;
  assign n2847 = n1292 & ~n2846 ;
  assign n2840 = \reg0_reg[11]/NET0131  & ~n1623 ;
  assign n2851 = n1607 & ~n2639 ;
  assign n2852 = ~n2840 & ~n2851 ;
  assign n2853 = ~n2847 & n2852 ;
  assign n2854 = ~n2850 & n2853 ;
  assign n2855 = ~n2844 & n2854 ;
  assign n2856 = n1386 & ~n2855 ;
  assign n2857 = ~n2839 & ~n2856 ;
  assign n2858 = \state_reg[0]/NET0131  & ~n2857 ;
  assign n2859 = ~n2838 & ~n2858 ;
  assign n2860 = \reg2_reg[20]/NET0131  & ~n1426 ;
  assign n2861 = \reg2_reg[20]/NET0131  & n1388 ;
  assign n2863 = \reg2_reg[20]/NET0131  & ~n1396 ;
  assign n2864 = n1396 & ~n2434 ;
  assign n2865 = ~n2863 & ~n2864 ;
  assign n2866 = n1190 & ~n2865 ;
  assign n2870 = n1396 & ~n2449 ;
  assign n2871 = ~n2863 & ~n2870 ;
  assign n2872 = n1292 & ~n2871 ;
  assign n2867 = n1396 & n2443 ;
  assign n2868 = ~n2863 & ~n2867 ;
  assign n2869 = n1370 & ~n2868 ;
  assign n2873 = n1396 & n2454 ;
  assign n2874 = ~n2863 & ~n2873 ;
  assign n2875 = n1326 & ~n2874 ;
  assign n2877 = \reg2_reg[20]/NET0131  & ~n1414 ;
  assign n2862 = n1396 & n2587 ;
  assign n2876 = n847 & n1331 ;
  assign n2878 = ~n2862 & ~n2876 ;
  assign n2879 = ~n2877 & n2878 ;
  assign n2880 = ~n2875 & n2879 ;
  assign n2881 = ~n2869 & n2880 ;
  assign n2882 = ~n2872 & n2881 ;
  assign n2883 = ~n2866 & n2882 ;
  assign n2884 = n1386 & ~n2883 ;
  assign n2885 = ~n2861 & ~n2884 ;
  assign n2886 = \state_reg[0]/NET0131  & ~n2885 ;
  assign n2887 = ~n2860 & ~n2886 ;
  assign n2888 = \reg0_reg[12]/NET0131  & ~n1426 ;
  assign n2889 = \reg0_reg[12]/NET0131  & n1388 ;
  assign n2891 = \reg0_reg[12]/NET0131  & ~n1607 ;
  assign n2892 = n1607 & n1939 ;
  assign n2893 = ~n2891 & ~n2892 ;
  assign n2894 = n1190 & ~n2893 ;
  assign n2898 = n1607 & ~n1954 ;
  assign n2899 = ~n2891 & ~n2898 ;
  assign n2900 = n1292 & ~n2899 ;
  assign n2895 = n1607 & n1948 ;
  assign n2896 = ~n2891 & ~n2895 ;
  assign n2897 = n1370 & ~n2896 ;
  assign n2901 = n1607 & n1960 ;
  assign n2902 = ~n2891 & ~n2901 ;
  assign n2903 = n1326 & ~n2902 ;
  assign n2890 = n1607 & n2651 ;
  assign n2904 = \reg0_reg[12]/NET0131  & ~n2142 ;
  assign n2905 = ~n2890 & ~n2904 ;
  assign n2906 = ~n2903 & n2905 ;
  assign n2907 = ~n2897 & n2906 ;
  assign n2908 = ~n2900 & n2907 ;
  assign n2909 = ~n2894 & n2908 ;
  assign n2910 = n1386 & ~n2909 ;
  assign n2911 = ~n2889 & ~n2910 ;
  assign n2912 = \state_reg[0]/NET0131  & ~n2911 ;
  assign n2913 = ~n2888 & ~n2912 ;
  assign n2914 = \reg2_reg[24]/NET0131  & ~n1426 ;
  assign n2915 = \reg2_reg[24]/NET0131  & n1388 ;
  assign n2916 = \reg2_reg[24]/NET0131  & ~n1396 ;
  assign n2917 = n1396 & ~n1987 ;
  assign n2918 = ~n2916 & ~n2917 ;
  assign n2919 = n1190 & ~n2918 ;
  assign n2920 = n1396 & ~n1997 ;
  assign n2921 = ~n2916 & ~n2920 ;
  assign n2922 = n1370 & ~n2921 ;
  assign n2931 = \reg2_reg[24]/NET0131  & ~n1414 ;
  assign n2929 = n1396 & n2139 ;
  assign n2930 = n437 & n1331 ;
  assign n2932 = ~n2929 & ~n2930 ;
  assign n2933 = ~n2931 & n2932 ;
  assign n2934 = ~n2922 & n2933 ;
  assign n2935 = ~n2919 & n2934 ;
  assign n2923 = n1396 & n2007 ;
  assign n2924 = ~n2916 & ~n2923 ;
  assign n2925 = n1326 & ~n2924 ;
  assign n2926 = n1396 & ~n2021 ;
  assign n2927 = ~n2916 & ~n2926 ;
  assign n2928 = n1292 & ~n2927 ;
  assign n2936 = ~n2925 & ~n2928 ;
  assign n2937 = n2935 & n2936 ;
  assign n2938 = n1386 & ~n2937 ;
  assign n2939 = ~n2915 & ~n2938 ;
  assign n2940 = \state_reg[0]/NET0131  & ~n2939 ;
  assign n2941 = ~n2914 & ~n2940 ;
  assign n2943 = n291 & n1388 ;
  assign n2954 = ~n1077 & n1551 ;
  assign n2953 = n1077 & ~n1551 ;
  assign n2955 = n1190 & ~n2953 ;
  assign n2956 = ~n2954 & n2955 ;
  assign n2945 = n530 & ~n1959 ;
  assign n2946 = ~n530 & n1959 ;
  assign n2947 = ~n2945 & ~n2946 ;
  assign n2948 = n1326 & ~n2947 ;
  assign n2950 = ~n1077 & ~n1486 ;
  assign n2949 = n1077 & n1486 ;
  assign n2951 = n1292 & ~n2949 ;
  assign n2952 = ~n2950 & n2951 ;
  assign n2957 = ~n2948 & ~n2952 ;
  assign n2958 = ~n2956 & n2957 ;
  assign n2959 = n1169 & ~n2958 ;
  assign n2964 = n498 & ~n1944 ;
  assign n2965 = ~n2243 & ~n2964 ;
  assign n2966 = ~n338 & ~n2965 ;
  assign n2967 = n338 & n541 ;
  assign n2968 = ~n2966 & ~n2967 ;
  assign n2969 = n1169 & ~n2968 ;
  assign n2970 = ~n291 & ~n1169 ;
  assign n2971 = n1370 & ~n2970 ;
  assign n2972 = ~n2969 & n2971 ;
  assign n2944 = ~n530 & ~n1332 ;
  assign n2960 = ~n1326 & n2732 ;
  assign n2961 = ~n1169 & ~n2960 ;
  assign n2962 = n1375 & ~n2961 ;
  assign n2963 = n291 & ~n2962 ;
  assign n2973 = ~n2944 & ~n2963 ;
  assign n2974 = ~n2972 & n2973 ;
  assign n2975 = ~n2959 & n2974 ;
  assign n2976 = n1386 & ~n2975 ;
  assign n2977 = ~n2943 & ~n2976 ;
  assign n2978 = \state_reg[0]/NET0131  & ~n2977 ;
  assign n2942 = n291 & n311 ;
  assign n2979 = \reg3_reg[13]/NET0131  & ~\state_reg[0]/NET0131  ;
  assign n2980 = ~n2942 & ~n2979 ;
  assign n2981 = ~n2978 & n2980 ;
  assign n2984 = n857 & n1388 ;
  assign n2987 = n857 & ~n1169 ;
  assign n2988 = n827 & ~n2316 ;
  assign n2989 = ~n827 & n2316 ;
  assign n2990 = ~n2988 & ~n2989 ;
  assign n2991 = ~n338 & ~n2990 ;
  assign n2992 = n338 & n887 ;
  assign n2993 = ~n2991 & ~n2992 ;
  assign n2994 = n1169 & n2993 ;
  assign n2995 = ~n2987 & ~n2994 ;
  assign n2996 = n1370 & ~n2995 ;
  assign n3013 = n871 & ~n2325 ;
  assign n3014 = ~n1310 & ~n3013 ;
  assign n3015 = n1169 & n3014 ;
  assign n3016 = ~n2987 & ~n3015 ;
  assign n3017 = n1326 & ~n3016 ;
  assign n2985 = n871 & ~n1332 ;
  assign n2986 = n857 & ~n1375 ;
  assign n3018 = ~n2985 & ~n2986 ;
  assign n3019 = ~n3017 & n3018 ;
  assign n3020 = ~n2996 & n3019 ;
  assign n2997 = n1557 & n2740 ;
  assign n2998 = n2737 & ~n2997 ;
  assign n2999 = n1043 & ~n2998 ;
  assign n3000 = ~n1043 & n2998 ;
  assign n3001 = ~n2999 & ~n3000 ;
  assign n3002 = n1169 & ~n3001 ;
  assign n3003 = ~n2987 & ~n3002 ;
  assign n3004 = n1190 & ~n3003 ;
  assign n3005 = n1455 & ~n1486 ;
  assign n3006 = n1493 & ~n3005 ;
  assign n3007 = n1043 & ~n3006 ;
  assign n3008 = ~n1043 & n3006 ;
  assign n3009 = ~n3007 & ~n3008 ;
  assign n3010 = n1169 & n3009 ;
  assign n3011 = ~n2987 & ~n3010 ;
  assign n3012 = n1292 & ~n3011 ;
  assign n3021 = ~n3004 & ~n3012 ;
  assign n3022 = n3020 & n3021 ;
  assign n3023 = n1386 & ~n3022 ;
  assign n3024 = ~n2984 & ~n3023 ;
  assign n3025 = \state_reg[0]/NET0131  & ~n3024 ;
  assign n2982 = \reg3_reg[17]/NET0131  & ~\state_reg[0]/NET0131  ;
  assign n2983 = n311 & n857 ;
  assign n3026 = ~n2982 & ~n2983 ;
  assign n3027 = ~n3025 & n3026 ;
  assign n3029 = ~n725 & ~n1332 ;
  assign n3030 = ~n743 & ~n1532 ;
  assign n3032 = n1067 & ~n3030 ;
  assign n3031 = ~n1067 & n3030 ;
  assign n3033 = n1190 & ~n3031 ;
  assign n3034 = ~n3032 & n3033 ;
  assign n3037 = ~n1066 & n1470 ;
  assign n3035 = ~n1222 & ~n1469 ;
  assign n3036 = ~n1067 & ~n3035 ;
  assign n3038 = n1292 & ~n3036 ;
  assign n3039 = ~n3037 & n3038 ;
  assign n3040 = ~n725 & ~n1295 ;
  assign n3041 = ~n1296 & n1326 ;
  assign n3042 = ~n3040 & n3041 ;
  assign n3043 = ~n3039 & ~n3042 ;
  assign n3044 = ~n3034 & n3043 ;
  assign n3045 = n708 & ~n1337 ;
  assign n3046 = ~n708 & n1337 ;
  assign n3047 = ~n3045 & ~n3046 ;
  assign n3048 = ~n338 & ~n3047 ;
  assign n3049 = n338 & n735 ;
  assign n3050 = n1370 & ~n3049 ;
  assign n3051 = ~n3048 & n3050 ;
  assign n3052 = n3044 & ~n3051 ;
  assign n3053 = n1169 & ~n3052 ;
  assign n3054 = ~n3029 & ~n3053 ;
  assign n3055 = ~n1385 & ~n3054 ;
  assign n3056 = ~n1169 & ~n2732 ;
  assign n3057 = ~n1385 & ~n3056 ;
  assign n3058 = n2345 & n3057 ;
  assign n3059 = ~\reg3_reg[3]/NET0131  & ~n3058 ;
  assign n3060 = ~n3055 & ~n3059 ;
  assign n3061 = n1426 & ~n3060 ;
  assign n3028 = \reg3_reg[3]/NET0131  & ~\state_reg[0]/NET0131  ;
  assign n3062 = ~\reg3_reg[3]/NET0131  & n311 ;
  assign n3063 = ~n3028 & ~n3062 ;
  assign n3064 = ~n3061 & n3063 ;
  assign n3067 = n275 & n1388 ;
  assign n3069 = n275 & ~n1169 ;
  assign n3070 = ~n661 & n1339 ;
  assign n3071 = n661 & ~n1339 ;
  assign n3072 = ~n3070 & ~n3071 ;
  assign n3073 = ~n338 & ~n3072 ;
  assign n3074 = n338 & n708 ;
  assign n3075 = ~n3073 & ~n3074 ;
  assign n3076 = n1169 & n3075 ;
  assign n3077 = ~n3069 & ~n3076 ;
  assign n3078 = n1370 & ~n3077 ;
  assign n3085 = ~n1215 & ~n1472 ;
  assign n3086 = n1039 & ~n3085 ;
  assign n3087 = ~n1039 & n3085 ;
  assign n3088 = ~n3086 & ~n3087 ;
  assign n3089 = n1169 & ~n3088 ;
  assign n3090 = ~n3069 & ~n3089 ;
  assign n3091 = n1292 & ~n3090 ;
  assign n3079 = n1039 & n1536 ;
  assign n3080 = ~n1039 & ~n1536 ;
  assign n3081 = ~n3079 & ~n3080 ;
  assign n3082 = n1169 & n3081 ;
  assign n3083 = ~n3069 & ~n3082 ;
  assign n3084 = n1190 & ~n3083 ;
  assign n3092 = n690 & ~n1297 ;
  assign n3093 = ~n1298 & ~n3092 ;
  assign n3094 = n1169 & n3093 ;
  assign n3095 = ~n3069 & ~n3094 ;
  assign n3096 = n1326 & ~n3095 ;
  assign n3068 = n690 & ~n1332 ;
  assign n3097 = n275 & ~n1375 ;
  assign n3098 = ~n3068 & ~n3097 ;
  assign n3099 = ~n3096 & n3098 ;
  assign n3100 = ~n3084 & n3099 ;
  assign n3101 = ~n3091 & n3100 ;
  assign n3102 = ~n3078 & n3101 ;
  assign n3103 = n1386 & ~n3102 ;
  assign n3104 = ~n3067 & ~n3103 ;
  assign n3105 = \state_reg[0]/NET0131  & ~n3104 ;
  assign n3065 = \reg3_reg[5]/NET0131  & ~\state_reg[0]/NET0131  ;
  assign n3066 = n275 & n311 ;
  assign n3106 = ~n3065 & ~n3066 ;
  assign n3107 = ~n3105 & n3106 ;
  assign n3110 = n611 & n1388 ;
  assign n3127 = ~n618 & n2355 ;
  assign n3128 = n592 & ~n3127 ;
  assign n3129 = ~n592 & n3127 ;
  assign n3130 = ~n3128 & ~n3129 ;
  assign n3131 = ~n338 & ~n3130 ;
  assign n3126 = n338 & n628 ;
  assign n3132 = n1370 & ~n3126 ;
  assign n3133 = ~n3131 & n3132 ;
  assign n3113 = ~n635 & n1300 ;
  assign n3114 = ~n609 & ~n3113 ;
  assign n3115 = ~n1302 & n1326 ;
  assign n3116 = ~n3114 & n3115 ;
  assign n3118 = ~n1057 & ~n1482 ;
  assign n3117 = n1057 & n1482 ;
  assign n3119 = n1292 & ~n3117 ;
  assign n3120 = ~n3118 & n3119 ;
  assign n3121 = ~n3116 & ~n3120 ;
  assign n3123 = n1057 & ~n2739 ;
  assign n3122 = ~n1057 & n2739 ;
  assign n3124 = n1190 & ~n3122 ;
  assign n3125 = ~n3123 & n3124 ;
  assign n3134 = n3121 & ~n3125 ;
  assign n3135 = ~n3133 & n3134 ;
  assign n3136 = n1169 & ~n3135 ;
  assign n3111 = ~n609 & ~n1332 ;
  assign n3112 = n611 & ~n2286 ;
  assign n3137 = ~n3111 & ~n3112 ;
  assign n3138 = ~n3136 & n3137 ;
  assign n3139 = n1386 & ~n3138 ;
  assign n3140 = ~n3110 & ~n3139 ;
  assign n3141 = \state_reg[0]/NET0131  & ~n3140 ;
  assign n3108 = \reg3_reg[9]/NET0131  & ~\state_reg[0]/NET0131  ;
  assign n3109 = n311 & n611 ;
  assign n3142 = ~n3108 & ~n3109 ;
  assign n3143 = ~n3141 & n3142 ;
  assign n3144 = n482 & n1388 ;
  assign n3145 = n482 & ~n1169 ;
  assign n3146 = ~n2262 & n2504 ;
  assign n3147 = n2509 & ~n3146 ;
  assign n3148 = n2501 & ~n3147 ;
  assign n3149 = n2513 & ~n3148 ;
  assign n3150 = n1070 & n3149 ;
  assign n3151 = ~n1070 & ~n3149 ;
  assign n3152 = ~n3150 & ~n3151 ;
  assign n3153 = n1169 & ~n3152 ;
  assign n3154 = ~n3145 & ~n3153 ;
  assign n3155 = n1292 & ~n3154 ;
  assign n3156 = n2471 & n2474 ;
  assign n3157 = ~n2275 & n3156 ;
  assign n3158 = ~n2470 & n2474 ;
  assign n3159 = n2480 & ~n3158 ;
  assign n3160 = ~n3157 & n3159 ;
  assign n3161 = n1070 & n3160 ;
  assign n3162 = ~n1070 & ~n3160 ;
  assign n3163 = ~n3161 & ~n3162 ;
  assign n3164 = n1169 & n3163 ;
  assign n3165 = ~n3145 & ~n3164 ;
  assign n3166 = n1190 & ~n3165 ;
  assign n3167 = n1354 & n2401 ;
  assign n3168 = n474 & ~n3167 ;
  assign n3169 = ~n1992 & ~n3168 ;
  assign n3170 = ~n338 & ~n3169 ;
  assign n3171 = n338 & n840 ;
  assign n3172 = ~n3170 & ~n3171 ;
  assign n3173 = n1169 & n3172 ;
  assign n3174 = ~n3145 & ~n3173 ;
  assign n3175 = n1370 & ~n3174 ;
  assign n3177 = n476 & ~n2003 ;
  assign n3178 = n1326 & ~n2004 ;
  assign n3179 = ~n3177 & n3178 ;
  assign n3180 = n1169 & n3179 ;
  assign n3176 = n482 & ~n2345 ;
  assign n3181 = n476 & ~n1332 ;
  assign n3182 = ~n3176 & ~n3181 ;
  assign n3183 = ~n3180 & n3182 ;
  assign n3184 = ~n3175 & n3183 ;
  assign n3185 = ~n3166 & n3184 ;
  assign n3186 = ~n3155 & n3185 ;
  assign n3187 = n1386 & ~n3186 ;
  assign n3188 = ~n3144 & ~n3187 ;
  assign n3189 = \state_reg[0]/NET0131  & ~n3188 ;
  assign n3190 = \reg3_reg[22]/NET0131  & ~\state_reg[0]/NET0131  ;
  assign n3191 = n311 & n482 ;
  assign n3192 = ~n3190 & ~n3191 ;
  assign n3193 = ~n3189 & n3192 ;
  assign n3194 = \reg2_reg[30]/NET0131  & ~n2561 ;
  assign n3195 = n367 & n1328 ;
  assign n3196 = n367 & ~n1433 ;
  assign n3197 = ~n2549 & ~n3196 ;
  assign n3198 = n1326 & n3197 ;
  assign n3199 = ~n3195 & ~n3198 ;
  assign n3200 = ~n2548 & n3199 ;
  assign n3201 = n1396 & ~n3200 ;
  assign n3202 = ~n1449 & ~n3201 ;
  assign n3203 = n1717 & ~n3202 ;
  assign n3204 = ~n3194 & ~n3203 ;
  assign n3205 = \reg2_reg[7]/NET0131  & ~n1426 ;
  assign n3206 = \reg2_reg[7]/NET0131  & n1388 ;
  assign n3210 = \reg2_reg[7]/NET0131  & ~n1396 ;
  assign n3214 = n1396 & n2350 ;
  assign n3215 = ~n3210 & ~n3214 ;
  assign n3216 = n1190 & ~n3215 ;
  assign n3211 = n1396 & n2359 ;
  assign n3212 = ~n3210 & ~n3211 ;
  assign n3213 = n1370 & ~n3212 ;
  assign n3217 = n1396 & ~n2365 ;
  assign n3218 = ~n3210 & ~n3217 ;
  assign n3219 = n1292 & ~n3218 ;
  assign n3207 = n679 & n1328 ;
  assign n3208 = ~n2372 & ~n3207 ;
  assign n3209 = n1396 & ~n3208 ;
  assign n3220 = n666 & n1331 ;
  assign n3221 = \reg2_reg[7]/NET0131  & ~n2208 ;
  assign n3222 = ~n3220 & ~n3221 ;
  assign n3223 = ~n3209 & n3222 ;
  assign n3224 = ~n3219 & n3223 ;
  assign n3225 = ~n3213 & n3224 ;
  assign n3226 = ~n3216 & n3225 ;
  assign n3227 = n1386 & ~n3226 ;
  assign n3228 = ~n3206 & ~n3227 ;
  assign n3229 = \state_reg[0]/NET0131  & ~n3228 ;
  assign n3230 = ~n3205 & ~n3229 ;
  assign n3231 = ~n1291 & ~n1369 ;
  assign n3232 = ~n1607 & ~n3231 ;
  assign n3233 = n1717 & ~n3232 ;
  assign n3234 = n1623 & n3233 ;
  assign n3235 = \reg0_reg[14]/NET0131  & ~n3234 ;
  assign n3236 = ~n504 & n1328 ;
  assign n3237 = n2282 & ~n3236 ;
  assign n3238 = n2621 & ~n3237 ;
  assign n3239 = ~n3235 & ~n3238 ;
  assign n3240 = \reg0_reg[16]/NET0131  & ~n1426 ;
  assign n3241 = \reg0_reg[16]/NET0131  & n1388 ;
  assign n3243 = \reg0_reg[16]/NET0131  & ~n1607 ;
  assign n3247 = n1607 & n2311 ;
  assign n3248 = ~n3243 & ~n3247 ;
  assign n3249 = n1190 & ~n3248 ;
  assign n3244 = n1607 & n2305 ;
  assign n3245 = ~n3243 & ~n3244 ;
  assign n3246 = n1292 & ~n3245 ;
  assign n3250 = n1607 & n2320 ;
  assign n3251 = ~n3243 & ~n3250 ;
  assign n3252 = n1370 & ~n3251 ;
  assign n3242 = \reg0_reg[16]/NET0131  & ~n1623 ;
  assign n3253 = n878 & n1328 ;
  assign n3254 = n1326 & n2326 ;
  assign n3255 = ~n3253 & ~n3254 ;
  assign n3256 = n1607 & ~n3255 ;
  assign n3257 = ~n3242 & ~n3256 ;
  assign n3258 = ~n3252 & n3257 ;
  assign n3259 = ~n3246 & n3258 ;
  assign n3260 = ~n3249 & n3259 ;
  assign n3261 = n1386 & ~n3260 ;
  assign n3262 = ~n3241 & ~n3261 ;
  assign n3263 = \state_reg[0]/NET0131  & ~n3262 ;
  assign n3264 = ~n3240 & ~n3263 ;
  assign n3266 = \reg0_reg[19]/NET0131  & ~n1607 ;
  assign n3267 = n1607 & n2391 ;
  assign n3268 = ~n3266 & ~n3267 ;
  assign n3269 = n1292 & ~n3268 ;
  assign n3270 = n1607 & ~n2397 ;
  assign n3271 = ~n3266 & ~n3270 ;
  assign n3272 = n1190 & ~n3271 ;
  assign n3265 = \reg0_reg[19]/NET0131  & ~n1624 ;
  assign n3274 = n1370 & n2406 ;
  assign n3273 = n1326 & n2413 ;
  assign n3275 = ~n797 & n1328 ;
  assign n3276 = ~n3273 & ~n3275 ;
  assign n3277 = ~n3274 & n3276 ;
  assign n3278 = n1607 & ~n3277 ;
  assign n3279 = ~n3265 & ~n3278 ;
  assign n3280 = ~n3272 & n3279 ;
  assign n3281 = ~n3269 & n3280 ;
  assign n3282 = n1386 & ~n3281 ;
  assign n3283 = \reg0_reg[19]/NET0131  & n1388 ;
  assign n3284 = ~n3282 & ~n3283 ;
  assign n3285 = \state_reg[0]/NET0131  & ~n3284 ;
  assign n3286 = \reg0_reg[19]/NET0131  & ~n1426 ;
  assign n3287 = ~n3285 & ~n3286 ;
  assign n3289 = \reg0_reg[25]/NET0131  & ~n1607 ;
  assign n3290 = n2621 & ~n2748 ;
  assign n3291 = ~n3289 & ~n3290 ;
  assign n3292 = n1190 & ~n3291 ;
  assign n3288 = n2621 & ~n2774 ;
  assign n3293 = n1292 & ~n1607 ;
  assign n3294 = n1717 & ~n3293 ;
  assign n3295 = n1624 & n3294 ;
  assign n3296 = \reg0_reg[25]/NET0131  & ~n3295 ;
  assign n3297 = ~n3288 & ~n3296 ;
  assign n3298 = ~n3292 & n3297 ;
  assign n3299 = \reg0_reg[30]/NET0131  & ~n3234 ;
  assign n3300 = n2621 & ~n3199 ;
  assign n3301 = ~n3299 & ~n3300 ;
  assign n3302 = \reg0_reg[31]/NET0131  & ~n3234 ;
  assign n3303 = ~n2555 & n2621 ;
  assign n3304 = ~n3302 & ~n3303 ;
  assign n3305 = \reg0_reg[7]/NET0131  & ~n1426 ;
  assign n3306 = \reg0_reg[7]/NET0131  & n1388 ;
  assign n3308 = \reg0_reg[7]/NET0131  & ~n1607 ;
  assign n3312 = n1607 & n2359 ;
  assign n3313 = ~n3308 & ~n3312 ;
  assign n3314 = n1370 & ~n3313 ;
  assign n3309 = n1607 & n2350 ;
  assign n3310 = ~n3308 & ~n3309 ;
  assign n3311 = n1190 & ~n3310 ;
  assign n3315 = n1607 & ~n2365 ;
  assign n3316 = ~n3308 & ~n3315 ;
  assign n3317 = n1292 & ~n3316 ;
  assign n3307 = \reg0_reg[7]/NET0131  & ~n1623 ;
  assign n3318 = n1607 & ~n3208 ;
  assign n3319 = ~n3307 & ~n3318 ;
  assign n3320 = ~n3317 & n3319 ;
  assign n3321 = ~n3311 & n3320 ;
  assign n3322 = ~n3314 & n3321 ;
  assign n3323 = n1386 & ~n3322 ;
  assign n3324 = ~n3306 & ~n3323 ;
  assign n3325 = \state_reg[0]/NET0131  & ~n3324 ;
  assign n3326 = ~n3305 & ~n3325 ;
  assign n3327 = \reg0_reg[8]/NET0131  & ~n1426 ;
  assign n3328 = \reg0_reg[8]/NET0131  & n1388 ;
  assign n3330 = \reg0_reg[8]/NET0131  & ~n1607 ;
  assign n3339 = n979 & n1035 ;
  assign n3340 = ~n979 & ~n1035 ;
  assign n3341 = ~n3339 & ~n3340 ;
  assign n3342 = n1607 & n3341 ;
  assign n3343 = ~n3330 & ~n3342 ;
  assign n3344 = n1190 & ~n3343 ;
  assign n3331 = n618 & ~n2355 ;
  assign n3332 = ~n3127 & ~n3331 ;
  assign n3333 = ~n338 & ~n3332 ;
  assign n3334 = n338 & n671 ;
  assign n3335 = ~n3333 & ~n3334 ;
  assign n3336 = n1607 & n3335 ;
  assign n3337 = ~n3330 & ~n3336 ;
  assign n3338 = n1370 & ~n3337 ;
  assign n3345 = n1035 & n1239 ;
  assign n3346 = ~n1035 & ~n1239 ;
  assign n3347 = ~n3345 & ~n3346 ;
  assign n3348 = n1607 & ~n3347 ;
  assign n3349 = ~n3330 & ~n3348 ;
  assign n3350 = n1292 & ~n3349 ;
  assign n3329 = \reg0_reg[8]/NET0131  & ~n1623 ;
  assign n3351 = n635 & n1328 ;
  assign n3352 = n635 & ~n1300 ;
  assign n3353 = n1326 & ~n3113 ;
  assign n3354 = ~n3352 & n3353 ;
  assign n3355 = ~n3351 & ~n3354 ;
  assign n3356 = n1607 & ~n3355 ;
  assign n3357 = ~n3329 & ~n3356 ;
  assign n3358 = ~n3350 & n3357 ;
  assign n3359 = ~n3338 & n3358 ;
  assign n3360 = ~n3344 & n3359 ;
  assign n3361 = n1386 & ~n3360 ;
  assign n3362 = ~n3328 & ~n3361 ;
  assign n3363 = \state_reg[0]/NET0131  & ~n3362 ;
  assign n3364 = ~n3327 & ~n3363 ;
  assign n3365 = ~n1635 & ~n3231 ;
  assign n3366 = n1717 & ~n3365 ;
  assign n3367 = n1646 & n3366 ;
  assign n3368 = \reg1_reg[14]/NET0131  & ~n3367 ;
  assign n3369 = n1635 & n1717 ;
  assign n3370 = ~n3237 & n3369 ;
  assign n3371 = ~n3368 & ~n3370 ;
  assign n3372 = \reg1_reg[16]/NET0131  & ~n1426 ;
  assign n3373 = \reg1_reg[16]/NET0131  & n1388 ;
  assign n3375 = \reg1_reg[16]/NET0131  & ~n1635 ;
  assign n3379 = n1635 & n2311 ;
  assign n3380 = ~n3375 & ~n3379 ;
  assign n3381 = n1190 & ~n3380 ;
  assign n3376 = n1635 & n2305 ;
  assign n3377 = ~n3375 & ~n3376 ;
  assign n3378 = n1292 & ~n3377 ;
  assign n3382 = n1635 & n2320 ;
  assign n3383 = ~n3375 & ~n3382 ;
  assign n3384 = n1370 & ~n3383 ;
  assign n3374 = \reg1_reg[16]/NET0131  & ~n1646 ;
  assign n3385 = n1635 & ~n3255 ;
  assign n3386 = ~n3374 & ~n3385 ;
  assign n3387 = ~n3384 & n3386 ;
  assign n3388 = ~n3378 & n3387 ;
  assign n3389 = ~n3381 & n3388 ;
  assign n3390 = n1386 & ~n3389 ;
  assign n3391 = ~n3373 & ~n3390 ;
  assign n3392 = \state_reg[0]/NET0131  & ~n3391 ;
  assign n3393 = ~n3372 & ~n3392 ;
  assign n3394 = \reg1_reg[19]/NET0131  & ~n1426 ;
  assign n3396 = \reg1_reg[19]/NET0131  & ~n1635 ;
  assign n3397 = n1635 & n2391 ;
  assign n3398 = ~n3396 & ~n3397 ;
  assign n3399 = n1292 & ~n3398 ;
  assign n3400 = n1635 & ~n2397 ;
  assign n3401 = ~n3396 & ~n3400 ;
  assign n3402 = n1190 & ~n3401 ;
  assign n3395 = \reg1_reg[19]/NET0131  & ~n1647 ;
  assign n3403 = n1635 & ~n3277 ;
  assign n3404 = ~n3395 & ~n3403 ;
  assign n3405 = ~n3402 & n3404 ;
  assign n3406 = ~n3399 & n3405 ;
  assign n3407 = n1386 & ~n3406 ;
  assign n3408 = \reg1_reg[19]/NET0131  & n1388 ;
  assign n3409 = ~n3407 & ~n3408 ;
  assign n3410 = \state_reg[0]/NET0131  & ~n3409 ;
  assign n3411 = ~n3394 & ~n3410 ;
  assign n3412 = ~n2620 & n3369 ;
  assign n3414 = ~n1635 & ~n2531 ;
  assign n3415 = n2667 & ~n3414 ;
  assign n3413 = n1190 & ~n1635 ;
  assign n3416 = n1717 & ~n3413 ;
  assign n3417 = n3415 & n3416 ;
  assign n3418 = \reg1_reg[26]/NET0131  & ~n3417 ;
  assign n3419 = ~n3412 & ~n3418 ;
  assign n3422 = \reg1_reg[30]/NET0131  & ~n1635 ;
  assign n3423 = n3197 & n3369 ;
  assign n3424 = ~n3422 & ~n3423 ;
  assign n3425 = n1326 & ~n3424 ;
  assign n3420 = n2667 & n3366 ;
  assign n3421 = \reg1_reg[30]/NET0131  & ~n3420 ;
  assign n3426 = ~n2548 & ~n3195 ;
  assign n3427 = n3369 & ~n3426 ;
  assign n3428 = ~n3421 & ~n3427 ;
  assign n3429 = ~n3425 & n3428 ;
  assign n3430 = \reg1_reg[31]/NET0131  & ~n3367 ;
  assign n3431 = ~n2555 & n3369 ;
  assign n3432 = ~n3430 & ~n3431 ;
  assign n3433 = \reg1_reg[7]/NET0131  & ~n1426 ;
  assign n3434 = \reg1_reg[7]/NET0131  & n1388 ;
  assign n3436 = \reg1_reg[7]/NET0131  & ~n1635 ;
  assign n3440 = n1635 & n2359 ;
  assign n3441 = ~n3436 & ~n3440 ;
  assign n3442 = n1370 & ~n3441 ;
  assign n3437 = n1635 & n2350 ;
  assign n3438 = ~n3436 & ~n3437 ;
  assign n3439 = n1190 & ~n3438 ;
  assign n3443 = n1635 & ~n2365 ;
  assign n3444 = ~n3436 & ~n3443 ;
  assign n3445 = n1292 & ~n3444 ;
  assign n3435 = \reg1_reg[7]/NET0131  & ~n1646 ;
  assign n3446 = n1635 & ~n3208 ;
  assign n3447 = ~n3435 & ~n3446 ;
  assign n3448 = ~n3445 & n3447 ;
  assign n3449 = ~n3439 & n3448 ;
  assign n3450 = ~n3442 & n3449 ;
  assign n3451 = n1386 & ~n3450 ;
  assign n3452 = ~n3434 & ~n3451 ;
  assign n3453 = \state_reg[0]/NET0131  & ~n3452 ;
  assign n3454 = ~n3433 & ~n3453 ;
  assign n3455 = n1190 & ~n1396 ;
  assign n3456 = n1717 & ~n3455 ;
  assign n3457 = \reg2_reg[14]/NET0131  & ~n3456 ;
  assign n3459 = n1396 & ~n3237 ;
  assign n3458 = n493 & n1331 ;
  assign n3460 = n1131 & ~n1291 ;
  assign n3461 = ~n1396 & n3460 ;
  assign n3462 = n1414 & ~n3461 ;
  assign n3463 = ~n2573 & n3462 ;
  assign n3464 = \reg2_reg[14]/NET0131  & ~n3463 ;
  assign n3465 = ~n3458 & ~n3464 ;
  assign n3466 = ~n3459 & n3465 ;
  assign n3467 = n1717 & ~n3466 ;
  assign n3468 = ~n3457 & ~n3467 ;
  assign n3469 = \reg2_reg[16]/NET0131  & ~n1426 ;
  assign n3470 = \reg2_reg[16]/NET0131  & n1388 ;
  assign n3472 = \reg2_reg[16]/NET0131  & ~n1396 ;
  assign n3476 = n1396 & n2311 ;
  assign n3477 = ~n3472 & ~n3476 ;
  assign n3478 = n1190 & ~n3477 ;
  assign n3473 = n1396 & n2305 ;
  assign n3474 = ~n3472 & ~n3473 ;
  assign n3475 = n1292 & ~n3474 ;
  assign n3481 = n1396 & n2320 ;
  assign n3482 = ~n3472 & ~n3481 ;
  assign n3483 = n1370 & ~n3482 ;
  assign n3480 = n1396 & ~n3255 ;
  assign n3471 = n880 & n1331 ;
  assign n3479 = \reg2_reg[16]/NET0131  & ~n2208 ;
  assign n3484 = ~n3471 & ~n3479 ;
  assign n3485 = ~n3480 & n3484 ;
  assign n3486 = ~n3483 & n3485 ;
  assign n3487 = ~n3475 & n3486 ;
  assign n3488 = ~n3478 & n3487 ;
  assign n3489 = n1386 & ~n3488 ;
  assign n3490 = ~n3470 & ~n3489 ;
  assign n3491 = \state_reg[0]/NET0131  & ~n3490 ;
  assign n3492 = ~n3469 & ~n3491 ;
  assign n3493 = \reg2_reg[19]/NET0131  & ~n1426 ;
  assign n3494 = \reg2_reg[19]/NET0131  & n1388 ;
  assign n3497 = \reg2_reg[19]/NET0131  & ~n1396 ;
  assign n3498 = n1396 & n2391 ;
  assign n3499 = ~n3497 & ~n3498 ;
  assign n3500 = n1292 & ~n3499 ;
  assign n3501 = n1396 & ~n2397 ;
  assign n3502 = ~n3497 & ~n3501 ;
  assign n3503 = n1190 & ~n3502 ;
  assign n3504 = n1396 & ~n3277 ;
  assign n3495 = n802 & n1331 ;
  assign n3496 = \reg2_reg[19]/NET0131  & ~n3462 ;
  assign n3505 = ~n3495 & ~n3496 ;
  assign n3506 = ~n3504 & n3505 ;
  assign n3507 = ~n3503 & n3506 ;
  assign n3508 = ~n3500 & n3507 ;
  assign n3509 = n1386 & ~n3508 ;
  assign n3510 = ~n3494 & ~n3509 ;
  assign n3511 = \state_reg[0]/NET0131  & ~n3510 ;
  assign n3512 = ~n3493 & ~n3511 ;
  assign n3513 = \reg2_reg[25]/NET0131  & ~n1426 ;
  assign n3514 = \reg2_reg[25]/NET0131  & n1388 ;
  assign n3515 = \reg2_reg[25]/NET0131  & ~n1396 ;
  assign n3516 = n1396 & ~n2748 ;
  assign n3517 = ~n3515 & ~n3516 ;
  assign n3518 = n1190 & ~n3517 ;
  assign n3520 = n1396 & ~n2767 ;
  assign n3521 = ~n3515 & ~n3520 ;
  assign n3522 = n1292 & ~n3521 ;
  assign n3523 = n1396 & n2754 ;
  assign n3524 = ~n3515 & ~n3523 ;
  assign n3525 = n1370 & ~n3524 ;
  assign n3526 = n1396 & n2770 ;
  assign n3527 = ~n3515 & ~n3526 ;
  assign n3528 = n1326 & ~n3527 ;
  assign n3519 = \reg2_reg[25]/NET0131  & ~n1414 ;
  assign n3529 = n1396 & n2756 ;
  assign n3530 = n422 & n1331 ;
  assign n3531 = ~n3529 & ~n3530 ;
  assign n3532 = ~n3519 & n3531 ;
  assign n3533 = ~n3528 & n3532 ;
  assign n3534 = ~n3525 & n3533 ;
  assign n3535 = ~n3522 & n3534 ;
  assign n3536 = ~n3518 & n3535 ;
  assign n3537 = n1386 & ~n3536 ;
  assign n3538 = ~n3514 & ~n3537 ;
  assign n3539 = \state_reg[0]/NET0131  & ~n3538 ;
  assign n3540 = ~n3513 & ~n3539 ;
  assign n3541 = \reg3_reg[1]/NET0131  & ~n1426 ;
  assign n3542 = \reg3_reg[1]/NET0131  & n1388 ;
  assign n3544 = \reg3_reg[1]/NET0131  & ~n1169 ;
  assign n3553 = n1064 & n1218 ;
  assign n3554 = ~n1064 & ~n1218 ;
  assign n3555 = ~n3553 & ~n3554 ;
  assign n3562 = ~n771 & ~n3555 ;
  assign n3563 = n771 & n1064 ;
  assign n3564 = ~n3562 & ~n3563 ;
  assign n3565 = n1169 & n3564 ;
  assign n3566 = ~n3544 & ~n3565 ;
  assign n3567 = n1190 & ~n3566 ;
  assign n3545 = n735 & ~n1335 ;
  assign n3546 = ~n1336 & ~n3545 ;
  assign n3547 = ~n338 & ~n3546 ;
  assign n3548 = n338 & n768 ;
  assign n3549 = ~n3547 & ~n3548 ;
  assign n3550 = n1169 & n3549 ;
  assign n3551 = ~n3544 & ~n3550 ;
  assign n3552 = n1370 & ~n3551 ;
  assign n3556 = n1169 & ~n3555 ;
  assign n3557 = ~n3544 & ~n3556 ;
  assign n3558 = n1292 & ~n3557 ;
  assign n3568 = ~n759 & ~n771 ;
  assign n3569 = ~n1294 & ~n3568 ;
  assign n3570 = n1169 & n3569 ;
  assign n3571 = ~n3544 & ~n3570 ;
  assign n3572 = n1326 & ~n3571 ;
  assign n3559 = ~n759 & n1169 ;
  assign n3560 = ~n3544 & ~n3559 ;
  assign n3561 = n1328 & ~n3560 ;
  assign n3543 = \reg3_reg[1]/NET0131  & n1373 ;
  assign n3573 = ~n759 & n1331 ;
  assign n3574 = ~n3543 & ~n3573 ;
  assign n3575 = ~n3561 & n3574 ;
  assign n3576 = ~n3572 & n3575 ;
  assign n3577 = ~n3558 & n3576 ;
  assign n3578 = ~n3552 & n3577 ;
  assign n3579 = ~n3567 & n3578 ;
  assign n3580 = n1386 & ~n3579 ;
  assign n3581 = ~n3542 & ~n3580 ;
  assign n3582 = \state_reg[0]/NET0131  & ~n3581 ;
  assign n3583 = ~n3541 & ~n3582 ;
  assign n3584 = \reg3_reg[2]/NET0131  & ~n1426 ;
  assign n3585 = \reg3_reg[2]/NET0131  & n1388 ;
  assign n3590 = n718 & ~n1336 ;
  assign n3591 = ~n1337 & ~n3590 ;
  assign n3592 = ~n338 & ~n3591 ;
  assign n3593 = n338 & n752 ;
  assign n3594 = n1370 & ~n3593 ;
  assign n3595 = ~n3592 & n3594 ;
  assign n3587 = ~n1091 & ~n1221 ;
  assign n3586 = n1091 & n1221 ;
  assign n3588 = n1292 & ~n3586 ;
  assign n3589 = ~n3587 & n3588 ;
  assign n3597 = n967 & n1091 ;
  assign n3596 = ~n967 & ~n1091 ;
  assign n3598 = n1190 & ~n3596 ;
  assign n3599 = ~n3597 & n3598 ;
  assign n3600 = ~n3589 & ~n3599 ;
  assign n3601 = ~n3595 & n3600 ;
  assign n3602 = n1169 & ~n3601 ;
  assign n3603 = ~n742 & n1331 ;
  assign n3604 = \reg3_reg[2]/NET0131  & ~n1169 ;
  assign n3605 = ~n742 & ~n1294 ;
  assign n3606 = ~n1295 & ~n3605 ;
  assign n3607 = n1169 & n3606 ;
  assign n3608 = ~n3604 & ~n3607 ;
  assign n3609 = n1326 & ~n3608 ;
  assign n3616 = ~n3603 & ~n3609 ;
  assign n3610 = ~n1169 & ~n3231 ;
  assign n3611 = ~n1373 & ~n3610 ;
  assign n3612 = \reg3_reg[2]/NET0131  & ~n3611 ;
  assign n3613 = ~n742 & n1169 ;
  assign n3614 = ~n3604 & ~n3613 ;
  assign n3615 = n1328 & ~n3614 ;
  assign n3617 = ~n3612 & ~n3615 ;
  assign n3618 = n3616 & n3617 ;
  assign n3619 = ~n3602 & n3618 ;
  assign n3620 = n1386 & ~n3619 ;
  assign n3621 = ~n3585 & ~n3620 ;
  assign n3622 = \state_reg[0]/NET0131  & ~n3621 ;
  assign n3623 = ~n3584 & ~n3622 ;
  assign n3626 = n701 & n1388 ;
  assign n3628 = n701 & ~n1169 ;
  assign n3629 = n338 & ~n718 ;
  assign n3630 = n281 & ~n3046 ;
  assign n3631 = ~n338 & ~n1339 ;
  assign n3632 = ~n3630 & n3631 ;
  assign n3633 = ~n3629 & ~n3632 ;
  assign n3634 = n1169 & ~n3633 ;
  assign n3635 = ~n3628 & ~n3634 ;
  assign n3636 = n1370 & ~n3635 ;
  assign n3643 = ~n971 & n1031 ;
  assign n3644 = n971 & ~n1031 ;
  assign n3645 = ~n3643 & ~n3644 ;
  assign n3646 = n1169 & n3645 ;
  assign n3647 = ~n3628 & ~n3646 ;
  assign n3648 = n1190 & ~n3647 ;
  assign n3637 = n1031 & ~n1228 ;
  assign n3638 = ~n1031 & n1228 ;
  assign n3639 = ~n3637 & ~n3638 ;
  assign n3640 = n1169 & ~n3639 ;
  assign n3641 = ~n3628 & ~n3640 ;
  assign n3642 = n1292 & ~n3641 ;
  assign n3649 = ~n699 & ~n1296 ;
  assign n3650 = ~n1297 & ~n3649 ;
  assign n3651 = n1169 & n3650 ;
  assign n3652 = ~n3628 & ~n3651 ;
  assign n3653 = n1326 & ~n3652 ;
  assign n3627 = ~n699 & ~n1332 ;
  assign n3654 = n701 & ~n1375 ;
  assign n3655 = ~n3627 & ~n3654 ;
  assign n3656 = ~n3653 & n3655 ;
  assign n3657 = ~n3642 & n3656 ;
  assign n3658 = ~n3648 & n3657 ;
  assign n3659 = ~n3636 & n3658 ;
  assign n3660 = n1386 & ~n3659 ;
  assign n3661 = ~n3626 & ~n3660 ;
  assign n3662 = \state_reg[0]/NET0131  & ~n3661 ;
  assign n3624 = \reg3_reg[4]/NET0131  & ~\state_reg[0]/NET0131  ;
  assign n3625 = n311 & n701 ;
  assign n3663 = ~n3624 & ~n3625 ;
  assign n3664 = ~n3662 & n3663 ;
  assign n3667 = n656 & n1388 ;
  assign n3669 = n656 & ~n1169 ;
  assign n3670 = ~n975 & n1027 ;
  assign n3671 = n975 & ~n1027 ;
  assign n3672 = ~n3670 & ~n3671 ;
  assign n3673 = n1169 & n3672 ;
  assign n3674 = ~n3669 & ~n3673 ;
  assign n3675 = n1190 & ~n3674 ;
  assign n3690 = ~n652 & ~n1298 ;
  assign n3691 = ~n2369 & ~n3690 ;
  assign n3692 = n1169 & n3691 ;
  assign n3693 = ~n3669 & ~n3692 ;
  assign n3694 = n1326 & ~n3693 ;
  assign n3668 = ~n652 & ~n1332 ;
  assign n3695 = n656 & ~n1375 ;
  assign n3696 = ~n3668 & ~n3695 ;
  assign n3697 = ~n3694 & n3696 ;
  assign n3698 = ~n3675 & n3697 ;
  assign n3676 = ~n281 & n338 ;
  assign n3677 = n671 & ~n3070 ;
  assign n3678 = ~n338 & ~n1341 ;
  assign n3679 = ~n3677 & n3678 ;
  assign n3680 = ~n3676 & ~n3679 ;
  assign n3681 = n1169 & ~n3680 ;
  assign n3682 = ~n3669 & ~n3681 ;
  assign n3683 = n1370 & ~n3682 ;
  assign n3684 = n1027 & ~n2254 ;
  assign n3685 = ~n1027 & n2254 ;
  assign n3686 = ~n3684 & ~n3685 ;
  assign n3687 = n1169 & ~n3686 ;
  assign n3688 = ~n3669 & ~n3687 ;
  assign n3689 = n1292 & ~n3688 ;
  assign n3699 = ~n3683 & ~n3689 ;
  assign n3700 = n3698 & n3699 ;
  assign n3701 = n1386 & ~n3700 ;
  assign n3702 = ~n3667 & ~n3701 ;
  assign n3703 = \state_reg[0]/NET0131  & ~n3702 ;
  assign n3665 = \reg3_reg[6]/NET0131  & ~\state_reg[0]/NET0131  ;
  assign n3666 = n311 & n656 ;
  assign n3704 = ~n3665 & ~n3666 ;
  assign n3705 = ~n3703 & n3704 ;
  assign n3708 = n621 & n1388 ;
  assign n3710 = n621 & ~n1169 ;
  assign n3714 = n1169 & n3335 ;
  assign n3715 = ~n3710 & ~n3714 ;
  assign n3716 = n1370 & ~n3715 ;
  assign n3711 = n1169 & n3341 ;
  assign n3712 = ~n3710 & ~n3711 ;
  assign n3713 = n1190 & ~n3712 ;
  assign n3717 = n1169 & ~n3347 ;
  assign n3718 = ~n3710 & ~n3717 ;
  assign n3719 = n1292 & ~n3718 ;
  assign n3709 = n1169 & n3354 ;
  assign n3720 = n621 & ~n2345 ;
  assign n3721 = n635 & ~n1332 ;
  assign n3722 = ~n3720 & ~n3721 ;
  assign n3723 = ~n3709 & n3722 ;
  assign n3724 = ~n3719 & n3723 ;
  assign n3725 = ~n3713 & n3724 ;
  assign n3726 = ~n3716 & n3725 ;
  assign n3727 = n1386 & ~n3726 ;
  assign n3728 = ~n3708 & ~n3727 ;
  assign n3729 = \state_reg[0]/NET0131  & ~n3728 ;
  assign n3706 = \reg3_reg[8]/NET0131  & ~\state_reg[0]/NET0131  ;
  assign n3707 = n311 & n621 ;
  assign n3730 = ~n3706 & ~n3707 ;
  assign n3731 = ~n3729 & n3730 ;
  assign n3732 = \reg3_reg[10]/NET0131  & ~\state_reg[0]/NET0131  ;
  assign n3735 = n585 & ~n1169 ;
  assign n3736 = n581 & ~n3129 ;
  assign n3737 = ~n1345 & ~n3736 ;
  assign n3738 = ~n338 & ~n3737 ;
  assign n3739 = n338 & n618 ;
  assign n3740 = ~n3738 & ~n3739 ;
  assign n3741 = n1169 & n3740 ;
  assign n3742 = ~n3735 & ~n3741 ;
  assign n3743 = n1370 & ~n3742 ;
  assign n3744 = n1056 & n2270 ;
  assign n3745 = ~n1056 & ~n2270 ;
  assign n3746 = ~n3744 & ~n3745 ;
  assign n3747 = n1169 & n3746 ;
  assign n3748 = ~n3735 & ~n3747 ;
  assign n3749 = n1190 & ~n3748 ;
  assign n3750 = n1056 & n2259 ;
  assign n3751 = ~n1056 & ~n2259 ;
  assign n3752 = ~n3750 & ~n3751 ;
  assign n3753 = n1169 & ~n3752 ;
  assign n3754 = ~n3735 & ~n3753 ;
  assign n3755 = n1292 & ~n3754 ;
  assign n3756 = n601 & ~n1302 ;
  assign n3757 = n1326 & ~n1914 ;
  assign n3758 = ~n3756 & n3757 ;
  assign n3759 = n1169 & n3758 ;
  assign n3760 = n601 & ~n1332 ;
  assign n3734 = n585 & ~n2345 ;
  assign n3761 = n1386 & ~n3734 ;
  assign n3762 = ~n3760 & n3761 ;
  assign n3763 = ~n3759 & n3762 ;
  assign n3764 = ~n3755 & n3763 ;
  assign n3765 = ~n3749 & n3764 ;
  assign n3766 = ~n3743 & n3765 ;
  assign n3733 = ~n585 & ~n1386 ;
  assign n3767 = \state_reg[0]/NET0131  & ~n3733 ;
  assign n3768 = ~n3766 & n3767 ;
  assign n3769 = ~n3732 & ~n3768 ;
  assign n3770 = \reg3_reg[18]/NET0131  & ~\state_reg[0]/NET0131  ;
  assign n3773 = n823 & ~n1169 ;
  assign n3774 = n1090 & n2473 ;
  assign n3775 = ~n1090 & ~n2473 ;
  assign n3776 = ~n3774 & ~n3775 ;
  assign n3777 = n1169 & n3776 ;
  assign n3778 = ~n3773 & ~n3777 ;
  assign n3779 = n1190 & ~n3778 ;
  assign n3786 = n806 & ~n2989 ;
  assign n3787 = ~n1353 & ~n3786 ;
  assign n3788 = ~n338 & ~n3787 ;
  assign n3789 = n338 & n862 ;
  assign n3790 = ~n3788 & ~n3789 ;
  assign n3791 = n1169 & n3790 ;
  assign n3792 = ~n3773 & ~n3791 ;
  assign n3793 = n1370 & ~n3792 ;
  assign n3780 = n1090 & n3147 ;
  assign n3781 = ~n1090 & ~n3147 ;
  assign n3782 = ~n3780 & ~n3781 ;
  assign n3783 = n1169 & ~n3782 ;
  assign n3784 = ~n3773 & ~n3783 ;
  assign n3785 = n1292 & ~n3784 ;
  assign n3794 = n817 & ~n1310 ;
  assign n3795 = n1326 & ~n2410 ;
  assign n3796 = ~n3794 & n3795 ;
  assign n3797 = n1169 & n3796 ;
  assign n3798 = n817 & ~n1332 ;
  assign n3772 = n823 & ~n2345 ;
  assign n3799 = n1386 & ~n3772 ;
  assign n3800 = ~n3798 & n3799 ;
  assign n3801 = ~n3797 & n3800 ;
  assign n3802 = ~n3785 & n3801 ;
  assign n3803 = ~n3793 & n3802 ;
  assign n3804 = ~n3779 & n3803 ;
  assign n3771 = ~n823 & ~n1386 ;
  assign n3805 = \state_reg[0]/NET0131  & ~n3771 ;
  assign n3806 = ~n3804 & n3805 ;
  assign n3807 = ~n3770 & ~n3806 ;
  assign n3810 = n836 & n1388 ;
  assign n3812 = n836 & ~n1169 ;
  assign n3813 = n486 & ~n2439 ;
  assign n3814 = ~n3167 & ~n3813 ;
  assign n3815 = ~n338 & ~n3814 ;
  assign n3816 = n338 & n851 ;
  assign n3817 = ~n3815 & ~n3816 ;
  assign n3818 = n1169 & n3817 ;
  assign n3819 = ~n3812 & ~n3818 ;
  assign n3820 = n1370 & ~n3819 ;
  assign n3827 = n1047 & n1502 ;
  assign n3828 = ~n1047 & ~n1502 ;
  assign n3829 = ~n3827 & ~n3828 ;
  assign n3830 = n1169 & ~n3829 ;
  assign n3831 = ~n3812 & ~n3830 ;
  assign n3832 = n1292 & ~n3831 ;
  assign n3821 = n1047 & ~n1572 ;
  assign n3822 = ~n1047 & n1572 ;
  assign n3823 = ~n3821 & ~n3822 ;
  assign n3824 = n1169 & ~n3823 ;
  assign n3825 = ~n3812 & ~n3824 ;
  assign n3826 = n1190 & ~n3825 ;
  assign n3833 = n830 & ~n1313 ;
  assign n3834 = ~n2003 & ~n3833 ;
  assign n3835 = n1169 & n3834 ;
  assign n3836 = ~n3812 & ~n3835 ;
  assign n3837 = n1326 & ~n3836 ;
  assign n3811 = n830 & ~n1332 ;
  assign n3838 = n836 & ~n1375 ;
  assign n3839 = ~n3811 & ~n3838 ;
  assign n3840 = ~n3837 & n3839 ;
  assign n3841 = ~n3826 & n3840 ;
  assign n3842 = ~n3832 & n3841 ;
  assign n3843 = ~n3820 & n3842 ;
  assign n3844 = n1386 & ~n3843 ;
  assign n3845 = ~n3810 & ~n3844 ;
  assign n3846 = \state_reg[0]/NET0131  & ~n3845 ;
  assign n3808 = \reg3_reg[21]/NET0131  & ~\state_reg[0]/NET0131  ;
  assign n3809 = n311 & n836 ;
  assign n3847 = ~n3808 & ~n3809 ;
  assign n3848 = ~n3846 & n3847 ;
  assign n3849 = \reg2_reg[5]/NET0131  & ~n1426 ;
  assign n3850 = \reg2_reg[5]/NET0131  & n1388 ;
  assign n3853 = \reg2_reg[5]/NET0131  & ~n1396 ;
  assign n3854 = n1396 & n3075 ;
  assign n3855 = ~n3853 & ~n3854 ;
  assign n3856 = n1370 & ~n3855 ;
  assign n3860 = n1396 & ~n3088 ;
  assign n3861 = ~n3853 & ~n3860 ;
  assign n3862 = n1292 & ~n3861 ;
  assign n3857 = n1396 & n3081 ;
  assign n3858 = ~n3853 & ~n3857 ;
  assign n3859 = n1190 & ~n3858 ;
  assign n3863 = n1396 & n3093 ;
  assign n3864 = ~n3853 & ~n3863 ;
  assign n3865 = n1326 & ~n3864 ;
  assign n3867 = \reg2_reg[5]/NET0131  & ~n1414 ;
  assign n3851 = n690 & n1328 ;
  assign n3852 = n1396 & n3851 ;
  assign n3866 = n275 & n1331 ;
  assign n3868 = ~n3852 & ~n3866 ;
  assign n3869 = ~n3867 & n3868 ;
  assign n3870 = ~n3865 & n3869 ;
  assign n3871 = ~n3859 & n3870 ;
  assign n3872 = ~n3862 & n3871 ;
  assign n3873 = ~n3856 & n3872 ;
  assign n3874 = n1386 & ~n3873 ;
  assign n3875 = ~n3850 & ~n3874 ;
  assign n3876 = \state_reg[0]/NET0131  & ~n3875 ;
  assign n3877 = ~n3849 & ~n3876 ;
  assign n3878 = \reg0_reg[17]/NET0131  & ~n1426 ;
  assign n3879 = \reg0_reg[17]/NET0131  & n1388 ;
  assign n3880 = \reg0_reg[17]/NET0131  & ~n1607 ;
  assign n3881 = n1607 & n2993 ;
  assign n3882 = ~n3880 & ~n3881 ;
  assign n3883 = n1370 & ~n3882 ;
  assign n3884 = \reg0_reg[17]/NET0131  & ~n1623 ;
  assign n3888 = n871 & n1328 ;
  assign n3889 = n1326 & n3014 ;
  assign n3890 = ~n3888 & ~n3889 ;
  assign n3891 = n1607 & ~n3890 ;
  assign n3895 = ~n3884 & ~n3891 ;
  assign n3896 = ~n3883 & n3895 ;
  assign n3885 = n1607 & ~n3001 ;
  assign n3886 = ~n3880 & ~n3885 ;
  assign n3887 = n1190 & ~n3886 ;
  assign n3892 = n1607 & n3009 ;
  assign n3893 = ~n3880 & ~n3892 ;
  assign n3894 = n1292 & ~n3893 ;
  assign n3897 = ~n3887 & ~n3894 ;
  assign n3898 = n3896 & n3897 ;
  assign n3899 = n1386 & ~n3898 ;
  assign n3900 = ~n3879 & ~n3899 ;
  assign n3901 = \state_reg[0]/NET0131  & ~n3900 ;
  assign n3902 = ~n3878 & ~n3901 ;
  assign n3903 = \reg0_reg[1]/NET0131  & ~n1426 ;
  assign n3904 = \reg0_reg[1]/NET0131  & n1388 ;
  assign n3906 = \reg0_reg[1]/NET0131  & ~n1607 ;
  assign n3916 = n1607 & n3564 ;
  assign n3917 = ~n3906 & ~n3916 ;
  assign n3918 = n1190 & ~n3917 ;
  assign n3907 = n1607 & n3549 ;
  assign n3908 = ~n3906 & ~n3907 ;
  assign n3909 = n1370 & ~n3908 ;
  assign n3910 = n1607 & ~n3555 ;
  assign n3911 = ~n3906 & ~n3910 ;
  assign n3912 = n1292 & ~n3911 ;
  assign n3919 = ~n759 & n1607 ;
  assign n3920 = ~n3906 & ~n3919 ;
  assign n3921 = n1328 & ~n3920 ;
  assign n3905 = \reg0_reg[1]/NET0131  & ~n1620 ;
  assign n3913 = n1607 & n3569 ;
  assign n3914 = ~n3906 & ~n3913 ;
  assign n3915 = n1326 & ~n3914 ;
  assign n3922 = ~n3905 & ~n3915 ;
  assign n3923 = ~n3921 & n3922 ;
  assign n3924 = ~n3912 & n3923 ;
  assign n3925 = ~n3909 & n3924 ;
  assign n3926 = ~n3918 & n3925 ;
  assign n3927 = n1386 & ~n3926 ;
  assign n3928 = ~n3904 & ~n3927 ;
  assign n3929 = \state_reg[0]/NET0131  & ~n3928 ;
  assign n3930 = ~n3903 & ~n3929 ;
  assign n3940 = \reg0_reg[21]/NET0131  & ~n1607 ;
  assign n3941 = n2621 & n3817 ;
  assign n3942 = ~n3940 & ~n3941 ;
  assign n3943 = n1370 & ~n3942 ;
  assign n3931 = \reg0_reg[21]/NET0131  & ~n2616 ;
  assign n3933 = n1190 & ~n3823 ;
  assign n3932 = n1292 & ~n3829 ;
  assign n3934 = n830 & n1328 ;
  assign n3935 = n1326 & n3834 ;
  assign n3936 = ~n3934 & ~n3935 ;
  assign n3937 = ~n3932 & n3936 ;
  assign n3938 = ~n3933 & n3937 ;
  assign n3939 = n2621 & ~n3938 ;
  assign n3944 = ~n3931 & ~n3939 ;
  assign n3945 = ~n3943 & n3944 ;
  assign n3946 = \reg0_reg[22]/NET0131  & ~n1426 ;
  assign n3947 = \reg0_reg[22]/NET0131  & n1388 ;
  assign n3948 = \reg0_reg[22]/NET0131  & ~n1607 ;
  assign n3949 = n1607 & ~n3152 ;
  assign n3950 = ~n3948 & ~n3949 ;
  assign n3951 = n1292 & ~n3950 ;
  assign n3952 = n1607 & n3163 ;
  assign n3953 = ~n3948 & ~n3952 ;
  assign n3954 = n1190 & ~n3953 ;
  assign n3955 = n1370 & n3172 ;
  assign n3956 = n476 & n1328 ;
  assign n3957 = ~n3179 & ~n3956 ;
  assign n3958 = ~n3955 & n3957 ;
  assign n3959 = n1607 & ~n3958 ;
  assign n3960 = \reg0_reg[22]/NET0131  & ~n1624 ;
  assign n3961 = ~n3959 & ~n3960 ;
  assign n3962 = ~n3954 & n3961 ;
  assign n3963 = ~n3951 & n3962 ;
  assign n3964 = n1386 & ~n3963 ;
  assign n3965 = ~n3947 & ~n3964 ;
  assign n3966 = \state_reg[0]/NET0131  & ~n3965 ;
  assign n3967 = ~n3946 & ~n3966 ;
  assign n3968 = n3234 & ~n3595 ;
  assign n3969 = \reg0_reg[2]/NET0131  & ~n3968 ;
  assign n3970 = n1326 & n3606 ;
  assign n3971 = ~n742 & n1328 ;
  assign n3972 = ~n3970 & ~n3971 ;
  assign n3973 = n3601 & n3972 ;
  assign n3974 = n2621 & ~n3973 ;
  assign n3975 = ~n3969 & ~n3974 ;
  assign n3976 = ~n725 & n1328 ;
  assign n3977 = n3044 & ~n3976 ;
  assign n3978 = n2621 & ~n3977 ;
  assign n3979 = \reg0_reg[3]/NET0131  & ~n2616 ;
  assign n3980 = ~n3978 & ~n3979 ;
  assign n3981 = \reg0_reg[5]/NET0131  & ~n1426 ;
  assign n3982 = \reg0_reg[5]/NET0131  & n1388 ;
  assign n3984 = \reg0_reg[5]/NET0131  & ~n1607 ;
  assign n3985 = n1607 & n3075 ;
  assign n3986 = ~n3984 & ~n3985 ;
  assign n3987 = n1370 & ~n3986 ;
  assign n3991 = n1607 & ~n3088 ;
  assign n3992 = ~n3984 & ~n3991 ;
  assign n3993 = n1292 & ~n3992 ;
  assign n3988 = n1607 & n3081 ;
  assign n3989 = ~n3984 & ~n3988 ;
  assign n3990 = n1190 & ~n3989 ;
  assign n3994 = n1607 & n3093 ;
  assign n3995 = ~n3984 & ~n3994 ;
  assign n3996 = n1326 & ~n3995 ;
  assign n3983 = \reg0_reg[5]/NET0131  & ~n2142 ;
  assign n3997 = n1607 & n3851 ;
  assign n3998 = ~n3983 & ~n3997 ;
  assign n3999 = ~n3996 & n3998 ;
  assign n4000 = ~n3990 & n3999 ;
  assign n4001 = ~n3993 & n4000 ;
  assign n4002 = ~n3987 & n4001 ;
  assign n4003 = n1386 & ~n4002 ;
  assign n4004 = ~n3982 & ~n4003 ;
  assign n4005 = \state_reg[0]/NET0131  & ~n4004 ;
  assign n4006 = ~n3981 & ~n4005 ;
  assign n4007 = n1370 & n2968 ;
  assign n4008 = ~n530 & n1328 ;
  assign n4009 = ~n4007 & ~n4008 ;
  assign n4010 = n2958 & n4009 ;
  assign n4011 = n3369 & ~n4010 ;
  assign n4012 = n1635 & n2947 ;
  assign n4013 = n1326 & ~n4012 ;
  assign n4014 = n3420 & ~n4013 ;
  assign n4015 = \reg1_reg[13]/NET0131  & ~n4014 ;
  assign n4016 = ~n4011 & ~n4015 ;
  assign n4017 = \reg1_reg[17]/NET0131  & ~n1426 ;
  assign n4018 = \reg1_reg[17]/NET0131  & n1388 ;
  assign n4019 = \reg1_reg[17]/NET0131  & ~n1635 ;
  assign n4020 = n1635 & n2993 ;
  assign n4021 = ~n4019 & ~n4020 ;
  assign n4022 = n1370 & ~n4021 ;
  assign n4023 = \reg1_reg[17]/NET0131  & ~n1646 ;
  assign n4027 = n1635 & ~n3890 ;
  assign n4031 = ~n4023 & ~n4027 ;
  assign n4032 = ~n4022 & n4031 ;
  assign n4024 = n1635 & ~n3001 ;
  assign n4025 = ~n4019 & ~n4024 ;
  assign n4026 = n1190 & ~n4025 ;
  assign n4028 = n1635 & n3009 ;
  assign n4029 = ~n4019 & ~n4028 ;
  assign n4030 = n1292 & ~n4029 ;
  assign n4033 = ~n4026 & ~n4030 ;
  assign n4034 = n4032 & n4033 ;
  assign n4035 = n1386 & ~n4034 ;
  assign n4036 = ~n4018 & ~n4035 ;
  assign n4037 = \state_reg[0]/NET0131  & ~n4036 ;
  assign n4038 = ~n4017 & ~n4037 ;
  assign n4039 = \reg1_reg[1]/NET0131  & ~n1426 ;
  assign n4040 = \reg1_reg[1]/NET0131  & n1388 ;
  assign n4042 = \reg1_reg[1]/NET0131  & ~n1635 ;
  assign n4052 = n1635 & n3564 ;
  assign n4053 = ~n4042 & ~n4052 ;
  assign n4054 = n1190 & ~n4053 ;
  assign n4043 = n1635 & n3549 ;
  assign n4044 = ~n4042 & ~n4043 ;
  assign n4045 = n1370 & ~n4044 ;
  assign n4046 = n1635 & ~n3555 ;
  assign n4047 = ~n4042 & ~n4046 ;
  assign n4048 = n1292 & ~n4047 ;
  assign n4055 = ~n759 & n1635 ;
  assign n4056 = ~n4042 & ~n4055 ;
  assign n4057 = n1328 & ~n4056 ;
  assign n4041 = \reg1_reg[1]/NET0131  & ~n1620 ;
  assign n4049 = n1635 & n3569 ;
  assign n4050 = ~n4042 & ~n4049 ;
  assign n4051 = n1326 & ~n4050 ;
  assign n4058 = ~n4041 & ~n4051 ;
  assign n4059 = ~n4057 & n4058 ;
  assign n4060 = ~n4048 & n4059 ;
  assign n4061 = ~n4045 & n4060 ;
  assign n4062 = ~n4054 & n4061 ;
  assign n4063 = n1386 & ~n4062 ;
  assign n4064 = ~n4040 & ~n4063 ;
  assign n4065 = \state_reg[0]/NET0131  & ~n4064 ;
  assign n4066 = ~n4039 & ~n4065 ;
  assign n4067 = \reg1_reg[22]/NET0131  & ~n1426 ;
  assign n4068 = \reg1_reg[22]/NET0131  & n1388 ;
  assign n4069 = \reg1_reg[22]/NET0131  & ~n1635 ;
  assign n4070 = n1635 & ~n3152 ;
  assign n4071 = ~n4069 & ~n4070 ;
  assign n4072 = n1292 & ~n4071 ;
  assign n4073 = n1635 & n3163 ;
  assign n4074 = ~n4069 & ~n4073 ;
  assign n4075 = n1190 & ~n4074 ;
  assign n4076 = n1635 & ~n3958 ;
  assign n4077 = \reg1_reg[22]/NET0131  & ~n1647 ;
  assign n4078 = ~n4076 & ~n4077 ;
  assign n4079 = ~n4075 & n4078 ;
  assign n4080 = ~n4072 & n4079 ;
  assign n4081 = n1386 & ~n4080 ;
  assign n4082 = ~n4068 & ~n4081 ;
  assign n4083 = \state_reg[0]/NET0131  & ~n4082 ;
  assign n4084 = ~n4067 & ~n4083 ;
  assign n4085 = \reg1_reg[2]/NET0131  & ~n3367 ;
  assign n4086 = n3369 & ~n3973 ;
  assign n4087 = ~n4085 & ~n4086 ;
  assign n4088 = \reg0_reg[10]/NET0131  & ~n1426 ;
  assign n4089 = \reg0_reg[10]/NET0131  & n1388 ;
  assign n4091 = \reg0_reg[10]/NET0131  & ~n1607 ;
  assign n4092 = n1607 & n3740 ;
  assign n4093 = ~n4091 & ~n4092 ;
  assign n4094 = n1370 & ~n4093 ;
  assign n4095 = n1607 & n3746 ;
  assign n4096 = ~n4091 & ~n4095 ;
  assign n4097 = n1190 & ~n4096 ;
  assign n4090 = \reg0_reg[10]/NET0131  & ~n2613 ;
  assign n4099 = n1292 & ~n3752 ;
  assign n4098 = n601 & n1328 ;
  assign n4100 = ~n3758 & ~n4098 ;
  assign n4101 = ~n4099 & n4100 ;
  assign n4102 = n1607 & ~n4101 ;
  assign n4103 = ~n4090 & ~n4102 ;
  assign n4104 = ~n4097 & n4103 ;
  assign n4105 = ~n4094 & n4104 ;
  assign n4106 = n1386 & ~n4105 ;
  assign n4107 = ~n4089 & ~n4106 ;
  assign n4108 = \state_reg[0]/NET0131  & ~n4107 ;
  assign n4109 = ~n4088 & ~n4108 ;
  assign n4110 = \reg1_reg[3]/NET0131  & ~n3417 ;
  assign n4111 = n3369 & ~n3977 ;
  assign n4112 = ~n4110 & ~n4111 ;
  assign n4113 = \reg1_reg[5]/NET0131  & ~n1426 ;
  assign n4114 = \reg1_reg[5]/NET0131  & n1388 ;
  assign n4116 = \reg1_reg[5]/NET0131  & ~n1635 ;
  assign n4117 = n1635 & n3075 ;
  assign n4118 = ~n4116 & ~n4117 ;
  assign n4119 = n1370 & ~n4118 ;
  assign n4123 = n1635 & ~n3088 ;
  assign n4124 = ~n4116 & ~n4123 ;
  assign n4125 = n1292 & ~n4124 ;
  assign n4120 = n1635 & n3081 ;
  assign n4121 = ~n4116 & ~n4120 ;
  assign n4122 = n1190 & ~n4121 ;
  assign n4126 = n1635 & n3093 ;
  assign n4127 = ~n4116 & ~n4126 ;
  assign n4128 = n1326 & ~n4127 ;
  assign n4115 = \reg1_reg[5]/NET0131  & ~n2667 ;
  assign n4129 = n1635 & n3851 ;
  assign n4130 = ~n4115 & ~n4129 ;
  assign n4131 = ~n4128 & n4130 ;
  assign n4132 = ~n4122 & n4131 ;
  assign n4133 = ~n4125 & n4132 ;
  assign n4134 = ~n4119 & n4133 ;
  assign n4135 = n1386 & ~n4134 ;
  assign n4136 = ~n4114 & ~n4135 ;
  assign n4137 = \state_reg[0]/NET0131  & ~n4136 ;
  assign n4138 = ~n4113 & ~n4137 ;
  assign n4139 = n291 & n1331 ;
  assign n4140 = n1396 & ~n4010 ;
  assign n4141 = ~n4139 & ~n4140 ;
  assign n4142 = n1717 & ~n4141 ;
  assign n4143 = n325 & ~n1396 ;
  assign n4144 = n1717 & ~n4143 ;
  assign n4145 = n2208 & n4144 ;
  assign n4146 = \reg2_reg[13]/NET0131  & ~n4145 ;
  assign n4147 = ~n4142 & ~n4146 ;
  assign n4148 = \reg2_reg[17]/NET0131  & ~n1426 ;
  assign n4149 = \reg2_reg[17]/NET0131  & n1388 ;
  assign n4153 = \reg2_reg[17]/NET0131  & ~n1396 ;
  assign n4154 = n1396 & ~n3001 ;
  assign n4155 = ~n4153 & ~n4154 ;
  assign n4156 = n1190 & ~n4155 ;
  assign n4152 = n1396 & ~n3890 ;
  assign n4150 = n857 & n1331 ;
  assign n4151 = \reg2_reg[17]/NET0131  & ~n2208 ;
  assign n4163 = ~n4150 & ~n4151 ;
  assign n4164 = ~n4152 & n4163 ;
  assign n4165 = ~n4156 & n4164 ;
  assign n4157 = n1396 & n2993 ;
  assign n4158 = ~n4153 & ~n4157 ;
  assign n4159 = n1370 & ~n4158 ;
  assign n4160 = n1396 & n3009 ;
  assign n4161 = ~n4153 & ~n4160 ;
  assign n4162 = n1292 & ~n4161 ;
  assign n4166 = ~n4159 & ~n4162 ;
  assign n4167 = n4165 & n4166 ;
  assign n4168 = n1386 & ~n4167 ;
  assign n4169 = ~n4149 & ~n4168 ;
  assign n4170 = \state_reg[0]/NET0131  & ~n4169 ;
  assign n4171 = ~n4148 & ~n4170 ;
  assign n4172 = \reg2_reg[22]/NET0131  & ~n1426 ;
  assign n4173 = \reg2_reg[22]/NET0131  & n1388 ;
  assign n4174 = \reg2_reg[22]/NET0131  & ~n1396 ;
  assign n4175 = n1396 & ~n3152 ;
  assign n4176 = ~n4174 & ~n4175 ;
  assign n4177 = n1292 & ~n4176 ;
  assign n4178 = n1396 & n3163 ;
  assign n4179 = ~n4174 & ~n4178 ;
  assign n4180 = n1190 & ~n4179 ;
  assign n4181 = n1396 & ~n3958 ;
  assign n4182 = \reg2_reg[22]/NET0131  & ~n2209 ;
  assign n4183 = n482 & n1331 ;
  assign n4184 = ~n4182 & ~n4183 ;
  assign n4185 = ~n4181 & n4184 ;
  assign n4186 = ~n4180 & n4185 ;
  assign n4187 = ~n4177 & n4186 ;
  assign n4188 = n1386 & ~n4187 ;
  assign n4189 = ~n4173 & ~n4188 ;
  assign n4190 = \state_reg[0]/NET0131  & ~n4189 ;
  assign n4191 = ~n4172 & ~n4190 ;
  assign n4192 = n1396 & ~n3973 ;
  assign n4193 = \reg3_reg[2]/NET0131  & n1331 ;
  assign n4194 = ~n4192 & ~n4193 ;
  assign n4195 = n1717 & ~n4194 ;
  assign n4196 = n2574 & n3456 ;
  assign n4197 = \reg2_reg[2]/NET0131  & ~n4196 ;
  assign n4198 = ~n4195 & ~n4197 ;
  assign n4199 = n2621 & ~n4010 ;
  assign n4200 = ~n1607 & ~n2284 ;
  assign n4201 = n1717 & ~n4200 ;
  assign n4202 = n2142 & n4201 ;
  assign n4203 = \reg0_reg[13]/NET0131  & ~n4202 ;
  assign n4204 = ~n4199 & ~n4203 ;
  assign n4205 = \reg2_reg[4]/NET0131  & ~n1426 ;
  assign n4206 = \reg2_reg[4]/NET0131  & n1388 ;
  assign n4209 = \reg2_reg[4]/NET0131  & ~n1396 ;
  assign n4210 = n1396 & ~n3633 ;
  assign n4211 = ~n4209 & ~n4210 ;
  assign n4212 = n1370 & ~n4211 ;
  assign n4216 = n1396 & n3645 ;
  assign n4217 = ~n4209 & ~n4216 ;
  assign n4218 = n1190 & ~n4217 ;
  assign n4213 = n1396 & ~n3639 ;
  assign n4214 = ~n4209 & ~n4213 ;
  assign n4215 = n1292 & ~n4214 ;
  assign n4219 = n1396 & n3650 ;
  assign n4220 = ~n4209 & ~n4219 ;
  assign n4221 = n1326 & ~n4220 ;
  assign n4223 = \reg2_reg[4]/NET0131  & ~n1414 ;
  assign n4207 = ~n699 & n1328 ;
  assign n4208 = n1396 & n4207 ;
  assign n4222 = n701 & n1331 ;
  assign n4224 = ~n4208 & ~n4222 ;
  assign n4225 = ~n4223 & n4224 ;
  assign n4226 = ~n4221 & n4225 ;
  assign n4227 = ~n4215 & n4226 ;
  assign n4228 = ~n4218 & n4227 ;
  assign n4229 = ~n4212 & n4228 ;
  assign n4230 = n1386 & ~n4229 ;
  assign n4231 = ~n4206 & ~n4230 ;
  assign n4232 = \state_reg[0]/NET0131  & ~n4231 ;
  assign n4233 = ~n4205 & ~n4232 ;
  assign n4234 = \reg2_reg[6]/NET0131  & ~n1426 ;
  assign n4235 = \reg2_reg[6]/NET0131  & n1388 ;
  assign n4238 = \reg2_reg[6]/NET0131  & ~n1396 ;
  assign n4239 = n1396 & ~n3680 ;
  assign n4240 = ~n4238 & ~n4239 ;
  assign n4241 = n1370 & ~n4240 ;
  assign n4248 = n1396 & n3691 ;
  assign n4249 = ~n4238 & ~n4248 ;
  assign n4250 = n1326 & ~n4249 ;
  assign n4252 = \reg2_reg[6]/NET0131  & ~n1414 ;
  assign n4236 = ~n652 & n1328 ;
  assign n4237 = n1396 & n4236 ;
  assign n4251 = n656 & n1331 ;
  assign n4253 = ~n4237 & ~n4251 ;
  assign n4254 = ~n4252 & n4253 ;
  assign n4255 = ~n4250 & n4254 ;
  assign n4256 = ~n4241 & n4255 ;
  assign n4242 = n1396 & ~n3686 ;
  assign n4243 = ~n4238 & ~n4242 ;
  assign n4244 = n1292 & ~n4243 ;
  assign n4245 = n1396 & n3672 ;
  assign n4246 = ~n4238 & ~n4245 ;
  assign n4247 = n1190 & ~n4246 ;
  assign n4257 = ~n4244 & ~n4247 ;
  assign n4258 = n4256 & n4257 ;
  assign n4259 = n1386 & ~n4258 ;
  assign n4260 = ~n4235 & ~n4259 ;
  assign n4261 = \state_reg[0]/NET0131  & ~n4260 ;
  assign n4262 = ~n4234 & ~n4261 ;
  assign n4263 = \reg2_reg[8]/NET0131  & ~n1426 ;
  assign n4264 = \reg2_reg[8]/NET0131  & n1388 ;
  assign n4266 = \reg2_reg[8]/NET0131  & ~n1396 ;
  assign n4270 = n1396 & n3341 ;
  assign n4271 = ~n4266 & ~n4270 ;
  assign n4272 = n1190 & ~n4271 ;
  assign n4267 = n1396 & n3335 ;
  assign n4268 = ~n4266 & ~n4267 ;
  assign n4269 = n1370 & ~n4268 ;
  assign n4273 = n1396 & ~n3347 ;
  assign n4274 = ~n4266 & ~n4273 ;
  assign n4275 = n1292 & ~n4274 ;
  assign n4265 = n1396 & ~n3355 ;
  assign n4276 = n621 & n1331 ;
  assign n4277 = \reg2_reg[8]/NET0131  & ~n2208 ;
  assign n4278 = ~n4276 & ~n4277 ;
  assign n4279 = ~n4265 & n4278 ;
  assign n4280 = ~n4275 & n4279 ;
  assign n4281 = ~n4269 & n4280 ;
  assign n4282 = ~n4272 & n4281 ;
  assign n4283 = n1386 & ~n4282 ;
  assign n4284 = ~n4264 & ~n4283 ;
  assign n4285 = \state_reg[0]/NET0131  & ~n4284 ;
  assign n4286 = ~n4263 & ~n4285 ;
  assign n4287 = ~n609 & n1328 ;
  assign n4288 = n3121 & ~n4287 ;
  assign n4289 = ~n3125 & n4288 ;
  assign n4290 = n1396 & ~n4289 ;
  assign n4291 = n611 & n1331 ;
  assign n4292 = ~n4290 & ~n4291 ;
  assign n4293 = n1717 & ~n4292 ;
  assign n4294 = \reg2_reg[9]/NET0131  & ~n4196 ;
  assign n4295 = ~n4293 & ~n4294 ;
  assign n4296 = ~n2614 & n3295 ;
  assign n4297 = \reg0_reg[18]/NET0131  & ~n4296 ;
  assign n4298 = n1190 & n3776 ;
  assign n4300 = n1292 & ~n3782 ;
  assign n4299 = n1370 & n3790 ;
  assign n4301 = n817 & n1328 ;
  assign n4302 = ~n3796 & ~n4301 ;
  assign n4303 = ~n4299 & n4302 ;
  assign n4304 = ~n4300 & n4303 ;
  assign n4305 = ~n4298 & n4304 ;
  assign n4306 = n2621 & ~n4305 ;
  assign n4307 = ~n4297 & ~n4306 ;
  assign n4308 = \reg0_reg[4]/NET0131  & ~n1426 ;
  assign n4309 = \reg0_reg[4]/NET0131  & n1388 ;
  assign n4311 = \reg0_reg[4]/NET0131  & ~n1607 ;
  assign n4312 = n1607 & ~n3633 ;
  assign n4313 = ~n4311 & ~n4312 ;
  assign n4314 = n1370 & ~n4313 ;
  assign n4318 = n1607 & ~n3639 ;
  assign n4319 = ~n4311 & ~n4318 ;
  assign n4320 = n1292 & ~n4319 ;
  assign n4315 = n1607 & n3645 ;
  assign n4316 = ~n4311 & ~n4315 ;
  assign n4317 = n1190 & ~n4316 ;
  assign n4321 = n1607 & n3650 ;
  assign n4322 = ~n4311 & ~n4321 ;
  assign n4323 = n1326 & ~n4322 ;
  assign n4310 = \reg0_reg[4]/NET0131  & ~n2142 ;
  assign n4324 = n1607 & n4207 ;
  assign n4325 = ~n4310 & ~n4324 ;
  assign n4326 = ~n4323 & n4325 ;
  assign n4327 = ~n4317 & n4326 ;
  assign n4328 = ~n4320 & n4327 ;
  assign n4329 = ~n4314 & n4328 ;
  assign n4330 = n1386 & ~n4329 ;
  assign n4331 = ~n4309 & ~n4330 ;
  assign n4332 = \state_reg[0]/NET0131  & ~n4331 ;
  assign n4333 = ~n4308 & ~n4332 ;
  assign n4334 = \reg0_reg[6]/NET0131  & ~n1426 ;
  assign n4335 = \reg0_reg[6]/NET0131  & n1388 ;
  assign n4337 = \reg0_reg[6]/NET0131  & ~n1607 ;
  assign n4338 = n1607 & n3672 ;
  assign n4339 = ~n4337 & ~n4338 ;
  assign n4340 = n1190 & ~n4339 ;
  assign n4347 = n1607 & n3691 ;
  assign n4348 = ~n4337 & ~n4347 ;
  assign n4349 = n1326 & ~n4348 ;
  assign n4336 = \reg0_reg[6]/NET0131  & ~n2142 ;
  assign n4350 = n1607 & n4236 ;
  assign n4351 = ~n4336 & ~n4350 ;
  assign n4352 = ~n4349 & n4351 ;
  assign n4353 = ~n4340 & n4352 ;
  assign n4341 = n1607 & ~n3680 ;
  assign n4342 = ~n4337 & ~n4341 ;
  assign n4343 = n1370 & ~n4342 ;
  assign n4344 = n1607 & ~n3686 ;
  assign n4345 = ~n4337 & ~n4344 ;
  assign n4346 = n1292 & ~n4345 ;
  assign n4354 = ~n4343 & ~n4346 ;
  assign n4355 = n4353 & n4354 ;
  assign n4356 = n1386 & ~n4355 ;
  assign n4357 = ~n4335 & ~n4356 ;
  assign n4358 = \state_reg[0]/NET0131  & ~n4357 ;
  assign n4359 = ~n4334 & ~n4358 ;
  assign n4360 = n2621 & ~n4289 ;
  assign n4361 = \reg0_reg[9]/NET0131  & ~n2616 ;
  assign n4362 = ~n4360 & ~n4361 ;
  assign n4363 = \reg1_reg[10]/NET0131  & ~n1426 ;
  assign n4364 = \reg1_reg[10]/NET0131  & n1388 ;
  assign n4366 = \reg1_reg[10]/NET0131  & ~n1635 ;
  assign n4367 = n1635 & n3740 ;
  assign n4368 = ~n4366 & ~n4367 ;
  assign n4369 = n1370 & ~n4368 ;
  assign n4370 = n1635 & n3746 ;
  assign n4371 = ~n4366 & ~n4370 ;
  assign n4372 = n1190 & ~n4371 ;
  assign n4365 = \reg1_reg[10]/NET0131  & ~n3415 ;
  assign n4373 = n1635 & ~n4101 ;
  assign n4374 = ~n4365 & ~n4373 ;
  assign n4375 = ~n4372 & n4374 ;
  assign n4376 = ~n4369 & n4375 ;
  assign n4377 = n1386 & ~n4376 ;
  assign n4378 = ~n4364 & ~n4377 ;
  assign n4379 = \state_reg[0]/NET0131  & ~n4378 ;
  assign n4380 = ~n4363 & ~n4379 ;
  assign n4381 = \reg1_reg[18]/NET0131  & ~n1426 ;
  assign n4382 = \reg1_reg[18]/NET0131  & n1388 ;
  assign n4383 = n1635 & ~n4305 ;
  assign n4384 = \reg1_reg[18]/NET0131  & ~n2734 ;
  assign n4385 = ~n4383 & ~n4384 ;
  assign n4386 = n1386 & ~n4385 ;
  assign n4387 = ~n4382 & ~n4386 ;
  assign n4388 = \state_reg[0]/NET0131  & ~n4387 ;
  assign n4389 = ~n4381 & ~n4388 ;
  assign n4390 = n3369 & ~n3938 ;
  assign n4391 = \reg1_reg[21]/NET0131  & ~n3417 ;
  assign n4392 = ~n4390 & ~n4391 ;
  assign n4393 = \reg1_reg[4]/NET0131  & ~n1426 ;
  assign n4394 = \reg1_reg[4]/NET0131  & n1388 ;
  assign n4396 = \reg1_reg[4]/NET0131  & ~n1635 ;
  assign n4397 = n1635 & ~n3633 ;
  assign n4398 = ~n4396 & ~n4397 ;
  assign n4399 = n1370 & ~n4398 ;
  assign n4403 = n1635 & ~n3639 ;
  assign n4404 = ~n4396 & ~n4403 ;
  assign n4405 = n1292 & ~n4404 ;
  assign n4400 = n1635 & n3645 ;
  assign n4401 = ~n4396 & ~n4400 ;
  assign n4402 = n1190 & ~n4401 ;
  assign n4406 = n1635 & n3650 ;
  assign n4407 = ~n4396 & ~n4406 ;
  assign n4408 = n1326 & ~n4407 ;
  assign n4395 = \reg1_reg[4]/NET0131  & ~n2667 ;
  assign n4409 = n1635 & n4207 ;
  assign n4410 = ~n4395 & ~n4409 ;
  assign n4411 = ~n4408 & n4410 ;
  assign n4412 = ~n4402 & n4411 ;
  assign n4413 = ~n4405 & n4412 ;
  assign n4414 = ~n4399 & n4413 ;
  assign n4415 = n1386 & ~n4414 ;
  assign n4416 = ~n4394 & ~n4415 ;
  assign n4417 = \state_reg[0]/NET0131  & ~n4416 ;
  assign n4418 = ~n4393 & ~n4417 ;
  assign n4419 = \reg1_reg[6]/NET0131  & ~n1426 ;
  assign n4420 = \reg1_reg[6]/NET0131  & n1388 ;
  assign n4422 = \reg1_reg[6]/NET0131  & ~n1635 ;
  assign n4423 = n1635 & ~n3680 ;
  assign n4424 = ~n4422 & ~n4423 ;
  assign n4425 = n1370 & ~n4424 ;
  assign n4432 = n1635 & n3691 ;
  assign n4433 = ~n4422 & ~n4432 ;
  assign n4434 = n1326 & ~n4433 ;
  assign n4421 = \reg1_reg[6]/NET0131  & ~n2667 ;
  assign n4435 = n1635 & n4236 ;
  assign n4436 = ~n4421 & ~n4435 ;
  assign n4437 = ~n4434 & n4436 ;
  assign n4438 = ~n4425 & n4437 ;
  assign n4426 = n1635 & n3672 ;
  assign n4427 = ~n4422 & ~n4426 ;
  assign n4428 = n1190 & ~n4427 ;
  assign n4429 = n1635 & ~n3686 ;
  assign n4430 = ~n4422 & ~n4429 ;
  assign n4431 = n1292 & ~n4430 ;
  assign n4439 = ~n4428 & ~n4431 ;
  assign n4440 = n4438 & n4439 ;
  assign n4441 = n1386 & ~n4440 ;
  assign n4442 = ~n4420 & ~n4441 ;
  assign n4443 = \state_reg[0]/NET0131  & ~n4442 ;
  assign n4444 = ~n4419 & ~n4443 ;
  assign n4445 = \reg1_reg[8]/NET0131  & ~n1426 ;
  assign n4446 = \reg1_reg[8]/NET0131  & n1388 ;
  assign n4448 = \reg1_reg[8]/NET0131  & ~n1635 ;
  assign n4452 = n1635 & n3341 ;
  assign n4453 = ~n4448 & ~n4452 ;
  assign n4454 = n1190 & ~n4453 ;
  assign n4449 = n1635 & n3335 ;
  assign n4450 = ~n4448 & ~n4449 ;
  assign n4451 = n1370 & ~n4450 ;
  assign n4455 = n1635 & ~n3347 ;
  assign n4456 = ~n4448 & ~n4455 ;
  assign n4457 = n1292 & ~n4456 ;
  assign n4447 = \reg1_reg[8]/NET0131  & ~n1646 ;
  assign n4458 = n1635 & ~n3355 ;
  assign n4459 = ~n4447 & ~n4458 ;
  assign n4460 = ~n4457 & n4459 ;
  assign n4461 = ~n4451 & n4460 ;
  assign n4462 = ~n4454 & n4461 ;
  assign n4463 = n1386 & ~n4462 ;
  assign n4464 = ~n4446 & ~n4463 ;
  assign n4465 = \state_reg[0]/NET0131  & ~n4464 ;
  assign n4466 = ~n4445 & ~n4465 ;
  assign n4467 = \reg1_reg[9]/NET0131  & ~n3417 ;
  assign n4468 = n3369 & ~n4289 ;
  assign n4469 = ~n4467 & ~n4468 ;
  assign n4470 = \reg2_reg[10]/NET0131  & ~n1426 ;
  assign n4471 = \reg2_reg[10]/NET0131  & n1388 ;
  assign n4473 = \reg2_reg[10]/NET0131  & ~n1396 ;
  assign n4474 = n1396 & n3740 ;
  assign n4475 = ~n4473 & ~n4474 ;
  assign n4476 = n1370 & ~n4475 ;
  assign n4478 = n1396 & n3746 ;
  assign n4479 = ~n4473 & ~n4478 ;
  assign n4480 = n1190 & ~n4479 ;
  assign n4472 = n1396 & ~n4101 ;
  assign n4477 = n585 & n1331 ;
  assign n4481 = \reg2_reg[10]/NET0131  & ~n2574 ;
  assign n4482 = ~n4477 & ~n4481 ;
  assign n4483 = ~n4472 & n4482 ;
  assign n4484 = ~n4480 & n4483 ;
  assign n4485 = ~n4476 & n4484 ;
  assign n4486 = n1386 & ~n4485 ;
  assign n4487 = ~n4471 & ~n4486 ;
  assign n4488 = \state_reg[0]/NET0131  & ~n4487 ;
  assign n4489 = ~n4470 & ~n4488 ;
  assign n4490 = \reg2_reg[18]/NET0131  & ~n1426 ;
  assign n4491 = \reg2_reg[18]/NET0131  & n1388 ;
  assign n4492 = n1396 & ~n4304 ;
  assign n4496 = n1396 & ~n3776 ;
  assign n4495 = ~\reg2_reg[18]/NET0131  & ~n1396 ;
  assign n4497 = n1190 & ~n4495 ;
  assign n4498 = ~n4496 & n4497 ;
  assign n4493 = n823 & n1331 ;
  assign n4494 = \reg2_reg[18]/NET0131  & ~n2575 ;
  assign n4499 = ~n4493 & ~n4494 ;
  assign n4500 = ~n4498 & n4499 ;
  assign n4501 = ~n4492 & n4500 ;
  assign n4502 = n1386 & ~n4501 ;
  assign n4503 = ~n4491 & ~n4502 ;
  assign n4504 = \state_reg[0]/NET0131  & ~n4503 ;
  assign n4505 = ~n4490 & ~n4504 ;
  assign n4506 = \reg2_reg[1]/NET0131  & ~n1426 ;
  assign n4507 = \reg2_reg[1]/NET0131  & n1388 ;
  assign n4509 = \reg2_reg[1]/NET0131  & ~n1396 ;
  assign n4519 = n1396 & n3564 ;
  assign n4520 = ~n4509 & ~n4519 ;
  assign n4521 = n1190 & ~n4520 ;
  assign n4510 = n1396 & n3549 ;
  assign n4511 = ~n4509 & ~n4510 ;
  assign n4512 = n1370 & ~n4511 ;
  assign n4513 = n1396 & ~n3555 ;
  assign n4514 = ~n4509 & ~n4513 ;
  assign n4515 = n1292 & ~n4514 ;
  assign n4522 = n1396 & n3569 ;
  assign n4523 = ~n4509 & ~n4522 ;
  assign n4524 = n1326 & ~n4523 ;
  assign n4516 = ~n759 & n1396 ;
  assign n4517 = ~n4509 & ~n4516 ;
  assign n4518 = n1328 & ~n4517 ;
  assign n4508 = \reg3_reg[1]/NET0131  & n1331 ;
  assign n4525 = \reg2_reg[1]/NET0131  & n1373 ;
  assign n4526 = ~n4508 & ~n4525 ;
  assign n4527 = ~n4518 & n4526 ;
  assign n4528 = ~n4524 & n4527 ;
  assign n4529 = ~n4515 & n4528 ;
  assign n4530 = ~n4512 & n4529 ;
  assign n4531 = ~n4521 & n4530 ;
  assign n4532 = n1386 & ~n4531 ;
  assign n4533 = ~n4507 & ~n4532 ;
  assign n4534 = \state_reg[0]/NET0131  & ~n4533 ;
  assign n4535 = ~n4506 & ~n4534 ;
  assign n4536 = \reg2_reg[21]/NET0131  & ~n1426 ;
  assign n4537 = \reg2_reg[21]/NET0131  & n1388 ;
  assign n4539 = \reg2_reg[21]/NET0131  & ~n1396 ;
  assign n4540 = n1396 & n3817 ;
  assign n4541 = ~n4539 & ~n4540 ;
  assign n4542 = n1370 & ~n4541 ;
  assign n4546 = n1396 & ~n3829 ;
  assign n4547 = ~n4539 & ~n4546 ;
  assign n4548 = n1292 & ~n4547 ;
  assign n4543 = n1396 & ~n3823 ;
  assign n4544 = ~n4539 & ~n4543 ;
  assign n4545 = n1190 & ~n4544 ;
  assign n4549 = n1396 & ~n3936 ;
  assign n4538 = n836 & n1331 ;
  assign n4550 = \reg2_reg[21]/NET0131  & ~n2208 ;
  assign n4551 = ~n4538 & ~n4550 ;
  assign n4552 = ~n4549 & n4551 ;
  assign n4553 = ~n4545 & n4552 ;
  assign n4554 = ~n4548 & n4553 ;
  assign n4555 = ~n4542 & n4554 ;
  assign n4556 = n1386 & ~n4555 ;
  assign n4557 = ~n4537 & ~n4556 ;
  assign n4558 = \state_reg[0]/NET0131  & ~n4557 ;
  assign n4559 = ~n4536 & ~n4558 ;
  assign n4560 = \reg1_reg[0]/NET0131  & ~n1426 ;
  assign n4561 = \reg1_reg[0]/NET0131  & n1388 ;
  assign n4563 = \reg1_reg[0]/NET0131  & ~n1635 ;
  assign n4570 = n752 & ~n1334 ;
  assign n4571 = ~n338 & ~n1335 ;
  assign n4572 = ~n4570 & n4571 ;
  assign n4573 = n1635 & n4572 ;
  assign n4574 = ~n4563 & ~n4573 ;
  assign n4575 = n1370 & ~n4574 ;
  assign n4567 = ~n1032 & n1635 ;
  assign n4568 = ~n4563 & ~n4567 ;
  assign n4569 = ~n2732 & ~n4568 ;
  assign n4562 = \reg1_reg[0]/NET0131  & ~n1620 ;
  assign n4564 = ~n771 & n1635 ;
  assign n4565 = ~n4563 & ~n4564 ;
  assign n4566 = ~n1621 & ~n4565 ;
  assign n4576 = ~n4562 & ~n4566 ;
  assign n4577 = ~n4569 & n4576 ;
  assign n4578 = ~n4575 & n4577 ;
  assign n4579 = n1386 & ~n4578 ;
  assign n4580 = ~n4561 & ~n4579 ;
  assign n4581 = \state_reg[0]/NET0131  & ~n4580 ;
  assign n4582 = ~n4560 & ~n4581 ;
  assign n4583 = \reg2_reg[0]/NET0131  & ~n1426 ;
  assign n4584 = \reg2_reg[0]/NET0131  & n1388 ;
  assign n4586 = \reg2_reg[0]/NET0131  & ~n1396 ;
  assign n4593 = n1396 & n4572 ;
  assign n4594 = ~n4586 & ~n4593 ;
  assign n4595 = n1370 & ~n4594 ;
  assign n4590 = ~n1032 & n1396 ;
  assign n4591 = ~n4586 & ~n4590 ;
  assign n4592 = ~n2732 & ~n4591 ;
  assign n4587 = ~n771 & n1396 ;
  assign n4588 = ~n4586 & ~n4587 ;
  assign n4589 = ~n1621 & ~n4588 ;
  assign n4585 = \reg3_reg[0]/NET0131  & n1331 ;
  assign n4596 = \reg2_reg[0]/NET0131  & n1373 ;
  assign n4597 = ~n4585 & ~n4596 ;
  assign n4598 = ~n4589 & n4597 ;
  assign n4599 = ~n4592 & n4598 ;
  assign n4600 = ~n4595 & n4599 ;
  assign n4601 = n1386 & ~n4600 ;
  assign n4602 = ~n4584 & ~n4601 ;
  assign n4603 = \state_reg[0]/NET0131  & ~n4602 ;
  assign n4604 = ~n4583 & ~n4603 ;
  assign n4605 = \reg0_reg[0]/NET0131  & ~n1426 ;
  assign n4606 = \reg0_reg[0]/NET0131  & n1388 ;
  assign n4608 = \reg0_reg[0]/NET0131  & ~n1607 ;
  assign n4615 = n1607 & n4572 ;
  assign n4616 = ~n4608 & ~n4615 ;
  assign n4617 = n1370 & ~n4616 ;
  assign n4612 = ~n771 & n1607 ;
  assign n4613 = ~n4608 & ~n4612 ;
  assign n4614 = ~n1621 & ~n4613 ;
  assign n4607 = \reg0_reg[0]/NET0131  & ~n1620 ;
  assign n4609 = ~n1032 & n1607 ;
  assign n4610 = ~n4608 & ~n4609 ;
  assign n4611 = ~n2732 & ~n4610 ;
  assign n4618 = ~n4607 & ~n4611 ;
  assign n4619 = ~n4614 & n4618 ;
  assign n4620 = ~n4617 & n4619 ;
  assign n4621 = n1386 & ~n4620 ;
  assign n4622 = ~n4606 & ~n4621 ;
  assign n4623 = \state_reg[0]/NET0131  & ~n4622 ;
  assign n4624 = ~n4605 & ~n4623 ;
  assign n4681 = \reg2_reg[11]/NET0131  & ~n570 ;
  assign n4682 = ~\reg2_reg[11]/NET0131  & n570 ;
  assign n4683 = ~n4681 & ~n4682 ;
  assign n4684 = ~\reg2_reg[7]/NET0131  & ~n676 ;
  assign n4685 = \reg2_reg[6]/NET0131  & ~n650 ;
  assign n4686 = ~\reg2_reg[6]/NET0131  & n650 ;
  assign n4687 = \reg2_reg[5]/NET0131  & n687 ;
  assign n4688 = ~\reg2_reg[5]/NET0131  & ~n687 ;
  assign n4689 = \reg2_reg[4]/NET0131  & ~n697 ;
  assign n4690 = ~\reg2_reg[4]/NET0131  & n697 ;
  assign n4691 = \reg2_reg[3]/NET0131  & n722 ;
  assign n4692 = ~\reg2_reg[3]/NET0131  & ~n722 ;
  assign n4693 = \reg2_reg[2]/NET0131  & ~n740 ;
  assign n4694 = ~\reg2_reg[2]/NET0131  & n740 ;
  assign n4695 = \reg2_reg[1]/NET0131  & ~n756 ;
  assign n4696 = ~\reg2_reg[1]/NET0131  & n756 ;
  assign n4697 = \IR_reg[0]/NET0131  & \reg2_reg[0]/NET0131  ;
  assign n4698 = ~n4696 & n4697 ;
  assign n4699 = ~n4695 & ~n4698 ;
  assign n4700 = ~n4694 & ~n4699 ;
  assign n4701 = ~n4693 & ~n4700 ;
  assign n4702 = ~n4692 & ~n4701 ;
  assign n4703 = ~n4691 & ~n4702 ;
  assign n4704 = ~n4690 & ~n4703 ;
  assign n4705 = ~n4689 & ~n4704 ;
  assign n4706 = ~n4688 & ~n4705 ;
  assign n4707 = ~n4687 & ~n4706 ;
  assign n4708 = ~n4686 & ~n4707 ;
  assign n4709 = ~n4685 & ~n4708 ;
  assign n4710 = ~n4684 & ~n4709 ;
  assign n4711 = \reg2_reg[7]/NET0131  & n676 ;
  assign n4712 = \reg2_reg[8]/NET0131  & n632 ;
  assign n4713 = ~n4711 & ~n4712 ;
  assign n4714 = ~n4710 & n4713 ;
  assign n4715 = ~\reg2_reg[9]/NET0131  & n607 ;
  assign n4716 = ~\reg2_reg[8]/NET0131  & ~n632 ;
  assign n4717 = ~n4715 & ~n4716 ;
  assign n4718 = ~n4714 & n4717 ;
  assign n4719 = \reg2_reg[9]/NET0131  & ~n607 ;
  assign n4720 = \reg2_reg[10]/NET0131  & n598 ;
  assign n4721 = ~n4719 & ~n4720 ;
  assign n4722 = ~n4718 & n4721 ;
  assign n4723 = ~\reg2_reg[10]/NET0131  & ~n598 ;
  assign n4724 = ~n4722 & ~n4723 ;
  assign n4726 = n4683 & n4724 ;
  assign n4680 = n332 & n338 ;
  assign n4725 = ~n4683 & ~n4724 ;
  assign n4727 = n4680 & ~n4725 ;
  assign n4728 = ~n4726 & n4727 ;
  assign n4666 = \reg1_reg[11]/NET0131  & ~n570 ;
  assign n4625 = ~\reg1_reg[10]/NET0131  & ~n598 ;
  assign n4626 = \reg1_reg[6]/NET0131  & ~n650 ;
  assign n4627 = \reg1_reg[5]/NET0131  & n687 ;
  assign n4628 = ~\reg1_reg[5]/NET0131  & ~n687 ;
  assign n4629 = \reg1_reg[4]/NET0131  & ~n697 ;
  assign n4630 = ~\reg1_reg[4]/NET0131  & n697 ;
  assign n4631 = \reg1_reg[3]/NET0131  & n722 ;
  assign n4632 = ~\reg1_reg[3]/NET0131  & ~n722 ;
  assign n4633 = \reg1_reg[2]/NET0131  & ~n740 ;
  assign n4634 = ~\reg1_reg[2]/NET0131  & n740 ;
  assign n4635 = \reg1_reg[1]/NET0131  & ~n756 ;
  assign n4636 = ~\reg1_reg[1]/NET0131  & n756 ;
  assign n4637 = \IR_reg[0]/NET0131  & \reg1_reg[0]/NET0131  ;
  assign n4638 = ~n4636 & n4637 ;
  assign n4639 = ~n4635 & ~n4638 ;
  assign n4640 = ~n4634 & ~n4639 ;
  assign n4641 = ~n4633 & ~n4640 ;
  assign n4642 = ~n4632 & ~n4641 ;
  assign n4643 = ~n4631 & ~n4642 ;
  assign n4644 = ~n4630 & ~n4643 ;
  assign n4645 = ~n4629 & ~n4644 ;
  assign n4646 = ~n4628 & ~n4645 ;
  assign n4647 = ~n4627 & ~n4646 ;
  assign n4648 = ~n4626 & n4647 ;
  assign n4649 = ~\reg1_reg[7]/NET0131  & ~n676 ;
  assign n4650 = ~\reg1_reg[6]/NET0131  & n650 ;
  assign n4651 = ~n4649 & ~n4650 ;
  assign n4652 = ~n4648 & n4651 ;
  assign n4653 = \reg1_reg[8]/NET0131  & n632 ;
  assign n4654 = \reg1_reg[7]/NET0131  & n676 ;
  assign n4655 = ~n4653 & ~n4654 ;
  assign n4656 = ~n4652 & n4655 ;
  assign n4657 = ~\reg1_reg[9]/NET0131  & n607 ;
  assign n4658 = ~\reg1_reg[8]/NET0131  & ~n632 ;
  assign n4659 = ~n4657 & ~n4658 ;
  assign n4660 = ~n4656 & n4659 ;
  assign n4661 = \reg1_reg[9]/NET0131  & ~n607 ;
  assign n4662 = \reg1_reg[10]/NET0131  & n598 ;
  assign n4663 = ~n4661 & ~n4662 ;
  assign n4664 = ~n4660 & n4663 ;
  assign n4665 = ~n4625 & ~n4664 ;
  assign n4667 = ~\reg1_reg[11]/NET0131  & n570 ;
  assign n4671 = n4665 & ~n4667 ;
  assign n4672 = ~n4666 & n4671 ;
  assign n4668 = ~n4666 & ~n4667 ;
  assign n4669 = ~n4665 & ~n4668 ;
  assign n4670 = ~n332 & n338 ;
  assign n4673 = ~n4669 & n4670 ;
  assign n4674 = ~n4672 & n4673 ;
  assign n4675 = ~n332 & ~n1388 ;
  assign n4677 = n570 & ~n4675 ;
  assign n4676 = ~\addr[11]_pad  & n4675 ;
  assign n4678 = ~n338 & ~n4676 ;
  assign n4679 = ~n4677 & n4678 ;
  assign n4729 = ~n4674 & ~n4679 ;
  assign n4730 = ~n4728 & n4729 ;
  assign n4731 = \state_reg[0]/NET0131  & ~n4730 ;
  assign n4732 = ~n1888 & ~n4731 ;
  assign n4755 = \reg2_reg[12]/NET0131  & n548 ;
  assign n4756 = ~\reg2_reg[12]/NET0131  & ~n548 ;
  assign n4757 = ~n4755 & ~n4756 ;
  assign n4758 = ~n4710 & ~n4711 ;
  assign n4759 = ~n4716 & ~n4758 ;
  assign n4760 = ~n4712 & ~n4719 ;
  assign n4761 = ~n4759 & n4760 ;
  assign n4762 = ~n4715 & ~n4761 ;
  assign n4763 = ~n4723 & n4762 ;
  assign n4764 = ~n4681 & ~n4720 ;
  assign n4765 = ~n4763 & n4764 ;
  assign n4766 = ~n4682 & ~n4765 ;
  assign n4768 = n4757 & n4766 ;
  assign n4767 = ~n4757 & ~n4766 ;
  assign n4769 = n4680 & ~n4767 ;
  assign n4770 = ~n4768 & n4769 ;
  assign n4733 = \reg1_reg[12]/NET0131  & n548 ;
  assign n4734 = ~\reg1_reg[12]/NET0131  & ~n548 ;
  assign n4735 = ~n4733 & ~n4734 ;
  assign n4736 = ~n4648 & ~n4650 ;
  assign n4737 = ~n4654 & ~n4736 ;
  assign n4738 = ~n4649 & ~n4737 ;
  assign n4739 = ~n4658 & n4738 ;
  assign n4740 = ~n4653 & ~n4661 ;
  assign n4741 = ~n4739 & n4740 ;
  assign n4742 = ~n4657 & ~n4741 ;
  assign n4743 = ~n4625 & n4742 ;
  assign n4744 = ~n4662 & ~n4666 ;
  assign n4745 = ~n4743 & n4744 ;
  assign n4746 = ~n4667 & ~n4745 ;
  assign n4748 = n4735 & n4746 ;
  assign n4747 = ~n4735 & ~n4746 ;
  assign n4749 = n4670 & ~n4747 ;
  assign n4750 = ~n4748 & n4749 ;
  assign n4752 = ~\addr[12]_pad  & n4675 ;
  assign n4751 = ~n548 & ~n4675 ;
  assign n4753 = ~n338 & ~n4751 ;
  assign n4754 = ~n4752 & n4753 ;
  assign n4771 = ~n4750 & ~n4754 ;
  assign n4772 = ~n4770 & n4771 ;
  assign n4773 = \state_reg[0]/NET0131  & ~n4772 ;
  assign n4774 = ~n1932 & ~n4773 ;
  assign n4799 = \reg1_reg[15]/NET0131  & n519 ;
  assign n4802 = ~\reg1_reg[13]/NET0131  & ~n527 ;
  assign n4803 = ~n4734 & ~n4802 ;
  assign n4804 = ~n4666 & ~n4733 ;
  assign n4805 = ~n4671 & n4804 ;
  assign n4806 = n4803 & ~n4805 ;
  assign n4807 = \reg1_reg[13]/NET0131  & n527 ;
  assign n4808 = \reg1_reg[14]/NET0131  & n501 ;
  assign n4809 = ~n4807 & ~n4808 ;
  assign n4810 = ~n4806 & n4809 ;
  assign n4800 = ~\reg1_reg[15]/NET0131  & ~n519 ;
  assign n4811 = ~\reg1_reg[14]/NET0131  & ~n501 ;
  assign n4814 = ~n4800 & ~n4811 ;
  assign n4815 = ~n4810 & n4814 ;
  assign n4816 = ~n4799 & n4815 ;
  assign n4801 = ~n4799 & ~n4800 ;
  assign n4812 = ~n4810 & ~n4811 ;
  assign n4813 = ~n4801 & ~n4812 ;
  assign n4817 = n4670 & ~n4813 ;
  assign n4818 = ~n4816 & n4817 ;
  assign n4775 = ~\reg2_reg[15]/NET0131  & ~n519 ;
  assign n4776 = \reg2_reg[15]/NET0131  & n519 ;
  assign n4777 = ~n4775 & ~n4776 ;
  assign n4778 = ~\reg2_reg[14]/NET0131  & ~n501 ;
  assign n4779 = ~\reg2_reg[13]/NET0131  & ~n527 ;
  assign n4780 = ~n4756 & ~n4779 ;
  assign n4781 = ~n4682 & ~n4723 ;
  assign n4782 = ~n4722 & n4781 ;
  assign n4783 = ~n4681 & ~n4755 ;
  assign n4784 = ~n4782 & n4783 ;
  assign n4785 = n4780 & ~n4784 ;
  assign n4786 = \reg2_reg[14]/NET0131  & n501 ;
  assign n4787 = \reg2_reg[13]/NET0131  & n527 ;
  assign n4788 = ~n4786 & ~n4787 ;
  assign n4789 = ~n4785 & n4788 ;
  assign n4790 = ~n4778 & ~n4789 ;
  assign n4792 = ~n4777 & ~n4790 ;
  assign n4791 = n4777 & n4790 ;
  assign n4793 = n4680 & ~n4791 ;
  assign n4794 = ~n4792 & n4793 ;
  assign n4796 = ~\addr[15]_pad  & n4675 ;
  assign n4795 = ~n519 & ~n4675 ;
  assign n4797 = ~n338 & ~n4795 ;
  assign n4798 = ~n4796 & n4797 ;
  assign n4819 = ~n4794 & ~n4798 ;
  assign n4820 = ~n4818 & n4819 ;
  assign n4821 = \state_reg[0]/NET0131  & ~n4820 ;
  assign n4822 = ~n1719 & ~n4821 ;
  assign n4839 = ~\reg2_reg[17]/NET0131  & ~n868 ;
  assign n4840 = \reg2_reg[17]/NET0131  & n868 ;
  assign n4841 = ~n4839 & ~n4840 ;
  assign n4842 = \reg2_reg[16]/NET0131  & n875 ;
  assign n4843 = ~n4776 & ~n4790 ;
  assign n4844 = ~\reg2_reg[16]/NET0131  & ~n875 ;
  assign n4845 = ~n4775 & ~n4844 ;
  assign n4846 = ~n4843 & n4845 ;
  assign n4847 = ~n4842 & ~n4846 ;
  assign n4849 = n4841 & ~n4847 ;
  assign n4848 = ~n4841 & n4847 ;
  assign n4850 = n4680 & ~n4848 ;
  assign n4851 = ~n4849 & n4850 ;
  assign n4823 = ~\reg1_reg[17]/NET0131  & ~n868 ;
  assign n4824 = \reg1_reg[17]/NET0131  & n868 ;
  assign n4825 = ~n4823 & ~n4824 ;
  assign n4826 = ~\reg1_reg[16]/NET0131  & ~n875 ;
  assign n4827 = \reg1_reg[16]/NET0131  & n875 ;
  assign n4828 = ~n4799 & ~n4827 ;
  assign n4829 = ~n4815 & n4828 ;
  assign n4830 = ~n4826 & ~n4829 ;
  assign n4832 = n4825 & n4830 ;
  assign n4831 = ~n4825 & ~n4830 ;
  assign n4833 = n4670 & ~n4831 ;
  assign n4834 = ~n4832 & n4833 ;
  assign n4836 = ~\addr[17]_pad  & n4675 ;
  assign n4835 = ~n868 & ~n4675 ;
  assign n4837 = ~n338 & ~n4835 ;
  assign n4838 = ~n4836 & n4837 ;
  assign n4852 = ~n4834 & ~n4838 ;
  assign n4853 = ~n4851 & n4852 ;
  assign n4854 = \state_reg[0]/NET0131  & ~n4853 ;
  assign n4855 = ~n2982 & ~n4854 ;
  assign n4867 = ~\addr[5]_pad  & n4675 ;
  assign n4866 = ~n687 & ~n4675 ;
  assign n4868 = ~n338 & ~n4866 ;
  assign n4869 = ~n4867 & n4868 ;
  assign n4856 = ~n4687 & ~n4688 ;
  assign n4858 = ~n4705 & n4856 ;
  assign n4857 = n4705 & ~n4856 ;
  assign n4859 = n4680 & ~n4857 ;
  assign n4860 = ~n4858 & n4859 ;
  assign n4861 = ~n4627 & ~n4628 ;
  assign n4863 = ~n4645 & n4861 ;
  assign n4862 = n4645 & ~n4861 ;
  assign n4864 = n4670 & ~n4862 ;
  assign n4865 = ~n4863 & n4864 ;
  assign n4870 = ~n4860 & ~n4865 ;
  assign n4871 = ~n4869 & n4870 ;
  assign n4872 = \state_reg[0]/NET0131  & ~n4871 ;
  assign n4873 = ~n3065 & ~n4872 ;
  assign n4883 = ~n4685 & ~n4686 ;
  assign n4885 = ~n4707 & n4883 ;
  assign n4884 = n4707 & ~n4883 ;
  assign n4886 = n4680 & ~n4884 ;
  assign n4887 = ~n4885 & n4886 ;
  assign n4874 = ~n4626 & ~n4650 ;
  assign n4876 = ~n4647 & n4874 ;
  assign n4875 = n4647 & ~n4874 ;
  assign n4877 = n4670 & ~n4875 ;
  assign n4878 = ~n4876 & n4877 ;
  assign n4880 = n650 & ~n4675 ;
  assign n4879 = ~\addr[6]_pad  & n4675 ;
  assign n4881 = ~n338 & ~n4879 ;
  assign n4882 = ~n4880 & n4881 ;
  assign n4888 = ~n4878 & ~n4882 ;
  assign n4889 = ~n4887 & n4888 ;
  assign n4890 = \state_reg[0]/NET0131  & ~n4889 ;
  assign n4891 = ~n3665 & ~n4890 ;
  assign n4901 = ~n4684 & ~n4711 ;
  assign n4903 = ~n4709 & n4901 ;
  assign n4902 = n4709 & ~n4901 ;
  assign n4904 = n4680 & ~n4902 ;
  assign n4905 = ~n4903 & n4904 ;
  assign n4892 = ~n4649 & ~n4654 ;
  assign n4894 = n4736 & n4892 ;
  assign n4893 = ~n4736 & ~n4892 ;
  assign n4895 = n4670 & ~n4893 ;
  assign n4896 = ~n4894 & n4895 ;
  assign n4898 = ~\addr[7]_pad  & n4675 ;
  assign n4897 = ~n676 & ~n4675 ;
  assign n4899 = ~n338 & ~n4897 ;
  assign n4900 = ~n4898 & n4899 ;
  assign n4906 = ~n4896 & ~n4900 ;
  assign n4907 = ~n4905 & n4906 ;
  assign n4908 = \state_reg[0]/NET0131  & ~n4907 ;
  assign n4909 = ~n2341 & ~n4908 ;
  assign n4919 = ~n4712 & ~n4716 ;
  assign n4921 = ~n4758 & n4919 ;
  assign n4920 = n4758 & ~n4919 ;
  assign n4922 = n4680 & ~n4920 ;
  assign n4923 = ~n4921 & n4922 ;
  assign n4911 = ~\addr[8]_pad  & n4675 ;
  assign n4910 = ~n632 & ~n4675 ;
  assign n4912 = ~n338 & ~n4910 ;
  assign n4913 = ~n4911 & n4912 ;
  assign n4914 = ~n4653 & ~n4658 ;
  assign n4916 = n4738 & n4914 ;
  assign n4915 = ~n4738 & ~n4914 ;
  assign n4917 = n4670 & ~n4915 ;
  assign n4918 = ~n4916 & n4917 ;
  assign n4924 = ~n4913 & ~n4918 ;
  assign n4925 = ~n4923 & n4924 ;
  assign n4926 = \state_reg[0]/NET0131  & ~n4925 ;
  assign n4927 = ~n3706 & ~n4926 ;
  assign n4939 = ~n4715 & ~n4719 ;
  assign n4940 = ~n4712 & ~n4939 ;
  assign n4941 = ~n4759 & n4940 ;
  assign n4938 = n4718 & ~n4719 ;
  assign n4942 = n4680 & ~n4938 ;
  assign n4943 = ~n4941 & n4942 ;
  assign n4931 = n4660 & ~n4661 ;
  assign n4928 = ~n4657 & ~n4661 ;
  assign n4929 = ~n4656 & ~n4658 ;
  assign n4930 = ~n4928 & ~n4929 ;
  assign n4932 = n4670 & ~n4930 ;
  assign n4933 = ~n4931 & n4932 ;
  assign n4935 = n607 & ~n4675 ;
  assign n4934 = ~\addr[9]_pad  & n4675 ;
  assign n4936 = ~n338 & ~n4934 ;
  assign n4937 = ~n4935 & n4936 ;
  assign n4944 = ~n4933 & ~n4937 ;
  assign n4945 = ~n4943 & n4944 ;
  assign n4946 = \state_reg[0]/NET0131  & ~n4945 ;
  assign n4947 = ~n3108 & ~n4946 ;
  assign n4961 = ~n4778 & ~n4786 ;
  assign n4962 = n4766 & n4780 ;
  assign n4963 = n4755 & ~n4779 ;
  assign n4964 = ~n4787 & ~n4963 ;
  assign n4965 = ~n4962 & n4964 ;
  assign n4967 = n4961 & ~n4965 ;
  assign n4966 = ~n4961 & n4965 ;
  assign n4968 = n4680 & ~n4966 ;
  assign n4969 = ~n4967 & n4968 ;
  assign n4948 = ~n4808 & ~n4811 ;
  assign n4949 = n4746 & n4803 ;
  assign n4950 = n4733 & ~n4802 ;
  assign n4951 = ~n4807 & ~n4950 ;
  assign n4952 = ~n4949 & n4951 ;
  assign n4954 = n4948 & ~n4952 ;
  assign n4953 = ~n4948 & n4952 ;
  assign n4955 = n4670 & ~n4953 ;
  assign n4956 = ~n4954 & n4955 ;
  assign n4958 = ~\addr[14]_pad  & n4675 ;
  assign n4957 = ~n501 & ~n4675 ;
  assign n4959 = ~n338 & ~n4957 ;
  assign n4960 = ~n4958 & n4959 ;
  assign n4970 = ~n4956 & ~n4960 ;
  assign n4971 = ~n4969 & n4970 ;
  assign n4972 = \state_reg[0]/NET0131  & ~n4971 ;
  assign n4973 = ~n2293 & ~n4972 ;
  assign n4983 = ~n4720 & ~n4723 ;
  assign n4985 = n4762 & n4983 ;
  assign n4984 = ~n4762 & ~n4983 ;
  assign n4986 = n4680 & ~n4984 ;
  assign n4987 = ~n4985 & n4986 ;
  assign n4975 = ~\addr[10]_pad  & n4675 ;
  assign n4974 = ~n598 & ~n4675 ;
  assign n4976 = ~n338 & ~n4974 ;
  assign n4977 = ~n4975 & n4976 ;
  assign n4978 = ~n4625 & ~n4662 ;
  assign n4980 = n4742 & n4978 ;
  assign n4979 = ~n4742 & ~n4978 ;
  assign n4981 = n4670 & ~n4979 ;
  assign n4982 = ~n4980 & n4981 ;
  assign n4988 = ~n4977 & ~n4982 ;
  assign n4989 = ~n4987 & n4988 ;
  assign n4990 = \state_reg[0]/NET0131  & ~n4989 ;
  assign n4991 = ~n3732 & ~n4990 ;
  assign n5005 = n4806 & ~n4807 ;
  assign n5002 = ~n4802 & ~n4807 ;
  assign n5003 = ~n4734 & ~n4805 ;
  assign n5004 = ~n5002 & ~n5003 ;
  assign n5006 = n4670 & ~n5004 ;
  assign n5007 = ~n5005 & n5006 ;
  assign n4995 = n4785 & ~n4787 ;
  assign n4992 = ~n4779 & ~n4787 ;
  assign n4993 = ~n4756 & ~n4784 ;
  assign n4994 = ~n4992 & ~n4993 ;
  assign n4996 = n4680 & ~n4994 ;
  assign n4997 = ~n4995 & n4996 ;
  assign n4999 = ~\addr[13]_pad  & n4675 ;
  assign n4998 = ~n527 & ~n4675 ;
  assign n5000 = ~n338 & ~n4998 ;
  assign n5001 = ~n4999 & n5000 ;
  assign n5008 = ~n4997 & ~n5001 ;
  assign n5009 = ~n5007 & n5008 ;
  assign n5010 = \state_reg[0]/NET0131  & ~n5009 ;
  assign n5011 = ~n2979 & ~n5010 ;
  assign n5031 = \reg2_reg[18]/NET0131  & n814 ;
  assign n5032 = ~\reg2_reg[18]/NET0131  & ~n814 ;
  assign n5033 = ~n5031 & ~n5032 ;
  assign n5034 = ~n4778 & ~n4965 ;
  assign n5035 = ~n4776 & ~n4786 ;
  assign n5036 = ~n5034 & n5035 ;
  assign n5037 = ~n4775 & ~n5036 ;
  assign n5038 = ~n4844 & n5037 ;
  assign n5039 = ~n4840 & ~n4842 ;
  assign n5040 = ~n5038 & n5039 ;
  assign n5041 = ~n4839 & ~n5040 ;
  assign n5043 = n5033 & n5041 ;
  assign n5042 = ~n5033 & ~n5041 ;
  assign n5044 = n4680 & ~n5042 ;
  assign n5045 = ~n5043 & n5044 ;
  assign n5012 = \reg1_reg[18]/NET0131  & n814 ;
  assign n5013 = ~\reg1_reg[18]/NET0131  & ~n814 ;
  assign n5014 = ~n5012 & ~n5013 ;
  assign n5015 = n4814 & ~n4952 ;
  assign n5016 = ~n4800 & n4808 ;
  assign n5017 = ~n4799 & ~n5016 ;
  assign n5018 = ~n5015 & n5017 ;
  assign n5019 = ~n4826 & ~n5018 ;
  assign n5020 = ~n4824 & ~n4827 ;
  assign n5021 = ~n5019 & n5020 ;
  assign n5022 = ~n4823 & ~n5021 ;
  assign n5024 = n5014 & n5022 ;
  assign n5023 = ~n5014 & ~n5022 ;
  assign n5025 = n4670 & ~n5023 ;
  assign n5026 = ~n5024 & n5025 ;
  assign n5028 = ~\addr[18]_pad  & n4675 ;
  assign n5027 = ~n814 & ~n4675 ;
  assign n5029 = ~n338 & ~n5027 ;
  assign n5030 = ~n5028 & n5029 ;
  assign n5046 = ~n5026 & ~n5030 ;
  assign n5047 = ~n5045 & n5046 ;
  assign n5048 = \state_reg[0]/NET0131  & ~n5047 ;
  assign n5049 = ~n3770 & ~n5048 ;
  assign n5065 = ~n4824 & ~n4830 ;
  assign n5066 = ~n4823 & ~n5013 ;
  assign n5067 = ~n5065 & n5066 ;
  assign n5068 = ~n5012 & ~n5067 ;
  assign n5069 = \reg1_reg[19]/NET0131  & ~n5068 ;
  assign n5070 = ~\reg1_reg[19]/NET0131  & n5068 ;
  assign n5071 = ~n5069 & ~n5070 ;
  assign n5073 = ~n794 & ~n5071 ;
  assign n5072 = n794 & n5071 ;
  assign n5074 = n4670 & ~n5072 ;
  assign n5075 = ~n5073 & n5074 ;
  assign n5050 = ~n4840 & n4847 ;
  assign n5051 = ~n4839 & ~n5032 ;
  assign n5052 = ~n5050 & n5051 ;
  assign n5053 = ~n5031 & ~n5052 ;
  assign n5054 = ~\reg2_reg[19]/NET0131  & ~n794 ;
  assign n5055 = \reg2_reg[19]/NET0131  & n794 ;
  assign n5056 = ~n5054 & ~n5055 ;
  assign n5058 = ~n5053 & n5056 ;
  assign n5057 = n5053 & ~n5056 ;
  assign n5059 = n4680 & ~n5057 ;
  assign n5060 = ~n5058 & n5059 ;
  assign n5062 = ~\addr[19]_pad  & n4675 ;
  assign n5061 = ~n794 & ~n4675 ;
  assign n5063 = ~n338 & ~n5061 ;
  assign n5064 = ~n5062 & n5063 ;
  assign n5076 = ~n5060 & ~n5064 ;
  assign n5077 = ~n5075 & n5076 ;
  assign n5078 = \state_reg[0]/NET0131  & ~n5077 ;
  assign n5079 = ~n2385 & ~n5078 ;
  assign n5089 = ~n4842 & ~n4844 ;
  assign n5091 = n5037 & n5089 ;
  assign n5090 = ~n5037 & ~n5089 ;
  assign n5092 = n4680 & ~n5090 ;
  assign n5093 = ~n5091 & n5092 ;
  assign n5081 = ~\addr[16]_pad  & n4675 ;
  assign n5080 = ~n875 & ~n4675 ;
  assign n5082 = ~n338 & ~n5080 ;
  assign n5083 = ~n5081 & n5082 ;
  assign n5084 = ~n4826 & ~n4827 ;
  assign n5086 = ~n5018 & n5084 ;
  assign n5085 = n5018 & ~n5084 ;
  assign n5087 = n4670 & ~n5085 ;
  assign n5088 = ~n5086 & n5087 ;
  assign n5094 = ~n5083 & ~n5088 ;
  assign n5095 = ~n5093 & n5094 ;
  assign n5096 = \state_reg[0]/NET0131  & ~n5095 ;
  assign n5097 = ~n2297 & ~n5096 ;
  assign n5098 = \reg3_reg[1]/NET0131  & ~\state_reg[0]/NET0131  ;
  assign n5102 = n756 & n1388 ;
  assign n5101 = ~\addr[1]_pad  & ~n1388 ;
  assign n5103 = n339 & ~n5101 ;
  assign n5104 = ~n5102 & n5103 ;
  assign n5110 = ~n4695 & ~n4696 ;
  assign n5111 = ~n4697 & ~n5110 ;
  assign n5112 = n4697 & n5110 ;
  assign n5113 = ~n5111 & ~n5112 ;
  assign n5114 = n4680 & n5113 ;
  assign n5099 = n332 & ~n338 ;
  assign n5100 = ~n756 & n5099 ;
  assign n5105 = ~n4635 & ~n4636 ;
  assign n5106 = n4637 & n5105 ;
  assign n5107 = ~n4637 & ~n5105 ;
  assign n5108 = ~n5106 & ~n5107 ;
  assign n5109 = n4670 & n5108 ;
  assign n5115 = ~n5100 & ~n5109 ;
  assign n5116 = ~n5114 & n5115 ;
  assign n5117 = ~n5104 & n5116 ;
  assign n5118 = \state_reg[0]/NET0131  & ~n5117 ;
  assign n5119 = ~n5098 & ~n5118 ;
  assign n5120 = \reg3_reg[2]/NET0131  & ~\state_reg[0]/NET0131  ;
  assign n5123 = n740 & n1388 ;
  assign n5122 = ~\addr[2]_pad  & ~n1388 ;
  assign n5124 = n339 & ~n5122 ;
  assign n5125 = ~n5123 & n5124 ;
  assign n5131 = ~n4633 & ~n4634 ;
  assign n5132 = n4639 & ~n5131 ;
  assign n5133 = ~n4639 & n5131 ;
  assign n5134 = ~n5132 & ~n5133 ;
  assign n5135 = n4670 & n5134 ;
  assign n5121 = ~n740 & n5099 ;
  assign n5126 = ~n4693 & ~n4694 ;
  assign n5127 = ~n4699 & n5126 ;
  assign n5128 = n4699 & ~n5126 ;
  assign n5129 = ~n5127 & ~n5128 ;
  assign n5130 = n4680 & n5129 ;
  assign n5136 = ~n5121 & ~n5130 ;
  assign n5137 = ~n5135 & n5136 ;
  assign n5138 = ~n5125 & n5137 ;
  assign n5139 = \state_reg[0]/NET0131  & ~n5138 ;
  assign n5140 = ~n5120 & ~n5139 ;
  assign n5143 = ~n722 & n1388 ;
  assign n5142 = ~\addr[3]_pad  & ~n1388 ;
  assign n5144 = n339 & ~n5142 ;
  assign n5145 = ~n5143 & n5144 ;
  assign n5151 = ~n4691 & ~n4692 ;
  assign n5152 = n4701 & ~n5151 ;
  assign n5153 = ~n4701 & n5151 ;
  assign n5154 = ~n5152 & ~n5153 ;
  assign n5155 = n4680 & n5154 ;
  assign n5141 = n722 & n5099 ;
  assign n5146 = ~n4631 & ~n4632 ;
  assign n5147 = ~n4641 & n5146 ;
  assign n5148 = n4641 & ~n5146 ;
  assign n5149 = ~n5147 & ~n5148 ;
  assign n5150 = n4670 & n5149 ;
  assign n5156 = ~n5141 & ~n5150 ;
  assign n5157 = ~n5155 & n5156 ;
  assign n5158 = ~n5145 & n5157 ;
  assign n5159 = \state_reg[0]/NET0131  & ~n5158 ;
  assign n5160 = ~n3028 & ~n5159 ;
  assign n5163 = n697 & n1388 ;
  assign n5162 = ~\addr[4]_pad  & ~n1388 ;
  assign n5164 = n339 & ~n5162 ;
  assign n5165 = ~n5163 & n5164 ;
  assign n5171 = ~n4689 & ~n4690 ;
  assign n5173 = ~n4703 & n5171 ;
  assign n5172 = n4703 & ~n5171 ;
  assign n5174 = n4680 & ~n5172 ;
  assign n5175 = ~n5173 & n5174 ;
  assign n5161 = ~n697 & n5099 ;
  assign n5166 = ~n4629 & ~n4630 ;
  assign n5168 = ~n4643 & n5166 ;
  assign n5167 = n4643 & ~n5166 ;
  assign n5169 = n4670 & ~n5167 ;
  assign n5170 = ~n5168 & n5169 ;
  assign n5176 = ~n5161 & ~n5170 ;
  assign n5177 = ~n5175 & n5176 ;
  assign n5178 = ~n5165 & n5177 ;
  assign n5179 = \state_reg[0]/NET0131  & ~n5178 ;
  assign n5180 = ~n3624 & ~n5179 ;
  assign n5181 = \reg3_reg[0]/NET0131  & ~\state_reg[0]/NET0131  ;
  assign n5184 = ~\IR_reg[0]/NET0131  & n1388 ;
  assign n5183 = ~\addr[0]_pad  & ~n1388 ;
  assign n5185 = n339 & ~n5183 ;
  assign n5186 = ~n5184 & n5185 ;
  assign n5190 = ~\IR_reg[0]/NET0131  & ~\reg2_reg[0]/NET0131  ;
  assign n5191 = ~n4697 & ~n5190 ;
  assign n5192 = n4680 & n5191 ;
  assign n5182 = \IR_reg[0]/NET0131  & n5099 ;
  assign n5187 = ~\IR_reg[0]/NET0131  & ~\reg1_reg[0]/NET0131  ;
  assign n5188 = ~n4637 & ~n5187 ;
  assign n5189 = n4670 & n5188 ;
  assign n5193 = ~n5182 & ~n5189 ;
  assign n5194 = ~n5192 & n5193 ;
  assign n5195 = ~n5186 & n5194 ;
  assign n5196 = \state_reg[0]/NET0131  & ~n5195 ;
  assign n5197 = ~n5181 & ~n5196 ;
  assign n5198 = ~n339 & ~n1388 ;
  assign n5199 = \state_reg[0]/NET0131  & ~n5198 ;
  assign n5200 = \state_reg[0]/NET0131  & n1388 ;
  assign n5201 = \state_reg[0]/NET0131  & n332 ;
  assign n5202 = \datai[27]_pad  & ~\state_reg[0]/NET0131  ;
  assign n5203 = ~n5201 & ~n5202 ;
  assign n5204 = \state_reg[0]/NET0131  & n247 ;
  assign n5205 = \datai[30]_pad  & ~\state_reg[0]/NET0131  ;
  assign n5206 = ~n5204 & ~n5205 ;
  assign n5207 = \datai[31]_pad  & ~\state_reg[0]/NET0131  ;
  assign n5208 = ~\IR_reg[30]/NET0131  & \IR_reg[31]/NET0131  ;
  assign n5209 = \state_reg[0]/NET0131  & n5208 ;
  assign n5210 = n240 & n5209 ;
  assign n5211 = n328 & n5210 ;
  assign n5212 = ~n5207 & ~n5211 ;
  assign n5213 = \state_reg[0]/NET0131  & n266 ;
  assign n5214 = \datai[29]_pad  & ~\state_reg[0]/NET0131  ;
  assign n5215 = ~n5213 & ~n5214 ;
  assign n5216 = \state_reg[0]/NET0131  & n338 ;
  assign n5217 = \datai[28]_pad  & ~\state_reg[0]/NET0131  ;
  assign n5218 = ~n5216 & ~n5217 ;
  assign n5219 = \state_reg[0]/NET0131  & n794 ;
  assign n5220 = \datai[19]_pad  & ~\state_reg[0]/NET0131  ;
  assign n5221 = ~n5219 & ~n5220 ;
  assign n5222 = \state_reg[0]/NET0131  & n325 ;
  assign n5223 = \datai[22]_pad  & ~\state_reg[0]/NET0131  ;
  assign n5224 = ~n5222 & ~n5223 ;
  assign n5225 = \state_reg[0]/NET0131  & n317 ;
  assign n5226 = \datai[21]_pad  & ~\state_reg[0]/NET0131  ;
  assign n5227 = ~n5225 & ~n5226 ;
  assign n5228 = \state_reg[0]/NET0131  & n868 ;
  assign n5229 = \datai[17]_pad  & ~\state_reg[0]/NET0131  ;
  assign n5230 = ~n5228 & ~n5229 ;
  assign n5231 = \datai[23]_pad  & ~\state_reg[0]/NET0131  ;
  assign n5232 = ~n311 & ~n5231 ;
  assign n5233 = \state_reg[0]/NET0131  & n1144 ;
  assign n5234 = \datai[24]_pad  & ~\state_reg[0]/NET0131  ;
  assign n5235 = ~n5233 & ~n5234 ;
  assign n5236 = \state_reg[0]/NET0131  & n519 ;
  assign n5237 = \datai[15]_pad  & ~\state_reg[0]/NET0131  ;
  assign n5238 = ~n5236 & ~n5237 ;
  assign n5239 = \datai[20]_pad  & ~\state_reg[0]/NET0131  ;
  assign n5240 = \state_reg[0]/NET0131  & ~n932 ;
  assign n5241 = ~n5239 & ~n5240 ;
  assign n5242 = \state_reg[0]/NET0131  & ~n570 ;
  assign n5243 = \datai[11]_pad  & ~\state_reg[0]/NET0131  ;
  assign n5244 = ~n5242 & ~n5243 ;
  assign n5245 = \state_reg[0]/NET0131  & n1157 ;
  assign n5246 = \datai[25]_pad  & ~\state_reg[0]/NET0131  ;
  assign n5247 = ~n5245 & ~n5246 ;
  assign n5248 = \state_reg[0]/NET0131  & n814 ;
  assign n5249 = \datai[18]_pad  & ~\state_reg[0]/NET0131  ;
  assign n5250 = ~n5248 & ~n5249 ;
  assign n5251 = \state_reg[0]/NET0131  & n1149 ;
  assign n5252 = \datai[26]_pad  & ~\state_reg[0]/NET0131  ;
  assign n5253 = ~n5251 & ~n5252 ;
  assign n5254 = \state_reg[0]/NET0131  & n501 ;
  assign n5255 = \datai[14]_pad  & ~\state_reg[0]/NET0131  ;
  assign n5256 = ~n5254 & ~n5255 ;
  assign n5257 = \state_reg[0]/NET0131  & ~n875 ;
  assign n5258 = ~\datai[16]_pad  & ~\state_reg[0]/NET0131  ;
  assign n5259 = ~n5257 & ~n5258 ;
  assign n5260 = \state_reg[0]/NET0131  & n527 ;
  assign n5261 = \datai[13]_pad  & ~\state_reg[0]/NET0131  ;
  assign n5262 = ~n5260 & ~n5261 ;
  assign n5263 = \state_reg[0]/NET0131  & n676 ;
  assign n5264 = \datai[7]_pad  & ~\state_reg[0]/NET0131  ;
  assign n5265 = ~n5263 & ~n5264 ;
  assign n5266 = \state_reg[0]/NET0131  & n548 ;
  assign n5267 = \datai[12]_pad  & ~\state_reg[0]/NET0131  ;
  assign n5268 = ~n5266 & ~n5267 ;
  assign n5269 = \state_reg[0]/NET0131  & ~n607 ;
  assign n5270 = \datai[9]_pad  & ~\state_reg[0]/NET0131  ;
  assign n5271 = ~n5269 & ~n5270 ;
  assign n5272 = \state_reg[0]/NET0131  & n598 ;
  assign n5273 = \datai[10]_pad  & ~\state_reg[0]/NET0131  ;
  assign n5274 = ~n5272 & ~n5273 ;
  assign n5275 = \state_reg[0]/NET0131  & n632 ;
  assign n5276 = \datai[8]_pad  & ~\state_reg[0]/NET0131  ;
  assign n5277 = ~n5275 & ~n5276 ;
  assign n5278 = \state_reg[0]/NET0131  & n687 ;
  assign n5279 = \datai[5]_pad  & ~\state_reg[0]/NET0131  ;
  assign n5280 = ~n5278 & ~n5279 ;
  assign n5281 = \datai[6]_pad  & ~\state_reg[0]/NET0131  ;
  assign n5282 = \state_reg[0]/NET0131  & ~n650 ;
  assign n5283 = ~n5281 & ~n5282 ;
  assign n5284 = \state_reg[0]/NET0131  & n722 ;
  assign n5285 = \datai[3]_pad  & ~\state_reg[0]/NET0131  ;
  assign n5286 = ~n5284 & ~n5285 ;
  assign n5287 = \state_reg[0]/NET0131  & ~n697 ;
  assign n5288 = \datai[4]_pad  & ~\state_reg[0]/NET0131  ;
  assign n5289 = ~n5287 & ~n5288 ;
  assign n5290 = \state_reg[0]/NET0131  & ~n756 ;
  assign n5291 = \datai[1]_pad  & ~\state_reg[0]/NET0131  ;
  assign n5292 = ~n5290 & ~n5291 ;
  assign n5293 = \datai[2]_pad  & ~\state_reg[0]/NET0131  ;
  assign n5294 = \state_reg[0]/NET0131  & ~n740 ;
  assign n5295 = ~n5293 & ~n5294 ;
  assign n5298 = n410 & ~n1169 ;
  assign n5299 = n1169 & ~n1743 ;
  assign n5300 = ~n5298 & ~n5299 ;
  assign n5301 = n1292 & ~n5300 ;
  assign n5302 = n1169 & ~n1767 ;
  assign n5303 = ~n5298 & ~n5302 ;
  assign n5304 = n1190 & ~n5303 ;
  assign n5305 = n1169 & n1777 ;
  assign n5306 = ~n5298 & ~n5305 ;
  assign n5307 = n1370 & ~n5306 ;
  assign n5308 = n1169 & n1811 ;
  assign n5297 = n410 & ~n2345 ;
  assign n5309 = n405 & ~n1332 ;
  assign n5310 = ~n5297 & ~n5309 ;
  assign n5311 = ~n5308 & n5310 ;
  assign n5312 = ~n5307 & n5311 ;
  assign n5313 = ~n5304 & n5312 ;
  assign n5314 = ~n5301 & n5313 ;
  assign n5315 = n1717 & ~n5314 ;
  assign n5296 = n410 & n1657 ;
  assign n5316 = \reg3_reg[27]/NET0131  & ~\state_reg[0]/NET0131  ;
  assign n5317 = ~n5296 & ~n5316 ;
  assign n5318 = ~n5315 & n5317 ;
  assign n5319 = \reg3_reg[0]/NET0131  & ~n1426 ;
  assign n5320 = \reg3_reg[0]/NET0131  & n1388 ;
  assign n5322 = \reg3_reg[0]/NET0131  & ~n1169 ;
  assign n5329 = n1169 & n4572 ;
  assign n5330 = ~n5322 & ~n5329 ;
  assign n5331 = n1370 & ~n5330 ;
  assign n5326 = ~n1032 & n1169 ;
  assign n5327 = ~n5322 & ~n5326 ;
  assign n5328 = ~n2732 & ~n5327 ;
  assign n5323 = ~n771 & n1169 ;
  assign n5324 = ~n5322 & ~n5323 ;
  assign n5325 = ~n1621 & ~n5324 ;
  assign n5321 = \reg3_reg[0]/NET0131  & n1373 ;
  assign n5332 = ~n771 & n1331 ;
  assign n5333 = ~n5321 & ~n5332 ;
  assign n5334 = ~n5325 & n5333 ;
  assign n5335 = ~n5328 & n5334 ;
  assign n5336 = ~n5331 & n5335 ;
  assign n5337 = n1386 & ~n5336 ;
  assign n5338 = ~n5320 & ~n5337 ;
  assign n5339 = \state_reg[0]/NET0131  & ~n5338 ;
  assign n5340 = ~n5319 & ~n5339 ;
  assign n5341 = ~\reg3_reg[3]/NET0131  & n1331 ;
  assign n5342 = ~n3051 & n3977 ;
  assign n5343 = n1396 & ~n5342 ;
  assign n5344 = ~n5341 & ~n5343 ;
  assign n5345 = n1717 & ~n5344 ;
  assign n5346 = ~n2206 & n4196 ;
  assign n5347 = \reg2_reg[3]/NET0131  & ~n5346 ;
  assign n5348 = ~n5345 & ~n5347 ;
  assign n5351 = n422 & ~n1169 ;
  assign n5352 = n1169 & ~n2748 ;
  assign n5353 = ~n5351 & ~n5352 ;
  assign n5354 = n1190 & ~n5353 ;
  assign n5355 = n1169 & ~n2767 ;
  assign n5356 = ~n5351 & ~n5355 ;
  assign n5357 = n1292 & ~n5356 ;
  assign n5358 = n1169 & n2754 ;
  assign n5359 = ~n5351 & ~n5358 ;
  assign n5360 = n1370 & ~n5359 ;
  assign n5361 = n1169 & n2771 ;
  assign n5350 = n422 & ~n2345 ;
  assign n5362 = n417 & ~n1332 ;
  assign n5363 = ~n5350 & ~n5362 ;
  assign n5364 = ~n5361 & n5363 ;
  assign n5365 = ~n5360 & n5364 ;
  assign n5366 = ~n5357 & n5365 ;
  assign n5367 = ~n5354 & n5366 ;
  assign n5368 = n1717 & ~n5367 ;
  assign n5349 = n422 & n1657 ;
  assign n5369 = \reg3_reg[25]/NET0131  & ~\state_reg[0]/NET0131  ;
  assign n5370 = ~n5349 & ~n5369 ;
  assign n5371 = ~n5368 & n5370 ;
  assign \_al_n0  = 1'b0 ;
  assign \_al_n1  = ~1'b0 ;
  assign \g29_dup/_0_  = ~n281 ;
  assign \g33_dup47063/_0_  = ~n298 ;
  assign \g36117/_0_  = ~n1139 ;
  assign \g36132/_0_  = ~n1395 ;
  assign \g36133/_0_  = ~n1428 ;
  assign \g36134/_0_  = ~n1605 ;
  assign \g36135/_0_  = ~n1633 ;
  assign \g36136/_0_  = ~n1656 ;
  assign \g36153/_0_  = ~n1721 ;
  assign \g36154/_0_  = ~n1801 ;
  assign \g36155/_0_  = ~n1823 ;
  assign \g36156/_0_  = ~n1847 ;
  assign \g36157/_0_  = ~n1865 ;
  assign \g36158/_0_  = ~n1887 ;
  assign \g36186/_0_  = ~n1931 ;
  assign \g36187/_0_  = ~n1974 ;
  assign \g36193/_0_  = ~n2034 ;
  assign \g36197/_0_  = ~n2083 ;
  assign \g36198/_0_  = ~n2106 ;
  assign \g36199/_0_  = ~n2129 ;
  assign \g36200/_0_  = ~n2158 ;
  assign \g36201/_0_  = ~n2176 ;
  assign \g36202/_0_  = ~n2194 ;
  assign \g36203/_0_  = ~n2218 ;
  assign \g36204/_0_  = ~n2238 ;
  assign \g36239/_0_  = ~n2295 ;
  assign \g36240/_0_  = ~n2340 ;
  assign \g36242/_0_  = ~n2384 ;
  assign \g36246/_0_  = ~n2426 ;
  assign \g36255/_0_  = ~n2468 ;
  assign \g36259/_0_  = ~n2545 ;
  assign \g36260/_0_  = ~n2563 ;
  assign \g36261/_0_  = ~n2584 ;
  assign \g36262/_0_  = ~n2611 ;
  assign \g36263/_0_  = ~n2623 ;
  assign \g36264/_0_  = ~n2648 ;
  assign \g36265/_0_  = ~n2677 ;
  assign \g36266/_0_  = ~n2703 ;
  assign \g36267/_0_  = ~n2729 ;
  assign \g36268/_0_  = ~n2781 ;
  assign \g36269/_0_  = ~n2809 ;
  assign \g36270/_0_  = ~n2837 ;
  assign \g36271/_0_  = ~n2859 ;
  assign \g36272/_0_  = ~n2887 ;
  assign \g36273/_0_  = ~n2913 ;
  assign \g36274/_0_  = ~n2941 ;
  assign \g36321/_0_  = ~n2981 ;
  assign \g36322/_0_  = ~n3027 ;
  assign \g36323/_0_  = ~n3064 ;
  assign \g36324/_0_  = ~n3107 ;
  assign \g36325/_0_  = ~n3143 ;
  assign \g36341/_0_  = ~n3193 ;
  assign \g36343/_0_  = ~n3204 ;
  assign \g36344/_0_  = ~n3230 ;
  assign \g36345/_0_  = ~n3239 ;
  assign \g36346/_0_  = ~n3264 ;
  assign \g36347/_0_  = ~n3287 ;
  assign \g36348/_0_  = ~n3298 ;
  assign \g36349/_0_  = ~n3301 ;
  assign \g36350/_0_  = ~n3304 ;
  assign \g36351/_0_  = ~n3326 ;
  assign \g36352/_0_  = ~n3364 ;
  assign \g36353/_0_  = ~n3371 ;
  assign \g36354/_0_  = ~n3393 ;
  assign \g36355/_0_  = ~n3411 ;
  assign \g36356/_0_  = ~n3419 ;
  assign \g36357/_0_  = ~n3429 ;
  assign \g36358/_0_  = ~n3432 ;
  assign \g36359/_0_  = ~n3454 ;
  assign \g36360/_0_  = ~n3468 ;
  assign \g36361/_0_  = ~n3492 ;
  assign \g36362/_0_  = ~n3512 ;
  assign \g36363/_0_  = ~n3540 ;
  assign \g36410/_0_  = ~n3583 ;
  assign \g36413/_0_  = ~n3623 ;
  assign \g36414/_0_  = ~n3664 ;
  assign \g36415/_0_  = ~n3705 ;
  assign \g36416/_0_  = ~n3731 ;
  assign \g36424/_0_  = ~n3769 ;
  assign \g36425/_0_  = ~n3807 ;
  assign \g36452/_0_  = ~n3848 ;
  assign \g36455/_0_  = ~n3877 ;
  assign \g36456/_0_  = ~n3902 ;
  assign \g36457/_0_  = ~n3930 ;
  assign \g36458/_0_  = ~n3945 ;
  assign \g36459/_0_  = ~n3967 ;
  assign \g36460/_0_  = ~n3975 ;
  assign \g36461/_0_  = ~n3980 ;
  assign \g36462/_0_  = ~n4006 ;
  assign \g36463/_0_  = ~n4016 ;
  assign \g36464/_0_  = ~n4038 ;
  assign \g36465/_0_  = ~n4066 ;
  assign \g36466/_0_  = ~n4084 ;
  assign \g36467/_0_  = ~n4087 ;
  assign \g36468/_0_  = ~n4109 ;
  assign \g36469/_0_  = ~n4112 ;
  assign \g36470/_0_  = ~n4138 ;
  assign \g36471/_0_  = ~n4147 ;
  assign \g36472/_0_  = ~n4171 ;
  assign \g36473/_0_  = ~n4191 ;
  assign \g36557/_0_  = ~n4198 ;
  assign \g36558/_0_  = ~n4204 ;
  assign \g36559/_0_  = ~n4233 ;
  assign \g36560/_0_  = ~n4262 ;
  assign \g36561/_0_  = ~n4286 ;
  assign \g36562/_0_  = ~n4295 ;
  assign \g36563/_0_  = ~n4307 ;
  assign \g36564/_0_  = ~n4333 ;
  assign \g36565/_0_  = ~n4359 ;
  assign \g36566/_0_  = ~n4362 ;
  assign \g36567/_0_  = ~n4380 ;
  assign \g36568/_0_  = ~n4389 ;
  assign \g36569/_0_  = ~n4392 ;
  assign \g36570/_0_  = ~n4418 ;
  assign \g36571/_0_  = ~n4444 ;
  assign \g36572/_0_  = ~n4466 ;
  assign \g36573/_0_  = ~n4469 ;
  assign \g36574/_0_  = ~n4489 ;
  assign \g36575/_0_  = ~n4505 ;
  assign \g36576/_0_  = ~n4535 ;
  assign \g36577/_0_  = ~n4559 ;
  assign \g36672/_0_  = ~n4582 ;
  assign \g36673/_0_  = ~n4604 ;
  assign \g36674/_0_  = ~n4624 ;
  assign \g38/_0_  = ~n708 ;
  assign \g38_dup47616/_1_  = ~n441 ;
  assign \g39789/u3_syn_4  = n1717 ;
  assign \g40089/_0_  = ~n4732 ;
  assign \g40090/_0_  = ~n4774 ;
  assign \g40092/_0_  = ~n4822 ;
  assign \g40093/_0_  = ~n4855 ;
  assign \g40095/_0_  = ~n4873 ;
  assign \g40096/_0_  = ~n4891 ;
  assign \g40097/_0_  = ~n4909 ;
  assign \g40098/_0_  = ~n4927 ;
  assign \g40099/_0_  = ~n4947 ;
  assign \g40100/_0_  = ~n4973 ;
  assign \g40105/_0_  = ~n4991 ;
  assign \g40106/_0_  = ~n5011 ;
  assign \g40108/_0_  = ~n5049 ;
  assign \g40109/_0_  = ~n5079 ;
  assign \g40219/_0_  = ~n5097 ;
  assign \g40220/_0_  = ~n5119 ;
  assign \g40221/_0_  = ~n5140 ;
  assign \g40222/_0_  = ~n5160 ;
  assign \g40223/_0_  = ~n5180 ;
  assign \g40228/_0_  = ~n5197 ;
  assign \g40434/_0_  = n1164 ;
  assign \g40495/_0_  = ~n5199 ;
  assign \g40760/_0_  = n1168 ;
  assign \g41149/u3_syn_4  = n5200 ;
  assign \g42397/_0_  = ~n364 ;
  assign \g42487/_0_  = ~n383 ;
  assign \g42553/_0_  = ~n373 ;
  assign \g43089/_0_  = ~n862 ;
  assign \g43163/_0_  = ~n454 ;
  assign \g43169/_0_  = ~n474 ;
  assign \g43180/_0_  = ~n414 ;
  assign \g43189_dup/_0_  = ~n515 ;
  assign \g43196/_0_  = ~n581 ;
  assign \g43217/_0_  = ~n887 ;
  assign \g43236/_0_  = ~n718 ;
  assign \g43251/_0_  = ~n401 ;
  assign \g43256/_0_  = ~n541 ;
  assign \g43272/_0_  = ~n827 ;
  assign \g43277/_0_  = ~n752 ;
  assign \g43324/_0_  = ~n768 ;
  assign \g43341/_0_  = ~n498 ;
  assign \g43350/_0_  = ~n661 ;
  assign \g43360/_0_  = ~n671 ;
  assign \g44419/_3_  = ~n5203 ;
  assign \g44452/_3_  = ~n5206 ;
  assign \g44514/_3_  = ~n5212 ;
  assign \g44515/_3_  = ~n5215 ;
  assign \g44516/_3_  = ~n5218 ;
  assign \g44583/_3_  = ~n5221 ;
  assign \g44586/_3_  = ~n5224 ;
  assign \g44587/_3_  = ~n5227 ;
  assign \g44588/_3_  = ~n5230 ;
  assign \g44589/_3_  = ~n5232 ;
  assign \g44590/_3_  = ~n5235 ;
  assign \g44591/_3_  = ~n5238 ;
  assign \g44679/_0_  = ~n5241 ;
  assign \g44680/_3_  = ~n5244 ;
  assign \g44681/_3_  = ~n5247 ;
  assign \g44682/_3_  = ~n5250 ;
  assign \g44686/_3_  = ~n5253 ;
  assign \g44687/_3_  = ~n5256 ;
  assign \g44688/_3_  = n5259 ;
  assign \g44689/_3_  = ~n5262 ;
  assign \g44771/_3_  = ~n5265 ;
  assign \g44785/_3_  = ~n5268 ;
  assign \g44795/_3_  = ~n5271 ;
  assign \g44796/_3_  = ~n5274 ;
  assign \g44906/_3_  = ~n5277 ;
  assign \g44968/_3_  = ~n5280 ;
  assign \g44984/_3_  = ~n5283 ;
  assign \g45042/_3_  = ~n5286 ;
  assign \g45044/_3_  = ~n5289 ;
  assign \g45115/_3_  = ~n5292 ;
  assign \g45116/_3_  = ~n5295 ;
  assign \g46478/_1_  = ~n735 ;
  assign \g46505/_0_  = ~n5318 ;
  assign \g46519/_0_  = ~n426 ;
  assign \g46696/_0_  = ~n5340 ;
  assign \g47017/_2_  = ~n592 ;
  assign \g47072_dup/_0_  = ~n628 ;
  assign \g47395/_0_  = ~n840 ;
  assign \g47397/_0_  = ~n486 ;
  assign \g47401/_0_  = ~n851 ;
  assign \g47404/_0_  = ~n806 ;
  assign \g47458/_0_  = ~n5348 ;
  assign \g47540/_0_  = ~n5371 ;
  assign \g47791/_0_  = ~n618 ;
  assign \state_reg[0]/NET0131_syn_2  = ~\state_reg[0]/NET0131  ;
endmodule
