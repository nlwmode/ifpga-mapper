module top (\DATA_0_0_pad , \DATA_0_10_pad , \DATA_0_11_pad , \DATA_0_12_pad , \DATA_0_13_pad , \DATA_0_14_pad , \DATA_0_15_pad , \DATA_0_16_pad , \DATA_0_17_pad , \DATA_0_18_pad , \DATA_0_19_pad , \DATA_0_1_pad , \DATA_0_20_pad , \DATA_0_21_pad , \DATA_0_22_pad , \DATA_0_23_pad , \DATA_0_24_pad , \DATA_0_25_pad , \DATA_0_26_pad , \DATA_0_27_pad , \DATA_0_28_pad , \DATA_0_29_pad , \DATA_0_2_pad , \DATA_0_30_pad , \DATA_0_31_pad , \DATA_0_3_pad , \DATA_0_4_pad , \DATA_0_5_pad , \DATA_0_6_pad , \DATA_0_7_pad , \DATA_0_8_pad , \DATA_0_9_pad , RESET_pad, \TM0_pad , \TM1_pad , \WX10829_reg/NET0131 , \WX10831_reg/NET0131 , \WX10833_reg/NET0131 , \WX10835_reg/NET0131 , \WX10837_reg/NET0131 , \WX10839_reg/NET0131 , \WX10841_reg/NET0131 , \WX10843_reg/NET0131 , \WX10845_reg/NET0131 , \WX10847_reg/NET0131 , \WX10849_reg/NET0131 , \WX10851_reg/NET0131 , \WX10853_reg/NET0131 , \WX10855_reg/NET0131 , \WX10857_reg/NET0131 , \WX10859_reg/NET0131 , \WX10861_reg/NET0131 , \WX10863_reg/NET0131 , \WX10865_reg/NET0131 , \WX10867_reg/NET0131 , \WX10869_reg/NET0131 , \WX10871_reg/NET0131 , \WX10873_reg/NET0131 , \WX10875_reg/NET0131 , \WX10877_reg/NET0131 , \WX10879_reg/NET0131 , \WX10881_reg/NET0131 , \WX10883_reg/NET0131 , \WX10885_reg/NET0131 , \WX10887_reg/NET0131 , \WX10889_reg/NET0131 , \WX10891_reg/NET0131 , \WX10989_reg/NET0131 , \WX10991_reg/NET0131 , \WX10993_reg/NET0131 , \WX10995_reg/NET0131 , \WX10997_reg/NET0131 , \WX10999_reg/NET0131 , \WX11001_reg/NET0131 , \WX11003_reg/NET0131 , \WX11005_reg/NET0131 , \WX11007_reg/NET0131 , \WX11009_reg/NET0131 , \WX11011_reg/NET0131 , \WX11013_reg/NET0131 , \WX11015_reg/NET0131 , \WX11017_reg/NET0131 , \WX11019_reg/NET0131 , \WX11021_reg/NET0131 , \WX11023_reg/NET0131 , \WX11025_reg/NET0131 , \WX11027_reg/NET0131 , \WX11029_reg/NET0131 , \WX11031_reg/NET0131 , \WX11033_reg/NET0131 , \WX11035_reg/NET0131 , \WX11037_reg/NET0131 , \WX11039_reg/NET0131 , \WX11041_reg/NET0131 , \WX11043_reg/NET0131 , \WX11045_reg/NET0131 , \WX11047_reg/NET0131 , \WX11049_reg/NET0131 , \WX11051_reg/NET0131 , \WX11053_reg/NET0131 , \WX11055_reg/NET0131 , \WX11057_reg/NET0131 , \WX11059_reg/NET0131 , \WX11061_reg/NET0131 , \WX11063_reg/NET0131 , \WX11065_reg/NET0131 , \WX11067_reg/NET0131 , \WX11069_reg/NET0131 , \WX11071_reg/NET0131 , \WX11073_reg/NET0131 , \WX11075_reg/NET0131 , \WX11077_reg/NET0131 , \WX11079_reg/NET0131 , \WX11081_reg/NET0131 , \WX11083_reg/NET0131 , \WX11085_reg/NET0131 , \WX11087_reg/NET0131 , \WX11089_reg/NET0131 , \WX11091_reg/NET0131 , \WX11093_reg/NET0131 , \WX11095_reg/NET0131 , \WX11097_reg/NET0131 , \WX11099_reg/NET0131 , \WX11101_reg/NET0131 , \WX11103_reg/NET0131 , \WX11105_reg/NET0131 , \WX11107_reg/NET0131 , \WX11109_reg/NET0131 , \WX11111_reg/NET0131 , \WX11113_reg/NET0131 , \WX11115_reg/NET0131 , \WX11117_reg/NET0131 , \WX11119_reg/NET0131 , \WX11121_reg/NET0131 , \WX11123_reg/NET0131 , \WX11125_reg/NET0131 , \WX11127_reg/NET0131 , \WX11129_reg/NET0131 , \WX11131_reg/NET0131 , \WX11133_reg/NET0131 , \WX11135_reg/NET0131 , \WX11137_reg/NET0131 , \WX11139_reg/NET0131 , \WX11141_reg/NET0131 , \WX11143_reg/NET0131 , \WX11145_reg/NET0131 , \WX11147_reg/NET0131 , \WX11149_reg/NET0131 , \WX11151_reg/NET0131 , \WX11153_reg/NET0131 , \WX11155_reg/NET0131 , \WX11157_reg/NET0131 , \WX11159_reg/NET0131 , \WX11161_reg/NET0131 , \WX11163_reg/NET0131 , \WX11165_reg/NET0131 , \WX11167_reg/NET0131 , \WX11169_reg/NET0131 , \WX11171_reg/NET0131 , \WX11173_reg/NET0131 , \WX11175_reg/NET0131 , \WX11177_reg/NET0131 , \WX11179_reg/NET0131 , \WX11181_reg/NET0131 , \WX11183_reg/NET0131 , \WX11185_reg/NET0131 , \WX11187_reg/NET0131 , \WX11189_reg/NET0131 , \WX11191_reg/NET0131 , \WX11193_reg/NET0131 , \WX11195_reg/NET0131 , \WX11197_reg/NET0131 , \WX11199_reg/NET0131 , \WX11201_reg/NET0131 , \WX11203_reg/NET0131 , \WX11205_reg/NET0131 , \WX11207_reg/NET0131 , \WX11209_reg/NET0131 , \WX11211_reg/NET0131 , \WX11213_reg/NET0131 , \WX11215_reg/NET0131 , \WX11217_reg/NET0131 , \WX11219_reg/NET0131 , \WX11221_reg/NET0131 , \WX11223_reg/NET0131 , \WX11225_reg/NET0131 , \WX11227_reg/NET0131 , \WX11229_reg/NET0131 , \WX11231_reg/NET0131 , \WX11233_reg/NET0131 , \WX11235_reg/NET0131 , \WX11237_reg/NET0131 , \WX11239_reg/NET0131 , \WX11241_reg/NET0131 , \WX11243_reg/NET0131 , \WX1938_reg/NET0131 , \WX1940_reg/NET0131 , \WX1942_reg/NET0131 , \WX1944_reg/NET0131 , \WX1946_reg/NET0131 , \WX1948_reg/NET0131 , \WX1950_reg/NET0131 , \WX1952_reg/NET0131 , \WX1954_reg/NET0131 , \WX1956_reg/NET0131 , \WX1958_reg/NET0131 , \WX1960_reg/NET0131 , \WX1962_reg/NET0131 , \WX1964_reg/NET0131 , \WX1966_reg/NET0131 , \WX1968_reg/NET0131 , \WX1970_reg/NET0131 , \WX1972_reg/NET0131 , \WX1974_reg/NET0131 , \WX1976_reg/NET0131 , \WX1978_reg/NET0131 , \WX1980_reg/NET0131 , \WX1982_reg/NET0131 , \WX1984_reg/NET0131 , \WX1986_reg/NET0131 , \WX1988_reg/NET0131 , \WX1990_reg/NET0131 , \WX1992_reg/NET0131 , \WX1994_reg/NET0131 , \WX1996_reg/NET0131 , \WX1998_reg/NET0131 , \WX2000_reg/NET0131 , \WX2002_reg/NET0131 , \WX2004_reg/NET0131 , \WX2006_reg/NET0131 , \WX2008_reg/NET0131 , \WX2010_reg/NET0131 , \WX2012_reg/NET0131 , \WX2014_reg/NET0131 , \WX2016_reg/NET0131 , \WX2018_reg/NET0131 , \WX2020_reg/NET0131 , \WX2022_reg/NET0131 , \WX2024_reg/NET0131 , \WX2026_reg/NET0131 , \WX2028_reg/NET0131 , \WX2030_reg/NET0131 , \WX2032_reg/NET0131 , \WX2034_reg/NET0131 , \WX2036_reg/NET0131 , \WX2038_reg/NET0131 , \WX2040_reg/NET0131 , \WX2042_reg/NET0131 , \WX2044_reg/NET0131 , \WX2046_reg/NET0131 , \WX2048_reg/NET0131 , \WX2050_reg/NET0131 , \WX2052_reg/NET0131 , \WX2054_reg/NET0131 , \WX2056_reg/NET0131 , \WX2058_reg/NET0131 , \WX2060_reg/NET0131 , \WX2062_reg/NET0131 , \WX2064_reg/NET0131 , \WX2066_reg/NET0131 , \WX2068_reg/NET0131 , \WX2070_reg/NET0131 , \WX2072_reg/NET0131 , \WX2074_reg/NET0131 , \WX2076_reg/NET0131 , \WX2078_reg/NET0131 , \WX2080_reg/NET0131 , \WX2082_reg/NET0131 , \WX2084_reg/NET0131 , \WX2086_reg/NET0131 , \WX2088_reg/NET0131 , \WX2090_reg/NET0131 , \WX2092_reg/NET0131 , \WX2094_reg/NET0131 , \WX2096_reg/NET0131 , \WX2098_reg/NET0131 , \WX2100_reg/NET0131 , \WX2102_reg/NET0131 , \WX2104_reg/NET0131 , \WX2106_reg/NET0131 , \WX2108_reg/NET0131 , \WX2110_reg/NET0131 , \WX2112_reg/NET0131 , \WX2114_reg/NET0131 , \WX2116_reg/NET0131 , \WX2118_reg/NET0131 , \WX2120_reg/NET0131 , \WX2122_reg/NET0131 , \WX2124_reg/NET0131 , \WX2126_reg/NET0131 , \WX2128_reg/NET0131 , \WX2130_reg/NET0131 , \WX2132_reg/NET0131 , \WX2134_reg/NET0131 , \WX2136_reg/NET0131 , \WX2138_reg/NET0131 , \WX2140_reg/NET0131 , \WX2142_reg/NET0131 , \WX2144_reg/NET0131 , \WX2146_reg/NET0131 , \WX2148_reg/NET0131 , \WX2150_reg/NET0131 , \WX2152_reg/NET0131 , \WX2154_reg/NET0131 , \WX2156_reg/NET0131 , \WX2158_reg/NET0131 , \WX2160_reg/NET0131 , \WX2162_reg/NET0131 , \WX2164_reg/NET0131 , \WX2166_reg/NET0131 , \WX2168_reg/NET0131 , \WX2170_reg/NET0131 , \WX2172_reg/NET0131 , \WX2174_reg/NET0131 , \WX2176_reg/NET0131 , \WX2178_reg/NET0131 , \WX2180_reg/NET0131 , \WX2182_reg/NET0131 , \WX2184_reg/NET0131 , \WX2186_reg/NET0131 , \WX2188_reg/NET0131 , \WX2190_reg/NET0131 , \WX2192_reg/NET0131 , \WX3231_reg/NET0131 , \WX3233_reg/NET0131 , \WX3235_reg/NET0131 , \WX3237_reg/NET0131 , \WX3239_reg/NET0131 , \WX3241_reg/NET0131 , \WX3243_reg/NET0131 , \WX3245_reg/NET0131 , \WX3247_reg/NET0131 , \WX3249_reg/NET0131 , \WX3251_reg/NET0131 , \WX3253_reg/NET0131 , \WX3255_reg/NET0131 , \WX3257_reg/NET0131 , \WX3259_reg/NET0131 , \WX3261_reg/NET0131 , \WX3263_reg/NET0131 , \WX3265_reg/NET0131 , \WX3267_reg/NET0131 , \WX3269_reg/NET0131 , \WX3271_reg/NET0131 , \WX3273_reg/NET0131 , \WX3275_reg/NET0131 , \WX3277_reg/NET0131 , \WX3279_reg/NET0131 , \WX3281_reg/NET0131 , \WX3283_reg/NET0131 , \WX3285_reg/NET0131 , \WX3287_reg/NET0131 , \WX3289_reg/NET0131 , \WX3291_reg/NET0131 , \WX3293_reg/NET0131 , \WX3295_reg/NET0131 , \WX3297_reg/NET0131 , \WX3299_reg/NET0131 , \WX3301_reg/NET0131 , \WX3303_reg/NET0131 , \WX3305_reg/NET0131 , \WX3307_reg/NET0131 , \WX3309_reg/NET0131 , \WX3311_reg/NET0131 , \WX3313_reg/NET0131 , \WX3315_reg/NET0131 , \WX3317_reg/NET0131 , \WX3319_reg/NET0131 , \WX3321_reg/NET0131 , \WX3323_reg/NET0131 , \WX3325_reg/NET0131 , \WX3327_reg/NET0131 , \WX3329_reg/NET0131 , \WX3331_reg/NET0131 , \WX3333_reg/NET0131 , \WX3335_reg/NET0131 , \WX3337_reg/NET0131 , \WX3339_reg/NET0131 , \WX3341_reg/NET0131 , \WX3343_reg/NET0131 , \WX3345_reg/NET0131 , \WX3347_reg/NET0131 , \WX3349_reg/NET0131 , \WX3351_reg/NET0131 , \WX3353_reg/NET0131 , \WX3355_reg/NET0131 , \WX3357_reg/NET0131 , \WX3359_reg/NET0131 , \WX3361_reg/NET0131 , \WX3363_reg/NET0131 , \WX3365_reg/NET0131 , \WX3367_reg/NET0131 , \WX3369_reg/NET0131 , \WX3371_reg/NET0131 , \WX3373_reg/NET0131 , \WX3375_reg/NET0131 , \WX3377_reg/NET0131 , \WX3379_reg/NET0131 , \WX3381_reg/NET0131 , \WX3383_reg/NET0131 , \WX3385_reg/NET0131 , \WX3387_reg/NET0131 , \WX3389_reg/NET0131 , \WX3391_reg/NET0131 , \WX3393_reg/NET0131 , \WX3395_reg/NET0131 , \WX3397_reg/NET0131 , \WX3399_reg/NET0131 , \WX3401_reg/NET0131 , \WX3403_reg/NET0131 , \WX3405_reg/NET0131 , \WX3407_reg/NET0131 , \WX3409_reg/NET0131 , \WX3411_reg/NET0131 , \WX3413_reg/NET0131 , \WX3415_reg/NET0131 , \WX3417_reg/NET0131 , \WX3419_reg/NET0131 , \WX3421_reg/NET0131 , \WX3423_reg/NET0131 , \WX3425_reg/NET0131 , \WX3427_reg/NET0131 , \WX3429_reg/NET0131 , \WX3431_reg/NET0131 , \WX3433_reg/NET0131 , \WX3435_reg/NET0131 , \WX3437_reg/NET0131 , \WX3439_reg/NET0131 , \WX3441_reg/NET0131 , \WX3443_reg/NET0131 , \WX3445_reg/NET0131 , \WX3447_reg/NET0131 , \WX3449_reg/NET0131 , \WX3451_reg/NET0131 , \WX3453_reg/NET0131 , \WX3455_reg/NET0131 , \WX3457_reg/NET0131 , \WX3459_reg/NET0131 , \WX3461_reg/NET0131 , \WX3463_reg/NET0131 , \WX3465_reg/NET0131 , \WX3467_reg/NET0131 , \WX3469_reg/NET0131 , \WX3471_reg/NET0131 , \WX3473_reg/NET0131 , \WX3475_reg/NET0131 , \WX3477_reg/NET0131 , \WX3479_reg/NET0131 , \WX3481_reg/NET0131 , \WX3483_reg/NET0131 , \WX3485_reg/NET0131 , \WX4524_reg/NET0131 , \WX4526_reg/NET0131 , \WX4528_reg/NET0131 , \WX4530_reg/NET0131 , \WX4532_reg/NET0131 , \WX4534_reg/NET0131 , \WX4536_reg/NET0131 , \WX4538_reg/NET0131 , \WX4540_reg/NET0131 , \WX4542_reg/NET0131 , \WX4544_reg/NET0131 , \WX4546_reg/NET0131 , \WX4548_reg/NET0131 , \WX4550_reg/NET0131 , \WX4552_reg/NET0131 , \WX4554_reg/NET0131 , \WX4556_reg/NET0131 , \WX4558_reg/NET0131 , \WX4560_reg/NET0131 , \WX4562_reg/NET0131 , \WX4564_reg/NET0131 , \WX4566_reg/NET0131 , \WX4568_reg/NET0131 , \WX4570_reg/NET0131 , \WX4572_reg/NET0131 , \WX4574_reg/NET0131 , \WX4576_reg/NET0131 , \WX4578_reg/NET0131 , \WX4580_reg/NET0131 , \WX4582_reg/NET0131 , \WX4584_reg/NET0131 , \WX4586_reg/NET0131 , \WX4588_reg/NET0131 , \WX4590_reg/NET0131 , \WX4592_reg/NET0131 , \WX4594_reg/NET0131 , \WX4596_reg/NET0131 , \WX4598_reg/NET0131 , \WX4600_reg/NET0131 , \WX4602_reg/NET0131 , \WX4604_reg/NET0131 , \WX4606_reg/NET0131 , \WX4608_reg/NET0131 , \WX4610_reg/NET0131 , \WX4612_reg/NET0131 , \WX4614_reg/NET0131 , \WX4616_reg/NET0131 , \WX4618_reg/NET0131 , \WX4620_reg/NET0131 , \WX4622_reg/NET0131 , \WX4624_reg/NET0131 , \WX4626_reg/NET0131 , \WX4628_reg/NET0131 , \WX4630_reg/NET0131 , \WX4632_reg/NET0131 , \WX4634_reg/NET0131 , \WX4636_reg/NET0131 , \WX4638_reg/NET0131 , \WX4640_reg/NET0131 , \WX4642_reg/NET0131 , \WX4644_reg/NET0131 , \WX4646_reg/NET0131 , \WX4648_reg/NET0131 , \WX4650_reg/NET0131 , \WX4652_reg/NET0131 , \WX4654_reg/NET0131 , \WX4656_reg/NET0131 , \WX4658_reg/NET0131 , \WX4660_reg/NET0131 , \WX4662_reg/NET0131 , \WX4664_reg/NET0131 , \WX4666_reg/NET0131 , \WX4668_reg/NET0131 , \WX4670_reg/NET0131 , \WX4672_reg/NET0131 , \WX4674_reg/NET0131 , \WX4676_reg/NET0131 , \WX4678_reg/NET0131 , \WX4680_reg/NET0131 , \WX4682_reg/NET0131 , \WX4684_reg/NET0131 , \WX4686_reg/NET0131 , \WX4688_reg/NET0131 , \WX4690_reg/NET0131 , \WX4692_reg/NET0131 , \WX4694_reg/NET0131 , \WX4696_reg/NET0131 , \WX4698_reg/NET0131 , \WX4700_reg/NET0131 , \WX4702_reg/NET0131 , \WX4704_reg/NET0131 , \WX4706_reg/NET0131 , \WX4708_reg/NET0131 , \WX4710_reg/NET0131 , \WX4712_reg/NET0131 , \WX4714_reg/NET0131 , \WX4716_reg/NET0131 , \WX4718_reg/NET0131 , \WX4720_reg/NET0131 , \WX4722_reg/NET0131 , \WX4724_reg/NET0131 , \WX4726_reg/NET0131 , \WX4728_reg/NET0131 , \WX4730_reg/NET0131 , \WX4732_reg/NET0131 , \WX4734_reg/NET0131 , \WX4736_reg/NET0131 , \WX4738_reg/NET0131 , \WX4740_reg/NET0131 , \WX4742_reg/NET0131 , \WX4744_reg/NET0131 , \WX4746_reg/NET0131 , \WX4748_reg/NET0131 , \WX4750_reg/NET0131 , \WX4752_reg/NET0131 , \WX4754_reg/NET0131 , \WX4756_reg/NET0131 , \WX4758_reg/NET0131 , \WX4760_reg/NET0131 , \WX4762_reg/NET0131 , \WX4764_reg/NET0131 , \WX4766_reg/NET0131 , \WX4768_reg/NET0131 , \WX4770_reg/NET0131 , \WX4772_reg/NET0131 , \WX4774_reg/NET0131 , \WX4776_reg/NET0131 , \WX4778_reg/NET0131 , \WX5817_reg/NET0131 , \WX5819_reg/NET0131 , \WX5821_reg/NET0131 , \WX5823_reg/NET0131 , \WX5825_reg/NET0131 , \WX5827_reg/NET0131 , \WX5829_reg/NET0131 , \WX5831_reg/NET0131 , \WX5833_reg/NET0131 , \WX5835_reg/NET0131 , \WX5837_reg/NET0131 , \WX5839_reg/NET0131 , \WX5841_reg/NET0131 , \WX5843_reg/NET0131 , \WX5845_reg/NET0131 , \WX5847_reg/NET0131 , \WX5849_reg/NET0131 , \WX5851_reg/NET0131 , \WX5853_reg/NET0131 , \WX5855_reg/NET0131 , \WX5857_reg/NET0131 , \WX5859_reg/NET0131 , \WX5861_reg/NET0131 , \WX5863_reg/NET0131 , \WX5865_reg/NET0131 , \WX5867_reg/NET0131 , \WX5869_reg/NET0131 , \WX5871_reg/NET0131 , \WX5873_reg/NET0131 , \WX5875_reg/NET0131 , \WX5877_reg/NET0131 , \WX5879_reg/NET0131 , \WX5881_reg/NET0131 , \WX5883_reg/NET0131 , \WX5885_reg/NET0131 , \WX5887_reg/NET0131 , \WX5889_reg/NET0131 , \WX5891_reg/NET0131 , \WX5893_reg/NET0131 , \WX5895_reg/NET0131 , \WX5897_reg/NET0131 , \WX5899_reg/NET0131 , \WX5901_reg/NET0131 , \WX5903_reg/NET0131 , \WX5905_reg/NET0131 , \WX5907_reg/NET0131 , \WX5909_reg/NET0131 , \WX5911_reg/NET0131 , \WX5913_reg/NET0131 , \WX5915_reg/NET0131 , \WX5917_reg/NET0131 , \WX5919_reg/NET0131 , \WX5921_reg/NET0131 , \WX5923_reg/NET0131 , \WX5925_reg/NET0131 , \WX5927_reg/NET0131 , \WX5929_reg/NET0131 , \WX5931_reg/NET0131 , \WX5933_reg/NET0131 , \WX5935_reg/NET0131 , \WX5937_reg/NET0131 , \WX5939_reg/NET0131 , \WX5941_reg/NET0131 , \WX5943_reg/NET0131 , \WX5945_reg/NET0131 , \WX5947_reg/NET0131 , \WX5949_reg/NET0131 , \WX5951_reg/NET0131 , \WX5953_reg/NET0131 , \WX5955_reg/NET0131 , \WX5957_reg/NET0131 , \WX5959_reg/NET0131 , \WX5961_reg/NET0131 , \WX5963_reg/NET0131 , \WX5965_reg/NET0131 , \WX5967_reg/NET0131 , \WX5969_reg/NET0131 , \WX5971_reg/NET0131 , \WX5973_reg/NET0131 , \WX5975_reg/NET0131 , \WX5977_reg/NET0131 , \WX5979_reg/NET0131 , \WX5981_reg/NET0131 , \WX5983_reg/NET0131 , \WX5985_reg/NET0131 , \WX5987_reg/NET0131 , \WX5989_reg/NET0131 , \WX5991_reg/NET0131 , \WX5993_reg/NET0131 , \WX5995_reg/NET0131 , \WX5997_reg/NET0131 , \WX5999_reg/NET0131 , \WX6001_reg/NET0131 , \WX6003_reg/NET0131 , \WX6005_reg/NET0131 , \WX6007_reg/NET0131 , \WX6009_reg/NET0131 , \WX6011_reg/NET0131 , \WX6013_reg/NET0131 , \WX6015_reg/NET0131 , \WX6017_reg/NET0131 , \WX6019_reg/NET0131 , \WX6021_reg/NET0131 , \WX6023_reg/NET0131 , \WX6025_reg/NET0131 , \WX6027_reg/NET0131 , \WX6029_reg/NET0131 , \WX6031_reg/NET0131 , \WX6033_reg/NET0131 , \WX6035_reg/NET0131 , \WX6037_reg/NET0131 , \WX6039_reg/NET0131 , \WX6041_reg/NET0131 , \WX6043_reg/NET0131 , \WX6045_reg/NET0131 , \WX6047_reg/NET0131 , \WX6049_reg/NET0131 , \WX6051_reg/NET0131 , \WX6053_reg/NET0131 , \WX6055_reg/NET0131 , \WX6057_reg/NET0131 , \WX6059_reg/NET0131 , \WX6061_reg/NET0131 , \WX6063_reg/NET0131 , \WX6065_reg/NET0131 , \WX6067_reg/NET0131 , \WX6069_reg/NET0131 , \WX6071_reg/NET0131 , \WX645_reg/NET0131 , \WX647_reg/NET0131 , \WX649_reg/NET0131 , \WX651_reg/NET0131 , \WX653_reg/NET0131 , \WX655_reg/NET0131 , \WX657_reg/NET0131 , \WX659_reg/NET0131 , \WX661_reg/NET0131 , \WX663_reg/NET0131 , \WX665_reg/NET0131 , \WX667_reg/NET0131 , \WX669_reg/NET0131 , \WX671_reg/NET0131 , \WX673_reg/NET0131 , \WX675_reg/NET0131 , \WX677_reg/NET0131 , \WX679_reg/NET0131 , \WX681_reg/NET0131 , \WX683_reg/NET0131 , \WX685_reg/NET0131 , \WX687_reg/NET0131 , \WX689_reg/NET0131 , \WX691_reg/NET0131 , \WX693_reg/NET0131 , \WX695_reg/NET0131 , \WX697_reg/NET0131 , \WX699_reg/NET0131 , \WX701_reg/NET0131 , \WX703_reg/NET0131 , \WX705_reg/NET0131 , \WX707_reg/NET0131 , \WX709_reg/NET0131 , \WX7110_reg/NET0131 , \WX7112_reg/NET0131 , \WX7114_reg/NET0131 , \WX7116_reg/NET0131 , \WX7118_reg/NET0131 , \WX711_reg/NET0131 , \WX7120_reg/NET0131 , \WX7122_reg/NET0131 , \WX7124_reg/NET0131 , \WX7126_reg/NET0131 , \WX7128_reg/NET0131 , \WX7130_reg/NET0131 , \WX7132_reg/NET0131 , \WX7134_reg/NET0131 , \WX7136_reg/NET0131 , \WX7138_reg/NET0131 , \WX713_reg/NET0131 , \WX7140_reg/NET0131 , \WX7142_reg/NET0131 , \WX7144_reg/NET0131 , \WX7146_reg/NET0131 , \WX7148_reg/NET0131 , \WX7150_reg/NET0131 , \WX7152_reg/NET0131 , \WX7154_reg/NET0131 , \WX7156_reg/NET0131 , \WX7158_reg/NET0131 , \WX715_reg/NET0131 , \WX7160_reg/NET0131 , \WX7162_reg/NET0131 , \WX7164_reg/NET0131 , \WX7166_reg/NET0131 , \WX7168_reg/NET0131 , \WX7170_reg/NET0131 , \WX7172_reg/NET0131 , \WX7174_reg/NET0131 , \WX7176_reg/NET0131 , \WX7178_reg/NET0131 , \WX717_reg/NET0131 , \WX7180_reg/NET0131 , \WX7182_reg/NET0131 , \WX7184_reg/NET0131 , \WX7186_reg/NET0131 , \WX7188_reg/NET0131 , \WX7190_reg/NET0131 , \WX7192_reg/NET0131 , \WX7194_reg/NET0131 , \WX7196_reg/NET0131 , \WX7198_reg/NET0131 , \WX719_reg/NET0131 , \WX7200_reg/NET0131 , \WX7202_reg/NET0131 , \WX7204_reg/NET0131 , \WX7206_reg/NET0131 , \WX7208_reg/NET0131 , \WX7210_reg/NET0131 , \WX7212_reg/NET0131 , \WX7214_reg/NET0131 , \WX7216_reg/NET0131 , \WX7218_reg/NET0131 , \WX721_reg/NET0131 , \WX7220_reg/NET0131 , \WX7222_reg/NET0131 , \WX7224_reg/NET0131 , \WX7226_reg/NET0131 , \WX7228_reg/NET0131 , \WX7230_reg/NET0131 , \WX7232_reg/NET0131 , \WX7234_reg/NET0131 , \WX7236_reg/NET0131 , \WX7238_reg/NET0131 , \WX723_reg/NET0131 , \WX7240_reg/NET0131 , \WX7242_reg/NET0131 , \WX7244_reg/NET0131 , \WX7246_reg/NET0131 , \WX7248_reg/NET0131 , \WX7250_reg/NET0131 , \WX7252_reg/NET0131 , \WX7254_reg/NET0131 , \WX7256_reg/NET0131 , \WX7258_reg/NET0131 , \WX725_reg/NET0131 , \WX7260_reg/NET0131 , \WX7262_reg/NET0131 , \WX7264_reg/NET0131 , \WX7266_reg/NET0131 , \WX7268_reg/NET0131 , \WX7270_reg/NET0131 , \WX7272_reg/NET0131 , \WX7274_reg/NET0131 , \WX7276_reg/NET0131 , \WX7278_reg/NET0131 , \WX727_reg/NET0131 , \WX7280_reg/NET0131 , \WX7282_reg/NET0131 , \WX7284_reg/NET0131 , \WX7286_reg/NET0131 , \WX7288_reg/NET0131 , \WX7290_reg/NET0131 , \WX7292_reg/NET0131 , \WX7294_reg/NET0131 , \WX7296_reg/NET0131 , \WX7298_reg/NET0131 , \WX729_reg/NET0131 , \WX7300_reg/NET0131 , \WX7302_reg/NET0131 , \WX7304_reg/NET0131 , \WX7306_reg/NET0131 , \WX7308_reg/NET0131 , \WX7310_reg/NET0131 , \WX7312_reg/NET0131 , \WX7314_reg/NET0131 , \WX7316_reg/NET0131 , \WX7318_reg/NET0131 , \WX731_reg/NET0131 , \WX7320_reg/NET0131 , \WX7322_reg/NET0131 , \WX7324_reg/NET0131 , \WX7326_reg/NET0131 , \WX7328_reg/NET0131 , \WX7330_reg/NET0131 , \WX7332_reg/NET0131 , \WX7334_reg/NET0131 , \WX7336_reg/NET0131 , \WX7338_reg/NET0131 , \WX733_reg/NET0131 , \WX7340_reg/NET0131 , \WX7342_reg/NET0131 , \WX7344_reg/NET0131 , \WX7346_reg/NET0131 , \WX7348_reg/NET0131 , \WX7350_reg/NET0131 , \WX7352_reg/NET0131 , \WX7354_reg/NET0131 , \WX7356_reg/NET0131 , \WX7358_reg/NET0131 , \WX735_reg/NET0131 , \WX7360_reg/NET0131 , \WX7362_reg/NET0131 , \WX7364_reg/NET0131 , \WX737_reg/NET0131 , \WX739_reg/NET0131 , \WX741_reg/NET0131 , \WX743_reg/NET0131 , \WX745_reg/NET0131 , \WX747_reg/NET0131 , \WX749_reg/NET0131 , \WX751_reg/NET0131 , \WX753_reg/NET0131 , \WX755_reg/NET0131 , \WX757_reg/NET0131 , \WX759_reg/NET0131 , \WX761_reg/NET0131 , \WX763_reg/NET0131 , \WX765_reg/NET0131 , \WX767_reg/NET0131 , \WX769_reg/NET0131 , \WX771_reg/NET0131 , \WX773_reg/NET0131 , \WX775_reg/NET0131 , \WX777_reg/NET0131 , \WX779_reg/NET0131 , \WX781_reg/NET0131 , \WX783_reg/NET0131 , \WX785_reg/NET0131 , \WX787_reg/NET0131 , \WX789_reg/NET0131 , \WX791_reg/NET0131 , \WX793_reg/NET0131 , \WX795_reg/NET0131 , \WX797_reg/NET0131 , \WX799_reg/NET0131 , \WX801_reg/NET0131 , \WX803_reg/NET0131 , \WX805_reg/NET0131 , \WX807_reg/NET0131 , \WX809_reg/NET0131 , \WX811_reg/NET0131 , \WX813_reg/NET0131 , \WX815_reg/NET0131 , \WX817_reg/NET0131 , \WX819_reg/NET0131 , \WX821_reg/NET0131 , \WX823_reg/NET0131 , \WX825_reg/NET0131 , \WX827_reg/NET0131 , \WX829_reg/NET0131 , \WX831_reg/NET0131 , \WX833_reg/NET0131 , \WX835_reg/NET0131 , \WX837_reg/NET0131 , \WX839_reg/NET0131 , \WX8403_reg/NET0131 , \WX8405_reg/NET0131 , \WX8407_reg/NET0131 , \WX8409_reg/NET0131 , \WX8411_reg/NET0131 , \WX8413_reg/NET0131 , \WX8415_reg/NET0131 , \WX8417_reg/NET0131 , \WX8419_reg/NET0131 , \WX841_reg/NET0131 , \WX8421_reg/NET0131 , \WX8423_reg/NET0131 , \WX8425_reg/NET0131 , \WX8427_reg/NET0131 , \WX8429_reg/NET0131 , \WX8431_reg/NET0131 , \WX8433_reg/NET0131 , \WX8435_reg/NET0131 , \WX8437_reg/NET0131 , \WX8439_reg/NET0131 , \WX843_reg/NET0131 , \WX8441_reg/NET0131 , \WX8443_reg/NET0131 , \WX8445_reg/NET0131 , \WX8447_reg/NET0131 , \WX8449_reg/NET0131 , \WX8451_reg/NET0131 , \WX8453_reg/NET0131 , \WX8455_reg/NET0131 , \WX8457_reg/NET0131 , \WX8459_reg/NET0131 , \WX845_reg/NET0131 , \WX8461_reg/NET0131 , \WX8463_reg/NET0131 , \WX8465_reg/NET0131 , \WX8467_reg/NET0131 , \WX8469_reg/NET0131 , \WX8471_reg/NET0131 , \WX8473_reg/NET0131 , \WX8475_reg/NET0131 , \WX8477_reg/NET0131 , \WX8479_reg/NET0131 , \WX847_reg/NET0131 , \WX8481_reg/NET0131 , \WX8483_reg/NET0131 , \WX8485_reg/NET0131 , \WX8487_reg/NET0131 , \WX8489_reg/NET0131 , \WX8491_reg/NET0131 , \WX8493_reg/NET0131 , \WX8495_reg/NET0131 , \WX8497_reg/NET0131 , \WX8499_reg/NET0131 , \WX849_reg/NET0131 , \WX8501_reg/NET0131 , \WX8503_reg/NET0131 , \WX8505_reg/NET0131 , \WX8507_reg/NET0131 , \WX8509_reg/NET0131 , \WX8511_reg/NET0131 , \WX8513_reg/NET0131 , \WX8515_reg/NET0131 , \WX8517_reg/NET0131 , \WX8519_reg/NET0131 , \WX851_reg/NET0131 , \WX8521_reg/NET0131 , \WX8523_reg/NET0131 , \WX8525_reg/NET0131 , \WX8527_reg/NET0131 , \WX8529_reg/NET0131 , \WX8531_reg/NET0131 , \WX8533_reg/NET0131 , \WX8535_reg/NET0131 , \WX8537_reg/NET0131 , \WX8539_reg/NET0131 , \WX853_reg/NET0131 , \WX8541_reg/NET0131 , \WX8543_reg/NET0131 , \WX8545_reg/NET0131 , \WX8547_reg/NET0131 , \WX8549_reg/NET0131 , \WX8551_reg/NET0131 , \WX8553_reg/NET0131 , \WX8555_reg/NET0131 , \WX8557_reg/NET0131 , \WX8559_reg/NET0131 , \WX855_reg/NET0131 , \WX8561_reg/NET0131 , \WX8563_reg/NET0131 , \WX8565_reg/NET0131 , \WX8567_reg/NET0131 , \WX8569_reg/NET0131 , \WX8571_reg/NET0131 , \WX8573_reg/NET0131 , \WX8575_reg/NET0131 , \WX8577_reg/NET0131 , \WX8579_reg/NET0131 , \WX857_reg/NET0131 , \WX8581_reg/NET0131 , \WX8583_reg/NET0131 , \WX8585_reg/NET0131 , \WX8587_reg/NET0131 , \WX8589_reg/NET0131 , \WX8591_reg/NET0131 , \WX8593_reg/NET0131 , \WX8595_reg/NET0131 , \WX8597_reg/NET0131 , \WX8599_reg/NET0131 , \WX859_reg/NET0131 , \WX8601_reg/NET0131 , \WX8603_reg/NET0131 , \WX8605_reg/NET0131 , \WX8607_reg/NET0131 , \WX8609_reg/NET0131 , \WX8611_reg/NET0131 , \WX8613_reg/NET0131 , \WX8615_reg/NET0131 , \WX8617_reg/NET0131 , \WX8619_reg/NET0131 , \WX861_reg/NET0131 , \WX8621_reg/NET0131 , \WX8623_reg/NET0131 , \WX8625_reg/NET0131 , \WX8627_reg/NET0131 , \WX8629_reg/NET0131 , \WX8631_reg/NET0131 , \WX8633_reg/NET0131 , \WX8635_reg/NET0131 , \WX8637_reg/NET0131 , \WX8639_reg/NET0131 , \WX863_reg/NET0131 , \WX8641_reg/NET0131 , \WX8643_reg/NET0131 , \WX8645_reg/NET0131 , \WX8647_reg/NET0131 , \WX8649_reg/NET0131 , \WX8651_reg/NET0131 , \WX8653_reg/NET0131 , \WX8655_reg/NET0131 , \WX8657_reg/NET0131 , \WX865_reg/NET0131 , \WX867_reg/NET0131 , \WX869_reg/NET0131 , \WX871_reg/NET0131 , \WX873_reg/NET0131 , \WX875_reg/NET0131 , \WX877_reg/NET0131 , \WX879_reg/NET0131 , \WX881_reg/NET0131 , \WX883_reg/NET0131 , \WX885_reg/NET0131 , \WX887_reg/NET0131 , \WX889_reg/NET0131 , \WX891_reg/NET0131 , \WX893_reg/NET0131 , \WX895_reg/NET0131 , \WX897_reg/NET0131 , \WX899_reg/NET0131 , \WX9696_reg/NET0131 , \WX9698_reg/NET0131 , \WX9700_reg/NET0131 , \WX9702_reg/NET0131 , \WX9704_reg/NET0131 , \WX9706_reg/NET0131 , \WX9708_reg/NET0131 , \WX9710_reg/NET0131 , \WX9712_reg/NET0131 , \WX9714_reg/NET0131 , \WX9716_reg/NET0131 , \WX9718_reg/NET0131 , \WX9720_reg/NET0131 , \WX9722_reg/NET0131 , \WX9724_reg/NET0131 , \WX9726_reg/NET0131 , \WX9728_reg/NET0131 , \WX9730_reg/NET0131 , \WX9732_reg/NET0131 , \WX9734_reg/NET0131 , \WX9736_reg/NET0131 , \WX9738_reg/NET0131 , \WX9740_reg/NET0131 , \WX9742_reg/NET0131 , \WX9744_reg/NET0131 , \WX9746_reg/NET0131 , \WX9748_reg/NET0131 , \WX9750_reg/NET0131 , \WX9752_reg/NET0131 , \WX9754_reg/NET0131 , \WX9756_reg/NET0131 , \WX9758_reg/NET0131 , \WX9760_reg/NET0131 , \WX9762_reg/NET0131 , \WX9764_reg/NET0131 , \WX9766_reg/NET0131 , \WX9768_reg/NET0131 , \WX9770_reg/NET0131 , \WX9772_reg/NET0131 , \WX9774_reg/NET0131 , \WX9776_reg/NET0131 , \WX9778_reg/NET0131 , \WX9780_reg/NET0131 , \WX9782_reg/NET0131 , \WX9784_reg/NET0131 , \WX9786_reg/NET0131 , \WX9788_reg/NET0131 , \WX9790_reg/NET0131 , \WX9792_reg/NET0131 , \WX9794_reg/NET0131 , \WX9796_reg/NET0131 , \WX9798_reg/NET0131 , \WX9800_reg/NET0131 , \WX9802_reg/NET0131 , \WX9804_reg/NET0131 , \WX9806_reg/NET0131 , \WX9808_reg/NET0131 , \WX9810_reg/NET0131 , \WX9812_reg/NET0131 , \WX9814_reg/NET0131 , \WX9816_reg/NET0131 , \WX9818_reg/NET0131 , \WX9820_reg/NET0131 , \WX9822_reg/NET0131 , \WX9824_reg/NET0131 , \WX9826_reg/NET0131 , \WX9828_reg/NET0131 , \WX9830_reg/NET0131 , \WX9832_reg/NET0131 , \WX9834_reg/NET0131 , \WX9836_reg/NET0131 , \WX9838_reg/NET0131 , \WX9840_reg/NET0131 , \WX9842_reg/NET0131 , \WX9844_reg/NET0131 , \WX9846_reg/NET0131 , \WX9848_reg/NET0131 , \WX9850_reg/NET0131 , \WX9852_reg/NET0131 , \WX9854_reg/NET0131 , \WX9856_reg/NET0131 , \WX9858_reg/NET0131 , \WX9860_reg/NET0131 , \WX9862_reg/NET0131 , \WX9864_reg/NET0131 , \WX9866_reg/NET0131 , \WX9868_reg/NET0131 , \WX9870_reg/NET0131 , \WX9872_reg/NET0131 , \WX9874_reg/NET0131 , \WX9876_reg/NET0131 , \WX9878_reg/NET0131 , \WX9880_reg/NET0131 , \WX9882_reg/NET0131 , \WX9884_reg/NET0131 , \WX9886_reg/NET0131 , \WX9888_reg/NET0131 , \WX9890_reg/NET0131 , \WX9892_reg/NET0131 , \WX9894_reg/NET0131 , \WX9896_reg/NET0131 , \WX9898_reg/NET0131 , \WX9900_reg/NET0131 , \WX9902_reg/NET0131 , \WX9904_reg/NET0131 , \WX9906_reg/NET0131 , \WX9908_reg/NET0131 , \WX9910_reg/NET0131 , \WX9912_reg/NET0131 , \WX9914_reg/NET0131 , \WX9916_reg/NET0131 , \WX9918_reg/NET0131 , \WX9920_reg/NET0131 , \WX9922_reg/NET0131 , \WX9924_reg/NET0131 , \WX9926_reg/NET0131 , \WX9928_reg/NET0131 , \WX9930_reg/NET0131 , \WX9932_reg/NET0131 , \WX9934_reg/NET0131 , \WX9936_reg/NET0131 , \WX9938_reg/NET0131 , \WX9940_reg/NET0131 , \WX9942_reg/NET0131 , \WX9944_reg/NET0131 , \WX9946_reg/NET0131 , \WX9948_reg/NET0131 , \WX9950_reg/NET0131 , \_2077__reg/NET0131 , \_2078__reg/NET0131 , \_2079__reg/NET0131 , \_2080__reg/NET0131 , \_2081__reg/NET0131 , \_2082__reg/NET0131 , \_2083__reg/NET0131 , \_2084__reg/NET0131 , \_2085__reg/NET0131 , \_2086__reg/NET0131 , \_2087__reg/NET0131 , \_2088__reg/NET0131 , \_2089__reg/NET0131 , \_2090__reg/NET0131 , \_2091__reg/NET0131 , \_2092__reg/NET0131 , \_2093__reg/NET0131 , \_2094__reg/NET0131 , \_2095__reg/NET0131 , \_2096__reg/NET0131 , \_2097__reg/NET0131 , \_2098__reg/NET0131 , \_2099__reg/NET0131 , \_2100__reg/NET0131 , \_2101__reg/NET0131 , \_2102__reg/NET0131 , \_2103__reg/NET0131 , \_2104__reg/NET0131 , \_2105__reg/NET0131 , \_2106__reg/NET0131 , \_2107__reg/NET0131 , \_2108__reg/NET0131 , \_2109__reg/NET0131 , \_2110__reg/NET0131 , \_2111__reg/NET0131 , \_2112__reg/NET0131 , \_2113__reg/NET0131 , \_2114__reg/NET0131 , \_2115__reg/NET0131 , \_2116__reg/NET0131 , \_2117__reg/NET0131 , \_2118__reg/NET0131 , \_2119__reg/NET0131 , \_2120__reg/NET0131 , \_2121__reg/NET0131 , \_2122__reg/NET0131 , \_2123__reg/NET0131 , \_2124__reg/NET0131 , \_2125__reg/NET0131 , \_2126__reg/NET0131 , \_2127__reg/NET0131 , \_2128__reg/NET0131 , \_2129__reg/NET0131 , \_2130__reg/NET0131 , \_2131__reg/NET0131 , \_2132__reg/NET0131 , \_2133__reg/NET0131 , \_2134__reg/NET0131 , \_2135__reg/NET0131 , \_2136__reg/NET0131 , \_2137__reg/NET0131 , \_2138__reg/NET0131 , \_2139__reg/NET0131 , \_2140__reg/NET0131 , \_2141__reg/NET0131 , \_2142__reg/NET0131 , \_2143__reg/NET0131 , \_2144__reg/NET0131 , \_2145__reg/NET0131 , \_2146__reg/NET0131 , \_2147__reg/NET0131 , \_2148__reg/NET0131 , \_2149__reg/NET0131 , \_2150__reg/NET0131 , \_2151__reg/NET0131 , \_2152__reg/NET0131 , \_2153__reg/NET0131 , \_2154__reg/NET0131 , \_2155__reg/NET0131 , \_2156__reg/NET0131 , \_2157__reg/NET0131 , \_2158__reg/NET0131 , \_2159__reg/NET0131 , \_2160__reg/NET0131 , \_2161__reg/NET0131 , \_2162__reg/NET0131 , \_2163__reg/NET0131 , \_2164__reg/NET0131 , \_2165__reg/NET0131 , \_2166__reg/NET0131 , \_2167__reg/NET0131 , \_2168__reg/NET0131 , \_2169__reg/NET0131 , \_2170__reg/NET0131 , \_2171__reg/NET0131 , \_2172__reg/NET0131 , \_2173__reg/NET0131 , \_2174__reg/NET0131 , \_2175__reg/NET0131 , \_2176__reg/NET0131 , \_2177__reg/NET0131 , \_2178__reg/NET0131 , \_2179__reg/NET0131 , \_2180__reg/NET0131 , \_2181__reg/NET0131 , \_2182__reg/NET0131 , \_2183__reg/NET0131 , \_2184__reg/NET0131 , \_2185__reg/NET0131 , \_2186__reg/NET0131 , \_2187__reg/NET0131 , \_2188__reg/NET0131 , \_2189__reg/NET0131 , \_2190__reg/NET0131 , \_2191__reg/NET0131 , \_2192__reg/NET0131 , \_2193__reg/NET0131 , \_2194__reg/NET0131 , \_2195__reg/NET0131 , \_2196__reg/NET0131 , \_2197__reg/NET0131 , \_2198__reg/NET0131 , \_2199__reg/NET0131 , \_2200__reg/NET0131 , \_2201__reg/NET0131 , \_2202__reg/NET0131 , \_2203__reg/NET0131 , \_2204__reg/NET0131 , \_2205__reg/NET0131 , \_2206__reg/NET0131 , \_2207__reg/NET0131 , \_2208__reg/NET0131 , \_2209__reg/NET0131 , \_2210__reg/NET0131 , \_2211__reg/NET0131 , \_2212__reg/NET0131 , \_2213__reg/NET0131 , \_2214__reg/NET0131 , \_2215__reg/NET0131 , \_2216__reg/NET0131 , \_2217__reg/NET0131 , \_2218__reg/NET0131 , \_2219__reg/NET0131 , \_2220__reg/NET0131 , \_2221__reg/NET0131 , \_2222__reg/NET0131 , \_2223__reg/NET0131 , \_2224__reg/NET0131 , \_2225__reg/NET0131 , \_2226__reg/NET0131 , \_2227__reg/NET0131 , \_2228__reg/NET0131 , \_2229__reg/NET0131 , \_2230__reg/NET0131 , \_2231__reg/NET0131 , \_2232__reg/NET0131 , \_2233__reg/NET0131 , \_2234__reg/NET0131 , \_2235__reg/NET0131 , \_2236__reg/NET0131 , \_2237__reg/NET0131 , \_2238__reg/NET0131 , \_2239__reg/NET0131 , \_2240__reg/NET0131 , \_2241__reg/NET0131 , \_2242__reg/NET0131 , \_2243__reg/NET0131 , \_2244__reg/NET0131 , \_2245__reg/NET0131 , \_2246__reg/NET0131 , \_2247__reg/NET0131 , \_2248__reg/NET0131 , \_2249__reg/NET0131 , \_2250__reg/NET0131 , \_2251__reg/NET0131 , \_2252__reg/NET0131 , \_2253__reg/NET0131 , \_2254__reg/NET0131 , \_2255__reg/NET0131 , \_2256__reg/NET0131 , \_2257__reg/NET0131 , \_2258__reg/NET0131 , \_2259__reg/NET0131 , \_2260__reg/NET0131 , \_2261__reg/NET0131 , \_2262__reg/NET0131 , \_2263__reg/NET0131 , \_2264__reg/NET0131 , \_2265__reg/NET0131 , \_2266__reg/NET0131 , \_2267__reg/NET0131 , \_2268__reg/NET0131 , \_2269__reg/NET0131 , \_2270__reg/NET0131 , \_2271__reg/NET0131 , \_2272__reg/NET0131 , \_2273__reg/NET0131 , \_2274__reg/NET0131 , \_2275__reg/NET0131 , \_2276__reg/NET0131 , \_2277__reg/NET0131 , \_2278__reg/NET0131 , \_2279__reg/NET0131 , \_2280__reg/NET0131 , \_2281__reg/NET0131 , \_2282__reg/NET0131 , \_2283__reg/NET0131 , \_2284__reg/NET0131 , \_2285__reg/NET0131 , \_2286__reg/NET0131 , \_2287__reg/NET0131 , \_2288__reg/NET0131 , \_2289__reg/NET0131 , \_2290__reg/NET0131 , \_2291__reg/NET0131 , \_2292__reg/NET0131 , \_2293__reg/NET0131 , \_2294__reg/NET0131 , \_2295__reg/NET0131 , \_2296__reg/NET0131 , \_2297__reg/NET0131 , \_2298__reg/NET0131 , \_2299__reg/NET0131 , \_2300__reg/NET0131 , \_2301__reg/NET0131 , \_2302__reg/NET0131 , \_2303__reg/NET0131 , \_2304__reg/NET0131 , \_2305__reg/NET0131 , \_2306__reg/NET0131 , \_2307__reg/NET0131 , \_2308__reg/NET0131 , \_2309__reg/NET0131 , \_2310__reg/NET0131 , \_2311__reg/NET0131 , \_2312__reg/NET0131 , \_2313__reg/NET0131 , \_2314__reg/NET0131 , \_2315__reg/NET0131 , \_2316__reg/NET0131 , \_2317__reg/NET0131 , \_2318__reg/NET0131 , \_2319__reg/NET0131 , \_2320__reg/NET0131 , \_2321__reg/NET0131 , \_2322__reg/NET0131 , \_2323__reg/NET0131 , \_2324__reg/NET0131 , \_2325__reg/NET0131 , \_2326__reg/NET0131 , \_2327__reg/NET0131 , \_2328__reg/NET0131 , \_2329__reg/NET0131 , \_2330__reg/NET0131 , \_2331__reg/NET0131 , \_2332__reg/NET0131 , \_2333__reg/NET0131 , \_2334__reg/NET0131 , \_2335__reg/NET0131 , \_2336__reg/NET0131 , \_2337__reg/NET0131 , \_2338__reg/NET0131 , \_2339__reg/NET0131 , \_2340__reg/NET0131 , \_2341__reg/NET0131 , \_2342__reg/NET0131 , \_2343__reg/NET0131 , \_2344__reg/NET0131 , \_2345__reg/NET0131 , \_2346__reg/NET0131 , \_2347__reg/NET0131 , \_2348__reg/NET0131 , \_2349__reg/NET0131 , \_2350__reg/NET0131 , \_2351__reg/NET0131 , \_2352__reg/NET0131 , \_2353__reg/NET0131 , \_2354__reg/NET0131 , \_2355__reg/NET0131 , \_2356__reg/NET0131 , \_2357__reg/NET0131 , \_2358__reg/NET0131 , \_2359__reg/NET0131 , \_2360__reg/NET0131 , \_2361__reg/NET0131 , \_2362__reg/NET0131 , \_2363__reg/NET0131 , \_2364__reg/NET0131 , \DATA_9_0_pad , \DATA_9_10_pad , \DATA_9_11_pad , \DATA_9_12_pad , \DATA_9_13_pad , \DATA_9_14_pad , \DATA_9_15_pad , \DATA_9_16_pad , \DATA_9_17_pad , \DATA_9_18_pad , \DATA_9_19_pad , \DATA_9_1_pad , \DATA_9_20_pad , \DATA_9_21_pad , \DATA_9_22_pad , \DATA_9_23_pad , \DATA_9_24_pad , \DATA_9_25_pad , \DATA_9_26_pad , \DATA_9_27_pad , \DATA_9_28_pad , \DATA_9_29_pad , \DATA_9_2_pad , \DATA_9_30_pad , \DATA_9_31_pad , \DATA_9_3_pad , \DATA_9_4_pad , \DATA_9_5_pad , \DATA_9_6_pad , \DATA_9_7_pad , \DATA_9_8_pad , \DATA_9_9_pad , \_al_n0 , \_al_n1 , \g19/_0_ , \g35/_0_ , \g36/_0_ , \g40/_0_ , \g55780/_0_ , \g55783/_0_ , \g55795/_0_ , \g55796/_0_ , \g55797/_0_ , \g55798/_0_ , \g55799/_0_ , \g55800/_0_ , \g55801/_0_ , \g55802/_0_ , \g55803/_0_ , \g55834/_0_ , \g55835/_0_ , \g55836/_0_ , \g55837/_0_ , \g55838/_0_ , \g55839/_0_ , \g55840/_0_ , \g55841/_0_ , \g55842/_0_ , \g55856/_0_ , \g55894/_0_ , \g55895/_0_ , \g55896/_0_ , \g55897/_0_ , \g55898/_0_ , \g55899/_0_ , \g55900/_0_ , \g55901/_0_ , \g55902/_0_ , \g55916/_0_ , \g55953/_0_ , \g55954/_0_ , \g55955/_0_ , \g55956/_0_ , \g55957/_0_ , \g55958/_0_ , \g55959/_0_ , \g55960/_0_ , \g55961/_0_ , \g55975/_0_ , \g56012/_0_ , \g56013/_0_ , \g56014/_0_ , \g56015/_0_ , \g56016/_0_ , \g56017/_0_ , \g56018/_0_ , \g56019/_0_ , \g56020/_0_ , \g56034/_0_ , \g56071/_0_ , \g56072/_0_ , \g56073/_0_ , \g56074/_0_ , \g56075/_0_ , \g56076/_0_ , \g56077/_0_ , \g56078/_0_ , \g56079/_0_ , \g56093/_0_ , \g56130/_0_ , \g56131/_0_ , \g56132/_0_ , \g56133/_0_ , \g56134/_0_ , \g56135/_0_ , \g56136/_0_ , \g56137/_0_ , \g56138/_0_ , \g56152/_0_ , \g56189/_0_ , \g56190/_0_ , \g56191/_0_ , \g56192/_0_ , \g56193/_0_ , \g56194/_0_ , \g56195/_0_ , \g56196/_0_ , \g56197/_0_ , \g56211/_0_ , \g56248/_0_ , \g56249/_0_ , \g56250/_0_ , \g56251/_0_ , \g56252/_0_ , \g56253/_0_ , \g56254/_0_ , \g56255/_0_ , \g56256/_0_ , \g56270/_0_ , \g56307/_0_ , \g56308/_0_ , \g56309/_0_ , \g56310/_0_ , \g56311/_0_ , \g56312/_0_ , \g56313/_0_ , \g56314/_0_ , \g56315/_0_ , \g56329/_0_ , \g56366/_0_ , \g56367/_0_ , \g56368/_0_ , \g56369/_0_ , \g56370/_0_ , \g56371/_0_ , \g56372/_0_ , \g56373/_0_ , \g56374/_0_ , \g56388/_0_ , \g56425/_0_ , \g56426/_0_ , \g56427/_0_ , \g56428/_0_ , \g56429/_0_ , \g56430/_0_ , \g56431/_0_ , \g56432/_0_ , \g56433/_0_ , \g56447/_0_ , \g56484/_0_ , \g56485/_0_ , \g56486/_0_ , \g56487/_0_ , \g56488/_0_ , \g56489/_0_ , \g56490/_0_ , \g56491/_0_ , \g56492/_0_ , \g56507/_0_ , \g56543/_0_ , \g56544/_0_ , \g56545/_0_ , \g56546/_0_ , \g56547/_0_ , \g56548/_0_ , \g56549/_0_ , \g56551/_0_ , \g56567/_0_ , \g56602/_0_ , \g56603/_0_ , \g56604/_0_ , \g56605/_0_ , \g56606/_0_ , \g56607/_0_ , \g56608/_0_ , \g56610/_0_ , \g56627/_0_ , \g56661/_0_ , \g56662/_0_ , \g56663/_0_ , \g56664/_0_ , \g56665/_0_ , \g56666/_0_ , \g56667/_0_ , \g56668/_0_ , \g56686/_0_ , \g56720/_0_ , \g56721/_0_ , \g56722/_0_ , \g56723/_0_ , \g56724/_0_ , \g56725/_0_ , \g56726/_0_ , \g56727/_0_ , \g56728/_0_ , \g56745/_0_ , \g56779/_0_ , \g56780/_0_ , \g56781/_0_ , \g56782/_0_ , \g56783/_0_ , \g56784/_0_ , \g56785/_0_ , \g56804/_0_ , \g56838/_0_ , \g56839/_0_ , \g56840/_0_ , \g56841/_0_ , \g56842/_0_ , \g56843/_0_ , \g56844/_0_ , \g56845/_0_ , \g56846/_0_ , \g56863/_0_ , \g56897/_0_ , \g56898/_0_ , \g56899/_0_ , \g56900/_0_ , \g56901/_0_ , \g56902/_0_ , \g56903/_0_ , \g56905/_0_ , \g56921/_0_ , \g56956/_0_ , \g56957/_0_ , \g56958/_0_ , \g56959/_0_ , \g56960/_0_ , \g56961/_0_ , \g56962/_0_ , \g56964/_0_ , \g56980/_0_ , \g57015/_0_ , \g57016/_0_ , \g57017/_0_ , \g57018/_0_ , \g57019/_0_ , \g57020/_0_ , \g57021/_0_ , \g57023/_0_ , \g57040/_0_ , \g57074/_0_ , \g57075/_0_ , \g57076/_0_ , \g57077/_0_ , \g57078/_0_ , \g57079/_0_ , \g57080/_0_ , \g57081/_0_ , \g57099/_0_ , \g57133/_0_ , \g57134/_0_ , \g57135/_0_ , \g57136/_0_ , \g57137/_0_ , \g57138/_0_ , \g57139/_0_ , \g57140/_0_ , \g57141/_0_ , \g57159/_0_ , \g57193/_0_ , \g57195/_0_ , \g57196/_0_ , \g57197/_0_ , \g57198/_0_ , \g57199/_0_ , \g57200/_0_ , \g57202/_0_ , \g57219/_0_ , \g57254/_0_ , \g57255/_0_ , \g57256/_0_ , \g57257/_0_ , \g57258/_0_ , \g57259/_0_ , \g57260/_0_ , \g57262/_0_ , \g57263/_0_ , \g57285/_0_ , \g57318/_0_ , \g57319/_0_ , \g57320/_0_ , \g57321/_0_ , \g57322/_0_ , \g57323/_0_ , \g57324/_0_ , \g57325/_0_ , \g57326/_0_ , \g57328/_0_ , \g57329/_0_ , \g57330/_0_ , \g57350/_0_ , \g57387/_0_ , \g57388/_0_ , \g57390/_0_ , \g57391/_0_ , \g57392/_0_ , \g57393/_0_ , \g57395/_0_ , \g57396/_0_ , \g57439/_0_ , \g57476/_0_ , \g57477/_0_ , \g57478/_0_ , \g57479/_0_ , \g57480/_0_ , \g57481/_0_ , \g57482/_0_ , \g57483/_0_ , \g57484/_0_ , \g57485/_0_ , \g57486/_0_ , \g57487/_0_ , \g57488/_0_ , \g57489/_0_ , \g57490/_0_ , \g57491/_0_ , \g57492/_0_ , \g57493/_0_ , \g57494/_0_ , \g57495/_0_ , \g57496/_0_ , \g57497/_0_ , \g57498/_0_ , \g57499/_0_ , \g57500/_0_ , \g57501/_0_ , \g57502/_0_ , \g57503/_0_ , \g57504/_0_ , \g57505/_0_ , \g57524/_0_ , \g57537/_0_ , \g57541/_0_ , \g57543/_0_ , \g58163/_0_ , \g58572/_0_ , \g58573/_0_ , \g58574/_0_ , \g58575/_0_ , \g58576/_0_ , \g58577/_0_ , \g58578/_0_ , \g58579/_0_ , \g58580/_0_ , \g58581/_0_ , \g58582/_0_ , \g58583/_0_ , \g58584/_0_ , \g58585/_0_ , \g58586/_0_ , \g58587/_0_ , \g58588/_0_ , \g58589/_0_ , \g58590/_0_ , \g58591/_0_ , \g58592/_0_ , \g58593/_0_ , \g58594/_0_ , \g58595/_0_ , \g58596/_0_ , \g58597/_0_ , \g58598/_0_ , \g58600/_0_ , \g58602/_0_ , \g58604/_0_ , \g58615/_0_ , \g59240/_0_ , \g59241/_0_ , \g59242/_0_ , \g59243/_0_ , \g59244/_0_ , \g59245/_0_ , \g59246/_0_ , \g59247/_0_ , \g59248/_0_ , \g59249/_0_ , \g59250/_0_ , \g59251/_0_ , \g59252/_0_ , \g59253/_0_ , \g59254/_0_ , \g59255/_0_ , \g59256/_0_ , \g59257/_0_ , \g59258/_0_ , \g59259/_0_ , \g59260/_0_ , \g59261/_0_ , \g59262/_0_ , \g59263/_0_ , \g59264/_0_ , \g59265/_0_ , \g59266/_0_ , \g59267/_0_ , \g59268/_0_ , \g59269/_0_ , \g59270/_0_ , \g59271/_0_ , \g59272/_0_ , \g59273/_0_ , \g59274/_0_ , \g59275/_0_ , \g59276/_0_ , \g59277/_0_ , \g59278/_0_ , \g59279/_0_ , \g59280/_0_ , \g59281/_0_ , \g59282/_0_ , \g59283/_0_ , \g59284/_0_ , \g59285/_0_ , \g59286/_0_ , \g59287/_0_ , \g59288/_0_ , \g59289/_0_ , \g59290/_0_ , \g59291/_0_ , \g59292/_0_ , \g59293/_0_ , \g59294/_0_ , \g59295/_0_ , \g59296/_0_ , \g59297/_0_ , \g59298/_0_ , \g59299/_0_ , \g59300/_0_ , \g59301/_0_ , \g59302/_0_ , \g59303/_0_ , \g59304/_0_ , \g59305/_0_ , \g59306/_0_ , \g59307/_0_ , \g59308/_0_ , \g59309/_0_ , \g59310/_0_ , \g59311/_0_ , \g59312/_0_ , \g59313/_0_ , \g59314/_0_ , \g59315/_0_ , \g59316/_0_ , \g59317/_0_ , \g59318/_0_ , \g59319/_0_ , \g59320/_0_ , \g59321/_0_ , \g59322/_0_ , \g59323/_0_ , \g59324/_0_ , \g59325/_0_ , \g59326/_0_ , \g59327/_0_ , \g59328/_0_ , \g59329/_0_ , \g59330/_0_ , \g59331/_0_ , \g59332/_0_ , \g59333/_0_ , \g59334/_0_ , \g59335/_0_ , \g59336/_0_ , \g59337/_0_ , \g59338/_0_ , \g59339/_0_ , \g59340/_0_ , \g59341/_0_ , \g59342/_0_ , \g59343/_0_ , \g59344/_0_ , \g59345/_0_ , \g59346/_0_ , \g59347/_0_ , \g59348/_0_ , \g59349/_0_ , \g59350/_0_ , \g59351/_0_ , \g59352/_0_ , \g59353/_0_ , \g59354/_0_ , \g59355/_0_ , \g59356/_0_ , \g59357/_0_ , \g59358/_0_ , \g59359/_0_ , \g59360/_0_ , \g59361/_0_ , \g59362/_0_ , \g59363/_0_ , \g59364/_0_ , \g59365/_0_ , \g59366/_0_ , \g59367/_0_ , \g59368/_0_ , \g59369/_0_ , \g59370/_0_ , \g59371/_0_ , \g59372/_0_ , \g59373/_0_ , \g59374/_0_ , \g59375/_0_ , \g59376/_0_ , \g59377/_0_ , \g59378/_0_ , \g59379/_0_ , \g59380/_0_ , \g59381/_0_ , \g59382/_0_ , \g59383/_0_ , \g59384/_0_ , \g59385/_0_ , \g59386/_0_ , \g59387/_0_ , \g59388/_0_ , \g59389/_0_ , \g59390/_0_ , \g59391/_0_ , \g59392/_0_ , \g59393/_0_ , \g59394/_0_ , \g59395/_0_ , \g59396/_0_ , \g59397/_0_ , \g59398/_0_ , \g59399/_0_ , \g59400/_0_ , \g59401/_0_ , \g59402/_0_ , \g59403/_0_ , \g59404/_0_ , \g59405/_0_ , \g59406/_0_ , \g59407/_0_ , \g59408/_0_ , \g59409/_0_ , \g59410/_0_ , \g59411/_0_ , \g59412/_0_ , \g59413/_0_ , \g59414/_0_ , \g59415/_0_ , \g59416/_0_ , \g59417/_0_ , \g59418/_0_ , \g59419/_0_ , \g59420/_0_ , \g59421/_0_ , \g59422/_0_ , \g59423/_0_ , \g59424/_0_ , \g59425/_0_ , \g59426/_0_ , \g59427/_0_ , \g59428/_0_ , \g59429/_0_ , \g59430/_0_ , \g59431/_0_ , \g59432/_0_ , \g59433/_0_ , \g59434/_0_ , \g59435/_0_ , \g59436/_0_ , \g59437/_0_ , \g59438/_0_ , \g59439/_0_ , \g59440/_0_ , \g59441/_0_ , \g59442/_0_ , \g59443/_0_ , \g59444/_0_ , \g59445/_0_ , \g59446/_0_ , \g59447/_0_ , \g59448/_0_ , \g59449/_0_ , \g59450/_0_ , \g59451/_0_ , \g59452/_0_ , \g59453/_0_ , \g59454/_0_ , \g59455/_0_ , \g59456/_0_ , \g59457/_0_ , \g59458/_0_ , \g59459/_0_ , \g59460/_0_ , \g59461/_0_ , \g59462/_0_ , \g59463/_0_ , \g59464/_0_ , \g59465/_0_ , \g59466/_0_ , \g59467/_0_ , \g59468/_0_ , \g59469/_0_ , \g59470/_0_ , \g59471/_0_ , \g59472/_0_ , \g59473/_0_ , \g59474/_0_ , \g59475/_0_ , \g59476/_0_ , \g59477/_0_ , \g59478/_0_ , \g59479/_0_ , \g59480/_0_ , \g59481/_0_ , \g59482/_0_ , \g59483/_0_ , \g59484/_0_ , \g59485/_0_ , \g59486/_0_ , \g59487/_0_ , \g59488/_0_ , \g59489/_0_ , \g59490/_0_ , \g59491/_0_ , \g59492/_0_ , \g59493/_0_ , \g59494/_0_ , \g59495/_0_ , \g59496/_0_ , \g59497/_0_ , \g59498/_0_ , \g59500/_0_ , \g59503/_0_ , \g59512/_0_ , \g61336/_0_ , \g61521/_0_ , \g61523/_0_ , \g61524/_0_ , \g61526/_0_ , \g61527/_0_ , \g61528/_0_ , \g61529/_0_ , \g61530/_0_ , \g61531/_0_ , \g61532/_0_ , \g61533/_0_ , \g61535/_0_ , \g61537/_0_ , \g61539/_0_ , \g61540/_0_ , \g61541/_0_ , \g61542/_0_ , \g61546/_0_ , \g61550/_0_ , \g61551/_0_ , \g61552/_0_ , \g61554/_0_ , \g61555/_0_ , \g61556/_0_ , \g61558/_0_ , \g61559/_0_ , \g61561/_0_ , \g61562/_0_ , \g61563/_0_ , \g61564/_0_ , \g61565/_0_ , \g61566/_0_ , \g61568/_0_ , \g61570/_0_ , \g61571/_0_ , \g61572/_0_ , \g61573/_0_ , \g61577/_0_ , \g61578/_0_ , \g61579/_0_ , \g61580/_0_ , \g61581/_0_ , \g61582/_0_ , \g61583/_0_ , \g61584/_0_ , \g61585/_0_ , \g61586/_0_ , \g61587/_0_ , \g61588/_0_ , \g61589/_0_ , \g61591/_0_ , \g61592/_0_ , \g61594/_0_ , \g61595/_0_ , \g61596/_0_ , \g61597/_0_ , \g61598/_0_ , \g61599/_0_ , \g61600/_0_ , \g61601/_0_ , \g61605/_0_ , \g61606/_0_ , \g61607/_0_ , \g61608/_0_ , \g61609/_0_ , \g61610/_0_ , \g61611/_0_ , \g61612/_0_ , \g61613/_0_ , \g61615/_0_ , \g61616/_0_ , \g61617/_0_ , \g61618/_0_ , \g61619/_0_ , \g61620/_0_ , \g61621/_0_ , \g61623/_0_ , \g61624/_0_ , \g61625/_0_ , \g61626/_0_ , \g61627/_0_ , \g61629/_0_ , \g61630/_0_ , \g61631/_0_ , \g61632/_0_ , \g61633/_0_ , \g61634/_0_ , \g61636/_0_ , \g61638/_0_ , \g61639/_0_ , \g61640/_0_ , \g61641/_0_ , \g61642/_0_ , \g61644/_0_ , \g61647/_0_ , \g61648/_0_ , \g61649/_0_ , \g61650/_0_ , \g61653/_0_ , \g61654/_0_ , \g61655/_0_ , \g61656/_0_ , \g61658/_0_ , \g61661/_0_ , \g61662/_0_ , \g61663/_0_ , \g61664/_0_ , \g61666/_0_ , \g61667/_0_ , \g61668/_0_ , \g61670/_0_ , \g61671/_0_ , \g61672/_0_ , \g61673/_0_ , \g61675/_0_ , \g61676/_0_ , \g61680/_0_ , \g61681/_0_ , \g61682/_0_ , \g61683/_0_ , \g61684/_0_ , \g61686/_0_ , \g61687/_0_ , \g61688/_0_ , \g61689/_0_ , \g61690/_0_ , \g61691/_0_ , \g61693/_0_ , \g61694/_0_ , \g61696/_0_ , \g61697/_0_ , \g61698/_0_ , \g61699/_0_ , \g61700/_0_ , \g61701/_0_ , \g61702/_0_ , \g61703/_0_ , \g61704/_0_ , \g61705/_0_ , \g61706/_0_ , \g61707/_0_ , \g61708/_0_ , \g61711/_0_ , \g61712/_0_ , \g61714/_0_ , \g61716/_0_ , \g61717/_0_ , \g61719/_0_ , \g61720/_0_ , \g61721/_0_ , \g61724/_0_ , \g61725/_0_ , \g61728/_0_ , \g61729/_0_ , \g61731/_0_ , \g61732/_0_ , \g61733/_0_ , \g61736/_0_ , \g61737/_0_ , \g61739/_0_ , \g61740/_0_ , \g61741/_0_ , \g61743/_0_ , \g61744/_0_ , \g61745/_0_ , \g61746/_0_ , \g61747/_0_ , \g61748/_0_ , \g61749/_0_ , \g61750/_0_ , \g61751/_0_ , \g61752/_0_ , \g61753/_0_ , \g61754/_0_ , \g61755/_0_ , \g61757/_0_ , \g61758/_0_ , \g61759/_0_ , \g61760/_0_ , \g61761/_0_ , \g61762/_0_ , \g61763/_0_ , \g61764/_0_ , \g61765/_0_ , \g61766/_0_ , \g61767/_0_ , \g61768/_0_ , \g61769/_0_ , \g61770/_0_ , \g61771/_0_ , \g61772/_0_ , \g61773/_0_ , \g61774/_0_ , \g61775/_0_ , \g61776/_0_ , \g61777/_0_ , \g61778/_0_ , \g61780/_0_ , \g61781/_0_ , \g61783/_0_ , \g61784/_0_ , \g61786/_0_ , \g61787/_0_ , \g61790/_0_ , \g61791/_0_ , \g61794/_0_ , \g61795/_0_ , \g61796/_0_ , \g61797/_0_ , \g61798/_0_ , \g61799/_0_ , \g61800/_0_ , \g61801/_0_ , \g61802/_0_ , \g61803/_0_ , \g61805/_0_ , \g61806/_0_ , \g61807/_0_ , \g61808/_0_ , \g61809/_0_ , \g61810/_0_ , \g61811/_0_ , \g61812/_0_ , \g61813/_0_ , \g61816/_0_ , \g61817/_0_ , \g61818/_0_ , \g61820/_0_ , \g61822/_0_ , \g61823/_0_ , \g61825/_0_ , \g61826/_0_ , \g61827/_0_ , \g61828/_0_ , \g61829/_0_ , \g61832/_0_ , \g61834/_0_ , \g61835/_0_ , \g61837/_0_ , \g61838/_0_ , \g61839/_0_ , \g61840/_0_ , \g61844/_0_ , \g61847/_0_ , \g61848/_0_ , \g61849/_0_ , \g61850/_0_ , \g61851/_0_ , \g61853/_0_ , \g61854/_0_ , \g61855/_0_ , \g61856/_0_ , \g61858/_0_ , \g61859/_0_ , \g61861/_0_ , \g61862/_0_ , \g61863/_0_ , \g61864/_0_ , \g61865/_0_ , \g61866/_0_ , \g61867/_0_ , \g61868/_0_ , \g61869/_0_ , \g61870/_0_ , \g61871/_0_ , \g61873/_0_ , \g61874/_0_ , \g61875/_0_ , \g61877/_0_ , \g61878/_0_ , \g61879/_0_ , \g61880/_0_ , \g61881/_0_ , \g61883/_0_ , \g61884/_0_ , \g61886/_0_ , \g61887/_0_ , \g61890/_0_ , \g61891/_0_ , \g61892/_0_ , \g61893/_0_ , \g61894/_0_ , \g61895/_0_ , \g61900/_0_ , \g61901/_0_ , \g61902/_0_ , \g61904/_0_ , \g61905/_0_ , \g61906/_0_ , \g61907/_0_ , \g61914/_0_ , \g61915/_0_ , \g61917/_0_ , \g61919/_0_ , \g61921/_0_ , \g61924/_0_ , \g61925/_0_ , \g61926/_0_ , \g61927/_0_ , \g61928/_0_ , \g61929/_0_ , \g61930/_0_ , \g61931/_0_ , \g61932/_0_ , \g61933/_0_ , \g61934/_0_ , \g61935/_0_ , \g61936/_0_ , \g61937/_0_ , \g61938/_0_ , \g61939/_0_ , \g61943/_0_ , \g61944/_0_ , \g61945/_0_ , \g61947/_0_ , \g61948/_0_ , \g61949/_0_ , \g61950/_0_ , \g61951/_0_ , \g61952/_0_ , \g61953/_0_ , \g61955/_0_ , \g61956/_0_ , \g61957/_0_ , \g61958/_0_ , \g61959/_0_ , \g61960/_0_ , \g61961/_0_ , \g61962/_0_ , \g61963/_0_ , \g61964/_0_ , \g61965/_0_ , \g61966/_0_ , \g61967/_0_ , \g61968/_0_ , \g61969/_0_ , \g61970/_0_ , \g61971/_0_ , \g61972/_0_ , \g61973/_0_ , \g61974/_0_ , \g61976/_0_ , \g61978/_0_ , \g61980/_0_ , \g61981/_0_ , \g61982/_0_ , \g61983/_0_ , \g61984/_0_ , \g61985/_0_ , \g61986/_0_ , \g61987/_0_ , \g61988/_0_ , \g61989/_0_ , \g61990/_0_ , \g61992/_0_ , \g61994/_0_ , \g61995/_0_ , \g61996/_0_ , \g61997/_0_ , \g61998/_0_ , \g62000/_0_ , \g62001/_0_ , \g62002/_0_ , \g62003/_0_ , \g62004/_0_ , \g62005/_0_ , \g62007/_0_ , \g62008/_0_ , \g62009/_0_ , \g62010/_0_ , \g62011/_0_ , \g62012/_0_ , \g62013/_0_ , \g62014/_0_ , \g62015/_0_ , \g62016/_0_ , \g62017/_0_ , \g62018/_0_ , \g62019/_0_ , \g62020/_0_ , \g62021/_0_ , \g62022/_0_ , \g62023/_0_ , \g62024/_0_ , \g62025/_0_ , \g62026/_0_ , \g62027/_0_ , \g62030/_0_ , \g62033/_0_ , \g62034/_0_ , \g62036/_0_ , \g62038/_0_ , \g62041/_0_ , \g62042/_0_ , \g62043/_0_ , \g62044/_0_ , \g62045/_0_ , \g62046/_0_ , \g62047/_0_ , \g62048/_0_ , \g62050/_0_ , \g62051/_0_ , \g62052/_0_ , \g62055/_0_ , \g62057/_0_ , \g62058/_0_ , \g62059/_0_ , \g62060/_0_ , \g62061/_0_ , \g62062/_0_ , \g62064/_0_ , \g62065/_0_ , \g62066/_0_ , \g62067/_0_ , \g62068/_0_ , \g62072/_0_ , \g62073/_0_ , \g62074/_0_ , \g62075/_0_ , \g62076/_0_ , \g62077/_0_ , \g62078/_0_ , \g62080/_0_ , \g62081/_0_ , \g62082/_0_ , \g62084/_0_ , \g62085/_0_ , \g62086/_0_ , \g62087/_0_ , \g62088/_0_ , \g62089/_0_ , \g62090/_0_ , \g62091/_0_ , \g62092/_0_ , \g62094/_0_ , \g62096/_0_ , \g62097/_0_ , \g62098/_0_ , \g62099/_0_ , \g62100/_0_ , \g62101/_0_ , \g62102/_0_ , \g62104/_0_ , \g62106/_0_ , \g62107/_0_ , \g62108/_0_ , \g62110/_0_ , \g62112/_0_ , \g62113/_0_ , \g62114/_0_ , \g62116/_0_ , \g62117/_0_ , \g62118/_0_ , \g62119/_0_ , \g62120/_0_ , \g62121/_0_ , \g62122/_0_ , \g62124/_0_ , \g62126/_0_ , \g62127/_0_ , \g62128/_0_ , \g62129/_0_ , \g62130/_0_ , \g62131/_0_ , \g62132/_0_ , \g62133/_0_ , \g62135/_0_ , \g62136/_0_ , \g62137/_0_ , \g62138/_0_ , \g62140/_0_ , \g62143/_0_ , \g62144/_0_ , \g62149/_0_ , \g62150/_0_ , \g62151/_0_ , \g62153/_0_ , \g62155/_0_ , \g62156/_0_ , \g62158/_0_ , \g62160/_0_ , \g62161/_0_ , \g62162/_0_ , \g62164/_0_ , \g62165/_0_ , \g62166/_0_ , \g62167/_0_ , \g62168/_0_ , \g62169/_0_ , \g62172/_0_ , \g62173/_0_ , \g62175/_0_ , \g62176/_0_ , \g62177/_0_ , \g62178/_0_ , \g62179/_0_ , \g62180/_0_ , \g62181/_0_ , \g62182/_0_ , \g62183/_0_ , \g62184/_0_ , \g62185/_0_ , \g62186/_0_ , \g62188/_0_ , \g62189/_0_ , \g62190/_0_ , \g62191/_0_ , \g62193/_0_ , \g62194/_0_ , \g62195/_0_ , \g62196/_0_ , \g62197/_0_ , \g62200/_0_ , \g62201/_0_ , \g62202/_0_ , \g62203/_0_ , \g62205/_0_ , \g62206/_0_ , \g62207/_0_ , \g62208/_0_ , \g62209/_0_ , \g62210/_0_ , \g62211/_0_ , \g62215/_0_ , \g62218/_0_ , \g62219/_0_ , \g62221/_0_ , \g62222/_0_ , \g62223/_0_ , \g62224/_0_ , \g62225/_0_ , \g62226/_0_ , \g62229/_0_ , \g62230/_0_ , \g62231/_0_ , \g62233/_0_ , \g62236/_0_ , \g62237/_0_ , \g62238/_0_ , \g62240/_0_ , \g62241/_0_ , \g62243/_0_ , \g62244/_0_ , \g62245/_0_ , \g62247/_0_ , \g62248/_0_ , \g62250/_0_ , \g62252/_0_ , \g62253/_0_ , \g62255/_0_ , \g62256/_0_ , \g62257/_0_ , \g62258/_0_ , \g62259/_0_ , \g62260/_0_ , \g62261/_0_ , \g62262/_0_ , \g62263/_0_ , \g62264/_0_ , \g62265/_0_ , \g62267/_0_ , \g62269/_0_ , \g62270/_0_ , \g62272/_0_ , \g62274/_0_ , \g62277/_0_ , \g62279/_0_ , \g62280/_0_ , \g62281/_0_ , \g62283/_0_ , \g62284/_0_ , \g62285/_0_ , \g62286/_0_ , \g62288/_0_ , \g62289/_0_ , \g62290/_0_ , \g62294/_0_ , \g62295/_0_ , \g62296/_0_ , \g62297/_0_ , \g62298/_0_ , \g62299/_0_ , \g62303/_0_ , \g62305/_0_ , \g62306/_0_ , \g62307/_0_ , \g62309/_0_ , \g62311/_0_ , \g62312/_0_ , \g62313/_0_ , \g62314/_0_ , \g62315/_0_ , \g62316/_0_ , \g62317/_0_ , \g62318/_0_ , \g62319/_0_ , \g62320/_0_ , \g62322/_0_ , \g62324/_0_ , \g62325/_0_ , \g62326/_0_ , \g62327/_0_ , \g62329/_0_ , \g62330/_0_ , \g62331/_0_ , \g62332/_0_ , \g62333/_0_ , \g62335/_0_ , \g62336/_0_ , \g62338/_0_ , \g62341/_0_ , \g62342/_0_ , \g62344/_0_ , \g62345/_0_ , \g62348/_0_ , \g62349/_0_ , \g62350/_0_ , \g62353/_0_ , \g62354/_0_ , \g62355/_0_ , \g62356/_0_ , \g62359/_0_ , \g62362/_0_ , \g62363/_0_ , \g62364/_0_ , \g62365/_0_ , \g62366/_0_ , \g62367/_0_ , \g62368/_0_ , \g62369/_0_ , \g62370/_0_ , \g62371/_0_ , \g62372/_0_ , \g62373/_0_ , \g62374/_0_ , \g62376/_0_ , \g62467/_0_ , \g62468/_0_ , \g62469/_0_ , \g62470/_0_ , \g62471/_0_ , \g62472/_0_ , \g62473/_0_ , \g62474/_0_ , \g62475/_0_ , \g62478/_0_ , \g62480/_0_ , \g62481/_0_ , \g62482/_0_ , \g62483/_0_ , \g62484/_0_ , \g62485/_0_ , \g62486/_0_ , \g62487/_0_ , \g62488/_0_ , \g62489/_0_ , \g62490/_0_ , \g62491/_0_ , \g62492/_0_ , \g62493/_0_ , \g62494/_0_ , \g62495/_0_ , \g62496/_0_ , \g62497/_0_ , \g62498/_0_ , \g62499/_0_ , \g62500/_0_ , \g62501/_0_ , \g62502/_0_ , \g62503/_0_ , \g62504/_0_ , \g62509/_0_ , \g62510/_0_ , \g62511/_0_ , \g62512/_0_ , \g62513/_0_ , \g62514/_0_ , \g62515/_0_ , \g62516/_0_ , \g62517/_0_ , \g62518/_0_ , \g62519/_0_ , \g62520/_0_ , \g62521/_0_ , \g62523/_0_ , \g62526/_0_ , \g62528/_0_ , \g62529/_0_ , \g62531/_0_ , \g62532/_0_ , \g62533/_0_ , \g62534/_0_ , \g62535/_0_ , \g62536/_0_ , \g62537/_0_ , \g62539/_0_ , \g62540/_0_ , \g62541/_0_ , \g62542/_0_ , \g62543/_0_ , \g62544/_0_ , \g62545/_0_ , \g62547/_0_ , \g62548/_0_ , \g62549/_0_ , \g62550/_0_ , \g62551/_0_ , \g62552/_0_ , \g62553/_0_ , \g62554/_0_ , \g62555/_0_ , \g62556/_0_ , \g62557/_0_ , \g62560/_0_ , \g62562/_0_ , \g62563/_0_ , \g62564/_0_ , \g62565/_0_ , \g62566/_0_ , \g62567/_0_ , \g62569/_0_ , \g62570/_0_ , \g62571/_0_ , \g62572/_0_ , \g62573/_0_ , \g62574/_0_ , \g62576/_0_ , \g62577/_0_ , \g62581/_0_ , \g62582/_0_ , \g62584/_0_ , \g62585/_0_ , \g62586/_0_ , \g62588/_0_ , \g62589/_0_ , \g62593/_0_ , \g62594/_0_ , \g62595/_0_ , \g62596/_0_ , \g62597/_0_ , \g62598/_0_ , \g62599/_0_ , \g62600/_0_ , \g62601/_0_ , \g62602/_0_ , \g62603/_0_ , \g62604/_0_ , \g62605/_0_ , \g62606/_0_ , \g62607/_0_ , \g62608/_0_ , \g62609/_0_ , \g62610/_0_ , \g62612/_0_ , \g62613/_0_ , \g62614/_0_ , \g62615/_0_ , \g62617/_0_ , \g62618/_0_ , \g62620/_0_ , \g62621/_0_ , \g62622/_0_ , \g62624/_0_ , \g62625/_0_ , \g62626/_0_ , \g62627/_0_ , \g62629/_0_ , \g62630/_0_ , \g62632/_0_ , \g62633/_0_ , \g62635/_0_ , \g62636/_0_ , \g62637/_0_ , \g62638/_0_ , \g62640/_0_ , \g62641/_0_ , \g62642/_0_ , \g62643/_0_ , \g62644/_0_ , \g62646/_0_ , \g62647/_0_ , \g62649/_0_ , \g62650/_0_ , \g62651/_0_ , \g62653/_0_ , \g62655/_0_ , \g62656/_0_ , \g62657/_0_ , \g62658/_0_ , \g62660/_0_ , \g62661/_0_ , \g62662/_0_ , \g62663/_0_ , \g62664/_0_ , \g62665/_0_ , \g62667/_0_ , \g62669/_0_ , \g62670/_0_ , \g62671/_0_ , \g62672/_0_ , \g62674/_0_ , \g62675/_0_ , \g62676/_0_ , \g62677/_0_ , \g62678/_0_ , \g62679/_0_ , \g62680/_0_ , \g62681/_0_ , \g62682/_0_ , \g62684/_0_ , \g62685/_0_ , \g62686/_0_ , \g62687/_0_ , \g62690/_0_ , \g62693/_0_ , \g62698/_0_ , \g62699/_0_ , \g62700/_0_ , \g62701/_0_ , \g62702/_0_ , \g62703/_0_ , \g62704/_0_ , \g62709/_0_ , \g62710/_0_ , \g62711/_0_ , \g62714/_0_ , \g62715/_0_ , \g62717/_0_ , \g62718/_0_ , \g62719/_0_ , \g62720/_0_ , \g62721/_0_ , \g62723/_0_ , \g62725/_0_ , \g62726/_0_ , \g62729/_0_ , \g62731/_0_ , \g62733/_0_ , \g62738/_0_ , \g62741/_0_ , \g62742/_0_ , \g62744/_0_ , \g62745/_0_ , \g62746/_0_ , \g62747/_0_ , \g62748/_0_ , \g62749/_0_ , \g62753/_0_ , \g62755/_0_ , \g62756/_0_ , \g62758/_0_ , \g62759/_0_ , \g62760/_0_ , \g62761/_0_ , \g62763/_0_ , \g62766/_0_ , \g62767/_0_ , \g62768/_0_ , \g65554/_0_ , \g65561/_0_ , \g65569/_0_ , \g65580/_0_ , \g65599/_0_ , \g65606/_0_ , \g65636/_0_ , \g65864/_0_ );
	input \DATA_0_0_pad  ;
	input \DATA_0_10_pad  ;
	input \DATA_0_11_pad  ;
	input \DATA_0_12_pad  ;
	input \DATA_0_13_pad  ;
	input \DATA_0_14_pad  ;
	input \DATA_0_15_pad  ;
	input \DATA_0_16_pad  ;
	input \DATA_0_17_pad  ;
	input \DATA_0_18_pad  ;
	input \DATA_0_19_pad  ;
	input \DATA_0_1_pad  ;
	input \DATA_0_20_pad  ;
	input \DATA_0_21_pad  ;
	input \DATA_0_22_pad  ;
	input \DATA_0_23_pad  ;
	input \DATA_0_24_pad  ;
	input \DATA_0_25_pad  ;
	input \DATA_0_26_pad  ;
	input \DATA_0_27_pad  ;
	input \DATA_0_28_pad  ;
	input \DATA_0_29_pad  ;
	input \DATA_0_2_pad  ;
	input \DATA_0_30_pad  ;
	input \DATA_0_31_pad  ;
	input \DATA_0_3_pad  ;
	input \DATA_0_4_pad  ;
	input \DATA_0_5_pad  ;
	input \DATA_0_6_pad  ;
	input \DATA_0_7_pad  ;
	input \DATA_0_8_pad  ;
	input \DATA_0_9_pad  ;
	input RESET_pad ;
	input \TM0_pad  ;
	input \TM1_pad  ;
	input \WX10829_reg/NET0131  ;
	input \WX10831_reg/NET0131  ;
	input \WX10833_reg/NET0131  ;
	input \WX10835_reg/NET0131  ;
	input \WX10837_reg/NET0131  ;
	input \WX10839_reg/NET0131  ;
	input \WX10841_reg/NET0131  ;
	input \WX10843_reg/NET0131  ;
	input \WX10845_reg/NET0131  ;
	input \WX10847_reg/NET0131  ;
	input \WX10849_reg/NET0131  ;
	input \WX10851_reg/NET0131  ;
	input \WX10853_reg/NET0131  ;
	input \WX10855_reg/NET0131  ;
	input \WX10857_reg/NET0131  ;
	input \WX10859_reg/NET0131  ;
	input \WX10861_reg/NET0131  ;
	input \WX10863_reg/NET0131  ;
	input \WX10865_reg/NET0131  ;
	input \WX10867_reg/NET0131  ;
	input \WX10869_reg/NET0131  ;
	input \WX10871_reg/NET0131  ;
	input \WX10873_reg/NET0131  ;
	input \WX10875_reg/NET0131  ;
	input \WX10877_reg/NET0131  ;
	input \WX10879_reg/NET0131  ;
	input \WX10881_reg/NET0131  ;
	input \WX10883_reg/NET0131  ;
	input \WX10885_reg/NET0131  ;
	input \WX10887_reg/NET0131  ;
	input \WX10889_reg/NET0131  ;
	input \WX10891_reg/NET0131  ;
	input \WX10989_reg/NET0131  ;
	input \WX10991_reg/NET0131  ;
	input \WX10993_reg/NET0131  ;
	input \WX10995_reg/NET0131  ;
	input \WX10997_reg/NET0131  ;
	input \WX10999_reg/NET0131  ;
	input \WX11001_reg/NET0131  ;
	input \WX11003_reg/NET0131  ;
	input \WX11005_reg/NET0131  ;
	input \WX11007_reg/NET0131  ;
	input \WX11009_reg/NET0131  ;
	input \WX11011_reg/NET0131  ;
	input \WX11013_reg/NET0131  ;
	input \WX11015_reg/NET0131  ;
	input \WX11017_reg/NET0131  ;
	input \WX11019_reg/NET0131  ;
	input \WX11021_reg/NET0131  ;
	input \WX11023_reg/NET0131  ;
	input \WX11025_reg/NET0131  ;
	input \WX11027_reg/NET0131  ;
	input \WX11029_reg/NET0131  ;
	input \WX11031_reg/NET0131  ;
	input \WX11033_reg/NET0131  ;
	input \WX11035_reg/NET0131  ;
	input \WX11037_reg/NET0131  ;
	input \WX11039_reg/NET0131  ;
	input \WX11041_reg/NET0131  ;
	input \WX11043_reg/NET0131  ;
	input \WX11045_reg/NET0131  ;
	input \WX11047_reg/NET0131  ;
	input \WX11049_reg/NET0131  ;
	input \WX11051_reg/NET0131  ;
	input \WX11053_reg/NET0131  ;
	input \WX11055_reg/NET0131  ;
	input \WX11057_reg/NET0131  ;
	input \WX11059_reg/NET0131  ;
	input \WX11061_reg/NET0131  ;
	input \WX11063_reg/NET0131  ;
	input \WX11065_reg/NET0131  ;
	input \WX11067_reg/NET0131  ;
	input \WX11069_reg/NET0131  ;
	input \WX11071_reg/NET0131  ;
	input \WX11073_reg/NET0131  ;
	input \WX11075_reg/NET0131  ;
	input \WX11077_reg/NET0131  ;
	input \WX11079_reg/NET0131  ;
	input \WX11081_reg/NET0131  ;
	input \WX11083_reg/NET0131  ;
	input \WX11085_reg/NET0131  ;
	input \WX11087_reg/NET0131  ;
	input \WX11089_reg/NET0131  ;
	input \WX11091_reg/NET0131  ;
	input \WX11093_reg/NET0131  ;
	input \WX11095_reg/NET0131  ;
	input \WX11097_reg/NET0131  ;
	input \WX11099_reg/NET0131  ;
	input \WX11101_reg/NET0131  ;
	input \WX11103_reg/NET0131  ;
	input \WX11105_reg/NET0131  ;
	input \WX11107_reg/NET0131  ;
	input \WX11109_reg/NET0131  ;
	input \WX11111_reg/NET0131  ;
	input \WX11113_reg/NET0131  ;
	input \WX11115_reg/NET0131  ;
	input \WX11117_reg/NET0131  ;
	input \WX11119_reg/NET0131  ;
	input \WX11121_reg/NET0131  ;
	input \WX11123_reg/NET0131  ;
	input \WX11125_reg/NET0131  ;
	input \WX11127_reg/NET0131  ;
	input \WX11129_reg/NET0131  ;
	input \WX11131_reg/NET0131  ;
	input \WX11133_reg/NET0131  ;
	input \WX11135_reg/NET0131  ;
	input \WX11137_reg/NET0131  ;
	input \WX11139_reg/NET0131  ;
	input \WX11141_reg/NET0131  ;
	input \WX11143_reg/NET0131  ;
	input \WX11145_reg/NET0131  ;
	input \WX11147_reg/NET0131  ;
	input \WX11149_reg/NET0131  ;
	input \WX11151_reg/NET0131  ;
	input \WX11153_reg/NET0131  ;
	input \WX11155_reg/NET0131  ;
	input \WX11157_reg/NET0131  ;
	input \WX11159_reg/NET0131  ;
	input \WX11161_reg/NET0131  ;
	input \WX11163_reg/NET0131  ;
	input \WX11165_reg/NET0131  ;
	input \WX11167_reg/NET0131  ;
	input \WX11169_reg/NET0131  ;
	input \WX11171_reg/NET0131  ;
	input \WX11173_reg/NET0131  ;
	input \WX11175_reg/NET0131  ;
	input \WX11177_reg/NET0131  ;
	input \WX11179_reg/NET0131  ;
	input \WX11181_reg/NET0131  ;
	input \WX11183_reg/NET0131  ;
	input \WX11185_reg/NET0131  ;
	input \WX11187_reg/NET0131  ;
	input \WX11189_reg/NET0131  ;
	input \WX11191_reg/NET0131  ;
	input \WX11193_reg/NET0131  ;
	input \WX11195_reg/NET0131  ;
	input \WX11197_reg/NET0131  ;
	input \WX11199_reg/NET0131  ;
	input \WX11201_reg/NET0131  ;
	input \WX11203_reg/NET0131  ;
	input \WX11205_reg/NET0131  ;
	input \WX11207_reg/NET0131  ;
	input \WX11209_reg/NET0131  ;
	input \WX11211_reg/NET0131  ;
	input \WX11213_reg/NET0131  ;
	input \WX11215_reg/NET0131  ;
	input \WX11217_reg/NET0131  ;
	input \WX11219_reg/NET0131  ;
	input \WX11221_reg/NET0131  ;
	input \WX11223_reg/NET0131  ;
	input \WX11225_reg/NET0131  ;
	input \WX11227_reg/NET0131  ;
	input \WX11229_reg/NET0131  ;
	input \WX11231_reg/NET0131  ;
	input \WX11233_reg/NET0131  ;
	input \WX11235_reg/NET0131  ;
	input \WX11237_reg/NET0131  ;
	input \WX11239_reg/NET0131  ;
	input \WX11241_reg/NET0131  ;
	input \WX11243_reg/NET0131  ;
	input \WX1938_reg/NET0131  ;
	input \WX1940_reg/NET0131  ;
	input \WX1942_reg/NET0131  ;
	input \WX1944_reg/NET0131  ;
	input \WX1946_reg/NET0131  ;
	input \WX1948_reg/NET0131  ;
	input \WX1950_reg/NET0131  ;
	input \WX1952_reg/NET0131  ;
	input \WX1954_reg/NET0131  ;
	input \WX1956_reg/NET0131  ;
	input \WX1958_reg/NET0131  ;
	input \WX1960_reg/NET0131  ;
	input \WX1962_reg/NET0131  ;
	input \WX1964_reg/NET0131  ;
	input \WX1966_reg/NET0131  ;
	input \WX1968_reg/NET0131  ;
	input \WX1970_reg/NET0131  ;
	input \WX1972_reg/NET0131  ;
	input \WX1974_reg/NET0131  ;
	input \WX1976_reg/NET0131  ;
	input \WX1978_reg/NET0131  ;
	input \WX1980_reg/NET0131  ;
	input \WX1982_reg/NET0131  ;
	input \WX1984_reg/NET0131  ;
	input \WX1986_reg/NET0131  ;
	input \WX1988_reg/NET0131  ;
	input \WX1990_reg/NET0131  ;
	input \WX1992_reg/NET0131  ;
	input \WX1994_reg/NET0131  ;
	input \WX1996_reg/NET0131  ;
	input \WX1998_reg/NET0131  ;
	input \WX2000_reg/NET0131  ;
	input \WX2002_reg/NET0131  ;
	input \WX2004_reg/NET0131  ;
	input \WX2006_reg/NET0131  ;
	input \WX2008_reg/NET0131  ;
	input \WX2010_reg/NET0131  ;
	input \WX2012_reg/NET0131  ;
	input \WX2014_reg/NET0131  ;
	input \WX2016_reg/NET0131  ;
	input \WX2018_reg/NET0131  ;
	input \WX2020_reg/NET0131  ;
	input \WX2022_reg/NET0131  ;
	input \WX2024_reg/NET0131  ;
	input \WX2026_reg/NET0131  ;
	input \WX2028_reg/NET0131  ;
	input \WX2030_reg/NET0131  ;
	input \WX2032_reg/NET0131  ;
	input \WX2034_reg/NET0131  ;
	input \WX2036_reg/NET0131  ;
	input \WX2038_reg/NET0131  ;
	input \WX2040_reg/NET0131  ;
	input \WX2042_reg/NET0131  ;
	input \WX2044_reg/NET0131  ;
	input \WX2046_reg/NET0131  ;
	input \WX2048_reg/NET0131  ;
	input \WX2050_reg/NET0131  ;
	input \WX2052_reg/NET0131  ;
	input \WX2054_reg/NET0131  ;
	input \WX2056_reg/NET0131  ;
	input \WX2058_reg/NET0131  ;
	input \WX2060_reg/NET0131  ;
	input \WX2062_reg/NET0131  ;
	input \WX2064_reg/NET0131  ;
	input \WX2066_reg/NET0131  ;
	input \WX2068_reg/NET0131  ;
	input \WX2070_reg/NET0131  ;
	input \WX2072_reg/NET0131  ;
	input \WX2074_reg/NET0131  ;
	input \WX2076_reg/NET0131  ;
	input \WX2078_reg/NET0131  ;
	input \WX2080_reg/NET0131  ;
	input \WX2082_reg/NET0131  ;
	input \WX2084_reg/NET0131  ;
	input \WX2086_reg/NET0131  ;
	input \WX2088_reg/NET0131  ;
	input \WX2090_reg/NET0131  ;
	input \WX2092_reg/NET0131  ;
	input \WX2094_reg/NET0131  ;
	input \WX2096_reg/NET0131  ;
	input \WX2098_reg/NET0131  ;
	input \WX2100_reg/NET0131  ;
	input \WX2102_reg/NET0131  ;
	input \WX2104_reg/NET0131  ;
	input \WX2106_reg/NET0131  ;
	input \WX2108_reg/NET0131  ;
	input \WX2110_reg/NET0131  ;
	input \WX2112_reg/NET0131  ;
	input \WX2114_reg/NET0131  ;
	input \WX2116_reg/NET0131  ;
	input \WX2118_reg/NET0131  ;
	input \WX2120_reg/NET0131  ;
	input \WX2122_reg/NET0131  ;
	input \WX2124_reg/NET0131  ;
	input \WX2126_reg/NET0131  ;
	input \WX2128_reg/NET0131  ;
	input \WX2130_reg/NET0131  ;
	input \WX2132_reg/NET0131  ;
	input \WX2134_reg/NET0131  ;
	input \WX2136_reg/NET0131  ;
	input \WX2138_reg/NET0131  ;
	input \WX2140_reg/NET0131  ;
	input \WX2142_reg/NET0131  ;
	input \WX2144_reg/NET0131  ;
	input \WX2146_reg/NET0131  ;
	input \WX2148_reg/NET0131  ;
	input \WX2150_reg/NET0131  ;
	input \WX2152_reg/NET0131  ;
	input \WX2154_reg/NET0131  ;
	input \WX2156_reg/NET0131  ;
	input \WX2158_reg/NET0131  ;
	input \WX2160_reg/NET0131  ;
	input \WX2162_reg/NET0131  ;
	input \WX2164_reg/NET0131  ;
	input \WX2166_reg/NET0131  ;
	input \WX2168_reg/NET0131  ;
	input \WX2170_reg/NET0131  ;
	input \WX2172_reg/NET0131  ;
	input \WX2174_reg/NET0131  ;
	input \WX2176_reg/NET0131  ;
	input \WX2178_reg/NET0131  ;
	input \WX2180_reg/NET0131  ;
	input \WX2182_reg/NET0131  ;
	input \WX2184_reg/NET0131  ;
	input \WX2186_reg/NET0131  ;
	input \WX2188_reg/NET0131  ;
	input \WX2190_reg/NET0131  ;
	input \WX2192_reg/NET0131  ;
	input \WX3231_reg/NET0131  ;
	input \WX3233_reg/NET0131  ;
	input \WX3235_reg/NET0131  ;
	input \WX3237_reg/NET0131  ;
	input \WX3239_reg/NET0131  ;
	input \WX3241_reg/NET0131  ;
	input \WX3243_reg/NET0131  ;
	input \WX3245_reg/NET0131  ;
	input \WX3247_reg/NET0131  ;
	input \WX3249_reg/NET0131  ;
	input \WX3251_reg/NET0131  ;
	input \WX3253_reg/NET0131  ;
	input \WX3255_reg/NET0131  ;
	input \WX3257_reg/NET0131  ;
	input \WX3259_reg/NET0131  ;
	input \WX3261_reg/NET0131  ;
	input \WX3263_reg/NET0131  ;
	input \WX3265_reg/NET0131  ;
	input \WX3267_reg/NET0131  ;
	input \WX3269_reg/NET0131  ;
	input \WX3271_reg/NET0131  ;
	input \WX3273_reg/NET0131  ;
	input \WX3275_reg/NET0131  ;
	input \WX3277_reg/NET0131  ;
	input \WX3279_reg/NET0131  ;
	input \WX3281_reg/NET0131  ;
	input \WX3283_reg/NET0131  ;
	input \WX3285_reg/NET0131  ;
	input \WX3287_reg/NET0131  ;
	input \WX3289_reg/NET0131  ;
	input \WX3291_reg/NET0131  ;
	input \WX3293_reg/NET0131  ;
	input \WX3295_reg/NET0131  ;
	input \WX3297_reg/NET0131  ;
	input \WX3299_reg/NET0131  ;
	input \WX3301_reg/NET0131  ;
	input \WX3303_reg/NET0131  ;
	input \WX3305_reg/NET0131  ;
	input \WX3307_reg/NET0131  ;
	input \WX3309_reg/NET0131  ;
	input \WX3311_reg/NET0131  ;
	input \WX3313_reg/NET0131  ;
	input \WX3315_reg/NET0131  ;
	input \WX3317_reg/NET0131  ;
	input \WX3319_reg/NET0131  ;
	input \WX3321_reg/NET0131  ;
	input \WX3323_reg/NET0131  ;
	input \WX3325_reg/NET0131  ;
	input \WX3327_reg/NET0131  ;
	input \WX3329_reg/NET0131  ;
	input \WX3331_reg/NET0131  ;
	input \WX3333_reg/NET0131  ;
	input \WX3335_reg/NET0131  ;
	input \WX3337_reg/NET0131  ;
	input \WX3339_reg/NET0131  ;
	input \WX3341_reg/NET0131  ;
	input \WX3343_reg/NET0131  ;
	input \WX3345_reg/NET0131  ;
	input \WX3347_reg/NET0131  ;
	input \WX3349_reg/NET0131  ;
	input \WX3351_reg/NET0131  ;
	input \WX3353_reg/NET0131  ;
	input \WX3355_reg/NET0131  ;
	input \WX3357_reg/NET0131  ;
	input \WX3359_reg/NET0131  ;
	input \WX3361_reg/NET0131  ;
	input \WX3363_reg/NET0131  ;
	input \WX3365_reg/NET0131  ;
	input \WX3367_reg/NET0131  ;
	input \WX3369_reg/NET0131  ;
	input \WX3371_reg/NET0131  ;
	input \WX3373_reg/NET0131  ;
	input \WX3375_reg/NET0131  ;
	input \WX3377_reg/NET0131  ;
	input \WX3379_reg/NET0131  ;
	input \WX3381_reg/NET0131  ;
	input \WX3383_reg/NET0131  ;
	input \WX3385_reg/NET0131  ;
	input \WX3387_reg/NET0131  ;
	input \WX3389_reg/NET0131  ;
	input \WX3391_reg/NET0131  ;
	input \WX3393_reg/NET0131  ;
	input \WX3395_reg/NET0131  ;
	input \WX3397_reg/NET0131  ;
	input \WX3399_reg/NET0131  ;
	input \WX3401_reg/NET0131  ;
	input \WX3403_reg/NET0131  ;
	input \WX3405_reg/NET0131  ;
	input \WX3407_reg/NET0131  ;
	input \WX3409_reg/NET0131  ;
	input \WX3411_reg/NET0131  ;
	input \WX3413_reg/NET0131  ;
	input \WX3415_reg/NET0131  ;
	input \WX3417_reg/NET0131  ;
	input \WX3419_reg/NET0131  ;
	input \WX3421_reg/NET0131  ;
	input \WX3423_reg/NET0131  ;
	input \WX3425_reg/NET0131  ;
	input \WX3427_reg/NET0131  ;
	input \WX3429_reg/NET0131  ;
	input \WX3431_reg/NET0131  ;
	input \WX3433_reg/NET0131  ;
	input \WX3435_reg/NET0131  ;
	input \WX3437_reg/NET0131  ;
	input \WX3439_reg/NET0131  ;
	input \WX3441_reg/NET0131  ;
	input \WX3443_reg/NET0131  ;
	input \WX3445_reg/NET0131  ;
	input \WX3447_reg/NET0131  ;
	input \WX3449_reg/NET0131  ;
	input \WX3451_reg/NET0131  ;
	input \WX3453_reg/NET0131  ;
	input \WX3455_reg/NET0131  ;
	input \WX3457_reg/NET0131  ;
	input \WX3459_reg/NET0131  ;
	input \WX3461_reg/NET0131  ;
	input \WX3463_reg/NET0131  ;
	input \WX3465_reg/NET0131  ;
	input \WX3467_reg/NET0131  ;
	input \WX3469_reg/NET0131  ;
	input \WX3471_reg/NET0131  ;
	input \WX3473_reg/NET0131  ;
	input \WX3475_reg/NET0131  ;
	input \WX3477_reg/NET0131  ;
	input \WX3479_reg/NET0131  ;
	input \WX3481_reg/NET0131  ;
	input \WX3483_reg/NET0131  ;
	input \WX3485_reg/NET0131  ;
	input \WX4524_reg/NET0131  ;
	input \WX4526_reg/NET0131  ;
	input \WX4528_reg/NET0131  ;
	input \WX4530_reg/NET0131  ;
	input \WX4532_reg/NET0131  ;
	input \WX4534_reg/NET0131  ;
	input \WX4536_reg/NET0131  ;
	input \WX4538_reg/NET0131  ;
	input \WX4540_reg/NET0131  ;
	input \WX4542_reg/NET0131  ;
	input \WX4544_reg/NET0131  ;
	input \WX4546_reg/NET0131  ;
	input \WX4548_reg/NET0131  ;
	input \WX4550_reg/NET0131  ;
	input \WX4552_reg/NET0131  ;
	input \WX4554_reg/NET0131  ;
	input \WX4556_reg/NET0131  ;
	input \WX4558_reg/NET0131  ;
	input \WX4560_reg/NET0131  ;
	input \WX4562_reg/NET0131  ;
	input \WX4564_reg/NET0131  ;
	input \WX4566_reg/NET0131  ;
	input \WX4568_reg/NET0131  ;
	input \WX4570_reg/NET0131  ;
	input \WX4572_reg/NET0131  ;
	input \WX4574_reg/NET0131  ;
	input \WX4576_reg/NET0131  ;
	input \WX4578_reg/NET0131  ;
	input \WX4580_reg/NET0131  ;
	input \WX4582_reg/NET0131  ;
	input \WX4584_reg/NET0131  ;
	input \WX4586_reg/NET0131  ;
	input \WX4588_reg/NET0131  ;
	input \WX4590_reg/NET0131  ;
	input \WX4592_reg/NET0131  ;
	input \WX4594_reg/NET0131  ;
	input \WX4596_reg/NET0131  ;
	input \WX4598_reg/NET0131  ;
	input \WX4600_reg/NET0131  ;
	input \WX4602_reg/NET0131  ;
	input \WX4604_reg/NET0131  ;
	input \WX4606_reg/NET0131  ;
	input \WX4608_reg/NET0131  ;
	input \WX4610_reg/NET0131  ;
	input \WX4612_reg/NET0131  ;
	input \WX4614_reg/NET0131  ;
	input \WX4616_reg/NET0131  ;
	input \WX4618_reg/NET0131  ;
	input \WX4620_reg/NET0131  ;
	input \WX4622_reg/NET0131  ;
	input \WX4624_reg/NET0131  ;
	input \WX4626_reg/NET0131  ;
	input \WX4628_reg/NET0131  ;
	input \WX4630_reg/NET0131  ;
	input \WX4632_reg/NET0131  ;
	input \WX4634_reg/NET0131  ;
	input \WX4636_reg/NET0131  ;
	input \WX4638_reg/NET0131  ;
	input \WX4640_reg/NET0131  ;
	input \WX4642_reg/NET0131  ;
	input \WX4644_reg/NET0131  ;
	input \WX4646_reg/NET0131  ;
	input \WX4648_reg/NET0131  ;
	input \WX4650_reg/NET0131  ;
	input \WX4652_reg/NET0131  ;
	input \WX4654_reg/NET0131  ;
	input \WX4656_reg/NET0131  ;
	input \WX4658_reg/NET0131  ;
	input \WX4660_reg/NET0131  ;
	input \WX4662_reg/NET0131  ;
	input \WX4664_reg/NET0131  ;
	input \WX4666_reg/NET0131  ;
	input \WX4668_reg/NET0131  ;
	input \WX4670_reg/NET0131  ;
	input \WX4672_reg/NET0131  ;
	input \WX4674_reg/NET0131  ;
	input \WX4676_reg/NET0131  ;
	input \WX4678_reg/NET0131  ;
	input \WX4680_reg/NET0131  ;
	input \WX4682_reg/NET0131  ;
	input \WX4684_reg/NET0131  ;
	input \WX4686_reg/NET0131  ;
	input \WX4688_reg/NET0131  ;
	input \WX4690_reg/NET0131  ;
	input \WX4692_reg/NET0131  ;
	input \WX4694_reg/NET0131  ;
	input \WX4696_reg/NET0131  ;
	input \WX4698_reg/NET0131  ;
	input \WX4700_reg/NET0131  ;
	input \WX4702_reg/NET0131  ;
	input \WX4704_reg/NET0131  ;
	input \WX4706_reg/NET0131  ;
	input \WX4708_reg/NET0131  ;
	input \WX4710_reg/NET0131  ;
	input \WX4712_reg/NET0131  ;
	input \WX4714_reg/NET0131  ;
	input \WX4716_reg/NET0131  ;
	input \WX4718_reg/NET0131  ;
	input \WX4720_reg/NET0131  ;
	input \WX4722_reg/NET0131  ;
	input \WX4724_reg/NET0131  ;
	input \WX4726_reg/NET0131  ;
	input \WX4728_reg/NET0131  ;
	input \WX4730_reg/NET0131  ;
	input \WX4732_reg/NET0131  ;
	input \WX4734_reg/NET0131  ;
	input \WX4736_reg/NET0131  ;
	input \WX4738_reg/NET0131  ;
	input \WX4740_reg/NET0131  ;
	input \WX4742_reg/NET0131  ;
	input \WX4744_reg/NET0131  ;
	input \WX4746_reg/NET0131  ;
	input \WX4748_reg/NET0131  ;
	input \WX4750_reg/NET0131  ;
	input \WX4752_reg/NET0131  ;
	input \WX4754_reg/NET0131  ;
	input \WX4756_reg/NET0131  ;
	input \WX4758_reg/NET0131  ;
	input \WX4760_reg/NET0131  ;
	input \WX4762_reg/NET0131  ;
	input \WX4764_reg/NET0131  ;
	input \WX4766_reg/NET0131  ;
	input \WX4768_reg/NET0131  ;
	input \WX4770_reg/NET0131  ;
	input \WX4772_reg/NET0131  ;
	input \WX4774_reg/NET0131  ;
	input \WX4776_reg/NET0131  ;
	input \WX4778_reg/NET0131  ;
	input \WX5817_reg/NET0131  ;
	input \WX5819_reg/NET0131  ;
	input \WX5821_reg/NET0131  ;
	input \WX5823_reg/NET0131  ;
	input \WX5825_reg/NET0131  ;
	input \WX5827_reg/NET0131  ;
	input \WX5829_reg/NET0131  ;
	input \WX5831_reg/NET0131  ;
	input \WX5833_reg/NET0131  ;
	input \WX5835_reg/NET0131  ;
	input \WX5837_reg/NET0131  ;
	input \WX5839_reg/NET0131  ;
	input \WX5841_reg/NET0131  ;
	input \WX5843_reg/NET0131  ;
	input \WX5845_reg/NET0131  ;
	input \WX5847_reg/NET0131  ;
	input \WX5849_reg/NET0131  ;
	input \WX5851_reg/NET0131  ;
	input \WX5853_reg/NET0131  ;
	input \WX5855_reg/NET0131  ;
	input \WX5857_reg/NET0131  ;
	input \WX5859_reg/NET0131  ;
	input \WX5861_reg/NET0131  ;
	input \WX5863_reg/NET0131  ;
	input \WX5865_reg/NET0131  ;
	input \WX5867_reg/NET0131  ;
	input \WX5869_reg/NET0131  ;
	input \WX5871_reg/NET0131  ;
	input \WX5873_reg/NET0131  ;
	input \WX5875_reg/NET0131  ;
	input \WX5877_reg/NET0131  ;
	input \WX5879_reg/NET0131  ;
	input \WX5881_reg/NET0131  ;
	input \WX5883_reg/NET0131  ;
	input \WX5885_reg/NET0131  ;
	input \WX5887_reg/NET0131  ;
	input \WX5889_reg/NET0131  ;
	input \WX5891_reg/NET0131  ;
	input \WX5893_reg/NET0131  ;
	input \WX5895_reg/NET0131  ;
	input \WX5897_reg/NET0131  ;
	input \WX5899_reg/NET0131  ;
	input \WX5901_reg/NET0131  ;
	input \WX5903_reg/NET0131  ;
	input \WX5905_reg/NET0131  ;
	input \WX5907_reg/NET0131  ;
	input \WX5909_reg/NET0131  ;
	input \WX5911_reg/NET0131  ;
	input \WX5913_reg/NET0131  ;
	input \WX5915_reg/NET0131  ;
	input \WX5917_reg/NET0131  ;
	input \WX5919_reg/NET0131  ;
	input \WX5921_reg/NET0131  ;
	input \WX5923_reg/NET0131  ;
	input \WX5925_reg/NET0131  ;
	input \WX5927_reg/NET0131  ;
	input \WX5929_reg/NET0131  ;
	input \WX5931_reg/NET0131  ;
	input \WX5933_reg/NET0131  ;
	input \WX5935_reg/NET0131  ;
	input \WX5937_reg/NET0131  ;
	input \WX5939_reg/NET0131  ;
	input \WX5941_reg/NET0131  ;
	input \WX5943_reg/NET0131  ;
	input \WX5945_reg/NET0131  ;
	input \WX5947_reg/NET0131  ;
	input \WX5949_reg/NET0131  ;
	input \WX5951_reg/NET0131  ;
	input \WX5953_reg/NET0131  ;
	input \WX5955_reg/NET0131  ;
	input \WX5957_reg/NET0131  ;
	input \WX5959_reg/NET0131  ;
	input \WX5961_reg/NET0131  ;
	input \WX5963_reg/NET0131  ;
	input \WX5965_reg/NET0131  ;
	input \WX5967_reg/NET0131  ;
	input \WX5969_reg/NET0131  ;
	input \WX5971_reg/NET0131  ;
	input \WX5973_reg/NET0131  ;
	input \WX5975_reg/NET0131  ;
	input \WX5977_reg/NET0131  ;
	input \WX5979_reg/NET0131  ;
	input \WX5981_reg/NET0131  ;
	input \WX5983_reg/NET0131  ;
	input \WX5985_reg/NET0131  ;
	input \WX5987_reg/NET0131  ;
	input \WX5989_reg/NET0131  ;
	input \WX5991_reg/NET0131  ;
	input \WX5993_reg/NET0131  ;
	input \WX5995_reg/NET0131  ;
	input \WX5997_reg/NET0131  ;
	input \WX5999_reg/NET0131  ;
	input \WX6001_reg/NET0131  ;
	input \WX6003_reg/NET0131  ;
	input \WX6005_reg/NET0131  ;
	input \WX6007_reg/NET0131  ;
	input \WX6009_reg/NET0131  ;
	input \WX6011_reg/NET0131  ;
	input \WX6013_reg/NET0131  ;
	input \WX6015_reg/NET0131  ;
	input \WX6017_reg/NET0131  ;
	input \WX6019_reg/NET0131  ;
	input \WX6021_reg/NET0131  ;
	input \WX6023_reg/NET0131  ;
	input \WX6025_reg/NET0131  ;
	input \WX6027_reg/NET0131  ;
	input \WX6029_reg/NET0131  ;
	input \WX6031_reg/NET0131  ;
	input \WX6033_reg/NET0131  ;
	input \WX6035_reg/NET0131  ;
	input \WX6037_reg/NET0131  ;
	input \WX6039_reg/NET0131  ;
	input \WX6041_reg/NET0131  ;
	input \WX6043_reg/NET0131  ;
	input \WX6045_reg/NET0131  ;
	input \WX6047_reg/NET0131  ;
	input \WX6049_reg/NET0131  ;
	input \WX6051_reg/NET0131  ;
	input \WX6053_reg/NET0131  ;
	input \WX6055_reg/NET0131  ;
	input \WX6057_reg/NET0131  ;
	input \WX6059_reg/NET0131  ;
	input \WX6061_reg/NET0131  ;
	input \WX6063_reg/NET0131  ;
	input \WX6065_reg/NET0131  ;
	input \WX6067_reg/NET0131  ;
	input \WX6069_reg/NET0131  ;
	input \WX6071_reg/NET0131  ;
	input \WX645_reg/NET0131  ;
	input \WX647_reg/NET0131  ;
	input \WX649_reg/NET0131  ;
	input \WX651_reg/NET0131  ;
	input \WX653_reg/NET0131  ;
	input \WX655_reg/NET0131  ;
	input \WX657_reg/NET0131  ;
	input \WX659_reg/NET0131  ;
	input \WX661_reg/NET0131  ;
	input \WX663_reg/NET0131  ;
	input \WX665_reg/NET0131  ;
	input \WX667_reg/NET0131  ;
	input \WX669_reg/NET0131  ;
	input \WX671_reg/NET0131  ;
	input \WX673_reg/NET0131  ;
	input \WX675_reg/NET0131  ;
	input \WX677_reg/NET0131  ;
	input \WX679_reg/NET0131  ;
	input \WX681_reg/NET0131  ;
	input \WX683_reg/NET0131  ;
	input \WX685_reg/NET0131  ;
	input \WX687_reg/NET0131  ;
	input \WX689_reg/NET0131  ;
	input \WX691_reg/NET0131  ;
	input \WX693_reg/NET0131  ;
	input \WX695_reg/NET0131  ;
	input \WX697_reg/NET0131  ;
	input \WX699_reg/NET0131  ;
	input \WX701_reg/NET0131  ;
	input \WX703_reg/NET0131  ;
	input \WX705_reg/NET0131  ;
	input \WX707_reg/NET0131  ;
	input \WX709_reg/NET0131  ;
	input \WX7110_reg/NET0131  ;
	input \WX7112_reg/NET0131  ;
	input \WX7114_reg/NET0131  ;
	input \WX7116_reg/NET0131  ;
	input \WX7118_reg/NET0131  ;
	input \WX711_reg/NET0131  ;
	input \WX7120_reg/NET0131  ;
	input \WX7122_reg/NET0131  ;
	input \WX7124_reg/NET0131  ;
	input \WX7126_reg/NET0131  ;
	input \WX7128_reg/NET0131  ;
	input \WX7130_reg/NET0131  ;
	input \WX7132_reg/NET0131  ;
	input \WX7134_reg/NET0131  ;
	input \WX7136_reg/NET0131  ;
	input \WX7138_reg/NET0131  ;
	input \WX713_reg/NET0131  ;
	input \WX7140_reg/NET0131  ;
	input \WX7142_reg/NET0131  ;
	input \WX7144_reg/NET0131  ;
	input \WX7146_reg/NET0131  ;
	input \WX7148_reg/NET0131  ;
	input \WX7150_reg/NET0131  ;
	input \WX7152_reg/NET0131  ;
	input \WX7154_reg/NET0131  ;
	input \WX7156_reg/NET0131  ;
	input \WX7158_reg/NET0131  ;
	input \WX715_reg/NET0131  ;
	input \WX7160_reg/NET0131  ;
	input \WX7162_reg/NET0131  ;
	input \WX7164_reg/NET0131  ;
	input \WX7166_reg/NET0131  ;
	input \WX7168_reg/NET0131  ;
	input \WX7170_reg/NET0131  ;
	input \WX7172_reg/NET0131  ;
	input \WX7174_reg/NET0131  ;
	input \WX7176_reg/NET0131  ;
	input \WX7178_reg/NET0131  ;
	input \WX717_reg/NET0131  ;
	input \WX7180_reg/NET0131  ;
	input \WX7182_reg/NET0131  ;
	input \WX7184_reg/NET0131  ;
	input \WX7186_reg/NET0131  ;
	input \WX7188_reg/NET0131  ;
	input \WX7190_reg/NET0131  ;
	input \WX7192_reg/NET0131  ;
	input \WX7194_reg/NET0131  ;
	input \WX7196_reg/NET0131  ;
	input \WX7198_reg/NET0131  ;
	input \WX719_reg/NET0131  ;
	input \WX7200_reg/NET0131  ;
	input \WX7202_reg/NET0131  ;
	input \WX7204_reg/NET0131  ;
	input \WX7206_reg/NET0131  ;
	input \WX7208_reg/NET0131  ;
	input \WX7210_reg/NET0131  ;
	input \WX7212_reg/NET0131  ;
	input \WX7214_reg/NET0131  ;
	input \WX7216_reg/NET0131  ;
	input \WX7218_reg/NET0131  ;
	input \WX721_reg/NET0131  ;
	input \WX7220_reg/NET0131  ;
	input \WX7222_reg/NET0131  ;
	input \WX7224_reg/NET0131  ;
	input \WX7226_reg/NET0131  ;
	input \WX7228_reg/NET0131  ;
	input \WX7230_reg/NET0131  ;
	input \WX7232_reg/NET0131  ;
	input \WX7234_reg/NET0131  ;
	input \WX7236_reg/NET0131  ;
	input \WX7238_reg/NET0131  ;
	input \WX723_reg/NET0131  ;
	input \WX7240_reg/NET0131  ;
	input \WX7242_reg/NET0131  ;
	input \WX7244_reg/NET0131  ;
	input \WX7246_reg/NET0131  ;
	input \WX7248_reg/NET0131  ;
	input \WX7250_reg/NET0131  ;
	input \WX7252_reg/NET0131  ;
	input \WX7254_reg/NET0131  ;
	input \WX7256_reg/NET0131  ;
	input \WX7258_reg/NET0131  ;
	input \WX725_reg/NET0131  ;
	input \WX7260_reg/NET0131  ;
	input \WX7262_reg/NET0131  ;
	input \WX7264_reg/NET0131  ;
	input \WX7266_reg/NET0131  ;
	input \WX7268_reg/NET0131  ;
	input \WX7270_reg/NET0131  ;
	input \WX7272_reg/NET0131  ;
	input \WX7274_reg/NET0131  ;
	input \WX7276_reg/NET0131  ;
	input \WX7278_reg/NET0131  ;
	input \WX727_reg/NET0131  ;
	input \WX7280_reg/NET0131  ;
	input \WX7282_reg/NET0131  ;
	input \WX7284_reg/NET0131  ;
	input \WX7286_reg/NET0131  ;
	input \WX7288_reg/NET0131  ;
	input \WX7290_reg/NET0131  ;
	input \WX7292_reg/NET0131  ;
	input \WX7294_reg/NET0131  ;
	input \WX7296_reg/NET0131  ;
	input \WX7298_reg/NET0131  ;
	input \WX729_reg/NET0131  ;
	input \WX7300_reg/NET0131  ;
	input \WX7302_reg/NET0131  ;
	input \WX7304_reg/NET0131  ;
	input \WX7306_reg/NET0131  ;
	input \WX7308_reg/NET0131  ;
	input \WX7310_reg/NET0131  ;
	input \WX7312_reg/NET0131  ;
	input \WX7314_reg/NET0131  ;
	input \WX7316_reg/NET0131  ;
	input \WX7318_reg/NET0131  ;
	input \WX731_reg/NET0131  ;
	input \WX7320_reg/NET0131  ;
	input \WX7322_reg/NET0131  ;
	input \WX7324_reg/NET0131  ;
	input \WX7326_reg/NET0131  ;
	input \WX7328_reg/NET0131  ;
	input \WX7330_reg/NET0131  ;
	input \WX7332_reg/NET0131  ;
	input \WX7334_reg/NET0131  ;
	input \WX7336_reg/NET0131  ;
	input \WX7338_reg/NET0131  ;
	input \WX733_reg/NET0131  ;
	input \WX7340_reg/NET0131  ;
	input \WX7342_reg/NET0131  ;
	input \WX7344_reg/NET0131  ;
	input \WX7346_reg/NET0131  ;
	input \WX7348_reg/NET0131  ;
	input \WX7350_reg/NET0131  ;
	input \WX7352_reg/NET0131  ;
	input \WX7354_reg/NET0131  ;
	input \WX7356_reg/NET0131  ;
	input \WX7358_reg/NET0131  ;
	input \WX735_reg/NET0131  ;
	input \WX7360_reg/NET0131  ;
	input \WX7362_reg/NET0131  ;
	input \WX7364_reg/NET0131  ;
	input \WX737_reg/NET0131  ;
	input \WX739_reg/NET0131  ;
	input \WX741_reg/NET0131  ;
	input \WX743_reg/NET0131  ;
	input \WX745_reg/NET0131  ;
	input \WX747_reg/NET0131  ;
	input \WX749_reg/NET0131  ;
	input \WX751_reg/NET0131  ;
	input \WX753_reg/NET0131  ;
	input \WX755_reg/NET0131  ;
	input \WX757_reg/NET0131  ;
	input \WX759_reg/NET0131  ;
	input \WX761_reg/NET0131  ;
	input \WX763_reg/NET0131  ;
	input \WX765_reg/NET0131  ;
	input \WX767_reg/NET0131  ;
	input \WX769_reg/NET0131  ;
	input \WX771_reg/NET0131  ;
	input \WX773_reg/NET0131  ;
	input \WX775_reg/NET0131  ;
	input \WX777_reg/NET0131  ;
	input \WX779_reg/NET0131  ;
	input \WX781_reg/NET0131  ;
	input \WX783_reg/NET0131  ;
	input \WX785_reg/NET0131  ;
	input \WX787_reg/NET0131  ;
	input \WX789_reg/NET0131  ;
	input \WX791_reg/NET0131  ;
	input \WX793_reg/NET0131  ;
	input \WX795_reg/NET0131  ;
	input \WX797_reg/NET0131  ;
	input \WX799_reg/NET0131  ;
	input \WX801_reg/NET0131  ;
	input \WX803_reg/NET0131  ;
	input \WX805_reg/NET0131  ;
	input \WX807_reg/NET0131  ;
	input \WX809_reg/NET0131  ;
	input \WX811_reg/NET0131  ;
	input \WX813_reg/NET0131  ;
	input \WX815_reg/NET0131  ;
	input \WX817_reg/NET0131  ;
	input \WX819_reg/NET0131  ;
	input \WX821_reg/NET0131  ;
	input \WX823_reg/NET0131  ;
	input \WX825_reg/NET0131  ;
	input \WX827_reg/NET0131  ;
	input \WX829_reg/NET0131  ;
	input \WX831_reg/NET0131  ;
	input \WX833_reg/NET0131  ;
	input \WX835_reg/NET0131  ;
	input \WX837_reg/NET0131  ;
	input \WX839_reg/NET0131  ;
	input \WX8403_reg/NET0131  ;
	input \WX8405_reg/NET0131  ;
	input \WX8407_reg/NET0131  ;
	input \WX8409_reg/NET0131  ;
	input \WX8411_reg/NET0131  ;
	input \WX8413_reg/NET0131  ;
	input \WX8415_reg/NET0131  ;
	input \WX8417_reg/NET0131  ;
	input \WX8419_reg/NET0131  ;
	input \WX841_reg/NET0131  ;
	input \WX8421_reg/NET0131  ;
	input \WX8423_reg/NET0131  ;
	input \WX8425_reg/NET0131  ;
	input \WX8427_reg/NET0131  ;
	input \WX8429_reg/NET0131  ;
	input \WX8431_reg/NET0131  ;
	input \WX8433_reg/NET0131  ;
	input \WX8435_reg/NET0131  ;
	input \WX8437_reg/NET0131  ;
	input \WX8439_reg/NET0131  ;
	input \WX843_reg/NET0131  ;
	input \WX8441_reg/NET0131  ;
	input \WX8443_reg/NET0131  ;
	input \WX8445_reg/NET0131  ;
	input \WX8447_reg/NET0131  ;
	input \WX8449_reg/NET0131  ;
	input \WX8451_reg/NET0131  ;
	input \WX8453_reg/NET0131  ;
	input \WX8455_reg/NET0131  ;
	input \WX8457_reg/NET0131  ;
	input \WX8459_reg/NET0131  ;
	input \WX845_reg/NET0131  ;
	input \WX8461_reg/NET0131  ;
	input \WX8463_reg/NET0131  ;
	input \WX8465_reg/NET0131  ;
	input \WX8467_reg/NET0131  ;
	input \WX8469_reg/NET0131  ;
	input \WX8471_reg/NET0131  ;
	input \WX8473_reg/NET0131  ;
	input \WX8475_reg/NET0131  ;
	input \WX8477_reg/NET0131  ;
	input \WX8479_reg/NET0131  ;
	input \WX847_reg/NET0131  ;
	input \WX8481_reg/NET0131  ;
	input \WX8483_reg/NET0131  ;
	input \WX8485_reg/NET0131  ;
	input \WX8487_reg/NET0131  ;
	input \WX8489_reg/NET0131  ;
	input \WX8491_reg/NET0131  ;
	input \WX8493_reg/NET0131  ;
	input \WX8495_reg/NET0131  ;
	input \WX8497_reg/NET0131  ;
	input \WX8499_reg/NET0131  ;
	input \WX849_reg/NET0131  ;
	input \WX8501_reg/NET0131  ;
	input \WX8503_reg/NET0131  ;
	input \WX8505_reg/NET0131  ;
	input \WX8507_reg/NET0131  ;
	input \WX8509_reg/NET0131  ;
	input \WX8511_reg/NET0131  ;
	input \WX8513_reg/NET0131  ;
	input \WX8515_reg/NET0131  ;
	input \WX8517_reg/NET0131  ;
	input \WX8519_reg/NET0131  ;
	input \WX851_reg/NET0131  ;
	input \WX8521_reg/NET0131  ;
	input \WX8523_reg/NET0131  ;
	input \WX8525_reg/NET0131  ;
	input \WX8527_reg/NET0131  ;
	input \WX8529_reg/NET0131  ;
	input \WX8531_reg/NET0131  ;
	input \WX8533_reg/NET0131  ;
	input \WX8535_reg/NET0131  ;
	input \WX8537_reg/NET0131  ;
	input \WX8539_reg/NET0131  ;
	input \WX853_reg/NET0131  ;
	input \WX8541_reg/NET0131  ;
	input \WX8543_reg/NET0131  ;
	input \WX8545_reg/NET0131  ;
	input \WX8547_reg/NET0131  ;
	input \WX8549_reg/NET0131  ;
	input \WX8551_reg/NET0131  ;
	input \WX8553_reg/NET0131  ;
	input \WX8555_reg/NET0131  ;
	input \WX8557_reg/NET0131  ;
	input \WX8559_reg/NET0131  ;
	input \WX855_reg/NET0131  ;
	input \WX8561_reg/NET0131  ;
	input \WX8563_reg/NET0131  ;
	input \WX8565_reg/NET0131  ;
	input \WX8567_reg/NET0131  ;
	input \WX8569_reg/NET0131  ;
	input \WX8571_reg/NET0131  ;
	input \WX8573_reg/NET0131  ;
	input \WX8575_reg/NET0131  ;
	input \WX8577_reg/NET0131  ;
	input \WX8579_reg/NET0131  ;
	input \WX857_reg/NET0131  ;
	input \WX8581_reg/NET0131  ;
	input \WX8583_reg/NET0131  ;
	input \WX8585_reg/NET0131  ;
	input \WX8587_reg/NET0131  ;
	input \WX8589_reg/NET0131  ;
	input \WX8591_reg/NET0131  ;
	input \WX8593_reg/NET0131  ;
	input \WX8595_reg/NET0131  ;
	input \WX8597_reg/NET0131  ;
	input \WX8599_reg/NET0131  ;
	input \WX859_reg/NET0131  ;
	input \WX8601_reg/NET0131  ;
	input \WX8603_reg/NET0131  ;
	input \WX8605_reg/NET0131  ;
	input \WX8607_reg/NET0131  ;
	input \WX8609_reg/NET0131  ;
	input \WX8611_reg/NET0131  ;
	input \WX8613_reg/NET0131  ;
	input \WX8615_reg/NET0131  ;
	input \WX8617_reg/NET0131  ;
	input \WX8619_reg/NET0131  ;
	input \WX861_reg/NET0131  ;
	input \WX8621_reg/NET0131  ;
	input \WX8623_reg/NET0131  ;
	input \WX8625_reg/NET0131  ;
	input \WX8627_reg/NET0131  ;
	input \WX8629_reg/NET0131  ;
	input \WX8631_reg/NET0131  ;
	input \WX8633_reg/NET0131  ;
	input \WX8635_reg/NET0131  ;
	input \WX8637_reg/NET0131  ;
	input \WX8639_reg/NET0131  ;
	input \WX863_reg/NET0131  ;
	input \WX8641_reg/NET0131  ;
	input \WX8643_reg/NET0131  ;
	input \WX8645_reg/NET0131  ;
	input \WX8647_reg/NET0131  ;
	input \WX8649_reg/NET0131  ;
	input \WX8651_reg/NET0131  ;
	input \WX8653_reg/NET0131  ;
	input \WX8655_reg/NET0131  ;
	input \WX8657_reg/NET0131  ;
	input \WX865_reg/NET0131  ;
	input \WX867_reg/NET0131  ;
	input \WX869_reg/NET0131  ;
	input \WX871_reg/NET0131  ;
	input \WX873_reg/NET0131  ;
	input \WX875_reg/NET0131  ;
	input \WX877_reg/NET0131  ;
	input \WX879_reg/NET0131  ;
	input \WX881_reg/NET0131  ;
	input \WX883_reg/NET0131  ;
	input \WX885_reg/NET0131  ;
	input \WX887_reg/NET0131  ;
	input \WX889_reg/NET0131  ;
	input \WX891_reg/NET0131  ;
	input \WX893_reg/NET0131  ;
	input \WX895_reg/NET0131  ;
	input \WX897_reg/NET0131  ;
	input \WX899_reg/NET0131  ;
	input \WX9696_reg/NET0131  ;
	input \WX9698_reg/NET0131  ;
	input \WX9700_reg/NET0131  ;
	input \WX9702_reg/NET0131  ;
	input \WX9704_reg/NET0131  ;
	input \WX9706_reg/NET0131  ;
	input \WX9708_reg/NET0131  ;
	input \WX9710_reg/NET0131  ;
	input \WX9712_reg/NET0131  ;
	input \WX9714_reg/NET0131  ;
	input \WX9716_reg/NET0131  ;
	input \WX9718_reg/NET0131  ;
	input \WX9720_reg/NET0131  ;
	input \WX9722_reg/NET0131  ;
	input \WX9724_reg/NET0131  ;
	input \WX9726_reg/NET0131  ;
	input \WX9728_reg/NET0131  ;
	input \WX9730_reg/NET0131  ;
	input \WX9732_reg/NET0131  ;
	input \WX9734_reg/NET0131  ;
	input \WX9736_reg/NET0131  ;
	input \WX9738_reg/NET0131  ;
	input \WX9740_reg/NET0131  ;
	input \WX9742_reg/NET0131  ;
	input \WX9744_reg/NET0131  ;
	input \WX9746_reg/NET0131  ;
	input \WX9748_reg/NET0131  ;
	input \WX9750_reg/NET0131  ;
	input \WX9752_reg/NET0131  ;
	input \WX9754_reg/NET0131  ;
	input \WX9756_reg/NET0131  ;
	input \WX9758_reg/NET0131  ;
	input \WX9760_reg/NET0131  ;
	input \WX9762_reg/NET0131  ;
	input \WX9764_reg/NET0131  ;
	input \WX9766_reg/NET0131  ;
	input \WX9768_reg/NET0131  ;
	input \WX9770_reg/NET0131  ;
	input \WX9772_reg/NET0131  ;
	input \WX9774_reg/NET0131  ;
	input \WX9776_reg/NET0131  ;
	input \WX9778_reg/NET0131  ;
	input \WX9780_reg/NET0131  ;
	input \WX9782_reg/NET0131  ;
	input \WX9784_reg/NET0131  ;
	input \WX9786_reg/NET0131  ;
	input \WX9788_reg/NET0131  ;
	input \WX9790_reg/NET0131  ;
	input \WX9792_reg/NET0131  ;
	input \WX9794_reg/NET0131  ;
	input \WX9796_reg/NET0131  ;
	input \WX9798_reg/NET0131  ;
	input \WX9800_reg/NET0131  ;
	input \WX9802_reg/NET0131  ;
	input \WX9804_reg/NET0131  ;
	input \WX9806_reg/NET0131  ;
	input \WX9808_reg/NET0131  ;
	input \WX9810_reg/NET0131  ;
	input \WX9812_reg/NET0131  ;
	input \WX9814_reg/NET0131  ;
	input \WX9816_reg/NET0131  ;
	input \WX9818_reg/NET0131  ;
	input \WX9820_reg/NET0131  ;
	input \WX9822_reg/NET0131  ;
	input \WX9824_reg/NET0131  ;
	input \WX9826_reg/NET0131  ;
	input \WX9828_reg/NET0131  ;
	input \WX9830_reg/NET0131  ;
	input \WX9832_reg/NET0131  ;
	input \WX9834_reg/NET0131  ;
	input \WX9836_reg/NET0131  ;
	input \WX9838_reg/NET0131  ;
	input \WX9840_reg/NET0131  ;
	input \WX9842_reg/NET0131  ;
	input \WX9844_reg/NET0131  ;
	input \WX9846_reg/NET0131  ;
	input \WX9848_reg/NET0131  ;
	input \WX9850_reg/NET0131  ;
	input \WX9852_reg/NET0131  ;
	input \WX9854_reg/NET0131  ;
	input \WX9856_reg/NET0131  ;
	input \WX9858_reg/NET0131  ;
	input \WX9860_reg/NET0131  ;
	input \WX9862_reg/NET0131  ;
	input \WX9864_reg/NET0131  ;
	input \WX9866_reg/NET0131  ;
	input \WX9868_reg/NET0131  ;
	input \WX9870_reg/NET0131  ;
	input \WX9872_reg/NET0131  ;
	input \WX9874_reg/NET0131  ;
	input \WX9876_reg/NET0131  ;
	input \WX9878_reg/NET0131  ;
	input \WX9880_reg/NET0131  ;
	input \WX9882_reg/NET0131  ;
	input \WX9884_reg/NET0131  ;
	input \WX9886_reg/NET0131  ;
	input \WX9888_reg/NET0131  ;
	input \WX9890_reg/NET0131  ;
	input \WX9892_reg/NET0131  ;
	input \WX9894_reg/NET0131  ;
	input \WX9896_reg/NET0131  ;
	input \WX9898_reg/NET0131  ;
	input \WX9900_reg/NET0131  ;
	input \WX9902_reg/NET0131  ;
	input \WX9904_reg/NET0131  ;
	input \WX9906_reg/NET0131  ;
	input \WX9908_reg/NET0131  ;
	input \WX9910_reg/NET0131  ;
	input \WX9912_reg/NET0131  ;
	input \WX9914_reg/NET0131  ;
	input \WX9916_reg/NET0131  ;
	input \WX9918_reg/NET0131  ;
	input \WX9920_reg/NET0131  ;
	input \WX9922_reg/NET0131  ;
	input \WX9924_reg/NET0131  ;
	input \WX9926_reg/NET0131  ;
	input \WX9928_reg/NET0131  ;
	input \WX9930_reg/NET0131  ;
	input \WX9932_reg/NET0131  ;
	input \WX9934_reg/NET0131  ;
	input \WX9936_reg/NET0131  ;
	input \WX9938_reg/NET0131  ;
	input \WX9940_reg/NET0131  ;
	input \WX9942_reg/NET0131  ;
	input \WX9944_reg/NET0131  ;
	input \WX9946_reg/NET0131  ;
	input \WX9948_reg/NET0131  ;
	input \WX9950_reg/NET0131  ;
	input \_2077__reg/NET0131  ;
	input \_2078__reg/NET0131  ;
	input \_2079__reg/NET0131  ;
	input \_2080__reg/NET0131  ;
	input \_2081__reg/NET0131  ;
	input \_2082__reg/NET0131  ;
	input \_2083__reg/NET0131  ;
	input \_2084__reg/NET0131  ;
	input \_2085__reg/NET0131  ;
	input \_2086__reg/NET0131  ;
	input \_2087__reg/NET0131  ;
	input \_2088__reg/NET0131  ;
	input \_2089__reg/NET0131  ;
	input \_2090__reg/NET0131  ;
	input \_2091__reg/NET0131  ;
	input \_2092__reg/NET0131  ;
	input \_2093__reg/NET0131  ;
	input \_2094__reg/NET0131  ;
	input \_2095__reg/NET0131  ;
	input \_2096__reg/NET0131  ;
	input \_2097__reg/NET0131  ;
	input \_2098__reg/NET0131  ;
	input \_2099__reg/NET0131  ;
	input \_2100__reg/NET0131  ;
	input \_2101__reg/NET0131  ;
	input \_2102__reg/NET0131  ;
	input \_2103__reg/NET0131  ;
	input \_2104__reg/NET0131  ;
	input \_2105__reg/NET0131  ;
	input \_2106__reg/NET0131  ;
	input \_2107__reg/NET0131  ;
	input \_2108__reg/NET0131  ;
	input \_2109__reg/NET0131  ;
	input \_2110__reg/NET0131  ;
	input \_2111__reg/NET0131  ;
	input \_2112__reg/NET0131  ;
	input \_2113__reg/NET0131  ;
	input \_2114__reg/NET0131  ;
	input \_2115__reg/NET0131  ;
	input \_2116__reg/NET0131  ;
	input \_2117__reg/NET0131  ;
	input \_2118__reg/NET0131  ;
	input \_2119__reg/NET0131  ;
	input \_2120__reg/NET0131  ;
	input \_2121__reg/NET0131  ;
	input \_2122__reg/NET0131  ;
	input \_2123__reg/NET0131  ;
	input \_2124__reg/NET0131  ;
	input \_2125__reg/NET0131  ;
	input \_2126__reg/NET0131  ;
	input \_2127__reg/NET0131  ;
	input \_2128__reg/NET0131  ;
	input \_2129__reg/NET0131  ;
	input \_2130__reg/NET0131  ;
	input \_2131__reg/NET0131  ;
	input \_2132__reg/NET0131  ;
	input \_2133__reg/NET0131  ;
	input \_2134__reg/NET0131  ;
	input \_2135__reg/NET0131  ;
	input \_2136__reg/NET0131  ;
	input \_2137__reg/NET0131  ;
	input \_2138__reg/NET0131  ;
	input \_2139__reg/NET0131  ;
	input \_2140__reg/NET0131  ;
	input \_2141__reg/NET0131  ;
	input \_2142__reg/NET0131  ;
	input \_2143__reg/NET0131  ;
	input \_2144__reg/NET0131  ;
	input \_2145__reg/NET0131  ;
	input \_2146__reg/NET0131  ;
	input \_2147__reg/NET0131  ;
	input \_2148__reg/NET0131  ;
	input \_2149__reg/NET0131  ;
	input \_2150__reg/NET0131  ;
	input \_2151__reg/NET0131  ;
	input \_2152__reg/NET0131  ;
	input \_2153__reg/NET0131  ;
	input \_2154__reg/NET0131  ;
	input \_2155__reg/NET0131  ;
	input \_2156__reg/NET0131  ;
	input \_2157__reg/NET0131  ;
	input \_2158__reg/NET0131  ;
	input \_2159__reg/NET0131  ;
	input \_2160__reg/NET0131  ;
	input \_2161__reg/NET0131  ;
	input \_2162__reg/NET0131  ;
	input \_2163__reg/NET0131  ;
	input \_2164__reg/NET0131  ;
	input \_2165__reg/NET0131  ;
	input \_2166__reg/NET0131  ;
	input \_2167__reg/NET0131  ;
	input \_2168__reg/NET0131  ;
	input \_2169__reg/NET0131  ;
	input \_2170__reg/NET0131  ;
	input \_2171__reg/NET0131  ;
	input \_2172__reg/NET0131  ;
	input \_2173__reg/NET0131  ;
	input \_2174__reg/NET0131  ;
	input \_2175__reg/NET0131  ;
	input \_2176__reg/NET0131  ;
	input \_2177__reg/NET0131  ;
	input \_2178__reg/NET0131  ;
	input \_2179__reg/NET0131  ;
	input \_2180__reg/NET0131  ;
	input \_2181__reg/NET0131  ;
	input \_2182__reg/NET0131  ;
	input \_2183__reg/NET0131  ;
	input \_2184__reg/NET0131  ;
	input \_2185__reg/NET0131  ;
	input \_2186__reg/NET0131  ;
	input \_2187__reg/NET0131  ;
	input \_2188__reg/NET0131  ;
	input \_2189__reg/NET0131  ;
	input \_2190__reg/NET0131  ;
	input \_2191__reg/NET0131  ;
	input \_2192__reg/NET0131  ;
	input \_2193__reg/NET0131  ;
	input \_2194__reg/NET0131  ;
	input \_2195__reg/NET0131  ;
	input \_2196__reg/NET0131  ;
	input \_2197__reg/NET0131  ;
	input \_2198__reg/NET0131  ;
	input \_2199__reg/NET0131  ;
	input \_2200__reg/NET0131  ;
	input \_2201__reg/NET0131  ;
	input \_2202__reg/NET0131  ;
	input \_2203__reg/NET0131  ;
	input \_2204__reg/NET0131  ;
	input \_2205__reg/NET0131  ;
	input \_2206__reg/NET0131  ;
	input \_2207__reg/NET0131  ;
	input \_2208__reg/NET0131  ;
	input \_2209__reg/NET0131  ;
	input \_2210__reg/NET0131  ;
	input \_2211__reg/NET0131  ;
	input \_2212__reg/NET0131  ;
	input \_2213__reg/NET0131  ;
	input \_2214__reg/NET0131  ;
	input \_2215__reg/NET0131  ;
	input \_2216__reg/NET0131  ;
	input \_2217__reg/NET0131  ;
	input \_2218__reg/NET0131  ;
	input \_2219__reg/NET0131  ;
	input \_2220__reg/NET0131  ;
	input \_2221__reg/NET0131  ;
	input \_2222__reg/NET0131  ;
	input \_2223__reg/NET0131  ;
	input \_2224__reg/NET0131  ;
	input \_2225__reg/NET0131  ;
	input \_2226__reg/NET0131  ;
	input \_2227__reg/NET0131  ;
	input \_2228__reg/NET0131  ;
	input \_2229__reg/NET0131  ;
	input \_2230__reg/NET0131  ;
	input \_2231__reg/NET0131  ;
	input \_2232__reg/NET0131  ;
	input \_2233__reg/NET0131  ;
	input \_2234__reg/NET0131  ;
	input \_2235__reg/NET0131  ;
	input \_2236__reg/NET0131  ;
	input \_2237__reg/NET0131  ;
	input \_2238__reg/NET0131  ;
	input \_2239__reg/NET0131  ;
	input \_2240__reg/NET0131  ;
	input \_2241__reg/NET0131  ;
	input \_2242__reg/NET0131  ;
	input \_2243__reg/NET0131  ;
	input \_2244__reg/NET0131  ;
	input \_2245__reg/NET0131  ;
	input \_2246__reg/NET0131  ;
	input \_2247__reg/NET0131  ;
	input \_2248__reg/NET0131  ;
	input \_2249__reg/NET0131  ;
	input \_2250__reg/NET0131  ;
	input \_2251__reg/NET0131  ;
	input \_2252__reg/NET0131  ;
	input \_2253__reg/NET0131  ;
	input \_2254__reg/NET0131  ;
	input \_2255__reg/NET0131  ;
	input \_2256__reg/NET0131  ;
	input \_2257__reg/NET0131  ;
	input \_2258__reg/NET0131  ;
	input \_2259__reg/NET0131  ;
	input \_2260__reg/NET0131  ;
	input \_2261__reg/NET0131  ;
	input \_2262__reg/NET0131  ;
	input \_2263__reg/NET0131  ;
	input \_2264__reg/NET0131  ;
	input \_2265__reg/NET0131  ;
	input \_2266__reg/NET0131  ;
	input \_2267__reg/NET0131  ;
	input \_2268__reg/NET0131  ;
	input \_2269__reg/NET0131  ;
	input \_2270__reg/NET0131  ;
	input \_2271__reg/NET0131  ;
	input \_2272__reg/NET0131  ;
	input \_2273__reg/NET0131  ;
	input \_2274__reg/NET0131  ;
	input \_2275__reg/NET0131  ;
	input \_2276__reg/NET0131  ;
	input \_2277__reg/NET0131  ;
	input \_2278__reg/NET0131  ;
	input \_2279__reg/NET0131  ;
	input \_2280__reg/NET0131  ;
	input \_2281__reg/NET0131  ;
	input \_2282__reg/NET0131  ;
	input \_2283__reg/NET0131  ;
	input \_2284__reg/NET0131  ;
	input \_2285__reg/NET0131  ;
	input \_2286__reg/NET0131  ;
	input \_2287__reg/NET0131  ;
	input \_2288__reg/NET0131  ;
	input \_2289__reg/NET0131  ;
	input \_2290__reg/NET0131  ;
	input \_2291__reg/NET0131  ;
	input \_2292__reg/NET0131  ;
	input \_2293__reg/NET0131  ;
	input \_2294__reg/NET0131  ;
	input \_2295__reg/NET0131  ;
	input \_2296__reg/NET0131  ;
	input \_2297__reg/NET0131  ;
	input \_2298__reg/NET0131  ;
	input \_2299__reg/NET0131  ;
	input \_2300__reg/NET0131  ;
	input \_2301__reg/NET0131  ;
	input \_2302__reg/NET0131  ;
	input \_2303__reg/NET0131  ;
	input \_2304__reg/NET0131  ;
	input \_2305__reg/NET0131  ;
	input \_2306__reg/NET0131  ;
	input \_2307__reg/NET0131  ;
	input \_2308__reg/NET0131  ;
	input \_2309__reg/NET0131  ;
	input \_2310__reg/NET0131  ;
	input \_2311__reg/NET0131  ;
	input \_2312__reg/NET0131  ;
	input \_2313__reg/NET0131  ;
	input \_2314__reg/NET0131  ;
	input \_2315__reg/NET0131  ;
	input \_2316__reg/NET0131  ;
	input \_2317__reg/NET0131  ;
	input \_2318__reg/NET0131  ;
	input \_2319__reg/NET0131  ;
	input \_2320__reg/NET0131  ;
	input \_2321__reg/NET0131  ;
	input \_2322__reg/NET0131  ;
	input \_2323__reg/NET0131  ;
	input \_2324__reg/NET0131  ;
	input \_2325__reg/NET0131  ;
	input \_2326__reg/NET0131  ;
	input \_2327__reg/NET0131  ;
	input \_2328__reg/NET0131  ;
	input \_2329__reg/NET0131  ;
	input \_2330__reg/NET0131  ;
	input \_2331__reg/NET0131  ;
	input \_2332__reg/NET0131  ;
	input \_2333__reg/NET0131  ;
	input \_2334__reg/NET0131  ;
	input \_2335__reg/NET0131  ;
	input \_2336__reg/NET0131  ;
	input \_2337__reg/NET0131  ;
	input \_2338__reg/NET0131  ;
	input \_2339__reg/NET0131  ;
	input \_2340__reg/NET0131  ;
	input \_2341__reg/NET0131  ;
	input \_2342__reg/NET0131  ;
	input \_2343__reg/NET0131  ;
	input \_2344__reg/NET0131  ;
	input \_2345__reg/NET0131  ;
	input \_2346__reg/NET0131  ;
	input \_2347__reg/NET0131  ;
	input \_2348__reg/NET0131  ;
	input \_2349__reg/NET0131  ;
	input \_2350__reg/NET0131  ;
	input \_2351__reg/NET0131  ;
	input \_2352__reg/NET0131  ;
	input \_2353__reg/NET0131  ;
	input \_2354__reg/NET0131  ;
	input \_2355__reg/NET0131  ;
	input \_2356__reg/NET0131  ;
	input \_2357__reg/NET0131  ;
	input \_2358__reg/NET0131  ;
	input \_2359__reg/NET0131  ;
	input \_2360__reg/NET0131  ;
	input \_2361__reg/NET0131  ;
	input \_2362__reg/NET0131  ;
	input \_2363__reg/NET0131  ;
	input \_2364__reg/NET0131  ;
	output \DATA_9_0_pad  ;
	output \DATA_9_10_pad  ;
	output \DATA_9_11_pad  ;
	output \DATA_9_12_pad  ;
	output \DATA_9_13_pad  ;
	output \DATA_9_14_pad  ;
	output \DATA_9_15_pad  ;
	output \DATA_9_16_pad  ;
	output \DATA_9_17_pad  ;
	output \DATA_9_18_pad  ;
	output \DATA_9_19_pad  ;
	output \DATA_9_1_pad  ;
	output \DATA_9_20_pad  ;
	output \DATA_9_21_pad  ;
	output \DATA_9_22_pad  ;
	output \DATA_9_23_pad  ;
	output \DATA_9_24_pad  ;
	output \DATA_9_25_pad  ;
	output \DATA_9_26_pad  ;
	output \DATA_9_27_pad  ;
	output \DATA_9_28_pad  ;
	output \DATA_9_29_pad  ;
	output \DATA_9_2_pad  ;
	output \DATA_9_30_pad  ;
	output \DATA_9_31_pad  ;
	output \DATA_9_3_pad  ;
	output \DATA_9_4_pad  ;
	output \DATA_9_5_pad  ;
	output \DATA_9_6_pad  ;
	output \DATA_9_7_pad  ;
	output \DATA_9_8_pad  ;
	output \DATA_9_9_pad  ;
	output \_al_n0  ;
	output \_al_n1  ;
	output \g19/_0_  ;
	output \g35/_0_  ;
	output \g36/_0_  ;
	output \g40/_0_  ;
	output \g55780/_0_  ;
	output \g55783/_0_  ;
	output \g55795/_0_  ;
	output \g55796/_0_  ;
	output \g55797/_0_  ;
	output \g55798/_0_  ;
	output \g55799/_0_  ;
	output \g55800/_0_  ;
	output \g55801/_0_  ;
	output \g55802/_0_  ;
	output \g55803/_0_  ;
	output \g55834/_0_  ;
	output \g55835/_0_  ;
	output \g55836/_0_  ;
	output \g55837/_0_  ;
	output \g55838/_0_  ;
	output \g55839/_0_  ;
	output \g55840/_0_  ;
	output \g55841/_0_  ;
	output \g55842/_0_  ;
	output \g55856/_0_  ;
	output \g55894/_0_  ;
	output \g55895/_0_  ;
	output \g55896/_0_  ;
	output \g55897/_0_  ;
	output \g55898/_0_  ;
	output \g55899/_0_  ;
	output \g55900/_0_  ;
	output \g55901/_0_  ;
	output \g55902/_0_  ;
	output \g55916/_0_  ;
	output \g55953/_0_  ;
	output \g55954/_0_  ;
	output \g55955/_0_  ;
	output \g55956/_0_  ;
	output \g55957/_0_  ;
	output \g55958/_0_  ;
	output \g55959/_0_  ;
	output \g55960/_0_  ;
	output \g55961/_0_  ;
	output \g55975/_0_  ;
	output \g56012/_0_  ;
	output \g56013/_0_  ;
	output \g56014/_0_  ;
	output \g56015/_0_  ;
	output \g56016/_0_  ;
	output \g56017/_0_  ;
	output \g56018/_0_  ;
	output \g56019/_0_  ;
	output \g56020/_0_  ;
	output \g56034/_0_  ;
	output \g56071/_0_  ;
	output \g56072/_0_  ;
	output \g56073/_0_  ;
	output \g56074/_0_  ;
	output \g56075/_0_  ;
	output \g56076/_0_  ;
	output \g56077/_0_  ;
	output \g56078/_0_  ;
	output \g56079/_0_  ;
	output \g56093/_0_  ;
	output \g56130/_0_  ;
	output \g56131/_0_  ;
	output \g56132/_0_  ;
	output \g56133/_0_  ;
	output \g56134/_0_  ;
	output \g56135/_0_  ;
	output \g56136/_0_  ;
	output \g56137/_0_  ;
	output \g56138/_0_  ;
	output \g56152/_0_  ;
	output \g56189/_0_  ;
	output \g56190/_0_  ;
	output \g56191/_0_  ;
	output \g56192/_0_  ;
	output \g56193/_0_  ;
	output \g56194/_0_  ;
	output \g56195/_0_  ;
	output \g56196/_0_  ;
	output \g56197/_0_  ;
	output \g56211/_0_  ;
	output \g56248/_0_  ;
	output \g56249/_0_  ;
	output \g56250/_0_  ;
	output \g56251/_0_  ;
	output \g56252/_0_  ;
	output \g56253/_0_  ;
	output \g56254/_0_  ;
	output \g56255/_0_  ;
	output \g56256/_0_  ;
	output \g56270/_0_  ;
	output \g56307/_0_  ;
	output \g56308/_0_  ;
	output \g56309/_0_  ;
	output \g56310/_0_  ;
	output \g56311/_0_  ;
	output \g56312/_0_  ;
	output \g56313/_0_  ;
	output \g56314/_0_  ;
	output \g56315/_0_  ;
	output \g56329/_0_  ;
	output \g56366/_0_  ;
	output \g56367/_0_  ;
	output \g56368/_0_  ;
	output \g56369/_0_  ;
	output \g56370/_0_  ;
	output \g56371/_0_  ;
	output \g56372/_0_  ;
	output \g56373/_0_  ;
	output \g56374/_0_  ;
	output \g56388/_0_  ;
	output \g56425/_0_  ;
	output \g56426/_0_  ;
	output \g56427/_0_  ;
	output \g56428/_0_  ;
	output \g56429/_0_  ;
	output \g56430/_0_  ;
	output \g56431/_0_  ;
	output \g56432/_0_  ;
	output \g56433/_0_  ;
	output \g56447/_0_  ;
	output \g56484/_0_  ;
	output \g56485/_0_  ;
	output \g56486/_0_  ;
	output \g56487/_0_  ;
	output \g56488/_0_  ;
	output \g56489/_0_  ;
	output \g56490/_0_  ;
	output \g56491/_0_  ;
	output \g56492/_0_  ;
	output \g56507/_0_  ;
	output \g56543/_0_  ;
	output \g56544/_0_  ;
	output \g56545/_0_  ;
	output \g56546/_0_  ;
	output \g56547/_0_  ;
	output \g56548/_0_  ;
	output \g56549/_0_  ;
	output \g56551/_0_  ;
	output \g56567/_0_  ;
	output \g56602/_0_  ;
	output \g56603/_0_  ;
	output \g56604/_0_  ;
	output \g56605/_0_  ;
	output \g56606/_0_  ;
	output \g56607/_0_  ;
	output \g56608/_0_  ;
	output \g56610/_0_  ;
	output \g56627/_0_  ;
	output \g56661/_0_  ;
	output \g56662/_0_  ;
	output \g56663/_0_  ;
	output \g56664/_0_  ;
	output \g56665/_0_  ;
	output \g56666/_0_  ;
	output \g56667/_0_  ;
	output \g56668/_0_  ;
	output \g56686/_0_  ;
	output \g56720/_0_  ;
	output \g56721/_0_  ;
	output \g56722/_0_  ;
	output \g56723/_0_  ;
	output \g56724/_0_  ;
	output \g56725/_0_  ;
	output \g56726/_0_  ;
	output \g56727/_0_  ;
	output \g56728/_0_  ;
	output \g56745/_0_  ;
	output \g56779/_0_  ;
	output \g56780/_0_  ;
	output \g56781/_0_  ;
	output \g56782/_0_  ;
	output \g56783/_0_  ;
	output \g56784/_0_  ;
	output \g56785/_0_  ;
	output \g56804/_0_  ;
	output \g56838/_0_  ;
	output \g56839/_0_  ;
	output \g56840/_0_  ;
	output \g56841/_0_  ;
	output \g56842/_0_  ;
	output \g56843/_0_  ;
	output \g56844/_0_  ;
	output \g56845/_0_  ;
	output \g56846/_0_  ;
	output \g56863/_0_  ;
	output \g56897/_0_  ;
	output \g56898/_0_  ;
	output \g56899/_0_  ;
	output \g56900/_0_  ;
	output \g56901/_0_  ;
	output \g56902/_0_  ;
	output \g56903/_0_  ;
	output \g56905/_0_  ;
	output \g56921/_0_  ;
	output \g56956/_0_  ;
	output \g56957/_0_  ;
	output \g56958/_0_  ;
	output \g56959/_0_  ;
	output \g56960/_0_  ;
	output \g56961/_0_  ;
	output \g56962/_0_  ;
	output \g56964/_0_  ;
	output \g56980/_0_  ;
	output \g57015/_0_  ;
	output \g57016/_0_  ;
	output \g57017/_0_  ;
	output \g57018/_0_  ;
	output \g57019/_0_  ;
	output \g57020/_0_  ;
	output \g57021/_0_  ;
	output \g57023/_0_  ;
	output \g57040/_0_  ;
	output \g57074/_0_  ;
	output \g57075/_0_  ;
	output \g57076/_0_  ;
	output \g57077/_0_  ;
	output \g57078/_0_  ;
	output \g57079/_0_  ;
	output \g57080/_0_  ;
	output \g57081/_0_  ;
	output \g57099/_0_  ;
	output \g57133/_0_  ;
	output \g57134/_0_  ;
	output \g57135/_0_  ;
	output \g57136/_0_  ;
	output \g57137/_0_  ;
	output \g57138/_0_  ;
	output \g57139/_0_  ;
	output \g57140/_0_  ;
	output \g57141/_0_  ;
	output \g57159/_0_  ;
	output \g57193/_0_  ;
	output \g57195/_0_  ;
	output \g57196/_0_  ;
	output \g57197/_0_  ;
	output \g57198/_0_  ;
	output \g57199/_0_  ;
	output \g57200/_0_  ;
	output \g57202/_0_  ;
	output \g57219/_0_  ;
	output \g57254/_0_  ;
	output \g57255/_0_  ;
	output \g57256/_0_  ;
	output \g57257/_0_  ;
	output \g57258/_0_  ;
	output \g57259/_0_  ;
	output \g57260/_0_  ;
	output \g57262/_0_  ;
	output \g57263/_0_  ;
	output \g57285/_0_  ;
	output \g57318/_0_  ;
	output \g57319/_0_  ;
	output \g57320/_0_  ;
	output \g57321/_0_  ;
	output \g57322/_0_  ;
	output \g57323/_0_  ;
	output \g57324/_0_  ;
	output \g57325/_0_  ;
	output \g57326/_0_  ;
	output \g57328/_0_  ;
	output \g57329/_0_  ;
	output \g57330/_0_  ;
	output \g57350/_0_  ;
	output \g57387/_0_  ;
	output \g57388/_0_  ;
	output \g57390/_0_  ;
	output \g57391/_0_  ;
	output \g57392/_0_  ;
	output \g57393/_0_  ;
	output \g57395/_0_  ;
	output \g57396/_0_  ;
	output \g57439/_0_  ;
	output \g57476/_0_  ;
	output \g57477/_0_  ;
	output \g57478/_0_  ;
	output \g57479/_0_  ;
	output \g57480/_0_  ;
	output \g57481/_0_  ;
	output \g57482/_0_  ;
	output \g57483/_0_  ;
	output \g57484/_0_  ;
	output \g57485/_0_  ;
	output \g57486/_0_  ;
	output \g57487/_0_  ;
	output \g57488/_0_  ;
	output \g57489/_0_  ;
	output \g57490/_0_  ;
	output \g57491/_0_  ;
	output \g57492/_0_  ;
	output \g57493/_0_  ;
	output \g57494/_0_  ;
	output \g57495/_0_  ;
	output \g57496/_0_  ;
	output \g57497/_0_  ;
	output \g57498/_0_  ;
	output \g57499/_0_  ;
	output \g57500/_0_  ;
	output \g57501/_0_  ;
	output \g57502/_0_  ;
	output \g57503/_0_  ;
	output \g57504/_0_  ;
	output \g57505/_0_  ;
	output \g57524/_0_  ;
	output \g57537/_0_  ;
	output \g57541/_0_  ;
	output \g57543/_0_  ;
	output \g58163/_0_  ;
	output \g58572/_0_  ;
	output \g58573/_0_  ;
	output \g58574/_0_  ;
	output \g58575/_0_  ;
	output \g58576/_0_  ;
	output \g58577/_0_  ;
	output \g58578/_0_  ;
	output \g58579/_0_  ;
	output \g58580/_0_  ;
	output \g58581/_0_  ;
	output \g58582/_0_  ;
	output \g58583/_0_  ;
	output \g58584/_0_  ;
	output \g58585/_0_  ;
	output \g58586/_0_  ;
	output \g58587/_0_  ;
	output \g58588/_0_  ;
	output \g58589/_0_  ;
	output \g58590/_0_  ;
	output \g58591/_0_  ;
	output \g58592/_0_  ;
	output \g58593/_0_  ;
	output \g58594/_0_  ;
	output \g58595/_0_  ;
	output \g58596/_0_  ;
	output \g58597/_0_  ;
	output \g58598/_0_  ;
	output \g58600/_0_  ;
	output \g58602/_0_  ;
	output \g58604/_0_  ;
	output \g58615/_0_  ;
	output \g59240/_0_  ;
	output \g59241/_0_  ;
	output \g59242/_0_  ;
	output \g59243/_0_  ;
	output \g59244/_0_  ;
	output \g59245/_0_  ;
	output \g59246/_0_  ;
	output \g59247/_0_  ;
	output \g59248/_0_  ;
	output \g59249/_0_  ;
	output \g59250/_0_  ;
	output \g59251/_0_  ;
	output \g59252/_0_  ;
	output \g59253/_0_  ;
	output \g59254/_0_  ;
	output \g59255/_0_  ;
	output \g59256/_0_  ;
	output \g59257/_0_  ;
	output \g59258/_0_  ;
	output \g59259/_0_  ;
	output \g59260/_0_  ;
	output \g59261/_0_  ;
	output \g59262/_0_  ;
	output \g59263/_0_  ;
	output \g59264/_0_  ;
	output \g59265/_0_  ;
	output \g59266/_0_  ;
	output \g59267/_0_  ;
	output \g59268/_0_  ;
	output \g59269/_0_  ;
	output \g59270/_0_  ;
	output \g59271/_0_  ;
	output \g59272/_0_  ;
	output \g59273/_0_  ;
	output \g59274/_0_  ;
	output \g59275/_0_  ;
	output \g59276/_0_  ;
	output \g59277/_0_  ;
	output \g59278/_0_  ;
	output \g59279/_0_  ;
	output \g59280/_0_  ;
	output \g59281/_0_  ;
	output \g59282/_0_  ;
	output \g59283/_0_  ;
	output \g59284/_0_  ;
	output \g59285/_0_  ;
	output \g59286/_0_  ;
	output \g59287/_0_  ;
	output \g59288/_0_  ;
	output \g59289/_0_  ;
	output \g59290/_0_  ;
	output \g59291/_0_  ;
	output \g59292/_0_  ;
	output \g59293/_0_  ;
	output \g59294/_0_  ;
	output \g59295/_0_  ;
	output \g59296/_0_  ;
	output \g59297/_0_  ;
	output \g59298/_0_  ;
	output \g59299/_0_  ;
	output \g59300/_0_  ;
	output \g59301/_0_  ;
	output \g59302/_0_  ;
	output \g59303/_0_  ;
	output \g59304/_0_  ;
	output \g59305/_0_  ;
	output \g59306/_0_  ;
	output \g59307/_0_  ;
	output \g59308/_0_  ;
	output \g59309/_0_  ;
	output \g59310/_0_  ;
	output \g59311/_0_  ;
	output \g59312/_0_  ;
	output \g59313/_0_  ;
	output \g59314/_0_  ;
	output \g59315/_0_  ;
	output \g59316/_0_  ;
	output \g59317/_0_  ;
	output \g59318/_0_  ;
	output \g59319/_0_  ;
	output \g59320/_0_  ;
	output \g59321/_0_  ;
	output \g59322/_0_  ;
	output \g59323/_0_  ;
	output \g59324/_0_  ;
	output \g59325/_0_  ;
	output \g59326/_0_  ;
	output \g59327/_0_  ;
	output \g59328/_0_  ;
	output \g59329/_0_  ;
	output \g59330/_0_  ;
	output \g59331/_0_  ;
	output \g59332/_0_  ;
	output \g59333/_0_  ;
	output \g59334/_0_  ;
	output \g59335/_0_  ;
	output \g59336/_0_  ;
	output \g59337/_0_  ;
	output \g59338/_0_  ;
	output \g59339/_0_  ;
	output \g59340/_0_  ;
	output \g59341/_0_  ;
	output \g59342/_0_  ;
	output \g59343/_0_  ;
	output \g59344/_0_  ;
	output \g59345/_0_  ;
	output \g59346/_0_  ;
	output \g59347/_0_  ;
	output \g59348/_0_  ;
	output \g59349/_0_  ;
	output \g59350/_0_  ;
	output \g59351/_0_  ;
	output \g59352/_0_  ;
	output \g59353/_0_  ;
	output \g59354/_0_  ;
	output \g59355/_0_  ;
	output \g59356/_0_  ;
	output \g59357/_0_  ;
	output \g59358/_0_  ;
	output \g59359/_0_  ;
	output \g59360/_0_  ;
	output \g59361/_0_  ;
	output \g59362/_0_  ;
	output \g59363/_0_  ;
	output \g59364/_0_  ;
	output \g59365/_0_  ;
	output \g59366/_0_  ;
	output \g59367/_0_  ;
	output \g59368/_0_  ;
	output \g59369/_0_  ;
	output \g59370/_0_  ;
	output \g59371/_0_  ;
	output \g59372/_0_  ;
	output \g59373/_0_  ;
	output \g59374/_0_  ;
	output \g59375/_0_  ;
	output \g59376/_0_  ;
	output \g59377/_0_  ;
	output \g59378/_0_  ;
	output \g59379/_0_  ;
	output \g59380/_0_  ;
	output \g59381/_0_  ;
	output \g59382/_0_  ;
	output \g59383/_0_  ;
	output \g59384/_0_  ;
	output \g59385/_0_  ;
	output \g59386/_0_  ;
	output \g59387/_0_  ;
	output \g59388/_0_  ;
	output \g59389/_0_  ;
	output \g59390/_0_  ;
	output \g59391/_0_  ;
	output \g59392/_0_  ;
	output \g59393/_0_  ;
	output \g59394/_0_  ;
	output \g59395/_0_  ;
	output \g59396/_0_  ;
	output \g59397/_0_  ;
	output \g59398/_0_  ;
	output \g59399/_0_  ;
	output \g59400/_0_  ;
	output \g59401/_0_  ;
	output \g59402/_0_  ;
	output \g59403/_0_  ;
	output \g59404/_0_  ;
	output \g59405/_0_  ;
	output \g59406/_0_  ;
	output \g59407/_0_  ;
	output \g59408/_0_  ;
	output \g59409/_0_  ;
	output \g59410/_0_  ;
	output \g59411/_0_  ;
	output \g59412/_0_  ;
	output \g59413/_0_  ;
	output \g59414/_0_  ;
	output \g59415/_0_  ;
	output \g59416/_0_  ;
	output \g59417/_0_  ;
	output \g59418/_0_  ;
	output \g59419/_0_  ;
	output \g59420/_0_  ;
	output \g59421/_0_  ;
	output \g59422/_0_  ;
	output \g59423/_0_  ;
	output \g59424/_0_  ;
	output \g59425/_0_  ;
	output \g59426/_0_  ;
	output \g59427/_0_  ;
	output \g59428/_0_  ;
	output \g59429/_0_  ;
	output \g59430/_0_  ;
	output \g59431/_0_  ;
	output \g59432/_0_  ;
	output \g59433/_0_  ;
	output \g59434/_0_  ;
	output \g59435/_0_  ;
	output \g59436/_0_  ;
	output \g59437/_0_  ;
	output \g59438/_0_  ;
	output \g59439/_0_  ;
	output \g59440/_0_  ;
	output \g59441/_0_  ;
	output \g59442/_0_  ;
	output \g59443/_0_  ;
	output \g59444/_0_  ;
	output \g59445/_0_  ;
	output \g59446/_0_  ;
	output \g59447/_0_  ;
	output \g59448/_0_  ;
	output \g59449/_0_  ;
	output \g59450/_0_  ;
	output \g59451/_0_  ;
	output \g59452/_0_  ;
	output \g59453/_0_  ;
	output \g59454/_0_  ;
	output \g59455/_0_  ;
	output \g59456/_0_  ;
	output \g59457/_0_  ;
	output \g59458/_0_  ;
	output \g59459/_0_  ;
	output \g59460/_0_  ;
	output \g59461/_0_  ;
	output \g59462/_0_  ;
	output \g59463/_0_  ;
	output \g59464/_0_  ;
	output \g59465/_0_  ;
	output \g59466/_0_  ;
	output \g59467/_0_  ;
	output \g59468/_0_  ;
	output \g59469/_0_  ;
	output \g59470/_0_  ;
	output \g59471/_0_  ;
	output \g59472/_0_  ;
	output \g59473/_0_  ;
	output \g59474/_0_  ;
	output \g59475/_0_  ;
	output \g59476/_0_  ;
	output \g59477/_0_  ;
	output \g59478/_0_  ;
	output \g59479/_0_  ;
	output \g59480/_0_  ;
	output \g59481/_0_  ;
	output \g59482/_0_  ;
	output \g59483/_0_  ;
	output \g59484/_0_  ;
	output \g59485/_0_  ;
	output \g59486/_0_  ;
	output \g59487/_0_  ;
	output \g59488/_0_  ;
	output \g59489/_0_  ;
	output \g59490/_0_  ;
	output \g59491/_0_  ;
	output \g59492/_0_  ;
	output \g59493/_0_  ;
	output \g59494/_0_  ;
	output \g59495/_0_  ;
	output \g59496/_0_  ;
	output \g59497/_0_  ;
	output \g59498/_0_  ;
	output \g59500/_0_  ;
	output \g59503/_0_  ;
	output \g59512/_0_  ;
	output \g61336/_0_  ;
	output \g61521/_0_  ;
	output \g61523/_0_  ;
	output \g61524/_0_  ;
	output \g61526/_0_  ;
	output \g61527/_0_  ;
	output \g61528/_0_  ;
	output \g61529/_0_  ;
	output \g61530/_0_  ;
	output \g61531/_0_  ;
	output \g61532/_0_  ;
	output \g61533/_0_  ;
	output \g61535/_0_  ;
	output \g61537/_0_  ;
	output \g61539/_0_  ;
	output \g61540/_0_  ;
	output \g61541/_0_  ;
	output \g61542/_0_  ;
	output \g61546/_0_  ;
	output \g61550/_0_  ;
	output \g61551/_0_  ;
	output \g61552/_0_  ;
	output \g61554/_0_  ;
	output \g61555/_0_  ;
	output \g61556/_0_  ;
	output \g61558/_0_  ;
	output \g61559/_0_  ;
	output \g61561/_0_  ;
	output \g61562/_0_  ;
	output \g61563/_0_  ;
	output \g61564/_0_  ;
	output \g61565/_0_  ;
	output \g61566/_0_  ;
	output \g61568/_0_  ;
	output \g61570/_0_  ;
	output \g61571/_0_  ;
	output \g61572/_0_  ;
	output \g61573/_0_  ;
	output \g61577/_0_  ;
	output \g61578/_0_  ;
	output \g61579/_0_  ;
	output \g61580/_0_  ;
	output \g61581/_0_  ;
	output \g61582/_0_  ;
	output \g61583/_0_  ;
	output \g61584/_0_  ;
	output \g61585/_0_  ;
	output \g61586/_0_  ;
	output \g61587/_0_  ;
	output \g61588/_0_  ;
	output \g61589/_0_  ;
	output \g61591/_0_  ;
	output \g61592/_0_  ;
	output \g61594/_0_  ;
	output \g61595/_0_  ;
	output \g61596/_0_  ;
	output \g61597/_0_  ;
	output \g61598/_0_  ;
	output \g61599/_0_  ;
	output \g61600/_0_  ;
	output \g61601/_0_  ;
	output \g61605/_0_  ;
	output \g61606/_0_  ;
	output \g61607/_0_  ;
	output \g61608/_0_  ;
	output \g61609/_0_  ;
	output \g61610/_0_  ;
	output \g61611/_0_  ;
	output \g61612/_0_  ;
	output \g61613/_0_  ;
	output \g61615/_0_  ;
	output \g61616/_0_  ;
	output \g61617/_0_  ;
	output \g61618/_0_  ;
	output \g61619/_0_  ;
	output \g61620/_0_  ;
	output \g61621/_0_  ;
	output \g61623/_0_  ;
	output \g61624/_0_  ;
	output \g61625/_0_  ;
	output \g61626/_0_  ;
	output \g61627/_0_  ;
	output \g61629/_0_  ;
	output \g61630/_0_  ;
	output \g61631/_0_  ;
	output \g61632/_0_  ;
	output \g61633/_0_  ;
	output \g61634/_0_  ;
	output \g61636/_0_  ;
	output \g61638/_0_  ;
	output \g61639/_0_  ;
	output \g61640/_0_  ;
	output \g61641/_0_  ;
	output \g61642/_0_  ;
	output \g61644/_0_  ;
	output \g61647/_0_  ;
	output \g61648/_0_  ;
	output \g61649/_0_  ;
	output \g61650/_0_  ;
	output \g61653/_0_  ;
	output \g61654/_0_  ;
	output \g61655/_0_  ;
	output \g61656/_0_  ;
	output \g61658/_0_  ;
	output \g61661/_0_  ;
	output \g61662/_0_  ;
	output \g61663/_0_  ;
	output \g61664/_0_  ;
	output \g61666/_0_  ;
	output \g61667/_0_  ;
	output \g61668/_0_  ;
	output \g61670/_0_  ;
	output \g61671/_0_  ;
	output \g61672/_0_  ;
	output \g61673/_0_  ;
	output \g61675/_0_  ;
	output \g61676/_0_  ;
	output \g61680/_0_  ;
	output \g61681/_0_  ;
	output \g61682/_0_  ;
	output \g61683/_0_  ;
	output \g61684/_0_  ;
	output \g61686/_0_  ;
	output \g61687/_0_  ;
	output \g61688/_0_  ;
	output \g61689/_0_  ;
	output \g61690/_0_  ;
	output \g61691/_0_  ;
	output \g61693/_0_  ;
	output \g61694/_0_  ;
	output \g61696/_0_  ;
	output \g61697/_0_  ;
	output \g61698/_0_  ;
	output \g61699/_0_  ;
	output \g61700/_0_  ;
	output \g61701/_0_  ;
	output \g61702/_0_  ;
	output \g61703/_0_  ;
	output \g61704/_0_  ;
	output \g61705/_0_  ;
	output \g61706/_0_  ;
	output \g61707/_0_  ;
	output \g61708/_0_  ;
	output \g61711/_0_  ;
	output \g61712/_0_  ;
	output \g61714/_0_  ;
	output \g61716/_0_  ;
	output \g61717/_0_  ;
	output \g61719/_0_  ;
	output \g61720/_0_  ;
	output \g61721/_0_  ;
	output \g61724/_0_  ;
	output \g61725/_0_  ;
	output \g61728/_0_  ;
	output \g61729/_0_  ;
	output \g61731/_0_  ;
	output \g61732/_0_  ;
	output \g61733/_0_  ;
	output \g61736/_0_  ;
	output \g61737/_0_  ;
	output \g61739/_0_  ;
	output \g61740/_0_  ;
	output \g61741/_0_  ;
	output \g61743/_0_  ;
	output \g61744/_0_  ;
	output \g61745/_0_  ;
	output \g61746/_0_  ;
	output \g61747/_0_  ;
	output \g61748/_0_  ;
	output \g61749/_0_  ;
	output \g61750/_0_  ;
	output \g61751/_0_  ;
	output \g61752/_0_  ;
	output \g61753/_0_  ;
	output \g61754/_0_  ;
	output \g61755/_0_  ;
	output \g61757/_0_  ;
	output \g61758/_0_  ;
	output \g61759/_0_  ;
	output \g61760/_0_  ;
	output \g61761/_0_  ;
	output \g61762/_0_  ;
	output \g61763/_0_  ;
	output \g61764/_0_  ;
	output \g61765/_0_  ;
	output \g61766/_0_  ;
	output \g61767/_0_  ;
	output \g61768/_0_  ;
	output \g61769/_0_  ;
	output \g61770/_0_  ;
	output \g61771/_0_  ;
	output \g61772/_0_  ;
	output \g61773/_0_  ;
	output \g61774/_0_  ;
	output \g61775/_0_  ;
	output \g61776/_0_  ;
	output \g61777/_0_  ;
	output \g61778/_0_  ;
	output \g61780/_0_  ;
	output \g61781/_0_  ;
	output \g61783/_0_  ;
	output \g61784/_0_  ;
	output \g61786/_0_  ;
	output \g61787/_0_  ;
	output \g61790/_0_  ;
	output \g61791/_0_  ;
	output \g61794/_0_  ;
	output \g61795/_0_  ;
	output \g61796/_0_  ;
	output \g61797/_0_  ;
	output \g61798/_0_  ;
	output \g61799/_0_  ;
	output \g61800/_0_  ;
	output \g61801/_0_  ;
	output \g61802/_0_  ;
	output \g61803/_0_  ;
	output \g61805/_0_  ;
	output \g61806/_0_  ;
	output \g61807/_0_  ;
	output \g61808/_0_  ;
	output \g61809/_0_  ;
	output \g61810/_0_  ;
	output \g61811/_0_  ;
	output \g61812/_0_  ;
	output \g61813/_0_  ;
	output \g61816/_0_  ;
	output \g61817/_0_  ;
	output \g61818/_0_  ;
	output \g61820/_0_  ;
	output \g61822/_0_  ;
	output \g61823/_0_  ;
	output \g61825/_0_  ;
	output \g61826/_0_  ;
	output \g61827/_0_  ;
	output \g61828/_0_  ;
	output \g61829/_0_  ;
	output \g61832/_0_  ;
	output \g61834/_0_  ;
	output \g61835/_0_  ;
	output \g61837/_0_  ;
	output \g61838/_0_  ;
	output \g61839/_0_  ;
	output \g61840/_0_  ;
	output \g61844/_0_  ;
	output \g61847/_0_  ;
	output \g61848/_0_  ;
	output \g61849/_0_  ;
	output \g61850/_0_  ;
	output \g61851/_0_  ;
	output \g61853/_0_  ;
	output \g61854/_0_  ;
	output \g61855/_0_  ;
	output \g61856/_0_  ;
	output \g61858/_0_  ;
	output \g61859/_0_  ;
	output \g61861/_0_  ;
	output \g61862/_0_  ;
	output \g61863/_0_  ;
	output \g61864/_0_  ;
	output \g61865/_0_  ;
	output \g61866/_0_  ;
	output \g61867/_0_  ;
	output \g61868/_0_  ;
	output \g61869/_0_  ;
	output \g61870/_0_  ;
	output \g61871/_0_  ;
	output \g61873/_0_  ;
	output \g61874/_0_  ;
	output \g61875/_0_  ;
	output \g61877/_0_  ;
	output \g61878/_0_  ;
	output \g61879/_0_  ;
	output \g61880/_0_  ;
	output \g61881/_0_  ;
	output \g61883/_0_  ;
	output \g61884/_0_  ;
	output \g61886/_0_  ;
	output \g61887/_0_  ;
	output \g61890/_0_  ;
	output \g61891/_0_  ;
	output \g61892/_0_  ;
	output \g61893/_0_  ;
	output \g61894/_0_  ;
	output \g61895/_0_  ;
	output \g61900/_0_  ;
	output \g61901/_0_  ;
	output \g61902/_0_  ;
	output \g61904/_0_  ;
	output \g61905/_0_  ;
	output \g61906/_0_  ;
	output \g61907/_0_  ;
	output \g61914/_0_  ;
	output \g61915/_0_  ;
	output \g61917/_0_  ;
	output \g61919/_0_  ;
	output \g61921/_0_  ;
	output \g61924/_0_  ;
	output \g61925/_0_  ;
	output \g61926/_0_  ;
	output \g61927/_0_  ;
	output \g61928/_0_  ;
	output \g61929/_0_  ;
	output \g61930/_0_  ;
	output \g61931/_0_  ;
	output \g61932/_0_  ;
	output \g61933/_0_  ;
	output \g61934/_0_  ;
	output \g61935/_0_  ;
	output \g61936/_0_  ;
	output \g61937/_0_  ;
	output \g61938/_0_  ;
	output \g61939/_0_  ;
	output \g61943/_0_  ;
	output \g61944/_0_  ;
	output \g61945/_0_  ;
	output \g61947/_0_  ;
	output \g61948/_0_  ;
	output \g61949/_0_  ;
	output \g61950/_0_  ;
	output \g61951/_0_  ;
	output \g61952/_0_  ;
	output \g61953/_0_  ;
	output \g61955/_0_  ;
	output \g61956/_0_  ;
	output \g61957/_0_  ;
	output \g61958/_0_  ;
	output \g61959/_0_  ;
	output \g61960/_0_  ;
	output \g61961/_0_  ;
	output \g61962/_0_  ;
	output \g61963/_0_  ;
	output \g61964/_0_  ;
	output \g61965/_0_  ;
	output \g61966/_0_  ;
	output \g61967/_0_  ;
	output \g61968/_0_  ;
	output \g61969/_0_  ;
	output \g61970/_0_  ;
	output \g61971/_0_  ;
	output \g61972/_0_  ;
	output \g61973/_0_  ;
	output \g61974/_0_  ;
	output \g61976/_0_  ;
	output \g61978/_0_  ;
	output \g61980/_0_  ;
	output \g61981/_0_  ;
	output \g61982/_0_  ;
	output \g61983/_0_  ;
	output \g61984/_0_  ;
	output \g61985/_0_  ;
	output \g61986/_0_  ;
	output \g61987/_0_  ;
	output \g61988/_0_  ;
	output \g61989/_0_  ;
	output \g61990/_0_  ;
	output \g61992/_0_  ;
	output \g61994/_0_  ;
	output \g61995/_0_  ;
	output \g61996/_0_  ;
	output \g61997/_0_  ;
	output \g61998/_0_  ;
	output \g62000/_0_  ;
	output \g62001/_0_  ;
	output \g62002/_0_  ;
	output \g62003/_0_  ;
	output \g62004/_0_  ;
	output \g62005/_0_  ;
	output \g62007/_0_  ;
	output \g62008/_0_  ;
	output \g62009/_0_  ;
	output \g62010/_0_  ;
	output \g62011/_0_  ;
	output \g62012/_0_  ;
	output \g62013/_0_  ;
	output \g62014/_0_  ;
	output \g62015/_0_  ;
	output \g62016/_0_  ;
	output \g62017/_0_  ;
	output \g62018/_0_  ;
	output \g62019/_0_  ;
	output \g62020/_0_  ;
	output \g62021/_0_  ;
	output \g62022/_0_  ;
	output \g62023/_0_  ;
	output \g62024/_0_  ;
	output \g62025/_0_  ;
	output \g62026/_0_  ;
	output \g62027/_0_  ;
	output \g62030/_0_  ;
	output \g62033/_0_  ;
	output \g62034/_0_  ;
	output \g62036/_0_  ;
	output \g62038/_0_  ;
	output \g62041/_0_  ;
	output \g62042/_0_  ;
	output \g62043/_0_  ;
	output \g62044/_0_  ;
	output \g62045/_0_  ;
	output \g62046/_0_  ;
	output \g62047/_0_  ;
	output \g62048/_0_  ;
	output \g62050/_0_  ;
	output \g62051/_0_  ;
	output \g62052/_0_  ;
	output \g62055/_0_  ;
	output \g62057/_0_  ;
	output \g62058/_0_  ;
	output \g62059/_0_  ;
	output \g62060/_0_  ;
	output \g62061/_0_  ;
	output \g62062/_0_  ;
	output \g62064/_0_  ;
	output \g62065/_0_  ;
	output \g62066/_0_  ;
	output \g62067/_0_  ;
	output \g62068/_0_  ;
	output \g62072/_0_  ;
	output \g62073/_0_  ;
	output \g62074/_0_  ;
	output \g62075/_0_  ;
	output \g62076/_0_  ;
	output \g62077/_0_  ;
	output \g62078/_0_  ;
	output \g62080/_0_  ;
	output \g62081/_0_  ;
	output \g62082/_0_  ;
	output \g62084/_0_  ;
	output \g62085/_0_  ;
	output \g62086/_0_  ;
	output \g62087/_0_  ;
	output \g62088/_0_  ;
	output \g62089/_0_  ;
	output \g62090/_0_  ;
	output \g62091/_0_  ;
	output \g62092/_0_  ;
	output \g62094/_0_  ;
	output \g62096/_0_  ;
	output \g62097/_0_  ;
	output \g62098/_0_  ;
	output \g62099/_0_  ;
	output \g62100/_0_  ;
	output \g62101/_0_  ;
	output \g62102/_0_  ;
	output \g62104/_0_  ;
	output \g62106/_0_  ;
	output \g62107/_0_  ;
	output \g62108/_0_  ;
	output \g62110/_0_  ;
	output \g62112/_0_  ;
	output \g62113/_0_  ;
	output \g62114/_0_  ;
	output \g62116/_0_  ;
	output \g62117/_0_  ;
	output \g62118/_0_  ;
	output \g62119/_0_  ;
	output \g62120/_0_  ;
	output \g62121/_0_  ;
	output \g62122/_0_  ;
	output \g62124/_0_  ;
	output \g62126/_0_  ;
	output \g62127/_0_  ;
	output \g62128/_0_  ;
	output \g62129/_0_  ;
	output \g62130/_0_  ;
	output \g62131/_0_  ;
	output \g62132/_0_  ;
	output \g62133/_0_  ;
	output \g62135/_0_  ;
	output \g62136/_0_  ;
	output \g62137/_0_  ;
	output \g62138/_0_  ;
	output \g62140/_0_  ;
	output \g62143/_0_  ;
	output \g62144/_0_  ;
	output \g62149/_0_  ;
	output \g62150/_0_  ;
	output \g62151/_0_  ;
	output \g62153/_0_  ;
	output \g62155/_0_  ;
	output \g62156/_0_  ;
	output \g62158/_0_  ;
	output \g62160/_0_  ;
	output \g62161/_0_  ;
	output \g62162/_0_  ;
	output \g62164/_0_  ;
	output \g62165/_0_  ;
	output \g62166/_0_  ;
	output \g62167/_0_  ;
	output \g62168/_0_  ;
	output \g62169/_0_  ;
	output \g62172/_0_  ;
	output \g62173/_0_  ;
	output \g62175/_0_  ;
	output \g62176/_0_  ;
	output \g62177/_0_  ;
	output \g62178/_0_  ;
	output \g62179/_0_  ;
	output \g62180/_0_  ;
	output \g62181/_0_  ;
	output \g62182/_0_  ;
	output \g62183/_0_  ;
	output \g62184/_0_  ;
	output \g62185/_0_  ;
	output \g62186/_0_  ;
	output \g62188/_0_  ;
	output \g62189/_0_  ;
	output \g62190/_0_  ;
	output \g62191/_0_  ;
	output \g62193/_0_  ;
	output \g62194/_0_  ;
	output \g62195/_0_  ;
	output \g62196/_0_  ;
	output \g62197/_0_  ;
	output \g62200/_0_  ;
	output \g62201/_0_  ;
	output \g62202/_0_  ;
	output \g62203/_0_  ;
	output \g62205/_0_  ;
	output \g62206/_0_  ;
	output \g62207/_0_  ;
	output \g62208/_0_  ;
	output \g62209/_0_  ;
	output \g62210/_0_  ;
	output \g62211/_0_  ;
	output \g62215/_0_  ;
	output \g62218/_0_  ;
	output \g62219/_0_  ;
	output \g62221/_0_  ;
	output \g62222/_0_  ;
	output \g62223/_0_  ;
	output \g62224/_0_  ;
	output \g62225/_0_  ;
	output \g62226/_0_  ;
	output \g62229/_0_  ;
	output \g62230/_0_  ;
	output \g62231/_0_  ;
	output \g62233/_0_  ;
	output \g62236/_0_  ;
	output \g62237/_0_  ;
	output \g62238/_0_  ;
	output \g62240/_0_  ;
	output \g62241/_0_  ;
	output \g62243/_0_  ;
	output \g62244/_0_  ;
	output \g62245/_0_  ;
	output \g62247/_0_  ;
	output \g62248/_0_  ;
	output \g62250/_0_  ;
	output \g62252/_0_  ;
	output \g62253/_0_  ;
	output \g62255/_0_  ;
	output \g62256/_0_  ;
	output \g62257/_0_  ;
	output \g62258/_0_  ;
	output \g62259/_0_  ;
	output \g62260/_0_  ;
	output \g62261/_0_  ;
	output \g62262/_0_  ;
	output \g62263/_0_  ;
	output \g62264/_0_  ;
	output \g62265/_0_  ;
	output \g62267/_0_  ;
	output \g62269/_0_  ;
	output \g62270/_0_  ;
	output \g62272/_0_  ;
	output \g62274/_0_  ;
	output \g62277/_0_  ;
	output \g62279/_0_  ;
	output \g62280/_0_  ;
	output \g62281/_0_  ;
	output \g62283/_0_  ;
	output \g62284/_0_  ;
	output \g62285/_0_  ;
	output \g62286/_0_  ;
	output \g62288/_0_  ;
	output \g62289/_0_  ;
	output \g62290/_0_  ;
	output \g62294/_0_  ;
	output \g62295/_0_  ;
	output \g62296/_0_  ;
	output \g62297/_0_  ;
	output \g62298/_0_  ;
	output \g62299/_0_  ;
	output \g62303/_0_  ;
	output \g62305/_0_  ;
	output \g62306/_0_  ;
	output \g62307/_0_  ;
	output \g62309/_0_  ;
	output \g62311/_0_  ;
	output \g62312/_0_  ;
	output \g62313/_0_  ;
	output \g62314/_0_  ;
	output \g62315/_0_  ;
	output \g62316/_0_  ;
	output \g62317/_0_  ;
	output \g62318/_0_  ;
	output \g62319/_0_  ;
	output \g62320/_0_  ;
	output \g62322/_0_  ;
	output \g62324/_0_  ;
	output \g62325/_0_  ;
	output \g62326/_0_  ;
	output \g62327/_0_  ;
	output \g62329/_0_  ;
	output \g62330/_0_  ;
	output \g62331/_0_  ;
	output \g62332/_0_  ;
	output \g62333/_0_  ;
	output \g62335/_0_  ;
	output \g62336/_0_  ;
	output \g62338/_0_  ;
	output \g62341/_0_  ;
	output \g62342/_0_  ;
	output \g62344/_0_  ;
	output \g62345/_0_  ;
	output \g62348/_0_  ;
	output \g62349/_0_  ;
	output \g62350/_0_  ;
	output \g62353/_0_  ;
	output \g62354/_0_  ;
	output \g62355/_0_  ;
	output \g62356/_0_  ;
	output \g62359/_0_  ;
	output \g62362/_0_  ;
	output \g62363/_0_  ;
	output \g62364/_0_  ;
	output \g62365/_0_  ;
	output \g62366/_0_  ;
	output \g62367/_0_  ;
	output \g62368/_0_  ;
	output \g62369/_0_  ;
	output \g62370/_0_  ;
	output \g62371/_0_  ;
	output \g62372/_0_  ;
	output \g62373/_0_  ;
	output \g62374/_0_  ;
	output \g62376/_0_  ;
	output \g62467/_0_  ;
	output \g62468/_0_  ;
	output \g62469/_0_  ;
	output \g62470/_0_  ;
	output \g62471/_0_  ;
	output \g62472/_0_  ;
	output \g62473/_0_  ;
	output \g62474/_0_  ;
	output \g62475/_0_  ;
	output \g62478/_0_  ;
	output \g62480/_0_  ;
	output \g62481/_0_  ;
	output \g62482/_0_  ;
	output \g62483/_0_  ;
	output \g62484/_0_  ;
	output \g62485/_0_  ;
	output \g62486/_0_  ;
	output \g62487/_0_  ;
	output \g62488/_0_  ;
	output \g62489/_0_  ;
	output \g62490/_0_  ;
	output \g62491/_0_  ;
	output \g62492/_0_  ;
	output \g62493/_0_  ;
	output \g62494/_0_  ;
	output \g62495/_0_  ;
	output \g62496/_0_  ;
	output \g62497/_0_  ;
	output \g62498/_0_  ;
	output \g62499/_0_  ;
	output \g62500/_0_  ;
	output \g62501/_0_  ;
	output \g62502/_0_  ;
	output \g62503/_0_  ;
	output \g62504/_0_  ;
	output \g62509/_0_  ;
	output \g62510/_0_  ;
	output \g62511/_0_  ;
	output \g62512/_0_  ;
	output \g62513/_0_  ;
	output \g62514/_0_  ;
	output \g62515/_0_  ;
	output \g62516/_0_  ;
	output \g62517/_0_  ;
	output \g62518/_0_  ;
	output \g62519/_0_  ;
	output \g62520/_0_  ;
	output \g62521/_0_  ;
	output \g62523/_0_  ;
	output \g62526/_0_  ;
	output \g62528/_0_  ;
	output \g62529/_0_  ;
	output \g62531/_0_  ;
	output \g62532/_0_  ;
	output \g62533/_0_  ;
	output \g62534/_0_  ;
	output \g62535/_0_  ;
	output \g62536/_0_  ;
	output \g62537/_0_  ;
	output \g62539/_0_  ;
	output \g62540/_0_  ;
	output \g62541/_0_  ;
	output \g62542/_0_  ;
	output \g62543/_0_  ;
	output \g62544/_0_  ;
	output \g62545/_0_  ;
	output \g62547/_0_  ;
	output \g62548/_0_  ;
	output \g62549/_0_  ;
	output \g62550/_0_  ;
	output \g62551/_0_  ;
	output \g62552/_0_  ;
	output \g62553/_0_  ;
	output \g62554/_0_  ;
	output \g62555/_0_  ;
	output \g62556/_0_  ;
	output \g62557/_0_  ;
	output \g62560/_0_  ;
	output \g62562/_0_  ;
	output \g62563/_0_  ;
	output \g62564/_0_  ;
	output \g62565/_0_  ;
	output \g62566/_0_  ;
	output \g62567/_0_  ;
	output \g62569/_0_  ;
	output \g62570/_0_  ;
	output \g62571/_0_  ;
	output \g62572/_0_  ;
	output \g62573/_0_  ;
	output \g62574/_0_  ;
	output \g62576/_0_  ;
	output \g62577/_0_  ;
	output \g62581/_0_  ;
	output \g62582/_0_  ;
	output \g62584/_0_  ;
	output \g62585/_0_  ;
	output \g62586/_0_  ;
	output \g62588/_0_  ;
	output \g62589/_0_  ;
	output \g62593/_0_  ;
	output \g62594/_0_  ;
	output \g62595/_0_  ;
	output \g62596/_0_  ;
	output \g62597/_0_  ;
	output \g62598/_0_  ;
	output \g62599/_0_  ;
	output \g62600/_0_  ;
	output \g62601/_0_  ;
	output \g62602/_0_  ;
	output \g62603/_0_  ;
	output \g62604/_0_  ;
	output \g62605/_0_  ;
	output \g62606/_0_  ;
	output \g62607/_0_  ;
	output \g62608/_0_  ;
	output \g62609/_0_  ;
	output \g62610/_0_  ;
	output \g62612/_0_  ;
	output \g62613/_0_  ;
	output \g62614/_0_  ;
	output \g62615/_0_  ;
	output \g62617/_0_  ;
	output \g62618/_0_  ;
	output \g62620/_0_  ;
	output \g62621/_0_  ;
	output \g62622/_0_  ;
	output \g62624/_0_  ;
	output \g62625/_0_  ;
	output \g62626/_0_  ;
	output \g62627/_0_  ;
	output \g62629/_0_  ;
	output \g62630/_0_  ;
	output \g62632/_0_  ;
	output \g62633/_0_  ;
	output \g62635/_0_  ;
	output \g62636/_0_  ;
	output \g62637/_0_  ;
	output \g62638/_0_  ;
	output \g62640/_0_  ;
	output \g62641/_0_  ;
	output \g62642/_0_  ;
	output \g62643/_0_  ;
	output \g62644/_0_  ;
	output \g62646/_0_  ;
	output \g62647/_0_  ;
	output \g62649/_0_  ;
	output \g62650/_0_  ;
	output \g62651/_0_  ;
	output \g62653/_0_  ;
	output \g62655/_0_  ;
	output \g62656/_0_  ;
	output \g62657/_0_  ;
	output \g62658/_0_  ;
	output \g62660/_0_  ;
	output \g62661/_0_  ;
	output \g62662/_0_  ;
	output \g62663/_0_  ;
	output \g62664/_0_  ;
	output \g62665/_0_  ;
	output \g62667/_0_  ;
	output \g62669/_0_  ;
	output \g62670/_0_  ;
	output \g62671/_0_  ;
	output \g62672/_0_  ;
	output \g62674/_0_  ;
	output \g62675/_0_  ;
	output \g62676/_0_  ;
	output \g62677/_0_  ;
	output \g62678/_0_  ;
	output \g62679/_0_  ;
	output \g62680/_0_  ;
	output \g62681/_0_  ;
	output \g62682/_0_  ;
	output \g62684/_0_  ;
	output \g62685/_0_  ;
	output \g62686/_0_  ;
	output \g62687/_0_  ;
	output \g62690/_0_  ;
	output \g62693/_0_  ;
	output \g62698/_0_  ;
	output \g62699/_0_  ;
	output \g62700/_0_  ;
	output \g62701/_0_  ;
	output \g62702/_0_  ;
	output \g62703/_0_  ;
	output \g62704/_0_  ;
	output \g62709/_0_  ;
	output \g62710/_0_  ;
	output \g62711/_0_  ;
	output \g62714/_0_  ;
	output \g62715/_0_  ;
	output \g62717/_0_  ;
	output \g62718/_0_  ;
	output \g62719/_0_  ;
	output \g62720/_0_  ;
	output \g62721/_0_  ;
	output \g62723/_0_  ;
	output \g62725/_0_  ;
	output \g62726/_0_  ;
	output \g62729/_0_  ;
	output \g62731/_0_  ;
	output \g62733/_0_  ;
	output \g62738/_0_  ;
	output \g62741/_0_  ;
	output \g62742/_0_  ;
	output \g62744/_0_  ;
	output \g62745/_0_  ;
	output \g62746/_0_  ;
	output \g62747/_0_  ;
	output \g62748/_0_  ;
	output \g62749/_0_  ;
	output \g62753/_0_  ;
	output \g62755/_0_  ;
	output \g62756/_0_  ;
	output \g62758/_0_  ;
	output \g62759/_0_  ;
	output \g62760/_0_  ;
	output \g62761/_0_  ;
	output \g62763/_0_  ;
	output \g62766/_0_  ;
	output \g62767/_0_  ;
	output \g62768/_0_  ;
	output \g65554/_0_  ;
	output \g65561/_0_  ;
	output \g65569/_0_  ;
	output \g65580/_0_  ;
	output \g65599/_0_  ;
	output \g65606/_0_  ;
	output \g65636/_0_  ;
	output \g65864/_0_  ;
	wire _w4373_ ;
	wire _w4372_ ;
	wire _w4371_ ;
	wire _w4370_ ;
	wire _w4369_ ;
	wire _w4368_ ;
	wire _w4367_ ;
	wire _w4366_ ;
	wire _w4365_ ;
	wire _w4364_ ;
	wire _w4363_ ;
	wire _w4362_ ;
	wire _w4361_ ;
	wire _w4360_ ;
	wire _w4359_ ;
	wire _w4358_ ;
	wire _w4357_ ;
	wire _w4356_ ;
	wire _w4355_ ;
	wire _w4354_ ;
	wire _w4353_ ;
	wire _w4352_ ;
	wire _w4351_ ;
	wire _w4350_ ;
	wire _w4349_ ;
	wire _w4348_ ;
	wire _w4347_ ;
	wire _w4346_ ;
	wire _w4345_ ;
	wire _w4344_ ;
	wire _w4343_ ;
	wire _w4342_ ;
	wire _w4341_ ;
	wire _w4340_ ;
	wire _w4339_ ;
	wire _w4338_ ;
	wire _w4337_ ;
	wire _w4336_ ;
	wire _w4335_ ;
	wire _w4334_ ;
	wire _w4333_ ;
	wire _w4332_ ;
	wire _w4331_ ;
	wire _w4330_ ;
	wire _w4329_ ;
	wire _w4328_ ;
	wire _w4327_ ;
	wire _w4326_ ;
	wire _w4325_ ;
	wire _w4324_ ;
	wire _w4323_ ;
	wire _w4322_ ;
	wire _w4321_ ;
	wire _w4320_ ;
	wire _w4319_ ;
	wire _w4318_ ;
	wire _w4317_ ;
	wire _w4316_ ;
	wire _w4315_ ;
	wire _w4314_ ;
	wire _w4313_ ;
	wire _w4312_ ;
	wire _w4311_ ;
	wire _w4310_ ;
	wire _w4309_ ;
	wire _w4308_ ;
	wire _w4307_ ;
	wire _w4306_ ;
	wire _w4305_ ;
	wire _w4304_ ;
	wire _w4303_ ;
	wire _w4302_ ;
	wire _w4301_ ;
	wire _w4300_ ;
	wire _w4299_ ;
	wire _w4298_ ;
	wire _w4297_ ;
	wire _w4296_ ;
	wire _w4295_ ;
	wire _w4294_ ;
	wire _w4293_ ;
	wire _w4292_ ;
	wire _w4291_ ;
	wire _w4290_ ;
	wire _w4289_ ;
	wire _w4288_ ;
	wire _w4287_ ;
	wire _w4286_ ;
	wire _w4285_ ;
	wire _w4284_ ;
	wire _w4283_ ;
	wire _w4282_ ;
	wire _w4281_ ;
	wire _w4280_ ;
	wire _w4279_ ;
	wire _w4278_ ;
	wire _w4277_ ;
	wire _w4276_ ;
	wire _w4275_ ;
	wire _w4274_ ;
	wire _w4273_ ;
	wire _w4272_ ;
	wire _w4271_ ;
	wire _w4270_ ;
	wire _w4269_ ;
	wire _w4268_ ;
	wire _w4267_ ;
	wire _w4266_ ;
	wire _w4265_ ;
	wire _w4264_ ;
	wire _w4263_ ;
	wire _w4262_ ;
	wire _w4261_ ;
	wire _w4260_ ;
	wire _w4259_ ;
	wire _w4258_ ;
	wire _w4257_ ;
	wire _w4256_ ;
	wire _w4255_ ;
	wire _w4254_ ;
	wire _w4253_ ;
	wire _w4252_ ;
	wire _w4251_ ;
	wire _w4250_ ;
	wire _w4249_ ;
	wire _w4248_ ;
	wire _w4247_ ;
	wire _w4246_ ;
	wire _w4245_ ;
	wire _w4244_ ;
	wire _w4243_ ;
	wire _w4242_ ;
	wire _w4241_ ;
	wire _w4240_ ;
	wire _w4239_ ;
	wire _w4238_ ;
	wire _w4237_ ;
	wire _w4236_ ;
	wire _w4235_ ;
	wire _w4234_ ;
	wire _w4233_ ;
	wire _w4232_ ;
	wire _w4231_ ;
	wire _w4230_ ;
	wire _w4229_ ;
	wire _w4228_ ;
	wire _w4227_ ;
	wire _w4226_ ;
	wire _w4225_ ;
	wire _w4224_ ;
	wire _w4223_ ;
	wire _w4222_ ;
	wire _w4221_ ;
	wire _w4220_ ;
	wire _w4219_ ;
	wire _w4218_ ;
	wire _w4217_ ;
	wire _w4216_ ;
	wire _w4215_ ;
	wire _w4214_ ;
	wire _w4213_ ;
	wire _w4212_ ;
	wire _w4211_ ;
	wire _w4210_ ;
	wire _w4209_ ;
	wire _w4208_ ;
	wire _w4207_ ;
	wire _w4206_ ;
	wire _w4205_ ;
	wire _w4204_ ;
	wire _w4203_ ;
	wire _w4202_ ;
	wire _w4201_ ;
	wire _w4200_ ;
	wire _w4199_ ;
	wire _w4198_ ;
	wire _w4197_ ;
	wire _w4196_ ;
	wire _w4195_ ;
	wire _w4194_ ;
	wire _w4193_ ;
	wire _w4192_ ;
	wire _w4191_ ;
	wire _w4190_ ;
	wire _w4189_ ;
	wire _w4188_ ;
	wire _w4187_ ;
	wire _w4186_ ;
	wire _w4185_ ;
	wire _w4184_ ;
	wire _w4183_ ;
	wire _w4182_ ;
	wire _w4181_ ;
	wire _w4180_ ;
	wire _w4179_ ;
	wire _w4178_ ;
	wire _w4177_ ;
	wire _w4176_ ;
	wire _w4175_ ;
	wire _w4174_ ;
	wire _w4173_ ;
	wire _w4172_ ;
	wire _w4171_ ;
	wire _w4170_ ;
	wire _w4169_ ;
	wire _w4168_ ;
	wire _w4167_ ;
	wire _w4166_ ;
	wire _w4165_ ;
	wire _w4164_ ;
	wire _w4163_ ;
	wire _w4162_ ;
	wire _w4161_ ;
	wire _w4160_ ;
	wire _w4159_ ;
	wire _w4158_ ;
	wire _w4157_ ;
	wire _w4156_ ;
	wire _w4155_ ;
	wire _w4154_ ;
	wire _w4153_ ;
	wire _w4152_ ;
	wire _w4151_ ;
	wire _w4150_ ;
	wire _w4149_ ;
	wire _w4148_ ;
	wire _w4147_ ;
	wire _w4146_ ;
	wire _w4145_ ;
	wire _w4144_ ;
	wire _w4143_ ;
	wire _w4142_ ;
	wire _w4141_ ;
	wire _w4140_ ;
	wire _w4139_ ;
	wire _w4138_ ;
	wire _w4137_ ;
	wire _w4136_ ;
	wire _w4135_ ;
	wire _w4134_ ;
	wire _w4133_ ;
	wire _w4132_ ;
	wire _w4131_ ;
	wire _w4130_ ;
	wire _w4129_ ;
	wire _w4128_ ;
	wire _w4127_ ;
	wire _w4126_ ;
	wire _w4125_ ;
	wire _w4124_ ;
	wire _w4123_ ;
	wire _w4122_ ;
	wire _w4121_ ;
	wire _w4120_ ;
	wire _w4119_ ;
	wire _w4118_ ;
	wire _w4117_ ;
	wire _w4116_ ;
	wire _w4115_ ;
	wire _w4114_ ;
	wire _w4113_ ;
	wire _w4112_ ;
	wire _w4111_ ;
	wire _w4110_ ;
	wire _w4109_ ;
	wire _w4108_ ;
	wire _w4107_ ;
	wire _w4106_ ;
	wire _w4105_ ;
	wire _w4104_ ;
	wire _w4103_ ;
	wire _w4102_ ;
	wire _w4101_ ;
	wire _w4100_ ;
	wire _w4099_ ;
	wire _w4098_ ;
	wire _w4097_ ;
	wire _w4096_ ;
	wire _w4095_ ;
	wire _w4094_ ;
	wire _w4093_ ;
	wire _w4092_ ;
	wire _w4091_ ;
	wire _w4090_ ;
	wire _w4089_ ;
	wire _w4088_ ;
	wire _w4087_ ;
	wire _w4086_ ;
	wire _w4085_ ;
	wire _w4084_ ;
	wire _w4083_ ;
	wire _w4082_ ;
	wire _w4081_ ;
	wire _w4080_ ;
	wire _w4079_ ;
	wire _w4078_ ;
	wire _w4077_ ;
	wire _w4076_ ;
	wire _w4075_ ;
	wire _w4074_ ;
	wire _w4073_ ;
	wire _w4072_ ;
	wire _w4071_ ;
	wire _w4070_ ;
	wire _w4069_ ;
	wire _w4068_ ;
	wire _w4067_ ;
	wire _w4066_ ;
	wire _w4065_ ;
	wire _w4064_ ;
	wire _w4063_ ;
	wire _w4062_ ;
	wire _w4061_ ;
	wire _w4060_ ;
	wire _w4059_ ;
	wire _w4058_ ;
	wire _w4057_ ;
	wire _w4056_ ;
	wire _w4055_ ;
	wire _w4054_ ;
	wire _w4053_ ;
	wire _w4052_ ;
	wire _w4051_ ;
	wire _w4050_ ;
	wire _w4049_ ;
	wire _w4048_ ;
	wire _w4047_ ;
	wire _w4046_ ;
	wire _w4045_ ;
	wire _w4044_ ;
	wire _w4043_ ;
	wire _w4042_ ;
	wire _w4041_ ;
	wire _w4040_ ;
	wire _w4039_ ;
	wire _w4038_ ;
	wire _w4037_ ;
	wire _w4036_ ;
	wire _w4035_ ;
	wire _w4034_ ;
	wire _w4033_ ;
	wire _w4032_ ;
	wire _w4031_ ;
	wire _w4030_ ;
	wire _w4029_ ;
	wire _w4028_ ;
	wire _w4027_ ;
	wire _w4026_ ;
	wire _w4025_ ;
	wire _w4024_ ;
	wire _w4023_ ;
	wire _w4022_ ;
	wire _w4021_ ;
	wire _w4020_ ;
	wire _w4019_ ;
	wire _w4018_ ;
	wire _w4017_ ;
	wire _w4016_ ;
	wire _w4015_ ;
	wire _w4014_ ;
	wire _w4013_ ;
	wire _w4012_ ;
	wire _w4011_ ;
	wire _w4010_ ;
	wire _w4009_ ;
	wire _w4008_ ;
	wire _w4007_ ;
	wire _w4006_ ;
	wire _w4005_ ;
	wire _w4004_ ;
	wire _w4003_ ;
	wire _w4002_ ;
	wire _w4001_ ;
	wire _w4000_ ;
	wire _w3999_ ;
	wire _w3998_ ;
	wire _w3997_ ;
	wire _w3996_ ;
	wire _w3995_ ;
	wire _w3994_ ;
	wire _w3993_ ;
	wire _w3992_ ;
	wire _w3991_ ;
	wire _w3990_ ;
	wire _w3989_ ;
	wire _w3988_ ;
	wire _w3987_ ;
	wire _w3986_ ;
	wire _w3985_ ;
	wire _w3984_ ;
	wire _w3983_ ;
	wire _w3982_ ;
	wire _w3981_ ;
	wire _w3980_ ;
	wire _w3979_ ;
	wire _w3978_ ;
	wire _w3977_ ;
	wire _w3976_ ;
	wire _w3975_ ;
	wire _w3974_ ;
	wire _w3973_ ;
	wire _w3972_ ;
	wire _w3971_ ;
	wire _w3970_ ;
	wire _w3969_ ;
	wire _w3968_ ;
	wire _w3967_ ;
	wire _w3966_ ;
	wire _w3965_ ;
	wire _w3964_ ;
	wire _w3963_ ;
	wire _w3962_ ;
	wire _w3961_ ;
	wire _w3960_ ;
	wire _w3959_ ;
	wire _w3958_ ;
	wire _w3957_ ;
	wire _w3956_ ;
	wire _w3955_ ;
	wire _w3954_ ;
	wire _w3953_ ;
	wire _w3952_ ;
	wire _w3951_ ;
	wire _w3950_ ;
	wire _w3949_ ;
	wire _w3948_ ;
	wire _w3947_ ;
	wire _w3946_ ;
	wire _w3945_ ;
	wire _w3944_ ;
	wire _w3943_ ;
	wire _w3942_ ;
	wire _w3941_ ;
	wire _w3940_ ;
	wire _w3939_ ;
	wire _w3938_ ;
	wire _w3937_ ;
	wire _w3936_ ;
	wire _w3935_ ;
	wire _w3934_ ;
	wire _w3933_ ;
	wire _w3932_ ;
	wire _w3931_ ;
	wire _w3930_ ;
	wire _w3929_ ;
	wire _w3928_ ;
	wire _w3927_ ;
	wire _w3926_ ;
	wire _w3925_ ;
	wire _w3924_ ;
	wire _w3923_ ;
	wire _w3922_ ;
	wire _w3921_ ;
	wire _w3920_ ;
	wire _w3919_ ;
	wire _w3918_ ;
	wire _w3917_ ;
	wire _w3916_ ;
	wire _w3915_ ;
	wire _w3914_ ;
	wire _w3913_ ;
	wire _w3912_ ;
	wire _w3911_ ;
	wire _w3910_ ;
	wire _w3909_ ;
	wire _w3908_ ;
	wire _w3907_ ;
	wire _w3906_ ;
	wire _w3905_ ;
	wire _w3904_ ;
	wire _w3903_ ;
	wire _w3902_ ;
	wire _w3901_ ;
	wire _w3900_ ;
	wire _w3899_ ;
	wire _w3898_ ;
	wire _w3897_ ;
	wire _w3896_ ;
	wire _w3895_ ;
	wire _w3894_ ;
	wire _w3893_ ;
	wire _w3892_ ;
	wire _w3891_ ;
	wire _w3890_ ;
	wire _w3889_ ;
	wire _w3888_ ;
	wire _w3887_ ;
	wire _w3886_ ;
	wire _w3885_ ;
	wire _w3884_ ;
	wire _w3883_ ;
	wire _w3882_ ;
	wire _w3881_ ;
	wire _w3880_ ;
	wire _w3879_ ;
	wire _w3878_ ;
	wire _w3877_ ;
	wire _w3876_ ;
	wire _w3875_ ;
	wire _w3874_ ;
	wire _w3873_ ;
	wire _w3872_ ;
	wire _w3871_ ;
	wire _w3870_ ;
	wire _w3869_ ;
	wire _w3868_ ;
	wire _w3867_ ;
	wire _w3866_ ;
	wire _w2617_ ;
	wire _w2616_ ;
	wire _w2615_ ;
	wire _w2614_ ;
	wire _w2613_ ;
	wire _w2612_ ;
	wire _w2611_ ;
	wire _w2610_ ;
	wire _w2609_ ;
	wire _w2608_ ;
	wire _w2607_ ;
	wire _w2606_ ;
	wire _w2605_ ;
	wire _w2604_ ;
	wire _w2603_ ;
	wire _w2602_ ;
	wire _w2601_ ;
	wire _w2600_ ;
	wire _w2599_ ;
	wire _w2598_ ;
	wire _w2597_ ;
	wire _w2596_ ;
	wire _w2595_ ;
	wire _w2594_ ;
	wire _w2593_ ;
	wire _w2592_ ;
	wire _w2591_ ;
	wire _w2590_ ;
	wire _w2589_ ;
	wire _w2588_ ;
	wire _w2587_ ;
	wire _w2586_ ;
	wire _w2585_ ;
	wire _w2584_ ;
	wire _w2583_ ;
	wire _w2582_ ;
	wire _w2581_ ;
	wire _w2580_ ;
	wire _w2579_ ;
	wire _w2578_ ;
	wire _w2577_ ;
	wire _w2576_ ;
	wire _w2575_ ;
	wire _w2574_ ;
	wire _w2573_ ;
	wire _w2572_ ;
	wire _w2571_ ;
	wire _w2570_ ;
	wire _w2569_ ;
	wire _w2568_ ;
	wire _w2567_ ;
	wire _w2566_ ;
	wire _w2565_ ;
	wire _w2564_ ;
	wire _w2563_ ;
	wire _w2562_ ;
	wire _w2561_ ;
	wire _w2560_ ;
	wire _w2559_ ;
	wire _w2558_ ;
	wire _w2557_ ;
	wire _w2556_ ;
	wire _w2555_ ;
	wire _w2554_ ;
	wire _w2553_ ;
	wire _w2552_ ;
	wire _w2551_ ;
	wire _w2550_ ;
	wire _w2549_ ;
	wire _w2548_ ;
	wire _w2547_ ;
	wire _w2546_ ;
	wire _w2545_ ;
	wire _w2544_ ;
	wire _w2543_ ;
	wire _w2542_ ;
	wire _w2541_ ;
	wire _w2540_ ;
	wire _w2539_ ;
	wire _w2538_ ;
	wire _w2537_ ;
	wire _w2536_ ;
	wire _w2535_ ;
	wire _w2534_ ;
	wire _w2533_ ;
	wire _w2532_ ;
	wire _w2531_ ;
	wire _w2530_ ;
	wire _w2529_ ;
	wire _w2528_ ;
	wire _w2527_ ;
	wire _w2526_ ;
	wire _w2525_ ;
	wire _w2524_ ;
	wire _w2523_ ;
	wire _w2522_ ;
	wire _w2521_ ;
	wire _w2520_ ;
	wire _w2519_ ;
	wire _w2518_ ;
	wire _w2517_ ;
	wire _w2516_ ;
	wire _w2515_ ;
	wire _w2514_ ;
	wire _w2513_ ;
	wire _w2512_ ;
	wire _w2511_ ;
	wire _w2510_ ;
	wire _w2509_ ;
	wire _w2508_ ;
	wire _w2507_ ;
	wire _w2506_ ;
	wire _w2505_ ;
	wire _w2504_ ;
	wire _w2503_ ;
	wire _w2502_ ;
	wire _w2501_ ;
	wire _w2500_ ;
	wire _w2499_ ;
	wire _w2498_ ;
	wire _w2497_ ;
	wire _w2496_ ;
	wire _w2495_ ;
	wire _w2494_ ;
	wire _w2493_ ;
	wire _w2492_ ;
	wire _w2491_ ;
	wire _w2490_ ;
	wire _w2489_ ;
	wire _w2488_ ;
	wire _w2487_ ;
	wire _w2486_ ;
	wire _w2485_ ;
	wire _w2484_ ;
	wire _w2483_ ;
	wire _w2482_ ;
	wire _w2481_ ;
	wire _w2480_ ;
	wire _w2479_ ;
	wire _w2478_ ;
	wire _w2477_ ;
	wire _w2476_ ;
	wire _w2475_ ;
	wire _w2474_ ;
	wire _w2473_ ;
	wire _w2472_ ;
	wire _w2471_ ;
	wire _w2470_ ;
	wire _w2469_ ;
	wire _w2468_ ;
	wire _w2467_ ;
	wire _w2466_ ;
	wire _w2465_ ;
	wire _w2464_ ;
	wire _w2463_ ;
	wire _w2462_ ;
	wire _w2461_ ;
	wire _w2460_ ;
	wire _w2459_ ;
	wire _w2458_ ;
	wire _w2457_ ;
	wire _w2456_ ;
	wire _w2455_ ;
	wire _w2454_ ;
	wire _w2453_ ;
	wire _w2452_ ;
	wire _w2451_ ;
	wire _w2450_ ;
	wire _w2449_ ;
	wire _w2448_ ;
	wire _w2447_ ;
	wire _w2446_ ;
	wire _w2445_ ;
	wire _w2444_ ;
	wire _w2443_ ;
	wire _w2442_ ;
	wire _w2441_ ;
	wire _w2440_ ;
	wire _w2439_ ;
	wire _w2438_ ;
	wire _w2437_ ;
	wire _w2436_ ;
	wire _w2435_ ;
	wire _w2434_ ;
	wire _w2433_ ;
	wire _w2432_ ;
	wire _w2431_ ;
	wire _w2430_ ;
	wire _w2429_ ;
	wire _w2428_ ;
	wire _w2427_ ;
	wire _w2426_ ;
	wire _w2425_ ;
	wire _w2424_ ;
	wire _w2423_ ;
	wire _w2422_ ;
	wire _w2421_ ;
	wire _w2420_ ;
	wire _w2419_ ;
	wire _w2418_ ;
	wire _w2417_ ;
	wire _w2416_ ;
	wire _w2415_ ;
	wire _w2414_ ;
	wire _w2413_ ;
	wire _w2412_ ;
	wire _w2411_ ;
	wire _w2410_ ;
	wire _w2409_ ;
	wire _w2408_ ;
	wire _w2407_ ;
	wire _w2406_ ;
	wire _w2405_ ;
	wire _w2404_ ;
	wire _w2403_ ;
	wire _w2402_ ;
	wire _w2401_ ;
	wire _w2400_ ;
	wire _w2399_ ;
	wire _w2398_ ;
	wire _w2397_ ;
	wire _w2396_ ;
	wire _w2395_ ;
	wire _w2394_ ;
	wire _w2393_ ;
	wire _w2392_ ;
	wire _w2391_ ;
	wire _w2390_ ;
	wire _w2389_ ;
	wire _w2388_ ;
	wire _w2387_ ;
	wire _w2386_ ;
	wire _w2385_ ;
	wire _w2384_ ;
	wire _w2383_ ;
	wire _w2382_ ;
	wire _w2381_ ;
	wire _w2380_ ;
	wire _w2379_ ;
	wire _w2378_ ;
	wire _w2377_ ;
	wire _w2376_ ;
	wire _w2375_ ;
	wire _w2374_ ;
	wire _w2373_ ;
	wire _w2372_ ;
	wire _w2371_ ;
	wire _w2370_ ;
	wire _w2369_ ;
	wire _w2368_ ;
	wire _w2367_ ;
	wire _w2366_ ;
	wire _w2365_ ;
	wire _w2364_ ;
	wire _w2363_ ;
	wire _w2362_ ;
	wire _w2361_ ;
	wire _w2360_ ;
	wire _w2359_ ;
	wire _w2358_ ;
	wire _w2357_ ;
	wire _w2356_ ;
	wire _w2355_ ;
	wire _w2354_ ;
	wire _w2353_ ;
	wire _w2352_ ;
	wire _w2351_ ;
	wire _w2350_ ;
	wire _w2349_ ;
	wire _w2348_ ;
	wire _w2347_ ;
	wire _w2346_ ;
	wire _w2345_ ;
	wire _w2344_ ;
	wire _w2343_ ;
	wire _w2342_ ;
	wire _w2341_ ;
	wire _w2340_ ;
	wire _w2339_ ;
	wire _w2338_ ;
	wire _w2337_ ;
	wire _w2336_ ;
	wire _w2335_ ;
	wire _w2334_ ;
	wire _w2333_ ;
	wire _w2332_ ;
	wire _w2331_ ;
	wire _w2330_ ;
	wire _w2329_ ;
	wire _w2328_ ;
	wire _w2327_ ;
	wire _w2326_ ;
	wire _w2325_ ;
	wire _w2324_ ;
	wire _w2323_ ;
	wire _w2322_ ;
	wire _w2321_ ;
	wire _w2320_ ;
	wire _w2319_ ;
	wire _w2318_ ;
	wire _w2317_ ;
	wire _w2316_ ;
	wire _w2315_ ;
	wire _w2314_ ;
	wire _w2313_ ;
	wire _w2312_ ;
	wire _w2311_ ;
	wire _w2310_ ;
	wire _w2309_ ;
	wire _w2308_ ;
	wire _w2307_ ;
	wire _w2306_ ;
	wire _w2305_ ;
	wire _w2304_ ;
	wire _w2303_ ;
	wire _w2302_ ;
	wire _w2301_ ;
	wire _w2300_ ;
	wire _w2299_ ;
	wire _w2298_ ;
	wire _w2297_ ;
	wire _w2296_ ;
	wire _w2295_ ;
	wire _w2294_ ;
	wire _w2293_ ;
	wire _w2292_ ;
	wire _w2291_ ;
	wire _w2290_ ;
	wire _w2289_ ;
	wire _w2288_ ;
	wire _w2287_ ;
	wire _w2286_ ;
	wire _w2285_ ;
	wire _w2284_ ;
	wire _w2283_ ;
	wire _w2282_ ;
	wire _w2281_ ;
	wire _w2280_ ;
	wire _w2279_ ;
	wire _w2278_ ;
	wire _w2277_ ;
	wire _w2276_ ;
	wire _w2275_ ;
	wire _w2274_ ;
	wire _w2273_ ;
	wire _w2272_ ;
	wire _w2271_ ;
	wire _w2270_ ;
	wire _w2269_ ;
	wire _w2268_ ;
	wire _w2267_ ;
	wire _w2266_ ;
	wire _w2265_ ;
	wire _w2264_ ;
	wire _w2263_ ;
	wire _w2262_ ;
	wire _w2261_ ;
	wire _w2260_ ;
	wire _w2259_ ;
	wire _w2258_ ;
	wire _w2257_ ;
	wire _w2256_ ;
	wire _w2255_ ;
	wire _w2254_ ;
	wire _w2253_ ;
	wire _w2252_ ;
	wire _w2251_ ;
	wire _w2250_ ;
	wire _w2249_ ;
	wire _w2248_ ;
	wire _w2247_ ;
	wire _w2246_ ;
	wire _w2245_ ;
	wire _w2244_ ;
	wire _w2243_ ;
	wire _w2242_ ;
	wire _w2241_ ;
	wire _w2240_ ;
	wire _w2239_ ;
	wire _w2238_ ;
	wire _w2237_ ;
	wire _w2236_ ;
	wire _w2235_ ;
	wire _w2234_ ;
	wire _w2233_ ;
	wire _w2232_ ;
	wire _w2231_ ;
	wire _w2230_ ;
	wire _w2229_ ;
	wire _w2228_ ;
	wire _w2227_ ;
	wire _w2226_ ;
	wire _w2225_ ;
	wire _w2224_ ;
	wire _w2223_ ;
	wire _w2222_ ;
	wire _w2221_ ;
	wire _w2220_ ;
	wire _w2219_ ;
	wire _w2218_ ;
	wire _w2217_ ;
	wire _w2216_ ;
	wire _w2215_ ;
	wire _w2214_ ;
	wire _w2213_ ;
	wire _w2212_ ;
	wire _w2211_ ;
	wire _w2210_ ;
	wire _w2209_ ;
	wire _w2208_ ;
	wire _w2207_ ;
	wire _w2206_ ;
	wire _w2205_ ;
	wire _w2204_ ;
	wire _w2203_ ;
	wire _w2202_ ;
	wire _w2201_ ;
	wire _w2200_ ;
	wire _w2199_ ;
	wire _w2198_ ;
	wire _w2197_ ;
	wire _w2196_ ;
	wire _w2195_ ;
	wire _w2194_ ;
	wire _w2193_ ;
	wire _w2192_ ;
	wire _w2191_ ;
	wire _w2190_ ;
	wire _w2189_ ;
	wire _w2188_ ;
	wire _w2187_ ;
	wire _w2186_ ;
	wire _w2185_ ;
	wire _w2184_ ;
	wire _w2183_ ;
	wire _w2182_ ;
	wire _w2181_ ;
	wire _w2180_ ;
	wire _w2179_ ;
	wire _w2178_ ;
	wire _w2177_ ;
	wire _w2176_ ;
	wire _w2175_ ;
	wire _w2174_ ;
	wire _w2173_ ;
	wire _w2172_ ;
	wire _w2171_ ;
	wire _w2170_ ;
	wire _w2169_ ;
	wire _w2168_ ;
	wire _w2167_ ;
	wire _w2166_ ;
	wire _w2165_ ;
	wire _w2164_ ;
	wire _w2163_ ;
	wire _w2162_ ;
	wire _w2161_ ;
	wire _w2160_ ;
	wire _w2159_ ;
	wire _w2158_ ;
	wire _w2157_ ;
	wire _w2156_ ;
	wire _w2155_ ;
	wire _w2154_ ;
	wire _w2153_ ;
	wire _w2152_ ;
	wire _w2151_ ;
	wire _w2150_ ;
	wire _w2149_ ;
	wire _w2148_ ;
	wire _w2147_ ;
	wire _w2146_ ;
	wire _w2145_ ;
	wire _w2144_ ;
	wire _w2143_ ;
	wire _w2142_ ;
	wire _w2141_ ;
	wire _w2140_ ;
	wire _w2139_ ;
	wire _w2138_ ;
	wire _w2137_ ;
	wire _w2136_ ;
	wire _w2135_ ;
	wire _w2134_ ;
	wire _w2133_ ;
	wire _w2132_ ;
	wire _w2131_ ;
	wire _w2130_ ;
	wire _w2129_ ;
	wire _w2128_ ;
	wire _w2127_ ;
	wire _w2126_ ;
	wire _w2125_ ;
	wire _w2124_ ;
	wire _w2123_ ;
	wire _w2122_ ;
	wire _w2121_ ;
	wire _w2120_ ;
	wire _w2119_ ;
	wire _w2118_ ;
	wire _w2117_ ;
	wire _w2116_ ;
	wire _w2115_ ;
	wire _w2114_ ;
	wire _w2113_ ;
	wire _w2112_ ;
	wire _w2111_ ;
	wire _w2110_ ;
	wire _w2109_ ;
	wire _w2108_ ;
	wire _w2107_ ;
	wire _w2106_ ;
	wire _w2105_ ;
	wire _w2104_ ;
	wire _w2103_ ;
	wire _w2102_ ;
	wire _w2101_ ;
	wire _w2100_ ;
	wire _w2099_ ;
	wire _w2098_ ;
	wire _w2097_ ;
	wire _w2096_ ;
	wire _w2095_ ;
	wire _w2094_ ;
	wire _w2093_ ;
	wire _w2092_ ;
	wire _w2091_ ;
	wire _w2090_ ;
	wire _w2089_ ;
	wire _w2088_ ;
	wire _w2087_ ;
	wire _w2086_ ;
	wire _w2085_ ;
	wire _w2084_ ;
	wire _w2083_ ;
	wire _w2082_ ;
	wire _w2081_ ;
	wire _w2080_ ;
	wire _w2079_ ;
	wire _w2078_ ;
	wire _w2077_ ;
	wire _w2076_ ;
	wire _w2075_ ;
	wire _w2074_ ;
	wire _w2073_ ;
	wire _w2072_ ;
	wire _w2071_ ;
	wire _w2070_ ;
	wire _w2069_ ;
	wire _w2068_ ;
	wire _w2067_ ;
	wire _w2066_ ;
	wire _w2065_ ;
	wire _w2064_ ;
	wire _w2063_ ;
	wire _w2062_ ;
	wire _w2061_ ;
	wire _w2060_ ;
	wire _w2059_ ;
	wire _w2058_ ;
	wire _w2057_ ;
	wire _w2056_ ;
	wire _w2055_ ;
	wire _w2054_ ;
	wire _w2053_ ;
	wire _w2052_ ;
	wire _w2051_ ;
	wire _w2050_ ;
	wire _w1765_ ;
	wire _w1764_ ;
	wire _w1763_ ;
	wire _w1762_ ;
	wire _w1761_ ;
	wire _w1760_ ;
	wire _w1759_ ;
	wire _w1758_ ;
	wire _w1757_ ;
	wire _w1756_ ;
	wire _w1755_ ;
	wire _w1754_ ;
	wire _w1753_ ;
	wire _w1752_ ;
	wire _w1751_ ;
	wire _w1750_ ;
	wire _w1749_ ;
	wire _w1748_ ;
	wire _w1747_ ;
	wire _w1746_ ;
	wire _w1745_ ;
	wire _w1744_ ;
	wire _w1743_ ;
	wire _w1742_ ;
	wire _w1741_ ;
	wire _w1740_ ;
	wire _w1739_ ;
	wire _w1738_ ;
	wire _w1737_ ;
	wire _w1736_ ;
	wire _w1735_ ;
	wire _w1734_ ;
	wire _w1733_ ;
	wire _w1732_ ;
	wire _w1731_ ;
	wire _w1730_ ;
	wire _w1729_ ;
	wire _w1728_ ;
	wire _w1727_ ;
	wire _w1726_ ;
	wire _w1725_ ;
	wire _w1724_ ;
	wire _w1723_ ;
	wire _w1722_ ;
	wire _w1721_ ;
	wire _w1720_ ;
	wire _w1719_ ;
	wire _w1718_ ;
	wire _w1717_ ;
	wire _w1716_ ;
	wire _w1715_ ;
	wire _w1714_ ;
	wire _w1713_ ;
	wire _w1712_ ;
	wire _w1711_ ;
	wire _w1710_ ;
	wire _w1709_ ;
	wire _w1708_ ;
	wire _w1707_ ;
	wire _w1706_ ;
	wire _w1705_ ;
	wire _w1704_ ;
	wire _w1703_ ;
	wire _w1702_ ;
	wire _w1701_ ;
	wire _w1700_ ;
	wire _w1699_ ;
	wire _w1698_ ;
	wire _w1697_ ;
	wire _w1696_ ;
	wire _w1695_ ;
	wire _w1694_ ;
	wire _w1693_ ;
	wire _w1692_ ;
	wire _w1691_ ;
	wire _w1690_ ;
	wire _w1689_ ;
	wire _w1688_ ;
	wire _w1687_ ;
	wire _w1686_ ;
	wire _w1685_ ;
	wire _w1684_ ;
	wire _w1683_ ;
	wire _w1682_ ;
	wire _w1681_ ;
	wire _w1680_ ;
	wire _w1679_ ;
	wire _w1678_ ;
	wire _w1677_ ;
	wire _w1676_ ;
	wire _w1675_ ;
	wire _w1674_ ;
	wire _w1673_ ;
	wire _w1672_ ;
	wire _w1671_ ;
	wire _w1670_ ;
	wire _w1669_ ;
	wire _w1668_ ;
	wire _w1667_ ;
	wire _w1666_ ;
	wire _w1665_ ;
	wire _w1664_ ;
	wire _w1663_ ;
	wire _w1662_ ;
	wire _w1661_ ;
	wire _w1660_ ;
	wire _w1659_ ;
	wire _w1658_ ;
	wire _w1657_ ;
	wire _w1656_ ;
	wire _w1655_ ;
	wire _w1654_ ;
	wire _w1653_ ;
	wire _w1652_ ;
	wire _w1651_ ;
	wire _w1650_ ;
	wire _w1649_ ;
	wire _w1648_ ;
	wire _w1647_ ;
	wire _w1646_ ;
	wire _w1645_ ;
	wire _w1644_ ;
	wire _w1643_ ;
	wire _w1642_ ;
	wire _w1641_ ;
	wire _w1640_ ;
	wire _w1639_ ;
	wire _w1638_ ;
	wire _w1637_ ;
	wire _w1636_ ;
	wire _w1567_ ;
	wire _w1566_ ;
	wire _w1565_ ;
	wire _w1564_ ;
	wire _w1563_ ;
	wire _w1562_ ;
	wire _w1561_ ;
	wire _w1560_ ;
	wire _w1559_ ;
	wire _w1558_ ;
	wire _w1557_ ;
	wire _w1556_ ;
	wire _w1555_ ;
	wire _w1554_ ;
	wire _w1553_ ;
	wire _w1552_ ;
	wire _w1551_ ;
	wire _w1550_ ;
	wire _w1549_ ;
	wire _w1548_ ;
	wire _w1547_ ;
	wire _w1546_ ;
	wire _w1545_ ;
	wire _w1544_ ;
	wire _w1543_ ;
	wire _w1542_ ;
	wire _w1541_ ;
	wire _w1540_ ;
	wire _w1539_ ;
	wire _w1538_ ;
	wire _w1521_ ;
	wire _w1520_ ;
	wire _w1519_ ;
	wire _w1518_ ;
	wire _w1517_ ;
	wire _w1516_ ;
	wire _w1515_ ;
	wire _w1514_ ;
	wire _w1513_ ;
	wire _w1512_ ;
	wire _w1511_ ;
	wire _w1510_ ;
	wire _w1509_ ;
	wire _w1522_ ;
	wire _w1523_ ;
	wire _w1524_ ;
	wire _w1525_ ;
	wire _w1526_ ;
	wire _w1527_ ;
	wire _w1528_ ;
	wire _w1529_ ;
	wire _w1530_ ;
	wire _w1531_ ;
	wire _w1532_ ;
	wire _w1533_ ;
	wire _w1534_ ;
	wire _w1535_ ;
	wire _w1536_ ;
	wire _w1537_ ;
	wire _w1568_ ;
	wire _w1569_ ;
	wire _w1570_ ;
	wire _w1571_ ;
	wire _w1572_ ;
	wire _w1573_ ;
	wire _w1574_ ;
	wire _w1575_ ;
	wire _w1576_ ;
	wire _w1577_ ;
	wire _w1578_ ;
	wire _w1579_ ;
	wire _w1580_ ;
	wire _w1581_ ;
	wire _w1582_ ;
	wire _w1583_ ;
	wire _w1584_ ;
	wire _w1585_ ;
	wire _w1586_ ;
	wire _w1587_ ;
	wire _w1588_ ;
	wire _w1589_ ;
	wire _w1590_ ;
	wire _w1591_ ;
	wire _w1592_ ;
	wire _w1593_ ;
	wire _w1594_ ;
	wire _w1595_ ;
	wire _w1596_ ;
	wire _w1597_ ;
	wire _w1598_ ;
	wire _w1599_ ;
	wire _w1600_ ;
	wire _w1601_ ;
	wire _w1602_ ;
	wire _w1603_ ;
	wire _w1604_ ;
	wire _w1605_ ;
	wire _w1606_ ;
	wire _w1607_ ;
	wire _w1608_ ;
	wire _w1609_ ;
	wire _w1610_ ;
	wire _w1611_ ;
	wire _w1612_ ;
	wire _w1613_ ;
	wire _w1614_ ;
	wire _w1615_ ;
	wire _w1616_ ;
	wire _w1617_ ;
	wire _w1618_ ;
	wire _w1619_ ;
	wire _w1620_ ;
	wire _w1621_ ;
	wire _w1622_ ;
	wire _w1623_ ;
	wire _w1624_ ;
	wire _w1625_ ;
	wire _w1626_ ;
	wire _w1627_ ;
	wire _w1628_ ;
	wire _w1629_ ;
	wire _w1630_ ;
	wire _w1631_ ;
	wire _w1632_ ;
	wire _w1633_ ;
	wire _w1634_ ;
	wire _w1635_ ;
	wire _w1766_ ;
	wire _w1767_ ;
	wire _w1768_ ;
	wire _w1769_ ;
	wire _w1770_ ;
	wire _w1771_ ;
	wire _w1772_ ;
	wire _w1773_ ;
	wire _w1774_ ;
	wire _w1775_ ;
	wire _w1776_ ;
	wire _w1777_ ;
	wire _w1778_ ;
	wire _w1779_ ;
	wire _w1780_ ;
	wire _w1781_ ;
	wire _w1782_ ;
	wire _w1783_ ;
	wire _w1784_ ;
	wire _w1785_ ;
	wire _w1786_ ;
	wire _w1787_ ;
	wire _w1788_ ;
	wire _w1789_ ;
	wire _w1790_ ;
	wire _w1791_ ;
	wire _w1792_ ;
	wire _w1793_ ;
	wire _w1794_ ;
	wire _w1795_ ;
	wire _w1796_ ;
	wire _w1797_ ;
	wire _w1798_ ;
	wire _w1799_ ;
	wire _w1800_ ;
	wire _w1801_ ;
	wire _w1802_ ;
	wire _w1803_ ;
	wire _w1804_ ;
	wire _w1805_ ;
	wire _w1806_ ;
	wire _w1807_ ;
	wire _w1808_ ;
	wire _w1809_ ;
	wire _w1810_ ;
	wire _w1811_ ;
	wire _w1812_ ;
	wire _w1813_ ;
	wire _w1814_ ;
	wire _w1815_ ;
	wire _w1816_ ;
	wire _w1817_ ;
	wire _w1818_ ;
	wire _w1819_ ;
	wire _w1820_ ;
	wire _w1821_ ;
	wire _w1822_ ;
	wire _w1823_ ;
	wire _w1824_ ;
	wire _w1825_ ;
	wire _w1826_ ;
	wire _w1827_ ;
	wire _w1828_ ;
	wire _w1829_ ;
	wire _w1830_ ;
	wire _w1831_ ;
	wire _w1832_ ;
	wire _w1833_ ;
	wire _w1834_ ;
	wire _w1835_ ;
	wire _w1836_ ;
	wire _w1837_ ;
	wire _w1838_ ;
	wire _w1839_ ;
	wire _w1840_ ;
	wire _w1841_ ;
	wire _w1842_ ;
	wire _w1843_ ;
	wire _w1844_ ;
	wire _w1845_ ;
	wire _w1846_ ;
	wire _w1847_ ;
	wire _w1848_ ;
	wire _w1849_ ;
	wire _w1850_ ;
	wire _w1851_ ;
	wire _w1852_ ;
	wire _w1853_ ;
	wire _w1854_ ;
	wire _w1855_ ;
	wire _w1856_ ;
	wire _w1857_ ;
	wire _w1858_ ;
	wire _w1859_ ;
	wire _w1860_ ;
	wire _w1861_ ;
	wire _w1862_ ;
	wire _w1863_ ;
	wire _w1864_ ;
	wire _w1865_ ;
	wire _w1866_ ;
	wire _w1867_ ;
	wire _w1868_ ;
	wire _w1869_ ;
	wire _w1870_ ;
	wire _w1871_ ;
	wire _w1872_ ;
	wire _w1873_ ;
	wire _w1874_ ;
	wire _w1875_ ;
	wire _w1876_ ;
	wire _w1877_ ;
	wire _w1878_ ;
	wire _w1879_ ;
	wire _w1880_ ;
	wire _w1881_ ;
	wire _w1882_ ;
	wire _w1883_ ;
	wire _w1884_ ;
	wire _w1885_ ;
	wire _w1886_ ;
	wire _w1887_ ;
	wire _w1888_ ;
	wire _w1889_ ;
	wire _w1890_ ;
	wire _w1891_ ;
	wire _w1892_ ;
	wire _w1893_ ;
	wire _w1894_ ;
	wire _w1895_ ;
	wire _w1896_ ;
	wire _w1897_ ;
	wire _w1898_ ;
	wire _w1899_ ;
	wire _w1900_ ;
	wire _w1901_ ;
	wire _w1902_ ;
	wire _w1903_ ;
	wire _w1904_ ;
	wire _w1905_ ;
	wire _w1906_ ;
	wire _w1907_ ;
	wire _w1908_ ;
	wire _w1909_ ;
	wire _w1910_ ;
	wire _w1911_ ;
	wire _w1912_ ;
	wire _w1913_ ;
	wire _w1914_ ;
	wire _w1915_ ;
	wire _w1916_ ;
	wire _w1917_ ;
	wire _w1918_ ;
	wire _w1919_ ;
	wire _w1920_ ;
	wire _w1921_ ;
	wire _w1922_ ;
	wire _w1923_ ;
	wire _w1924_ ;
	wire _w1925_ ;
	wire _w1926_ ;
	wire _w1927_ ;
	wire _w1928_ ;
	wire _w1929_ ;
	wire _w1930_ ;
	wire _w1931_ ;
	wire _w1932_ ;
	wire _w1933_ ;
	wire _w1934_ ;
	wire _w1935_ ;
	wire _w1936_ ;
	wire _w1937_ ;
	wire _w1938_ ;
	wire _w1939_ ;
	wire _w1940_ ;
	wire _w1941_ ;
	wire _w1942_ ;
	wire _w1943_ ;
	wire _w1944_ ;
	wire _w1945_ ;
	wire _w1946_ ;
	wire _w1947_ ;
	wire _w1948_ ;
	wire _w1949_ ;
	wire _w1950_ ;
	wire _w1951_ ;
	wire _w1952_ ;
	wire _w1953_ ;
	wire _w1954_ ;
	wire _w1955_ ;
	wire _w1956_ ;
	wire _w1957_ ;
	wire _w1958_ ;
	wire _w1959_ ;
	wire _w1960_ ;
	wire _w1961_ ;
	wire _w1962_ ;
	wire _w1963_ ;
	wire _w1964_ ;
	wire _w1965_ ;
	wire _w1966_ ;
	wire _w1967_ ;
	wire _w1968_ ;
	wire _w1969_ ;
	wire _w1970_ ;
	wire _w1971_ ;
	wire _w1972_ ;
	wire _w1973_ ;
	wire _w1974_ ;
	wire _w1975_ ;
	wire _w1976_ ;
	wire _w1977_ ;
	wire _w1978_ ;
	wire _w1979_ ;
	wire _w1980_ ;
	wire _w1981_ ;
	wire _w1982_ ;
	wire _w1983_ ;
	wire _w1984_ ;
	wire _w1985_ ;
	wire _w1986_ ;
	wire _w1987_ ;
	wire _w1988_ ;
	wire _w1989_ ;
	wire _w1990_ ;
	wire _w1991_ ;
	wire _w1992_ ;
	wire _w1993_ ;
	wire _w1994_ ;
	wire _w1995_ ;
	wire _w1996_ ;
	wire _w1997_ ;
	wire _w1998_ ;
	wire _w1999_ ;
	wire _w2000_ ;
	wire _w2001_ ;
	wire _w2002_ ;
	wire _w2003_ ;
	wire _w2004_ ;
	wire _w2005_ ;
	wire _w2006_ ;
	wire _w2007_ ;
	wire _w2008_ ;
	wire _w2009_ ;
	wire _w2010_ ;
	wire _w2011_ ;
	wire _w2012_ ;
	wire _w2013_ ;
	wire _w2014_ ;
	wire _w2015_ ;
	wire _w2016_ ;
	wire _w2017_ ;
	wire _w2018_ ;
	wire _w2019_ ;
	wire _w2020_ ;
	wire _w2021_ ;
	wire _w2022_ ;
	wire _w2023_ ;
	wire _w2024_ ;
	wire _w2025_ ;
	wire _w2026_ ;
	wire _w2027_ ;
	wire _w2028_ ;
	wire _w2029_ ;
	wire _w2030_ ;
	wire _w2031_ ;
	wire _w2032_ ;
	wire _w2033_ ;
	wire _w2034_ ;
	wire _w2035_ ;
	wire _w2036_ ;
	wire _w2037_ ;
	wire _w2038_ ;
	wire _w2039_ ;
	wire _w2040_ ;
	wire _w2041_ ;
	wire _w2042_ ;
	wire _w2043_ ;
	wire _w2044_ ;
	wire _w2045_ ;
	wire _w2046_ ;
	wire _w2047_ ;
	wire _w2048_ ;
	wire _w2049_ ;
	wire _w2618_ ;
	wire _w2619_ ;
	wire _w2620_ ;
	wire _w2621_ ;
	wire _w2622_ ;
	wire _w2623_ ;
	wire _w2624_ ;
	wire _w2625_ ;
	wire _w2626_ ;
	wire _w2627_ ;
	wire _w2628_ ;
	wire _w2629_ ;
	wire _w2630_ ;
	wire _w2631_ ;
	wire _w2632_ ;
	wire _w2633_ ;
	wire _w2634_ ;
	wire _w2635_ ;
	wire _w2636_ ;
	wire _w2637_ ;
	wire _w2638_ ;
	wire _w2639_ ;
	wire _w2640_ ;
	wire _w2641_ ;
	wire _w2642_ ;
	wire _w2643_ ;
	wire _w2644_ ;
	wire _w2645_ ;
	wire _w2646_ ;
	wire _w2647_ ;
	wire _w2648_ ;
	wire _w2649_ ;
	wire _w2650_ ;
	wire _w2651_ ;
	wire _w2652_ ;
	wire _w2653_ ;
	wire _w2654_ ;
	wire _w2655_ ;
	wire _w2656_ ;
	wire _w2657_ ;
	wire _w2658_ ;
	wire _w2659_ ;
	wire _w2660_ ;
	wire _w2661_ ;
	wire _w2662_ ;
	wire _w2663_ ;
	wire _w2664_ ;
	wire _w2665_ ;
	wire _w2666_ ;
	wire _w2667_ ;
	wire _w2668_ ;
	wire _w2669_ ;
	wire _w2670_ ;
	wire _w2671_ ;
	wire _w2672_ ;
	wire _w2673_ ;
	wire _w2674_ ;
	wire _w2675_ ;
	wire _w2676_ ;
	wire _w2677_ ;
	wire _w2678_ ;
	wire _w2679_ ;
	wire _w2680_ ;
	wire _w2681_ ;
	wire _w2682_ ;
	wire _w2683_ ;
	wire _w2684_ ;
	wire _w2685_ ;
	wire _w2686_ ;
	wire _w2687_ ;
	wire _w2688_ ;
	wire _w2689_ ;
	wire _w2690_ ;
	wire _w2691_ ;
	wire _w2692_ ;
	wire _w2693_ ;
	wire _w2694_ ;
	wire _w2695_ ;
	wire _w2696_ ;
	wire _w2697_ ;
	wire _w2698_ ;
	wire _w2699_ ;
	wire _w2700_ ;
	wire _w2701_ ;
	wire _w2702_ ;
	wire _w2703_ ;
	wire _w2704_ ;
	wire _w2705_ ;
	wire _w2706_ ;
	wire _w2707_ ;
	wire _w2708_ ;
	wire _w2709_ ;
	wire _w2710_ ;
	wire _w2711_ ;
	wire _w2712_ ;
	wire _w2713_ ;
	wire _w2714_ ;
	wire _w2715_ ;
	wire _w2716_ ;
	wire _w2717_ ;
	wire _w2718_ ;
	wire _w2719_ ;
	wire _w2720_ ;
	wire _w2721_ ;
	wire _w2722_ ;
	wire _w2723_ ;
	wire _w2724_ ;
	wire _w2725_ ;
	wire _w2726_ ;
	wire _w2727_ ;
	wire _w2728_ ;
	wire _w2729_ ;
	wire _w2730_ ;
	wire _w2731_ ;
	wire _w2732_ ;
	wire _w2733_ ;
	wire _w2734_ ;
	wire _w2735_ ;
	wire _w2736_ ;
	wire _w2737_ ;
	wire _w2738_ ;
	wire _w2739_ ;
	wire _w2740_ ;
	wire _w2741_ ;
	wire _w2742_ ;
	wire _w2743_ ;
	wire _w2744_ ;
	wire _w2745_ ;
	wire _w2746_ ;
	wire _w2747_ ;
	wire _w2748_ ;
	wire _w2749_ ;
	wire _w2750_ ;
	wire _w2751_ ;
	wire _w2752_ ;
	wire _w2753_ ;
	wire _w2754_ ;
	wire _w2755_ ;
	wire _w2756_ ;
	wire _w2757_ ;
	wire _w2758_ ;
	wire _w2759_ ;
	wire _w2760_ ;
	wire _w2761_ ;
	wire _w2762_ ;
	wire _w2763_ ;
	wire _w2764_ ;
	wire _w2765_ ;
	wire _w2766_ ;
	wire _w2767_ ;
	wire _w2768_ ;
	wire _w2769_ ;
	wire _w2770_ ;
	wire _w2771_ ;
	wire _w2772_ ;
	wire _w2773_ ;
	wire _w2774_ ;
	wire _w2775_ ;
	wire _w2776_ ;
	wire _w2777_ ;
	wire _w2778_ ;
	wire _w2779_ ;
	wire _w2780_ ;
	wire _w2781_ ;
	wire _w2782_ ;
	wire _w2783_ ;
	wire _w2784_ ;
	wire _w2785_ ;
	wire _w2786_ ;
	wire _w2787_ ;
	wire _w2788_ ;
	wire _w2789_ ;
	wire _w2790_ ;
	wire _w2791_ ;
	wire _w2792_ ;
	wire _w2793_ ;
	wire _w2794_ ;
	wire _w2795_ ;
	wire _w2796_ ;
	wire _w2797_ ;
	wire _w2798_ ;
	wire _w2799_ ;
	wire _w2800_ ;
	wire _w2801_ ;
	wire _w2802_ ;
	wire _w2803_ ;
	wire _w2804_ ;
	wire _w2805_ ;
	wire _w2806_ ;
	wire _w2807_ ;
	wire _w2808_ ;
	wire _w2809_ ;
	wire _w2810_ ;
	wire _w2811_ ;
	wire _w2812_ ;
	wire _w2813_ ;
	wire _w2814_ ;
	wire _w2815_ ;
	wire _w2816_ ;
	wire _w2817_ ;
	wire _w2818_ ;
	wire _w2819_ ;
	wire _w2820_ ;
	wire _w2821_ ;
	wire _w2822_ ;
	wire _w2823_ ;
	wire _w2824_ ;
	wire _w2825_ ;
	wire _w2826_ ;
	wire _w2827_ ;
	wire _w2828_ ;
	wire _w2829_ ;
	wire _w2830_ ;
	wire _w2831_ ;
	wire _w2832_ ;
	wire _w2833_ ;
	wire _w2834_ ;
	wire _w2835_ ;
	wire _w2836_ ;
	wire _w2837_ ;
	wire _w2838_ ;
	wire _w2839_ ;
	wire _w2840_ ;
	wire _w2841_ ;
	wire _w2842_ ;
	wire _w2843_ ;
	wire _w2844_ ;
	wire _w2845_ ;
	wire _w2846_ ;
	wire _w2847_ ;
	wire _w2848_ ;
	wire _w2849_ ;
	wire _w2850_ ;
	wire _w2851_ ;
	wire _w2852_ ;
	wire _w2853_ ;
	wire _w2854_ ;
	wire _w2855_ ;
	wire _w2856_ ;
	wire _w2857_ ;
	wire _w2858_ ;
	wire _w2859_ ;
	wire _w2860_ ;
	wire _w2861_ ;
	wire _w2862_ ;
	wire _w2863_ ;
	wire _w2864_ ;
	wire _w2865_ ;
	wire _w2866_ ;
	wire _w2867_ ;
	wire _w2868_ ;
	wire _w2869_ ;
	wire _w2870_ ;
	wire _w2871_ ;
	wire _w2872_ ;
	wire _w2873_ ;
	wire _w2874_ ;
	wire _w2875_ ;
	wire _w2876_ ;
	wire _w2877_ ;
	wire _w2878_ ;
	wire _w2879_ ;
	wire _w2880_ ;
	wire _w2881_ ;
	wire _w2882_ ;
	wire _w2883_ ;
	wire _w2884_ ;
	wire _w2885_ ;
	wire _w2886_ ;
	wire _w2887_ ;
	wire _w2888_ ;
	wire _w2889_ ;
	wire _w2890_ ;
	wire _w2891_ ;
	wire _w2892_ ;
	wire _w2893_ ;
	wire _w2894_ ;
	wire _w2895_ ;
	wire _w2896_ ;
	wire _w2897_ ;
	wire _w2898_ ;
	wire _w2899_ ;
	wire _w2900_ ;
	wire _w2901_ ;
	wire _w2902_ ;
	wire _w2903_ ;
	wire _w2904_ ;
	wire _w2905_ ;
	wire _w2906_ ;
	wire _w2907_ ;
	wire _w2908_ ;
	wire _w2909_ ;
	wire _w2910_ ;
	wire _w2911_ ;
	wire _w2912_ ;
	wire _w2913_ ;
	wire _w2914_ ;
	wire _w2915_ ;
	wire _w2916_ ;
	wire _w2917_ ;
	wire _w2918_ ;
	wire _w2919_ ;
	wire _w2920_ ;
	wire _w2921_ ;
	wire _w2922_ ;
	wire _w2923_ ;
	wire _w2924_ ;
	wire _w2925_ ;
	wire _w2926_ ;
	wire _w2927_ ;
	wire _w2928_ ;
	wire _w2929_ ;
	wire _w2930_ ;
	wire _w2931_ ;
	wire _w2932_ ;
	wire _w2933_ ;
	wire _w2934_ ;
	wire _w2935_ ;
	wire _w2936_ ;
	wire _w2937_ ;
	wire _w2938_ ;
	wire _w2939_ ;
	wire _w2940_ ;
	wire _w2941_ ;
	wire _w2942_ ;
	wire _w2943_ ;
	wire _w2944_ ;
	wire _w2945_ ;
	wire _w2946_ ;
	wire _w2947_ ;
	wire _w2948_ ;
	wire _w2949_ ;
	wire _w2950_ ;
	wire _w2951_ ;
	wire _w2952_ ;
	wire _w2953_ ;
	wire _w2954_ ;
	wire _w2955_ ;
	wire _w2956_ ;
	wire _w2957_ ;
	wire _w2958_ ;
	wire _w2959_ ;
	wire _w2960_ ;
	wire _w2961_ ;
	wire _w2962_ ;
	wire _w2963_ ;
	wire _w2964_ ;
	wire _w2965_ ;
	wire _w2966_ ;
	wire _w2967_ ;
	wire _w2968_ ;
	wire _w2969_ ;
	wire _w2970_ ;
	wire _w2971_ ;
	wire _w2972_ ;
	wire _w2973_ ;
	wire _w2974_ ;
	wire _w2975_ ;
	wire _w2976_ ;
	wire _w2977_ ;
	wire _w2978_ ;
	wire _w2979_ ;
	wire _w2980_ ;
	wire _w2981_ ;
	wire _w2982_ ;
	wire _w2983_ ;
	wire _w2984_ ;
	wire _w2985_ ;
	wire _w2986_ ;
	wire _w2987_ ;
	wire _w2988_ ;
	wire _w2989_ ;
	wire _w2990_ ;
	wire _w2991_ ;
	wire _w2992_ ;
	wire _w2993_ ;
	wire _w2994_ ;
	wire _w2995_ ;
	wire _w2996_ ;
	wire _w2997_ ;
	wire _w2998_ ;
	wire _w2999_ ;
	wire _w3000_ ;
	wire _w3001_ ;
	wire _w3002_ ;
	wire _w3003_ ;
	wire _w3004_ ;
	wire _w3005_ ;
	wire _w3006_ ;
	wire _w3007_ ;
	wire _w3008_ ;
	wire _w3009_ ;
	wire _w3010_ ;
	wire _w3011_ ;
	wire _w3012_ ;
	wire _w3013_ ;
	wire _w3014_ ;
	wire _w3015_ ;
	wire _w3016_ ;
	wire _w3017_ ;
	wire _w3018_ ;
	wire _w3019_ ;
	wire _w3020_ ;
	wire _w3021_ ;
	wire _w3022_ ;
	wire _w3023_ ;
	wire _w3024_ ;
	wire _w3025_ ;
	wire _w3026_ ;
	wire _w3027_ ;
	wire _w3028_ ;
	wire _w3029_ ;
	wire _w3030_ ;
	wire _w3031_ ;
	wire _w3032_ ;
	wire _w3033_ ;
	wire _w3034_ ;
	wire _w3035_ ;
	wire _w3036_ ;
	wire _w3037_ ;
	wire _w3038_ ;
	wire _w3039_ ;
	wire _w3040_ ;
	wire _w3041_ ;
	wire _w3042_ ;
	wire _w3043_ ;
	wire _w3044_ ;
	wire _w3045_ ;
	wire _w3046_ ;
	wire _w3047_ ;
	wire _w3048_ ;
	wire _w3049_ ;
	wire _w3050_ ;
	wire _w3051_ ;
	wire _w3052_ ;
	wire _w3053_ ;
	wire _w3054_ ;
	wire _w3055_ ;
	wire _w3056_ ;
	wire _w3057_ ;
	wire _w3058_ ;
	wire _w3059_ ;
	wire _w3060_ ;
	wire _w3061_ ;
	wire _w3062_ ;
	wire _w3063_ ;
	wire _w3064_ ;
	wire _w3065_ ;
	wire _w3066_ ;
	wire _w3067_ ;
	wire _w3068_ ;
	wire _w3069_ ;
	wire _w3070_ ;
	wire _w3071_ ;
	wire _w3072_ ;
	wire _w3073_ ;
	wire _w3074_ ;
	wire _w3075_ ;
	wire _w3076_ ;
	wire _w3077_ ;
	wire _w3078_ ;
	wire _w3079_ ;
	wire _w3080_ ;
	wire _w3081_ ;
	wire _w3082_ ;
	wire _w3083_ ;
	wire _w3084_ ;
	wire _w3085_ ;
	wire _w3086_ ;
	wire _w3087_ ;
	wire _w3088_ ;
	wire _w3089_ ;
	wire _w3090_ ;
	wire _w3091_ ;
	wire _w3092_ ;
	wire _w3093_ ;
	wire _w3094_ ;
	wire _w3095_ ;
	wire _w3096_ ;
	wire _w3097_ ;
	wire _w3098_ ;
	wire _w3099_ ;
	wire _w3100_ ;
	wire _w3101_ ;
	wire _w3102_ ;
	wire _w3103_ ;
	wire _w3104_ ;
	wire _w3105_ ;
	wire _w3106_ ;
	wire _w3107_ ;
	wire _w3108_ ;
	wire _w3109_ ;
	wire _w3110_ ;
	wire _w3111_ ;
	wire _w3112_ ;
	wire _w3113_ ;
	wire _w3114_ ;
	wire _w3115_ ;
	wire _w3116_ ;
	wire _w3117_ ;
	wire _w3118_ ;
	wire _w3119_ ;
	wire _w3120_ ;
	wire _w3121_ ;
	wire _w3122_ ;
	wire _w3123_ ;
	wire _w3124_ ;
	wire _w3125_ ;
	wire _w3126_ ;
	wire _w3127_ ;
	wire _w3128_ ;
	wire _w3129_ ;
	wire _w3130_ ;
	wire _w3131_ ;
	wire _w3132_ ;
	wire _w3133_ ;
	wire _w3134_ ;
	wire _w3135_ ;
	wire _w3136_ ;
	wire _w3137_ ;
	wire _w3138_ ;
	wire _w3139_ ;
	wire _w3140_ ;
	wire _w3141_ ;
	wire _w3142_ ;
	wire _w3143_ ;
	wire _w3144_ ;
	wire _w3145_ ;
	wire _w3146_ ;
	wire _w3147_ ;
	wire _w3148_ ;
	wire _w3149_ ;
	wire _w3150_ ;
	wire _w3151_ ;
	wire _w3152_ ;
	wire _w3153_ ;
	wire _w3154_ ;
	wire _w3155_ ;
	wire _w3156_ ;
	wire _w3157_ ;
	wire _w3158_ ;
	wire _w3159_ ;
	wire _w3160_ ;
	wire _w3161_ ;
	wire _w3162_ ;
	wire _w3163_ ;
	wire _w3164_ ;
	wire _w3165_ ;
	wire _w3166_ ;
	wire _w3167_ ;
	wire _w3168_ ;
	wire _w3169_ ;
	wire _w3170_ ;
	wire _w3171_ ;
	wire _w3172_ ;
	wire _w3173_ ;
	wire _w3174_ ;
	wire _w3175_ ;
	wire _w3176_ ;
	wire _w3177_ ;
	wire _w3178_ ;
	wire _w3179_ ;
	wire _w3180_ ;
	wire _w3181_ ;
	wire _w3182_ ;
	wire _w3183_ ;
	wire _w3184_ ;
	wire _w3185_ ;
	wire _w3186_ ;
	wire _w3187_ ;
	wire _w3188_ ;
	wire _w3189_ ;
	wire _w3190_ ;
	wire _w3191_ ;
	wire _w3192_ ;
	wire _w3193_ ;
	wire _w3194_ ;
	wire _w3195_ ;
	wire _w3196_ ;
	wire _w3197_ ;
	wire _w3198_ ;
	wire _w3199_ ;
	wire _w3200_ ;
	wire _w3201_ ;
	wire _w3202_ ;
	wire _w3203_ ;
	wire _w3204_ ;
	wire _w3205_ ;
	wire _w3206_ ;
	wire _w3207_ ;
	wire _w3208_ ;
	wire _w3209_ ;
	wire _w3210_ ;
	wire _w3211_ ;
	wire _w3212_ ;
	wire _w3213_ ;
	wire _w3214_ ;
	wire _w3215_ ;
	wire _w3216_ ;
	wire _w3217_ ;
	wire _w3218_ ;
	wire _w3219_ ;
	wire _w3220_ ;
	wire _w3221_ ;
	wire _w3222_ ;
	wire _w3223_ ;
	wire _w3224_ ;
	wire _w3225_ ;
	wire _w3226_ ;
	wire _w3227_ ;
	wire _w3228_ ;
	wire _w3229_ ;
	wire _w3230_ ;
	wire _w3231_ ;
	wire _w3232_ ;
	wire _w3233_ ;
	wire _w3234_ ;
	wire _w3235_ ;
	wire _w3236_ ;
	wire _w3237_ ;
	wire _w3238_ ;
	wire _w3239_ ;
	wire _w3240_ ;
	wire _w3241_ ;
	wire _w3242_ ;
	wire _w3243_ ;
	wire _w3244_ ;
	wire _w3245_ ;
	wire _w3246_ ;
	wire _w3247_ ;
	wire _w3248_ ;
	wire _w3249_ ;
	wire _w3250_ ;
	wire _w3251_ ;
	wire _w3252_ ;
	wire _w3253_ ;
	wire _w3254_ ;
	wire _w3255_ ;
	wire _w3256_ ;
	wire _w3257_ ;
	wire _w3258_ ;
	wire _w3259_ ;
	wire _w3260_ ;
	wire _w3261_ ;
	wire _w3262_ ;
	wire _w3263_ ;
	wire _w3264_ ;
	wire _w3265_ ;
	wire _w3266_ ;
	wire _w3267_ ;
	wire _w3268_ ;
	wire _w3269_ ;
	wire _w3270_ ;
	wire _w3271_ ;
	wire _w3272_ ;
	wire _w3273_ ;
	wire _w3274_ ;
	wire _w3275_ ;
	wire _w3276_ ;
	wire _w3277_ ;
	wire _w3278_ ;
	wire _w3279_ ;
	wire _w3280_ ;
	wire _w3281_ ;
	wire _w3282_ ;
	wire _w3283_ ;
	wire _w3284_ ;
	wire _w3285_ ;
	wire _w3286_ ;
	wire _w3287_ ;
	wire _w3288_ ;
	wire _w3289_ ;
	wire _w3290_ ;
	wire _w3291_ ;
	wire _w3292_ ;
	wire _w3293_ ;
	wire _w3294_ ;
	wire _w3295_ ;
	wire _w3296_ ;
	wire _w3297_ ;
	wire _w3298_ ;
	wire _w3299_ ;
	wire _w3300_ ;
	wire _w3301_ ;
	wire _w3302_ ;
	wire _w3303_ ;
	wire _w3304_ ;
	wire _w3305_ ;
	wire _w3306_ ;
	wire _w3307_ ;
	wire _w3308_ ;
	wire _w3309_ ;
	wire _w3310_ ;
	wire _w3311_ ;
	wire _w3312_ ;
	wire _w3313_ ;
	wire _w3314_ ;
	wire _w3315_ ;
	wire _w3316_ ;
	wire _w3317_ ;
	wire _w3318_ ;
	wire _w3319_ ;
	wire _w3320_ ;
	wire _w3321_ ;
	wire _w3322_ ;
	wire _w3323_ ;
	wire _w3324_ ;
	wire _w3325_ ;
	wire _w3326_ ;
	wire _w3327_ ;
	wire _w3328_ ;
	wire _w3329_ ;
	wire _w3330_ ;
	wire _w3331_ ;
	wire _w3332_ ;
	wire _w3333_ ;
	wire _w3334_ ;
	wire _w3335_ ;
	wire _w3336_ ;
	wire _w3337_ ;
	wire _w3338_ ;
	wire _w3339_ ;
	wire _w3340_ ;
	wire _w3341_ ;
	wire _w3342_ ;
	wire _w3343_ ;
	wire _w3344_ ;
	wire _w3345_ ;
	wire _w3346_ ;
	wire _w3347_ ;
	wire _w3348_ ;
	wire _w3349_ ;
	wire _w3350_ ;
	wire _w3351_ ;
	wire _w3352_ ;
	wire _w3353_ ;
	wire _w3354_ ;
	wire _w3355_ ;
	wire _w3356_ ;
	wire _w3357_ ;
	wire _w3358_ ;
	wire _w3359_ ;
	wire _w3360_ ;
	wire _w3361_ ;
	wire _w3362_ ;
	wire _w3363_ ;
	wire _w3364_ ;
	wire _w3365_ ;
	wire _w3366_ ;
	wire _w3367_ ;
	wire _w3368_ ;
	wire _w3369_ ;
	wire _w3370_ ;
	wire _w3371_ ;
	wire _w3372_ ;
	wire _w3373_ ;
	wire _w3374_ ;
	wire _w3375_ ;
	wire _w3376_ ;
	wire _w3377_ ;
	wire _w3378_ ;
	wire _w3379_ ;
	wire _w3380_ ;
	wire _w3381_ ;
	wire _w3382_ ;
	wire _w3383_ ;
	wire _w3384_ ;
	wire _w3385_ ;
	wire _w3386_ ;
	wire _w3387_ ;
	wire _w3388_ ;
	wire _w3389_ ;
	wire _w3390_ ;
	wire _w3391_ ;
	wire _w3392_ ;
	wire _w3393_ ;
	wire _w3394_ ;
	wire _w3395_ ;
	wire _w3396_ ;
	wire _w3397_ ;
	wire _w3398_ ;
	wire _w3399_ ;
	wire _w3400_ ;
	wire _w3401_ ;
	wire _w3402_ ;
	wire _w3403_ ;
	wire _w3404_ ;
	wire _w3405_ ;
	wire _w3406_ ;
	wire _w3407_ ;
	wire _w3408_ ;
	wire _w3409_ ;
	wire _w3410_ ;
	wire _w3411_ ;
	wire _w3412_ ;
	wire _w3413_ ;
	wire _w3414_ ;
	wire _w3415_ ;
	wire _w3416_ ;
	wire _w3417_ ;
	wire _w3418_ ;
	wire _w3419_ ;
	wire _w3420_ ;
	wire _w3421_ ;
	wire _w3422_ ;
	wire _w3423_ ;
	wire _w3424_ ;
	wire _w3425_ ;
	wire _w3426_ ;
	wire _w3427_ ;
	wire _w3428_ ;
	wire _w3429_ ;
	wire _w3430_ ;
	wire _w3431_ ;
	wire _w3432_ ;
	wire _w3433_ ;
	wire _w3434_ ;
	wire _w3435_ ;
	wire _w3436_ ;
	wire _w3437_ ;
	wire _w3438_ ;
	wire _w3439_ ;
	wire _w3440_ ;
	wire _w3441_ ;
	wire _w3442_ ;
	wire _w3443_ ;
	wire _w3444_ ;
	wire _w3445_ ;
	wire _w3446_ ;
	wire _w3447_ ;
	wire _w3448_ ;
	wire _w3449_ ;
	wire _w3450_ ;
	wire _w3451_ ;
	wire _w3452_ ;
	wire _w3453_ ;
	wire _w3454_ ;
	wire _w3455_ ;
	wire _w3456_ ;
	wire _w3457_ ;
	wire _w3458_ ;
	wire _w3459_ ;
	wire _w3460_ ;
	wire _w3461_ ;
	wire _w3462_ ;
	wire _w3463_ ;
	wire _w3464_ ;
	wire _w3465_ ;
	wire _w3466_ ;
	wire _w3467_ ;
	wire _w3468_ ;
	wire _w3469_ ;
	wire _w3470_ ;
	wire _w3471_ ;
	wire _w3472_ ;
	wire _w3473_ ;
	wire _w3474_ ;
	wire _w3475_ ;
	wire _w3476_ ;
	wire _w3477_ ;
	wire _w3478_ ;
	wire _w3479_ ;
	wire _w3480_ ;
	wire _w3481_ ;
	wire _w3482_ ;
	wire _w3483_ ;
	wire _w3484_ ;
	wire _w3485_ ;
	wire _w3486_ ;
	wire _w3487_ ;
	wire _w3488_ ;
	wire _w3489_ ;
	wire _w3490_ ;
	wire _w3491_ ;
	wire _w3492_ ;
	wire _w3493_ ;
	wire _w3494_ ;
	wire _w3495_ ;
	wire _w3496_ ;
	wire _w3497_ ;
	wire _w3498_ ;
	wire _w3499_ ;
	wire _w3500_ ;
	wire _w3501_ ;
	wire _w3502_ ;
	wire _w3503_ ;
	wire _w3504_ ;
	wire _w3505_ ;
	wire _w3506_ ;
	wire _w3507_ ;
	wire _w3508_ ;
	wire _w3509_ ;
	wire _w3510_ ;
	wire _w3511_ ;
	wire _w3512_ ;
	wire _w3513_ ;
	wire _w3514_ ;
	wire _w3515_ ;
	wire _w3516_ ;
	wire _w3517_ ;
	wire _w3518_ ;
	wire _w3519_ ;
	wire _w3520_ ;
	wire _w3521_ ;
	wire _w3522_ ;
	wire _w3523_ ;
	wire _w3524_ ;
	wire _w3525_ ;
	wire _w3526_ ;
	wire _w3527_ ;
	wire _w3528_ ;
	wire _w3529_ ;
	wire _w3530_ ;
	wire _w3531_ ;
	wire _w3532_ ;
	wire _w3533_ ;
	wire _w3534_ ;
	wire _w3535_ ;
	wire _w3536_ ;
	wire _w3537_ ;
	wire _w3538_ ;
	wire _w3539_ ;
	wire _w3540_ ;
	wire _w3541_ ;
	wire _w3542_ ;
	wire _w3543_ ;
	wire _w3544_ ;
	wire _w3545_ ;
	wire _w3546_ ;
	wire _w3547_ ;
	wire _w3548_ ;
	wire _w3549_ ;
	wire _w3550_ ;
	wire _w3551_ ;
	wire _w3552_ ;
	wire _w3553_ ;
	wire _w3554_ ;
	wire _w3555_ ;
	wire _w3556_ ;
	wire _w3557_ ;
	wire _w3558_ ;
	wire _w3559_ ;
	wire _w3560_ ;
	wire _w3561_ ;
	wire _w3562_ ;
	wire _w3563_ ;
	wire _w3564_ ;
	wire _w3565_ ;
	wire _w3566_ ;
	wire _w3567_ ;
	wire _w3568_ ;
	wire _w3569_ ;
	wire _w3570_ ;
	wire _w3571_ ;
	wire _w3572_ ;
	wire _w3573_ ;
	wire _w3574_ ;
	wire _w3575_ ;
	wire _w3576_ ;
	wire _w3577_ ;
	wire _w3578_ ;
	wire _w3579_ ;
	wire _w3580_ ;
	wire _w3581_ ;
	wire _w3582_ ;
	wire _w3583_ ;
	wire _w3584_ ;
	wire _w3585_ ;
	wire _w3586_ ;
	wire _w3587_ ;
	wire _w3588_ ;
	wire _w3589_ ;
	wire _w3590_ ;
	wire _w3591_ ;
	wire _w3592_ ;
	wire _w3593_ ;
	wire _w3594_ ;
	wire _w3595_ ;
	wire _w3596_ ;
	wire _w3597_ ;
	wire _w3598_ ;
	wire _w3599_ ;
	wire _w3600_ ;
	wire _w3601_ ;
	wire _w3602_ ;
	wire _w3603_ ;
	wire _w3604_ ;
	wire _w3605_ ;
	wire _w3606_ ;
	wire _w3607_ ;
	wire _w3608_ ;
	wire _w3609_ ;
	wire _w3610_ ;
	wire _w3611_ ;
	wire _w3612_ ;
	wire _w3613_ ;
	wire _w3614_ ;
	wire _w3615_ ;
	wire _w3616_ ;
	wire _w3617_ ;
	wire _w3618_ ;
	wire _w3619_ ;
	wire _w3620_ ;
	wire _w3621_ ;
	wire _w3622_ ;
	wire _w3623_ ;
	wire _w3624_ ;
	wire _w3625_ ;
	wire _w3626_ ;
	wire _w3627_ ;
	wire _w3628_ ;
	wire _w3629_ ;
	wire _w3630_ ;
	wire _w3631_ ;
	wire _w3632_ ;
	wire _w3633_ ;
	wire _w3634_ ;
	wire _w3635_ ;
	wire _w3636_ ;
	wire _w3637_ ;
	wire _w3638_ ;
	wire _w3639_ ;
	wire _w3640_ ;
	wire _w3641_ ;
	wire _w3642_ ;
	wire _w3643_ ;
	wire _w3644_ ;
	wire _w3645_ ;
	wire _w3646_ ;
	wire _w3647_ ;
	wire _w3648_ ;
	wire _w3649_ ;
	wire _w3650_ ;
	wire _w3651_ ;
	wire _w3652_ ;
	wire _w3653_ ;
	wire _w3654_ ;
	wire _w3655_ ;
	wire _w3656_ ;
	wire _w3657_ ;
	wire _w3658_ ;
	wire _w3659_ ;
	wire _w3660_ ;
	wire _w3661_ ;
	wire _w3662_ ;
	wire _w3663_ ;
	wire _w3664_ ;
	wire _w3665_ ;
	wire _w3666_ ;
	wire _w3667_ ;
	wire _w3668_ ;
	wire _w3669_ ;
	wire _w3670_ ;
	wire _w3671_ ;
	wire _w3672_ ;
	wire _w3673_ ;
	wire _w3674_ ;
	wire _w3675_ ;
	wire _w3676_ ;
	wire _w3677_ ;
	wire _w3678_ ;
	wire _w3679_ ;
	wire _w3680_ ;
	wire _w3681_ ;
	wire _w3682_ ;
	wire _w3683_ ;
	wire _w3684_ ;
	wire _w3685_ ;
	wire _w3686_ ;
	wire _w3687_ ;
	wire _w3688_ ;
	wire _w3689_ ;
	wire _w3690_ ;
	wire _w3691_ ;
	wire _w3692_ ;
	wire _w3693_ ;
	wire _w3694_ ;
	wire _w3695_ ;
	wire _w3696_ ;
	wire _w3697_ ;
	wire _w3698_ ;
	wire _w3699_ ;
	wire _w3700_ ;
	wire _w3701_ ;
	wire _w3702_ ;
	wire _w3703_ ;
	wire _w3704_ ;
	wire _w3705_ ;
	wire _w3706_ ;
	wire _w3707_ ;
	wire _w3708_ ;
	wire _w3709_ ;
	wire _w3710_ ;
	wire _w3711_ ;
	wire _w3712_ ;
	wire _w3713_ ;
	wire _w3714_ ;
	wire _w3715_ ;
	wire _w3716_ ;
	wire _w3717_ ;
	wire _w3718_ ;
	wire _w3719_ ;
	wire _w3720_ ;
	wire _w3721_ ;
	wire _w3722_ ;
	wire _w3723_ ;
	wire _w3724_ ;
	wire _w3725_ ;
	wire _w3726_ ;
	wire _w3727_ ;
	wire _w3728_ ;
	wire _w3729_ ;
	wire _w3730_ ;
	wire _w3731_ ;
	wire _w3732_ ;
	wire _w3733_ ;
	wire _w3734_ ;
	wire _w3735_ ;
	wire _w3736_ ;
	wire _w3737_ ;
	wire _w3738_ ;
	wire _w3739_ ;
	wire _w3740_ ;
	wire _w3741_ ;
	wire _w3742_ ;
	wire _w3743_ ;
	wire _w3744_ ;
	wire _w3745_ ;
	wire _w3746_ ;
	wire _w3747_ ;
	wire _w3748_ ;
	wire _w3749_ ;
	wire _w3750_ ;
	wire _w3751_ ;
	wire _w3752_ ;
	wire _w3753_ ;
	wire _w3754_ ;
	wire _w3755_ ;
	wire _w3756_ ;
	wire _w3757_ ;
	wire _w3758_ ;
	wire _w3759_ ;
	wire _w3760_ ;
	wire _w3761_ ;
	wire _w3762_ ;
	wire _w3763_ ;
	wire _w3764_ ;
	wire _w3765_ ;
	wire _w3766_ ;
	wire _w3767_ ;
	wire _w3768_ ;
	wire _w3769_ ;
	wire _w3770_ ;
	wire _w3771_ ;
	wire _w3772_ ;
	wire _w3773_ ;
	wire _w3774_ ;
	wire _w3775_ ;
	wire _w3776_ ;
	wire _w3777_ ;
	wire _w3778_ ;
	wire _w3779_ ;
	wire _w3780_ ;
	wire _w3781_ ;
	wire _w3782_ ;
	wire _w3783_ ;
	wire _w3784_ ;
	wire _w3785_ ;
	wire _w3786_ ;
	wire _w3787_ ;
	wire _w3788_ ;
	wire _w3789_ ;
	wire _w3790_ ;
	wire _w3791_ ;
	wire _w3792_ ;
	wire _w3793_ ;
	wire _w3794_ ;
	wire _w3795_ ;
	wire _w3796_ ;
	wire _w3797_ ;
	wire _w3798_ ;
	wire _w3799_ ;
	wire _w3800_ ;
	wire _w3801_ ;
	wire _w3802_ ;
	wire _w3803_ ;
	wire _w3804_ ;
	wire _w3805_ ;
	wire _w3806_ ;
	wire _w3807_ ;
	wire _w3808_ ;
	wire _w3809_ ;
	wire _w3810_ ;
	wire _w3811_ ;
	wire _w3812_ ;
	wire _w3813_ ;
	wire _w3814_ ;
	wire _w3815_ ;
	wire _w3816_ ;
	wire _w3817_ ;
	wire _w3818_ ;
	wire _w3819_ ;
	wire _w3820_ ;
	wire _w3821_ ;
	wire _w3822_ ;
	wire _w3823_ ;
	wire _w3824_ ;
	wire _w3825_ ;
	wire _w3826_ ;
	wire _w3827_ ;
	wire _w3828_ ;
	wire _w3829_ ;
	wire _w3830_ ;
	wire _w3831_ ;
	wire _w3832_ ;
	wire _w3833_ ;
	wire _w3834_ ;
	wire _w3835_ ;
	wire _w3836_ ;
	wire _w3837_ ;
	wire _w3838_ ;
	wire _w3839_ ;
	wire _w3840_ ;
	wire _w3841_ ;
	wire _w3842_ ;
	wire _w3843_ ;
	wire _w3844_ ;
	wire _w3845_ ;
	wire _w3846_ ;
	wire _w3847_ ;
	wire _w3848_ ;
	wire _w3849_ ;
	wire _w3850_ ;
	wire _w3851_ ;
	wire _w3852_ ;
	wire _w3853_ ;
	wire _w3854_ ;
	wire _w3855_ ;
	wire _w3856_ ;
	wire _w3857_ ;
	wire _w3858_ ;
	wire _w3859_ ;
	wire _w3860_ ;
	wire _w3861_ ;
	wire _w3862_ ;
	wire _w3863_ ;
	wire _w3864_ ;
	wire _w3865_ ;
	LUT2 #(
		.INIT('h2)
	) name0 (
		\TM0_pad ,
		\WX10891_reg/NET0131 ,
		_w1509_
	);
	LUT4 #(
		.INIT('h6996)
	) name1 (
		\WX707_reg/NET0131 ,
		\WX771_reg/NET0131 ,
		\WX835_reg/NET0131 ,
		\WX899_reg/NET0131 ,
		_w1510_
	);
	LUT2 #(
		.INIT('h6)
	) name2 (
		_w1509_,
		_w1510_,
		_w1511_
	);
	LUT2 #(
		.INIT('h2)
	) name3 (
		\TM0_pad ,
		\WX10871_reg/NET0131 ,
		_w1512_
	);
	LUT4 #(
		.INIT('h6996)
	) name4 (
		\WX687_reg/NET0131 ,
		\WX751_reg/NET0131 ,
		\WX815_reg/NET0131 ,
		\WX879_reg/NET0131 ,
		_w1513_
	);
	LUT2 #(
		.INIT('h6)
	) name5 (
		_w1512_,
		_w1513_,
		_w1514_
	);
	LUT2 #(
		.INIT('h2)
	) name6 (
		\TM0_pad ,
		\WX10869_reg/NET0131 ,
		_w1515_
	);
	LUT4 #(
		.INIT('h6996)
	) name7 (
		\WX685_reg/NET0131 ,
		\WX749_reg/NET0131 ,
		\WX813_reg/NET0131 ,
		\WX877_reg/NET0131 ,
		_w1516_
	);
	LUT2 #(
		.INIT('h6)
	) name8 (
		_w1515_,
		_w1516_,
		_w1517_
	);
	LUT2 #(
		.INIT('h2)
	) name9 (
		\TM0_pad ,
		\WX10867_reg/NET0131 ,
		_w1518_
	);
	LUT4 #(
		.INIT('h6996)
	) name10 (
		\WX683_reg/NET0131 ,
		\WX747_reg/NET0131 ,
		\WX811_reg/NET0131 ,
		\WX875_reg/NET0131 ,
		_w1519_
	);
	LUT2 #(
		.INIT('h6)
	) name11 (
		_w1518_,
		_w1519_,
		_w1520_
	);
	LUT2 #(
		.INIT('h2)
	) name12 (
		\TM0_pad ,
		\WX10865_reg/NET0131 ,
		_w1521_
	);
	LUT4 #(
		.INIT('h6996)
	) name13 (
		\WX681_reg/NET0131 ,
		\WX745_reg/NET0131 ,
		\WX809_reg/NET0131 ,
		\WX873_reg/NET0131 ,
		_w1522_
	);
	LUT2 #(
		.INIT('h6)
	) name14 (
		_w1521_,
		_w1522_,
		_w1523_
	);
	LUT2 #(
		.INIT('h2)
	) name15 (
		\TM0_pad ,
		\WX10863_reg/NET0131 ,
		_w1524_
	);
	LUT4 #(
		.INIT('h6996)
	) name16 (
		\WX679_reg/NET0131 ,
		\WX743_reg/NET0131 ,
		\WX807_reg/NET0131 ,
		\WX871_reg/NET0131 ,
		_w1525_
	);
	LUT2 #(
		.INIT('h6)
	) name17 (
		_w1524_,
		_w1525_,
		_w1526_
	);
	LUT2 #(
		.INIT('h2)
	) name18 (
		\TM0_pad ,
		\WX10861_reg/NET0131 ,
		_w1527_
	);
	LUT4 #(
		.INIT('h6996)
	) name19 (
		\WX677_reg/NET0131 ,
		\WX741_reg/NET0131 ,
		\WX805_reg/NET0131 ,
		\WX869_reg/NET0131 ,
		_w1528_
	);
	LUT2 #(
		.INIT('h6)
	) name20 (
		_w1527_,
		_w1528_,
		_w1529_
	);
	LUT3 #(
		.INIT('h96)
	) name21 (
		\WX739_reg/NET0131 ,
		\WX803_reg/NET0131 ,
		\WX867_reg/NET0131 ,
		_w1530_
	);
	LUT4 #(
		.INIT('h6c93)
	) name22 (
		\TM0_pad ,
		\TM1_pad ,
		\WX10859_reg/NET0131 ,
		\WX675_reg/NET0131 ,
		_w1531_
	);
	LUT2 #(
		.INIT('h9)
	) name23 (
		_w1530_,
		_w1531_,
		_w1532_
	);
	LUT3 #(
		.INIT('h96)
	) name24 (
		\WX737_reg/NET0131 ,
		\WX801_reg/NET0131 ,
		\WX865_reg/NET0131 ,
		_w1533_
	);
	LUT4 #(
		.INIT('h6c93)
	) name25 (
		\TM0_pad ,
		\TM1_pad ,
		\WX10857_reg/NET0131 ,
		\WX673_reg/NET0131 ,
		_w1534_
	);
	LUT2 #(
		.INIT('h9)
	) name26 (
		_w1533_,
		_w1534_,
		_w1535_
	);
	LUT3 #(
		.INIT('h96)
	) name27 (
		\WX735_reg/NET0131 ,
		\WX799_reg/NET0131 ,
		\WX863_reg/NET0131 ,
		_w1536_
	);
	LUT4 #(
		.INIT('h6c93)
	) name28 (
		\TM0_pad ,
		\TM1_pad ,
		\WX10855_reg/NET0131 ,
		\WX671_reg/NET0131 ,
		_w1537_
	);
	LUT2 #(
		.INIT('h9)
	) name29 (
		_w1536_,
		_w1537_,
		_w1538_
	);
	LUT3 #(
		.INIT('h96)
	) name30 (
		\WX733_reg/NET0131 ,
		\WX797_reg/NET0131 ,
		\WX861_reg/NET0131 ,
		_w1539_
	);
	LUT4 #(
		.INIT('h6c93)
	) name31 (
		\TM0_pad ,
		\TM1_pad ,
		\WX10853_reg/NET0131 ,
		\WX669_reg/NET0131 ,
		_w1540_
	);
	LUT2 #(
		.INIT('h9)
	) name32 (
		_w1539_,
		_w1540_,
		_w1541_
	);
	LUT2 #(
		.INIT('h2)
	) name33 (
		\TM0_pad ,
		\WX10889_reg/NET0131 ,
		_w1542_
	);
	LUT4 #(
		.INIT('h6996)
	) name34 (
		\WX705_reg/NET0131 ,
		\WX769_reg/NET0131 ,
		\WX833_reg/NET0131 ,
		\WX897_reg/NET0131 ,
		_w1543_
	);
	LUT2 #(
		.INIT('h6)
	) name35 (
		_w1542_,
		_w1543_,
		_w1544_
	);
	LUT3 #(
		.INIT('h96)
	) name36 (
		\WX731_reg/NET0131 ,
		\WX795_reg/NET0131 ,
		\WX859_reg/NET0131 ,
		_w1545_
	);
	LUT4 #(
		.INIT('h6c93)
	) name37 (
		\TM0_pad ,
		\TM1_pad ,
		\WX10851_reg/NET0131 ,
		\WX667_reg/NET0131 ,
		_w1546_
	);
	LUT2 #(
		.INIT('h9)
	) name38 (
		_w1545_,
		_w1546_,
		_w1547_
	);
	LUT3 #(
		.INIT('h96)
	) name39 (
		\WX729_reg/NET0131 ,
		\WX793_reg/NET0131 ,
		\WX857_reg/NET0131 ,
		_w1548_
	);
	LUT4 #(
		.INIT('h6c93)
	) name40 (
		\TM0_pad ,
		\TM1_pad ,
		\WX10849_reg/NET0131 ,
		\WX665_reg/NET0131 ,
		_w1549_
	);
	LUT2 #(
		.INIT('h9)
	) name41 (
		_w1548_,
		_w1549_,
		_w1550_
	);
	LUT3 #(
		.INIT('h96)
	) name42 (
		\WX727_reg/NET0131 ,
		\WX791_reg/NET0131 ,
		\WX855_reg/NET0131 ,
		_w1551_
	);
	LUT4 #(
		.INIT('h6c93)
	) name43 (
		\TM0_pad ,
		\TM1_pad ,
		\WX10847_reg/NET0131 ,
		\WX663_reg/NET0131 ,
		_w1552_
	);
	LUT2 #(
		.INIT('h9)
	) name44 (
		_w1551_,
		_w1552_,
		_w1553_
	);
	LUT3 #(
		.INIT('h96)
	) name45 (
		\WX725_reg/NET0131 ,
		\WX789_reg/NET0131 ,
		\WX853_reg/NET0131 ,
		_w1554_
	);
	LUT4 #(
		.INIT('h6c93)
	) name46 (
		\TM0_pad ,
		\TM1_pad ,
		\WX10845_reg/NET0131 ,
		\WX661_reg/NET0131 ,
		_w1555_
	);
	LUT2 #(
		.INIT('h9)
	) name47 (
		_w1554_,
		_w1555_,
		_w1556_
	);
	LUT3 #(
		.INIT('h96)
	) name48 (
		\WX723_reg/NET0131 ,
		\WX787_reg/NET0131 ,
		\WX851_reg/NET0131 ,
		_w1557_
	);
	LUT4 #(
		.INIT('h6c93)
	) name49 (
		\TM0_pad ,
		\TM1_pad ,
		\WX10843_reg/NET0131 ,
		\WX659_reg/NET0131 ,
		_w1558_
	);
	LUT2 #(
		.INIT('h9)
	) name50 (
		_w1557_,
		_w1558_,
		_w1559_
	);
	LUT3 #(
		.INIT('h96)
	) name51 (
		\WX721_reg/NET0131 ,
		\WX785_reg/NET0131 ,
		\WX849_reg/NET0131 ,
		_w1560_
	);
	LUT4 #(
		.INIT('h6c93)
	) name52 (
		\TM0_pad ,
		\TM1_pad ,
		\WX10841_reg/NET0131 ,
		\WX657_reg/NET0131 ,
		_w1561_
	);
	LUT2 #(
		.INIT('h9)
	) name53 (
		_w1560_,
		_w1561_,
		_w1562_
	);
	LUT3 #(
		.INIT('h96)
	) name54 (
		\WX719_reg/NET0131 ,
		\WX783_reg/NET0131 ,
		\WX847_reg/NET0131 ,
		_w1563_
	);
	LUT4 #(
		.INIT('h6c93)
	) name55 (
		\TM0_pad ,
		\TM1_pad ,
		\WX10839_reg/NET0131 ,
		\WX655_reg/NET0131 ,
		_w1564_
	);
	LUT2 #(
		.INIT('h9)
	) name56 (
		_w1563_,
		_w1564_,
		_w1565_
	);
	LUT3 #(
		.INIT('h96)
	) name57 (
		\WX717_reg/NET0131 ,
		\WX781_reg/NET0131 ,
		\WX845_reg/NET0131 ,
		_w1566_
	);
	LUT4 #(
		.INIT('h6c93)
	) name58 (
		\TM0_pad ,
		\TM1_pad ,
		\WX10837_reg/NET0131 ,
		\WX653_reg/NET0131 ,
		_w1567_
	);
	LUT2 #(
		.INIT('h9)
	) name59 (
		_w1566_,
		_w1567_,
		_w1568_
	);
	LUT3 #(
		.INIT('h96)
	) name60 (
		\WX715_reg/NET0131 ,
		\WX779_reg/NET0131 ,
		\WX843_reg/NET0131 ,
		_w1569_
	);
	LUT4 #(
		.INIT('h6c93)
	) name61 (
		\TM0_pad ,
		\TM1_pad ,
		\WX10835_reg/NET0131 ,
		\WX651_reg/NET0131 ,
		_w1570_
	);
	LUT2 #(
		.INIT('h9)
	) name62 (
		_w1569_,
		_w1570_,
		_w1571_
	);
	LUT3 #(
		.INIT('h96)
	) name63 (
		\WX713_reg/NET0131 ,
		\WX777_reg/NET0131 ,
		\WX841_reg/NET0131 ,
		_w1572_
	);
	LUT4 #(
		.INIT('h6c93)
	) name64 (
		\TM0_pad ,
		\TM1_pad ,
		\WX10833_reg/NET0131 ,
		\WX649_reg/NET0131 ,
		_w1573_
	);
	LUT2 #(
		.INIT('h9)
	) name65 (
		_w1572_,
		_w1573_,
		_w1574_
	);
	LUT2 #(
		.INIT('h2)
	) name66 (
		\TM0_pad ,
		\WX10887_reg/NET0131 ,
		_w1575_
	);
	LUT4 #(
		.INIT('h6996)
	) name67 (
		\WX703_reg/NET0131 ,
		\WX767_reg/NET0131 ,
		\WX831_reg/NET0131 ,
		\WX895_reg/NET0131 ,
		_w1576_
	);
	LUT2 #(
		.INIT('h6)
	) name68 (
		_w1575_,
		_w1576_,
		_w1577_
	);
	LUT3 #(
		.INIT('h96)
	) name69 (
		\WX711_reg/NET0131 ,
		\WX775_reg/NET0131 ,
		\WX839_reg/NET0131 ,
		_w1578_
	);
	LUT4 #(
		.INIT('h6c93)
	) name70 (
		\TM0_pad ,
		\TM1_pad ,
		\WX10831_reg/NET0131 ,
		\WX647_reg/NET0131 ,
		_w1579_
	);
	LUT2 #(
		.INIT('h9)
	) name71 (
		_w1578_,
		_w1579_,
		_w1580_
	);
	LUT3 #(
		.INIT('h96)
	) name72 (
		\WX709_reg/NET0131 ,
		\WX773_reg/NET0131 ,
		\WX837_reg/NET0131 ,
		_w1581_
	);
	LUT4 #(
		.INIT('h6c93)
	) name73 (
		\TM0_pad ,
		\TM1_pad ,
		\WX10829_reg/NET0131 ,
		\WX645_reg/NET0131 ,
		_w1582_
	);
	LUT2 #(
		.INIT('h9)
	) name74 (
		_w1581_,
		_w1582_,
		_w1583_
	);
	LUT2 #(
		.INIT('h2)
	) name75 (
		\TM0_pad ,
		\WX10885_reg/NET0131 ,
		_w1584_
	);
	LUT4 #(
		.INIT('h6996)
	) name76 (
		\WX701_reg/NET0131 ,
		\WX765_reg/NET0131 ,
		\WX829_reg/NET0131 ,
		\WX893_reg/NET0131 ,
		_w1585_
	);
	LUT2 #(
		.INIT('h6)
	) name77 (
		_w1584_,
		_w1585_,
		_w1586_
	);
	LUT2 #(
		.INIT('h2)
	) name78 (
		\TM0_pad ,
		\WX10883_reg/NET0131 ,
		_w1587_
	);
	LUT4 #(
		.INIT('h6996)
	) name79 (
		\WX699_reg/NET0131 ,
		\WX763_reg/NET0131 ,
		\WX827_reg/NET0131 ,
		\WX891_reg/NET0131 ,
		_w1588_
	);
	LUT2 #(
		.INIT('h6)
	) name80 (
		_w1587_,
		_w1588_,
		_w1589_
	);
	LUT2 #(
		.INIT('h2)
	) name81 (
		\TM0_pad ,
		\WX10881_reg/NET0131 ,
		_w1590_
	);
	LUT4 #(
		.INIT('h6996)
	) name82 (
		\WX697_reg/NET0131 ,
		\WX761_reg/NET0131 ,
		\WX825_reg/NET0131 ,
		\WX889_reg/NET0131 ,
		_w1591_
	);
	LUT2 #(
		.INIT('h6)
	) name83 (
		_w1590_,
		_w1591_,
		_w1592_
	);
	LUT2 #(
		.INIT('h2)
	) name84 (
		\TM0_pad ,
		\WX10879_reg/NET0131 ,
		_w1593_
	);
	LUT4 #(
		.INIT('h6996)
	) name85 (
		\WX695_reg/NET0131 ,
		\WX759_reg/NET0131 ,
		\WX823_reg/NET0131 ,
		\WX887_reg/NET0131 ,
		_w1594_
	);
	LUT2 #(
		.INIT('h6)
	) name86 (
		_w1593_,
		_w1594_,
		_w1595_
	);
	LUT2 #(
		.INIT('h2)
	) name87 (
		\TM0_pad ,
		\WX10877_reg/NET0131 ,
		_w1596_
	);
	LUT4 #(
		.INIT('h6996)
	) name88 (
		\WX693_reg/NET0131 ,
		\WX757_reg/NET0131 ,
		\WX821_reg/NET0131 ,
		\WX885_reg/NET0131 ,
		_w1597_
	);
	LUT2 #(
		.INIT('h6)
	) name89 (
		_w1596_,
		_w1597_,
		_w1598_
	);
	LUT2 #(
		.INIT('h2)
	) name90 (
		\TM0_pad ,
		\WX10875_reg/NET0131 ,
		_w1599_
	);
	LUT4 #(
		.INIT('h6996)
	) name91 (
		\WX691_reg/NET0131 ,
		\WX755_reg/NET0131 ,
		\WX819_reg/NET0131 ,
		\WX883_reg/NET0131 ,
		_w1600_
	);
	LUT2 #(
		.INIT('h6)
	) name92 (
		_w1599_,
		_w1600_,
		_w1601_
	);
	LUT2 #(
		.INIT('h2)
	) name93 (
		\TM0_pad ,
		\WX10873_reg/NET0131 ,
		_w1602_
	);
	LUT4 #(
		.INIT('h6996)
	) name94 (
		\WX689_reg/NET0131 ,
		\WX753_reg/NET0131 ,
		\WX817_reg/NET0131 ,
		\WX881_reg/NET0131 ,
		_w1603_
	);
	LUT2 #(
		.INIT('h6)
	) name95 (
		_w1602_,
		_w1603_,
		_w1604_
	);
	LUT2 #(
		.INIT('h8)
	) name96 (
		RESET_pad,
		\TM1_pad ,
		_w1605_
	);
	LUT4 #(
		.INIT('ha020)
	) name97 (
		RESET_pad,
		\TM0_pad ,
		\TM1_pad ,
		\WX10861_reg/NET0131 ,
		_w1606_
	);
	LUT3 #(
		.INIT('he0)
	) name98 (
		\TM0_pad ,
		_w1528_,
		_w1606_,
		_w1607_
	);
	LUT2 #(
		.INIT('h9)
	) name99 (
		\WX2098_reg/NET0131 ,
		\WX2162_reg/NET0131 ,
		_w1608_
	);
	LUT2 #(
		.INIT('h9)
	) name100 (
		\WX1970_reg/NET0131 ,
		\WX2034_reg/NET0131 ,
		_w1609_
	);
	LUT4 #(
		.INIT('h0a02)
	) name101 (
		RESET_pad,
		\TM0_pad ,
		\TM1_pad ,
		\_2092__reg/NET0131 ,
		_w1610_
	);
	LUT4 #(
		.INIT('hbe00)
	) name102 (
		\TM0_pad ,
		_w1608_,
		_w1609_,
		_w1610_,
		_w1611_
	);
	LUT2 #(
		.INIT('he)
	) name103 (
		_w1607_,
		_w1611_,
		_w1612_
	);
	LUT3 #(
		.INIT('h96)
	) name104 (
		\WX9766_reg/NET0131 ,
		\WX9830_reg/NET0131 ,
		\WX9894_reg/NET0131 ,
		_w1613_
	);
	LUT2 #(
		.INIT('h9)
	) name105 (
		\TM1_pad ,
		\WX9702_reg/NET0131 ,
		_w1614_
	);
	LUT4 #(
		.INIT('h2772)
	) name106 (
		\TM0_pad ,
		\WX10835_reg/NET0131 ,
		_w1613_,
		_w1614_,
		_w1615_
	);
	LUT3 #(
		.INIT('h96)
	) name107 (
		\WX11059_reg/NET0131 ,
		\WX11123_reg/NET0131 ,
		\WX11187_reg/NET0131 ,
		_w1616_
	);
	LUT2 #(
		.INIT('h9)
	) name108 (
		\TM1_pad ,
		\WX10995_reg/NET0131 ,
		_w1617_
	);
	LUT4 #(
		.INIT('h2772)
	) name109 (
		\TM0_pad ,
		\_2329__reg/NET0131 ,
		_w1616_,
		_w1617_,
		_w1618_
	);
	LUT4 #(
		.INIT('h082a)
	) name110 (
		RESET_pad,
		\TM1_pad ,
		_w1615_,
		_w1618_,
		_w1619_
	);
	LUT4 #(
		.INIT('ha020)
	) name111 (
		RESET_pad,
		\TM0_pad ,
		\TM1_pad ,
		\WX10875_reg/NET0131 ,
		_w1620_
	);
	LUT2 #(
		.INIT('h9)
	) name112 (
		\WX11163_reg/NET0131 ,
		\WX11227_reg/NET0131 ,
		_w1621_
	);
	LUT2 #(
		.INIT('h9)
	) name113 (
		\WX11035_reg/NET0131 ,
		\WX11099_reg/NET0131 ,
		_w1622_
	);
	LUT4 #(
		.INIT('h8cc8)
	) name114 (
		\TM0_pad ,
		_w1620_,
		_w1621_,
		_w1622_,
		_w1623_
	);
	LUT2 #(
		.INIT('h2)
	) name115 (
		\TM0_pad ,
		\_2341__reg/NET0131 ,
		_w1624_
	);
	LUT4 #(
		.INIT('h00c8)
	) name116 (
		\DATA_0_8_pad ,
		RESET_pad,
		\TM0_pad ,
		\TM1_pad ,
		_w1625_
	);
	LUT2 #(
		.INIT('h4)
	) name117 (
		_w1624_,
		_w1625_,
		_w1626_
	);
	LUT2 #(
		.INIT('he)
	) name118 (
		_w1623_,
		_w1626_,
		_w1627_
	);
	LUT4 #(
		.INIT('ha020)
	) name119 (
		RESET_pad,
		\TM0_pad ,
		\TM1_pad ,
		\WX10865_reg/NET0131 ,
		_w1628_
	);
	LUT2 #(
		.INIT('h9)
	) name120 (
		\WX11153_reg/NET0131 ,
		\WX11217_reg/NET0131 ,
		_w1629_
	);
	LUT2 #(
		.INIT('h9)
	) name121 (
		\WX11025_reg/NET0131 ,
		\WX11089_reg/NET0131 ,
		_w1630_
	);
	LUT4 #(
		.INIT('h8cc8)
	) name122 (
		\TM0_pad ,
		_w1628_,
		_w1629_,
		_w1630_,
		_w1631_
	);
	LUT2 #(
		.INIT('h2)
	) name123 (
		\TM0_pad ,
		\_2346__reg/NET0131 ,
		_w1632_
	);
	LUT4 #(
		.INIT('h00c8)
	) name124 (
		\DATA_0_13_pad ,
		RESET_pad,
		\TM0_pad ,
		\TM1_pad ,
		_w1633_
	);
	LUT2 #(
		.INIT('h4)
	) name125 (
		_w1632_,
		_w1633_,
		_w1634_
	);
	LUT2 #(
		.INIT('he)
	) name126 (
		_w1631_,
		_w1634_,
		_w1635_
	);
	LUT4 #(
		.INIT('h2772)
	) name127 (
		\TM0_pad ,
		\WX10831_reg/NET0131 ,
		_w1578_,
		_w1579_,
		_w1636_
	);
	LUT3 #(
		.INIT('h96)
	) name128 (
		\WX2004_reg/NET0131 ,
		\WX2068_reg/NET0131 ,
		\WX2132_reg/NET0131 ,
		_w1637_
	);
	LUT2 #(
		.INIT('h9)
	) name129 (
		\TM1_pad ,
		\WX1940_reg/NET0131 ,
		_w1638_
	);
	LUT4 #(
		.INIT('h2772)
	) name130 (
		\TM0_pad ,
		\_2107__reg/NET0131 ,
		_w1637_,
		_w1638_,
		_w1639_
	);
	LUT4 #(
		.INIT('h082a)
	) name131 (
		RESET_pad,
		\TM1_pad ,
		_w1636_,
		_w1639_,
		_w1640_
	);
	LUT4 #(
		.INIT('h2772)
	) name132 (
		\TM0_pad ,
		\WX10833_reg/NET0131 ,
		_w1572_,
		_w1573_,
		_w1641_
	);
	LUT3 #(
		.INIT('h96)
	) name133 (
		\WX2006_reg/NET0131 ,
		\WX2070_reg/NET0131 ,
		\WX2134_reg/NET0131 ,
		_w1642_
	);
	LUT2 #(
		.INIT('h9)
	) name134 (
		\TM1_pad ,
		\WX1942_reg/NET0131 ,
		_w1643_
	);
	LUT4 #(
		.INIT('h2772)
	) name135 (
		\TM0_pad ,
		\_2106__reg/NET0131 ,
		_w1642_,
		_w1643_,
		_w1644_
	);
	LUT4 #(
		.INIT('h082a)
	) name136 (
		RESET_pad,
		\TM1_pad ,
		_w1641_,
		_w1644_,
		_w1645_
	);
	LUT2 #(
		.INIT('h9)
	) name137 (
		\WX3391_reg/NET0131 ,
		\WX3455_reg/NET0131 ,
		_w1646_
	);
	LUT2 #(
		.INIT('h9)
	) name138 (
		\WX3263_reg/NET0131 ,
		\WX3327_reg/NET0131 ,
		_w1647_
	);
	LUT4 #(
		.INIT('h8cc8)
	) name139 (
		\TM0_pad ,
		_w1606_,
		_w1646_,
		_w1647_,
		_w1648_
	);
	LUT2 #(
		.INIT('h9)
	) name140 (
		\WX4684_reg/NET0131 ,
		\WX4748_reg/NET0131 ,
		_w1649_
	);
	LUT2 #(
		.INIT('h9)
	) name141 (
		\WX4556_reg/NET0131 ,
		\WX4620_reg/NET0131 ,
		_w1650_
	);
	LUT4 #(
		.INIT('h0a02)
	) name142 (
		RESET_pad,
		\TM0_pad ,
		\TM1_pad ,
		\_2156__reg/NET0131 ,
		_w1651_
	);
	LUT4 #(
		.INIT('hbe00)
	) name143 (
		\TM0_pad ,
		_w1649_,
		_w1650_,
		_w1651_,
		_w1652_
	);
	LUT2 #(
		.INIT('he)
	) name144 (
		_w1648_,
		_w1652_,
		_w1653_
	);
	LUT3 #(
		.INIT('h96)
	) name145 (
		\WX3297_reg/NET0131 ,
		\WX3361_reg/NET0131 ,
		\WX3425_reg/NET0131 ,
		_w1654_
	);
	LUT2 #(
		.INIT('h9)
	) name146 (
		\TM1_pad ,
		\WX3233_reg/NET0131 ,
		_w1655_
	);
	LUT4 #(
		.INIT('h2772)
	) name147 (
		\TM0_pad ,
		\_2139__reg/NET0131 ,
		_w1654_,
		_w1655_,
		_w1656_
	);
	LUT4 #(
		.INIT('h2772)
	) name148 (
		\TM0_pad ,
		\WX10831_reg/NET0131 ,
		_w1637_,
		_w1638_,
		_w1657_
	);
	LUT4 #(
		.INIT('h028a)
	) name149 (
		RESET_pad,
		\TM1_pad ,
		_w1656_,
		_w1657_,
		_w1658_
	);
	LUT3 #(
		.INIT('h96)
	) name150 (
		\WX9784_reg/NET0131 ,
		\WX9848_reg/NET0131 ,
		\WX9912_reg/NET0131 ,
		_w1659_
	);
	LUT2 #(
		.INIT('h9)
	) name151 (
		\TM1_pad ,
		\WX9720_reg/NET0131 ,
		_w1660_
	);
	LUT4 #(
		.INIT('h2772)
	) name152 (
		\TM0_pad ,
		\_2288__reg/NET0131 ,
		_w1659_,
		_w1660_,
		_w1661_
	);
	LUT3 #(
		.INIT('h96)
	) name153 (
		\WX8491_reg/NET0131 ,
		\WX8555_reg/NET0131 ,
		\WX8619_reg/NET0131 ,
		_w1662_
	);
	LUT2 #(
		.INIT('h9)
	) name154 (
		\TM1_pad ,
		\WX8427_reg/NET0131 ,
		_w1663_
	);
	LUT4 #(
		.INIT('h2772)
	) name155 (
		\TM0_pad ,
		\WX10853_reg/NET0131 ,
		_w1662_,
		_w1663_,
		_w1664_
	);
	LUT4 #(
		.INIT('h028a)
	) name156 (
		RESET_pad,
		\TM1_pad ,
		_w1661_,
		_w1664_,
		_w1665_
	);
	LUT3 #(
		.INIT('h96)
	) name157 (
		\WX11075_reg/NET0131 ,
		\WX11139_reg/NET0131 ,
		\WX11203_reg/NET0131 ,
		_w1666_
	);
	LUT2 #(
		.INIT('h9)
	) name158 (
		\TM1_pad ,
		\WX11011_reg/NET0131 ,
		_w1667_
	);
	LUT4 #(
		.INIT('h2772)
	) name159 (
		\TM0_pad ,
		\_2321__reg/NET0131 ,
		_w1666_,
		_w1667_,
		_w1668_
	);
	LUT3 #(
		.INIT('h96)
	) name160 (
		\WX9782_reg/NET0131 ,
		\WX9846_reg/NET0131 ,
		\WX9910_reg/NET0131 ,
		_w1669_
	);
	LUT2 #(
		.INIT('h9)
	) name161 (
		\TM1_pad ,
		\WX9718_reg/NET0131 ,
		_w1670_
	);
	LUT4 #(
		.INIT('h2772)
	) name162 (
		\TM0_pad ,
		\WX10851_reg/NET0131 ,
		_w1669_,
		_w1670_,
		_w1671_
	);
	LUT4 #(
		.INIT('h028a)
	) name163 (
		RESET_pad,
		\TM1_pad ,
		_w1668_,
		_w1671_,
		_w1672_
	);
	LUT3 #(
		.INIT('h96)
	) name164 (
		\WX5911_reg/NET0131 ,
		\WX5975_reg/NET0131 ,
		\WX6039_reg/NET0131 ,
		_w1673_
	);
	LUT2 #(
		.INIT('h9)
	) name165 (
		\TM1_pad ,
		\WX5847_reg/NET0131 ,
		_w1674_
	);
	LUT4 #(
		.INIT('h2772)
	) name166 (
		\TM0_pad ,
		\_2189__reg/NET0131 ,
		_w1673_,
		_w1674_,
		_w1675_
	);
	LUT3 #(
		.INIT('h96)
	) name167 (
		\WX4618_reg/NET0131 ,
		\WX4682_reg/NET0131 ,
		\WX4746_reg/NET0131 ,
		_w1676_
	);
	LUT2 #(
		.INIT('h9)
	) name168 (
		\TM1_pad ,
		\WX4554_reg/NET0131 ,
		_w1677_
	);
	LUT4 #(
		.INIT('h2772)
	) name169 (
		\TM0_pad ,
		\WX10859_reg/NET0131 ,
		_w1676_,
		_w1677_,
		_w1678_
	);
	LUT4 #(
		.INIT('h028a)
	) name170 (
		RESET_pad,
		\TM1_pad ,
		_w1675_,
		_w1678_,
		_w1679_
	);
	LUT3 #(
		.INIT('h96)
	) name171 (
		\WX7202_reg/NET0131 ,
		\WX7266_reg/NET0131 ,
		\WX7330_reg/NET0131 ,
		_w1680_
	);
	LUT2 #(
		.INIT('h9)
	) name172 (
		\TM1_pad ,
		\WX7138_reg/NET0131 ,
		_w1681_
	);
	LUT4 #(
		.INIT('h2772)
	) name173 (
		\TM0_pad ,
		\_2222__reg/NET0131 ,
		_w1680_,
		_w1681_,
		_w1682_
	);
	LUT3 #(
		.INIT('h96)
	) name174 (
		\WX5909_reg/NET0131 ,
		\WX5973_reg/NET0131 ,
		\WX6037_reg/NET0131 ,
		_w1683_
	);
	LUT2 #(
		.INIT('h9)
	) name175 (
		\TM1_pad ,
		\WX5845_reg/NET0131 ,
		_w1684_
	);
	LUT4 #(
		.INIT('h2772)
	) name176 (
		\TM0_pad ,
		\WX10857_reg/NET0131 ,
		_w1683_,
		_w1684_,
		_w1685_
	);
	LUT4 #(
		.INIT('h028a)
	) name177 (
		RESET_pad,
		\TM1_pad ,
		_w1682_,
		_w1685_,
		_w1686_
	);
	LUT3 #(
		.INIT('h96)
	) name178 (
		\WX8493_reg/NET0131 ,
		\WX8557_reg/NET0131 ,
		\WX8621_reg/NET0131 ,
		_w1687_
	);
	LUT2 #(
		.INIT('h9)
	) name179 (
		\TM1_pad ,
		\WX8429_reg/NET0131 ,
		_w1688_
	);
	LUT4 #(
		.INIT('h2772)
	) name180 (
		\TM0_pad ,
		\_2255__reg/NET0131 ,
		_w1687_,
		_w1688_,
		_w1689_
	);
	LUT3 #(
		.INIT('h96)
	) name181 (
		\WX7200_reg/NET0131 ,
		\WX7264_reg/NET0131 ,
		\WX7328_reg/NET0131 ,
		_w1690_
	);
	LUT2 #(
		.INIT('h9)
	) name182 (
		\TM1_pad ,
		\WX7136_reg/NET0131 ,
		_w1691_
	);
	LUT4 #(
		.INIT('h2772)
	) name183 (
		\TM0_pad ,
		\WX10855_reg/NET0131 ,
		_w1690_,
		_w1691_,
		_w1692_
	);
	LUT4 #(
		.INIT('h028a)
	) name184 (
		RESET_pad,
		\TM1_pad ,
		_w1689_,
		_w1692_,
		_w1693_
	);
	LUT4 #(
		.INIT('h2772)
	) name185 (
		\TM0_pad ,
		\WX10835_reg/NET0131 ,
		_w1569_,
		_w1570_,
		_w1694_
	);
	LUT3 #(
		.INIT('h96)
	) name186 (
		\WX2008_reg/NET0131 ,
		\WX2072_reg/NET0131 ,
		\WX2136_reg/NET0131 ,
		_w1695_
	);
	LUT2 #(
		.INIT('h9)
	) name187 (
		\TM1_pad ,
		\WX1944_reg/NET0131 ,
		_w1696_
	);
	LUT4 #(
		.INIT('h2772)
	) name188 (
		\TM0_pad ,
		\_2105__reg/NET0131 ,
		_w1695_,
		_w1696_,
		_w1697_
	);
	LUT4 #(
		.INIT('h082a)
	) name189 (
		RESET_pad,
		\TM1_pad ,
		_w1694_,
		_w1697_,
		_w1698_
	);
	LUT3 #(
		.INIT('h96)
	) name190 (
		\WX11055_reg/NET0131 ,
		\WX11119_reg/NET0131 ,
		\WX11183_reg/NET0131 ,
		_w1699_
	);
	LUT2 #(
		.INIT('h9)
	) name191 (
		\TM1_pad ,
		\WX10991_reg/NET0131 ,
		_w1700_
	);
	LUT4 #(
		.INIT('h2772)
	) name192 (
		\TM0_pad ,
		\WX10831_reg/NET0131 ,
		_w1699_,
		_w1700_,
		_w1701_
	);
	LUT2 #(
		.INIT('h2)
	) name193 (
		\TM0_pad ,
		\_2363__reg/NET0131 ,
		_w1702_
	);
	LUT4 #(
		.INIT('h00c8)
	) name194 (
		\DATA_0_30_pad ,
		RESET_pad,
		\TM0_pad ,
		\TM1_pad ,
		_w1703_
	);
	LUT2 #(
		.INIT('h4)
	) name195 (
		_w1702_,
		_w1703_,
		_w1704_
	);
	LUT3 #(
		.INIT('hf2)
	) name196 (
		_w1605_,
		_w1701_,
		_w1704_,
		_w1705_
	);
	LUT4 #(
		.INIT('ha020)
	) name197 (
		RESET_pad,
		\TM0_pad ,
		\TM1_pad ,
		\WX10863_reg/NET0131 ,
		_w1706_
	);
	LUT2 #(
		.INIT('h9)
	) name198 (
		\WX3393_reg/NET0131 ,
		\WX3457_reg/NET0131 ,
		_w1707_
	);
	LUT2 #(
		.INIT('h9)
	) name199 (
		\WX3265_reg/NET0131 ,
		\WX3329_reg/NET0131 ,
		_w1708_
	);
	LUT4 #(
		.INIT('h8cc8)
	) name200 (
		\TM0_pad ,
		_w1706_,
		_w1707_,
		_w1708_,
		_w1709_
	);
	LUT2 #(
		.INIT('h9)
	) name201 (
		\WX4686_reg/NET0131 ,
		\WX4750_reg/NET0131 ,
		_w1710_
	);
	LUT2 #(
		.INIT('h9)
	) name202 (
		\WX4558_reg/NET0131 ,
		\WX4622_reg/NET0131 ,
		_w1711_
	);
	LUT4 #(
		.INIT('h0a02)
	) name203 (
		RESET_pad,
		\TM0_pad ,
		\TM1_pad ,
		\_2155__reg/NET0131 ,
		_w1712_
	);
	LUT4 #(
		.INIT('hbe00)
	) name204 (
		\TM0_pad ,
		_w1710_,
		_w1711_,
		_w1712_,
		_w1713_
	);
	LUT2 #(
		.INIT('he)
	) name205 (
		_w1709_,
		_w1713_,
		_w1714_
	);
	LUT3 #(
		.INIT('h96)
	) name206 (
		\WX9786_reg/NET0131 ,
		\WX9850_reg/NET0131 ,
		\WX9914_reg/NET0131 ,
		_w1715_
	);
	LUT2 #(
		.INIT('h9)
	) name207 (
		\TM1_pad ,
		\WX9722_reg/NET0131 ,
		_w1716_
	);
	LUT4 #(
		.INIT('h2772)
	) name208 (
		\TM0_pad ,
		\_2287__reg/NET0131 ,
		_w1715_,
		_w1716_,
		_w1717_
	);
	LUT4 #(
		.INIT('h2772)
	) name209 (
		\TM0_pad ,
		\WX10855_reg/NET0131 ,
		_w1687_,
		_w1688_,
		_w1718_
	);
	LUT4 #(
		.INIT('h028a)
	) name210 (
		RESET_pad,
		\TM1_pad ,
		_w1717_,
		_w1718_,
		_w1719_
	);
	LUT3 #(
		.INIT('h96)
	) name211 (
		\WX3299_reg/NET0131 ,
		\WX3363_reg/NET0131 ,
		\WX3427_reg/NET0131 ,
		_w1720_
	);
	LUT2 #(
		.INIT('h9)
	) name212 (
		\TM1_pad ,
		\WX3235_reg/NET0131 ,
		_w1721_
	);
	LUT4 #(
		.INIT('h2772)
	) name213 (
		\TM0_pad ,
		\_2138__reg/NET0131 ,
		_w1720_,
		_w1721_,
		_w1722_
	);
	LUT4 #(
		.INIT('h2772)
	) name214 (
		\TM0_pad ,
		\WX10833_reg/NET0131 ,
		_w1642_,
		_w1643_,
		_w1723_
	);
	LUT4 #(
		.INIT('h028a)
	) name215 (
		RESET_pad,
		\TM1_pad ,
		_w1722_,
		_w1723_,
		_w1724_
	);
	LUT3 #(
		.INIT('h96)
	) name216 (
		\WX11077_reg/NET0131 ,
		\WX11141_reg/NET0131 ,
		\WX11205_reg/NET0131 ,
		_w1725_
	);
	LUT2 #(
		.INIT('h9)
	) name217 (
		\TM1_pad ,
		\WX11013_reg/NET0131 ,
		_w1726_
	);
	LUT4 #(
		.INIT('h2772)
	) name218 (
		\TM0_pad ,
		\_2320__reg/NET0131 ,
		_w1725_,
		_w1726_,
		_w1727_
	);
	LUT4 #(
		.INIT('h2772)
	) name219 (
		\TM0_pad ,
		\WX10853_reg/NET0131 ,
		_w1659_,
		_w1660_,
		_w1728_
	);
	LUT4 #(
		.INIT('h028a)
	) name220 (
		RESET_pad,
		\TM1_pad ,
		_w1727_,
		_w1728_,
		_w1729_
	);
	LUT4 #(
		.INIT('h8cc8)
	) name221 (
		\TM0_pad ,
		_w1606_,
		_w1649_,
		_w1650_,
		_w1730_
	);
	LUT2 #(
		.INIT('h9)
	) name222 (
		\WX5977_reg/NET0131 ,
		\WX6041_reg/NET0131 ,
		_w1731_
	);
	LUT2 #(
		.INIT('h9)
	) name223 (
		\WX5849_reg/NET0131 ,
		\WX5913_reg/NET0131 ,
		_w1732_
	);
	LUT4 #(
		.INIT('h0a02)
	) name224 (
		RESET_pad,
		\TM0_pad ,
		\TM1_pad ,
		\_2188__reg/NET0131 ,
		_w1733_
	);
	LUT4 #(
		.INIT('hbe00)
	) name225 (
		\TM0_pad ,
		_w1731_,
		_w1732_,
		_w1733_,
		_w1734_
	);
	LUT2 #(
		.INIT('he)
	) name226 (
		_w1730_,
		_w1734_,
		_w1735_
	);
	LUT3 #(
		.INIT('h96)
	) name227 (
		\WX7204_reg/NET0131 ,
		\WX7268_reg/NET0131 ,
		\WX7332_reg/NET0131 ,
		_w1736_
	);
	LUT2 #(
		.INIT('h9)
	) name228 (
		\TM1_pad ,
		\WX7140_reg/NET0131 ,
		_w1737_
	);
	LUT4 #(
		.INIT('h2772)
	) name229 (
		\TM0_pad ,
		\_2221__reg/NET0131 ,
		_w1736_,
		_w1737_,
		_w1738_
	);
	LUT4 #(
		.INIT('h2772)
	) name230 (
		\TM0_pad ,
		\WX10859_reg/NET0131 ,
		_w1673_,
		_w1674_,
		_w1739_
	);
	LUT4 #(
		.INIT('h028a)
	) name231 (
		RESET_pad,
		\TM1_pad ,
		_w1738_,
		_w1739_,
		_w1740_
	);
	LUT3 #(
		.INIT('h96)
	) name232 (
		\WX8495_reg/NET0131 ,
		\WX8559_reg/NET0131 ,
		\WX8623_reg/NET0131 ,
		_w1741_
	);
	LUT2 #(
		.INIT('h9)
	) name233 (
		\TM1_pad ,
		\WX8431_reg/NET0131 ,
		_w1742_
	);
	LUT4 #(
		.INIT('h2772)
	) name234 (
		\TM0_pad ,
		\_2254__reg/NET0131 ,
		_w1741_,
		_w1742_,
		_w1743_
	);
	LUT4 #(
		.INIT('h2772)
	) name235 (
		\TM0_pad ,
		\WX10857_reg/NET0131 ,
		_w1680_,
		_w1681_,
		_w1744_
	);
	LUT4 #(
		.INIT('h028a)
	) name236 (
		RESET_pad,
		\TM1_pad ,
		_w1743_,
		_w1744_,
		_w1745_
	);
	LUT4 #(
		.INIT('h2772)
	) name237 (
		\TM0_pad ,
		\WX10837_reg/NET0131 ,
		_w1566_,
		_w1567_,
		_w1746_
	);
	LUT3 #(
		.INIT('h96)
	) name238 (
		\WX2010_reg/NET0131 ,
		\WX2074_reg/NET0131 ,
		\WX2138_reg/NET0131 ,
		_w1747_
	);
	LUT2 #(
		.INIT('h9)
	) name239 (
		\TM1_pad ,
		\WX1946_reg/NET0131 ,
		_w1748_
	);
	LUT4 #(
		.INIT('h2772)
	) name240 (
		\TM0_pad ,
		\_2104__reg/NET0131 ,
		_w1747_,
		_w1748_,
		_w1749_
	);
	LUT4 #(
		.INIT('h082a)
	) name241 (
		RESET_pad,
		\TM1_pad ,
		_w1746_,
		_w1749_,
		_w1750_
	);
	LUT3 #(
		.INIT('h96)
	) name242 (
		\WX11057_reg/NET0131 ,
		\WX11121_reg/NET0131 ,
		\WX11185_reg/NET0131 ,
		_w1751_
	);
	LUT2 #(
		.INIT('h9)
	) name243 (
		\TM1_pad ,
		\WX10993_reg/NET0131 ,
		_w1752_
	);
	LUT4 #(
		.INIT('h2772)
	) name244 (
		\TM0_pad ,
		\WX10833_reg/NET0131 ,
		_w1751_,
		_w1752_,
		_w1753_
	);
	LUT2 #(
		.INIT('h2)
	) name245 (
		\TM0_pad ,
		\_2362__reg/NET0131 ,
		_w1754_
	);
	LUT4 #(
		.INIT('h00c8)
	) name246 (
		\DATA_0_29_pad ,
		RESET_pad,
		\TM0_pad ,
		\TM1_pad ,
		_w1755_
	);
	LUT2 #(
		.INIT('h4)
	) name247 (
		_w1754_,
		_w1755_,
		_w1756_
	);
	LUT3 #(
		.INIT('hf2)
	) name248 (
		_w1605_,
		_w1753_,
		_w1756_,
		_w1757_
	);
	LUT2 #(
		.INIT('h8)
	) name249 (
		RESET_pad,
		\WX10831_reg/NET0131 ,
		_w1758_
	);
	LUT2 #(
		.INIT('h9)
	) name250 (
		\WX3395_reg/NET0131 ,
		\WX3459_reg/NET0131 ,
		_w1759_
	);
	LUT2 #(
		.INIT('h9)
	) name251 (
		\WX3267_reg/NET0131 ,
		\WX3331_reg/NET0131 ,
		_w1760_
	);
	LUT4 #(
		.INIT('h8cc8)
	) name252 (
		\TM0_pad ,
		_w1628_,
		_w1759_,
		_w1760_,
		_w1761_
	);
	LUT2 #(
		.INIT('h9)
	) name253 (
		\WX4688_reg/NET0131 ,
		\WX4752_reg/NET0131 ,
		_w1762_
	);
	LUT2 #(
		.INIT('h9)
	) name254 (
		\WX4560_reg/NET0131 ,
		\WX4624_reg/NET0131 ,
		_w1763_
	);
	LUT4 #(
		.INIT('h0a02)
	) name255 (
		RESET_pad,
		\TM0_pad ,
		\TM1_pad ,
		\_2154__reg/NET0131 ,
		_w1764_
	);
	LUT4 #(
		.INIT('hbe00)
	) name256 (
		\TM0_pad ,
		_w1762_,
		_w1763_,
		_w1764_,
		_w1765_
	);
	LUT2 #(
		.INIT('he)
	) name257 (
		_w1761_,
		_w1765_,
		_w1766_
	);
	LUT3 #(
		.INIT('h96)
	) name258 (
		\WX9788_reg/NET0131 ,
		\WX9852_reg/NET0131 ,
		\WX9916_reg/NET0131 ,
		_w1767_
	);
	LUT2 #(
		.INIT('h9)
	) name259 (
		\TM1_pad ,
		\WX9724_reg/NET0131 ,
		_w1768_
	);
	LUT4 #(
		.INIT('h2772)
	) name260 (
		\TM0_pad ,
		\_2286__reg/NET0131 ,
		_w1767_,
		_w1768_,
		_w1769_
	);
	LUT4 #(
		.INIT('h2772)
	) name261 (
		\TM0_pad ,
		\WX10857_reg/NET0131 ,
		_w1741_,
		_w1742_,
		_w1770_
	);
	LUT4 #(
		.INIT('h028a)
	) name262 (
		RESET_pad,
		\TM1_pad ,
		_w1769_,
		_w1770_,
		_w1771_
	);
	LUT3 #(
		.INIT('h96)
	) name263 (
		\WX3301_reg/NET0131 ,
		\WX3365_reg/NET0131 ,
		\WX3429_reg/NET0131 ,
		_w1772_
	);
	LUT2 #(
		.INIT('h9)
	) name264 (
		\TM1_pad ,
		\WX3237_reg/NET0131 ,
		_w1773_
	);
	LUT4 #(
		.INIT('h2772)
	) name265 (
		\TM0_pad ,
		\_2137__reg/NET0131 ,
		_w1772_,
		_w1773_,
		_w1774_
	);
	LUT4 #(
		.INIT('h2772)
	) name266 (
		\TM0_pad ,
		\WX10835_reg/NET0131 ,
		_w1695_,
		_w1696_,
		_w1775_
	);
	LUT4 #(
		.INIT('h028a)
	) name267 (
		RESET_pad,
		\TM1_pad ,
		_w1774_,
		_w1775_,
		_w1776_
	);
	LUT3 #(
		.INIT('h96)
	) name268 (
		\WX11079_reg/NET0131 ,
		\WX11143_reg/NET0131 ,
		\WX11207_reg/NET0131 ,
		_w1777_
	);
	LUT2 #(
		.INIT('h9)
	) name269 (
		\TM1_pad ,
		\WX11015_reg/NET0131 ,
		_w1778_
	);
	LUT4 #(
		.INIT('h2772)
	) name270 (
		\TM0_pad ,
		\_2319__reg/NET0131 ,
		_w1777_,
		_w1778_,
		_w1779_
	);
	LUT4 #(
		.INIT('h2772)
	) name271 (
		\TM0_pad ,
		\WX10855_reg/NET0131 ,
		_w1715_,
		_w1716_,
		_w1780_
	);
	LUT4 #(
		.INIT('h028a)
	) name272 (
		RESET_pad,
		\TM1_pad ,
		_w1779_,
		_w1780_,
		_w1781_
	);
	LUT4 #(
		.INIT('h8cc8)
	) name273 (
		\TM0_pad ,
		_w1706_,
		_w1710_,
		_w1711_,
		_w1782_
	);
	LUT2 #(
		.INIT('h9)
	) name274 (
		\WX5979_reg/NET0131 ,
		\WX6043_reg/NET0131 ,
		_w1783_
	);
	LUT2 #(
		.INIT('h9)
	) name275 (
		\WX5851_reg/NET0131 ,
		\WX5915_reg/NET0131 ,
		_w1784_
	);
	LUT4 #(
		.INIT('h0a02)
	) name276 (
		RESET_pad,
		\TM0_pad ,
		\TM1_pad ,
		\_2187__reg/NET0131 ,
		_w1785_
	);
	LUT4 #(
		.INIT('hbe00)
	) name277 (
		\TM0_pad ,
		_w1783_,
		_w1784_,
		_w1785_,
		_w1786_
	);
	LUT2 #(
		.INIT('he)
	) name278 (
		_w1782_,
		_w1786_,
		_w1787_
	);
	LUT4 #(
		.INIT('h8cc8)
	) name279 (
		\TM0_pad ,
		_w1606_,
		_w1731_,
		_w1732_,
		_w1788_
	);
	LUT2 #(
		.INIT('h9)
	) name280 (
		\WX7270_reg/NET0131 ,
		\WX7334_reg/NET0131 ,
		_w1789_
	);
	LUT2 #(
		.INIT('h9)
	) name281 (
		\WX7142_reg/NET0131 ,
		\WX7206_reg/NET0131 ,
		_w1790_
	);
	LUT4 #(
		.INIT('h0a02)
	) name282 (
		RESET_pad,
		\TM0_pad ,
		\TM1_pad ,
		\_2220__reg/NET0131 ,
		_w1791_
	);
	LUT4 #(
		.INIT('hbe00)
	) name283 (
		\TM0_pad ,
		_w1789_,
		_w1790_,
		_w1791_,
		_w1792_
	);
	LUT2 #(
		.INIT('he)
	) name284 (
		_w1788_,
		_w1792_,
		_w1793_
	);
	LUT3 #(
		.INIT('h96)
	) name285 (
		\WX8497_reg/NET0131 ,
		\WX8561_reg/NET0131 ,
		\WX8625_reg/NET0131 ,
		_w1794_
	);
	LUT2 #(
		.INIT('h9)
	) name286 (
		\TM1_pad ,
		\WX8433_reg/NET0131 ,
		_w1795_
	);
	LUT4 #(
		.INIT('h2772)
	) name287 (
		\TM0_pad ,
		\_2253__reg/NET0131 ,
		_w1794_,
		_w1795_,
		_w1796_
	);
	LUT4 #(
		.INIT('h2772)
	) name288 (
		\TM0_pad ,
		\WX10859_reg/NET0131 ,
		_w1736_,
		_w1737_,
		_w1797_
	);
	LUT4 #(
		.INIT('h028a)
	) name289 (
		RESET_pad,
		\TM1_pad ,
		_w1796_,
		_w1797_,
		_w1798_
	);
	LUT4 #(
		.INIT('h2772)
	) name290 (
		\TM0_pad ,
		\WX10839_reg/NET0131 ,
		_w1563_,
		_w1564_,
		_w1799_
	);
	LUT3 #(
		.INIT('h96)
	) name291 (
		\WX2012_reg/NET0131 ,
		\WX2076_reg/NET0131 ,
		\WX2140_reg/NET0131 ,
		_w1800_
	);
	LUT2 #(
		.INIT('h9)
	) name292 (
		\TM1_pad ,
		\WX1948_reg/NET0131 ,
		_w1801_
	);
	LUT4 #(
		.INIT('h2772)
	) name293 (
		\TM0_pad ,
		\_2103__reg/NET0131 ,
		_w1800_,
		_w1801_,
		_w1802_
	);
	LUT4 #(
		.INIT('h082a)
	) name294 (
		RESET_pad,
		\TM1_pad ,
		_w1799_,
		_w1802_,
		_w1803_
	);
	LUT4 #(
		.INIT('h2772)
	) name295 (
		\TM0_pad ,
		\WX10835_reg/NET0131 ,
		_w1616_,
		_w1617_,
		_w1804_
	);
	LUT2 #(
		.INIT('h2)
	) name296 (
		\TM0_pad ,
		\_2361__reg/NET0131 ,
		_w1805_
	);
	LUT4 #(
		.INIT('h00c8)
	) name297 (
		\DATA_0_28_pad ,
		RESET_pad,
		\TM0_pad ,
		\TM1_pad ,
		_w1806_
	);
	LUT2 #(
		.INIT('h4)
	) name298 (
		_w1805_,
		_w1806_,
		_w1807_
	);
	LUT3 #(
		.INIT('hf2)
	) name299 (
		_w1605_,
		_w1804_,
		_w1807_,
		_w1808_
	);
	LUT2 #(
		.INIT('h8)
	) name300 (
		RESET_pad,
		\WX10833_reg/NET0131 ,
		_w1809_
	);
	LUT4 #(
		.INIT('ha020)
	) name301 (
		RESET_pad,
		\TM0_pad ,
		\TM1_pad ,
		\WX10867_reg/NET0131 ,
		_w1810_
	);
	LUT2 #(
		.INIT('h9)
	) name302 (
		\WX3397_reg/NET0131 ,
		\WX3461_reg/NET0131 ,
		_w1811_
	);
	LUT2 #(
		.INIT('h9)
	) name303 (
		\WX3269_reg/NET0131 ,
		\WX3333_reg/NET0131 ,
		_w1812_
	);
	LUT4 #(
		.INIT('h8cc8)
	) name304 (
		\TM0_pad ,
		_w1810_,
		_w1811_,
		_w1812_,
		_w1813_
	);
	LUT2 #(
		.INIT('h9)
	) name305 (
		\WX4690_reg/NET0131 ,
		\WX4754_reg/NET0131 ,
		_w1814_
	);
	LUT2 #(
		.INIT('h9)
	) name306 (
		\WX4562_reg/NET0131 ,
		\WX4626_reg/NET0131 ,
		_w1815_
	);
	LUT4 #(
		.INIT('h0a02)
	) name307 (
		RESET_pad,
		\TM0_pad ,
		\TM1_pad ,
		\_2153__reg/NET0131 ,
		_w1816_
	);
	LUT4 #(
		.INIT('hbe00)
	) name308 (
		\TM0_pad ,
		_w1814_,
		_w1815_,
		_w1816_,
		_w1817_
	);
	LUT2 #(
		.INIT('he)
	) name309 (
		_w1813_,
		_w1817_,
		_w1818_
	);
	LUT3 #(
		.INIT('h96)
	) name310 (
		\WX9790_reg/NET0131 ,
		\WX9854_reg/NET0131 ,
		\WX9918_reg/NET0131 ,
		_w1819_
	);
	LUT2 #(
		.INIT('h9)
	) name311 (
		\TM1_pad ,
		\WX9726_reg/NET0131 ,
		_w1820_
	);
	LUT4 #(
		.INIT('h2772)
	) name312 (
		\TM0_pad ,
		\_2285__reg/NET0131 ,
		_w1819_,
		_w1820_,
		_w1821_
	);
	LUT4 #(
		.INIT('h2772)
	) name313 (
		\TM0_pad ,
		\WX10859_reg/NET0131 ,
		_w1794_,
		_w1795_,
		_w1822_
	);
	LUT4 #(
		.INIT('h028a)
	) name314 (
		RESET_pad,
		\TM1_pad ,
		_w1821_,
		_w1822_,
		_w1823_
	);
	LUT3 #(
		.INIT('h96)
	) name315 (
		\WX3303_reg/NET0131 ,
		\WX3367_reg/NET0131 ,
		\WX3431_reg/NET0131 ,
		_w1824_
	);
	LUT2 #(
		.INIT('h9)
	) name316 (
		\TM1_pad ,
		\WX3239_reg/NET0131 ,
		_w1825_
	);
	LUT4 #(
		.INIT('h2772)
	) name317 (
		\TM0_pad ,
		\_2136__reg/NET0131 ,
		_w1824_,
		_w1825_,
		_w1826_
	);
	LUT4 #(
		.INIT('h2772)
	) name318 (
		\TM0_pad ,
		\WX10837_reg/NET0131 ,
		_w1747_,
		_w1748_,
		_w1827_
	);
	LUT4 #(
		.INIT('h028a)
	) name319 (
		RESET_pad,
		\TM1_pad ,
		_w1826_,
		_w1827_,
		_w1828_
	);
	LUT3 #(
		.INIT('h96)
	) name320 (
		\WX11081_reg/NET0131 ,
		\WX11145_reg/NET0131 ,
		\WX11209_reg/NET0131 ,
		_w1829_
	);
	LUT2 #(
		.INIT('h9)
	) name321 (
		\TM1_pad ,
		\WX11017_reg/NET0131 ,
		_w1830_
	);
	LUT4 #(
		.INIT('h2772)
	) name322 (
		\TM0_pad ,
		\_2318__reg/NET0131 ,
		_w1829_,
		_w1830_,
		_w1831_
	);
	LUT4 #(
		.INIT('h2772)
	) name323 (
		\TM0_pad ,
		\WX10857_reg/NET0131 ,
		_w1767_,
		_w1768_,
		_w1832_
	);
	LUT4 #(
		.INIT('h028a)
	) name324 (
		RESET_pad,
		\TM1_pad ,
		_w1831_,
		_w1832_,
		_w1833_
	);
	LUT4 #(
		.INIT('h8cc8)
	) name325 (
		\TM0_pad ,
		_w1628_,
		_w1762_,
		_w1763_,
		_w1834_
	);
	LUT2 #(
		.INIT('h9)
	) name326 (
		\WX5981_reg/NET0131 ,
		\WX6045_reg/NET0131 ,
		_w1835_
	);
	LUT2 #(
		.INIT('h9)
	) name327 (
		\WX5853_reg/NET0131 ,
		\WX5917_reg/NET0131 ,
		_w1836_
	);
	LUT4 #(
		.INIT('h0a02)
	) name328 (
		RESET_pad,
		\TM0_pad ,
		\TM1_pad ,
		\_2186__reg/NET0131 ,
		_w1837_
	);
	LUT4 #(
		.INIT('hbe00)
	) name329 (
		\TM0_pad ,
		_w1835_,
		_w1836_,
		_w1837_,
		_w1838_
	);
	LUT2 #(
		.INIT('he)
	) name330 (
		_w1834_,
		_w1838_,
		_w1839_
	);
	LUT4 #(
		.INIT('h8cc8)
	) name331 (
		\TM0_pad ,
		_w1706_,
		_w1783_,
		_w1784_,
		_w1840_
	);
	LUT2 #(
		.INIT('h9)
	) name332 (
		\WX7272_reg/NET0131 ,
		\WX7336_reg/NET0131 ,
		_w1841_
	);
	LUT2 #(
		.INIT('h9)
	) name333 (
		\WX7144_reg/NET0131 ,
		\WX7208_reg/NET0131 ,
		_w1842_
	);
	LUT4 #(
		.INIT('h0a02)
	) name334 (
		RESET_pad,
		\TM0_pad ,
		\TM1_pad ,
		\_2219__reg/NET0131 ,
		_w1843_
	);
	LUT4 #(
		.INIT('hbe00)
	) name335 (
		\TM0_pad ,
		_w1841_,
		_w1842_,
		_w1843_,
		_w1844_
	);
	LUT2 #(
		.INIT('he)
	) name336 (
		_w1840_,
		_w1844_,
		_w1845_
	);
	LUT4 #(
		.INIT('h8cc8)
	) name337 (
		\TM0_pad ,
		_w1606_,
		_w1789_,
		_w1790_,
		_w1846_
	);
	LUT2 #(
		.INIT('h9)
	) name338 (
		\WX8563_reg/NET0131 ,
		\WX8627_reg/NET0131 ,
		_w1847_
	);
	LUT2 #(
		.INIT('h9)
	) name339 (
		\WX8435_reg/NET0131 ,
		\WX8499_reg/NET0131 ,
		_w1848_
	);
	LUT4 #(
		.INIT('h0a02)
	) name340 (
		RESET_pad,
		\TM0_pad ,
		\TM1_pad ,
		\_2252__reg/NET0131 ,
		_w1849_
	);
	LUT4 #(
		.INIT('hbe00)
	) name341 (
		\TM0_pad ,
		_w1847_,
		_w1848_,
		_w1849_,
		_w1850_
	);
	LUT2 #(
		.INIT('he)
	) name342 (
		_w1846_,
		_w1850_,
		_w1851_
	);
	LUT4 #(
		.INIT('h2772)
	) name343 (
		\TM0_pad ,
		\WX10841_reg/NET0131 ,
		_w1560_,
		_w1561_,
		_w1852_
	);
	LUT3 #(
		.INIT('h96)
	) name344 (
		\WX2014_reg/NET0131 ,
		\WX2078_reg/NET0131 ,
		\WX2142_reg/NET0131 ,
		_w1853_
	);
	LUT2 #(
		.INIT('h9)
	) name345 (
		\TM1_pad ,
		\WX1950_reg/NET0131 ,
		_w1854_
	);
	LUT4 #(
		.INIT('h2772)
	) name346 (
		\TM0_pad ,
		\_2102__reg/NET0131 ,
		_w1853_,
		_w1854_,
		_w1855_
	);
	LUT4 #(
		.INIT('h082a)
	) name347 (
		RESET_pad,
		\TM1_pad ,
		_w1852_,
		_w1855_,
		_w1856_
	);
	LUT3 #(
		.INIT('h96)
	) name348 (
		\WX11061_reg/NET0131 ,
		\WX11125_reg/NET0131 ,
		\WX11189_reg/NET0131 ,
		_w1857_
	);
	LUT2 #(
		.INIT('h9)
	) name349 (
		\TM1_pad ,
		\WX10997_reg/NET0131 ,
		_w1858_
	);
	LUT4 #(
		.INIT('h2772)
	) name350 (
		\TM0_pad ,
		\WX10837_reg/NET0131 ,
		_w1857_,
		_w1858_,
		_w1859_
	);
	LUT2 #(
		.INIT('h2)
	) name351 (
		\TM0_pad ,
		\_2360__reg/NET0131 ,
		_w1860_
	);
	LUT4 #(
		.INIT('h00c8)
	) name352 (
		\DATA_0_27_pad ,
		RESET_pad,
		\TM0_pad ,
		\TM1_pad ,
		_w1861_
	);
	LUT2 #(
		.INIT('h4)
	) name353 (
		_w1860_,
		_w1861_,
		_w1862_
	);
	LUT3 #(
		.INIT('hf2)
	) name354 (
		_w1605_,
		_w1859_,
		_w1862_,
		_w1863_
	);
	LUT2 #(
		.INIT('h8)
	) name355 (
		RESET_pad,
		\WX10835_reg/NET0131 ,
		_w1864_
	);
	LUT4 #(
		.INIT('ha020)
	) name356 (
		RESET_pad,
		\TM0_pad ,
		\TM1_pad ,
		\WX10869_reg/NET0131 ,
		_w1865_
	);
	LUT2 #(
		.INIT('h9)
	) name357 (
		\WX3399_reg/NET0131 ,
		\WX3463_reg/NET0131 ,
		_w1866_
	);
	LUT2 #(
		.INIT('h9)
	) name358 (
		\WX3271_reg/NET0131 ,
		\WX3335_reg/NET0131 ,
		_w1867_
	);
	LUT4 #(
		.INIT('h8cc8)
	) name359 (
		\TM0_pad ,
		_w1865_,
		_w1866_,
		_w1867_,
		_w1868_
	);
	LUT2 #(
		.INIT('h9)
	) name360 (
		\WX4692_reg/NET0131 ,
		\WX4756_reg/NET0131 ,
		_w1869_
	);
	LUT2 #(
		.INIT('h9)
	) name361 (
		\WX4564_reg/NET0131 ,
		\WX4628_reg/NET0131 ,
		_w1870_
	);
	LUT4 #(
		.INIT('h0a02)
	) name362 (
		RESET_pad,
		\TM0_pad ,
		\TM1_pad ,
		\_2152__reg/NET0131 ,
		_w1871_
	);
	LUT4 #(
		.INIT('hbe00)
	) name363 (
		\TM0_pad ,
		_w1869_,
		_w1870_,
		_w1871_,
		_w1872_
	);
	LUT2 #(
		.INIT('he)
	) name364 (
		_w1868_,
		_w1872_,
		_w1873_
	);
	LUT4 #(
		.INIT('h8cc8)
	) name365 (
		\TM0_pad ,
		_w1606_,
		_w1847_,
		_w1848_,
		_w1874_
	);
	LUT2 #(
		.INIT('h9)
	) name366 (
		\WX9856_reg/NET0131 ,
		\WX9920_reg/NET0131 ,
		_w1875_
	);
	LUT2 #(
		.INIT('h9)
	) name367 (
		\WX9728_reg/NET0131 ,
		\WX9792_reg/NET0131 ,
		_w1876_
	);
	LUT4 #(
		.INIT('h0a02)
	) name368 (
		RESET_pad,
		\TM0_pad ,
		\TM1_pad ,
		\_2284__reg/NET0131 ,
		_w1877_
	);
	LUT4 #(
		.INIT('hbe00)
	) name369 (
		\TM0_pad ,
		_w1875_,
		_w1876_,
		_w1877_,
		_w1878_
	);
	LUT2 #(
		.INIT('he)
	) name370 (
		_w1874_,
		_w1878_,
		_w1879_
	);
	LUT3 #(
		.INIT('h96)
	) name371 (
		\WX3305_reg/NET0131 ,
		\WX3369_reg/NET0131 ,
		\WX3433_reg/NET0131 ,
		_w1880_
	);
	LUT2 #(
		.INIT('h9)
	) name372 (
		\TM1_pad ,
		\WX3241_reg/NET0131 ,
		_w1881_
	);
	LUT4 #(
		.INIT('h2772)
	) name373 (
		\TM0_pad ,
		\_2135__reg/NET0131 ,
		_w1880_,
		_w1881_,
		_w1882_
	);
	LUT4 #(
		.INIT('h2772)
	) name374 (
		\TM0_pad ,
		\WX10839_reg/NET0131 ,
		_w1800_,
		_w1801_,
		_w1883_
	);
	LUT4 #(
		.INIT('h028a)
	) name375 (
		RESET_pad,
		\TM1_pad ,
		_w1882_,
		_w1883_,
		_w1884_
	);
	LUT3 #(
		.INIT('h96)
	) name376 (
		\WX11083_reg/NET0131 ,
		\WX11147_reg/NET0131 ,
		\WX11211_reg/NET0131 ,
		_w1885_
	);
	LUT2 #(
		.INIT('h9)
	) name377 (
		\TM1_pad ,
		\WX11019_reg/NET0131 ,
		_w1886_
	);
	LUT4 #(
		.INIT('h2772)
	) name378 (
		\TM0_pad ,
		\_2317__reg/NET0131 ,
		_w1885_,
		_w1886_,
		_w1887_
	);
	LUT4 #(
		.INIT('h2772)
	) name379 (
		\TM0_pad ,
		\WX10859_reg/NET0131 ,
		_w1819_,
		_w1820_,
		_w1888_
	);
	LUT4 #(
		.INIT('h028a)
	) name380 (
		RESET_pad,
		\TM1_pad ,
		_w1887_,
		_w1888_,
		_w1889_
	);
	LUT4 #(
		.INIT('h8cc8)
	) name381 (
		\TM0_pad ,
		_w1810_,
		_w1814_,
		_w1815_,
		_w1890_
	);
	LUT2 #(
		.INIT('h9)
	) name382 (
		\WX5983_reg/NET0131 ,
		\WX6047_reg/NET0131 ,
		_w1891_
	);
	LUT2 #(
		.INIT('h9)
	) name383 (
		\WX5855_reg/NET0131 ,
		\WX5919_reg/NET0131 ,
		_w1892_
	);
	LUT4 #(
		.INIT('h0a02)
	) name384 (
		RESET_pad,
		\TM0_pad ,
		\TM1_pad ,
		\_2185__reg/NET0131 ,
		_w1893_
	);
	LUT4 #(
		.INIT('hbe00)
	) name385 (
		\TM0_pad ,
		_w1891_,
		_w1892_,
		_w1893_,
		_w1894_
	);
	LUT2 #(
		.INIT('he)
	) name386 (
		_w1890_,
		_w1894_,
		_w1895_
	);
	LUT4 #(
		.INIT('h8cc8)
	) name387 (
		\TM0_pad ,
		_w1628_,
		_w1835_,
		_w1836_,
		_w1896_
	);
	LUT2 #(
		.INIT('h9)
	) name388 (
		\WX7274_reg/NET0131 ,
		\WX7338_reg/NET0131 ,
		_w1897_
	);
	LUT2 #(
		.INIT('h9)
	) name389 (
		\WX7146_reg/NET0131 ,
		\WX7210_reg/NET0131 ,
		_w1898_
	);
	LUT4 #(
		.INIT('h0a02)
	) name390 (
		RESET_pad,
		\TM0_pad ,
		\TM1_pad ,
		\_2218__reg/NET0131 ,
		_w1899_
	);
	LUT4 #(
		.INIT('hbe00)
	) name391 (
		\TM0_pad ,
		_w1897_,
		_w1898_,
		_w1899_,
		_w1900_
	);
	LUT2 #(
		.INIT('he)
	) name392 (
		_w1896_,
		_w1900_,
		_w1901_
	);
	LUT4 #(
		.INIT('h8cc8)
	) name393 (
		\TM0_pad ,
		_w1706_,
		_w1841_,
		_w1842_,
		_w1902_
	);
	LUT2 #(
		.INIT('h9)
	) name394 (
		\WX8565_reg/NET0131 ,
		\WX8629_reg/NET0131 ,
		_w1903_
	);
	LUT2 #(
		.INIT('h9)
	) name395 (
		\WX8437_reg/NET0131 ,
		\WX8501_reg/NET0131 ,
		_w1904_
	);
	LUT4 #(
		.INIT('h0a02)
	) name396 (
		RESET_pad,
		\TM0_pad ,
		\TM1_pad ,
		\_2251__reg/NET0131 ,
		_w1905_
	);
	LUT4 #(
		.INIT('hbe00)
	) name397 (
		\TM0_pad ,
		_w1903_,
		_w1904_,
		_w1905_,
		_w1906_
	);
	LUT2 #(
		.INIT('he)
	) name398 (
		_w1902_,
		_w1906_,
		_w1907_
	);
	LUT4 #(
		.INIT('h2772)
	) name399 (
		\TM0_pad ,
		\WX10843_reg/NET0131 ,
		_w1557_,
		_w1558_,
		_w1908_
	);
	LUT3 #(
		.INIT('h96)
	) name400 (
		\WX2016_reg/NET0131 ,
		\WX2080_reg/NET0131 ,
		\WX2144_reg/NET0131 ,
		_w1909_
	);
	LUT2 #(
		.INIT('h9)
	) name401 (
		\TM1_pad ,
		\WX1952_reg/NET0131 ,
		_w1910_
	);
	LUT4 #(
		.INIT('h2772)
	) name402 (
		\TM0_pad ,
		\_2101__reg/NET0131 ,
		_w1909_,
		_w1910_,
		_w1911_
	);
	LUT4 #(
		.INIT('h082a)
	) name403 (
		RESET_pad,
		\TM1_pad ,
		_w1908_,
		_w1911_,
		_w1912_
	);
	LUT3 #(
		.INIT('h96)
	) name404 (
		\WX11063_reg/NET0131 ,
		\WX11127_reg/NET0131 ,
		\WX11191_reg/NET0131 ,
		_w1913_
	);
	LUT2 #(
		.INIT('h9)
	) name405 (
		\TM1_pad ,
		\WX10999_reg/NET0131 ,
		_w1914_
	);
	LUT4 #(
		.INIT('h2772)
	) name406 (
		\TM0_pad ,
		\WX10839_reg/NET0131 ,
		_w1913_,
		_w1914_,
		_w1915_
	);
	LUT2 #(
		.INIT('h2)
	) name407 (
		\TM0_pad ,
		\_2359__reg/NET0131 ,
		_w1916_
	);
	LUT4 #(
		.INIT('h00c8)
	) name408 (
		\DATA_0_26_pad ,
		RESET_pad,
		\TM0_pad ,
		\TM1_pad ,
		_w1917_
	);
	LUT2 #(
		.INIT('h4)
	) name409 (
		_w1916_,
		_w1917_,
		_w1918_
	);
	LUT3 #(
		.INIT('hf2)
	) name410 (
		_w1605_,
		_w1915_,
		_w1918_,
		_w1919_
	);
	LUT2 #(
		.INIT('h8)
	) name411 (
		RESET_pad,
		\WX10837_reg/NET0131 ,
		_w1920_
	);
	LUT4 #(
		.INIT('ha020)
	) name412 (
		RESET_pad,
		\TM0_pad ,
		\TM1_pad ,
		\WX10871_reg/NET0131 ,
		_w1921_
	);
	LUT2 #(
		.INIT('h9)
	) name413 (
		\WX3401_reg/NET0131 ,
		\WX3465_reg/NET0131 ,
		_w1922_
	);
	LUT2 #(
		.INIT('h9)
	) name414 (
		\WX3273_reg/NET0131 ,
		\WX3337_reg/NET0131 ,
		_w1923_
	);
	LUT4 #(
		.INIT('h8cc8)
	) name415 (
		\TM0_pad ,
		_w1921_,
		_w1922_,
		_w1923_,
		_w1924_
	);
	LUT2 #(
		.INIT('h9)
	) name416 (
		\WX4694_reg/NET0131 ,
		\WX4758_reg/NET0131 ,
		_w1925_
	);
	LUT2 #(
		.INIT('h9)
	) name417 (
		\WX4566_reg/NET0131 ,
		\WX4630_reg/NET0131 ,
		_w1926_
	);
	LUT4 #(
		.INIT('h0a02)
	) name418 (
		RESET_pad,
		\TM0_pad ,
		\TM1_pad ,
		\_2151__reg/NET0131 ,
		_w1927_
	);
	LUT4 #(
		.INIT('hbe00)
	) name419 (
		\TM0_pad ,
		_w1925_,
		_w1926_,
		_w1927_,
		_w1928_
	);
	LUT2 #(
		.INIT('he)
	) name420 (
		_w1924_,
		_w1928_,
		_w1929_
	);
	LUT4 #(
		.INIT('h8cc8)
	) name421 (
		\TM0_pad ,
		_w1706_,
		_w1903_,
		_w1904_,
		_w1930_
	);
	LUT2 #(
		.INIT('h9)
	) name422 (
		\WX9858_reg/NET0131 ,
		\WX9922_reg/NET0131 ,
		_w1931_
	);
	LUT2 #(
		.INIT('h9)
	) name423 (
		\WX9730_reg/NET0131 ,
		\WX9794_reg/NET0131 ,
		_w1932_
	);
	LUT4 #(
		.INIT('h0a02)
	) name424 (
		RESET_pad,
		\TM0_pad ,
		\TM1_pad ,
		\_2283__reg/NET0131 ,
		_w1933_
	);
	LUT4 #(
		.INIT('hbe00)
	) name425 (
		\TM0_pad ,
		_w1931_,
		_w1932_,
		_w1933_,
		_w1934_
	);
	LUT2 #(
		.INIT('he)
	) name426 (
		_w1930_,
		_w1934_,
		_w1935_
	);
	LUT3 #(
		.INIT('h96)
	) name427 (
		\WX3307_reg/NET0131 ,
		\WX3371_reg/NET0131 ,
		\WX3435_reg/NET0131 ,
		_w1936_
	);
	LUT2 #(
		.INIT('h9)
	) name428 (
		\TM1_pad ,
		\WX3243_reg/NET0131 ,
		_w1937_
	);
	LUT4 #(
		.INIT('h2772)
	) name429 (
		\TM0_pad ,
		\_2134__reg/NET0131 ,
		_w1936_,
		_w1937_,
		_w1938_
	);
	LUT4 #(
		.INIT('h2772)
	) name430 (
		\TM0_pad ,
		\WX10841_reg/NET0131 ,
		_w1853_,
		_w1854_,
		_w1939_
	);
	LUT4 #(
		.INIT('h028a)
	) name431 (
		RESET_pad,
		\TM1_pad ,
		_w1938_,
		_w1939_,
		_w1940_
	);
	LUT4 #(
		.INIT('h8cc8)
	) name432 (
		\TM0_pad ,
		_w1606_,
		_w1875_,
		_w1876_,
		_w1941_
	);
	LUT2 #(
		.INIT('h9)
	) name433 (
		\WX11149_reg/NET0131 ,
		\WX11213_reg/NET0131 ,
		_w1942_
	);
	LUT2 #(
		.INIT('h9)
	) name434 (
		\WX11021_reg/NET0131 ,
		\WX11085_reg/NET0131 ,
		_w1943_
	);
	LUT4 #(
		.INIT('h0a02)
	) name435 (
		RESET_pad,
		\TM0_pad ,
		\TM1_pad ,
		\_2316__reg/NET0131 ,
		_w1944_
	);
	LUT4 #(
		.INIT('hbe00)
	) name436 (
		\TM0_pad ,
		_w1942_,
		_w1943_,
		_w1944_,
		_w1945_
	);
	LUT2 #(
		.INIT('he)
	) name437 (
		_w1941_,
		_w1945_,
		_w1946_
	);
	LUT4 #(
		.INIT('h8cc8)
	) name438 (
		\TM0_pad ,
		_w1865_,
		_w1869_,
		_w1870_,
		_w1947_
	);
	LUT2 #(
		.INIT('h9)
	) name439 (
		\WX5985_reg/NET0131 ,
		\WX6049_reg/NET0131 ,
		_w1948_
	);
	LUT2 #(
		.INIT('h9)
	) name440 (
		\WX5857_reg/NET0131 ,
		\WX5921_reg/NET0131 ,
		_w1949_
	);
	LUT4 #(
		.INIT('h0a02)
	) name441 (
		RESET_pad,
		\TM0_pad ,
		\TM1_pad ,
		\_2184__reg/NET0131 ,
		_w1950_
	);
	LUT4 #(
		.INIT('hbe00)
	) name442 (
		\TM0_pad ,
		_w1948_,
		_w1949_,
		_w1950_,
		_w1951_
	);
	LUT2 #(
		.INIT('he)
	) name443 (
		_w1947_,
		_w1951_,
		_w1952_
	);
	LUT4 #(
		.INIT('h8cc8)
	) name444 (
		\TM0_pad ,
		_w1810_,
		_w1891_,
		_w1892_,
		_w1953_
	);
	LUT2 #(
		.INIT('h9)
	) name445 (
		\WX7276_reg/NET0131 ,
		\WX7340_reg/NET0131 ,
		_w1954_
	);
	LUT2 #(
		.INIT('h9)
	) name446 (
		\WX7148_reg/NET0131 ,
		\WX7212_reg/NET0131 ,
		_w1955_
	);
	LUT4 #(
		.INIT('h0a02)
	) name447 (
		RESET_pad,
		\TM0_pad ,
		\TM1_pad ,
		\_2217__reg/NET0131 ,
		_w1956_
	);
	LUT4 #(
		.INIT('hbe00)
	) name448 (
		\TM0_pad ,
		_w1954_,
		_w1955_,
		_w1956_,
		_w1957_
	);
	LUT2 #(
		.INIT('he)
	) name449 (
		_w1953_,
		_w1957_,
		_w1958_
	);
	LUT4 #(
		.INIT('h8cc8)
	) name450 (
		\TM0_pad ,
		_w1628_,
		_w1897_,
		_w1898_,
		_w1959_
	);
	LUT2 #(
		.INIT('h9)
	) name451 (
		\WX8567_reg/NET0131 ,
		\WX8631_reg/NET0131 ,
		_w1960_
	);
	LUT2 #(
		.INIT('h9)
	) name452 (
		\WX8439_reg/NET0131 ,
		\WX8503_reg/NET0131 ,
		_w1961_
	);
	LUT4 #(
		.INIT('h0a02)
	) name453 (
		RESET_pad,
		\TM0_pad ,
		\TM1_pad ,
		\_2250__reg/NET0131 ,
		_w1962_
	);
	LUT4 #(
		.INIT('hbe00)
	) name454 (
		\TM0_pad ,
		_w1960_,
		_w1961_,
		_w1962_,
		_w1963_
	);
	LUT2 #(
		.INIT('he)
	) name455 (
		_w1959_,
		_w1963_,
		_w1964_
	);
	LUT4 #(
		.INIT('h2772)
	) name456 (
		\TM0_pad ,
		\WX10845_reg/NET0131 ,
		_w1554_,
		_w1555_,
		_w1965_
	);
	LUT3 #(
		.INIT('h96)
	) name457 (
		\WX2018_reg/NET0131 ,
		\WX2082_reg/NET0131 ,
		\WX2146_reg/NET0131 ,
		_w1966_
	);
	LUT2 #(
		.INIT('h9)
	) name458 (
		\TM1_pad ,
		\WX1954_reg/NET0131 ,
		_w1967_
	);
	LUT4 #(
		.INIT('h2772)
	) name459 (
		\TM0_pad ,
		\_2100__reg/NET0131 ,
		_w1966_,
		_w1967_,
		_w1968_
	);
	LUT4 #(
		.INIT('h082a)
	) name460 (
		RESET_pad,
		\TM1_pad ,
		_w1965_,
		_w1968_,
		_w1969_
	);
	LUT3 #(
		.INIT('h96)
	) name461 (
		\WX11065_reg/NET0131 ,
		\WX11129_reg/NET0131 ,
		\WX11193_reg/NET0131 ,
		_w1970_
	);
	LUT2 #(
		.INIT('h9)
	) name462 (
		\TM1_pad ,
		\WX11001_reg/NET0131 ,
		_w1971_
	);
	LUT4 #(
		.INIT('h2772)
	) name463 (
		\TM0_pad ,
		\WX10841_reg/NET0131 ,
		_w1970_,
		_w1971_,
		_w1972_
	);
	LUT2 #(
		.INIT('h2)
	) name464 (
		\TM0_pad ,
		\_2358__reg/NET0131 ,
		_w1973_
	);
	LUT4 #(
		.INIT('h00c8)
	) name465 (
		\DATA_0_25_pad ,
		RESET_pad,
		\TM0_pad ,
		\TM1_pad ,
		_w1974_
	);
	LUT2 #(
		.INIT('h4)
	) name466 (
		_w1973_,
		_w1974_,
		_w1975_
	);
	LUT3 #(
		.INIT('hf2)
	) name467 (
		_w1605_,
		_w1972_,
		_w1975_,
		_w1976_
	);
	LUT2 #(
		.INIT('h8)
	) name468 (
		RESET_pad,
		\WX10839_reg/NET0131 ,
		_w1977_
	);
	LUT4 #(
		.INIT('ha020)
	) name469 (
		RESET_pad,
		\TM0_pad ,
		\TM1_pad ,
		\WX10873_reg/NET0131 ,
		_w1978_
	);
	LUT2 #(
		.INIT('h9)
	) name470 (
		\WX3403_reg/NET0131 ,
		\WX3467_reg/NET0131 ,
		_w1979_
	);
	LUT2 #(
		.INIT('h9)
	) name471 (
		\WX3275_reg/NET0131 ,
		\WX3339_reg/NET0131 ,
		_w1980_
	);
	LUT4 #(
		.INIT('h8cc8)
	) name472 (
		\TM0_pad ,
		_w1978_,
		_w1979_,
		_w1980_,
		_w1981_
	);
	LUT2 #(
		.INIT('h9)
	) name473 (
		\WX4696_reg/NET0131 ,
		\WX4760_reg/NET0131 ,
		_w1982_
	);
	LUT2 #(
		.INIT('h9)
	) name474 (
		\WX4568_reg/NET0131 ,
		\WX4632_reg/NET0131 ,
		_w1983_
	);
	LUT4 #(
		.INIT('h0a02)
	) name475 (
		RESET_pad,
		\TM0_pad ,
		\TM1_pad ,
		\_2150__reg/NET0131 ,
		_w1984_
	);
	LUT4 #(
		.INIT('hbe00)
	) name476 (
		\TM0_pad ,
		_w1982_,
		_w1983_,
		_w1984_,
		_w1985_
	);
	LUT2 #(
		.INIT('he)
	) name477 (
		_w1981_,
		_w1985_,
		_w1986_
	);
	LUT4 #(
		.INIT('h8cc8)
	) name478 (
		\TM0_pad ,
		_w1628_,
		_w1960_,
		_w1961_,
		_w1987_
	);
	LUT2 #(
		.INIT('h9)
	) name479 (
		\WX9860_reg/NET0131 ,
		\WX9924_reg/NET0131 ,
		_w1988_
	);
	LUT2 #(
		.INIT('h9)
	) name480 (
		\WX9732_reg/NET0131 ,
		\WX9796_reg/NET0131 ,
		_w1989_
	);
	LUT4 #(
		.INIT('h0a02)
	) name481 (
		RESET_pad,
		\TM0_pad ,
		\TM1_pad ,
		\_2282__reg/NET0131 ,
		_w1990_
	);
	LUT4 #(
		.INIT('hbe00)
	) name482 (
		\TM0_pad ,
		_w1988_,
		_w1989_,
		_w1990_,
		_w1991_
	);
	LUT2 #(
		.INIT('he)
	) name483 (
		_w1987_,
		_w1991_,
		_w1992_
	);
	LUT4 #(
		.INIT('h8cc8)
	) name484 (
		\TM0_pad ,
		_w1706_,
		_w1931_,
		_w1932_,
		_w1993_
	);
	LUT2 #(
		.INIT('h9)
	) name485 (
		\WX11151_reg/NET0131 ,
		\WX11215_reg/NET0131 ,
		_w1994_
	);
	LUT2 #(
		.INIT('h9)
	) name486 (
		\WX11023_reg/NET0131 ,
		\WX11087_reg/NET0131 ,
		_w1995_
	);
	LUT4 #(
		.INIT('h0a02)
	) name487 (
		RESET_pad,
		\TM0_pad ,
		\TM1_pad ,
		\_2315__reg/NET0131 ,
		_w1996_
	);
	LUT4 #(
		.INIT('hbe00)
	) name488 (
		\TM0_pad ,
		_w1994_,
		_w1995_,
		_w1996_,
		_w1997_
	);
	LUT2 #(
		.INIT('he)
	) name489 (
		_w1993_,
		_w1997_,
		_w1998_
	);
	LUT3 #(
		.INIT('h96)
	) name490 (
		\WX3309_reg/NET0131 ,
		\WX3373_reg/NET0131 ,
		\WX3437_reg/NET0131 ,
		_w1999_
	);
	LUT2 #(
		.INIT('h9)
	) name491 (
		\TM1_pad ,
		\WX3245_reg/NET0131 ,
		_w2000_
	);
	LUT4 #(
		.INIT('h2772)
	) name492 (
		\TM0_pad ,
		\_2133__reg/NET0131 ,
		_w1999_,
		_w2000_,
		_w2001_
	);
	LUT4 #(
		.INIT('h2772)
	) name493 (
		\TM0_pad ,
		\WX10843_reg/NET0131 ,
		_w1909_,
		_w1910_,
		_w2002_
	);
	LUT4 #(
		.INIT('h028a)
	) name494 (
		RESET_pad,
		\TM1_pad ,
		_w2001_,
		_w2002_,
		_w2003_
	);
	LUT4 #(
		.INIT('h8cc8)
	) name495 (
		\TM0_pad ,
		_w1921_,
		_w1925_,
		_w1926_,
		_w2004_
	);
	LUT2 #(
		.INIT('h9)
	) name496 (
		\WX5987_reg/NET0131 ,
		\WX6051_reg/NET0131 ,
		_w2005_
	);
	LUT2 #(
		.INIT('h9)
	) name497 (
		\WX5859_reg/NET0131 ,
		\WX5923_reg/NET0131 ,
		_w2006_
	);
	LUT4 #(
		.INIT('h0a02)
	) name498 (
		RESET_pad,
		\TM0_pad ,
		\TM1_pad ,
		\_2183__reg/NET0131 ,
		_w2007_
	);
	LUT4 #(
		.INIT('hbe00)
	) name499 (
		\TM0_pad ,
		_w2005_,
		_w2006_,
		_w2007_,
		_w2008_
	);
	LUT2 #(
		.INIT('he)
	) name500 (
		_w2004_,
		_w2008_,
		_w2009_
	);
	LUT4 #(
		.INIT('h8cc8)
	) name501 (
		\TM0_pad ,
		_w1865_,
		_w1948_,
		_w1949_,
		_w2010_
	);
	LUT2 #(
		.INIT('h9)
	) name502 (
		\WX7278_reg/NET0131 ,
		\WX7342_reg/NET0131 ,
		_w2011_
	);
	LUT2 #(
		.INIT('h9)
	) name503 (
		\WX7150_reg/NET0131 ,
		\WX7214_reg/NET0131 ,
		_w2012_
	);
	LUT4 #(
		.INIT('h0a02)
	) name504 (
		RESET_pad,
		\TM0_pad ,
		\TM1_pad ,
		\_2216__reg/NET0131 ,
		_w2013_
	);
	LUT4 #(
		.INIT('hbe00)
	) name505 (
		\TM0_pad ,
		_w2011_,
		_w2012_,
		_w2013_,
		_w2014_
	);
	LUT2 #(
		.INIT('he)
	) name506 (
		_w2010_,
		_w2014_,
		_w2015_
	);
	LUT4 #(
		.INIT('h8cc8)
	) name507 (
		\TM0_pad ,
		_w1810_,
		_w1954_,
		_w1955_,
		_w2016_
	);
	LUT2 #(
		.INIT('h9)
	) name508 (
		\WX8569_reg/NET0131 ,
		\WX8633_reg/NET0131 ,
		_w2017_
	);
	LUT2 #(
		.INIT('h9)
	) name509 (
		\WX8441_reg/NET0131 ,
		\WX8505_reg/NET0131 ,
		_w2018_
	);
	LUT4 #(
		.INIT('h0a02)
	) name510 (
		RESET_pad,
		\TM0_pad ,
		\TM1_pad ,
		\_2249__reg/NET0131 ,
		_w2019_
	);
	LUT4 #(
		.INIT('hbe00)
	) name511 (
		\TM0_pad ,
		_w2017_,
		_w2018_,
		_w2019_,
		_w2020_
	);
	LUT2 #(
		.INIT('he)
	) name512 (
		_w2016_,
		_w2020_,
		_w2021_
	);
	LUT4 #(
		.INIT('h2772)
	) name513 (
		\TM0_pad ,
		\WX10847_reg/NET0131 ,
		_w1551_,
		_w1552_,
		_w2022_
	);
	LUT3 #(
		.INIT('h96)
	) name514 (
		\WX2020_reg/NET0131 ,
		\WX2084_reg/NET0131 ,
		\WX2148_reg/NET0131 ,
		_w2023_
	);
	LUT2 #(
		.INIT('h9)
	) name515 (
		\TM1_pad ,
		\WX1956_reg/NET0131 ,
		_w2024_
	);
	LUT4 #(
		.INIT('h2772)
	) name516 (
		\TM0_pad ,
		\_2099__reg/NET0131 ,
		_w2023_,
		_w2024_,
		_w2025_
	);
	LUT4 #(
		.INIT('h082a)
	) name517 (
		RESET_pad,
		\TM1_pad ,
		_w2022_,
		_w2025_,
		_w2026_
	);
	LUT3 #(
		.INIT('h96)
	) name518 (
		\WX11067_reg/NET0131 ,
		\WX11131_reg/NET0131 ,
		\WX11195_reg/NET0131 ,
		_w2027_
	);
	LUT2 #(
		.INIT('h9)
	) name519 (
		\TM1_pad ,
		\WX11003_reg/NET0131 ,
		_w2028_
	);
	LUT4 #(
		.INIT('h2772)
	) name520 (
		\TM0_pad ,
		\WX10843_reg/NET0131 ,
		_w2027_,
		_w2028_,
		_w2029_
	);
	LUT2 #(
		.INIT('h2)
	) name521 (
		\TM0_pad ,
		\_2357__reg/NET0131 ,
		_w2030_
	);
	LUT4 #(
		.INIT('h00c8)
	) name522 (
		\DATA_0_24_pad ,
		RESET_pad,
		\TM0_pad ,
		\TM1_pad ,
		_w2031_
	);
	LUT2 #(
		.INIT('h4)
	) name523 (
		_w2030_,
		_w2031_,
		_w2032_
	);
	LUT3 #(
		.INIT('hf2)
	) name524 (
		_w1605_,
		_w2029_,
		_w2032_,
		_w2033_
	);
	LUT2 #(
		.INIT('h8)
	) name525 (
		RESET_pad,
		\WX10841_reg/NET0131 ,
		_w2034_
	);
	LUT2 #(
		.INIT('h9)
	) name526 (
		\WX3405_reg/NET0131 ,
		\WX3469_reg/NET0131 ,
		_w2035_
	);
	LUT2 #(
		.INIT('h9)
	) name527 (
		\WX3277_reg/NET0131 ,
		\WX3341_reg/NET0131 ,
		_w2036_
	);
	LUT4 #(
		.INIT('h8cc8)
	) name528 (
		\TM0_pad ,
		_w1620_,
		_w2035_,
		_w2036_,
		_w2037_
	);
	LUT2 #(
		.INIT('h9)
	) name529 (
		\WX4698_reg/NET0131 ,
		\WX4762_reg/NET0131 ,
		_w2038_
	);
	LUT2 #(
		.INIT('h9)
	) name530 (
		\WX4570_reg/NET0131 ,
		\WX4634_reg/NET0131 ,
		_w2039_
	);
	LUT4 #(
		.INIT('h0a02)
	) name531 (
		RESET_pad,
		\TM0_pad ,
		\TM1_pad ,
		\_2149__reg/NET0131 ,
		_w2040_
	);
	LUT4 #(
		.INIT('hbe00)
	) name532 (
		\TM0_pad ,
		_w2038_,
		_w2039_,
		_w2040_,
		_w2041_
	);
	LUT2 #(
		.INIT('he)
	) name533 (
		_w2037_,
		_w2041_,
		_w2042_
	);
	LUT4 #(
		.INIT('h8cc8)
	) name534 (
		\TM0_pad ,
		_w1810_,
		_w2017_,
		_w2018_,
		_w2043_
	);
	LUT2 #(
		.INIT('h9)
	) name535 (
		\WX9862_reg/NET0131 ,
		\WX9926_reg/NET0131 ,
		_w2044_
	);
	LUT2 #(
		.INIT('h9)
	) name536 (
		\WX9734_reg/NET0131 ,
		\WX9798_reg/NET0131 ,
		_w2045_
	);
	LUT4 #(
		.INIT('h0a02)
	) name537 (
		RESET_pad,
		\TM0_pad ,
		\TM1_pad ,
		\_2281__reg/NET0131 ,
		_w2046_
	);
	LUT4 #(
		.INIT('hbe00)
	) name538 (
		\TM0_pad ,
		_w2044_,
		_w2045_,
		_w2046_,
		_w2047_
	);
	LUT2 #(
		.INIT('he)
	) name539 (
		_w2043_,
		_w2047_,
		_w2048_
	);
	LUT4 #(
		.INIT('h8cc8)
	) name540 (
		\TM0_pad ,
		_w1628_,
		_w1988_,
		_w1989_,
		_w2049_
	);
	LUT4 #(
		.INIT('h0a02)
	) name541 (
		RESET_pad,
		\TM0_pad ,
		\TM1_pad ,
		\_2314__reg/NET0131 ,
		_w2050_
	);
	LUT4 #(
		.INIT('hbe00)
	) name542 (
		\TM0_pad ,
		_w1629_,
		_w1630_,
		_w2050_,
		_w2051_
	);
	LUT2 #(
		.INIT('he)
	) name543 (
		_w2049_,
		_w2051_,
		_w2052_
	);
	LUT3 #(
		.INIT('h96)
	) name544 (
		\WX3311_reg/NET0131 ,
		\WX3375_reg/NET0131 ,
		\WX3439_reg/NET0131 ,
		_w2053_
	);
	LUT2 #(
		.INIT('h9)
	) name545 (
		\TM1_pad ,
		\WX3247_reg/NET0131 ,
		_w2054_
	);
	LUT4 #(
		.INIT('h2772)
	) name546 (
		\TM0_pad ,
		\_2132__reg/NET0131 ,
		_w2053_,
		_w2054_,
		_w2055_
	);
	LUT4 #(
		.INIT('h2772)
	) name547 (
		\TM0_pad ,
		\WX10845_reg/NET0131 ,
		_w1966_,
		_w1967_,
		_w2056_
	);
	LUT4 #(
		.INIT('h028a)
	) name548 (
		RESET_pad,
		\TM1_pad ,
		_w2055_,
		_w2056_,
		_w2057_
	);
	LUT4 #(
		.INIT('h8cc8)
	) name549 (
		\TM0_pad ,
		_w1978_,
		_w1982_,
		_w1983_,
		_w2058_
	);
	LUT2 #(
		.INIT('h9)
	) name550 (
		\WX5989_reg/NET0131 ,
		\WX6053_reg/NET0131 ,
		_w2059_
	);
	LUT2 #(
		.INIT('h9)
	) name551 (
		\WX5861_reg/NET0131 ,
		\WX5925_reg/NET0131 ,
		_w2060_
	);
	LUT4 #(
		.INIT('h0a02)
	) name552 (
		RESET_pad,
		\TM0_pad ,
		\TM1_pad ,
		\_2182__reg/NET0131 ,
		_w2061_
	);
	LUT4 #(
		.INIT('hbe00)
	) name553 (
		\TM0_pad ,
		_w2059_,
		_w2060_,
		_w2061_,
		_w2062_
	);
	LUT2 #(
		.INIT('he)
	) name554 (
		_w2058_,
		_w2062_,
		_w2063_
	);
	LUT4 #(
		.INIT('h8cc8)
	) name555 (
		\TM0_pad ,
		_w1921_,
		_w2005_,
		_w2006_,
		_w2064_
	);
	LUT2 #(
		.INIT('h9)
	) name556 (
		\WX7280_reg/NET0131 ,
		\WX7344_reg/NET0131 ,
		_w2065_
	);
	LUT2 #(
		.INIT('h9)
	) name557 (
		\WX7152_reg/NET0131 ,
		\WX7216_reg/NET0131 ,
		_w2066_
	);
	LUT4 #(
		.INIT('h0a02)
	) name558 (
		RESET_pad,
		\TM0_pad ,
		\TM1_pad ,
		\_2215__reg/NET0131 ,
		_w2067_
	);
	LUT4 #(
		.INIT('hbe00)
	) name559 (
		\TM0_pad ,
		_w2065_,
		_w2066_,
		_w2067_,
		_w2068_
	);
	LUT2 #(
		.INIT('he)
	) name560 (
		_w2064_,
		_w2068_,
		_w2069_
	);
	LUT4 #(
		.INIT('h8cc8)
	) name561 (
		\TM0_pad ,
		_w1865_,
		_w2011_,
		_w2012_,
		_w2070_
	);
	LUT2 #(
		.INIT('h9)
	) name562 (
		\WX8571_reg/NET0131 ,
		\WX8635_reg/NET0131 ,
		_w2071_
	);
	LUT2 #(
		.INIT('h9)
	) name563 (
		\WX8443_reg/NET0131 ,
		\WX8507_reg/NET0131 ,
		_w2072_
	);
	LUT4 #(
		.INIT('h0a02)
	) name564 (
		RESET_pad,
		\TM0_pad ,
		\TM1_pad ,
		\_2248__reg/NET0131 ,
		_w2073_
	);
	LUT4 #(
		.INIT('hbe00)
	) name565 (
		\TM0_pad ,
		_w2071_,
		_w2072_,
		_w2073_,
		_w2074_
	);
	LUT2 #(
		.INIT('he)
	) name566 (
		_w2070_,
		_w2074_,
		_w2075_
	);
	LUT4 #(
		.INIT('h2772)
	) name567 (
		\TM0_pad ,
		\WX10849_reg/NET0131 ,
		_w1548_,
		_w1549_,
		_w2076_
	);
	LUT3 #(
		.INIT('h96)
	) name568 (
		\WX2022_reg/NET0131 ,
		\WX2086_reg/NET0131 ,
		\WX2150_reg/NET0131 ,
		_w2077_
	);
	LUT2 #(
		.INIT('h9)
	) name569 (
		\TM1_pad ,
		\WX1958_reg/NET0131 ,
		_w2078_
	);
	LUT4 #(
		.INIT('h2772)
	) name570 (
		\TM0_pad ,
		\_2098__reg/NET0131 ,
		_w2077_,
		_w2078_,
		_w2079_
	);
	LUT4 #(
		.INIT('h082a)
	) name571 (
		RESET_pad,
		\TM1_pad ,
		_w2076_,
		_w2079_,
		_w2080_
	);
	LUT3 #(
		.INIT('h96)
	) name572 (
		\WX11069_reg/NET0131 ,
		\WX11133_reg/NET0131 ,
		\WX11197_reg/NET0131 ,
		_w2081_
	);
	LUT2 #(
		.INIT('h9)
	) name573 (
		\TM1_pad ,
		\WX11005_reg/NET0131 ,
		_w2082_
	);
	LUT4 #(
		.INIT('h2772)
	) name574 (
		\TM0_pad ,
		\WX10845_reg/NET0131 ,
		_w2081_,
		_w2082_,
		_w2083_
	);
	LUT2 #(
		.INIT('h2)
	) name575 (
		\TM0_pad ,
		\_2356__reg/NET0131 ,
		_w2084_
	);
	LUT4 #(
		.INIT('h00c8)
	) name576 (
		\DATA_0_23_pad ,
		RESET_pad,
		\TM0_pad ,
		\TM1_pad ,
		_w2085_
	);
	LUT2 #(
		.INIT('h4)
	) name577 (
		_w2084_,
		_w2085_,
		_w2086_
	);
	LUT3 #(
		.INIT('hf2)
	) name578 (
		_w1605_,
		_w2083_,
		_w2086_,
		_w2087_
	);
	LUT2 #(
		.INIT('h8)
	) name579 (
		RESET_pad,
		\WX10843_reg/NET0131 ,
		_w2088_
	);
	LUT4 #(
		.INIT('ha020)
	) name580 (
		RESET_pad,
		\TM0_pad ,
		\TM1_pad ,
		\WX10877_reg/NET0131 ,
		_w2089_
	);
	LUT2 #(
		.INIT('h9)
	) name581 (
		\WX3407_reg/NET0131 ,
		\WX3471_reg/NET0131 ,
		_w2090_
	);
	LUT2 #(
		.INIT('h9)
	) name582 (
		\WX3279_reg/NET0131 ,
		\WX3343_reg/NET0131 ,
		_w2091_
	);
	LUT4 #(
		.INIT('h8cc8)
	) name583 (
		\TM0_pad ,
		_w2089_,
		_w2090_,
		_w2091_,
		_w2092_
	);
	LUT2 #(
		.INIT('h9)
	) name584 (
		\WX4700_reg/NET0131 ,
		\WX4764_reg/NET0131 ,
		_w2093_
	);
	LUT2 #(
		.INIT('h9)
	) name585 (
		\WX4572_reg/NET0131 ,
		\WX4636_reg/NET0131 ,
		_w2094_
	);
	LUT4 #(
		.INIT('h0a02)
	) name586 (
		RESET_pad,
		\TM0_pad ,
		\TM1_pad ,
		\_2148__reg/NET0131 ,
		_w2095_
	);
	LUT4 #(
		.INIT('hbe00)
	) name587 (
		\TM0_pad ,
		_w2093_,
		_w2094_,
		_w2095_,
		_w2096_
	);
	LUT2 #(
		.INIT('he)
	) name588 (
		_w2092_,
		_w2096_,
		_w2097_
	);
	LUT4 #(
		.INIT('h8cc8)
	) name589 (
		\TM0_pad ,
		_w1865_,
		_w2071_,
		_w2072_,
		_w2098_
	);
	LUT2 #(
		.INIT('h9)
	) name590 (
		\WX9864_reg/NET0131 ,
		\WX9928_reg/NET0131 ,
		_w2099_
	);
	LUT2 #(
		.INIT('h9)
	) name591 (
		\WX9736_reg/NET0131 ,
		\WX9800_reg/NET0131 ,
		_w2100_
	);
	LUT4 #(
		.INIT('h0a02)
	) name592 (
		RESET_pad,
		\TM0_pad ,
		\TM1_pad ,
		\_2280__reg/NET0131 ,
		_w2101_
	);
	LUT4 #(
		.INIT('hbe00)
	) name593 (
		\TM0_pad ,
		_w2099_,
		_w2100_,
		_w2101_,
		_w2102_
	);
	LUT2 #(
		.INIT('he)
	) name594 (
		_w2098_,
		_w2102_,
		_w2103_
	);
	LUT4 #(
		.INIT('h8cc8)
	) name595 (
		\TM0_pad ,
		_w1810_,
		_w2044_,
		_w2045_,
		_w2104_
	);
	LUT2 #(
		.INIT('h9)
	) name596 (
		\WX11155_reg/NET0131 ,
		\WX11219_reg/NET0131 ,
		_w2105_
	);
	LUT2 #(
		.INIT('h9)
	) name597 (
		\WX11027_reg/NET0131 ,
		\WX11091_reg/NET0131 ,
		_w2106_
	);
	LUT4 #(
		.INIT('h0a02)
	) name598 (
		RESET_pad,
		\TM0_pad ,
		\TM1_pad ,
		\_2313__reg/NET0131 ,
		_w2107_
	);
	LUT4 #(
		.INIT('hbe00)
	) name599 (
		\TM0_pad ,
		_w2105_,
		_w2106_,
		_w2107_,
		_w2108_
	);
	LUT2 #(
		.INIT('he)
	) name600 (
		_w2104_,
		_w2108_,
		_w2109_
	);
	LUT3 #(
		.INIT('h96)
	) name601 (
		\WX3313_reg/NET0131 ,
		\WX3377_reg/NET0131 ,
		\WX3441_reg/NET0131 ,
		_w2110_
	);
	LUT2 #(
		.INIT('h9)
	) name602 (
		\TM1_pad ,
		\WX3249_reg/NET0131 ,
		_w2111_
	);
	LUT4 #(
		.INIT('h2772)
	) name603 (
		\TM0_pad ,
		\_2131__reg/NET0131 ,
		_w2110_,
		_w2111_,
		_w2112_
	);
	LUT4 #(
		.INIT('h2772)
	) name604 (
		\TM0_pad ,
		\WX10847_reg/NET0131 ,
		_w2023_,
		_w2024_,
		_w2113_
	);
	LUT4 #(
		.INIT('h028a)
	) name605 (
		RESET_pad,
		\TM1_pad ,
		_w2112_,
		_w2113_,
		_w2114_
	);
	LUT4 #(
		.INIT('h8cc8)
	) name606 (
		\TM0_pad ,
		_w1620_,
		_w2038_,
		_w2039_,
		_w2115_
	);
	LUT2 #(
		.INIT('h9)
	) name607 (
		\WX5991_reg/NET0131 ,
		\WX6055_reg/NET0131 ,
		_w2116_
	);
	LUT2 #(
		.INIT('h9)
	) name608 (
		\WX5863_reg/NET0131 ,
		\WX5927_reg/NET0131 ,
		_w2117_
	);
	LUT4 #(
		.INIT('h0a02)
	) name609 (
		RESET_pad,
		\TM0_pad ,
		\TM1_pad ,
		\_2181__reg/NET0131 ,
		_w2118_
	);
	LUT4 #(
		.INIT('hbe00)
	) name610 (
		\TM0_pad ,
		_w2116_,
		_w2117_,
		_w2118_,
		_w2119_
	);
	LUT2 #(
		.INIT('he)
	) name611 (
		_w2115_,
		_w2119_,
		_w2120_
	);
	LUT4 #(
		.INIT('h8cc8)
	) name612 (
		\TM0_pad ,
		_w1978_,
		_w2059_,
		_w2060_,
		_w2121_
	);
	LUT2 #(
		.INIT('h9)
	) name613 (
		\WX7282_reg/NET0131 ,
		\WX7346_reg/NET0131 ,
		_w2122_
	);
	LUT2 #(
		.INIT('h9)
	) name614 (
		\WX7154_reg/NET0131 ,
		\WX7218_reg/NET0131 ,
		_w2123_
	);
	LUT4 #(
		.INIT('h0a02)
	) name615 (
		RESET_pad,
		\TM0_pad ,
		\TM1_pad ,
		\_2214__reg/NET0131 ,
		_w2124_
	);
	LUT4 #(
		.INIT('hbe00)
	) name616 (
		\TM0_pad ,
		_w2122_,
		_w2123_,
		_w2124_,
		_w2125_
	);
	LUT2 #(
		.INIT('he)
	) name617 (
		_w2121_,
		_w2125_,
		_w2126_
	);
	LUT4 #(
		.INIT('h8cc8)
	) name618 (
		\TM0_pad ,
		_w1921_,
		_w2065_,
		_w2066_,
		_w2127_
	);
	LUT2 #(
		.INIT('h9)
	) name619 (
		\WX8573_reg/NET0131 ,
		\WX8637_reg/NET0131 ,
		_w2128_
	);
	LUT2 #(
		.INIT('h9)
	) name620 (
		\WX8445_reg/NET0131 ,
		\WX8509_reg/NET0131 ,
		_w2129_
	);
	LUT4 #(
		.INIT('h0a02)
	) name621 (
		RESET_pad,
		\TM0_pad ,
		\TM1_pad ,
		\_2247__reg/NET0131 ,
		_w2130_
	);
	LUT4 #(
		.INIT('hbe00)
	) name622 (
		\TM0_pad ,
		_w2128_,
		_w2129_,
		_w2130_,
		_w2131_
	);
	LUT2 #(
		.INIT('he)
	) name623 (
		_w2127_,
		_w2131_,
		_w2132_
	);
	LUT4 #(
		.INIT('h2772)
	) name624 (
		\TM0_pad ,
		\WX10851_reg/NET0131 ,
		_w1545_,
		_w1546_,
		_w2133_
	);
	LUT3 #(
		.INIT('h96)
	) name625 (
		\WX2024_reg/NET0131 ,
		\WX2088_reg/NET0131 ,
		\WX2152_reg/NET0131 ,
		_w2134_
	);
	LUT2 #(
		.INIT('h9)
	) name626 (
		\TM1_pad ,
		\WX1960_reg/NET0131 ,
		_w2135_
	);
	LUT4 #(
		.INIT('h2772)
	) name627 (
		\TM0_pad ,
		\_2097__reg/NET0131 ,
		_w2134_,
		_w2135_,
		_w2136_
	);
	LUT4 #(
		.INIT('h082a)
	) name628 (
		RESET_pad,
		\TM1_pad ,
		_w2133_,
		_w2136_,
		_w2137_
	);
	LUT3 #(
		.INIT('h96)
	) name629 (
		\WX11071_reg/NET0131 ,
		\WX11135_reg/NET0131 ,
		\WX11199_reg/NET0131 ,
		_w2138_
	);
	LUT2 #(
		.INIT('h9)
	) name630 (
		\TM1_pad ,
		\WX11007_reg/NET0131 ,
		_w2139_
	);
	LUT4 #(
		.INIT('h2772)
	) name631 (
		\TM0_pad ,
		\WX10847_reg/NET0131 ,
		_w2138_,
		_w2139_,
		_w2140_
	);
	LUT2 #(
		.INIT('h2)
	) name632 (
		\TM0_pad ,
		\_2355__reg/NET0131 ,
		_w2141_
	);
	LUT4 #(
		.INIT('h00c8)
	) name633 (
		\DATA_0_22_pad ,
		RESET_pad,
		\TM0_pad ,
		\TM1_pad ,
		_w2142_
	);
	LUT2 #(
		.INIT('h4)
	) name634 (
		_w2141_,
		_w2142_,
		_w2143_
	);
	LUT3 #(
		.INIT('hf2)
	) name635 (
		_w1605_,
		_w2140_,
		_w2143_,
		_w2144_
	);
	LUT2 #(
		.INIT('h8)
	) name636 (
		RESET_pad,
		\WX10845_reg/NET0131 ,
		_w2145_
	);
	LUT4 #(
		.INIT('ha020)
	) name637 (
		RESET_pad,
		\TM0_pad ,
		\TM1_pad ,
		\WX10879_reg/NET0131 ,
		_w2146_
	);
	LUT2 #(
		.INIT('h9)
	) name638 (
		\WX3409_reg/NET0131 ,
		\WX3473_reg/NET0131 ,
		_w2147_
	);
	LUT2 #(
		.INIT('h9)
	) name639 (
		\WX3281_reg/NET0131 ,
		\WX3345_reg/NET0131 ,
		_w2148_
	);
	LUT4 #(
		.INIT('h8cc8)
	) name640 (
		\TM0_pad ,
		_w2146_,
		_w2147_,
		_w2148_,
		_w2149_
	);
	LUT2 #(
		.INIT('h9)
	) name641 (
		\WX4702_reg/NET0131 ,
		\WX4766_reg/NET0131 ,
		_w2150_
	);
	LUT2 #(
		.INIT('h9)
	) name642 (
		\WX4574_reg/NET0131 ,
		\WX4638_reg/NET0131 ,
		_w2151_
	);
	LUT4 #(
		.INIT('h0a02)
	) name643 (
		RESET_pad,
		\TM0_pad ,
		\TM1_pad ,
		\_2147__reg/NET0131 ,
		_w2152_
	);
	LUT4 #(
		.INIT('hbe00)
	) name644 (
		\TM0_pad ,
		_w2150_,
		_w2151_,
		_w2152_,
		_w2153_
	);
	LUT2 #(
		.INIT('he)
	) name645 (
		_w2149_,
		_w2153_,
		_w2154_
	);
	LUT4 #(
		.INIT('h8cc8)
	) name646 (
		\TM0_pad ,
		_w1921_,
		_w2128_,
		_w2129_,
		_w2155_
	);
	LUT2 #(
		.INIT('h9)
	) name647 (
		\WX9866_reg/NET0131 ,
		\WX9930_reg/NET0131 ,
		_w2156_
	);
	LUT2 #(
		.INIT('h9)
	) name648 (
		\WX9738_reg/NET0131 ,
		\WX9802_reg/NET0131 ,
		_w2157_
	);
	LUT4 #(
		.INIT('h0a02)
	) name649 (
		RESET_pad,
		\TM0_pad ,
		\TM1_pad ,
		\_2279__reg/NET0131 ,
		_w2158_
	);
	LUT4 #(
		.INIT('hbe00)
	) name650 (
		\TM0_pad ,
		_w2156_,
		_w2157_,
		_w2158_,
		_w2159_
	);
	LUT2 #(
		.INIT('he)
	) name651 (
		_w2155_,
		_w2159_,
		_w2160_
	);
	LUT4 #(
		.INIT('h8cc8)
	) name652 (
		\TM0_pad ,
		_w1865_,
		_w2099_,
		_w2100_,
		_w2161_
	);
	LUT2 #(
		.INIT('h9)
	) name653 (
		\WX11157_reg/NET0131 ,
		\WX11221_reg/NET0131 ,
		_w2162_
	);
	LUT2 #(
		.INIT('h9)
	) name654 (
		\WX11029_reg/NET0131 ,
		\WX11093_reg/NET0131 ,
		_w2163_
	);
	LUT4 #(
		.INIT('h0a02)
	) name655 (
		RESET_pad,
		\TM0_pad ,
		\TM1_pad ,
		\_2312__reg/NET0131 ,
		_w2164_
	);
	LUT4 #(
		.INIT('hbe00)
	) name656 (
		\TM0_pad ,
		_w2162_,
		_w2163_,
		_w2164_,
		_w2165_
	);
	LUT2 #(
		.INIT('he)
	) name657 (
		_w2161_,
		_w2165_,
		_w2166_
	);
	LUT3 #(
		.INIT('h96)
	) name658 (
		\WX3315_reg/NET0131 ,
		\WX3379_reg/NET0131 ,
		\WX3443_reg/NET0131 ,
		_w2167_
	);
	LUT2 #(
		.INIT('h9)
	) name659 (
		\TM1_pad ,
		\WX3251_reg/NET0131 ,
		_w2168_
	);
	LUT4 #(
		.INIT('h2772)
	) name660 (
		\TM0_pad ,
		\_2130__reg/NET0131 ,
		_w2167_,
		_w2168_,
		_w2169_
	);
	LUT4 #(
		.INIT('h2772)
	) name661 (
		\TM0_pad ,
		\WX10849_reg/NET0131 ,
		_w2077_,
		_w2078_,
		_w2170_
	);
	LUT4 #(
		.INIT('h028a)
	) name662 (
		RESET_pad,
		\TM1_pad ,
		_w2169_,
		_w2170_,
		_w2171_
	);
	LUT4 #(
		.INIT('h8cc8)
	) name663 (
		\TM0_pad ,
		_w2089_,
		_w2093_,
		_w2094_,
		_w2172_
	);
	LUT2 #(
		.INIT('h9)
	) name664 (
		\WX5993_reg/NET0131 ,
		\WX6057_reg/NET0131 ,
		_w2173_
	);
	LUT2 #(
		.INIT('h9)
	) name665 (
		\WX5865_reg/NET0131 ,
		\WX5929_reg/NET0131 ,
		_w2174_
	);
	LUT4 #(
		.INIT('h0a02)
	) name666 (
		RESET_pad,
		\TM0_pad ,
		\TM1_pad ,
		\_2180__reg/NET0131 ,
		_w2175_
	);
	LUT4 #(
		.INIT('hbe00)
	) name667 (
		\TM0_pad ,
		_w2173_,
		_w2174_,
		_w2175_,
		_w2176_
	);
	LUT2 #(
		.INIT('he)
	) name668 (
		_w2172_,
		_w2176_,
		_w2177_
	);
	LUT4 #(
		.INIT('h8cc8)
	) name669 (
		\TM0_pad ,
		_w1620_,
		_w2116_,
		_w2117_,
		_w2178_
	);
	LUT2 #(
		.INIT('h9)
	) name670 (
		\WX7284_reg/NET0131 ,
		\WX7348_reg/NET0131 ,
		_w2179_
	);
	LUT2 #(
		.INIT('h9)
	) name671 (
		\WX7156_reg/NET0131 ,
		\WX7220_reg/NET0131 ,
		_w2180_
	);
	LUT4 #(
		.INIT('h0a02)
	) name672 (
		RESET_pad,
		\TM0_pad ,
		\TM1_pad ,
		\_2213__reg/NET0131 ,
		_w2181_
	);
	LUT4 #(
		.INIT('hbe00)
	) name673 (
		\TM0_pad ,
		_w2179_,
		_w2180_,
		_w2181_,
		_w2182_
	);
	LUT2 #(
		.INIT('he)
	) name674 (
		_w2178_,
		_w2182_,
		_w2183_
	);
	LUT4 #(
		.INIT('h8cc8)
	) name675 (
		\TM0_pad ,
		_w1978_,
		_w2122_,
		_w2123_,
		_w2184_
	);
	LUT2 #(
		.INIT('h9)
	) name676 (
		\WX8575_reg/NET0131 ,
		\WX8639_reg/NET0131 ,
		_w2185_
	);
	LUT2 #(
		.INIT('h9)
	) name677 (
		\WX8447_reg/NET0131 ,
		\WX8511_reg/NET0131 ,
		_w2186_
	);
	LUT4 #(
		.INIT('h0a02)
	) name678 (
		RESET_pad,
		\TM0_pad ,
		\TM1_pad ,
		\_2246__reg/NET0131 ,
		_w2187_
	);
	LUT4 #(
		.INIT('hbe00)
	) name679 (
		\TM0_pad ,
		_w2185_,
		_w2186_,
		_w2187_,
		_w2188_
	);
	LUT2 #(
		.INIT('he)
	) name680 (
		_w2184_,
		_w2188_,
		_w2189_
	);
	LUT4 #(
		.INIT('h2772)
	) name681 (
		\TM0_pad ,
		\WX10853_reg/NET0131 ,
		_w1539_,
		_w1540_,
		_w2190_
	);
	LUT3 #(
		.INIT('h96)
	) name682 (
		\WX2026_reg/NET0131 ,
		\WX2090_reg/NET0131 ,
		\WX2154_reg/NET0131 ,
		_w2191_
	);
	LUT2 #(
		.INIT('h9)
	) name683 (
		\TM1_pad ,
		\WX1962_reg/NET0131 ,
		_w2192_
	);
	LUT4 #(
		.INIT('h2772)
	) name684 (
		\TM0_pad ,
		\_2096__reg/NET0131 ,
		_w2191_,
		_w2192_,
		_w2193_
	);
	LUT4 #(
		.INIT('h082a)
	) name685 (
		RESET_pad,
		\TM1_pad ,
		_w2190_,
		_w2193_,
		_w2194_
	);
	LUT3 #(
		.INIT('h96)
	) name686 (
		\WX11073_reg/NET0131 ,
		\WX11137_reg/NET0131 ,
		\WX11201_reg/NET0131 ,
		_w2195_
	);
	LUT2 #(
		.INIT('h9)
	) name687 (
		\TM1_pad ,
		\WX11009_reg/NET0131 ,
		_w2196_
	);
	LUT4 #(
		.INIT('h2772)
	) name688 (
		\TM0_pad ,
		\WX10849_reg/NET0131 ,
		_w2195_,
		_w2196_,
		_w2197_
	);
	LUT2 #(
		.INIT('h2)
	) name689 (
		\TM0_pad ,
		\_2354__reg/NET0131 ,
		_w2198_
	);
	LUT4 #(
		.INIT('h00c8)
	) name690 (
		\DATA_0_21_pad ,
		RESET_pad,
		\TM0_pad ,
		\TM1_pad ,
		_w2199_
	);
	LUT2 #(
		.INIT('h4)
	) name691 (
		_w2198_,
		_w2199_,
		_w2200_
	);
	LUT3 #(
		.INIT('hf2)
	) name692 (
		_w1605_,
		_w2197_,
		_w2200_,
		_w2201_
	);
	LUT2 #(
		.INIT('h8)
	) name693 (
		RESET_pad,
		\WX10847_reg/NET0131 ,
		_w2202_
	);
	LUT4 #(
		.INIT('ha020)
	) name694 (
		RESET_pad,
		\TM0_pad ,
		\TM1_pad ,
		\WX10881_reg/NET0131 ,
		_w2203_
	);
	LUT2 #(
		.INIT('h9)
	) name695 (
		\WX3411_reg/NET0131 ,
		\WX3475_reg/NET0131 ,
		_w2204_
	);
	LUT2 #(
		.INIT('h9)
	) name696 (
		\WX3283_reg/NET0131 ,
		\WX3347_reg/NET0131 ,
		_w2205_
	);
	LUT4 #(
		.INIT('h8cc8)
	) name697 (
		\TM0_pad ,
		_w2203_,
		_w2204_,
		_w2205_,
		_w2206_
	);
	LUT2 #(
		.INIT('h9)
	) name698 (
		\WX4704_reg/NET0131 ,
		\WX4768_reg/NET0131 ,
		_w2207_
	);
	LUT2 #(
		.INIT('h9)
	) name699 (
		\WX4576_reg/NET0131 ,
		\WX4640_reg/NET0131 ,
		_w2208_
	);
	LUT4 #(
		.INIT('h0a02)
	) name700 (
		RESET_pad,
		\TM0_pad ,
		\TM1_pad ,
		\_2146__reg/NET0131 ,
		_w2209_
	);
	LUT4 #(
		.INIT('hbe00)
	) name701 (
		\TM0_pad ,
		_w2207_,
		_w2208_,
		_w2209_,
		_w2210_
	);
	LUT2 #(
		.INIT('he)
	) name702 (
		_w2206_,
		_w2210_,
		_w2211_
	);
	LUT4 #(
		.INIT('h8cc8)
	) name703 (
		\TM0_pad ,
		_w1978_,
		_w2185_,
		_w2186_,
		_w2212_
	);
	LUT2 #(
		.INIT('h9)
	) name704 (
		\WX9868_reg/NET0131 ,
		\WX9932_reg/NET0131 ,
		_w2213_
	);
	LUT2 #(
		.INIT('h9)
	) name705 (
		\WX9740_reg/NET0131 ,
		\WX9804_reg/NET0131 ,
		_w2214_
	);
	LUT4 #(
		.INIT('h0a02)
	) name706 (
		RESET_pad,
		\TM0_pad ,
		\TM1_pad ,
		\_2278__reg/NET0131 ,
		_w2215_
	);
	LUT4 #(
		.INIT('hbe00)
	) name707 (
		\TM0_pad ,
		_w2213_,
		_w2214_,
		_w2215_,
		_w2216_
	);
	LUT2 #(
		.INIT('he)
	) name708 (
		_w2212_,
		_w2216_,
		_w2217_
	);
	LUT4 #(
		.INIT('h8cc8)
	) name709 (
		\TM0_pad ,
		_w1921_,
		_w2156_,
		_w2157_,
		_w2218_
	);
	LUT2 #(
		.INIT('h9)
	) name710 (
		\WX11159_reg/NET0131 ,
		\WX11223_reg/NET0131 ,
		_w2219_
	);
	LUT2 #(
		.INIT('h9)
	) name711 (
		\WX11031_reg/NET0131 ,
		\WX11095_reg/NET0131 ,
		_w2220_
	);
	LUT4 #(
		.INIT('h0a02)
	) name712 (
		RESET_pad,
		\TM0_pad ,
		\TM1_pad ,
		\_2311__reg/NET0131 ,
		_w2221_
	);
	LUT4 #(
		.INIT('hbe00)
	) name713 (
		\TM0_pad ,
		_w2219_,
		_w2220_,
		_w2221_,
		_w2222_
	);
	LUT2 #(
		.INIT('he)
	) name714 (
		_w2218_,
		_w2222_,
		_w2223_
	);
	LUT3 #(
		.INIT('h96)
	) name715 (
		\WX3317_reg/NET0131 ,
		\WX3381_reg/NET0131 ,
		\WX3445_reg/NET0131 ,
		_w2224_
	);
	LUT2 #(
		.INIT('h9)
	) name716 (
		\TM1_pad ,
		\WX3253_reg/NET0131 ,
		_w2225_
	);
	LUT4 #(
		.INIT('h2772)
	) name717 (
		\TM0_pad ,
		\_2129__reg/NET0131 ,
		_w2224_,
		_w2225_,
		_w2226_
	);
	LUT4 #(
		.INIT('h2772)
	) name718 (
		\TM0_pad ,
		\WX10851_reg/NET0131 ,
		_w2134_,
		_w2135_,
		_w2227_
	);
	LUT4 #(
		.INIT('h028a)
	) name719 (
		RESET_pad,
		\TM1_pad ,
		_w2226_,
		_w2227_,
		_w2228_
	);
	LUT4 #(
		.INIT('h8cc8)
	) name720 (
		\TM0_pad ,
		_w2146_,
		_w2150_,
		_w2151_,
		_w2229_
	);
	LUT2 #(
		.INIT('h9)
	) name721 (
		\WX5995_reg/NET0131 ,
		\WX6059_reg/NET0131 ,
		_w2230_
	);
	LUT2 #(
		.INIT('h9)
	) name722 (
		\WX5867_reg/NET0131 ,
		\WX5931_reg/NET0131 ,
		_w2231_
	);
	LUT4 #(
		.INIT('h0a02)
	) name723 (
		RESET_pad,
		\TM0_pad ,
		\TM1_pad ,
		\_2179__reg/NET0131 ,
		_w2232_
	);
	LUT4 #(
		.INIT('hbe00)
	) name724 (
		\TM0_pad ,
		_w2230_,
		_w2231_,
		_w2232_,
		_w2233_
	);
	LUT2 #(
		.INIT('he)
	) name725 (
		_w2229_,
		_w2233_,
		_w2234_
	);
	LUT4 #(
		.INIT('h8cc8)
	) name726 (
		\TM0_pad ,
		_w2089_,
		_w2173_,
		_w2174_,
		_w2235_
	);
	LUT2 #(
		.INIT('h9)
	) name727 (
		\WX7286_reg/NET0131 ,
		\WX7350_reg/NET0131 ,
		_w2236_
	);
	LUT2 #(
		.INIT('h9)
	) name728 (
		\WX7158_reg/NET0131 ,
		\WX7222_reg/NET0131 ,
		_w2237_
	);
	LUT4 #(
		.INIT('h0a02)
	) name729 (
		RESET_pad,
		\TM0_pad ,
		\TM1_pad ,
		\_2212__reg/NET0131 ,
		_w2238_
	);
	LUT4 #(
		.INIT('hbe00)
	) name730 (
		\TM0_pad ,
		_w2236_,
		_w2237_,
		_w2238_,
		_w2239_
	);
	LUT2 #(
		.INIT('he)
	) name731 (
		_w2235_,
		_w2239_,
		_w2240_
	);
	LUT4 #(
		.INIT('h8cc8)
	) name732 (
		\TM0_pad ,
		_w1620_,
		_w2179_,
		_w2180_,
		_w2241_
	);
	LUT2 #(
		.INIT('h9)
	) name733 (
		\WX8577_reg/NET0131 ,
		\WX8641_reg/NET0131 ,
		_w2242_
	);
	LUT2 #(
		.INIT('h9)
	) name734 (
		\WX8449_reg/NET0131 ,
		\WX8513_reg/NET0131 ,
		_w2243_
	);
	LUT4 #(
		.INIT('h0a02)
	) name735 (
		RESET_pad,
		\TM0_pad ,
		\TM1_pad ,
		\_2245__reg/NET0131 ,
		_w2244_
	);
	LUT4 #(
		.INIT('hbe00)
	) name736 (
		\TM0_pad ,
		_w2242_,
		_w2243_,
		_w2244_,
		_w2245_
	);
	LUT2 #(
		.INIT('he)
	) name737 (
		_w2241_,
		_w2245_,
		_w2246_
	);
	LUT4 #(
		.INIT('h2772)
	) name738 (
		\TM0_pad ,
		\WX10855_reg/NET0131 ,
		_w1536_,
		_w1537_,
		_w2247_
	);
	LUT3 #(
		.INIT('h96)
	) name739 (
		\WX2028_reg/NET0131 ,
		\WX2092_reg/NET0131 ,
		\WX2156_reg/NET0131 ,
		_w2248_
	);
	LUT2 #(
		.INIT('h9)
	) name740 (
		\TM1_pad ,
		\WX1964_reg/NET0131 ,
		_w2249_
	);
	LUT4 #(
		.INIT('h2772)
	) name741 (
		\TM0_pad ,
		\_2095__reg/NET0131 ,
		_w2248_,
		_w2249_,
		_w2250_
	);
	LUT4 #(
		.INIT('h082a)
	) name742 (
		RESET_pad,
		\TM1_pad ,
		_w2247_,
		_w2250_,
		_w2251_
	);
	LUT4 #(
		.INIT('h2772)
	) name743 (
		\TM0_pad ,
		\WX10851_reg/NET0131 ,
		_w1666_,
		_w1667_,
		_w2252_
	);
	LUT2 #(
		.INIT('h2)
	) name744 (
		\TM0_pad ,
		\_2353__reg/NET0131 ,
		_w2253_
	);
	LUT4 #(
		.INIT('h00c8)
	) name745 (
		\DATA_0_20_pad ,
		RESET_pad,
		\TM0_pad ,
		\TM1_pad ,
		_w2254_
	);
	LUT2 #(
		.INIT('h4)
	) name746 (
		_w2253_,
		_w2254_,
		_w2255_
	);
	LUT3 #(
		.INIT('hf2)
	) name747 (
		_w1605_,
		_w2252_,
		_w2255_,
		_w2256_
	);
	LUT2 #(
		.INIT('h8)
	) name748 (
		RESET_pad,
		\WX10849_reg/NET0131 ,
		_w2257_
	);
	LUT4 #(
		.INIT('ha020)
	) name749 (
		RESET_pad,
		\TM0_pad ,
		\TM1_pad ,
		\WX10883_reg/NET0131 ,
		_w2258_
	);
	LUT2 #(
		.INIT('h9)
	) name750 (
		\WX3413_reg/NET0131 ,
		\WX3477_reg/NET0131 ,
		_w2259_
	);
	LUT2 #(
		.INIT('h9)
	) name751 (
		\WX3285_reg/NET0131 ,
		\WX3349_reg/NET0131 ,
		_w2260_
	);
	LUT4 #(
		.INIT('h8cc8)
	) name752 (
		\TM0_pad ,
		_w2258_,
		_w2259_,
		_w2260_,
		_w2261_
	);
	LUT2 #(
		.INIT('h9)
	) name753 (
		\WX4706_reg/NET0131 ,
		\WX4770_reg/NET0131 ,
		_w2262_
	);
	LUT2 #(
		.INIT('h9)
	) name754 (
		\WX4578_reg/NET0131 ,
		\WX4642_reg/NET0131 ,
		_w2263_
	);
	LUT4 #(
		.INIT('h0a02)
	) name755 (
		RESET_pad,
		\TM0_pad ,
		\TM1_pad ,
		\_2145__reg/NET0131 ,
		_w2264_
	);
	LUT4 #(
		.INIT('hbe00)
	) name756 (
		\TM0_pad ,
		_w2262_,
		_w2263_,
		_w2264_,
		_w2265_
	);
	LUT2 #(
		.INIT('he)
	) name757 (
		_w2261_,
		_w2265_,
		_w2266_
	);
	LUT4 #(
		.INIT('h8cc8)
	) name758 (
		\TM0_pad ,
		_w1620_,
		_w2242_,
		_w2243_,
		_w2267_
	);
	LUT2 #(
		.INIT('h9)
	) name759 (
		\WX9870_reg/NET0131 ,
		\WX9934_reg/NET0131 ,
		_w2268_
	);
	LUT2 #(
		.INIT('h9)
	) name760 (
		\WX9742_reg/NET0131 ,
		\WX9806_reg/NET0131 ,
		_w2269_
	);
	LUT4 #(
		.INIT('h0a02)
	) name761 (
		RESET_pad,
		\TM0_pad ,
		\TM1_pad ,
		\_2277__reg/NET0131 ,
		_w2270_
	);
	LUT4 #(
		.INIT('hbe00)
	) name762 (
		\TM0_pad ,
		_w2268_,
		_w2269_,
		_w2270_,
		_w2271_
	);
	LUT2 #(
		.INIT('he)
	) name763 (
		_w2267_,
		_w2271_,
		_w2272_
	);
	LUT4 #(
		.INIT('h8cc8)
	) name764 (
		\TM0_pad ,
		_w1978_,
		_w2213_,
		_w2214_,
		_w2273_
	);
	LUT2 #(
		.INIT('h9)
	) name765 (
		\WX11161_reg/NET0131 ,
		\WX11225_reg/NET0131 ,
		_w2274_
	);
	LUT2 #(
		.INIT('h9)
	) name766 (
		\WX11033_reg/NET0131 ,
		\WX11097_reg/NET0131 ,
		_w2275_
	);
	LUT4 #(
		.INIT('h0a02)
	) name767 (
		RESET_pad,
		\TM0_pad ,
		\TM1_pad ,
		\_2310__reg/NET0131 ,
		_w2276_
	);
	LUT4 #(
		.INIT('hbe00)
	) name768 (
		\TM0_pad ,
		_w2274_,
		_w2275_,
		_w2276_,
		_w2277_
	);
	LUT2 #(
		.INIT('he)
	) name769 (
		_w2273_,
		_w2277_,
		_w2278_
	);
	LUT3 #(
		.INIT('h96)
	) name770 (
		\WX3319_reg/NET0131 ,
		\WX3383_reg/NET0131 ,
		\WX3447_reg/NET0131 ,
		_w2279_
	);
	LUT2 #(
		.INIT('h9)
	) name771 (
		\TM1_pad ,
		\WX3255_reg/NET0131 ,
		_w2280_
	);
	LUT4 #(
		.INIT('h2772)
	) name772 (
		\TM0_pad ,
		\_2128__reg/NET0131 ,
		_w2279_,
		_w2280_,
		_w2281_
	);
	LUT4 #(
		.INIT('h2772)
	) name773 (
		\TM0_pad ,
		\WX10853_reg/NET0131 ,
		_w2191_,
		_w2192_,
		_w2282_
	);
	LUT4 #(
		.INIT('h028a)
	) name774 (
		RESET_pad,
		\TM1_pad ,
		_w2281_,
		_w2282_,
		_w2283_
	);
	LUT4 #(
		.INIT('h8cc8)
	) name775 (
		\TM0_pad ,
		_w2203_,
		_w2207_,
		_w2208_,
		_w2284_
	);
	LUT2 #(
		.INIT('h9)
	) name776 (
		\WX5997_reg/NET0131 ,
		\WX6061_reg/NET0131 ,
		_w2285_
	);
	LUT2 #(
		.INIT('h9)
	) name777 (
		\WX5869_reg/NET0131 ,
		\WX5933_reg/NET0131 ,
		_w2286_
	);
	LUT4 #(
		.INIT('h0a02)
	) name778 (
		RESET_pad,
		\TM0_pad ,
		\TM1_pad ,
		\_2178__reg/NET0131 ,
		_w2287_
	);
	LUT4 #(
		.INIT('hbe00)
	) name779 (
		\TM0_pad ,
		_w2285_,
		_w2286_,
		_w2287_,
		_w2288_
	);
	LUT2 #(
		.INIT('he)
	) name780 (
		_w2284_,
		_w2288_,
		_w2289_
	);
	LUT4 #(
		.INIT('h8cc8)
	) name781 (
		\TM0_pad ,
		_w2146_,
		_w2230_,
		_w2231_,
		_w2290_
	);
	LUT2 #(
		.INIT('h9)
	) name782 (
		\WX7288_reg/NET0131 ,
		\WX7352_reg/NET0131 ,
		_w2291_
	);
	LUT2 #(
		.INIT('h9)
	) name783 (
		\WX7160_reg/NET0131 ,
		\WX7224_reg/NET0131 ,
		_w2292_
	);
	LUT4 #(
		.INIT('h0a02)
	) name784 (
		RESET_pad,
		\TM0_pad ,
		\TM1_pad ,
		\_2211__reg/NET0131 ,
		_w2293_
	);
	LUT4 #(
		.INIT('hbe00)
	) name785 (
		\TM0_pad ,
		_w2291_,
		_w2292_,
		_w2293_,
		_w2294_
	);
	LUT2 #(
		.INIT('he)
	) name786 (
		_w2290_,
		_w2294_,
		_w2295_
	);
	LUT4 #(
		.INIT('h8cc8)
	) name787 (
		\TM0_pad ,
		_w2089_,
		_w2236_,
		_w2237_,
		_w2296_
	);
	LUT2 #(
		.INIT('h9)
	) name788 (
		\WX8579_reg/NET0131 ,
		\WX8643_reg/NET0131 ,
		_w2297_
	);
	LUT2 #(
		.INIT('h9)
	) name789 (
		\WX8451_reg/NET0131 ,
		\WX8515_reg/NET0131 ,
		_w2298_
	);
	LUT4 #(
		.INIT('h0a02)
	) name790 (
		RESET_pad,
		\TM0_pad ,
		\TM1_pad ,
		\_2244__reg/NET0131 ,
		_w2299_
	);
	LUT4 #(
		.INIT('hbe00)
	) name791 (
		\TM0_pad ,
		_w2297_,
		_w2298_,
		_w2299_,
		_w2300_
	);
	LUT2 #(
		.INIT('he)
	) name792 (
		_w2296_,
		_w2300_,
		_w2301_
	);
	LUT3 #(
		.INIT('h96)
	) name793 (
		\WX2030_reg/NET0131 ,
		\WX2094_reg/NET0131 ,
		\WX2158_reg/NET0131 ,
		_w2302_
	);
	LUT2 #(
		.INIT('h9)
	) name794 (
		\TM1_pad ,
		\WX1966_reg/NET0131 ,
		_w2303_
	);
	LUT4 #(
		.INIT('h2772)
	) name795 (
		\TM0_pad ,
		\_2094__reg/NET0131 ,
		_w2302_,
		_w2303_,
		_w2304_
	);
	LUT4 #(
		.INIT('h2772)
	) name796 (
		\TM0_pad ,
		\WX10857_reg/NET0131 ,
		_w1533_,
		_w1534_,
		_w2305_
	);
	LUT4 #(
		.INIT('h028a)
	) name797 (
		RESET_pad,
		\TM1_pad ,
		_w2304_,
		_w2305_,
		_w2306_
	);
	LUT4 #(
		.INIT('h2772)
	) name798 (
		\TM0_pad ,
		\WX10853_reg/NET0131 ,
		_w1725_,
		_w1726_,
		_w2307_
	);
	LUT2 #(
		.INIT('h2)
	) name799 (
		\TM0_pad ,
		\_2352__reg/NET0131 ,
		_w2308_
	);
	LUT4 #(
		.INIT('h00c8)
	) name800 (
		\DATA_0_19_pad ,
		RESET_pad,
		\TM0_pad ,
		\TM1_pad ,
		_w2309_
	);
	LUT2 #(
		.INIT('h4)
	) name801 (
		_w2308_,
		_w2309_,
		_w2310_
	);
	LUT3 #(
		.INIT('hf2)
	) name802 (
		_w1605_,
		_w2307_,
		_w2310_,
		_w2311_
	);
	LUT2 #(
		.INIT('h8)
	) name803 (
		RESET_pad,
		\WX10851_reg/NET0131 ,
		_w2312_
	);
	LUT4 #(
		.INIT('ha020)
	) name804 (
		RESET_pad,
		\TM0_pad ,
		\TM1_pad ,
		\WX10885_reg/NET0131 ,
		_w2313_
	);
	LUT2 #(
		.INIT('h9)
	) name805 (
		\WX3415_reg/NET0131 ,
		\WX3479_reg/NET0131 ,
		_w2314_
	);
	LUT2 #(
		.INIT('h9)
	) name806 (
		\WX3287_reg/NET0131 ,
		\WX3351_reg/NET0131 ,
		_w2315_
	);
	LUT4 #(
		.INIT('h8cc8)
	) name807 (
		\TM0_pad ,
		_w2313_,
		_w2314_,
		_w2315_,
		_w2316_
	);
	LUT2 #(
		.INIT('h9)
	) name808 (
		\WX4708_reg/NET0131 ,
		\WX4772_reg/NET0131 ,
		_w2317_
	);
	LUT2 #(
		.INIT('h9)
	) name809 (
		\WX4580_reg/NET0131 ,
		\WX4644_reg/NET0131 ,
		_w2318_
	);
	LUT4 #(
		.INIT('h0a02)
	) name810 (
		RESET_pad,
		\TM0_pad ,
		\TM1_pad ,
		\_2144__reg/NET0131 ,
		_w2319_
	);
	LUT4 #(
		.INIT('hbe00)
	) name811 (
		\TM0_pad ,
		_w2317_,
		_w2318_,
		_w2319_,
		_w2320_
	);
	LUT2 #(
		.INIT('he)
	) name812 (
		_w2316_,
		_w2320_,
		_w2321_
	);
	LUT4 #(
		.INIT('h8cc8)
	) name813 (
		\TM0_pad ,
		_w2089_,
		_w2297_,
		_w2298_,
		_w2322_
	);
	LUT2 #(
		.INIT('h9)
	) name814 (
		\WX9872_reg/NET0131 ,
		\WX9936_reg/NET0131 ,
		_w2323_
	);
	LUT2 #(
		.INIT('h9)
	) name815 (
		\WX9744_reg/NET0131 ,
		\WX9808_reg/NET0131 ,
		_w2324_
	);
	LUT4 #(
		.INIT('h0a02)
	) name816 (
		RESET_pad,
		\TM0_pad ,
		\TM1_pad ,
		\_2276__reg/NET0131 ,
		_w2325_
	);
	LUT4 #(
		.INIT('hbe00)
	) name817 (
		\TM0_pad ,
		_w2323_,
		_w2324_,
		_w2325_,
		_w2326_
	);
	LUT2 #(
		.INIT('he)
	) name818 (
		_w2322_,
		_w2326_,
		_w2327_
	);
	LUT4 #(
		.INIT('h8cc8)
	) name819 (
		\TM0_pad ,
		_w1620_,
		_w2268_,
		_w2269_,
		_w2328_
	);
	LUT4 #(
		.INIT('h0a02)
	) name820 (
		RESET_pad,
		\TM0_pad ,
		\TM1_pad ,
		\_2309__reg/NET0131 ,
		_w2329_
	);
	LUT4 #(
		.INIT('hbe00)
	) name821 (
		\TM0_pad ,
		_w1621_,
		_w1622_,
		_w2329_,
		_w2330_
	);
	LUT2 #(
		.INIT('he)
	) name822 (
		_w2328_,
		_w2330_,
		_w2331_
	);
	LUT3 #(
		.INIT('h96)
	) name823 (
		\WX3321_reg/NET0131 ,
		\WX3385_reg/NET0131 ,
		\WX3449_reg/NET0131 ,
		_w2332_
	);
	LUT2 #(
		.INIT('h9)
	) name824 (
		\TM1_pad ,
		\WX3257_reg/NET0131 ,
		_w2333_
	);
	LUT4 #(
		.INIT('h2772)
	) name825 (
		\TM0_pad ,
		\_2127__reg/NET0131 ,
		_w2332_,
		_w2333_,
		_w2334_
	);
	LUT4 #(
		.INIT('h2772)
	) name826 (
		\TM0_pad ,
		\WX10855_reg/NET0131 ,
		_w2248_,
		_w2249_,
		_w2335_
	);
	LUT4 #(
		.INIT('h028a)
	) name827 (
		RESET_pad,
		\TM1_pad ,
		_w2334_,
		_w2335_,
		_w2336_
	);
	LUT4 #(
		.INIT('h8cc8)
	) name828 (
		\TM0_pad ,
		_w2258_,
		_w2262_,
		_w2263_,
		_w2337_
	);
	LUT2 #(
		.INIT('h9)
	) name829 (
		\WX5999_reg/NET0131 ,
		\WX6063_reg/NET0131 ,
		_w2338_
	);
	LUT2 #(
		.INIT('h9)
	) name830 (
		\WX5871_reg/NET0131 ,
		\WX5935_reg/NET0131 ,
		_w2339_
	);
	LUT4 #(
		.INIT('h0a02)
	) name831 (
		RESET_pad,
		\TM0_pad ,
		\TM1_pad ,
		\_2177__reg/NET0131 ,
		_w2340_
	);
	LUT4 #(
		.INIT('hbe00)
	) name832 (
		\TM0_pad ,
		_w2338_,
		_w2339_,
		_w2340_,
		_w2341_
	);
	LUT2 #(
		.INIT('he)
	) name833 (
		_w2337_,
		_w2341_,
		_w2342_
	);
	LUT4 #(
		.INIT('h8cc8)
	) name834 (
		\TM0_pad ,
		_w2203_,
		_w2285_,
		_w2286_,
		_w2343_
	);
	LUT2 #(
		.INIT('h9)
	) name835 (
		\WX7290_reg/NET0131 ,
		\WX7354_reg/NET0131 ,
		_w2344_
	);
	LUT2 #(
		.INIT('h9)
	) name836 (
		\WX7162_reg/NET0131 ,
		\WX7226_reg/NET0131 ,
		_w2345_
	);
	LUT4 #(
		.INIT('h0a02)
	) name837 (
		RESET_pad,
		\TM0_pad ,
		\TM1_pad ,
		\_2210__reg/NET0131 ,
		_w2346_
	);
	LUT4 #(
		.INIT('hbe00)
	) name838 (
		\TM0_pad ,
		_w2344_,
		_w2345_,
		_w2346_,
		_w2347_
	);
	LUT2 #(
		.INIT('he)
	) name839 (
		_w2343_,
		_w2347_,
		_w2348_
	);
	LUT4 #(
		.INIT('h8cc8)
	) name840 (
		\TM0_pad ,
		_w2146_,
		_w2291_,
		_w2292_,
		_w2349_
	);
	LUT2 #(
		.INIT('h9)
	) name841 (
		\WX8581_reg/NET0131 ,
		\WX8645_reg/NET0131 ,
		_w2350_
	);
	LUT2 #(
		.INIT('h9)
	) name842 (
		\WX8453_reg/NET0131 ,
		\WX8517_reg/NET0131 ,
		_w2351_
	);
	LUT4 #(
		.INIT('h0a02)
	) name843 (
		RESET_pad,
		\TM0_pad ,
		\TM1_pad ,
		\_2243__reg/NET0131 ,
		_w2352_
	);
	LUT4 #(
		.INIT('hbe00)
	) name844 (
		\TM0_pad ,
		_w2350_,
		_w2351_,
		_w2352_,
		_w2353_
	);
	LUT2 #(
		.INIT('he)
	) name845 (
		_w2349_,
		_w2353_,
		_w2354_
	);
	LUT4 #(
		.INIT('h2772)
	) name846 (
		\TM0_pad ,
		\WX10859_reg/NET0131 ,
		_w1530_,
		_w1531_,
		_w2355_
	);
	LUT3 #(
		.INIT('h96)
	) name847 (
		\WX2032_reg/NET0131 ,
		\WX2096_reg/NET0131 ,
		\WX2160_reg/NET0131 ,
		_w2356_
	);
	LUT2 #(
		.INIT('h9)
	) name848 (
		\TM1_pad ,
		\WX1968_reg/NET0131 ,
		_w2357_
	);
	LUT4 #(
		.INIT('h2772)
	) name849 (
		\TM0_pad ,
		\_2093__reg/NET0131 ,
		_w2356_,
		_w2357_,
		_w2358_
	);
	LUT4 #(
		.INIT('h082a)
	) name850 (
		RESET_pad,
		\TM1_pad ,
		_w2355_,
		_w2358_,
		_w2359_
	);
	LUT4 #(
		.INIT('h2772)
	) name851 (
		\TM0_pad ,
		\WX10855_reg/NET0131 ,
		_w1777_,
		_w1778_,
		_w2360_
	);
	LUT2 #(
		.INIT('h2)
	) name852 (
		\TM0_pad ,
		\_2351__reg/NET0131 ,
		_w2361_
	);
	LUT4 #(
		.INIT('h00c8)
	) name853 (
		\DATA_0_18_pad ,
		RESET_pad,
		\TM0_pad ,
		\TM1_pad ,
		_w2362_
	);
	LUT2 #(
		.INIT('h4)
	) name854 (
		_w2361_,
		_w2362_,
		_w2363_
	);
	LUT3 #(
		.INIT('hf2)
	) name855 (
		_w1605_,
		_w2360_,
		_w2363_,
		_w2364_
	);
	LUT2 #(
		.INIT('h8)
	) name856 (
		RESET_pad,
		\WX10853_reg/NET0131 ,
		_w2365_
	);
	LUT4 #(
		.INIT('ha020)
	) name857 (
		RESET_pad,
		\TM0_pad ,
		\TM1_pad ,
		\WX10887_reg/NET0131 ,
		_w2366_
	);
	LUT2 #(
		.INIT('h9)
	) name858 (
		\WX3417_reg/NET0131 ,
		\WX3481_reg/NET0131 ,
		_w2367_
	);
	LUT2 #(
		.INIT('h9)
	) name859 (
		\WX3289_reg/NET0131 ,
		\WX3353_reg/NET0131 ,
		_w2368_
	);
	LUT4 #(
		.INIT('h8cc8)
	) name860 (
		\TM0_pad ,
		_w2366_,
		_w2367_,
		_w2368_,
		_w2369_
	);
	LUT2 #(
		.INIT('h9)
	) name861 (
		\WX4710_reg/NET0131 ,
		\WX4774_reg/NET0131 ,
		_w2370_
	);
	LUT2 #(
		.INIT('h9)
	) name862 (
		\WX4582_reg/NET0131 ,
		\WX4646_reg/NET0131 ,
		_w2371_
	);
	LUT4 #(
		.INIT('h0a02)
	) name863 (
		RESET_pad,
		\TM0_pad ,
		\TM1_pad ,
		\_2143__reg/NET0131 ,
		_w2372_
	);
	LUT4 #(
		.INIT('hbe00)
	) name864 (
		\TM0_pad ,
		_w2370_,
		_w2371_,
		_w2372_,
		_w2373_
	);
	LUT2 #(
		.INIT('he)
	) name865 (
		_w2369_,
		_w2373_,
		_w2374_
	);
	LUT4 #(
		.INIT('h8cc8)
	) name866 (
		\TM0_pad ,
		_w2146_,
		_w2350_,
		_w2351_,
		_w2375_
	);
	LUT2 #(
		.INIT('h9)
	) name867 (
		\WX9874_reg/NET0131 ,
		\WX9938_reg/NET0131 ,
		_w2376_
	);
	LUT2 #(
		.INIT('h9)
	) name868 (
		\WX9746_reg/NET0131 ,
		\WX9810_reg/NET0131 ,
		_w2377_
	);
	LUT4 #(
		.INIT('h0a02)
	) name869 (
		RESET_pad,
		\TM0_pad ,
		\TM1_pad ,
		\_2275__reg/NET0131 ,
		_w2378_
	);
	LUT4 #(
		.INIT('hbe00)
	) name870 (
		\TM0_pad ,
		_w2376_,
		_w2377_,
		_w2378_,
		_w2379_
	);
	LUT2 #(
		.INIT('he)
	) name871 (
		_w2375_,
		_w2379_,
		_w2380_
	);
	LUT4 #(
		.INIT('h8cc8)
	) name872 (
		\TM0_pad ,
		_w2089_,
		_w2323_,
		_w2324_,
		_w2381_
	);
	LUT2 #(
		.INIT('h9)
	) name873 (
		\WX11165_reg/NET0131 ,
		\WX11229_reg/NET0131 ,
		_w2382_
	);
	LUT2 #(
		.INIT('h9)
	) name874 (
		\WX11037_reg/NET0131 ,
		\WX11101_reg/NET0131 ,
		_w2383_
	);
	LUT4 #(
		.INIT('h0a02)
	) name875 (
		RESET_pad,
		\TM0_pad ,
		\TM1_pad ,
		\_2308__reg/NET0131 ,
		_w2384_
	);
	LUT4 #(
		.INIT('hbe00)
	) name876 (
		\TM0_pad ,
		_w2382_,
		_w2383_,
		_w2384_,
		_w2385_
	);
	LUT2 #(
		.INIT('he)
	) name877 (
		_w2381_,
		_w2385_,
		_w2386_
	);
	LUT4 #(
		.INIT('h8cc8)
	) name878 (
		\TM0_pad ,
		_w2313_,
		_w2317_,
		_w2318_,
		_w2387_
	);
	LUT2 #(
		.INIT('h9)
	) name879 (
		\WX6001_reg/NET0131 ,
		\WX6065_reg/NET0131 ,
		_w2388_
	);
	LUT2 #(
		.INIT('h9)
	) name880 (
		\WX5873_reg/NET0131 ,
		\WX5937_reg/NET0131 ,
		_w2389_
	);
	LUT4 #(
		.INIT('h0a02)
	) name881 (
		RESET_pad,
		\TM0_pad ,
		\TM1_pad ,
		\_2176__reg/NET0131 ,
		_w2390_
	);
	LUT4 #(
		.INIT('hbe00)
	) name882 (
		\TM0_pad ,
		_w2388_,
		_w2389_,
		_w2390_,
		_w2391_
	);
	LUT2 #(
		.INIT('he)
	) name883 (
		_w2387_,
		_w2391_,
		_w2392_
	);
	LUT3 #(
		.INIT('h96)
	) name884 (
		\WX3323_reg/NET0131 ,
		\WX3387_reg/NET0131 ,
		\WX3451_reg/NET0131 ,
		_w2393_
	);
	LUT2 #(
		.INIT('h9)
	) name885 (
		\TM1_pad ,
		\WX3259_reg/NET0131 ,
		_w2394_
	);
	LUT4 #(
		.INIT('h2772)
	) name886 (
		\TM0_pad ,
		\_2126__reg/NET0131 ,
		_w2393_,
		_w2394_,
		_w2395_
	);
	LUT4 #(
		.INIT('h2772)
	) name887 (
		\TM0_pad ,
		\WX10857_reg/NET0131 ,
		_w2302_,
		_w2303_,
		_w2396_
	);
	LUT4 #(
		.INIT('h028a)
	) name888 (
		RESET_pad,
		\TM1_pad ,
		_w2395_,
		_w2396_,
		_w2397_
	);
	LUT4 #(
		.INIT('h8cc8)
	) name889 (
		\TM0_pad ,
		_w2258_,
		_w2338_,
		_w2339_,
		_w2398_
	);
	LUT2 #(
		.INIT('h9)
	) name890 (
		\WX7292_reg/NET0131 ,
		\WX7356_reg/NET0131 ,
		_w2399_
	);
	LUT2 #(
		.INIT('h9)
	) name891 (
		\WX7164_reg/NET0131 ,
		\WX7228_reg/NET0131 ,
		_w2400_
	);
	LUT4 #(
		.INIT('h0a02)
	) name892 (
		RESET_pad,
		\TM0_pad ,
		\TM1_pad ,
		\_2209__reg/NET0131 ,
		_w2401_
	);
	LUT4 #(
		.INIT('hbe00)
	) name893 (
		\TM0_pad ,
		_w2399_,
		_w2400_,
		_w2401_,
		_w2402_
	);
	LUT2 #(
		.INIT('he)
	) name894 (
		_w2398_,
		_w2402_,
		_w2403_
	);
	LUT4 #(
		.INIT('h8cc8)
	) name895 (
		\TM0_pad ,
		_w2203_,
		_w2344_,
		_w2345_,
		_w2404_
	);
	LUT2 #(
		.INIT('h9)
	) name896 (
		\WX8583_reg/NET0131 ,
		\WX8647_reg/NET0131 ,
		_w2405_
	);
	LUT2 #(
		.INIT('h9)
	) name897 (
		\WX8455_reg/NET0131 ,
		\WX8519_reg/NET0131 ,
		_w2406_
	);
	LUT4 #(
		.INIT('h0a02)
	) name898 (
		RESET_pad,
		\TM0_pad ,
		\TM1_pad ,
		\_2242__reg/NET0131 ,
		_w2407_
	);
	LUT4 #(
		.INIT('hbe00)
	) name899 (
		\TM0_pad ,
		_w2405_,
		_w2406_,
		_w2407_,
		_w2408_
	);
	LUT2 #(
		.INIT('he)
	) name900 (
		_w2404_,
		_w2408_,
		_w2409_
	);
	LUT4 #(
		.INIT('h2772)
	) name901 (
		\TM0_pad ,
		\WX10857_reg/NET0131 ,
		_w1829_,
		_w1830_,
		_w2410_
	);
	LUT2 #(
		.INIT('h2)
	) name902 (
		\TM0_pad ,
		\_2350__reg/NET0131 ,
		_w2411_
	);
	LUT4 #(
		.INIT('h00c8)
	) name903 (
		\DATA_0_17_pad ,
		RESET_pad,
		\TM0_pad ,
		\TM1_pad ,
		_w2412_
	);
	LUT2 #(
		.INIT('h4)
	) name904 (
		_w2411_,
		_w2412_,
		_w2413_
	);
	LUT3 #(
		.INIT('hf2)
	) name905 (
		_w1605_,
		_w2410_,
		_w2413_,
		_w2414_
	);
	LUT2 #(
		.INIT('h8)
	) name906 (
		RESET_pad,
		\WX10855_reg/NET0131 ,
		_w2415_
	);
	LUT4 #(
		.INIT('h8cc8)
	) name907 (
		\TM0_pad ,
		_w2258_,
		_w2399_,
		_w2400_,
		_w2416_
	);
	LUT2 #(
		.INIT('h9)
	) name908 (
		\WX8585_reg/NET0131 ,
		\WX8649_reg/NET0131 ,
		_w2417_
	);
	LUT2 #(
		.INIT('h9)
	) name909 (
		\WX8457_reg/NET0131 ,
		\WX8521_reg/NET0131 ,
		_w2418_
	);
	LUT4 #(
		.INIT('h0a02)
	) name910 (
		RESET_pad,
		\TM0_pad ,
		\TM1_pad ,
		\_2241__reg/NET0131 ,
		_w2419_
	);
	LUT4 #(
		.INIT('hbe00)
	) name911 (
		\TM0_pad ,
		_w2417_,
		_w2418_,
		_w2419_,
		_w2420_
	);
	LUT2 #(
		.INIT('he)
	) name912 (
		_w2416_,
		_w2420_,
		_w2421_
	);
	LUT4 #(
		.INIT('ha020)
	) name913 (
		RESET_pad,
		\TM0_pad ,
		\TM1_pad ,
		\WX10889_reg/NET0131 ,
		_w2422_
	);
	LUT2 #(
		.INIT('h9)
	) name914 (
		\WX3419_reg/NET0131 ,
		\WX3483_reg/NET0131 ,
		_w2423_
	);
	LUT2 #(
		.INIT('h9)
	) name915 (
		\WX3291_reg/NET0131 ,
		\WX3355_reg/NET0131 ,
		_w2424_
	);
	LUT4 #(
		.INIT('h8cc8)
	) name916 (
		\TM0_pad ,
		_w2422_,
		_w2423_,
		_w2424_,
		_w2425_
	);
	LUT2 #(
		.INIT('h9)
	) name917 (
		\WX4712_reg/NET0131 ,
		\WX4776_reg/NET0131 ,
		_w2426_
	);
	LUT2 #(
		.INIT('h9)
	) name918 (
		\WX4584_reg/NET0131 ,
		\WX4648_reg/NET0131 ,
		_w2427_
	);
	LUT4 #(
		.INIT('h0a02)
	) name919 (
		RESET_pad,
		\TM0_pad ,
		\TM1_pad ,
		\_2142__reg/NET0131 ,
		_w2428_
	);
	LUT4 #(
		.INIT('hbe00)
	) name920 (
		\TM0_pad ,
		_w2426_,
		_w2427_,
		_w2428_,
		_w2429_
	);
	LUT2 #(
		.INIT('he)
	) name921 (
		_w2425_,
		_w2429_,
		_w2430_
	);
	LUT4 #(
		.INIT('h8cc8)
	) name922 (
		\TM0_pad ,
		_w2203_,
		_w2405_,
		_w2406_,
		_w2431_
	);
	LUT2 #(
		.INIT('h9)
	) name923 (
		\WX9876_reg/NET0131 ,
		\WX9940_reg/NET0131 ,
		_w2432_
	);
	LUT2 #(
		.INIT('h9)
	) name924 (
		\WX9748_reg/NET0131 ,
		\WX9812_reg/NET0131 ,
		_w2433_
	);
	LUT4 #(
		.INIT('h0a02)
	) name925 (
		RESET_pad,
		\TM0_pad ,
		\TM1_pad ,
		\_2274__reg/NET0131 ,
		_w2434_
	);
	LUT4 #(
		.INIT('hbe00)
	) name926 (
		\TM0_pad ,
		_w2432_,
		_w2433_,
		_w2434_,
		_w2435_
	);
	LUT2 #(
		.INIT('he)
	) name927 (
		_w2431_,
		_w2435_,
		_w2436_
	);
	LUT4 #(
		.INIT('h8cc8)
	) name928 (
		\TM0_pad ,
		_w2146_,
		_w2376_,
		_w2377_,
		_w2437_
	);
	LUT2 #(
		.INIT('h9)
	) name929 (
		\WX11167_reg/NET0131 ,
		\WX11231_reg/NET0131 ,
		_w2438_
	);
	LUT2 #(
		.INIT('h9)
	) name930 (
		\WX11039_reg/NET0131 ,
		\WX11103_reg/NET0131 ,
		_w2439_
	);
	LUT4 #(
		.INIT('h0a02)
	) name931 (
		RESET_pad,
		\TM0_pad ,
		\TM1_pad ,
		\_2307__reg/NET0131 ,
		_w2440_
	);
	LUT4 #(
		.INIT('hbe00)
	) name932 (
		\TM0_pad ,
		_w2438_,
		_w2439_,
		_w2440_,
		_w2441_
	);
	LUT2 #(
		.INIT('he)
	) name933 (
		_w2437_,
		_w2441_,
		_w2442_
	);
	LUT4 #(
		.INIT('h8cc8)
	) name934 (
		\TM0_pad ,
		_w2366_,
		_w2370_,
		_w2371_,
		_w2443_
	);
	LUT2 #(
		.INIT('h9)
	) name935 (
		\WX6003_reg/NET0131 ,
		\WX6067_reg/NET0131 ,
		_w2444_
	);
	LUT2 #(
		.INIT('h9)
	) name936 (
		\WX5875_reg/NET0131 ,
		\WX5939_reg/NET0131 ,
		_w2445_
	);
	LUT4 #(
		.INIT('h0a02)
	) name937 (
		RESET_pad,
		\TM0_pad ,
		\TM1_pad ,
		\_2175__reg/NET0131 ,
		_w2446_
	);
	LUT4 #(
		.INIT('hbe00)
	) name938 (
		\TM0_pad ,
		_w2444_,
		_w2445_,
		_w2446_,
		_w2447_
	);
	LUT2 #(
		.INIT('he)
	) name939 (
		_w2443_,
		_w2447_,
		_w2448_
	);
	LUT3 #(
		.INIT('h96)
	) name940 (
		\WX3325_reg/NET0131 ,
		\WX3389_reg/NET0131 ,
		\WX3453_reg/NET0131 ,
		_w2449_
	);
	LUT2 #(
		.INIT('h9)
	) name941 (
		\TM1_pad ,
		\WX3261_reg/NET0131 ,
		_w2450_
	);
	LUT4 #(
		.INIT('h2772)
	) name942 (
		\TM0_pad ,
		\_2125__reg/NET0131 ,
		_w2449_,
		_w2450_,
		_w2451_
	);
	LUT4 #(
		.INIT('h2772)
	) name943 (
		\TM0_pad ,
		\WX10859_reg/NET0131 ,
		_w2356_,
		_w2357_,
		_w2452_
	);
	LUT4 #(
		.INIT('h028a)
	) name944 (
		RESET_pad,
		\TM1_pad ,
		_w2451_,
		_w2452_,
		_w2453_
	);
	LUT4 #(
		.INIT('h8cc8)
	) name945 (
		\TM0_pad ,
		_w2313_,
		_w2388_,
		_w2389_,
		_w2454_
	);
	LUT2 #(
		.INIT('h9)
	) name946 (
		\WX7294_reg/NET0131 ,
		\WX7358_reg/NET0131 ,
		_w2455_
	);
	LUT2 #(
		.INIT('h9)
	) name947 (
		\WX7166_reg/NET0131 ,
		\WX7230_reg/NET0131 ,
		_w2456_
	);
	LUT4 #(
		.INIT('h0a02)
	) name948 (
		RESET_pad,
		\TM0_pad ,
		\TM1_pad ,
		\_2208__reg/NET0131 ,
		_w2457_
	);
	LUT4 #(
		.INIT('hbe00)
	) name949 (
		\TM0_pad ,
		_w2455_,
		_w2456_,
		_w2457_,
		_w2458_
	);
	LUT2 #(
		.INIT('he)
	) name950 (
		_w2454_,
		_w2458_,
		_w2459_
	);
	LUT4 #(
		.INIT('h2772)
	) name951 (
		\TM0_pad ,
		\WX10859_reg/NET0131 ,
		_w1885_,
		_w1886_,
		_w2460_
	);
	LUT2 #(
		.INIT('h2)
	) name952 (
		\TM0_pad ,
		\_2349__reg/NET0131 ,
		_w2461_
	);
	LUT4 #(
		.INIT('h00c8)
	) name953 (
		\DATA_0_16_pad ,
		RESET_pad,
		\TM0_pad ,
		\TM1_pad ,
		_w2462_
	);
	LUT2 #(
		.INIT('h4)
	) name954 (
		_w2461_,
		_w2462_,
		_w2463_
	);
	LUT3 #(
		.INIT('hf2)
	) name955 (
		_w1605_,
		_w2460_,
		_w2463_,
		_w2464_
	);
	LUT2 #(
		.INIT('h8)
	) name956 (
		RESET_pad,
		\WX10857_reg/NET0131 ,
		_w2465_
	);
	LUT4 #(
		.INIT('h8cc8)
	) name957 (
		\TM0_pad ,
		_w2313_,
		_w2455_,
		_w2456_,
		_w2466_
	);
	LUT2 #(
		.INIT('h9)
	) name958 (
		\WX8587_reg/NET0131 ,
		\WX8651_reg/NET0131 ,
		_w2467_
	);
	LUT2 #(
		.INIT('h9)
	) name959 (
		\WX8459_reg/NET0131 ,
		\WX8523_reg/NET0131 ,
		_w2468_
	);
	LUT4 #(
		.INIT('h0a02)
	) name960 (
		RESET_pad,
		\TM0_pad ,
		\TM1_pad ,
		\_2240__reg/NET0131 ,
		_w2469_
	);
	LUT4 #(
		.INIT('hbe00)
	) name961 (
		\TM0_pad ,
		_w2467_,
		_w2468_,
		_w2469_,
		_w2470_
	);
	LUT2 #(
		.INIT('he)
	) name962 (
		_w2466_,
		_w2470_,
		_w2471_
	);
	LUT4 #(
		.INIT('ha020)
	) name963 (
		RESET_pad,
		\TM0_pad ,
		\TM1_pad ,
		\WX10891_reg/NET0131 ,
		_w2472_
	);
	LUT2 #(
		.INIT('h9)
	) name964 (
		\WX3421_reg/NET0131 ,
		\WX3485_reg/NET0131 ,
		_w2473_
	);
	LUT2 #(
		.INIT('h9)
	) name965 (
		\WX3293_reg/NET0131 ,
		\WX3357_reg/NET0131 ,
		_w2474_
	);
	LUT4 #(
		.INIT('h8cc8)
	) name966 (
		\TM0_pad ,
		_w2472_,
		_w2473_,
		_w2474_,
		_w2475_
	);
	LUT2 #(
		.INIT('h9)
	) name967 (
		\WX4714_reg/NET0131 ,
		\WX4778_reg/NET0131 ,
		_w2476_
	);
	LUT2 #(
		.INIT('h9)
	) name968 (
		\WX4586_reg/NET0131 ,
		\WX4650_reg/NET0131 ,
		_w2477_
	);
	LUT4 #(
		.INIT('h0a02)
	) name969 (
		RESET_pad,
		\TM0_pad ,
		\TM1_pad ,
		\_2141__reg/NET0131 ,
		_w2478_
	);
	LUT4 #(
		.INIT('hbe00)
	) name970 (
		\TM0_pad ,
		_w2476_,
		_w2477_,
		_w2478_,
		_w2479_
	);
	LUT2 #(
		.INIT('he)
	) name971 (
		_w2475_,
		_w2479_,
		_w2480_
	);
	LUT4 #(
		.INIT('h8cc8)
	) name972 (
		\TM0_pad ,
		_w2258_,
		_w2417_,
		_w2418_,
		_w2481_
	);
	LUT2 #(
		.INIT('h9)
	) name973 (
		\WX9878_reg/NET0131 ,
		\WX9942_reg/NET0131 ,
		_w2482_
	);
	LUT2 #(
		.INIT('h9)
	) name974 (
		\WX9750_reg/NET0131 ,
		\WX9814_reg/NET0131 ,
		_w2483_
	);
	LUT4 #(
		.INIT('h0a02)
	) name975 (
		RESET_pad,
		\TM0_pad ,
		\TM1_pad ,
		\_2273__reg/NET0131 ,
		_w2484_
	);
	LUT4 #(
		.INIT('hbe00)
	) name976 (
		\TM0_pad ,
		_w2482_,
		_w2483_,
		_w2484_,
		_w2485_
	);
	LUT2 #(
		.INIT('he)
	) name977 (
		_w2481_,
		_w2485_,
		_w2486_
	);
	LUT4 #(
		.INIT('h8cc8)
	) name978 (
		\TM0_pad ,
		_w2203_,
		_w2432_,
		_w2433_,
		_w2487_
	);
	LUT2 #(
		.INIT('h9)
	) name979 (
		\WX11169_reg/NET0131 ,
		\WX11233_reg/NET0131 ,
		_w2488_
	);
	LUT2 #(
		.INIT('h9)
	) name980 (
		\WX11041_reg/NET0131 ,
		\WX11105_reg/NET0131 ,
		_w2489_
	);
	LUT4 #(
		.INIT('h0a02)
	) name981 (
		RESET_pad,
		\TM0_pad ,
		\TM1_pad ,
		\_2306__reg/NET0131 ,
		_w2490_
	);
	LUT4 #(
		.INIT('hbe00)
	) name982 (
		\TM0_pad ,
		_w2488_,
		_w2489_,
		_w2490_,
		_w2491_
	);
	LUT2 #(
		.INIT('he)
	) name983 (
		_w2487_,
		_w2491_,
		_w2492_
	);
	LUT4 #(
		.INIT('h8cc8)
	) name984 (
		\TM0_pad ,
		_w2422_,
		_w2426_,
		_w2427_,
		_w2493_
	);
	LUT2 #(
		.INIT('h9)
	) name985 (
		\WX6005_reg/NET0131 ,
		\WX6069_reg/NET0131 ,
		_w2494_
	);
	LUT2 #(
		.INIT('h9)
	) name986 (
		\WX5877_reg/NET0131 ,
		\WX5941_reg/NET0131 ,
		_w2495_
	);
	LUT4 #(
		.INIT('h0a02)
	) name987 (
		RESET_pad,
		\TM0_pad ,
		\TM1_pad ,
		\_2174__reg/NET0131 ,
		_w2496_
	);
	LUT4 #(
		.INIT('hbe00)
	) name988 (
		\TM0_pad ,
		_w2494_,
		_w2495_,
		_w2496_,
		_w2497_
	);
	LUT2 #(
		.INIT('he)
	) name989 (
		_w2493_,
		_w2497_,
		_w2498_
	);
	LUT4 #(
		.INIT('h8cc8)
	) name990 (
		\TM0_pad ,
		_w1606_,
		_w1608_,
		_w1609_,
		_w2499_
	);
	LUT4 #(
		.INIT('h0a02)
	) name991 (
		RESET_pad,
		\TM0_pad ,
		\TM1_pad ,
		\_2124__reg/NET0131 ,
		_w2500_
	);
	LUT4 #(
		.INIT('hbe00)
	) name992 (
		\TM0_pad ,
		_w1646_,
		_w1647_,
		_w2500_,
		_w2501_
	);
	LUT2 #(
		.INIT('he)
	) name993 (
		_w2499_,
		_w2501_,
		_w2502_
	);
	LUT4 #(
		.INIT('h8cc8)
	) name994 (
		\TM0_pad ,
		_w2366_,
		_w2444_,
		_w2445_,
		_w2503_
	);
	LUT2 #(
		.INIT('h9)
	) name995 (
		\WX7296_reg/NET0131 ,
		\WX7360_reg/NET0131 ,
		_w2504_
	);
	LUT2 #(
		.INIT('h9)
	) name996 (
		\WX7168_reg/NET0131 ,
		\WX7232_reg/NET0131 ,
		_w2505_
	);
	LUT4 #(
		.INIT('h0a02)
	) name997 (
		RESET_pad,
		\TM0_pad ,
		\TM1_pad ,
		\_2207__reg/NET0131 ,
		_w2506_
	);
	LUT4 #(
		.INIT('hbe00)
	) name998 (
		\TM0_pad ,
		_w2504_,
		_w2505_,
		_w2506_,
		_w2507_
	);
	LUT2 #(
		.INIT('he)
	) name999 (
		_w2503_,
		_w2507_,
		_w2508_
	);
	LUT3 #(
		.INIT('he0)
	) name1000 (
		\TM0_pad ,
		_w1522_,
		_w1628_,
		_w2509_
	);
	LUT2 #(
		.INIT('h9)
	) name1001 (
		\WX2102_reg/NET0131 ,
		\WX2166_reg/NET0131 ,
		_w2510_
	);
	LUT2 #(
		.INIT('h9)
	) name1002 (
		\WX1974_reg/NET0131 ,
		\WX2038_reg/NET0131 ,
		_w2511_
	);
	LUT4 #(
		.INIT('h0a02)
	) name1003 (
		RESET_pad,
		\TM0_pad ,
		\TM1_pad ,
		\_2090__reg/NET0131 ,
		_w2512_
	);
	LUT4 #(
		.INIT('hbe00)
	) name1004 (
		\TM0_pad ,
		_w2510_,
		_w2511_,
		_w2512_,
		_w2513_
	);
	LUT2 #(
		.INIT('he)
	) name1005 (
		_w2509_,
		_w2513_,
		_w2514_
	);
	LUT2 #(
		.INIT('h8)
	) name1006 (
		RESET_pad,
		\WX10859_reg/NET0131 ,
		_w2515_
	);
	LUT4 #(
		.INIT('h8cc8)
	) name1007 (
		\TM0_pad ,
		_w2366_,
		_w2504_,
		_w2505_,
		_w2516_
	);
	LUT2 #(
		.INIT('h9)
	) name1008 (
		\WX8589_reg/NET0131 ,
		\WX8653_reg/NET0131 ,
		_w2517_
	);
	LUT2 #(
		.INIT('h9)
	) name1009 (
		\WX8461_reg/NET0131 ,
		\WX8525_reg/NET0131 ,
		_w2518_
	);
	LUT4 #(
		.INIT('h0a02)
	) name1010 (
		RESET_pad,
		\TM0_pad ,
		\TM1_pad ,
		\_2239__reg/NET0131 ,
		_w2519_
	);
	LUT4 #(
		.INIT('hbe00)
	) name1011 (
		\TM0_pad ,
		_w2517_,
		_w2518_,
		_w2519_,
		_w2520_
	);
	LUT2 #(
		.INIT('he)
	) name1012 (
		_w2516_,
		_w2520_,
		_w2521_
	);
	LUT4 #(
		.INIT('h8cc8)
	) name1013 (
		\TM0_pad ,
		_w2313_,
		_w2467_,
		_w2468_,
		_w2522_
	);
	LUT2 #(
		.INIT('h9)
	) name1014 (
		\WX9880_reg/NET0131 ,
		\WX9944_reg/NET0131 ,
		_w2523_
	);
	LUT2 #(
		.INIT('h9)
	) name1015 (
		\WX9752_reg/NET0131 ,
		\WX9816_reg/NET0131 ,
		_w2524_
	);
	LUT4 #(
		.INIT('h0a02)
	) name1016 (
		RESET_pad,
		\TM0_pad ,
		\TM1_pad ,
		\_2272__reg/NET0131 ,
		_w2525_
	);
	LUT4 #(
		.INIT('hbe00)
	) name1017 (
		\TM0_pad ,
		_w2523_,
		_w2524_,
		_w2525_,
		_w2526_
	);
	LUT2 #(
		.INIT('he)
	) name1018 (
		_w2522_,
		_w2526_,
		_w2527_
	);
	LUT4 #(
		.INIT('h8cc8)
	) name1019 (
		\TM0_pad ,
		_w2258_,
		_w2482_,
		_w2483_,
		_w2528_
	);
	LUT2 #(
		.INIT('h9)
	) name1020 (
		\WX11171_reg/NET0131 ,
		\WX11235_reg/NET0131 ,
		_w2529_
	);
	LUT2 #(
		.INIT('h9)
	) name1021 (
		\WX11043_reg/NET0131 ,
		\WX11107_reg/NET0131 ,
		_w2530_
	);
	LUT4 #(
		.INIT('h0a02)
	) name1022 (
		RESET_pad,
		\TM0_pad ,
		\TM1_pad ,
		\_2305__reg/NET0131 ,
		_w2531_
	);
	LUT4 #(
		.INIT('hbe00)
	) name1023 (
		\TM0_pad ,
		_w2529_,
		_w2530_,
		_w2531_,
		_w2532_
	);
	LUT2 #(
		.INIT('he)
	) name1024 (
		_w2528_,
		_w2532_,
		_w2533_
	);
	LUT4 #(
		.INIT('h8cc8)
	) name1025 (
		\TM0_pad ,
		_w2472_,
		_w2476_,
		_w2477_,
		_w2534_
	);
	LUT2 #(
		.INIT('h9)
	) name1026 (
		\WX6007_reg/NET0131 ,
		\WX6071_reg/NET0131 ,
		_w2535_
	);
	LUT2 #(
		.INIT('h9)
	) name1027 (
		\WX5879_reg/NET0131 ,
		\WX5943_reg/NET0131 ,
		_w2536_
	);
	LUT4 #(
		.INIT('h0a02)
	) name1028 (
		RESET_pad,
		\TM0_pad ,
		\TM1_pad ,
		\_2173__reg/NET0131 ,
		_w2537_
	);
	LUT4 #(
		.INIT('hbe00)
	) name1029 (
		\TM0_pad ,
		_w2535_,
		_w2536_,
		_w2537_,
		_w2538_
	);
	LUT2 #(
		.INIT('he)
	) name1030 (
		_w2534_,
		_w2538_,
		_w2539_
	);
	LUT2 #(
		.INIT('h9)
	) name1031 (
		\WX2100_reg/NET0131 ,
		\WX2164_reg/NET0131 ,
		_w2540_
	);
	LUT2 #(
		.INIT('h9)
	) name1032 (
		\WX1972_reg/NET0131 ,
		\WX2036_reg/NET0131 ,
		_w2541_
	);
	LUT4 #(
		.INIT('h8cc8)
	) name1033 (
		\TM0_pad ,
		_w1706_,
		_w2540_,
		_w2541_,
		_w2542_
	);
	LUT4 #(
		.INIT('h0a02)
	) name1034 (
		RESET_pad,
		\TM0_pad ,
		\TM1_pad ,
		\_2123__reg/NET0131 ,
		_w2543_
	);
	LUT4 #(
		.INIT('hbe00)
	) name1035 (
		\TM0_pad ,
		_w1707_,
		_w1708_,
		_w2543_,
		_w2544_
	);
	LUT2 #(
		.INIT('he)
	) name1036 (
		_w2542_,
		_w2544_,
		_w2545_
	);
	LUT4 #(
		.INIT('h8cc8)
	) name1037 (
		\TM0_pad ,
		_w2422_,
		_w2494_,
		_w2495_,
		_w2546_
	);
	LUT2 #(
		.INIT('h9)
	) name1038 (
		\WX7298_reg/NET0131 ,
		\WX7362_reg/NET0131 ,
		_w2547_
	);
	LUT2 #(
		.INIT('h9)
	) name1039 (
		\WX7170_reg/NET0131 ,
		\WX7234_reg/NET0131 ,
		_w2548_
	);
	LUT4 #(
		.INIT('h0a02)
	) name1040 (
		RESET_pad,
		\TM0_pad ,
		\TM1_pad ,
		\_2206__reg/NET0131 ,
		_w2549_
	);
	LUT4 #(
		.INIT('hbe00)
	) name1041 (
		\TM0_pad ,
		_w2547_,
		_w2548_,
		_w2549_,
		_w2550_
	);
	LUT2 #(
		.INIT('he)
	) name1042 (
		_w2546_,
		_w2550_,
		_w2551_
	);
	LUT3 #(
		.INIT('h96)
	) name1043 (
		\WX4588_reg/NET0131 ,
		\WX4652_reg/NET0131 ,
		\WX4716_reg/NET0131 ,
		_w2552_
	);
	LUT2 #(
		.INIT('h9)
	) name1044 (
		\TM1_pad ,
		\WX4524_reg/NET0131 ,
		_w2553_
	);
	LUT4 #(
		.INIT('h2772)
	) name1045 (
		\TM0_pad ,
		\_2172__reg/NET0131 ,
		_w2552_,
		_w2553_,
		_w2554_
	);
	LUT3 #(
		.INIT('h96)
	) name1046 (
		\WX3295_reg/NET0131 ,
		\WX3359_reg/NET0131 ,
		\WX3423_reg/NET0131 ,
		_w2555_
	);
	LUT2 #(
		.INIT('h9)
	) name1047 (
		\TM1_pad ,
		\WX3231_reg/NET0131 ,
		_w2556_
	);
	LUT4 #(
		.INIT('h2772)
	) name1048 (
		\TM0_pad ,
		\WX10829_reg/NET0131 ,
		_w2555_,
		_w2556_,
		_w2557_
	);
	LUT4 #(
		.INIT('h028a)
	) name1049 (
		RESET_pad,
		\TM1_pad ,
		_w2554_,
		_w2557_,
		_w2558_
	);
	LUT3 #(
		.INIT('he0)
	) name1050 (
		\TM0_pad ,
		_w1519_,
		_w1810_,
		_w2559_
	);
	LUT2 #(
		.INIT('h9)
	) name1051 (
		\WX2104_reg/NET0131 ,
		\WX2168_reg/NET0131 ,
		_w2560_
	);
	LUT2 #(
		.INIT('h9)
	) name1052 (
		\WX1976_reg/NET0131 ,
		\WX2040_reg/NET0131 ,
		_w2561_
	);
	LUT4 #(
		.INIT('h0a02)
	) name1053 (
		RESET_pad,
		\TM0_pad ,
		\TM1_pad ,
		\_2089__reg/NET0131 ,
		_w2562_
	);
	LUT4 #(
		.INIT('hbe00)
	) name1054 (
		\TM0_pad ,
		_w2560_,
		_w2561_,
		_w2562_,
		_w2563_
	);
	LUT2 #(
		.INIT('he)
	) name1055 (
		_w2559_,
		_w2563_,
		_w2564_
	);
	LUT4 #(
		.INIT('h8cc8)
	) name1056 (
		\TM0_pad ,
		_w1706_,
		_w1994_,
		_w1995_,
		_w2565_
	);
	LUT2 #(
		.INIT('h2)
	) name1057 (
		\TM0_pad ,
		\_2347__reg/NET0131 ,
		_w2566_
	);
	LUT4 #(
		.INIT('h00c8)
	) name1058 (
		\DATA_0_14_pad ,
		RESET_pad,
		\TM0_pad ,
		\TM1_pad ,
		_w2567_
	);
	LUT2 #(
		.INIT('h4)
	) name1059 (
		_w2566_,
		_w2567_,
		_w2568_
	);
	LUT2 #(
		.INIT('he)
	) name1060 (
		_w2565_,
		_w2568_,
		_w2569_
	);
	LUT2 #(
		.INIT('h8)
	) name1061 (
		RESET_pad,
		\WX10861_reg/NET0131 ,
		_w2570_
	);
	LUT4 #(
		.INIT('h8cc8)
	) name1062 (
		\TM0_pad ,
		_w2422_,
		_w2547_,
		_w2548_,
		_w2571_
	);
	LUT2 #(
		.INIT('h9)
	) name1063 (
		\WX8591_reg/NET0131 ,
		\WX8655_reg/NET0131 ,
		_w2572_
	);
	LUT2 #(
		.INIT('h9)
	) name1064 (
		\WX8463_reg/NET0131 ,
		\WX8527_reg/NET0131 ,
		_w2573_
	);
	LUT4 #(
		.INIT('h0a02)
	) name1065 (
		RESET_pad,
		\TM0_pad ,
		\TM1_pad ,
		\_2238__reg/NET0131 ,
		_w2574_
	);
	LUT4 #(
		.INIT('hbe00)
	) name1066 (
		\TM0_pad ,
		_w2572_,
		_w2573_,
		_w2574_,
		_w2575_
	);
	LUT2 #(
		.INIT('he)
	) name1067 (
		_w2571_,
		_w2575_,
		_w2576_
	);
	LUT4 #(
		.INIT('h8cc8)
	) name1068 (
		\TM0_pad ,
		_w2366_,
		_w2517_,
		_w2518_,
		_w2577_
	);
	LUT2 #(
		.INIT('h9)
	) name1069 (
		\WX9882_reg/NET0131 ,
		\WX9946_reg/NET0131 ,
		_w2578_
	);
	LUT2 #(
		.INIT('h9)
	) name1070 (
		\WX9754_reg/NET0131 ,
		\WX9818_reg/NET0131 ,
		_w2579_
	);
	LUT4 #(
		.INIT('h0a02)
	) name1071 (
		RESET_pad,
		\TM0_pad ,
		\TM1_pad ,
		\_2271__reg/NET0131 ,
		_w2580_
	);
	LUT4 #(
		.INIT('hbe00)
	) name1072 (
		\TM0_pad ,
		_w2578_,
		_w2579_,
		_w2580_,
		_w2581_
	);
	LUT2 #(
		.INIT('he)
	) name1073 (
		_w2577_,
		_w2581_,
		_w2582_
	);
	LUT3 #(
		.INIT('h96)
	) name1074 (
		\WX5881_reg/NET0131 ,
		\WX5945_reg/NET0131 ,
		\WX6009_reg/NET0131 ,
		_w2583_
	);
	LUT2 #(
		.INIT('h9)
	) name1075 (
		\TM1_pad ,
		\WX5817_reg/NET0131 ,
		_w2584_
	);
	LUT4 #(
		.INIT('h2772)
	) name1076 (
		\TM0_pad ,
		\_2204__reg/NET0131 ,
		_w2583_,
		_w2584_,
		_w2585_
	);
	LUT4 #(
		.INIT('h2772)
	) name1077 (
		\TM0_pad ,
		\WX10829_reg/NET0131 ,
		_w2552_,
		_w2553_,
		_w2586_
	);
	LUT4 #(
		.INIT('h028a)
	) name1078 (
		RESET_pad,
		\TM1_pad ,
		_w2585_,
		_w2586_,
		_w2587_
	);
	LUT4 #(
		.INIT('h8cc8)
	) name1079 (
		\TM0_pad ,
		_w2313_,
		_w2523_,
		_w2524_,
		_w2588_
	);
	LUT2 #(
		.INIT('h9)
	) name1080 (
		\WX11173_reg/NET0131 ,
		\WX11237_reg/NET0131 ,
		_w2589_
	);
	LUT2 #(
		.INIT('h9)
	) name1081 (
		\WX11045_reg/NET0131 ,
		\WX11109_reg/NET0131 ,
		_w2590_
	);
	LUT4 #(
		.INIT('h0a02)
	) name1082 (
		RESET_pad,
		\TM0_pad ,
		\TM1_pad ,
		\_2304__reg/NET0131 ,
		_w2591_
	);
	LUT4 #(
		.INIT('hbe00)
	) name1083 (
		\TM0_pad ,
		_w2589_,
		_w2590_,
		_w2591_,
		_w2592_
	);
	LUT2 #(
		.INIT('he)
	) name1084 (
		_w2588_,
		_w2592_,
		_w2593_
	);
	LUT4 #(
		.INIT('h8cc8)
	) name1085 (
		\TM0_pad ,
		_w1628_,
		_w2510_,
		_w2511_,
		_w2594_
	);
	LUT4 #(
		.INIT('h0a02)
	) name1086 (
		RESET_pad,
		\TM0_pad ,
		\TM1_pad ,
		\_2122__reg/NET0131 ,
		_w2595_
	);
	LUT4 #(
		.INIT('hbe00)
	) name1087 (
		\TM0_pad ,
		_w1759_,
		_w1760_,
		_w2595_,
		_w2596_
	);
	LUT2 #(
		.INIT('he)
	) name1088 (
		_w2594_,
		_w2596_,
		_w2597_
	);
	LUT4 #(
		.INIT('h8cc8)
	) name1089 (
		\TM0_pad ,
		_w2472_,
		_w2535_,
		_w2536_,
		_w2598_
	);
	LUT2 #(
		.INIT('h9)
	) name1090 (
		\WX7300_reg/NET0131 ,
		\WX7364_reg/NET0131 ,
		_w2599_
	);
	LUT2 #(
		.INIT('h9)
	) name1091 (
		\WX7172_reg/NET0131 ,
		\WX7236_reg/NET0131 ,
		_w2600_
	);
	LUT4 #(
		.INIT('h0a02)
	) name1092 (
		RESET_pad,
		\TM0_pad ,
		\TM1_pad ,
		\_2205__reg/NET0131 ,
		_w2601_
	);
	LUT4 #(
		.INIT('hbe00)
	) name1093 (
		\TM0_pad ,
		_w2599_,
		_w2600_,
		_w2601_,
		_w2602_
	);
	LUT2 #(
		.INIT('he)
	) name1094 (
		_w2598_,
		_w2602_,
		_w2603_
	);
	LUT3 #(
		.INIT('h96)
	) name1095 (
		\WX4590_reg/NET0131 ,
		\WX4654_reg/NET0131 ,
		\WX4718_reg/NET0131 ,
		_w2604_
	);
	LUT2 #(
		.INIT('h9)
	) name1096 (
		\TM1_pad ,
		\WX4526_reg/NET0131 ,
		_w2605_
	);
	LUT4 #(
		.INIT('h2772)
	) name1097 (
		\TM0_pad ,
		\_2171__reg/NET0131 ,
		_w2604_,
		_w2605_,
		_w2606_
	);
	LUT4 #(
		.INIT('h2772)
	) name1098 (
		\TM0_pad ,
		\WX10831_reg/NET0131 ,
		_w1654_,
		_w1655_,
		_w2607_
	);
	LUT4 #(
		.INIT('h028a)
	) name1099 (
		RESET_pad,
		\TM1_pad ,
		_w2606_,
		_w2607_,
		_w2608_
	);
	LUT2 #(
		.INIT('h8)
	) name1100 (
		RESET_pad,
		\WX10863_reg/NET0131 ,
		_w2609_
	);
	LUT4 #(
		.INIT('h8cc8)
	) name1101 (
		\TM0_pad ,
		_w2472_,
		_w2599_,
		_w2600_,
		_w2610_
	);
	LUT2 #(
		.INIT('h9)
	) name1102 (
		\WX8593_reg/NET0131 ,
		\WX8657_reg/NET0131 ,
		_w2611_
	);
	LUT2 #(
		.INIT('h9)
	) name1103 (
		\WX8465_reg/NET0131 ,
		\WX8529_reg/NET0131 ,
		_w2612_
	);
	LUT4 #(
		.INIT('h0a02)
	) name1104 (
		RESET_pad,
		\TM0_pad ,
		\TM1_pad ,
		\_2237__reg/NET0131 ,
		_w2613_
	);
	LUT4 #(
		.INIT('hbe00)
	) name1105 (
		\TM0_pad ,
		_w2611_,
		_w2612_,
		_w2613_,
		_w2614_
	);
	LUT2 #(
		.INIT('he)
	) name1106 (
		_w2610_,
		_w2614_,
		_w2615_
	);
	LUT4 #(
		.INIT('h8cc8)
	) name1107 (
		\TM0_pad ,
		_w2422_,
		_w2572_,
		_w2573_,
		_w2616_
	);
	LUT2 #(
		.INIT('h9)
	) name1108 (
		\WX9884_reg/NET0131 ,
		\WX9948_reg/NET0131 ,
		_w2617_
	);
	LUT2 #(
		.INIT('h9)
	) name1109 (
		\WX9756_reg/NET0131 ,
		\WX9820_reg/NET0131 ,
		_w2618_
	);
	LUT4 #(
		.INIT('h0a02)
	) name1110 (
		RESET_pad,
		\TM0_pad ,
		\TM1_pad ,
		\_2270__reg/NET0131 ,
		_w2619_
	);
	LUT4 #(
		.INIT('hbe00)
	) name1111 (
		\TM0_pad ,
		_w2617_,
		_w2618_,
		_w2619_,
		_w2620_
	);
	LUT2 #(
		.INIT('he)
	) name1112 (
		_w2616_,
		_w2620_,
		_w2621_
	);
	LUT3 #(
		.INIT('h96)
	) name1113 (
		\WX5883_reg/NET0131 ,
		\WX5947_reg/NET0131 ,
		\WX6011_reg/NET0131 ,
		_w2622_
	);
	LUT2 #(
		.INIT('h9)
	) name1114 (
		\TM1_pad ,
		\WX5819_reg/NET0131 ,
		_w2623_
	);
	LUT4 #(
		.INIT('h2772)
	) name1115 (
		\TM0_pad ,
		\_2203__reg/NET0131 ,
		_w2622_,
		_w2623_,
		_w2624_
	);
	LUT4 #(
		.INIT('h2772)
	) name1116 (
		\TM0_pad ,
		\WX10831_reg/NET0131 ,
		_w2604_,
		_w2605_,
		_w2625_
	);
	LUT4 #(
		.INIT('h028a)
	) name1117 (
		RESET_pad,
		\TM1_pad ,
		_w2624_,
		_w2625_,
		_w2626_
	);
	LUT4 #(
		.INIT('h8cc8)
	) name1118 (
		\TM0_pad ,
		_w2366_,
		_w2578_,
		_w2579_,
		_w2627_
	);
	LUT2 #(
		.INIT('h9)
	) name1119 (
		\WX11175_reg/NET0131 ,
		\WX11239_reg/NET0131 ,
		_w2628_
	);
	LUT2 #(
		.INIT('h9)
	) name1120 (
		\WX11047_reg/NET0131 ,
		\WX11111_reg/NET0131 ,
		_w2629_
	);
	LUT4 #(
		.INIT('h0a02)
	) name1121 (
		RESET_pad,
		\TM0_pad ,
		\TM1_pad ,
		\_2303__reg/NET0131 ,
		_w2630_
	);
	LUT4 #(
		.INIT('hbe00)
	) name1122 (
		\TM0_pad ,
		_w2628_,
		_w2629_,
		_w2630_,
		_w2631_
	);
	LUT2 #(
		.INIT('he)
	) name1123 (
		_w2627_,
		_w2631_,
		_w2632_
	);
	LUT3 #(
		.INIT('h96)
	) name1124 (
		\WX7174_reg/NET0131 ,
		\WX7238_reg/NET0131 ,
		\WX7302_reg/NET0131 ,
		_w2633_
	);
	LUT2 #(
		.INIT('h9)
	) name1125 (
		\TM1_pad ,
		\WX7110_reg/NET0131 ,
		_w2634_
	);
	LUT4 #(
		.INIT('h2772)
	) name1126 (
		\TM0_pad ,
		\_2236__reg/NET0131 ,
		_w2633_,
		_w2634_,
		_w2635_
	);
	LUT4 #(
		.INIT('h2772)
	) name1127 (
		\TM0_pad ,
		\WX10829_reg/NET0131 ,
		_w2583_,
		_w2584_,
		_w2636_
	);
	LUT4 #(
		.INIT('h028a)
	) name1128 (
		RESET_pad,
		\TM1_pad ,
		_w2635_,
		_w2636_,
		_w2637_
	);
	LUT4 #(
		.INIT('h8cc8)
	) name1129 (
		\TM0_pad ,
		_w1810_,
		_w2560_,
		_w2561_,
		_w2638_
	);
	LUT4 #(
		.INIT('h0a02)
	) name1130 (
		RESET_pad,
		\TM0_pad ,
		\TM1_pad ,
		\_2121__reg/NET0131 ,
		_w2639_
	);
	LUT4 #(
		.INIT('hbe00)
	) name1131 (
		\TM0_pad ,
		_w1811_,
		_w1812_,
		_w2639_,
		_w2640_
	);
	LUT2 #(
		.INIT('he)
	) name1132 (
		_w2638_,
		_w2640_,
		_w2641_
	);
	LUT3 #(
		.INIT('h96)
	) name1133 (
		\WX4592_reg/NET0131 ,
		\WX4656_reg/NET0131 ,
		\WX4720_reg/NET0131 ,
		_w2642_
	);
	LUT2 #(
		.INIT('h9)
	) name1134 (
		\TM1_pad ,
		\WX4528_reg/NET0131 ,
		_w2643_
	);
	LUT4 #(
		.INIT('h2772)
	) name1135 (
		\TM0_pad ,
		\_2170__reg/NET0131 ,
		_w2642_,
		_w2643_,
		_w2644_
	);
	LUT4 #(
		.INIT('h2772)
	) name1136 (
		\TM0_pad ,
		\WX10833_reg/NET0131 ,
		_w1720_,
		_w1721_,
		_w2645_
	);
	LUT4 #(
		.INIT('h028a)
	) name1137 (
		RESET_pad,
		\TM1_pad ,
		_w2644_,
		_w2645_,
		_w2646_
	);
	LUT3 #(
		.INIT('he0)
	) name1138 (
		\TM0_pad ,
		_w1513_,
		_w1921_,
		_w2647_
	);
	LUT2 #(
		.INIT('h9)
	) name1139 (
		\WX2108_reg/NET0131 ,
		\WX2172_reg/NET0131 ,
		_w2648_
	);
	LUT2 #(
		.INIT('h9)
	) name1140 (
		\WX1980_reg/NET0131 ,
		\WX2044_reg/NET0131 ,
		_w2649_
	);
	LUT4 #(
		.INIT('h0a02)
	) name1141 (
		RESET_pad,
		\TM0_pad ,
		\TM1_pad ,
		\_2087__reg/NET0131 ,
		_w2650_
	);
	LUT4 #(
		.INIT('hbe00)
	) name1142 (
		\TM0_pad ,
		_w2648_,
		_w2649_,
		_w2650_,
		_w2651_
	);
	LUT2 #(
		.INIT('he)
	) name1143 (
		_w2647_,
		_w2651_,
		_w2652_
	);
	LUT4 #(
		.INIT('h8cc8)
	) name1144 (
		\TM0_pad ,
		_w1810_,
		_w2105_,
		_w2106_,
		_w2653_
	);
	LUT2 #(
		.INIT('h2)
	) name1145 (
		\TM0_pad ,
		\_2345__reg/NET0131 ,
		_w2654_
	);
	LUT4 #(
		.INIT('h00c8)
	) name1146 (
		\DATA_0_12_pad ,
		RESET_pad,
		\TM0_pad ,
		\TM1_pad ,
		_w2655_
	);
	LUT2 #(
		.INIT('h4)
	) name1147 (
		_w2654_,
		_w2655_,
		_w2656_
	);
	LUT2 #(
		.INIT('he)
	) name1148 (
		_w2653_,
		_w2656_,
		_w2657_
	);
	LUT2 #(
		.INIT('h8)
	) name1149 (
		RESET_pad,
		\WX10865_reg/NET0131 ,
		_w2658_
	);
	LUT4 #(
		.INIT('h8cc8)
	) name1150 (
		\TM0_pad ,
		_w2472_,
		_w2611_,
		_w2612_,
		_w2659_
	);
	LUT2 #(
		.INIT('h9)
	) name1151 (
		\WX9886_reg/NET0131 ,
		\WX9950_reg/NET0131 ,
		_w2660_
	);
	LUT2 #(
		.INIT('h9)
	) name1152 (
		\WX9758_reg/NET0131 ,
		\WX9822_reg/NET0131 ,
		_w2661_
	);
	LUT4 #(
		.INIT('h0a02)
	) name1153 (
		RESET_pad,
		\TM0_pad ,
		\TM1_pad ,
		\_2269__reg/NET0131 ,
		_w2662_
	);
	LUT4 #(
		.INIT('hbe00)
	) name1154 (
		\TM0_pad ,
		_w2660_,
		_w2661_,
		_w2662_,
		_w2663_
	);
	LUT2 #(
		.INIT('he)
	) name1155 (
		_w2659_,
		_w2663_,
		_w2664_
	);
	LUT3 #(
		.INIT('h96)
	) name1156 (
		\WX5885_reg/NET0131 ,
		\WX5949_reg/NET0131 ,
		\WX6013_reg/NET0131 ,
		_w2665_
	);
	LUT2 #(
		.INIT('h9)
	) name1157 (
		\TM1_pad ,
		\WX5821_reg/NET0131 ,
		_w2666_
	);
	LUT4 #(
		.INIT('h2772)
	) name1158 (
		\TM0_pad ,
		\_2202__reg/NET0131 ,
		_w2665_,
		_w2666_,
		_w2667_
	);
	LUT4 #(
		.INIT('h2772)
	) name1159 (
		\TM0_pad ,
		\WX10833_reg/NET0131 ,
		_w2642_,
		_w2643_,
		_w2668_
	);
	LUT4 #(
		.INIT('h028a)
	) name1160 (
		RESET_pad,
		\TM1_pad ,
		_w2667_,
		_w2668_,
		_w2669_
	);
	LUT4 #(
		.INIT('h8cc8)
	) name1161 (
		\TM0_pad ,
		_w2422_,
		_w2617_,
		_w2618_,
		_w2670_
	);
	LUT2 #(
		.INIT('h9)
	) name1162 (
		\WX11177_reg/NET0131 ,
		\WX11241_reg/NET0131 ,
		_w2671_
	);
	LUT2 #(
		.INIT('h9)
	) name1163 (
		\WX11049_reg/NET0131 ,
		\WX11113_reg/NET0131 ,
		_w2672_
	);
	LUT4 #(
		.INIT('h0a02)
	) name1164 (
		RESET_pad,
		\TM0_pad ,
		\TM1_pad ,
		\_2302__reg/NET0131 ,
		_w2673_
	);
	LUT4 #(
		.INIT('hbe00)
	) name1165 (
		\TM0_pad ,
		_w2671_,
		_w2672_,
		_w2673_,
		_w2674_
	);
	LUT2 #(
		.INIT('he)
	) name1166 (
		_w2670_,
		_w2674_,
		_w2675_
	);
	LUT3 #(
		.INIT('h69)
	) name1167 (
		\TM1_pad ,
		\WX7112_reg/NET0131 ,
		\WX7176_reg/NET0131 ,
		_w2676_
	);
	LUT2 #(
		.INIT('h9)
	) name1168 (
		\WX7240_reg/NET0131 ,
		\WX7304_reg/NET0131 ,
		_w2677_
	);
	LUT4 #(
		.INIT('h7227)
	) name1169 (
		\TM0_pad ,
		\_2235__reg/NET0131 ,
		_w2676_,
		_w2677_,
		_w2678_
	);
	LUT4 #(
		.INIT('h2772)
	) name1170 (
		\TM0_pad ,
		\WX10831_reg/NET0131 ,
		_w2622_,
		_w2623_,
		_w2679_
	);
	LUT4 #(
		.INIT('h028a)
	) name1171 (
		RESET_pad,
		\TM1_pad ,
		_w2678_,
		_w2679_,
		_w2680_
	);
	LUT2 #(
		.INIT('h9)
	) name1172 (
		\WX2106_reg/NET0131 ,
		\WX2170_reg/NET0131 ,
		_w2681_
	);
	LUT2 #(
		.INIT('h9)
	) name1173 (
		\WX1978_reg/NET0131 ,
		\WX2042_reg/NET0131 ,
		_w2682_
	);
	LUT4 #(
		.INIT('h8cc8)
	) name1174 (
		\TM0_pad ,
		_w1865_,
		_w2681_,
		_w2682_,
		_w2683_
	);
	LUT4 #(
		.INIT('h0a02)
	) name1175 (
		RESET_pad,
		\TM0_pad ,
		\TM1_pad ,
		\_2120__reg/NET0131 ,
		_w2684_
	);
	LUT4 #(
		.INIT('hbe00)
	) name1176 (
		\TM0_pad ,
		_w1866_,
		_w1867_,
		_w2684_,
		_w2685_
	);
	LUT2 #(
		.INIT('he)
	) name1177 (
		_w2683_,
		_w2685_,
		_w2686_
	);
	LUT3 #(
		.INIT('h96)
	) name1178 (
		\WX8467_reg/NET0131 ,
		\WX8531_reg/NET0131 ,
		\WX8595_reg/NET0131 ,
		_w2687_
	);
	LUT2 #(
		.INIT('h9)
	) name1179 (
		\TM1_pad ,
		\WX8403_reg/NET0131 ,
		_w2688_
	);
	LUT4 #(
		.INIT('h2772)
	) name1180 (
		\TM0_pad ,
		\_2268__reg/NET0131 ,
		_w2687_,
		_w2688_,
		_w2689_
	);
	LUT4 #(
		.INIT('h2772)
	) name1181 (
		\TM0_pad ,
		\WX10829_reg/NET0131 ,
		_w2633_,
		_w2634_,
		_w2690_
	);
	LUT4 #(
		.INIT('h028a)
	) name1182 (
		RESET_pad,
		\TM1_pad ,
		_w2689_,
		_w2690_,
		_w2691_
	);
	LUT3 #(
		.INIT('h96)
	) name1183 (
		\WX4594_reg/NET0131 ,
		\WX4658_reg/NET0131 ,
		\WX4722_reg/NET0131 ,
		_w2692_
	);
	LUT2 #(
		.INIT('h9)
	) name1184 (
		\TM1_pad ,
		\WX4530_reg/NET0131 ,
		_w2693_
	);
	LUT4 #(
		.INIT('h2772)
	) name1185 (
		\TM0_pad ,
		\_2169__reg/NET0131 ,
		_w2692_,
		_w2693_,
		_w2694_
	);
	LUT4 #(
		.INIT('h2772)
	) name1186 (
		\TM0_pad ,
		\WX10835_reg/NET0131 ,
		_w1772_,
		_w1773_,
		_w2695_
	);
	LUT4 #(
		.INIT('h028a)
	) name1187 (
		RESET_pad,
		\TM1_pad ,
		_w2694_,
		_w2695_,
		_w2696_
	);
	LUT4 #(
		.INIT('h8cc8)
	) name1188 (
		\TM0_pad ,
		_w1865_,
		_w2162_,
		_w2163_,
		_w2697_
	);
	LUT2 #(
		.INIT('h2)
	) name1189 (
		\TM0_pad ,
		\_2344__reg/NET0131 ,
		_w2698_
	);
	LUT4 #(
		.INIT('h00c8)
	) name1190 (
		\DATA_0_11_pad ,
		RESET_pad,
		\TM0_pad ,
		\TM1_pad ,
		_w2699_
	);
	LUT2 #(
		.INIT('h4)
	) name1191 (
		_w2698_,
		_w2699_,
		_w2700_
	);
	LUT2 #(
		.INIT('he)
	) name1192 (
		_w2697_,
		_w2700_,
		_w2701_
	);
	LUT2 #(
		.INIT('h8)
	) name1193 (
		RESET_pad,
		\WX10867_reg/NET0131 ,
		_w2702_
	);
	LUT3 #(
		.INIT('h96)
	) name1194 (
		\WX9760_reg/NET0131 ,
		\WX9824_reg/NET0131 ,
		\WX9888_reg/NET0131 ,
		_w2703_
	);
	LUT2 #(
		.INIT('h9)
	) name1195 (
		\TM1_pad ,
		\WX9696_reg/NET0131 ,
		_w2704_
	);
	LUT4 #(
		.INIT('h2772)
	) name1196 (
		\TM0_pad ,
		\_2300__reg/NET0131 ,
		_w2703_,
		_w2704_,
		_w2705_
	);
	LUT4 #(
		.INIT('h2772)
	) name1197 (
		\TM0_pad ,
		\WX10829_reg/NET0131 ,
		_w2687_,
		_w2688_,
		_w2706_
	);
	LUT4 #(
		.INIT('h028a)
	) name1198 (
		RESET_pad,
		\TM1_pad ,
		_w2705_,
		_w2706_,
		_w2707_
	);
	LUT3 #(
		.INIT('h96)
	) name1199 (
		\WX5887_reg/NET0131 ,
		\WX5951_reg/NET0131 ,
		\WX6015_reg/NET0131 ,
		_w2708_
	);
	LUT2 #(
		.INIT('h9)
	) name1200 (
		\TM1_pad ,
		\WX5823_reg/NET0131 ,
		_w2709_
	);
	LUT4 #(
		.INIT('h2772)
	) name1201 (
		\TM0_pad ,
		\_2201__reg/NET0131 ,
		_w2708_,
		_w2709_,
		_w2710_
	);
	LUT4 #(
		.INIT('h2772)
	) name1202 (
		\TM0_pad ,
		\WX10835_reg/NET0131 ,
		_w2692_,
		_w2693_,
		_w2711_
	);
	LUT4 #(
		.INIT('h028a)
	) name1203 (
		RESET_pad,
		\TM1_pad ,
		_w2710_,
		_w2711_,
		_w2712_
	);
	LUT4 #(
		.INIT('h8cc8)
	) name1204 (
		\TM0_pad ,
		_w2472_,
		_w2660_,
		_w2661_,
		_w2713_
	);
	LUT2 #(
		.INIT('h9)
	) name1205 (
		\WX11179_reg/NET0131 ,
		\WX11243_reg/NET0131 ,
		_w2714_
	);
	LUT2 #(
		.INIT('h9)
	) name1206 (
		\WX11051_reg/NET0131 ,
		\WX11115_reg/NET0131 ,
		_w2715_
	);
	LUT4 #(
		.INIT('h0a02)
	) name1207 (
		RESET_pad,
		\TM0_pad ,
		\TM1_pad ,
		\_2301__reg/NET0131 ,
		_w2716_
	);
	LUT4 #(
		.INIT('hbe00)
	) name1208 (
		\TM0_pad ,
		_w2714_,
		_w2715_,
		_w2716_,
		_w2717_
	);
	LUT2 #(
		.INIT('he)
	) name1209 (
		_w2713_,
		_w2717_,
		_w2718_
	);
	LUT3 #(
		.INIT('h96)
	) name1210 (
		\WX7178_reg/NET0131 ,
		\WX7242_reg/NET0131 ,
		\WX7306_reg/NET0131 ,
		_w2719_
	);
	LUT2 #(
		.INIT('h9)
	) name1211 (
		\TM1_pad ,
		\WX7114_reg/NET0131 ,
		_w2720_
	);
	LUT4 #(
		.INIT('h2772)
	) name1212 (
		\TM0_pad ,
		\_2234__reg/NET0131 ,
		_w2719_,
		_w2720_,
		_w2721_
	);
	LUT4 #(
		.INIT('h2772)
	) name1213 (
		\TM0_pad ,
		\WX10833_reg/NET0131 ,
		_w2665_,
		_w2666_,
		_w2722_
	);
	LUT4 #(
		.INIT('h028a)
	) name1214 (
		RESET_pad,
		\TM1_pad ,
		_w2721_,
		_w2722_,
		_w2723_
	);
	LUT4 #(
		.INIT('h8cc8)
	) name1215 (
		\TM0_pad ,
		_w1921_,
		_w2648_,
		_w2649_,
		_w2724_
	);
	LUT4 #(
		.INIT('h0a02)
	) name1216 (
		RESET_pad,
		\TM0_pad ,
		\TM1_pad ,
		\_2119__reg/NET0131 ,
		_w2725_
	);
	LUT4 #(
		.INIT('hbe00)
	) name1217 (
		\TM0_pad ,
		_w1922_,
		_w1923_,
		_w2725_,
		_w2726_
	);
	LUT2 #(
		.INIT('he)
	) name1218 (
		_w2724_,
		_w2726_,
		_w2727_
	);
	LUT3 #(
		.INIT('h96)
	) name1219 (
		\WX8469_reg/NET0131 ,
		\WX8533_reg/NET0131 ,
		\WX8597_reg/NET0131 ,
		_w2728_
	);
	LUT2 #(
		.INIT('h9)
	) name1220 (
		\TM1_pad ,
		\WX8405_reg/NET0131 ,
		_w2729_
	);
	LUT4 #(
		.INIT('h2772)
	) name1221 (
		\TM0_pad ,
		\_2267__reg/NET0131 ,
		_w2728_,
		_w2729_,
		_w2730_
	);
	LUT4 #(
		.INIT('h7227)
	) name1222 (
		\TM0_pad ,
		\WX10831_reg/NET0131 ,
		_w2676_,
		_w2677_,
		_w2731_
	);
	LUT4 #(
		.INIT('h028a)
	) name1223 (
		RESET_pad,
		\TM1_pad ,
		_w2730_,
		_w2731_,
		_w2732_
	);
	LUT3 #(
		.INIT('h96)
	) name1224 (
		\WX4596_reg/NET0131 ,
		\WX4660_reg/NET0131 ,
		\WX4724_reg/NET0131 ,
		_w2733_
	);
	LUT2 #(
		.INIT('h9)
	) name1225 (
		\TM1_pad ,
		\WX4532_reg/NET0131 ,
		_w2734_
	);
	LUT4 #(
		.INIT('h2772)
	) name1226 (
		\TM0_pad ,
		\_2168__reg/NET0131 ,
		_w2733_,
		_w2734_,
		_w2735_
	);
	LUT4 #(
		.INIT('h2772)
	) name1227 (
		\TM0_pad ,
		\WX10837_reg/NET0131 ,
		_w1824_,
		_w1825_,
		_w2736_
	);
	LUT4 #(
		.INIT('h028a)
	) name1228 (
		RESET_pad,
		\TM1_pad ,
		_w2735_,
		_w2736_,
		_w2737_
	);
	LUT4 #(
		.INIT('h8cc8)
	) name1229 (
		\TM0_pad ,
		_w1921_,
		_w2219_,
		_w2220_,
		_w2738_
	);
	LUT2 #(
		.INIT('h2)
	) name1230 (
		\TM0_pad ,
		\_2343__reg/NET0131 ,
		_w2739_
	);
	LUT4 #(
		.INIT('h00c8)
	) name1231 (
		\DATA_0_10_pad ,
		RESET_pad,
		\TM0_pad ,
		\TM1_pad ,
		_w2740_
	);
	LUT2 #(
		.INIT('h4)
	) name1232 (
		_w2739_,
		_w2740_,
		_w2741_
	);
	LUT2 #(
		.INIT('he)
	) name1233 (
		_w2738_,
		_w2741_,
		_w2742_
	);
	LUT2 #(
		.INIT('h8)
	) name1234 (
		RESET_pad,
		\WX10869_reg/NET0131 ,
		_w2743_
	);
	LUT3 #(
		.INIT('h96)
	) name1235 (
		\WX9762_reg/NET0131 ,
		\WX9826_reg/NET0131 ,
		\WX9890_reg/NET0131 ,
		_w2744_
	);
	LUT2 #(
		.INIT('h9)
	) name1236 (
		\TM1_pad ,
		\WX9698_reg/NET0131 ,
		_w2745_
	);
	LUT4 #(
		.INIT('h2772)
	) name1237 (
		\TM0_pad ,
		\_2299__reg/NET0131 ,
		_w2744_,
		_w2745_,
		_w2746_
	);
	LUT4 #(
		.INIT('h2772)
	) name1238 (
		\TM0_pad ,
		\WX10831_reg/NET0131 ,
		_w2728_,
		_w2729_,
		_w2747_
	);
	LUT4 #(
		.INIT('h028a)
	) name1239 (
		RESET_pad,
		\TM1_pad ,
		_w2746_,
		_w2747_,
		_w2748_
	);
	LUT3 #(
		.INIT('h69)
	) name1240 (
		\TM1_pad ,
		\WX10989_reg/NET0131 ,
		\WX11053_reg/NET0131 ,
		_w2749_
	);
	LUT2 #(
		.INIT('h9)
	) name1241 (
		\WX11117_reg/NET0131 ,
		\WX11181_reg/NET0131 ,
		_w2750_
	);
	LUT4 #(
		.INIT('h7227)
	) name1242 (
		\TM0_pad ,
		\_2332__reg/NET0131 ,
		_w2749_,
		_w2750_,
		_w2751_
	);
	LUT4 #(
		.INIT('h2772)
	) name1243 (
		\TM0_pad ,
		\WX10829_reg/NET0131 ,
		_w2703_,
		_w2704_,
		_w2752_
	);
	LUT4 #(
		.INIT('h028a)
	) name1244 (
		RESET_pad,
		\TM1_pad ,
		_w2751_,
		_w2752_,
		_w2753_
	);
	LUT3 #(
		.INIT('h96)
	) name1245 (
		\WX5889_reg/NET0131 ,
		\WX5953_reg/NET0131 ,
		\WX6017_reg/NET0131 ,
		_w2754_
	);
	LUT2 #(
		.INIT('h9)
	) name1246 (
		\TM1_pad ,
		\WX5825_reg/NET0131 ,
		_w2755_
	);
	LUT4 #(
		.INIT('h2772)
	) name1247 (
		\TM0_pad ,
		\_2200__reg/NET0131 ,
		_w2754_,
		_w2755_,
		_w2756_
	);
	LUT4 #(
		.INIT('h2772)
	) name1248 (
		\TM0_pad ,
		\WX10837_reg/NET0131 ,
		_w2733_,
		_w2734_,
		_w2757_
	);
	LUT4 #(
		.INIT('h028a)
	) name1249 (
		RESET_pad,
		\TM1_pad ,
		_w2756_,
		_w2757_,
		_w2758_
	);
	LUT3 #(
		.INIT('h96)
	) name1250 (
		\WX7180_reg/NET0131 ,
		\WX7244_reg/NET0131 ,
		\WX7308_reg/NET0131 ,
		_w2759_
	);
	LUT2 #(
		.INIT('h9)
	) name1251 (
		\TM1_pad ,
		\WX7116_reg/NET0131 ,
		_w2760_
	);
	LUT4 #(
		.INIT('h2772)
	) name1252 (
		\TM0_pad ,
		\_2233__reg/NET0131 ,
		_w2759_,
		_w2760_,
		_w2761_
	);
	LUT4 #(
		.INIT('h2772)
	) name1253 (
		\TM0_pad ,
		\WX10835_reg/NET0131 ,
		_w2708_,
		_w2709_,
		_w2762_
	);
	LUT4 #(
		.INIT('h028a)
	) name1254 (
		RESET_pad,
		\TM1_pad ,
		_w2761_,
		_w2762_,
		_w2763_
	);
	LUT2 #(
		.INIT('h9)
	) name1255 (
		\WX2110_reg/NET0131 ,
		\WX2174_reg/NET0131 ,
		_w2764_
	);
	LUT2 #(
		.INIT('h9)
	) name1256 (
		\WX1982_reg/NET0131 ,
		\WX2046_reg/NET0131 ,
		_w2765_
	);
	LUT4 #(
		.INIT('h8cc8)
	) name1257 (
		\TM0_pad ,
		_w1978_,
		_w2764_,
		_w2765_,
		_w2766_
	);
	LUT4 #(
		.INIT('h0a02)
	) name1258 (
		RESET_pad,
		\TM0_pad ,
		\TM1_pad ,
		\_2118__reg/NET0131 ,
		_w2767_
	);
	LUT4 #(
		.INIT('hbe00)
	) name1259 (
		\TM0_pad ,
		_w1979_,
		_w1980_,
		_w2767_,
		_w2768_
	);
	LUT2 #(
		.INIT('he)
	) name1260 (
		_w2766_,
		_w2768_,
		_w2769_
	);
	LUT3 #(
		.INIT('h96)
	) name1261 (
		\WX8471_reg/NET0131 ,
		\WX8535_reg/NET0131 ,
		\WX8599_reg/NET0131 ,
		_w2770_
	);
	LUT2 #(
		.INIT('h9)
	) name1262 (
		\TM1_pad ,
		\WX8407_reg/NET0131 ,
		_w2771_
	);
	LUT4 #(
		.INIT('h2772)
	) name1263 (
		\TM0_pad ,
		\_2266__reg/NET0131 ,
		_w2770_,
		_w2771_,
		_w2772_
	);
	LUT4 #(
		.INIT('h2772)
	) name1264 (
		\TM0_pad ,
		\WX10833_reg/NET0131 ,
		_w2719_,
		_w2720_,
		_w2773_
	);
	LUT4 #(
		.INIT('h028a)
	) name1265 (
		RESET_pad,
		\TM1_pad ,
		_w2772_,
		_w2773_,
		_w2774_
	);
	LUT3 #(
		.INIT('h96)
	) name1266 (
		\WX4598_reg/NET0131 ,
		\WX4662_reg/NET0131 ,
		\WX4726_reg/NET0131 ,
		_w2775_
	);
	LUT2 #(
		.INIT('h9)
	) name1267 (
		\TM1_pad ,
		\WX4534_reg/NET0131 ,
		_w2776_
	);
	LUT4 #(
		.INIT('h2772)
	) name1268 (
		\TM0_pad ,
		\_2167__reg/NET0131 ,
		_w2775_,
		_w2776_,
		_w2777_
	);
	LUT4 #(
		.INIT('h2772)
	) name1269 (
		\TM0_pad ,
		\WX10839_reg/NET0131 ,
		_w1880_,
		_w1881_,
		_w2778_
	);
	LUT4 #(
		.INIT('h028a)
	) name1270 (
		RESET_pad,
		\TM1_pad ,
		_w2777_,
		_w2778_,
		_w2779_
	);
	LUT4 #(
		.INIT('h8cc8)
	) name1271 (
		\TM0_pad ,
		_w1978_,
		_w2274_,
		_w2275_,
		_w2780_
	);
	LUT2 #(
		.INIT('h2)
	) name1272 (
		\TM0_pad ,
		\_2342__reg/NET0131 ,
		_w2781_
	);
	LUT4 #(
		.INIT('h00c8)
	) name1273 (
		\DATA_0_9_pad ,
		RESET_pad,
		\TM0_pad ,
		\TM1_pad ,
		_w2782_
	);
	LUT2 #(
		.INIT('h4)
	) name1274 (
		_w2781_,
		_w2782_,
		_w2783_
	);
	LUT2 #(
		.INIT('he)
	) name1275 (
		_w2780_,
		_w2783_,
		_w2784_
	);
	LUT2 #(
		.INIT('h8)
	) name1276 (
		RESET_pad,
		\WX10871_reg/NET0131 ,
		_w2785_
	);
	LUT3 #(
		.INIT('h96)
	) name1277 (
		\WX9764_reg/NET0131 ,
		\WX9828_reg/NET0131 ,
		\WX9892_reg/NET0131 ,
		_w2786_
	);
	LUT2 #(
		.INIT('h9)
	) name1278 (
		\TM1_pad ,
		\WX9700_reg/NET0131 ,
		_w2787_
	);
	LUT4 #(
		.INIT('h2772)
	) name1279 (
		\TM0_pad ,
		\_2298__reg/NET0131 ,
		_w2786_,
		_w2787_,
		_w2788_
	);
	LUT4 #(
		.INIT('h2772)
	) name1280 (
		\TM0_pad ,
		\WX10833_reg/NET0131 ,
		_w2770_,
		_w2771_,
		_w2789_
	);
	LUT4 #(
		.INIT('h028a)
	) name1281 (
		RESET_pad,
		\TM1_pad ,
		_w2788_,
		_w2789_,
		_w2790_
	);
	LUT4 #(
		.INIT('h2772)
	) name1282 (
		\TM0_pad ,
		\_2331__reg/NET0131 ,
		_w1699_,
		_w1700_,
		_w2791_
	);
	LUT4 #(
		.INIT('h2772)
	) name1283 (
		\TM0_pad ,
		\WX10831_reg/NET0131 ,
		_w2744_,
		_w2745_,
		_w2792_
	);
	LUT4 #(
		.INIT('h028a)
	) name1284 (
		RESET_pad,
		\TM1_pad ,
		_w2791_,
		_w2792_,
		_w2793_
	);
	LUT3 #(
		.INIT('h96)
	) name1285 (
		\WX5891_reg/NET0131 ,
		\WX5955_reg/NET0131 ,
		\WX6019_reg/NET0131 ,
		_w2794_
	);
	LUT2 #(
		.INIT('h9)
	) name1286 (
		\TM1_pad ,
		\WX5827_reg/NET0131 ,
		_w2795_
	);
	LUT4 #(
		.INIT('h2772)
	) name1287 (
		\TM0_pad ,
		\_2199__reg/NET0131 ,
		_w2794_,
		_w2795_,
		_w2796_
	);
	LUT4 #(
		.INIT('h2772)
	) name1288 (
		\TM0_pad ,
		\WX10839_reg/NET0131 ,
		_w2775_,
		_w2776_,
		_w2797_
	);
	LUT4 #(
		.INIT('h028a)
	) name1289 (
		RESET_pad,
		\TM1_pad ,
		_w2796_,
		_w2797_,
		_w2798_
	);
	LUT3 #(
		.INIT('h96)
	) name1290 (
		\WX7182_reg/NET0131 ,
		\WX7246_reg/NET0131 ,
		\WX7310_reg/NET0131 ,
		_w2799_
	);
	LUT2 #(
		.INIT('h9)
	) name1291 (
		\TM1_pad ,
		\WX7118_reg/NET0131 ,
		_w2800_
	);
	LUT4 #(
		.INIT('h2772)
	) name1292 (
		\TM0_pad ,
		\_2232__reg/NET0131 ,
		_w2799_,
		_w2800_,
		_w2801_
	);
	LUT4 #(
		.INIT('h2772)
	) name1293 (
		\TM0_pad ,
		\WX10837_reg/NET0131 ,
		_w2754_,
		_w2755_,
		_w2802_
	);
	LUT4 #(
		.INIT('h028a)
	) name1294 (
		RESET_pad,
		\TM1_pad ,
		_w2801_,
		_w2802_,
		_w2803_
	);
	LUT2 #(
		.INIT('h9)
	) name1295 (
		\WX2112_reg/NET0131 ,
		\WX2176_reg/NET0131 ,
		_w2804_
	);
	LUT2 #(
		.INIT('h9)
	) name1296 (
		\WX1984_reg/NET0131 ,
		\WX2048_reg/NET0131 ,
		_w2805_
	);
	LUT4 #(
		.INIT('h8cc8)
	) name1297 (
		\TM0_pad ,
		_w1620_,
		_w2804_,
		_w2805_,
		_w2806_
	);
	LUT4 #(
		.INIT('h0a02)
	) name1298 (
		RESET_pad,
		\TM0_pad ,
		\TM1_pad ,
		\_2117__reg/NET0131 ,
		_w2807_
	);
	LUT4 #(
		.INIT('hbe00)
	) name1299 (
		\TM0_pad ,
		_w2035_,
		_w2036_,
		_w2807_,
		_w2808_
	);
	LUT2 #(
		.INIT('he)
	) name1300 (
		_w2806_,
		_w2808_,
		_w2809_
	);
	LUT3 #(
		.INIT('h96)
	) name1301 (
		\WX8473_reg/NET0131 ,
		\WX8537_reg/NET0131 ,
		\WX8601_reg/NET0131 ,
		_w2810_
	);
	LUT2 #(
		.INIT('h9)
	) name1302 (
		\TM1_pad ,
		\WX8409_reg/NET0131 ,
		_w2811_
	);
	LUT4 #(
		.INIT('h2772)
	) name1303 (
		\TM0_pad ,
		\_2265__reg/NET0131 ,
		_w2810_,
		_w2811_,
		_w2812_
	);
	LUT4 #(
		.INIT('h2772)
	) name1304 (
		\TM0_pad ,
		\WX10835_reg/NET0131 ,
		_w2759_,
		_w2760_,
		_w2813_
	);
	LUT4 #(
		.INIT('h028a)
	) name1305 (
		RESET_pad,
		\TM1_pad ,
		_w2812_,
		_w2813_,
		_w2814_
	);
	LUT3 #(
		.INIT('h96)
	) name1306 (
		\WX4600_reg/NET0131 ,
		\WX4664_reg/NET0131 ,
		\WX4728_reg/NET0131 ,
		_w2815_
	);
	LUT2 #(
		.INIT('h9)
	) name1307 (
		\TM1_pad ,
		\WX4536_reg/NET0131 ,
		_w2816_
	);
	LUT4 #(
		.INIT('h2772)
	) name1308 (
		\TM0_pad ,
		\_2166__reg/NET0131 ,
		_w2815_,
		_w2816_,
		_w2817_
	);
	LUT4 #(
		.INIT('h2772)
	) name1309 (
		\TM0_pad ,
		\WX10841_reg/NET0131 ,
		_w1936_,
		_w1937_,
		_w2818_
	);
	LUT4 #(
		.INIT('h028a)
	) name1310 (
		RESET_pad,
		\TM1_pad ,
		_w2817_,
		_w2818_,
		_w2819_
	);
	LUT3 #(
		.INIT('he0)
	) name1311 (
		\TM0_pad ,
		_w1594_,
		_w2146_,
		_w2820_
	);
	LUT2 #(
		.INIT('h9)
	) name1312 (
		\WX2116_reg/NET0131 ,
		\WX2180_reg/NET0131 ,
		_w2821_
	);
	LUT2 #(
		.INIT('h9)
	) name1313 (
		\WX1988_reg/NET0131 ,
		\WX2052_reg/NET0131 ,
		_w2822_
	);
	LUT4 #(
		.INIT('h0a02)
	) name1314 (
		RESET_pad,
		\TM0_pad ,
		\TM1_pad ,
		\_2083__reg/NET0131 ,
		_w2823_
	);
	LUT4 #(
		.INIT('hbe00)
	) name1315 (
		\TM0_pad ,
		_w2821_,
		_w2822_,
		_w2823_,
		_w2824_
	);
	LUT2 #(
		.INIT('he)
	) name1316 (
		_w2820_,
		_w2824_,
		_w2825_
	);
	LUT2 #(
		.INIT('h8)
	) name1317 (
		RESET_pad,
		\WX10873_reg/NET0131 ,
		_w2826_
	);
	LUT4 #(
		.INIT('h2772)
	) name1318 (
		\TM0_pad ,
		\_2297__reg/NET0131 ,
		_w1613_,
		_w1614_,
		_w2827_
	);
	LUT4 #(
		.INIT('h2772)
	) name1319 (
		\TM0_pad ,
		\WX10835_reg/NET0131 ,
		_w2810_,
		_w2811_,
		_w2828_
	);
	LUT4 #(
		.INIT('h028a)
	) name1320 (
		RESET_pad,
		\TM1_pad ,
		_w2827_,
		_w2828_,
		_w2829_
	);
	LUT4 #(
		.INIT('h2772)
	) name1321 (
		\TM0_pad ,
		\_2330__reg/NET0131 ,
		_w1751_,
		_w1752_,
		_w2830_
	);
	LUT4 #(
		.INIT('h2772)
	) name1322 (
		\TM0_pad ,
		\WX10833_reg/NET0131 ,
		_w2786_,
		_w2787_,
		_w2831_
	);
	LUT4 #(
		.INIT('h028a)
	) name1323 (
		RESET_pad,
		\TM1_pad ,
		_w2830_,
		_w2831_,
		_w2832_
	);
	LUT3 #(
		.INIT('h96)
	) name1324 (
		\WX5893_reg/NET0131 ,
		\WX5957_reg/NET0131 ,
		\WX6021_reg/NET0131 ,
		_w2833_
	);
	LUT2 #(
		.INIT('h9)
	) name1325 (
		\TM1_pad ,
		\WX5829_reg/NET0131 ,
		_w2834_
	);
	LUT4 #(
		.INIT('h2772)
	) name1326 (
		\TM0_pad ,
		\_2198__reg/NET0131 ,
		_w2833_,
		_w2834_,
		_w2835_
	);
	LUT4 #(
		.INIT('h2772)
	) name1327 (
		\TM0_pad ,
		\WX10841_reg/NET0131 ,
		_w2815_,
		_w2816_,
		_w2836_
	);
	LUT4 #(
		.INIT('h028a)
	) name1328 (
		RESET_pad,
		\TM1_pad ,
		_w2835_,
		_w2836_,
		_w2837_
	);
	LUT3 #(
		.INIT('h96)
	) name1329 (
		\WX7184_reg/NET0131 ,
		\WX7248_reg/NET0131 ,
		\WX7312_reg/NET0131 ,
		_w2838_
	);
	LUT2 #(
		.INIT('h9)
	) name1330 (
		\TM1_pad ,
		\WX7120_reg/NET0131 ,
		_w2839_
	);
	LUT4 #(
		.INIT('h2772)
	) name1331 (
		\TM0_pad ,
		\_2231__reg/NET0131 ,
		_w2838_,
		_w2839_,
		_w2840_
	);
	LUT4 #(
		.INIT('h2772)
	) name1332 (
		\TM0_pad ,
		\WX10839_reg/NET0131 ,
		_w2794_,
		_w2795_,
		_w2841_
	);
	LUT4 #(
		.INIT('h028a)
	) name1333 (
		RESET_pad,
		\TM1_pad ,
		_w2840_,
		_w2841_,
		_w2842_
	);
	LUT2 #(
		.INIT('h9)
	) name1334 (
		\WX2114_reg/NET0131 ,
		\WX2178_reg/NET0131 ,
		_w2843_
	);
	LUT2 #(
		.INIT('h9)
	) name1335 (
		\WX1986_reg/NET0131 ,
		\WX2050_reg/NET0131 ,
		_w2844_
	);
	LUT4 #(
		.INIT('h8cc8)
	) name1336 (
		\TM0_pad ,
		_w2089_,
		_w2843_,
		_w2844_,
		_w2845_
	);
	LUT4 #(
		.INIT('h0a02)
	) name1337 (
		RESET_pad,
		\TM0_pad ,
		\TM1_pad ,
		\_2116__reg/NET0131 ,
		_w2846_
	);
	LUT4 #(
		.INIT('hbe00)
	) name1338 (
		\TM0_pad ,
		_w2090_,
		_w2091_,
		_w2846_,
		_w2847_
	);
	LUT2 #(
		.INIT('he)
	) name1339 (
		_w2845_,
		_w2847_,
		_w2848_
	);
	LUT3 #(
		.INIT('h96)
	) name1340 (
		\WX8475_reg/NET0131 ,
		\WX8539_reg/NET0131 ,
		\WX8603_reg/NET0131 ,
		_w2849_
	);
	LUT2 #(
		.INIT('h9)
	) name1341 (
		\TM1_pad ,
		\WX8411_reg/NET0131 ,
		_w2850_
	);
	LUT4 #(
		.INIT('h2772)
	) name1342 (
		\TM0_pad ,
		\_2264__reg/NET0131 ,
		_w2849_,
		_w2850_,
		_w2851_
	);
	LUT4 #(
		.INIT('h2772)
	) name1343 (
		\TM0_pad ,
		\WX10837_reg/NET0131 ,
		_w2799_,
		_w2800_,
		_w2852_
	);
	LUT4 #(
		.INIT('h028a)
	) name1344 (
		RESET_pad,
		\TM1_pad ,
		_w2851_,
		_w2852_,
		_w2853_
	);
	LUT3 #(
		.INIT('h96)
	) name1345 (
		\WX4602_reg/NET0131 ,
		\WX4666_reg/NET0131 ,
		\WX4730_reg/NET0131 ,
		_w2854_
	);
	LUT2 #(
		.INIT('h9)
	) name1346 (
		\TM1_pad ,
		\WX4538_reg/NET0131 ,
		_w2855_
	);
	LUT4 #(
		.INIT('h2772)
	) name1347 (
		\TM0_pad ,
		\_2165__reg/NET0131 ,
		_w2854_,
		_w2855_,
		_w2856_
	);
	LUT4 #(
		.INIT('h2772)
	) name1348 (
		\TM0_pad ,
		\WX10843_reg/NET0131 ,
		_w1999_,
		_w2000_,
		_w2857_
	);
	LUT4 #(
		.INIT('h028a)
	) name1349 (
		RESET_pad,
		\TM1_pad ,
		_w2856_,
		_w2857_,
		_w2858_
	);
	LUT3 #(
		.INIT('he0)
	) name1350 (
		\TM0_pad ,
		_w1591_,
		_w2203_,
		_w2859_
	);
	LUT2 #(
		.INIT('h9)
	) name1351 (
		\WX2118_reg/NET0131 ,
		\WX2182_reg/NET0131 ,
		_w2860_
	);
	LUT2 #(
		.INIT('h9)
	) name1352 (
		\WX1990_reg/NET0131 ,
		\WX2054_reg/NET0131 ,
		_w2861_
	);
	LUT4 #(
		.INIT('h0a02)
	) name1353 (
		RESET_pad,
		\TM0_pad ,
		\TM1_pad ,
		\_2082__reg/NET0131 ,
		_w2862_
	);
	LUT4 #(
		.INIT('hbe00)
	) name1354 (
		\TM0_pad ,
		_w2860_,
		_w2861_,
		_w2862_,
		_w2863_
	);
	LUT2 #(
		.INIT('he)
	) name1355 (
		_w2859_,
		_w2863_,
		_w2864_
	);
	LUT4 #(
		.INIT('h8cc8)
	) name1356 (
		\TM0_pad ,
		_w2089_,
		_w2382_,
		_w2383_,
		_w2865_
	);
	LUT2 #(
		.INIT('h2)
	) name1357 (
		\TM0_pad ,
		\_2340__reg/NET0131 ,
		_w2866_
	);
	LUT4 #(
		.INIT('h00c8)
	) name1358 (
		\DATA_0_7_pad ,
		RESET_pad,
		\TM0_pad ,
		\TM1_pad ,
		_w2867_
	);
	LUT2 #(
		.INIT('h4)
	) name1359 (
		_w2866_,
		_w2867_,
		_w2868_
	);
	LUT2 #(
		.INIT('he)
	) name1360 (
		_w2865_,
		_w2868_,
		_w2869_
	);
	LUT2 #(
		.INIT('h8)
	) name1361 (
		RESET_pad,
		\WX10875_reg/NET0131 ,
		_w2870_
	);
	LUT3 #(
		.INIT('h96)
	) name1362 (
		\WX9768_reg/NET0131 ,
		\WX9832_reg/NET0131 ,
		\WX9896_reg/NET0131 ,
		_w2871_
	);
	LUT2 #(
		.INIT('h9)
	) name1363 (
		\TM1_pad ,
		\WX9704_reg/NET0131 ,
		_w2872_
	);
	LUT4 #(
		.INIT('h2772)
	) name1364 (
		\TM0_pad ,
		\_2296__reg/NET0131 ,
		_w2871_,
		_w2872_,
		_w2873_
	);
	LUT4 #(
		.INIT('h2772)
	) name1365 (
		\TM0_pad ,
		\WX10837_reg/NET0131 ,
		_w2849_,
		_w2850_,
		_w2874_
	);
	LUT4 #(
		.INIT('h028a)
	) name1366 (
		RESET_pad,
		\TM1_pad ,
		_w2873_,
		_w2874_,
		_w2875_
	);
	LUT3 #(
		.INIT('h96)
	) name1367 (
		\WX5895_reg/NET0131 ,
		\WX5959_reg/NET0131 ,
		\WX6023_reg/NET0131 ,
		_w2876_
	);
	LUT2 #(
		.INIT('h9)
	) name1368 (
		\TM1_pad ,
		\WX5831_reg/NET0131 ,
		_w2877_
	);
	LUT4 #(
		.INIT('h2772)
	) name1369 (
		\TM0_pad ,
		\_2197__reg/NET0131 ,
		_w2876_,
		_w2877_,
		_w2878_
	);
	LUT4 #(
		.INIT('h2772)
	) name1370 (
		\TM0_pad ,
		\WX10843_reg/NET0131 ,
		_w2854_,
		_w2855_,
		_w2879_
	);
	LUT4 #(
		.INIT('h028a)
	) name1371 (
		RESET_pad,
		\TM1_pad ,
		_w2878_,
		_w2879_,
		_w2880_
	);
	LUT3 #(
		.INIT('h96)
	) name1372 (
		\WX7186_reg/NET0131 ,
		\WX7250_reg/NET0131 ,
		\WX7314_reg/NET0131 ,
		_w2881_
	);
	LUT2 #(
		.INIT('h9)
	) name1373 (
		\TM1_pad ,
		\WX7122_reg/NET0131 ,
		_w2882_
	);
	LUT4 #(
		.INIT('h2772)
	) name1374 (
		\TM0_pad ,
		\_2230__reg/NET0131 ,
		_w2881_,
		_w2882_,
		_w2883_
	);
	LUT4 #(
		.INIT('h2772)
	) name1375 (
		\TM0_pad ,
		\WX10841_reg/NET0131 ,
		_w2833_,
		_w2834_,
		_w2884_
	);
	LUT4 #(
		.INIT('h028a)
	) name1376 (
		RESET_pad,
		\TM1_pad ,
		_w2883_,
		_w2884_,
		_w2885_
	);
	LUT4 #(
		.INIT('h8cc8)
	) name1377 (
		\TM0_pad ,
		_w2146_,
		_w2821_,
		_w2822_,
		_w2886_
	);
	LUT4 #(
		.INIT('h0a02)
	) name1378 (
		RESET_pad,
		\TM0_pad ,
		\TM1_pad ,
		\_2115__reg/NET0131 ,
		_w2887_
	);
	LUT4 #(
		.INIT('hbe00)
	) name1379 (
		\TM0_pad ,
		_w2147_,
		_w2148_,
		_w2887_,
		_w2888_
	);
	LUT2 #(
		.INIT('he)
	) name1380 (
		_w2886_,
		_w2888_,
		_w2889_
	);
	LUT3 #(
		.INIT('h96)
	) name1381 (
		\WX8477_reg/NET0131 ,
		\WX8541_reg/NET0131 ,
		\WX8605_reg/NET0131 ,
		_w2890_
	);
	LUT2 #(
		.INIT('h9)
	) name1382 (
		\TM1_pad ,
		\WX8413_reg/NET0131 ,
		_w2891_
	);
	LUT4 #(
		.INIT('h2772)
	) name1383 (
		\TM0_pad ,
		\_2263__reg/NET0131 ,
		_w2890_,
		_w2891_,
		_w2892_
	);
	LUT4 #(
		.INIT('h2772)
	) name1384 (
		\TM0_pad ,
		\WX10839_reg/NET0131 ,
		_w2838_,
		_w2839_,
		_w2893_
	);
	LUT4 #(
		.INIT('h028a)
	) name1385 (
		RESET_pad,
		\TM1_pad ,
		_w2892_,
		_w2893_,
		_w2894_
	);
	LUT3 #(
		.INIT('h96)
	) name1386 (
		\WX4604_reg/NET0131 ,
		\WX4668_reg/NET0131 ,
		\WX4732_reg/NET0131 ,
		_w2895_
	);
	LUT2 #(
		.INIT('h9)
	) name1387 (
		\TM1_pad ,
		\WX4540_reg/NET0131 ,
		_w2896_
	);
	LUT4 #(
		.INIT('h2772)
	) name1388 (
		\TM0_pad ,
		\_2164__reg/NET0131 ,
		_w2895_,
		_w2896_,
		_w2897_
	);
	LUT4 #(
		.INIT('h2772)
	) name1389 (
		\TM0_pad ,
		\WX10845_reg/NET0131 ,
		_w2053_,
		_w2054_,
		_w2898_
	);
	LUT4 #(
		.INIT('h028a)
	) name1390 (
		RESET_pad,
		\TM1_pad ,
		_w2897_,
		_w2898_,
		_w2899_
	);
	LUT4 #(
		.INIT('h2772)
	) name1391 (
		\TM0_pad ,
		\WX10829_reg/NET0131 ,
		_w1581_,
		_w1582_,
		_w2900_
	);
	LUT3 #(
		.INIT('h69)
	) name1392 (
		\TM1_pad ,
		\WX1938_reg/NET0131 ,
		\WX2002_reg/NET0131 ,
		_w2901_
	);
	LUT2 #(
		.INIT('h9)
	) name1393 (
		\WX2066_reg/NET0131 ,
		\WX2130_reg/NET0131 ,
		_w2902_
	);
	LUT4 #(
		.INIT('h7227)
	) name1394 (
		\TM0_pad ,
		\_2108__reg/NET0131 ,
		_w2901_,
		_w2902_,
		_w2903_
	);
	LUT4 #(
		.INIT('h082a)
	) name1395 (
		RESET_pad,
		\TM1_pad ,
		_w2900_,
		_w2903_,
		_w2904_
	);
	LUT4 #(
		.INIT('h8cc8)
	) name1396 (
		\TM0_pad ,
		_w2146_,
		_w2438_,
		_w2439_,
		_w2905_
	);
	LUT2 #(
		.INIT('h2)
	) name1397 (
		\TM0_pad ,
		\_2339__reg/NET0131 ,
		_w2906_
	);
	LUT4 #(
		.INIT('h00c8)
	) name1398 (
		\DATA_0_6_pad ,
		RESET_pad,
		\TM0_pad ,
		\TM1_pad ,
		_w2907_
	);
	LUT2 #(
		.INIT('h4)
	) name1399 (
		_w2906_,
		_w2907_,
		_w2908_
	);
	LUT2 #(
		.INIT('he)
	) name1400 (
		_w2905_,
		_w2908_,
		_w2909_
	);
	LUT2 #(
		.INIT('h8)
	) name1401 (
		RESET_pad,
		\WX10877_reg/NET0131 ,
		_w2910_
	);
	LUT3 #(
		.INIT('h96)
	) name1402 (
		\WX4606_reg/NET0131 ,
		\WX4670_reg/NET0131 ,
		\WX4734_reg/NET0131 ,
		_w2911_
	);
	LUT2 #(
		.INIT('h9)
	) name1403 (
		\TM1_pad ,
		\WX4542_reg/NET0131 ,
		_w2912_
	);
	LUT4 #(
		.INIT('h2772)
	) name1404 (
		\TM0_pad ,
		\_2163__reg/NET0131 ,
		_w2911_,
		_w2912_,
		_w2913_
	);
	LUT4 #(
		.INIT('h2772)
	) name1405 (
		\TM0_pad ,
		\WX10847_reg/NET0131 ,
		_w2110_,
		_w2111_,
		_w2914_
	);
	LUT4 #(
		.INIT('h028a)
	) name1406 (
		RESET_pad,
		\TM1_pad ,
		_w2913_,
		_w2914_,
		_w2915_
	);
	LUT3 #(
		.INIT('h96)
	) name1407 (
		\WX9770_reg/NET0131 ,
		\WX9834_reg/NET0131 ,
		\WX9898_reg/NET0131 ,
		_w2916_
	);
	LUT2 #(
		.INIT('h9)
	) name1408 (
		\TM1_pad ,
		\WX9706_reg/NET0131 ,
		_w2917_
	);
	LUT4 #(
		.INIT('h2772)
	) name1409 (
		\TM0_pad ,
		\_2295__reg/NET0131 ,
		_w2916_,
		_w2917_,
		_w2918_
	);
	LUT4 #(
		.INIT('h2772)
	) name1410 (
		\TM0_pad ,
		\WX10839_reg/NET0131 ,
		_w2890_,
		_w2891_,
		_w2919_
	);
	LUT4 #(
		.INIT('h028a)
	) name1411 (
		RESET_pad,
		\TM1_pad ,
		_w2918_,
		_w2919_,
		_w2920_
	);
	LUT4 #(
		.INIT('h2772)
	) name1412 (
		\TM0_pad ,
		\_2328__reg/NET0131 ,
		_w1857_,
		_w1858_,
		_w2921_
	);
	LUT4 #(
		.INIT('h2772)
	) name1413 (
		\TM0_pad ,
		\WX10837_reg/NET0131 ,
		_w2871_,
		_w2872_,
		_w2922_
	);
	LUT4 #(
		.INIT('h028a)
	) name1414 (
		RESET_pad,
		\TM1_pad ,
		_w2921_,
		_w2922_,
		_w2923_
	);
	LUT3 #(
		.INIT('h96)
	) name1415 (
		\WX5897_reg/NET0131 ,
		\WX5961_reg/NET0131 ,
		\WX6025_reg/NET0131 ,
		_w2924_
	);
	LUT2 #(
		.INIT('h9)
	) name1416 (
		\TM1_pad ,
		\WX5833_reg/NET0131 ,
		_w2925_
	);
	LUT4 #(
		.INIT('h2772)
	) name1417 (
		\TM0_pad ,
		\_2196__reg/NET0131 ,
		_w2924_,
		_w2925_,
		_w2926_
	);
	LUT4 #(
		.INIT('h2772)
	) name1418 (
		\TM0_pad ,
		\WX10845_reg/NET0131 ,
		_w2895_,
		_w2896_,
		_w2927_
	);
	LUT4 #(
		.INIT('h028a)
	) name1419 (
		RESET_pad,
		\TM1_pad ,
		_w2926_,
		_w2927_,
		_w2928_
	);
	LUT3 #(
		.INIT('h96)
	) name1420 (
		\WX7188_reg/NET0131 ,
		\WX7252_reg/NET0131 ,
		\WX7316_reg/NET0131 ,
		_w2929_
	);
	LUT2 #(
		.INIT('h9)
	) name1421 (
		\TM1_pad ,
		\WX7124_reg/NET0131 ,
		_w2930_
	);
	LUT4 #(
		.INIT('h2772)
	) name1422 (
		\TM0_pad ,
		\_2229__reg/NET0131 ,
		_w2929_,
		_w2930_,
		_w2931_
	);
	LUT4 #(
		.INIT('h2772)
	) name1423 (
		\TM0_pad ,
		\WX10843_reg/NET0131 ,
		_w2876_,
		_w2877_,
		_w2932_
	);
	LUT4 #(
		.INIT('h028a)
	) name1424 (
		RESET_pad,
		\TM1_pad ,
		_w2931_,
		_w2932_,
		_w2933_
	);
	LUT4 #(
		.INIT('h8cc8)
	) name1425 (
		\TM0_pad ,
		_w2203_,
		_w2860_,
		_w2861_,
		_w2934_
	);
	LUT4 #(
		.INIT('h0a02)
	) name1426 (
		RESET_pad,
		\TM0_pad ,
		\TM1_pad ,
		\_2114__reg/NET0131 ,
		_w2935_
	);
	LUT4 #(
		.INIT('hbe00)
	) name1427 (
		\TM0_pad ,
		_w2204_,
		_w2205_,
		_w2935_,
		_w2936_
	);
	LUT2 #(
		.INIT('he)
	) name1428 (
		_w2934_,
		_w2936_,
		_w2937_
	);
	LUT3 #(
		.INIT('h96)
	) name1429 (
		\WX8479_reg/NET0131 ,
		\WX8543_reg/NET0131 ,
		\WX8607_reg/NET0131 ,
		_w2938_
	);
	LUT2 #(
		.INIT('h9)
	) name1430 (
		\TM1_pad ,
		\WX8415_reg/NET0131 ,
		_w2939_
	);
	LUT4 #(
		.INIT('h2772)
	) name1431 (
		\TM0_pad ,
		\_2262__reg/NET0131 ,
		_w2938_,
		_w2939_,
		_w2940_
	);
	LUT4 #(
		.INIT('h2772)
	) name1432 (
		\TM0_pad ,
		\WX10841_reg/NET0131 ,
		_w2881_,
		_w2882_,
		_w2941_
	);
	LUT4 #(
		.INIT('h028a)
	) name1433 (
		RESET_pad,
		\TM1_pad ,
		_w2940_,
		_w2941_,
		_w2942_
	);
	LUT3 #(
		.INIT('he0)
	) name1434 (
		\TM0_pad ,
		_w1585_,
		_w2313_,
		_w2943_
	);
	LUT2 #(
		.INIT('h9)
	) name1435 (
		\WX2122_reg/NET0131 ,
		\WX2186_reg/NET0131 ,
		_w2944_
	);
	LUT2 #(
		.INIT('h9)
	) name1436 (
		\WX1994_reg/NET0131 ,
		\WX2058_reg/NET0131 ,
		_w2945_
	);
	LUT4 #(
		.INIT('h0a02)
	) name1437 (
		RESET_pad,
		\TM0_pad ,
		\TM1_pad ,
		\_2080__reg/NET0131 ,
		_w2946_
	);
	LUT4 #(
		.INIT('hbe00)
	) name1438 (
		\TM0_pad ,
		_w2944_,
		_w2945_,
		_w2946_,
		_w2947_
	);
	LUT2 #(
		.INIT('he)
	) name1439 (
		_w2943_,
		_w2947_,
		_w2948_
	);
	LUT4 #(
		.INIT('h8cc8)
	) name1440 (
		\TM0_pad ,
		_w2203_,
		_w2488_,
		_w2489_,
		_w2949_
	);
	LUT2 #(
		.INIT('h2)
	) name1441 (
		\TM0_pad ,
		\_2338__reg/NET0131 ,
		_w2950_
	);
	LUT4 #(
		.INIT('h00c8)
	) name1442 (
		\DATA_0_5_pad ,
		RESET_pad,
		\TM0_pad ,
		\TM1_pad ,
		_w2951_
	);
	LUT2 #(
		.INIT('h4)
	) name1443 (
		_w2950_,
		_w2951_,
		_w2952_
	);
	LUT2 #(
		.INIT('he)
	) name1444 (
		_w2949_,
		_w2952_,
		_w2953_
	);
	LUT2 #(
		.INIT('h8)
	) name1445 (
		RESET_pad,
		\WX10879_reg/NET0131 ,
		_w2954_
	);
	LUT3 #(
		.INIT('h96)
	) name1446 (
		\WX4608_reg/NET0131 ,
		\WX4672_reg/NET0131 ,
		\WX4736_reg/NET0131 ,
		_w2955_
	);
	LUT2 #(
		.INIT('h9)
	) name1447 (
		\TM1_pad ,
		\WX4544_reg/NET0131 ,
		_w2956_
	);
	LUT4 #(
		.INIT('h2772)
	) name1448 (
		\TM0_pad ,
		\_2162__reg/NET0131 ,
		_w2955_,
		_w2956_,
		_w2957_
	);
	LUT4 #(
		.INIT('h2772)
	) name1449 (
		\TM0_pad ,
		\WX10849_reg/NET0131 ,
		_w2167_,
		_w2168_,
		_w2958_
	);
	LUT4 #(
		.INIT('h028a)
	) name1450 (
		RESET_pad,
		\TM1_pad ,
		_w2957_,
		_w2958_,
		_w2959_
	);
	LUT3 #(
		.INIT('h96)
	) name1451 (
		\WX9772_reg/NET0131 ,
		\WX9836_reg/NET0131 ,
		\WX9900_reg/NET0131 ,
		_w2960_
	);
	LUT2 #(
		.INIT('h9)
	) name1452 (
		\TM1_pad ,
		\WX9708_reg/NET0131 ,
		_w2961_
	);
	LUT4 #(
		.INIT('h2772)
	) name1453 (
		\TM0_pad ,
		\_2294__reg/NET0131 ,
		_w2960_,
		_w2961_,
		_w2962_
	);
	LUT4 #(
		.INIT('h2772)
	) name1454 (
		\TM0_pad ,
		\WX10841_reg/NET0131 ,
		_w2938_,
		_w2939_,
		_w2963_
	);
	LUT4 #(
		.INIT('h028a)
	) name1455 (
		RESET_pad,
		\TM1_pad ,
		_w2962_,
		_w2963_,
		_w2964_
	);
	LUT4 #(
		.INIT('h2772)
	) name1456 (
		\TM0_pad ,
		\_2140__reg/NET0131 ,
		_w2555_,
		_w2556_,
		_w2965_
	);
	LUT4 #(
		.INIT('h7227)
	) name1457 (
		\TM0_pad ,
		\WX10829_reg/NET0131 ,
		_w2901_,
		_w2902_,
		_w2966_
	);
	LUT4 #(
		.INIT('h028a)
	) name1458 (
		RESET_pad,
		\TM1_pad ,
		_w2965_,
		_w2966_,
		_w2967_
	);
	LUT4 #(
		.INIT('h2772)
	) name1459 (
		\TM0_pad ,
		\_2327__reg/NET0131 ,
		_w1913_,
		_w1914_,
		_w2968_
	);
	LUT4 #(
		.INIT('h2772)
	) name1460 (
		\TM0_pad ,
		\WX10839_reg/NET0131 ,
		_w2916_,
		_w2917_,
		_w2969_
	);
	LUT4 #(
		.INIT('h028a)
	) name1461 (
		RESET_pad,
		\TM1_pad ,
		_w2968_,
		_w2969_,
		_w2970_
	);
	LUT3 #(
		.INIT('h96)
	) name1462 (
		\WX5899_reg/NET0131 ,
		\WX5963_reg/NET0131 ,
		\WX6027_reg/NET0131 ,
		_w2971_
	);
	LUT2 #(
		.INIT('h9)
	) name1463 (
		\TM1_pad ,
		\WX5835_reg/NET0131 ,
		_w2972_
	);
	LUT4 #(
		.INIT('h2772)
	) name1464 (
		\TM0_pad ,
		\_2195__reg/NET0131 ,
		_w2971_,
		_w2972_,
		_w2973_
	);
	LUT4 #(
		.INIT('h2772)
	) name1465 (
		\TM0_pad ,
		\WX10847_reg/NET0131 ,
		_w2911_,
		_w2912_,
		_w2974_
	);
	LUT4 #(
		.INIT('h028a)
	) name1466 (
		RESET_pad,
		\TM1_pad ,
		_w2973_,
		_w2974_,
		_w2975_
	);
	LUT3 #(
		.INIT('h96)
	) name1467 (
		\WX7190_reg/NET0131 ,
		\WX7254_reg/NET0131 ,
		\WX7318_reg/NET0131 ,
		_w2976_
	);
	LUT2 #(
		.INIT('h9)
	) name1468 (
		\TM1_pad ,
		\WX7126_reg/NET0131 ,
		_w2977_
	);
	LUT4 #(
		.INIT('h2772)
	) name1469 (
		\TM0_pad ,
		\_2228__reg/NET0131 ,
		_w2976_,
		_w2977_,
		_w2978_
	);
	LUT4 #(
		.INIT('h2772)
	) name1470 (
		\TM0_pad ,
		\WX10845_reg/NET0131 ,
		_w2924_,
		_w2925_,
		_w2979_
	);
	LUT4 #(
		.INIT('h028a)
	) name1471 (
		RESET_pad,
		\TM1_pad ,
		_w2978_,
		_w2979_,
		_w2980_
	);
	LUT2 #(
		.INIT('h9)
	) name1472 (
		\WX2120_reg/NET0131 ,
		\WX2184_reg/NET0131 ,
		_w2981_
	);
	LUT2 #(
		.INIT('h9)
	) name1473 (
		\WX1992_reg/NET0131 ,
		\WX2056_reg/NET0131 ,
		_w2982_
	);
	LUT4 #(
		.INIT('h8cc8)
	) name1474 (
		\TM0_pad ,
		_w2258_,
		_w2981_,
		_w2982_,
		_w2983_
	);
	LUT4 #(
		.INIT('h0a02)
	) name1475 (
		RESET_pad,
		\TM0_pad ,
		\TM1_pad ,
		\_2113__reg/NET0131 ,
		_w2984_
	);
	LUT4 #(
		.INIT('hbe00)
	) name1476 (
		\TM0_pad ,
		_w2259_,
		_w2260_,
		_w2984_,
		_w2985_
	);
	LUT2 #(
		.INIT('he)
	) name1477 (
		_w2983_,
		_w2985_,
		_w2986_
	);
	LUT3 #(
		.INIT('h96)
	) name1478 (
		\WX8481_reg/NET0131 ,
		\WX8545_reg/NET0131 ,
		\WX8609_reg/NET0131 ,
		_w2987_
	);
	LUT2 #(
		.INIT('h9)
	) name1479 (
		\TM1_pad ,
		\WX8417_reg/NET0131 ,
		_w2988_
	);
	LUT4 #(
		.INIT('h2772)
	) name1480 (
		\TM0_pad ,
		\_2261__reg/NET0131 ,
		_w2987_,
		_w2988_,
		_w2989_
	);
	LUT4 #(
		.INIT('h2772)
	) name1481 (
		\TM0_pad ,
		\WX10843_reg/NET0131 ,
		_w2929_,
		_w2930_,
		_w2990_
	);
	LUT4 #(
		.INIT('h028a)
	) name1482 (
		RESET_pad,
		\TM1_pad ,
		_w2989_,
		_w2990_,
		_w2991_
	);
	LUT3 #(
		.INIT('he0)
	) name1483 (
		\TM0_pad ,
		_w1576_,
		_w2366_,
		_w2992_
	);
	LUT2 #(
		.INIT('h9)
	) name1484 (
		\WX2124_reg/NET0131 ,
		\WX2188_reg/NET0131 ,
		_w2993_
	);
	LUT2 #(
		.INIT('h9)
	) name1485 (
		\WX1996_reg/NET0131 ,
		\WX2060_reg/NET0131 ,
		_w2994_
	);
	LUT4 #(
		.INIT('h0a02)
	) name1486 (
		RESET_pad,
		\TM0_pad ,
		\TM1_pad ,
		\_2079__reg/NET0131 ,
		_w2995_
	);
	LUT4 #(
		.INIT('hbe00)
	) name1487 (
		\TM0_pad ,
		_w2993_,
		_w2994_,
		_w2995_,
		_w2996_
	);
	LUT2 #(
		.INIT('he)
	) name1488 (
		_w2992_,
		_w2996_,
		_w2997_
	);
	LUT3 #(
		.INIT('he0)
	) name1489 (
		\TM0_pad ,
		_w1510_,
		_w2472_,
		_w2998_
	);
	LUT2 #(
		.INIT('h9)
	) name1490 (
		\WX2128_reg/NET0131 ,
		\WX2192_reg/NET0131 ,
		_w2999_
	);
	LUT2 #(
		.INIT('h9)
	) name1491 (
		\WX2000_reg/NET0131 ,
		\WX2064_reg/NET0131 ,
		_w3000_
	);
	LUT4 #(
		.INIT('h0a02)
	) name1492 (
		RESET_pad,
		\TM0_pad ,
		\TM1_pad ,
		\_2077__reg/NET0131 ,
		_w3001_
	);
	LUT4 #(
		.INIT('hbe00)
	) name1493 (
		\TM0_pad ,
		_w2999_,
		_w3000_,
		_w3001_,
		_w3002_
	);
	LUT2 #(
		.INIT('he)
	) name1494 (
		_w2998_,
		_w3002_,
		_w3003_
	);
	LUT4 #(
		.INIT('h7227)
	) name1495 (
		\TM0_pad ,
		\WX10829_reg/NET0131 ,
		_w2749_,
		_w2750_,
		_w3004_
	);
	LUT2 #(
		.INIT('h2)
	) name1496 (
		\TM0_pad ,
		\_2364__reg/NET0131 ,
		_w3005_
	);
	LUT4 #(
		.INIT('h00c8)
	) name1497 (
		\DATA_0_31_pad ,
		RESET_pad,
		\TM0_pad ,
		\TM1_pad ,
		_w3006_
	);
	LUT2 #(
		.INIT('h4)
	) name1498 (
		_w3005_,
		_w3006_,
		_w3007_
	);
	LUT3 #(
		.INIT('hf2)
	) name1499 (
		_w1605_,
		_w3004_,
		_w3007_,
		_w3008_
	);
	LUT4 #(
		.INIT('h8cc8)
	) name1500 (
		\TM0_pad ,
		_w2258_,
		_w2529_,
		_w2530_,
		_w3009_
	);
	LUT2 #(
		.INIT('h2)
	) name1501 (
		\TM0_pad ,
		\_2337__reg/NET0131 ,
		_w3010_
	);
	LUT4 #(
		.INIT('h00c8)
	) name1502 (
		\DATA_0_4_pad ,
		RESET_pad,
		\TM0_pad ,
		\TM1_pad ,
		_w3011_
	);
	LUT2 #(
		.INIT('h4)
	) name1503 (
		_w3010_,
		_w3011_,
		_w3012_
	);
	LUT2 #(
		.INIT('he)
	) name1504 (
		_w3009_,
		_w3012_,
		_w3013_
	);
	LUT2 #(
		.INIT('h8)
	) name1505 (
		RESET_pad,
		\WX10881_reg/NET0131 ,
		_w3014_
	);
	LUT3 #(
		.INIT('h96)
	) name1506 (
		\WX4610_reg/NET0131 ,
		\WX4674_reg/NET0131 ,
		\WX4738_reg/NET0131 ,
		_w3015_
	);
	LUT2 #(
		.INIT('h9)
	) name1507 (
		\TM1_pad ,
		\WX4546_reg/NET0131 ,
		_w3016_
	);
	LUT4 #(
		.INIT('h2772)
	) name1508 (
		\TM0_pad ,
		\_2161__reg/NET0131 ,
		_w3015_,
		_w3016_,
		_w3017_
	);
	LUT4 #(
		.INIT('h2772)
	) name1509 (
		\TM0_pad ,
		\WX10851_reg/NET0131 ,
		_w2224_,
		_w2225_,
		_w3018_
	);
	LUT4 #(
		.INIT('h028a)
	) name1510 (
		RESET_pad,
		\TM1_pad ,
		_w3017_,
		_w3018_,
		_w3019_
	);
	LUT3 #(
		.INIT('h96)
	) name1511 (
		\WX9774_reg/NET0131 ,
		\WX9838_reg/NET0131 ,
		\WX9902_reg/NET0131 ,
		_w3020_
	);
	LUT2 #(
		.INIT('h9)
	) name1512 (
		\TM1_pad ,
		\WX9710_reg/NET0131 ,
		_w3021_
	);
	LUT4 #(
		.INIT('h2772)
	) name1513 (
		\TM0_pad ,
		\_2293__reg/NET0131 ,
		_w3020_,
		_w3021_,
		_w3022_
	);
	LUT4 #(
		.INIT('h2772)
	) name1514 (
		\TM0_pad ,
		\WX10843_reg/NET0131 ,
		_w2987_,
		_w2988_,
		_w3023_
	);
	LUT4 #(
		.INIT('h028a)
	) name1515 (
		RESET_pad,
		\TM1_pad ,
		_w3022_,
		_w3023_,
		_w3024_
	);
	LUT4 #(
		.INIT('h2772)
	) name1516 (
		\TM0_pad ,
		\_2326__reg/NET0131 ,
		_w1970_,
		_w1971_,
		_w3025_
	);
	LUT4 #(
		.INIT('h2772)
	) name1517 (
		\TM0_pad ,
		\WX10841_reg/NET0131 ,
		_w2960_,
		_w2961_,
		_w3026_
	);
	LUT4 #(
		.INIT('h028a)
	) name1518 (
		RESET_pad,
		\TM1_pad ,
		_w3025_,
		_w3026_,
		_w3027_
	);
	LUT3 #(
		.INIT('h96)
	) name1519 (
		\WX5901_reg/NET0131 ,
		\WX5965_reg/NET0131 ,
		\WX6029_reg/NET0131 ,
		_w3028_
	);
	LUT2 #(
		.INIT('h9)
	) name1520 (
		\TM1_pad ,
		\WX5837_reg/NET0131 ,
		_w3029_
	);
	LUT4 #(
		.INIT('h2772)
	) name1521 (
		\TM0_pad ,
		\_2194__reg/NET0131 ,
		_w3028_,
		_w3029_,
		_w3030_
	);
	LUT4 #(
		.INIT('h2772)
	) name1522 (
		\TM0_pad ,
		\WX10849_reg/NET0131 ,
		_w2955_,
		_w2956_,
		_w3031_
	);
	LUT4 #(
		.INIT('h028a)
	) name1523 (
		RESET_pad,
		\TM1_pad ,
		_w3030_,
		_w3031_,
		_w3032_
	);
	LUT3 #(
		.INIT('h96)
	) name1524 (
		\WX7192_reg/NET0131 ,
		\WX7256_reg/NET0131 ,
		\WX7320_reg/NET0131 ,
		_w3033_
	);
	LUT2 #(
		.INIT('h9)
	) name1525 (
		\TM1_pad ,
		\WX7128_reg/NET0131 ,
		_w3034_
	);
	LUT4 #(
		.INIT('h2772)
	) name1526 (
		\TM0_pad ,
		\_2227__reg/NET0131 ,
		_w3033_,
		_w3034_,
		_w3035_
	);
	LUT4 #(
		.INIT('h2772)
	) name1527 (
		\TM0_pad ,
		\WX10847_reg/NET0131 ,
		_w2971_,
		_w2972_,
		_w3036_
	);
	LUT4 #(
		.INIT('h028a)
	) name1528 (
		RESET_pad,
		\TM1_pad ,
		_w3035_,
		_w3036_,
		_w3037_
	);
	LUT4 #(
		.INIT('h8cc8)
	) name1529 (
		\TM0_pad ,
		_w2313_,
		_w2944_,
		_w2945_,
		_w3038_
	);
	LUT4 #(
		.INIT('h0a02)
	) name1530 (
		RESET_pad,
		\TM0_pad ,
		\TM1_pad ,
		\_2112__reg/NET0131 ,
		_w3039_
	);
	LUT4 #(
		.INIT('hbe00)
	) name1531 (
		\TM0_pad ,
		_w2314_,
		_w2315_,
		_w3039_,
		_w3040_
	);
	LUT2 #(
		.INIT('he)
	) name1532 (
		_w3038_,
		_w3040_,
		_w3041_
	);
	LUT3 #(
		.INIT('h96)
	) name1533 (
		\WX8483_reg/NET0131 ,
		\WX8547_reg/NET0131 ,
		\WX8611_reg/NET0131 ,
		_w3042_
	);
	LUT2 #(
		.INIT('h9)
	) name1534 (
		\TM1_pad ,
		\WX8419_reg/NET0131 ,
		_w3043_
	);
	LUT4 #(
		.INIT('h2772)
	) name1535 (
		\TM0_pad ,
		\_2260__reg/NET0131 ,
		_w3042_,
		_w3043_,
		_w3044_
	);
	LUT4 #(
		.INIT('h2772)
	) name1536 (
		\TM0_pad ,
		\WX10845_reg/NET0131 ,
		_w2976_,
		_w2977_,
		_w3045_
	);
	LUT4 #(
		.INIT('h028a)
	) name1537 (
		RESET_pad,
		\TM1_pad ,
		_w3044_,
		_w3045_,
		_w3046_
	);
	LUT4 #(
		.INIT('h8cc8)
	) name1538 (
		\TM0_pad ,
		_w2313_,
		_w2589_,
		_w2590_,
		_w3047_
	);
	LUT2 #(
		.INIT('h2)
	) name1539 (
		\TM0_pad ,
		\_2336__reg/NET0131 ,
		_w3048_
	);
	LUT4 #(
		.INIT('h00c8)
	) name1540 (
		\DATA_0_3_pad ,
		RESET_pad,
		\TM0_pad ,
		\TM1_pad ,
		_w3049_
	);
	LUT2 #(
		.INIT('h4)
	) name1541 (
		_w3048_,
		_w3049_,
		_w3050_
	);
	LUT2 #(
		.INIT('he)
	) name1542 (
		_w3047_,
		_w3050_,
		_w3051_
	);
	LUT2 #(
		.INIT('h8)
	) name1543 (
		RESET_pad,
		\WX10883_reg/NET0131 ,
		_w3052_
	);
	LUT3 #(
		.INIT('h69)
	) name1544 (
		\TM1_pad ,
		\WX4548_reg/NET0131 ,
		\WX4612_reg/NET0131 ,
		_w3053_
	);
	LUT2 #(
		.INIT('h9)
	) name1545 (
		\WX4676_reg/NET0131 ,
		\WX4740_reg/NET0131 ,
		_w3054_
	);
	LUT4 #(
		.INIT('h7227)
	) name1546 (
		\TM0_pad ,
		\_2160__reg/NET0131 ,
		_w3053_,
		_w3054_,
		_w3055_
	);
	LUT4 #(
		.INIT('h2772)
	) name1547 (
		\TM0_pad ,
		\WX10853_reg/NET0131 ,
		_w2279_,
		_w2280_,
		_w3056_
	);
	LUT4 #(
		.INIT('h028a)
	) name1548 (
		RESET_pad,
		\TM1_pad ,
		_w3055_,
		_w3056_,
		_w3057_
	);
	LUT3 #(
		.INIT('h96)
	) name1549 (
		\WX4614_reg/NET0131 ,
		\WX4678_reg/NET0131 ,
		\WX4742_reg/NET0131 ,
		_w3058_
	);
	LUT2 #(
		.INIT('h9)
	) name1550 (
		\TM1_pad ,
		\WX4550_reg/NET0131 ,
		_w3059_
	);
	LUT4 #(
		.INIT('h2772)
	) name1551 (
		\TM0_pad ,
		\_2159__reg/NET0131 ,
		_w3058_,
		_w3059_,
		_w3060_
	);
	LUT4 #(
		.INIT('h2772)
	) name1552 (
		\TM0_pad ,
		\WX10855_reg/NET0131 ,
		_w2332_,
		_w2333_,
		_w3061_
	);
	LUT4 #(
		.INIT('h028a)
	) name1553 (
		RESET_pad,
		\TM1_pad ,
		_w3060_,
		_w3061_,
		_w3062_
	);
	LUT3 #(
		.INIT('h96)
	) name1554 (
		\WX4616_reg/NET0131 ,
		\WX4680_reg/NET0131 ,
		\WX4744_reg/NET0131 ,
		_w3063_
	);
	LUT2 #(
		.INIT('h9)
	) name1555 (
		\TM1_pad ,
		\WX4552_reg/NET0131 ,
		_w3064_
	);
	LUT4 #(
		.INIT('h2772)
	) name1556 (
		\TM0_pad ,
		\_2158__reg/NET0131 ,
		_w3063_,
		_w3064_,
		_w3065_
	);
	LUT4 #(
		.INIT('h2772)
	) name1557 (
		\TM0_pad ,
		\WX10857_reg/NET0131 ,
		_w2393_,
		_w2394_,
		_w3066_
	);
	LUT4 #(
		.INIT('h028a)
	) name1558 (
		RESET_pad,
		\TM1_pad ,
		_w3065_,
		_w3066_,
		_w3067_
	);
	LUT4 #(
		.INIT('h2772)
	) name1559 (
		\TM0_pad ,
		\_2157__reg/NET0131 ,
		_w1676_,
		_w1677_,
		_w3068_
	);
	LUT4 #(
		.INIT('h2772)
	) name1560 (
		\TM0_pad ,
		\WX10859_reg/NET0131 ,
		_w2449_,
		_w2450_,
		_w3069_
	);
	LUT4 #(
		.INIT('h028a)
	) name1561 (
		RESET_pad,
		\TM1_pad ,
		_w3068_,
		_w3069_,
		_w3070_
	);
	LUT3 #(
		.INIT('h96)
	) name1562 (
		\WX9776_reg/NET0131 ,
		\WX9840_reg/NET0131 ,
		\WX9904_reg/NET0131 ,
		_w3071_
	);
	LUT2 #(
		.INIT('h9)
	) name1563 (
		\TM1_pad ,
		\WX9712_reg/NET0131 ,
		_w3072_
	);
	LUT4 #(
		.INIT('h2772)
	) name1564 (
		\TM0_pad ,
		\_2292__reg/NET0131 ,
		_w3071_,
		_w3072_,
		_w3073_
	);
	LUT4 #(
		.INIT('h2772)
	) name1565 (
		\TM0_pad ,
		\WX10845_reg/NET0131 ,
		_w3042_,
		_w3043_,
		_w3074_
	);
	LUT4 #(
		.INIT('h028a)
	) name1566 (
		RESET_pad,
		\TM1_pad ,
		_w3073_,
		_w3074_,
		_w3075_
	);
	LUT3 #(
		.INIT('h96)
	) name1567 (
		\WX9778_reg/NET0131 ,
		\WX9842_reg/NET0131 ,
		\WX9906_reg/NET0131 ,
		_w3076_
	);
	LUT2 #(
		.INIT('h9)
	) name1568 (
		\TM1_pad ,
		\WX9714_reg/NET0131 ,
		_w3077_
	);
	LUT4 #(
		.INIT('h2772)
	) name1569 (
		\TM0_pad ,
		\_2291__reg/NET0131 ,
		_w3076_,
		_w3077_,
		_w3078_
	);
	LUT3 #(
		.INIT('h96)
	) name1570 (
		\WX8485_reg/NET0131 ,
		\WX8549_reg/NET0131 ,
		\WX8613_reg/NET0131 ,
		_w3079_
	);
	LUT2 #(
		.INIT('h9)
	) name1571 (
		\TM1_pad ,
		\WX8421_reg/NET0131 ,
		_w3080_
	);
	LUT4 #(
		.INIT('h2772)
	) name1572 (
		\TM0_pad ,
		\WX10847_reg/NET0131 ,
		_w3079_,
		_w3080_,
		_w3081_
	);
	LUT4 #(
		.INIT('h028a)
	) name1573 (
		RESET_pad,
		\TM1_pad ,
		_w3078_,
		_w3081_,
		_w3082_
	);
	LUT3 #(
		.INIT('h96)
	) name1574 (
		\WX9780_reg/NET0131 ,
		\WX9844_reg/NET0131 ,
		\WX9908_reg/NET0131 ,
		_w3083_
	);
	LUT2 #(
		.INIT('h9)
	) name1575 (
		\TM1_pad ,
		\WX9716_reg/NET0131 ,
		_w3084_
	);
	LUT4 #(
		.INIT('h2772)
	) name1576 (
		\TM0_pad ,
		\_2290__reg/NET0131 ,
		_w3083_,
		_w3084_,
		_w3085_
	);
	LUT3 #(
		.INIT('h96)
	) name1577 (
		\WX8487_reg/NET0131 ,
		\WX8551_reg/NET0131 ,
		\WX8615_reg/NET0131 ,
		_w3086_
	);
	LUT2 #(
		.INIT('h9)
	) name1578 (
		\TM1_pad ,
		\WX8423_reg/NET0131 ,
		_w3087_
	);
	LUT4 #(
		.INIT('h2772)
	) name1579 (
		\TM0_pad ,
		\WX10849_reg/NET0131 ,
		_w3086_,
		_w3087_,
		_w3088_
	);
	LUT4 #(
		.INIT('h028a)
	) name1580 (
		RESET_pad,
		\TM1_pad ,
		_w3085_,
		_w3088_,
		_w3089_
	);
	LUT4 #(
		.INIT('h2772)
	) name1581 (
		\TM0_pad ,
		\_2289__reg/NET0131 ,
		_w1669_,
		_w1670_,
		_w3090_
	);
	LUT3 #(
		.INIT('h96)
	) name1582 (
		\WX8489_reg/NET0131 ,
		\WX8553_reg/NET0131 ,
		\WX8617_reg/NET0131 ,
		_w3091_
	);
	LUT2 #(
		.INIT('h9)
	) name1583 (
		\TM1_pad ,
		\WX8425_reg/NET0131 ,
		_w3092_
	);
	LUT4 #(
		.INIT('h2772)
	) name1584 (
		\TM0_pad ,
		\WX10851_reg/NET0131 ,
		_w3091_,
		_w3092_,
		_w3093_
	);
	LUT4 #(
		.INIT('h028a)
	) name1585 (
		RESET_pad,
		\TM1_pad ,
		_w3090_,
		_w3093_,
		_w3094_
	);
	LUT4 #(
		.INIT('h2772)
	) name1586 (
		\TM0_pad ,
		\_2325__reg/NET0131 ,
		_w2027_,
		_w2028_,
		_w3095_
	);
	LUT4 #(
		.INIT('h2772)
	) name1587 (
		\TM0_pad ,
		\WX10843_reg/NET0131 ,
		_w3020_,
		_w3021_,
		_w3096_
	);
	LUT4 #(
		.INIT('h028a)
	) name1588 (
		RESET_pad,
		\TM1_pad ,
		_w3095_,
		_w3096_,
		_w3097_
	);
	LUT4 #(
		.INIT('h2772)
	) name1589 (
		\TM0_pad ,
		\_2324__reg/NET0131 ,
		_w2081_,
		_w2082_,
		_w3098_
	);
	LUT4 #(
		.INIT('h2772)
	) name1590 (
		\TM0_pad ,
		\WX10845_reg/NET0131 ,
		_w3071_,
		_w3072_,
		_w3099_
	);
	LUT4 #(
		.INIT('h028a)
	) name1591 (
		RESET_pad,
		\TM1_pad ,
		_w3098_,
		_w3099_,
		_w3100_
	);
	LUT4 #(
		.INIT('h2772)
	) name1592 (
		\TM0_pad ,
		\_2323__reg/NET0131 ,
		_w2138_,
		_w2139_,
		_w3101_
	);
	LUT4 #(
		.INIT('h2772)
	) name1593 (
		\TM0_pad ,
		\WX10847_reg/NET0131 ,
		_w3076_,
		_w3077_,
		_w3102_
	);
	LUT4 #(
		.INIT('h028a)
	) name1594 (
		RESET_pad,
		\TM1_pad ,
		_w3101_,
		_w3102_,
		_w3103_
	);
	LUT4 #(
		.INIT('h2772)
	) name1595 (
		\TM0_pad ,
		\_2322__reg/NET0131 ,
		_w2195_,
		_w2196_,
		_w3104_
	);
	LUT4 #(
		.INIT('h2772)
	) name1596 (
		\TM0_pad ,
		\WX10849_reg/NET0131 ,
		_w3083_,
		_w3084_,
		_w3105_
	);
	LUT4 #(
		.INIT('h028a)
	) name1597 (
		RESET_pad,
		\TM1_pad ,
		_w3104_,
		_w3105_,
		_w3106_
	);
	LUT3 #(
		.INIT('h96)
	) name1598 (
		\WX5903_reg/NET0131 ,
		\WX5967_reg/NET0131 ,
		\WX6031_reg/NET0131 ,
		_w3107_
	);
	LUT2 #(
		.INIT('h9)
	) name1599 (
		\TM1_pad ,
		\WX5839_reg/NET0131 ,
		_w3108_
	);
	LUT4 #(
		.INIT('h2772)
	) name1600 (
		\TM0_pad ,
		\_2193__reg/NET0131 ,
		_w3107_,
		_w3108_,
		_w3109_
	);
	LUT4 #(
		.INIT('h2772)
	) name1601 (
		\TM0_pad ,
		\WX10851_reg/NET0131 ,
		_w3015_,
		_w3016_,
		_w3110_
	);
	LUT4 #(
		.INIT('h028a)
	) name1602 (
		RESET_pad,
		\TM1_pad ,
		_w3109_,
		_w3110_,
		_w3111_
	);
	LUT3 #(
		.INIT('h96)
	) name1603 (
		\WX5905_reg/NET0131 ,
		\WX5969_reg/NET0131 ,
		\WX6033_reg/NET0131 ,
		_w3112_
	);
	LUT2 #(
		.INIT('h9)
	) name1604 (
		\TM1_pad ,
		\WX5841_reg/NET0131 ,
		_w3113_
	);
	LUT4 #(
		.INIT('h2772)
	) name1605 (
		\TM0_pad ,
		\_2192__reg/NET0131 ,
		_w3112_,
		_w3113_,
		_w3114_
	);
	LUT4 #(
		.INIT('h7227)
	) name1606 (
		\TM0_pad ,
		\WX10853_reg/NET0131 ,
		_w3053_,
		_w3054_,
		_w3115_
	);
	LUT4 #(
		.INIT('h028a)
	) name1607 (
		RESET_pad,
		\TM1_pad ,
		_w3114_,
		_w3115_,
		_w3116_
	);
	LUT3 #(
		.INIT('h96)
	) name1608 (
		\WX5907_reg/NET0131 ,
		\WX5971_reg/NET0131 ,
		\WX6035_reg/NET0131 ,
		_w3117_
	);
	LUT2 #(
		.INIT('h9)
	) name1609 (
		\TM1_pad ,
		\WX5843_reg/NET0131 ,
		_w3118_
	);
	LUT4 #(
		.INIT('h2772)
	) name1610 (
		\TM0_pad ,
		\_2191__reg/NET0131 ,
		_w3117_,
		_w3118_,
		_w3119_
	);
	LUT4 #(
		.INIT('h2772)
	) name1611 (
		\TM0_pad ,
		\WX10855_reg/NET0131 ,
		_w3058_,
		_w3059_,
		_w3120_
	);
	LUT4 #(
		.INIT('h028a)
	) name1612 (
		RESET_pad,
		\TM1_pad ,
		_w3119_,
		_w3120_,
		_w3121_
	);
	LUT4 #(
		.INIT('h2772)
	) name1613 (
		\TM0_pad ,
		\_2190__reg/NET0131 ,
		_w1683_,
		_w1684_,
		_w3122_
	);
	LUT4 #(
		.INIT('h2772)
	) name1614 (
		\TM0_pad ,
		\WX10857_reg/NET0131 ,
		_w3063_,
		_w3064_,
		_w3123_
	);
	LUT4 #(
		.INIT('h028a)
	) name1615 (
		RESET_pad,
		\TM1_pad ,
		_w3122_,
		_w3123_,
		_w3124_
	);
	LUT3 #(
		.INIT('h96)
	) name1616 (
		\WX7194_reg/NET0131 ,
		\WX7258_reg/NET0131 ,
		\WX7322_reg/NET0131 ,
		_w3125_
	);
	LUT2 #(
		.INIT('h9)
	) name1617 (
		\TM1_pad ,
		\WX7130_reg/NET0131 ,
		_w3126_
	);
	LUT4 #(
		.INIT('h2772)
	) name1618 (
		\TM0_pad ,
		\_2226__reg/NET0131 ,
		_w3125_,
		_w3126_,
		_w3127_
	);
	LUT4 #(
		.INIT('h2772)
	) name1619 (
		\TM0_pad ,
		\WX10849_reg/NET0131 ,
		_w3028_,
		_w3029_,
		_w3128_
	);
	LUT4 #(
		.INIT('h028a)
	) name1620 (
		RESET_pad,
		\TM1_pad ,
		_w3127_,
		_w3128_,
		_w3129_
	);
	LUT3 #(
		.INIT('h96)
	) name1621 (
		\WX7196_reg/NET0131 ,
		\WX7260_reg/NET0131 ,
		\WX7324_reg/NET0131 ,
		_w3130_
	);
	LUT2 #(
		.INIT('h9)
	) name1622 (
		\TM1_pad ,
		\WX7132_reg/NET0131 ,
		_w3131_
	);
	LUT4 #(
		.INIT('h2772)
	) name1623 (
		\TM0_pad ,
		\_2225__reg/NET0131 ,
		_w3130_,
		_w3131_,
		_w3132_
	);
	LUT4 #(
		.INIT('h2772)
	) name1624 (
		\TM0_pad ,
		\WX10851_reg/NET0131 ,
		_w3107_,
		_w3108_,
		_w3133_
	);
	LUT4 #(
		.INIT('h028a)
	) name1625 (
		RESET_pad,
		\TM1_pad ,
		_w3132_,
		_w3133_,
		_w3134_
	);
	LUT3 #(
		.INIT('h96)
	) name1626 (
		\WX7198_reg/NET0131 ,
		\WX7262_reg/NET0131 ,
		\WX7326_reg/NET0131 ,
		_w3135_
	);
	LUT2 #(
		.INIT('h9)
	) name1627 (
		\TM1_pad ,
		\WX7134_reg/NET0131 ,
		_w3136_
	);
	LUT4 #(
		.INIT('h2772)
	) name1628 (
		\TM0_pad ,
		\_2224__reg/NET0131 ,
		_w3135_,
		_w3136_,
		_w3137_
	);
	LUT4 #(
		.INIT('h2772)
	) name1629 (
		\TM0_pad ,
		\WX10853_reg/NET0131 ,
		_w3112_,
		_w3113_,
		_w3138_
	);
	LUT4 #(
		.INIT('h028a)
	) name1630 (
		RESET_pad,
		\TM1_pad ,
		_w3137_,
		_w3138_,
		_w3139_
	);
	LUT4 #(
		.INIT('h2772)
	) name1631 (
		\TM0_pad ,
		\_2223__reg/NET0131 ,
		_w1690_,
		_w1691_,
		_w3140_
	);
	LUT4 #(
		.INIT('h2772)
	) name1632 (
		\TM0_pad ,
		\WX10855_reg/NET0131 ,
		_w3117_,
		_w3118_,
		_w3141_
	);
	LUT4 #(
		.INIT('h028a)
	) name1633 (
		RESET_pad,
		\TM1_pad ,
		_w3140_,
		_w3141_,
		_w3142_
	);
	LUT4 #(
		.INIT('h8cc8)
	) name1634 (
		\TM0_pad ,
		_w2366_,
		_w2993_,
		_w2994_,
		_w3143_
	);
	LUT4 #(
		.INIT('h0a02)
	) name1635 (
		RESET_pad,
		\TM0_pad ,
		\TM1_pad ,
		\_2111__reg/NET0131 ,
		_w3144_
	);
	LUT4 #(
		.INIT('hbe00)
	) name1636 (
		\TM0_pad ,
		_w2367_,
		_w2368_,
		_w3144_,
		_w3145_
	);
	LUT2 #(
		.INIT('he)
	) name1637 (
		_w3143_,
		_w3145_,
		_w3146_
	);
	LUT2 #(
		.INIT('h9)
	) name1638 (
		\WX2126_reg/NET0131 ,
		\WX2190_reg/NET0131 ,
		_w3147_
	);
	LUT2 #(
		.INIT('h9)
	) name1639 (
		\WX1998_reg/NET0131 ,
		\WX2062_reg/NET0131 ,
		_w3148_
	);
	LUT4 #(
		.INIT('h8cc8)
	) name1640 (
		\TM0_pad ,
		_w2422_,
		_w3147_,
		_w3148_,
		_w3149_
	);
	LUT4 #(
		.INIT('h0a02)
	) name1641 (
		RESET_pad,
		\TM0_pad ,
		\TM1_pad ,
		\_2110__reg/NET0131 ,
		_w3150_
	);
	LUT4 #(
		.INIT('hbe00)
	) name1642 (
		\TM0_pad ,
		_w2423_,
		_w2424_,
		_w3150_,
		_w3151_
	);
	LUT2 #(
		.INIT('he)
	) name1643 (
		_w3149_,
		_w3151_,
		_w3152_
	);
	LUT4 #(
		.INIT('h8cc8)
	) name1644 (
		\TM0_pad ,
		_w2472_,
		_w2999_,
		_w3000_,
		_w3153_
	);
	LUT4 #(
		.INIT('h0a02)
	) name1645 (
		RESET_pad,
		\TM0_pad ,
		\TM1_pad ,
		\_2109__reg/NET0131 ,
		_w3154_
	);
	LUT4 #(
		.INIT('hbe00)
	) name1646 (
		\TM0_pad ,
		_w2473_,
		_w2474_,
		_w3154_,
		_w3155_
	);
	LUT2 #(
		.INIT('he)
	) name1647 (
		_w3153_,
		_w3155_,
		_w3156_
	);
	LUT4 #(
		.INIT('h2772)
	) name1648 (
		\TM0_pad ,
		\_2259__reg/NET0131 ,
		_w3079_,
		_w3080_,
		_w3157_
	);
	LUT4 #(
		.INIT('h2772)
	) name1649 (
		\TM0_pad ,
		\WX10847_reg/NET0131 ,
		_w3033_,
		_w3034_,
		_w3158_
	);
	LUT4 #(
		.INIT('h028a)
	) name1650 (
		RESET_pad,
		\TM1_pad ,
		_w3157_,
		_w3158_,
		_w3159_
	);
	LUT4 #(
		.INIT('h2772)
	) name1651 (
		\TM0_pad ,
		\_2258__reg/NET0131 ,
		_w3086_,
		_w3087_,
		_w3160_
	);
	LUT4 #(
		.INIT('h2772)
	) name1652 (
		\TM0_pad ,
		\WX10849_reg/NET0131 ,
		_w3125_,
		_w3126_,
		_w3161_
	);
	LUT4 #(
		.INIT('h028a)
	) name1653 (
		RESET_pad,
		\TM1_pad ,
		_w3160_,
		_w3161_,
		_w3162_
	);
	LUT4 #(
		.INIT('h2772)
	) name1654 (
		\TM0_pad ,
		\_2257__reg/NET0131 ,
		_w3091_,
		_w3092_,
		_w3163_
	);
	LUT4 #(
		.INIT('h2772)
	) name1655 (
		\TM0_pad ,
		\WX10851_reg/NET0131 ,
		_w3130_,
		_w3131_,
		_w3164_
	);
	LUT4 #(
		.INIT('h028a)
	) name1656 (
		RESET_pad,
		\TM1_pad ,
		_w3163_,
		_w3164_,
		_w3165_
	);
	LUT4 #(
		.INIT('h2772)
	) name1657 (
		\TM0_pad ,
		\_2256__reg/NET0131 ,
		_w1662_,
		_w1663_,
		_w3166_
	);
	LUT4 #(
		.INIT('h2772)
	) name1658 (
		\TM0_pad ,
		\WX10853_reg/NET0131 ,
		_w3135_,
		_w3136_,
		_w3167_
	);
	LUT4 #(
		.INIT('h028a)
	) name1659 (
		RESET_pad,
		\TM1_pad ,
		_w3166_,
		_w3167_,
		_w3168_
	);
	LUT4 #(
		.INIT('h8cc8)
	) name1660 (
		\TM0_pad ,
		_w2366_,
		_w2628_,
		_w2629_,
		_w3169_
	);
	LUT2 #(
		.INIT('h2)
	) name1661 (
		\TM0_pad ,
		\_2335__reg/NET0131 ,
		_w3170_
	);
	LUT4 #(
		.INIT('h00c8)
	) name1662 (
		\DATA_0_2_pad ,
		RESET_pad,
		\TM0_pad ,
		\TM1_pad ,
		_w3171_
	);
	LUT2 #(
		.INIT('h4)
	) name1663 (
		_w3170_,
		_w3171_,
		_w3172_
	);
	LUT2 #(
		.INIT('he)
	) name1664 (
		_w3169_,
		_w3172_,
		_w3173_
	);
	LUT4 #(
		.INIT('h8cc8)
	) name1665 (
		\TM0_pad ,
		_w2422_,
		_w2671_,
		_w2672_,
		_w3174_
	);
	LUT2 #(
		.INIT('h2)
	) name1666 (
		\TM0_pad ,
		\_2334__reg/NET0131 ,
		_w3175_
	);
	LUT4 #(
		.INIT('h00c8)
	) name1667 (
		\DATA_0_1_pad ,
		RESET_pad,
		\TM0_pad ,
		\TM1_pad ,
		_w3176_
	);
	LUT2 #(
		.INIT('h4)
	) name1668 (
		_w3175_,
		_w3176_,
		_w3177_
	);
	LUT2 #(
		.INIT('he)
	) name1669 (
		_w3174_,
		_w3177_,
		_w3178_
	);
	LUT4 #(
		.INIT('h8cc8)
	) name1670 (
		\TM0_pad ,
		_w2472_,
		_w2714_,
		_w2715_,
		_w3179_
	);
	LUT2 #(
		.INIT('h2)
	) name1671 (
		\TM0_pad ,
		\_2333__reg/NET0131 ,
		_w3180_
	);
	LUT4 #(
		.INIT('h00c8)
	) name1672 (
		\DATA_0_0_pad ,
		RESET_pad,
		\TM0_pad ,
		\TM1_pad ,
		_w3181_
	);
	LUT2 #(
		.INIT('h4)
	) name1673 (
		_w3180_,
		_w3181_,
		_w3182_
	);
	LUT2 #(
		.INIT('he)
	) name1674 (
		_w3179_,
		_w3182_,
		_w3183_
	);
	LUT2 #(
		.INIT('h8)
	) name1675 (
		RESET_pad,
		\WX10885_reg/NET0131 ,
		_w3184_
	);
	LUT3 #(
		.INIT('h82)
	) name1676 (
		RESET_pad,
		\WX837_reg/NET0131 ,
		\_2107__reg/NET0131 ,
		_w3185_
	);
	LUT3 #(
		.INIT('h82)
	) name1677 (
		RESET_pad,
		\WX2130_reg/NET0131 ,
		\_2139__reg/NET0131 ,
		_w3186_
	);
	LUT3 #(
		.INIT('h82)
	) name1678 (
		RESET_pad,
		\WX11181_reg/NET0131 ,
		\_2363__reg/NET0131 ,
		_w3187_
	);
	LUT2 #(
		.INIT('h8)
	) name1679 (
		RESET_pad,
		\WX10887_reg/NET0131 ,
		_w3188_
	);
	LUT4 #(
		.INIT('h2882)
	) name1680 (
		RESET_pad,
		\WX891_reg/NET0131 ,
		\_2080__reg/NET0131 ,
		\_2108__reg/NET0131 ,
		_w3189_
	);
	LUT4 #(
		.INIT('h2882)
	) name1681 (
		RESET_pad,
		\WX877_reg/NET0131 ,
		\_2087__reg/NET0131 ,
		\_2108__reg/NET0131 ,
		_w3190_
	);
	LUT4 #(
		.INIT('h2882)
	) name1682 (
		RESET_pad,
		\WX867_reg/NET0131 ,
		\_2092__reg/NET0131 ,
		\_2108__reg/NET0131 ,
		_w3191_
	);
	LUT4 #(
		.INIT('h2882)
	) name1683 (
		RESET_pad,
		\WX2184_reg/NET0131 ,
		\_2112__reg/NET0131 ,
		\_2140__reg/NET0131 ,
		_w3192_
	);
	LUT4 #(
		.INIT('h2882)
	) name1684 (
		RESET_pad,
		\WX2170_reg/NET0131 ,
		\_2119__reg/NET0131 ,
		\_2140__reg/NET0131 ,
		_w3193_
	);
	LUT4 #(
		.INIT('h2882)
	) name1685 (
		RESET_pad,
		\WX2160_reg/NET0131 ,
		\_2124__reg/NET0131 ,
		\_2140__reg/NET0131 ,
		_w3194_
	);
	LUT4 #(
		.INIT('h2882)
	) name1686 (
		RESET_pad,
		\WX3477_reg/NET0131 ,
		\_2144__reg/NET0131 ,
		\_2172__reg/NET0131 ,
		_w3195_
	);
	LUT4 #(
		.INIT('h2882)
	) name1687 (
		RESET_pad,
		\WX3463_reg/NET0131 ,
		\_2151__reg/NET0131 ,
		\_2172__reg/NET0131 ,
		_w3196_
	);
	LUT4 #(
		.INIT('h2882)
	) name1688 (
		RESET_pad,
		\WX3453_reg/NET0131 ,
		\_2156__reg/NET0131 ,
		\_2172__reg/NET0131 ,
		_w3197_
	);
	LUT4 #(
		.INIT('h2882)
	) name1689 (
		RESET_pad,
		\WX4770_reg/NET0131 ,
		\_2176__reg/NET0131 ,
		\_2204__reg/NET0131 ,
		_w3198_
	);
	LUT4 #(
		.INIT('h2882)
	) name1690 (
		RESET_pad,
		\WX4756_reg/NET0131 ,
		\_2183__reg/NET0131 ,
		\_2204__reg/NET0131 ,
		_w3199_
	);
	LUT4 #(
		.INIT('h2882)
	) name1691 (
		RESET_pad,
		\WX4746_reg/NET0131 ,
		\_2188__reg/NET0131 ,
		\_2204__reg/NET0131 ,
		_w3200_
	);
	LUT4 #(
		.INIT('h2882)
	) name1692 (
		RESET_pad,
		\WX6063_reg/NET0131 ,
		\_2208__reg/NET0131 ,
		\_2236__reg/NET0131 ,
		_w3201_
	);
	LUT4 #(
		.INIT('h2882)
	) name1693 (
		RESET_pad,
		\WX6049_reg/NET0131 ,
		\_2215__reg/NET0131 ,
		\_2236__reg/NET0131 ,
		_w3202_
	);
	LUT4 #(
		.INIT('h2882)
	) name1694 (
		RESET_pad,
		\WX6039_reg/NET0131 ,
		\_2220__reg/NET0131 ,
		\_2236__reg/NET0131 ,
		_w3203_
	);
	LUT4 #(
		.INIT('h2882)
	) name1695 (
		RESET_pad,
		\WX7356_reg/NET0131 ,
		\_2240__reg/NET0131 ,
		\_2268__reg/NET0131 ,
		_w3204_
	);
	LUT4 #(
		.INIT('h2882)
	) name1696 (
		RESET_pad,
		\WX7342_reg/NET0131 ,
		\_2247__reg/NET0131 ,
		\_2268__reg/NET0131 ,
		_w3205_
	);
	LUT4 #(
		.INIT('h2882)
	) name1697 (
		RESET_pad,
		\WX7332_reg/NET0131 ,
		\_2252__reg/NET0131 ,
		\_2268__reg/NET0131 ,
		_w3206_
	);
	LUT4 #(
		.INIT('h2882)
	) name1698 (
		RESET_pad,
		\WX8649_reg/NET0131 ,
		\_2272__reg/NET0131 ,
		\_2300__reg/NET0131 ,
		_w3207_
	);
	LUT4 #(
		.INIT('h2882)
	) name1699 (
		RESET_pad,
		\WX8635_reg/NET0131 ,
		\_2279__reg/NET0131 ,
		\_2300__reg/NET0131 ,
		_w3208_
	);
	LUT4 #(
		.INIT('h2882)
	) name1700 (
		RESET_pad,
		\WX8625_reg/NET0131 ,
		\_2284__reg/NET0131 ,
		\_2300__reg/NET0131 ,
		_w3209_
	);
	LUT4 #(
		.INIT('h2882)
	) name1701 (
		RESET_pad,
		\WX9942_reg/NET0131 ,
		\_2304__reg/NET0131 ,
		\_2332__reg/NET0131 ,
		_w3210_
	);
	LUT4 #(
		.INIT('h2882)
	) name1702 (
		RESET_pad,
		\WX9928_reg/NET0131 ,
		\_2311__reg/NET0131 ,
		\_2332__reg/NET0131 ,
		_w3211_
	);
	LUT4 #(
		.INIT('h2882)
	) name1703 (
		RESET_pad,
		\WX9918_reg/NET0131 ,
		\_2316__reg/NET0131 ,
		\_2332__reg/NET0131 ,
		_w3212_
	);
	LUT4 #(
		.INIT('h2882)
	) name1704 (
		RESET_pad,
		\WX11235_reg/NET0131 ,
		\_2336__reg/NET0131 ,
		\_2364__reg/NET0131 ,
		_w3213_
	);
	LUT4 #(
		.INIT('h2882)
	) name1705 (
		RESET_pad,
		\WX11221_reg/NET0131 ,
		\_2343__reg/NET0131 ,
		\_2364__reg/NET0131 ,
		_w3214_
	);
	LUT4 #(
		.INIT('h2882)
	) name1706 (
		RESET_pad,
		\WX11211_reg/NET0131 ,
		\_2348__reg/NET0131 ,
		\_2364__reg/NET0131 ,
		_w3215_
	);
	LUT2 #(
		.INIT('h8)
	) name1707 (
		RESET_pad,
		\WX11117_reg/NET0131 ,
		_w3216_
	);
	LUT2 #(
		.INIT('h8)
	) name1708 (
		RESET_pad,
		\WX773_reg/NET0131 ,
		_w3217_
	);
	LUT2 #(
		.INIT('h8)
	) name1709 (
		RESET_pad,
		\WX10889_reg/NET0131 ,
		_w3218_
	);
	LUT2 #(
		.INIT('h8)
	) name1710 (
		RESET_pad,
		\WX2066_reg/NET0131 ,
		_w3219_
	);
	LUT3 #(
		.INIT('h82)
	) name1711 (
		RESET_pad,
		\WX3475_reg/NET0131 ,
		\_2145__reg/NET0131 ,
		_w3220_
	);
	LUT3 #(
		.INIT('h82)
	) name1712 (
		RESET_pad,
		\WX3427_reg/NET0131 ,
		\_2169__reg/NET0131 ,
		_w3221_
	);
	LUT3 #(
		.INIT('h82)
	) name1713 (
		RESET_pad,
		\WX2132_reg/NET0131 ,
		\_2138__reg/NET0131 ,
		_w3222_
	);
	LUT3 #(
		.INIT('h82)
	) name1714 (
		RESET_pad,
		\WX11215_reg/NET0131 ,
		\_2346__reg/NET0131 ,
		_w3223_
	);
	LUT3 #(
		.INIT('h82)
	) name1715 (
		RESET_pad,
		\WX8599_reg/NET0131 ,
		\_2297__reg/NET0131 ,
		_w3224_
	);
	LUT3 #(
		.INIT('h82)
	) name1716 (
		RESET_pad,
		\WX6043_reg/NET0131 ,
		\_2218__reg/NET0131 ,
		_w3225_
	);
	LUT3 #(
		.INIT('h82)
	) name1717 (
		RESET_pad,
		\WX3461_reg/NET0131 ,
		\_2152__reg/NET0131 ,
		_w3226_
	);
	LUT3 #(
		.INIT('h82)
	) name1718 (
		RESET_pad,
		\WX857_reg/NET0131 ,
		\_2097__reg/NET0131 ,
		_w3227_
	);
	LUT3 #(
		.INIT('h82)
	) name1719 (
		RESET_pad,
		\WX9934_reg/NET0131 ,
		\_2308__reg/NET0131 ,
		_w3228_
	);
	LUT3 #(
		.INIT('h82)
	) name1720 (
		RESET_pad,
		\WX7312_reg/NET0131 ,
		\_2262__reg/NET0131 ,
		_w3229_
	);
	LUT3 #(
		.INIT('h82)
	) name1721 (
		RESET_pad,
		\WX7338_reg/NET0131 ,
		\_2249__reg/NET0131 ,
		_w3230_
	);
	LUT3 #(
		.INIT('h82)
	) name1722 (
		RESET_pad,
		\WX8605_reg/NET0131 ,
		\_2294__reg/NET0131 ,
		_w3231_
	);
	LUT3 #(
		.INIT('h82)
	) name1723 (
		RESET_pad,
		\WX8601_reg/NET0131 ,
		\_2296__reg/NET0131 ,
		_w3232_
	);
	LUT3 #(
		.INIT('h82)
	) name1724 (
		RESET_pad,
		\WX8603_reg/NET0131 ,
		\_2295__reg/NET0131 ,
		_w3233_
	);
	LUT3 #(
		.INIT('h82)
	) name1725 (
		RESET_pad,
		\WX6037_reg/NET0131 ,
		\_2221__reg/NET0131 ,
		_w3234_
	);
	LUT3 #(
		.INIT('h82)
	) name1726 (
		RESET_pad,
		\WX8619_reg/NET0131 ,
		\_2287__reg/NET0131 ,
		_w3235_
	);
	LUT3 #(
		.INIT('h82)
	) name1727 (
		RESET_pad,
		\WX7362_reg/NET0131 ,
		\_2237__reg/NET0131 ,
		_w3236_
	);
	LUT3 #(
		.INIT('h82)
	) name1728 (
		RESET_pad,
		\WX3425_reg/NET0131 ,
		\_2170__reg/NET0131 ,
		_w3237_
	);
	LUT3 #(
		.INIT('h82)
	) name1729 (
		RESET_pad,
		\WX4728_reg/NET0131 ,
		\_2197__reg/NET0131 ,
		_w3238_
	);
	LUT3 #(
		.INIT('h82)
	) name1730 (
		RESET_pad,
		\WX3485_reg/NET0131 ,
		\_2172__reg/NET0131 ,
		_w3239_
	);
	LUT3 #(
		.INIT('h82)
	) name1731 (
		RESET_pad,
		\WX7328_reg/NET0131 ,
		\_2254__reg/NET0131 ,
		_w3240_
	);
	LUT3 #(
		.INIT('h82)
	) name1732 (
		RESET_pad,
		\WX9930_reg/NET0131 ,
		\_2310__reg/NET0131 ,
		_w3241_
	);
	LUT3 #(
		.INIT('h82)
	) name1733 (
		RESET_pad,
		\WX2148_reg/NET0131 ,
		\_2130__reg/NET0131 ,
		_w3242_
	);
	LUT3 #(
		.INIT('h82)
	) name1734 (
		RESET_pad,
		\WX7340_reg/NET0131 ,
		\_2248__reg/NET0131 ,
		_w3243_
	);
	LUT3 #(
		.INIT('h82)
	) name1735 (
		RESET_pad,
		\WX6061_reg/NET0131 ,
		\_2209__reg/NET0131 ,
		_w3244_
	);
	LUT3 #(
		.INIT('h82)
	) name1736 (
		RESET_pad,
		\WX8657_reg/NET0131 ,
		\_2300__reg/NET0131 ,
		_w3245_
	);
	LUT3 #(
		.INIT('h82)
	) name1737 (
		RESET_pad,
		\WX2172_reg/NET0131 ,
		\_2118__reg/NET0131 ,
		_w3246_
	);
	LUT3 #(
		.INIT('h82)
	) name1738 (
		RESET_pad,
		\WX8607_reg/NET0131 ,
		\_2293__reg/NET0131 ,
		_w3247_
	);
	LUT3 #(
		.INIT('h82)
	) name1739 (
		RESET_pad,
		\WX899_reg/NET0131 ,
		\_2108__reg/NET0131 ,
		_w3248_
	);
	LUT3 #(
		.INIT('h82)
	) name1740 (
		RESET_pad,
		\WX897_reg/NET0131 ,
		\_2077__reg/NET0131 ,
		_w3249_
	);
	LUT3 #(
		.INIT('h82)
	) name1741 (
		RESET_pad,
		\WX895_reg/NET0131 ,
		\_2078__reg/NET0131 ,
		_w3250_
	);
	LUT3 #(
		.INIT('h82)
	) name1742 (
		RESET_pad,
		\WX893_reg/NET0131 ,
		\_2079__reg/NET0131 ,
		_w3251_
	);
	LUT3 #(
		.INIT('h82)
	) name1743 (
		RESET_pad,
		\WX889_reg/NET0131 ,
		\_2081__reg/NET0131 ,
		_w3252_
	);
	LUT3 #(
		.INIT('h82)
	) name1744 (
		RESET_pad,
		\WX887_reg/NET0131 ,
		\_2082__reg/NET0131 ,
		_w3253_
	);
	LUT3 #(
		.INIT('h82)
	) name1745 (
		RESET_pad,
		\WX883_reg/NET0131 ,
		\_2084__reg/NET0131 ,
		_w3254_
	);
	LUT3 #(
		.INIT('h82)
	) name1746 (
		RESET_pad,
		\WX881_reg/NET0131 ,
		\_2085__reg/NET0131 ,
		_w3255_
	);
	LUT3 #(
		.INIT('h82)
	) name1747 (
		RESET_pad,
		\WX875_reg/NET0131 ,
		\_2088__reg/NET0131 ,
		_w3256_
	);
	LUT3 #(
		.INIT('h82)
	) name1748 (
		RESET_pad,
		\WX873_reg/NET0131 ,
		\_2089__reg/NET0131 ,
		_w3257_
	);
	LUT3 #(
		.INIT('h82)
	) name1749 (
		RESET_pad,
		\WX869_reg/NET0131 ,
		\_2091__reg/NET0131 ,
		_w3258_
	);
	LUT3 #(
		.INIT('h82)
	) name1750 (
		RESET_pad,
		\WX865_reg/NET0131 ,
		\_2093__reg/NET0131 ,
		_w3259_
	);
	LUT3 #(
		.INIT('h82)
	) name1751 (
		RESET_pad,
		\WX863_reg/NET0131 ,
		\_2094__reg/NET0131 ,
		_w3260_
	);
	LUT3 #(
		.INIT('h82)
	) name1752 (
		RESET_pad,
		\WX855_reg/NET0131 ,
		\_2098__reg/NET0131 ,
		_w3261_
	);
	LUT3 #(
		.INIT('h82)
	) name1753 (
		RESET_pad,
		\WX851_reg/NET0131 ,
		\_2100__reg/NET0131 ,
		_w3262_
	);
	LUT3 #(
		.INIT('h82)
	) name1754 (
		RESET_pad,
		\WX845_reg/NET0131 ,
		\_2103__reg/NET0131 ,
		_w3263_
	);
	LUT3 #(
		.INIT('h82)
	) name1755 (
		RESET_pad,
		\WX843_reg/NET0131 ,
		\_2104__reg/NET0131 ,
		_w3264_
	);
	LUT3 #(
		.INIT('h82)
	) name1756 (
		RESET_pad,
		\WX841_reg/NET0131 ,
		\_2105__reg/NET0131 ,
		_w3265_
	);
	LUT3 #(
		.INIT('h82)
	) name1757 (
		RESET_pad,
		\WX839_reg/NET0131 ,
		\_2106__reg/NET0131 ,
		_w3266_
	);
	LUT3 #(
		.INIT('h82)
	) name1758 (
		RESET_pad,
		\WX2192_reg/NET0131 ,
		\_2140__reg/NET0131 ,
		_w3267_
	);
	LUT3 #(
		.INIT('h82)
	) name1759 (
		RESET_pad,
		\WX2190_reg/NET0131 ,
		\_2109__reg/NET0131 ,
		_w3268_
	);
	LUT3 #(
		.INIT('h82)
	) name1760 (
		RESET_pad,
		\WX2188_reg/NET0131 ,
		\_2110__reg/NET0131 ,
		_w3269_
	);
	LUT3 #(
		.INIT('h82)
	) name1761 (
		RESET_pad,
		\WX2186_reg/NET0131 ,
		\_2111__reg/NET0131 ,
		_w3270_
	);
	LUT3 #(
		.INIT('h82)
	) name1762 (
		RESET_pad,
		\WX2182_reg/NET0131 ,
		\_2113__reg/NET0131 ,
		_w3271_
	);
	LUT3 #(
		.INIT('h82)
	) name1763 (
		RESET_pad,
		\WX2180_reg/NET0131 ,
		\_2114__reg/NET0131 ,
		_w3272_
	);
	LUT3 #(
		.INIT('h82)
	) name1764 (
		RESET_pad,
		\WX2174_reg/NET0131 ,
		\_2117__reg/NET0131 ,
		_w3273_
	);
	LUT3 #(
		.INIT('h82)
	) name1765 (
		RESET_pad,
		\WX2168_reg/NET0131 ,
		\_2120__reg/NET0131 ,
		_w3274_
	);
	LUT3 #(
		.INIT('h82)
	) name1766 (
		RESET_pad,
		\WX2166_reg/NET0131 ,
		\_2121__reg/NET0131 ,
		_w3275_
	);
	LUT3 #(
		.INIT('h82)
	) name1767 (
		RESET_pad,
		\WX2164_reg/NET0131 ,
		\_2122__reg/NET0131 ,
		_w3276_
	);
	LUT3 #(
		.INIT('h82)
	) name1768 (
		RESET_pad,
		\WX2162_reg/NET0131 ,
		\_2123__reg/NET0131 ,
		_w3277_
	);
	LUT3 #(
		.INIT('h82)
	) name1769 (
		RESET_pad,
		\WX2158_reg/NET0131 ,
		\_2125__reg/NET0131 ,
		_w3278_
	);
	LUT3 #(
		.INIT('h82)
	) name1770 (
		RESET_pad,
		\WX2156_reg/NET0131 ,
		\_2126__reg/NET0131 ,
		_w3279_
	);
	LUT3 #(
		.INIT('h82)
	) name1771 (
		RESET_pad,
		\WX2154_reg/NET0131 ,
		\_2127__reg/NET0131 ,
		_w3280_
	);
	LUT3 #(
		.INIT('h82)
	) name1772 (
		RESET_pad,
		\WX2146_reg/NET0131 ,
		\_2131__reg/NET0131 ,
		_w3281_
	);
	LUT3 #(
		.INIT('h82)
	) name1773 (
		RESET_pad,
		\WX2144_reg/NET0131 ,
		\_2132__reg/NET0131 ,
		_w3282_
	);
	LUT3 #(
		.INIT('h82)
	) name1774 (
		RESET_pad,
		\WX2142_reg/NET0131 ,
		\_2133__reg/NET0131 ,
		_w3283_
	);
	LUT3 #(
		.INIT('h82)
	) name1775 (
		RESET_pad,
		\WX2138_reg/NET0131 ,
		\_2135__reg/NET0131 ,
		_w3284_
	);
	LUT3 #(
		.INIT('h82)
	) name1776 (
		RESET_pad,
		\WX2134_reg/NET0131 ,
		\_2137__reg/NET0131 ,
		_w3285_
	);
	LUT3 #(
		.INIT('h82)
	) name1777 (
		RESET_pad,
		\WX7348_reg/NET0131 ,
		\_2244__reg/NET0131 ,
		_w3286_
	);
	LUT3 #(
		.INIT('h82)
	) name1778 (
		RESET_pad,
		\WX3483_reg/NET0131 ,
		\_2141__reg/NET0131 ,
		_w3287_
	);
	LUT3 #(
		.INIT('h82)
	) name1779 (
		RESET_pad,
		\WX3481_reg/NET0131 ,
		\_2142__reg/NET0131 ,
		_w3288_
	);
	LUT3 #(
		.INIT('h82)
	) name1780 (
		RESET_pad,
		\WX3479_reg/NET0131 ,
		\_2143__reg/NET0131 ,
		_w3289_
	);
	LUT3 #(
		.INIT('h82)
	) name1781 (
		RESET_pad,
		\WX3473_reg/NET0131 ,
		\_2146__reg/NET0131 ,
		_w3290_
	);
	LUT3 #(
		.INIT('h82)
	) name1782 (
		RESET_pad,
		\WX3471_reg/NET0131 ,
		\_2147__reg/NET0131 ,
		_w3291_
	);
	LUT3 #(
		.INIT('h82)
	) name1783 (
		RESET_pad,
		\WX3469_reg/NET0131 ,
		\_2148__reg/NET0131 ,
		_w3292_
	);
	LUT3 #(
		.INIT('h82)
	) name1784 (
		RESET_pad,
		\WX3465_reg/NET0131 ,
		\_2150__reg/NET0131 ,
		_w3293_
	);
	LUT3 #(
		.INIT('h82)
	) name1785 (
		RESET_pad,
		\WX3459_reg/NET0131 ,
		\_2153__reg/NET0131 ,
		_w3294_
	);
	LUT3 #(
		.INIT('h82)
	) name1786 (
		RESET_pad,
		\WX3457_reg/NET0131 ,
		\_2154__reg/NET0131 ,
		_w3295_
	);
	LUT3 #(
		.INIT('h82)
	) name1787 (
		RESET_pad,
		\WX3455_reg/NET0131 ,
		\_2155__reg/NET0131 ,
		_w3296_
	);
	LUT3 #(
		.INIT('h82)
	) name1788 (
		RESET_pad,
		\WX3451_reg/NET0131 ,
		\_2157__reg/NET0131 ,
		_w3297_
	);
	LUT3 #(
		.INIT('h82)
	) name1789 (
		RESET_pad,
		\WX3449_reg/NET0131 ,
		\_2158__reg/NET0131 ,
		_w3298_
	);
	LUT3 #(
		.INIT('h82)
	) name1790 (
		RESET_pad,
		\WX3445_reg/NET0131 ,
		\_2160__reg/NET0131 ,
		_w3299_
	);
	LUT3 #(
		.INIT('h82)
	) name1791 (
		RESET_pad,
		\WX3443_reg/NET0131 ,
		\_2161__reg/NET0131 ,
		_w3300_
	);
	LUT3 #(
		.INIT('h82)
	) name1792 (
		RESET_pad,
		\WX3441_reg/NET0131 ,
		\_2162__reg/NET0131 ,
		_w3301_
	);
	LUT3 #(
		.INIT('h82)
	) name1793 (
		RESET_pad,
		\WX3439_reg/NET0131 ,
		\_2163__reg/NET0131 ,
		_w3302_
	);
	LUT3 #(
		.INIT('h82)
	) name1794 (
		RESET_pad,
		\WX3437_reg/NET0131 ,
		\_2164__reg/NET0131 ,
		_w3303_
	);
	LUT3 #(
		.INIT('h82)
	) name1795 (
		RESET_pad,
		\WX3435_reg/NET0131 ,
		\_2165__reg/NET0131 ,
		_w3304_
	);
	LUT3 #(
		.INIT('h82)
	) name1796 (
		RESET_pad,
		\WX3433_reg/NET0131 ,
		\_2166__reg/NET0131 ,
		_w3305_
	);
	LUT3 #(
		.INIT('h82)
	) name1797 (
		RESET_pad,
		\WX3431_reg/NET0131 ,
		\_2167__reg/NET0131 ,
		_w3306_
	);
	LUT3 #(
		.INIT('h82)
	) name1798 (
		RESET_pad,
		\WX3429_reg/NET0131 ,
		\_2168__reg/NET0131 ,
		_w3307_
	);
	LUT3 #(
		.INIT('h82)
	) name1799 (
		RESET_pad,
		\WX3423_reg/NET0131 ,
		\_2171__reg/NET0131 ,
		_w3308_
	);
	LUT3 #(
		.INIT('h82)
	) name1800 (
		RESET_pad,
		\WX4778_reg/NET0131 ,
		\_2204__reg/NET0131 ,
		_w3309_
	);
	LUT3 #(
		.INIT('h82)
	) name1801 (
		RESET_pad,
		\WX4776_reg/NET0131 ,
		\_2173__reg/NET0131 ,
		_w3310_
	);
	LUT3 #(
		.INIT('h82)
	) name1802 (
		RESET_pad,
		\WX4774_reg/NET0131 ,
		\_2174__reg/NET0131 ,
		_w3311_
	);
	LUT3 #(
		.INIT('h82)
	) name1803 (
		RESET_pad,
		\WX4772_reg/NET0131 ,
		\_2175__reg/NET0131 ,
		_w3312_
	);
	LUT3 #(
		.INIT('h82)
	) name1804 (
		RESET_pad,
		\WX7316_reg/NET0131 ,
		\_2260__reg/NET0131 ,
		_w3313_
	);
	LUT3 #(
		.INIT('h82)
	) name1805 (
		RESET_pad,
		\WX4768_reg/NET0131 ,
		\_2177__reg/NET0131 ,
		_w3314_
	);
	LUT3 #(
		.INIT('h82)
	) name1806 (
		RESET_pad,
		\WX4766_reg/NET0131 ,
		\_2178__reg/NET0131 ,
		_w3315_
	);
	LUT3 #(
		.INIT('h82)
	) name1807 (
		RESET_pad,
		\WX4764_reg/NET0131 ,
		\_2179__reg/NET0131 ,
		_w3316_
	);
	LUT3 #(
		.INIT('h82)
	) name1808 (
		RESET_pad,
		\WX4760_reg/NET0131 ,
		\_2181__reg/NET0131 ,
		_w3317_
	);
	LUT3 #(
		.INIT('h82)
	) name1809 (
		RESET_pad,
		\WX4758_reg/NET0131 ,
		\_2182__reg/NET0131 ,
		_w3318_
	);
	LUT3 #(
		.INIT('h82)
	) name1810 (
		RESET_pad,
		\WX4754_reg/NET0131 ,
		\_2184__reg/NET0131 ,
		_w3319_
	);
	LUT3 #(
		.INIT('h82)
	) name1811 (
		RESET_pad,
		\WX4752_reg/NET0131 ,
		\_2185__reg/NET0131 ,
		_w3320_
	);
	LUT3 #(
		.INIT('h82)
	) name1812 (
		RESET_pad,
		\WX4750_reg/NET0131 ,
		\_2186__reg/NET0131 ,
		_w3321_
	);
	LUT3 #(
		.INIT('h82)
	) name1813 (
		RESET_pad,
		\WX4748_reg/NET0131 ,
		\_2187__reg/NET0131 ,
		_w3322_
	);
	LUT3 #(
		.INIT('h82)
	) name1814 (
		RESET_pad,
		\WX4744_reg/NET0131 ,
		\_2189__reg/NET0131 ,
		_w3323_
	);
	LUT3 #(
		.INIT('h82)
	) name1815 (
		RESET_pad,
		\WX4742_reg/NET0131 ,
		\_2190__reg/NET0131 ,
		_w3324_
	);
	LUT3 #(
		.INIT('h82)
	) name1816 (
		RESET_pad,
		\WX4740_reg/NET0131 ,
		\_2191__reg/NET0131 ,
		_w3325_
	);
	LUT3 #(
		.INIT('h82)
	) name1817 (
		RESET_pad,
		\WX4738_reg/NET0131 ,
		\_2192__reg/NET0131 ,
		_w3326_
	);
	LUT3 #(
		.INIT('h82)
	) name1818 (
		RESET_pad,
		\WX4736_reg/NET0131 ,
		\_2193__reg/NET0131 ,
		_w3327_
	);
	LUT3 #(
		.INIT('h82)
	) name1819 (
		RESET_pad,
		\WX4734_reg/NET0131 ,
		\_2194__reg/NET0131 ,
		_w3328_
	);
	LUT3 #(
		.INIT('h82)
	) name1820 (
		RESET_pad,
		\WX4732_reg/NET0131 ,
		\_2195__reg/NET0131 ,
		_w3329_
	);
	LUT3 #(
		.INIT('h82)
	) name1821 (
		RESET_pad,
		\WX4730_reg/NET0131 ,
		\_2196__reg/NET0131 ,
		_w3330_
	);
	LUT3 #(
		.INIT('h82)
	) name1822 (
		RESET_pad,
		\WX4724_reg/NET0131 ,
		\_2199__reg/NET0131 ,
		_w3331_
	);
	LUT3 #(
		.INIT('h82)
	) name1823 (
		RESET_pad,
		\WX4722_reg/NET0131 ,
		\_2200__reg/NET0131 ,
		_w3332_
	);
	LUT3 #(
		.INIT('h82)
	) name1824 (
		RESET_pad,
		\WX4720_reg/NET0131 ,
		\_2201__reg/NET0131 ,
		_w3333_
	);
	LUT3 #(
		.INIT('h82)
	) name1825 (
		RESET_pad,
		\WX4718_reg/NET0131 ,
		\_2202__reg/NET0131 ,
		_w3334_
	);
	LUT3 #(
		.INIT('h82)
	) name1826 (
		RESET_pad,
		\WX4716_reg/NET0131 ,
		\_2203__reg/NET0131 ,
		_w3335_
	);
	LUT3 #(
		.INIT('h82)
	) name1827 (
		RESET_pad,
		\WX6071_reg/NET0131 ,
		\_2236__reg/NET0131 ,
		_w3336_
	);
	LUT3 #(
		.INIT('h82)
	) name1828 (
		RESET_pad,
		\WX6067_reg/NET0131 ,
		\_2206__reg/NET0131 ,
		_w3337_
	);
	LUT3 #(
		.INIT('h82)
	) name1829 (
		RESET_pad,
		\WX6065_reg/NET0131 ,
		\_2207__reg/NET0131 ,
		_w3338_
	);
	LUT3 #(
		.INIT('h82)
	) name1830 (
		RESET_pad,
		\WX6059_reg/NET0131 ,
		\_2210__reg/NET0131 ,
		_w3339_
	);
	LUT3 #(
		.INIT('h82)
	) name1831 (
		RESET_pad,
		\WX6057_reg/NET0131 ,
		\_2211__reg/NET0131 ,
		_w3340_
	);
	LUT3 #(
		.INIT('h82)
	) name1832 (
		RESET_pad,
		\WX6055_reg/NET0131 ,
		\_2212__reg/NET0131 ,
		_w3341_
	);
	LUT3 #(
		.INIT('h82)
	) name1833 (
		RESET_pad,
		\WX6053_reg/NET0131 ,
		\_2213__reg/NET0131 ,
		_w3342_
	);
	LUT3 #(
		.INIT('h82)
	) name1834 (
		RESET_pad,
		\WX6051_reg/NET0131 ,
		\_2214__reg/NET0131 ,
		_w3343_
	);
	LUT3 #(
		.INIT('h82)
	) name1835 (
		RESET_pad,
		\WX6047_reg/NET0131 ,
		\_2216__reg/NET0131 ,
		_w3344_
	);
	LUT3 #(
		.INIT('h82)
	) name1836 (
		RESET_pad,
		\WX6045_reg/NET0131 ,
		\_2217__reg/NET0131 ,
		_w3345_
	);
	LUT3 #(
		.INIT('h82)
	) name1837 (
		RESET_pad,
		\WX6035_reg/NET0131 ,
		\_2222__reg/NET0131 ,
		_w3346_
	);
	LUT3 #(
		.INIT('h82)
	) name1838 (
		RESET_pad,
		\WX6033_reg/NET0131 ,
		\_2223__reg/NET0131 ,
		_w3347_
	);
	LUT3 #(
		.INIT('h82)
	) name1839 (
		RESET_pad,
		\WX6031_reg/NET0131 ,
		\_2224__reg/NET0131 ,
		_w3348_
	);
	LUT3 #(
		.INIT('h82)
	) name1840 (
		RESET_pad,
		\WX6029_reg/NET0131 ,
		\_2225__reg/NET0131 ,
		_w3349_
	);
	LUT3 #(
		.INIT('h82)
	) name1841 (
		RESET_pad,
		\WX6023_reg/NET0131 ,
		\_2228__reg/NET0131 ,
		_w3350_
	);
	LUT3 #(
		.INIT('h82)
	) name1842 (
		RESET_pad,
		\WX6021_reg/NET0131 ,
		\_2229__reg/NET0131 ,
		_w3351_
	);
	LUT3 #(
		.INIT('h82)
	) name1843 (
		RESET_pad,
		\WX6019_reg/NET0131 ,
		\_2230__reg/NET0131 ,
		_w3352_
	);
	LUT3 #(
		.INIT('h82)
	) name1844 (
		RESET_pad,
		\WX6015_reg/NET0131 ,
		\_2232__reg/NET0131 ,
		_w3353_
	);
	LUT3 #(
		.INIT('h82)
	) name1845 (
		RESET_pad,
		\WX6011_reg/NET0131 ,
		\_2234__reg/NET0131 ,
		_w3354_
	);
	LUT3 #(
		.INIT('h82)
	) name1846 (
		RESET_pad,
		\WX6009_reg/NET0131 ,
		\_2235__reg/NET0131 ,
		_w3355_
	);
	LUT3 #(
		.INIT('h82)
	) name1847 (
		RESET_pad,
		\WX7364_reg/NET0131 ,
		\_2268__reg/NET0131 ,
		_w3356_
	);
	LUT3 #(
		.INIT('h82)
	) name1848 (
		RESET_pad,
		\WX7360_reg/NET0131 ,
		\_2238__reg/NET0131 ,
		_w3357_
	);
	LUT3 #(
		.INIT('h82)
	) name1849 (
		RESET_pad,
		\WX7358_reg/NET0131 ,
		\_2239__reg/NET0131 ,
		_w3358_
	);
	LUT3 #(
		.INIT('h82)
	) name1850 (
		RESET_pad,
		\WX7354_reg/NET0131 ,
		\_2241__reg/NET0131 ,
		_w3359_
	);
	LUT3 #(
		.INIT('h82)
	) name1851 (
		RESET_pad,
		\WX7352_reg/NET0131 ,
		\_2242__reg/NET0131 ,
		_w3360_
	);
	LUT3 #(
		.INIT('h82)
	) name1852 (
		RESET_pad,
		\WX6025_reg/NET0131 ,
		\_2227__reg/NET0131 ,
		_w3361_
	);
	LUT3 #(
		.INIT('h82)
	) name1853 (
		RESET_pad,
		\WX8647_reg/NET0131 ,
		\_2273__reg/NET0131 ,
		_w3362_
	);
	LUT3 #(
		.INIT('h82)
	) name1854 (
		RESET_pad,
		\WX7336_reg/NET0131 ,
		\_2250__reg/NET0131 ,
		_w3363_
	);
	LUT3 #(
		.INIT('h82)
	) name1855 (
		RESET_pad,
		\WX7330_reg/NET0131 ,
		\_2253__reg/NET0131 ,
		_w3364_
	);
	LUT3 #(
		.INIT('h82)
	) name1856 (
		RESET_pad,
		\WX7326_reg/NET0131 ,
		\_2255__reg/NET0131 ,
		_w3365_
	);
	LUT3 #(
		.INIT('h82)
	) name1857 (
		RESET_pad,
		\WX7322_reg/NET0131 ,
		\_2257__reg/NET0131 ,
		_w3366_
	);
	LUT3 #(
		.INIT('h82)
	) name1858 (
		RESET_pad,
		\WX7320_reg/NET0131 ,
		\_2258__reg/NET0131 ,
		_w3367_
	);
	LUT3 #(
		.INIT('h82)
	) name1859 (
		RESET_pad,
		\WX7318_reg/NET0131 ,
		\_2259__reg/NET0131 ,
		_w3368_
	);
	LUT3 #(
		.INIT('h82)
	) name1860 (
		RESET_pad,
		\WX6069_reg/NET0131 ,
		\_2205__reg/NET0131 ,
		_w3369_
	);
	LUT3 #(
		.INIT('h82)
	) name1861 (
		RESET_pad,
		\WX7314_reg/NET0131 ,
		\_2261__reg/NET0131 ,
		_w3370_
	);
	LUT3 #(
		.INIT('h82)
	) name1862 (
		RESET_pad,
		\WX6017_reg/NET0131 ,
		\_2231__reg/NET0131 ,
		_w3371_
	);
	LUT3 #(
		.INIT('h82)
	) name1863 (
		RESET_pad,
		\WX6027_reg/NET0131 ,
		\_2226__reg/NET0131 ,
		_w3372_
	);
	LUT3 #(
		.INIT('h82)
	) name1864 (
		RESET_pad,
		\WX7306_reg/NET0131 ,
		\_2265__reg/NET0131 ,
		_w3373_
	);
	LUT3 #(
		.INIT('h82)
	) name1865 (
		RESET_pad,
		\WX7302_reg/NET0131 ,
		\_2267__reg/NET0131 ,
		_w3374_
	);
	LUT3 #(
		.INIT('h82)
	) name1866 (
		RESET_pad,
		\WX8655_reg/NET0131 ,
		\_2269__reg/NET0131 ,
		_w3375_
	);
	LUT3 #(
		.INIT('h82)
	) name1867 (
		RESET_pad,
		\WX8653_reg/NET0131 ,
		\_2270__reg/NET0131 ,
		_w3376_
	);
	LUT3 #(
		.INIT('h82)
	) name1868 (
		RESET_pad,
		\WX8651_reg/NET0131 ,
		\_2271__reg/NET0131 ,
		_w3377_
	);
	LUT3 #(
		.INIT('h82)
	) name1869 (
		RESET_pad,
		\WX8645_reg/NET0131 ,
		\_2274__reg/NET0131 ,
		_w3378_
	);
	LUT3 #(
		.INIT('h82)
	) name1870 (
		RESET_pad,
		\WX8641_reg/NET0131 ,
		\_2276__reg/NET0131 ,
		_w3379_
	);
	LUT3 #(
		.INIT('h82)
	) name1871 (
		RESET_pad,
		\WX8637_reg/NET0131 ,
		\_2278__reg/NET0131 ,
		_w3380_
	);
	LUT3 #(
		.INIT('h82)
	) name1872 (
		RESET_pad,
		\WX8631_reg/NET0131 ,
		\_2281__reg/NET0131 ,
		_w3381_
	);
	LUT3 #(
		.INIT('h82)
	) name1873 (
		RESET_pad,
		\WX8629_reg/NET0131 ,
		\_2282__reg/NET0131 ,
		_w3382_
	);
	LUT3 #(
		.INIT('h82)
	) name1874 (
		RESET_pad,
		\WX8627_reg/NET0131 ,
		\_2283__reg/NET0131 ,
		_w3383_
	);
	LUT3 #(
		.INIT('h82)
	) name1875 (
		RESET_pad,
		\WX8621_reg/NET0131 ,
		\_2286__reg/NET0131 ,
		_w3384_
	);
	LUT3 #(
		.INIT('h82)
	) name1876 (
		RESET_pad,
		\WX8617_reg/NET0131 ,
		\_2288__reg/NET0131 ,
		_w3385_
	);
	LUT3 #(
		.INIT('h82)
	) name1877 (
		RESET_pad,
		\WX8615_reg/NET0131 ,
		\_2289__reg/NET0131 ,
		_w3386_
	);
	LUT3 #(
		.INIT('h82)
	) name1878 (
		RESET_pad,
		\WX8613_reg/NET0131 ,
		\_2290__reg/NET0131 ,
		_w3387_
	);
	LUT3 #(
		.INIT('h82)
	) name1879 (
		RESET_pad,
		\WX8611_reg/NET0131 ,
		\_2291__reg/NET0131 ,
		_w3388_
	);
	LUT3 #(
		.INIT('h82)
	) name1880 (
		RESET_pad,
		\WX8609_reg/NET0131 ,
		\_2292__reg/NET0131 ,
		_w3389_
	);
	LUT3 #(
		.INIT('h82)
	) name1881 (
		RESET_pad,
		\WX8597_reg/NET0131 ,
		\_2298__reg/NET0131 ,
		_w3390_
	);
	LUT3 #(
		.INIT('h82)
	) name1882 (
		RESET_pad,
		\WX8595_reg/NET0131 ,
		\_2299__reg/NET0131 ,
		_w3391_
	);
	LUT3 #(
		.INIT('h82)
	) name1883 (
		RESET_pad,
		\WX9950_reg/NET0131 ,
		\_2332__reg/NET0131 ,
		_w3392_
	);
	LUT3 #(
		.INIT('h82)
	) name1884 (
		RESET_pad,
		\WX9948_reg/NET0131 ,
		\_2301__reg/NET0131 ,
		_w3393_
	);
	LUT3 #(
		.INIT('h82)
	) name1885 (
		RESET_pad,
		\WX9946_reg/NET0131 ,
		\_2302__reg/NET0131 ,
		_w3394_
	);
	LUT3 #(
		.INIT('h82)
	) name1886 (
		RESET_pad,
		\WX9940_reg/NET0131 ,
		\_2305__reg/NET0131 ,
		_w3395_
	);
	LUT3 #(
		.INIT('h82)
	) name1887 (
		RESET_pad,
		\WX9938_reg/NET0131 ,
		\_2306__reg/NET0131 ,
		_w3396_
	);
	LUT3 #(
		.INIT('h82)
	) name1888 (
		RESET_pad,
		\WX9932_reg/NET0131 ,
		\_2309__reg/NET0131 ,
		_w3397_
	);
	LUT3 #(
		.INIT('h82)
	) name1889 (
		RESET_pad,
		\WX9926_reg/NET0131 ,
		\_2312__reg/NET0131 ,
		_w3398_
	);
	LUT3 #(
		.INIT('h82)
	) name1890 (
		RESET_pad,
		\WX9922_reg/NET0131 ,
		\_2314__reg/NET0131 ,
		_w3399_
	);
	LUT3 #(
		.INIT('h82)
	) name1891 (
		RESET_pad,
		\WX9920_reg/NET0131 ,
		\_2315__reg/NET0131 ,
		_w3400_
	);
	LUT3 #(
		.INIT('h82)
	) name1892 (
		RESET_pad,
		\WX9916_reg/NET0131 ,
		\_2317__reg/NET0131 ,
		_w3401_
	);
	LUT3 #(
		.INIT('h82)
	) name1893 (
		RESET_pad,
		\WX9914_reg/NET0131 ,
		\_2318__reg/NET0131 ,
		_w3402_
	);
	LUT3 #(
		.INIT('h82)
	) name1894 (
		RESET_pad,
		\WX9912_reg/NET0131 ,
		\_2319__reg/NET0131 ,
		_w3403_
	);
	LUT3 #(
		.INIT('h82)
	) name1895 (
		RESET_pad,
		\WX9910_reg/NET0131 ,
		\_2320__reg/NET0131 ,
		_w3404_
	);
	LUT3 #(
		.INIT('h82)
	) name1896 (
		RESET_pad,
		\WX9908_reg/NET0131 ,
		\_2321__reg/NET0131 ,
		_w3405_
	);
	LUT3 #(
		.INIT('h82)
	) name1897 (
		RESET_pad,
		\WX9906_reg/NET0131 ,
		\_2322__reg/NET0131 ,
		_w3406_
	);
	LUT3 #(
		.INIT('h82)
	) name1898 (
		RESET_pad,
		\WX9904_reg/NET0131 ,
		\_2323__reg/NET0131 ,
		_w3407_
	);
	LUT3 #(
		.INIT('h82)
	) name1899 (
		RESET_pad,
		\WX9902_reg/NET0131 ,
		\_2324__reg/NET0131 ,
		_w3408_
	);
	LUT3 #(
		.INIT('h82)
	) name1900 (
		RESET_pad,
		\WX9900_reg/NET0131 ,
		\_2325__reg/NET0131 ,
		_w3409_
	);
	LUT3 #(
		.INIT('h82)
	) name1901 (
		RESET_pad,
		\WX9898_reg/NET0131 ,
		\_2326__reg/NET0131 ,
		_w3410_
	);
	LUT3 #(
		.INIT('h82)
	) name1902 (
		RESET_pad,
		\WX9896_reg/NET0131 ,
		\_2327__reg/NET0131 ,
		_w3411_
	);
	LUT3 #(
		.INIT('h82)
	) name1903 (
		RESET_pad,
		\WX9894_reg/NET0131 ,
		\_2328__reg/NET0131 ,
		_w3412_
	);
	LUT3 #(
		.INIT('h82)
	) name1904 (
		RESET_pad,
		\WX9892_reg/NET0131 ,
		\_2329__reg/NET0131 ,
		_w3413_
	);
	LUT3 #(
		.INIT('h82)
	) name1905 (
		RESET_pad,
		\WX9888_reg/NET0131 ,
		\_2331__reg/NET0131 ,
		_w3414_
	);
	LUT3 #(
		.INIT('h82)
	) name1906 (
		RESET_pad,
		\WX11243_reg/NET0131 ,
		\_2364__reg/NET0131 ,
		_w3415_
	);
	LUT3 #(
		.INIT('h82)
	) name1907 (
		RESET_pad,
		\WX11241_reg/NET0131 ,
		\_2333__reg/NET0131 ,
		_w3416_
	);
	LUT3 #(
		.INIT('h82)
	) name1908 (
		RESET_pad,
		\WX11239_reg/NET0131 ,
		\_2334__reg/NET0131 ,
		_w3417_
	);
	LUT3 #(
		.INIT('h82)
	) name1909 (
		RESET_pad,
		\WX11237_reg/NET0131 ,
		\_2335__reg/NET0131 ,
		_w3418_
	);
	LUT3 #(
		.INIT('h82)
	) name1910 (
		RESET_pad,
		\WX11233_reg/NET0131 ,
		\_2337__reg/NET0131 ,
		_w3419_
	);
	LUT3 #(
		.INIT('h82)
	) name1911 (
		RESET_pad,
		\WX11231_reg/NET0131 ,
		\_2338__reg/NET0131 ,
		_w3420_
	);
	LUT3 #(
		.INIT('h82)
	) name1912 (
		RESET_pad,
		\WX11229_reg/NET0131 ,
		\_2339__reg/NET0131 ,
		_w3421_
	);
	LUT3 #(
		.INIT('h82)
	) name1913 (
		RESET_pad,
		\WX11227_reg/NET0131 ,
		\_2340__reg/NET0131 ,
		_w3422_
	);
	LUT3 #(
		.INIT('h82)
	) name1914 (
		RESET_pad,
		\WX11225_reg/NET0131 ,
		\_2341__reg/NET0131 ,
		_w3423_
	);
	LUT3 #(
		.INIT('h82)
	) name1915 (
		RESET_pad,
		\WX11223_reg/NET0131 ,
		\_2342__reg/NET0131 ,
		_w3424_
	);
	LUT3 #(
		.INIT('h82)
	) name1916 (
		RESET_pad,
		\WX11219_reg/NET0131 ,
		\_2344__reg/NET0131 ,
		_w3425_
	);
	LUT3 #(
		.INIT('h82)
	) name1917 (
		RESET_pad,
		\WX11217_reg/NET0131 ,
		\_2345__reg/NET0131 ,
		_w3426_
	);
	LUT3 #(
		.INIT('h82)
	) name1918 (
		RESET_pad,
		\WX11213_reg/NET0131 ,
		\_2347__reg/NET0131 ,
		_w3427_
	);
	LUT3 #(
		.INIT('h82)
	) name1919 (
		RESET_pad,
		\WX11209_reg/NET0131 ,
		\_2349__reg/NET0131 ,
		_w3428_
	);
	LUT3 #(
		.INIT('h82)
	) name1920 (
		RESET_pad,
		\WX11207_reg/NET0131 ,
		\_2350__reg/NET0131 ,
		_w3429_
	);
	LUT3 #(
		.INIT('h82)
	) name1921 (
		RESET_pad,
		\WX11205_reg/NET0131 ,
		\_2351__reg/NET0131 ,
		_w3430_
	);
	LUT3 #(
		.INIT('h82)
	) name1922 (
		RESET_pad,
		\WX11203_reg/NET0131 ,
		\_2352__reg/NET0131 ,
		_w3431_
	);
	LUT3 #(
		.INIT('h82)
	) name1923 (
		RESET_pad,
		\WX11201_reg/NET0131 ,
		\_2353__reg/NET0131 ,
		_w3432_
	);
	LUT3 #(
		.INIT('h82)
	) name1924 (
		RESET_pad,
		\WX11199_reg/NET0131 ,
		\_2354__reg/NET0131 ,
		_w3433_
	);
	LUT3 #(
		.INIT('h82)
	) name1925 (
		RESET_pad,
		\WX11197_reg/NET0131 ,
		\_2355__reg/NET0131 ,
		_w3434_
	);
	LUT3 #(
		.INIT('h82)
	) name1926 (
		RESET_pad,
		\WX11195_reg/NET0131 ,
		\_2356__reg/NET0131 ,
		_w3435_
	);
	LUT3 #(
		.INIT('h82)
	) name1927 (
		RESET_pad,
		\WX11193_reg/NET0131 ,
		\_2357__reg/NET0131 ,
		_w3436_
	);
	LUT3 #(
		.INIT('h82)
	) name1928 (
		RESET_pad,
		\WX11191_reg/NET0131 ,
		\_2358__reg/NET0131 ,
		_w3437_
	);
	LUT3 #(
		.INIT('h82)
	) name1929 (
		RESET_pad,
		\WX11189_reg/NET0131 ,
		\_2359__reg/NET0131 ,
		_w3438_
	);
	LUT3 #(
		.INIT('h82)
	) name1930 (
		RESET_pad,
		\WX11187_reg/NET0131 ,
		\_2360__reg/NET0131 ,
		_w3439_
	);
	LUT3 #(
		.INIT('h82)
	) name1931 (
		RESET_pad,
		\WX11183_reg/NET0131 ,
		\_2362__reg/NET0131 ,
		_w3440_
	);
	LUT3 #(
		.INIT('h82)
	) name1932 (
		RESET_pad,
		\WX2150_reg/NET0131 ,
		\_2129__reg/NET0131 ,
		_w3441_
	);
	LUT3 #(
		.INIT('h82)
	) name1933 (
		RESET_pad,
		\WX7304_reg/NET0131 ,
		\_2266__reg/NET0131 ,
		_w3442_
	);
	LUT3 #(
		.INIT('h82)
	) name1934 (
		RESET_pad,
		\WX2136_reg/NET0131 ,
		\_2136__reg/NET0131 ,
		_w3443_
	);
	LUT3 #(
		.INIT('h82)
	) name1935 (
		RESET_pad,
		\WX3467_reg/NET0131 ,
		\_2149__reg/NET0131 ,
		_w3444_
	);
	LUT3 #(
		.INIT('h82)
	) name1936 (
		RESET_pad,
		\WX8633_reg/NET0131 ,
		\_2280__reg/NET0131 ,
		_w3445_
	);
	LUT3 #(
		.INIT('h82)
	) name1937 (
		RESET_pad,
		\WX853_reg/NET0131 ,
		\_2099__reg/NET0131 ,
		_w3446_
	);
	LUT3 #(
		.INIT('h82)
	) name1938 (
		RESET_pad,
		\WX859_reg/NET0131 ,
		\_2096__reg/NET0131 ,
		_w3447_
	);
	LUT3 #(
		.INIT('h82)
	) name1939 (
		RESET_pad,
		\WX7310_reg/NET0131 ,
		\_2263__reg/NET0131 ,
		_w3448_
	);
	LUT3 #(
		.INIT('h82)
	) name1940 (
		RESET_pad,
		\WX9936_reg/NET0131 ,
		\_2307__reg/NET0131 ,
		_w3449_
	);
	LUT3 #(
		.INIT('h82)
	) name1941 (
		RESET_pad,
		\WX849_reg/NET0131 ,
		\_2101__reg/NET0131 ,
		_w3450_
	);
	LUT3 #(
		.INIT('h82)
	) name1942 (
		RESET_pad,
		\WX2140_reg/NET0131 ,
		\_2134__reg/NET0131 ,
		_w3451_
	);
	LUT3 #(
		.INIT('h82)
	) name1943 (
		RESET_pad,
		\WX2178_reg/NET0131 ,
		\_2115__reg/NET0131 ,
		_w3452_
	);
	LUT3 #(
		.INIT('h82)
	) name1944 (
		RESET_pad,
		\WX8623_reg/NET0131 ,
		\_2285__reg/NET0131 ,
		_w3453_
	);
	LUT3 #(
		.INIT('h82)
	) name1945 (
		RESET_pad,
		\WX2176_reg/NET0131 ,
		\_2116__reg/NET0131 ,
		_w3454_
	);
	LUT3 #(
		.INIT('h82)
	) name1946 (
		RESET_pad,
		\WX7346_reg/NET0131 ,
		\_2245__reg/NET0131 ,
		_w3455_
	);
	LUT3 #(
		.INIT('h82)
	) name1947 (
		RESET_pad,
		\WX6041_reg/NET0131 ,
		\_2219__reg/NET0131 ,
		_w3456_
	);
	LUT3 #(
		.INIT('h82)
	) name1948 (
		RESET_pad,
		\WX7350_reg/NET0131 ,
		\_2243__reg/NET0131 ,
		_w3457_
	);
	LUT3 #(
		.INIT('h82)
	) name1949 (
		RESET_pad,
		\WX4762_reg/NET0131 ,
		\_2180__reg/NET0131 ,
		_w3458_
	);
	LUT3 #(
		.INIT('h82)
	) name1950 (
		RESET_pad,
		\WX871_reg/NET0131 ,
		\_2090__reg/NET0131 ,
		_w3459_
	);
	LUT3 #(
		.INIT('h82)
	) name1951 (
		RESET_pad,
		\WX885_reg/NET0131 ,
		\_2083__reg/NET0131 ,
		_w3460_
	);
	LUT3 #(
		.INIT('h82)
	) name1952 (
		RESET_pad,
		\WX11185_reg/NET0131 ,
		\_2361__reg/NET0131 ,
		_w3461_
	);
	LUT3 #(
		.INIT('h82)
	) name1953 (
		RESET_pad,
		\WX9890_reg/NET0131 ,
		\_2330__reg/NET0131 ,
		_w3462_
	);
	LUT3 #(
		.INIT('h82)
	) name1954 (
		RESET_pad,
		\WX9944_reg/NET0131 ,
		\_2303__reg/NET0131 ,
		_w3463_
	);
	LUT3 #(
		.INIT('h82)
	) name1955 (
		RESET_pad,
		\WX7344_reg/NET0131 ,
		\_2246__reg/NET0131 ,
		_w3464_
	);
	LUT3 #(
		.INIT('h82)
	) name1956 (
		RESET_pad,
		\WX7324_reg/NET0131 ,
		\_2256__reg/NET0131 ,
		_w3465_
	);
	LUT3 #(
		.INIT('h82)
	) name1957 (
		RESET_pad,
		\WX6013_reg/NET0131 ,
		\_2233__reg/NET0131 ,
		_w3466_
	);
	LUT3 #(
		.INIT('h82)
	) name1958 (
		RESET_pad,
		\WX2152_reg/NET0131 ,
		\_2128__reg/NET0131 ,
		_w3467_
	);
	LUT3 #(
		.INIT('h82)
	) name1959 (
		RESET_pad,
		\WX847_reg/NET0131 ,
		\_2102__reg/NET0131 ,
		_w3468_
	);
	LUT3 #(
		.INIT('h82)
	) name1960 (
		RESET_pad,
		\WX3447_reg/NET0131 ,
		\_2159__reg/NET0131 ,
		_w3469_
	);
	LUT3 #(
		.INIT('h82)
	) name1961 (
		RESET_pad,
		\WX9924_reg/NET0131 ,
		\_2313__reg/NET0131 ,
		_w3470_
	);
	LUT3 #(
		.INIT('h82)
	) name1962 (
		RESET_pad,
		\WX861_reg/NET0131 ,
		\_2095__reg/NET0131 ,
		_w3471_
	);
	LUT3 #(
		.INIT('h82)
	) name1963 (
		RESET_pad,
		\WX8639_reg/NET0131 ,
		\_2277__reg/NET0131 ,
		_w3472_
	);
	LUT3 #(
		.INIT('h82)
	) name1964 (
		RESET_pad,
		\WX7308_reg/NET0131 ,
		\_2264__reg/NET0131 ,
		_w3473_
	);
	LUT3 #(
		.INIT('h82)
	) name1965 (
		RESET_pad,
		\WX879_reg/NET0131 ,
		\_2086__reg/NET0131 ,
		_w3474_
	);
	LUT3 #(
		.INIT('h82)
	) name1966 (
		RESET_pad,
		\WX7334_reg/NET0131 ,
		\_2251__reg/NET0131 ,
		_w3475_
	);
	LUT3 #(
		.INIT('h82)
	) name1967 (
		RESET_pad,
		\WX8643_reg/NET0131 ,
		\_2275__reg/NET0131 ,
		_w3476_
	);
	LUT3 #(
		.INIT('h82)
	) name1968 (
		RESET_pad,
		\WX4726_reg/NET0131 ,
		\_2198__reg/NET0131 ,
		_w3477_
	);
	LUT2 #(
		.INIT('h8)
	) name1969 (
		RESET_pad,
		\WX11053_reg/NET0131 ,
		_w3478_
	);
	LUT2 #(
		.INIT('h8)
	) name1970 (
		RESET_pad,
		\WX709_reg/NET0131 ,
		_w3479_
	);
	LUT2 #(
		.INIT('h8)
	) name1971 (
		RESET_pad,
		\WX10891_reg/NET0131 ,
		_w3480_
	);
	LUT2 #(
		.INIT('h8)
	) name1972 (
		RESET_pad,
		\WX2002_reg/NET0131 ,
		_w3481_
	);
	LUT2 #(
		.INIT('h2)
	) name1973 (
		RESET_pad,
		\WX10829_reg/NET0131 ,
		_w3482_
	);
	LUT2 #(
		.INIT('h8)
	) name1974 (
		RESET_pad,
		\WX11059_reg/NET0131 ,
		_w3483_
	);
	LUT2 #(
		.INIT('h8)
	) name1975 (
		RESET_pad,
		\WX3271_reg/NET0131 ,
		_w3484_
	);
	LUT2 #(
		.INIT('h8)
	) name1976 (
		RESET_pad,
		\WX11033_reg/NET0131 ,
		_w3485_
	);
	LUT2 #(
		.INIT('h8)
	) name1977 (
		RESET_pad,
		\WX7252_reg/NET0131 ,
		_w3486_
	);
	LUT2 #(
		.INIT('h8)
	) name1978 (
		RESET_pad,
		\WX3257_reg/NET0131 ,
		_w3487_
	);
	LUT2 #(
		.INIT('h8)
	) name1979 (
		RESET_pad,
		\WX3403_reg/NET0131 ,
		_w3488_
	);
	LUT2 #(
		.INIT('h8)
	) name1980 (
		RESET_pad,
		\WX11115_reg/NET0131 ,
		_w3489_
	);
	LUT2 #(
		.INIT('h8)
	) name1981 (
		RESET_pad,
		\WX11049_reg/NET0131 ,
		_w3490_
	);
	LUT2 #(
		.INIT('h8)
	) name1982 (
		RESET_pad,
		\WX9714_reg/NET0131 ,
		_w3491_
	);
	LUT2 #(
		.INIT('h8)
	) name1983 (
		RESET_pad,
		\WX2004_reg/NET0131 ,
		_w3492_
	);
	LUT2 #(
		.INIT('h8)
	) name1984 (
		RESET_pad,
		\WX11037_reg/NET0131 ,
		_w3493_
	);
	LUT2 #(
		.INIT('h8)
	) name1985 (
		RESET_pad,
		\WX9852_reg/NET0131 ,
		_w3494_
	);
	LUT2 #(
		.INIT('h8)
	) name1986 (
		RESET_pad,
		\WX9702_reg/NET0131 ,
		_w3495_
	);
	LUT2 #(
		.INIT('h8)
	) name1987 (
		RESET_pad,
		\WX9876_reg/NET0131 ,
		_w3496_
	);
	LUT2 #(
		.INIT('h8)
	) name1988 (
		RESET_pad,
		\WX11121_reg/NET0131 ,
		_w3497_
	);
	LUT2 #(
		.INIT('h8)
	) name1989 (
		RESET_pad,
		\WX7114_reg/NET0131 ,
		_w3498_
	);
	LUT2 #(
		.INIT('h8)
	) name1990 (
		RESET_pad,
		\WX1986_reg/NET0131 ,
		_w3499_
	);
	LUT2 #(
		.INIT('h8)
	) name1991 (
		RESET_pad,
		\WX9802_reg/NET0131 ,
		_w3500_
	);
	LUT2 #(
		.INIT('h8)
	) name1992 (
		RESET_pad,
		\WX9824_reg/NET0131 ,
		_w3501_
	);
	LUT2 #(
		.INIT('h8)
	) name1993 (
		RESET_pad,
		\WX7220_reg/NET0131 ,
		_w3502_
	);
	LUT2 #(
		.INIT('h8)
	) name1994 (
		RESET_pad,
		\WX9806_reg/NET0131 ,
		_w3503_
	);
	LUT2 #(
		.INIT('h8)
	) name1995 (
		RESET_pad,
		\WX11073_reg/NET0131 ,
		_w3504_
	);
	LUT2 #(
		.INIT('h8)
	) name1996 (
		RESET_pad,
		\WX9878_reg/NET0131 ,
		_w3505_
	);
	LUT2 #(
		.INIT('h8)
	) name1997 (
		RESET_pad,
		\WX11111_reg/NET0131 ,
		_w3506_
	);
	LUT2 #(
		.INIT('h8)
	) name1998 (
		RESET_pad,
		\WX11169_reg/NET0131 ,
		_w3507_
	);
	LUT2 #(
		.INIT('h8)
	) name1999 (
		RESET_pad,
		\WX1998_reg/NET0131 ,
		_w3508_
	);
	LUT2 #(
		.INIT('h8)
	) name2000 (
		RESET_pad,
		\WX9850_reg/NET0131 ,
		_w3509_
	);
	LUT2 #(
		.INIT('h8)
	) name2001 (
		RESET_pad,
		\WX11079_reg/NET0131 ,
		_w3510_
	);
	LUT2 #(
		.INIT('h8)
	) name2002 (
		RESET_pad,
		\WX7110_reg/NET0131 ,
		_w3511_
	);
	LUT2 #(
		.INIT('h8)
	) name2003 (
		RESET_pad,
		\WX7240_reg/NET0131 ,
		_w3512_
	);
	LUT2 #(
		.INIT('h8)
	) name2004 (
		RESET_pad,
		\WX1954_reg/NET0131 ,
		_w3513_
	);
	LUT2 #(
		.INIT('h8)
	) name2005 (
		RESET_pad,
		\WX11081_reg/NET0131 ,
		_w3514_
	);
	LUT2 #(
		.INIT('h8)
	) name2006 (
		RESET_pad,
		\WX11083_reg/NET0131 ,
		_w3515_
	);
	LUT2 #(
		.INIT('h8)
	) name2007 (
		RESET_pad,
		\WX3339_reg/NET0131 ,
		_w3516_
	);
	LUT2 #(
		.INIT('h8)
	) name2008 (
		RESET_pad,
		\WX8491_reg/NET0131 ,
		_w3517_
	);
	LUT2 #(
		.INIT('h8)
	) name2009 (
		RESET_pad,
		\WX11175_reg/NET0131 ,
		_w3518_
	);
	LUT2 #(
		.INIT('h8)
	) name2010 (
		RESET_pad,
		\WX11089_reg/NET0131 ,
		_w3519_
	);
	LUT2 #(
		.INIT('h8)
	) name2011 (
		RESET_pad,
		\WX9770_reg/NET0131 ,
		_w3520_
	);
	LUT2 #(
		.INIT('h8)
	) name2012 (
		RESET_pad,
		\WX2068_reg/NET0131 ,
		_w3521_
	);
	LUT2 #(
		.INIT('h8)
	) name2013 (
		RESET_pad,
		\WX823_reg/NET0131 ,
		_w3522_
	);
	LUT2 #(
		.INIT('h8)
	) name2014 (
		RESET_pad,
		\WX5941_reg/NET0131 ,
		_w3523_
	);
	LUT2 #(
		.INIT('h8)
	) name2015 (
		RESET_pad,
		\WX11093_reg/NET0131 ,
		_w3524_
	);
	LUT2 #(
		.INIT('h8)
	) name2016 (
		RESET_pad,
		\WX5919_reg/NET0131 ,
		_w3525_
	);
	LUT2 #(
		.INIT('h8)
	) name2017 (
		RESET_pad,
		\WX7160_reg/NET0131 ,
		_w3526_
	);
	LUT2 #(
		.INIT('h8)
	) name2018 (
		RESET_pad,
		\WX791_reg/NET0131 ,
		_w3527_
	);
	LUT2 #(
		.INIT('h8)
	) name2019 (
		RESET_pad,
		\WX11095_reg/NET0131 ,
		_w3528_
	);
	LUT2 #(
		.INIT('h8)
	) name2020 (
		RESET_pad,
		\WX3349_reg/NET0131 ,
		_w3529_
	);
	LUT2 #(
		.INIT('h8)
	) name2021 (
		RESET_pad,
		\WX9708_reg/NET0131 ,
		_w3530_
	);
	LUT2 #(
		.INIT('h8)
	) name2022 (
		RESET_pad,
		\WX769_reg/NET0131 ,
		_w3531_
	);
	LUT2 #(
		.INIT('h8)
	) name2023 (
		RESET_pad,
		\WX11153_reg/NET0131 ,
		_w3532_
	);
	LUT2 #(
		.INIT('h8)
	) name2024 (
		RESET_pad,
		\WX7182_reg/NET0131 ,
		_w3533_
	);
	LUT2 #(
		.INIT('h8)
	) name2025 (
		RESET_pad,
		\WX7238_reg/NET0131 ,
		_w3534_
	);
	LUT2 #(
		.INIT('h8)
	) name2026 (
		RESET_pad,
		\WX11103_reg/NET0131 ,
		_w3535_
	);
	LUT2 #(
		.INIT('h8)
	) name2027 (
		RESET_pad,
		\WX5925_reg/NET0131 ,
		_w3536_
	);
	LUT2 #(
		.INIT('h8)
	) name2028 (
		RESET_pad,
		\WX7196_reg/NET0131 ,
		_w3537_
	);
	LUT2 #(
		.INIT('h8)
	) name2029 (
		RESET_pad,
		\WX7204_reg/NET0131 ,
		_w3538_
	);
	LUT2 #(
		.INIT('h8)
	) name2030 (
		RESET_pad,
		\WX3279_reg/NET0131 ,
		_w3539_
	);
	LUT2 #(
		.INIT('h8)
	) name2031 (
		RESET_pad,
		\WX5953_reg/NET0131 ,
		_w3540_
	);
	LUT2 #(
		.INIT('h8)
	) name2032 (
		RESET_pad,
		\WX3285_reg/NET0131 ,
		_w3541_
	);
	LUT2 #(
		.INIT('h8)
	) name2033 (
		RESET_pad,
		\WX4594_reg/NET0131 ,
		_w3542_
	);
	LUT2 #(
		.INIT('h8)
	) name2034 (
		RESET_pad,
		\WX777_reg/NET0131 ,
		_w3543_
	);
	LUT2 #(
		.INIT('h8)
	) name2035 (
		RESET_pad,
		\WX7164_reg/NET0131 ,
		_w3544_
	);
	LUT2 #(
		.INIT('h8)
	) name2036 (
		RESET_pad,
		\WX11167_reg/NET0131 ,
		_w3545_
	);
	LUT2 #(
		.INIT('h8)
	) name2037 (
		RESET_pad,
		\WX719_reg/NET0131 ,
		_w3546_
	);
	LUT2 #(
		.INIT('h8)
	) name2038 (
		RESET_pad,
		\WX707_reg/NET0131 ,
		_w3547_
	);
	LUT2 #(
		.INIT('h8)
	) name2039 (
		RESET_pad,
		\WX7294_reg/NET0131 ,
		_w3548_
	);
	LUT2 #(
		.INIT('h8)
	) name2040 (
		RESET_pad,
		\WX11113_reg/NET0131 ,
		_w3549_
	);
	LUT2 #(
		.INIT('h8)
	) name2041 (
		RESET_pad,
		\WX1988_reg/NET0131 ,
		_w3550_
	);
	LUT2 #(
		.INIT('h8)
	) name2042 (
		RESET_pad,
		\WX7234_reg/NET0131 ,
		_w3551_
	);
	LUT2 #(
		.INIT('h8)
	) name2043 (
		RESET_pad,
		\WX9712_reg/NET0131 ,
		_w3552_
	);
	LUT2 #(
		.INIT('h8)
	) name2044 (
		RESET_pad,
		\WX5929_reg/NET0131 ,
		_w3553_
	);
	LUT2 #(
		.INIT('h8)
	) name2045 (
		RESET_pad,
		\WX7244_reg/NET0131 ,
		_w3554_
	);
	LUT2 #(
		.INIT('h8)
	) name2046 (
		RESET_pad,
		\WX7248_reg/NET0131 ,
		_w3555_
	);
	LUT2 #(
		.INIT('h8)
	) name2047 (
		RESET_pad,
		\WX9882_reg/NET0131 ,
		_w3556_
	);
	LUT2 #(
		.INIT('h8)
	) name2048 (
		RESET_pad,
		\WX4550_reg/NET0131 ,
		_w3557_
	);
	LUT2 #(
		.INIT('h8)
	) name2049 (
		RESET_pad,
		\WX665_reg/NET0131 ,
		_w3558_
	);
	LUT2 #(
		.INIT('h8)
	) name2050 (
		RESET_pad,
		\WX7232_reg/NET0131 ,
		_w3559_
	);
	LUT2 #(
		.INIT('h8)
	) name2051 (
		RESET_pad,
		\WX705_reg/NET0131 ,
		_w3560_
	);
	LUT2 #(
		.INIT('h8)
	) name2052 (
		RESET_pad,
		\WX2064_reg/NET0131 ,
		_w3561_
	);
	LUT2 #(
		.INIT('h8)
	) name2053 (
		RESET_pad,
		\WX5927_reg/NET0131 ,
		_w3562_
	);
	LUT2 #(
		.INIT('h8)
	) name2054 (
		RESET_pad,
		\WX9822_reg/NET0131 ,
		_w3563_
	);
	LUT2 #(
		.INIT('h8)
	) name2055 (
		RESET_pad,
		\WX7276_reg/NET0131 ,
		_w3564_
	);
	LUT2 #(
		.INIT('h8)
	) name2056 (
		RESET_pad,
		\WX3277_reg/NET0131 ,
		_w3565_
	);
	LUT2 #(
		.INIT('h8)
	) name2057 (
		RESET_pad,
		\WX7284_reg/NET0131 ,
		_w3566_
	);
	LUT2 #(
		.INIT('h8)
	) name2058 (
		RESET_pad,
		\WX11177_reg/NET0131 ,
		_w3567_
	);
	LUT2 #(
		.INIT('h8)
	) name2059 (
		RESET_pad,
		\WX645_reg/NET0131 ,
		_w3568_
	);
	LUT2 #(
		.INIT('h8)
	) name2060 (
		RESET_pad,
		\WX11133_reg/NET0131 ,
		_w3569_
	);
	LUT2 #(
		.INIT('h8)
	) name2061 (
		RESET_pad,
		\WX1992_reg/NET0131 ,
		_w3570_
	);
	LUT2 #(
		.INIT('h8)
	) name2062 (
		RESET_pad,
		\WX11135_reg/NET0131 ,
		_w3571_
	);
	LUT2 #(
		.INIT('h8)
	) name2063 (
		RESET_pad,
		\WX11137_reg/NET0131 ,
		_w3572_
	);
	LUT2 #(
		.INIT('h8)
	) name2064 (
		RESET_pad,
		\WX2072_reg/NET0131 ,
		_w3573_
	);
	LUT2 #(
		.INIT('h8)
	) name2065 (
		RESET_pad,
		\WX11161_reg/NET0131 ,
		_w3574_
	);
	LUT2 #(
		.INIT('h8)
	) name2066 (
		RESET_pad,
		\WX5933_reg/NET0131 ,
		_w3575_
	);
	LUT2 #(
		.INIT('h8)
	) name2067 (
		RESET_pad,
		\WX3379_reg/NET0131 ,
		_w3576_
	);
	LUT2 #(
		.INIT('h8)
	) name2068 (
		RESET_pad,
		\WX4556_reg/NET0131 ,
		_w3577_
	);
	LUT2 #(
		.INIT('h8)
	) name2069 (
		RESET_pad,
		\WX11143_reg/NET0131 ,
		_w3578_
	);
	LUT2 #(
		.INIT('h8)
	) name2070 (
		RESET_pad,
		\WX9750_reg/NET0131 ,
		_w3579_
	);
	LUT2 #(
		.INIT('h8)
	) name2071 (
		RESET_pad,
		\WX9786_reg/NET0131 ,
		_w3580_
	);
	LUT2 #(
		.INIT('h8)
	) name2072 (
		RESET_pad,
		\WX7230_reg/NET0131 ,
		_w3581_
	);
	LUT2 #(
		.INIT('h8)
	) name2073 (
		RESET_pad,
		\WX3237_reg/NET0131 ,
		_w3582_
	);
	LUT2 #(
		.INIT('h8)
	) name2074 (
		RESET_pad,
		\WX11041_reg/NET0131 ,
		_w3583_
	);
	LUT2 #(
		.INIT('h8)
	) name2075 (
		RESET_pad,
		\WX5939_reg/NET0131 ,
		_w3584_
	);
	LUT2 #(
		.INIT('h8)
	) name2076 (
		RESET_pad,
		\WX9716_reg/NET0131 ,
		_w3585_
	);
	LUT2 #(
		.INIT('h8)
	) name2077 (
		RESET_pad,
		\WX5871_reg/NET0131 ,
		_w3586_
	);
	LUT2 #(
		.INIT('h8)
	) name2078 (
		RESET_pad,
		\WX757_reg/NET0131 ,
		_w3587_
	);
	LUT2 #(
		.INIT('h8)
	) name2079 (
		RESET_pad,
		\WX11045_reg/NET0131 ,
		_w3588_
	);
	LUT2 #(
		.INIT('h8)
	) name2080 (
		RESET_pad,
		\WX9744_reg/NET0131 ,
		_w3589_
	);
	LUT2 #(
		.INIT('h8)
	) name2081 (
		RESET_pad,
		\WX9762_reg/NET0131 ,
		_w3590_
	);
	LUT2 #(
		.INIT('h8)
	) name2082 (
		RESET_pad,
		\WX4558_reg/NET0131 ,
		_w3591_
	);
	LUT2 #(
		.INIT('h8)
	) name2083 (
		RESET_pad,
		\WX3273_reg/NET0131 ,
		_w3592_
	);
	LUT2 #(
		.INIT('h8)
	) name2084 (
		RESET_pad,
		\WX5945_reg/NET0131 ,
		_w3593_
	);
	LUT2 #(
		.INIT('h8)
	) name2085 (
		RESET_pad,
		\WX9860_reg/NET0131 ,
		_w3594_
	);
	LUT2 #(
		.INIT('h8)
	) name2086 (
		RESET_pad,
		\WX7228_reg/NET0131 ,
		_w3595_
	);
	LUT2 #(
		.INIT('h8)
	) name2087 (
		RESET_pad,
		\WX7226_reg/NET0131 ,
		_w3596_
	);
	LUT2 #(
		.INIT('h8)
	) name2088 (
		RESET_pad,
		\WX4542_reg/NET0131 ,
		_w3597_
	);
	LUT2 #(
		.INIT('h8)
	) name2089 (
		RESET_pad,
		\WX9808_reg/NET0131 ,
		_w3598_
	);
	LUT2 #(
		.INIT('h8)
	) name2090 (
		RESET_pad,
		\WX11109_reg/NET0131 ,
		_w3599_
	);
	LUT2 #(
		.INIT('h8)
	) name2091 (
		RESET_pad,
		\WX8423_reg/NET0131 ,
		_w3600_
	);
	LUT2 #(
		.INIT('h8)
	) name2092 (
		RESET_pad,
		\WX3327_reg/NET0131 ,
		_w3601_
	);
	LUT2 #(
		.INIT('h8)
	) name2093 (
		RESET_pad,
		\WX807_reg/NET0131 ,
		_w3602_
	);
	LUT2 #(
		.INIT('h8)
	) name2094 (
		RESET_pad,
		\WX8533_reg/NET0131 ,
		_w3603_
	);
	LUT2 #(
		.INIT('h8)
	) name2095 (
		RESET_pad,
		\WX7222_reg/NET0131 ,
		_w3604_
	);
	LUT2 #(
		.INIT('h8)
	) name2096 (
		RESET_pad,
		\WX9856_reg/NET0131 ,
		_w3605_
	);
	LUT2 #(
		.INIT('h8)
	) name2097 (
		RESET_pad,
		\WX1984_reg/NET0131 ,
		_w3606_
	);
	LUT2 #(
		.INIT('h8)
	) name2098 (
		RESET_pad,
		\WX7118_reg/NET0131 ,
		_w3607_
	);
	LUT2 #(
		.INIT('h8)
	) name2099 (
		RESET_pad,
		\WX7218_reg/NET0131 ,
		_w3608_
	);
	LUT2 #(
		.INIT('h8)
	) name2100 (
		RESET_pad,
		\WX7224_reg/NET0131 ,
		_w3609_
	);
	LUT2 #(
		.INIT('h8)
	) name2101 (
		RESET_pad,
		\WX4544_reg/NET0131 ,
		_w3610_
	);
	LUT2 #(
		.INIT('h8)
	) name2102 (
		RESET_pad,
		\WX4560_reg/NET0131 ,
		_w3611_
	);
	LUT2 #(
		.INIT('h8)
	) name2103 (
		RESET_pad,
		\WX667_reg/NET0131 ,
		_w3612_
	);
	LUT2 #(
		.INIT('h8)
	) name2104 (
		RESET_pad,
		\WX7214_reg/NET0131 ,
		_w3613_
	);
	LUT2 #(
		.INIT('h8)
	) name2105 (
		RESET_pad,
		\WX3319_reg/NET0131 ,
		_w3614_
	);
	LUT2 #(
		.INIT('h8)
	) name2106 (
		RESET_pad,
		\WX663_reg/NET0131 ,
		_w3615_
	);
	LUT2 #(
		.INIT('h8)
	) name2107 (
		RESET_pad,
		\WX4598_reg/NET0131 ,
		_w3616_
	);
	LUT2 #(
		.INIT('h8)
	) name2108 (
		RESET_pad,
		\WX9820_reg/NET0131 ,
		_w3617_
	);
	LUT2 #(
		.INIT('h8)
	) name2109 (
		RESET_pad,
		\WX5979_reg/NET0131 ,
		_w3618_
	);
	LUT2 #(
		.INIT('h8)
	) name2110 (
		RESET_pad,
		\WX11107_reg/NET0131 ,
		_w3619_
	);
	LUT2 #(
		.INIT('h8)
	) name2111 (
		RESET_pad,
		\WX9698_reg/NET0131 ,
		_w3620_
	);
	LUT2 #(
		.INIT('h8)
	) name2112 (
		RESET_pad,
		\WX7198_reg/NET0131 ,
		_w3621_
	);
	LUT2 #(
		.INIT('h8)
	) name2113 (
		RESET_pad,
		\WX3365_reg/NET0131 ,
		_w3622_
	);
	LUT2 #(
		.INIT('h8)
	) name2114 (
		RESET_pad,
		\WX11131_reg/NET0131 ,
		_w3623_
	);
	LUT2 #(
		.INIT('h8)
	) name2115 (
		RESET_pad,
		\WX3361_reg/NET0131 ,
		_w3624_
	);
	LUT2 #(
		.INIT('h8)
	) name2116 (
		RESET_pad,
		\WX11163_reg/NET0131 ,
		_w3625_
	);
	LUT2 #(
		.INIT('h8)
	) name2117 (
		RESET_pad,
		\WX8517_reg/NET0131 ,
		_w3626_
	);
	LUT2 #(
		.INIT('h8)
	) name2118 (
		RESET_pad,
		\WX9772_reg/NET0131 ,
		_w3627_
	);
	LUT2 #(
		.INIT('h8)
	) name2119 (
		RESET_pad,
		\WX11105_reg/NET0131 ,
		_w3628_
	);
	LUT2 #(
		.INIT('h8)
	) name2120 (
		RESET_pad,
		\WX11123_reg/NET0131 ,
		_w3629_
	);
	LUT2 #(
		.INIT('h8)
	) name2121 (
		RESET_pad,
		\WX3351_reg/NET0131 ,
		_w3630_
	);
	LUT2 #(
		.INIT('h8)
	) name2122 (
		RESET_pad,
		\WX4562_reg/NET0131 ,
		_w3631_
	);
	LUT2 #(
		.INIT('h8)
	) name2123 (
		RESET_pad,
		\WX4540_reg/NET0131 ,
		_w3632_
	);
	LUT2 #(
		.INIT('h8)
	) name2124 (
		RESET_pad,
		\WX5879_reg/NET0131 ,
		_w3633_
	);
	LUT2 #(
		.INIT('h8)
	) name2125 (
		RESET_pad,
		\WX5875_reg/NET0131 ,
		_w3634_
	);
	LUT2 #(
		.INIT('h8)
	) name2126 (
		RESET_pad,
		\WX5991_reg/NET0131 ,
		_w3635_
	);
	LUT2 #(
		.INIT('h8)
	) name2127 (
		RESET_pad,
		\WX2056_reg/NET0131 ,
		_w3636_
	);
	LUT2 #(
		.INIT('h8)
	) name2128 (
		RESET_pad,
		\WX3263_reg/NET0131 ,
		_w3637_
	);
	LUT2 #(
		.INIT('h8)
	) name2129 (
		RESET_pad,
		\WX7166_reg/NET0131 ,
		_w3638_
	);
	LUT2 #(
		.INIT('h8)
	) name2130 (
		RESET_pad,
		\WX7190_reg/NET0131 ,
		_w3639_
	);
	LUT2 #(
		.INIT('h8)
	) name2131 (
		RESET_pad,
		\WX1972_reg/NET0131 ,
		_w3640_
	);
	LUT2 #(
		.INIT('h8)
	) name2132 (
		RESET_pad,
		\WX661_reg/NET0131 ,
		_w3641_
	);
	LUT2 #(
		.INIT('h8)
	) name2133 (
		RESET_pad,
		\WX9774_reg/NET0131 ,
		_w3642_
	);
	LUT2 #(
		.INIT('h8)
	) name2134 (
		RESET_pad,
		\WX1994_reg/NET0131 ,
		_w3643_
	);
	LUT2 #(
		.INIT('h8)
	) name2135 (
		RESET_pad,
		\WX7256_reg/NET0131 ,
		_w3644_
	);
	LUT2 #(
		.INIT('h8)
	) name2136 (
		RESET_pad,
		\WX5985_reg/NET0131 ,
		_w3645_
	);
	LUT2 #(
		.INIT('h8)
	) name2137 (
		RESET_pad,
		\WX7192_reg/NET0131 ,
		_w3646_
	);
	LUT2 #(
		.INIT('h8)
	) name2138 (
		RESET_pad,
		\WX7194_reg/NET0131 ,
		_w3647_
	);
	LUT2 #(
		.INIT('h8)
	) name2139 (
		RESET_pad,
		\WX8445_reg/NET0131 ,
		_w3648_
	);
	LUT2 #(
		.INIT('h8)
	) name2140 (
		RESET_pad,
		\WX5999_reg/NET0131 ,
		_w3649_
	);
	LUT2 #(
		.INIT('h8)
	) name2141 (
		RESET_pad,
		\WX1966_reg/NET0131 ,
		_w3650_
	);
	LUT2 #(
		.INIT('h8)
	) name2142 (
		RESET_pad,
		\WX9726_reg/NET0131 ,
		_w3651_
	);
	LUT2 #(
		.INIT('h8)
	) name2143 (
		RESET_pad,
		\WX9704_reg/NET0131 ,
		_w3652_
	);
	LUT2 #(
		.INIT('h8)
	) name2144 (
		RESET_pad,
		\WX7186_reg/NET0131 ,
		_w3653_
	);
	LUT2 #(
		.INIT('h8)
	) name2145 (
		RESET_pad,
		\WX8441_reg/NET0131 ,
		_w3654_
	);
	LUT2 #(
		.INIT('h8)
	) name2146 (
		RESET_pad,
		\WX5923_reg/NET0131 ,
		_w3655_
	);
	LUT2 #(
		.INIT('h8)
	) name2147 (
		RESET_pad,
		\WX2128_reg/NET0131 ,
		_w3656_
	);
	LUT2 #(
		.INIT('h8)
	) name2148 (
		RESET_pad,
		\WX2126_reg/NET0131 ,
		_w3657_
	);
	LUT2 #(
		.INIT('h8)
	) name2149 (
		RESET_pad,
		\WX7180_reg/NET0131 ,
		_w3658_
	);
	LUT2 #(
		.INIT('h8)
	) name2150 (
		RESET_pad,
		\WX721_reg/NET0131 ,
		_w3659_
	);
	LUT2 #(
		.INIT('h8)
	) name2151 (
		RESET_pad,
		\WX7278_reg/NET0131 ,
		_w3660_
	);
	LUT2 #(
		.INIT('h8)
	) name2152 (
		RESET_pad,
		\WX835_reg/NET0131 ,
		_w3661_
	);
	LUT2 #(
		.INIT('h8)
	) name2153 (
		RESET_pad,
		\WX5997_reg/NET0131 ,
		_w3662_
	);
	LUT2 #(
		.INIT('h8)
	) name2154 (
		RESET_pad,
		\WX3363_reg/NET0131 ,
		_w3663_
	);
	LUT2 #(
		.INIT('h8)
	) name2155 (
		RESET_pad,
		\WX5921_reg/NET0131 ,
		_w3664_
	);
	LUT2 #(
		.INIT('h8)
	) name2156 (
		RESET_pad,
		\WX659_reg/NET0131 ,
		_w3665_
	);
	LUT2 #(
		.INIT('h8)
	) name2157 (
		RESET_pad,
		\WX3259_reg/NET0131 ,
		_w3666_
	);
	LUT2 #(
		.INIT('h8)
	) name2158 (
		RESET_pad,
		\WX9780_reg/NET0131 ,
		_w3667_
	);
	LUT2 #(
		.INIT('h8)
	) name2159 (
		RESET_pad,
		\WX1956_reg/NET0131 ,
		_w3668_
	);
	LUT2 #(
		.INIT('h8)
	) name2160 (
		RESET_pad,
		\WX11099_reg/NET0131 ,
		_w3669_
	);
	LUT2 #(
		.INIT('h8)
	) name2161 (
		RESET_pad,
		\WX2088_reg/NET0131 ,
		_w3670_
	);
	LUT2 #(
		.INIT('h8)
	) name2162 (
		RESET_pad,
		\WX9800_reg/NET0131 ,
		_w3671_
	);
	LUT2 #(
		.INIT('h8)
	) name2163 (
		RESET_pad,
		\WX767_reg/NET0131 ,
		_w3672_
	);
	LUT2 #(
		.INIT('h8)
	) name2164 (
		RESET_pad,
		\WX7280_reg/NET0131 ,
		_w3673_
	);
	LUT2 #(
		.INIT('h8)
	) name2165 (
		RESET_pad,
		\WX8519_reg/NET0131 ,
		_w3674_
	);
	LUT2 #(
		.INIT('h8)
	) name2166 (
		RESET_pad,
		\WX771_reg/NET0131 ,
		_w3675_
	);
	LUT2 #(
		.INIT('h8)
	) name2167 (
		RESET_pad,
		\WX781_reg/NET0131 ,
		_w3676_
	);
	LUT2 #(
		.INIT('h8)
	) name2168 (
		RESET_pad,
		\WX1958_reg/NET0131 ,
		_w3677_
	);
	LUT2 #(
		.INIT('h8)
	) name2169 (
		RESET_pad,
		\WX3289_reg/NET0131 ,
		_w3678_
	);
	LUT2 #(
		.INIT('h8)
	) name2170 (
		RESET_pad,
		\WX4638_reg/NET0131 ,
		_w3679_
	);
	LUT2 #(
		.INIT('h8)
	) name2171 (
		RESET_pad,
		\WX687_reg/NET0131 ,
		_w3680_
	);
	LUT2 #(
		.INIT('h8)
	) name2172 (
		RESET_pad,
		\WX2112_reg/NET0131 ,
		_w3681_
	);
	LUT2 #(
		.INIT('h8)
	) name2173 (
		RESET_pad,
		\WX9730_reg/NET0131 ,
		_w3682_
	);
	LUT2 #(
		.INIT('h8)
	) name2174 (
		RESET_pad,
		\WX9754_reg/NET0131 ,
		_w3683_
	);
	LUT2 #(
		.INIT('h8)
	) name2175 (
		RESET_pad,
		\WX787_reg/NET0131 ,
		_w3684_
	);
	LUT2 #(
		.INIT('h8)
	) name2176 (
		RESET_pad,
		\WX731_reg/NET0131 ,
		_w3685_
	);
	LUT2 #(
		.INIT('h8)
	) name2177 (
		RESET_pad,
		\WX3415_reg/NET0131 ,
		_w3686_
	);
	LUT2 #(
		.INIT('h8)
	) name2178 (
		RESET_pad,
		\WX3255_reg/NET0131 ,
		_w3687_
	);
	LUT2 #(
		.INIT('h8)
	) name2179 (
		RESET_pad,
		\WX2122_reg/NET0131 ,
		_w3688_
	);
	LUT2 #(
		.INIT('h8)
	) name2180 (
		RESET_pad,
		\WX8529_reg/NET0131 ,
		_w3689_
	);
	LUT2 #(
		.INIT('h8)
	) name2181 (
		RESET_pad,
		\WX9832_reg/NET0131 ,
		_w3690_
	);
	LUT2 #(
		.INIT('h8)
	) name2182 (
		RESET_pad,
		\WX8449_reg/NET0131 ,
		_w3691_
	);
	LUT2 #(
		.INIT('h8)
	) name2183 (
		RESET_pad,
		\WX727_reg/NET0131 ,
		_w3692_
	);
	LUT2 #(
		.INIT('h8)
	) name2184 (
		RESET_pad,
		\WX7158_reg/NET0131 ,
		_w3693_
	);
	LUT2 #(
		.INIT('h8)
	) name2185 (
		RESET_pad,
		\WX11011_reg/NET0131 ,
		_w3694_
	);
	LUT2 #(
		.INIT('h8)
	) name2186 (
		RESET_pad,
		\WX7152_reg/NET0131 ,
		_w3695_
	);
	LUT2 #(
		.INIT('h8)
	) name2187 (
		RESET_pad,
		\WX4676_reg/NET0131 ,
		_w3696_
	);
	LUT2 #(
		.INIT('h8)
	) name2188 (
		RESET_pad,
		\WX7156_reg/NET0131 ,
		_w3697_
	);
	LUT2 #(
		.INIT('h8)
	) name2189 (
		RESET_pad,
		\WX7154_reg/NET0131 ,
		_w3698_
	);
	LUT2 #(
		.INIT('h8)
	) name2190 (
		RESET_pad,
		\WX657_reg/NET0131 ,
		_w3699_
	);
	LUT2 #(
		.INIT('h8)
	) name2191 (
		RESET_pad,
		\WX9816_reg/NET0131 ,
		_w3700_
	);
	LUT2 #(
		.INIT('h8)
	) name2192 (
		RESET_pad,
		\WX831_reg/NET0131 ,
		_w3701_
	);
	LUT2 #(
		.INIT('h8)
	) name2193 (
		RESET_pad,
		\WX7134_reg/NET0131 ,
		_w3702_
	);
	LUT2 #(
		.INIT('h8)
	) name2194 (
		RESET_pad,
		\WX7246_reg/NET0131 ,
		_w3703_
	);
	LUT2 #(
		.INIT('h8)
	) name2195 (
		RESET_pad,
		\WX7144_reg/NET0131 ,
		_w3704_
	);
	LUT2 #(
		.INIT('h8)
	) name2196 (
		RESET_pad,
		\WX9736_reg/NET0131 ,
		_w3705_
	);
	LUT2 #(
		.INIT('h8)
	) name2197 (
		RESET_pad,
		\WX1946_reg/NET0131 ,
		_w3706_
	);
	LUT2 #(
		.INIT('h8)
	) name2198 (
		RESET_pad,
		\WX7150_reg/NET0131 ,
		_w3707_
	);
	LUT2 #(
		.INIT('h8)
	) name2199 (
		RESET_pad,
		\WX2000_reg/NET0131 ,
		_w3708_
	);
	LUT2 #(
		.INIT('h8)
	) name2200 (
		RESET_pad,
		\WX761_reg/NET0131 ,
		_w3709_
	);
	LUT2 #(
		.INIT('h8)
	) name2201 (
		RESET_pad,
		\WX9842_reg/NET0131 ,
		_w3710_
	);
	LUT2 #(
		.INIT('h8)
	) name2202 (
		RESET_pad,
		\WX819_reg/NET0131 ,
		_w3711_
	);
	LUT2 #(
		.INIT('h8)
	) name2203 (
		RESET_pad,
		\WX7148_reg/NET0131 ,
		_w3712_
	);
	LUT2 #(
		.INIT('h8)
	) name2204 (
		RESET_pad,
		\WX3321_reg/NET0131 ,
		_w3713_
	);
	LUT2 #(
		.INIT('h8)
	) name2205 (
		RESET_pad,
		\WX4634_reg/NET0131 ,
		_w3714_
	);
	LUT2 #(
		.INIT('h8)
	) name2206 (
		RESET_pad,
		\WX11087_reg/NET0131 ,
		_w3715_
	);
	LUT2 #(
		.INIT('h8)
	) name2207 (
		RESET_pad,
		\WX7124_reg/NET0131 ,
		_w3716_
	);
	LUT2 #(
		.INIT('h8)
	) name2208 (
		RESET_pad,
		\WX3301_reg/NET0131 ,
		_w3717_
	);
	LUT2 #(
		.INIT('h8)
	) name2209 (
		RESET_pad,
		\WX3409_reg/NET0131 ,
		_w3718_
	);
	LUT2 #(
		.INIT('h8)
	) name2210 (
		RESET_pad,
		\WX9778_reg/NET0131 ,
		_w3719_
	);
	LUT2 #(
		.INIT('h8)
	) name2211 (
		RESET_pad,
		\WX7272_reg/NET0131 ,
		_w3720_
	);
	LUT2 #(
		.INIT('h8)
	) name2212 (
		RESET_pad,
		\WX7138_reg/NET0131 ,
		_w3721_
	);
	LUT2 #(
		.INIT('h8)
	) name2213 (
		RESET_pad,
		\WX2118_reg/NET0131 ,
		_w3722_
	);
	LUT2 #(
		.INIT('h8)
	) name2214 (
		RESET_pad,
		\WX4626_reg/NET0131 ,
		_w3723_
	);
	LUT2 #(
		.INIT('h8)
	) name2215 (
		RESET_pad,
		\WX5949_reg/NET0131 ,
		_w3724_
	);
	LUT2 #(
		.INIT('h8)
	) name2216 (
		RESET_pad,
		\WX693_reg/NET0131 ,
		_w3725_
	);
	LUT2 #(
		.INIT('h8)
	) name2217 (
		RESET_pad,
		\WX3265_reg/NET0131 ,
		_w3726_
	);
	LUT2 #(
		.INIT('h8)
	) name2218 (
		RESET_pad,
		\WX11141_reg/NET0131 ,
		_w3727_
	);
	LUT2 #(
		.INIT('h8)
	) name2219 (
		RESET_pad,
		\WX5947_reg/NET0131 ,
		_w3728_
	);
	LUT2 #(
		.INIT('h8)
	) name2220 (
		RESET_pad,
		\WX2114_reg/NET0131 ,
		_w3729_
	);
	LUT2 #(
		.INIT('h8)
	) name2221 (
		RESET_pad,
		\WX4584_reg/NET0131 ,
		_w3730_
	);
	LUT2 #(
		.INIT('h8)
	) name2222 (
		RESET_pad,
		\WX735_reg/NET0131 ,
		_w3731_
	);
	LUT2 #(
		.INIT('h8)
	) name2223 (
		RESET_pad,
		\WX3267_reg/NET0131 ,
		_w3732_
	);
	LUT2 #(
		.INIT('h8)
	) name2224 (
		RESET_pad,
		\WX7120_reg/NET0131 ,
		_w3733_
	);
	LUT2 #(
		.INIT('h8)
	) name2225 (
		RESET_pad,
		\WX7132_reg/NET0131 ,
		_w3734_
	);
	LUT2 #(
		.INIT('h8)
	) name2226 (
		RESET_pad,
		\WX3357_reg/NET0131 ,
		_w3735_
	);
	LUT2 #(
		.INIT('h8)
	) name2227 (
		RESET_pad,
		\WX3281_reg/NET0131 ,
		_w3736_
	);
	LUT2 #(
		.INIT('h8)
	) name2228 (
		RESET_pad,
		\WX3247_reg/NET0131 ,
		_w3737_
	);
	LUT2 #(
		.INIT('h8)
	) name2229 (
		RESET_pad,
		\WX9798_reg/NET0131 ,
		_w3738_
	);
	LUT2 #(
		.INIT('h8)
	) name2230 (
		RESET_pad,
		\WX11119_reg/NET0131 ,
		_w3739_
	);
	LUT2 #(
		.INIT('h8)
	) name2231 (
		RESET_pad,
		\WX7126_reg/NET0131 ,
		_w3740_
	);
	LUT2 #(
		.INIT('h8)
	) name2232 (
		RESET_pad,
		\WX5937_reg/NET0131 ,
		_w3741_
	);
	LUT2 #(
		.INIT('h8)
	) name2233 (
		RESET_pad,
		\WX7128_reg/NET0131 ,
		_w3742_
	);
	LUT2 #(
		.INIT('h8)
	) name2234 (
		RESET_pad,
		\WX3347_reg/NET0131 ,
		_w3743_
	);
	LUT2 #(
		.INIT('h8)
	) name2235 (
		RESET_pad,
		\WX2060_reg/NET0131 ,
		_w3744_
	);
	LUT2 #(
		.INIT('h8)
	) name2236 (
		RESET_pad,
		\WX7130_reg/NET0131 ,
		_w3745_
	);
	LUT2 #(
		.INIT('h8)
	) name2237 (
		RESET_pad,
		\WX9742_reg/NET0131 ,
		_w3746_
	);
	LUT2 #(
		.INIT('h8)
	) name2238 (
		RESET_pad,
		\WX11085_reg/NET0131 ,
		_w3747_
	);
	LUT2 #(
		.INIT('h8)
	) name2239 (
		RESET_pad,
		\WX11043_reg/NET0131 ,
		_w3748_
	);
	LUT2 #(
		.INIT('h8)
	) name2240 (
		RESET_pad,
		\WX3283_reg/NET0131 ,
		_w3749_
	);
	LUT2 #(
		.INIT('h8)
	) name2241 (
		RESET_pad,
		\WX755_reg/NET0131 ,
		_w3750_
	);
	LUT2 #(
		.INIT('h8)
	) name2242 (
		RESET_pad,
		\WX8447_reg/NET0131 ,
		_w3751_
	);
	LUT2 #(
		.INIT('h8)
	) name2243 (
		RESET_pad,
		\WX669_reg/NET0131 ,
		_w3752_
	);
	LUT2 #(
		.INIT('h8)
	) name2244 (
		RESET_pad,
		\WX4564_reg/NET0131 ,
		_w3753_
	);
	LUT2 #(
		.INIT('h8)
	) name2245 (
		RESET_pad,
		\WX685_reg/NET0131 ,
		_w3754_
	);
	LUT2 #(
		.INIT('h8)
	) name2246 (
		RESET_pad,
		\WX11067_reg/NET0131 ,
		_w3755_
	);
	LUT2 #(
		.INIT('h8)
	) name2247 (
		RESET_pad,
		\WX8453_reg/NET0131 ,
		_w3756_
	);
	LUT2 #(
		.INIT('h8)
	) name2248 (
		RESET_pad,
		\WX4538_reg/NET0131 ,
		_w3757_
	);
	LUT2 #(
		.INIT('h8)
	) name2249 (
		RESET_pad,
		\WX5959_reg/NET0131 ,
		_w3758_
	);
	LUT2 #(
		.INIT('h8)
	) name2250 (
		RESET_pad,
		\WX3355_reg/NET0131 ,
		_w3759_
	);
	LUT2 #(
		.INIT('h8)
	) name2251 (
		RESET_pad,
		\WX4588_reg/NET0131 ,
		_w3760_
	);
	LUT2 #(
		.INIT('h8)
	) name2252 (
		RESET_pad,
		\WX9724_reg/NET0131 ,
		_w3761_
	);
	LUT2 #(
		.INIT('h8)
	) name2253 (
		RESET_pad,
		\WX5965_reg/NET0131 ,
		_w3762_
	);
	LUT2 #(
		.INIT('h8)
	) name2254 (
		RESET_pad,
		\WX11147_reg/NET0131 ,
		_w3763_
	);
	LUT2 #(
		.INIT('h8)
	) name2255 (
		RESET_pad,
		\WX7122_reg/NET0131 ,
		_w3764_
	);
	LUT2 #(
		.INIT('h8)
	) name2256 (
		RESET_pad,
		\WX695_reg/NET0131 ,
		_w3765_
	);
	LUT2 #(
		.INIT('h8)
	) name2257 (
		RESET_pad,
		\WX4636_reg/NET0131 ,
		_w3766_
	);
	LUT2 #(
		.INIT('h8)
	) name2258 (
		RESET_pad,
		\WX4628_reg/NET0131 ,
		_w3767_
	);
	LUT2 #(
		.INIT('h8)
	) name2259 (
		RESET_pad,
		\WX8551_reg/NET0131 ,
		_w3768_
	);
	LUT2 #(
		.INIT('h8)
	) name2260 (
		RESET_pad,
		\WX9872_reg/NET0131 ,
		_w3769_
	);
	LUT2 #(
		.INIT('h8)
	) name2261 (
		RESET_pad,
		\WX5861_reg/NET0131 ,
		_w3770_
	);
	LUT2 #(
		.INIT('h8)
	) name2262 (
		RESET_pad,
		\WX8407_reg/NET0131 ,
		_w3771_
	);
	LUT2 #(
		.INIT('h8)
	) name2263 (
		RESET_pad,
		\WX8547_reg/NET0131 ,
		_w3772_
	);
	LUT2 #(
		.INIT('h8)
	) name2264 (
		RESET_pad,
		\WX9862_reg/NET0131 ,
		_w3773_
	);
	LUT2 #(
		.INIT('h8)
	) name2265 (
		RESET_pad,
		\WX4570_reg/NET0131 ,
		_w3774_
	);
	LUT2 #(
		.INIT('h8)
	) name2266 (
		RESET_pad,
		\WX11027_reg/NET0131 ,
		_w3775_
	);
	LUT2 #(
		.INIT('h8)
	) name2267 (
		RESET_pad,
		\WX11139_reg/NET0131 ,
		_w3776_
	);
	LUT2 #(
		.INIT('h8)
	) name2268 (
		RESET_pad,
		\WX4652_reg/NET0131 ,
		_w3777_
	);
	LUT2 #(
		.INIT('h8)
	) name2269 (
		RESET_pad,
		\WX729_reg/NET0131 ,
		_w3778_
	);
	LUT2 #(
		.INIT('h8)
	) name2270 (
		RESET_pad,
		\WX5957_reg/NET0131 ,
		_w3779_
	);
	LUT2 #(
		.INIT('h8)
	) name2271 (
		RESET_pad,
		\WX3287_reg/NET0131 ,
		_w3780_
	);
	LUT2 #(
		.INIT('h8)
	) name2272 (
		RESET_pad,
		\WX801_reg/NET0131 ,
		_w3781_
	);
	LUT2 #(
		.INIT('h8)
	) name2273 (
		RESET_pad,
		\WX805_reg/NET0131 ,
		_w3782_
	);
	LUT2 #(
		.INIT('h8)
	) name2274 (
		RESET_pad,
		\WX11149_reg/NET0131 ,
		_w3783_
	);
	LUT2 #(
		.INIT('h8)
	) name2275 (
		RESET_pad,
		\WX691_reg/NET0131 ,
		_w3784_
	);
	LUT2 #(
		.INIT('h8)
	) name2276 (
		RESET_pad,
		\WX8557_reg/NET0131 ,
		_w3785_
	);
	LUT2 #(
		.INIT('h8)
	) name2277 (
		RESET_pad,
		\WX9722_reg/NET0131 ,
		_w3786_
	);
	LUT2 #(
		.INIT('h8)
	) name2278 (
		RESET_pad,
		\WX9840_reg/NET0131 ,
		_w3787_
	);
	LUT2 #(
		.INIT('h8)
	) name2279 (
		RESET_pad,
		\WX9764_reg/NET0131 ,
		_w3788_
	);
	LUT2 #(
		.INIT('h8)
	) name2280 (
		RESET_pad,
		\WX2076_reg/NET0131 ,
		_w3789_
	);
	LUT2 #(
		.INIT('h8)
	) name2281 (
		RESET_pad,
		\WX7116_reg/NET0131 ,
		_w3790_
	);
	LUT2 #(
		.INIT('h8)
	) name2282 (
		RESET_pad,
		\WX9796_reg/NET0131 ,
		_w3791_
	);
	LUT2 #(
		.INIT('h8)
	) name2283 (
		RESET_pad,
		\WX9776_reg/NET0131 ,
		_w3792_
	);
	LUT2 #(
		.INIT('h8)
	) name2284 (
		RESET_pad,
		\WX11071_reg/NET0131 ,
		_w3793_
	);
	LUT2 #(
		.INIT('h8)
	) name2285 (
		RESET_pad,
		\WX9760_reg/NET0131 ,
		_w3794_
	);
	LUT2 #(
		.INIT('h8)
	) name2286 (
		RESET_pad,
		\WX4576_reg/NET0131 ,
		_w3795_
	);
	LUT2 #(
		.INIT('h8)
	) name2287 (
		RESET_pad,
		\WX803_reg/NET0131 ,
		_w3796_
	);
	LUT2 #(
		.INIT('h8)
	) name2288 (
		RESET_pad,
		\WX3395_reg/NET0131 ,
		_w3797_
	);
	LUT2 #(
		.INIT('h8)
	) name2289 (
		RESET_pad,
		\WX4526_reg/NET0131 ,
		_w3798_
	);
	LUT2 #(
		.INIT('h8)
	) name2290 (
		RESET_pad,
		\WX9790_reg/NET0131 ,
		_w3799_
	);
	LUT2 #(
		.INIT('h8)
	) name2291 (
		RESET_pad,
		\WX9768_reg/NET0131 ,
		_w3800_
	);
	LUT2 #(
		.INIT('h8)
	) name2292 (
		RESET_pad,
		\WX653_reg/NET0131 ,
		_w3801_
	);
	LUT2 #(
		.INIT('h8)
	) name2293 (
		RESET_pad,
		\WX4662_reg/NET0131 ,
		_w3802_
	);
	LUT2 #(
		.INIT('h8)
	) name2294 (
		RESET_pad,
		\WX4580_reg/NET0131 ,
		_w3803_
	);
	LUT2 #(
		.INIT('h8)
	) name2295 (
		RESET_pad,
		\WX9728_reg/NET0131 ,
		_w3804_
	);
	LUT2 #(
		.INIT('h8)
	) name2296 (
		RESET_pad,
		\WX9718_reg/NET0131 ,
		_w3805_
	);
	LUT2 #(
		.INIT('h8)
	) name2297 (
		RESET_pad,
		\WX3405_reg/NET0131 ,
		_w3806_
	);
	LUT2 #(
		.INIT('h8)
	) name2298 (
		RESET_pad,
		\WX3245_reg/NET0131 ,
		_w3807_
	);
	LUT2 #(
		.INIT('h8)
	) name2299 (
		RESET_pad,
		\WX2010_reg/NET0131 ,
		_w3808_
	);
	LUT2 #(
		.INIT('h8)
	) name2300 (
		RESET_pad,
		\WX4682_reg/NET0131 ,
		_w3809_
	);
	LUT2 #(
		.INIT('h8)
	) name2301 (
		RESET_pad,
		\WX8589_reg/NET0131 ,
		_w3810_
	);
	LUT2 #(
		.INIT('h8)
	) name2302 (
		RESET_pad,
		\WX4688_reg/NET0131 ,
		_w3811_
	);
	LUT2 #(
		.INIT('h8)
	) name2303 (
		RESET_pad,
		\WX9706_reg/NET0131 ,
		_w3812_
	);
	LUT2 #(
		.INIT('h8)
	) name2304 (
		RESET_pad,
		\WX4690_reg/NET0131 ,
		_w3813_
	);
	LUT2 #(
		.INIT('h8)
	) name2305 (
		RESET_pad,
		\WX3243_reg/NET0131 ,
		_w3814_
	);
	LUT2 #(
		.INIT('h8)
	) name2306 (
		RESET_pad,
		\WX3241_reg/NET0131 ,
		_w3815_
	);
	LUT2 #(
		.INIT('h8)
	) name2307 (
		RESET_pad,
		\WX4698_reg/NET0131 ,
		_w3816_
	);
	LUT2 #(
		.INIT('h8)
	) name2308 (
		RESET_pad,
		\WX8591_reg/NET0131 ,
		_w3817_
	);
	LUT2 #(
		.INIT('h8)
	) name2309 (
		RESET_pad,
		\WX3239_reg/NET0131 ,
		_w3818_
	);
	LUT2 #(
		.INIT('h8)
	) name2310 (
		RESET_pad,
		\WX4704_reg/NET0131 ,
		_w3819_
	);
	LUT2 #(
		.INIT('h8)
	) name2311 (
		RESET_pad,
		\WX8583_reg/NET0131 ,
		_w3820_
	);
	LUT2 #(
		.INIT('h8)
	) name2312 (
		RESET_pad,
		\WX11029_reg/NET0131 ,
		_w3821_
	);
	LUT2 #(
		.INIT('h8)
	) name2313 (
		RESET_pad,
		\WX4712_reg/NET0131 ,
		_w3822_
	);
	LUT2 #(
		.INIT('h8)
	) name2314 (
		RESET_pad,
		\WX743_reg/NET0131 ,
		_w3823_
	);
	LUT2 #(
		.INIT('h8)
	) name2315 (
		RESET_pad,
		\WX8565_reg/NET0131 ,
		_w3824_
	);
	LUT2 #(
		.INIT('h8)
	) name2316 (
		RESET_pad,
		\WX8579_reg/NET0131 ,
		_w3825_
	);
	LUT2 #(
		.INIT('h8)
	) name2317 (
		RESET_pad,
		\WX3383_reg/NET0131 ,
		_w3826_
	);
	LUT2 #(
		.INIT('h8)
	) name2318 (
		RESET_pad,
		\WX8559_reg/NET0131 ,
		_w3827_
	);
	LUT2 #(
		.INIT('h8)
	) name2319 (
		RESET_pad,
		\WX2104_reg/NET0131 ,
		_w3828_
	);
	LUT2 #(
		.INIT('h8)
	) name2320 (
		RESET_pad,
		\WX4678_reg/NET0131 ,
		_w3829_
	);
	LUT2 #(
		.INIT('h8)
	) name2321 (
		RESET_pad,
		\WX689_reg/NET0131 ,
		_w3830_
	);
	LUT2 #(
		.INIT('h8)
	) name2322 (
		RESET_pad,
		\WX3233_reg/NET0131 ,
		_w3831_
	);
	LUT2 #(
		.INIT('h8)
	) name2323 (
		RESET_pad,
		\WX3393_reg/NET0131 ,
		_w3832_
	);
	LUT2 #(
		.INIT('h8)
	) name2324 (
		RESET_pad,
		\WX8455_reg/NET0131 ,
		_w3833_
	);
	LUT2 #(
		.INIT('h8)
	) name2325 (
		RESET_pad,
		\WX3235_reg/NET0131 ,
		_w3834_
	);
	LUT2 #(
		.INIT('h8)
	) name2326 (
		RESET_pad,
		\WX739_reg/NET0131 ,
		_w3835_
	);
	LUT2 #(
		.INIT('h8)
	) name2327 (
		RESET_pad,
		\WX8567_reg/NET0131 ,
		_w3836_
	);
	LUT2 #(
		.INIT('h8)
	) name2328 (
		RESET_pad,
		\WX8573_reg/NET0131 ,
		_w3837_
	);
	LUT2 #(
		.INIT('h8)
	) name2329 (
		RESET_pad,
		\WX3391_reg/NET0131 ,
		_w3838_
	);
	LUT2 #(
		.INIT('h8)
	) name2330 (
		RESET_pad,
		\WX10995_reg/NET0131 ,
		_w3839_
	);
	LUT2 #(
		.INIT('h8)
	) name2331 (
		RESET_pad,
		\WX8571_reg/NET0131 ,
		_w3840_
	);
	LUT2 #(
		.INIT('h8)
	) name2332 (
		RESET_pad,
		\WX2108_reg/NET0131 ,
		_w3841_
	);
	LUT2 #(
		.INIT('h8)
	) name2333 (
		RESET_pad,
		\WX2008_reg/NET0131 ,
		_w3842_
	);
	LUT2 #(
		.INIT('h8)
	) name2334 (
		RESET_pad,
		\WX7242_reg/NET0131 ,
		_w3843_
	);
	LUT2 #(
		.INIT('h8)
	) name2335 (
		RESET_pad,
		\WX11015_reg/NET0131 ,
		_w3844_
	);
	LUT2 #(
		.INIT('h8)
	) name2336 (
		RESET_pad,
		\WX9864_reg/NET0131 ,
		_w3845_
	);
	LUT2 #(
		.INIT('h8)
	) name2337 (
		RESET_pad,
		\WX3385_reg/NET0131 ,
		_w3846_
	);
	LUT2 #(
		.INIT('h8)
	) name2338 (
		RESET_pad,
		\WX4710_reg/NET0131 ,
		_w3847_
	);
	LUT2 #(
		.INIT('h8)
	) name2339 (
		RESET_pad,
		\WX779_reg/NET0131 ,
		_w3848_
	);
	LUT2 #(
		.INIT('h8)
	) name2340 (
		RESET_pad,
		\WX753_reg/NET0131 ,
		_w3849_
	);
	LUT2 #(
		.INIT('h8)
	) name2341 (
		RESET_pad,
		\WX733_reg/NET0131 ,
		_w3850_
	);
	LUT2 #(
		.INIT('h8)
	) name2342 (
		RESET_pad,
		\WX2012_reg/NET0131 ,
		_w3851_
	);
	LUT2 #(
		.INIT('h8)
	) name2343 (
		RESET_pad,
		\WX2086_reg/NET0131 ,
		_w3852_
	);
	LUT2 #(
		.INIT('h8)
	) name2344 (
		RESET_pad,
		\WX4680_reg/NET0131 ,
		_w3853_
	);
	LUT2 #(
		.INIT('h8)
	) name2345 (
		RESET_pad,
		\WX4696_reg/NET0131 ,
		_w3854_
	);
	LUT2 #(
		.INIT('h8)
	) name2346 (
		RESET_pad,
		\WX8561_reg/NET0131 ,
		_w3855_
	);
	LUT2 #(
		.INIT('h8)
	) name2347 (
		RESET_pad,
		\WX11077_reg/NET0131 ,
		_w3856_
	);
	LUT2 #(
		.INIT('h8)
	) name2348 (
		RESET_pad,
		\WX2106_reg/NET0131 ,
		_w3857_
	);
	LUT2 #(
		.INIT('h8)
	) name2349 (
		RESET_pad,
		\WX4686_reg/NET0131 ,
		_w3858_
	);
	LUT2 #(
		.INIT('h8)
	) name2350 (
		RESET_pad,
		\WX3335_reg/NET0131 ,
		_w3859_
	);
	LUT2 #(
		.INIT('h8)
	) name2351 (
		RESET_pad,
		\WX4666_reg/NET0131 ,
		_w3860_
	);
	LUT2 #(
		.INIT('h8)
	) name2352 (
		RESET_pad,
		\WX9830_reg/NET0131 ,
		_w3861_
	);
	LUT2 #(
		.INIT('h8)
	) name2353 (
		RESET_pad,
		\WX9788_reg/NET0131 ,
		_w3862_
	);
	LUT2 #(
		.INIT('h8)
	) name2354 (
		RESET_pad,
		\WX4674_reg/NET0131 ,
		_w3863_
	);
	LUT2 #(
		.INIT('h8)
	) name2355 (
		RESET_pad,
		\WX9838_reg/NET0131 ,
		_w3864_
	);
	LUT2 #(
		.INIT('h8)
	) name2356 (
		RESET_pad,
		\WX4670_reg/NET0131 ,
		_w3865_
	);
	LUT2 #(
		.INIT('h8)
	) name2357 (
		RESET_pad,
		\WX3253_reg/NET0131 ,
		_w3866_
	);
	LUT2 #(
		.INIT('h8)
	) name2358 (
		RESET_pad,
		\WX4664_reg/NET0131 ,
		_w3867_
	);
	LUT2 #(
		.INIT('h8)
	) name2359 (
		RESET_pad,
		\WX7296_reg/NET0131 ,
		_w3868_
	);
	LUT2 #(
		.INIT('h8)
	) name2360 (
		RESET_pad,
		\WX4660_reg/NET0131 ,
		_w3869_
	);
	LUT2 #(
		.INIT('h8)
	) name2361 (
		RESET_pad,
		\WX9696_reg/NET0131 ,
		_w3870_
	);
	LUT2 #(
		.INIT('h8)
	) name2362 (
		RESET_pad,
		\WX4566_reg/NET0131 ,
		_w3871_
	);
	LUT2 #(
		.INIT('h8)
	) name2363 (
		RESET_pad,
		\WX11001_reg/NET0131 ,
		_w3872_
	);
	LUT2 #(
		.INIT('h8)
	) name2364 (
		RESET_pad,
		\WX9812_reg/NET0131 ,
		_w3873_
	);
	LUT2 #(
		.INIT('h8)
	) name2365 (
		RESET_pad,
		\WX4620_reg/NET0131 ,
		_w3874_
	);
	LUT2 #(
		.INIT('h8)
	) name2366 (
		RESET_pad,
		\WX3407_reg/NET0131 ,
		_w3875_
	);
	LUT2 #(
		.INIT('h8)
	) name2367 (
		RESET_pad,
		\WX821_reg/NET0131 ,
		_w3876_
	);
	LUT2 #(
		.INIT('h8)
	) name2368 (
		RESET_pad,
		\WX8531_reg/NET0131 ,
		_w3877_
	);
	LUT2 #(
		.INIT('h8)
	) name2369 (
		RESET_pad,
		\WX2102_reg/NET0131 ,
		_w3878_
	);
	LUT2 #(
		.INIT('h8)
	) name2370 (
		RESET_pad,
		\WX649_reg/NET0131 ,
		_w3879_
	);
	LUT2 #(
		.INIT('h8)
	) name2371 (
		RESET_pad,
		\WX829_reg/NET0131 ,
		_w3880_
	);
	LUT2 #(
		.INIT('h8)
	) name2372 (
		RESET_pad,
		\WX8555_reg/NET0131 ,
		_w3881_
	);
	LUT2 #(
		.INIT('h8)
	) name2373 (
		RESET_pad,
		\WX3295_reg/NET0131 ,
		_w3882_
	);
	LUT2 #(
		.INIT('h8)
	) name2374 (
		RESET_pad,
		\WX2100_reg/NET0131 ,
		_w3883_
	);
	LUT2 #(
		.INIT('h8)
	) name2375 (
		RESET_pad,
		\WX825_reg/NET0131 ,
		_w3884_
	);
	LUT2 #(
		.INIT('h8)
	) name2376 (
		RESET_pad,
		\WX11017_reg/NET0131 ,
		_w3885_
	);
	LUT2 #(
		.INIT('h8)
	) name2377 (
		RESET_pad,
		\WX5951_reg/NET0131 ,
		_w3886_
	);
	LUT2 #(
		.INIT('h8)
	) name2378 (
		RESET_pad,
		\WX2098_reg/NET0131 ,
		_w3887_
	);
	LUT2 #(
		.INIT('h8)
	) name2379 (
		RESET_pad,
		\WX3297_reg/NET0131 ,
		_w3888_
	);
	LUT2 #(
		.INIT('h8)
	) name2380 (
		RESET_pad,
		\WX5849_reg/NET0131 ,
		_w3889_
	);
	LUT2 #(
		.INIT('h8)
	) name2381 (
		RESET_pad,
		\WX8553_reg/NET0131 ,
		_w3890_
	);
	LUT2 #(
		.INIT('h8)
	) name2382 (
		RESET_pad,
		\WX2016_reg/NET0131 ,
		_w3891_
	);
	LUT2 #(
		.INIT('h8)
	) name2383 (
		RESET_pad,
		\WX11063_reg/NET0131 ,
		_w3892_
	);
	LUT2 #(
		.INIT('h8)
	) name2384 (
		RESET_pad,
		\WX9700_reg/NET0131 ,
		_w3893_
	);
	LUT2 #(
		.INIT('h8)
	) name2385 (
		RESET_pad,
		\WX8463_reg/NET0131 ,
		_w3894_
	);
	LUT2 #(
		.INIT('h8)
	) name2386 (
		RESET_pad,
		\WX2096_reg/NET0131 ,
		_w3895_
	);
	LUT2 #(
		.INIT('h8)
	) name2387 (
		RESET_pad,
		\WX3331_reg/NET0131 ,
		_w3896_
	);
	LUT2 #(
		.INIT('h8)
	) name2388 (
		RESET_pad,
		\WX3299_reg/NET0131 ,
		_w3897_
	);
	LUT2 #(
		.INIT('h8)
	) name2389 (
		RESET_pad,
		\WX8549_reg/NET0131 ,
		_w3898_
	);
	LUT2 #(
		.INIT('h8)
	) name2390 (
		RESET_pad,
		\WX795_reg/NET0131 ,
		_w3899_
	);
	LUT2 #(
		.INIT('h8)
	) name2391 (
		RESET_pad,
		\WX3375_reg/NET0131 ,
		_w3900_
	);
	LUT2 #(
		.INIT('h8)
	) name2392 (
		RESET_pad,
		\WX5859_reg/NET0131 ,
		_w3901_
	);
	LUT2 #(
		.INIT('h8)
	) name2393 (
		RESET_pad,
		\WX4548_reg/NET0131 ,
		_w3902_
	);
	LUT2 #(
		.INIT('h8)
	) name2394 (
		RESET_pad,
		\WX3419_reg/NET0131 ,
		_w3903_
	);
	LUT2 #(
		.INIT('h8)
	) name2395 (
		RESET_pad,
		\WX8545_reg/NET0131 ,
		_w3904_
	);
	LUT2 #(
		.INIT('h8)
	) name2396 (
		RESET_pad,
		\WX4622_reg/NET0131 ,
		_w3905_
	);
	LUT2 #(
		.INIT('h8)
	) name2397 (
		RESET_pad,
		\WX8539_reg/NET0131 ,
		_w3906_
	);
	LUT2 #(
		.INIT('h8)
	) name2398 (
		RESET_pad,
		\WX2094_reg/NET0131 ,
		_w3907_
	);
	LUT2 #(
		.INIT('h8)
	) name2399 (
		RESET_pad,
		\WX2048_reg/NET0131 ,
		_w3908_
	);
	LUT2 #(
		.INIT('h8)
	) name2400 (
		RESET_pad,
		\WX723_reg/NET0131 ,
		_w3909_
	);
	LUT2 #(
		.INIT('h8)
	) name2401 (
		RESET_pad,
		\WX4600_reg/NET0131 ,
		_w3910_
	);
	LUT2 #(
		.INIT('h8)
	) name2402 (
		RESET_pad,
		\WX4602_reg/NET0131 ,
		_w3911_
	);
	LUT2 #(
		.INIT('h8)
	) name2403 (
		RESET_pad,
		\WX8405_reg/NET0131 ,
		_w3912_
	);
	LUT2 #(
		.INIT('h8)
	) name2404 (
		RESET_pad,
		\WX4650_reg/NET0131 ,
		_w3913_
	);
	LUT2 #(
		.INIT('h8)
	) name2405 (
		RESET_pad,
		\WX8543_reg/NET0131 ,
		_w3914_
	);
	LUT2 #(
		.INIT('h8)
	) name2406 (
		RESET_pad,
		\WX10997_reg/NET0131 ,
		_w3915_
	);
	LUT2 #(
		.INIT('h8)
	) name2407 (
		RESET_pad,
		\WX7282_reg/NET0131 ,
		_w3916_
	);
	LUT2 #(
		.INIT('h8)
	) name2408 (
		RESET_pad,
		\WX9884_reg/NET0131 ,
		_w3917_
	);
	LUT2 #(
		.INIT('h8)
	) name2409 (
		RESET_pad,
		\WX5899_reg/NET0131 ,
		_w3918_
	);
	LUT2 #(
		.INIT('h8)
	) name2410 (
		RESET_pad,
		\WX3369_reg/NET0131 ,
		_w3919_
	);
	LUT2 #(
		.INIT('h8)
	) name2411 (
		RESET_pad,
		\WX4616_reg/NET0131 ,
		_w3920_
	);
	LUT2 #(
		.INIT('h8)
	) name2412 (
		RESET_pad,
		\WX8457_reg/NET0131 ,
		_w3921_
	);
	LUT2 #(
		.INIT('h8)
	) name2413 (
		RESET_pad,
		\WX5855_reg/NET0131 ,
		_w3922_
	);
	LUT2 #(
		.INIT('h8)
	) name2414 (
		RESET_pad,
		\WX8435_reg/NET0131 ,
		_w3923_
	);
	LUT2 #(
		.INIT('h8)
	) name2415 (
		RESET_pad,
		\WX759_reg/NET0131 ,
		_w3924_
	);
	LUT2 #(
		.INIT('h8)
	) name2416 (
		RESET_pad,
		\WX8537_reg/NET0131 ,
		_w3925_
	);
	LUT2 #(
		.INIT('h8)
	) name2417 (
		RESET_pad,
		\WX9854_reg/NET0131 ,
		_w3926_
	);
	LUT2 #(
		.INIT('h8)
	) name2418 (
		RESET_pad,
		\WX10999_reg/NET0131 ,
		_w3927_
	);
	LUT2 #(
		.INIT('h8)
	) name2419 (
		RESET_pad,
		\WX7250_reg/NET0131 ,
		_w3928_
	);
	LUT2 #(
		.INIT('h8)
	) name2420 (
		RESET_pad,
		\WX1978_reg/NET0131 ,
		_w3929_
	);
	LUT2 #(
		.INIT('h8)
	) name2421 (
		RESET_pad,
		\WX651_reg/NET0131 ,
		_w3930_
	);
	LUT2 #(
		.INIT('h8)
	) name2422 (
		RESET_pad,
		\WX3387_reg/NET0131 ,
		_w3931_
	);
	LUT2 #(
		.INIT('h8)
	) name2423 (
		RESET_pad,
		\WX681_reg/NET0131 ,
		_w3932_
	);
	LUT2 #(
		.INIT('h8)
	) name2424 (
		RESET_pad,
		\WX8535_reg/NET0131 ,
		_w3933_
	);
	LUT2 #(
		.INIT('h8)
	) name2425 (
		RESET_pad,
		\WX7212_reg/NET0131 ,
		_w3934_
	);
	LUT2 #(
		.INIT('h8)
	) name2426 (
		RESET_pad,
		\WX5981_reg/NET0131 ,
		_w3935_
	);
	LUT2 #(
		.INIT('h8)
	) name2427 (
		RESET_pad,
		\WX4586_reg/NET0131 ,
		_w3936_
	);
	LUT2 #(
		.INIT('h8)
	) name2428 (
		RESET_pad,
		\WX4656_reg/NET0131 ,
		_w3937_
	);
	LUT2 #(
		.INIT('h8)
	) name2429 (
		RESET_pad,
		\WX3333_reg/NET0131 ,
		_w3938_
	);
	LUT2 #(
		.INIT('h8)
	) name2430 (
		RESET_pad,
		\WX9826_reg/NET0131 ,
		_w3939_
	);
	LUT2 #(
		.INIT('h8)
	) name2431 (
		RESET_pad,
		\WX2092_reg/NET0131 ,
		_w3940_
	);
	LUT2 #(
		.INIT('h8)
	) name2432 (
		RESET_pad,
		\WX4624_reg/NET0131 ,
		_w3941_
	);
	LUT2 #(
		.INIT('h8)
	) name2433 (
		RESET_pad,
		\WX7136_reg/NET0131 ,
		_w3942_
	);
	LUT2 #(
		.INIT('h8)
	) name2434 (
		RESET_pad,
		\WX7268_reg/NET0131 ,
		_w3943_
	);
	LUT2 #(
		.INIT('h8)
	) name2435 (
		RESET_pad,
		\WX4642_reg/NET0131 ,
		_w3944_
	);
	LUT2 #(
		.INIT('h8)
	) name2436 (
		RESET_pad,
		\WX8409_reg/NET0131 ,
		_w3945_
	);
	LUT2 #(
		.INIT('h8)
	) name2437 (
		RESET_pad,
		\WX4618_reg/NET0131 ,
		_w3946_
	);
	LUT2 #(
		.INIT('h8)
	) name2438 (
		RESET_pad,
		\WX4612_reg/NET0131 ,
		_w3947_
	);
	LUT2 #(
		.INIT('h8)
	) name2439 (
		RESET_pad,
		\WX7292_reg/NET0131 ,
		_w3948_
	);
	LUT2 #(
		.INIT('h8)
	) name2440 (
		RESET_pad,
		\WX3231_reg/NET0131 ,
		_w3949_
	);
	LUT2 #(
		.INIT('h8)
	) name2441 (
		RESET_pad,
		\WX8489_reg/NET0131 ,
		_w3950_
	);
	LUT2 #(
		.INIT('h8)
	) name2442 (
		RESET_pad,
		\WX3305_reg/NET0131 ,
		_w3951_
	);
	LUT2 #(
		.INIT('h8)
	) name2443 (
		RESET_pad,
		\WX8525_reg/NET0131 ,
		_w3952_
	);
	LUT2 #(
		.INIT('h8)
	) name2444 (
		RESET_pad,
		\WX11159_reg/NET0131 ,
		_w3953_
	);
	LUT2 #(
		.INIT('h8)
	) name2445 (
		RESET_pad,
		\WX3367_reg/NET0131 ,
		_w3954_
	);
	LUT2 #(
		.INIT('h8)
	) name2446 (
		RESET_pad,
		\WX11061_reg/NET0131 ,
		_w3955_
	);
	LUT2 #(
		.INIT('h8)
	) name2447 (
		RESET_pad,
		\WX8569_reg/NET0131 ,
		_w3956_
	);
	LUT2 #(
		.INIT('h8)
	) name2448 (
		RESET_pad,
		\WX11125_reg/NET0131 ,
		_w3957_
	);
	LUT2 #(
		.INIT('h8)
	) name2449 (
		RESET_pad,
		\WX809_reg/NET0131 ,
		_w3958_
	);
	LUT2 #(
		.INIT('h8)
	) name2450 (
		RESET_pad,
		\WX683_reg/NET0131 ,
		_w3959_
	);
	LUT2 #(
		.INIT('h8)
	) name2451 (
		RESET_pad,
		\WX8413_reg/NET0131 ,
		_w3960_
	);
	LUT2 #(
		.INIT('h8)
	) name2452 (
		RESET_pad,
		\WX2062_reg/NET0131 ,
		_w3961_
	);
	LUT2 #(
		.INIT('h8)
	) name2453 (
		RESET_pad,
		\WX9758_reg/NET0131 ,
		_w3962_
	);
	LUT2 #(
		.INIT('h8)
	) name2454 (
		RESET_pad,
		\WX3397_reg/NET0131 ,
		_w3963_
	);
	LUT2 #(
		.INIT('h8)
	) name2455 (
		RESET_pad,
		\WX7300_reg/NET0131 ,
		_w3964_
	);
	LUT2 #(
		.INIT('h8)
	) name2456 (
		RESET_pad,
		\WX6003_reg/NET0131 ,
		_w3965_
	);
	LUT2 #(
		.INIT('h8)
	) name2457 (
		RESET_pad,
		\WX4646_reg/NET0131 ,
		_w3966_
	);
	LUT2 #(
		.INIT('h8)
	) name2458 (
		RESET_pad,
		\WX9880_reg/NET0131 ,
		_w3967_
	);
	LUT2 #(
		.INIT('h8)
	) name2459 (
		RESET_pad,
		\WX7258_reg/NET0131 ,
		_w3968_
	);
	LUT2 #(
		.INIT('h8)
	) name2460 (
		RESET_pad,
		\WX8593_reg/NET0131 ,
		_w3969_
	);
	LUT2 #(
		.INIT('h8)
	) name2461 (
		RESET_pad,
		\WX11057_reg/NET0131 ,
		_w3970_
	);
	LUT2 #(
		.INIT('h8)
	) name2462 (
		RESET_pad,
		\WX675_reg/NET0131 ,
		_w3971_
	);
	LUT2 #(
		.INIT('h8)
	) name2463 (
		RESET_pad,
		\WX3371_reg/NET0131 ,
		_w3972_
	);
	LUT2 #(
		.INIT('h8)
	) name2464 (
		RESET_pad,
		\WX783_reg/NET0131 ,
		_w3973_
	);
	LUT2 #(
		.INIT('h8)
	) name2465 (
		RESET_pad,
		\WX8411_reg/NET0131 ,
		_w3974_
	);
	LUT2 #(
		.INIT('h8)
	) name2466 (
		RESET_pad,
		\WX9836_reg/NET0131 ,
		_w3975_
	);
	LUT2 #(
		.INIT('h8)
	) name2467 (
		RESET_pad,
		\WX11055_reg/NET0131 ,
		_w3976_
	);
	LUT2 #(
		.INIT('h8)
	) name2468 (
		RESET_pad,
		\WX8467_reg/NET0131 ,
		_w3977_
	);
	LUT2 #(
		.INIT('h8)
	) name2469 (
		RESET_pad,
		\WX817_reg/NET0131 ,
		_w3978_
	);
	LUT2 #(
		.INIT('h8)
	) name2470 (
		RESET_pad,
		\WX9870_reg/NET0131 ,
		_w3979_
	);
	LUT2 #(
		.INIT('h8)
	) name2471 (
		RESET_pad,
		\WX7262_reg/NET0131 ,
		_w3980_
	);
	LUT2 #(
		.INIT('h8)
	) name2472 (
		RESET_pad,
		\WX7264_reg/NET0131 ,
		_w3981_
	);
	LUT2 #(
		.INIT('h8)
	) name2473 (
		RESET_pad,
		\WX4604_reg/NET0131 ,
		_w3982_
	);
	LUT2 #(
		.INIT('h8)
	) name2474 (
		RESET_pad,
		\WX9804_reg/NET0131 ,
		_w3983_
	);
	LUT2 #(
		.INIT('h8)
	) name2475 (
		RESET_pad,
		\WX8429_reg/NET0131 ,
		_w3984_
	);
	LUT2 #(
		.INIT('h8)
	) name2476 (
		RESET_pad,
		\WX815_reg/NET0131 ,
		_w3985_
	);
	LUT2 #(
		.INIT('h8)
	) name2477 (
		RESET_pad,
		\WX5877_reg/NET0131 ,
		_w3986_
	);
	LUT2 #(
		.INIT('h8)
	) name2478 (
		RESET_pad,
		\WX6001_reg/NET0131 ,
		_w3987_
	);
	LUT2 #(
		.INIT('h8)
	) name2479 (
		RESET_pad,
		\WX8521_reg/NET0131 ,
		_w3988_
	);
	LUT2 #(
		.INIT('h8)
	) name2480 (
		RESET_pad,
		\WX7270_reg/NET0131 ,
		_w3989_
	);
	LUT2 #(
		.INIT('h8)
	) name2481 (
		RESET_pad,
		\WX677_reg/NET0131 ,
		_w3990_
	);
	LUT2 #(
		.INIT('h8)
	) name2482 (
		RESET_pad,
		\WX5989_reg/NET0131 ,
		_w3991_
	);
	LUT2 #(
		.INIT('h8)
	) name2483 (
		RESET_pad,
		\WX5993_reg/NET0131 ,
		_w3992_
	);
	LUT2 #(
		.INIT('h8)
	) name2484 (
		RESET_pad,
		\WX3303_reg/NET0131 ,
		_w3993_
	);
	LUT2 #(
		.INIT('h8)
	) name2485 (
		RESET_pad,
		\WX7142_reg/NET0131 ,
		_w3994_
	);
	LUT2 #(
		.INIT('h8)
	) name2486 (
		RESET_pad,
		\WX793_reg/NET0131 ,
		_w3995_
	);
	LUT2 #(
		.INIT('h8)
	) name2487 (
		RESET_pad,
		\WX9756_reg/NET0131 ,
		_w3996_
	);
	LUT2 #(
		.INIT('h8)
	) name2488 (
		RESET_pad,
		\WX7260_reg/NET0131 ,
		_w3997_
	);
	LUT2 #(
		.INIT('h8)
	) name2489 (
		RESET_pad,
		\WX5903_reg/NET0131 ,
		_w3998_
	);
	LUT2 #(
		.INIT('h8)
	) name2490 (
		RESET_pad,
		\WX11065_reg/NET0131 ,
		_w3999_
	);
	LUT2 #(
		.INIT('h8)
	) name2491 (
		RESET_pad,
		\WX4534_reg/NET0131 ,
		_w4000_
	);
	LUT2 #(
		.INIT('h8)
	) name2492 (
		RESET_pad,
		\WX4546_reg/NET0131 ,
		_w4001_
	);
	LUT2 #(
		.INIT('h8)
	) name2493 (
		RESET_pad,
		\WX2074_reg/NET0131 ,
		_w4002_
	);
	LUT2 #(
		.INIT('h8)
	) name2494 (
		RESET_pad,
		\WX8483_reg/NET0131 ,
		_w4003_
	);
	LUT2 #(
		.INIT('h8)
	) name2495 (
		RESET_pad,
		\WX3307_reg/NET0131 ,
		_w4004_
	);
	LUT2 #(
		.INIT('h8)
	) name2496 (
		RESET_pad,
		\WX9866_reg/NET0131 ,
		_w4005_
	);
	LUT2 #(
		.INIT('h8)
	) name2497 (
		RESET_pad,
		\WX4610_reg/NET0131 ,
		_w4006_
	);
	LUT2 #(
		.INIT('h8)
	) name2498 (
		RESET_pad,
		\WX4582_reg/NET0131 ,
		_w4007_
	);
	LUT2 #(
		.INIT('h8)
	) name2499 (
		RESET_pad,
		\WX5987_reg/NET0131 ,
		_w4008_
	);
	LUT2 #(
		.INIT('h8)
	) name2500 (
		RESET_pad,
		\WX11051_reg/NET0131 ,
		_w4009_
	);
	LUT2 #(
		.INIT('h8)
	) name2501 (
		RESET_pad,
		\WX4640_reg/NET0131 ,
		_w4010_
	);
	LUT2 #(
		.INIT('h8)
	) name2502 (
		RESET_pad,
		\WX655_reg/NET0131 ,
		_w4011_
	);
	LUT2 #(
		.INIT('h8)
	) name2503 (
		RESET_pad,
		\WX4596_reg/NET0131 ,
		_w4012_
	);
	LUT2 #(
		.INIT('h8)
	) name2504 (
		RESET_pad,
		\WX673_reg/NET0131 ,
		_w4013_
	);
	LUT2 #(
		.INIT('h8)
	) name2505 (
		RESET_pad,
		\WX4592_reg/NET0131 ,
		_w4014_
	);
	LUT2 #(
		.INIT('h8)
	) name2506 (
		RESET_pad,
		\WX7298_reg/NET0131 ,
		_w4015_
	);
	LUT2 #(
		.INIT('h8)
	) name2507 (
		RESET_pad,
		\WX2078_reg/NET0131 ,
		_w4016_
	);
	LUT2 #(
		.INIT('h8)
	) name2508 (
		RESET_pad,
		\WX2038_reg/NET0131 ,
		_w4017_
	);
	LUT2 #(
		.INIT('h8)
	) name2509 (
		RESET_pad,
		\WX11003_reg/NET0131 ,
		_w4018_
	);
	LUT2 #(
		.INIT('h8)
	) name2510 (
		RESET_pad,
		\WX5881_reg/NET0131 ,
		_w4019_
	);
	LUT2 #(
		.INIT('h8)
	) name2511 (
		RESET_pad,
		\WX4644_reg/NET0131 ,
		_w4020_
	);
	LUT2 #(
		.INIT('h8)
	) name2512 (
		RESET_pad,
		\WX2120_reg/NET0131 ,
		_w4021_
	);
	LUT2 #(
		.INIT('h8)
	) name2513 (
		RESET_pad,
		\WX4654_reg/NET0131 ,
		_w4022_
	);
	LUT2 #(
		.INIT('h8)
	) name2514 (
		RESET_pad,
		\WX3353_reg/NET0131 ,
		_w4023_
	);
	LUT2 #(
		.INIT('h8)
	) name2515 (
		RESET_pad,
		\WX5983_reg/NET0131 ,
		_w4024_
	);
	LUT2 #(
		.INIT('h8)
	) name2516 (
		RESET_pad,
		\WX4572_reg/NET0131 ,
		_w4025_
	);
	LUT2 #(
		.INIT('h8)
	) name2517 (
		RESET_pad,
		\WX8427_reg/NET0131 ,
		_w4026_
	);
	LUT2 #(
		.INIT('h8)
	) name2518 (
		RESET_pad,
		\WX4684_reg/NET0131 ,
		_w4027_
	);
	LUT2 #(
		.INIT('h8)
	) name2519 (
		RESET_pad,
		\WX4694_reg/NET0131 ,
		_w4028_
	);
	LUT2 #(
		.INIT('h8)
	) name2520 (
		RESET_pad,
		\WX833_reg/NET0131 ,
		_w4029_
	);
	LUT2 #(
		.INIT('h8)
	) name2521 (
		RESET_pad,
		\WX9886_reg/NET0131 ,
		_w4030_
	);
	LUT2 #(
		.INIT('h8)
	) name2522 (
		RESET_pad,
		\WX4552_reg/NET0131 ,
		_w4031_
	);
	LUT2 #(
		.INIT('h8)
	) name2523 (
		RESET_pad,
		\WX4606_reg/NET0131 ,
		_w4032_
	);
	LUT2 #(
		.INIT('h8)
	) name2524 (
		RESET_pad,
		\WX4536_reg/NET0131 ,
		_w4033_
	);
	LUT2 #(
		.INIT('h8)
	) name2525 (
		RESET_pad,
		\WX7140_reg/NET0131 ,
		_w4034_
	);
	LUT2 #(
		.INIT('h8)
	) name2526 (
		RESET_pad,
		\WX5975_reg/NET0131 ,
		_w4035_
	);
	LUT2 #(
		.INIT('h8)
	) name2527 (
		RESET_pad,
		\WX2110_reg/NET0131 ,
		_w4036_
	);
	LUT2 #(
		.INIT('h8)
	) name2528 (
		RESET_pad,
		\WX7274_reg/NET0131 ,
		_w4037_
	);
	LUT2 #(
		.INIT('h8)
	) name2529 (
		RESET_pad,
		\WX5977_reg/NET0131 ,
		_w4038_
	);
	LUT2 #(
		.INIT('h8)
	) name2530 (
		RESET_pad,
		\WX3417_reg/NET0131 ,
		_w4039_
	);
	LUT2 #(
		.INIT('h8)
	) name2531 (
		RESET_pad,
		\WX8507_reg/NET0131 ,
		_w4040_
	);
	LUT2 #(
		.INIT('h8)
	) name2532 (
		RESET_pad,
		\WX9720_reg/NET0131 ,
		_w4041_
	);
	LUT2 #(
		.INIT('h8)
	) name2533 (
		RESET_pad,
		\WX5971_reg/NET0131 ,
		_w4042_
	);
	LUT2 #(
		.INIT('h8)
	) name2534 (
		RESET_pad,
		\WX5967_reg/NET0131 ,
		_w4043_
	);
	LUT2 #(
		.INIT('h8)
	) name2535 (
		RESET_pad,
		\WX7146_reg/NET0131 ,
		_w4044_
	);
	LUT2 #(
		.INIT('h8)
	) name2536 (
		RESET_pad,
		\WX8541_reg/NET0131 ,
		_w4045_
	);
	LUT2 #(
		.INIT('h8)
	) name2537 (
		RESET_pad,
		\WX5969_reg/NET0131 ,
		_w4046_
	);
	LUT2 #(
		.INIT('h8)
	) name2538 (
		RESET_pad,
		\WX3373_reg/NET0131 ,
		_w4047_
	);
	LUT2 #(
		.INIT('h8)
	) name2539 (
		RESET_pad,
		\WX5963_reg/NET0131 ,
		_w4048_
	);
	LUT2 #(
		.INIT('h8)
	) name2540 (
		RESET_pad,
		\WX8513_reg/NET0131 ,
		_w4049_
	);
	LUT2 #(
		.INIT('h8)
	) name2541 (
		RESET_pad,
		\WX8509_reg/NET0131 ,
		_w4050_
	);
	LUT2 #(
		.INIT('h8)
	) name2542 (
		RESET_pad,
		\WX8433_reg/NET0131 ,
		_w4051_
	);
	LUT2 #(
		.INIT('h8)
	) name2543 (
		RESET_pad,
		\WX11047_reg/NET0131 ,
		_w4052_
	);
	LUT2 #(
		.INIT('h8)
	) name2544 (
		RESET_pad,
		\WX1942_reg/NET0131 ,
		_w4053_
	);
	LUT2 #(
		.INIT('h8)
	) name2545 (
		RESET_pad,
		\WX5961_reg/NET0131 ,
		_w4054_
	);
	LUT2 #(
		.INIT('h8)
	) name2546 (
		RESET_pad,
		\WX8511_reg/NET0131 ,
		_w4055_
	);
	LUT2 #(
		.INIT('h8)
	) name2547 (
		RESET_pad,
		\WX8431_reg/NET0131 ,
		_w4056_
	);
	LUT2 #(
		.INIT('h8)
	) name2548 (
		RESET_pad,
		\WX7286_reg/NET0131 ,
		_w4057_
	);
	LUT2 #(
		.INIT('h8)
	) name2549 (
		RESET_pad,
		\WX7288_reg/NET0131 ,
		_w4058_
	);
	LUT2 #(
		.INIT('h8)
	) name2550 (
		RESET_pad,
		\WX3343_reg/NET0131 ,
		_w4059_
	);
	LUT2 #(
		.INIT('h8)
	) name2551 (
		RESET_pad,
		\WX7112_reg/NET0131 ,
		_w4060_
	);
	LUT2 #(
		.INIT('h8)
	) name2552 (
		RESET_pad,
		\WX9766_reg/NET0131 ,
		_w4061_
	);
	LUT2 #(
		.INIT('h8)
	) name2553 (
		RESET_pad,
		\WX3315_reg/NET0131 ,
		_w4062_
	);
	LUT2 #(
		.INIT('h8)
	) name2554 (
		RESET_pad,
		\WX2070_reg/NET0131 ,
		_w4063_
	);
	LUT2 #(
		.INIT('h8)
	) name2555 (
		RESET_pad,
		\WX11091_reg/NET0131 ,
		_w4064_
	);
	LUT2 #(
		.INIT('h8)
	) name2556 (
		RESET_pad,
		\WX3377_reg/NET0131 ,
		_w4065_
	);
	LUT2 #(
		.INIT('h8)
	) name2557 (
		RESET_pad,
		\WX5943_reg/NET0131 ,
		_w4066_
	);
	LUT2 #(
		.INIT('h8)
	) name2558 (
		RESET_pad,
		\WX8479_reg/NET0131 ,
		_w4067_
	);
	LUT2 #(
		.INIT('h8)
	) name2559 (
		RESET_pad,
		\WX1948_reg/NET0131 ,
		_w4068_
	);
	LUT2 #(
		.INIT('h8)
	) name2560 (
		RESET_pad,
		\WX747_reg/NET0131 ,
		_w4069_
	);
	LUT2 #(
		.INIT('h8)
	) name2561 (
		RESET_pad,
		\WX8439_reg/NET0131 ,
		_w4070_
	);
	LUT2 #(
		.INIT('h8)
	) name2562 (
		RESET_pad,
		\WX9738_reg/NET0131 ,
		_w4071_
	);
	LUT2 #(
		.INIT('h8)
	) name2563 (
		RESET_pad,
		\WX9858_reg/NET0131 ,
		_w4072_
	);
	LUT2 #(
		.INIT('h8)
	) name2564 (
		RESET_pad,
		\WX7216_reg/NET0131 ,
		_w4073_
	);
	LUT2 #(
		.INIT('h8)
	) name2565 (
		RESET_pad,
		\WX2022_reg/NET0131 ,
		_w4074_
	);
	LUT2 #(
		.INIT('h8)
	) name2566 (
		RESET_pad,
		\WX4702_reg/NET0131 ,
		_w4075_
	);
	LUT2 #(
		.INIT('h8)
	) name2567 (
		RESET_pad,
		\WX4524_reg/NET0131 ,
		_w4076_
	);
	LUT2 #(
		.INIT('h8)
	) name2568 (
		RESET_pad,
		\WX5853_reg/NET0131 ,
		_w4077_
	);
	LUT2 #(
		.INIT('h8)
	) name2569 (
		RESET_pad,
		\WX5889_reg/NET0131 ,
		_w4078_
	);
	LUT2 #(
		.INIT('h8)
	) name2570 (
		RESET_pad,
		\WX8477_reg/NET0131 ,
		_w4079_
	);
	LUT2 #(
		.INIT('h8)
	) name2571 (
		RESET_pad,
		\WX4608_reg/NET0131 ,
		_w4080_
	);
	LUT2 #(
		.INIT('h8)
	) name2572 (
		RESET_pad,
		\WX5915_reg/NET0131 ,
		_w4081_
	);
	LUT2 #(
		.INIT('h8)
	) name2573 (
		RESET_pad,
		\WX8495_reg/NET0131 ,
		_w4082_
	);
	LUT2 #(
		.INIT('h8)
	) name2574 (
		RESET_pad,
		\WX3313_reg/NET0131 ,
		_w4083_
	);
	LUT2 #(
		.INIT('h8)
	) name2575 (
		RESET_pad,
		\WX8437_reg/NET0131 ,
		_w4084_
	);
	LUT2 #(
		.INIT('h8)
	) name2576 (
		RESET_pad,
		\WX5935_reg/NET0131 ,
		_w4085_
	);
	LUT2 #(
		.INIT('h8)
	) name2577 (
		RESET_pad,
		\WX715_reg/NET0131 ,
		_w4086_
	);
	LUT2 #(
		.INIT('h8)
	) name2578 (
		RESET_pad,
		\WX8501_reg/NET0131 ,
		_w4087_
	);
	LUT2 #(
		.INIT('h8)
	) name2579 (
		RESET_pad,
		\WX11009_reg/NET0131 ,
		_w4088_
	);
	LUT2 #(
		.INIT('h8)
	) name2580 (
		RESET_pad,
		\WX5931_reg/NET0131 ,
		_w4089_
	);
	LUT2 #(
		.INIT('h8)
	) name2581 (
		RESET_pad,
		\WX4590_reg/NET0131 ,
		_w4090_
	);
	LUT2 #(
		.INIT('h8)
	) name2582 (
		RESET_pad,
		\WX2124_reg/NET0131 ,
		_w4091_
	);
	LUT2 #(
		.INIT('h8)
	) name2583 (
		RESET_pad,
		\WX775_reg/NET0131 ,
		_w4092_
	);
	LUT2 #(
		.INIT('h8)
	) name2584 (
		RESET_pad,
		\WX9792_reg/NET0131 ,
		_w4093_
	);
	LUT2 #(
		.INIT('h8)
	) name2585 (
		RESET_pad,
		\WX811_reg/NET0131 ,
		_w4094_
	);
	LUT2 #(
		.INIT('h8)
	) name2586 (
		RESET_pad,
		\WX8499_reg/NET0131 ,
		_w4095_
	);
	LUT2 #(
		.INIT('h8)
	) name2587 (
		RESET_pad,
		\WX10991_reg/NET0131 ,
		_w4096_
	);
	LUT2 #(
		.INIT('h8)
	) name2588 (
		RESET_pad,
		\WX7162_reg/NET0131 ,
		_w4097_
	);
	LUT2 #(
		.INIT('h8)
	) name2589 (
		RESET_pad,
		\WX3411_reg/NET0131 ,
		_w4098_
	);
	LUT2 #(
		.INIT('h8)
	) name2590 (
		RESET_pad,
		\WX8497_reg/NET0131 ,
		_w4099_
	);
	LUT2 #(
		.INIT('h8)
	) name2591 (
		RESET_pad,
		\WX703_reg/NET0131 ,
		_w4100_
	);
	LUT2 #(
		.INIT('h8)
	) name2592 (
		RESET_pad,
		\WX5917_reg/NET0131 ,
		_w4101_
	);
	LUT2 #(
		.INIT('h8)
	) name2593 (
		RESET_pad,
		\WX11157_reg/NET0131 ,
		_w4102_
	);
	LUT2 #(
		.INIT('h8)
	) name2594 (
		RESET_pad,
		\WX1970_reg/NET0131 ,
		_w4103_
	);
	LUT2 #(
		.INIT('h8)
	) name2595 (
		RESET_pad,
		\WX1974_reg/NET0131 ,
		_w4104_
	);
	LUT2 #(
		.INIT('h8)
	) name2596 (
		RESET_pad,
		\WX8493_reg/NET0131 ,
		_w4105_
	);
	LUT2 #(
		.INIT('h8)
	) name2597 (
		RESET_pad,
		\WX9828_reg/NET0131 ,
		_w4106_
	);
	LUT2 #(
		.INIT('h8)
	) name2598 (
		RESET_pad,
		\WX5911_reg/NET0131 ,
		_w4107_
	);
	LUT2 #(
		.INIT('h8)
	) name2599 (
		RESET_pad,
		\WX797_reg/NET0131 ,
		_w4108_
	);
	LUT2 #(
		.INIT('h8)
	) name2600 (
		RESET_pad,
		\WX1962_reg/NET0131 ,
		_w4109_
	);
	LUT2 #(
		.INIT('h8)
	) name2601 (
		RESET_pad,
		\WX2040_reg/NET0131 ,
		_w4110_
	);
	LUT2 #(
		.INIT('h8)
	) name2602 (
		RESET_pad,
		\WX827_reg/NET0131 ,
		_w4111_
	);
	LUT2 #(
		.INIT('h8)
	) name2603 (
		RESET_pad,
		\WX8487_reg/NET0131 ,
		_w4112_
	);
	LUT2 #(
		.INIT('h8)
	) name2604 (
		RESET_pad,
		\WX5913_reg/NET0131 ,
		_w4113_
	);
	LUT2 #(
		.INIT('h8)
	) name2605 (
		RESET_pad,
		\WX1952_reg/NET0131 ,
		_w4114_
	);
	LUT2 #(
		.INIT('h8)
	) name2606 (
		RESET_pad,
		\WX5905_reg/NET0131 ,
		_w4115_
	);
	LUT2 #(
		.INIT('h8)
	) name2607 (
		RESET_pad,
		\WX3345_reg/NET0131 ,
		_w4116_
	);
	LUT2 #(
		.INIT('h8)
	) name2608 (
		RESET_pad,
		\WX9748_reg/NET0131 ,
		_w4117_
	);
	LUT2 #(
		.INIT('h8)
	) name2609 (
		RESET_pad,
		\WX2058_reg/NET0131 ,
		_w4118_
	);
	LUT2 #(
		.INIT('h8)
	) name2610 (
		RESET_pad,
		\WX5907_reg/NET0131 ,
		_w4119_
	);
	LUT2 #(
		.INIT('h8)
	) name2611 (
		RESET_pad,
		\WX3249_reg/NET0131 ,
		_w4120_
	);
	LUT2 #(
		.INIT('h8)
	) name2612 (
		RESET_pad,
		\WX1944_reg/NET0131 ,
		_w4121_
	);
	LUT2 #(
		.INIT('h8)
	) name2613 (
		RESET_pad,
		\WX4630_reg/NET0131 ,
		_w4122_
	);
	LUT2 #(
		.INIT('h8)
	) name2614 (
		RESET_pad,
		\WX5895_reg/NET0131 ,
		_w4123_
	);
	LUT2 #(
		.INIT('h8)
	) name2615 (
		RESET_pad,
		\WX5887_reg/NET0131 ,
		_w4124_
	);
	LUT2 #(
		.INIT('h8)
	) name2616 (
		RESET_pad,
		\WX1938_reg/NET0131 ,
		_w4125_
	);
	LUT2 #(
		.INIT('h8)
	) name2617 (
		RESET_pad,
		\WX1940_reg/NET0131 ,
		_w4126_
	);
	LUT2 #(
		.INIT('h8)
	) name2618 (
		RESET_pad,
		\WX8403_reg/NET0131 ,
		_w4127_
	);
	LUT2 #(
		.INIT('h8)
	) name2619 (
		RESET_pad,
		\WX725_reg/NET0131 ,
		_w4128_
	);
	LUT2 #(
		.INIT('h8)
	) name2620 (
		RESET_pad,
		\WX5897_reg/NET0131 ,
		_w4129_
	);
	LUT2 #(
		.INIT('h8)
	) name2621 (
		RESET_pad,
		\WX11173_reg/NET0131 ,
		_w4130_
	);
	LUT2 #(
		.INIT('h8)
	) name2622 (
		RESET_pad,
		\WX8425_reg/NET0131 ,
		_w4131_
	);
	LUT2 #(
		.INIT('h8)
	) name2623 (
		RESET_pad,
		\WX7170_reg/NET0131 ,
		_w4132_
	);
	LUT2 #(
		.INIT('h8)
	) name2624 (
		RESET_pad,
		\WX8465_reg/NET0131 ,
		_w4133_
	);
	LUT2 #(
		.INIT('h8)
	) name2625 (
		RESET_pad,
		\WX4530_reg/NET0131 ,
		_w4134_
	);
	LUT2 #(
		.INIT('h8)
	) name2626 (
		RESET_pad,
		\WX7172_reg/NET0131 ,
		_w4135_
	);
	LUT2 #(
		.INIT('h8)
	) name2627 (
		RESET_pad,
		\WX5893_reg/NET0131 ,
		_w4136_
	);
	LUT2 #(
		.INIT('h8)
	) name2628 (
		RESET_pad,
		\WX785_reg/NET0131 ,
		_w4137_
	);
	LUT2 #(
		.INIT('h8)
	) name2629 (
		RESET_pad,
		\WX2050_reg/NET0131 ,
		_w4138_
	);
	LUT2 #(
		.INIT('h8)
	) name2630 (
		RESET_pad,
		\WX8585_reg/NET0131 ,
		_w4139_
	);
	LUT2 #(
		.INIT('h8)
	) name2631 (
		RESET_pad,
		\WX8587_reg/NET0131 ,
		_w4140_
	);
	LUT2 #(
		.INIT('h8)
	) name2632 (
		RESET_pad,
		\WX5891_reg/NET0131 ,
		_w4141_
	);
	LUT2 #(
		.INIT('h8)
	) name2633 (
		RESET_pad,
		\WX671_reg/NET0131 ,
		_w4142_
	);
	LUT2 #(
		.INIT('h8)
	) name2634 (
		RESET_pad,
		\WX2028_reg/NET0131 ,
		_w4143_
	);
	LUT2 #(
		.INIT('h8)
	) name2635 (
		RESET_pad,
		\WX11097_reg/NET0131 ,
		_w4144_
	);
	LUT2 #(
		.INIT('h8)
	) name2636 (
		RESET_pad,
		\WX2116_reg/NET0131 ,
		_w4145_
	);
	LUT2 #(
		.INIT('h8)
	) name2637 (
		RESET_pad,
		\WX11151_reg/NET0131 ,
		_w4146_
	);
	LUT2 #(
		.INIT('h8)
	) name2638 (
		RESET_pad,
		\WX679_reg/NET0131 ,
		_w4147_
	);
	LUT2 #(
		.INIT('h8)
	) name2639 (
		RESET_pad,
		\WX2024_reg/NET0131 ,
		_w4148_
	);
	LUT2 #(
		.INIT('h8)
	) name2640 (
		RESET_pad,
		\WX4706_reg/NET0131 ,
		_w4149_
	);
	LUT2 #(
		.INIT('h8)
	) name2641 (
		RESET_pad,
		\WX7168_reg/NET0131 ,
		_w4150_
	);
	LUT2 #(
		.INIT('h8)
	) name2642 (
		RESET_pad,
		\WX4554_reg/NET0131 ,
		_w4151_
	);
	LUT2 #(
		.INIT('h8)
	) name2643 (
		RESET_pad,
		\WX8421_reg/NET0131 ,
		_w4152_
	);
	LUT2 #(
		.INIT('h8)
	) name2644 (
		RESET_pad,
		\WX2090_reg/NET0131 ,
		_w4153_
	);
	LUT2 #(
		.INIT('h8)
	) name2645 (
		RESET_pad,
		\WX9784_reg/NET0131 ,
		_w4154_
	);
	LUT2 #(
		.INIT('h8)
	) name2646 (
		RESET_pad,
		\WX4714_reg/NET0131 ,
		_w4155_
	);
	LUT2 #(
		.INIT('h8)
	) name2647 (
		RESET_pad,
		\WX11013_reg/NET0131 ,
		_w4156_
	);
	LUT2 #(
		.INIT('h8)
	) name2648 (
		RESET_pad,
		\WX2052_reg/NET0131 ,
		_w4157_
	);
	LUT2 #(
		.INIT('h8)
	) name2649 (
		RESET_pad,
		\WX8417_reg/NET0131 ,
		_w4158_
	);
	LUT2 #(
		.INIT('h8)
	) name2650 (
		RESET_pad,
		\WX3341_reg/NET0131 ,
		_w4159_
	);
	LUT2 #(
		.INIT('h8)
	) name2651 (
		RESET_pad,
		\WX5883_reg/NET0131 ,
		_w4160_
	);
	LUT2 #(
		.INIT('h8)
	) name2652 (
		RESET_pad,
		\WX3323_reg/NET0131 ,
		_w4161_
	);
	LUT2 #(
		.INIT('h8)
	) name2653 (
		RESET_pad,
		\WX9868_reg/NET0131 ,
		_w4162_
	);
	LUT2 #(
		.INIT('h8)
	) name2654 (
		RESET_pad,
		\WX8461_reg/NET0131 ,
		_w4163_
	);
	LUT2 #(
		.INIT('h8)
	) name2655 (
		RESET_pad,
		\WX3329_reg/NET0131 ,
		_w4164_
	);
	LUT2 #(
		.INIT('h8)
	) name2656 (
		RESET_pad,
		\WX11171_reg/NET0131 ,
		_w4165_
	);
	LUT2 #(
		.INIT('h8)
	) name2657 (
		RESET_pad,
		\WX9734_reg/NET0131 ,
		_w4166_
	);
	LUT2 #(
		.INIT('h8)
	) name2658 (
		RESET_pad,
		\WX7176_reg/NET0131 ,
		_w4167_
	);
	LUT2 #(
		.INIT('h8)
	) name2659 (
		RESET_pad,
		\WX2018_reg/NET0131 ,
		_w4168_
	);
	LUT2 #(
		.INIT('h8)
	) name2660 (
		RESET_pad,
		\WX9834_reg/NET0131 ,
		_w4169_
	);
	LUT2 #(
		.INIT('h8)
	) name2661 (
		RESET_pad,
		\WX3401_reg/NET0131 ,
		_w4170_
	);
	LUT2 #(
		.INIT('h8)
	) name2662 (
		RESET_pad,
		\WX2006_reg/NET0131 ,
		_w4171_
	);
	LUT2 #(
		.INIT('h8)
	) name2663 (
		RESET_pad,
		\WX3337_reg/NET0131 ,
		_w4172_
	);
	LUT2 #(
		.INIT('h8)
	) name2664 (
		RESET_pad,
		\WX8503_reg/NET0131 ,
		_w4173_
	);
	LUT2 #(
		.INIT('h8)
	) name2665 (
		RESET_pad,
		\WX5867_reg/NET0131 ,
		_w4174_
	);
	LUT2 #(
		.INIT('h8)
	) name2666 (
		RESET_pad,
		\WX6005_reg/NET0131 ,
		_w4175_
	);
	LUT2 #(
		.INIT('h8)
	) name2667 (
		RESET_pad,
		\WX11025_reg/NET0131 ,
		_w4176_
	);
	LUT2 #(
		.INIT('h8)
	) name2668 (
		RESET_pad,
		\WX1990_reg/NET0131 ,
		_w4177_
	);
	LUT2 #(
		.INIT('h8)
	) name2669 (
		RESET_pad,
		\WX5831_reg/NET0131 ,
		_w4178_
	);
	LUT2 #(
		.INIT('h8)
	) name2670 (
		RESET_pad,
		\WX5955_reg/NET0131 ,
		_w4179_
	);
	LUT2 #(
		.INIT('h8)
	) name2671 (
		RESET_pad,
		\WX8523_reg/NET0131 ,
		_w4180_
	);
	LUT2 #(
		.INIT('h8)
	) name2672 (
		RESET_pad,
		\WX2084_reg/NET0131 ,
		_w4181_
	);
	LUT2 #(
		.INIT('h8)
	) name2673 (
		RESET_pad,
		\WX789_reg/NET0131 ,
		_w4182_
	);
	LUT2 #(
		.INIT('h8)
	) name2674 (
		RESET_pad,
		\WX3381_reg/NET0131 ,
		_w4183_
	);
	LUT2 #(
		.INIT('h8)
	) name2675 (
		RESET_pad,
		\WX5865_reg/NET0131 ,
		_w4184_
	);
	LUT2 #(
		.INIT('h8)
	) name2676 (
		RESET_pad,
		\WX5885_reg/NET0131 ,
		_w4185_
	);
	LUT2 #(
		.INIT('h8)
	) name2677 (
		RESET_pad,
		\WX9794_reg/NET0131 ,
		_w4186_
	);
	LUT2 #(
		.INIT('h8)
	) name2678 (
		RESET_pad,
		\WX5819_reg/NET0131 ,
		_w4187_
	);
	LUT2 #(
		.INIT('h8)
	) name2679 (
		RESET_pad,
		\WX5863_reg/NET0131 ,
		_w4188_
	);
	LUT2 #(
		.INIT('h8)
	) name2680 (
		RESET_pad,
		\WX2042_reg/NET0131 ,
		_w4189_
	);
	LUT2 #(
		.INIT('h8)
	) name2681 (
		RESET_pad,
		\WX7178_reg/NET0131 ,
		_w4190_
	);
	LUT2 #(
		.INIT('h8)
	) name2682 (
		RESET_pad,
		\WX813_reg/NET0131 ,
		_w4191_
	);
	LUT2 #(
		.INIT('h8)
	) name2683 (
		RESET_pad,
		\WX5821_reg/NET0131 ,
		_w4192_
	);
	LUT2 #(
		.INIT('h8)
	) name2684 (
		RESET_pad,
		\WX5851_reg/NET0131 ,
		_w4193_
	);
	LUT2 #(
		.INIT('h8)
	) name2685 (
		RESET_pad,
		\WX8473_reg/NET0131 ,
		_w4194_
	);
	LUT2 #(
		.INIT('h8)
	) name2686 (
		RESET_pad,
		\WX4578_reg/NET0131 ,
		_w4195_
	);
	LUT2 #(
		.INIT('h8)
	) name2687 (
		RESET_pad,
		\WX3421_reg/NET0131 ,
		_w4196_
	);
	LUT2 #(
		.INIT('h8)
	) name2688 (
		RESET_pad,
		\WX9732_reg/NET0131 ,
		_w4197_
	);
	LUT2 #(
		.INIT('h8)
	) name2689 (
		RESET_pad,
		\WX11127_reg/NET0131 ,
		_w4198_
	);
	LUT2 #(
		.INIT('h8)
	) name2690 (
		RESET_pad,
		\WX5847_reg/NET0131 ,
		_w4199_
	);
	LUT2 #(
		.INIT('h8)
	) name2691 (
		RESET_pad,
		\WX8469_reg/NET0131 ,
		_w4200_
	);
	LUT2 #(
		.INIT('h8)
	) name2692 (
		RESET_pad,
		\WX763_reg/NET0131 ,
		_w4201_
	);
	LUT2 #(
		.INIT('h8)
	) name2693 (
		RESET_pad,
		\WX2036_reg/NET0131 ,
		_w4202_
	);
	LUT2 #(
		.INIT('h8)
	) name2694 (
		RESET_pad,
		\WX8475_reg/NET0131 ,
		_w4203_
	);
	LUT2 #(
		.INIT('h8)
	) name2695 (
		RESET_pad,
		\WX11021_reg/NET0131 ,
		_w4204_
	);
	LUT2 #(
		.INIT('h8)
	) name2696 (
		RESET_pad,
		\WX5901_reg/NET0131 ,
		_w4205_
	);
	LUT2 #(
		.INIT('h8)
	) name2697 (
		RESET_pad,
		\WX11005_reg/NET0131 ,
		_w4206_
	);
	LUT2 #(
		.INIT('h8)
	) name2698 (
		RESET_pad,
		\WX3275_reg/NET0131 ,
		_w4207_
	);
	LUT2 #(
		.INIT('h8)
	) name2699 (
		RESET_pad,
		\WX4632_reg/NET0131 ,
		_w4208_
	);
	LUT2 #(
		.INIT('h8)
	) name2700 (
		RESET_pad,
		\WX5841_reg/NET0131 ,
		_w4209_
	);
	LUT2 #(
		.INIT('h8)
	) name2701 (
		RESET_pad,
		\WX5973_reg/NET0131 ,
		_w4210_
	);
	LUT2 #(
		.INIT('h8)
	) name2702 (
		RESET_pad,
		\WX11019_reg/NET0131 ,
		_w4211_
	);
	LUT2 #(
		.INIT('h8)
	) name2703 (
		RESET_pad,
		\WX5829_reg/NET0131 ,
		_w4212_
	);
	LUT2 #(
		.INIT('h8)
	) name2704 (
		RESET_pad,
		\WX647_reg/NET0131 ,
		_w4213_
	);
	LUT2 #(
		.INIT('h8)
	) name2705 (
		RESET_pad,
		\WX5833_reg/NET0131 ,
		_w4214_
	);
	LUT2 #(
		.INIT('h8)
	) name2706 (
		RESET_pad,
		\WX5995_reg/NET0131 ,
		_w4215_
	);
	LUT2 #(
		.INIT('h8)
	) name2707 (
		RESET_pad,
		\WX3261_reg/NET0131 ,
		_w4216_
	);
	LUT2 #(
		.INIT('h8)
	) name2708 (
		RESET_pad,
		\WX7184_reg/NET0131 ,
		_w4217_
	);
	LUT2 #(
		.INIT('h8)
	) name2709 (
		RESET_pad,
		\WX11165_reg/NET0131 ,
		_w4218_
	);
	LUT2 #(
		.INIT('h8)
	) name2710 (
		RESET_pad,
		\WX8419_reg/NET0131 ,
		_w4219_
	);
	LUT2 #(
		.INIT('h8)
	) name2711 (
		RESET_pad,
		\WX697_reg/NET0131 ,
		_w4220_
	);
	LUT2 #(
		.INIT('h8)
	) name2712 (
		RESET_pad,
		\WX5823_reg/NET0131 ,
		_w4221_
	);
	LUT2 #(
		.INIT('h8)
	) name2713 (
		RESET_pad,
		\WX5857_reg/NET0131 ,
		_w4222_
	);
	LUT2 #(
		.INIT('h8)
	) name2714 (
		RESET_pad,
		\WX717_reg/NET0131 ,
		_w4223_
	);
	LUT2 #(
		.INIT('h8)
	) name2715 (
		RESET_pad,
		\WX4528_reg/NET0131 ,
		_w4224_
	);
	LUT2 #(
		.INIT('h8)
	) name2716 (
		RESET_pad,
		\WX5843_reg/NET0131 ,
		_w4225_
	);
	LUT2 #(
		.INIT('h8)
	) name2717 (
		RESET_pad,
		\WX5827_reg/NET0131 ,
		_w4226_
	);
	LUT2 #(
		.INIT('h8)
	) name2718 (
		RESET_pad,
		\WX7254_reg/NET0131 ,
		_w4227_
	);
	LUT2 #(
		.INIT('h8)
	) name2719 (
		RESET_pad,
		\WX5835_reg/NET0131 ,
		_w4228_
	);
	LUT2 #(
		.INIT('h8)
	) name2720 (
		RESET_pad,
		\WX737_reg/NET0131 ,
		_w4229_
	);
	LUT2 #(
		.INIT('h8)
	) name2721 (
		RESET_pad,
		\WX3293_reg/NET0131 ,
		_w4230_
	);
	LUT2 #(
		.INIT('h8)
	) name2722 (
		RESET_pad,
		\WX9846_reg/NET0131 ,
		_w4231_
	);
	LUT2 #(
		.INIT('h8)
	) name2723 (
		RESET_pad,
		\WX1964_reg/NET0131 ,
		_w4232_
	);
	LUT2 #(
		.INIT('h8)
	) name2724 (
		RESET_pad,
		\WX9814_reg/NET0131 ,
		_w4233_
	);
	LUT2 #(
		.INIT('h8)
	) name2725 (
		RESET_pad,
		\WX8505_reg/NET0131 ,
		_w4234_
	);
	LUT2 #(
		.INIT('h8)
	) name2726 (
		RESET_pad,
		\WX4658_reg/NET0131 ,
		_w4235_
	);
	LUT2 #(
		.INIT('h8)
	) name2727 (
		RESET_pad,
		\WX5825_reg/NET0131 ,
		_w4236_
	);
	LUT2 #(
		.INIT('h8)
	) name2728 (
		RESET_pad,
		\WX7188_reg/NET0131 ,
		_w4237_
	);
	LUT2 #(
		.INIT('h8)
	) name2729 (
		RESET_pad,
		\WX3399_reg/NET0131 ,
		_w4238_
	);
	LUT2 #(
		.INIT('h8)
	) name2730 (
		RESET_pad,
		\WX2034_reg/NET0131 ,
		_w4239_
	);
	LUT2 #(
		.INIT('h8)
	) name2731 (
		RESET_pad,
		\WX8471_reg/NET0131 ,
		_w4240_
	);
	LUT2 #(
		.INIT('h8)
	) name2732 (
		RESET_pad,
		\WX1968_reg/NET0131 ,
		_w4241_
	);
	LUT2 #(
		.INIT('h8)
	) name2733 (
		RESET_pad,
		\WX7290_reg/NET0131 ,
		_w4242_
	);
	LUT2 #(
		.INIT('h8)
	) name2734 (
		RESET_pad,
		\WX11101_reg/NET0131 ,
		_w4243_
	);
	LUT2 #(
		.INIT('h8)
	) name2735 (
		RESET_pad,
		\WX5837_reg/NET0131 ,
		_w4244_
	);
	LUT2 #(
		.INIT('h8)
	) name2736 (
		RESET_pad,
		\WX8459_reg/NET0131 ,
		_w4245_
	);
	LUT2 #(
		.INIT('h8)
	) name2737 (
		RESET_pad,
		\WX5817_reg/NET0131 ,
		_w4246_
	);
	LUT2 #(
		.INIT('h8)
	) name2738 (
		RESET_pad,
		\WX4668_reg/NET0131 ,
		_w4247_
	);
	LUT2 #(
		.INIT('h8)
	) name2739 (
		RESET_pad,
		\WX4614_reg/NET0131 ,
		_w4248_
	);
	LUT2 #(
		.INIT('h8)
	) name2740 (
		RESET_pad,
		\WX4672_reg/NET0131 ,
		_w4249_
	);
	LUT2 #(
		.INIT('h8)
	) name2741 (
		RESET_pad,
		\WX9844_reg/NET0131 ,
		_w4250_
	);
	LUT2 #(
		.INIT('h8)
	) name2742 (
		RESET_pad,
		\WX4648_reg/NET0131 ,
		_w4251_
	);
	LUT2 #(
		.INIT('h8)
	) name2743 (
		RESET_pad,
		\WX3325_reg/NET0131 ,
		_w4252_
	);
	LUT2 #(
		.INIT('h8)
	) name2744 (
		RESET_pad,
		\WX713_reg/NET0131 ,
		_w4253_
	);
	LUT2 #(
		.INIT('h8)
	) name2745 (
		RESET_pad,
		\WX11069_reg/NET0131 ,
		_w4254_
	);
	LUT2 #(
		.INIT('h8)
	) name2746 (
		RESET_pad,
		\WX9746_reg/NET0131 ,
		_w4255_
	);
	LUT2 #(
		.INIT('h8)
	) name2747 (
		RESET_pad,
		\WX9874_reg/NET0131 ,
		_w4256_
	);
	LUT2 #(
		.INIT('h8)
	) name2748 (
		RESET_pad,
		\WX8451_reg/NET0131 ,
		_w4257_
	);
	LUT2 #(
		.INIT('h8)
	) name2749 (
		RESET_pad,
		\WX1950_reg/NET0131 ,
		_w4258_
	);
	LUT2 #(
		.INIT('h8)
	) name2750 (
		RESET_pad,
		\WX5909_reg/NET0131 ,
		_w4259_
	);
	LUT2 #(
		.INIT('h8)
	) name2751 (
		RESET_pad,
		\WX8515_reg/NET0131 ,
		_w4260_
	);
	LUT2 #(
		.INIT('h8)
	) name2752 (
		RESET_pad,
		\WX1960_reg/NET0131 ,
		_w4261_
	);
	LUT2 #(
		.INIT('h8)
	) name2753 (
		RESET_pad,
		\WX7236_reg/NET0131 ,
		_w4262_
	);
	LUT2 #(
		.INIT('h8)
	) name2754 (
		RESET_pad,
		\WX4700_reg/NET0131 ,
		_w4263_
	);
	LUT2 #(
		.INIT('h8)
	) name2755 (
		RESET_pad,
		\WX4692_reg/NET0131 ,
		_w4264_
	);
	LUT2 #(
		.INIT('h8)
	) name2756 (
		RESET_pad,
		\WX1976_reg/NET0131 ,
		_w4265_
	);
	LUT2 #(
		.INIT('h8)
	) name2757 (
		RESET_pad,
		\WX1980_reg/NET0131 ,
		_w4266_
	);
	LUT2 #(
		.INIT('h8)
	) name2758 (
		RESET_pad,
		\WX8443_reg/NET0131 ,
		_w4267_
	);
	LUT2 #(
		.INIT('h8)
	) name2759 (
		RESET_pad,
		\WX1996_reg/NET0131 ,
		_w4268_
	);
	LUT2 #(
		.INIT('h8)
	) name2760 (
		RESET_pad,
		\WX2032_reg/NET0131 ,
		_w4269_
	);
	LUT2 #(
		.INIT('h8)
	) name2761 (
		RESET_pad,
		\WX9848_reg/NET0131 ,
		_w4270_
	);
	LUT2 #(
		.INIT('h8)
	) name2762 (
		RESET_pad,
		\WX11023_reg/NET0131 ,
		_w4271_
	);
	LUT2 #(
		.INIT('h8)
	) name2763 (
		RESET_pad,
		\WX3317_reg/NET0131 ,
		_w4272_
	);
	LUT2 #(
		.INIT('h8)
	) name2764 (
		RESET_pad,
		\WX9740_reg/NET0131 ,
		_w4273_
	);
	LUT2 #(
		.INIT('h8)
	) name2765 (
		RESET_pad,
		\WX2014_reg/NET0131 ,
		_w4274_
	);
	LUT2 #(
		.INIT('h8)
	) name2766 (
		RESET_pad,
		\WX11155_reg/NET0131 ,
		_w4275_
	);
	LUT2 #(
		.INIT('h8)
	) name2767 (
		RESET_pad,
		\WX2020_reg/NET0131 ,
		_w4276_
	);
	LUT2 #(
		.INIT('h8)
	) name2768 (
		RESET_pad,
		\WX6007_reg/NET0131 ,
		_w4277_
	);
	LUT2 #(
		.INIT('h8)
	) name2769 (
		RESET_pad,
		\WX4708_reg/NET0131 ,
		_w4278_
	);
	LUT2 #(
		.INIT('h8)
	) name2770 (
		RESET_pad,
		\WX2044_reg/NET0131 ,
		_w4279_
	);
	LUT2 #(
		.INIT('h8)
	) name2771 (
		RESET_pad,
		\WX2046_reg/NET0131 ,
		_w4280_
	);
	LUT2 #(
		.INIT('h8)
	) name2772 (
		RESET_pad,
		\WX3359_reg/NET0131 ,
		_w4281_
	);
	LUT2 #(
		.INIT('h8)
	) name2773 (
		RESET_pad,
		\WX2054_reg/NET0131 ,
		_w4282_
	);
	LUT2 #(
		.INIT('h8)
	) name2774 (
		RESET_pad,
		\WX5869_reg/NET0131 ,
		_w4283_
	);
	LUT2 #(
		.INIT('h8)
	) name2775 (
		RESET_pad,
		\WX11179_reg/NET0131 ,
		_w4284_
	);
	LUT2 #(
		.INIT('h8)
	) name2776 (
		RESET_pad,
		\WX11129_reg/NET0131 ,
		_w4285_
	);
	LUT2 #(
		.INIT('h8)
	) name2777 (
		RESET_pad,
		\WX11145_reg/NET0131 ,
		_w4286_
	);
	LUT2 #(
		.INIT('h8)
	) name2778 (
		RESET_pad,
		\WX699_reg/NET0131 ,
		_w4287_
	);
	LUT2 #(
		.INIT('h8)
	) name2779 (
		RESET_pad,
		\WX2080_reg/NET0131 ,
		_w4288_
	);
	LUT2 #(
		.INIT('h8)
	) name2780 (
		RESET_pad,
		\WX2082_reg/NET0131 ,
		_w4289_
	);
	LUT2 #(
		.INIT('h8)
	) name2781 (
		RESET_pad,
		\WX2030_reg/NET0131 ,
		_w4290_
	);
	LUT2 #(
		.INIT('h8)
	) name2782 (
		RESET_pad,
		\WX11075_reg/NET0131 ,
		_w4291_
	);
	LUT2 #(
		.INIT('h8)
	) name2783 (
		RESET_pad,
		\WX3311_reg/NET0131 ,
		_w4292_
	);
	LUT2 #(
		.INIT('h8)
	) name2784 (
		RESET_pad,
		\WX9818_reg/NET0131 ,
		_w4293_
	);
	LUT2 #(
		.INIT('h8)
	) name2785 (
		RESET_pad,
		\WX701_reg/NET0131 ,
		_w4294_
	);
	LUT2 #(
		.INIT('h8)
	) name2786 (
		RESET_pad,
		\WX2026_reg/NET0131 ,
		_w4295_
	);
	LUT2 #(
		.INIT('h8)
	) name2787 (
		RESET_pad,
		\WX5839_reg/NET0131 ,
		_w4296_
	);
	LUT2 #(
		.INIT('h8)
	) name2788 (
		RESET_pad,
		\WX11007_reg/NET0131 ,
		_w4297_
	);
	LUT2 #(
		.INIT('h8)
	) name2789 (
		RESET_pad,
		\WX8563_reg/NET0131 ,
		_w4298_
	);
	LUT2 #(
		.INIT('h8)
	) name2790 (
		RESET_pad,
		\WX3309_reg/NET0131 ,
		_w4299_
	);
	LUT2 #(
		.INIT('h8)
	) name2791 (
		RESET_pad,
		\WX9710_reg/NET0131 ,
		_w4300_
	);
	LUT2 #(
		.INIT('h8)
	) name2792 (
		RESET_pad,
		\WX4574_reg/NET0131 ,
		_w4301_
	);
	LUT2 #(
		.INIT('h8)
	) name2793 (
		RESET_pad,
		\WX7202_reg/NET0131 ,
		_w4302_
	);
	LUT2 #(
		.INIT('h8)
	) name2794 (
		RESET_pad,
		\WX8415_reg/NET0131 ,
		_w4303_
	);
	LUT2 #(
		.INIT('h8)
	) name2795 (
		RESET_pad,
		\WX9810_reg/NET0131 ,
		_w4304_
	);
	LUT2 #(
		.INIT('h8)
	) name2796 (
		RESET_pad,
		\WX3269_reg/NET0131 ,
		_w4305_
	);
	LUT2 #(
		.INIT('h8)
	) name2797 (
		RESET_pad,
		\WX7200_reg/NET0131 ,
		_w4306_
	);
	LUT2 #(
		.INIT('h8)
	) name2798 (
		RESET_pad,
		\WX9752_reg/NET0131 ,
		_w4307_
	);
	LUT2 #(
		.INIT('h8)
	) name2799 (
		RESET_pad,
		\WX7174_reg/NET0131 ,
		_w4308_
	);
	LUT2 #(
		.INIT('h8)
	) name2800 (
		RESET_pad,
		\WX3389_reg/NET0131 ,
		_w4309_
	);
	LUT2 #(
		.INIT('h8)
	) name2801 (
		RESET_pad,
		\WX8581_reg/NET0131 ,
		_w4310_
	);
	LUT2 #(
		.INIT('h8)
	) name2802 (
		RESET_pad,
		\WX5845_reg/NET0131 ,
		_w4311_
	);
	LUT2 #(
		.INIT('h8)
	) name2803 (
		RESET_pad,
		\WX5873_reg/NET0131 ,
		_w4312_
	);
	LUT2 #(
		.INIT('h8)
	) name2804 (
		RESET_pad,
		\WX9782_reg/NET0131 ,
		_w4313_
	);
	LUT2 #(
		.INIT('h8)
	) name2805 (
		RESET_pad,
		\WX7208_reg/NET0131 ,
		_w4314_
	);
	LUT2 #(
		.INIT('h8)
	) name2806 (
		RESET_pad,
		\WX8485_reg/NET0131 ,
		_w4315_
	);
	LUT2 #(
		.INIT('h8)
	) name2807 (
		RESET_pad,
		\WX8575_reg/NET0131 ,
		_w4316_
	);
	LUT2 #(
		.INIT('h8)
	) name2808 (
		RESET_pad,
		\WX8481_reg/NET0131 ,
		_w4317_
	);
	LUT2 #(
		.INIT('h8)
	) name2809 (
		RESET_pad,
		\WX4532_reg/NET0131 ,
		_w4318_
	);
	LUT2 #(
		.INIT('h8)
	) name2810 (
		RESET_pad,
		\WX11031_reg/NET0131 ,
		_w4319_
	);
	LUT2 #(
		.INIT('h8)
	) name2811 (
		RESET_pad,
		\WX7210_reg/NET0131 ,
		_w4320_
	);
	LUT2 #(
		.INIT('h8)
	) name2812 (
		RESET_pad,
		\WX7206_reg/NET0131 ,
		_w4321_
	);
	LUT2 #(
		.INIT('h8)
	) name2813 (
		RESET_pad,
		\WX10989_reg/NET0131 ,
		_w4322_
	);
	LUT2 #(
		.INIT('h8)
	) name2814 (
		RESET_pad,
		\WX765_reg/NET0131 ,
		_w4323_
	);
	LUT2 #(
		.INIT('h8)
	) name2815 (
		RESET_pad,
		\WX799_reg/NET0131 ,
		_w4324_
	);
	LUT2 #(
		.INIT('h8)
	) name2816 (
		RESET_pad,
		\WX711_reg/NET0131 ,
		_w4325_
	);
	LUT2 #(
		.INIT('h8)
	) name2817 (
		RESET_pad,
		\WX751_reg/NET0131 ,
		_w4326_
	);
	LUT2 #(
		.INIT('h8)
	) name2818 (
		RESET_pad,
		\WX10993_reg/NET0131 ,
		_w4327_
	);
	LUT2 #(
		.INIT('h8)
	) name2819 (
		RESET_pad,
		\WX3413_reg/NET0131 ,
		_w4328_
	);
	LUT2 #(
		.INIT('h8)
	) name2820 (
		RESET_pad,
		\WX8577_reg/NET0131 ,
		_w4329_
	);
	LUT2 #(
		.INIT('h8)
	) name2821 (
		RESET_pad,
		\WX3291_reg/NET0131 ,
		_w4330_
	);
	LUT2 #(
		.INIT('h8)
	) name2822 (
		RESET_pad,
		\WX741_reg/NET0131 ,
		_w4331_
	);
	LUT2 #(
		.INIT('h8)
	) name2823 (
		RESET_pad,
		\WX749_reg/NET0131 ,
		_w4332_
	);
	LUT2 #(
		.INIT('h8)
	) name2824 (
		RESET_pad,
		\WX7266_reg/NET0131 ,
		_w4333_
	);
	LUT2 #(
		.INIT('h8)
	) name2825 (
		RESET_pad,
		\WX4568_reg/NET0131 ,
		_w4334_
	);
	LUT2 #(
		.INIT('h8)
	) name2826 (
		RESET_pad,
		\WX8527_reg/NET0131 ,
		_w4335_
	);
	LUT2 #(
		.INIT('h8)
	) name2827 (
		RESET_pad,
		\WX1982_reg/NET0131 ,
		_w4336_
	);
	LUT2 #(
		.INIT('h8)
	) name2828 (
		RESET_pad,
		\WX11035_reg/NET0131 ,
		_w4337_
	);
	LUT2 #(
		.INIT('h8)
	) name2829 (
		RESET_pad,
		\WX11039_reg/NET0131 ,
		_w4338_
	);
	LUT2 #(
		.INIT('h8)
	) name2830 (
		RESET_pad,
		\WX3251_reg/NET0131 ,
		_w4339_
	);
	LUT2 #(
		.INIT('h8)
	) name2831 (
		RESET_pad,
		\WX745_reg/NET0131 ,
		_w4340_
	);
	LUT3 #(
		.INIT('he0)
	) name2832 (
		\TM0_pad ,
		_w1516_,
		_w1865_,
		_w4341_
	);
	LUT4 #(
		.INIT('h0a02)
	) name2833 (
		RESET_pad,
		\TM0_pad ,
		\TM1_pad ,
		\_2088__reg/NET0131 ,
		_w4342_
	);
	LUT4 #(
		.INIT('hbe00)
	) name2834 (
		\TM0_pad ,
		_w2681_,
		_w2682_,
		_w4342_,
		_w4343_
	);
	LUT2 #(
		.INIT('he)
	) name2835 (
		_w4341_,
		_w4343_,
		_w4344_
	);
	LUT3 #(
		.INIT('he0)
	) name2836 (
		\TM0_pad ,
		_w1600_,
		_w1620_,
		_w4345_
	);
	LUT4 #(
		.INIT('h0a02)
	) name2837 (
		RESET_pad,
		\TM0_pad ,
		\TM1_pad ,
		\_2085__reg/NET0131 ,
		_w4346_
	);
	LUT4 #(
		.INIT('hbe00)
	) name2838 (
		\TM0_pad ,
		_w2804_,
		_w2805_,
		_w4346_,
		_w4347_
	);
	LUT2 #(
		.INIT('he)
	) name2839 (
		_w4345_,
		_w4347_,
		_w4348_
	);
	LUT3 #(
		.INIT('he0)
	) name2840 (
		\TM0_pad ,
		_w1588_,
		_w2258_,
		_w4349_
	);
	LUT4 #(
		.INIT('h0a02)
	) name2841 (
		RESET_pad,
		\TM0_pad ,
		\TM1_pad ,
		\_2081__reg/NET0131 ,
		_w4350_
	);
	LUT4 #(
		.INIT('hbe00)
	) name2842 (
		\TM0_pad ,
		_w2981_,
		_w2982_,
		_w4350_,
		_w4351_
	);
	LUT2 #(
		.INIT('he)
	) name2843 (
		_w4349_,
		_w4351_,
		_w4352_
	);
	LUT3 #(
		.INIT('he0)
	) name2844 (
		\TM0_pad ,
		_w1525_,
		_w1706_,
		_w4353_
	);
	LUT4 #(
		.INIT('h0a02)
	) name2845 (
		RESET_pad,
		\TM0_pad ,
		\TM1_pad ,
		\_2091__reg/NET0131 ,
		_w4354_
	);
	LUT4 #(
		.INIT('hbe00)
	) name2846 (
		\TM0_pad ,
		_w2540_,
		_w2541_,
		_w4354_,
		_w4355_
	);
	LUT2 #(
		.INIT('he)
	) name2847 (
		_w4353_,
		_w4355_,
		_w4356_
	);
	LUT3 #(
		.INIT('he0)
	) name2848 (
		\TM0_pad ,
		_w1603_,
		_w1978_,
		_w4357_
	);
	LUT4 #(
		.INIT('h0a02)
	) name2849 (
		RESET_pad,
		\TM0_pad ,
		\TM1_pad ,
		\_2086__reg/NET0131 ,
		_w4358_
	);
	LUT4 #(
		.INIT('hbe00)
	) name2850 (
		\TM0_pad ,
		_w2764_,
		_w2765_,
		_w4358_,
		_w4359_
	);
	LUT2 #(
		.INIT('he)
	) name2851 (
		_w4357_,
		_w4359_,
		_w4360_
	);
	LUT3 #(
		.INIT('he0)
	) name2852 (
		\TM0_pad ,
		_w1597_,
		_w2089_,
		_w4361_
	);
	LUT4 #(
		.INIT('h0a02)
	) name2853 (
		RESET_pad,
		\TM0_pad ,
		\TM1_pad ,
		\_2084__reg/NET0131 ,
		_w4362_
	);
	LUT4 #(
		.INIT('hbe00)
	) name2854 (
		\TM0_pad ,
		_w2843_,
		_w2844_,
		_w4362_,
		_w4363_
	);
	LUT2 #(
		.INIT('he)
	) name2855 (
		_w4361_,
		_w4363_,
		_w4364_
	);
	LUT3 #(
		.INIT('he0)
	) name2856 (
		\TM0_pad ,
		_w1543_,
		_w2422_,
		_w4365_
	);
	LUT4 #(
		.INIT('h0a02)
	) name2857 (
		RESET_pad,
		\TM0_pad ,
		\TM1_pad ,
		\_2078__reg/NET0131 ,
		_w4366_
	);
	LUT4 #(
		.INIT('hbe00)
	) name2858 (
		\TM0_pad ,
		_w3147_,
		_w3148_,
		_w4366_,
		_w4367_
	);
	LUT2 #(
		.INIT('he)
	) name2859 (
		_w4365_,
		_w4367_,
		_w4368_
	);
	LUT4 #(
		.INIT('h8cc8)
	) name2860 (
		\TM0_pad ,
		_w1606_,
		_w1942_,
		_w1943_,
		_w4369_
	);
	LUT2 #(
		.INIT('h2)
	) name2861 (
		\TM0_pad ,
		\_2348__reg/NET0131 ,
		_w4370_
	);
	LUT4 #(
		.INIT('h00c8)
	) name2862 (
		\DATA_0_15_pad ,
		RESET_pad,
		\TM0_pad ,
		\TM1_pad ,
		_w4371_
	);
	LUT2 #(
		.INIT('h4)
	) name2863 (
		_w4370_,
		_w4371_,
		_w4372_
	);
	LUT2 #(
		.INIT('he)
	) name2864 (
		_w4369_,
		_w4372_,
		_w4373_
	);
	assign \DATA_9_0_pad  = _w1511_ ;
	assign \DATA_9_10_pad  = _w1514_ ;
	assign \DATA_9_11_pad  = _w1517_ ;
	assign \DATA_9_12_pad  = _w1520_ ;
	assign \DATA_9_13_pad  = _w1523_ ;
	assign \DATA_9_14_pad  = _w1526_ ;
	assign \DATA_9_15_pad  = _w1529_ ;
	assign \DATA_9_16_pad  = _w1532_ ;
	assign \DATA_9_17_pad  = _w1535_ ;
	assign \DATA_9_18_pad  = _w1538_ ;
	assign \DATA_9_19_pad  = _w1541_ ;
	assign \DATA_9_1_pad  = _w1544_ ;
	assign \DATA_9_20_pad  = _w1547_ ;
	assign \DATA_9_21_pad  = _w1550_ ;
	assign \DATA_9_22_pad  = _w1553_ ;
	assign \DATA_9_23_pad  = _w1556_ ;
	assign \DATA_9_24_pad  = _w1559_ ;
	assign \DATA_9_25_pad  = _w1562_ ;
	assign \DATA_9_26_pad  = _w1565_ ;
	assign \DATA_9_27_pad  = _w1568_ ;
	assign \DATA_9_28_pad  = _w1571_ ;
	assign \DATA_9_29_pad  = _w1574_ ;
	assign \DATA_9_2_pad  = _w1577_ ;
	assign \DATA_9_30_pad  = _w1580_ ;
	assign \DATA_9_31_pad  = _w1583_ ;
	assign \DATA_9_3_pad  = _w1586_ ;
	assign \DATA_9_4_pad  = _w1589_ ;
	assign \DATA_9_5_pad  = _w1592_ ;
	assign \DATA_9_6_pad  = _w1595_ ;
	assign \DATA_9_7_pad  = _w1598_ ;
	assign \DATA_9_8_pad  = _w1601_ ;
	assign \DATA_9_9_pad  = _w1604_ ;
	assign \_al_n0  = 1'b0;
	assign \_al_n1  = 1'b1;
	assign \g19/_0_  = _w1612_ ;
	assign \g35/_0_  = _w1619_ ;
	assign \g36/_0_  = _w1627_ ;
	assign \g40/_0_  = _w1635_ ;
	assign \g55780/_0_  = _w1640_ ;
	assign \g55783/_0_  = _w1645_ ;
	assign \g55795/_0_  = _w1653_ ;
	assign \g55796/_0_  = _w1658_ ;
	assign \g55797/_0_  = _w1665_ ;
	assign \g55798/_0_  = _w1672_ ;
	assign \g55799/_0_  = _w1679_ ;
	assign \g55800/_0_  = _w1686_ ;
	assign \g55801/_0_  = _w1693_ ;
	assign \g55802/_0_  = _w1698_ ;
	assign \g55803/_0_  = _w1705_ ;
	assign \g55834/_0_  = _w1714_ ;
	assign \g55835/_0_  = _w1719_ ;
	assign \g55836/_0_  = _w1724_ ;
	assign \g55837/_0_  = _w1729_ ;
	assign \g55838/_0_  = _w1735_ ;
	assign \g55839/_0_  = _w1740_ ;
	assign \g55840/_0_  = _w1745_ ;
	assign \g55841/_0_  = _w1750_ ;
	assign \g55842/_0_  = _w1757_ ;
	assign \g55856/_0_  = _w1758_ ;
	assign \g55894/_0_  = _w1766_ ;
	assign \g55895/_0_  = _w1771_ ;
	assign \g55896/_0_  = _w1776_ ;
	assign \g55897/_0_  = _w1781_ ;
	assign \g55898/_0_  = _w1787_ ;
	assign \g55899/_0_  = _w1793_ ;
	assign \g55900/_0_  = _w1798_ ;
	assign \g55901/_0_  = _w1803_ ;
	assign \g55902/_0_  = _w1808_ ;
	assign \g55916/_0_  = _w1809_ ;
	assign \g55953/_0_  = _w1818_ ;
	assign \g55954/_0_  = _w1823_ ;
	assign \g55955/_0_  = _w1828_ ;
	assign \g55956/_0_  = _w1833_ ;
	assign \g55957/_0_  = _w1839_ ;
	assign \g55958/_0_  = _w1845_ ;
	assign \g55959/_0_  = _w1851_ ;
	assign \g55960/_0_  = _w1856_ ;
	assign \g55961/_0_  = _w1863_ ;
	assign \g55975/_0_  = _w1864_ ;
	assign \g56012/_0_  = _w1873_ ;
	assign \g56013/_0_  = _w1879_ ;
	assign \g56014/_0_  = _w1884_ ;
	assign \g56015/_0_  = _w1889_ ;
	assign \g56016/_0_  = _w1895_ ;
	assign \g56017/_0_  = _w1901_ ;
	assign \g56018/_0_  = _w1907_ ;
	assign \g56019/_0_  = _w1912_ ;
	assign \g56020/_0_  = _w1919_ ;
	assign \g56034/_0_  = _w1920_ ;
	assign \g56071/_0_  = _w1929_ ;
	assign \g56072/_0_  = _w1935_ ;
	assign \g56073/_0_  = _w1940_ ;
	assign \g56074/_0_  = _w1946_ ;
	assign \g56075/_0_  = _w1952_ ;
	assign \g56076/_0_  = _w1958_ ;
	assign \g56077/_0_  = _w1964_ ;
	assign \g56078/_0_  = _w1969_ ;
	assign \g56079/_0_  = _w1976_ ;
	assign \g56093/_0_  = _w1977_ ;
	assign \g56130/_0_  = _w1986_ ;
	assign \g56131/_0_  = _w1992_ ;
	assign \g56132/_0_  = _w1998_ ;
	assign \g56133/_0_  = _w2003_ ;
	assign \g56134/_0_  = _w2009_ ;
	assign \g56135/_0_  = _w2015_ ;
	assign \g56136/_0_  = _w2021_ ;
	assign \g56137/_0_  = _w2026_ ;
	assign \g56138/_0_  = _w2033_ ;
	assign \g56152/_0_  = _w2034_ ;
	assign \g56189/_0_  = _w2042_ ;
	assign \g56190/_0_  = _w2048_ ;
	assign \g56191/_0_  = _w2052_ ;
	assign \g56192/_0_  = _w2057_ ;
	assign \g56193/_0_  = _w2063_ ;
	assign \g56194/_0_  = _w2069_ ;
	assign \g56195/_0_  = _w2075_ ;
	assign \g56196/_0_  = _w2080_ ;
	assign \g56197/_0_  = _w2087_ ;
	assign \g56211/_0_  = _w2088_ ;
	assign \g56248/_0_  = _w2097_ ;
	assign \g56249/_0_  = _w2103_ ;
	assign \g56250/_0_  = _w2109_ ;
	assign \g56251/_0_  = _w2114_ ;
	assign \g56252/_0_  = _w2120_ ;
	assign \g56253/_0_  = _w2126_ ;
	assign \g56254/_0_  = _w2132_ ;
	assign \g56255/_0_  = _w2137_ ;
	assign \g56256/_0_  = _w2144_ ;
	assign \g56270/_0_  = _w2145_ ;
	assign \g56307/_0_  = _w2154_ ;
	assign \g56308/_0_  = _w2160_ ;
	assign \g56309/_0_  = _w2166_ ;
	assign \g56310/_0_  = _w2171_ ;
	assign \g56311/_0_  = _w2177_ ;
	assign \g56312/_0_  = _w2183_ ;
	assign \g56313/_0_  = _w2189_ ;
	assign \g56314/_0_  = _w2194_ ;
	assign \g56315/_0_  = _w2201_ ;
	assign \g56329/_0_  = _w2202_ ;
	assign \g56366/_0_  = _w2211_ ;
	assign \g56367/_0_  = _w2217_ ;
	assign \g56368/_0_  = _w2223_ ;
	assign \g56369/_0_  = _w2228_ ;
	assign \g56370/_0_  = _w2234_ ;
	assign \g56371/_0_  = _w2240_ ;
	assign \g56372/_0_  = _w2246_ ;
	assign \g56373/_0_  = _w2251_ ;
	assign \g56374/_0_  = _w2256_ ;
	assign \g56388/_0_  = _w2257_ ;
	assign \g56425/_0_  = _w2266_ ;
	assign \g56426/_0_  = _w2272_ ;
	assign \g56427/_0_  = _w2278_ ;
	assign \g56428/_0_  = _w2283_ ;
	assign \g56429/_0_  = _w2289_ ;
	assign \g56430/_0_  = _w2295_ ;
	assign \g56431/_0_  = _w2301_ ;
	assign \g56432/_0_  = _w2306_ ;
	assign \g56433/_0_  = _w2311_ ;
	assign \g56447/_0_  = _w2312_ ;
	assign \g56484/_0_  = _w2321_ ;
	assign \g56485/_0_  = _w2327_ ;
	assign \g56486/_0_  = _w2331_ ;
	assign \g56487/_0_  = _w2336_ ;
	assign \g56488/_0_  = _w2342_ ;
	assign \g56489/_0_  = _w2348_ ;
	assign \g56490/_0_  = _w2354_ ;
	assign \g56491/_0_  = _w2359_ ;
	assign \g56492/_0_  = _w2364_ ;
	assign \g56507/_0_  = _w2365_ ;
	assign \g56543/_0_  = _w2374_ ;
	assign \g56544/_0_  = _w2380_ ;
	assign \g56545/_0_  = _w2386_ ;
	assign \g56546/_0_  = _w2392_ ;
	assign \g56547/_0_  = _w2397_ ;
	assign \g56548/_0_  = _w2403_ ;
	assign \g56549/_0_  = _w2409_ ;
	assign \g56551/_0_  = _w2414_ ;
	assign \g56567/_0_  = _w2415_ ;
	assign \g56602/_0_  = _w2421_ ;
	assign \g56603/_0_  = _w2430_ ;
	assign \g56604/_0_  = _w2436_ ;
	assign \g56605/_0_  = _w2442_ ;
	assign \g56606/_0_  = _w2448_ ;
	assign \g56607/_0_  = _w2453_ ;
	assign \g56608/_0_  = _w2459_ ;
	assign \g56610/_0_  = _w2464_ ;
	assign \g56627/_0_  = _w2465_ ;
	assign \g56661/_0_  = _w2471_ ;
	assign \g56662/_0_  = _w2480_ ;
	assign \g56663/_0_  = _w2486_ ;
	assign \g56664/_0_  = _w2492_ ;
	assign \g56665/_0_  = _w2498_ ;
	assign \g56666/_0_  = _w2502_ ;
	assign \g56667/_0_  = _w2508_ ;
	assign \g56668/_0_  = _w2514_ ;
	assign \g56686/_0_  = _w2515_ ;
	assign \g56720/_0_  = _w2521_ ;
	assign \g56721/_0_  = _w2527_ ;
	assign \g56722/_0_  = _w2533_ ;
	assign \g56723/_0_  = _w2539_ ;
	assign \g56724/_0_  = _w2545_ ;
	assign \g56725/_0_  = _w2551_ ;
	assign \g56726/_0_  = _w2558_ ;
	assign \g56727/_0_  = _w2564_ ;
	assign \g56728/_0_  = _w2569_ ;
	assign \g56745/_0_  = _w2570_ ;
	assign \g56779/_0_  = _w2576_ ;
	assign \g56780/_0_  = _w2582_ ;
	assign \g56781/_0_  = _w2587_ ;
	assign \g56782/_0_  = _w2593_ ;
	assign \g56783/_0_  = _w2597_ ;
	assign \g56784/_0_  = _w2603_ ;
	assign \g56785/_0_  = _w2608_ ;
	assign \g56804/_0_  = _w2609_ ;
	assign \g56838/_0_  = _w2615_ ;
	assign \g56839/_0_  = _w2621_ ;
	assign \g56840/_0_  = _w2626_ ;
	assign \g56841/_0_  = _w2632_ ;
	assign \g56842/_0_  = _w2637_ ;
	assign \g56843/_0_  = _w2641_ ;
	assign \g56844/_0_  = _w2646_ ;
	assign \g56845/_0_  = _w2652_ ;
	assign \g56846/_0_  = _w2657_ ;
	assign \g56863/_0_  = _w2658_ ;
	assign \g56897/_0_  = _w2664_ ;
	assign \g56898/_0_  = _w2669_ ;
	assign \g56899/_0_  = _w2675_ ;
	assign \g56900/_0_  = _w2680_ ;
	assign \g56901/_0_  = _w2686_ ;
	assign \g56902/_0_  = _w2691_ ;
	assign \g56903/_0_  = _w2696_ ;
	assign \g56905/_0_  = _w2701_ ;
	assign \g56921/_0_  = _w2702_ ;
	assign \g56956/_0_  = _w2707_ ;
	assign \g56957/_0_  = _w2712_ ;
	assign \g56958/_0_  = _w2718_ ;
	assign \g56959/_0_  = _w2723_ ;
	assign \g56960/_0_  = _w2727_ ;
	assign \g56961/_0_  = _w2732_ ;
	assign \g56962/_0_  = _w2737_ ;
	assign \g56964/_0_  = _w2742_ ;
	assign \g56980/_0_  = _w2743_ ;
	assign \g57015/_0_  = _w2748_ ;
	assign \g57016/_0_  = _w2753_ ;
	assign \g57017/_0_  = _w2758_ ;
	assign \g57018/_0_  = _w2763_ ;
	assign \g57019/_0_  = _w2769_ ;
	assign \g57020/_0_  = _w2774_ ;
	assign \g57021/_0_  = _w2779_ ;
	assign \g57023/_0_  = _w2784_ ;
	assign \g57040/_0_  = _w2785_ ;
	assign \g57074/_0_  = _w2790_ ;
	assign \g57075/_0_  = _w2793_ ;
	assign \g57076/_0_  = _w2798_ ;
	assign \g57077/_0_  = _w2803_ ;
	assign \g57078/_0_  = _w2809_ ;
	assign \g57079/_0_  = _w2814_ ;
	assign \g57080/_0_  = _w2819_ ;
	assign \g57081/_0_  = _w2825_ ;
	assign \g57099/_0_  = _w2826_ ;
	assign \g57133/_0_  = _w2829_ ;
	assign \g57134/_0_  = _w2832_ ;
	assign \g57135/_0_  = _w2837_ ;
	assign \g57136/_0_  = _w2842_ ;
	assign \g57137/_0_  = _w2848_ ;
	assign \g57138/_0_  = _w2853_ ;
	assign \g57139/_0_  = _w2858_ ;
	assign \g57140/_0_  = _w2864_ ;
	assign \g57141/_0_  = _w2869_ ;
	assign \g57159/_0_  = _w2870_ ;
	assign \g57193/_0_  = _w2875_ ;
	assign \g57195/_0_  = _w2880_ ;
	assign \g57196/_0_  = _w2885_ ;
	assign \g57197/_0_  = _w2889_ ;
	assign \g57198/_0_  = _w2894_ ;
	assign \g57199/_0_  = _w2899_ ;
	assign \g57200/_0_  = _w2904_ ;
	assign \g57202/_0_  = _w2909_ ;
	assign \g57219/_0_  = _w2910_ ;
	assign \g57254/_0_  = _w2915_ ;
	assign \g57255/_0_  = _w2920_ ;
	assign \g57256/_0_  = _w2923_ ;
	assign \g57257/_0_  = _w2928_ ;
	assign \g57258/_0_  = _w2933_ ;
	assign \g57259/_0_  = _w2937_ ;
	assign \g57260/_0_  = _w2942_ ;
	assign \g57262/_0_  = _w2948_ ;
	assign \g57263/_0_  = _w2953_ ;
	assign \g57285/_0_  = _w2954_ ;
	assign \g57318/_0_  = _w2959_ ;
	assign \g57319/_0_  = _w2964_ ;
	assign \g57320/_0_  = _w2967_ ;
	assign \g57321/_0_  = _w2970_ ;
	assign \g57322/_0_  = _w2975_ ;
	assign \g57323/_0_  = _w2980_ ;
	assign \g57324/_0_  = _w2986_ ;
	assign \g57325/_0_  = _w2991_ ;
	assign \g57326/_0_  = _w2997_ ;
	assign \g57328/_0_  = _w3003_ ;
	assign \g57329/_0_  = _w3008_ ;
	assign \g57330/_0_  = _w3013_ ;
	assign \g57350/_0_  = _w3014_ ;
	assign \g57387/_0_  = _w3019_ ;
	assign \g57388/_0_  = _w3024_ ;
	assign \g57390/_0_  = _w3027_ ;
	assign \g57391/_0_  = _w3032_ ;
	assign \g57392/_0_  = _w3037_ ;
	assign \g57393/_0_  = _w3041_ ;
	assign \g57395/_0_  = _w3046_ ;
	assign \g57396/_0_  = _w3051_ ;
	assign \g57439/_0_  = _w3052_ ;
	assign \g57476/_0_  = _w3057_ ;
	assign \g57477/_0_  = _w3062_ ;
	assign \g57478/_0_  = _w3067_ ;
	assign \g57479/_0_  = _w3070_ ;
	assign \g57480/_0_  = _w3075_ ;
	assign \g57481/_0_  = _w3082_ ;
	assign \g57482/_0_  = _w3089_ ;
	assign \g57483/_0_  = _w3094_ ;
	assign \g57484/_0_  = _w3097_ ;
	assign \g57485/_0_  = _w3100_ ;
	assign \g57486/_0_  = _w3103_ ;
	assign \g57487/_0_  = _w3106_ ;
	assign \g57488/_0_  = _w3111_ ;
	assign \g57489/_0_  = _w3116_ ;
	assign \g57490/_0_  = _w3121_ ;
	assign \g57491/_0_  = _w3124_ ;
	assign \g57492/_0_  = _w3129_ ;
	assign \g57493/_0_  = _w3134_ ;
	assign \g57494/_0_  = _w3139_ ;
	assign \g57495/_0_  = _w3142_ ;
	assign \g57496/_0_  = _w3146_ ;
	assign \g57497/_0_  = _w3152_ ;
	assign \g57498/_0_  = _w3156_ ;
	assign \g57499/_0_  = _w3159_ ;
	assign \g57500/_0_  = _w3162_ ;
	assign \g57501/_0_  = _w3165_ ;
	assign \g57502/_0_  = _w3168_ ;
	assign \g57503/_0_  = _w3173_ ;
	assign \g57504/_0_  = _w3178_ ;
	assign \g57505/_0_  = _w3183_ ;
	assign \g57524/_0_  = _w3184_ ;
	assign \g57537/_0_  = _w3185_ ;
	assign \g57541/_0_  = _w3186_ ;
	assign \g57543/_0_  = _w3187_ ;
	assign \g58163/_0_  = _w3188_ ;
	assign \g58572/_0_  = _w3189_ ;
	assign \g58573/_0_  = _w3190_ ;
	assign \g58574/_0_  = _w3191_ ;
	assign \g58575/_0_  = _w3192_ ;
	assign \g58576/_0_  = _w3193_ ;
	assign \g58577/_0_  = _w3194_ ;
	assign \g58578/_0_  = _w3195_ ;
	assign \g58579/_0_  = _w3196_ ;
	assign \g58580/_0_  = _w3197_ ;
	assign \g58581/_0_  = _w3198_ ;
	assign \g58582/_0_  = _w3199_ ;
	assign \g58583/_0_  = _w3200_ ;
	assign \g58584/_0_  = _w3201_ ;
	assign \g58585/_0_  = _w3202_ ;
	assign \g58586/_0_  = _w3203_ ;
	assign \g58587/_0_  = _w3204_ ;
	assign \g58588/_0_  = _w3205_ ;
	assign \g58589/_0_  = _w3206_ ;
	assign \g58590/_0_  = _w3207_ ;
	assign \g58591/_0_  = _w3208_ ;
	assign \g58592/_0_  = _w3209_ ;
	assign \g58593/_0_  = _w3210_ ;
	assign \g58594/_0_  = _w3211_ ;
	assign \g58595/_0_  = _w3212_ ;
	assign \g58596/_0_  = _w3213_ ;
	assign \g58597/_0_  = _w3214_ ;
	assign \g58598/_0_  = _w3215_ ;
	assign \g58600/_0_  = _w3216_ ;
	assign \g58602/_0_  = _w3217_ ;
	assign \g58604/_0_  = _w3218_ ;
	assign \g58615/_0_  = _w3219_ ;
	assign \g59240/_0_  = _w3220_ ;
	assign \g59241/_0_  = _w3221_ ;
	assign \g59242/_0_  = _w3222_ ;
	assign \g59243/_0_  = _w3223_ ;
	assign \g59244/_0_  = _w3224_ ;
	assign \g59245/_0_  = _w3225_ ;
	assign \g59246/_0_  = _w3226_ ;
	assign \g59247/_0_  = _w3227_ ;
	assign \g59248/_0_  = _w3228_ ;
	assign \g59249/_0_  = _w3229_ ;
	assign \g59250/_0_  = _w3230_ ;
	assign \g59251/_0_  = _w3231_ ;
	assign \g59252/_0_  = _w3232_ ;
	assign \g59253/_0_  = _w3233_ ;
	assign \g59254/_0_  = _w3234_ ;
	assign \g59255/_0_  = _w3235_ ;
	assign \g59256/_0_  = _w3236_ ;
	assign \g59257/_0_  = _w3237_ ;
	assign \g59258/_0_  = _w3238_ ;
	assign \g59259/_0_  = _w3239_ ;
	assign \g59260/_0_  = _w3240_ ;
	assign \g59261/_0_  = _w3241_ ;
	assign \g59262/_0_  = _w3242_ ;
	assign \g59263/_0_  = _w3243_ ;
	assign \g59264/_0_  = _w3244_ ;
	assign \g59265/_0_  = _w3245_ ;
	assign \g59266/_0_  = _w3246_ ;
	assign \g59267/_0_  = _w3247_ ;
	assign \g59268/_0_  = _w3248_ ;
	assign \g59269/_0_  = _w3249_ ;
	assign \g59270/_0_  = _w3250_ ;
	assign \g59271/_0_  = _w3251_ ;
	assign \g59272/_0_  = _w3252_ ;
	assign \g59273/_0_  = _w3253_ ;
	assign \g59274/_0_  = _w3254_ ;
	assign \g59275/_0_  = _w3255_ ;
	assign \g59276/_0_  = _w3256_ ;
	assign \g59277/_0_  = _w3257_ ;
	assign \g59278/_0_  = _w3258_ ;
	assign \g59279/_0_  = _w3259_ ;
	assign \g59280/_0_  = _w3260_ ;
	assign \g59281/_0_  = _w3261_ ;
	assign \g59282/_0_  = _w3262_ ;
	assign \g59283/_0_  = _w3263_ ;
	assign \g59284/_0_  = _w3264_ ;
	assign \g59285/_0_  = _w3265_ ;
	assign \g59286/_0_  = _w3266_ ;
	assign \g59287/_0_  = _w3267_ ;
	assign \g59288/_0_  = _w3268_ ;
	assign \g59289/_0_  = _w3269_ ;
	assign \g59290/_0_  = _w3270_ ;
	assign \g59291/_0_  = _w3271_ ;
	assign \g59292/_0_  = _w3272_ ;
	assign \g59293/_0_  = _w3273_ ;
	assign \g59294/_0_  = _w3274_ ;
	assign \g59295/_0_  = _w3275_ ;
	assign \g59296/_0_  = _w3276_ ;
	assign \g59297/_0_  = _w3277_ ;
	assign \g59298/_0_  = _w3278_ ;
	assign \g59299/_0_  = _w3279_ ;
	assign \g59300/_0_  = _w3280_ ;
	assign \g59301/_0_  = _w3281_ ;
	assign \g59302/_0_  = _w3282_ ;
	assign \g59303/_0_  = _w3283_ ;
	assign \g59304/_0_  = _w3284_ ;
	assign \g59305/_0_  = _w3285_ ;
	assign \g59306/_0_  = _w3286_ ;
	assign \g59307/_0_  = _w3287_ ;
	assign \g59308/_0_  = _w3288_ ;
	assign \g59309/_0_  = _w3289_ ;
	assign \g59310/_0_  = _w3290_ ;
	assign \g59311/_0_  = _w3291_ ;
	assign \g59312/_0_  = _w3292_ ;
	assign \g59313/_0_  = _w3293_ ;
	assign \g59314/_0_  = _w3294_ ;
	assign \g59315/_0_  = _w3295_ ;
	assign \g59316/_0_  = _w3296_ ;
	assign \g59317/_0_  = _w3297_ ;
	assign \g59318/_0_  = _w3298_ ;
	assign \g59319/_0_  = _w3299_ ;
	assign \g59320/_0_  = _w3300_ ;
	assign \g59321/_0_  = _w3301_ ;
	assign \g59322/_0_  = _w3302_ ;
	assign \g59323/_0_  = _w3303_ ;
	assign \g59324/_0_  = _w3304_ ;
	assign \g59325/_0_  = _w3305_ ;
	assign \g59326/_0_  = _w3306_ ;
	assign \g59327/_0_  = _w3307_ ;
	assign \g59328/_0_  = _w3308_ ;
	assign \g59329/_0_  = _w3309_ ;
	assign \g59330/_0_  = _w3310_ ;
	assign \g59331/_0_  = _w3311_ ;
	assign \g59332/_0_  = _w3312_ ;
	assign \g59333/_0_  = _w3313_ ;
	assign \g59334/_0_  = _w3314_ ;
	assign \g59335/_0_  = _w3315_ ;
	assign \g59336/_0_  = _w3316_ ;
	assign \g59337/_0_  = _w3317_ ;
	assign \g59338/_0_  = _w3318_ ;
	assign \g59339/_0_  = _w3319_ ;
	assign \g59340/_0_  = _w3320_ ;
	assign \g59341/_0_  = _w3321_ ;
	assign \g59342/_0_  = _w3322_ ;
	assign \g59343/_0_  = _w3323_ ;
	assign \g59344/_0_  = _w3324_ ;
	assign \g59345/_0_  = _w3325_ ;
	assign \g59346/_0_  = _w3326_ ;
	assign \g59347/_0_  = _w3327_ ;
	assign \g59348/_0_  = _w3328_ ;
	assign \g59349/_0_  = _w3329_ ;
	assign \g59350/_0_  = _w3330_ ;
	assign \g59351/_0_  = _w3331_ ;
	assign \g59352/_0_  = _w3332_ ;
	assign \g59353/_0_  = _w3333_ ;
	assign \g59354/_0_  = _w3334_ ;
	assign \g59355/_0_  = _w3335_ ;
	assign \g59356/_0_  = _w3336_ ;
	assign \g59357/_0_  = _w3337_ ;
	assign \g59358/_0_  = _w3338_ ;
	assign \g59359/_0_  = _w3339_ ;
	assign \g59360/_0_  = _w3340_ ;
	assign \g59361/_0_  = _w3341_ ;
	assign \g59362/_0_  = _w3342_ ;
	assign \g59363/_0_  = _w3343_ ;
	assign \g59364/_0_  = _w3344_ ;
	assign \g59365/_0_  = _w3345_ ;
	assign \g59366/_0_  = _w3346_ ;
	assign \g59367/_0_  = _w3347_ ;
	assign \g59368/_0_  = _w3348_ ;
	assign \g59369/_0_  = _w3349_ ;
	assign \g59370/_0_  = _w3350_ ;
	assign \g59371/_0_  = _w3351_ ;
	assign \g59372/_0_  = _w3352_ ;
	assign \g59373/_0_  = _w3353_ ;
	assign \g59374/_0_  = _w3354_ ;
	assign \g59375/_0_  = _w3355_ ;
	assign \g59376/_0_  = _w3356_ ;
	assign \g59377/_0_  = _w3357_ ;
	assign \g59378/_0_  = _w3358_ ;
	assign \g59379/_0_  = _w3359_ ;
	assign \g59380/_0_  = _w3360_ ;
	assign \g59381/_0_  = _w3361_ ;
	assign \g59382/_0_  = _w3362_ ;
	assign \g59383/_0_  = _w3363_ ;
	assign \g59384/_0_  = _w3364_ ;
	assign \g59385/_0_  = _w3365_ ;
	assign \g59386/_0_  = _w3366_ ;
	assign \g59387/_0_  = _w3367_ ;
	assign \g59388/_0_  = _w3368_ ;
	assign \g59389/_0_  = _w3369_ ;
	assign \g59390/_0_  = _w3370_ ;
	assign \g59391/_0_  = _w3371_ ;
	assign \g59392/_0_  = _w3372_ ;
	assign \g59393/_0_  = _w3373_ ;
	assign \g59394/_0_  = _w3374_ ;
	assign \g59395/_0_  = _w3375_ ;
	assign \g59396/_0_  = _w3376_ ;
	assign \g59397/_0_  = _w3377_ ;
	assign \g59398/_0_  = _w3378_ ;
	assign \g59399/_0_  = _w3379_ ;
	assign \g59400/_0_  = _w3380_ ;
	assign \g59401/_0_  = _w3381_ ;
	assign \g59402/_0_  = _w3382_ ;
	assign \g59403/_0_  = _w3383_ ;
	assign \g59404/_0_  = _w3384_ ;
	assign \g59405/_0_  = _w3385_ ;
	assign \g59406/_0_  = _w3386_ ;
	assign \g59407/_0_  = _w3387_ ;
	assign \g59408/_0_  = _w3388_ ;
	assign \g59409/_0_  = _w3389_ ;
	assign \g59410/_0_  = _w3390_ ;
	assign \g59411/_0_  = _w3391_ ;
	assign \g59412/_0_  = _w3392_ ;
	assign \g59413/_0_  = _w3393_ ;
	assign \g59414/_0_  = _w3394_ ;
	assign \g59415/_0_  = _w3395_ ;
	assign \g59416/_0_  = _w3396_ ;
	assign \g59417/_0_  = _w3397_ ;
	assign \g59418/_0_  = _w3398_ ;
	assign \g59419/_0_  = _w3399_ ;
	assign \g59420/_0_  = _w3400_ ;
	assign \g59421/_0_  = _w3401_ ;
	assign \g59422/_0_  = _w3402_ ;
	assign \g59423/_0_  = _w3403_ ;
	assign \g59424/_0_  = _w3404_ ;
	assign \g59425/_0_  = _w3405_ ;
	assign \g59426/_0_  = _w3406_ ;
	assign \g59427/_0_  = _w3407_ ;
	assign \g59428/_0_  = _w3408_ ;
	assign \g59429/_0_  = _w3409_ ;
	assign \g59430/_0_  = _w3410_ ;
	assign \g59431/_0_  = _w3411_ ;
	assign \g59432/_0_  = _w3412_ ;
	assign \g59433/_0_  = _w3413_ ;
	assign \g59434/_0_  = _w3414_ ;
	assign \g59435/_0_  = _w3415_ ;
	assign \g59436/_0_  = _w3416_ ;
	assign \g59437/_0_  = _w3417_ ;
	assign \g59438/_0_  = _w3418_ ;
	assign \g59439/_0_  = _w3419_ ;
	assign \g59440/_0_  = _w3420_ ;
	assign \g59441/_0_  = _w3421_ ;
	assign \g59442/_0_  = _w3422_ ;
	assign \g59443/_0_  = _w3423_ ;
	assign \g59444/_0_  = _w3424_ ;
	assign \g59445/_0_  = _w3425_ ;
	assign \g59446/_0_  = _w3426_ ;
	assign \g59447/_0_  = _w3427_ ;
	assign \g59448/_0_  = _w3428_ ;
	assign \g59449/_0_  = _w3429_ ;
	assign \g59450/_0_  = _w3430_ ;
	assign \g59451/_0_  = _w3431_ ;
	assign \g59452/_0_  = _w3432_ ;
	assign \g59453/_0_  = _w3433_ ;
	assign \g59454/_0_  = _w3434_ ;
	assign \g59455/_0_  = _w3435_ ;
	assign \g59456/_0_  = _w3436_ ;
	assign \g59457/_0_  = _w3437_ ;
	assign \g59458/_0_  = _w3438_ ;
	assign \g59459/_0_  = _w3439_ ;
	assign \g59460/_0_  = _w3440_ ;
	assign \g59461/_0_  = _w3441_ ;
	assign \g59462/_0_  = _w3442_ ;
	assign \g59463/_0_  = _w3443_ ;
	assign \g59464/_0_  = _w3444_ ;
	assign \g59465/_0_  = _w3445_ ;
	assign \g59466/_0_  = _w3446_ ;
	assign \g59467/_0_  = _w3447_ ;
	assign \g59468/_0_  = _w3448_ ;
	assign \g59469/_0_  = _w3449_ ;
	assign \g59470/_0_  = _w3450_ ;
	assign \g59471/_0_  = _w3451_ ;
	assign \g59472/_0_  = _w3452_ ;
	assign \g59473/_0_  = _w3453_ ;
	assign \g59474/_0_  = _w3454_ ;
	assign \g59475/_0_  = _w3455_ ;
	assign \g59476/_0_  = _w3456_ ;
	assign \g59477/_0_  = _w3457_ ;
	assign \g59478/_0_  = _w3458_ ;
	assign \g59479/_0_  = _w3459_ ;
	assign \g59480/_0_  = _w3460_ ;
	assign \g59481/_0_  = _w3461_ ;
	assign \g59482/_0_  = _w3462_ ;
	assign \g59483/_0_  = _w3463_ ;
	assign \g59484/_0_  = _w3464_ ;
	assign \g59485/_0_  = _w3465_ ;
	assign \g59486/_0_  = _w3466_ ;
	assign \g59487/_0_  = _w3467_ ;
	assign \g59488/_0_  = _w3468_ ;
	assign \g59489/_0_  = _w3469_ ;
	assign \g59490/_0_  = _w3470_ ;
	assign \g59491/_0_  = _w3471_ ;
	assign \g59492/_0_  = _w3472_ ;
	assign \g59493/_0_  = _w3473_ ;
	assign \g59494/_0_  = _w3474_ ;
	assign \g59495/_0_  = _w3475_ ;
	assign \g59496/_0_  = _w3476_ ;
	assign \g59497/_0_  = _w3477_ ;
	assign \g59498/_0_  = _w3478_ ;
	assign \g59500/_0_  = _w3479_ ;
	assign \g59503/_0_  = _w3480_ ;
	assign \g59512/_0_  = _w3481_ ;
	assign \g61336/_0_  = _w3482_ ;
	assign \g61521/_0_  = _w3483_ ;
	assign \g61523/_0_  = _w3484_ ;
	assign \g61524/_0_  = _w3485_ ;
	assign \g61526/_0_  = _w3486_ ;
	assign \g61527/_0_  = _w3487_ ;
	assign \g61528/_0_  = _w3488_ ;
	assign \g61529/_0_  = _w3489_ ;
	assign \g61530/_0_  = _w3490_ ;
	assign \g61531/_0_  = _w3491_ ;
	assign \g61532/_0_  = _w3492_ ;
	assign \g61533/_0_  = _w3493_ ;
	assign \g61535/_0_  = _w3494_ ;
	assign \g61537/_0_  = _w3495_ ;
	assign \g61539/_0_  = _w3496_ ;
	assign \g61540/_0_  = _w3497_ ;
	assign \g61541/_0_  = _w3498_ ;
	assign \g61542/_0_  = _w3499_ ;
	assign \g61546/_0_  = _w3500_ ;
	assign \g61550/_0_  = _w3501_ ;
	assign \g61551/_0_  = _w3502_ ;
	assign \g61552/_0_  = _w3503_ ;
	assign \g61554/_0_  = _w3504_ ;
	assign \g61555/_0_  = _w3505_ ;
	assign \g61556/_0_  = _w3506_ ;
	assign \g61558/_0_  = _w3507_ ;
	assign \g61559/_0_  = _w3508_ ;
	assign \g61561/_0_  = _w3509_ ;
	assign \g61562/_0_  = _w3510_ ;
	assign \g61563/_0_  = _w3511_ ;
	assign \g61564/_0_  = _w3512_ ;
	assign \g61565/_0_  = _w3513_ ;
	assign \g61566/_0_  = _w3514_ ;
	assign \g61568/_0_  = _w3515_ ;
	assign \g61570/_0_  = _w3516_ ;
	assign \g61571/_0_  = _w3517_ ;
	assign \g61572/_0_  = _w3518_ ;
	assign \g61573/_0_  = _w3519_ ;
	assign \g61577/_0_  = _w3520_ ;
	assign \g61578/_0_  = _w3521_ ;
	assign \g61579/_0_  = _w3522_ ;
	assign \g61580/_0_  = _w3523_ ;
	assign \g61581/_0_  = _w3524_ ;
	assign \g61582/_0_  = _w3525_ ;
	assign \g61583/_0_  = _w3526_ ;
	assign \g61584/_0_  = _w3527_ ;
	assign \g61585/_0_  = _w3528_ ;
	assign \g61586/_0_  = _w3529_ ;
	assign \g61587/_0_  = _w3530_ ;
	assign \g61588/_0_  = _w3531_ ;
	assign \g61589/_0_  = _w3532_ ;
	assign \g61591/_0_  = _w3533_ ;
	assign \g61592/_0_  = _w3534_ ;
	assign \g61594/_0_  = _w3535_ ;
	assign \g61595/_0_  = _w3536_ ;
	assign \g61596/_0_  = _w3537_ ;
	assign \g61597/_0_  = _w3538_ ;
	assign \g61598/_0_  = _w3539_ ;
	assign \g61599/_0_  = _w3540_ ;
	assign \g61600/_0_  = _w3541_ ;
	assign \g61601/_0_  = _w3542_ ;
	assign \g61605/_0_  = _w3543_ ;
	assign \g61606/_0_  = _w3544_ ;
	assign \g61607/_0_  = _w3545_ ;
	assign \g61608/_0_  = _w3546_ ;
	assign \g61609/_0_  = _w3547_ ;
	assign \g61610/_0_  = _w3548_ ;
	assign \g61611/_0_  = _w3549_ ;
	assign \g61612/_0_  = _w3550_ ;
	assign \g61613/_0_  = _w3551_ ;
	assign \g61615/_0_  = _w3552_ ;
	assign \g61616/_0_  = _w3553_ ;
	assign \g61617/_0_  = _w3554_ ;
	assign \g61618/_0_  = _w3555_ ;
	assign \g61619/_0_  = _w3556_ ;
	assign \g61620/_0_  = _w3557_ ;
	assign \g61621/_0_  = _w3558_ ;
	assign \g61623/_0_  = _w3559_ ;
	assign \g61624/_0_  = _w3560_ ;
	assign \g61625/_0_  = _w3561_ ;
	assign \g61626/_0_  = _w3562_ ;
	assign \g61627/_0_  = _w3563_ ;
	assign \g61629/_0_  = _w3564_ ;
	assign \g61630/_0_  = _w3565_ ;
	assign \g61631/_0_  = _w3566_ ;
	assign \g61632/_0_  = _w3567_ ;
	assign \g61633/_0_  = _w3568_ ;
	assign \g61634/_0_  = _w3569_ ;
	assign \g61636/_0_  = _w3570_ ;
	assign \g61638/_0_  = _w3571_ ;
	assign \g61639/_0_  = _w3572_ ;
	assign \g61640/_0_  = _w3573_ ;
	assign \g61641/_0_  = _w3574_ ;
	assign \g61642/_0_  = _w3575_ ;
	assign \g61644/_0_  = _w3576_ ;
	assign \g61647/_0_  = _w3577_ ;
	assign \g61648/_0_  = _w3578_ ;
	assign \g61649/_0_  = _w3579_ ;
	assign \g61650/_0_  = _w3580_ ;
	assign \g61653/_0_  = _w3581_ ;
	assign \g61654/_0_  = _w3582_ ;
	assign \g61655/_0_  = _w3583_ ;
	assign \g61656/_0_  = _w3584_ ;
	assign \g61658/_0_  = _w3585_ ;
	assign \g61661/_0_  = _w3586_ ;
	assign \g61662/_0_  = _w3587_ ;
	assign \g61663/_0_  = _w3588_ ;
	assign \g61664/_0_  = _w3589_ ;
	assign \g61666/_0_  = _w3590_ ;
	assign \g61667/_0_  = _w3591_ ;
	assign \g61668/_0_  = _w3592_ ;
	assign \g61670/_0_  = _w3593_ ;
	assign \g61671/_0_  = _w3594_ ;
	assign \g61672/_0_  = _w3595_ ;
	assign \g61673/_0_  = _w3596_ ;
	assign \g61675/_0_  = _w3597_ ;
	assign \g61676/_0_  = _w3598_ ;
	assign \g61680/_0_  = _w3599_ ;
	assign \g61681/_0_  = _w3600_ ;
	assign \g61682/_0_  = _w3601_ ;
	assign \g61683/_0_  = _w3602_ ;
	assign \g61684/_0_  = _w3603_ ;
	assign \g61686/_0_  = _w3604_ ;
	assign \g61687/_0_  = _w3605_ ;
	assign \g61688/_0_  = _w3606_ ;
	assign \g61689/_0_  = _w3607_ ;
	assign \g61690/_0_  = _w3608_ ;
	assign \g61691/_0_  = _w3609_ ;
	assign \g61693/_0_  = _w3610_ ;
	assign \g61694/_0_  = _w3611_ ;
	assign \g61696/_0_  = _w3612_ ;
	assign \g61697/_0_  = _w3613_ ;
	assign \g61698/_0_  = _w3614_ ;
	assign \g61699/_0_  = _w3615_ ;
	assign \g61700/_0_  = _w3616_ ;
	assign \g61701/_0_  = _w3617_ ;
	assign \g61702/_0_  = _w3618_ ;
	assign \g61703/_0_  = _w3619_ ;
	assign \g61704/_0_  = _w3620_ ;
	assign \g61705/_0_  = _w3621_ ;
	assign \g61706/_0_  = _w3622_ ;
	assign \g61707/_0_  = _w3623_ ;
	assign \g61708/_0_  = _w3624_ ;
	assign \g61711/_0_  = _w3625_ ;
	assign \g61712/_0_  = _w3626_ ;
	assign \g61714/_0_  = _w3627_ ;
	assign \g61716/_0_  = _w3628_ ;
	assign \g61717/_0_  = _w3629_ ;
	assign \g61719/_0_  = _w3630_ ;
	assign \g61720/_0_  = _w3631_ ;
	assign \g61721/_0_  = _w3632_ ;
	assign \g61724/_0_  = _w3633_ ;
	assign \g61725/_0_  = _w3634_ ;
	assign \g61728/_0_  = _w3635_ ;
	assign \g61729/_0_  = _w3636_ ;
	assign \g61731/_0_  = _w3637_ ;
	assign \g61732/_0_  = _w3638_ ;
	assign \g61733/_0_  = _w3639_ ;
	assign \g61736/_0_  = _w3640_ ;
	assign \g61737/_0_  = _w3641_ ;
	assign \g61739/_0_  = _w3642_ ;
	assign \g61740/_0_  = _w3643_ ;
	assign \g61741/_0_  = _w3644_ ;
	assign \g61743/_0_  = _w3645_ ;
	assign \g61744/_0_  = _w3646_ ;
	assign \g61745/_0_  = _w3647_ ;
	assign \g61746/_0_  = _w3648_ ;
	assign \g61747/_0_  = _w3649_ ;
	assign \g61748/_0_  = _w3650_ ;
	assign \g61749/_0_  = _w3651_ ;
	assign \g61750/_0_  = _w3652_ ;
	assign \g61751/_0_  = _w3653_ ;
	assign \g61752/_0_  = _w3654_ ;
	assign \g61753/_0_  = _w3655_ ;
	assign \g61754/_0_  = _w3656_ ;
	assign \g61755/_0_  = _w3657_ ;
	assign \g61757/_0_  = _w3658_ ;
	assign \g61758/_0_  = _w3659_ ;
	assign \g61759/_0_  = _w3660_ ;
	assign \g61760/_0_  = _w3661_ ;
	assign \g61761/_0_  = _w3662_ ;
	assign \g61762/_0_  = _w3663_ ;
	assign \g61763/_0_  = _w3664_ ;
	assign \g61764/_0_  = _w3665_ ;
	assign \g61765/_0_  = _w3666_ ;
	assign \g61766/_0_  = _w3667_ ;
	assign \g61767/_0_  = _w3668_ ;
	assign \g61768/_0_  = _w3669_ ;
	assign \g61769/_0_  = _w3670_ ;
	assign \g61770/_0_  = _w3671_ ;
	assign \g61771/_0_  = _w3672_ ;
	assign \g61772/_0_  = _w3673_ ;
	assign \g61773/_0_  = _w3674_ ;
	assign \g61774/_0_  = _w3675_ ;
	assign \g61775/_0_  = _w3676_ ;
	assign \g61776/_0_  = _w3677_ ;
	assign \g61777/_0_  = _w3678_ ;
	assign \g61778/_0_  = _w3679_ ;
	assign \g61780/_0_  = _w3680_ ;
	assign \g61781/_0_  = _w3681_ ;
	assign \g61783/_0_  = _w3682_ ;
	assign \g61784/_0_  = _w3683_ ;
	assign \g61786/_0_  = _w3684_ ;
	assign \g61787/_0_  = _w3685_ ;
	assign \g61790/_0_  = _w3686_ ;
	assign \g61791/_0_  = _w3687_ ;
	assign \g61794/_0_  = _w3688_ ;
	assign \g61795/_0_  = _w3689_ ;
	assign \g61796/_0_  = _w3690_ ;
	assign \g61797/_0_  = _w3691_ ;
	assign \g61798/_0_  = _w3692_ ;
	assign \g61799/_0_  = _w3693_ ;
	assign \g61800/_0_  = _w3694_ ;
	assign \g61801/_0_  = _w3695_ ;
	assign \g61802/_0_  = _w3696_ ;
	assign \g61803/_0_  = _w3697_ ;
	assign \g61805/_0_  = _w3698_ ;
	assign \g61806/_0_  = _w3699_ ;
	assign \g61807/_0_  = _w3700_ ;
	assign \g61808/_0_  = _w3701_ ;
	assign \g61809/_0_  = _w3702_ ;
	assign \g61810/_0_  = _w3703_ ;
	assign \g61811/_0_  = _w3704_ ;
	assign \g61812/_0_  = _w3705_ ;
	assign \g61813/_0_  = _w3706_ ;
	assign \g61816/_0_  = _w3707_ ;
	assign \g61817/_0_  = _w3708_ ;
	assign \g61818/_0_  = _w3709_ ;
	assign \g61820/_0_  = _w3710_ ;
	assign \g61822/_0_  = _w3711_ ;
	assign \g61823/_0_  = _w3712_ ;
	assign \g61825/_0_  = _w3713_ ;
	assign \g61826/_0_  = _w3714_ ;
	assign \g61827/_0_  = _w3715_ ;
	assign \g61828/_0_  = _w3716_ ;
	assign \g61829/_0_  = _w3717_ ;
	assign \g61832/_0_  = _w3718_ ;
	assign \g61834/_0_  = _w3719_ ;
	assign \g61835/_0_  = _w3720_ ;
	assign \g61837/_0_  = _w3721_ ;
	assign \g61838/_0_  = _w3722_ ;
	assign \g61839/_0_  = _w3723_ ;
	assign \g61840/_0_  = _w3724_ ;
	assign \g61844/_0_  = _w3725_ ;
	assign \g61847/_0_  = _w3726_ ;
	assign \g61848/_0_  = _w3727_ ;
	assign \g61849/_0_  = _w3728_ ;
	assign \g61850/_0_  = _w3729_ ;
	assign \g61851/_0_  = _w3730_ ;
	assign \g61853/_0_  = _w3731_ ;
	assign \g61854/_0_  = _w3732_ ;
	assign \g61855/_0_  = _w3733_ ;
	assign \g61856/_0_  = _w3734_ ;
	assign \g61858/_0_  = _w3735_ ;
	assign \g61859/_0_  = _w3736_ ;
	assign \g61861/_0_  = _w3737_ ;
	assign \g61862/_0_  = _w3738_ ;
	assign \g61863/_0_  = _w3739_ ;
	assign \g61864/_0_  = _w3740_ ;
	assign \g61865/_0_  = _w3741_ ;
	assign \g61866/_0_  = _w3742_ ;
	assign \g61867/_0_  = _w3743_ ;
	assign \g61868/_0_  = _w3744_ ;
	assign \g61869/_0_  = _w3745_ ;
	assign \g61870/_0_  = _w3746_ ;
	assign \g61871/_0_  = _w3747_ ;
	assign \g61873/_0_  = _w3748_ ;
	assign \g61874/_0_  = _w3749_ ;
	assign \g61875/_0_  = _w3750_ ;
	assign \g61877/_0_  = _w3751_ ;
	assign \g61878/_0_  = _w3752_ ;
	assign \g61879/_0_  = _w3753_ ;
	assign \g61880/_0_  = _w3754_ ;
	assign \g61881/_0_  = _w3755_ ;
	assign \g61883/_0_  = _w3756_ ;
	assign \g61884/_0_  = _w3757_ ;
	assign \g61886/_0_  = _w3758_ ;
	assign \g61887/_0_  = _w3759_ ;
	assign \g61890/_0_  = _w3760_ ;
	assign \g61891/_0_  = _w3761_ ;
	assign \g61892/_0_  = _w3762_ ;
	assign \g61893/_0_  = _w3763_ ;
	assign \g61894/_0_  = _w3764_ ;
	assign \g61895/_0_  = _w3765_ ;
	assign \g61900/_0_  = _w3766_ ;
	assign \g61901/_0_  = _w3767_ ;
	assign \g61902/_0_  = _w3768_ ;
	assign \g61904/_0_  = _w3769_ ;
	assign \g61905/_0_  = _w3770_ ;
	assign \g61906/_0_  = _w3771_ ;
	assign \g61907/_0_  = _w3772_ ;
	assign \g61914/_0_  = _w3773_ ;
	assign \g61915/_0_  = _w3774_ ;
	assign \g61917/_0_  = _w3775_ ;
	assign \g61919/_0_  = _w3776_ ;
	assign \g61921/_0_  = _w3777_ ;
	assign \g61924/_0_  = _w3778_ ;
	assign \g61925/_0_  = _w3779_ ;
	assign \g61926/_0_  = _w3780_ ;
	assign \g61927/_0_  = _w3781_ ;
	assign \g61928/_0_  = _w3782_ ;
	assign \g61929/_0_  = _w3783_ ;
	assign \g61930/_0_  = _w3784_ ;
	assign \g61931/_0_  = _w3785_ ;
	assign \g61932/_0_  = _w3786_ ;
	assign \g61933/_0_  = _w3787_ ;
	assign \g61934/_0_  = _w3788_ ;
	assign \g61935/_0_  = _w3789_ ;
	assign \g61936/_0_  = _w3790_ ;
	assign \g61937/_0_  = _w3791_ ;
	assign \g61938/_0_  = _w3792_ ;
	assign \g61939/_0_  = _w3793_ ;
	assign \g61943/_0_  = _w3794_ ;
	assign \g61944/_0_  = _w3795_ ;
	assign \g61945/_0_  = _w3796_ ;
	assign \g61947/_0_  = _w3797_ ;
	assign \g61948/_0_  = _w3798_ ;
	assign \g61949/_0_  = _w3799_ ;
	assign \g61950/_0_  = _w3800_ ;
	assign \g61951/_0_  = _w3801_ ;
	assign \g61952/_0_  = _w3802_ ;
	assign \g61953/_0_  = _w3803_ ;
	assign \g61955/_0_  = _w3804_ ;
	assign \g61956/_0_  = _w3805_ ;
	assign \g61957/_0_  = _w3806_ ;
	assign \g61958/_0_  = _w3807_ ;
	assign \g61959/_0_  = _w3808_ ;
	assign \g61960/_0_  = _w3809_ ;
	assign \g61961/_0_  = _w3810_ ;
	assign \g61962/_0_  = _w3811_ ;
	assign \g61963/_0_  = _w3812_ ;
	assign \g61964/_0_  = _w3813_ ;
	assign \g61965/_0_  = _w3814_ ;
	assign \g61966/_0_  = _w3815_ ;
	assign \g61967/_0_  = _w3816_ ;
	assign \g61968/_0_  = _w3817_ ;
	assign \g61969/_0_  = _w3818_ ;
	assign \g61970/_0_  = _w3819_ ;
	assign \g61971/_0_  = _w3820_ ;
	assign \g61972/_0_  = _w3821_ ;
	assign \g61973/_0_  = _w3822_ ;
	assign \g61974/_0_  = _w3823_ ;
	assign \g61976/_0_  = _w3824_ ;
	assign \g61978/_0_  = _w3825_ ;
	assign \g61980/_0_  = _w3826_ ;
	assign \g61981/_0_  = _w3827_ ;
	assign \g61982/_0_  = _w3828_ ;
	assign \g61983/_0_  = _w3829_ ;
	assign \g61984/_0_  = _w3830_ ;
	assign \g61985/_0_  = _w3831_ ;
	assign \g61986/_0_  = _w3832_ ;
	assign \g61987/_0_  = _w3833_ ;
	assign \g61988/_0_  = _w3834_ ;
	assign \g61989/_0_  = _w3835_ ;
	assign \g61990/_0_  = _w3836_ ;
	assign \g61992/_0_  = _w3837_ ;
	assign \g61994/_0_  = _w3838_ ;
	assign \g61995/_0_  = _w3839_ ;
	assign \g61996/_0_  = _w3840_ ;
	assign \g61997/_0_  = _w3841_ ;
	assign \g61998/_0_  = _w3842_ ;
	assign \g62000/_0_  = _w3843_ ;
	assign \g62001/_0_  = _w3844_ ;
	assign \g62002/_0_  = _w3845_ ;
	assign \g62003/_0_  = _w3846_ ;
	assign \g62004/_0_  = _w3847_ ;
	assign \g62005/_0_  = _w3848_ ;
	assign \g62007/_0_  = _w3849_ ;
	assign \g62008/_0_  = _w3850_ ;
	assign \g62009/_0_  = _w3851_ ;
	assign \g62010/_0_  = _w3852_ ;
	assign \g62011/_0_  = _w3853_ ;
	assign \g62012/_0_  = _w3854_ ;
	assign \g62013/_0_  = _w3855_ ;
	assign \g62014/_0_  = _w3856_ ;
	assign \g62015/_0_  = _w3857_ ;
	assign \g62016/_0_  = _w3858_ ;
	assign \g62017/_0_  = _w3859_ ;
	assign \g62018/_0_  = _w3860_ ;
	assign \g62019/_0_  = _w3861_ ;
	assign \g62020/_0_  = _w3862_ ;
	assign \g62021/_0_  = _w3863_ ;
	assign \g62022/_0_  = _w3864_ ;
	assign \g62023/_0_  = _w3865_ ;
	assign \g62024/_0_  = _w3866_ ;
	assign \g62025/_0_  = _w3867_ ;
	assign \g62026/_0_  = _w3868_ ;
	assign \g62027/_0_  = _w3869_ ;
	assign \g62030/_0_  = _w3870_ ;
	assign \g62033/_0_  = _w3871_ ;
	assign \g62034/_0_  = _w3872_ ;
	assign \g62036/_0_  = _w3873_ ;
	assign \g62038/_0_  = _w3874_ ;
	assign \g62041/_0_  = _w3875_ ;
	assign \g62042/_0_  = _w3876_ ;
	assign \g62043/_0_  = _w3877_ ;
	assign \g62044/_0_  = _w3878_ ;
	assign \g62045/_0_  = _w3879_ ;
	assign \g62046/_0_  = _w3880_ ;
	assign \g62047/_0_  = _w3881_ ;
	assign \g62048/_0_  = _w3882_ ;
	assign \g62050/_0_  = _w3883_ ;
	assign \g62051/_0_  = _w3884_ ;
	assign \g62052/_0_  = _w3885_ ;
	assign \g62055/_0_  = _w3886_ ;
	assign \g62057/_0_  = _w3887_ ;
	assign \g62058/_0_  = _w3888_ ;
	assign \g62059/_0_  = _w3889_ ;
	assign \g62060/_0_  = _w3890_ ;
	assign \g62061/_0_  = _w3891_ ;
	assign \g62062/_0_  = _w3892_ ;
	assign \g62064/_0_  = _w3893_ ;
	assign \g62065/_0_  = _w3894_ ;
	assign \g62066/_0_  = _w3895_ ;
	assign \g62067/_0_  = _w3896_ ;
	assign \g62068/_0_  = _w3897_ ;
	assign \g62072/_0_  = _w3898_ ;
	assign \g62073/_0_  = _w3899_ ;
	assign \g62074/_0_  = _w3900_ ;
	assign \g62075/_0_  = _w3901_ ;
	assign \g62076/_0_  = _w3902_ ;
	assign \g62077/_0_  = _w3903_ ;
	assign \g62078/_0_  = _w3904_ ;
	assign \g62080/_0_  = _w3905_ ;
	assign \g62081/_0_  = _w3906_ ;
	assign \g62082/_0_  = _w3907_ ;
	assign \g62084/_0_  = _w3908_ ;
	assign \g62085/_0_  = _w3909_ ;
	assign \g62086/_0_  = _w3910_ ;
	assign \g62087/_0_  = _w3911_ ;
	assign \g62088/_0_  = _w3912_ ;
	assign \g62089/_0_  = _w3913_ ;
	assign \g62090/_0_  = _w3914_ ;
	assign \g62091/_0_  = _w3915_ ;
	assign \g62092/_0_  = _w3916_ ;
	assign \g62094/_0_  = _w3917_ ;
	assign \g62096/_0_  = _w3918_ ;
	assign \g62097/_0_  = _w3919_ ;
	assign \g62098/_0_  = _w3920_ ;
	assign \g62099/_0_  = _w3921_ ;
	assign \g62100/_0_  = _w3922_ ;
	assign \g62101/_0_  = _w3923_ ;
	assign \g62102/_0_  = _w3924_ ;
	assign \g62104/_0_  = _w3925_ ;
	assign \g62106/_0_  = _w3926_ ;
	assign \g62107/_0_  = _w3927_ ;
	assign \g62108/_0_  = _w3928_ ;
	assign \g62110/_0_  = _w3929_ ;
	assign \g62112/_0_  = _w3930_ ;
	assign \g62113/_0_  = _w3931_ ;
	assign \g62114/_0_  = _w3932_ ;
	assign \g62116/_0_  = _w3933_ ;
	assign \g62117/_0_  = _w3934_ ;
	assign \g62118/_0_  = _w3935_ ;
	assign \g62119/_0_  = _w3936_ ;
	assign \g62120/_0_  = _w3937_ ;
	assign \g62121/_0_  = _w3938_ ;
	assign \g62122/_0_  = _w3939_ ;
	assign \g62124/_0_  = _w3940_ ;
	assign \g62126/_0_  = _w3941_ ;
	assign \g62127/_0_  = _w3942_ ;
	assign \g62128/_0_  = _w3943_ ;
	assign \g62129/_0_  = _w3944_ ;
	assign \g62130/_0_  = _w3945_ ;
	assign \g62131/_0_  = _w3946_ ;
	assign \g62132/_0_  = _w3947_ ;
	assign \g62133/_0_  = _w3948_ ;
	assign \g62135/_0_  = _w3949_ ;
	assign \g62136/_0_  = _w3950_ ;
	assign \g62137/_0_  = _w3951_ ;
	assign \g62138/_0_  = _w3952_ ;
	assign \g62140/_0_  = _w3953_ ;
	assign \g62143/_0_  = _w3954_ ;
	assign \g62144/_0_  = _w3955_ ;
	assign \g62149/_0_  = _w3956_ ;
	assign \g62150/_0_  = _w3957_ ;
	assign \g62151/_0_  = _w3958_ ;
	assign \g62153/_0_  = _w3959_ ;
	assign \g62155/_0_  = _w3960_ ;
	assign \g62156/_0_  = _w3961_ ;
	assign \g62158/_0_  = _w3962_ ;
	assign \g62160/_0_  = _w3963_ ;
	assign \g62161/_0_  = _w3964_ ;
	assign \g62162/_0_  = _w3965_ ;
	assign \g62164/_0_  = _w3966_ ;
	assign \g62165/_0_  = _w3967_ ;
	assign \g62166/_0_  = _w3968_ ;
	assign \g62167/_0_  = _w3969_ ;
	assign \g62168/_0_  = _w3970_ ;
	assign \g62169/_0_  = _w3971_ ;
	assign \g62172/_0_  = _w3972_ ;
	assign \g62173/_0_  = _w3973_ ;
	assign \g62175/_0_  = _w3974_ ;
	assign \g62176/_0_  = _w3975_ ;
	assign \g62177/_0_  = _w3976_ ;
	assign \g62178/_0_  = _w3977_ ;
	assign \g62179/_0_  = _w3978_ ;
	assign \g62180/_0_  = _w3979_ ;
	assign \g62181/_0_  = _w3980_ ;
	assign \g62182/_0_  = _w3981_ ;
	assign \g62183/_0_  = _w3982_ ;
	assign \g62184/_0_  = _w3983_ ;
	assign \g62185/_0_  = _w3984_ ;
	assign \g62186/_0_  = _w3985_ ;
	assign \g62188/_0_  = _w3986_ ;
	assign \g62189/_0_  = _w3987_ ;
	assign \g62190/_0_  = _w3988_ ;
	assign \g62191/_0_  = _w3989_ ;
	assign \g62193/_0_  = _w3990_ ;
	assign \g62194/_0_  = _w3991_ ;
	assign \g62195/_0_  = _w3992_ ;
	assign \g62196/_0_  = _w3993_ ;
	assign \g62197/_0_  = _w3994_ ;
	assign \g62200/_0_  = _w3995_ ;
	assign \g62201/_0_  = _w3996_ ;
	assign \g62202/_0_  = _w3997_ ;
	assign \g62203/_0_  = _w3998_ ;
	assign \g62205/_0_  = _w3999_ ;
	assign \g62206/_0_  = _w4000_ ;
	assign \g62207/_0_  = _w4001_ ;
	assign \g62208/_0_  = _w4002_ ;
	assign \g62209/_0_  = _w4003_ ;
	assign \g62210/_0_  = _w4004_ ;
	assign \g62211/_0_  = _w4005_ ;
	assign \g62215/_0_  = _w4006_ ;
	assign \g62218/_0_  = _w4007_ ;
	assign \g62219/_0_  = _w4008_ ;
	assign \g62221/_0_  = _w4009_ ;
	assign \g62222/_0_  = _w4010_ ;
	assign \g62223/_0_  = _w4011_ ;
	assign \g62224/_0_  = _w4012_ ;
	assign \g62225/_0_  = _w4013_ ;
	assign \g62226/_0_  = _w4014_ ;
	assign \g62229/_0_  = _w4015_ ;
	assign \g62230/_0_  = _w4016_ ;
	assign \g62231/_0_  = _w4017_ ;
	assign \g62233/_0_  = _w4018_ ;
	assign \g62236/_0_  = _w4019_ ;
	assign \g62237/_0_  = _w4020_ ;
	assign \g62238/_0_  = _w4021_ ;
	assign \g62240/_0_  = _w4022_ ;
	assign \g62241/_0_  = _w4023_ ;
	assign \g62243/_0_  = _w4024_ ;
	assign \g62244/_0_  = _w4025_ ;
	assign \g62245/_0_  = _w4026_ ;
	assign \g62247/_0_  = _w4027_ ;
	assign \g62248/_0_  = _w4028_ ;
	assign \g62250/_0_  = _w4029_ ;
	assign \g62252/_0_  = _w4030_ ;
	assign \g62253/_0_  = _w4031_ ;
	assign \g62255/_0_  = _w4032_ ;
	assign \g62256/_0_  = _w4033_ ;
	assign \g62257/_0_  = _w4034_ ;
	assign \g62258/_0_  = _w4035_ ;
	assign \g62259/_0_  = _w4036_ ;
	assign \g62260/_0_  = _w4037_ ;
	assign \g62261/_0_  = _w4038_ ;
	assign \g62262/_0_  = _w4039_ ;
	assign \g62263/_0_  = _w4040_ ;
	assign \g62264/_0_  = _w4041_ ;
	assign \g62265/_0_  = _w4042_ ;
	assign \g62267/_0_  = _w4043_ ;
	assign \g62269/_0_  = _w4044_ ;
	assign \g62270/_0_  = _w4045_ ;
	assign \g62272/_0_  = _w4046_ ;
	assign \g62274/_0_  = _w4047_ ;
	assign \g62277/_0_  = _w4048_ ;
	assign \g62279/_0_  = _w4049_ ;
	assign \g62280/_0_  = _w4050_ ;
	assign \g62281/_0_  = _w4051_ ;
	assign \g62283/_0_  = _w4052_ ;
	assign \g62284/_0_  = _w4053_ ;
	assign \g62285/_0_  = _w4054_ ;
	assign \g62286/_0_  = _w4055_ ;
	assign \g62288/_0_  = _w4056_ ;
	assign \g62289/_0_  = _w4057_ ;
	assign \g62290/_0_  = _w4058_ ;
	assign \g62294/_0_  = _w4059_ ;
	assign \g62295/_0_  = _w4060_ ;
	assign \g62296/_0_  = _w4061_ ;
	assign \g62297/_0_  = _w4062_ ;
	assign \g62298/_0_  = _w4063_ ;
	assign \g62299/_0_  = _w4064_ ;
	assign \g62303/_0_  = _w4065_ ;
	assign \g62305/_0_  = _w4066_ ;
	assign \g62306/_0_  = _w4067_ ;
	assign \g62307/_0_  = _w4068_ ;
	assign \g62309/_0_  = _w4069_ ;
	assign \g62311/_0_  = _w4070_ ;
	assign \g62312/_0_  = _w4071_ ;
	assign \g62313/_0_  = _w4072_ ;
	assign \g62314/_0_  = _w4073_ ;
	assign \g62315/_0_  = _w4074_ ;
	assign \g62316/_0_  = _w4075_ ;
	assign \g62317/_0_  = _w4076_ ;
	assign \g62318/_0_  = _w4077_ ;
	assign \g62319/_0_  = _w4078_ ;
	assign \g62320/_0_  = _w4079_ ;
	assign \g62322/_0_  = _w4080_ ;
	assign \g62324/_0_  = _w4081_ ;
	assign \g62325/_0_  = _w4082_ ;
	assign \g62326/_0_  = _w4083_ ;
	assign \g62327/_0_  = _w4084_ ;
	assign \g62329/_0_  = _w4085_ ;
	assign \g62330/_0_  = _w4086_ ;
	assign \g62331/_0_  = _w4087_ ;
	assign \g62332/_0_  = _w4088_ ;
	assign \g62333/_0_  = _w4089_ ;
	assign \g62335/_0_  = _w4090_ ;
	assign \g62336/_0_  = _w4091_ ;
	assign \g62338/_0_  = _w4092_ ;
	assign \g62341/_0_  = _w4093_ ;
	assign \g62342/_0_  = _w4094_ ;
	assign \g62344/_0_  = _w4095_ ;
	assign \g62345/_0_  = _w4096_ ;
	assign \g62348/_0_  = _w4097_ ;
	assign \g62349/_0_  = _w4098_ ;
	assign \g62350/_0_  = _w4099_ ;
	assign \g62353/_0_  = _w4100_ ;
	assign \g62354/_0_  = _w4101_ ;
	assign \g62355/_0_  = _w4102_ ;
	assign \g62356/_0_  = _w4103_ ;
	assign \g62359/_0_  = _w4104_ ;
	assign \g62362/_0_  = _w4105_ ;
	assign \g62363/_0_  = _w4106_ ;
	assign \g62364/_0_  = _w4107_ ;
	assign \g62365/_0_  = _w4108_ ;
	assign \g62366/_0_  = _w4109_ ;
	assign \g62367/_0_  = _w4110_ ;
	assign \g62368/_0_  = _w4111_ ;
	assign \g62369/_0_  = _w4112_ ;
	assign \g62370/_0_  = _w4113_ ;
	assign \g62371/_0_  = _w4114_ ;
	assign \g62372/_0_  = _w4115_ ;
	assign \g62373/_0_  = _w4116_ ;
	assign \g62374/_0_  = _w4117_ ;
	assign \g62376/_0_  = _w4118_ ;
	assign \g62467/_0_  = _w4119_ ;
	assign \g62468/_0_  = _w4120_ ;
	assign \g62469/_0_  = _w4121_ ;
	assign \g62470/_0_  = _w4122_ ;
	assign \g62471/_0_  = _w4123_ ;
	assign \g62472/_0_  = _w4124_ ;
	assign \g62473/_0_  = _w4125_ ;
	assign \g62474/_0_  = _w4126_ ;
	assign \g62475/_0_  = _w4127_ ;
	assign \g62478/_0_  = _w4128_ ;
	assign \g62480/_0_  = _w4129_ ;
	assign \g62481/_0_  = _w4130_ ;
	assign \g62482/_0_  = _w4131_ ;
	assign \g62483/_0_  = _w4132_ ;
	assign \g62484/_0_  = _w4133_ ;
	assign \g62485/_0_  = _w4134_ ;
	assign \g62486/_0_  = _w4135_ ;
	assign \g62487/_0_  = _w4136_ ;
	assign \g62488/_0_  = _w4137_ ;
	assign \g62489/_0_  = _w4138_ ;
	assign \g62490/_0_  = _w4139_ ;
	assign \g62491/_0_  = _w4140_ ;
	assign \g62492/_0_  = _w4141_ ;
	assign \g62493/_0_  = _w4142_ ;
	assign \g62494/_0_  = _w4143_ ;
	assign \g62495/_0_  = _w4144_ ;
	assign \g62496/_0_  = _w4145_ ;
	assign \g62497/_0_  = _w4146_ ;
	assign \g62498/_0_  = _w4147_ ;
	assign \g62499/_0_  = _w4148_ ;
	assign \g62500/_0_  = _w4149_ ;
	assign \g62501/_0_  = _w4150_ ;
	assign \g62502/_0_  = _w4151_ ;
	assign \g62503/_0_  = _w4152_ ;
	assign \g62504/_0_  = _w4153_ ;
	assign \g62509/_0_  = _w4154_ ;
	assign \g62510/_0_  = _w4155_ ;
	assign \g62511/_0_  = _w4156_ ;
	assign \g62512/_0_  = _w4157_ ;
	assign \g62513/_0_  = _w4158_ ;
	assign \g62514/_0_  = _w4159_ ;
	assign \g62515/_0_  = _w4160_ ;
	assign \g62516/_0_  = _w4161_ ;
	assign \g62517/_0_  = _w4162_ ;
	assign \g62518/_0_  = _w4163_ ;
	assign \g62519/_0_  = _w4164_ ;
	assign \g62520/_0_  = _w4165_ ;
	assign \g62521/_0_  = _w4166_ ;
	assign \g62523/_0_  = _w4167_ ;
	assign \g62526/_0_  = _w4168_ ;
	assign \g62528/_0_  = _w4169_ ;
	assign \g62529/_0_  = _w4170_ ;
	assign \g62531/_0_  = _w4171_ ;
	assign \g62532/_0_  = _w4172_ ;
	assign \g62533/_0_  = _w4173_ ;
	assign \g62534/_0_  = _w4174_ ;
	assign \g62535/_0_  = _w4175_ ;
	assign \g62536/_0_  = _w4176_ ;
	assign \g62537/_0_  = _w4177_ ;
	assign \g62539/_0_  = _w4178_ ;
	assign \g62540/_0_  = _w4179_ ;
	assign \g62541/_0_  = _w4180_ ;
	assign \g62542/_0_  = _w4181_ ;
	assign \g62543/_0_  = _w4182_ ;
	assign \g62544/_0_  = _w4183_ ;
	assign \g62545/_0_  = _w4184_ ;
	assign \g62547/_0_  = _w4185_ ;
	assign \g62548/_0_  = _w4186_ ;
	assign \g62549/_0_  = _w4187_ ;
	assign \g62550/_0_  = _w4188_ ;
	assign \g62551/_0_  = _w4189_ ;
	assign \g62552/_0_  = _w4190_ ;
	assign \g62553/_0_  = _w4191_ ;
	assign \g62554/_0_  = _w4192_ ;
	assign \g62555/_0_  = _w4193_ ;
	assign \g62556/_0_  = _w4194_ ;
	assign \g62557/_0_  = _w4195_ ;
	assign \g62560/_0_  = _w4196_ ;
	assign \g62562/_0_  = _w4197_ ;
	assign \g62563/_0_  = _w4198_ ;
	assign \g62564/_0_  = _w4199_ ;
	assign \g62565/_0_  = _w4200_ ;
	assign \g62566/_0_  = _w4201_ ;
	assign \g62567/_0_  = _w4202_ ;
	assign \g62569/_0_  = _w4203_ ;
	assign \g62570/_0_  = _w4204_ ;
	assign \g62571/_0_  = _w4205_ ;
	assign \g62572/_0_  = _w4206_ ;
	assign \g62573/_0_  = _w4207_ ;
	assign \g62574/_0_  = _w4208_ ;
	assign \g62576/_0_  = _w4209_ ;
	assign \g62577/_0_  = _w4210_ ;
	assign \g62581/_0_  = _w4211_ ;
	assign \g62582/_0_  = _w4212_ ;
	assign \g62584/_0_  = _w4213_ ;
	assign \g62585/_0_  = _w4214_ ;
	assign \g62586/_0_  = _w4215_ ;
	assign \g62588/_0_  = _w4216_ ;
	assign \g62589/_0_  = _w4217_ ;
	assign \g62593/_0_  = _w4218_ ;
	assign \g62594/_0_  = _w4219_ ;
	assign \g62595/_0_  = _w4220_ ;
	assign \g62596/_0_  = _w4221_ ;
	assign \g62597/_0_  = _w4222_ ;
	assign \g62598/_0_  = _w4223_ ;
	assign \g62599/_0_  = _w4224_ ;
	assign \g62600/_0_  = _w4225_ ;
	assign \g62601/_0_  = _w4226_ ;
	assign \g62602/_0_  = _w4227_ ;
	assign \g62603/_0_  = _w4228_ ;
	assign \g62604/_0_  = _w4229_ ;
	assign \g62605/_0_  = _w4230_ ;
	assign \g62606/_0_  = _w4231_ ;
	assign \g62607/_0_  = _w4232_ ;
	assign \g62608/_0_  = _w4233_ ;
	assign \g62609/_0_  = _w4234_ ;
	assign \g62610/_0_  = _w4235_ ;
	assign \g62612/_0_  = _w4236_ ;
	assign \g62613/_0_  = _w4237_ ;
	assign \g62614/_0_  = _w4238_ ;
	assign \g62615/_0_  = _w4239_ ;
	assign \g62617/_0_  = _w4240_ ;
	assign \g62618/_0_  = _w4241_ ;
	assign \g62620/_0_  = _w4242_ ;
	assign \g62621/_0_  = _w4243_ ;
	assign \g62622/_0_  = _w4244_ ;
	assign \g62624/_0_  = _w4245_ ;
	assign \g62625/_0_  = _w4246_ ;
	assign \g62626/_0_  = _w4247_ ;
	assign \g62627/_0_  = _w4248_ ;
	assign \g62629/_0_  = _w4249_ ;
	assign \g62630/_0_  = _w4250_ ;
	assign \g62632/_0_  = _w4251_ ;
	assign \g62633/_0_  = _w4252_ ;
	assign \g62635/_0_  = _w4253_ ;
	assign \g62636/_0_  = _w4254_ ;
	assign \g62637/_0_  = _w4255_ ;
	assign \g62638/_0_  = _w4256_ ;
	assign \g62640/_0_  = _w4257_ ;
	assign \g62641/_0_  = _w4258_ ;
	assign \g62642/_0_  = _w4259_ ;
	assign \g62643/_0_  = _w4260_ ;
	assign \g62644/_0_  = _w4261_ ;
	assign \g62646/_0_  = _w4262_ ;
	assign \g62647/_0_  = _w4263_ ;
	assign \g62649/_0_  = _w4264_ ;
	assign \g62650/_0_  = _w4265_ ;
	assign \g62651/_0_  = _w4266_ ;
	assign \g62653/_0_  = _w4267_ ;
	assign \g62655/_0_  = _w4268_ ;
	assign \g62656/_0_  = _w4269_ ;
	assign \g62657/_0_  = _w4270_ ;
	assign \g62658/_0_  = _w4271_ ;
	assign \g62660/_0_  = _w4272_ ;
	assign \g62661/_0_  = _w4273_ ;
	assign \g62662/_0_  = _w4274_ ;
	assign \g62663/_0_  = _w4275_ ;
	assign \g62664/_0_  = _w4276_ ;
	assign \g62665/_0_  = _w4277_ ;
	assign \g62667/_0_  = _w4278_ ;
	assign \g62669/_0_  = _w4279_ ;
	assign \g62670/_0_  = _w4280_ ;
	assign \g62671/_0_  = _w4281_ ;
	assign \g62672/_0_  = _w4282_ ;
	assign \g62674/_0_  = _w4283_ ;
	assign \g62675/_0_  = _w4284_ ;
	assign \g62676/_0_  = _w4285_ ;
	assign \g62677/_0_  = _w4286_ ;
	assign \g62678/_0_  = _w4287_ ;
	assign \g62679/_0_  = _w4288_ ;
	assign \g62680/_0_  = _w4289_ ;
	assign \g62681/_0_  = _w4290_ ;
	assign \g62682/_0_  = _w4291_ ;
	assign \g62684/_0_  = _w4292_ ;
	assign \g62685/_0_  = _w4293_ ;
	assign \g62686/_0_  = _w4294_ ;
	assign \g62687/_0_  = _w4295_ ;
	assign \g62690/_0_  = _w4296_ ;
	assign \g62693/_0_  = _w4297_ ;
	assign \g62698/_0_  = _w4298_ ;
	assign \g62699/_0_  = _w4299_ ;
	assign \g62700/_0_  = _w4300_ ;
	assign \g62701/_0_  = _w4301_ ;
	assign \g62702/_0_  = _w4302_ ;
	assign \g62703/_0_  = _w4303_ ;
	assign \g62704/_0_  = _w4304_ ;
	assign \g62709/_0_  = _w4305_ ;
	assign \g62710/_0_  = _w4306_ ;
	assign \g62711/_0_  = _w4307_ ;
	assign \g62714/_0_  = _w4308_ ;
	assign \g62715/_0_  = _w4309_ ;
	assign \g62717/_0_  = _w4310_ ;
	assign \g62718/_0_  = _w4311_ ;
	assign \g62719/_0_  = _w4312_ ;
	assign \g62720/_0_  = _w4313_ ;
	assign \g62721/_0_  = _w4314_ ;
	assign \g62723/_0_  = _w4315_ ;
	assign \g62725/_0_  = _w4316_ ;
	assign \g62726/_0_  = _w4317_ ;
	assign \g62729/_0_  = _w4318_ ;
	assign \g62731/_0_  = _w4319_ ;
	assign \g62733/_0_  = _w4320_ ;
	assign \g62738/_0_  = _w4321_ ;
	assign \g62741/_0_  = _w4322_ ;
	assign \g62742/_0_  = _w4323_ ;
	assign \g62744/_0_  = _w4324_ ;
	assign \g62745/_0_  = _w4325_ ;
	assign \g62746/_0_  = _w4326_ ;
	assign \g62747/_0_  = _w4327_ ;
	assign \g62748/_0_  = _w4328_ ;
	assign \g62749/_0_  = _w4329_ ;
	assign \g62753/_0_  = _w4330_ ;
	assign \g62755/_0_  = _w4331_ ;
	assign \g62756/_0_  = _w4332_ ;
	assign \g62758/_0_  = _w4333_ ;
	assign \g62759/_0_  = _w4334_ ;
	assign \g62760/_0_  = _w4335_ ;
	assign \g62761/_0_  = _w4336_ ;
	assign \g62763/_0_  = _w4337_ ;
	assign \g62766/_0_  = _w4338_ ;
	assign \g62767/_0_  = _w4339_ ;
	assign \g62768/_0_  = _w4340_ ;
	assign \g65554/_0_  = _w4344_ ;
	assign \g65561/_0_  = _w4348_ ;
	assign \g65569/_0_  = _w4352_ ;
	assign \g65580/_0_  = _w4356_ ;
	assign \g65599/_0_  = _w4360_ ;
	assign \g65606/_0_  = _w4364_ ;
	assign \g65636/_0_  = _w4368_ ;
	assign \g65864/_0_  = _w4373_ ;
endmodule;