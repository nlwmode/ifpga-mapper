module top (a_pad, b_pad, c_pad, d_pad, e_pad, f_pad, g_pad, h_pad, i_pad, j_pad, k_pad, l_pad, m_pad, n_pad);
	input a_pad ;
	input b_pad ;
	input c_pad ;
	input d_pad ;
	input e_pad ;
	input f_pad ;
	input g_pad ;
	input h_pad ;
	input i_pad ;
	input j_pad ;
	input k_pad ;
	output l_pad ;
	output m_pad ;
	output n_pad ;
	wire _w42_ ;
	wire _w41_ ;
	wire _w24_ ;
	wire _w23_ ;
	wire _w22_ ;
	wire _w21_ ;
	wire _w20_ ;
	wire _w19_ ;
	wire _w18_ ;
	wire _w17_ ;
	wire _w16_ ;
	wire _w15_ ;
	wire _w14_ ;
	wire _w13_ ;
	wire _w12_ ;
	wire _w25_ ;
	wire _w26_ ;
	wire _w27_ ;
	wire _w28_ ;
	wire _w29_ ;
	wire _w30_ ;
	wire _w31_ ;
	wire _w32_ ;
	wire _w33_ ;
	wire _w34_ ;
	wire _w35_ ;
	wire _w36_ ;
	wire _w37_ ;
	wire _w38_ ;
	wire _w39_ ;
	wire _w40_ ;
	LUT2 #(
		.INIT('h4)
	) name0 (
		f_pad,
		g_pad,
		_w12_
	);
	LUT2 #(
		.INIT('h4)
	) name1 (
		h_pad,
		i_pad,
		_w13_
	);
	LUT2 #(
		.INIT('h4)
	) name2 (
		j_pad,
		k_pad,
		_w14_
	);
	LUT2 #(
		.INIT('h1)
	) name3 (
		_w13_,
		_w14_,
		_w15_
	);
	LUT2 #(
		.INIT('h2)
	) name4 (
		h_pad,
		i_pad,
		_w16_
	);
	LUT2 #(
		.INIT('h2)
	) name5 (
		f_pad,
		g_pad,
		_w17_
	);
	LUT2 #(
		.INIT('h1)
	) name6 (
		_w16_,
		_w17_,
		_w18_
	);
	LUT2 #(
		.INIT('h4)
	) name7 (
		_w15_,
		_w18_,
		_w19_
	);
	LUT2 #(
		.INIT('h1)
	) name8 (
		_w12_,
		_w19_,
		_w20_
	);
	LUT2 #(
		.INIT('h1)
	) name9 (
		d_pad,
		e_pad,
		_w21_
	);
	LUT2 #(
		.INIT('h8)
	) name10 (
		d_pad,
		e_pad,
		_w22_
	);
	LUT2 #(
		.INIT('h1)
	) name11 (
		_w21_,
		_w22_,
		_w23_
	);
	LUT2 #(
		.INIT('h2)
	) name12 (
		b_pad,
		_w23_,
		_w24_
	);
	LUT2 #(
		.INIT('h4)
	) name13 (
		_w20_,
		_w24_,
		_w25_
	);
	LUT2 #(
		.INIT('h2)
	) name14 (
		b_pad,
		d_pad,
		_w26_
	);
	LUT2 #(
		.INIT('h8)
	) name15 (
		e_pad,
		_w26_,
		_w27_
	);
	LUT2 #(
		.INIT('h1)
	) name16 (
		a_pad,
		_w27_,
		_w28_
	);
	LUT2 #(
		.INIT('h4)
	) name17 (
		_w25_,
		_w28_,
		_w29_
	);
	LUT2 #(
		.INIT('h1)
	) name18 (
		_w12_,
		_w13_,
		_w30_
	);
	LUT2 #(
		.INIT('h2)
	) name19 (
		j_pad,
		k_pad,
		_w31_
	);
	LUT2 #(
		.INIT('h2)
	) name20 (
		_w18_,
		_w31_,
		_w32_
	);
	LUT2 #(
		.INIT('h4)
	) name21 (
		_w14_,
		_w30_,
		_w33_
	);
	LUT2 #(
		.INIT('h8)
	) name22 (
		_w24_,
		_w33_,
		_w34_
	);
	LUT2 #(
		.INIT('h8)
	) name23 (
		_w32_,
		_w34_,
		_w35_
	);
	LUT2 #(
		.INIT('h8)
	) name24 (
		b_pad,
		d_pad,
		_w36_
	);
	LUT2 #(
		.INIT('h4)
	) name25 (
		e_pad,
		_w36_,
		_w37_
	);
	LUT2 #(
		.INIT('h1)
	) name26 (
		_w17_,
		_w30_,
		_w38_
	);
	LUT2 #(
		.INIT('h2)
	) name27 (
		_w24_,
		_w32_,
		_w39_
	);
	LUT2 #(
		.INIT('h4)
	) name28 (
		_w38_,
		_w39_,
		_w40_
	);
	LUT2 #(
		.INIT('h1)
	) name29 (
		c_pad,
		_w37_,
		_w41_
	);
	LUT2 #(
		.INIT('h4)
	) name30 (
		_w40_,
		_w41_,
		_w42_
	);
	assign l_pad = _w29_ ;
	assign m_pad = _w35_ ;
	assign n_pad = _w42_ ;
endmodule;