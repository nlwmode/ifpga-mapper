module top (\ac97_reset_pad_o__pad , \dma_ack_i[0]_pad , \dma_ack_i[1]_pad , \dma_ack_i[2]_pad , \dma_ack_i[3]_pad , \dma_ack_i[4]_pad , \dma_ack_i[5]_pad , \dma_ack_i[6]_pad , \dma_ack_i[7]_pad , \dma_ack_i[8]_pad , \dma_req_o[0]_pad , \dma_req_o[1]_pad , \dma_req_o[2]_pad , \dma_req_o[3]_pad , \dma_req_o[4]_pad , \dma_req_o[5]_pad , \dma_req_o[6]_pad , \dma_req_o[7]_pad , \dma_req_o[8]_pad , \in_valid_s_reg[0]/NET0131 , \in_valid_s_reg[1]/NET0131 , \in_valid_s_reg[2]/NET0131 , suspended_o_pad, \u0_slt0_r_reg[0]/P0001 , \u0_slt0_r_reg[10]/P0001 , \u0_slt0_r_reg[11]/P0001 , \u0_slt0_r_reg[12]/P0001 , \u0_slt0_r_reg[13]/P0001 , \u0_slt0_r_reg[14]/P0001 , \u0_slt0_r_reg[1]/P0001 , \u0_slt0_r_reg[2]/P0001 , \u0_slt0_r_reg[3]/P0001 , \u0_slt0_r_reg[4]/P0001 , \u0_slt0_r_reg[5]/P0001 , \u0_slt0_r_reg[6]/P0001 , \u0_slt0_r_reg[7]/P0001 , \u0_slt0_r_reg[8]/P0001 , \u0_slt0_r_reg[9]/P0001 , \u0_slt1_r_reg[0]/P0001 , \u0_slt1_r_reg[10]/P0001 , \u0_slt1_r_reg[11]/P0001 , \u0_slt1_r_reg[12]/P0001 , \u0_slt1_r_reg[13]/P0001 , \u0_slt1_r_reg[14]/P0001 , \u0_slt1_r_reg[15]/P0001 , \u0_slt1_r_reg[16]/P0001 , \u0_slt1_r_reg[17]/P0001 , \u0_slt1_r_reg[18]/P0001 , \u0_slt1_r_reg[19]/P0001 , \u0_slt1_r_reg[1]/P0001 , \u0_slt1_r_reg[2]/P0001 , \u0_slt1_r_reg[3]/P0001 , \u0_slt1_r_reg[4]/P0001 , \u0_slt1_r_reg[5]/P0001 , \u0_slt1_r_reg[6]/P0001 , \u0_slt1_r_reg[7]/P0001 , \u0_slt1_r_reg[8]/P0001 , \u0_slt1_r_reg[9]/P0001 , \u0_slt2_r_reg[0]/P0001 , \u0_slt2_r_reg[10]/P0001 , \u0_slt2_r_reg[11]/P0001 , \u0_slt2_r_reg[12]/P0001 , \u0_slt2_r_reg[13]/P0001 , \u0_slt2_r_reg[14]/P0001 , \u0_slt2_r_reg[15]/P0001 , \u0_slt2_r_reg[16]/P0001 , \u0_slt2_r_reg[17]/P0001 , \u0_slt2_r_reg[18]/P0001 , \u0_slt2_r_reg[19]/P0001 , \u0_slt2_r_reg[1]/P0001 , \u0_slt2_r_reg[2]/P0001 , \u0_slt2_r_reg[3]/P0001 , \u0_slt2_r_reg[4]/P0001 , \u0_slt2_r_reg[5]/P0001 , \u0_slt2_r_reg[6]/P0001 , \u0_slt2_r_reg[7]/P0001 , \u0_slt2_r_reg[8]/P0001 , \u0_slt2_r_reg[9]/P0001 , \u0_slt3_r_reg[0]/P0001 , \u0_slt3_r_reg[10]/P0001 , \u0_slt3_r_reg[11]/P0001 , \u0_slt3_r_reg[12]/P0001 , \u0_slt3_r_reg[13]/P0001 , \u0_slt3_r_reg[14]/P0001 , \u0_slt3_r_reg[15]/P0001 , \u0_slt3_r_reg[16]/P0001 , \u0_slt3_r_reg[17]/P0001 , \u0_slt3_r_reg[18]/P0001 , \u0_slt3_r_reg[19]/P0001 , \u0_slt3_r_reg[1]/P0001 , \u0_slt3_r_reg[2]/P0001 , \u0_slt3_r_reg[3]/P0001 , \u0_slt3_r_reg[4]/P0001 , \u0_slt3_r_reg[5]/P0001 , \u0_slt3_r_reg[6]/P0001 , \u0_slt3_r_reg[7]/P0001 , \u0_slt3_r_reg[8]/P0001 , \u0_slt3_r_reg[9]/P0001 , \u0_slt4_r_reg[0]/P0001 , \u0_slt4_r_reg[10]/P0001 , \u0_slt4_r_reg[11]/P0001 , \u0_slt4_r_reg[12]/P0001 , \u0_slt4_r_reg[13]/P0001 , \u0_slt4_r_reg[14]/P0001 , \u0_slt4_r_reg[15]/P0001 , \u0_slt4_r_reg[16]/P0001 , \u0_slt4_r_reg[17]/P0001 , \u0_slt4_r_reg[18]/P0001 , \u0_slt4_r_reg[19]/P0001 , \u0_slt4_r_reg[1]/P0001 , \u0_slt4_r_reg[2]/P0001 , \u0_slt4_r_reg[3]/P0001 , \u0_slt4_r_reg[4]/P0001 , \u0_slt4_r_reg[5]/P0001 , \u0_slt4_r_reg[6]/P0001 , \u0_slt4_r_reg[7]/P0001 , \u0_slt4_r_reg[8]/P0001 , \u0_slt4_r_reg[9]/P0001 , \u0_slt5_r_reg[0]/P0001 , \u0_slt5_r_reg[10]/P0001 , \u0_slt5_r_reg[11]/P0001 , \u0_slt5_r_reg[12]/P0001 , \u0_slt5_r_reg[13]/P0001 , \u0_slt5_r_reg[14]/P0001 , \u0_slt5_r_reg[15]/P0001 , \u0_slt5_r_reg[16]/P0001 , \u0_slt5_r_reg[17]/P0001 , \u0_slt5_r_reg[18]/P0001 , \u0_slt5_r_reg[19]/P0001 , \u0_slt5_r_reg[1]/P0001 , \u0_slt5_r_reg[2]/P0001 , \u0_slt5_r_reg[3]/P0001 , \u0_slt5_r_reg[4]/P0001 , \u0_slt5_r_reg[5]/P0001 , \u0_slt5_r_reg[6]/P0001 , \u0_slt5_r_reg[7]/P0001 , \u0_slt5_r_reg[8]/P0001 , \u0_slt5_r_reg[9]/P0001 , \u0_slt6_r_reg[0]/P0001 , \u0_slt6_r_reg[10]/P0001 , \u0_slt6_r_reg[11]/P0001 , \u0_slt6_r_reg[12]/P0001 , \u0_slt6_r_reg[13]/P0001 , \u0_slt6_r_reg[14]/P0001 , \u0_slt6_r_reg[15]/P0001 , \u0_slt6_r_reg[16]/P0001 , \u0_slt6_r_reg[17]/P0001 , \u0_slt6_r_reg[18]/P0001 , \u0_slt6_r_reg[19]/P0001 , \u0_slt6_r_reg[1]/P0001 , \u0_slt6_r_reg[2]/P0001 , \u0_slt6_r_reg[3]/P0001 , \u0_slt6_r_reg[4]/P0001 , \u0_slt6_r_reg[5]/P0001 , \u0_slt6_r_reg[6]/P0001 , \u0_slt6_r_reg[7]/P0001 , \u0_slt6_r_reg[8]/P0001 , \u0_slt6_r_reg[9]/P0001 , \u0_slt7_r_reg[0]/P0001 , \u0_slt7_r_reg[10]/P0001 , \u0_slt7_r_reg[11]/P0001 , \u0_slt7_r_reg[12]/P0001 , \u0_slt7_r_reg[13]/P0001 , \u0_slt7_r_reg[14]/P0001 , \u0_slt7_r_reg[15]/P0001 , \u0_slt7_r_reg[16]/P0001 , \u0_slt7_r_reg[17]/P0001 , \u0_slt7_r_reg[18]/P0001 , \u0_slt7_r_reg[19]/P0001 , \u0_slt7_r_reg[1]/P0001 , \u0_slt7_r_reg[2]/P0001 , \u0_slt7_r_reg[3]/P0001 , \u0_slt7_r_reg[4]/P0001 , \u0_slt7_r_reg[5]/P0001 , \u0_slt7_r_reg[6]/P0001 , \u0_slt7_r_reg[7]/P0001 , \u0_slt7_r_reg[8]/P0001 , \u0_slt7_r_reg[9]/P0001 , \u0_slt8_r_reg[0]/P0001 , \u0_slt8_r_reg[10]/P0001 , \u0_slt8_r_reg[11]/P0001 , \u0_slt8_r_reg[12]/P0001 , \u0_slt8_r_reg[13]/P0001 , \u0_slt8_r_reg[14]/P0001 , \u0_slt8_r_reg[15]/P0001 , \u0_slt8_r_reg[16]/P0001 , \u0_slt8_r_reg[17]/P0001 , \u0_slt8_r_reg[18]/P0001 , \u0_slt8_r_reg[19]/P0001 , \u0_slt8_r_reg[1]/P0001 , \u0_slt8_r_reg[2]/P0001 , \u0_slt8_r_reg[3]/P0001 , \u0_slt8_r_reg[4]/P0001 , \u0_slt8_r_reg[5]/P0001 , \u0_slt8_r_reg[6]/P0001 , \u0_slt8_r_reg[7]/P0001 , \u0_slt8_r_reg[8]/P0001 , \u0_slt8_r_reg[9]/P0001 , \u0_slt9_r_reg[0]/P0001 , \u0_slt9_r_reg[10]/P0001 , \u0_slt9_r_reg[11]/P0001 , \u0_slt9_r_reg[12]/P0001 , \u0_slt9_r_reg[13]/P0001 , \u0_slt9_r_reg[14]/P0001 , \u0_slt9_r_reg[15]/P0001 , \u0_slt9_r_reg[16]/P0001 , \u0_slt9_r_reg[17]/P0001 , \u0_slt9_r_reg[18]/P0001 , \u0_slt9_r_reg[19]/P0001 , \u0_slt9_r_reg[1]/P0001 , \u0_slt9_r_reg[2]/P0001 , \u0_slt9_r_reg[3]/P0001 , \u0_slt9_r_reg[4]/P0001 , \u0_slt9_r_reg[5]/P0001 , \u0_slt9_r_reg[6]/P0001 , \u0_slt9_r_reg[7]/P0001 , \u0_slt9_r_reg[8]/P0001 , \u0_slt9_r_reg[9]/P0001 , \u10_din_tmp1_reg[0]/P0001 , \u10_din_tmp1_reg[10]/P0001 , \u10_din_tmp1_reg[11]/P0001 , \u10_din_tmp1_reg[12]/P0001 , \u10_din_tmp1_reg[13]/P0001 , \u10_din_tmp1_reg[14]/P0001 , \u10_din_tmp1_reg[15]/P0001 , \u10_din_tmp1_reg[1]/P0001 , \u10_din_tmp1_reg[2]/P0001 , \u10_din_tmp1_reg[3]/P0001 , \u10_din_tmp1_reg[4]/P0001 , \u10_din_tmp1_reg[5]/P0001 , \u10_din_tmp1_reg[6]/P0001 , \u10_din_tmp1_reg[7]/P0001 , \u10_din_tmp1_reg[8]/P0001 , \u10_din_tmp1_reg[9]/P0001 , \u10_dout_reg[0]/P0001 , \u10_dout_reg[10]/P0001 , \u10_dout_reg[11]/P0001 , \u10_dout_reg[12]/P0001 , \u10_dout_reg[13]/P0001 , \u10_dout_reg[14]/P0001 , \u10_dout_reg[15]/P0001 , \u10_dout_reg[16]/P0001 , \u10_dout_reg[17]/P0001 , \u10_dout_reg[18]/P0001 , \u10_dout_reg[19]/P0001 , \u10_dout_reg[1]/P0001 , \u10_dout_reg[20]/P0001 , \u10_dout_reg[21]/P0001 , \u10_dout_reg[22]/P0001 , \u10_dout_reg[23]/P0001 , \u10_dout_reg[24]/P0001 , \u10_dout_reg[25]/P0001 , \u10_dout_reg[26]/P0001 , \u10_dout_reg[27]/P0001 , \u10_dout_reg[28]/P0001 , \u10_dout_reg[29]/P0001 , \u10_dout_reg[2]/P0001 , \u10_dout_reg[30]/P0001 , \u10_dout_reg[31]/P0001 , \u10_dout_reg[3]/P0001 , \u10_dout_reg[4]/P0001 , \u10_dout_reg[5]/P0001 , \u10_dout_reg[6]/P0001 , \u10_dout_reg[7]/P0001 , \u10_dout_reg[8]/P0001 , \u10_dout_reg[9]/P0001 , \u10_empty_reg/P0001 , \u10_full_reg/NET0131 , \u10_mem_reg[0][0]/P0001 , \u10_mem_reg[0][10]/P0001 , \u10_mem_reg[0][11]/P0001 , \u10_mem_reg[0][12]/P0001 , \u10_mem_reg[0][13]/P0001 , \u10_mem_reg[0][14]/P0001 , \u10_mem_reg[0][15]/P0001 , \u10_mem_reg[0][16]/P0001 , \u10_mem_reg[0][17]/P0001 , \u10_mem_reg[0][18]/P0001 , \u10_mem_reg[0][19]/P0001 , \u10_mem_reg[0][1]/P0001 , \u10_mem_reg[0][20]/P0001 , \u10_mem_reg[0][21]/P0001 , \u10_mem_reg[0][22]/P0001 , \u10_mem_reg[0][23]/P0001 , \u10_mem_reg[0][24]/P0001 , \u10_mem_reg[0][25]/P0001 , \u10_mem_reg[0][26]/P0001 , \u10_mem_reg[0][27]/P0001 , \u10_mem_reg[0][28]/P0001 , \u10_mem_reg[0][29]/P0001 , \u10_mem_reg[0][2]/P0001 , \u10_mem_reg[0][30]/P0001 , \u10_mem_reg[0][31]/P0001 , \u10_mem_reg[0][3]/P0001 , \u10_mem_reg[0][4]/P0001 , \u10_mem_reg[0][5]/P0001 , \u10_mem_reg[0][6]/P0001 , \u10_mem_reg[0][7]/P0001 , \u10_mem_reg[0][8]/P0001 , \u10_mem_reg[0][9]/P0001 , \u10_mem_reg[1][0]/P0001 , \u10_mem_reg[1][10]/P0001 , \u10_mem_reg[1][11]/P0001 , \u10_mem_reg[1][12]/P0001 , \u10_mem_reg[1][13]/P0001 , \u10_mem_reg[1][14]/P0001 , \u10_mem_reg[1][15]/P0001 , \u10_mem_reg[1][16]/P0001 , \u10_mem_reg[1][17]/P0001 , \u10_mem_reg[1][18]/P0001 , \u10_mem_reg[1][19]/P0001 , \u10_mem_reg[1][1]/P0001 , \u10_mem_reg[1][20]/P0001 , \u10_mem_reg[1][21]/P0001 , \u10_mem_reg[1][22]/P0001 , \u10_mem_reg[1][23]/P0001 , \u10_mem_reg[1][24]/P0001 , \u10_mem_reg[1][25]/P0001 , \u10_mem_reg[1][26]/P0001 , \u10_mem_reg[1][27]/P0001 , \u10_mem_reg[1][28]/P0001 , \u10_mem_reg[1][29]/P0001 , \u10_mem_reg[1][2]/P0001 , \u10_mem_reg[1][30]/P0001 , \u10_mem_reg[1][31]/P0001 , \u10_mem_reg[1][3]/P0001 , \u10_mem_reg[1][4]/P0001 , \u10_mem_reg[1][5]/P0001 , \u10_mem_reg[1][6]/P0001 , \u10_mem_reg[1][7]/P0001 , \u10_mem_reg[1][8]/P0001 , \u10_mem_reg[1][9]/P0001 , \u10_mem_reg[2][0]/P0001 , \u10_mem_reg[2][10]/P0001 , \u10_mem_reg[2][11]/P0001 , \u10_mem_reg[2][12]/P0001 , \u10_mem_reg[2][13]/P0001 , \u10_mem_reg[2][14]/P0001 , \u10_mem_reg[2][15]/P0001 , \u10_mem_reg[2][16]/P0001 , \u10_mem_reg[2][17]/P0001 , \u10_mem_reg[2][18]/P0001 , \u10_mem_reg[2][19]/P0001 , \u10_mem_reg[2][1]/P0001 , \u10_mem_reg[2][20]/P0001 , \u10_mem_reg[2][21]/P0001 , \u10_mem_reg[2][22]/P0001 , \u10_mem_reg[2][23]/P0001 , \u10_mem_reg[2][24]/P0001 , \u10_mem_reg[2][25]/P0001 , \u10_mem_reg[2][26]/P0001 , \u10_mem_reg[2][27]/P0001 , \u10_mem_reg[2][28]/P0001 , \u10_mem_reg[2][29]/P0001 , \u10_mem_reg[2][2]/P0001 , \u10_mem_reg[2][30]/P0001 , \u10_mem_reg[2][31]/P0001 , \u10_mem_reg[2][3]/P0001 , \u10_mem_reg[2][4]/P0001 , \u10_mem_reg[2][5]/P0001 , \u10_mem_reg[2][6]/P0001 , \u10_mem_reg[2][7]/P0001 , \u10_mem_reg[2][8]/P0001 , \u10_mem_reg[2][9]/P0001 , \u10_mem_reg[3][0]/P0001 , \u10_mem_reg[3][10]/P0001 , \u10_mem_reg[3][11]/P0001 , \u10_mem_reg[3][12]/P0001 , \u10_mem_reg[3][13]/P0001 , \u10_mem_reg[3][14]/P0001 , \u10_mem_reg[3][15]/P0001 , \u10_mem_reg[3][16]/P0001 , \u10_mem_reg[3][17]/P0001 , \u10_mem_reg[3][18]/P0001 , \u10_mem_reg[3][19]/P0001 , \u10_mem_reg[3][1]/P0001 , \u10_mem_reg[3][20]/P0001 , \u10_mem_reg[3][21]/P0001 , \u10_mem_reg[3][22]/P0001 , \u10_mem_reg[3][23]/P0001 , \u10_mem_reg[3][24]/P0001 , \u10_mem_reg[3][25]/P0001 , \u10_mem_reg[3][26]/P0001 , \u10_mem_reg[3][27]/P0001 , \u10_mem_reg[3][28]/P0001 , \u10_mem_reg[3][29]/P0001 , \u10_mem_reg[3][2]/P0001 , \u10_mem_reg[3][30]/P0001 , \u10_mem_reg[3][31]/P0001 , \u10_mem_reg[3][3]/P0001 , \u10_mem_reg[3][4]/P0001 , \u10_mem_reg[3][5]/P0001 , \u10_mem_reg[3][6]/P0001 , \u10_mem_reg[3][7]/P0001 , \u10_mem_reg[3][8]/P0001 , \u10_mem_reg[3][9]/P0001 , \u10_rp_reg[0]/P0001 , \u10_rp_reg[1]/P0001 , \u10_rp_reg[2]/P0001 , \u10_status_reg[0]/P0001 , \u10_status_reg[1]/P0001 , \u10_wp_reg[0]/NET0131 , \u10_wp_reg[1]/P0001 , \u10_wp_reg[2]/P0001 , \u10_wp_reg[3]/P0001 , \u11_din_tmp1_reg[0]/P0001 , \u11_din_tmp1_reg[10]/P0001 , \u11_din_tmp1_reg[11]/P0001 , \u11_din_tmp1_reg[12]/P0001 , \u11_din_tmp1_reg[13]/P0001 , \u11_din_tmp1_reg[14]/P0001 , \u11_din_tmp1_reg[15]/P0001 , \u11_din_tmp1_reg[1]/P0001 , \u11_din_tmp1_reg[2]/P0001 , \u11_din_tmp1_reg[3]/P0001 , \u11_din_tmp1_reg[4]/P0001 , \u11_din_tmp1_reg[5]/P0001 , \u11_din_tmp1_reg[6]/P0001 , \u11_din_tmp1_reg[7]/P0001 , \u11_din_tmp1_reg[8]/P0001 , \u11_din_tmp1_reg[9]/P0001 , \u11_dout_reg[0]/P0001 , \u11_dout_reg[10]/P0001 , \u11_dout_reg[11]/P0001 , \u11_dout_reg[12]/P0001 , \u11_dout_reg[13]/P0001 , \u11_dout_reg[14]/P0001 , \u11_dout_reg[15]/P0001 , \u11_dout_reg[16]/P0001 , \u11_dout_reg[17]/P0001 , \u11_dout_reg[18]/P0001 , \u11_dout_reg[19]/P0001 , \u11_dout_reg[1]/P0001 , \u11_dout_reg[20]/P0001 , \u11_dout_reg[21]/P0001 , \u11_dout_reg[22]/P0001 , \u11_dout_reg[23]/P0001 , \u11_dout_reg[24]/P0001 , \u11_dout_reg[25]/P0001 , \u11_dout_reg[26]/P0001 , \u11_dout_reg[27]/P0001 , \u11_dout_reg[28]/P0001 , \u11_dout_reg[29]/P0001 , \u11_dout_reg[2]/P0001 , \u11_dout_reg[30]/P0001 , \u11_dout_reg[31]/P0001 , \u11_dout_reg[3]/P0001 , \u11_dout_reg[4]/P0001 , \u11_dout_reg[5]/P0001 , \u11_dout_reg[6]/P0001 , \u11_dout_reg[7]/P0001 , \u11_dout_reg[8]/P0001 , \u11_dout_reg[9]/P0001 , \u11_empty_reg/P0001 , \u11_full_reg/NET0131 , \u11_mem_reg[0][0]/P0001 , \u11_mem_reg[0][10]/P0001 , \u11_mem_reg[0][11]/P0001 , \u11_mem_reg[0][12]/P0001 , \u11_mem_reg[0][13]/P0001 , \u11_mem_reg[0][14]/P0001 , \u11_mem_reg[0][15]/P0001 , \u11_mem_reg[0][16]/P0001 , \u11_mem_reg[0][17]/P0001 , \u11_mem_reg[0][18]/P0001 , \u11_mem_reg[0][19]/P0001 , \u11_mem_reg[0][1]/P0001 , \u11_mem_reg[0][20]/P0001 , \u11_mem_reg[0][21]/P0001 , \u11_mem_reg[0][22]/P0001 , \u11_mem_reg[0][23]/P0001 , \u11_mem_reg[0][24]/P0001 , \u11_mem_reg[0][25]/P0001 , \u11_mem_reg[0][26]/P0001 , \u11_mem_reg[0][27]/P0001 , \u11_mem_reg[0][28]/P0001 , \u11_mem_reg[0][29]/P0001 , \u11_mem_reg[0][2]/P0001 , \u11_mem_reg[0][30]/P0001 , \u11_mem_reg[0][31]/P0001 , \u11_mem_reg[0][3]/P0001 , \u11_mem_reg[0][4]/P0001 , \u11_mem_reg[0][5]/P0001 , \u11_mem_reg[0][6]/P0001 , \u11_mem_reg[0][7]/P0001 , \u11_mem_reg[0][8]/P0001 , \u11_mem_reg[0][9]/P0001 , \u11_mem_reg[1][0]/P0001 , \u11_mem_reg[1][10]/P0001 , \u11_mem_reg[1][11]/P0001 , \u11_mem_reg[1][12]/P0001 , \u11_mem_reg[1][13]/P0001 , \u11_mem_reg[1][14]/P0001 , \u11_mem_reg[1][15]/P0001 , \u11_mem_reg[1][16]/P0001 , \u11_mem_reg[1][17]/P0001 , \u11_mem_reg[1][18]/P0001 , \u11_mem_reg[1][19]/P0001 , \u11_mem_reg[1][1]/P0001 , \u11_mem_reg[1][20]/P0001 , \u11_mem_reg[1][21]/P0001 , \u11_mem_reg[1][22]/P0001 , \u11_mem_reg[1][23]/P0001 , \u11_mem_reg[1][24]/P0001 , \u11_mem_reg[1][25]/P0001 , \u11_mem_reg[1][26]/P0001 , \u11_mem_reg[1][27]/P0001 , \u11_mem_reg[1][28]/P0001 , \u11_mem_reg[1][29]/P0001 , \u11_mem_reg[1][2]/P0001 , \u11_mem_reg[1][30]/P0001 , \u11_mem_reg[1][31]/P0001 , \u11_mem_reg[1][3]/P0001 , \u11_mem_reg[1][4]/P0001 , \u11_mem_reg[1][5]/P0001 , \u11_mem_reg[1][6]/P0001 , \u11_mem_reg[1][7]/P0001 , \u11_mem_reg[1][8]/P0001 , \u11_mem_reg[1][9]/P0001 , \u11_mem_reg[2][0]/P0001 , \u11_mem_reg[2][10]/P0001 , \u11_mem_reg[2][11]/P0001 , \u11_mem_reg[2][12]/P0001 , \u11_mem_reg[2][13]/P0001 , \u11_mem_reg[2][14]/P0001 , \u11_mem_reg[2][15]/P0001 , \u11_mem_reg[2][16]/P0001 , \u11_mem_reg[2][17]/P0001 , \u11_mem_reg[2][18]/P0001 , \u11_mem_reg[2][19]/P0001 , \u11_mem_reg[2][1]/P0001 , \u11_mem_reg[2][20]/P0001 , \u11_mem_reg[2][21]/P0001 , \u11_mem_reg[2][22]/P0001 , \u11_mem_reg[2][23]/P0001 , \u11_mem_reg[2][24]/P0001 , \u11_mem_reg[2][25]/P0001 , \u11_mem_reg[2][26]/P0001 , \u11_mem_reg[2][27]/P0001 , \u11_mem_reg[2][28]/P0001 , \u11_mem_reg[2][29]/P0001 , \u11_mem_reg[2][2]/P0001 , \u11_mem_reg[2][30]/P0001 , \u11_mem_reg[2][31]/P0001 , \u11_mem_reg[2][3]/P0001 , \u11_mem_reg[2][4]/P0001 , \u11_mem_reg[2][5]/P0001 , \u11_mem_reg[2][6]/P0001 , \u11_mem_reg[2][7]/P0001 , \u11_mem_reg[2][8]/P0001 , \u11_mem_reg[2][9]/P0001 , \u11_mem_reg[3][0]/P0001 , \u11_mem_reg[3][10]/P0001 , \u11_mem_reg[3][11]/P0001 , \u11_mem_reg[3][12]/P0001 , \u11_mem_reg[3][13]/P0001 , \u11_mem_reg[3][14]/P0001 , \u11_mem_reg[3][15]/P0001 , \u11_mem_reg[3][16]/P0001 , \u11_mem_reg[3][17]/P0001 , \u11_mem_reg[3][18]/P0001 , \u11_mem_reg[3][19]/P0001 , \u11_mem_reg[3][1]/P0001 , \u11_mem_reg[3][20]/P0001 , \u11_mem_reg[3][21]/P0001 , \u11_mem_reg[3][22]/P0001 , \u11_mem_reg[3][23]/P0001 , \u11_mem_reg[3][24]/P0001 , \u11_mem_reg[3][25]/P0001 , \u11_mem_reg[3][26]/P0001 , \u11_mem_reg[3][27]/P0001 , \u11_mem_reg[3][28]/P0001 , \u11_mem_reg[3][29]/P0001 , \u11_mem_reg[3][2]/P0001 , \u11_mem_reg[3][30]/P0001 , \u11_mem_reg[3][31]/P0001 , \u11_mem_reg[3][3]/P0001 , \u11_mem_reg[3][4]/P0001 , \u11_mem_reg[3][5]/P0001 , \u11_mem_reg[3][6]/P0001 , \u11_mem_reg[3][7]/P0001 , \u11_mem_reg[3][8]/P0001 , \u11_mem_reg[3][9]/P0001 , \u11_rp_reg[0]/P0001 , \u11_rp_reg[1]/P0001 , \u11_rp_reg[2]/P0001 , \u11_status_reg[0]/P0001 , \u11_status_reg[1]/P0001 , \u11_wp_reg[0]/NET0131 , \u11_wp_reg[1]/P0001 , \u11_wp_reg[2]/P0001 , \u11_wp_reg[3]/P0001 , \u12_dout_reg[0]/P0001 , \u12_dout_reg[10]/P0001 , \u12_dout_reg[11]/P0001 , \u12_dout_reg[12]/P0001 , \u12_dout_reg[13]/P0001 , \u12_dout_reg[14]/P0001 , \u12_dout_reg[15]/P0001 , \u12_dout_reg[16]/P0001 , \u12_dout_reg[17]/P0001 , \u12_dout_reg[18]/P0001 , \u12_dout_reg[19]/P0001 , \u12_dout_reg[1]/P0001 , \u12_dout_reg[20]/P0001 , \u12_dout_reg[21]/P0001 , \u12_dout_reg[22]/P0001 , \u12_dout_reg[23]/P0001 , \u12_dout_reg[24]/P0001 , \u12_dout_reg[25]/P0001 , \u12_dout_reg[26]/P0001 , \u12_dout_reg[27]/P0001 , \u12_dout_reg[28]/P0001 , \u12_dout_reg[29]/P0001 , \u12_dout_reg[2]/P0001 , \u12_dout_reg[30]/P0001 , \u12_dout_reg[31]/P0001 , \u12_dout_reg[3]/P0001 , \u12_dout_reg[4]/P0001 , \u12_dout_reg[5]/P0001 , \u12_dout_reg[6]/P0001 , \u12_dout_reg[7]/P0001 , \u12_dout_reg[8]/P0001 , \u12_dout_reg[9]/P0001 , \u12_i3_re_reg/NET0131 , \u12_i4_re_reg/P0001 , \u12_i6_re_reg/NET0131 , \u12_o3_we_reg/P0001 , \u12_o4_we_reg/P0001 , \u12_o6_we_reg/P0001 , \u12_o7_we_reg/P0001 , \u12_o8_we_reg/P0001 , \u12_o9_we_reg/P0001 , \u12_re1_reg/P0001 , \u12_re2_reg/NET0131 , \u12_rf_we_reg/P0001 , \u12_we1_reg/P0001 , \u12_we2_reg/P0001 , \u13_ac97_rst_force_reg/P0001 , \u13_crac_dout_r_reg[0]/P0001 , \u13_crac_dout_r_reg[10]/P0001 , \u13_crac_dout_r_reg[11]/P0001 , \u13_crac_dout_r_reg[12]/P0001 , \u13_crac_dout_r_reg[13]/P0001 , \u13_crac_dout_r_reg[14]/P0001 , \u13_crac_dout_r_reg[15]/P0001 , \u13_crac_dout_r_reg[1]/P0001 , \u13_crac_dout_r_reg[2]/P0001 , \u13_crac_dout_r_reg[3]/P0001 , \u13_crac_dout_r_reg[4]/P0001 , \u13_crac_dout_r_reg[5]/P0001 , \u13_crac_dout_r_reg[6]/P0001 , \u13_crac_dout_r_reg[7]/P0001 , \u13_crac_dout_r_reg[8]/P0001 , \u13_crac_dout_r_reg[9]/P0001 , \u13_crac_r_reg[0]/NET0131 , \u13_crac_r_reg[1]/NET0131 , \u13_crac_r_reg[2]/NET0131 , \u13_crac_r_reg[3]/NET0131 , \u13_crac_r_reg[4]/NET0131 , \u13_crac_r_reg[5]/NET0131 , \u13_crac_r_reg[6]/NET0131 , \u13_crac_r_reg[7]/NET0131 , \u13_icc_r_reg[0]/NET0131 , \u13_icc_r_reg[10]/NET0131 , \u13_icc_r_reg[11]/NET0131 , \u13_icc_r_reg[12]/NET0131 , \u13_icc_r_reg[13]/NET0131 , \u13_icc_r_reg[14]/NET0131 , \u13_icc_r_reg[15]/NET0131 , \u13_icc_r_reg[16]/NET0131 , \u13_icc_r_reg[17]/NET0131 , \u13_icc_r_reg[18]/NET0131 , \u13_icc_r_reg[19]/NET0131 , \u13_icc_r_reg[1]/NET0131 , \u13_icc_r_reg[20]/NET0131 , \u13_icc_r_reg[21]/NET0131 , \u13_icc_r_reg[22]/NET0131 , \u13_icc_r_reg[23]/NET0131 , \u13_icc_r_reg[2]/NET0131 , \u13_icc_r_reg[3]/NET0131 , \u13_icc_r_reg[4]/NET0131 , \u13_icc_r_reg[5]/NET0131 , \u13_icc_r_reg[6]/NET0131 , \u13_icc_r_reg[7]/NET0131 , \u13_icc_r_reg[8]/NET0131 , \u13_icc_r_reg[9]/NET0131 , \u13_intm_r_reg[0]/NET0131 , \u13_intm_r_reg[10]/NET0131 , \u13_intm_r_reg[11]/NET0131 , \u13_intm_r_reg[12]/NET0131 , \u13_intm_r_reg[13]/NET0131 , \u13_intm_r_reg[14]/NET0131 , \u13_intm_r_reg[15]/NET0131 , \u13_intm_r_reg[16]/NET0131 , \u13_intm_r_reg[17]/NET0131 , \u13_intm_r_reg[18]/NET0131 , \u13_intm_r_reg[19]/NET0131 , \u13_intm_r_reg[1]/NET0131 , \u13_intm_r_reg[20]/NET0131 , \u13_intm_r_reg[21]/NET0131 , \u13_intm_r_reg[22]/NET0131 , \u13_intm_r_reg[23]/NET0131 , \u13_intm_r_reg[24]/NET0131 , \u13_intm_r_reg[25]/NET0131 , \u13_intm_r_reg[26]/NET0131 , \u13_intm_r_reg[27]/NET0131 , \u13_intm_r_reg[28]/NET0131 , \u13_intm_r_reg[2]/NET0131 , \u13_intm_r_reg[3]/NET0131 , \u13_intm_r_reg[4]/NET0131 , \u13_intm_r_reg[5]/NET0131 , \u13_intm_r_reg[6]/NET0131 , \u13_intm_r_reg[7]/NET0131 , \u13_intm_r_reg[8]/NET0131 , \u13_intm_r_reg[9]/NET0131 , \u13_ints_r_reg[0]/NET0131 , \u13_ints_r_reg[10]/NET0131 , \u13_ints_r_reg[11]/NET0131 , \u13_ints_r_reg[12]/NET0131 , \u13_ints_r_reg[13]/NET0131 , \u13_ints_r_reg[14]/NET0131 , \u13_ints_r_reg[15]/NET0131 , \u13_ints_r_reg[16]/NET0131 , \u13_ints_r_reg[17]/NET0131 , \u13_ints_r_reg[18]/NET0131 , \u13_ints_r_reg[19]/NET0131 , \u13_ints_r_reg[1]/NET0131 , \u13_ints_r_reg[20]/NET0131 , \u13_ints_r_reg[21]/NET0131 , \u13_ints_r_reg[22]/NET0131 , \u13_ints_r_reg[23]/NET0131 , \u13_ints_r_reg[24]/NET0131 , \u13_ints_r_reg[25]/NET0131 , \u13_ints_r_reg[26]/NET0131 , \u13_ints_r_reg[27]/NET0131 , \u13_ints_r_reg[28]/NET0131 , \u13_ints_r_reg[2]/NET0131 , \u13_ints_r_reg[3]/NET0131 , \u13_ints_r_reg[4]/NET0131 , \u13_ints_r_reg[5]/NET0131 , \u13_ints_r_reg[6]/NET0131 , \u13_ints_r_reg[7]/NET0131 , \u13_ints_r_reg[8]/NET0131 , \u13_ints_r_reg[9]/NET0131 , \u13_occ0_r_reg[0]/NET0131 , \u13_occ0_r_reg[10]/NET0131 , \u13_occ0_r_reg[11]/NET0131 , \u13_occ0_r_reg[12]/NET0131 , \u13_occ0_r_reg[13]/NET0131 , \u13_occ0_r_reg[14]/NET0131 , \u13_occ0_r_reg[15]/NET0131 , \u13_occ0_r_reg[16]/NET0131 , \u13_occ0_r_reg[17]/NET0131 , \u13_occ0_r_reg[18]/NET0131 , \u13_occ0_r_reg[19]/NET0131 , \u13_occ0_r_reg[1]/NET0131 , \u13_occ0_r_reg[20]/NET0131 , \u13_occ0_r_reg[21]/NET0131 , \u13_occ0_r_reg[22]/NET0131 , \u13_occ0_r_reg[23]/NET0131 , \u13_occ0_r_reg[24]/NET0131 , \u13_occ0_r_reg[25]/NET0131 , \u13_occ0_r_reg[26]/NET0131 , \u13_occ0_r_reg[27]/NET0131 , \u13_occ0_r_reg[28]/NET0131 , \u13_occ0_r_reg[29]/NET0131 , \u13_occ0_r_reg[2]/NET0131 , \u13_occ0_r_reg[30]/NET0131 , \u13_occ0_r_reg[31]/NET0131 , \u13_occ0_r_reg[3]/NET0131 , \u13_occ0_r_reg[4]/NET0131 , \u13_occ0_r_reg[5]/NET0131 , \u13_occ0_r_reg[6]/NET0131 , \u13_occ0_r_reg[7]/NET0131 , \u13_occ0_r_reg[8]/NET0131 , \u13_occ0_r_reg[9]/NET0131 , \u13_occ1_r_reg[0]/NET0131 , \u13_occ1_r_reg[10]/NET0131 , \u13_occ1_r_reg[11]/NET0131 , \u13_occ1_r_reg[12]/NET0131 , \u13_occ1_r_reg[13]/NET0131 , \u13_occ1_r_reg[14]/NET0131 , \u13_occ1_r_reg[15]/NET0131 , \u13_occ1_r_reg[1]/NET0131 , \u13_occ1_r_reg[2]/NET0131 , \u13_occ1_r_reg[3]/NET0131 , \u13_occ1_r_reg[4]/NET0131 , \u13_occ1_r_reg[5]/NET0131 , \u13_occ1_r_reg[6]/NET0131 , \u13_occ1_r_reg[7]/NET0131 , \u13_occ1_r_reg[8]/NET0131 , \u13_occ1_r_reg[9]/NET0131 , \u13_resume_req_reg/P0001 , \u14_crac_valid_r_reg/P0001 , \u14_crac_wr_r_reg/P0001 , \u14_u0_en_out_l2_reg/P0001 , \u14_u0_en_out_l_reg/NET0131 , \u14_u0_full_empty_r_reg/P0001 , \u14_u1_en_out_l2_reg/P0001 , \u14_u1_en_out_l_reg/NET0131 , \u14_u1_full_empty_r_reg/P0001 , \u14_u2_en_out_l2_reg/P0001 , \u14_u2_en_out_l_reg/NET0131 , \u14_u2_full_empty_r_reg/P0001 , \u14_u3_en_out_l2_reg/P0001 , \u14_u3_en_out_l_reg/NET0131 , \u14_u3_full_empty_r_reg/P0001 , \u14_u4_en_out_l2_reg/P0001 , \u14_u4_en_out_l_reg/NET0131 , \u14_u4_full_empty_r_reg/P0001 , \u14_u5_en_out_l2_reg/P0001 , \u14_u5_en_out_l_reg/NET0131 , \u14_u5_full_empty_r_reg/P0001 , \u14_u6_en_out_l2_reg/P0001 , \u14_u6_en_out_l_reg/NET0131 , \u14_u6_full_empty_r_reg/P0001 , \u14_u7_en_out_l2_reg/P0001 , \u14_u7_en_out_l_reg/NET0131 , \u14_u7_full_empty_r_reg/P0001 , \u14_u8_en_out_l2_reg/P0001 , \u14_u8_en_out_l_reg/NET0131 , \u14_u8_full_empty_r_reg/P0001 , \u15_crac_din_reg[0]/NET0131 , \u15_crac_din_reg[10]/NET0131 , \u15_crac_din_reg[11]/NET0131 , \u15_crac_din_reg[12]/NET0131 , \u15_crac_din_reg[13]/NET0131 , \u15_crac_din_reg[14]/NET0131 , \u15_crac_din_reg[15]/NET0131 , \u15_crac_din_reg[1]/NET0131 , \u15_crac_din_reg[2]/NET0131 , \u15_crac_din_reg[3]/NET0131 , \u15_crac_din_reg[4]/NET0131 , \u15_crac_din_reg[5]/NET0131 , \u15_crac_din_reg[6]/NET0131 , \u15_crac_din_reg[7]/NET0131 , \u15_crac_din_reg[8]/NET0131 , \u15_crac_din_reg[9]/NET0131 , \u15_crac_rd_done_reg/P0001 , \u15_crac_rd_reg/NET0131 , \u15_crac_we_r_reg/P0001 , \u15_crac_wr_reg/NET0131 , \u15_rdd1_reg/NET0131 , \u15_rdd2_reg/NET0131 , \u15_rdd3_reg/NET0131 , \u15_valid_r_reg/P0001 , \u16_u0_dma_req_r1_reg/P0001 , \u16_u1_dma_req_r1_reg/P0001 , \u16_u2_dma_req_r1_reg/P0001 , \u16_u3_dma_req_r1_reg/P0001 , \u16_u4_dma_req_r1_reg/P0001 , \u16_u5_dma_req_r1_reg/P0001 , \u16_u6_dma_req_r1_reg/P0001 , \u16_u7_dma_req_r1_reg/P0001 , \u16_u8_dma_req_r1_reg/P0001 , \u17_int_set_reg[0]/NET0131 , \u17_int_set_reg[1]/NET0131 , \u17_int_set_reg[2]/NET0131 , \u18_int_set_reg[0]/NET0131 , \u18_int_set_reg[1]/NET0131 , \u18_int_set_reg[2]/NET0131 , \u19_int_set_reg[0]/NET0131 , \u19_int_set_reg[1]/NET0131 , \u19_int_set_reg[2]/NET0131 , \u1_slt0_reg[11]/P0001 , \u1_slt0_reg[12]/P0001 , \u1_slt0_reg[15]/P0001 , \u1_slt0_reg[9]/P0001 , \u1_slt1_reg[10]/P0001 , \u1_slt1_reg[11]/P0001 , \u1_slt1_reg[5]/P0001 , \u1_slt1_reg[6]/P0001 , \u1_slt1_reg[7]/P0001 , \u1_slt1_reg[8]/P0001 , \u1_slt3_reg[0]/P0001 , \u1_slt3_reg[10]/P0001 , \u1_slt3_reg[11]/P0001 , \u1_slt3_reg[12]/P0001 , \u1_slt3_reg[13]/P0001 , \u1_slt3_reg[14]/P0001 , \u1_slt3_reg[15]/P0001 , \u1_slt3_reg[16]/P0001 , \u1_slt3_reg[17]/P0001 , \u1_slt3_reg[18]/P0001 , \u1_slt3_reg[19]/P0001 , \u1_slt3_reg[1]/P0001 , \u1_slt3_reg[2]/P0001 , \u1_slt3_reg[3]/P0001 , \u1_slt3_reg[4]/P0001 , \u1_slt3_reg[5]/P0001 , \u1_slt3_reg[6]/P0001 , \u1_slt3_reg[7]/P0001 , \u1_slt3_reg[8]/P0001 , \u1_slt3_reg[9]/P0001 , \u1_slt4_reg[0]/P0001 , \u1_slt4_reg[10]/P0001 , \u1_slt4_reg[11]/P0001 , \u1_slt4_reg[12]/P0001 , \u1_slt4_reg[13]/P0001 , \u1_slt4_reg[14]/P0001 , \u1_slt4_reg[15]/P0001 , \u1_slt4_reg[16]/P0001 , \u1_slt4_reg[17]/P0001 , \u1_slt4_reg[18]/P0001 , \u1_slt4_reg[19]/P0001 , \u1_slt4_reg[1]/P0001 , \u1_slt4_reg[2]/P0001 , \u1_slt4_reg[3]/P0001 , \u1_slt4_reg[4]/P0001 , \u1_slt4_reg[5]/P0001 , \u1_slt4_reg[6]/P0001 , \u1_slt4_reg[7]/P0001 , \u1_slt4_reg[8]/P0001 , \u1_slt4_reg[9]/P0001 , \u1_slt6_reg[0]/P0001 , \u1_slt6_reg[10]/P0001 , \u1_slt6_reg[11]/P0001 , \u1_slt6_reg[12]/P0001 , \u1_slt6_reg[13]/P0001 , \u1_slt6_reg[14]/P0001 , \u1_slt6_reg[15]/P0001 , \u1_slt6_reg[16]/P0001 , \u1_slt6_reg[17]/P0001 , \u1_slt6_reg[18]/P0001 , \u1_slt6_reg[19]/P0001 , \u1_slt6_reg[1]/P0001 , \u1_slt6_reg[2]/P0001 , \u1_slt6_reg[3]/P0001 , \u1_slt6_reg[4]/P0001 , \u1_slt6_reg[5]/P0001 , \u1_slt6_reg[6]/P0001 , \u1_slt6_reg[7]/P0001 , \u1_slt6_reg[8]/P0001 , \u1_slt6_reg[9]/P0001 , \u1_sr_reg[10]/P0001 , \u1_sr_reg[11]/P0001 , \u1_sr_reg[12]/P0001 , \u1_sr_reg[15]/P0001 , \u1_sr_reg[5]/P0001 , \u1_sr_reg[6]/P0001 , \u1_sr_reg[7]/P0001 , \u1_sr_reg[8]/P0001 , \u1_sr_reg[9]/P0001 , \u20_int_set_reg[0]/NET0131 , \u20_int_set_reg[1]/NET0131 , \u20_int_set_reg[2]/NET0131 , \u21_int_set_reg[0]/NET0131 , \u21_int_set_reg[1]/NET0131 , \u21_int_set_reg[2]/NET0131 , \u22_int_set_reg[0]/NET0131 , \u22_int_set_reg[1]/NET0131 , \u22_int_set_reg[2]/NET0131 , \u23_int_set_reg[0]/NET0131 , \u23_int_set_reg[1]/NET0131 , \u23_int_set_reg[2]/NET0131 , \u24_int_set_reg[0]/NET0131 , \u24_int_set_reg[1]/NET0131 , \u24_int_set_reg[2]/NET0131 , \u25_int_set_reg[0]/NET0131 , \u25_int_set_reg[1]/NET0131 , \u25_int_set_reg[2]/NET0131 , \u26_cnt_reg[0]/NET0131 , \u26_cnt_reg[1]/NET0131 , \u26_cnt_reg[2]/NET0131 , \u26_ps_cnt_reg[0]/NET0131 , \u26_ps_cnt_reg[1]/NET0131 , \u26_ps_cnt_reg[2]/NET0131 , \u26_ps_cnt_reg[3]/NET0131 , \u26_ps_cnt_reg[4]/NET0131 , \u26_ps_cnt_reg[5]/NET0131 , \u2_bit_clk_e_reg/P0001 , \u2_bit_clk_r1_reg/P0001 , \u2_bit_clk_r_reg/P0001 , \u2_cnt_reg[0]/NET0131 , \u2_cnt_reg[1]/NET0131 , \u2_cnt_reg[2]/NET0131 , \u2_cnt_reg[3]/NET0131 , \u2_cnt_reg[4]/NET0131 , \u2_cnt_reg[5]/NET0131 , \u2_cnt_reg[6]/NET0131 , \u2_cnt_reg[7]/NET0131 , \u2_ld_reg/P0001 , \u2_out_le_reg[0]/P0001 , \u2_out_le_reg[1]/P0001 , \u2_res_cnt_reg[0]/P0001 , \u2_res_cnt_reg[1]/P0001 , \u2_res_cnt_reg[2]/P0001 , \u2_res_cnt_reg[3]/P0001 , \u2_sync_beat_reg/P0001 , \u2_sync_resume_reg/NET0131 , \u2_to_cnt_reg[0]/NET0131 , \u2_to_cnt_reg[1]/NET0131 , \u2_to_cnt_reg[2]/NET0131 , \u2_to_cnt_reg[3]/NET0131 , \u2_to_cnt_reg[4]/NET0131 , \u2_to_cnt_reg[5]/NET0131 , \u3_dout_reg[0]/P0001 , \u3_dout_reg[10]/P0001 , \u3_dout_reg[11]/P0001 , \u3_dout_reg[12]/P0001 , \u3_dout_reg[13]/P0001 , \u3_dout_reg[14]/P0001 , \u3_dout_reg[15]/P0001 , \u3_dout_reg[16]/P0001 , \u3_dout_reg[17]/P0001 , \u3_dout_reg[18]/P0001 , \u3_dout_reg[19]/P0001 , \u3_dout_reg[1]/P0001 , \u3_dout_reg[2]/P0001 , \u3_dout_reg[3]/P0001 , \u3_dout_reg[4]/P0001 , \u3_dout_reg[5]/P0001 , \u3_dout_reg[6]/P0001 , \u3_dout_reg[7]/P0001 , \u3_dout_reg[8]/P0001 , \u3_dout_reg[9]/P0001 , \u3_empty_reg/NET0131 , \u3_mem_reg[0][0]/NET0131 , \u3_mem_reg[0][10]/NET0131 , \u3_mem_reg[0][11]/NET0131 , \u3_mem_reg[0][12]/NET0131 , \u3_mem_reg[0][13]/NET0131 , \u3_mem_reg[0][14]/NET0131 , \u3_mem_reg[0][15]/NET0131 , \u3_mem_reg[0][16]/NET0131 , \u3_mem_reg[0][17]/NET0131 , \u3_mem_reg[0][18]/NET0131 , \u3_mem_reg[0][19]/NET0131 , \u3_mem_reg[0][1]/NET0131 , \u3_mem_reg[0][20]/NET0131 , \u3_mem_reg[0][21]/NET0131 , \u3_mem_reg[0][22]/NET0131 , \u3_mem_reg[0][23]/NET0131 , \u3_mem_reg[0][24]/NET0131 , \u3_mem_reg[0][25]/NET0131 , \u3_mem_reg[0][26]/NET0131 , \u3_mem_reg[0][27]/NET0131 , \u3_mem_reg[0][28]/NET0131 , \u3_mem_reg[0][29]/NET0131 , \u3_mem_reg[0][2]/NET0131 , \u3_mem_reg[0][30]/NET0131 , \u3_mem_reg[0][31]/NET0131 , \u3_mem_reg[0][3]/NET0131 , \u3_mem_reg[0][4]/NET0131 , \u3_mem_reg[0][5]/NET0131 , \u3_mem_reg[0][6]/NET0131 , \u3_mem_reg[0][7]/NET0131 , \u3_mem_reg[0][8]/NET0131 , \u3_mem_reg[0][9]/NET0131 , \u3_mem_reg[1][0]/NET0131 , \u3_mem_reg[1][10]/NET0131 , \u3_mem_reg[1][11]/NET0131 , \u3_mem_reg[1][12]/NET0131 , \u3_mem_reg[1][13]/NET0131 , \u3_mem_reg[1][14]/NET0131 , \u3_mem_reg[1][15]/NET0131 , \u3_mem_reg[1][16]/NET0131 , \u3_mem_reg[1][17]/NET0131 , \u3_mem_reg[1][18]/NET0131 , \u3_mem_reg[1][19]/NET0131 , \u3_mem_reg[1][1]/NET0131 , \u3_mem_reg[1][20]/NET0131 , \u3_mem_reg[1][21]/NET0131 , \u3_mem_reg[1][22]/NET0131 , \u3_mem_reg[1][23]/NET0131 , \u3_mem_reg[1][24]/NET0131 , \u3_mem_reg[1][25]/NET0131 , \u3_mem_reg[1][26]/NET0131 , \u3_mem_reg[1][27]/NET0131 , \u3_mem_reg[1][28]/NET0131 , \u3_mem_reg[1][29]/NET0131 , \u3_mem_reg[1][2]/NET0131 , \u3_mem_reg[1][30]/NET0131 , \u3_mem_reg[1][31]/NET0131 , \u3_mem_reg[1][3]/NET0131 , \u3_mem_reg[1][4]/NET0131 , \u3_mem_reg[1][5]/NET0131 , \u3_mem_reg[1][6]/NET0131 , \u3_mem_reg[1][7]/NET0131 , \u3_mem_reg[1][8]/NET0131 , \u3_mem_reg[1][9]/NET0131 , \u3_mem_reg[2][0]/NET0131 , \u3_mem_reg[2][10]/NET0131 , \u3_mem_reg[2][11]/NET0131 , \u3_mem_reg[2][12]/NET0131 , \u3_mem_reg[2][13]/NET0131 , \u3_mem_reg[2][14]/NET0131 , \u3_mem_reg[2][15]/NET0131 , \u3_mem_reg[2][16]/NET0131 , \u3_mem_reg[2][17]/NET0131 , \u3_mem_reg[2][18]/NET0131 , \u3_mem_reg[2][19]/NET0131 , \u3_mem_reg[2][1]/NET0131 , \u3_mem_reg[2][20]/NET0131 , \u3_mem_reg[2][21]/NET0131 , \u3_mem_reg[2][22]/NET0131 , \u3_mem_reg[2][23]/NET0131 , \u3_mem_reg[2][24]/NET0131 , \u3_mem_reg[2][25]/NET0131 , \u3_mem_reg[2][26]/NET0131 , \u3_mem_reg[2][27]/NET0131 , \u3_mem_reg[2][28]/NET0131 , \u3_mem_reg[2][29]/NET0131 , \u3_mem_reg[2][2]/NET0131 , \u3_mem_reg[2][30]/NET0131 , \u3_mem_reg[2][31]/NET0131 , \u3_mem_reg[2][3]/NET0131 , \u3_mem_reg[2][4]/NET0131 , \u3_mem_reg[2][5]/NET0131 , \u3_mem_reg[2][6]/NET0131 , \u3_mem_reg[2][7]/NET0131 , \u3_mem_reg[2][8]/NET0131 , \u3_mem_reg[2][9]/NET0131 , \u3_mem_reg[3][0]/NET0131 , \u3_mem_reg[3][10]/NET0131 , \u3_mem_reg[3][11]/NET0131 , \u3_mem_reg[3][12]/NET0131 , \u3_mem_reg[3][13]/NET0131 , \u3_mem_reg[3][14]/NET0131 , \u3_mem_reg[3][15]/NET0131 , \u3_mem_reg[3][16]/NET0131 , \u3_mem_reg[3][17]/NET0131 , \u3_mem_reg[3][18]/NET0131 , \u3_mem_reg[3][19]/NET0131 , \u3_mem_reg[3][1]/NET0131 , \u3_mem_reg[3][20]/NET0131 , \u3_mem_reg[3][21]/NET0131 , \u3_mem_reg[3][22]/NET0131 , \u3_mem_reg[3][23]/NET0131 , \u3_mem_reg[3][24]/NET0131 , \u3_mem_reg[3][25]/NET0131 , \u3_mem_reg[3][26]/NET0131 , \u3_mem_reg[3][27]/NET0131 , \u3_mem_reg[3][28]/NET0131 , \u3_mem_reg[3][29]/NET0131 , \u3_mem_reg[3][2]/NET0131 , \u3_mem_reg[3][30]/NET0131 , \u3_mem_reg[3][31]/NET0131 , \u3_mem_reg[3][3]/NET0131 , \u3_mem_reg[3][4]/NET0131 , \u3_mem_reg[3][5]/NET0131 , \u3_mem_reg[3][6]/NET0131 , \u3_mem_reg[3][7]/NET0131 , \u3_mem_reg[3][8]/NET0131 , \u3_mem_reg[3][9]/NET0131 , \u3_rp_reg[0]/P0001 , \u3_rp_reg[1]/NET0131 , \u3_rp_reg[2]/NET0131 , \u3_rp_reg[3]/NET0131 , \u3_status_reg[0]/P0001 , \u3_status_reg[1]/P0001 , \u3_wp_reg[0]/P0001 , \u3_wp_reg[1]/NET0131 , \u3_wp_reg[2]/P0001 , \u4_dout_reg[0]/P0001 , \u4_dout_reg[10]/P0001 , \u4_dout_reg[11]/P0001 , \u4_dout_reg[12]/P0001 , \u4_dout_reg[13]/P0001 , \u4_dout_reg[14]/P0001 , \u4_dout_reg[15]/P0001 , \u4_dout_reg[16]/P0001 , \u4_dout_reg[17]/P0001 , \u4_dout_reg[18]/P0001 , \u4_dout_reg[19]/P0001 , \u4_dout_reg[1]/P0001 , \u4_dout_reg[2]/P0001 , \u4_dout_reg[3]/P0001 , \u4_dout_reg[4]/P0001 , \u4_dout_reg[5]/P0001 , \u4_dout_reg[6]/P0001 , \u4_dout_reg[7]/P0001 , \u4_dout_reg[8]/P0001 , \u4_dout_reg[9]/P0001 , \u4_empty_reg/NET0131 , \u4_mem_reg[0][0]/NET0131 , \u4_mem_reg[0][10]/NET0131 , \u4_mem_reg[0][11]/NET0131 , \u4_mem_reg[0][12]/NET0131 , \u4_mem_reg[0][13]/NET0131 , \u4_mem_reg[0][14]/NET0131 , \u4_mem_reg[0][15]/NET0131 , \u4_mem_reg[0][16]/NET0131 , \u4_mem_reg[0][17]/NET0131 , \u4_mem_reg[0][18]/NET0131 , \u4_mem_reg[0][19]/NET0131 , \u4_mem_reg[0][1]/NET0131 , \u4_mem_reg[0][20]/NET0131 , \u4_mem_reg[0][21]/NET0131 , \u4_mem_reg[0][22]/NET0131 , \u4_mem_reg[0][23]/NET0131 , \u4_mem_reg[0][24]/NET0131 , \u4_mem_reg[0][25]/NET0131 , \u4_mem_reg[0][26]/NET0131 , \u4_mem_reg[0][27]/NET0131 , \u4_mem_reg[0][28]/NET0131 , \u4_mem_reg[0][29]/NET0131 , \u4_mem_reg[0][2]/NET0131 , \u4_mem_reg[0][30]/NET0131 , \u4_mem_reg[0][31]/NET0131 , \u4_mem_reg[0][3]/NET0131 , \u4_mem_reg[0][4]/NET0131 , \u4_mem_reg[0][5]/NET0131 , \u4_mem_reg[0][6]/NET0131 , \u4_mem_reg[0][7]/NET0131 , \u4_mem_reg[0][8]/NET0131 , \u4_mem_reg[0][9]/NET0131 , \u4_mem_reg[1][0]/NET0131 , \u4_mem_reg[1][10]/NET0131 , \u4_mem_reg[1][11]/NET0131 , \u4_mem_reg[1][12]/NET0131 , \u4_mem_reg[1][13]/NET0131 , \u4_mem_reg[1][14]/NET0131 , \u4_mem_reg[1][15]/NET0131 , \u4_mem_reg[1][16]/NET0131 , \u4_mem_reg[1][17]/NET0131 , \u4_mem_reg[1][18]/NET0131 , \u4_mem_reg[1][19]/NET0131 , \u4_mem_reg[1][1]/NET0131 , \u4_mem_reg[1][20]/NET0131 , \u4_mem_reg[1][21]/NET0131 , \u4_mem_reg[1][22]/NET0131 , \u4_mem_reg[1][23]/NET0131 , \u4_mem_reg[1][24]/NET0131 , \u4_mem_reg[1][25]/NET0131 , \u4_mem_reg[1][26]/NET0131 , \u4_mem_reg[1][27]/NET0131 , \u4_mem_reg[1][28]/NET0131 , \u4_mem_reg[1][29]/NET0131 , \u4_mem_reg[1][2]/NET0131 , \u4_mem_reg[1][30]/NET0131 , \u4_mem_reg[1][31]/NET0131 , \u4_mem_reg[1][3]/NET0131 , \u4_mem_reg[1][4]/NET0131 , \u4_mem_reg[1][5]/NET0131 , \u4_mem_reg[1][6]/NET0131 , \u4_mem_reg[1][7]/NET0131 , \u4_mem_reg[1][8]/NET0131 , \u4_mem_reg[1][9]/NET0131 , \u4_mem_reg[2][0]/NET0131 , \u4_mem_reg[2][10]/NET0131 , \u4_mem_reg[2][11]/NET0131 , \u4_mem_reg[2][12]/NET0131 , \u4_mem_reg[2][13]/NET0131 , \u4_mem_reg[2][14]/NET0131 , \u4_mem_reg[2][15]/NET0131 , \u4_mem_reg[2][16]/NET0131 , \u4_mem_reg[2][17]/NET0131 , \u4_mem_reg[2][18]/NET0131 , \u4_mem_reg[2][19]/NET0131 , \u4_mem_reg[2][1]/NET0131 , \u4_mem_reg[2][20]/NET0131 , \u4_mem_reg[2][21]/NET0131 , \u4_mem_reg[2][22]/NET0131 , \u4_mem_reg[2][23]/NET0131 , \u4_mem_reg[2][24]/NET0131 , \u4_mem_reg[2][25]/NET0131 , \u4_mem_reg[2][26]/NET0131 , \u4_mem_reg[2][27]/NET0131 , \u4_mem_reg[2][28]/NET0131 , \u4_mem_reg[2][29]/NET0131 , \u4_mem_reg[2][2]/NET0131 , \u4_mem_reg[2][30]/NET0131 , \u4_mem_reg[2][31]/NET0131 , \u4_mem_reg[2][3]/NET0131 , \u4_mem_reg[2][4]/NET0131 , \u4_mem_reg[2][5]/NET0131 , \u4_mem_reg[2][6]/NET0131 , \u4_mem_reg[2][7]/NET0131 , \u4_mem_reg[2][8]/NET0131 , \u4_mem_reg[2][9]/NET0131 , \u4_mem_reg[3][0]/NET0131 , \u4_mem_reg[3][10]/NET0131 , \u4_mem_reg[3][11]/NET0131 , \u4_mem_reg[3][12]/NET0131 , \u4_mem_reg[3][13]/NET0131 , \u4_mem_reg[3][14]/NET0131 , \u4_mem_reg[3][15]/NET0131 , \u4_mem_reg[3][16]/NET0131 , \u4_mem_reg[3][17]/NET0131 , \u4_mem_reg[3][18]/NET0131 , \u4_mem_reg[3][19]/NET0131 , \u4_mem_reg[3][1]/NET0131 , \u4_mem_reg[3][20]/NET0131 , \u4_mem_reg[3][21]/NET0131 , \u4_mem_reg[3][22]/NET0131 , \u4_mem_reg[3][23]/NET0131 , \u4_mem_reg[3][24]/NET0131 , \u4_mem_reg[3][25]/NET0131 , \u4_mem_reg[3][26]/NET0131 , \u4_mem_reg[3][27]/NET0131 , \u4_mem_reg[3][28]/NET0131 , \u4_mem_reg[3][29]/NET0131 , \u4_mem_reg[3][2]/NET0131 , \u4_mem_reg[3][30]/NET0131 , \u4_mem_reg[3][31]/NET0131 , \u4_mem_reg[3][3]/NET0131 , \u4_mem_reg[3][4]/NET0131 , \u4_mem_reg[3][5]/NET0131 , \u4_mem_reg[3][6]/NET0131 , \u4_mem_reg[3][7]/NET0131 , \u4_mem_reg[3][8]/NET0131 , \u4_mem_reg[3][9]/NET0131 , \u4_rp_reg[0]/P0001 , \u4_rp_reg[1]/NET0131 , \u4_rp_reg[2]/NET0131 , \u4_rp_reg[3]/NET0131 , \u4_status_reg[0]/P0001 , \u4_status_reg[1]/P0001 , \u4_wp_reg[0]/P0001 , \u4_wp_reg[1]/NET0131 , \u4_wp_reg[2]/P0001 , \u5_dout_reg[0]/P0001 , \u5_dout_reg[10]/P0001 , \u5_dout_reg[11]/P0001 , \u5_dout_reg[12]/P0001 , \u5_dout_reg[13]/P0001 , \u5_dout_reg[14]/P0001 , \u5_dout_reg[15]/P0001 , \u5_dout_reg[16]/P0001 , \u5_dout_reg[17]/P0001 , \u5_dout_reg[18]/P0001 , \u5_dout_reg[19]/P0001 , \u5_dout_reg[1]/P0001 , \u5_dout_reg[2]/P0001 , \u5_dout_reg[3]/P0001 , \u5_dout_reg[4]/P0001 , \u5_dout_reg[5]/P0001 , \u5_dout_reg[6]/P0001 , \u5_dout_reg[7]/P0001 , \u5_dout_reg[8]/P0001 , \u5_dout_reg[9]/P0001 , \u5_empty_reg/NET0131 , \u5_mem_reg[0][0]/NET0131 , \u5_mem_reg[0][10]/NET0131 , \u5_mem_reg[0][11]/NET0131 , \u5_mem_reg[0][12]/NET0131 , \u5_mem_reg[0][13]/NET0131 , \u5_mem_reg[0][14]/NET0131 , \u5_mem_reg[0][15]/NET0131 , \u5_mem_reg[0][16]/NET0131 , \u5_mem_reg[0][17]/NET0131 , \u5_mem_reg[0][18]/NET0131 , \u5_mem_reg[0][19]/NET0131 , \u5_mem_reg[0][1]/NET0131 , \u5_mem_reg[0][20]/NET0131 , \u5_mem_reg[0][21]/NET0131 , \u5_mem_reg[0][22]/NET0131 , \u5_mem_reg[0][23]/NET0131 , \u5_mem_reg[0][24]/NET0131 , \u5_mem_reg[0][25]/NET0131 , \u5_mem_reg[0][26]/NET0131 , \u5_mem_reg[0][27]/NET0131 , \u5_mem_reg[0][28]/NET0131 , \u5_mem_reg[0][29]/NET0131 , \u5_mem_reg[0][2]/NET0131 , \u5_mem_reg[0][30]/NET0131 , \u5_mem_reg[0][31]/NET0131 , \u5_mem_reg[0][3]/NET0131 , \u5_mem_reg[0][4]/NET0131 , \u5_mem_reg[0][5]/NET0131 , \u5_mem_reg[0][6]/NET0131 , \u5_mem_reg[0][7]/NET0131 , \u5_mem_reg[0][8]/NET0131 , \u5_mem_reg[0][9]/NET0131 , \u5_mem_reg[1][0]/NET0131 , \u5_mem_reg[1][10]/NET0131 , \u5_mem_reg[1][11]/NET0131 , \u5_mem_reg[1][12]/NET0131 , \u5_mem_reg[1][13]/NET0131 , \u5_mem_reg[1][14]/NET0131 , \u5_mem_reg[1][15]/NET0131 , \u5_mem_reg[1][16]/NET0131 , \u5_mem_reg[1][17]/NET0131 , \u5_mem_reg[1][18]/NET0131 , \u5_mem_reg[1][19]/NET0131 , \u5_mem_reg[1][1]/NET0131 , \u5_mem_reg[1][20]/NET0131 , \u5_mem_reg[1][21]/NET0131 , \u5_mem_reg[1][22]/NET0131 , \u5_mem_reg[1][23]/NET0131 , \u5_mem_reg[1][24]/NET0131 , \u5_mem_reg[1][25]/NET0131 , \u5_mem_reg[1][26]/NET0131 , \u5_mem_reg[1][27]/NET0131 , \u5_mem_reg[1][28]/NET0131 , \u5_mem_reg[1][29]/NET0131 , \u5_mem_reg[1][2]/NET0131 , \u5_mem_reg[1][30]/NET0131 , \u5_mem_reg[1][31]/NET0131 , \u5_mem_reg[1][3]/NET0131 , \u5_mem_reg[1][4]/NET0131 , \u5_mem_reg[1][5]/NET0131 , \u5_mem_reg[1][6]/NET0131 , \u5_mem_reg[1][7]/NET0131 , \u5_mem_reg[1][8]/NET0131 , \u5_mem_reg[1][9]/NET0131 , \u5_mem_reg[2][0]/NET0131 , \u5_mem_reg[2][10]/NET0131 , \u5_mem_reg[2][11]/NET0131 , \u5_mem_reg[2][12]/NET0131 , \u5_mem_reg[2][13]/NET0131 , \u5_mem_reg[2][14]/NET0131 , \u5_mem_reg[2][15]/NET0131 , \u5_mem_reg[2][16]/NET0131 , \u5_mem_reg[2][17]/NET0131 , \u5_mem_reg[2][18]/NET0131 , \u5_mem_reg[2][19]/NET0131 , \u5_mem_reg[2][1]/NET0131 , \u5_mem_reg[2][20]/NET0131 , \u5_mem_reg[2][21]/NET0131 , \u5_mem_reg[2][22]/NET0131 , \u5_mem_reg[2][23]/NET0131 , \u5_mem_reg[2][24]/NET0131 , \u5_mem_reg[2][25]/NET0131 , \u5_mem_reg[2][26]/NET0131 , \u5_mem_reg[2][27]/NET0131 , \u5_mem_reg[2][28]/NET0131 , \u5_mem_reg[2][29]/NET0131 , \u5_mem_reg[2][2]/NET0131 , \u5_mem_reg[2][30]/NET0131 , \u5_mem_reg[2][31]/NET0131 , \u5_mem_reg[2][3]/NET0131 , \u5_mem_reg[2][4]/NET0131 , \u5_mem_reg[2][5]/NET0131 , \u5_mem_reg[2][6]/NET0131 , \u5_mem_reg[2][7]/NET0131 , \u5_mem_reg[2][8]/NET0131 , \u5_mem_reg[2][9]/NET0131 , \u5_mem_reg[3][0]/NET0131 , \u5_mem_reg[3][10]/NET0131 , \u5_mem_reg[3][11]/NET0131 , \u5_mem_reg[3][12]/NET0131 , \u5_mem_reg[3][13]/NET0131 , \u5_mem_reg[3][14]/NET0131 , \u5_mem_reg[3][15]/NET0131 , \u5_mem_reg[3][16]/NET0131 , \u5_mem_reg[3][17]/NET0131 , \u5_mem_reg[3][18]/NET0131 , \u5_mem_reg[3][19]/NET0131 , \u5_mem_reg[3][1]/NET0131 , \u5_mem_reg[3][20]/NET0131 , \u5_mem_reg[3][21]/NET0131 , \u5_mem_reg[3][22]/NET0131 , \u5_mem_reg[3][23]/NET0131 , \u5_mem_reg[3][24]/NET0131 , \u5_mem_reg[3][25]/NET0131 , \u5_mem_reg[3][26]/NET0131 , \u5_mem_reg[3][27]/NET0131 , \u5_mem_reg[3][28]/NET0131 , \u5_mem_reg[3][29]/NET0131 , \u5_mem_reg[3][2]/NET0131 , \u5_mem_reg[3][30]/NET0131 , \u5_mem_reg[3][31]/NET0131 , \u5_mem_reg[3][3]/NET0131 , \u5_mem_reg[3][4]/NET0131 , \u5_mem_reg[3][5]/NET0131 , \u5_mem_reg[3][6]/NET0131 , \u5_mem_reg[3][7]/NET0131 , \u5_mem_reg[3][8]/NET0131 , \u5_mem_reg[3][9]/NET0131 , \u5_rp_reg[0]/P0001 , \u5_rp_reg[1]/NET0131 , \u5_rp_reg[2]/NET0131 , \u5_rp_reg[3]/NET0131 , \u5_status_reg[0]/P0001 , \u5_status_reg[1]/P0001 , \u5_wp_reg[0]/P0001 , \u5_wp_reg[1]/NET0131 , \u5_wp_reg[2]/P0001 , \u6_dout_reg[0]/P0001 , \u6_dout_reg[10]/P0001 , \u6_dout_reg[11]/P0001 , \u6_dout_reg[12]/P0001 , \u6_dout_reg[13]/P0001 , \u6_dout_reg[14]/P0001 , \u6_dout_reg[15]/P0001 , \u6_dout_reg[16]/P0001 , \u6_dout_reg[17]/P0001 , \u6_dout_reg[18]/P0001 , \u6_dout_reg[19]/P0001 , \u6_dout_reg[1]/P0001 , \u6_dout_reg[2]/P0001 , \u6_dout_reg[3]/P0001 , \u6_dout_reg[4]/P0001 , \u6_dout_reg[5]/P0001 , \u6_dout_reg[6]/P0001 , \u6_dout_reg[7]/P0001 , \u6_dout_reg[8]/P0001 , \u6_dout_reg[9]/P0001 , \u6_empty_reg/NET0131 , \u6_mem_reg[0][0]/NET0131 , \u6_mem_reg[0][10]/NET0131 , \u6_mem_reg[0][11]/NET0131 , \u6_mem_reg[0][12]/NET0131 , \u6_mem_reg[0][13]/NET0131 , \u6_mem_reg[0][14]/NET0131 , \u6_mem_reg[0][15]/NET0131 , \u6_mem_reg[0][16]/NET0131 , \u6_mem_reg[0][17]/NET0131 , \u6_mem_reg[0][18]/NET0131 , \u6_mem_reg[0][19]/NET0131 , \u6_mem_reg[0][1]/NET0131 , \u6_mem_reg[0][20]/NET0131 , \u6_mem_reg[0][21]/NET0131 , \u6_mem_reg[0][22]/NET0131 , \u6_mem_reg[0][23]/NET0131 , \u6_mem_reg[0][24]/NET0131 , \u6_mem_reg[0][25]/NET0131 , \u6_mem_reg[0][26]/NET0131 , \u6_mem_reg[0][27]/NET0131 , \u6_mem_reg[0][28]/NET0131 , \u6_mem_reg[0][29]/NET0131 , \u6_mem_reg[0][2]/NET0131 , \u6_mem_reg[0][30]/NET0131 , \u6_mem_reg[0][31]/NET0131 , \u6_mem_reg[0][3]/NET0131 , \u6_mem_reg[0][4]/NET0131 , \u6_mem_reg[0][5]/NET0131 , \u6_mem_reg[0][6]/NET0131 , \u6_mem_reg[0][7]/NET0131 , \u6_mem_reg[0][8]/NET0131 , \u6_mem_reg[0][9]/NET0131 , \u6_mem_reg[1][0]/NET0131 , \u6_mem_reg[1][10]/NET0131 , \u6_mem_reg[1][11]/NET0131 , \u6_mem_reg[1][12]/NET0131 , \u6_mem_reg[1][13]/NET0131 , \u6_mem_reg[1][14]/NET0131 , \u6_mem_reg[1][15]/NET0131 , \u6_mem_reg[1][16]/NET0131 , \u6_mem_reg[1][17]/NET0131 , \u6_mem_reg[1][18]/NET0131 , \u6_mem_reg[1][19]/NET0131 , \u6_mem_reg[1][1]/NET0131 , \u6_mem_reg[1][20]/NET0131 , \u6_mem_reg[1][21]/NET0131 , \u6_mem_reg[1][22]/NET0131 , \u6_mem_reg[1][23]/NET0131 , \u6_mem_reg[1][24]/NET0131 , \u6_mem_reg[1][25]/NET0131 , \u6_mem_reg[1][26]/NET0131 , \u6_mem_reg[1][27]/NET0131 , \u6_mem_reg[1][28]/NET0131 , \u6_mem_reg[1][29]/NET0131 , \u6_mem_reg[1][2]/NET0131 , \u6_mem_reg[1][30]/NET0131 , \u6_mem_reg[1][31]/NET0131 , \u6_mem_reg[1][3]/NET0131 , \u6_mem_reg[1][4]/NET0131 , \u6_mem_reg[1][5]/NET0131 , \u6_mem_reg[1][6]/NET0131 , \u6_mem_reg[1][7]/NET0131 , \u6_mem_reg[1][8]/NET0131 , \u6_mem_reg[1][9]/NET0131 , \u6_mem_reg[2][0]/NET0131 , \u6_mem_reg[2][10]/NET0131 , \u6_mem_reg[2][11]/NET0131 , \u6_mem_reg[2][12]/NET0131 , \u6_mem_reg[2][13]/NET0131 , \u6_mem_reg[2][14]/NET0131 , \u6_mem_reg[2][15]/NET0131 , \u6_mem_reg[2][16]/NET0131 , \u6_mem_reg[2][17]/NET0131 , \u6_mem_reg[2][18]/NET0131 , \u6_mem_reg[2][19]/NET0131 , \u6_mem_reg[2][1]/NET0131 , \u6_mem_reg[2][20]/NET0131 , \u6_mem_reg[2][21]/NET0131 , \u6_mem_reg[2][22]/NET0131 , \u6_mem_reg[2][23]/NET0131 , \u6_mem_reg[2][24]/NET0131 , \u6_mem_reg[2][25]/NET0131 , \u6_mem_reg[2][26]/NET0131 , \u6_mem_reg[2][27]/NET0131 , \u6_mem_reg[2][28]/NET0131 , \u6_mem_reg[2][29]/NET0131 , \u6_mem_reg[2][2]/NET0131 , \u6_mem_reg[2][30]/NET0131 , \u6_mem_reg[2][31]/NET0131 , \u6_mem_reg[2][3]/NET0131 , \u6_mem_reg[2][4]/NET0131 , \u6_mem_reg[2][5]/NET0131 , \u6_mem_reg[2][6]/NET0131 , \u6_mem_reg[2][7]/NET0131 , \u6_mem_reg[2][8]/NET0131 , \u6_mem_reg[2][9]/NET0131 , \u6_mem_reg[3][0]/NET0131 , \u6_mem_reg[3][10]/NET0131 , \u6_mem_reg[3][11]/NET0131 , \u6_mem_reg[3][12]/NET0131 , \u6_mem_reg[3][13]/NET0131 , \u6_mem_reg[3][14]/NET0131 , \u6_mem_reg[3][15]/NET0131 , \u6_mem_reg[3][16]/NET0131 , \u6_mem_reg[3][17]/NET0131 , \u6_mem_reg[3][18]/NET0131 , \u6_mem_reg[3][19]/NET0131 , \u6_mem_reg[3][1]/NET0131 , \u6_mem_reg[3][20]/NET0131 , \u6_mem_reg[3][21]/NET0131 , \u6_mem_reg[3][22]/NET0131 , \u6_mem_reg[3][23]/NET0131 , \u6_mem_reg[3][24]/NET0131 , \u6_mem_reg[3][25]/NET0131 , \u6_mem_reg[3][26]/NET0131 , \u6_mem_reg[3][27]/NET0131 , \u6_mem_reg[3][28]/NET0131 , \u6_mem_reg[3][29]/NET0131 , \u6_mem_reg[3][2]/NET0131 , \u6_mem_reg[3][30]/NET0131 , \u6_mem_reg[3][31]/NET0131 , \u6_mem_reg[3][3]/NET0131 , \u6_mem_reg[3][4]/NET0131 , \u6_mem_reg[3][5]/NET0131 , \u6_mem_reg[3][6]/NET0131 , \u6_mem_reg[3][7]/NET0131 , \u6_mem_reg[3][8]/NET0131 , \u6_mem_reg[3][9]/NET0131 , \u6_rp_reg[0]/P0001 , \u6_rp_reg[1]/NET0131 , \u6_rp_reg[2]/NET0131 , \u6_rp_reg[3]/NET0131 , \u6_status_reg[0]/P0001 , \u6_status_reg[1]/P0001 , \u6_wp_reg[0]/P0001 , \u6_wp_reg[1]/NET0131 , \u6_wp_reg[2]/P0001 , \u7_dout_reg[0]/P0001 , \u7_dout_reg[10]/P0001 , \u7_dout_reg[11]/P0001 , \u7_dout_reg[12]/P0001 , \u7_dout_reg[13]/P0001 , \u7_dout_reg[14]/P0001 , \u7_dout_reg[15]/P0001 , \u7_dout_reg[16]/P0001 , \u7_dout_reg[17]/P0001 , \u7_dout_reg[18]/P0001 , \u7_dout_reg[19]/P0001 , \u7_dout_reg[1]/P0001 , \u7_dout_reg[2]/P0001 , \u7_dout_reg[3]/P0001 , \u7_dout_reg[4]/P0001 , \u7_dout_reg[5]/P0001 , \u7_dout_reg[6]/P0001 , \u7_dout_reg[7]/P0001 , \u7_dout_reg[8]/P0001 , \u7_dout_reg[9]/P0001 , \u7_empty_reg/NET0131 , \u7_mem_reg[0][0]/NET0131 , \u7_mem_reg[0][10]/NET0131 , \u7_mem_reg[0][11]/NET0131 , \u7_mem_reg[0][12]/NET0131 , \u7_mem_reg[0][13]/NET0131 , \u7_mem_reg[0][14]/NET0131 , \u7_mem_reg[0][15]/NET0131 , \u7_mem_reg[0][16]/NET0131 , \u7_mem_reg[0][17]/NET0131 , \u7_mem_reg[0][18]/NET0131 , \u7_mem_reg[0][19]/NET0131 , \u7_mem_reg[0][1]/NET0131 , \u7_mem_reg[0][20]/NET0131 , \u7_mem_reg[0][21]/NET0131 , \u7_mem_reg[0][22]/NET0131 , \u7_mem_reg[0][23]/NET0131 , \u7_mem_reg[0][24]/NET0131 , \u7_mem_reg[0][25]/NET0131 , \u7_mem_reg[0][26]/NET0131 , \u7_mem_reg[0][27]/NET0131 , \u7_mem_reg[0][28]/NET0131 , \u7_mem_reg[0][29]/NET0131 , \u7_mem_reg[0][2]/NET0131 , \u7_mem_reg[0][30]/NET0131 , \u7_mem_reg[0][31]/NET0131 , \u7_mem_reg[0][3]/NET0131 , \u7_mem_reg[0][4]/NET0131 , \u7_mem_reg[0][5]/NET0131 , \u7_mem_reg[0][6]/NET0131 , \u7_mem_reg[0][7]/NET0131 , \u7_mem_reg[0][8]/NET0131 , \u7_mem_reg[0][9]/NET0131 , \u7_mem_reg[1][0]/NET0131 , \u7_mem_reg[1][10]/NET0131 , \u7_mem_reg[1][11]/NET0131 , \u7_mem_reg[1][12]/NET0131 , \u7_mem_reg[1][13]/NET0131 , \u7_mem_reg[1][14]/NET0131 , \u7_mem_reg[1][15]/NET0131 , \u7_mem_reg[1][16]/NET0131 , \u7_mem_reg[1][17]/NET0131 , \u7_mem_reg[1][18]/NET0131 , \u7_mem_reg[1][19]/NET0131 , \u7_mem_reg[1][1]/NET0131 , \u7_mem_reg[1][20]/NET0131 , \u7_mem_reg[1][21]/NET0131 , \u7_mem_reg[1][22]/NET0131 , \u7_mem_reg[1][23]/NET0131 , \u7_mem_reg[1][24]/NET0131 , \u7_mem_reg[1][25]/NET0131 , \u7_mem_reg[1][26]/NET0131 , \u7_mem_reg[1][27]/NET0131 , \u7_mem_reg[1][28]/NET0131 , \u7_mem_reg[1][29]/NET0131 , \u7_mem_reg[1][2]/NET0131 , \u7_mem_reg[1][30]/NET0131 , \u7_mem_reg[1][31]/NET0131 , \u7_mem_reg[1][3]/NET0131 , \u7_mem_reg[1][4]/NET0131 , \u7_mem_reg[1][5]/NET0131 , \u7_mem_reg[1][6]/NET0131 , \u7_mem_reg[1][7]/NET0131 , \u7_mem_reg[1][8]/NET0131 , \u7_mem_reg[1][9]/NET0131 , \u7_mem_reg[2][0]/NET0131 , \u7_mem_reg[2][10]/NET0131 , \u7_mem_reg[2][11]/NET0131 , \u7_mem_reg[2][12]/NET0131 , \u7_mem_reg[2][13]/NET0131 , \u7_mem_reg[2][14]/NET0131 , \u7_mem_reg[2][15]/NET0131 , \u7_mem_reg[2][16]/NET0131 , \u7_mem_reg[2][17]/NET0131 , \u7_mem_reg[2][18]/NET0131 , \u7_mem_reg[2][19]/NET0131 , \u7_mem_reg[2][1]/NET0131 , \u7_mem_reg[2][20]/NET0131 , \u7_mem_reg[2][21]/NET0131 , \u7_mem_reg[2][22]/NET0131 , \u7_mem_reg[2][23]/NET0131 , \u7_mem_reg[2][24]/NET0131 , \u7_mem_reg[2][25]/NET0131 , \u7_mem_reg[2][26]/NET0131 , \u7_mem_reg[2][27]/NET0131 , \u7_mem_reg[2][28]/NET0131 , \u7_mem_reg[2][29]/NET0131 , \u7_mem_reg[2][2]/NET0131 , \u7_mem_reg[2][30]/NET0131 , \u7_mem_reg[2][31]/NET0131 , \u7_mem_reg[2][3]/NET0131 , \u7_mem_reg[2][4]/NET0131 , \u7_mem_reg[2][5]/NET0131 , \u7_mem_reg[2][6]/NET0131 , \u7_mem_reg[2][7]/NET0131 , \u7_mem_reg[2][8]/NET0131 , \u7_mem_reg[2][9]/NET0131 , \u7_mem_reg[3][0]/NET0131 , \u7_mem_reg[3][10]/NET0131 , \u7_mem_reg[3][11]/NET0131 , \u7_mem_reg[3][12]/NET0131 , \u7_mem_reg[3][13]/NET0131 , \u7_mem_reg[3][14]/NET0131 , \u7_mem_reg[3][15]/NET0131 , \u7_mem_reg[3][16]/NET0131 , \u7_mem_reg[3][17]/NET0131 , \u7_mem_reg[3][18]/NET0131 , \u7_mem_reg[3][19]/NET0131 , \u7_mem_reg[3][1]/NET0131 , \u7_mem_reg[3][20]/NET0131 , \u7_mem_reg[3][21]/NET0131 , \u7_mem_reg[3][22]/NET0131 , \u7_mem_reg[3][23]/NET0131 , \u7_mem_reg[3][24]/NET0131 , \u7_mem_reg[3][25]/NET0131 , \u7_mem_reg[3][26]/NET0131 , \u7_mem_reg[3][27]/NET0131 , \u7_mem_reg[3][28]/NET0131 , \u7_mem_reg[3][29]/NET0131 , \u7_mem_reg[3][2]/NET0131 , \u7_mem_reg[3][30]/NET0131 , \u7_mem_reg[3][31]/NET0131 , \u7_mem_reg[3][3]/NET0131 , \u7_mem_reg[3][4]/NET0131 , \u7_mem_reg[3][5]/NET0131 , \u7_mem_reg[3][6]/NET0131 , \u7_mem_reg[3][7]/NET0131 , \u7_mem_reg[3][8]/NET0131 , \u7_mem_reg[3][9]/NET0131 , \u7_rp_reg[0]/P0001 , \u7_rp_reg[1]/NET0131 , \u7_rp_reg[2]/NET0131 , \u7_rp_reg[3]/NET0131 , \u7_status_reg[0]/P0001 , \u7_status_reg[1]/P0001 , \u7_wp_reg[0]/P0001 , \u7_wp_reg[1]/NET0131 , \u7_wp_reg[2]/P0001 , \u8_dout_reg[0]/P0001 , \u8_dout_reg[10]/P0001 , \u8_dout_reg[11]/P0001 , \u8_dout_reg[12]/P0001 , \u8_dout_reg[13]/P0001 , \u8_dout_reg[14]/P0001 , \u8_dout_reg[15]/P0001 , \u8_dout_reg[16]/P0001 , \u8_dout_reg[17]/P0001 , \u8_dout_reg[18]/P0001 , \u8_dout_reg[19]/P0001 , \u8_dout_reg[1]/P0001 , \u8_dout_reg[2]/P0001 , \u8_dout_reg[3]/P0001 , \u8_dout_reg[4]/P0001 , \u8_dout_reg[5]/P0001 , \u8_dout_reg[6]/P0001 , \u8_dout_reg[7]/P0001 , \u8_dout_reg[8]/P0001 , \u8_dout_reg[9]/P0001 , \u8_empty_reg/NET0131 , \u8_mem_reg[0][0]/NET0131 , \u8_mem_reg[0][10]/NET0131 , \u8_mem_reg[0][11]/NET0131 , \u8_mem_reg[0][12]/NET0131 , \u8_mem_reg[0][13]/NET0131 , \u8_mem_reg[0][14]/NET0131 , \u8_mem_reg[0][15]/NET0131 , \u8_mem_reg[0][16]/NET0131 , \u8_mem_reg[0][17]/NET0131 , \u8_mem_reg[0][18]/NET0131 , \u8_mem_reg[0][19]/NET0131 , \u8_mem_reg[0][1]/NET0131 , \u8_mem_reg[0][20]/NET0131 , \u8_mem_reg[0][21]/NET0131 , \u8_mem_reg[0][22]/NET0131 , \u8_mem_reg[0][23]/NET0131 , \u8_mem_reg[0][24]/NET0131 , \u8_mem_reg[0][25]/NET0131 , \u8_mem_reg[0][26]/NET0131 , \u8_mem_reg[0][27]/NET0131 , \u8_mem_reg[0][28]/NET0131 , \u8_mem_reg[0][29]/NET0131 , \u8_mem_reg[0][2]/NET0131 , \u8_mem_reg[0][30]/NET0131 , \u8_mem_reg[0][31]/NET0131 , \u8_mem_reg[0][3]/NET0131 , \u8_mem_reg[0][4]/NET0131 , \u8_mem_reg[0][5]/NET0131 , \u8_mem_reg[0][6]/NET0131 , \u8_mem_reg[0][7]/NET0131 , \u8_mem_reg[0][8]/NET0131 , \u8_mem_reg[0][9]/NET0131 , \u8_mem_reg[1][0]/NET0131 , \u8_mem_reg[1][10]/NET0131 , \u8_mem_reg[1][11]/NET0131 , \u8_mem_reg[1][12]/NET0131 , \u8_mem_reg[1][13]/NET0131 , \u8_mem_reg[1][14]/NET0131 , \u8_mem_reg[1][15]/NET0131 , \u8_mem_reg[1][16]/NET0131 , \u8_mem_reg[1][17]/NET0131 , \u8_mem_reg[1][18]/NET0131 , \u8_mem_reg[1][19]/NET0131 , \u8_mem_reg[1][1]/NET0131 , \u8_mem_reg[1][20]/NET0131 , \u8_mem_reg[1][21]/NET0131 , \u8_mem_reg[1][22]/NET0131 , \u8_mem_reg[1][23]/NET0131 , \u8_mem_reg[1][24]/NET0131 , \u8_mem_reg[1][25]/NET0131 , \u8_mem_reg[1][26]/NET0131 , \u8_mem_reg[1][27]/NET0131 , \u8_mem_reg[1][28]/NET0131 , \u8_mem_reg[1][29]/NET0131 , \u8_mem_reg[1][2]/NET0131 , \u8_mem_reg[1][30]/NET0131 , \u8_mem_reg[1][31]/NET0131 , \u8_mem_reg[1][3]/NET0131 , \u8_mem_reg[1][4]/NET0131 , \u8_mem_reg[1][5]/NET0131 , \u8_mem_reg[1][6]/NET0131 , \u8_mem_reg[1][7]/NET0131 , \u8_mem_reg[1][8]/NET0131 , \u8_mem_reg[1][9]/NET0131 , \u8_mem_reg[2][0]/NET0131 , \u8_mem_reg[2][10]/NET0131 , \u8_mem_reg[2][11]/NET0131 , \u8_mem_reg[2][12]/NET0131 , \u8_mem_reg[2][13]/NET0131 , \u8_mem_reg[2][14]/NET0131 , \u8_mem_reg[2][15]/NET0131 , \u8_mem_reg[2][16]/NET0131 , \u8_mem_reg[2][17]/NET0131 , \u8_mem_reg[2][18]/NET0131 , \u8_mem_reg[2][19]/NET0131 , \u8_mem_reg[2][1]/NET0131 , \u8_mem_reg[2][20]/NET0131 , \u8_mem_reg[2][21]/NET0131 , \u8_mem_reg[2][22]/NET0131 , \u8_mem_reg[2][23]/NET0131 , \u8_mem_reg[2][24]/NET0131 , \u8_mem_reg[2][25]/NET0131 , \u8_mem_reg[2][26]/NET0131 , \u8_mem_reg[2][27]/NET0131 , \u8_mem_reg[2][28]/NET0131 , \u8_mem_reg[2][29]/NET0131 , \u8_mem_reg[2][2]/NET0131 , \u8_mem_reg[2][30]/NET0131 , \u8_mem_reg[2][31]/NET0131 , \u8_mem_reg[2][3]/NET0131 , \u8_mem_reg[2][4]/NET0131 , \u8_mem_reg[2][5]/NET0131 , \u8_mem_reg[2][6]/NET0131 , \u8_mem_reg[2][7]/NET0131 , \u8_mem_reg[2][8]/NET0131 , \u8_mem_reg[2][9]/NET0131 , \u8_mem_reg[3][0]/NET0131 , \u8_mem_reg[3][10]/NET0131 , \u8_mem_reg[3][11]/NET0131 , \u8_mem_reg[3][12]/NET0131 , \u8_mem_reg[3][13]/NET0131 , \u8_mem_reg[3][14]/NET0131 , \u8_mem_reg[3][15]/NET0131 , \u8_mem_reg[3][16]/NET0131 , \u8_mem_reg[3][17]/NET0131 , \u8_mem_reg[3][18]/NET0131 , \u8_mem_reg[3][19]/NET0131 , \u8_mem_reg[3][1]/NET0131 , \u8_mem_reg[3][20]/NET0131 , \u8_mem_reg[3][21]/NET0131 , \u8_mem_reg[3][22]/NET0131 , \u8_mem_reg[3][23]/NET0131 , \u8_mem_reg[3][24]/NET0131 , \u8_mem_reg[3][25]/NET0131 , \u8_mem_reg[3][26]/NET0131 , \u8_mem_reg[3][27]/NET0131 , \u8_mem_reg[3][28]/NET0131 , \u8_mem_reg[3][29]/NET0131 , \u8_mem_reg[3][2]/NET0131 , \u8_mem_reg[3][30]/NET0131 , \u8_mem_reg[3][31]/NET0131 , \u8_mem_reg[3][3]/NET0131 , \u8_mem_reg[3][4]/NET0131 , \u8_mem_reg[3][5]/NET0131 , \u8_mem_reg[3][6]/NET0131 , \u8_mem_reg[3][7]/NET0131 , \u8_mem_reg[3][8]/NET0131 , \u8_mem_reg[3][9]/NET0131 , \u8_rp_reg[0]/P0001 , \u8_rp_reg[1]/NET0131 , \u8_rp_reg[2]/NET0131 , \u8_rp_reg[3]/NET0131 , \u8_status_reg[0]/P0001 , \u8_status_reg[1]/P0001 , \u8_wp_reg[0]/P0001 , \u8_wp_reg[1]/NET0131 , \u8_wp_reg[2]/P0001 , \u9_din_tmp1_reg[0]/P0001 , \u9_din_tmp1_reg[10]/P0001 , \u9_din_tmp1_reg[11]/P0001 , \u9_din_tmp1_reg[12]/P0001 , \u9_din_tmp1_reg[13]/P0001 , \u9_din_tmp1_reg[14]/P0001 , \u9_din_tmp1_reg[15]/P0001 , \u9_din_tmp1_reg[1]/P0001 , \u9_din_tmp1_reg[2]/P0001 , \u9_din_tmp1_reg[3]/P0001 , \u9_din_tmp1_reg[4]/P0001 , \u9_din_tmp1_reg[5]/P0001 , \u9_din_tmp1_reg[6]/P0001 , \u9_din_tmp1_reg[7]/P0001 , \u9_din_tmp1_reg[8]/P0001 , \u9_din_tmp1_reg[9]/P0001 , \u9_dout_reg[0]/P0001 , \u9_dout_reg[10]/P0001 , \u9_dout_reg[11]/P0001 , \u9_dout_reg[12]/P0001 , \u9_dout_reg[13]/P0001 , \u9_dout_reg[14]/P0001 , \u9_dout_reg[15]/P0001 , \u9_dout_reg[16]/P0001 , \u9_dout_reg[17]/P0001 , \u9_dout_reg[18]/P0001 , \u9_dout_reg[19]/P0001 , \u9_dout_reg[1]/P0001 , \u9_dout_reg[20]/P0001 , \u9_dout_reg[21]/P0001 , \u9_dout_reg[22]/P0001 , \u9_dout_reg[23]/P0001 , \u9_dout_reg[24]/P0001 , \u9_dout_reg[25]/P0001 , \u9_dout_reg[26]/P0001 , \u9_dout_reg[27]/P0001 , \u9_dout_reg[28]/P0001 , \u9_dout_reg[29]/P0001 , \u9_dout_reg[2]/P0001 , \u9_dout_reg[30]/P0001 , \u9_dout_reg[31]/P0001 , \u9_dout_reg[3]/P0001 , \u9_dout_reg[4]/P0001 , \u9_dout_reg[5]/P0001 , \u9_dout_reg[6]/P0001 , \u9_dout_reg[7]/P0001 , \u9_dout_reg[8]/P0001 , \u9_dout_reg[9]/P0001 , \u9_empty_reg/P0001 , \u9_full_reg/NET0131 , \u9_mem_reg[0][0]/P0001 , \u9_mem_reg[0][10]/P0001 , \u9_mem_reg[0][11]/P0001 , \u9_mem_reg[0][12]/P0001 , \u9_mem_reg[0][13]/P0001 , \u9_mem_reg[0][14]/P0001 , \u9_mem_reg[0][15]/P0001 , \u9_mem_reg[0][16]/P0001 , \u9_mem_reg[0][17]/P0001 , \u9_mem_reg[0][18]/P0001 , \u9_mem_reg[0][19]/P0001 , \u9_mem_reg[0][1]/P0001 , \u9_mem_reg[0][20]/P0001 , \u9_mem_reg[0][21]/P0001 , \u9_mem_reg[0][22]/P0001 , \u9_mem_reg[0][23]/P0001 , \u9_mem_reg[0][24]/P0001 , \u9_mem_reg[0][25]/P0001 , \u9_mem_reg[0][26]/P0001 , \u9_mem_reg[0][27]/P0001 , \u9_mem_reg[0][28]/P0001 , \u9_mem_reg[0][29]/P0001 , \u9_mem_reg[0][2]/P0001 , \u9_mem_reg[0][30]/P0001 , \u9_mem_reg[0][31]/P0001 , \u9_mem_reg[0][3]/P0001 , \u9_mem_reg[0][4]/P0001 , \u9_mem_reg[0][5]/P0001 , \u9_mem_reg[0][6]/P0001 , \u9_mem_reg[0][7]/P0001 , \u9_mem_reg[0][8]/P0001 , \u9_mem_reg[0][9]/P0001 , \u9_mem_reg[1][0]/P0001 , \u9_mem_reg[1][10]/P0001 , \u9_mem_reg[1][11]/P0001 , \u9_mem_reg[1][12]/P0001 , \u9_mem_reg[1][13]/P0001 , \u9_mem_reg[1][14]/P0001 , \u9_mem_reg[1][15]/P0001 , \u9_mem_reg[1][16]/P0001 , \u9_mem_reg[1][17]/P0001 , \u9_mem_reg[1][18]/P0001 , \u9_mem_reg[1][19]/P0001 , \u9_mem_reg[1][1]/P0001 , \u9_mem_reg[1][20]/P0001 , \u9_mem_reg[1][21]/P0001 , \u9_mem_reg[1][22]/P0001 , \u9_mem_reg[1][23]/P0001 , \u9_mem_reg[1][24]/P0001 , \u9_mem_reg[1][25]/P0001 , \u9_mem_reg[1][26]/P0001 , \u9_mem_reg[1][27]/P0001 , \u9_mem_reg[1][28]/P0001 , \u9_mem_reg[1][29]/P0001 , \u9_mem_reg[1][2]/P0001 , \u9_mem_reg[1][30]/P0001 , \u9_mem_reg[1][31]/P0001 , \u9_mem_reg[1][3]/P0001 , \u9_mem_reg[1][4]/P0001 , \u9_mem_reg[1][5]/P0001 , \u9_mem_reg[1][6]/P0001 , \u9_mem_reg[1][7]/P0001 , \u9_mem_reg[1][8]/P0001 , \u9_mem_reg[1][9]/P0001 , \u9_mem_reg[2][0]/P0001 , \u9_mem_reg[2][10]/P0001 , \u9_mem_reg[2][11]/P0001 , \u9_mem_reg[2][12]/P0001 , \u9_mem_reg[2][13]/P0001 , \u9_mem_reg[2][14]/P0001 , \u9_mem_reg[2][15]/P0001 , \u9_mem_reg[2][16]/P0001 , \u9_mem_reg[2][17]/P0001 , \u9_mem_reg[2][18]/P0001 , \u9_mem_reg[2][19]/P0001 , \u9_mem_reg[2][1]/P0001 , \u9_mem_reg[2][20]/P0001 , \u9_mem_reg[2][21]/P0001 , \u9_mem_reg[2][22]/P0001 , \u9_mem_reg[2][23]/P0001 , \u9_mem_reg[2][24]/P0001 , \u9_mem_reg[2][25]/P0001 , \u9_mem_reg[2][26]/P0001 , \u9_mem_reg[2][27]/P0001 , \u9_mem_reg[2][28]/P0001 , \u9_mem_reg[2][29]/P0001 , \u9_mem_reg[2][2]/P0001 , \u9_mem_reg[2][30]/P0001 , \u9_mem_reg[2][31]/P0001 , \u9_mem_reg[2][3]/P0001 , \u9_mem_reg[2][4]/P0001 , \u9_mem_reg[2][5]/P0001 , \u9_mem_reg[2][6]/P0001 , \u9_mem_reg[2][7]/P0001 , \u9_mem_reg[2][8]/P0001 , \u9_mem_reg[2][9]/P0001 , \u9_mem_reg[3][0]/P0001 , \u9_mem_reg[3][10]/P0001 , \u9_mem_reg[3][11]/P0001 , \u9_mem_reg[3][12]/P0001 , \u9_mem_reg[3][13]/P0001 , \u9_mem_reg[3][14]/P0001 , \u9_mem_reg[3][15]/P0001 , \u9_mem_reg[3][16]/P0001 , \u9_mem_reg[3][17]/P0001 , \u9_mem_reg[3][18]/P0001 , \u9_mem_reg[3][19]/P0001 , \u9_mem_reg[3][1]/P0001 , \u9_mem_reg[3][20]/P0001 , \u9_mem_reg[3][21]/P0001 , \u9_mem_reg[3][22]/P0001 , \u9_mem_reg[3][23]/P0001 , \u9_mem_reg[3][24]/P0001 , \u9_mem_reg[3][25]/P0001 , \u9_mem_reg[3][26]/P0001 , \u9_mem_reg[3][27]/P0001 , \u9_mem_reg[3][28]/P0001 , \u9_mem_reg[3][29]/P0001 , \u9_mem_reg[3][2]/P0001 , \u9_mem_reg[3][30]/P0001 , \u9_mem_reg[3][31]/P0001 , \u9_mem_reg[3][3]/P0001 , \u9_mem_reg[3][4]/P0001 , \u9_mem_reg[3][5]/P0001 , \u9_mem_reg[3][6]/P0001 , \u9_mem_reg[3][7]/P0001 , \u9_mem_reg[3][8]/P0001 , \u9_mem_reg[3][9]/P0001 , \u9_rp_reg[0]/P0001 , \u9_rp_reg[1]/P0001 , \u9_rp_reg[2]/P0001 , \u9_status_reg[0]/P0001 , \u9_status_reg[1]/P0001 , \u9_wp_reg[0]/NET0131 , \u9_wp_reg[1]/P0001 , \u9_wp_reg[2]/P0001 , \u9_wp_reg[3]/P0001 , \valid_s_reg/NET0131 , wb_ack_o_pad, \wb_addr_i[29]_pad , \wb_addr_i[2]_pad , \wb_addr_i[30]_pad , \wb_addr_i[31]_pad , \wb_addr_i[3]_pad , \wb_addr_i[4]_pad , \wb_addr_i[5]_pad , \wb_addr_i[6]_pad , wb_cyc_i_pad, wb_stb_i_pad, wb_we_i_pad, \_al_n1 , \g16/_0_ , \g23/_0_ , \g29500/_0_ , \g29503/_3_ , \g29505/_3_ , \g29507/_3_ , \g29509/_3_ , \g29511/_0_ , \g29513/_3_ , \g29515/_3_ , \g29517/_3_ , \g29519/_0_ , \g29522/_0_ , \g29524/_0_ , \g29526/_0_ , \g29528/_0_ , \g29530/_0_ , \g29532/_0_ , \g29534/_3_ , \g29536/_3_ , \g29538/_3_ , \g29540/_3_ , \g29542/_3_ , \g29544/_3_ , \g29546/_3_ , \g29548/_3_ , \g29550/_0_ , \g29552/_0_ , \g29554/_0_ , \g29556/_0_ , \g29558/_0_ , \g29560/_0_ , \g29562/_0_ , \g29564/_0_ , \g29566/_0_ , \g29568/_0_ , \g29570/_0_ , \g29572/_0_ , \g29574/_3_ , \g29576/_3_ , \g29578/_3_ , \g29580/_3_ , \g29582/_3_ , \g29584/_3_ , \g29586/_3_ , \g29588/_3_ , \g29590/_3_ , \g29592/_3_ , \g29594/_3_ , \g29596/_3_ , \g29598/_3_ , \g29600/_3_ , \g29602/_3_ , \g29604/_3_ , \g29606/_0_ , \g29608/_0_ , \g29610/_0_ , \g29612/_0_ , \g29614/_3_ , \g29616/_3_ , \g29618/_3_ , \g29620/_3_ , \g29622/_3_ , \g29624/_3_ , \g29626/_3_ , \g29628/_3_ , \g29630/_3_ , \g29632/_3_ , \g29634/_3_ , \g29636/_3_ , \g29638/_3_ , \g29640/_3_ , \g29642/_3_ , \g29644/_3_ , \g29646/_3_ , \g29648/_3_ , \g29650/_3_ , \g29652/_3_ , \g29654/_3_ , \g29656/_3_ , \g29658/_3_ , \g29660/_3_ , \g29662/_3_ , \g29664/_3_ , \g29666/_3_ , \g29668/_3_ , \g29670/_3_ , \g29672/_3_ , \g29674/_3_ , \g29676/_3_ , \g29678/_3_ , \g29680/_3_ , \g29682/_3_ , \g29684/_3_ , \g29686/_3_ , \g29688/_3_ , \g29690/_3_ , \g29692/_3_ , \g29694/_0_ , \g29696/_0_ , \g29698/_0_ , \g29700/_0_ , \g29702/_0_ , \g29704/_0_ , \g29706/_0_ , \g29708/_0_ , \g29710/_0_ , \g29712/_0_ , \g29714/_0_ , \g29716/_0_ , \g29718/_0_ , \g29720/_0_ , \g29722/_0_ , \g29724/_0_ , \g29726/_0_ , \g29728/_0_ , \g29730/_0_ , \g29732/_0_ , \g29734/_3_ , \g29736/_3_ , \g29738/_3_ , \g29740/_3_ , \g29742/_3_ , \g29744/_3_ , \g29746/_3_ , \g29748/_3_ , \g29750/_3_ , \g29752/_3_ , \g29754/_3_ , \g29756/_3_ , \g29758/_3_ , \g29760/_3_ , \g29762/_3_ , \g29764/_3_ , \g29766/_3_ , \g29768/_3_ , \g29770/_3_ , \g29772/_3_ , \g29774/_3_ , \g29776/_3_ , \g29778/_3_ , \g29780/_3_ , \g29782/_3_ , \g29784/_3_ , \g29786/_3_ , \g29788/_3_ , \g29790/_3_ , \g29792/_3_ , \g29794/_3_ , \g29796/_3_ , \g29798/_3_ , \g29800/_3_ , \g29802/_3_ , \g29804/_3_ , \g29806/_3_ , \g29808/_3_ , \g29810/_3_ , \g29812/_3_ , \g29814/_3_ , \g29816/_3_ , \g29818/_3_ , \g29820/_3_ , \g29822/_3_ , \g29824/_3_ , \g29826/_3_ , \g29828/_3_ , \g29830/_3_ , \g29832/_3_ , \g29834/_3_ , \g29836/_3_ , \g29838/_3_ , \g29840/_3_ , \g29842/_3_ , \g29844/_3_ , \g29846/_3_ , \g29848/_3_ , \g29850/_3_ , \g29852/_3_ , \g29854/_3_ , \g29856/_3_ , \g29858/_3_ , \g29860/_3_ , \g29862/_3_ , \g29864/_3_ , \g29866/_3_ , \g29868/_3_ , \g29870/_3_ , \g29872/_3_ , \g29874/_3_ , \g29876/_3_ , \g29878/_3_ , \g29880/_3_ , \g29904/_0_ , \g29905/_0_ , \g29906/_0_ , \g29907/_0_ , \g29908/_0_ , \g29909/_0_ , \g29914/_3_ , \g29952/_0_ , \g29953/_0_ , \g29954/_0_ , \g29955/_0_ , \g29956/_0_ , \g29957/_0_ , \g29975/_0_ , \g29976/_0_ , \g29977/_0_ , \g29978/_0_ , \g29979/_0_ , \g29980/_0_ , \g29989/_3_ , \g30020/_0_ , \g30021/_0_ , \g30045/_0_ , \g30046/_0_ , \g30047/_0_ , \g30048/_0_ , \g30049/_0_ , \g30050/_0_ , \g30051/_0_ , \g30052/_0_ , \g30053/_0_ , \g30054/_0_ , \g30062/_0_ , \g30063/_0_ , \g30064/_0_ , \g30065/_0_ , \g30066/_0_ , \g30067/_0_ , \g30068/_0_ , \g30069/_0_ , \g30070/_0_ , \g30071/_0_ , \g30072/_0_ , \g30073/_0_ , \g30074/_0_ , \g30075/_0_ , \g30136/_3_ , \g30707/_0_ , \g30708/_0_ , \g30711/_0_ , \g30714/_0_ , \g30715/_0_ , \g30720/_0_ , \g30725/_0_ , \g30741/_0_ , \g30742/_0_ , \g30743/_0_ , \g30744/_0_ , \g30745/_0_ , \g30746/_0_ , \g30747/_0_ , \g30748/_0_ , \g30749/_0_ , \g30750/_0_ , \g30751/_0_ , \g30752/_0_ , \g30789/_0_ , \g30790/_0_ , \g30791/_0_ , \g30792/_0_ , \g30793/_0_ , \g30794/_0_ , \g30795/_0_ , \g30796/_0_ , \g30797/_0_ , \g30798/_0_ , \g30799/_0_ , \g30800/_0_ , \g30801/_0_ , \g30802/_0_ , \g30803/_0_ , \g30804/_0_ , \g30805/_0_ , \g30806/_0_ , \g30807/_0_ , \g30808/_0_ , \g30809/_0_ , \g30810/_0_ , \g30811/_0_ , \g30812/_0_ , \g30813/_0_ , \g30814/_0_ , \g30815/_0_ , \g30816/_0_ , \g30817/_0_ , \g30818/_0_ , \g30819/_0_ , \g30820/_0_ , \g30821/_0_ , \g30822/_0_ , \g30823/_0_ , \g30824/_0_ , \g30825/_0_ , \g30826/_0_ , \g30827/_0_ , \g30828/_0_ , \g30829/_0_ , \g30830/_0_ , \g30831/_0_ , \g30832/_0_ , \g30833/_0_ , \g30834/_0_ , \g30835/_0_ , \g30836/_0_ , \g30837/_0_ , \g30838/_0_ , \g30839/_0_ , \g30840/_0_ , \g30841/_0_ , \g30842/_0_ , \g30843/_0_ , \g30844/_0_ , \g30845/_0_ , \g30846/_0_ , \g30847/_0_ , \g30848/_0_ , \g30849/_0_ , \g30850/_0_ , \g30851/_0_ , \g30852/_0_ , \g30853/_0_ , \g30854/_0_ , \g30855/_0_ , \g30856/_0_ , \g30857/_0_ , \g30858/_0_ , \g30859/_0_ , \g30860/_0_ , \g30861/_0_ , \g30862/_0_ , \g30863/_0_ , \g30864/_0_ , \g30865/_0_ , \g30866/_0_ , \g30867/_0_ , \g30868/_0_ , \g30869/_0_ , \g30870/_0_ , \g30871/_0_ , \g30872/_0_ , \g30873/_0_ , \g30874/_0_ , \g30875/_0_ , \g30876/_0_ , \g30877/_0_ , \g30878/_0_ , \g30879/_0_ , \g30880/_0_ , \g30881/_0_ , \g30882/_0_ , \g30883/_0_ , \g30884/_0_ , \g30885/_0_ , \g30886/_0_ , \g30887/_0_ , \g30888/_0_ , \g30889/_0_ , \g30890/_0_ , \g30891/_0_ , \g30892/_0_ , \g30893/_0_ , \g30894/_0_ , \g30895/_0_ , \g30896/_0_ , \g30897/_0_ , \g30898/_0_ , \g30899/_0_ , \g30900/_0_ , \g30901/_0_ , \g30902/_0_ , \g30906/_0_ , \g30907/_0_ , \g30908/_0_ , \g30909/_0_ , \g30910/_0_ , \g30911/_0_ , \g30918/_0_ , \g30919/_0_ , \g30920/_0_ , \g30921/_0_ , \g30922/_0_ , \g30923/_0_ , \g30924/_0_ , \g30925/_0_ , \g30926/_0_ , \g30946/_0_ , \g30947/_0_ , \g30948/_0_ , \g30949/_0_ , \g30950/_0_ , \g30951/_0_ , \g30952/_0_ , \g30953/_0_ , \g30954/_0_ , \g30955/_0_ , \g30956/_0_ , \g30957/_0_ , \g30958/_0_ , \g30959/_0_ , \g30960/_0_ , \g30961/_0_ , \g30962/_0_ , \g30963/_0_ , \g30964/_0_ , \g30965/_0_ , \g30966/_0_ , \g30967/_0_ , \g30968/_0_ , \g30969/_0_ , \g30970/_0_ , \g30971/_0_ , \g30972/_0_ , \g30973/_0_ , \g30974/_0_ , \g30975/_0_ , \g30976/_0_ , \g30977/_0_ , \g30978/_0_ , \g30979/_0_ , \g30980/_0_ , \g30981/_0_ , \g30982/_0_ , \g30983/_0_ , \g30984/_0_ , \g30985/_0_ , \g30986/_0_ , \g30987/_0_ , \g30988/_0_ , \g30989/_0_ , \g30990/_0_ , \g30991/_0_ , \g30992/_0_ , \g30993/_0_ , \g30994/_0_ , \g30995/_0_ , \g30996/_0_ , \g30997/_0_ , \g30998/_0_ , \g30999/_0_ , \g31000/_0_ , \g31001/_0_ , \g31002/_0_ , \g31003/_0_ , \g31004/_0_ , \g31005/_0_ , \g31006/_0_ , \g31007/_0_ , \g31008/_0_ , \g31009/_0_ , \g31010/_0_ , \g31011/_0_ , \g31012/_0_ , \g31013/_0_ , \g31014/_0_ , \g31015/_0_ , \g31016/_0_ , \g31017/_0_ , \g31018/_0_ , \g31019/_0_ , \g31020/_0_ , \g31021/_0_ , \g31022/_0_ , \g31023/_0_ , \g31024/_0_ , \g31025/_0_ , \g31026/_0_ , \g31027/_0_ , \g31028/_0_ , \g31029/_0_ , \g31030/_0_ , \g31031/_0_ , \g31032/_0_ , \g31033/_0_ , \g31034/_0_ , \g31035/_0_ , \g31036/_0_ , \g31037/_0_ , \g31038/_0_ , \g31039/_0_ , \g31040/_0_ , \g31041/_0_ , \g31042/_0_ , \g31043/_0_ , \g31044/_0_ , \g31045/_0_ , \g31046/_0_ , \g31047/_0_ , \g31048/_0_ , \g31049/_0_ , \g31050/_0_ , \g31051/_0_ , \g31052/_0_ , \g31053/_0_ , \g31054/_0_ , \g31055/_0_ , \g31056/_0_ , \g31057/_0_ , \g31058/_0_ , \g31059/_0_ , \g31060/_0_ , \g31061/_0_ , \g31062/_0_ , \g31063/_0_ , \g31064/_0_ , \g31065/_0_ , \g31066/_0_ , \g31067/_0_ , \g31068/_0_ , \g31069/_0_ , \g31070/_0_ , \g31071/_0_ , \g31072/_0_ , \g31073/_0_ , \g31074/_0_ , \g31075/_0_ , \g31076/_0_ , \g31077/_0_ , \g31084/u3_syn_4 , \g31085/u3_syn_4 , \g31096/u3_syn_4 , \g31115/u3_syn_4 , \g31136/u3_syn_4 , \g31158/u3_syn_4 , \g31176/u3_syn_4 , \g31193/u3_syn_4 , \g31195/u3_syn_4 , \g31247/u3_syn_4 , \g31280/u3_syn_4 , \g31285/u3_syn_4 , \g31568/_0_ , \g31631/_0_ , \g31672/_0_ , \g31731/_0_ , \g31732/_0_ , \g31742/_2_ , \g31744/_2_ , \g31746/_2_ , \g31748/_2_ , \g31751/_2_ , \g31754/_2_ , \g31756/_2_ , \g31758/_2_ , \g31760/_2_ , \g31761/_0_ , \g31789/_0_ , \g31807/_3_ , \g31825/_3_ , \g32607/_0_ , \g32608/_0_ , \g32609/_0_ , \g32610/_0_ , \g32611/_0_ , \g32612/_0_ , \g32613/_0_ , \g32614/_0_ , \g32615/_0_ , \g32616/_0_ , \g32617/_0_ , \g32618/_0_ , \g32645/_0__syn_2 , \g32687/_0__syn_2 , \g32749/_0__syn_2 , \g32757/_0_ , \g32758/_0_ , \g32759/_0_ , \g32760/_0_ , \g32761/_0_ , \g32762/_0_ , \g32763/_0_ , \g32764/_0_ , \g32765/_0_ , \g32769/_0_ , \g32835/_1_ , \g32839/_0_ , \g32844/_0_ , \g32901/_1_ , \g32902/_0_ , \g32963/_1_ , \g32972/_0_ , \g32977/_0_ , \g32979/_0_ , \g32980/_0_ , \g32981/_0_ , \g32982/_0_ , \g32983/_0_ , \g32987/_0_ , \g33018/_0_ , \g33019/_0_ , \g33088/_0_ , \g33261/_0_ , \g33264/_0_ , \g33275/_0_ , \g33276/_0_ , \g33277/_0_ , \g33371/_0_ , \g33382/_0_ , \g33401/_0_ , \g33402/_0_ , \g33403/_0_ , \g33404/_0_ , \g33405/_0_ , \g33406/_0_ , \g33407/_0_ , \g33408/_0_ , \g33409/_0_ , \g33410/_0_ , \g33411/_0_ , \g33412/_0_ , \g33413/_0_ , \g33414/_0_ , \g33415/_0_ , \g33416/_0_ , \g33417/_0_ , \g33418/_0_ , \g33419/_0_ , \g33420/_0_ , \g33421/_0_ , \g33422/_0_ , \g33423/_0_ , \g33424/_0_ , \g33425/_0_ , \g33426/_0_ , \g33427/_0_ , \g33428/_0_ , \g33429/_0_ , \g33430/_0_ , \g33431/_0_ , \g33432/_0_ , \g33433/_0_ , \g33434/_0_ , \g33435/_0_ , \g33436/_0_ , \g33437/_0_ , \g33438/_0_ , \g33439/_0_ , \g33440/_0_ , \g33441/_0_ , \g33442/_0_ , \g33443/_0_ , \g33444/_0_ , \g33445/_0_ , \g33446/_0_ , \g33447/_0_ , \g33448/_0_ , \g33449/_0_ , \g33450/_0_ , \g33451/_0_ , \g33452/_0_ , \g33453/_0_ , \g33454/_0_ , \g33455/_0_ , \g33456/_0_ , \g33457/_0_ , \g33458/_0_ , \g33459/_0_ , \g33460/_0_ , \g33461/_0_ , \g33462/_0_ , \g33463/_0_ , \g33464/_0_ , \g33465/_0_ , \g33466/_0_ , \g33467/_0_ , \g33468/_0_ , \g33469/_0_ , \g33470/_0_ , \g33471/_0_ , \g33472/_0_ , \g33473/_0_ , \g33474/_0_ , \g33475/_0_ , \g33476/_0_ , \g33477/_0_ , \g33478/_0_ , \g33479/_0_ , \g33480/_0_ , \g33481/_0_ , \g33482/_0_ , \g33483/_0_ , \g33484/_0_ , \g33485/_0_ , \g33486/_0_ , \g33487/_0_ , \g33488/_0_ , \g33489/_0_ , \g33490/_0_ , \g33491/_0_ , \g33492/_0_ , \g33493/_0_ , \g33494/_0_ , \g33495/_0_ , \g33496/_0_ , \g33497/_0_ , \g33498/_0_ , \g33499/_0_ , \g33500/_0_ , \g33501/_0_ , \g33502/_0_ , \g33503/_0_ , \g33504/_0_ , \g33505/_0_ , \g33506/_0_ , \g33507/_0_ , \g33508/_0_ , \g33509/_0_ , \g33510/_0_ , \g33511/_0_ , \g33512/_0_ , \g33513/_0_ , \g33514/_0_ , \g33515/_0_ , \g33516/_0_ , \g33517/_0_ , \g33518/_0_ , \g33519/_0_ , \g33520/_0_ , \g33521/_0_ , \g33522/_0_ , \g33523/_0_ , \g33524/_0_ , \g33525/_0_ , \g33526/_0_ , \g33527/_0_ , \g33528/_0_ , \g33529/_0_ , \g33530/_0_ , \g33531/_0_ , \g33532/_0_ , \g33533/_0_ , \g33534/_0_ , \g33535/_0_ , \g33536/_0_ , \g33537/_0_ , \g33538/_0_ , \g33539/_0_ , \g33540/_0_ , \g33541/_0_ , \g33542/_0_ , \g33543/_0_ , \g33544/_0_ , \g33545/_0_ , \g33546/_0_ , \g33547/_0_ , \g33548/_0_ , \g33549/_0_ , \g33550/_0_ , \g33551/_0_ , \g33552/_0_ , \g33553/_0_ , \g33554/_0_ , \g33555/_0_ , \g33556/_0_ , \g33557/_0_ , \g33558/_0_ , \g33559/_0_ , \g33560/_0_ , \g33561/_0_ , \g33562/_0_ , \g33563/_0_ , \g33564/_0_ , \g33565/_0_ , \g33566/_0_ , \g33567/_0_ , \g33568/_0_ , \g33569/_0_ , \g33570/_0_ , \g33571/_0_ , \g33572/_0_ , \g33573/_0_ , \g33574/_0_ , \g33575/_0_ , \g33576/_0_ , \g33577/_0_ , \g33578/_0_ , \g33579/_0_ , \g33580/_0_ , \g33581/_0_ , \g33582/_0_ , \g33583/_0_ , \g33584/_0_ , \g33585/_0_ , \g33586/_0_ , \g33587/_0_ , \g33588/_0_ , \g33589/_0_ , \g33590/_0_ , \g33591/_0_ , \g33592/_0_ , \g33593/_0_ , \g33594/_0_ , \g33595/_0_ , \g33596/_0_ , \g33597/_0_ , \g33598/_0_ , \g33599/_0_ , \g33600/_0_ , \g33601/_0_ , \g33602/_0_ , \g33603/_0_ , \g33604/_0_ , \g33605/_0_ , \g33606/_0_ , \g33607/_0_ , \g33608/_0_ , \g33609/_0_ , \g33610/_0_ , \g33611/_0_ , \g33612/_0_ , \g33613/_0_ , \g33614/_0_ , \g33615/_0_ , \g33616/_0_ , \g33617/_0_ , \g33618/_0_ , \g33619/_0_ , \g33620/_0_ , \g33621/_0_ , \g33622/_0_ , \g33623/_0_ , \g33624/_0_ , \g33625/_0_ , \g33626/_0_ , \g33627/_0_ , \g33628/_0_ , \g33629/_0_ , \g33630/_0_ , \g33631/_0_ , \g33632/_0_ , \g33633/_0_ , \g33634/_0_ , \g33635/_0_ , \g33636/_0_ , \g33637/_0_ , \g33638/_0_ , \g33639/_0_ , \g33640/_0_ , \g33641/_0_ , \g33642/_0_ , \g33643/_0_ , \g33644/_0_ , \g33645/_0_ , \g33646/_0_ , \g33647/_0_ , \g33648/_0_ , \g33649/_0_ , \g33650/_0_ , \g33651/_0_ , \g33652/_0_ , \g33653/_0_ , \g33654/_0_ , \g33655/_0_ , \g33656/_0_ , \g33657/_0_ , \g33658/_0_ , \g33659/_0_ , \g33660/_0_ , \g33661/_0_ , \g33662/_0_ , \g33663/_0_ , \g33664/_0_ , \g33665/_0_ , \g33666/_0_ , \g33667/_0_ , \g33668/_0_ , \g33669/_0_ , \g33670/_0_ , \g33671/_0_ , \g33672/_0_ , \g33673/_0_ , \g33674/_0_ , \g33675/_0_ , \g33676/_0_ , \g33677/_0_ , \g33678/_0_ , \g33679/_0_ , \g33680/_0_ , \g33681/_0_ , \g33682/_0_ , \g33683/_0_ , \g33684/_0_ , \g33685/_0_ , \g33686/_0_ , \g33687/_0_ , \g33688/_0_ , \g33689/_0_ , \g33690/_0_ , \g33691/_0_ , \g33692/_0_ , \g33693/_0_ , \g33694/_0_ , \g33695/_0_ , \g33696/_0_ , \g33697/_0_ , \g33698/_0_ , \g33699/_0_ , \g33700/_0_ , \g33701/_0_ , \g33702/_0_ , \g33703/_0_ , \g33704/_0_ , \g33705/_0_ , \g33706/_0_ , \g33707/_0_ , \g33708/_0_ , \g33709/_0_ , \g33710/_0_ , \g33711/_0_ , \g33712/_0_ , \g33713/_0_ , \g33714/_0_ , \g33715/_0_ , \g33716/_0_ , \g33717/_0_ , \g33718/_0_ , \g33719/_0_ , \g33720/_0_ , \g33721/_0_ , \g33722/_0_ , \g33723/_0_ , \g33724/_0_ , \g33725/_0_ , \g33726/_0_ , \g33727/_0_ , \g33728/_0_ , \g33729/_0_ , \g33730/_0_ , \g33731/_0_ , \g33732/_0_ , \g33733/_0_ , \g33734/_0_ , \g33735/_0_ , \g33736/_0_ , \g33737/_0_ , \g33738/_0_ , \g33739/_0_ , \g33740/_0_ , \g33741/_0_ , \g33742/_0_ , \g33743/_0_ , \g33744/_0_ , \g33745/_0_ , \g33746/_0_ , \g33747/_0_ , \g33748/_0_ , \g33749/_0_ , \g33750/_0_ , \g33751/_0_ , \g33752/_0_ , \g33753/_0_ , \g33754/_0_ , \g33755/_0_ , \g33756/_0_ , \g33757/_0_ , \g33758/_0_ , \g33759/_0_ , \g33760/_0_ , \g33761/_0_ , \g33762/_0_ , \g33763/_0_ , \g33764/_0_ , \g33765/_0_ , \g33766/_0_ , \g33767/_0_ , \g33768/_0_ , \g33769/_0_ , \g33770/_0_ , \g33771/_0_ , \g33772/_0_ , \g33773/_0_ , \g33774/_0_ , \g33775/_0_ , \g33776/_0_ , \g33777/_0_ , \g33778/_0_ , \g33779/_0_ , \g33780/_0_ , \g33781/_0_ , \g33782/_0_ , \g33783/_0_ , \g33784/_0_ , \g33785/_0_ , \g33786/_0_ , \g33787/_0_ , \g33788/_0_ , \g33789/_0_ , \g33790/_0_ , \g33791/_0_ , \g33792/_0_ , \g33793/_0_ , \g33794/_0_ , \g33795/_0_ , \g33796/_0_ , \g33797/_0_ , \g33798/_0_ , \g33799/_0_ , \g33800/_0_ , \g33801/_0_ , \g33802/_0_ , \g33803/_0_ , \g33804/_0_ , \g33805/_0_ , \g33806/_0_ , \g33807/_0_ , \g33808/_0_ , \g33809/_0_ , \g33810/_0_ , \g33811/_0_ , \g33812/_0_ , \g33813/_0_ , \g33814/_0_ , \g33815/_0_ , \g33816/_0_ , \g33817/_0_ , \g33818/_0_ , \g33819/_0_ , \g33820/_0_ , \g33821/_0_ , \g33822/_0_ , \g33823/_0_ , \g33824/_0_ , \g33825/_0_ , \g33826/_0_ , \g33827/_0_ , \g33828/_0_ , \g33829/_0_ , \g33830/_0_ , \g33831/_0_ , \g33832/_0_ , \g33833/_0_ , \g33834/_0_ , \g33835/_0_ , \g33836/_0_ , \g33837/_0_ , \g33838/_0_ , \g33839/_0_ , \g33840/_0_ , \g33841/_0_ , \g33842/_0_ , \g33843/_0_ , \g33844/_0_ , \g33845/_0_ , \g33846/_0_ , \g33847/_0_ , \g33848/_0_ , \g33849/_0_ , \g33850/_0_ , \g33851/_0_ , \g33852/_0_ , \g33853/_0_ , \g33854/_0_ , \g33855/_0_ , \g33856/_0_ , \g33857/_0_ , \g33858/_0_ , \g33859/_0_ , \g33860/_0_ , \g33861/_0_ , \g33862/_0_ , \g33863/_0_ , \g33864/_0_ , \g33865/_0_ , \g33866/_0_ , \g33867/_0_ , \g33868/_0_ , \g33869/_0_ , \g33870/_0_ , \g33871/_0_ , \g33872/_0_ , \g33873/_0_ , \g33874/_0_ , \g33875/_0_ , \g33876/_0_ , \g33877/_0_ , \g33878/_0_ , \g33879/_0_ , \g33880/_0_ , \g33881/_0_ , \g33882/_0_ , \g33883/_0_ , \g33884/_0_ , \g33885/_0_ , \g33886/_0_ , \g33887/_0_ , \g33888/_0_ , \g33889/_0_ , \g33890/_0_ , \g33891/_0_ , \g33892/_0_ , \g33893/_0_ , \g33894/_0_ , \g33895/_0_ , \g33896/_0_ , \g33897/_0_ , \g33898/_0_ , \g33899/_0_ , \g33900/_0_ , \g33901/_0_ , \g33902/_0_ , \g33903/_0_ , \g33904/_0_ , \g33905/_0_ , \g33906/_0_ , \g33907/_0_ , \g33908/_0_ , \g33909/_0_ , \g33910/_0_ , \g33911/_0_ , \g33912/_0_ , \g33913/_0_ , \g33914/_0_ , \g33915/_0_ , \g33916/_0_ , \g33917/_0_ , \g33918/_0_ , \g33919/_0_ , \g33920/_0_ , \g33921/_0_ , \g33922/_0_ , \g33923/_0_ , \g33924/_0_ , \g33925/_0_ , \g33926/_0_ , \g33927/_0_ , \g33928/_0_ , \g33929/_0_ , \g33930/_0_ , \g33931/_0_ , \g33932/_0_ , \g33933/_0_ , \g33934/_0_ , \g33935/_0_ , \g33936/_0_ , \g33937/_0_ , \g33938/_0_ , \g33939/_0_ , \g33940/_0_ , \g33941/_0_ , \g33942/_0_ , \g33943/_0_ , \g33944/_0_ , \g33945/_0_ , \g33946/_0_ , \g33947/_0_ , \g33948/_0_ , \g33949/_0_ , \g33950/_0_ , \g33951/_0_ , \g33952/_0_ , \g33953/_0_ , \g33954/_0_ , \g33955/_0_ , \g33956/_0_ , \g33957/_0_ , \g33958/_0_ , \g33959/_0_ , \g33960/_0_ , \g33961/_0_ , \g33962/_0_ , \g33963/_0_ , \g33964/_0_ , \g33965/_0_ , \g33966/_0_ , \g33967/_0_ , \g33968/_0_ , \g33969/_0_ , \g33970/_0_ , \g33971/_0_ , \g33972/_0_ , \g33973/_0_ , \g33974/_0_ , \g33975/_0_ , \g33976/_0_ , \g33977/u3_syn_4 , \g33981/u3_syn_4 , \g34014/u3_syn_4 , \g34047/u3_syn_4 , \g34084/u3_syn_4 , \g34123/u3_syn_4 , \g34306/_0_ , \g34316/_0_ , \g34324/_0_ , \g34326/_0_ , \g34328/_0_ , \g34331/_0_ , \g34333/_0_ , \g34344/_0_ , \g34347/_0_ , \g34351/_0_ , \g34361/_0_ , \g34368/_0_ , \g34377/_0_ , \g34385/_0_ , \g34393/_0_ , \g34414/_1_ , \g34451/_1_ , \g34476/_1_ , \g34487/_0_ , \g34490/_1_ , \g34715/_0_ , \g34878/_0_ , \g34882/_0_ , \g34883/_0_ , \g34893/_0_ , \g34896/_0_ , \g34898/_0_ , \g34899/_0_ , \g34916/_3_ , \g35264/_0_ , \g35265/_0_ , \g35266/_0_ , \g35267/_0_ , \g35268/_0_ , \g35269/_0_ , \g35270/_0_ , \g35271/_0_ , \g35272/_0_ , \g35273/_0_ , \g35274/_0_ , \g35275/_0_ , \g35276/_0_ , \g35277/_0_ , \g35278/_0_ , \g35279/_0_ , \g35283/_0_ , \g35287/_0_ , \g35294/_0_ , \g35300/_0_ , \g35304/_0_ , \g35308/_0_ , \g35312/_0_ , \g35316/_0_ , \g35318/_0_ , \g35326/_0_ , \g35334/_0_ , \g35336/_0_ , \g35337/_0_ , \g35338/_0_ , \g35357/_0_ , \g35358/_0_ , \g35359/_0_ , \g35419/_0_ , \g35438/_0_ , \g35439/_0_ , \g35440/_0_ , \g35441/_0_ , \g35442/_0_ , \g35444/_0_ , \g35445/_0_ , \g35446/_0_ , \g35447/_0_ , \g35448/_0_ , \g35449/_0_ , \g35450/_0_ , \g35451/_0_ , \g35452/_0_ , \g35463/_0_ , \g35464/_0_ , \g35466/_0_ , \g35485/_2_ , \g35495/_0_ , \g35496/_0_ , \g35499/_0_ , \g35500/_0_ , \g35501/_0_ , \g35502/_0_ , \g35563/_0_ , \g35633/_0_ , \g35717/_0_ , \g35718/_0_ , \g35719/_0_ , \g35809/_0_ , \g35810/_0_ , \g35811/_0_ , \g35812/_0_ , \g35813/_0_ , \g35814/_0_ , \g35815/_0_ , \g35816/_0_ , \g35817/_0_ , \g35818/_0_ , \g35819/_0_ , \g35820/_0_ , \g35821/_0_ , \g35822/_0_ , \g35823/_0_ , \g35824/_0_ , \g35825/_0_ , \g35826/_0_ , \g35827/_0_ , \g35830/_0_ , \g35833/_0_ , \g35835/_0_ , \g35836/_0_ , \g35837/_0_ , \g35839/_0_ , \g35840/_0_ , \g35841/_0_ , \g35843/_0_ , \g35844/_0_ , \g35845/_0_ , \g35853/_0_ , \g35854/_0_ , \g35855/_0_ , \g35856/_0_ , \g36306/_0_ , \g36414/_0_ , \g36415/_0_ , \g36449/_0_ , \g36550/_0_ , \g36551/_0_ , \g36553/_0_ , \g36560/_0_ , \g36562/_3_ , \g36563/_0_ , \g36612/_0_ , \g36614/_2_ , \g36695/_0_ , \g36784/_0_ , \g36785/_0_ , \g36786/_0_ , \g36787/_0_ , \g36788/_0_ , \g36789/_0_ , \g36790/_0_ , \g36791/_0_ , \g36792/_0_ , \g36793/_0_ , \g36794/_0_ , \g36796/_0_ , \g36797/_0_ , \g36798/_0_ , \g36799/_0_ , \g36800/_0_ , \g36801/_0_ , \g36802/_0_ , \g36803/_0_ , \g36804/_0_ , \g36805/_0_ , \g36806/_0_ , \g36807/_0_ , \g36808/_0_ , \g36809/_0_ , \g36810/_0_ , \g36811/_0_ , \g36813/_0_ , \g36814/_0_ , \g36815/_0_ , \g36820/_0_ , \g36825/_0_ , \g36832/_0_ , \g36846/_0_ , \g36855/_0_ , \g36857/_0_ , \g36859/_0_ , \g36860/_0_ , \g36861/_0_ , \g36862/_0_ , \g36863/_0_ , \g36864/_0_ , \g36867/_0_ , \g36870/_0_ , \g36871/_0_ , \g36877/_0_ , \g36879/_0_ , \g36892/_0_ , \g36893/_0_ , \g36901/_0_ , \g36909/_0_ , \g36914/_0_ , \g36919/_0_ , \g36922/_0_ , \g36923/_0_ , \g36927/_0_ , \g36930/_0_ , \g36931/_0_ , \g36933/_0_ , \g36934/_0_ , \g36935/_0_ , \g36936/_0_ , \g36937/_0_ , \g36938/_0_ , \g36939/_0_ , \g36940/_0_ , \g36941/_0_ , \g36943/_0_ , \g36944/_0_ , \g36945/_0_ , \g36946/_0_ , \g36947/_0_ , \g36948/_0_ , \g36949/_0_ , \g36950/_0_ , \g36951/_0_ , \g36952/_0_ , \g36953/_0_ , \g36954/_0_ , \g36957/_0_ , \g36958/_0_ , \g36959/_0_ , \g36960/_0_ , \g36961/_0_ , \g36962/_0_ , \g36963/_0_ , \g36970/_0_ , \g36977/_0_ , \g36986/_0_ , \g36991/_0_ , \g36994/_0_ , \g37015/_0_ , \g37057/_0_ , \g37073/_0_ , \g37128/_0_ , \g37129/_0_ , \g37138/_0_ , \g37139/_0_ , \g37140/_0_ , \g37141/_0_ , \g37142/_0_ , \g37143/_0_ , \g37144/_0_ , \g37145/_0_ , \g37146/_0_ , \g37147/_0_ , \g37148/_0_ , \g37149/_0_ , \g37150/_0_ , \g37151/_0_ , \g37152/_0_ , \g37153/_0_ , \g37154/_0_ , \g37155/_0_ , \g37156/_0_ , \g37157/_0_ , \g37158/_0_ , \g37159/_0_ , \g37160/_0_ , \g37161/_0_ , \g37162/_0_ , \g37163/_0_ , \g37164/_0_ , \g37165/_0_ , \g37166/_0_ , \g37167/_0_ , \g37168/_0_ , \g37169/_0_ , \g37170/_0_ , \g37171/_0_ , \g37172/_0_ , \g37173/_0_ , \g37174/_0_ , \g37175/_0_ , \g37176/_0_ , \g37177/_0_ , \g37178/_0_ , \g37179/_0_ , \g37180/_0_ , \g37181/_0_ , \g37182/_0_ , \g37183/_0_ , \g37184/_0_ , \g37185/_0_ , \g37187/_0_ , \g37188/_0_ , \g37190/_0_ , \g37191/_0_ , \g37192/_0_ , \g37193/_0_ , \g37194/_0_ , \g37372/_3_ , \g37377/_0_ , \g37378/_0_ , \g37379/_0_ , \g37380/_0_ , \g37381/_0_ , \g37382/_0_ , \g37383/_0_ , \g37384/_0_ , \g37385/_0_ , \g37386/_0_ , \g37387/_0_ , \g37388/_0_ , \g37389/_0_ , \g37390/_0_ , \g37391/_0_ , \g37392/_0_ , \g37393/_0_ , \g37394/_0_ , \g37395/_0_ , \g37396/_0_ , \g37397/_0_ , \g37398/_0_ , \g37399/_0_ , \g37400/_0_ , \g37401/_0_ , \g37402/_0_ , \g37403/_0_ , \g37404/_0_ , \g37405/_0_ , \g37406/_0_ , \g37407/_0_ , \g37408/_0_ , \g37409/_0_ , \g37410/_0_ , \g37411/_0_ , \g37412/_0_ , \g37413/_0_ , \g37576/_3_ , \g37590/_2_ , \g40278/_0_ , \g40379/_0_ , \g40389/_2_ , \g40390/_2_ , \g40391/_0_ , \g40393/_2_ , \g40395/_0_ , \g40397/_0_ , \g40400/_0_ , \g40402/_0_ , \g45458/_0_ , \g45675/_0_ , \g45677/_0_ , \g45678/_0_ , \g45682/_0_ , sync_pad_o_pad, \u14_u0_full_empty_r_reg/P0001_reg_syn_3 , \u14_u1_full_empty_r_reg/P0001_reg_syn_3 , \u14_u2_full_empty_r_reg/P0001_reg_syn_3 , \u14_u3_full_empty_r_reg/P0001_reg_syn_3 , \u14_u4_full_empty_r_reg/P0001_reg_syn_3 , \u14_u5_full_empty_r_reg/P0001_reg_syn_3 , \u14_u6_full_empty_r_reg/P0001_reg_syn_3 , \u14_u7_full_empty_r_reg/P0001_reg_syn_3 , \u14_u8_full_empty_r_reg/P0001_reg_syn_3 , \u1_slt0_reg[11]/P0001_reg_syn_3 , \u1_slt0_reg[12]/P0001_reg_syn_3 , \u1_slt0_reg[15]/P0001_reg_syn_3 , \u1_slt0_reg[9]/P0001_reg_syn_3 , \u1_slt1_reg[10]/P0001_reg_syn_3 , \u1_slt1_reg[11]/P0001_reg_syn_3 , \u1_slt1_reg[5]/P0001_reg_syn_3 , \u1_slt1_reg[6]/P0001_reg_syn_3 , \u1_slt1_reg[7]/P0001_reg_syn_3 , \u1_slt1_reg[8]/P0001_reg_syn_3 , wb_err_o_pad);
	input \ac97_reset_pad_o__pad  ;
	input \dma_ack_i[0]_pad  ;
	input \dma_ack_i[1]_pad  ;
	input \dma_ack_i[2]_pad  ;
	input \dma_ack_i[3]_pad  ;
	input \dma_ack_i[4]_pad  ;
	input \dma_ack_i[5]_pad  ;
	input \dma_ack_i[6]_pad  ;
	input \dma_ack_i[7]_pad  ;
	input \dma_ack_i[8]_pad  ;
	input \dma_req_o[0]_pad  ;
	input \dma_req_o[1]_pad  ;
	input \dma_req_o[2]_pad  ;
	input \dma_req_o[3]_pad  ;
	input \dma_req_o[4]_pad  ;
	input \dma_req_o[5]_pad  ;
	input \dma_req_o[6]_pad  ;
	input \dma_req_o[7]_pad  ;
	input \dma_req_o[8]_pad  ;
	input \in_valid_s_reg[0]/NET0131  ;
	input \in_valid_s_reg[1]/NET0131  ;
	input \in_valid_s_reg[2]/NET0131  ;
	input suspended_o_pad ;
	input \u0_slt0_r_reg[0]/P0001  ;
	input \u0_slt0_r_reg[10]/P0001  ;
	input \u0_slt0_r_reg[11]/P0001  ;
	input \u0_slt0_r_reg[12]/P0001  ;
	input \u0_slt0_r_reg[13]/P0001  ;
	input \u0_slt0_r_reg[14]/P0001  ;
	input \u0_slt0_r_reg[1]/P0001  ;
	input \u0_slt0_r_reg[2]/P0001  ;
	input \u0_slt0_r_reg[3]/P0001  ;
	input \u0_slt0_r_reg[4]/P0001  ;
	input \u0_slt0_r_reg[5]/P0001  ;
	input \u0_slt0_r_reg[6]/P0001  ;
	input \u0_slt0_r_reg[7]/P0001  ;
	input \u0_slt0_r_reg[8]/P0001  ;
	input \u0_slt0_r_reg[9]/P0001  ;
	input \u0_slt1_r_reg[0]/P0001  ;
	input \u0_slt1_r_reg[10]/P0001  ;
	input \u0_slt1_r_reg[11]/P0001  ;
	input \u0_slt1_r_reg[12]/P0001  ;
	input \u0_slt1_r_reg[13]/P0001  ;
	input \u0_slt1_r_reg[14]/P0001  ;
	input \u0_slt1_r_reg[15]/P0001  ;
	input \u0_slt1_r_reg[16]/P0001  ;
	input \u0_slt1_r_reg[17]/P0001  ;
	input \u0_slt1_r_reg[18]/P0001  ;
	input \u0_slt1_r_reg[19]/P0001  ;
	input \u0_slt1_r_reg[1]/P0001  ;
	input \u0_slt1_r_reg[2]/P0001  ;
	input \u0_slt1_r_reg[3]/P0001  ;
	input \u0_slt1_r_reg[4]/P0001  ;
	input \u0_slt1_r_reg[5]/P0001  ;
	input \u0_slt1_r_reg[6]/P0001  ;
	input \u0_slt1_r_reg[7]/P0001  ;
	input \u0_slt1_r_reg[8]/P0001  ;
	input \u0_slt1_r_reg[9]/P0001  ;
	input \u0_slt2_r_reg[0]/P0001  ;
	input \u0_slt2_r_reg[10]/P0001  ;
	input \u0_slt2_r_reg[11]/P0001  ;
	input \u0_slt2_r_reg[12]/P0001  ;
	input \u0_slt2_r_reg[13]/P0001  ;
	input \u0_slt2_r_reg[14]/P0001  ;
	input \u0_slt2_r_reg[15]/P0001  ;
	input \u0_slt2_r_reg[16]/P0001  ;
	input \u0_slt2_r_reg[17]/P0001  ;
	input \u0_slt2_r_reg[18]/P0001  ;
	input \u0_slt2_r_reg[19]/P0001  ;
	input \u0_slt2_r_reg[1]/P0001  ;
	input \u0_slt2_r_reg[2]/P0001  ;
	input \u0_slt2_r_reg[3]/P0001  ;
	input \u0_slt2_r_reg[4]/P0001  ;
	input \u0_slt2_r_reg[5]/P0001  ;
	input \u0_slt2_r_reg[6]/P0001  ;
	input \u0_slt2_r_reg[7]/P0001  ;
	input \u0_slt2_r_reg[8]/P0001  ;
	input \u0_slt2_r_reg[9]/P0001  ;
	input \u0_slt3_r_reg[0]/P0001  ;
	input \u0_slt3_r_reg[10]/P0001  ;
	input \u0_slt3_r_reg[11]/P0001  ;
	input \u0_slt3_r_reg[12]/P0001  ;
	input \u0_slt3_r_reg[13]/P0001  ;
	input \u0_slt3_r_reg[14]/P0001  ;
	input \u0_slt3_r_reg[15]/P0001  ;
	input \u0_slt3_r_reg[16]/P0001  ;
	input \u0_slt3_r_reg[17]/P0001  ;
	input \u0_slt3_r_reg[18]/P0001  ;
	input \u0_slt3_r_reg[19]/P0001  ;
	input \u0_slt3_r_reg[1]/P0001  ;
	input \u0_slt3_r_reg[2]/P0001  ;
	input \u0_slt3_r_reg[3]/P0001  ;
	input \u0_slt3_r_reg[4]/P0001  ;
	input \u0_slt3_r_reg[5]/P0001  ;
	input \u0_slt3_r_reg[6]/P0001  ;
	input \u0_slt3_r_reg[7]/P0001  ;
	input \u0_slt3_r_reg[8]/P0001  ;
	input \u0_slt3_r_reg[9]/P0001  ;
	input \u0_slt4_r_reg[0]/P0001  ;
	input \u0_slt4_r_reg[10]/P0001  ;
	input \u0_slt4_r_reg[11]/P0001  ;
	input \u0_slt4_r_reg[12]/P0001  ;
	input \u0_slt4_r_reg[13]/P0001  ;
	input \u0_slt4_r_reg[14]/P0001  ;
	input \u0_slt4_r_reg[15]/P0001  ;
	input \u0_slt4_r_reg[16]/P0001  ;
	input \u0_slt4_r_reg[17]/P0001  ;
	input \u0_slt4_r_reg[18]/P0001  ;
	input \u0_slt4_r_reg[19]/P0001  ;
	input \u0_slt4_r_reg[1]/P0001  ;
	input \u0_slt4_r_reg[2]/P0001  ;
	input \u0_slt4_r_reg[3]/P0001  ;
	input \u0_slt4_r_reg[4]/P0001  ;
	input \u0_slt4_r_reg[5]/P0001  ;
	input \u0_slt4_r_reg[6]/P0001  ;
	input \u0_slt4_r_reg[7]/P0001  ;
	input \u0_slt4_r_reg[8]/P0001  ;
	input \u0_slt4_r_reg[9]/P0001  ;
	input \u0_slt5_r_reg[0]/P0001  ;
	input \u0_slt5_r_reg[10]/P0001  ;
	input \u0_slt5_r_reg[11]/P0001  ;
	input \u0_slt5_r_reg[12]/P0001  ;
	input \u0_slt5_r_reg[13]/P0001  ;
	input \u0_slt5_r_reg[14]/P0001  ;
	input \u0_slt5_r_reg[15]/P0001  ;
	input \u0_slt5_r_reg[16]/P0001  ;
	input \u0_slt5_r_reg[17]/P0001  ;
	input \u0_slt5_r_reg[18]/P0001  ;
	input \u0_slt5_r_reg[19]/P0001  ;
	input \u0_slt5_r_reg[1]/P0001  ;
	input \u0_slt5_r_reg[2]/P0001  ;
	input \u0_slt5_r_reg[3]/P0001  ;
	input \u0_slt5_r_reg[4]/P0001  ;
	input \u0_slt5_r_reg[5]/P0001  ;
	input \u0_slt5_r_reg[6]/P0001  ;
	input \u0_slt5_r_reg[7]/P0001  ;
	input \u0_slt5_r_reg[8]/P0001  ;
	input \u0_slt5_r_reg[9]/P0001  ;
	input \u0_slt6_r_reg[0]/P0001  ;
	input \u0_slt6_r_reg[10]/P0001  ;
	input \u0_slt6_r_reg[11]/P0001  ;
	input \u0_slt6_r_reg[12]/P0001  ;
	input \u0_slt6_r_reg[13]/P0001  ;
	input \u0_slt6_r_reg[14]/P0001  ;
	input \u0_slt6_r_reg[15]/P0001  ;
	input \u0_slt6_r_reg[16]/P0001  ;
	input \u0_slt6_r_reg[17]/P0001  ;
	input \u0_slt6_r_reg[18]/P0001  ;
	input \u0_slt6_r_reg[19]/P0001  ;
	input \u0_slt6_r_reg[1]/P0001  ;
	input \u0_slt6_r_reg[2]/P0001  ;
	input \u0_slt6_r_reg[3]/P0001  ;
	input \u0_slt6_r_reg[4]/P0001  ;
	input \u0_slt6_r_reg[5]/P0001  ;
	input \u0_slt6_r_reg[6]/P0001  ;
	input \u0_slt6_r_reg[7]/P0001  ;
	input \u0_slt6_r_reg[8]/P0001  ;
	input \u0_slt6_r_reg[9]/P0001  ;
	input \u0_slt7_r_reg[0]/P0001  ;
	input \u0_slt7_r_reg[10]/P0001  ;
	input \u0_slt7_r_reg[11]/P0001  ;
	input \u0_slt7_r_reg[12]/P0001  ;
	input \u0_slt7_r_reg[13]/P0001  ;
	input \u0_slt7_r_reg[14]/P0001  ;
	input \u0_slt7_r_reg[15]/P0001  ;
	input \u0_slt7_r_reg[16]/P0001  ;
	input \u0_slt7_r_reg[17]/P0001  ;
	input \u0_slt7_r_reg[18]/P0001  ;
	input \u0_slt7_r_reg[19]/P0001  ;
	input \u0_slt7_r_reg[1]/P0001  ;
	input \u0_slt7_r_reg[2]/P0001  ;
	input \u0_slt7_r_reg[3]/P0001  ;
	input \u0_slt7_r_reg[4]/P0001  ;
	input \u0_slt7_r_reg[5]/P0001  ;
	input \u0_slt7_r_reg[6]/P0001  ;
	input \u0_slt7_r_reg[7]/P0001  ;
	input \u0_slt7_r_reg[8]/P0001  ;
	input \u0_slt7_r_reg[9]/P0001  ;
	input \u0_slt8_r_reg[0]/P0001  ;
	input \u0_slt8_r_reg[10]/P0001  ;
	input \u0_slt8_r_reg[11]/P0001  ;
	input \u0_slt8_r_reg[12]/P0001  ;
	input \u0_slt8_r_reg[13]/P0001  ;
	input \u0_slt8_r_reg[14]/P0001  ;
	input \u0_slt8_r_reg[15]/P0001  ;
	input \u0_slt8_r_reg[16]/P0001  ;
	input \u0_slt8_r_reg[17]/P0001  ;
	input \u0_slt8_r_reg[18]/P0001  ;
	input \u0_slt8_r_reg[19]/P0001  ;
	input \u0_slt8_r_reg[1]/P0001  ;
	input \u0_slt8_r_reg[2]/P0001  ;
	input \u0_slt8_r_reg[3]/P0001  ;
	input \u0_slt8_r_reg[4]/P0001  ;
	input \u0_slt8_r_reg[5]/P0001  ;
	input \u0_slt8_r_reg[6]/P0001  ;
	input \u0_slt8_r_reg[7]/P0001  ;
	input \u0_slt8_r_reg[8]/P0001  ;
	input \u0_slt8_r_reg[9]/P0001  ;
	input \u0_slt9_r_reg[0]/P0001  ;
	input \u0_slt9_r_reg[10]/P0001  ;
	input \u0_slt9_r_reg[11]/P0001  ;
	input \u0_slt9_r_reg[12]/P0001  ;
	input \u0_slt9_r_reg[13]/P0001  ;
	input \u0_slt9_r_reg[14]/P0001  ;
	input \u0_slt9_r_reg[15]/P0001  ;
	input \u0_slt9_r_reg[16]/P0001  ;
	input \u0_slt9_r_reg[17]/P0001  ;
	input \u0_slt9_r_reg[18]/P0001  ;
	input \u0_slt9_r_reg[19]/P0001  ;
	input \u0_slt9_r_reg[1]/P0001  ;
	input \u0_slt9_r_reg[2]/P0001  ;
	input \u0_slt9_r_reg[3]/P0001  ;
	input \u0_slt9_r_reg[4]/P0001  ;
	input \u0_slt9_r_reg[5]/P0001  ;
	input \u0_slt9_r_reg[6]/P0001  ;
	input \u0_slt9_r_reg[7]/P0001  ;
	input \u0_slt9_r_reg[8]/P0001  ;
	input \u0_slt9_r_reg[9]/P0001  ;
	input \u10_din_tmp1_reg[0]/P0001  ;
	input \u10_din_tmp1_reg[10]/P0001  ;
	input \u10_din_tmp1_reg[11]/P0001  ;
	input \u10_din_tmp1_reg[12]/P0001  ;
	input \u10_din_tmp1_reg[13]/P0001  ;
	input \u10_din_tmp1_reg[14]/P0001  ;
	input \u10_din_tmp1_reg[15]/P0001  ;
	input \u10_din_tmp1_reg[1]/P0001  ;
	input \u10_din_tmp1_reg[2]/P0001  ;
	input \u10_din_tmp1_reg[3]/P0001  ;
	input \u10_din_tmp1_reg[4]/P0001  ;
	input \u10_din_tmp1_reg[5]/P0001  ;
	input \u10_din_tmp1_reg[6]/P0001  ;
	input \u10_din_tmp1_reg[7]/P0001  ;
	input \u10_din_tmp1_reg[8]/P0001  ;
	input \u10_din_tmp1_reg[9]/P0001  ;
	input \u10_dout_reg[0]/P0001  ;
	input \u10_dout_reg[10]/P0001  ;
	input \u10_dout_reg[11]/P0001  ;
	input \u10_dout_reg[12]/P0001  ;
	input \u10_dout_reg[13]/P0001  ;
	input \u10_dout_reg[14]/P0001  ;
	input \u10_dout_reg[15]/P0001  ;
	input \u10_dout_reg[16]/P0001  ;
	input \u10_dout_reg[17]/P0001  ;
	input \u10_dout_reg[18]/P0001  ;
	input \u10_dout_reg[19]/P0001  ;
	input \u10_dout_reg[1]/P0001  ;
	input \u10_dout_reg[20]/P0001  ;
	input \u10_dout_reg[21]/P0001  ;
	input \u10_dout_reg[22]/P0001  ;
	input \u10_dout_reg[23]/P0001  ;
	input \u10_dout_reg[24]/P0001  ;
	input \u10_dout_reg[25]/P0001  ;
	input \u10_dout_reg[26]/P0001  ;
	input \u10_dout_reg[27]/P0001  ;
	input \u10_dout_reg[28]/P0001  ;
	input \u10_dout_reg[29]/P0001  ;
	input \u10_dout_reg[2]/P0001  ;
	input \u10_dout_reg[30]/P0001  ;
	input \u10_dout_reg[31]/P0001  ;
	input \u10_dout_reg[3]/P0001  ;
	input \u10_dout_reg[4]/P0001  ;
	input \u10_dout_reg[5]/P0001  ;
	input \u10_dout_reg[6]/P0001  ;
	input \u10_dout_reg[7]/P0001  ;
	input \u10_dout_reg[8]/P0001  ;
	input \u10_dout_reg[9]/P0001  ;
	input \u10_empty_reg/P0001  ;
	input \u10_full_reg/NET0131  ;
	input \u10_mem_reg[0][0]/P0001  ;
	input \u10_mem_reg[0][10]/P0001  ;
	input \u10_mem_reg[0][11]/P0001  ;
	input \u10_mem_reg[0][12]/P0001  ;
	input \u10_mem_reg[0][13]/P0001  ;
	input \u10_mem_reg[0][14]/P0001  ;
	input \u10_mem_reg[0][15]/P0001  ;
	input \u10_mem_reg[0][16]/P0001  ;
	input \u10_mem_reg[0][17]/P0001  ;
	input \u10_mem_reg[0][18]/P0001  ;
	input \u10_mem_reg[0][19]/P0001  ;
	input \u10_mem_reg[0][1]/P0001  ;
	input \u10_mem_reg[0][20]/P0001  ;
	input \u10_mem_reg[0][21]/P0001  ;
	input \u10_mem_reg[0][22]/P0001  ;
	input \u10_mem_reg[0][23]/P0001  ;
	input \u10_mem_reg[0][24]/P0001  ;
	input \u10_mem_reg[0][25]/P0001  ;
	input \u10_mem_reg[0][26]/P0001  ;
	input \u10_mem_reg[0][27]/P0001  ;
	input \u10_mem_reg[0][28]/P0001  ;
	input \u10_mem_reg[0][29]/P0001  ;
	input \u10_mem_reg[0][2]/P0001  ;
	input \u10_mem_reg[0][30]/P0001  ;
	input \u10_mem_reg[0][31]/P0001  ;
	input \u10_mem_reg[0][3]/P0001  ;
	input \u10_mem_reg[0][4]/P0001  ;
	input \u10_mem_reg[0][5]/P0001  ;
	input \u10_mem_reg[0][6]/P0001  ;
	input \u10_mem_reg[0][7]/P0001  ;
	input \u10_mem_reg[0][8]/P0001  ;
	input \u10_mem_reg[0][9]/P0001  ;
	input \u10_mem_reg[1][0]/P0001  ;
	input \u10_mem_reg[1][10]/P0001  ;
	input \u10_mem_reg[1][11]/P0001  ;
	input \u10_mem_reg[1][12]/P0001  ;
	input \u10_mem_reg[1][13]/P0001  ;
	input \u10_mem_reg[1][14]/P0001  ;
	input \u10_mem_reg[1][15]/P0001  ;
	input \u10_mem_reg[1][16]/P0001  ;
	input \u10_mem_reg[1][17]/P0001  ;
	input \u10_mem_reg[1][18]/P0001  ;
	input \u10_mem_reg[1][19]/P0001  ;
	input \u10_mem_reg[1][1]/P0001  ;
	input \u10_mem_reg[1][20]/P0001  ;
	input \u10_mem_reg[1][21]/P0001  ;
	input \u10_mem_reg[1][22]/P0001  ;
	input \u10_mem_reg[1][23]/P0001  ;
	input \u10_mem_reg[1][24]/P0001  ;
	input \u10_mem_reg[1][25]/P0001  ;
	input \u10_mem_reg[1][26]/P0001  ;
	input \u10_mem_reg[1][27]/P0001  ;
	input \u10_mem_reg[1][28]/P0001  ;
	input \u10_mem_reg[1][29]/P0001  ;
	input \u10_mem_reg[1][2]/P0001  ;
	input \u10_mem_reg[1][30]/P0001  ;
	input \u10_mem_reg[1][31]/P0001  ;
	input \u10_mem_reg[1][3]/P0001  ;
	input \u10_mem_reg[1][4]/P0001  ;
	input \u10_mem_reg[1][5]/P0001  ;
	input \u10_mem_reg[1][6]/P0001  ;
	input \u10_mem_reg[1][7]/P0001  ;
	input \u10_mem_reg[1][8]/P0001  ;
	input \u10_mem_reg[1][9]/P0001  ;
	input \u10_mem_reg[2][0]/P0001  ;
	input \u10_mem_reg[2][10]/P0001  ;
	input \u10_mem_reg[2][11]/P0001  ;
	input \u10_mem_reg[2][12]/P0001  ;
	input \u10_mem_reg[2][13]/P0001  ;
	input \u10_mem_reg[2][14]/P0001  ;
	input \u10_mem_reg[2][15]/P0001  ;
	input \u10_mem_reg[2][16]/P0001  ;
	input \u10_mem_reg[2][17]/P0001  ;
	input \u10_mem_reg[2][18]/P0001  ;
	input \u10_mem_reg[2][19]/P0001  ;
	input \u10_mem_reg[2][1]/P0001  ;
	input \u10_mem_reg[2][20]/P0001  ;
	input \u10_mem_reg[2][21]/P0001  ;
	input \u10_mem_reg[2][22]/P0001  ;
	input \u10_mem_reg[2][23]/P0001  ;
	input \u10_mem_reg[2][24]/P0001  ;
	input \u10_mem_reg[2][25]/P0001  ;
	input \u10_mem_reg[2][26]/P0001  ;
	input \u10_mem_reg[2][27]/P0001  ;
	input \u10_mem_reg[2][28]/P0001  ;
	input \u10_mem_reg[2][29]/P0001  ;
	input \u10_mem_reg[2][2]/P0001  ;
	input \u10_mem_reg[2][30]/P0001  ;
	input \u10_mem_reg[2][31]/P0001  ;
	input \u10_mem_reg[2][3]/P0001  ;
	input \u10_mem_reg[2][4]/P0001  ;
	input \u10_mem_reg[2][5]/P0001  ;
	input \u10_mem_reg[2][6]/P0001  ;
	input \u10_mem_reg[2][7]/P0001  ;
	input \u10_mem_reg[2][8]/P0001  ;
	input \u10_mem_reg[2][9]/P0001  ;
	input \u10_mem_reg[3][0]/P0001  ;
	input \u10_mem_reg[3][10]/P0001  ;
	input \u10_mem_reg[3][11]/P0001  ;
	input \u10_mem_reg[3][12]/P0001  ;
	input \u10_mem_reg[3][13]/P0001  ;
	input \u10_mem_reg[3][14]/P0001  ;
	input \u10_mem_reg[3][15]/P0001  ;
	input \u10_mem_reg[3][16]/P0001  ;
	input \u10_mem_reg[3][17]/P0001  ;
	input \u10_mem_reg[3][18]/P0001  ;
	input \u10_mem_reg[3][19]/P0001  ;
	input \u10_mem_reg[3][1]/P0001  ;
	input \u10_mem_reg[3][20]/P0001  ;
	input \u10_mem_reg[3][21]/P0001  ;
	input \u10_mem_reg[3][22]/P0001  ;
	input \u10_mem_reg[3][23]/P0001  ;
	input \u10_mem_reg[3][24]/P0001  ;
	input \u10_mem_reg[3][25]/P0001  ;
	input \u10_mem_reg[3][26]/P0001  ;
	input \u10_mem_reg[3][27]/P0001  ;
	input \u10_mem_reg[3][28]/P0001  ;
	input \u10_mem_reg[3][29]/P0001  ;
	input \u10_mem_reg[3][2]/P0001  ;
	input \u10_mem_reg[3][30]/P0001  ;
	input \u10_mem_reg[3][31]/P0001  ;
	input \u10_mem_reg[3][3]/P0001  ;
	input \u10_mem_reg[3][4]/P0001  ;
	input \u10_mem_reg[3][5]/P0001  ;
	input \u10_mem_reg[3][6]/P0001  ;
	input \u10_mem_reg[3][7]/P0001  ;
	input \u10_mem_reg[3][8]/P0001  ;
	input \u10_mem_reg[3][9]/P0001  ;
	input \u10_rp_reg[0]/P0001  ;
	input \u10_rp_reg[1]/P0001  ;
	input \u10_rp_reg[2]/P0001  ;
	input \u10_status_reg[0]/P0001  ;
	input \u10_status_reg[1]/P0001  ;
	input \u10_wp_reg[0]/NET0131  ;
	input \u10_wp_reg[1]/P0001  ;
	input \u10_wp_reg[2]/P0001  ;
	input \u10_wp_reg[3]/P0001  ;
	input \u11_din_tmp1_reg[0]/P0001  ;
	input \u11_din_tmp1_reg[10]/P0001  ;
	input \u11_din_tmp1_reg[11]/P0001  ;
	input \u11_din_tmp1_reg[12]/P0001  ;
	input \u11_din_tmp1_reg[13]/P0001  ;
	input \u11_din_tmp1_reg[14]/P0001  ;
	input \u11_din_tmp1_reg[15]/P0001  ;
	input \u11_din_tmp1_reg[1]/P0001  ;
	input \u11_din_tmp1_reg[2]/P0001  ;
	input \u11_din_tmp1_reg[3]/P0001  ;
	input \u11_din_tmp1_reg[4]/P0001  ;
	input \u11_din_tmp1_reg[5]/P0001  ;
	input \u11_din_tmp1_reg[6]/P0001  ;
	input \u11_din_tmp1_reg[7]/P0001  ;
	input \u11_din_tmp1_reg[8]/P0001  ;
	input \u11_din_tmp1_reg[9]/P0001  ;
	input \u11_dout_reg[0]/P0001  ;
	input \u11_dout_reg[10]/P0001  ;
	input \u11_dout_reg[11]/P0001  ;
	input \u11_dout_reg[12]/P0001  ;
	input \u11_dout_reg[13]/P0001  ;
	input \u11_dout_reg[14]/P0001  ;
	input \u11_dout_reg[15]/P0001  ;
	input \u11_dout_reg[16]/P0001  ;
	input \u11_dout_reg[17]/P0001  ;
	input \u11_dout_reg[18]/P0001  ;
	input \u11_dout_reg[19]/P0001  ;
	input \u11_dout_reg[1]/P0001  ;
	input \u11_dout_reg[20]/P0001  ;
	input \u11_dout_reg[21]/P0001  ;
	input \u11_dout_reg[22]/P0001  ;
	input \u11_dout_reg[23]/P0001  ;
	input \u11_dout_reg[24]/P0001  ;
	input \u11_dout_reg[25]/P0001  ;
	input \u11_dout_reg[26]/P0001  ;
	input \u11_dout_reg[27]/P0001  ;
	input \u11_dout_reg[28]/P0001  ;
	input \u11_dout_reg[29]/P0001  ;
	input \u11_dout_reg[2]/P0001  ;
	input \u11_dout_reg[30]/P0001  ;
	input \u11_dout_reg[31]/P0001  ;
	input \u11_dout_reg[3]/P0001  ;
	input \u11_dout_reg[4]/P0001  ;
	input \u11_dout_reg[5]/P0001  ;
	input \u11_dout_reg[6]/P0001  ;
	input \u11_dout_reg[7]/P0001  ;
	input \u11_dout_reg[8]/P0001  ;
	input \u11_dout_reg[9]/P0001  ;
	input \u11_empty_reg/P0001  ;
	input \u11_full_reg/NET0131  ;
	input \u11_mem_reg[0][0]/P0001  ;
	input \u11_mem_reg[0][10]/P0001  ;
	input \u11_mem_reg[0][11]/P0001  ;
	input \u11_mem_reg[0][12]/P0001  ;
	input \u11_mem_reg[0][13]/P0001  ;
	input \u11_mem_reg[0][14]/P0001  ;
	input \u11_mem_reg[0][15]/P0001  ;
	input \u11_mem_reg[0][16]/P0001  ;
	input \u11_mem_reg[0][17]/P0001  ;
	input \u11_mem_reg[0][18]/P0001  ;
	input \u11_mem_reg[0][19]/P0001  ;
	input \u11_mem_reg[0][1]/P0001  ;
	input \u11_mem_reg[0][20]/P0001  ;
	input \u11_mem_reg[0][21]/P0001  ;
	input \u11_mem_reg[0][22]/P0001  ;
	input \u11_mem_reg[0][23]/P0001  ;
	input \u11_mem_reg[0][24]/P0001  ;
	input \u11_mem_reg[0][25]/P0001  ;
	input \u11_mem_reg[0][26]/P0001  ;
	input \u11_mem_reg[0][27]/P0001  ;
	input \u11_mem_reg[0][28]/P0001  ;
	input \u11_mem_reg[0][29]/P0001  ;
	input \u11_mem_reg[0][2]/P0001  ;
	input \u11_mem_reg[0][30]/P0001  ;
	input \u11_mem_reg[0][31]/P0001  ;
	input \u11_mem_reg[0][3]/P0001  ;
	input \u11_mem_reg[0][4]/P0001  ;
	input \u11_mem_reg[0][5]/P0001  ;
	input \u11_mem_reg[0][6]/P0001  ;
	input \u11_mem_reg[0][7]/P0001  ;
	input \u11_mem_reg[0][8]/P0001  ;
	input \u11_mem_reg[0][9]/P0001  ;
	input \u11_mem_reg[1][0]/P0001  ;
	input \u11_mem_reg[1][10]/P0001  ;
	input \u11_mem_reg[1][11]/P0001  ;
	input \u11_mem_reg[1][12]/P0001  ;
	input \u11_mem_reg[1][13]/P0001  ;
	input \u11_mem_reg[1][14]/P0001  ;
	input \u11_mem_reg[1][15]/P0001  ;
	input \u11_mem_reg[1][16]/P0001  ;
	input \u11_mem_reg[1][17]/P0001  ;
	input \u11_mem_reg[1][18]/P0001  ;
	input \u11_mem_reg[1][19]/P0001  ;
	input \u11_mem_reg[1][1]/P0001  ;
	input \u11_mem_reg[1][20]/P0001  ;
	input \u11_mem_reg[1][21]/P0001  ;
	input \u11_mem_reg[1][22]/P0001  ;
	input \u11_mem_reg[1][23]/P0001  ;
	input \u11_mem_reg[1][24]/P0001  ;
	input \u11_mem_reg[1][25]/P0001  ;
	input \u11_mem_reg[1][26]/P0001  ;
	input \u11_mem_reg[1][27]/P0001  ;
	input \u11_mem_reg[1][28]/P0001  ;
	input \u11_mem_reg[1][29]/P0001  ;
	input \u11_mem_reg[1][2]/P0001  ;
	input \u11_mem_reg[1][30]/P0001  ;
	input \u11_mem_reg[1][31]/P0001  ;
	input \u11_mem_reg[1][3]/P0001  ;
	input \u11_mem_reg[1][4]/P0001  ;
	input \u11_mem_reg[1][5]/P0001  ;
	input \u11_mem_reg[1][6]/P0001  ;
	input \u11_mem_reg[1][7]/P0001  ;
	input \u11_mem_reg[1][8]/P0001  ;
	input \u11_mem_reg[1][9]/P0001  ;
	input \u11_mem_reg[2][0]/P0001  ;
	input \u11_mem_reg[2][10]/P0001  ;
	input \u11_mem_reg[2][11]/P0001  ;
	input \u11_mem_reg[2][12]/P0001  ;
	input \u11_mem_reg[2][13]/P0001  ;
	input \u11_mem_reg[2][14]/P0001  ;
	input \u11_mem_reg[2][15]/P0001  ;
	input \u11_mem_reg[2][16]/P0001  ;
	input \u11_mem_reg[2][17]/P0001  ;
	input \u11_mem_reg[2][18]/P0001  ;
	input \u11_mem_reg[2][19]/P0001  ;
	input \u11_mem_reg[2][1]/P0001  ;
	input \u11_mem_reg[2][20]/P0001  ;
	input \u11_mem_reg[2][21]/P0001  ;
	input \u11_mem_reg[2][22]/P0001  ;
	input \u11_mem_reg[2][23]/P0001  ;
	input \u11_mem_reg[2][24]/P0001  ;
	input \u11_mem_reg[2][25]/P0001  ;
	input \u11_mem_reg[2][26]/P0001  ;
	input \u11_mem_reg[2][27]/P0001  ;
	input \u11_mem_reg[2][28]/P0001  ;
	input \u11_mem_reg[2][29]/P0001  ;
	input \u11_mem_reg[2][2]/P0001  ;
	input \u11_mem_reg[2][30]/P0001  ;
	input \u11_mem_reg[2][31]/P0001  ;
	input \u11_mem_reg[2][3]/P0001  ;
	input \u11_mem_reg[2][4]/P0001  ;
	input \u11_mem_reg[2][5]/P0001  ;
	input \u11_mem_reg[2][6]/P0001  ;
	input \u11_mem_reg[2][7]/P0001  ;
	input \u11_mem_reg[2][8]/P0001  ;
	input \u11_mem_reg[2][9]/P0001  ;
	input \u11_mem_reg[3][0]/P0001  ;
	input \u11_mem_reg[3][10]/P0001  ;
	input \u11_mem_reg[3][11]/P0001  ;
	input \u11_mem_reg[3][12]/P0001  ;
	input \u11_mem_reg[3][13]/P0001  ;
	input \u11_mem_reg[3][14]/P0001  ;
	input \u11_mem_reg[3][15]/P0001  ;
	input \u11_mem_reg[3][16]/P0001  ;
	input \u11_mem_reg[3][17]/P0001  ;
	input \u11_mem_reg[3][18]/P0001  ;
	input \u11_mem_reg[3][19]/P0001  ;
	input \u11_mem_reg[3][1]/P0001  ;
	input \u11_mem_reg[3][20]/P0001  ;
	input \u11_mem_reg[3][21]/P0001  ;
	input \u11_mem_reg[3][22]/P0001  ;
	input \u11_mem_reg[3][23]/P0001  ;
	input \u11_mem_reg[3][24]/P0001  ;
	input \u11_mem_reg[3][25]/P0001  ;
	input \u11_mem_reg[3][26]/P0001  ;
	input \u11_mem_reg[3][27]/P0001  ;
	input \u11_mem_reg[3][28]/P0001  ;
	input \u11_mem_reg[3][29]/P0001  ;
	input \u11_mem_reg[3][2]/P0001  ;
	input \u11_mem_reg[3][30]/P0001  ;
	input \u11_mem_reg[3][31]/P0001  ;
	input \u11_mem_reg[3][3]/P0001  ;
	input \u11_mem_reg[3][4]/P0001  ;
	input \u11_mem_reg[3][5]/P0001  ;
	input \u11_mem_reg[3][6]/P0001  ;
	input \u11_mem_reg[3][7]/P0001  ;
	input \u11_mem_reg[3][8]/P0001  ;
	input \u11_mem_reg[3][9]/P0001  ;
	input \u11_rp_reg[0]/P0001  ;
	input \u11_rp_reg[1]/P0001  ;
	input \u11_rp_reg[2]/P0001  ;
	input \u11_status_reg[0]/P0001  ;
	input \u11_status_reg[1]/P0001  ;
	input \u11_wp_reg[0]/NET0131  ;
	input \u11_wp_reg[1]/P0001  ;
	input \u11_wp_reg[2]/P0001  ;
	input \u11_wp_reg[3]/P0001  ;
	input \u12_dout_reg[0]/P0001  ;
	input \u12_dout_reg[10]/P0001  ;
	input \u12_dout_reg[11]/P0001  ;
	input \u12_dout_reg[12]/P0001  ;
	input \u12_dout_reg[13]/P0001  ;
	input \u12_dout_reg[14]/P0001  ;
	input \u12_dout_reg[15]/P0001  ;
	input \u12_dout_reg[16]/P0001  ;
	input \u12_dout_reg[17]/P0001  ;
	input \u12_dout_reg[18]/P0001  ;
	input \u12_dout_reg[19]/P0001  ;
	input \u12_dout_reg[1]/P0001  ;
	input \u12_dout_reg[20]/P0001  ;
	input \u12_dout_reg[21]/P0001  ;
	input \u12_dout_reg[22]/P0001  ;
	input \u12_dout_reg[23]/P0001  ;
	input \u12_dout_reg[24]/P0001  ;
	input \u12_dout_reg[25]/P0001  ;
	input \u12_dout_reg[26]/P0001  ;
	input \u12_dout_reg[27]/P0001  ;
	input \u12_dout_reg[28]/P0001  ;
	input \u12_dout_reg[29]/P0001  ;
	input \u12_dout_reg[2]/P0001  ;
	input \u12_dout_reg[30]/P0001  ;
	input \u12_dout_reg[31]/P0001  ;
	input \u12_dout_reg[3]/P0001  ;
	input \u12_dout_reg[4]/P0001  ;
	input \u12_dout_reg[5]/P0001  ;
	input \u12_dout_reg[6]/P0001  ;
	input \u12_dout_reg[7]/P0001  ;
	input \u12_dout_reg[8]/P0001  ;
	input \u12_dout_reg[9]/P0001  ;
	input \u12_i3_re_reg/NET0131  ;
	input \u12_i4_re_reg/P0001  ;
	input \u12_i6_re_reg/NET0131  ;
	input \u12_o3_we_reg/P0001  ;
	input \u12_o4_we_reg/P0001  ;
	input \u12_o6_we_reg/P0001  ;
	input \u12_o7_we_reg/P0001  ;
	input \u12_o8_we_reg/P0001  ;
	input \u12_o9_we_reg/P0001  ;
	input \u12_re1_reg/P0001  ;
	input \u12_re2_reg/NET0131  ;
	input \u12_rf_we_reg/P0001  ;
	input \u12_we1_reg/P0001  ;
	input \u12_we2_reg/P0001  ;
	input \u13_ac97_rst_force_reg/P0001  ;
	input \u13_crac_dout_r_reg[0]/P0001  ;
	input \u13_crac_dout_r_reg[10]/P0001  ;
	input \u13_crac_dout_r_reg[11]/P0001  ;
	input \u13_crac_dout_r_reg[12]/P0001  ;
	input \u13_crac_dout_r_reg[13]/P0001  ;
	input \u13_crac_dout_r_reg[14]/P0001  ;
	input \u13_crac_dout_r_reg[15]/P0001  ;
	input \u13_crac_dout_r_reg[1]/P0001  ;
	input \u13_crac_dout_r_reg[2]/P0001  ;
	input \u13_crac_dout_r_reg[3]/P0001  ;
	input \u13_crac_dout_r_reg[4]/P0001  ;
	input \u13_crac_dout_r_reg[5]/P0001  ;
	input \u13_crac_dout_r_reg[6]/P0001  ;
	input \u13_crac_dout_r_reg[7]/P0001  ;
	input \u13_crac_dout_r_reg[8]/P0001  ;
	input \u13_crac_dout_r_reg[9]/P0001  ;
	input \u13_crac_r_reg[0]/NET0131  ;
	input \u13_crac_r_reg[1]/NET0131  ;
	input \u13_crac_r_reg[2]/NET0131  ;
	input \u13_crac_r_reg[3]/NET0131  ;
	input \u13_crac_r_reg[4]/NET0131  ;
	input \u13_crac_r_reg[5]/NET0131  ;
	input \u13_crac_r_reg[6]/NET0131  ;
	input \u13_crac_r_reg[7]/NET0131  ;
	input \u13_icc_r_reg[0]/NET0131  ;
	input \u13_icc_r_reg[10]/NET0131  ;
	input \u13_icc_r_reg[11]/NET0131  ;
	input \u13_icc_r_reg[12]/NET0131  ;
	input \u13_icc_r_reg[13]/NET0131  ;
	input \u13_icc_r_reg[14]/NET0131  ;
	input \u13_icc_r_reg[15]/NET0131  ;
	input \u13_icc_r_reg[16]/NET0131  ;
	input \u13_icc_r_reg[17]/NET0131  ;
	input \u13_icc_r_reg[18]/NET0131  ;
	input \u13_icc_r_reg[19]/NET0131  ;
	input \u13_icc_r_reg[1]/NET0131  ;
	input \u13_icc_r_reg[20]/NET0131  ;
	input \u13_icc_r_reg[21]/NET0131  ;
	input \u13_icc_r_reg[22]/NET0131  ;
	input \u13_icc_r_reg[23]/NET0131  ;
	input \u13_icc_r_reg[2]/NET0131  ;
	input \u13_icc_r_reg[3]/NET0131  ;
	input \u13_icc_r_reg[4]/NET0131  ;
	input \u13_icc_r_reg[5]/NET0131  ;
	input \u13_icc_r_reg[6]/NET0131  ;
	input \u13_icc_r_reg[7]/NET0131  ;
	input \u13_icc_r_reg[8]/NET0131  ;
	input \u13_icc_r_reg[9]/NET0131  ;
	input \u13_intm_r_reg[0]/NET0131  ;
	input \u13_intm_r_reg[10]/NET0131  ;
	input \u13_intm_r_reg[11]/NET0131  ;
	input \u13_intm_r_reg[12]/NET0131  ;
	input \u13_intm_r_reg[13]/NET0131  ;
	input \u13_intm_r_reg[14]/NET0131  ;
	input \u13_intm_r_reg[15]/NET0131  ;
	input \u13_intm_r_reg[16]/NET0131  ;
	input \u13_intm_r_reg[17]/NET0131  ;
	input \u13_intm_r_reg[18]/NET0131  ;
	input \u13_intm_r_reg[19]/NET0131  ;
	input \u13_intm_r_reg[1]/NET0131  ;
	input \u13_intm_r_reg[20]/NET0131  ;
	input \u13_intm_r_reg[21]/NET0131  ;
	input \u13_intm_r_reg[22]/NET0131  ;
	input \u13_intm_r_reg[23]/NET0131  ;
	input \u13_intm_r_reg[24]/NET0131  ;
	input \u13_intm_r_reg[25]/NET0131  ;
	input \u13_intm_r_reg[26]/NET0131  ;
	input \u13_intm_r_reg[27]/NET0131  ;
	input \u13_intm_r_reg[28]/NET0131  ;
	input \u13_intm_r_reg[2]/NET0131  ;
	input \u13_intm_r_reg[3]/NET0131  ;
	input \u13_intm_r_reg[4]/NET0131  ;
	input \u13_intm_r_reg[5]/NET0131  ;
	input \u13_intm_r_reg[6]/NET0131  ;
	input \u13_intm_r_reg[7]/NET0131  ;
	input \u13_intm_r_reg[8]/NET0131  ;
	input \u13_intm_r_reg[9]/NET0131  ;
	input \u13_ints_r_reg[0]/NET0131  ;
	input \u13_ints_r_reg[10]/NET0131  ;
	input \u13_ints_r_reg[11]/NET0131  ;
	input \u13_ints_r_reg[12]/NET0131  ;
	input \u13_ints_r_reg[13]/NET0131  ;
	input \u13_ints_r_reg[14]/NET0131  ;
	input \u13_ints_r_reg[15]/NET0131  ;
	input \u13_ints_r_reg[16]/NET0131  ;
	input \u13_ints_r_reg[17]/NET0131  ;
	input \u13_ints_r_reg[18]/NET0131  ;
	input \u13_ints_r_reg[19]/NET0131  ;
	input \u13_ints_r_reg[1]/NET0131  ;
	input \u13_ints_r_reg[20]/NET0131  ;
	input \u13_ints_r_reg[21]/NET0131  ;
	input \u13_ints_r_reg[22]/NET0131  ;
	input \u13_ints_r_reg[23]/NET0131  ;
	input \u13_ints_r_reg[24]/NET0131  ;
	input \u13_ints_r_reg[25]/NET0131  ;
	input \u13_ints_r_reg[26]/NET0131  ;
	input \u13_ints_r_reg[27]/NET0131  ;
	input \u13_ints_r_reg[28]/NET0131  ;
	input \u13_ints_r_reg[2]/NET0131  ;
	input \u13_ints_r_reg[3]/NET0131  ;
	input \u13_ints_r_reg[4]/NET0131  ;
	input \u13_ints_r_reg[5]/NET0131  ;
	input \u13_ints_r_reg[6]/NET0131  ;
	input \u13_ints_r_reg[7]/NET0131  ;
	input \u13_ints_r_reg[8]/NET0131  ;
	input \u13_ints_r_reg[9]/NET0131  ;
	input \u13_occ0_r_reg[0]/NET0131  ;
	input \u13_occ0_r_reg[10]/NET0131  ;
	input \u13_occ0_r_reg[11]/NET0131  ;
	input \u13_occ0_r_reg[12]/NET0131  ;
	input \u13_occ0_r_reg[13]/NET0131  ;
	input \u13_occ0_r_reg[14]/NET0131  ;
	input \u13_occ0_r_reg[15]/NET0131  ;
	input \u13_occ0_r_reg[16]/NET0131  ;
	input \u13_occ0_r_reg[17]/NET0131  ;
	input \u13_occ0_r_reg[18]/NET0131  ;
	input \u13_occ0_r_reg[19]/NET0131  ;
	input \u13_occ0_r_reg[1]/NET0131  ;
	input \u13_occ0_r_reg[20]/NET0131  ;
	input \u13_occ0_r_reg[21]/NET0131  ;
	input \u13_occ0_r_reg[22]/NET0131  ;
	input \u13_occ0_r_reg[23]/NET0131  ;
	input \u13_occ0_r_reg[24]/NET0131  ;
	input \u13_occ0_r_reg[25]/NET0131  ;
	input \u13_occ0_r_reg[26]/NET0131  ;
	input \u13_occ0_r_reg[27]/NET0131  ;
	input \u13_occ0_r_reg[28]/NET0131  ;
	input \u13_occ0_r_reg[29]/NET0131  ;
	input \u13_occ0_r_reg[2]/NET0131  ;
	input \u13_occ0_r_reg[30]/NET0131  ;
	input \u13_occ0_r_reg[31]/NET0131  ;
	input \u13_occ0_r_reg[3]/NET0131  ;
	input \u13_occ0_r_reg[4]/NET0131  ;
	input \u13_occ0_r_reg[5]/NET0131  ;
	input \u13_occ0_r_reg[6]/NET0131  ;
	input \u13_occ0_r_reg[7]/NET0131  ;
	input \u13_occ0_r_reg[8]/NET0131  ;
	input \u13_occ0_r_reg[9]/NET0131  ;
	input \u13_occ1_r_reg[0]/NET0131  ;
	input \u13_occ1_r_reg[10]/NET0131  ;
	input \u13_occ1_r_reg[11]/NET0131  ;
	input \u13_occ1_r_reg[12]/NET0131  ;
	input \u13_occ1_r_reg[13]/NET0131  ;
	input \u13_occ1_r_reg[14]/NET0131  ;
	input \u13_occ1_r_reg[15]/NET0131  ;
	input \u13_occ1_r_reg[1]/NET0131  ;
	input \u13_occ1_r_reg[2]/NET0131  ;
	input \u13_occ1_r_reg[3]/NET0131  ;
	input \u13_occ1_r_reg[4]/NET0131  ;
	input \u13_occ1_r_reg[5]/NET0131  ;
	input \u13_occ1_r_reg[6]/NET0131  ;
	input \u13_occ1_r_reg[7]/NET0131  ;
	input \u13_occ1_r_reg[8]/NET0131  ;
	input \u13_occ1_r_reg[9]/NET0131  ;
	input \u13_resume_req_reg/P0001  ;
	input \u14_crac_valid_r_reg/P0001  ;
	input \u14_crac_wr_r_reg/P0001  ;
	input \u14_u0_en_out_l2_reg/P0001  ;
	input \u14_u0_en_out_l_reg/NET0131  ;
	input \u14_u0_full_empty_r_reg/P0001  ;
	input \u14_u1_en_out_l2_reg/P0001  ;
	input \u14_u1_en_out_l_reg/NET0131  ;
	input \u14_u1_full_empty_r_reg/P0001  ;
	input \u14_u2_en_out_l2_reg/P0001  ;
	input \u14_u2_en_out_l_reg/NET0131  ;
	input \u14_u2_full_empty_r_reg/P0001  ;
	input \u14_u3_en_out_l2_reg/P0001  ;
	input \u14_u3_en_out_l_reg/NET0131  ;
	input \u14_u3_full_empty_r_reg/P0001  ;
	input \u14_u4_en_out_l2_reg/P0001  ;
	input \u14_u4_en_out_l_reg/NET0131  ;
	input \u14_u4_full_empty_r_reg/P0001  ;
	input \u14_u5_en_out_l2_reg/P0001  ;
	input \u14_u5_en_out_l_reg/NET0131  ;
	input \u14_u5_full_empty_r_reg/P0001  ;
	input \u14_u6_en_out_l2_reg/P0001  ;
	input \u14_u6_en_out_l_reg/NET0131  ;
	input \u14_u6_full_empty_r_reg/P0001  ;
	input \u14_u7_en_out_l2_reg/P0001  ;
	input \u14_u7_en_out_l_reg/NET0131  ;
	input \u14_u7_full_empty_r_reg/P0001  ;
	input \u14_u8_en_out_l2_reg/P0001  ;
	input \u14_u8_en_out_l_reg/NET0131  ;
	input \u14_u8_full_empty_r_reg/P0001  ;
	input \u15_crac_din_reg[0]/NET0131  ;
	input \u15_crac_din_reg[10]/NET0131  ;
	input \u15_crac_din_reg[11]/NET0131  ;
	input \u15_crac_din_reg[12]/NET0131  ;
	input \u15_crac_din_reg[13]/NET0131  ;
	input \u15_crac_din_reg[14]/NET0131  ;
	input \u15_crac_din_reg[15]/NET0131  ;
	input \u15_crac_din_reg[1]/NET0131  ;
	input \u15_crac_din_reg[2]/NET0131  ;
	input \u15_crac_din_reg[3]/NET0131  ;
	input \u15_crac_din_reg[4]/NET0131  ;
	input \u15_crac_din_reg[5]/NET0131  ;
	input \u15_crac_din_reg[6]/NET0131  ;
	input \u15_crac_din_reg[7]/NET0131  ;
	input \u15_crac_din_reg[8]/NET0131  ;
	input \u15_crac_din_reg[9]/NET0131  ;
	input \u15_crac_rd_done_reg/P0001  ;
	input \u15_crac_rd_reg/NET0131  ;
	input \u15_crac_we_r_reg/P0001  ;
	input \u15_crac_wr_reg/NET0131  ;
	input \u15_rdd1_reg/NET0131  ;
	input \u15_rdd2_reg/NET0131  ;
	input \u15_rdd3_reg/NET0131  ;
	input \u15_valid_r_reg/P0001  ;
	input \u16_u0_dma_req_r1_reg/P0001  ;
	input \u16_u1_dma_req_r1_reg/P0001  ;
	input \u16_u2_dma_req_r1_reg/P0001  ;
	input \u16_u3_dma_req_r1_reg/P0001  ;
	input \u16_u4_dma_req_r1_reg/P0001  ;
	input \u16_u5_dma_req_r1_reg/P0001  ;
	input \u16_u6_dma_req_r1_reg/P0001  ;
	input \u16_u7_dma_req_r1_reg/P0001  ;
	input \u16_u8_dma_req_r1_reg/P0001  ;
	input \u17_int_set_reg[0]/NET0131  ;
	input \u17_int_set_reg[1]/NET0131  ;
	input \u17_int_set_reg[2]/NET0131  ;
	input \u18_int_set_reg[0]/NET0131  ;
	input \u18_int_set_reg[1]/NET0131  ;
	input \u18_int_set_reg[2]/NET0131  ;
	input \u19_int_set_reg[0]/NET0131  ;
	input \u19_int_set_reg[1]/NET0131  ;
	input \u19_int_set_reg[2]/NET0131  ;
	input \u1_slt0_reg[11]/P0001  ;
	input \u1_slt0_reg[12]/P0001  ;
	input \u1_slt0_reg[15]/P0001  ;
	input \u1_slt0_reg[9]/P0001  ;
	input \u1_slt1_reg[10]/P0001  ;
	input \u1_slt1_reg[11]/P0001  ;
	input \u1_slt1_reg[5]/P0001  ;
	input \u1_slt1_reg[6]/P0001  ;
	input \u1_slt1_reg[7]/P0001  ;
	input \u1_slt1_reg[8]/P0001  ;
	input \u1_slt3_reg[0]/P0001  ;
	input \u1_slt3_reg[10]/P0001  ;
	input \u1_slt3_reg[11]/P0001  ;
	input \u1_slt3_reg[12]/P0001  ;
	input \u1_slt3_reg[13]/P0001  ;
	input \u1_slt3_reg[14]/P0001  ;
	input \u1_slt3_reg[15]/P0001  ;
	input \u1_slt3_reg[16]/P0001  ;
	input \u1_slt3_reg[17]/P0001  ;
	input \u1_slt3_reg[18]/P0001  ;
	input \u1_slt3_reg[19]/P0001  ;
	input \u1_slt3_reg[1]/P0001  ;
	input \u1_slt3_reg[2]/P0001  ;
	input \u1_slt3_reg[3]/P0001  ;
	input \u1_slt3_reg[4]/P0001  ;
	input \u1_slt3_reg[5]/P0001  ;
	input \u1_slt3_reg[6]/P0001  ;
	input \u1_slt3_reg[7]/P0001  ;
	input \u1_slt3_reg[8]/P0001  ;
	input \u1_slt3_reg[9]/P0001  ;
	input \u1_slt4_reg[0]/P0001  ;
	input \u1_slt4_reg[10]/P0001  ;
	input \u1_slt4_reg[11]/P0001  ;
	input \u1_slt4_reg[12]/P0001  ;
	input \u1_slt4_reg[13]/P0001  ;
	input \u1_slt4_reg[14]/P0001  ;
	input \u1_slt4_reg[15]/P0001  ;
	input \u1_slt4_reg[16]/P0001  ;
	input \u1_slt4_reg[17]/P0001  ;
	input \u1_slt4_reg[18]/P0001  ;
	input \u1_slt4_reg[19]/P0001  ;
	input \u1_slt4_reg[1]/P0001  ;
	input \u1_slt4_reg[2]/P0001  ;
	input \u1_slt4_reg[3]/P0001  ;
	input \u1_slt4_reg[4]/P0001  ;
	input \u1_slt4_reg[5]/P0001  ;
	input \u1_slt4_reg[6]/P0001  ;
	input \u1_slt4_reg[7]/P0001  ;
	input \u1_slt4_reg[8]/P0001  ;
	input \u1_slt4_reg[9]/P0001  ;
	input \u1_slt6_reg[0]/P0001  ;
	input \u1_slt6_reg[10]/P0001  ;
	input \u1_slt6_reg[11]/P0001  ;
	input \u1_slt6_reg[12]/P0001  ;
	input \u1_slt6_reg[13]/P0001  ;
	input \u1_slt6_reg[14]/P0001  ;
	input \u1_slt6_reg[15]/P0001  ;
	input \u1_slt6_reg[16]/P0001  ;
	input \u1_slt6_reg[17]/P0001  ;
	input \u1_slt6_reg[18]/P0001  ;
	input \u1_slt6_reg[19]/P0001  ;
	input \u1_slt6_reg[1]/P0001  ;
	input \u1_slt6_reg[2]/P0001  ;
	input \u1_slt6_reg[3]/P0001  ;
	input \u1_slt6_reg[4]/P0001  ;
	input \u1_slt6_reg[5]/P0001  ;
	input \u1_slt6_reg[6]/P0001  ;
	input \u1_slt6_reg[7]/P0001  ;
	input \u1_slt6_reg[8]/P0001  ;
	input \u1_slt6_reg[9]/P0001  ;
	input \u1_sr_reg[10]/P0001  ;
	input \u1_sr_reg[11]/P0001  ;
	input \u1_sr_reg[12]/P0001  ;
	input \u1_sr_reg[15]/P0001  ;
	input \u1_sr_reg[5]/P0001  ;
	input \u1_sr_reg[6]/P0001  ;
	input \u1_sr_reg[7]/P0001  ;
	input \u1_sr_reg[8]/P0001  ;
	input \u1_sr_reg[9]/P0001  ;
	input \u20_int_set_reg[0]/NET0131  ;
	input \u20_int_set_reg[1]/NET0131  ;
	input \u20_int_set_reg[2]/NET0131  ;
	input \u21_int_set_reg[0]/NET0131  ;
	input \u21_int_set_reg[1]/NET0131  ;
	input \u21_int_set_reg[2]/NET0131  ;
	input \u22_int_set_reg[0]/NET0131  ;
	input \u22_int_set_reg[1]/NET0131  ;
	input \u22_int_set_reg[2]/NET0131  ;
	input \u23_int_set_reg[0]/NET0131  ;
	input \u23_int_set_reg[1]/NET0131  ;
	input \u23_int_set_reg[2]/NET0131  ;
	input \u24_int_set_reg[0]/NET0131  ;
	input \u24_int_set_reg[1]/NET0131  ;
	input \u24_int_set_reg[2]/NET0131  ;
	input \u25_int_set_reg[0]/NET0131  ;
	input \u25_int_set_reg[1]/NET0131  ;
	input \u25_int_set_reg[2]/NET0131  ;
	input \u26_cnt_reg[0]/NET0131  ;
	input \u26_cnt_reg[1]/NET0131  ;
	input \u26_cnt_reg[2]/NET0131  ;
	input \u26_ps_cnt_reg[0]/NET0131  ;
	input \u26_ps_cnt_reg[1]/NET0131  ;
	input \u26_ps_cnt_reg[2]/NET0131  ;
	input \u26_ps_cnt_reg[3]/NET0131  ;
	input \u26_ps_cnt_reg[4]/NET0131  ;
	input \u26_ps_cnt_reg[5]/NET0131  ;
	input \u2_bit_clk_e_reg/P0001  ;
	input \u2_bit_clk_r1_reg/P0001  ;
	input \u2_bit_clk_r_reg/P0001  ;
	input \u2_cnt_reg[0]/NET0131  ;
	input \u2_cnt_reg[1]/NET0131  ;
	input \u2_cnt_reg[2]/NET0131  ;
	input \u2_cnt_reg[3]/NET0131  ;
	input \u2_cnt_reg[4]/NET0131  ;
	input \u2_cnt_reg[5]/NET0131  ;
	input \u2_cnt_reg[6]/NET0131  ;
	input \u2_cnt_reg[7]/NET0131  ;
	input \u2_ld_reg/P0001  ;
	input \u2_out_le_reg[0]/P0001  ;
	input \u2_out_le_reg[1]/P0001  ;
	input \u2_res_cnt_reg[0]/P0001  ;
	input \u2_res_cnt_reg[1]/P0001  ;
	input \u2_res_cnt_reg[2]/P0001  ;
	input \u2_res_cnt_reg[3]/P0001  ;
	input \u2_sync_beat_reg/P0001  ;
	input \u2_sync_resume_reg/NET0131  ;
	input \u2_to_cnt_reg[0]/NET0131  ;
	input \u2_to_cnt_reg[1]/NET0131  ;
	input \u2_to_cnt_reg[2]/NET0131  ;
	input \u2_to_cnt_reg[3]/NET0131  ;
	input \u2_to_cnt_reg[4]/NET0131  ;
	input \u2_to_cnt_reg[5]/NET0131  ;
	input \u3_dout_reg[0]/P0001  ;
	input \u3_dout_reg[10]/P0001  ;
	input \u3_dout_reg[11]/P0001  ;
	input \u3_dout_reg[12]/P0001  ;
	input \u3_dout_reg[13]/P0001  ;
	input \u3_dout_reg[14]/P0001  ;
	input \u3_dout_reg[15]/P0001  ;
	input \u3_dout_reg[16]/P0001  ;
	input \u3_dout_reg[17]/P0001  ;
	input \u3_dout_reg[18]/P0001  ;
	input \u3_dout_reg[19]/P0001  ;
	input \u3_dout_reg[1]/P0001  ;
	input \u3_dout_reg[2]/P0001  ;
	input \u3_dout_reg[3]/P0001  ;
	input \u3_dout_reg[4]/P0001  ;
	input \u3_dout_reg[5]/P0001  ;
	input \u3_dout_reg[6]/P0001  ;
	input \u3_dout_reg[7]/P0001  ;
	input \u3_dout_reg[8]/P0001  ;
	input \u3_dout_reg[9]/P0001  ;
	input \u3_empty_reg/NET0131  ;
	input \u3_mem_reg[0][0]/NET0131  ;
	input \u3_mem_reg[0][10]/NET0131  ;
	input \u3_mem_reg[0][11]/NET0131  ;
	input \u3_mem_reg[0][12]/NET0131  ;
	input \u3_mem_reg[0][13]/NET0131  ;
	input \u3_mem_reg[0][14]/NET0131  ;
	input \u3_mem_reg[0][15]/NET0131  ;
	input \u3_mem_reg[0][16]/NET0131  ;
	input \u3_mem_reg[0][17]/NET0131  ;
	input \u3_mem_reg[0][18]/NET0131  ;
	input \u3_mem_reg[0][19]/NET0131  ;
	input \u3_mem_reg[0][1]/NET0131  ;
	input \u3_mem_reg[0][20]/NET0131  ;
	input \u3_mem_reg[0][21]/NET0131  ;
	input \u3_mem_reg[0][22]/NET0131  ;
	input \u3_mem_reg[0][23]/NET0131  ;
	input \u3_mem_reg[0][24]/NET0131  ;
	input \u3_mem_reg[0][25]/NET0131  ;
	input \u3_mem_reg[0][26]/NET0131  ;
	input \u3_mem_reg[0][27]/NET0131  ;
	input \u3_mem_reg[0][28]/NET0131  ;
	input \u3_mem_reg[0][29]/NET0131  ;
	input \u3_mem_reg[0][2]/NET0131  ;
	input \u3_mem_reg[0][30]/NET0131  ;
	input \u3_mem_reg[0][31]/NET0131  ;
	input \u3_mem_reg[0][3]/NET0131  ;
	input \u3_mem_reg[0][4]/NET0131  ;
	input \u3_mem_reg[0][5]/NET0131  ;
	input \u3_mem_reg[0][6]/NET0131  ;
	input \u3_mem_reg[0][7]/NET0131  ;
	input \u3_mem_reg[0][8]/NET0131  ;
	input \u3_mem_reg[0][9]/NET0131  ;
	input \u3_mem_reg[1][0]/NET0131  ;
	input \u3_mem_reg[1][10]/NET0131  ;
	input \u3_mem_reg[1][11]/NET0131  ;
	input \u3_mem_reg[1][12]/NET0131  ;
	input \u3_mem_reg[1][13]/NET0131  ;
	input \u3_mem_reg[1][14]/NET0131  ;
	input \u3_mem_reg[1][15]/NET0131  ;
	input \u3_mem_reg[1][16]/NET0131  ;
	input \u3_mem_reg[1][17]/NET0131  ;
	input \u3_mem_reg[1][18]/NET0131  ;
	input \u3_mem_reg[1][19]/NET0131  ;
	input \u3_mem_reg[1][1]/NET0131  ;
	input \u3_mem_reg[1][20]/NET0131  ;
	input \u3_mem_reg[1][21]/NET0131  ;
	input \u3_mem_reg[1][22]/NET0131  ;
	input \u3_mem_reg[1][23]/NET0131  ;
	input \u3_mem_reg[1][24]/NET0131  ;
	input \u3_mem_reg[1][25]/NET0131  ;
	input \u3_mem_reg[1][26]/NET0131  ;
	input \u3_mem_reg[1][27]/NET0131  ;
	input \u3_mem_reg[1][28]/NET0131  ;
	input \u3_mem_reg[1][29]/NET0131  ;
	input \u3_mem_reg[1][2]/NET0131  ;
	input \u3_mem_reg[1][30]/NET0131  ;
	input \u3_mem_reg[1][31]/NET0131  ;
	input \u3_mem_reg[1][3]/NET0131  ;
	input \u3_mem_reg[1][4]/NET0131  ;
	input \u3_mem_reg[1][5]/NET0131  ;
	input \u3_mem_reg[1][6]/NET0131  ;
	input \u3_mem_reg[1][7]/NET0131  ;
	input \u3_mem_reg[1][8]/NET0131  ;
	input \u3_mem_reg[1][9]/NET0131  ;
	input \u3_mem_reg[2][0]/NET0131  ;
	input \u3_mem_reg[2][10]/NET0131  ;
	input \u3_mem_reg[2][11]/NET0131  ;
	input \u3_mem_reg[2][12]/NET0131  ;
	input \u3_mem_reg[2][13]/NET0131  ;
	input \u3_mem_reg[2][14]/NET0131  ;
	input \u3_mem_reg[2][15]/NET0131  ;
	input \u3_mem_reg[2][16]/NET0131  ;
	input \u3_mem_reg[2][17]/NET0131  ;
	input \u3_mem_reg[2][18]/NET0131  ;
	input \u3_mem_reg[2][19]/NET0131  ;
	input \u3_mem_reg[2][1]/NET0131  ;
	input \u3_mem_reg[2][20]/NET0131  ;
	input \u3_mem_reg[2][21]/NET0131  ;
	input \u3_mem_reg[2][22]/NET0131  ;
	input \u3_mem_reg[2][23]/NET0131  ;
	input \u3_mem_reg[2][24]/NET0131  ;
	input \u3_mem_reg[2][25]/NET0131  ;
	input \u3_mem_reg[2][26]/NET0131  ;
	input \u3_mem_reg[2][27]/NET0131  ;
	input \u3_mem_reg[2][28]/NET0131  ;
	input \u3_mem_reg[2][29]/NET0131  ;
	input \u3_mem_reg[2][2]/NET0131  ;
	input \u3_mem_reg[2][30]/NET0131  ;
	input \u3_mem_reg[2][31]/NET0131  ;
	input \u3_mem_reg[2][3]/NET0131  ;
	input \u3_mem_reg[2][4]/NET0131  ;
	input \u3_mem_reg[2][5]/NET0131  ;
	input \u3_mem_reg[2][6]/NET0131  ;
	input \u3_mem_reg[2][7]/NET0131  ;
	input \u3_mem_reg[2][8]/NET0131  ;
	input \u3_mem_reg[2][9]/NET0131  ;
	input \u3_mem_reg[3][0]/NET0131  ;
	input \u3_mem_reg[3][10]/NET0131  ;
	input \u3_mem_reg[3][11]/NET0131  ;
	input \u3_mem_reg[3][12]/NET0131  ;
	input \u3_mem_reg[3][13]/NET0131  ;
	input \u3_mem_reg[3][14]/NET0131  ;
	input \u3_mem_reg[3][15]/NET0131  ;
	input \u3_mem_reg[3][16]/NET0131  ;
	input \u3_mem_reg[3][17]/NET0131  ;
	input \u3_mem_reg[3][18]/NET0131  ;
	input \u3_mem_reg[3][19]/NET0131  ;
	input \u3_mem_reg[3][1]/NET0131  ;
	input \u3_mem_reg[3][20]/NET0131  ;
	input \u3_mem_reg[3][21]/NET0131  ;
	input \u3_mem_reg[3][22]/NET0131  ;
	input \u3_mem_reg[3][23]/NET0131  ;
	input \u3_mem_reg[3][24]/NET0131  ;
	input \u3_mem_reg[3][25]/NET0131  ;
	input \u3_mem_reg[3][26]/NET0131  ;
	input \u3_mem_reg[3][27]/NET0131  ;
	input \u3_mem_reg[3][28]/NET0131  ;
	input \u3_mem_reg[3][29]/NET0131  ;
	input \u3_mem_reg[3][2]/NET0131  ;
	input \u3_mem_reg[3][30]/NET0131  ;
	input \u3_mem_reg[3][31]/NET0131  ;
	input \u3_mem_reg[3][3]/NET0131  ;
	input \u3_mem_reg[3][4]/NET0131  ;
	input \u3_mem_reg[3][5]/NET0131  ;
	input \u3_mem_reg[3][6]/NET0131  ;
	input \u3_mem_reg[3][7]/NET0131  ;
	input \u3_mem_reg[3][8]/NET0131  ;
	input \u3_mem_reg[3][9]/NET0131  ;
	input \u3_rp_reg[0]/P0001  ;
	input \u3_rp_reg[1]/NET0131  ;
	input \u3_rp_reg[2]/NET0131  ;
	input \u3_rp_reg[3]/NET0131  ;
	input \u3_status_reg[0]/P0001  ;
	input \u3_status_reg[1]/P0001  ;
	input \u3_wp_reg[0]/P0001  ;
	input \u3_wp_reg[1]/NET0131  ;
	input \u3_wp_reg[2]/P0001  ;
	input \u4_dout_reg[0]/P0001  ;
	input \u4_dout_reg[10]/P0001  ;
	input \u4_dout_reg[11]/P0001  ;
	input \u4_dout_reg[12]/P0001  ;
	input \u4_dout_reg[13]/P0001  ;
	input \u4_dout_reg[14]/P0001  ;
	input \u4_dout_reg[15]/P0001  ;
	input \u4_dout_reg[16]/P0001  ;
	input \u4_dout_reg[17]/P0001  ;
	input \u4_dout_reg[18]/P0001  ;
	input \u4_dout_reg[19]/P0001  ;
	input \u4_dout_reg[1]/P0001  ;
	input \u4_dout_reg[2]/P0001  ;
	input \u4_dout_reg[3]/P0001  ;
	input \u4_dout_reg[4]/P0001  ;
	input \u4_dout_reg[5]/P0001  ;
	input \u4_dout_reg[6]/P0001  ;
	input \u4_dout_reg[7]/P0001  ;
	input \u4_dout_reg[8]/P0001  ;
	input \u4_dout_reg[9]/P0001  ;
	input \u4_empty_reg/NET0131  ;
	input \u4_mem_reg[0][0]/NET0131  ;
	input \u4_mem_reg[0][10]/NET0131  ;
	input \u4_mem_reg[0][11]/NET0131  ;
	input \u4_mem_reg[0][12]/NET0131  ;
	input \u4_mem_reg[0][13]/NET0131  ;
	input \u4_mem_reg[0][14]/NET0131  ;
	input \u4_mem_reg[0][15]/NET0131  ;
	input \u4_mem_reg[0][16]/NET0131  ;
	input \u4_mem_reg[0][17]/NET0131  ;
	input \u4_mem_reg[0][18]/NET0131  ;
	input \u4_mem_reg[0][19]/NET0131  ;
	input \u4_mem_reg[0][1]/NET0131  ;
	input \u4_mem_reg[0][20]/NET0131  ;
	input \u4_mem_reg[0][21]/NET0131  ;
	input \u4_mem_reg[0][22]/NET0131  ;
	input \u4_mem_reg[0][23]/NET0131  ;
	input \u4_mem_reg[0][24]/NET0131  ;
	input \u4_mem_reg[0][25]/NET0131  ;
	input \u4_mem_reg[0][26]/NET0131  ;
	input \u4_mem_reg[0][27]/NET0131  ;
	input \u4_mem_reg[0][28]/NET0131  ;
	input \u4_mem_reg[0][29]/NET0131  ;
	input \u4_mem_reg[0][2]/NET0131  ;
	input \u4_mem_reg[0][30]/NET0131  ;
	input \u4_mem_reg[0][31]/NET0131  ;
	input \u4_mem_reg[0][3]/NET0131  ;
	input \u4_mem_reg[0][4]/NET0131  ;
	input \u4_mem_reg[0][5]/NET0131  ;
	input \u4_mem_reg[0][6]/NET0131  ;
	input \u4_mem_reg[0][7]/NET0131  ;
	input \u4_mem_reg[0][8]/NET0131  ;
	input \u4_mem_reg[0][9]/NET0131  ;
	input \u4_mem_reg[1][0]/NET0131  ;
	input \u4_mem_reg[1][10]/NET0131  ;
	input \u4_mem_reg[1][11]/NET0131  ;
	input \u4_mem_reg[1][12]/NET0131  ;
	input \u4_mem_reg[1][13]/NET0131  ;
	input \u4_mem_reg[1][14]/NET0131  ;
	input \u4_mem_reg[1][15]/NET0131  ;
	input \u4_mem_reg[1][16]/NET0131  ;
	input \u4_mem_reg[1][17]/NET0131  ;
	input \u4_mem_reg[1][18]/NET0131  ;
	input \u4_mem_reg[1][19]/NET0131  ;
	input \u4_mem_reg[1][1]/NET0131  ;
	input \u4_mem_reg[1][20]/NET0131  ;
	input \u4_mem_reg[1][21]/NET0131  ;
	input \u4_mem_reg[1][22]/NET0131  ;
	input \u4_mem_reg[1][23]/NET0131  ;
	input \u4_mem_reg[1][24]/NET0131  ;
	input \u4_mem_reg[1][25]/NET0131  ;
	input \u4_mem_reg[1][26]/NET0131  ;
	input \u4_mem_reg[1][27]/NET0131  ;
	input \u4_mem_reg[1][28]/NET0131  ;
	input \u4_mem_reg[1][29]/NET0131  ;
	input \u4_mem_reg[1][2]/NET0131  ;
	input \u4_mem_reg[1][30]/NET0131  ;
	input \u4_mem_reg[1][31]/NET0131  ;
	input \u4_mem_reg[1][3]/NET0131  ;
	input \u4_mem_reg[1][4]/NET0131  ;
	input \u4_mem_reg[1][5]/NET0131  ;
	input \u4_mem_reg[1][6]/NET0131  ;
	input \u4_mem_reg[1][7]/NET0131  ;
	input \u4_mem_reg[1][8]/NET0131  ;
	input \u4_mem_reg[1][9]/NET0131  ;
	input \u4_mem_reg[2][0]/NET0131  ;
	input \u4_mem_reg[2][10]/NET0131  ;
	input \u4_mem_reg[2][11]/NET0131  ;
	input \u4_mem_reg[2][12]/NET0131  ;
	input \u4_mem_reg[2][13]/NET0131  ;
	input \u4_mem_reg[2][14]/NET0131  ;
	input \u4_mem_reg[2][15]/NET0131  ;
	input \u4_mem_reg[2][16]/NET0131  ;
	input \u4_mem_reg[2][17]/NET0131  ;
	input \u4_mem_reg[2][18]/NET0131  ;
	input \u4_mem_reg[2][19]/NET0131  ;
	input \u4_mem_reg[2][1]/NET0131  ;
	input \u4_mem_reg[2][20]/NET0131  ;
	input \u4_mem_reg[2][21]/NET0131  ;
	input \u4_mem_reg[2][22]/NET0131  ;
	input \u4_mem_reg[2][23]/NET0131  ;
	input \u4_mem_reg[2][24]/NET0131  ;
	input \u4_mem_reg[2][25]/NET0131  ;
	input \u4_mem_reg[2][26]/NET0131  ;
	input \u4_mem_reg[2][27]/NET0131  ;
	input \u4_mem_reg[2][28]/NET0131  ;
	input \u4_mem_reg[2][29]/NET0131  ;
	input \u4_mem_reg[2][2]/NET0131  ;
	input \u4_mem_reg[2][30]/NET0131  ;
	input \u4_mem_reg[2][31]/NET0131  ;
	input \u4_mem_reg[2][3]/NET0131  ;
	input \u4_mem_reg[2][4]/NET0131  ;
	input \u4_mem_reg[2][5]/NET0131  ;
	input \u4_mem_reg[2][6]/NET0131  ;
	input \u4_mem_reg[2][7]/NET0131  ;
	input \u4_mem_reg[2][8]/NET0131  ;
	input \u4_mem_reg[2][9]/NET0131  ;
	input \u4_mem_reg[3][0]/NET0131  ;
	input \u4_mem_reg[3][10]/NET0131  ;
	input \u4_mem_reg[3][11]/NET0131  ;
	input \u4_mem_reg[3][12]/NET0131  ;
	input \u4_mem_reg[3][13]/NET0131  ;
	input \u4_mem_reg[3][14]/NET0131  ;
	input \u4_mem_reg[3][15]/NET0131  ;
	input \u4_mem_reg[3][16]/NET0131  ;
	input \u4_mem_reg[3][17]/NET0131  ;
	input \u4_mem_reg[3][18]/NET0131  ;
	input \u4_mem_reg[3][19]/NET0131  ;
	input \u4_mem_reg[3][1]/NET0131  ;
	input \u4_mem_reg[3][20]/NET0131  ;
	input \u4_mem_reg[3][21]/NET0131  ;
	input \u4_mem_reg[3][22]/NET0131  ;
	input \u4_mem_reg[3][23]/NET0131  ;
	input \u4_mem_reg[3][24]/NET0131  ;
	input \u4_mem_reg[3][25]/NET0131  ;
	input \u4_mem_reg[3][26]/NET0131  ;
	input \u4_mem_reg[3][27]/NET0131  ;
	input \u4_mem_reg[3][28]/NET0131  ;
	input \u4_mem_reg[3][29]/NET0131  ;
	input \u4_mem_reg[3][2]/NET0131  ;
	input \u4_mem_reg[3][30]/NET0131  ;
	input \u4_mem_reg[3][31]/NET0131  ;
	input \u4_mem_reg[3][3]/NET0131  ;
	input \u4_mem_reg[3][4]/NET0131  ;
	input \u4_mem_reg[3][5]/NET0131  ;
	input \u4_mem_reg[3][6]/NET0131  ;
	input \u4_mem_reg[3][7]/NET0131  ;
	input \u4_mem_reg[3][8]/NET0131  ;
	input \u4_mem_reg[3][9]/NET0131  ;
	input \u4_rp_reg[0]/P0001  ;
	input \u4_rp_reg[1]/NET0131  ;
	input \u4_rp_reg[2]/NET0131  ;
	input \u4_rp_reg[3]/NET0131  ;
	input \u4_status_reg[0]/P0001  ;
	input \u4_status_reg[1]/P0001  ;
	input \u4_wp_reg[0]/P0001  ;
	input \u4_wp_reg[1]/NET0131  ;
	input \u4_wp_reg[2]/P0001  ;
	input \u5_dout_reg[0]/P0001  ;
	input \u5_dout_reg[10]/P0001  ;
	input \u5_dout_reg[11]/P0001  ;
	input \u5_dout_reg[12]/P0001  ;
	input \u5_dout_reg[13]/P0001  ;
	input \u5_dout_reg[14]/P0001  ;
	input \u5_dout_reg[15]/P0001  ;
	input \u5_dout_reg[16]/P0001  ;
	input \u5_dout_reg[17]/P0001  ;
	input \u5_dout_reg[18]/P0001  ;
	input \u5_dout_reg[19]/P0001  ;
	input \u5_dout_reg[1]/P0001  ;
	input \u5_dout_reg[2]/P0001  ;
	input \u5_dout_reg[3]/P0001  ;
	input \u5_dout_reg[4]/P0001  ;
	input \u5_dout_reg[5]/P0001  ;
	input \u5_dout_reg[6]/P0001  ;
	input \u5_dout_reg[7]/P0001  ;
	input \u5_dout_reg[8]/P0001  ;
	input \u5_dout_reg[9]/P0001  ;
	input \u5_empty_reg/NET0131  ;
	input \u5_mem_reg[0][0]/NET0131  ;
	input \u5_mem_reg[0][10]/NET0131  ;
	input \u5_mem_reg[0][11]/NET0131  ;
	input \u5_mem_reg[0][12]/NET0131  ;
	input \u5_mem_reg[0][13]/NET0131  ;
	input \u5_mem_reg[0][14]/NET0131  ;
	input \u5_mem_reg[0][15]/NET0131  ;
	input \u5_mem_reg[0][16]/NET0131  ;
	input \u5_mem_reg[0][17]/NET0131  ;
	input \u5_mem_reg[0][18]/NET0131  ;
	input \u5_mem_reg[0][19]/NET0131  ;
	input \u5_mem_reg[0][1]/NET0131  ;
	input \u5_mem_reg[0][20]/NET0131  ;
	input \u5_mem_reg[0][21]/NET0131  ;
	input \u5_mem_reg[0][22]/NET0131  ;
	input \u5_mem_reg[0][23]/NET0131  ;
	input \u5_mem_reg[0][24]/NET0131  ;
	input \u5_mem_reg[0][25]/NET0131  ;
	input \u5_mem_reg[0][26]/NET0131  ;
	input \u5_mem_reg[0][27]/NET0131  ;
	input \u5_mem_reg[0][28]/NET0131  ;
	input \u5_mem_reg[0][29]/NET0131  ;
	input \u5_mem_reg[0][2]/NET0131  ;
	input \u5_mem_reg[0][30]/NET0131  ;
	input \u5_mem_reg[0][31]/NET0131  ;
	input \u5_mem_reg[0][3]/NET0131  ;
	input \u5_mem_reg[0][4]/NET0131  ;
	input \u5_mem_reg[0][5]/NET0131  ;
	input \u5_mem_reg[0][6]/NET0131  ;
	input \u5_mem_reg[0][7]/NET0131  ;
	input \u5_mem_reg[0][8]/NET0131  ;
	input \u5_mem_reg[0][9]/NET0131  ;
	input \u5_mem_reg[1][0]/NET0131  ;
	input \u5_mem_reg[1][10]/NET0131  ;
	input \u5_mem_reg[1][11]/NET0131  ;
	input \u5_mem_reg[1][12]/NET0131  ;
	input \u5_mem_reg[1][13]/NET0131  ;
	input \u5_mem_reg[1][14]/NET0131  ;
	input \u5_mem_reg[1][15]/NET0131  ;
	input \u5_mem_reg[1][16]/NET0131  ;
	input \u5_mem_reg[1][17]/NET0131  ;
	input \u5_mem_reg[1][18]/NET0131  ;
	input \u5_mem_reg[1][19]/NET0131  ;
	input \u5_mem_reg[1][1]/NET0131  ;
	input \u5_mem_reg[1][20]/NET0131  ;
	input \u5_mem_reg[1][21]/NET0131  ;
	input \u5_mem_reg[1][22]/NET0131  ;
	input \u5_mem_reg[1][23]/NET0131  ;
	input \u5_mem_reg[1][24]/NET0131  ;
	input \u5_mem_reg[1][25]/NET0131  ;
	input \u5_mem_reg[1][26]/NET0131  ;
	input \u5_mem_reg[1][27]/NET0131  ;
	input \u5_mem_reg[1][28]/NET0131  ;
	input \u5_mem_reg[1][29]/NET0131  ;
	input \u5_mem_reg[1][2]/NET0131  ;
	input \u5_mem_reg[1][30]/NET0131  ;
	input \u5_mem_reg[1][31]/NET0131  ;
	input \u5_mem_reg[1][3]/NET0131  ;
	input \u5_mem_reg[1][4]/NET0131  ;
	input \u5_mem_reg[1][5]/NET0131  ;
	input \u5_mem_reg[1][6]/NET0131  ;
	input \u5_mem_reg[1][7]/NET0131  ;
	input \u5_mem_reg[1][8]/NET0131  ;
	input \u5_mem_reg[1][9]/NET0131  ;
	input \u5_mem_reg[2][0]/NET0131  ;
	input \u5_mem_reg[2][10]/NET0131  ;
	input \u5_mem_reg[2][11]/NET0131  ;
	input \u5_mem_reg[2][12]/NET0131  ;
	input \u5_mem_reg[2][13]/NET0131  ;
	input \u5_mem_reg[2][14]/NET0131  ;
	input \u5_mem_reg[2][15]/NET0131  ;
	input \u5_mem_reg[2][16]/NET0131  ;
	input \u5_mem_reg[2][17]/NET0131  ;
	input \u5_mem_reg[2][18]/NET0131  ;
	input \u5_mem_reg[2][19]/NET0131  ;
	input \u5_mem_reg[2][1]/NET0131  ;
	input \u5_mem_reg[2][20]/NET0131  ;
	input \u5_mem_reg[2][21]/NET0131  ;
	input \u5_mem_reg[2][22]/NET0131  ;
	input \u5_mem_reg[2][23]/NET0131  ;
	input \u5_mem_reg[2][24]/NET0131  ;
	input \u5_mem_reg[2][25]/NET0131  ;
	input \u5_mem_reg[2][26]/NET0131  ;
	input \u5_mem_reg[2][27]/NET0131  ;
	input \u5_mem_reg[2][28]/NET0131  ;
	input \u5_mem_reg[2][29]/NET0131  ;
	input \u5_mem_reg[2][2]/NET0131  ;
	input \u5_mem_reg[2][30]/NET0131  ;
	input \u5_mem_reg[2][31]/NET0131  ;
	input \u5_mem_reg[2][3]/NET0131  ;
	input \u5_mem_reg[2][4]/NET0131  ;
	input \u5_mem_reg[2][5]/NET0131  ;
	input \u5_mem_reg[2][6]/NET0131  ;
	input \u5_mem_reg[2][7]/NET0131  ;
	input \u5_mem_reg[2][8]/NET0131  ;
	input \u5_mem_reg[2][9]/NET0131  ;
	input \u5_mem_reg[3][0]/NET0131  ;
	input \u5_mem_reg[3][10]/NET0131  ;
	input \u5_mem_reg[3][11]/NET0131  ;
	input \u5_mem_reg[3][12]/NET0131  ;
	input \u5_mem_reg[3][13]/NET0131  ;
	input \u5_mem_reg[3][14]/NET0131  ;
	input \u5_mem_reg[3][15]/NET0131  ;
	input \u5_mem_reg[3][16]/NET0131  ;
	input \u5_mem_reg[3][17]/NET0131  ;
	input \u5_mem_reg[3][18]/NET0131  ;
	input \u5_mem_reg[3][19]/NET0131  ;
	input \u5_mem_reg[3][1]/NET0131  ;
	input \u5_mem_reg[3][20]/NET0131  ;
	input \u5_mem_reg[3][21]/NET0131  ;
	input \u5_mem_reg[3][22]/NET0131  ;
	input \u5_mem_reg[3][23]/NET0131  ;
	input \u5_mem_reg[3][24]/NET0131  ;
	input \u5_mem_reg[3][25]/NET0131  ;
	input \u5_mem_reg[3][26]/NET0131  ;
	input \u5_mem_reg[3][27]/NET0131  ;
	input \u5_mem_reg[3][28]/NET0131  ;
	input \u5_mem_reg[3][29]/NET0131  ;
	input \u5_mem_reg[3][2]/NET0131  ;
	input \u5_mem_reg[3][30]/NET0131  ;
	input \u5_mem_reg[3][31]/NET0131  ;
	input \u5_mem_reg[3][3]/NET0131  ;
	input \u5_mem_reg[3][4]/NET0131  ;
	input \u5_mem_reg[3][5]/NET0131  ;
	input \u5_mem_reg[3][6]/NET0131  ;
	input \u5_mem_reg[3][7]/NET0131  ;
	input \u5_mem_reg[3][8]/NET0131  ;
	input \u5_mem_reg[3][9]/NET0131  ;
	input \u5_rp_reg[0]/P0001  ;
	input \u5_rp_reg[1]/NET0131  ;
	input \u5_rp_reg[2]/NET0131  ;
	input \u5_rp_reg[3]/NET0131  ;
	input \u5_status_reg[0]/P0001  ;
	input \u5_status_reg[1]/P0001  ;
	input \u5_wp_reg[0]/P0001  ;
	input \u5_wp_reg[1]/NET0131  ;
	input \u5_wp_reg[2]/P0001  ;
	input \u6_dout_reg[0]/P0001  ;
	input \u6_dout_reg[10]/P0001  ;
	input \u6_dout_reg[11]/P0001  ;
	input \u6_dout_reg[12]/P0001  ;
	input \u6_dout_reg[13]/P0001  ;
	input \u6_dout_reg[14]/P0001  ;
	input \u6_dout_reg[15]/P0001  ;
	input \u6_dout_reg[16]/P0001  ;
	input \u6_dout_reg[17]/P0001  ;
	input \u6_dout_reg[18]/P0001  ;
	input \u6_dout_reg[19]/P0001  ;
	input \u6_dout_reg[1]/P0001  ;
	input \u6_dout_reg[2]/P0001  ;
	input \u6_dout_reg[3]/P0001  ;
	input \u6_dout_reg[4]/P0001  ;
	input \u6_dout_reg[5]/P0001  ;
	input \u6_dout_reg[6]/P0001  ;
	input \u6_dout_reg[7]/P0001  ;
	input \u6_dout_reg[8]/P0001  ;
	input \u6_dout_reg[9]/P0001  ;
	input \u6_empty_reg/NET0131  ;
	input \u6_mem_reg[0][0]/NET0131  ;
	input \u6_mem_reg[0][10]/NET0131  ;
	input \u6_mem_reg[0][11]/NET0131  ;
	input \u6_mem_reg[0][12]/NET0131  ;
	input \u6_mem_reg[0][13]/NET0131  ;
	input \u6_mem_reg[0][14]/NET0131  ;
	input \u6_mem_reg[0][15]/NET0131  ;
	input \u6_mem_reg[0][16]/NET0131  ;
	input \u6_mem_reg[0][17]/NET0131  ;
	input \u6_mem_reg[0][18]/NET0131  ;
	input \u6_mem_reg[0][19]/NET0131  ;
	input \u6_mem_reg[0][1]/NET0131  ;
	input \u6_mem_reg[0][20]/NET0131  ;
	input \u6_mem_reg[0][21]/NET0131  ;
	input \u6_mem_reg[0][22]/NET0131  ;
	input \u6_mem_reg[0][23]/NET0131  ;
	input \u6_mem_reg[0][24]/NET0131  ;
	input \u6_mem_reg[0][25]/NET0131  ;
	input \u6_mem_reg[0][26]/NET0131  ;
	input \u6_mem_reg[0][27]/NET0131  ;
	input \u6_mem_reg[0][28]/NET0131  ;
	input \u6_mem_reg[0][29]/NET0131  ;
	input \u6_mem_reg[0][2]/NET0131  ;
	input \u6_mem_reg[0][30]/NET0131  ;
	input \u6_mem_reg[0][31]/NET0131  ;
	input \u6_mem_reg[0][3]/NET0131  ;
	input \u6_mem_reg[0][4]/NET0131  ;
	input \u6_mem_reg[0][5]/NET0131  ;
	input \u6_mem_reg[0][6]/NET0131  ;
	input \u6_mem_reg[0][7]/NET0131  ;
	input \u6_mem_reg[0][8]/NET0131  ;
	input \u6_mem_reg[0][9]/NET0131  ;
	input \u6_mem_reg[1][0]/NET0131  ;
	input \u6_mem_reg[1][10]/NET0131  ;
	input \u6_mem_reg[1][11]/NET0131  ;
	input \u6_mem_reg[1][12]/NET0131  ;
	input \u6_mem_reg[1][13]/NET0131  ;
	input \u6_mem_reg[1][14]/NET0131  ;
	input \u6_mem_reg[1][15]/NET0131  ;
	input \u6_mem_reg[1][16]/NET0131  ;
	input \u6_mem_reg[1][17]/NET0131  ;
	input \u6_mem_reg[1][18]/NET0131  ;
	input \u6_mem_reg[1][19]/NET0131  ;
	input \u6_mem_reg[1][1]/NET0131  ;
	input \u6_mem_reg[1][20]/NET0131  ;
	input \u6_mem_reg[1][21]/NET0131  ;
	input \u6_mem_reg[1][22]/NET0131  ;
	input \u6_mem_reg[1][23]/NET0131  ;
	input \u6_mem_reg[1][24]/NET0131  ;
	input \u6_mem_reg[1][25]/NET0131  ;
	input \u6_mem_reg[1][26]/NET0131  ;
	input \u6_mem_reg[1][27]/NET0131  ;
	input \u6_mem_reg[1][28]/NET0131  ;
	input \u6_mem_reg[1][29]/NET0131  ;
	input \u6_mem_reg[1][2]/NET0131  ;
	input \u6_mem_reg[1][30]/NET0131  ;
	input \u6_mem_reg[1][31]/NET0131  ;
	input \u6_mem_reg[1][3]/NET0131  ;
	input \u6_mem_reg[1][4]/NET0131  ;
	input \u6_mem_reg[1][5]/NET0131  ;
	input \u6_mem_reg[1][6]/NET0131  ;
	input \u6_mem_reg[1][7]/NET0131  ;
	input \u6_mem_reg[1][8]/NET0131  ;
	input \u6_mem_reg[1][9]/NET0131  ;
	input \u6_mem_reg[2][0]/NET0131  ;
	input \u6_mem_reg[2][10]/NET0131  ;
	input \u6_mem_reg[2][11]/NET0131  ;
	input \u6_mem_reg[2][12]/NET0131  ;
	input \u6_mem_reg[2][13]/NET0131  ;
	input \u6_mem_reg[2][14]/NET0131  ;
	input \u6_mem_reg[2][15]/NET0131  ;
	input \u6_mem_reg[2][16]/NET0131  ;
	input \u6_mem_reg[2][17]/NET0131  ;
	input \u6_mem_reg[2][18]/NET0131  ;
	input \u6_mem_reg[2][19]/NET0131  ;
	input \u6_mem_reg[2][1]/NET0131  ;
	input \u6_mem_reg[2][20]/NET0131  ;
	input \u6_mem_reg[2][21]/NET0131  ;
	input \u6_mem_reg[2][22]/NET0131  ;
	input \u6_mem_reg[2][23]/NET0131  ;
	input \u6_mem_reg[2][24]/NET0131  ;
	input \u6_mem_reg[2][25]/NET0131  ;
	input \u6_mem_reg[2][26]/NET0131  ;
	input \u6_mem_reg[2][27]/NET0131  ;
	input \u6_mem_reg[2][28]/NET0131  ;
	input \u6_mem_reg[2][29]/NET0131  ;
	input \u6_mem_reg[2][2]/NET0131  ;
	input \u6_mem_reg[2][30]/NET0131  ;
	input \u6_mem_reg[2][31]/NET0131  ;
	input \u6_mem_reg[2][3]/NET0131  ;
	input \u6_mem_reg[2][4]/NET0131  ;
	input \u6_mem_reg[2][5]/NET0131  ;
	input \u6_mem_reg[2][6]/NET0131  ;
	input \u6_mem_reg[2][7]/NET0131  ;
	input \u6_mem_reg[2][8]/NET0131  ;
	input \u6_mem_reg[2][9]/NET0131  ;
	input \u6_mem_reg[3][0]/NET0131  ;
	input \u6_mem_reg[3][10]/NET0131  ;
	input \u6_mem_reg[3][11]/NET0131  ;
	input \u6_mem_reg[3][12]/NET0131  ;
	input \u6_mem_reg[3][13]/NET0131  ;
	input \u6_mem_reg[3][14]/NET0131  ;
	input \u6_mem_reg[3][15]/NET0131  ;
	input \u6_mem_reg[3][16]/NET0131  ;
	input \u6_mem_reg[3][17]/NET0131  ;
	input \u6_mem_reg[3][18]/NET0131  ;
	input \u6_mem_reg[3][19]/NET0131  ;
	input \u6_mem_reg[3][1]/NET0131  ;
	input \u6_mem_reg[3][20]/NET0131  ;
	input \u6_mem_reg[3][21]/NET0131  ;
	input \u6_mem_reg[3][22]/NET0131  ;
	input \u6_mem_reg[3][23]/NET0131  ;
	input \u6_mem_reg[3][24]/NET0131  ;
	input \u6_mem_reg[3][25]/NET0131  ;
	input \u6_mem_reg[3][26]/NET0131  ;
	input \u6_mem_reg[3][27]/NET0131  ;
	input \u6_mem_reg[3][28]/NET0131  ;
	input \u6_mem_reg[3][29]/NET0131  ;
	input \u6_mem_reg[3][2]/NET0131  ;
	input \u6_mem_reg[3][30]/NET0131  ;
	input \u6_mem_reg[3][31]/NET0131  ;
	input \u6_mem_reg[3][3]/NET0131  ;
	input \u6_mem_reg[3][4]/NET0131  ;
	input \u6_mem_reg[3][5]/NET0131  ;
	input \u6_mem_reg[3][6]/NET0131  ;
	input \u6_mem_reg[3][7]/NET0131  ;
	input \u6_mem_reg[3][8]/NET0131  ;
	input \u6_mem_reg[3][9]/NET0131  ;
	input \u6_rp_reg[0]/P0001  ;
	input \u6_rp_reg[1]/NET0131  ;
	input \u6_rp_reg[2]/NET0131  ;
	input \u6_rp_reg[3]/NET0131  ;
	input \u6_status_reg[0]/P0001  ;
	input \u6_status_reg[1]/P0001  ;
	input \u6_wp_reg[0]/P0001  ;
	input \u6_wp_reg[1]/NET0131  ;
	input \u6_wp_reg[2]/P0001  ;
	input \u7_dout_reg[0]/P0001  ;
	input \u7_dout_reg[10]/P0001  ;
	input \u7_dout_reg[11]/P0001  ;
	input \u7_dout_reg[12]/P0001  ;
	input \u7_dout_reg[13]/P0001  ;
	input \u7_dout_reg[14]/P0001  ;
	input \u7_dout_reg[15]/P0001  ;
	input \u7_dout_reg[16]/P0001  ;
	input \u7_dout_reg[17]/P0001  ;
	input \u7_dout_reg[18]/P0001  ;
	input \u7_dout_reg[19]/P0001  ;
	input \u7_dout_reg[1]/P0001  ;
	input \u7_dout_reg[2]/P0001  ;
	input \u7_dout_reg[3]/P0001  ;
	input \u7_dout_reg[4]/P0001  ;
	input \u7_dout_reg[5]/P0001  ;
	input \u7_dout_reg[6]/P0001  ;
	input \u7_dout_reg[7]/P0001  ;
	input \u7_dout_reg[8]/P0001  ;
	input \u7_dout_reg[9]/P0001  ;
	input \u7_empty_reg/NET0131  ;
	input \u7_mem_reg[0][0]/NET0131  ;
	input \u7_mem_reg[0][10]/NET0131  ;
	input \u7_mem_reg[0][11]/NET0131  ;
	input \u7_mem_reg[0][12]/NET0131  ;
	input \u7_mem_reg[0][13]/NET0131  ;
	input \u7_mem_reg[0][14]/NET0131  ;
	input \u7_mem_reg[0][15]/NET0131  ;
	input \u7_mem_reg[0][16]/NET0131  ;
	input \u7_mem_reg[0][17]/NET0131  ;
	input \u7_mem_reg[0][18]/NET0131  ;
	input \u7_mem_reg[0][19]/NET0131  ;
	input \u7_mem_reg[0][1]/NET0131  ;
	input \u7_mem_reg[0][20]/NET0131  ;
	input \u7_mem_reg[0][21]/NET0131  ;
	input \u7_mem_reg[0][22]/NET0131  ;
	input \u7_mem_reg[0][23]/NET0131  ;
	input \u7_mem_reg[0][24]/NET0131  ;
	input \u7_mem_reg[0][25]/NET0131  ;
	input \u7_mem_reg[0][26]/NET0131  ;
	input \u7_mem_reg[0][27]/NET0131  ;
	input \u7_mem_reg[0][28]/NET0131  ;
	input \u7_mem_reg[0][29]/NET0131  ;
	input \u7_mem_reg[0][2]/NET0131  ;
	input \u7_mem_reg[0][30]/NET0131  ;
	input \u7_mem_reg[0][31]/NET0131  ;
	input \u7_mem_reg[0][3]/NET0131  ;
	input \u7_mem_reg[0][4]/NET0131  ;
	input \u7_mem_reg[0][5]/NET0131  ;
	input \u7_mem_reg[0][6]/NET0131  ;
	input \u7_mem_reg[0][7]/NET0131  ;
	input \u7_mem_reg[0][8]/NET0131  ;
	input \u7_mem_reg[0][9]/NET0131  ;
	input \u7_mem_reg[1][0]/NET0131  ;
	input \u7_mem_reg[1][10]/NET0131  ;
	input \u7_mem_reg[1][11]/NET0131  ;
	input \u7_mem_reg[1][12]/NET0131  ;
	input \u7_mem_reg[1][13]/NET0131  ;
	input \u7_mem_reg[1][14]/NET0131  ;
	input \u7_mem_reg[1][15]/NET0131  ;
	input \u7_mem_reg[1][16]/NET0131  ;
	input \u7_mem_reg[1][17]/NET0131  ;
	input \u7_mem_reg[1][18]/NET0131  ;
	input \u7_mem_reg[1][19]/NET0131  ;
	input \u7_mem_reg[1][1]/NET0131  ;
	input \u7_mem_reg[1][20]/NET0131  ;
	input \u7_mem_reg[1][21]/NET0131  ;
	input \u7_mem_reg[1][22]/NET0131  ;
	input \u7_mem_reg[1][23]/NET0131  ;
	input \u7_mem_reg[1][24]/NET0131  ;
	input \u7_mem_reg[1][25]/NET0131  ;
	input \u7_mem_reg[1][26]/NET0131  ;
	input \u7_mem_reg[1][27]/NET0131  ;
	input \u7_mem_reg[1][28]/NET0131  ;
	input \u7_mem_reg[1][29]/NET0131  ;
	input \u7_mem_reg[1][2]/NET0131  ;
	input \u7_mem_reg[1][30]/NET0131  ;
	input \u7_mem_reg[1][31]/NET0131  ;
	input \u7_mem_reg[1][3]/NET0131  ;
	input \u7_mem_reg[1][4]/NET0131  ;
	input \u7_mem_reg[1][5]/NET0131  ;
	input \u7_mem_reg[1][6]/NET0131  ;
	input \u7_mem_reg[1][7]/NET0131  ;
	input \u7_mem_reg[1][8]/NET0131  ;
	input \u7_mem_reg[1][9]/NET0131  ;
	input \u7_mem_reg[2][0]/NET0131  ;
	input \u7_mem_reg[2][10]/NET0131  ;
	input \u7_mem_reg[2][11]/NET0131  ;
	input \u7_mem_reg[2][12]/NET0131  ;
	input \u7_mem_reg[2][13]/NET0131  ;
	input \u7_mem_reg[2][14]/NET0131  ;
	input \u7_mem_reg[2][15]/NET0131  ;
	input \u7_mem_reg[2][16]/NET0131  ;
	input \u7_mem_reg[2][17]/NET0131  ;
	input \u7_mem_reg[2][18]/NET0131  ;
	input \u7_mem_reg[2][19]/NET0131  ;
	input \u7_mem_reg[2][1]/NET0131  ;
	input \u7_mem_reg[2][20]/NET0131  ;
	input \u7_mem_reg[2][21]/NET0131  ;
	input \u7_mem_reg[2][22]/NET0131  ;
	input \u7_mem_reg[2][23]/NET0131  ;
	input \u7_mem_reg[2][24]/NET0131  ;
	input \u7_mem_reg[2][25]/NET0131  ;
	input \u7_mem_reg[2][26]/NET0131  ;
	input \u7_mem_reg[2][27]/NET0131  ;
	input \u7_mem_reg[2][28]/NET0131  ;
	input \u7_mem_reg[2][29]/NET0131  ;
	input \u7_mem_reg[2][2]/NET0131  ;
	input \u7_mem_reg[2][30]/NET0131  ;
	input \u7_mem_reg[2][31]/NET0131  ;
	input \u7_mem_reg[2][3]/NET0131  ;
	input \u7_mem_reg[2][4]/NET0131  ;
	input \u7_mem_reg[2][5]/NET0131  ;
	input \u7_mem_reg[2][6]/NET0131  ;
	input \u7_mem_reg[2][7]/NET0131  ;
	input \u7_mem_reg[2][8]/NET0131  ;
	input \u7_mem_reg[2][9]/NET0131  ;
	input \u7_mem_reg[3][0]/NET0131  ;
	input \u7_mem_reg[3][10]/NET0131  ;
	input \u7_mem_reg[3][11]/NET0131  ;
	input \u7_mem_reg[3][12]/NET0131  ;
	input \u7_mem_reg[3][13]/NET0131  ;
	input \u7_mem_reg[3][14]/NET0131  ;
	input \u7_mem_reg[3][15]/NET0131  ;
	input \u7_mem_reg[3][16]/NET0131  ;
	input \u7_mem_reg[3][17]/NET0131  ;
	input \u7_mem_reg[3][18]/NET0131  ;
	input \u7_mem_reg[3][19]/NET0131  ;
	input \u7_mem_reg[3][1]/NET0131  ;
	input \u7_mem_reg[3][20]/NET0131  ;
	input \u7_mem_reg[3][21]/NET0131  ;
	input \u7_mem_reg[3][22]/NET0131  ;
	input \u7_mem_reg[3][23]/NET0131  ;
	input \u7_mem_reg[3][24]/NET0131  ;
	input \u7_mem_reg[3][25]/NET0131  ;
	input \u7_mem_reg[3][26]/NET0131  ;
	input \u7_mem_reg[3][27]/NET0131  ;
	input \u7_mem_reg[3][28]/NET0131  ;
	input \u7_mem_reg[3][29]/NET0131  ;
	input \u7_mem_reg[3][2]/NET0131  ;
	input \u7_mem_reg[3][30]/NET0131  ;
	input \u7_mem_reg[3][31]/NET0131  ;
	input \u7_mem_reg[3][3]/NET0131  ;
	input \u7_mem_reg[3][4]/NET0131  ;
	input \u7_mem_reg[3][5]/NET0131  ;
	input \u7_mem_reg[3][6]/NET0131  ;
	input \u7_mem_reg[3][7]/NET0131  ;
	input \u7_mem_reg[3][8]/NET0131  ;
	input \u7_mem_reg[3][9]/NET0131  ;
	input \u7_rp_reg[0]/P0001  ;
	input \u7_rp_reg[1]/NET0131  ;
	input \u7_rp_reg[2]/NET0131  ;
	input \u7_rp_reg[3]/NET0131  ;
	input \u7_status_reg[0]/P0001  ;
	input \u7_status_reg[1]/P0001  ;
	input \u7_wp_reg[0]/P0001  ;
	input \u7_wp_reg[1]/NET0131  ;
	input \u7_wp_reg[2]/P0001  ;
	input \u8_dout_reg[0]/P0001  ;
	input \u8_dout_reg[10]/P0001  ;
	input \u8_dout_reg[11]/P0001  ;
	input \u8_dout_reg[12]/P0001  ;
	input \u8_dout_reg[13]/P0001  ;
	input \u8_dout_reg[14]/P0001  ;
	input \u8_dout_reg[15]/P0001  ;
	input \u8_dout_reg[16]/P0001  ;
	input \u8_dout_reg[17]/P0001  ;
	input \u8_dout_reg[18]/P0001  ;
	input \u8_dout_reg[19]/P0001  ;
	input \u8_dout_reg[1]/P0001  ;
	input \u8_dout_reg[2]/P0001  ;
	input \u8_dout_reg[3]/P0001  ;
	input \u8_dout_reg[4]/P0001  ;
	input \u8_dout_reg[5]/P0001  ;
	input \u8_dout_reg[6]/P0001  ;
	input \u8_dout_reg[7]/P0001  ;
	input \u8_dout_reg[8]/P0001  ;
	input \u8_dout_reg[9]/P0001  ;
	input \u8_empty_reg/NET0131  ;
	input \u8_mem_reg[0][0]/NET0131  ;
	input \u8_mem_reg[0][10]/NET0131  ;
	input \u8_mem_reg[0][11]/NET0131  ;
	input \u8_mem_reg[0][12]/NET0131  ;
	input \u8_mem_reg[0][13]/NET0131  ;
	input \u8_mem_reg[0][14]/NET0131  ;
	input \u8_mem_reg[0][15]/NET0131  ;
	input \u8_mem_reg[0][16]/NET0131  ;
	input \u8_mem_reg[0][17]/NET0131  ;
	input \u8_mem_reg[0][18]/NET0131  ;
	input \u8_mem_reg[0][19]/NET0131  ;
	input \u8_mem_reg[0][1]/NET0131  ;
	input \u8_mem_reg[0][20]/NET0131  ;
	input \u8_mem_reg[0][21]/NET0131  ;
	input \u8_mem_reg[0][22]/NET0131  ;
	input \u8_mem_reg[0][23]/NET0131  ;
	input \u8_mem_reg[0][24]/NET0131  ;
	input \u8_mem_reg[0][25]/NET0131  ;
	input \u8_mem_reg[0][26]/NET0131  ;
	input \u8_mem_reg[0][27]/NET0131  ;
	input \u8_mem_reg[0][28]/NET0131  ;
	input \u8_mem_reg[0][29]/NET0131  ;
	input \u8_mem_reg[0][2]/NET0131  ;
	input \u8_mem_reg[0][30]/NET0131  ;
	input \u8_mem_reg[0][31]/NET0131  ;
	input \u8_mem_reg[0][3]/NET0131  ;
	input \u8_mem_reg[0][4]/NET0131  ;
	input \u8_mem_reg[0][5]/NET0131  ;
	input \u8_mem_reg[0][6]/NET0131  ;
	input \u8_mem_reg[0][7]/NET0131  ;
	input \u8_mem_reg[0][8]/NET0131  ;
	input \u8_mem_reg[0][9]/NET0131  ;
	input \u8_mem_reg[1][0]/NET0131  ;
	input \u8_mem_reg[1][10]/NET0131  ;
	input \u8_mem_reg[1][11]/NET0131  ;
	input \u8_mem_reg[1][12]/NET0131  ;
	input \u8_mem_reg[1][13]/NET0131  ;
	input \u8_mem_reg[1][14]/NET0131  ;
	input \u8_mem_reg[1][15]/NET0131  ;
	input \u8_mem_reg[1][16]/NET0131  ;
	input \u8_mem_reg[1][17]/NET0131  ;
	input \u8_mem_reg[1][18]/NET0131  ;
	input \u8_mem_reg[1][19]/NET0131  ;
	input \u8_mem_reg[1][1]/NET0131  ;
	input \u8_mem_reg[1][20]/NET0131  ;
	input \u8_mem_reg[1][21]/NET0131  ;
	input \u8_mem_reg[1][22]/NET0131  ;
	input \u8_mem_reg[1][23]/NET0131  ;
	input \u8_mem_reg[1][24]/NET0131  ;
	input \u8_mem_reg[1][25]/NET0131  ;
	input \u8_mem_reg[1][26]/NET0131  ;
	input \u8_mem_reg[1][27]/NET0131  ;
	input \u8_mem_reg[1][28]/NET0131  ;
	input \u8_mem_reg[1][29]/NET0131  ;
	input \u8_mem_reg[1][2]/NET0131  ;
	input \u8_mem_reg[1][30]/NET0131  ;
	input \u8_mem_reg[1][31]/NET0131  ;
	input \u8_mem_reg[1][3]/NET0131  ;
	input \u8_mem_reg[1][4]/NET0131  ;
	input \u8_mem_reg[1][5]/NET0131  ;
	input \u8_mem_reg[1][6]/NET0131  ;
	input \u8_mem_reg[1][7]/NET0131  ;
	input \u8_mem_reg[1][8]/NET0131  ;
	input \u8_mem_reg[1][9]/NET0131  ;
	input \u8_mem_reg[2][0]/NET0131  ;
	input \u8_mem_reg[2][10]/NET0131  ;
	input \u8_mem_reg[2][11]/NET0131  ;
	input \u8_mem_reg[2][12]/NET0131  ;
	input \u8_mem_reg[2][13]/NET0131  ;
	input \u8_mem_reg[2][14]/NET0131  ;
	input \u8_mem_reg[2][15]/NET0131  ;
	input \u8_mem_reg[2][16]/NET0131  ;
	input \u8_mem_reg[2][17]/NET0131  ;
	input \u8_mem_reg[2][18]/NET0131  ;
	input \u8_mem_reg[2][19]/NET0131  ;
	input \u8_mem_reg[2][1]/NET0131  ;
	input \u8_mem_reg[2][20]/NET0131  ;
	input \u8_mem_reg[2][21]/NET0131  ;
	input \u8_mem_reg[2][22]/NET0131  ;
	input \u8_mem_reg[2][23]/NET0131  ;
	input \u8_mem_reg[2][24]/NET0131  ;
	input \u8_mem_reg[2][25]/NET0131  ;
	input \u8_mem_reg[2][26]/NET0131  ;
	input \u8_mem_reg[2][27]/NET0131  ;
	input \u8_mem_reg[2][28]/NET0131  ;
	input \u8_mem_reg[2][29]/NET0131  ;
	input \u8_mem_reg[2][2]/NET0131  ;
	input \u8_mem_reg[2][30]/NET0131  ;
	input \u8_mem_reg[2][31]/NET0131  ;
	input \u8_mem_reg[2][3]/NET0131  ;
	input \u8_mem_reg[2][4]/NET0131  ;
	input \u8_mem_reg[2][5]/NET0131  ;
	input \u8_mem_reg[2][6]/NET0131  ;
	input \u8_mem_reg[2][7]/NET0131  ;
	input \u8_mem_reg[2][8]/NET0131  ;
	input \u8_mem_reg[2][9]/NET0131  ;
	input \u8_mem_reg[3][0]/NET0131  ;
	input \u8_mem_reg[3][10]/NET0131  ;
	input \u8_mem_reg[3][11]/NET0131  ;
	input \u8_mem_reg[3][12]/NET0131  ;
	input \u8_mem_reg[3][13]/NET0131  ;
	input \u8_mem_reg[3][14]/NET0131  ;
	input \u8_mem_reg[3][15]/NET0131  ;
	input \u8_mem_reg[3][16]/NET0131  ;
	input \u8_mem_reg[3][17]/NET0131  ;
	input \u8_mem_reg[3][18]/NET0131  ;
	input \u8_mem_reg[3][19]/NET0131  ;
	input \u8_mem_reg[3][1]/NET0131  ;
	input \u8_mem_reg[3][20]/NET0131  ;
	input \u8_mem_reg[3][21]/NET0131  ;
	input \u8_mem_reg[3][22]/NET0131  ;
	input \u8_mem_reg[3][23]/NET0131  ;
	input \u8_mem_reg[3][24]/NET0131  ;
	input \u8_mem_reg[3][25]/NET0131  ;
	input \u8_mem_reg[3][26]/NET0131  ;
	input \u8_mem_reg[3][27]/NET0131  ;
	input \u8_mem_reg[3][28]/NET0131  ;
	input \u8_mem_reg[3][29]/NET0131  ;
	input \u8_mem_reg[3][2]/NET0131  ;
	input \u8_mem_reg[3][30]/NET0131  ;
	input \u8_mem_reg[3][31]/NET0131  ;
	input \u8_mem_reg[3][3]/NET0131  ;
	input \u8_mem_reg[3][4]/NET0131  ;
	input \u8_mem_reg[3][5]/NET0131  ;
	input \u8_mem_reg[3][6]/NET0131  ;
	input \u8_mem_reg[3][7]/NET0131  ;
	input \u8_mem_reg[3][8]/NET0131  ;
	input \u8_mem_reg[3][9]/NET0131  ;
	input \u8_rp_reg[0]/P0001  ;
	input \u8_rp_reg[1]/NET0131  ;
	input \u8_rp_reg[2]/NET0131  ;
	input \u8_rp_reg[3]/NET0131  ;
	input \u8_status_reg[0]/P0001  ;
	input \u8_status_reg[1]/P0001  ;
	input \u8_wp_reg[0]/P0001  ;
	input \u8_wp_reg[1]/NET0131  ;
	input \u8_wp_reg[2]/P0001  ;
	input \u9_din_tmp1_reg[0]/P0001  ;
	input \u9_din_tmp1_reg[10]/P0001  ;
	input \u9_din_tmp1_reg[11]/P0001  ;
	input \u9_din_tmp1_reg[12]/P0001  ;
	input \u9_din_tmp1_reg[13]/P0001  ;
	input \u9_din_tmp1_reg[14]/P0001  ;
	input \u9_din_tmp1_reg[15]/P0001  ;
	input \u9_din_tmp1_reg[1]/P0001  ;
	input \u9_din_tmp1_reg[2]/P0001  ;
	input \u9_din_tmp1_reg[3]/P0001  ;
	input \u9_din_tmp1_reg[4]/P0001  ;
	input \u9_din_tmp1_reg[5]/P0001  ;
	input \u9_din_tmp1_reg[6]/P0001  ;
	input \u9_din_tmp1_reg[7]/P0001  ;
	input \u9_din_tmp1_reg[8]/P0001  ;
	input \u9_din_tmp1_reg[9]/P0001  ;
	input \u9_dout_reg[0]/P0001  ;
	input \u9_dout_reg[10]/P0001  ;
	input \u9_dout_reg[11]/P0001  ;
	input \u9_dout_reg[12]/P0001  ;
	input \u9_dout_reg[13]/P0001  ;
	input \u9_dout_reg[14]/P0001  ;
	input \u9_dout_reg[15]/P0001  ;
	input \u9_dout_reg[16]/P0001  ;
	input \u9_dout_reg[17]/P0001  ;
	input \u9_dout_reg[18]/P0001  ;
	input \u9_dout_reg[19]/P0001  ;
	input \u9_dout_reg[1]/P0001  ;
	input \u9_dout_reg[20]/P0001  ;
	input \u9_dout_reg[21]/P0001  ;
	input \u9_dout_reg[22]/P0001  ;
	input \u9_dout_reg[23]/P0001  ;
	input \u9_dout_reg[24]/P0001  ;
	input \u9_dout_reg[25]/P0001  ;
	input \u9_dout_reg[26]/P0001  ;
	input \u9_dout_reg[27]/P0001  ;
	input \u9_dout_reg[28]/P0001  ;
	input \u9_dout_reg[29]/P0001  ;
	input \u9_dout_reg[2]/P0001  ;
	input \u9_dout_reg[30]/P0001  ;
	input \u9_dout_reg[31]/P0001  ;
	input \u9_dout_reg[3]/P0001  ;
	input \u9_dout_reg[4]/P0001  ;
	input \u9_dout_reg[5]/P0001  ;
	input \u9_dout_reg[6]/P0001  ;
	input \u9_dout_reg[7]/P0001  ;
	input \u9_dout_reg[8]/P0001  ;
	input \u9_dout_reg[9]/P0001  ;
	input \u9_empty_reg/P0001  ;
	input \u9_full_reg/NET0131  ;
	input \u9_mem_reg[0][0]/P0001  ;
	input \u9_mem_reg[0][10]/P0001  ;
	input \u9_mem_reg[0][11]/P0001  ;
	input \u9_mem_reg[0][12]/P0001  ;
	input \u9_mem_reg[0][13]/P0001  ;
	input \u9_mem_reg[0][14]/P0001  ;
	input \u9_mem_reg[0][15]/P0001  ;
	input \u9_mem_reg[0][16]/P0001  ;
	input \u9_mem_reg[0][17]/P0001  ;
	input \u9_mem_reg[0][18]/P0001  ;
	input \u9_mem_reg[0][19]/P0001  ;
	input \u9_mem_reg[0][1]/P0001  ;
	input \u9_mem_reg[0][20]/P0001  ;
	input \u9_mem_reg[0][21]/P0001  ;
	input \u9_mem_reg[0][22]/P0001  ;
	input \u9_mem_reg[0][23]/P0001  ;
	input \u9_mem_reg[0][24]/P0001  ;
	input \u9_mem_reg[0][25]/P0001  ;
	input \u9_mem_reg[0][26]/P0001  ;
	input \u9_mem_reg[0][27]/P0001  ;
	input \u9_mem_reg[0][28]/P0001  ;
	input \u9_mem_reg[0][29]/P0001  ;
	input \u9_mem_reg[0][2]/P0001  ;
	input \u9_mem_reg[0][30]/P0001  ;
	input \u9_mem_reg[0][31]/P0001  ;
	input \u9_mem_reg[0][3]/P0001  ;
	input \u9_mem_reg[0][4]/P0001  ;
	input \u9_mem_reg[0][5]/P0001  ;
	input \u9_mem_reg[0][6]/P0001  ;
	input \u9_mem_reg[0][7]/P0001  ;
	input \u9_mem_reg[0][8]/P0001  ;
	input \u9_mem_reg[0][9]/P0001  ;
	input \u9_mem_reg[1][0]/P0001  ;
	input \u9_mem_reg[1][10]/P0001  ;
	input \u9_mem_reg[1][11]/P0001  ;
	input \u9_mem_reg[1][12]/P0001  ;
	input \u9_mem_reg[1][13]/P0001  ;
	input \u9_mem_reg[1][14]/P0001  ;
	input \u9_mem_reg[1][15]/P0001  ;
	input \u9_mem_reg[1][16]/P0001  ;
	input \u9_mem_reg[1][17]/P0001  ;
	input \u9_mem_reg[1][18]/P0001  ;
	input \u9_mem_reg[1][19]/P0001  ;
	input \u9_mem_reg[1][1]/P0001  ;
	input \u9_mem_reg[1][20]/P0001  ;
	input \u9_mem_reg[1][21]/P0001  ;
	input \u9_mem_reg[1][22]/P0001  ;
	input \u9_mem_reg[1][23]/P0001  ;
	input \u9_mem_reg[1][24]/P0001  ;
	input \u9_mem_reg[1][25]/P0001  ;
	input \u9_mem_reg[1][26]/P0001  ;
	input \u9_mem_reg[1][27]/P0001  ;
	input \u9_mem_reg[1][28]/P0001  ;
	input \u9_mem_reg[1][29]/P0001  ;
	input \u9_mem_reg[1][2]/P0001  ;
	input \u9_mem_reg[1][30]/P0001  ;
	input \u9_mem_reg[1][31]/P0001  ;
	input \u9_mem_reg[1][3]/P0001  ;
	input \u9_mem_reg[1][4]/P0001  ;
	input \u9_mem_reg[1][5]/P0001  ;
	input \u9_mem_reg[1][6]/P0001  ;
	input \u9_mem_reg[1][7]/P0001  ;
	input \u9_mem_reg[1][8]/P0001  ;
	input \u9_mem_reg[1][9]/P0001  ;
	input \u9_mem_reg[2][0]/P0001  ;
	input \u9_mem_reg[2][10]/P0001  ;
	input \u9_mem_reg[2][11]/P0001  ;
	input \u9_mem_reg[2][12]/P0001  ;
	input \u9_mem_reg[2][13]/P0001  ;
	input \u9_mem_reg[2][14]/P0001  ;
	input \u9_mem_reg[2][15]/P0001  ;
	input \u9_mem_reg[2][16]/P0001  ;
	input \u9_mem_reg[2][17]/P0001  ;
	input \u9_mem_reg[2][18]/P0001  ;
	input \u9_mem_reg[2][19]/P0001  ;
	input \u9_mem_reg[2][1]/P0001  ;
	input \u9_mem_reg[2][20]/P0001  ;
	input \u9_mem_reg[2][21]/P0001  ;
	input \u9_mem_reg[2][22]/P0001  ;
	input \u9_mem_reg[2][23]/P0001  ;
	input \u9_mem_reg[2][24]/P0001  ;
	input \u9_mem_reg[2][25]/P0001  ;
	input \u9_mem_reg[2][26]/P0001  ;
	input \u9_mem_reg[2][27]/P0001  ;
	input \u9_mem_reg[2][28]/P0001  ;
	input \u9_mem_reg[2][29]/P0001  ;
	input \u9_mem_reg[2][2]/P0001  ;
	input \u9_mem_reg[2][30]/P0001  ;
	input \u9_mem_reg[2][31]/P0001  ;
	input \u9_mem_reg[2][3]/P0001  ;
	input \u9_mem_reg[2][4]/P0001  ;
	input \u9_mem_reg[2][5]/P0001  ;
	input \u9_mem_reg[2][6]/P0001  ;
	input \u9_mem_reg[2][7]/P0001  ;
	input \u9_mem_reg[2][8]/P0001  ;
	input \u9_mem_reg[2][9]/P0001  ;
	input \u9_mem_reg[3][0]/P0001  ;
	input \u9_mem_reg[3][10]/P0001  ;
	input \u9_mem_reg[3][11]/P0001  ;
	input \u9_mem_reg[3][12]/P0001  ;
	input \u9_mem_reg[3][13]/P0001  ;
	input \u9_mem_reg[3][14]/P0001  ;
	input \u9_mem_reg[3][15]/P0001  ;
	input \u9_mem_reg[3][16]/P0001  ;
	input \u9_mem_reg[3][17]/P0001  ;
	input \u9_mem_reg[3][18]/P0001  ;
	input \u9_mem_reg[3][19]/P0001  ;
	input \u9_mem_reg[3][1]/P0001  ;
	input \u9_mem_reg[3][20]/P0001  ;
	input \u9_mem_reg[3][21]/P0001  ;
	input \u9_mem_reg[3][22]/P0001  ;
	input \u9_mem_reg[3][23]/P0001  ;
	input \u9_mem_reg[3][24]/P0001  ;
	input \u9_mem_reg[3][25]/P0001  ;
	input \u9_mem_reg[3][26]/P0001  ;
	input \u9_mem_reg[3][27]/P0001  ;
	input \u9_mem_reg[3][28]/P0001  ;
	input \u9_mem_reg[3][29]/P0001  ;
	input \u9_mem_reg[3][2]/P0001  ;
	input \u9_mem_reg[3][30]/P0001  ;
	input \u9_mem_reg[3][31]/P0001  ;
	input \u9_mem_reg[3][3]/P0001  ;
	input \u9_mem_reg[3][4]/P0001  ;
	input \u9_mem_reg[3][5]/P0001  ;
	input \u9_mem_reg[3][6]/P0001  ;
	input \u9_mem_reg[3][7]/P0001  ;
	input \u9_mem_reg[3][8]/P0001  ;
	input \u9_mem_reg[3][9]/P0001  ;
	input \u9_rp_reg[0]/P0001  ;
	input \u9_rp_reg[1]/P0001  ;
	input \u9_rp_reg[2]/P0001  ;
	input \u9_status_reg[0]/P0001  ;
	input \u9_status_reg[1]/P0001  ;
	input \u9_wp_reg[0]/NET0131  ;
	input \u9_wp_reg[1]/P0001  ;
	input \u9_wp_reg[2]/P0001  ;
	input \u9_wp_reg[3]/P0001  ;
	input \valid_s_reg/NET0131  ;
	input wb_ack_o_pad ;
	input \wb_addr_i[29]_pad  ;
	input \wb_addr_i[2]_pad  ;
	input \wb_addr_i[30]_pad  ;
	input \wb_addr_i[31]_pad  ;
	input \wb_addr_i[3]_pad  ;
	input \wb_addr_i[4]_pad  ;
	input \wb_addr_i[5]_pad  ;
	input \wb_addr_i[6]_pad  ;
	input wb_cyc_i_pad ;
	input wb_stb_i_pad ;
	input wb_we_i_pad ;
	output \_al_n1  ;
	output \g16/_0_  ;
	output \g23/_0_  ;
	output \g29500/_0_  ;
	output \g29503/_3_  ;
	output \g29505/_3_  ;
	output \g29507/_3_  ;
	output \g29509/_3_  ;
	output \g29511/_0_  ;
	output \g29513/_3_  ;
	output \g29515/_3_  ;
	output \g29517/_3_  ;
	output \g29519/_0_  ;
	output \g29522/_0_  ;
	output \g29524/_0_  ;
	output \g29526/_0_  ;
	output \g29528/_0_  ;
	output \g29530/_0_  ;
	output \g29532/_0_  ;
	output \g29534/_3_  ;
	output \g29536/_3_  ;
	output \g29538/_3_  ;
	output \g29540/_3_  ;
	output \g29542/_3_  ;
	output \g29544/_3_  ;
	output \g29546/_3_  ;
	output \g29548/_3_  ;
	output \g29550/_0_  ;
	output \g29552/_0_  ;
	output \g29554/_0_  ;
	output \g29556/_0_  ;
	output \g29558/_0_  ;
	output \g29560/_0_  ;
	output \g29562/_0_  ;
	output \g29564/_0_  ;
	output \g29566/_0_  ;
	output \g29568/_0_  ;
	output \g29570/_0_  ;
	output \g29572/_0_  ;
	output \g29574/_3_  ;
	output \g29576/_3_  ;
	output \g29578/_3_  ;
	output \g29580/_3_  ;
	output \g29582/_3_  ;
	output \g29584/_3_  ;
	output \g29586/_3_  ;
	output \g29588/_3_  ;
	output \g29590/_3_  ;
	output \g29592/_3_  ;
	output \g29594/_3_  ;
	output \g29596/_3_  ;
	output \g29598/_3_  ;
	output \g29600/_3_  ;
	output \g29602/_3_  ;
	output \g29604/_3_  ;
	output \g29606/_0_  ;
	output \g29608/_0_  ;
	output \g29610/_0_  ;
	output \g29612/_0_  ;
	output \g29614/_3_  ;
	output \g29616/_3_  ;
	output \g29618/_3_  ;
	output \g29620/_3_  ;
	output \g29622/_3_  ;
	output \g29624/_3_  ;
	output \g29626/_3_  ;
	output \g29628/_3_  ;
	output \g29630/_3_  ;
	output \g29632/_3_  ;
	output \g29634/_3_  ;
	output \g29636/_3_  ;
	output \g29638/_3_  ;
	output \g29640/_3_  ;
	output \g29642/_3_  ;
	output \g29644/_3_  ;
	output \g29646/_3_  ;
	output \g29648/_3_  ;
	output \g29650/_3_  ;
	output \g29652/_3_  ;
	output \g29654/_3_  ;
	output \g29656/_3_  ;
	output \g29658/_3_  ;
	output \g29660/_3_  ;
	output \g29662/_3_  ;
	output \g29664/_3_  ;
	output \g29666/_3_  ;
	output \g29668/_3_  ;
	output \g29670/_3_  ;
	output \g29672/_3_  ;
	output \g29674/_3_  ;
	output \g29676/_3_  ;
	output \g29678/_3_  ;
	output \g29680/_3_  ;
	output \g29682/_3_  ;
	output \g29684/_3_  ;
	output \g29686/_3_  ;
	output \g29688/_3_  ;
	output \g29690/_3_  ;
	output \g29692/_3_  ;
	output \g29694/_0_  ;
	output \g29696/_0_  ;
	output \g29698/_0_  ;
	output \g29700/_0_  ;
	output \g29702/_0_  ;
	output \g29704/_0_  ;
	output \g29706/_0_  ;
	output \g29708/_0_  ;
	output \g29710/_0_  ;
	output \g29712/_0_  ;
	output \g29714/_0_  ;
	output \g29716/_0_  ;
	output \g29718/_0_  ;
	output \g29720/_0_  ;
	output \g29722/_0_  ;
	output \g29724/_0_  ;
	output \g29726/_0_  ;
	output \g29728/_0_  ;
	output \g29730/_0_  ;
	output \g29732/_0_  ;
	output \g29734/_3_  ;
	output \g29736/_3_  ;
	output \g29738/_3_  ;
	output \g29740/_3_  ;
	output \g29742/_3_  ;
	output \g29744/_3_  ;
	output \g29746/_3_  ;
	output \g29748/_3_  ;
	output \g29750/_3_  ;
	output \g29752/_3_  ;
	output \g29754/_3_  ;
	output \g29756/_3_  ;
	output \g29758/_3_  ;
	output \g29760/_3_  ;
	output \g29762/_3_  ;
	output \g29764/_3_  ;
	output \g29766/_3_  ;
	output \g29768/_3_  ;
	output \g29770/_3_  ;
	output \g29772/_3_  ;
	output \g29774/_3_  ;
	output \g29776/_3_  ;
	output \g29778/_3_  ;
	output \g29780/_3_  ;
	output \g29782/_3_  ;
	output \g29784/_3_  ;
	output \g29786/_3_  ;
	output \g29788/_3_  ;
	output \g29790/_3_  ;
	output \g29792/_3_  ;
	output \g29794/_3_  ;
	output \g29796/_3_  ;
	output \g29798/_3_  ;
	output \g29800/_3_  ;
	output \g29802/_3_  ;
	output \g29804/_3_  ;
	output \g29806/_3_  ;
	output \g29808/_3_  ;
	output \g29810/_3_  ;
	output \g29812/_3_  ;
	output \g29814/_3_  ;
	output \g29816/_3_  ;
	output \g29818/_3_  ;
	output \g29820/_3_  ;
	output \g29822/_3_  ;
	output \g29824/_3_  ;
	output \g29826/_3_  ;
	output \g29828/_3_  ;
	output \g29830/_3_  ;
	output \g29832/_3_  ;
	output \g29834/_3_  ;
	output \g29836/_3_  ;
	output \g29838/_3_  ;
	output \g29840/_3_  ;
	output \g29842/_3_  ;
	output \g29844/_3_  ;
	output \g29846/_3_  ;
	output \g29848/_3_  ;
	output \g29850/_3_  ;
	output \g29852/_3_  ;
	output \g29854/_3_  ;
	output \g29856/_3_  ;
	output \g29858/_3_  ;
	output \g29860/_3_  ;
	output \g29862/_3_  ;
	output \g29864/_3_  ;
	output \g29866/_3_  ;
	output \g29868/_3_  ;
	output \g29870/_3_  ;
	output \g29872/_3_  ;
	output \g29874/_3_  ;
	output \g29876/_3_  ;
	output \g29878/_3_  ;
	output \g29880/_3_  ;
	output \g29904/_0_  ;
	output \g29905/_0_  ;
	output \g29906/_0_  ;
	output \g29907/_0_  ;
	output \g29908/_0_  ;
	output \g29909/_0_  ;
	output \g29914/_3_  ;
	output \g29952/_0_  ;
	output \g29953/_0_  ;
	output \g29954/_0_  ;
	output \g29955/_0_  ;
	output \g29956/_0_  ;
	output \g29957/_0_  ;
	output \g29975/_0_  ;
	output \g29976/_0_  ;
	output \g29977/_0_  ;
	output \g29978/_0_  ;
	output \g29979/_0_  ;
	output \g29980/_0_  ;
	output \g29989/_3_  ;
	output \g30020/_0_  ;
	output \g30021/_0_  ;
	output \g30045/_0_  ;
	output \g30046/_0_  ;
	output \g30047/_0_  ;
	output \g30048/_0_  ;
	output \g30049/_0_  ;
	output \g30050/_0_  ;
	output \g30051/_0_  ;
	output \g30052/_0_  ;
	output \g30053/_0_  ;
	output \g30054/_0_  ;
	output \g30062/_0_  ;
	output \g30063/_0_  ;
	output \g30064/_0_  ;
	output \g30065/_0_  ;
	output \g30066/_0_  ;
	output \g30067/_0_  ;
	output \g30068/_0_  ;
	output \g30069/_0_  ;
	output \g30070/_0_  ;
	output \g30071/_0_  ;
	output \g30072/_0_  ;
	output \g30073/_0_  ;
	output \g30074/_0_  ;
	output \g30075/_0_  ;
	output \g30136/_3_  ;
	output \g30707/_0_  ;
	output \g30708/_0_  ;
	output \g30711/_0_  ;
	output \g30714/_0_  ;
	output \g30715/_0_  ;
	output \g30720/_0_  ;
	output \g30725/_0_  ;
	output \g30741/_0_  ;
	output \g30742/_0_  ;
	output \g30743/_0_  ;
	output \g30744/_0_  ;
	output \g30745/_0_  ;
	output \g30746/_0_  ;
	output \g30747/_0_  ;
	output \g30748/_0_  ;
	output \g30749/_0_  ;
	output \g30750/_0_  ;
	output \g30751/_0_  ;
	output \g30752/_0_  ;
	output \g30789/_0_  ;
	output \g30790/_0_  ;
	output \g30791/_0_  ;
	output \g30792/_0_  ;
	output \g30793/_0_  ;
	output \g30794/_0_  ;
	output \g30795/_0_  ;
	output \g30796/_0_  ;
	output \g30797/_0_  ;
	output \g30798/_0_  ;
	output \g30799/_0_  ;
	output \g30800/_0_  ;
	output \g30801/_0_  ;
	output \g30802/_0_  ;
	output \g30803/_0_  ;
	output \g30804/_0_  ;
	output \g30805/_0_  ;
	output \g30806/_0_  ;
	output \g30807/_0_  ;
	output \g30808/_0_  ;
	output \g30809/_0_  ;
	output \g30810/_0_  ;
	output \g30811/_0_  ;
	output \g30812/_0_  ;
	output \g30813/_0_  ;
	output \g30814/_0_  ;
	output \g30815/_0_  ;
	output \g30816/_0_  ;
	output \g30817/_0_  ;
	output \g30818/_0_  ;
	output \g30819/_0_  ;
	output \g30820/_0_  ;
	output \g30821/_0_  ;
	output \g30822/_0_  ;
	output \g30823/_0_  ;
	output \g30824/_0_  ;
	output \g30825/_0_  ;
	output \g30826/_0_  ;
	output \g30827/_0_  ;
	output \g30828/_0_  ;
	output \g30829/_0_  ;
	output \g30830/_0_  ;
	output \g30831/_0_  ;
	output \g30832/_0_  ;
	output \g30833/_0_  ;
	output \g30834/_0_  ;
	output \g30835/_0_  ;
	output \g30836/_0_  ;
	output \g30837/_0_  ;
	output \g30838/_0_  ;
	output \g30839/_0_  ;
	output \g30840/_0_  ;
	output \g30841/_0_  ;
	output \g30842/_0_  ;
	output \g30843/_0_  ;
	output \g30844/_0_  ;
	output \g30845/_0_  ;
	output \g30846/_0_  ;
	output \g30847/_0_  ;
	output \g30848/_0_  ;
	output \g30849/_0_  ;
	output \g30850/_0_  ;
	output \g30851/_0_  ;
	output \g30852/_0_  ;
	output \g30853/_0_  ;
	output \g30854/_0_  ;
	output \g30855/_0_  ;
	output \g30856/_0_  ;
	output \g30857/_0_  ;
	output \g30858/_0_  ;
	output \g30859/_0_  ;
	output \g30860/_0_  ;
	output \g30861/_0_  ;
	output \g30862/_0_  ;
	output \g30863/_0_  ;
	output \g30864/_0_  ;
	output \g30865/_0_  ;
	output \g30866/_0_  ;
	output \g30867/_0_  ;
	output \g30868/_0_  ;
	output \g30869/_0_  ;
	output \g30870/_0_  ;
	output \g30871/_0_  ;
	output \g30872/_0_  ;
	output \g30873/_0_  ;
	output \g30874/_0_  ;
	output \g30875/_0_  ;
	output \g30876/_0_  ;
	output \g30877/_0_  ;
	output \g30878/_0_  ;
	output \g30879/_0_  ;
	output \g30880/_0_  ;
	output \g30881/_0_  ;
	output \g30882/_0_  ;
	output \g30883/_0_  ;
	output \g30884/_0_  ;
	output \g30885/_0_  ;
	output \g30886/_0_  ;
	output \g30887/_0_  ;
	output \g30888/_0_  ;
	output \g30889/_0_  ;
	output \g30890/_0_  ;
	output \g30891/_0_  ;
	output \g30892/_0_  ;
	output \g30893/_0_  ;
	output \g30894/_0_  ;
	output \g30895/_0_  ;
	output \g30896/_0_  ;
	output \g30897/_0_  ;
	output \g30898/_0_  ;
	output \g30899/_0_  ;
	output \g30900/_0_  ;
	output \g30901/_0_  ;
	output \g30902/_0_  ;
	output \g30906/_0_  ;
	output \g30907/_0_  ;
	output \g30908/_0_  ;
	output \g30909/_0_  ;
	output \g30910/_0_  ;
	output \g30911/_0_  ;
	output \g30918/_0_  ;
	output \g30919/_0_  ;
	output \g30920/_0_  ;
	output \g30921/_0_  ;
	output \g30922/_0_  ;
	output \g30923/_0_  ;
	output \g30924/_0_  ;
	output \g30925/_0_  ;
	output \g30926/_0_  ;
	output \g30946/_0_  ;
	output \g30947/_0_  ;
	output \g30948/_0_  ;
	output \g30949/_0_  ;
	output \g30950/_0_  ;
	output \g30951/_0_  ;
	output \g30952/_0_  ;
	output \g30953/_0_  ;
	output \g30954/_0_  ;
	output \g30955/_0_  ;
	output \g30956/_0_  ;
	output \g30957/_0_  ;
	output \g30958/_0_  ;
	output \g30959/_0_  ;
	output \g30960/_0_  ;
	output \g30961/_0_  ;
	output \g30962/_0_  ;
	output \g30963/_0_  ;
	output \g30964/_0_  ;
	output \g30965/_0_  ;
	output \g30966/_0_  ;
	output \g30967/_0_  ;
	output \g30968/_0_  ;
	output \g30969/_0_  ;
	output \g30970/_0_  ;
	output \g30971/_0_  ;
	output \g30972/_0_  ;
	output \g30973/_0_  ;
	output \g30974/_0_  ;
	output \g30975/_0_  ;
	output \g30976/_0_  ;
	output \g30977/_0_  ;
	output \g30978/_0_  ;
	output \g30979/_0_  ;
	output \g30980/_0_  ;
	output \g30981/_0_  ;
	output \g30982/_0_  ;
	output \g30983/_0_  ;
	output \g30984/_0_  ;
	output \g30985/_0_  ;
	output \g30986/_0_  ;
	output \g30987/_0_  ;
	output \g30988/_0_  ;
	output \g30989/_0_  ;
	output \g30990/_0_  ;
	output \g30991/_0_  ;
	output \g30992/_0_  ;
	output \g30993/_0_  ;
	output \g30994/_0_  ;
	output \g30995/_0_  ;
	output \g30996/_0_  ;
	output \g30997/_0_  ;
	output \g30998/_0_  ;
	output \g30999/_0_  ;
	output \g31000/_0_  ;
	output \g31001/_0_  ;
	output \g31002/_0_  ;
	output \g31003/_0_  ;
	output \g31004/_0_  ;
	output \g31005/_0_  ;
	output \g31006/_0_  ;
	output \g31007/_0_  ;
	output \g31008/_0_  ;
	output \g31009/_0_  ;
	output \g31010/_0_  ;
	output \g31011/_0_  ;
	output \g31012/_0_  ;
	output \g31013/_0_  ;
	output \g31014/_0_  ;
	output \g31015/_0_  ;
	output \g31016/_0_  ;
	output \g31017/_0_  ;
	output \g31018/_0_  ;
	output \g31019/_0_  ;
	output \g31020/_0_  ;
	output \g31021/_0_  ;
	output \g31022/_0_  ;
	output \g31023/_0_  ;
	output \g31024/_0_  ;
	output \g31025/_0_  ;
	output \g31026/_0_  ;
	output \g31027/_0_  ;
	output \g31028/_0_  ;
	output \g31029/_0_  ;
	output \g31030/_0_  ;
	output \g31031/_0_  ;
	output \g31032/_0_  ;
	output \g31033/_0_  ;
	output \g31034/_0_  ;
	output \g31035/_0_  ;
	output \g31036/_0_  ;
	output \g31037/_0_  ;
	output \g31038/_0_  ;
	output \g31039/_0_  ;
	output \g31040/_0_  ;
	output \g31041/_0_  ;
	output \g31042/_0_  ;
	output \g31043/_0_  ;
	output \g31044/_0_  ;
	output \g31045/_0_  ;
	output \g31046/_0_  ;
	output \g31047/_0_  ;
	output \g31048/_0_  ;
	output \g31049/_0_  ;
	output \g31050/_0_  ;
	output \g31051/_0_  ;
	output \g31052/_0_  ;
	output \g31053/_0_  ;
	output \g31054/_0_  ;
	output \g31055/_0_  ;
	output \g31056/_0_  ;
	output \g31057/_0_  ;
	output \g31058/_0_  ;
	output \g31059/_0_  ;
	output \g31060/_0_  ;
	output \g31061/_0_  ;
	output \g31062/_0_  ;
	output \g31063/_0_  ;
	output \g31064/_0_  ;
	output \g31065/_0_  ;
	output \g31066/_0_  ;
	output \g31067/_0_  ;
	output \g31068/_0_  ;
	output \g31069/_0_  ;
	output \g31070/_0_  ;
	output \g31071/_0_  ;
	output \g31072/_0_  ;
	output \g31073/_0_  ;
	output \g31074/_0_  ;
	output \g31075/_0_  ;
	output \g31076/_0_  ;
	output \g31077/_0_  ;
	output \g31084/u3_syn_4  ;
	output \g31085/u3_syn_4  ;
	output \g31096/u3_syn_4  ;
	output \g31115/u3_syn_4  ;
	output \g31136/u3_syn_4  ;
	output \g31158/u3_syn_4  ;
	output \g31176/u3_syn_4  ;
	output \g31193/u3_syn_4  ;
	output \g31195/u3_syn_4  ;
	output \g31247/u3_syn_4  ;
	output \g31280/u3_syn_4  ;
	output \g31285/u3_syn_4  ;
	output \g31568/_0_  ;
	output \g31631/_0_  ;
	output \g31672/_0_  ;
	output \g31731/_0_  ;
	output \g31732/_0_  ;
	output \g31742/_2_  ;
	output \g31744/_2_  ;
	output \g31746/_2_  ;
	output \g31748/_2_  ;
	output \g31751/_2_  ;
	output \g31754/_2_  ;
	output \g31756/_2_  ;
	output \g31758/_2_  ;
	output \g31760/_2_  ;
	output \g31761/_0_  ;
	output \g31789/_0_  ;
	output \g31807/_3_  ;
	output \g31825/_3_  ;
	output \g32607/_0_  ;
	output \g32608/_0_  ;
	output \g32609/_0_  ;
	output \g32610/_0_  ;
	output \g32611/_0_  ;
	output \g32612/_0_  ;
	output \g32613/_0_  ;
	output \g32614/_0_  ;
	output \g32615/_0_  ;
	output \g32616/_0_  ;
	output \g32617/_0_  ;
	output \g32618/_0_  ;
	output \g32645/_0__syn_2  ;
	output \g32687/_0__syn_2  ;
	output \g32749/_0__syn_2  ;
	output \g32757/_0_  ;
	output \g32758/_0_  ;
	output \g32759/_0_  ;
	output \g32760/_0_  ;
	output \g32761/_0_  ;
	output \g32762/_0_  ;
	output \g32763/_0_  ;
	output \g32764/_0_  ;
	output \g32765/_0_  ;
	output \g32769/_0_  ;
	output \g32835/_1_  ;
	output \g32839/_0_  ;
	output \g32844/_0_  ;
	output \g32901/_1_  ;
	output \g32902/_0_  ;
	output \g32963/_1_  ;
	output \g32972/_0_  ;
	output \g32977/_0_  ;
	output \g32979/_0_  ;
	output \g32980/_0_  ;
	output \g32981/_0_  ;
	output \g32982/_0_  ;
	output \g32983/_0_  ;
	output \g32987/_0_  ;
	output \g33018/_0_  ;
	output \g33019/_0_  ;
	output \g33088/_0_  ;
	output \g33261/_0_  ;
	output \g33264/_0_  ;
	output \g33275/_0_  ;
	output \g33276/_0_  ;
	output \g33277/_0_  ;
	output \g33371/_0_  ;
	output \g33382/_0_  ;
	output \g33401/_0_  ;
	output \g33402/_0_  ;
	output \g33403/_0_  ;
	output \g33404/_0_  ;
	output \g33405/_0_  ;
	output \g33406/_0_  ;
	output \g33407/_0_  ;
	output \g33408/_0_  ;
	output \g33409/_0_  ;
	output \g33410/_0_  ;
	output \g33411/_0_  ;
	output \g33412/_0_  ;
	output \g33413/_0_  ;
	output \g33414/_0_  ;
	output \g33415/_0_  ;
	output \g33416/_0_  ;
	output \g33417/_0_  ;
	output \g33418/_0_  ;
	output \g33419/_0_  ;
	output \g33420/_0_  ;
	output \g33421/_0_  ;
	output \g33422/_0_  ;
	output \g33423/_0_  ;
	output \g33424/_0_  ;
	output \g33425/_0_  ;
	output \g33426/_0_  ;
	output \g33427/_0_  ;
	output \g33428/_0_  ;
	output \g33429/_0_  ;
	output \g33430/_0_  ;
	output \g33431/_0_  ;
	output \g33432/_0_  ;
	output \g33433/_0_  ;
	output \g33434/_0_  ;
	output \g33435/_0_  ;
	output \g33436/_0_  ;
	output \g33437/_0_  ;
	output \g33438/_0_  ;
	output \g33439/_0_  ;
	output \g33440/_0_  ;
	output \g33441/_0_  ;
	output \g33442/_0_  ;
	output \g33443/_0_  ;
	output \g33444/_0_  ;
	output \g33445/_0_  ;
	output \g33446/_0_  ;
	output \g33447/_0_  ;
	output \g33448/_0_  ;
	output \g33449/_0_  ;
	output \g33450/_0_  ;
	output \g33451/_0_  ;
	output \g33452/_0_  ;
	output \g33453/_0_  ;
	output \g33454/_0_  ;
	output \g33455/_0_  ;
	output \g33456/_0_  ;
	output \g33457/_0_  ;
	output \g33458/_0_  ;
	output \g33459/_0_  ;
	output \g33460/_0_  ;
	output \g33461/_0_  ;
	output \g33462/_0_  ;
	output \g33463/_0_  ;
	output \g33464/_0_  ;
	output \g33465/_0_  ;
	output \g33466/_0_  ;
	output \g33467/_0_  ;
	output \g33468/_0_  ;
	output \g33469/_0_  ;
	output \g33470/_0_  ;
	output \g33471/_0_  ;
	output \g33472/_0_  ;
	output \g33473/_0_  ;
	output \g33474/_0_  ;
	output \g33475/_0_  ;
	output \g33476/_0_  ;
	output \g33477/_0_  ;
	output \g33478/_0_  ;
	output \g33479/_0_  ;
	output \g33480/_0_  ;
	output \g33481/_0_  ;
	output \g33482/_0_  ;
	output \g33483/_0_  ;
	output \g33484/_0_  ;
	output \g33485/_0_  ;
	output \g33486/_0_  ;
	output \g33487/_0_  ;
	output \g33488/_0_  ;
	output \g33489/_0_  ;
	output \g33490/_0_  ;
	output \g33491/_0_  ;
	output \g33492/_0_  ;
	output \g33493/_0_  ;
	output \g33494/_0_  ;
	output \g33495/_0_  ;
	output \g33496/_0_  ;
	output \g33497/_0_  ;
	output \g33498/_0_  ;
	output \g33499/_0_  ;
	output \g33500/_0_  ;
	output \g33501/_0_  ;
	output \g33502/_0_  ;
	output \g33503/_0_  ;
	output \g33504/_0_  ;
	output \g33505/_0_  ;
	output \g33506/_0_  ;
	output \g33507/_0_  ;
	output \g33508/_0_  ;
	output \g33509/_0_  ;
	output \g33510/_0_  ;
	output \g33511/_0_  ;
	output \g33512/_0_  ;
	output \g33513/_0_  ;
	output \g33514/_0_  ;
	output \g33515/_0_  ;
	output \g33516/_0_  ;
	output \g33517/_0_  ;
	output \g33518/_0_  ;
	output \g33519/_0_  ;
	output \g33520/_0_  ;
	output \g33521/_0_  ;
	output \g33522/_0_  ;
	output \g33523/_0_  ;
	output \g33524/_0_  ;
	output \g33525/_0_  ;
	output \g33526/_0_  ;
	output \g33527/_0_  ;
	output \g33528/_0_  ;
	output \g33529/_0_  ;
	output \g33530/_0_  ;
	output \g33531/_0_  ;
	output \g33532/_0_  ;
	output \g33533/_0_  ;
	output \g33534/_0_  ;
	output \g33535/_0_  ;
	output \g33536/_0_  ;
	output \g33537/_0_  ;
	output \g33538/_0_  ;
	output \g33539/_0_  ;
	output \g33540/_0_  ;
	output \g33541/_0_  ;
	output \g33542/_0_  ;
	output \g33543/_0_  ;
	output \g33544/_0_  ;
	output \g33545/_0_  ;
	output \g33546/_0_  ;
	output \g33547/_0_  ;
	output \g33548/_0_  ;
	output \g33549/_0_  ;
	output \g33550/_0_  ;
	output \g33551/_0_  ;
	output \g33552/_0_  ;
	output \g33553/_0_  ;
	output \g33554/_0_  ;
	output \g33555/_0_  ;
	output \g33556/_0_  ;
	output \g33557/_0_  ;
	output \g33558/_0_  ;
	output \g33559/_0_  ;
	output \g33560/_0_  ;
	output \g33561/_0_  ;
	output \g33562/_0_  ;
	output \g33563/_0_  ;
	output \g33564/_0_  ;
	output \g33565/_0_  ;
	output \g33566/_0_  ;
	output \g33567/_0_  ;
	output \g33568/_0_  ;
	output \g33569/_0_  ;
	output \g33570/_0_  ;
	output \g33571/_0_  ;
	output \g33572/_0_  ;
	output \g33573/_0_  ;
	output \g33574/_0_  ;
	output \g33575/_0_  ;
	output \g33576/_0_  ;
	output \g33577/_0_  ;
	output \g33578/_0_  ;
	output \g33579/_0_  ;
	output \g33580/_0_  ;
	output \g33581/_0_  ;
	output \g33582/_0_  ;
	output \g33583/_0_  ;
	output \g33584/_0_  ;
	output \g33585/_0_  ;
	output \g33586/_0_  ;
	output \g33587/_0_  ;
	output \g33588/_0_  ;
	output \g33589/_0_  ;
	output \g33590/_0_  ;
	output \g33591/_0_  ;
	output \g33592/_0_  ;
	output \g33593/_0_  ;
	output \g33594/_0_  ;
	output \g33595/_0_  ;
	output \g33596/_0_  ;
	output \g33597/_0_  ;
	output \g33598/_0_  ;
	output \g33599/_0_  ;
	output \g33600/_0_  ;
	output \g33601/_0_  ;
	output \g33602/_0_  ;
	output \g33603/_0_  ;
	output \g33604/_0_  ;
	output \g33605/_0_  ;
	output \g33606/_0_  ;
	output \g33607/_0_  ;
	output \g33608/_0_  ;
	output \g33609/_0_  ;
	output \g33610/_0_  ;
	output \g33611/_0_  ;
	output \g33612/_0_  ;
	output \g33613/_0_  ;
	output \g33614/_0_  ;
	output \g33615/_0_  ;
	output \g33616/_0_  ;
	output \g33617/_0_  ;
	output \g33618/_0_  ;
	output \g33619/_0_  ;
	output \g33620/_0_  ;
	output \g33621/_0_  ;
	output \g33622/_0_  ;
	output \g33623/_0_  ;
	output \g33624/_0_  ;
	output \g33625/_0_  ;
	output \g33626/_0_  ;
	output \g33627/_0_  ;
	output \g33628/_0_  ;
	output \g33629/_0_  ;
	output \g33630/_0_  ;
	output \g33631/_0_  ;
	output \g33632/_0_  ;
	output \g33633/_0_  ;
	output \g33634/_0_  ;
	output \g33635/_0_  ;
	output \g33636/_0_  ;
	output \g33637/_0_  ;
	output \g33638/_0_  ;
	output \g33639/_0_  ;
	output \g33640/_0_  ;
	output \g33641/_0_  ;
	output \g33642/_0_  ;
	output \g33643/_0_  ;
	output \g33644/_0_  ;
	output \g33645/_0_  ;
	output \g33646/_0_  ;
	output \g33647/_0_  ;
	output \g33648/_0_  ;
	output \g33649/_0_  ;
	output \g33650/_0_  ;
	output \g33651/_0_  ;
	output \g33652/_0_  ;
	output \g33653/_0_  ;
	output \g33654/_0_  ;
	output \g33655/_0_  ;
	output \g33656/_0_  ;
	output \g33657/_0_  ;
	output \g33658/_0_  ;
	output \g33659/_0_  ;
	output \g33660/_0_  ;
	output \g33661/_0_  ;
	output \g33662/_0_  ;
	output \g33663/_0_  ;
	output \g33664/_0_  ;
	output \g33665/_0_  ;
	output \g33666/_0_  ;
	output \g33667/_0_  ;
	output \g33668/_0_  ;
	output \g33669/_0_  ;
	output \g33670/_0_  ;
	output \g33671/_0_  ;
	output \g33672/_0_  ;
	output \g33673/_0_  ;
	output \g33674/_0_  ;
	output \g33675/_0_  ;
	output \g33676/_0_  ;
	output \g33677/_0_  ;
	output \g33678/_0_  ;
	output \g33679/_0_  ;
	output \g33680/_0_  ;
	output \g33681/_0_  ;
	output \g33682/_0_  ;
	output \g33683/_0_  ;
	output \g33684/_0_  ;
	output \g33685/_0_  ;
	output \g33686/_0_  ;
	output \g33687/_0_  ;
	output \g33688/_0_  ;
	output \g33689/_0_  ;
	output \g33690/_0_  ;
	output \g33691/_0_  ;
	output \g33692/_0_  ;
	output \g33693/_0_  ;
	output \g33694/_0_  ;
	output \g33695/_0_  ;
	output \g33696/_0_  ;
	output \g33697/_0_  ;
	output \g33698/_0_  ;
	output \g33699/_0_  ;
	output \g33700/_0_  ;
	output \g33701/_0_  ;
	output \g33702/_0_  ;
	output \g33703/_0_  ;
	output \g33704/_0_  ;
	output \g33705/_0_  ;
	output \g33706/_0_  ;
	output \g33707/_0_  ;
	output \g33708/_0_  ;
	output \g33709/_0_  ;
	output \g33710/_0_  ;
	output \g33711/_0_  ;
	output \g33712/_0_  ;
	output \g33713/_0_  ;
	output \g33714/_0_  ;
	output \g33715/_0_  ;
	output \g33716/_0_  ;
	output \g33717/_0_  ;
	output \g33718/_0_  ;
	output \g33719/_0_  ;
	output \g33720/_0_  ;
	output \g33721/_0_  ;
	output \g33722/_0_  ;
	output \g33723/_0_  ;
	output \g33724/_0_  ;
	output \g33725/_0_  ;
	output \g33726/_0_  ;
	output \g33727/_0_  ;
	output \g33728/_0_  ;
	output \g33729/_0_  ;
	output \g33730/_0_  ;
	output \g33731/_0_  ;
	output \g33732/_0_  ;
	output \g33733/_0_  ;
	output \g33734/_0_  ;
	output \g33735/_0_  ;
	output \g33736/_0_  ;
	output \g33737/_0_  ;
	output \g33738/_0_  ;
	output \g33739/_0_  ;
	output \g33740/_0_  ;
	output \g33741/_0_  ;
	output \g33742/_0_  ;
	output \g33743/_0_  ;
	output \g33744/_0_  ;
	output \g33745/_0_  ;
	output \g33746/_0_  ;
	output \g33747/_0_  ;
	output \g33748/_0_  ;
	output \g33749/_0_  ;
	output \g33750/_0_  ;
	output \g33751/_0_  ;
	output \g33752/_0_  ;
	output \g33753/_0_  ;
	output \g33754/_0_  ;
	output \g33755/_0_  ;
	output \g33756/_0_  ;
	output \g33757/_0_  ;
	output \g33758/_0_  ;
	output \g33759/_0_  ;
	output \g33760/_0_  ;
	output \g33761/_0_  ;
	output \g33762/_0_  ;
	output \g33763/_0_  ;
	output \g33764/_0_  ;
	output \g33765/_0_  ;
	output \g33766/_0_  ;
	output \g33767/_0_  ;
	output \g33768/_0_  ;
	output \g33769/_0_  ;
	output \g33770/_0_  ;
	output \g33771/_0_  ;
	output \g33772/_0_  ;
	output \g33773/_0_  ;
	output \g33774/_0_  ;
	output \g33775/_0_  ;
	output \g33776/_0_  ;
	output \g33777/_0_  ;
	output \g33778/_0_  ;
	output \g33779/_0_  ;
	output \g33780/_0_  ;
	output \g33781/_0_  ;
	output \g33782/_0_  ;
	output \g33783/_0_  ;
	output \g33784/_0_  ;
	output \g33785/_0_  ;
	output \g33786/_0_  ;
	output \g33787/_0_  ;
	output \g33788/_0_  ;
	output \g33789/_0_  ;
	output \g33790/_0_  ;
	output \g33791/_0_  ;
	output \g33792/_0_  ;
	output \g33793/_0_  ;
	output \g33794/_0_  ;
	output \g33795/_0_  ;
	output \g33796/_0_  ;
	output \g33797/_0_  ;
	output \g33798/_0_  ;
	output \g33799/_0_  ;
	output \g33800/_0_  ;
	output \g33801/_0_  ;
	output \g33802/_0_  ;
	output \g33803/_0_  ;
	output \g33804/_0_  ;
	output \g33805/_0_  ;
	output \g33806/_0_  ;
	output \g33807/_0_  ;
	output \g33808/_0_  ;
	output \g33809/_0_  ;
	output \g33810/_0_  ;
	output \g33811/_0_  ;
	output \g33812/_0_  ;
	output \g33813/_0_  ;
	output \g33814/_0_  ;
	output \g33815/_0_  ;
	output \g33816/_0_  ;
	output \g33817/_0_  ;
	output \g33818/_0_  ;
	output \g33819/_0_  ;
	output \g33820/_0_  ;
	output \g33821/_0_  ;
	output \g33822/_0_  ;
	output \g33823/_0_  ;
	output \g33824/_0_  ;
	output \g33825/_0_  ;
	output \g33826/_0_  ;
	output \g33827/_0_  ;
	output \g33828/_0_  ;
	output \g33829/_0_  ;
	output \g33830/_0_  ;
	output \g33831/_0_  ;
	output \g33832/_0_  ;
	output \g33833/_0_  ;
	output \g33834/_0_  ;
	output \g33835/_0_  ;
	output \g33836/_0_  ;
	output \g33837/_0_  ;
	output \g33838/_0_  ;
	output \g33839/_0_  ;
	output \g33840/_0_  ;
	output \g33841/_0_  ;
	output \g33842/_0_  ;
	output \g33843/_0_  ;
	output \g33844/_0_  ;
	output \g33845/_0_  ;
	output \g33846/_0_  ;
	output \g33847/_0_  ;
	output \g33848/_0_  ;
	output \g33849/_0_  ;
	output \g33850/_0_  ;
	output \g33851/_0_  ;
	output \g33852/_0_  ;
	output \g33853/_0_  ;
	output \g33854/_0_  ;
	output \g33855/_0_  ;
	output \g33856/_0_  ;
	output \g33857/_0_  ;
	output \g33858/_0_  ;
	output \g33859/_0_  ;
	output \g33860/_0_  ;
	output \g33861/_0_  ;
	output \g33862/_0_  ;
	output \g33863/_0_  ;
	output \g33864/_0_  ;
	output \g33865/_0_  ;
	output \g33866/_0_  ;
	output \g33867/_0_  ;
	output \g33868/_0_  ;
	output \g33869/_0_  ;
	output \g33870/_0_  ;
	output \g33871/_0_  ;
	output \g33872/_0_  ;
	output \g33873/_0_  ;
	output \g33874/_0_  ;
	output \g33875/_0_  ;
	output \g33876/_0_  ;
	output \g33877/_0_  ;
	output \g33878/_0_  ;
	output \g33879/_0_  ;
	output \g33880/_0_  ;
	output \g33881/_0_  ;
	output \g33882/_0_  ;
	output \g33883/_0_  ;
	output \g33884/_0_  ;
	output \g33885/_0_  ;
	output \g33886/_0_  ;
	output \g33887/_0_  ;
	output \g33888/_0_  ;
	output \g33889/_0_  ;
	output \g33890/_0_  ;
	output \g33891/_0_  ;
	output \g33892/_0_  ;
	output \g33893/_0_  ;
	output \g33894/_0_  ;
	output \g33895/_0_  ;
	output \g33896/_0_  ;
	output \g33897/_0_  ;
	output \g33898/_0_  ;
	output \g33899/_0_  ;
	output \g33900/_0_  ;
	output \g33901/_0_  ;
	output \g33902/_0_  ;
	output \g33903/_0_  ;
	output \g33904/_0_  ;
	output \g33905/_0_  ;
	output \g33906/_0_  ;
	output \g33907/_0_  ;
	output \g33908/_0_  ;
	output \g33909/_0_  ;
	output \g33910/_0_  ;
	output \g33911/_0_  ;
	output \g33912/_0_  ;
	output \g33913/_0_  ;
	output \g33914/_0_  ;
	output \g33915/_0_  ;
	output \g33916/_0_  ;
	output \g33917/_0_  ;
	output \g33918/_0_  ;
	output \g33919/_0_  ;
	output \g33920/_0_  ;
	output \g33921/_0_  ;
	output \g33922/_0_  ;
	output \g33923/_0_  ;
	output \g33924/_0_  ;
	output \g33925/_0_  ;
	output \g33926/_0_  ;
	output \g33927/_0_  ;
	output \g33928/_0_  ;
	output \g33929/_0_  ;
	output \g33930/_0_  ;
	output \g33931/_0_  ;
	output \g33932/_0_  ;
	output \g33933/_0_  ;
	output \g33934/_0_  ;
	output \g33935/_0_  ;
	output \g33936/_0_  ;
	output \g33937/_0_  ;
	output \g33938/_0_  ;
	output \g33939/_0_  ;
	output \g33940/_0_  ;
	output \g33941/_0_  ;
	output \g33942/_0_  ;
	output \g33943/_0_  ;
	output \g33944/_0_  ;
	output \g33945/_0_  ;
	output \g33946/_0_  ;
	output \g33947/_0_  ;
	output \g33948/_0_  ;
	output \g33949/_0_  ;
	output \g33950/_0_  ;
	output \g33951/_0_  ;
	output \g33952/_0_  ;
	output \g33953/_0_  ;
	output \g33954/_0_  ;
	output \g33955/_0_  ;
	output \g33956/_0_  ;
	output \g33957/_0_  ;
	output \g33958/_0_  ;
	output \g33959/_0_  ;
	output \g33960/_0_  ;
	output \g33961/_0_  ;
	output \g33962/_0_  ;
	output \g33963/_0_  ;
	output \g33964/_0_  ;
	output \g33965/_0_  ;
	output \g33966/_0_  ;
	output \g33967/_0_  ;
	output \g33968/_0_  ;
	output \g33969/_0_  ;
	output \g33970/_0_  ;
	output \g33971/_0_  ;
	output \g33972/_0_  ;
	output \g33973/_0_  ;
	output \g33974/_0_  ;
	output \g33975/_0_  ;
	output \g33976/_0_  ;
	output \g33977/u3_syn_4  ;
	output \g33981/u3_syn_4  ;
	output \g34014/u3_syn_4  ;
	output \g34047/u3_syn_4  ;
	output \g34084/u3_syn_4  ;
	output \g34123/u3_syn_4  ;
	output \g34306/_0_  ;
	output \g34316/_0_  ;
	output \g34324/_0_  ;
	output \g34326/_0_  ;
	output \g34328/_0_  ;
	output \g34331/_0_  ;
	output \g34333/_0_  ;
	output \g34344/_0_  ;
	output \g34347/_0_  ;
	output \g34351/_0_  ;
	output \g34361/_0_  ;
	output \g34368/_0_  ;
	output \g34377/_0_  ;
	output \g34385/_0_  ;
	output \g34393/_0_  ;
	output \g34414/_1_  ;
	output \g34451/_1_  ;
	output \g34476/_1_  ;
	output \g34487/_0_  ;
	output \g34490/_1_  ;
	output \g34715/_0_  ;
	output \g34878/_0_  ;
	output \g34882/_0_  ;
	output \g34883/_0_  ;
	output \g34893/_0_  ;
	output \g34896/_0_  ;
	output \g34898/_0_  ;
	output \g34899/_0_  ;
	output \g34916/_3_  ;
	output \g35264/_0_  ;
	output \g35265/_0_  ;
	output \g35266/_0_  ;
	output \g35267/_0_  ;
	output \g35268/_0_  ;
	output \g35269/_0_  ;
	output \g35270/_0_  ;
	output \g35271/_0_  ;
	output \g35272/_0_  ;
	output \g35273/_0_  ;
	output \g35274/_0_  ;
	output \g35275/_0_  ;
	output \g35276/_0_  ;
	output \g35277/_0_  ;
	output \g35278/_0_  ;
	output \g35279/_0_  ;
	output \g35283/_0_  ;
	output \g35287/_0_  ;
	output \g35294/_0_  ;
	output \g35300/_0_  ;
	output \g35304/_0_  ;
	output \g35308/_0_  ;
	output \g35312/_0_  ;
	output \g35316/_0_  ;
	output \g35318/_0_  ;
	output \g35326/_0_  ;
	output \g35334/_0_  ;
	output \g35336/_0_  ;
	output \g35337/_0_  ;
	output \g35338/_0_  ;
	output \g35357/_0_  ;
	output \g35358/_0_  ;
	output \g35359/_0_  ;
	output \g35419/_0_  ;
	output \g35438/_0_  ;
	output \g35439/_0_  ;
	output \g35440/_0_  ;
	output \g35441/_0_  ;
	output \g35442/_0_  ;
	output \g35444/_0_  ;
	output \g35445/_0_  ;
	output \g35446/_0_  ;
	output \g35447/_0_  ;
	output \g35448/_0_  ;
	output \g35449/_0_  ;
	output \g35450/_0_  ;
	output \g35451/_0_  ;
	output \g35452/_0_  ;
	output \g35463/_0_  ;
	output \g35464/_0_  ;
	output \g35466/_0_  ;
	output \g35485/_2_  ;
	output \g35495/_0_  ;
	output \g35496/_0_  ;
	output \g35499/_0_  ;
	output \g35500/_0_  ;
	output \g35501/_0_  ;
	output \g35502/_0_  ;
	output \g35563/_0_  ;
	output \g35633/_0_  ;
	output \g35717/_0_  ;
	output \g35718/_0_  ;
	output \g35719/_0_  ;
	output \g35809/_0_  ;
	output \g35810/_0_  ;
	output \g35811/_0_  ;
	output \g35812/_0_  ;
	output \g35813/_0_  ;
	output \g35814/_0_  ;
	output \g35815/_0_  ;
	output \g35816/_0_  ;
	output \g35817/_0_  ;
	output \g35818/_0_  ;
	output \g35819/_0_  ;
	output \g35820/_0_  ;
	output \g35821/_0_  ;
	output \g35822/_0_  ;
	output \g35823/_0_  ;
	output \g35824/_0_  ;
	output \g35825/_0_  ;
	output \g35826/_0_  ;
	output \g35827/_0_  ;
	output \g35830/_0_  ;
	output \g35833/_0_  ;
	output \g35835/_0_  ;
	output \g35836/_0_  ;
	output \g35837/_0_  ;
	output \g35839/_0_  ;
	output \g35840/_0_  ;
	output \g35841/_0_  ;
	output \g35843/_0_  ;
	output \g35844/_0_  ;
	output \g35845/_0_  ;
	output \g35853/_0_  ;
	output \g35854/_0_  ;
	output \g35855/_0_  ;
	output \g35856/_0_  ;
	output \g36306/_0_  ;
	output \g36414/_0_  ;
	output \g36415/_0_  ;
	output \g36449/_0_  ;
	output \g36550/_0_  ;
	output \g36551/_0_  ;
	output \g36553/_0_  ;
	output \g36560/_0_  ;
	output \g36562/_3_  ;
	output \g36563/_0_  ;
	output \g36612/_0_  ;
	output \g36614/_2_  ;
	output \g36695/_0_  ;
	output \g36784/_0_  ;
	output \g36785/_0_  ;
	output \g36786/_0_  ;
	output \g36787/_0_  ;
	output \g36788/_0_  ;
	output \g36789/_0_  ;
	output \g36790/_0_  ;
	output \g36791/_0_  ;
	output \g36792/_0_  ;
	output \g36793/_0_  ;
	output \g36794/_0_  ;
	output \g36796/_0_  ;
	output \g36797/_0_  ;
	output \g36798/_0_  ;
	output \g36799/_0_  ;
	output \g36800/_0_  ;
	output \g36801/_0_  ;
	output \g36802/_0_  ;
	output \g36803/_0_  ;
	output \g36804/_0_  ;
	output \g36805/_0_  ;
	output \g36806/_0_  ;
	output \g36807/_0_  ;
	output \g36808/_0_  ;
	output \g36809/_0_  ;
	output \g36810/_0_  ;
	output \g36811/_0_  ;
	output \g36813/_0_  ;
	output \g36814/_0_  ;
	output \g36815/_0_  ;
	output \g36820/_0_  ;
	output \g36825/_0_  ;
	output \g36832/_0_  ;
	output \g36846/_0_  ;
	output \g36855/_0_  ;
	output \g36857/_0_  ;
	output \g36859/_0_  ;
	output \g36860/_0_  ;
	output \g36861/_0_  ;
	output \g36862/_0_  ;
	output \g36863/_0_  ;
	output \g36864/_0_  ;
	output \g36867/_0_  ;
	output \g36870/_0_  ;
	output \g36871/_0_  ;
	output \g36877/_0_  ;
	output \g36879/_0_  ;
	output \g36892/_0_  ;
	output \g36893/_0_  ;
	output \g36901/_0_  ;
	output \g36909/_0_  ;
	output \g36914/_0_  ;
	output \g36919/_0_  ;
	output \g36922/_0_  ;
	output \g36923/_0_  ;
	output \g36927/_0_  ;
	output \g36930/_0_  ;
	output \g36931/_0_  ;
	output \g36933/_0_  ;
	output \g36934/_0_  ;
	output \g36935/_0_  ;
	output \g36936/_0_  ;
	output \g36937/_0_  ;
	output \g36938/_0_  ;
	output \g36939/_0_  ;
	output \g36940/_0_  ;
	output \g36941/_0_  ;
	output \g36943/_0_  ;
	output \g36944/_0_  ;
	output \g36945/_0_  ;
	output \g36946/_0_  ;
	output \g36947/_0_  ;
	output \g36948/_0_  ;
	output \g36949/_0_  ;
	output \g36950/_0_  ;
	output \g36951/_0_  ;
	output \g36952/_0_  ;
	output \g36953/_0_  ;
	output \g36954/_0_  ;
	output \g36957/_0_  ;
	output \g36958/_0_  ;
	output \g36959/_0_  ;
	output \g36960/_0_  ;
	output \g36961/_0_  ;
	output \g36962/_0_  ;
	output \g36963/_0_  ;
	output \g36970/_0_  ;
	output \g36977/_0_  ;
	output \g36986/_0_  ;
	output \g36991/_0_  ;
	output \g36994/_0_  ;
	output \g37015/_0_  ;
	output \g37057/_0_  ;
	output \g37073/_0_  ;
	output \g37128/_0_  ;
	output \g37129/_0_  ;
	output \g37138/_0_  ;
	output \g37139/_0_  ;
	output \g37140/_0_  ;
	output \g37141/_0_  ;
	output \g37142/_0_  ;
	output \g37143/_0_  ;
	output \g37144/_0_  ;
	output \g37145/_0_  ;
	output \g37146/_0_  ;
	output \g37147/_0_  ;
	output \g37148/_0_  ;
	output \g37149/_0_  ;
	output \g37150/_0_  ;
	output \g37151/_0_  ;
	output \g37152/_0_  ;
	output \g37153/_0_  ;
	output \g37154/_0_  ;
	output \g37155/_0_  ;
	output \g37156/_0_  ;
	output \g37157/_0_  ;
	output \g37158/_0_  ;
	output \g37159/_0_  ;
	output \g37160/_0_  ;
	output \g37161/_0_  ;
	output \g37162/_0_  ;
	output \g37163/_0_  ;
	output \g37164/_0_  ;
	output \g37165/_0_  ;
	output \g37166/_0_  ;
	output \g37167/_0_  ;
	output \g37168/_0_  ;
	output \g37169/_0_  ;
	output \g37170/_0_  ;
	output \g37171/_0_  ;
	output \g37172/_0_  ;
	output \g37173/_0_  ;
	output \g37174/_0_  ;
	output \g37175/_0_  ;
	output \g37176/_0_  ;
	output \g37177/_0_  ;
	output \g37178/_0_  ;
	output \g37179/_0_  ;
	output \g37180/_0_  ;
	output \g37181/_0_  ;
	output \g37182/_0_  ;
	output \g37183/_0_  ;
	output \g37184/_0_  ;
	output \g37185/_0_  ;
	output \g37187/_0_  ;
	output \g37188/_0_  ;
	output \g37190/_0_  ;
	output \g37191/_0_  ;
	output \g37192/_0_  ;
	output \g37193/_0_  ;
	output \g37194/_0_  ;
	output \g37372/_3_  ;
	output \g37377/_0_  ;
	output \g37378/_0_  ;
	output \g37379/_0_  ;
	output \g37380/_0_  ;
	output \g37381/_0_  ;
	output \g37382/_0_  ;
	output \g37383/_0_  ;
	output \g37384/_0_  ;
	output \g37385/_0_  ;
	output \g37386/_0_  ;
	output \g37387/_0_  ;
	output \g37388/_0_  ;
	output \g37389/_0_  ;
	output \g37390/_0_  ;
	output \g37391/_0_  ;
	output \g37392/_0_  ;
	output \g37393/_0_  ;
	output \g37394/_0_  ;
	output \g37395/_0_  ;
	output \g37396/_0_  ;
	output \g37397/_0_  ;
	output \g37398/_0_  ;
	output \g37399/_0_  ;
	output \g37400/_0_  ;
	output \g37401/_0_  ;
	output \g37402/_0_  ;
	output \g37403/_0_  ;
	output \g37404/_0_  ;
	output \g37405/_0_  ;
	output \g37406/_0_  ;
	output \g37407/_0_  ;
	output \g37408/_0_  ;
	output \g37409/_0_  ;
	output \g37410/_0_  ;
	output \g37411/_0_  ;
	output \g37412/_0_  ;
	output \g37413/_0_  ;
	output \g37576/_3_  ;
	output \g37590/_2_  ;
	output \g40278/_0_  ;
	output \g40379/_0_  ;
	output \g40389/_2_  ;
	output \g40390/_2_  ;
	output \g40391/_0_  ;
	output \g40393/_2_  ;
	output \g40395/_0_  ;
	output \g40397/_0_  ;
	output \g40400/_0_  ;
	output \g40402/_0_  ;
	output \g45458/_0_  ;
	output \g45675/_0_  ;
	output \g45677/_0_  ;
	output \g45678/_0_  ;
	output \g45682/_0_  ;
	output sync_pad_o_pad ;
	output \u14_u0_full_empty_r_reg/P0001_reg_syn_3  ;
	output \u14_u1_full_empty_r_reg/P0001_reg_syn_3  ;
	output \u14_u2_full_empty_r_reg/P0001_reg_syn_3  ;
	output \u14_u3_full_empty_r_reg/P0001_reg_syn_3  ;
	output \u14_u4_full_empty_r_reg/P0001_reg_syn_3  ;
	output \u14_u5_full_empty_r_reg/P0001_reg_syn_3  ;
	output \u14_u6_full_empty_r_reg/P0001_reg_syn_3  ;
	output \u14_u7_full_empty_r_reg/P0001_reg_syn_3  ;
	output \u14_u8_full_empty_r_reg/P0001_reg_syn_3  ;
	output \u1_slt0_reg[11]/P0001_reg_syn_3  ;
	output \u1_slt0_reg[12]/P0001_reg_syn_3  ;
	output \u1_slt0_reg[15]/P0001_reg_syn_3  ;
	output \u1_slt0_reg[9]/P0001_reg_syn_3  ;
	output \u1_slt1_reg[10]/P0001_reg_syn_3  ;
	output \u1_slt1_reg[11]/P0001_reg_syn_3  ;
	output \u1_slt1_reg[5]/P0001_reg_syn_3  ;
	output \u1_slt1_reg[6]/P0001_reg_syn_3  ;
	output \u1_slt1_reg[7]/P0001_reg_syn_3  ;
	output \u1_slt1_reg[8]/P0001_reg_syn_3  ;
	output wb_err_o_pad ;
	wire _w7143_ ;
	wire _w7142_ ;
	wire _w7141_ ;
	wire _w7140_ ;
	wire _w7139_ ;
	wire _w7138_ ;
	wire _w7137_ ;
	wire _w7136_ ;
	wire _w7135_ ;
	wire _w7134_ ;
	wire _w7133_ ;
	wire _w7132_ ;
	wire _w7131_ ;
	wire _w7130_ ;
	wire _w7129_ ;
	wire _w7128_ ;
	wire _w7127_ ;
	wire _w7126_ ;
	wire _w7125_ ;
	wire _w7124_ ;
	wire _w7123_ ;
	wire _w7122_ ;
	wire _w7121_ ;
	wire _w7120_ ;
	wire _w7119_ ;
	wire _w7118_ ;
	wire _w7117_ ;
	wire _w7116_ ;
	wire _w7115_ ;
	wire _w7114_ ;
	wire _w7113_ ;
	wire _w7112_ ;
	wire _w7111_ ;
	wire _w7110_ ;
	wire _w7109_ ;
	wire _w7108_ ;
	wire _w7107_ ;
	wire _w7106_ ;
	wire _w7105_ ;
	wire _w7104_ ;
	wire _w7103_ ;
	wire _w7102_ ;
	wire _w7101_ ;
	wire _w7100_ ;
	wire _w7099_ ;
	wire _w7098_ ;
	wire _w7097_ ;
	wire _w7096_ ;
	wire _w7095_ ;
	wire _w7094_ ;
	wire _w7093_ ;
	wire _w7092_ ;
	wire _w7091_ ;
	wire _w7090_ ;
	wire _w7089_ ;
	wire _w7088_ ;
	wire _w7087_ ;
	wire _w7086_ ;
	wire _w7085_ ;
	wire _w7084_ ;
	wire _w7083_ ;
	wire _w7082_ ;
	wire _w7081_ ;
	wire _w7080_ ;
	wire _w7079_ ;
	wire _w7078_ ;
	wire _w7077_ ;
	wire _w7076_ ;
	wire _w7075_ ;
	wire _w7074_ ;
	wire _w7073_ ;
	wire _w7072_ ;
	wire _w7071_ ;
	wire _w7070_ ;
	wire _w7069_ ;
	wire _w7068_ ;
	wire _w7067_ ;
	wire _w7066_ ;
	wire _w7065_ ;
	wire _w7064_ ;
	wire _w7063_ ;
	wire _w7062_ ;
	wire _w7061_ ;
	wire _w7060_ ;
	wire _w7059_ ;
	wire _w7058_ ;
	wire _w7057_ ;
	wire _w7056_ ;
	wire _w7055_ ;
	wire _w7054_ ;
	wire _w7053_ ;
	wire _w7052_ ;
	wire _w7051_ ;
	wire _w7050_ ;
	wire _w7049_ ;
	wire _w7048_ ;
	wire _w7047_ ;
	wire _w7046_ ;
	wire _w7045_ ;
	wire _w7044_ ;
	wire _w7043_ ;
	wire _w7042_ ;
	wire _w7041_ ;
	wire _w7040_ ;
	wire _w7039_ ;
	wire _w7038_ ;
	wire _w7037_ ;
	wire _w7036_ ;
	wire _w7035_ ;
	wire _w7034_ ;
	wire _w7033_ ;
	wire _w7032_ ;
	wire _w7031_ ;
	wire _w7030_ ;
	wire _w7029_ ;
	wire _w7028_ ;
	wire _w7027_ ;
	wire _w7026_ ;
	wire _w7025_ ;
	wire _w7024_ ;
	wire _w7023_ ;
	wire _w7022_ ;
	wire _w7021_ ;
	wire _w7020_ ;
	wire _w7019_ ;
	wire _w7018_ ;
	wire _w7017_ ;
	wire _w7016_ ;
	wire _w7015_ ;
	wire _w7014_ ;
	wire _w7013_ ;
	wire _w7012_ ;
	wire _w7011_ ;
	wire _w7010_ ;
	wire _w7009_ ;
	wire _w7008_ ;
	wire _w7007_ ;
	wire _w7006_ ;
	wire _w7005_ ;
	wire _w7004_ ;
	wire _w7003_ ;
	wire _w7002_ ;
	wire _w7001_ ;
	wire _w7000_ ;
	wire _w6999_ ;
	wire _w6998_ ;
	wire _w6997_ ;
	wire _w6996_ ;
	wire _w6995_ ;
	wire _w6994_ ;
	wire _w6993_ ;
	wire _w6992_ ;
	wire _w6991_ ;
	wire _w6990_ ;
	wire _w6989_ ;
	wire _w6988_ ;
	wire _w6987_ ;
	wire _w6986_ ;
	wire _w6985_ ;
	wire _w6984_ ;
	wire _w6983_ ;
	wire _w6982_ ;
	wire _w6981_ ;
	wire _w6980_ ;
	wire _w6979_ ;
	wire _w6978_ ;
	wire _w6977_ ;
	wire _w6976_ ;
	wire _w6975_ ;
	wire _w6974_ ;
	wire _w6973_ ;
	wire _w6972_ ;
	wire _w6971_ ;
	wire _w6970_ ;
	wire _w6969_ ;
	wire _w6968_ ;
	wire _w6967_ ;
	wire _w6966_ ;
	wire _w6965_ ;
	wire _w6964_ ;
	wire _w6963_ ;
	wire _w6962_ ;
	wire _w6961_ ;
	wire _w6960_ ;
	wire _w6959_ ;
	wire _w6958_ ;
	wire _w6957_ ;
	wire _w6956_ ;
	wire _w6955_ ;
	wire _w6954_ ;
	wire _w6953_ ;
	wire _w6952_ ;
	wire _w6951_ ;
	wire _w6950_ ;
	wire _w6949_ ;
	wire _w6948_ ;
	wire _w6947_ ;
	wire _w6946_ ;
	wire _w6945_ ;
	wire _w6944_ ;
	wire _w6943_ ;
	wire _w6942_ ;
	wire _w6941_ ;
	wire _w6940_ ;
	wire _w6939_ ;
	wire _w6938_ ;
	wire _w6937_ ;
	wire _w6936_ ;
	wire _w6935_ ;
	wire _w6934_ ;
	wire _w6933_ ;
	wire _w6932_ ;
	wire _w6931_ ;
	wire _w6930_ ;
	wire _w6929_ ;
	wire _w6928_ ;
	wire _w6927_ ;
	wire _w6926_ ;
	wire _w6925_ ;
	wire _w6924_ ;
	wire _w6923_ ;
	wire _w6922_ ;
	wire _w6921_ ;
	wire _w6920_ ;
	wire _w6919_ ;
	wire _w6918_ ;
	wire _w6917_ ;
	wire _w6916_ ;
	wire _w6915_ ;
	wire _w6914_ ;
	wire _w6913_ ;
	wire _w6912_ ;
	wire _w6911_ ;
	wire _w6910_ ;
	wire _w6909_ ;
	wire _w6908_ ;
	wire _w6907_ ;
	wire _w6906_ ;
	wire _w6905_ ;
	wire _w6904_ ;
	wire _w6903_ ;
	wire _w6902_ ;
	wire _w6901_ ;
	wire _w6900_ ;
	wire _w6899_ ;
	wire _w6898_ ;
	wire _w6897_ ;
	wire _w6896_ ;
	wire _w6895_ ;
	wire _w6894_ ;
	wire _w6893_ ;
	wire _w6892_ ;
	wire _w6891_ ;
	wire _w6890_ ;
	wire _w6889_ ;
	wire _w6888_ ;
	wire _w6887_ ;
	wire _w6886_ ;
	wire _w6885_ ;
	wire _w6884_ ;
	wire _w6883_ ;
	wire _w6882_ ;
	wire _w6881_ ;
	wire _w6880_ ;
	wire _w6879_ ;
	wire _w6878_ ;
	wire _w6877_ ;
	wire _w6876_ ;
	wire _w6875_ ;
	wire _w6874_ ;
	wire _w6873_ ;
	wire _w6872_ ;
	wire _w6871_ ;
	wire _w6870_ ;
	wire _w6869_ ;
	wire _w6868_ ;
	wire _w6867_ ;
	wire _w6866_ ;
	wire _w6865_ ;
	wire _w6864_ ;
	wire _w6863_ ;
	wire _w6862_ ;
	wire _w6861_ ;
	wire _w6860_ ;
	wire _w6859_ ;
	wire _w6858_ ;
	wire _w6857_ ;
	wire _w6856_ ;
	wire _w6855_ ;
	wire _w6854_ ;
	wire _w6853_ ;
	wire _w6852_ ;
	wire _w6851_ ;
	wire _w6850_ ;
	wire _w6849_ ;
	wire _w6848_ ;
	wire _w6847_ ;
	wire _w6846_ ;
	wire _w6845_ ;
	wire _w6844_ ;
	wire _w6843_ ;
	wire _w6842_ ;
	wire _w6841_ ;
	wire _w6840_ ;
	wire _w6839_ ;
	wire _w6838_ ;
	wire _w6837_ ;
	wire _w6836_ ;
	wire _w6835_ ;
	wire _w6834_ ;
	wire _w6833_ ;
	wire _w6832_ ;
	wire _w6831_ ;
	wire _w6830_ ;
	wire _w6829_ ;
	wire _w6828_ ;
	wire _w6827_ ;
	wire _w6826_ ;
	wire _w6825_ ;
	wire _w6824_ ;
	wire _w6823_ ;
	wire _w6822_ ;
	wire _w6821_ ;
	wire _w6820_ ;
	wire _w6819_ ;
	wire _w6818_ ;
	wire _w6817_ ;
	wire _w6816_ ;
	wire _w6815_ ;
	wire _w6814_ ;
	wire _w6813_ ;
	wire _w6812_ ;
	wire _w6811_ ;
	wire _w6810_ ;
	wire _w6809_ ;
	wire _w6808_ ;
	wire _w6807_ ;
	wire _w6806_ ;
	wire _w6805_ ;
	wire _w6804_ ;
	wire _w6803_ ;
	wire _w6802_ ;
	wire _w6801_ ;
	wire _w6800_ ;
	wire _w6799_ ;
	wire _w6798_ ;
	wire _w6797_ ;
	wire _w6796_ ;
	wire _w6795_ ;
	wire _w6794_ ;
	wire _w6793_ ;
	wire _w6792_ ;
	wire _w6791_ ;
	wire _w6790_ ;
	wire _w6789_ ;
	wire _w6788_ ;
	wire _w6787_ ;
	wire _w6786_ ;
	wire _w6785_ ;
	wire _w6784_ ;
	wire _w6783_ ;
	wire _w6782_ ;
	wire _w6781_ ;
	wire _w6780_ ;
	wire _w6779_ ;
	wire _w6778_ ;
	wire _w6777_ ;
	wire _w6776_ ;
	wire _w6775_ ;
	wire _w6774_ ;
	wire _w6773_ ;
	wire _w6772_ ;
	wire _w6771_ ;
	wire _w6770_ ;
	wire _w6769_ ;
	wire _w6768_ ;
	wire _w6767_ ;
	wire _w6766_ ;
	wire _w6765_ ;
	wire _w6764_ ;
	wire _w6763_ ;
	wire _w6762_ ;
	wire _w6761_ ;
	wire _w6760_ ;
	wire _w6759_ ;
	wire _w6758_ ;
	wire _w6757_ ;
	wire _w6756_ ;
	wire _w6755_ ;
	wire _w6754_ ;
	wire _w6753_ ;
	wire _w6752_ ;
	wire _w6751_ ;
	wire _w6750_ ;
	wire _w6749_ ;
	wire _w6748_ ;
	wire _w6747_ ;
	wire _w6746_ ;
	wire _w6745_ ;
	wire _w6744_ ;
	wire _w6743_ ;
	wire _w6742_ ;
	wire _w6741_ ;
	wire _w6740_ ;
	wire _w6739_ ;
	wire _w6738_ ;
	wire _w6737_ ;
	wire _w6736_ ;
	wire _w6735_ ;
	wire _w6734_ ;
	wire _w6733_ ;
	wire _w6732_ ;
	wire _w6731_ ;
	wire _w6730_ ;
	wire _w6729_ ;
	wire _w6728_ ;
	wire _w6727_ ;
	wire _w6726_ ;
	wire _w6725_ ;
	wire _w6724_ ;
	wire _w6723_ ;
	wire _w6722_ ;
	wire _w6721_ ;
	wire _w6720_ ;
	wire _w6719_ ;
	wire _w6718_ ;
	wire _w6717_ ;
	wire _w6716_ ;
	wire _w6715_ ;
	wire _w6714_ ;
	wire _w6713_ ;
	wire _w6712_ ;
	wire _w6711_ ;
	wire _w6710_ ;
	wire _w6709_ ;
	wire _w6708_ ;
	wire _w6707_ ;
	wire _w6706_ ;
	wire _w6705_ ;
	wire _w6704_ ;
	wire _w6703_ ;
	wire _w6702_ ;
	wire _w6701_ ;
	wire _w6700_ ;
	wire _w6699_ ;
	wire _w6698_ ;
	wire _w6697_ ;
	wire _w6696_ ;
	wire _w6695_ ;
	wire _w6694_ ;
	wire _w6693_ ;
	wire _w6692_ ;
	wire _w6691_ ;
	wire _w6690_ ;
	wire _w6689_ ;
	wire _w6688_ ;
	wire _w6687_ ;
	wire _w6686_ ;
	wire _w6685_ ;
	wire _w6684_ ;
	wire _w6683_ ;
	wire _w6682_ ;
	wire _w6681_ ;
	wire _w6680_ ;
	wire _w6679_ ;
	wire _w6678_ ;
	wire _w6677_ ;
	wire _w6676_ ;
	wire _w6675_ ;
	wire _w6674_ ;
	wire _w6673_ ;
	wire _w6672_ ;
	wire _w6671_ ;
	wire _w6670_ ;
	wire _w6669_ ;
	wire _w6668_ ;
	wire _w6667_ ;
	wire _w6666_ ;
	wire _w6665_ ;
	wire _w6664_ ;
	wire _w6663_ ;
	wire _w6662_ ;
	wire _w6661_ ;
	wire _w6660_ ;
	wire _w6659_ ;
	wire _w6658_ ;
	wire _w6657_ ;
	wire _w6656_ ;
	wire _w6655_ ;
	wire _w6654_ ;
	wire _w6653_ ;
	wire _w6652_ ;
	wire _w6651_ ;
	wire _w6650_ ;
	wire _w6649_ ;
	wire _w6648_ ;
	wire _w6647_ ;
	wire _w6646_ ;
	wire _w6645_ ;
	wire _w6644_ ;
	wire _w6643_ ;
	wire _w6642_ ;
	wire _w6641_ ;
	wire _w6640_ ;
	wire _w6639_ ;
	wire _w6638_ ;
	wire _w6637_ ;
	wire _w6636_ ;
	wire _w6635_ ;
	wire _w6634_ ;
	wire _w6633_ ;
	wire _w6632_ ;
	wire _w6631_ ;
	wire _w6630_ ;
	wire _w6629_ ;
	wire _w6628_ ;
	wire _w6627_ ;
	wire _w6626_ ;
	wire _w6625_ ;
	wire _w6624_ ;
	wire _w6623_ ;
	wire _w6622_ ;
	wire _w6621_ ;
	wire _w6620_ ;
	wire _w6619_ ;
	wire _w6618_ ;
	wire _w6617_ ;
	wire _w6616_ ;
	wire _w6615_ ;
	wire _w6614_ ;
	wire _w6613_ ;
	wire _w6612_ ;
	wire _w6611_ ;
	wire _w6610_ ;
	wire _w6609_ ;
	wire _w6608_ ;
	wire _w6607_ ;
	wire _w6606_ ;
	wire _w6605_ ;
	wire _w6604_ ;
	wire _w6603_ ;
	wire _w6602_ ;
	wire _w6601_ ;
	wire _w6600_ ;
	wire _w6599_ ;
	wire _w6598_ ;
	wire _w6597_ ;
	wire _w6596_ ;
	wire _w6595_ ;
	wire _w6594_ ;
	wire _w6593_ ;
	wire _w6592_ ;
	wire _w6591_ ;
	wire _w6590_ ;
	wire _w6589_ ;
	wire _w6588_ ;
	wire _w6587_ ;
	wire _w6586_ ;
	wire _w6585_ ;
	wire _w6584_ ;
	wire _w6583_ ;
	wire _w6582_ ;
	wire _w6581_ ;
	wire _w6580_ ;
	wire _w6579_ ;
	wire _w6578_ ;
	wire _w6577_ ;
	wire _w6576_ ;
	wire _w6575_ ;
	wire _w6574_ ;
	wire _w6573_ ;
	wire _w6572_ ;
	wire _w6571_ ;
	wire _w6570_ ;
	wire _w6569_ ;
	wire _w6568_ ;
	wire _w6567_ ;
	wire _w6566_ ;
	wire _w6565_ ;
	wire _w6564_ ;
	wire _w6563_ ;
	wire _w6562_ ;
	wire _w6561_ ;
	wire _w6560_ ;
	wire _w6559_ ;
	wire _w6558_ ;
	wire _w6557_ ;
	wire _w6556_ ;
	wire _w6555_ ;
	wire _w6554_ ;
	wire _w6553_ ;
	wire _w6552_ ;
	wire _w6551_ ;
	wire _w6550_ ;
	wire _w6549_ ;
	wire _w6548_ ;
	wire _w6547_ ;
	wire _w6546_ ;
	wire _w6545_ ;
	wire _w6544_ ;
	wire _w6543_ ;
	wire _w6542_ ;
	wire _w6541_ ;
	wire _w6540_ ;
	wire _w6539_ ;
	wire _w6538_ ;
	wire _w6537_ ;
	wire _w6536_ ;
	wire _w6535_ ;
	wire _w6534_ ;
	wire _w6533_ ;
	wire _w6532_ ;
	wire _w6531_ ;
	wire _w6530_ ;
	wire _w6529_ ;
	wire _w6528_ ;
	wire _w6527_ ;
	wire _w6526_ ;
	wire _w6525_ ;
	wire _w6524_ ;
	wire _w6523_ ;
	wire _w6522_ ;
	wire _w6521_ ;
	wire _w6520_ ;
	wire _w6519_ ;
	wire _w6518_ ;
	wire _w6517_ ;
	wire _w6516_ ;
	wire _w6515_ ;
	wire _w6514_ ;
	wire _w6513_ ;
	wire _w6512_ ;
	wire _w6511_ ;
	wire _w6510_ ;
	wire _w6509_ ;
	wire _w6508_ ;
	wire _w6507_ ;
	wire _w6506_ ;
	wire _w6505_ ;
	wire _w6504_ ;
	wire _w6503_ ;
	wire _w6502_ ;
	wire _w6501_ ;
	wire _w6500_ ;
	wire _w6499_ ;
	wire _w6498_ ;
	wire _w6497_ ;
	wire _w6496_ ;
	wire _w6495_ ;
	wire _w6494_ ;
	wire _w6493_ ;
	wire _w6492_ ;
	wire _w6491_ ;
	wire _w6490_ ;
	wire _w6489_ ;
	wire _w6488_ ;
	wire _w6487_ ;
	wire _w6486_ ;
	wire _w6485_ ;
	wire _w6484_ ;
	wire _w6483_ ;
	wire _w6482_ ;
	wire _w6481_ ;
	wire _w6480_ ;
	wire _w6479_ ;
	wire _w6478_ ;
	wire _w6477_ ;
	wire _w6476_ ;
	wire _w6475_ ;
	wire _w6474_ ;
	wire _w6473_ ;
	wire _w6472_ ;
	wire _w6471_ ;
	wire _w6470_ ;
	wire _w6469_ ;
	wire _w6468_ ;
	wire _w6467_ ;
	wire _w6466_ ;
	wire _w6465_ ;
	wire _w6464_ ;
	wire _w6463_ ;
	wire _w6462_ ;
	wire _w6461_ ;
	wire _w6460_ ;
	wire _w6459_ ;
	wire _w6458_ ;
	wire _w6457_ ;
	wire _w6456_ ;
	wire _w6455_ ;
	wire _w6454_ ;
	wire _w6453_ ;
	wire _w6452_ ;
	wire _w6451_ ;
	wire _w6450_ ;
	wire _w6449_ ;
	wire _w6448_ ;
	wire _w6447_ ;
	wire _w6446_ ;
	wire _w6445_ ;
	wire _w6444_ ;
	wire _w6443_ ;
	wire _w6442_ ;
	wire _w6441_ ;
	wire _w6440_ ;
	wire _w6439_ ;
	wire _w6438_ ;
	wire _w6437_ ;
	wire _w6436_ ;
	wire _w6435_ ;
	wire _w6434_ ;
	wire _w6433_ ;
	wire _w6432_ ;
	wire _w6431_ ;
	wire _w6430_ ;
	wire _w6429_ ;
	wire _w6428_ ;
	wire _w6427_ ;
	wire _w6426_ ;
	wire _w6425_ ;
	wire _w6424_ ;
	wire _w6423_ ;
	wire _w6422_ ;
	wire _w6421_ ;
	wire _w6420_ ;
	wire _w6419_ ;
	wire _w6418_ ;
	wire _w6417_ ;
	wire _w6416_ ;
	wire _w6415_ ;
	wire _w6414_ ;
	wire _w6413_ ;
	wire _w6412_ ;
	wire _w6411_ ;
	wire _w6410_ ;
	wire _w6409_ ;
	wire _w6408_ ;
	wire _w6407_ ;
	wire _w6406_ ;
	wire _w6405_ ;
	wire _w6404_ ;
	wire _w6403_ ;
	wire _w6402_ ;
	wire _w6401_ ;
	wire _w6400_ ;
	wire _w6399_ ;
	wire _w6398_ ;
	wire _w6397_ ;
	wire _w6396_ ;
	wire _w6395_ ;
	wire _w6394_ ;
	wire _w6393_ ;
	wire _w6392_ ;
	wire _w6391_ ;
	wire _w6390_ ;
	wire _w6389_ ;
	wire _w6388_ ;
	wire _w6387_ ;
	wire _w6386_ ;
	wire _w6385_ ;
	wire _w6384_ ;
	wire _w6383_ ;
	wire _w6382_ ;
	wire _w6381_ ;
	wire _w6380_ ;
	wire _w6379_ ;
	wire _w6378_ ;
	wire _w6377_ ;
	wire _w6376_ ;
	wire _w6375_ ;
	wire _w6374_ ;
	wire _w6373_ ;
	wire _w6372_ ;
	wire _w6371_ ;
	wire _w6370_ ;
	wire _w6369_ ;
	wire _w6368_ ;
	wire _w6367_ ;
	wire _w6366_ ;
	wire _w6365_ ;
	wire _w6364_ ;
	wire _w6363_ ;
	wire _w6362_ ;
	wire _w6361_ ;
	wire _w6360_ ;
	wire _w6359_ ;
	wire _w6358_ ;
	wire _w6357_ ;
	wire _w6356_ ;
	wire _w6355_ ;
	wire _w6354_ ;
	wire _w6353_ ;
	wire _w6352_ ;
	wire _w6351_ ;
	wire _w6350_ ;
	wire _w6349_ ;
	wire _w6348_ ;
	wire _w6347_ ;
	wire _w6346_ ;
	wire _w6345_ ;
	wire _w6344_ ;
	wire _w6343_ ;
	wire _w6342_ ;
	wire _w6341_ ;
	wire _w6340_ ;
	wire _w6339_ ;
	wire _w6338_ ;
	wire _w6337_ ;
	wire _w6336_ ;
	wire _w6335_ ;
	wire _w6334_ ;
	wire _w6333_ ;
	wire _w6332_ ;
	wire _w6331_ ;
	wire _w6330_ ;
	wire _w6329_ ;
	wire _w6328_ ;
	wire _w6327_ ;
	wire _w6326_ ;
	wire _w6325_ ;
	wire _w6324_ ;
	wire _w6323_ ;
	wire _w6322_ ;
	wire _w6321_ ;
	wire _w6320_ ;
	wire _w6319_ ;
	wire _w6318_ ;
	wire _w6317_ ;
	wire _w6316_ ;
	wire _w6315_ ;
	wire _w6314_ ;
	wire _w6313_ ;
	wire _w6312_ ;
	wire _w6311_ ;
	wire _w6310_ ;
	wire _w6309_ ;
	wire _w6308_ ;
	wire _w6307_ ;
	wire _w6306_ ;
	wire _w6305_ ;
	wire _w6304_ ;
	wire _w6303_ ;
	wire _w6302_ ;
	wire _w6301_ ;
	wire _w6300_ ;
	wire _w6299_ ;
	wire _w6298_ ;
	wire _w6297_ ;
	wire _w6296_ ;
	wire _w6295_ ;
	wire _w6294_ ;
	wire _w6293_ ;
	wire _w6292_ ;
	wire _w6291_ ;
	wire _w6290_ ;
	wire _w6289_ ;
	wire _w6288_ ;
	wire _w6287_ ;
	wire _w6286_ ;
	wire _w6285_ ;
	wire _w6284_ ;
	wire _w6283_ ;
	wire _w6282_ ;
	wire _w6281_ ;
	wire _w6280_ ;
	wire _w6279_ ;
	wire _w6278_ ;
	wire _w6277_ ;
	wire _w6276_ ;
	wire _w6275_ ;
	wire _w6274_ ;
	wire _w6273_ ;
	wire _w6272_ ;
	wire _w6271_ ;
	wire _w6270_ ;
	wire _w6269_ ;
	wire _w6268_ ;
	wire _w6267_ ;
	wire _w6266_ ;
	wire _w6265_ ;
	wire _w6264_ ;
	wire _w6263_ ;
	wire _w6262_ ;
	wire _w6261_ ;
	wire _w6260_ ;
	wire _w6259_ ;
	wire _w6258_ ;
	wire _w6257_ ;
	wire _w6256_ ;
	wire _w6255_ ;
	wire _w6254_ ;
	wire _w6253_ ;
	wire _w6252_ ;
	wire _w6251_ ;
	wire _w6250_ ;
	wire _w6249_ ;
	wire _w6248_ ;
	wire _w6247_ ;
	wire _w6246_ ;
	wire _w6245_ ;
	wire _w6244_ ;
	wire _w6243_ ;
	wire _w6242_ ;
	wire _w6241_ ;
	wire _w6240_ ;
	wire _w6239_ ;
	wire _w6238_ ;
	wire _w6237_ ;
	wire _w6236_ ;
	wire _w6235_ ;
	wire _w6234_ ;
	wire _w6233_ ;
	wire _w6232_ ;
	wire _w6231_ ;
	wire _w6230_ ;
	wire _w6229_ ;
	wire _w6228_ ;
	wire _w6227_ ;
	wire _w6226_ ;
	wire _w6225_ ;
	wire _w6224_ ;
	wire _w6223_ ;
	wire _w6222_ ;
	wire _w6221_ ;
	wire _w6220_ ;
	wire _w6219_ ;
	wire _w6218_ ;
	wire _w6217_ ;
	wire _w6216_ ;
	wire _w6215_ ;
	wire _w6214_ ;
	wire _w6213_ ;
	wire _w6212_ ;
	wire _w6211_ ;
	wire _w6210_ ;
	wire _w6209_ ;
	wire _w6208_ ;
	wire _w6207_ ;
	wire _w6206_ ;
	wire _w6205_ ;
	wire _w6204_ ;
	wire _w6203_ ;
	wire _w6202_ ;
	wire _w6201_ ;
	wire _w6200_ ;
	wire _w6199_ ;
	wire _w6198_ ;
	wire _w6197_ ;
	wire _w6196_ ;
	wire _w6195_ ;
	wire _w6194_ ;
	wire _w6193_ ;
	wire _w6192_ ;
	wire _w6191_ ;
	wire _w6190_ ;
	wire _w6189_ ;
	wire _w6188_ ;
	wire _w6187_ ;
	wire _w6186_ ;
	wire _w6185_ ;
	wire _w6184_ ;
	wire _w6183_ ;
	wire _w6182_ ;
	wire _w6181_ ;
	wire _w6180_ ;
	wire _w6179_ ;
	wire _w6178_ ;
	wire _w6177_ ;
	wire _w6176_ ;
	wire _w6175_ ;
	wire _w6174_ ;
	wire _w6173_ ;
	wire _w6172_ ;
	wire _w6171_ ;
	wire _w6170_ ;
	wire _w6169_ ;
	wire _w6168_ ;
	wire _w6167_ ;
	wire _w6166_ ;
	wire _w6165_ ;
	wire _w6164_ ;
	wire _w6163_ ;
	wire _w6162_ ;
	wire _w6161_ ;
	wire _w6160_ ;
	wire _w6159_ ;
	wire _w6158_ ;
	wire _w6157_ ;
	wire _w6156_ ;
	wire _w6155_ ;
	wire _w6154_ ;
	wire _w6153_ ;
	wire _w6152_ ;
	wire _w6151_ ;
	wire _w6150_ ;
	wire _w6149_ ;
	wire _w6148_ ;
	wire _w6147_ ;
	wire _w6146_ ;
	wire _w6145_ ;
	wire _w6144_ ;
	wire _w6143_ ;
	wire _w6142_ ;
	wire _w6141_ ;
	wire _w6140_ ;
	wire _w6139_ ;
	wire _w6138_ ;
	wire _w6137_ ;
	wire _w6136_ ;
	wire _w6135_ ;
	wire _w6134_ ;
	wire _w6133_ ;
	wire _w6132_ ;
	wire _w6131_ ;
	wire _w6130_ ;
	wire _w6129_ ;
	wire _w6128_ ;
	wire _w6127_ ;
	wire _w6126_ ;
	wire _w6125_ ;
	wire _w6124_ ;
	wire _w6123_ ;
	wire _w6122_ ;
	wire _w6121_ ;
	wire _w6120_ ;
	wire _w6119_ ;
	wire _w6118_ ;
	wire _w6117_ ;
	wire _w6116_ ;
	wire _w6115_ ;
	wire _w6114_ ;
	wire _w6113_ ;
	wire _w6112_ ;
	wire _w6111_ ;
	wire _w6110_ ;
	wire _w6109_ ;
	wire _w6108_ ;
	wire _w6107_ ;
	wire _w6106_ ;
	wire _w6105_ ;
	wire _w6104_ ;
	wire _w6103_ ;
	wire _w6102_ ;
	wire _w6101_ ;
	wire _w6100_ ;
	wire _w6099_ ;
	wire _w6098_ ;
	wire _w6097_ ;
	wire _w6096_ ;
	wire _w6095_ ;
	wire _w6094_ ;
	wire _w6093_ ;
	wire _w6092_ ;
	wire _w6091_ ;
	wire _w6090_ ;
	wire _w6089_ ;
	wire _w6088_ ;
	wire _w6087_ ;
	wire _w6086_ ;
	wire _w6085_ ;
	wire _w6084_ ;
	wire _w6083_ ;
	wire _w6082_ ;
	wire _w6081_ ;
	wire _w6080_ ;
	wire _w6079_ ;
	wire _w6078_ ;
	wire _w6077_ ;
	wire _w6076_ ;
	wire _w6075_ ;
	wire _w6074_ ;
	wire _w6073_ ;
	wire _w6072_ ;
	wire _w6071_ ;
	wire _w6070_ ;
	wire _w6069_ ;
	wire _w6068_ ;
	wire _w6067_ ;
	wire _w6066_ ;
	wire _w6065_ ;
	wire _w6064_ ;
	wire _w6063_ ;
	wire _w6062_ ;
	wire _w6061_ ;
	wire _w6060_ ;
	wire _w6059_ ;
	wire _w6058_ ;
	wire _w6057_ ;
	wire _w6056_ ;
	wire _w6055_ ;
	wire _w6054_ ;
	wire _w6053_ ;
	wire _w6052_ ;
	wire _w6051_ ;
	wire _w6050_ ;
	wire _w6049_ ;
	wire _w6048_ ;
	wire _w6047_ ;
	wire _w6046_ ;
	wire _w6045_ ;
	wire _w6044_ ;
	wire _w6043_ ;
	wire _w6042_ ;
	wire _w6041_ ;
	wire _w6040_ ;
	wire _w6039_ ;
	wire _w6038_ ;
	wire _w6037_ ;
	wire _w6036_ ;
	wire _w6035_ ;
	wire _w6034_ ;
	wire _w6033_ ;
	wire _w6032_ ;
	wire _w6031_ ;
	wire _w6030_ ;
	wire _w6029_ ;
	wire _w6028_ ;
	wire _w6027_ ;
	wire _w6026_ ;
	wire _w6025_ ;
	wire _w6024_ ;
	wire _w6023_ ;
	wire _w6022_ ;
	wire _w6021_ ;
	wire _w6020_ ;
	wire _w6019_ ;
	wire _w6018_ ;
	wire _w6017_ ;
	wire _w6016_ ;
	wire _w6015_ ;
	wire _w6014_ ;
	wire _w6013_ ;
	wire _w6012_ ;
	wire _w6011_ ;
	wire _w6010_ ;
	wire _w6009_ ;
	wire _w6008_ ;
	wire _w6007_ ;
	wire _w6006_ ;
	wire _w6005_ ;
	wire _w6004_ ;
	wire _w6003_ ;
	wire _w6002_ ;
	wire _w6001_ ;
	wire _w6000_ ;
	wire _w5999_ ;
	wire _w5998_ ;
	wire _w5997_ ;
	wire _w5996_ ;
	wire _w5995_ ;
	wire _w5994_ ;
	wire _w5993_ ;
	wire _w5992_ ;
	wire _w5991_ ;
	wire _w5990_ ;
	wire _w5989_ ;
	wire _w5988_ ;
	wire _w5987_ ;
	wire _w5986_ ;
	wire _w5985_ ;
	wire _w5984_ ;
	wire _w5983_ ;
	wire _w5982_ ;
	wire _w5981_ ;
	wire _w5980_ ;
	wire _w5979_ ;
	wire _w5978_ ;
	wire _w5977_ ;
	wire _w5976_ ;
	wire _w5975_ ;
	wire _w5974_ ;
	wire _w5973_ ;
	wire _w5972_ ;
	wire _w5971_ ;
	wire _w5970_ ;
	wire _w5969_ ;
	wire _w5968_ ;
	wire _w5967_ ;
	wire _w5966_ ;
	wire _w5965_ ;
	wire _w5964_ ;
	wire _w5963_ ;
	wire _w5962_ ;
	wire _w5961_ ;
	wire _w5960_ ;
	wire _w5959_ ;
	wire _w5958_ ;
	wire _w5957_ ;
	wire _w5956_ ;
	wire _w5955_ ;
	wire _w5954_ ;
	wire _w5953_ ;
	wire _w5952_ ;
	wire _w5951_ ;
	wire _w5950_ ;
	wire _w5949_ ;
	wire _w5948_ ;
	wire _w5947_ ;
	wire _w5946_ ;
	wire _w5945_ ;
	wire _w5944_ ;
	wire _w5943_ ;
	wire _w5942_ ;
	wire _w5941_ ;
	wire _w5940_ ;
	wire _w5939_ ;
	wire _w5938_ ;
	wire _w5937_ ;
	wire _w5936_ ;
	wire _w5935_ ;
	wire _w5934_ ;
	wire _w5933_ ;
	wire _w5932_ ;
	wire _w5931_ ;
	wire _w5930_ ;
	wire _w5929_ ;
	wire _w5928_ ;
	wire _w5927_ ;
	wire _w5926_ ;
	wire _w5925_ ;
	wire _w5924_ ;
	wire _w5923_ ;
	wire _w5922_ ;
	wire _w5921_ ;
	wire _w5920_ ;
	wire _w5919_ ;
	wire _w5918_ ;
	wire _w5917_ ;
	wire _w5916_ ;
	wire _w5915_ ;
	wire _w5914_ ;
	wire _w5913_ ;
	wire _w5912_ ;
	wire _w5911_ ;
	wire _w5910_ ;
	wire _w5909_ ;
	wire _w5908_ ;
	wire _w5907_ ;
	wire _w5906_ ;
	wire _w5905_ ;
	wire _w5904_ ;
	wire _w5903_ ;
	wire _w5902_ ;
	wire _w5901_ ;
	wire _w5900_ ;
	wire _w5899_ ;
	wire _w5898_ ;
	wire _w5897_ ;
	wire _w5896_ ;
	wire _w5895_ ;
	wire _w5894_ ;
	wire _w5893_ ;
	wire _w5892_ ;
	wire _w5891_ ;
	wire _w5890_ ;
	wire _w5889_ ;
	wire _w5888_ ;
	wire _w5887_ ;
	wire _w5886_ ;
	wire _w5885_ ;
	wire _w5884_ ;
	wire _w5883_ ;
	wire _w5882_ ;
	wire _w5881_ ;
	wire _w5880_ ;
	wire _w5879_ ;
	wire _w5878_ ;
	wire _w5877_ ;
	wire _w5876_ ;
	wire _w5875_ ;
	wire _w5874_ ;
	wire _w5873_ ;
	wire _w5872_ ;
	wire _w5871_ ;
	wire _w5870_ ;
	wire _w5869_ ;
	wire _w5868_ ;
	wire _w5867_ ;
	wire _w5866_ ;
	wire _w5865_ ;
	wire _w5864_ ;
	wire _w5863_ ;
	wire _w5862_ ;
	wire _w5861_ ;
	wire _w5860_ ;
	wire _w5859_ ;
	wire _w5858_ ;
	wire _w5857_ ;
	wire _w5856_ ;
	wire _w5855_ ;
	wire _w5854_ ;
	wire _w5853_ ;
	wire _w5852_ ;
	wire _w5851_ ;
	wire _w5850_ ;
	wire _w5849_ ;
	wire _w5848_ ;
	wire _w5847_ ;
	wire _w5846_ ;
	wire _w5845_ ;
	wire _w5844_ ;
	wire _w5843_ ;
	wire _w5842_ ;
	wire _w5841_ ;
	wire _w5840_ ;
	wire _w5839_ ;
	wire _w5838_ ;
	wire _w5837_ ;
	wire _w5836_ ;
	wire _w5835_ ;
	wire _w5834_ ;
	wire _w5833_ ;
	wire _w5832_ ;
	wire _w5831_ ;
	wire _w5830_ ;
	wire _w5829_ ;
	wire _w5828_ ;
	wire _w5827_ ;
	wire _w5826_ ;
	wire _w5825_ ;
	wire _w5824_ ;
	wire _w5823_ ;
	wire _w5822_ ;
	wire _w5821_ ;
	wire _w5820_ ;
	wire _w5819_ ;
	wire _w5818_ ;
	wire _w5817_ ;
	wire _w5816_ ;
	wire _w5815_ ;
	wire _w5814_ ;
	wire _w5813_ ;
	wire _w5812_ ;
	wire _w5811_ ;
	wire _w5810_ ;
	wire _w5809_ ;
	wire _w5808_ ;
	wire _w5807_ ;
	wire _w5806_ ;
	wire _w5805_ ;
	wire _w5804_ ;
	wire _w5803_ ;
	wire _w5802_ ;
	wire _w5801_ ;
	wire _w5800_ ;
	wire _w5799_ ;
	wire _w5798_ ;
	wire _w5797_ ;
	wire _w5796_ ;
	wire _w5795_ ;
	wire _w5794_ ;
	wire _w5793_ ;
	wire _w5792_ ;
	wire _w5791_ ;
	wire _w5790_ ;
	wire _w5789_ ;
	wire _w5788_ ;
	wire _w5787_ ;
	wire _w5786_ ;
	wire _w5785_ ;
	wire _w5784_ ;
	wire _w5783_ ;
	wire _w5782_ ;
	wire _w5781_ ;
	wire _w5780_ ;
	wire _w5779_ ;
	wire _w5778_ ;
	wire _w5777_ ;
	wire _w5776_ ;
	wire _w5775_ ;
	wire _w5774_ ;
	wire _w5773_ ;
	wire _w5772_ ;
	wire _w5771_ ;
	wire _w5770_ ;
	wire _w5769_ ;
	wire _w5768_ ;
	wire _w5767_ ;
	wire _w5766_ ;
	wire _w5765_ ;
	wire _w5764_ ;
	wire _w5763_ ;
	wire _w5762_ ;
	wire _w5761_ ;
	wire _w5760_ ;
	wire _w5759_ ;
	wire _w5758_ ;
	wire _w5757_ ;
	wire _w5756_ ;
	wire _w5755_ ;
	wire _w5754_ ;
	wire _w5753_ ;
	wire _w5752_ ;
	wire _w5751_ ;
	wire _w5750_ ;
	wire _w5749_ ;
	wire _w5748_ ;
	wire _w5747_ ;
	wire _w5746_ ;
	wire _w5745_ ;
	wire _w5744_ ;
	wire _w5743_ ;
	wire _w5742_ ;
	wire _w5741_ ;
	wire _w5740_ ;
	wire _w5739_ ;
	wire _w5738_ ;
	wire _w5737_ ;
	wire _w5736_ ;
	wire _w5735_ ;
	wire _w5734_ ;
	wire _w5733_ ;
	wire _w5732_ ;
	wire _w5731_ ;
	wire _w5730_ ;
	wire _w5729_ ;
	wire _w5728_ ;
	wire _w5727_ ;
	wire _w5726_ ;
	wire _w5725_ ;
	wire _w5724_ ;
	wire _w5723_ ;
	wire _w5722_ ;
	wire _w5721_ ;
	wire _w5720_ ;
	wire _w5719_ ;
	wire _w5718_ ;
	wire _w5717_ ;
	wire _w5716_ ;
	wire _w5715_ ;
	wire _w5714_ ;
	wire _w5713_ ;
	wire _w5712_ ;
	wire _w5711_ ;
	wire _w5710_ ;
	wire _w5709_ ;
	wire _w5708_ ;
	wire _w5707_ ;
	wire _w5706_ ;
	wire _w5705_ ;
	wire _w5704_ ;
	wire _w5703_ ;
	wire _w5702_ ;
	wire _w5701_ ;
	wire _w5700_ ;
	wire _w5699_ ;
	wire _w5698_ ;
	wire _w5697_ ;
	wire _w5696_ ;
	wire _w5695_ ;
	wire _w5694_ ;
	wire _w5693_ ;
	wire _w5692_ ;
	wire _w5691_ ;
	wire _w5690_ ;
	wire _w5689_ ;
	wire _w5688_ ;
	wire _w5687_ ;
	wire _w5686_ ;
	wire _w5685_ ;
	wire _w5684_ ;
	wire _w5683_ ;
	wire _w5682_ ;
	wire _w5681_ ;
	wire _w5680_ ;
	wire _w5679_ ;
	wire _w5678_ ;
	wire _w5677_ ;
	wire _w5676_ ;
	wire _w5675_ ;
	wire _w5674_ ;
	wire _w5673_ ;
	wire _w5672_ ;
	wire _w5671_ ;
	wire _w5670_ ;
	wire _w5669_ ;
	wire _w5668_ ;
	wire _w5667_ ;
	wire _w5666_ ;
	wire _w5665_ ;
	wire _w5664_ ;
	wire _w5663_ ;
	wire _w5662_ ;
	wire _w5661_ ;
	wire _w5660_ ;
	wire _w5659_ ;
	wire _w5658_ ;
	wire _w5657_ ;
	wire _w5656_ ;
	wire _w5655_ ;
	wire _w5654_ ;
	wire _w5653_ ;
	wire _w5652_ ;
	wire _w5651_ ;
	wire _w5650_ ;
	wire _w5649_ ;
	wire _w5648_ ;
	wire _w5647_ ;
	wire _w5646_ ;
	wire _w5645_ ;
	wire _w5644_ ;
	wire _w5643_ ;
	wire _w5642_ ;
	wire _w5641_ ;
	wire _w5640_ ;
	wire _w5639_ ;
	wire _w5638_ ;
	wire _w5637_ ;
	wire _w5636_ ;
	wire _w5635_ ;
	wire _w5634_ ;
	wire _w5633_ ;
	wire _w5632_ ;
	wire _w5631_ ;
	wire _w5630_ ;
	wire _w5629_ ;
	wire _w5628_ ;
	wire _w5627_ ;
	wire _w5626_ ;
	wire _w5625_ ;
	wire _w5624_ ;
	wire _w5623_ ;
	wire _w5622_ ;
	wire _w5621_ ;
	wire _w5620_ ;
	wire _w5619_ ;
	wire _w5618_ ;
	wire _w5617_ ;
	wire _w5616_ ;
	wire _w5615_ ;
	wire _w5614_ ;
	wire _w5613_ ;
	wire _w5612_ ;
	wire _w5611_ ;
	wire _w5610_ ;
	wire _w5609_ ;
	wire _w5608_ ;
	wire _w5607_ ;
	wire _w5606_ ;
	wire _w5605_ ;
	wire _w5604_ ;
	wire _w5603_ ;
	wire _w5602_ ;
	wire _w5601_ ;
	wire _w5600_ ;
	wire _w5599_ ;
	wire _w5598_ ;
	wire _w5597_ ;
	wire _w5596_ ;
	wire _w5595_ ;
	wire _w5594_ ;
	wire _w5593_ ;
	wire _w5592_ ;
	wire _w5591_ ;
	wire _w5590_ ;
	wire _w5589_ ;
	wire _w5588_ ;
	wire _w5587_ ;
	wire _w5586_ ;
	wire _w5585_ ;
	wire _w5584_ ;
	wire _w5583_ ;
	wire _w5582_ ;
	wire _w5581_ ;
	wire _w5580_ ;
	wire _w5579_ ;
	wire _w5578_ ;
	wire _w5577_ ;
	wire _w5576_ ;
	wire _w5575_ ;
	wire _w5574_ ;
	wire _w5573_ ;
	wire _w5572_ ;
	wire _w5571_ ;
	wire _w5570_ ;
	wire _w5569_ ;
	wire _w5568_ ;
	wire _w5567_ ;
	wire _w5566_ ;
	wire _w5565_ ;
	wire _w5564_ ;
	wire _w5563_ ;
	wire _w5562_ ;
	wire _w5561_ ;
	wire _w5560_ ;
	wire _w5559_ ;
	wire _w5558_ ;
	wire _w5557_ ;
	wire _w5556_ ;
	wire _w5555_ ;
	wire _w5554_ ;
	wire _w5553_ ;
	wire _w5552_ ;
	wire _w5551_ ;
	wire _w5550_ ;
	wire _w5549_ ;
	wire _w5548_ ;
	wire _w5547_ ;
	wire _w5546_ ;
	wire _w5545_ ;
	wire _w5544_ ;
	wire _w5543_ ;
	wire _w5542_ ;
	wire _w5541_ ;
	wire _w5540_ ;
	wire _w5539_ ;
	wire _w5538_ ;
	wire _w5537_ ;
	wire _w5536_ ;
	wire _w5535_ ;
	wire _w5534_ ;
	wire _w5533_ ;
	wire _w5532_ ;
	wire _w5531_ ;
	wire _w5530_ ;
	wire _w5529_ ;
	wire _w5528_ ;
	wire _w5527_ ;
	wire _w5526_ ;
	wire _w5525_ ;
	wire _w5524_ ;
	wire _w5523_ ;
	wire _w5522_ ;
	wire _w5521_ ;
	wire _w5520_ ;
	wire _w5519_ ;
	wire _w5518_ ;
	wire _w5517_ ;
	wire _w5516_ ;
	wire _w5515_ ;
	wire _w5514_ ;
	wire _w5513_ ;
	wire _w5512_ ;
	wire _w5511_ ;
	wire _w5510_ ;
	wire _w5509_ ;
	wire _w5508_ ;
	wire _w5507_ ;
	wire _w5506_ ;
	wire _w5505_ ;
	wire _w5504_ ;
	wire _w5503_ ;
	wire _w5502_ ;
	wire _w5501_ ;
	wire _w5500_ ;
	wire _w5499_ ;
	wire _w5498_ ;
	wire _w5497_ ;
	wire _w5496_ ;
	wire _w5495_ ;
	wire _w5494_ ;
	wire _w5493_ ;
	wire _w5492_ ;
	wire _w5491_ ;
	wire _w5490_ ;
	wire _w5489_ ;
	wire _w5488_ ;
	wire _w5487_ ;
	wire _w5486_ ;
	wire _w5485_ ;
	wire _w5484_ ;
	wire _w5483_ ;
	wire _w5482_ ;
	wire _w5481_ ;
	wire _w5480_ ;
	wire _w5479_ ;
	wire _w5478_ ;
	wire _w5477_ ;
	wire _w5476_ ;
	wire _w5475_ ;
	wire _w5474_ ;
	wire _w5473_ ;
	wire _w5472_ ;
	wire _w5471_ ;
	wire _w5470_ ;
	wire _w5469_ ;
	wire _w5468_ ;
	wire _w5467_ ;
	wire _w5466_ ;
	wire _w5465_ ;
	wire _w5464_ ;
	wire _w5463_ ;
	wire _w5462_ ;
	wire _w5461_ ;
	wire _w5460_ ;
	wire _w5459_ ;
	wire _w5458_ ;
	wire _w5457_ ;
	wire _w5456_ ;
	wire _w5455_ ;
	wire _w5454_ ;
	wire _w5453_ ;
	wire _w5452_ ;
	wire _w5451_ ;
	wire _w5450_ ;
	wire _w5449_ ;
	wire _w5448_ ;
	wire _w5447_ ;
	wire _w5446_ ;
	wire _w5445_ ;
	wire _w5444_ ;
	wire _w5443_ ;
	wire _w5442_ ;
	wire _w5441_ ;
	wire _w5440_ ;
	wire _w5439_ ;
	wire _w5438_ ;
	wire _w5437_ ;
	wire _w5436_ ;
	wire _w5435_ ;
	wire _w5434_ ;
	wire _w5433_ ;
	wire _w5432_ ;
	wire _w5431_ ;
	wire _w5430_ ;
	wire _w5429_ ;
	wire _w5428_ ;
	wire _w5427_ ;
	wire _w5426_ ;
	wire _w5425_ ;
	wire _w5424_ ;
	wire _w5423_ ;
	wire _w5422_ ;
	wire _w5421_ ;
	wire _w5420_ ;
	wire _w5419_ ;
	wire _w5418_ ;
	wire _w5417_ ;
	wire _w5416_ ;
	wire _w5415_ ;
	wire _w5414_ ;
	wire _w5413_ ;
	wire _w5412_ ;
	wire _w5411_ ;
	wire _w5410_ ;
	wire _w5409_ ;
	wire _w5408_ ;
	wire _w5407_ ;
	wire _w5406_ ;
	wire _w5405_ ;
	wire _w5404_ ;
	wire _w5403_ ;
	wire _w5402_ ;
	wire _w5401_ ;
	wire _w5400_ ;
	wire _w5399_ ;
	wire _w5398_ ;
	wire _w5397_ ;
	wire _w5396_ ;
	wire _w5395_ ;
	wire _w5394_ ;
	wire _w5393_ ;
	wire _w5392_ ;
	wire _w5391_ ;
	wire _w5390_ ;
	wire _w5389_ ;
	wire _w5388_ ;
	wire _w5387_ ;
	wire _w5386_ ;
	wire _w5385_ ;
	wire _w5384_ ;
	wire _w5383_ ;
	wire _w5382_ ;
	wire _w5381_ ;
	wire _w5380_ ;
	wire _w5379_ ;
	wire _w5378_ ;
	wire _w5377_ ;
	wire _w5376_ ;
	wire _w5375_ ;
	wire _w5374_ ;
	wire _w5373_ ;
	wire _w5372_ ;
	wire _w5371_ ;
	wire _w5370_ ;
	wire _w5369_ ;
	wire _w5368_ ;
	wire _w5367_ ;
	wire _w5366_ ;
	wire _w5365_ ;
	wire _w5364_ ;
	wire _w5363_ ;
	wire _w5362_ ;
	wire _w5361_ ;
	wire _w5360_ ;
	wire _w5359_ ;
	wire _w5358_ ;
	wire _w5357_ ;
	wire _w5356_ ;
	wire _w5355_ ;
	wire _w5354_ ;
	wire _w5353_ ;
	wire _w5352_ ;
	wire _w5351_ ;
	wire _w5350_ ;
	wire _w5349_ ;
	wire _w5348_ ;
	wire _w5347_ ;
	wire _w5346_ ;
	wire _w5345_ ;
	wire _w5344_ ;
	wire _w5343_ ;
	wire _w5342_ ;
	wire _w5341_ ;
	wire _w5340_ ;
	wire _w5339_ ;
	wire _w5338_ ;
	wire _w5337_ ;
	wire _w5336_ ;
	wire _w5335_ ;
	wire _w5334_ ;
	wire _w5333_ ;
	wire _w5332_ ;
	wire _w5331_ ;
	wire _w5330_ ;
	wire _w5329_ ;
	wire _w5328_ ;
	wire _w5327_ ;
	wire _w5326_ ;
	wire _w5325_ ;
	wire _w5324_ ;
	wire _w5323_ ;
	wire _w5322_ ;
	wire _w5321_ ;
	wire _w5320_ ;
	wire _w5319_ ;
	wire _w5318_ ;
	wire _w5317_ ;
	wire _w5316_ ;
	wire _w5315_ ;
	wire _w5314_ ;
	wire _w5313_ ;
	wire _w5312_ ;
	wire _w5311_ ;
	wire _w5310_ ;
	wire _w5309_ ;
	wire _w5308_ ;
	wire _w5307_ ;
	wire _w5306_ ;
	wire _w5305_ ;
	wire _w5304_ ;
	wire _w5303_ ;
	wire _w5302_ ;
	wire _w5301_ ;
	wire _w5300_ ;
	wire _w5299_ ;
	wire _w5298_ ;
	wire _w5297_ ;
	wire _w5296_ ;
	wire _w5295_ ;
	wire _w5294_ ;
	wire _w5293_ ;
	wire _w5292_ ;
	wire _w5291_ ;
	wire _w5290_ ;
	wire _w5289_ ;
	wire _w5288_ ;
	wire _w5287_ ;
	wire _w5286_ ;
	wire _w5285_ ;
	wire _w5284_ ;
	wire _w5283_ ;
	wire _w5282_ ;
	wire _w5281_ ;
	wire _w5280_ ;
	wire _w5279_ ;
	wire _w5278_ ;
	wire _w5277_ ;
	wire _w5276_ ;
	wire _w5275_ ;
	wire _w5274_ ;
	wire _w5273_ ;
	wire _w5272_ ;
	wire _w5271_ ;
	wire _w5270_ ;
	wire _w5269_ ;
	wire _w5268_ ;
	wire _w5267_ ;
	wire _w5266_ ;
	wire _w5265_ ;
	wire _w5264_ ;
	wire _w5263_ ;
	wire _w5262_ ;
	wire _w5261_ ;
	wire _w5260_ ;
	wire _w5259_ ;
	wire _w5258_ ;
	wire _w5257_ ;
	wire _w5256_ ;
	wire _w5255_ ;
	wire _w5254_ ;
	wire _w5253_ ;
	wire _w5252_ ;
	wire _w5251_ ;
	wire _w5250_ ;
	wire _w5249_ ;
	wire _w5248_ ;
	wire _w5247_ ;
	wire _w5246_ ;
	wire _w5245_ ;
	wire _w5244_ ;
	wire _w5243_ ;
	wire _w5242_ ;
	wire _w5241_ ;
	wire _w5240_ ;
	wire _w5239_ ;
	wire _w5238_ ;
	wire _w5237_ ;
	wire _w5236_ ;
	wire _w5235_ ;
	wire _w5234_ ;
	wire _w5233_ ;
	wire _w5232_ ;
	wire _w5231_ ;
	wire _w5230_ ;
	wire _w5229_ ;
	wire _w5228_ ;
	wire _w5227_ ;
	wire _w5226_ ;
	wire _w5225_ ;
	wire _w5224_ ;
	wire _w5223_ ;
	wire _w5222_ ;
	wire _w5221_ ;
	wire _w5220_ ;
	wire _w5219_ ;
	wire _w5218_ ;
	wire _w5217_ ;
	wire _w5216_ ;
	wire _w5215_ ;
	wire _w5214_ ;
	wire _w5213_ ;
	wire _w5212_ ;
	wire _w5211_ ;
	wire _w5210_ ;
	wire _w5209_ ;
	wire _w5208_ ;
	wire _w5207_ ;
	wire _w5206_ ;
	wire _w5205_ ;
	wire _w5204_ ;
	wire _w5203_ ;
	wire _w5202_ ;
	wire _w5201_ ;
	wire _w5200_ ;
	wire _w5199_ ;
	wire _w5198_ ;
	wire _w5197_ ;
	wire _w5196_ ;
	wire _w5195_ ;
	wire _w5194_ ;
	wire _w5193_ ;
	wire _w5192_ ;
	wire _w5191_ ;
	wire _w5190_ ;
	wire _w5189_ ;
	wire _w5188_ ;
	wire _w5187_ ;
	wire _w5186_ ;
	wire _w5185_ ;
	wire _w5184_ ;
	wire _w5183_ ;
	wire _w5182_ ;
	wire _w5181_ ;
	wire _w5180_ ;
	wire _w5179_ ;
	wire _w5178_ ;
	wire _w5177_ ;
	wire _w5176_ ;
	wire _w5175_ ;
	wire _w5174_ ;
	wire _w5173_ ;
	wire _w5172_ ;
	wire _w5171_ ;
	wire _w5170_ ;
	wire _w5169_ ;
	wire _w5168_ ;
	wire _w5167_ ;
	wire _w5166_ ;
	wire _w5165_ ;
	wire _w5164_ ;
	wire _w5163_ ;
	wire _w5162_ ;
	wire _w5161_ ;
	wire _w5160_ ;
	wire _w5159_ ;
	wire _w5158_ ;
	wire _w5157_ ;
	wire _w5156_ ;
	wire _w5155_ ;
	wire _w5154_ ;
	wire _w5153_ ;
	wire _w5152_ ;
	wire _w5151_ ;
	wire _w5150_ ;
	wire _w5149_ ;
	wire _w5148_ ;
	wire _w5147_ ;
	wire _w5146_ ;
	wire _w5145_ ;
	wire _w5144_ ;
	wire _w5143_ ;
	wire _w5142_ ;
	wire _w5141_ ;
	wire _w5140_ ;
	wire _w5139_ ;
	wire _w5138_ ;
	wire _w5137_ ;
	wire _w5136_ ;
	wire _w5135_ ;
	wire _w5134_ ;
	wire _w5133_ ;
	wire _w5132_ ;
	wire _w5131_ ;
	wire _w5130_ ;
	wire _w5129_ ;
	wire _w5128_ ;
	wire _w5127_ ;
	wire _w5126_ ;
	wire _w5125_ ;
	wire _w5124_ ;
	wire _w5123_ ;
	wire _w5122_ ;
	wire _w5121_ ;
	wire _w5120_ ;
	wire _w5119_ ;
	wire _w5118_ ;
	wire _w5117_ ;
	wire _w5116_ ;
	wire _w5115_ ;
	wire _w5114_ ;
	wire _w5113_ ;
	wire _w5112_ ;
	wire _w5111_ ;
	wire _w5110_ ;
	wire _w5109_ ;
	wire _w5108_ ;
	wire _w5107_ ;
	wire _w5106_ ;
	wire _w5105_ ;
	wire _w5104_ ;
	wire _w5103_ ;
	wire _w5102_ ;
	wire _w5101_ ;
	wire _w5100_ ;
	wire _w5099_ ;
	wire _w5098_ ;
	wire _w5097_ ;
	wire _w5096_ ;
	wire _w5095_ ;
	wire _w5094_ ;
	wire _w5093_ ;
	wire _w5092_ ;
	wire _w5091_ ;
	wire _w5090_ ;
	wire _w5089_ ;
	wire _w5088_ ;
	wire _w5087_ ;
	wire _w5086_ ;
	wire _w5085_ ;
	wire _w5084_ ;
	wire _w5083_ ;
	wire _w5082_ ;
	wire _w5081_ ;
	wire _w5080_ ;
	wire _w5079_ ;
	wire _w5078_ ;
	wire _w5077_ ;
	wire _w5076_ ;
	wire _w5075_ ;
	wire _w5074_ ;
	wire _w5073_ ;
	wire _w5072_ ;
	wire _w5071_ ;
	wire _w5070_ ;
	wire _w5069_ ;
	wire _w5068_ ;
	wire _w5067_ ;
	wire _w5066_ ;
	wire _w5065_ ;
	wire _w5064_ ;
	wire _w5063_ ;
	wire _w5062_ ;
	wire _w5061_ ;
	wire _w5060_ ;
	wire _w5059_ ;
	wire _w5058_ ;
	wire _w5057_ ;
	wire _w5056_ ;
	wire _w5055_ ;
	wire _w5054_ ;
	wire _w5053_ ;
	wire _w5052_ ;
	wire _w5051_ ;
	wire _w5050_ ;
	wire _w5049_ ;
	wire _w5048_ ;
	wire _w5047_ ;
	wire _w5046_ ;
	wire _w5045_ ;
	wire _w5044_ ;
	wire _w5043_ ;
	wire _w5042_ ;
	wire _w5041_ ;
	wire _w5040_ ;
	wire _w5039_ ;
	wire _w5038_ ;
	wire _w5037_ ;
	wire _w5036_ ;
	wire _w5035_ ;
	wire _w5034_ ;
	wire _w5033_ ;
	wire _w5032_ ;
	wire _w5031_ ;
	wire _w5030_ ;
	wire _w5029_ ;
	wire _w5028_ ;
	wire _w5027_ ;
	wire _w5026_ ;
	wire _w5025_ ;
	wire _w5024_ ;
	wire _w5023_ ;
	wire _w5022_ ;
	wire _w5021_ ;
	wire _w5020_ ;
	wire _w5019_ ;
	wire _w5018_ ;
	wire _w5017_ ;
	wire _w5016_ ;
	wire _w5015_ ;
	wire _w5014_ ;
	wire _w5013_ ;
	wire _w5012_ ;
	wire _w5011_ ;
	wire _w5010_ ;
	wire _w5009_ ;
	wire _w5008_ ;
	wire _w5007_ ;
	wire _w5006_ ;
	wire _w5005_ ;
	wire _w5004_ ;
	wire _w5003_ ;
	wire _w5002_ ;
	wire _w5001_ ;
	wire _w5000_ ;
	wire _w4999_ ;
	wire _w4998_ ;
	wire _w4997_ ;
	wire _w4996_ ;
	wire _w4995_ ;
	wire _w4994_ ;
	wire _w4993_ ;
	wire _w4992_ ;
	wire _w4991_ ;
	wire _w4990_ ;
	wire _w4989_ ;
	wire _w4988_ ;
	wire _w4987_ ;
	wire _w4986_ ;
	wire _w4985_ ;
	wire _w4984_ ;
	wire _w4983_ ;
	wire _w4982_ ;
	wire _w4981_ ;
	wire _w4980_ ;
	wire _w4979_ ;
	wire _w4978_ ;
	wire _w4977_ ;
	wire _w4976_ ;
	wire _w4975_ ;
	wire _w4974_ ;
	wire _w4973_ ;
	wire _w4972_ ;
	wire _w4971_ ;
	wire _w4970_ ;
	wire _w4969_ ;
	wire _w4968_ ;
	wire _w4967_ ;
	wire _w4966_ ;
	wire _w4965_ ;
	wire _w4964_ ;
	wire _w4963_ ;
	wire _w4962_ ;
	wire _w4961_ ;
	wire _w4960_ ;
	wire _w4959_ ;
	wire _w4958_ ;
	wire _w4957_ ;
	wire _w4956_ ;
	wire _w4955_ ;
	wire _w4954_ ;
	wire _w4953_ ;
	wire _w4952_ ;
	wire _w4951_ ;
	wire _w4950_ ;
	wire _w4949_ ;
	wire _w4948_ ;
	wire _w4947_ ;
	wire _w4946_ ;
	wire _w4945_ ;
	wire _w4944_ ;
	wire _w4943_ ;
	wire _w4942_ ;
	wire _w4941_ ;
	wire _w4940_ ;
	wire _w4939_ ;
	wire _w4938_ ;
	wire _w4937_ ;
	wire _w4936_ ;
	wire _w4935_ ;
	wire _w4934_ ;
	wire _w4933_ ;
	wire _w4932_ ;
	wire _w4931_ ;
	wire _w4930_ ;
	wire _w4929_ ;
	wire _w4928_ ;
	wire _w4927_ ;
	wire _w4926_ ;
	wire _w4925_ ;
	wire _w4924_ ;
	wire _w4923_ ;
	wire _w4922_ ;
	wire _w4921_ ;
	wire _w4920_ ;
	wire _w4919_ ;
	wire _w4918_ ;
	wire _w4917_ ;
	wire _w4916_ ;
	wire _w4915_ ;
	wire _w4914_ ;
	wire _w4913_ ;
	wire _w4912_ ;
	wire _w4911_ ;
	wire _w4910_ ;
	wire _w4909_ ;
	wire _w4908_ ;
	wire _w4907_ ;
	wire _w4906_ ;
	wire _w4905_ ;
	wire _w4904_ ;
	wire _w4903_ ;
	wire _w4902_ ;
	wire _w4901_ ;
	wire _w4900_ ;
	wire _w4899_ ;
	wire _w4898_ ;
	wire _w4897_ ;
	wire _w4896_ ;
	wire _w4895_ ;
	wire _w4894_ ;
	wire _w4893_ ;
	wire _w4892_ ;
	wire _w4891_ ;
	wire _w4890_ ;
	wire _w4889_ ;
	wire _w4888_ ;
	wire _w4887_ ;
	wire _w4886_ ;
	wire _w4885_ ;
	wire _w4884_ ;
	wire _w4883_ ;
	wire _w4882_ ;
	wire _w4881_ ;
	wire _w4880_ ;
	wire _w4879_ ;
	wire _w4878_ ;
	wire _w4877_ ;
	wire _w4876_ ;
	wire _w4875_ ;
	wire _w4874_ ;
	wire _w4873_ ;
	wire _w4872_ ;
	wire _w4871_ ;
	wire _w4870_ ;
	wire _w4869_ ;
	wire _w4868_ ;
	wire _w4867_ ;
	wire _w4866_ ;
	wire _w4865_ ;
	wire _w4864_ ;
	wire _w4863_ ;
	wire _w4862_ ;
	wire _w4861_ ;
	wire _w4860_ ;
	wire _w4859_ ;
	wire _w4858_ ;
	wire _w4857_ ;
	wire _w4856_ ;
	wire _w4855_ ;
	wire _w4854_ ;
	wire _w4853_ ;
	wire _w4852_ ;
	wire _w4851_ ;
	wire _w4850_ ;
	wire _w4849_ ;
	wire _w4848_ ;
	wire _w4847_ ;
	wire _w4846_ ;
	wire _w4845_ ;
	wire _w4844_ ;
	wire _w4843_ ;
	wire _w4842_ ;
	wire _w4841_ ;
	wire _w4840_ ;
	wire _w4839_ ;
	wire _w4838_ ;
	wire _w4837_ ;
	wire _w4836_ ;
	wire _w4835_ ;
	wire _w4834_ ;
	wire _w4833_ ;
	wire _w4832_ ;
	wire _w4831_ ;
	wire _w4830_ ;
	wire _w4829_ ;
	wire _w4828_ ;
	wire _w4827_ ;
	wire _w4826_ ;
	wire _w4825_ ;
	wire _w4824_ ;
	wire _w4823_ ;
	wire _w4822_ ;
	wire _w4821_ ;
	wire _w4820_ ;
	wire _w4819_ ;
	wire _w4818_ ;
	wire _w4817_ ;
	wire _w4816_ ;
	wire _w4815_ ;
	wire _w4814_ ;
	wire _w4813_ ;
	wire _w4812_ ;
	wire _w4811_ ;
	wire _w4810_ ;
	wire _w4809_ ;
	wire _w4808_ ;
	wire _w4807_ ;
	wire _w4806_ ;
	wire _w4805_ ;
	wire _w4804_ ;
	wire _w4803_ ;
	wire _w4802_ ;
	wire _w4801_ ;
	wire _w4800_ ;
	wire _w4799_ ;
	wire _w4798_ ;
	wire _w4797_ ;
	wire _w4796_ ;
	wire _w4795_ ;
	wire _w4794_ ;
	wire _w4793_ ;
	wire _w4792_ ;
	wire _w4791_ ;
	wire _w4790_ ;
	wire _w4789_ ;
	wire _w4788_ ;
	wire _w4787_ ;
	wire _w4786_ ;
	wire _w4785_ ;
	wire _w4784_ ;
	wire _w4783_ ;
	wire _w4782_ ;
	wire _w4781_ ;
	wire _w4780_ ;
	wire _w4779_ ;
	wire _w4778_ ;
	wire _w4777_ ;
	wire _w4776_ ;
	wire _w4775_ ;
	wire _w4774_ ;
	wire _w4773_ ;
	wire _w4772_ ;
	wire _w4771_ ;
	wire _w4770_ ;
	wire _w4769_ ;
	wire _w4768_ ;
	wire _w4767_ ;
	wire _w4766_ ;
	wire _w4765_ ;
	wire _w4764_ ;
	wire _w4763_ ;
	wire _w4762_ ;
	wire _w4761_ ;
	wire _w4760_ ;
	wire _w4759_ ;
	wire _w4758_ ;
	wire _w4757_ ;
	wire _w4756_ ;
	wire _w4755_ ;
	wire _w4754_ ;
	wire _w4753_ ;
	wire _w4752_ ;
	wire _w4751_ ;
	wire _w4750_ ;
	wire _w4749_ ;
	wire _w4748_ ;
	wire _w4747_ ;
	wire _w4746_ ;
	wire _w4745_ ;
	wire _w4744_ ;
	wire _w4743_ ;
	wire _w4742_ ;
	wire _w4741_ ;
	wire _w4740_ ;
	wire _w4739_ ;
	wire _w4738_ ;
	wire _w4737_ ;
	wire _w4736_ ;
	wire _w4735_ ;
	wire _w4734_ ;
	wire _w4733_ ;
	wire _w4732_ ;
	wire _w4731_ ;
	wire _w4730_ ;
	wire _w4729_ ;
	wire _w4728_ ;
	wire _w4727_ ;
	wire _w4726_ ;
	wire _w4725_ ;
	wire _w4724_ ;
	wire _w4723_ ;
	wire _w4722_ ;
	wire _w4721_ ;
	wire _w4720_ ;
	wire _w4719_ ;
	wire _w4718_ ;
	wire _w4717_ ;
	wire _w4716_ ;
	wire _w4715_ ;
	wire _w4714_ ;
	wire _w4713_ ;
	wire _w4712_ ;
	wire _w4711_ ;
	wire _w4710_ ;
	wire _w4709_ ;
	wire _w4708_ ;
	wire _w4707_ ;
	wire _w4706_ ;
	wire _w4705_ ;
	wire _w4704_ ;
	wire _w4703_ ;
	wire _w4702_ ;
	wire _w4701_ ;
	wire _w4700_ ;
	wire _w4699_ ;
	wire _w4698_ ;
	wire _w4697_ ;
	wire _w4696_ ;
	wire _w4695_ ;
	wire _w4694_ ;
	wire _w4693_ ;
	wire _w4692_ ;
	wire _w4691_ ;
	wire _w4690_ ;
	wire _w4689_ ;
	wire _w4688_ ;
	wire _w4687_ ;
	wire _w4686_ ;
	wire _w4685_ ;
	wire _w4684_ ;
	wire _w4683_ ;
	wire _w4682_ ;
	wire _w4681_ ;
	wire _w4680_ ;
	wire _w4679_ ;
	wire _w4678_ ;
	wire _w4677_ ;
	wire _w4676_ ;
	wire _w4675_ ;
	wire _w4674_ ;
	wire _w4673_ ;
	wire _w4672_ ;
	wire _w4671_ ;
	wire _w4670_ ;
	wire _w4669_ ;
	wire _w4668_ ;
	wire _w4667_ ;
	wire _w4666_ ;
	wire _w4665_ ;
	wire _w4664_ ;
	wire _w4663_ ;
	wire _w4662_ ;
	wire _w4661_ ;
	wire _w4660_ ;
	wire _w4659_ ;
	wire _w4658_ ;
	wire _w4657_ ;
	wire _w4656_ ;
	wire _w4655_ ;
	wire _w4654_ ;
	wire _w4653_ ;
	wire _w4652_ ;
	wire _w4651_ ;
	wire _w4650_ ;
	wire _w4649_ ;
	wire _w4648_ ;
	wire _w4647_ ;
	wire _w4646_ ;
	wire _w4645_ ;
	wire _w4644_ ;
	wire _w4643_ ;
	wire _w4642_ ;
	wire _w4641_ ;
	wire _w4640_ ;
	wire _w4639_ ;
	wire _w4638_ ;
	wire _w4637_ ;
	wire _w4636_ ;
	wire _w4635_ ;
	wire _w4634_ ;
	wire _w4633_ ;
	wire _w4632_ ;
	wire _w4631_ ;
	wire _w4630_ ;
	wire _w4629_ ;
	wire _w4628_ ;
	wire _w4627_ ;
	wire _w4626_ ;
	wire _w4625_ ;
	wire _w4624_ ;
	wire _w4623_ ;
	wire _w4622_ ;
	wire _w4621_ ;
	wire _w4620_ ;
	wire _w4619_ ;
	wire _w4618_ ;
	wire _w4617_ ;
	wire _w4616_ ;
	wire _w4615_ ;
	wire _w4614_ ;
	wire _w4613_ ;
	wire _w4612_ ;
	wire _w4611_ ;
	wire _w4610_ ;
	wire _w4609_ ;
	wire _w4608_ ;
	wire _w4607_ ;
	wire _w4606_ ;
	wire _w4605_ ;
	wire _w4604_ ;
	wire _w4603_ ;
	wire _w4602_ ;
	wire _w4601_ ;
	wire _w4600_ ;
	wire _w4599_ ;
	wire _w4598_ ;
	wire _w4597_ ;
	wire _w4596_ ;
	wire _w4595_ ;
	wire _w4594_ ;
	wire _w4593_ ;
	wire _w4592_ ;
	wire _w4591_ ;
	wire _w4590_ ;
	wire _w4589_ ;
	wire _w4588_ ;
	wire _w4587_ ;
	wire _w4586_ ;
	wire _w4585_ ;
	wire _w4584_ ;
	wire _w4583_ ;
	wire _w4582_ ;
	wire _w4581_ ;
	wire _w4580_ ;
	wire _w4579_ ;
	wire _w4578_ ;
	wire _w4577_ ;
	wire _w4576_ ;
	wire _w4575_ ;
	wire _w4574_ ;
	wire _w4573_ ;
	wire _w4572_ ;
	wire _w4571_ ;
	wire _w4570_ ;
	wire _w4569_ ;
	wire _w4568_ ;
	wire _w4567_ ;
	wire _w4566_ ;
	wire _w4565_ ;
	wire _w4564_ ;
	wire _w4563_ ;
	wire _w4562_ ;
	wire _w4561_ ;
	wire _w4560_ ;
	wire _w4559_ ;
	wire _w4558_ ;
	wire _w4557_ ;
	wire _w4556_ ;
	wire _w4555_ ;
	wire _w4554_ ;
	wire _w4553_ ;
	wire _w4552_ ;
	wire _w4551_ ;
	wire _w4550_ ;
	wire _w4549_ ;
	wire _w4548_ ;
	wire _w4547_ ;
	wire _w4546_ ;
	wire _w4545_ ;
	wire _w4544_ ;
	wire _w4543_ ;
	wire _w4542_ ;
	wire _w4541_ ;
	wire _w4540_ ;
	wire _w4539_ ;
	wire _w4538_ ;
	wire _w4537_ ;
	wire _w4536_ ;
	wire _w4535_ ;
	wire _w4534_ ;
	wire _w4533_ ;
	wire _w4532_ ;
	wire _w4531_ ;
	wire _w4530_ ;
	wire _w4529_ ;
	wire _w4528_ ;
	wire _w4527_ ;
	wire _w4526_ ;
	wire _w4525_ ;
	wire _w4524_ ;
	wire _w4523_ ;
	wire _w4522_ ;
	wire _w4521_ ;
	wire _w4520_ ;
	wire _w4519_ ;
	wire _w4518_ ;
	wire _w4517_ ;
	wire _w4516_ ;
	wire _w4515_ ;
	wire _w4514_ ;
	wire _w4513_ ;
	wire _w4512_ ;
	wire _w4511_ ;
	wire _w4510_ ;
	wire _w4509_ ;
	wire _w4508_ ;
	wire _w4507_ ;
	wire _w4506_ ;
	wire _w4505_ ;
	wire _w4504_ ;
	wire _w3255_ ;
	wire _w3254_ ;
	wire _w3253_ ;
	wire _w3252_ ;
	wire _w3251_ ;
	wire _w3250_ ;
	wire _w3249_ ;
	wire _w3248_ ;
	wire _w3247_ ;
	wire _w3246_ ;
	wire _w3245_ ;
	wire _w3244_ ;
	wire _w3243_ ;
	wire _w3242_ ;
	wire _w3241_ ;
	wire _w3240_ ;
	wire _w3239_ ;
	wire _w3238_ ;
	wire _w3237_ ;
	wire _w3236_ ;
	wire _w3235_ ;
	wire _w3234_ ;
	wire _w3233_ ;
	wire _w3232_ ;
	wire _w3231_ ;
	wire _w3230_ ;
	wire _w3229_ ;
	wire _w3228_ ;
	wire _w3227_ ;
	wire _w3226_ ;
	wire _w3225_ ;
	wire _w3224_ ;
	wire _w3223_ ;
	wire _w3222_ ;
	wire _w3221_ ;
	wire _w3220_ ;
	wire _w3219_ ;
	wire _w3218_ ;
	wire _w3217_ ;
	wire _w3216_ ;
	wire _w3215_ ;
	wire _w3214_ ;
	wire _w3213_ ;
	wire _w3212_ ;
	wire _w3211_ ;
	wire _w3210_ ;
	wire _w3209_ ;
	wire _w3208_ ;
	wire _w3207_ ;
	wire _w3206_ ;
	wire _w3205_ ;
	wire _w3204_ ;
	wire _w3203_ ;
	wire _w3202_ ;
	wire _w3201_ ;
	wire _w3200_ ;
	wire _w3199_ ;
	wire _w3198_ ;
	wire _w3197_ ;
	wire _w3196_ ;
	wire _w3195_ ;
	wire _w3194_ ;
	wire _w3193_ ;
	wire _w3192_ ;
	wire _w3191_ ;
	wire _w3190_ ;
	wire _w3189_ ;
	wire _w3188_ ;
	wire _w3187_ ;
	wire _w3186_ ;
	wire _w3185_ ;
	wire _w3184_ ;
	wire _w3183_ ;
	wire _w3182_ ;
	wire _w3181_ ;
	wire _w3180_ ;
	wire _w3179_ ;
	wire _w3178_ ;
	wire _w3177_ ;
	wire _w3176_ ;
	wire _w3175_ ;
	wire _w3174_ ;
	wire _w3173_ ;
	wire _w3172_ ;
	wire _w3171_ ;
	wire _w3170_ ;
	wire _w3169_ ;
	wire _w3168_ ;
	wire _w3167_ ;
	wire _w3166_ ;
	wire _w3165_ ;
	wire _w3164_ ;
	wire _w3163_ ;
	wire _w3162_ ;
	wire _w3161_ ;
	wire _w3160_ ;
	wire _w3159_ ;
	wire _w3158_ ;
	wire _w3157_ ;
	wire _w3156_ ;
	wire _w3155_ ;
	wire _w3154_ ;
	wire _w3153_ ;
	wire _w3152_ ;
	wire _w3151_ ;
	wire _w3150_ ;
	wire _w3149_ ;
	wire _w3148_ ;
	wire _w3147_ ;
	wire _w3146_ ;
	wire _w3145_ ;
	wire _w3144_ ;
	wire _w3143_ ;
	wire _w3142_ ;
	wire _w3141_ ;
	wire _w3140_ ;
	wire _w3139_ ;
	wire _w3138_ ;
	wire _w3137_ ;
	wire _w3136_ ;
	wire _w3135_ ;
	wire _w3134_ ;
	wire _w3133_ ;
	wire _w3132_ ;
	wire _w3131_ ;
	wire _w3130_ ;
	wire _w3129_ ;
	wire _w3128_ ;
	wire _w3127_ ;
	wire _w3126_ ;
	wire _w3125_ ;
	wire _w3124_ ;
	wire _w3123_ ;
	wire _w3122_ ;
	wire _w3121_ ;
	wire _w3120_ ;
	wire _w3119_ ;
	wire _w3118_ ;
	wire _w3117_ ;
	wire _w3116_ ;
	wire _w3115_ ;
	wire _w3114_ ;
	wire _w3113_ ;
	wire _w3112_ ;
	wire _w3111_ ;
	wire _w3110_ ;
	wire _w3109_ ;
	wire _w3108_ ;
	wire _w3107_ ;
	wire _w3106_ ;
	wire _w3105_ ;
	wire _w3104_ ;
	wire _w3103_ ;
	wire _w3102_ ;
	wire _w3101_ ;
	wire _w3100_ ;
	wire _w3099_ ;
	wire _w3098_ ;
	wire _w3097_ ;
	wire _w3096_ ;
	wire _w3095_ ;
	wire _w3094_ ;
	wire _w3093_ ;
	wire _w3092_ ;
	wire _w3091_ ;
	wire _w3090_ ;
	wire _w3089_ ;
	wire _w3088_ ;
	wire _w3087_ ;
	wire _w3086_ ;
	wire _w3085_ ;
	wire _w3084_ ;
	wire _w3083_ ;
	wire _w3082_ ;
	wire _w3081_ ;
	wire _w3080_ ;
	wire _w3079_ ;
	wire _w3078_ ;
	wire _w3077_ ;
	wire _w3076_ ;
	wire _w3075_ ;
	wire _w3074_ ;
	wire _w3073_ ;
	wire _w3072_ ;
	wire _w3071_ ;
	wire _w3070_ ;
	wire _w3069_ ;
	wire _w3068_ ;
	wire _w3067_ ;
	wire _w3066_ ;
	wire _w3065_ ;
	wire _w3064_ ;
	wire _w3063_ ;
	wire _w3062_ ;
	wire _w3061_ ;
	wire _w3060_ ;
	wire _w3059_ ;
	wire _w3058_ ;
	wire _w3057_ ;
	wire _w3056_ ;
	wire _w3055_ ;
	wire _w3054_ ;
	wire _w3053_ ;
	wire _w3052_ ;
	wire _w3051_ ;
	wire _w3050_ ;
	wire _w3049_ ;
	wire _w3048_ ;
	wire _w3047_ ;
	wire _w3046_ ;
	wire _w3045_ ;
	wire _w3044_ ;
	wire _w3043_ ;
	wire _w3042_ ;
	wire _w3041_ ;
	wire _w3040_ ;
	wire _w3039_ ;
	wire _w3038_ ;
	wire _w3037_ ;
	wire _w3036_ ;
	wire _w3035_ ;
	wire _w3034_ ;
	wire _w3033_ ;
	wire _w3032_ ;
	wire _w3031_ ;
	wire _w3030_ ;
	wire _w3029_ ;
	wire _w3028_ ;
	wire _w3027_ ;
	wire _w3026_ ;
	wire _w3025_ ;
	wire _w3024_ ;
	wire _w3023_ ;
	wire _w3022_ ;
	wire _w3021_ ;
	wire _w3020_ ;
	wire _w3019_ ;
	wire _w3018_ ;
	wire _w3017_ ;
	wire _w3016_ ;
	wire _w3015_ ;
	wire _w3014_ ;
	wire _w3013_ ;
	wire _w3012_ ;
	wire _w3011_ ;
	wire _w3010_ ;
	wire _w3009_ ;
	wire _w3008_ ;
	wire _w3007_ ;
	wire _w3006_ ;
	wire _w3005_ ;
	wire _w3004_ ;
	wire _w3003_ ;
	wire _w3002_ ;
	wire _w3001_ ;
	wire _w3000_ ;
	wire _w2999_ ;
	wire _w2998_ ;
	wire _w2997_ ;
	wire _w2996_ ;
	wire _w2995_ ;
	wire _w2994_ ;
	wire _w2993_ ;
	wire _w2992_ ;
	wire _w2991_ ;
	wire _w2990_ ;
	wire _w2989_ ;
	wire _w2988_ ;
	wire _w2987_ ;
	wire _w2986_ ;
	wire _w2985_ ;
	wire _w2984_ ;
	wire _w2983_ ;
	wire _w2982_ ;
	wire _w2981_ ;
	wire _w2980_ ;
	wire _w2979_ ;
	wire _w2978_ ;
	wire _w2977_ ;
	wire _w2976_ ;
	wire _w2975_ ;
	wire _w2974_ ;
	wire _w2973_ ;
	wire _w2972_ ;
	wire _w2971_ ;
	wire _w2970_ ;
	wire _w2969_ ;
	wire _w2968_ ;
	wire _w2967_ ;
	wire _w2966_ ;
	wire _w2965_ ;
	wire _w2964_ ;
	wire _w2963_ ;
	wire _w2962_ ;
	wire _w2961_ ;
	wire _w2960_ ;
	wire _w2959_ ;
	wire _w2958_ ;
	wire _w2957_ ;
	wire _w2956_ ;
	wire _w2955_ ;
	wire _w2954_ ;
	wire _w2953_ ;
	wire _w2952_ ;
	wire _w2951_ ;
	wire _w2950_ ;
	wire _w2949_ ;
	wire _w2948_ ;
	wire _w2947_ ;
	wire _w2946_ ;
	wire _w2945_ ;
	wire _w2944_ ;
	wire _w2943_ ;
	wire _w2942_ ;
	wire _w2941_ ;
	wire _w2940_ ;
	wire _w2939_ ;
	wire _w2938_ ;
	wire _w2937_ ;
	wire _w2936_ ;
	wire _w2935_ ;
	wire _w2934_ ;
	wire _w2933_ ;
	wire _w2932_ ;
	wire _w2931_ ;
	wire _w2930_ ;
	wire _w2929_ ;
	wire _w2928_ ;
	wire _w2927_ ;
	wire _w2926_ ;
	wire _w2925_ ;
	wire _w2924_ ;
	wire _w2923_ ;
	wire _w2922_ ;
	wire _w2921_ ;
	wire _w2920_ ;
	wire _w2919_ ;
	wire _w2918_ ;
	wire _w2917_ ;
	wire _w2916_ ;
	wire _w2915_ ;
	wire _w2914_ ;
	wire _w2913_ ;
	wire _w2912_ ;
	wire _w2911_ ;
	wire _w2910_ ;
	wire _w2909_ ;
	wire _w2908_ ;
	wire _w2907_ ;
	wire _w2906_ ;
	wire _w2905_ ;
	wire _w2904_ ;
	wire _w2903_ ;
	wire _w2902_ ;
	wire _w2901_ ;
	wire _w2900_ ;
	wire _w2899_ ;
	wire _w2898_ ;
	wire _w2897_ ;
	wire _w2896_ ;
	wire _w2895_ ;
	wire _w2894_ ;
	wire _w2893_ ;
	wire _w2892_ ;
	wire _w2891_ ;
	wire _w2890_ ;
	wire _w2889_ ;
	wire _w2888_ ;
	wire _w2887_ ;
	wire _w2886_ ;
	wire _w2885_ ;
	wire _w2884_ ;
	wire _w2883_ ;
	wire _w2882_ ;
	wire _w2881_ ;
	wire _w2880_ ;
	wire _w2879_ ;
	wire _w2878_ ;
	wire _w2877_ ;
	wire _w2876_ ;
	wire _w2875_ ;
	wire _w2874_ ;
	wire _w2873_ ;
	wire _w2872_ ;
	wire _w2871_ ;
	wire _w2870_ ;
	wire _w2869_ ;
	wire _w2868_ ;
	wire _w2867_ ;
	wire _w2866_ ;
	wire _w2865_ ;
	wire _w2864_ ;
	wire _w2863_ ;
	wire _w2862_ ;
	wire _w2861_ ;
	wire _w2860_ ;
	wire _w2859_ ;
	wire _w2858_ ;
	wire _w2857_ ;
	wire _w2856_ ;
	wire _w2855_ ;
	wire _w2854_ ;
	wire _w2853_ ;
	wire _w2852_ ;
	wire _w2851_ ;
	wire _w2850_ ;
	wire _w2849_ ;
	wire _w2848_ ;
	wire _w2847_ ;
	wire _w2846_ ;
	wire _w2845_ ;
	wire _w2844_ ;
	wire _w2843_ ;
	wire _w2842_ ;
	wire _w2841_ ;
	wire _w2840_ ;
	wire _w2839_ ;
	wire _w2838_ ;
	wire _w2837_ ;
	wire _w2836_ ;
	wire _w2835_ ;
	wire _w2834_ ;
	wire _w2833_ ;
	wire _w2832_ ;
	wire _w2831_ ;
	wire _w2830_ ;
	wire _w2829_ ;
	wire _w2828_ ;
	wire _w2827_ ;
	wire _w2826_ ;
	wire _w2825_ ;
	wire _w2824_ ;
	wire _w2823_ ;
	wire _w2822_ ;
	wire _w2821_ ;
	wire _w2820_ ;
	wire _w2819_ ;
	wire _w2818_ ;
	wire _w2817_ ;
	wire _w2816_ ;
	wire _w2815_ ;
	wire _w2814_ ;
	wire _w2813_ ;
	wire _w2812_ ;
	wire _w2811_ ;
	wire _w2810_ ;
	wire _w2809_ ;
	wire _w2808_ ;
	wire _w2807_ ;
	wire _w2806_ ;
	wire _w2805_ ;
	wire _w2804_ ;
	wire _w2803_ ;
	wire _w2802_ ;
	wire _w2801_ ;
	wire _w2800_ ;
	wire _w2799_ ;
	wire _w2798_ ;
	wire _w2797_ ;
	wire _w2796_ ;
	wire _w2795_ ;
	wire _w2794_ ;
	wire _w2793_ ;
	wire _w2792_ ;
	wire _w2791_ ;
	wire _w2790_ ;
	wire _w2789_ ;
	wire _w2788_ ;
	wire _w2787_ ;
	wire _w2786_ ;
	wire _w2785_ ;
	wire _w2784_ ;
	wire _w2783_ ;
	wire _w2782_ ;
	wire _w2781_ ;
	wire _w2780_ ;
	wire _w2779_ ;
	wire _w2778_ ;
	wire _w2777_ ;
	wire _w2776_ ;
	wire _w2775_ ;
	wire _w2774_ ;
	wire _w2773_ ;
	wire _w2772_ ;
	wire _w2771_ ;
	wire _w2770_ ;
	wire _w2769_ ;
	wire _w2768_ ;
	wire _w2767_ ;
	wire _w2766_ ;
	wire _w2765_ ;
	wire _w2764_ ;
	wire _w2763_ ;
	wire _w2762_ ;
	wire _w2761_ ;
	wire _w2760_ ;
	wire _w2759_ ;
	wire _w2758_ ;
	wire _w2757_ ;
	wire _w2756_ ;
	wire _w2755_ ;
	wire _w2754_ ;
	wire _w2753_ ;
	wire _w2752_ ;
	wire _w2751_ ;
	wire _w2750_ ;
	wire _w2749_ ;
	wire _w2748_ ;
	wire _w2747_ ;
	wire _w2746_ ;
	wire _w2745_ ;
	wire _w2744_ ;
	wire _w2743_ ;
	wire _w2742_ ;
	wire _w2741_ ;
	wire _w2740_ ;
	wire _w2739_ ;
	wire _w2738_ ;
	wire _w2737_ ;
	wire _w2736_ ;
	wire _w2735_ ;
	wire _w2734_ ;
	wire _w2733_ ;
	wire _w2732_ ;
	wire _w2731_ ;
	wire _w2730_ ;
	wire _w2729_ ;
	wire _w2728_ ;
	wire _w2727_ ;
	wire _w2726_ ;
	wire _w2725_ ;
	wire _w2724_ ;
	wire _w2723_ ;
	wire _w2722_ ;
	wire _w2721_ ;
	wire _w2720_ ;
	wire _w2719_ ;
	wire _w2718_ ;
	wire _w2717_ ;
	wire _w2716_ ;
	wire _w2715_ ;
	wire _w2714_ ;
	wire _w2713_ ;
	wire _w2712_ ;
	wire _w2711_ ;
	wire _w2710_ ;
	wire _w2709_ ;
	wire _w2708_ ;
	wire _w2707_ ;
	wire _w2706_ ;
	wire _w2705_ ;
	wire _w2704_ ;
	wire _w2703_ ;
	wire _w2702_ ;
	wire _w2701_ ;
	wire _w2700_ ;
	wire _w2699_ ;
	wire _w2698_ ;
	wire _w2697_ ;
	wire _w2696_ ;
	wire _w2695_ ;
	wire _w2694_ ;
	wire _w2693_ ;
	wire _w2692_ ;
	wire _w2691_ ;
	wire _w2690_ ;
	wire _w2689_ ;
	wire _w2688_ ;
	wire _w2403_ ;
	wire _w2402_ ;
	wire _w2401_ ;
	wire _w2400_ ;
	wire _w2399_ ;
	wire _w2398_ ;
	wire _w2397_ ;
	wire _w2396_ ;
	wire _w2395_ ;
	wire _w2394_ ;
	wire _w2393_ ;
	wire _w2392_ ;
	wire _w2391_ ;
	wire _w2390_ ;
	wire _w2389_ ;
	wire _w2388_ ;
	wire _w2387_ ;
	wire _w2386_ ;
	wire _w2385_ ;
	wire _w2384_ ;
	wire _w2383_ ;
	wire _w2382_ ;
	wire _w2381_ ;
	wire _w2380_ ;
	wire _w2379_ ;
	wire _w2378_ ;
	wire _w2377_ ;
	wire _w2376_ ;
	wire _w2375_ ;
	wire _w2374_ ;
	wire _w2373_ ;
	wire _w2372_ ;
	wire _w2371_ ;
	wire _w2370_ ;
	wire _w2369_ ;
	wire _w2368_ ;
	wire _w2367_ ;
	wire _w2366_ ;
	wire _w2365_ ;
	wire _w2364_ ;
	wire _w2363_ ;
	wire _w2362_ ;
	wire _w2361_ ;
	wire _w2360_ ;
	wire _w2359_ ;
	wire _w2358_ ;
	wire _w2357_ ;
	wire _w2356_ ;
	wire _w2355_ ;
	wire _w2354_ ;
	wire _w2353_ ;
	wire _w2352_ ;
	wire _w2351_ ;
	wire _w2350_ ;
	wire _w2349_ ;
	wire _w2348_ ;
	wire _w2347_ ;
	wire _w2346_ ;
	wire _w2345_ ;
	wire _w2344_ ;
	wire _w2343_ ;
	wire _w2342_ ;
	wire _w2341_ ;
	wire _w2340_ ;
	wire _w2339_ ;
	wire _w2338_ ;
	wire _w2337_ ;
	wire _w2336_ ;
	wire _w2335_ ;
	wire _w2334_ ;
	wire _w2333_ ;
	wire _w2332_ ;
	wire _w2331_ ;
	wire _w2330_ ;
	wire _w2329_ ;
	wire _w2328_ ;
	wire _w2327_ ;
	wire _w2326_ ;
	wire _w2325_ ;
	wire _w2324_ ;
	wire _w2323_ ;
	wire _w2322_ ;
	wire _w2321_ ;
	wire _w2320_ ;
	wire _w2319_ ;
	wire _w2318_ ;
	wire _w2317_ ;
	wire _w2316_ ;
	wire _w2315_ ;
	wire _w2314_ ;
	wire _w2313_ ;
	wire _w2312_ ;
	wire _w2311_ ;
	wire _w2310_ ;
	wire _w2309_ ;
	wire _w2308_ ;
	wire _w2307_ ;
	wire _w2306_ ;
	wire _w2305_ ;
	wire _w2304_ ;
	wire _w2303_ ;
	wire _w2302_ ;
	wire _w2301_ ;
	wire _w2300_ ;
	wire _w2299_ ;
	wire _w2298_ ;
	wire _w2297_ ;
	wire _w2296_ ;
	wire _w2295_ ;
	wire _w2294_ ;
	wire _w2293_ ;
	wire _w2292_ ;
	wire _w2291_ ;
	wire _w2290_ ;
	wire _w2289_ ;
	wire _w2288_ ;
	wire _w2287_ ;
	wire _w2286_ ;
	wire _w2285_ ;
	wire _w2284_ ;
	wire _w2283_ ;
	wire _w2282_ ;
	wire _w2281_ ;
	wire _w2280_ ;
	wire _w2279_ ;
	wire _w2278_ ;
	wire _w2277_ ;
	wire _w2276_ ;
	wire _w2275_ ;
	wire _w2274_ ;
	wire _w2205_ ;
	wire _w2204_ ;
	wire _w2203_ ;
	wire _w2202_ ;
	wire _w2201_ ;
	wire _w2200_ ;
	wire _w2199_ ;
	wire _w2198_ ;
	wire _w2197_ ;
	wire _w2196_ ;
	wire _w2195_ ;
	wire _w2194_ ;
	wire _w2193_ ;
	wire _w2192_ ;
	wire _w2191_ ;
	wire _w2190_ ;
	wire _w2189_ ;
	wire _w2188_ ;
	wire _w2187_ ;
	wire _w2186_ ;
	wire _w2185_ ;
	wire _w2184_ ;
	wire _w2183_ ;
	wire _w2182_ ;
	wire _w2181_ ;
	wire _w2180_ ;
	wire _w2179_ ;
	wire _w2178_ ;
	wire _w2177_ ;
	wire _w2176_ ;
	wire _w2159_ ;
	wire _w2158_ ;
	wire _w2157_ ;
	wire _w2156_ ;
	wire _w2155_ ;
	wire _w2154_ ;
	wire _w2153_ ;
	wire _w2152_ ;
	wire _w2151_ ;
	wire _w2150_ ;
	wire _w2149_ ;
	wire _w2148_ ;
	wire _w2147_ ;
	wire _w2160_ ;
	wire _w2161_ ;
	wire _w2162_ ;
	wire _w2163_ ;
	wire _w2164_ ;
	wire _w2165_ ;
	wire _w2166_ ;
	wire _w2167_ ;
	wire _w2168_ ;
	wire _w2169_ ;
	wire _w2170_ ;
	wire _w2171_ ;
	wire _w2172_ ;
	wire _w2173_ ;
	wire _w2174_ ;
	wire _w2175_ ;
	wire _w2206_ ;
	wire _w2207_ ;
	wire _w2208_ ;
	wire _w2209_ ;
	wire _w2210_ ;
	wire _w2211_ ;
	wire _w2212_ ;
	wire _w2213_ ;
	wire _w2214_ ;
	wire _w2215_ ;
	wire _w2216_ ;
	wire _w2217_ ;
	wire _w2218_ ;
	wire _w2219_ ;
	wire _w2220_ ;
	wire _w2221_ ;
	wire _w2222_ ;
	wire _w2223_ ;
	wire _w2224_ ;
	wire _w2225_ ;
	wire _w2226_ ;
	wire _w2227_ ;
	wire _w2228_ ;
	wire _w2229_ ;
	wire _w2230_ ;
	wire _w2231_ ;
	wire _w2232_ ;
	wire _w2233_ ;
	wire _w2234_ ;
	wire _w2235_ ;
	wire _w2236_ ;
	wire _w2237_ ;
	wire _w2238_ ;
	wire _w2239_ ;
	wire _w2240_ ;
	wire _w2241_ ;
	wire _w2242_ ;
	wire _w2243_ ;
	wire _w2244_ ;
	wire _w2245_ ;
	wire _w2246_ ;
	wire _w2247_ ;
	wire _w2248_ ;
	wire _w2249_ ;
	wire _w2250_ ;
	wire _w2251_ ;
	wire _w2252_ ;
	wire _w2253_ ;
	wire _w2254_ ;
	wire _w2255_ ;
	wire _w2256_ ;
	wire _w2257_ ;
	wire _w2258_ ;
	wire _w2259_ ;
	wire _w2260_ ;
	wire _w2261_ ;
	wire _w2262_ ;
	wire _w2263_ ;
	wire _w2264_ ;
	wire _w2265_ ;
	wire _w2266_ ;
	wire _w2267_ ;
	wire _w2268_ ;
	wire _w2269_ ;
	wire _w2270_ ;
	wire _w2271_ ;
	wire _w2272_ ;
	wire _w2273_ ;
	wire _w2404_ ;
	wire _w2405_ ;
	wire _w2406_ ;
	wire _w2407_ ;
	wire _w2408_ ;
	wire _w2409_ ;
	wire _w2410_ ;
	wire _w2411_ ;
	wire _w2412_ ;
	wire _w2413_ ;
	wire _w2414_ ;
	wire _w2415_ ;
	wire _w2416_ ;
	wire _w2417_ ;
	wire _w2418_ ;
	wire _w2419_ ;
	wire _w2420_ ;
	wire _w2421_ ;
	wire _w2422_ ;
	wire _w2423_ ;
	wire _w2424_ ;
	wire _w2425_ ;
	wire _w2426_ ;
	wire _w2427_ ;
	wire _w2428_ ;
	wire _w2429_ ;
	wire _w2430_ ;
	wire _w2431_ ;
	wire _w2432_ ;
	wire _w2433_ ;
	wire _w2434_ ;
	wire _w2435_ ;
	wire _w2436_ ;
	wire _w2437_ ;
	wire _w2438_ ;
	wire _w2439_ ;
	wire _w2440_ ;
	wire _w2441_ ;
	wire _w2442_ ;
	wire _w2443_ ;
	wire _w2444_ ;
	wire _w2445_ ;
	wire _w2446_ ;
	wire _w2447_ ;
	wire _w2448_ ;
	wire _w2449_ ;
	wire _w2450_ ;
	wire _w2451_ ;
	wire _w2452_ ;
	wire _w2453_ ;
	wire _w2454_ ;
	wire _w2455_ ;
	wire _w2456_ ;
	wire _w2457_ ;
	wire _w2458_ ;
	wire _w2459_ ;
	wire _w2460_ ;
	wire _w2461_ ;
	wire _w2462_ ;
	wire _w2463_ ;
	wire _w2464_ ;
	wire _w2465_ ;
	wire _w2466_ ;
	wire _w2467_ ;
	wire _w2468_ ;
	wire _w2469_ ;
	wire _w2470_ ;
	wire _w2471_ ;
	wire _w2472_ ;
	wire _w2473_ ;
	wire _w2474_ ;
	wire _w2475_ ;
	wire _w2476_ ;
	wire _w2477_ ;
	wire _w2478_ ;
	wire _w2479_ ;
	wire _w2480_ ;
	wire _w2481_ ;
	wire _w2482_ ;
	wire _w2483_ ;
	wire _w2484_ ;
	wire _w2485_ ;
	wire _w2486_ ;
	wire _w2487_ ;
	wire _w2488_ ;
	wire _w2489_ ;
	wire _w2490_ ;
	wire _w2491_ ;
	wire _w2492_ ;
	wire _w2493_ ;
	wire _w2494_ ;
	wire _w2495_ ;
	wire _w2496_ ;
	wire _w2497_ ;
	wire _w2498_ ;
	wire _w2499_ ;
	wire _w2500_ ;
	wire _w2501_ ;
	wire _w2502_ ;
	wire _w2503_ ;
	wire _w2504_ ;
	wire _w2505_ ;
	wire _w2506_ ;
	wire _w2507_ ;
	wire _w2508_ ;
	wire _w2509_ ;
	wire _w2510_ ;
	wire _w2511_ ;
	wire _w2512_ ;
	wire _w2513_ ;
	wire _w2514_ ;
	wire _w2515_ ;
	wire _w2516_ ;
	wire _w2517_ ;
	wire _w2518_ ;
	wire _w2519_ ;
	wire _w2520_ ;
	wire _w2521_ ;
	wire _w2522_ ;
	wire _w2523_ ;
	wire _w2524_ ;
	wire _w2525_ ;
	wire _w2526_ ;
	wire _w2527_ ;
	wire _w2528_ ;
	wire _w2529_ ;
	wire _w2530_ ;
	wire _w2531_ ;
	wire _w2532_ ;
	wire _w2533_ ;
	wire _w2534_ ;
	wire _w2535_ ;
	wire _w2536_ ;
	wire _w2537_ ;
	wire _w2538_ ;
	wire _w2539_ ;
	wire _w2540_ ;
	wire _w2541_ ;
	wire _w2542_ ;
	wire _w2543_ ;
	wire _w2544_ ;
	wire _w2545_ ;
	wire _w2546_ ;
	wire _w2547_ ;
	wire _w2548_ ;
	wire _w2549_ ;
	wire _w2550_ ;
	wire _w2551_ ;
	wire _w2552_ ;
	wire _w2553_ ;
	wire _w2554_ ;
	wire _w2555_ ;
	wire _w2556_ ;
	wire _w2557_ ;
	wire _w2558_ ;
	wire _w2559_ ;
	wire _w2560_ ;
	wire _w2561_ ;
	wire _w2562_ ;
	wire _w2563_ ;
	wire _w2564_ ;
	wire _w2565_ ;
	wire _w2566_ ;
	wire _w2567_ ;
	wire _w2568_ ;
	wire _w2569_ ;
	wire _w2570_ ;
	wire _w2571_ ;
	wire _w2572_ ;
	wire _w2573_ ;
	wire _w2574_ ;
	wire _w2575_ ;
	wire _w2576_ ;
	wire _w2577_ ;
	wire _w2578_ ;
	wire _w2579_ ;
	wire _w2580_ ;
	wire _w2581_ ;
	wire _w2582_ ;
	wire _w2583_ ;
	wire _w2584_ ;
	wire _w2585_ ;
	wire _w2586_ ;
	wire _w2587_ ;
	wire _w2588_ ;
	wire _w2589_ ;
	wire _w2590_ ;
	wire _w2591_ ;
	wire _w2592_ ;
	wire _w2593_ ;
	wire _w2594_ ;
	wire _w2595_ ;
	wire _w2596_ ;
	wire _w2597_ ;
	wire _w2598_ ;
	wire _w2599_ ;
	wire _w2600_ ;
	wire _w2601_ ;
	wire _w2602_ ;
	wire _w2603_ ;
	wire _w2604_ ;
	wire _w2605_ ;
	wire _w2606_ ;
	wire _w2607_ ;
	wire _w2608_ ;
	wire _w2609_ ;
	wire _w2610_ ;
	wire _w2611_ ;
	wire _w2612_ ;
	wire _w2613_ ;
	wire _w2614_ ;
	wire _w2615_ ;
	wire _w2616_ ;
	wire _w2617_ ;
	wire _w2618_ ;
	wire _w2619_ ;
	wire _w2620_ ;
	wire _w2621_ ;
	wire _w2622_ ;
	wire _w2623_ ;
	wire _w2624_ ;
	wire _w2625_ ;
	wire _w2626_ ;
	wire _w2627_ ;
	wire _w2628_ ;
	wire _w2629_ ;
	wire _w2630_ ;
	wire _w2631_ ;
	wire _w2632_ ;
	wire _w2633_ ;
	wire _w2634_ ;
	wire _w2635_ ;
	wire _w2636_ ;
	wire _w2637_ ;
	wire _w2638_ ;
	wire _w2639_ ;
	wire _w2640_ ;
	wire _w2641_ ;
	wire _w2642_ ;
	wire _w2643_ ;
	wire _w2644_ ;
	wire _w2645_ ;
	wire _w2646_ ;
	wire _w2647_ ;
	wire _w2648_ ;
	wire _w2649_ ;
	wire _w2650_ ;
	wire _w2651_ ;
	wire _w2652_ ;
	wire _w2653_ ;
	wire _w2654_ ;
	wire _w2655_ ;
	wire _w2656_ ;
	wire _w2657_ ;
	wire _w2658_ ;
	wire _w2659_ ;
	wire _w2660_ ;
	wire _w2661_ ;
	wire _w2662_ ;
	wire _w2663_ ;
	wire _w2664_ ;
	wire _w2665_ ;
	wire _w2666_ ;
	wire _w2667_ ;
	wire _w2668_ ;
	wire _w2669_ ;
	wire _w2670_ ;
	wire _w2671_ ;
	wire _w2672_ ;
	wire _w2673_ ;
	wire _w2674_ ;
	wire _w2675_ ;
	wire _w2676_ ;
	wire _w2677_ ;
	wire _w2678_ ;
	wire _w2679_ ;
	wire _w2680_ ;
	wire _w2681_ ;
	wire _w2682_ ;
	wire _w2683_ ;
	wire _w2684_ ;
	wire _w2685_ ;
	wire _w2686_ ;
	wire _w2687_ ;
	wire _w3256_ ;
	wire _w3257_ ;
	wire _w3258_ ;
	wire _w3259_ ;
	wire _w3260_ ;
	wire _w3261_ ;
	wire _w3262_ ;
	wire _w3263_ ;
	wire _w3264_ ;
	wire _w3265_ ;
	wire _w3266_ ;
	wire _w3267_ ;
	wire _w3268_ ;
	wire _w3269_ ;
	wire _w3270_ ;
	wire _w3271_ ;
	wire _w3272_ ;
	wire _w3273_ ;
	wire _w3274_ ;
	wire _w3275_ ;
	wire _w3276_ ;
	wire _w3277_ ;
	wire _w3278_ ;
	wire _w3279_ ;
	wire _w3280_ ;
	wire _w3281_ ;
	wire _w3282_ ;
	wire _w3283_ ;
	wire _w3284_ ;
	wire _w3285_ ;
	wire _w3286_ ;
	wire _w3287_ ;
	wire _w3288_ ;
	wire _w3289_ ;
	wire _w3290_ ;
	wire _w3291_ ;
	wire _w3292_ ;
	wire _w3293_ ;
	wire _w3294_ ;
	wire _w3295_ ;
	wire _w3296_ ;
	wire _w3297_ ;
	wire _w3298_ ;
	wire _w3299_ ;
	wire _w3300_ ;
	wire _w3301_ ;
	wire _w3302_ ;
	wire _w3303_ ;
	wire _w3304_ ;
	wire _w3305_ ;
	wire _w3306_ ;
	wire _w3307_ ;
	wire _w3308_ ;
	wire _w3309_ ;
	wire _w3310_ ;
	wire _w3311_ ;
	wire _w3312_ ;
	wire _w3313_ ;
	wire _w3314_ ;
	wire _w3315_ ;
	wire _w3316_ ;
	wire _w3317_ ;
	wire _w3318_ ;
	wire _w3319_ ;
	wire _w3320_ ;
	wire _w3321_ ;
	wire _w3322_ ;
	wire _w3323_ ;
	wire _w3324_ ;
	wire _w3325_ ;
	wire _w3326_ ;
	wire _w3327_ ;
	wire _w3328_ ;
	wire _w3329_ ;
	wire _w3330_ ;
	wire _w3331_ ;
	wire _w3332_ ;
	wire _w3333_ ;
	wire _w3334_ ;
	wire _w3335_ ;
	wire _w3336_ ;
	wire _w3337_ ;
	wire _w3338_ ;
	wire _w3339_ ;
	wire _w3340_ ;
	wire _w3341_ ;
	wire _w3342_ ;
	wire _w3343_ ;
	wire _w3344_ ;
	wire _w3345_ ;
	wire _w3346_ ;
	wire _w3347_ ;
	wire _w3348_ ;
	wire _w3349_ ;
	wire _w3350_ ;
	wire _w3351_ ;
	wire _w3352_ ;
	wire _w3353_ ;
	wire _w3354_ ;
	wire _w3355_ ;
	wire _w3356_ ;
	wire _w3357_ ;
	wire _w3358_ ;
	wire _w3359_ ;
	wire _w3360_ ;
	wire _w3361_ ;
	wire _w3362_ ;
	wire _w3363_ ;
	wire _w3364_ ;
	wire _w3365_ ;
	wire _w3366_ ;
	wire _w3367_ ;
	wire _w3368_ ;
	wire _w3369_ ;
	wire _w3370_ ;
	wire _w3371_ ;
	wire _w3372_ ;
	wire _w3373_ ;
	wire _w3374_ ;
	wire _w3375_ ;
	wire _w3376_ ;
	wire _w3377_ ;
	wire _w3378_ ;
	wire _w3379_ ;
	wire _w3380_ ;
	wire _w3381_ ;
	wire _w3382_ ;
	wire _w3383_ ;
	wire _w3384_ ;
	wire _w3385_ ;
	wire _w3386_ ;
	wire _w3387_ ;
	wire _w3388_ ;
	wire _w3389_ ;
	wire _w3390_ ;
	wire _w3391_ ;
	wire _w3392_ ;
	wire _w3393_ ;
	wire _w3394_ ;
	wire _w3395_ ;
	wire _w3396_ ;
	wire _w3397_ ;
	wire _w3398_ ;
	wire _w3399_ ;
	wire _w3400_ ;
	wire _w3401_ ;
	wire _w3402_ ;
	wire _w3403_ ;
	wire _w3404_ ;
	wire _w3405_ ;
	wire _w3406_ ;
	wire _w3407_ ;
	wire _w3408_ ;
	wire _w3409_ ;
	wire _w3410_ ;
	wire _w3411_ ;
	wire _w3412_ ;
	wire _w3413_ ;
	wire _w3414_ ;
	wire _w3415_ ;
	wire _w3416_ ;
	wire _w3417_ ;
	wire _w3418_ ;
	wire _w3419_ ;
	wire _w3420_ ;
	wire _w3421_ ;
	wire _w3422_ ;
	wire _w3423_ ;
	wire _w3424_ ;
	wire _w3425_ ;
	wire _w3426_ ;
	wire _w3427_ ;
	wire _w3428_ ;
	wire _w3429_ ;
	wire _w3430_ ;
	wire _w3431_ ;
	wire _w3432_ ;
	wire _w3433_ ;
	wire _w3434_ ;
	wire _w3435_ ;
	wire _w3436_ ;
	wire _w3437_ ;
	wire _w3438_ ;
	wire _w3439_ ;
	wire _w3440_ ;
	wire _w3441_ ;
	wire _w3442_ ;
	wire _w3443_ ;
	wire _w3444_ ;
	wire _w3445_ ;
	wire _w3446_ ;
	wire _w3447_ ;
	wire _w3448_ ;
	wire _w3449_ ;
	wire _w3450_ ;
	wire _w3451_ ;
	wire _w3452_ ;
	wire _w3453_ ;
	wire _w3454_ ;
	wire _w3455_ ;
	wire _w3456_ ;
	wire _w3457_ ;
	wire _w3458_ ;
	wire _w3459_ ;
	wire _w3460_ ;
	wire _w3461_ ;
	wire _w3462_ ;
	wire _w3463_ ;
	wire _w3464_ ;
	wire _w3465_ ;
	wire _w3466_ ;
	wire _w3467_ ;
	wire _w3468_ ;
	wire _w3469_ ;
	wire _w3470_ ;
	wire _w3471_ ;
	wire _w3472_ ;
	wire _w3473_ ;
	wire _w3474_ ;
	wire _w3475_ ;
	wire _w3476_ ;
	wire _w3477_ ;
	wire _w3478_ ;
	wire _w3479_ ;
	wire _w3480_ ;
	wire _w3481_ ;
	wire _w3482_ ;
	wire _w3483_ ;
	wire _w3484_ ;
	wire _w3485_ ;
	wire _w3486_ ;
	wire _w3487_ ;
	wire _w3488_ ;
	wire _w3489_ ;
	wire _w3490_ ;
	wire _w3491_ ;
	wire _w3492_ ;
	wire _w3493_ ;
	wire _w3494_ ;
	wire _w3495_ ;
	wire _w3496_ ;
	wire _w3497_ ;
	wire _w3498_ ;
	wire _w3499_ ;
	wire _w3500_ ;
	wire _w3501_ ;
	wire _w3502_ ;
	wire _w3503_ ;
	wire _w3504_ ;
	wire _w3505_ ;
	wire _w3506_ ;
	wire _w3507_ ;
	wire _w3508_ ;
	wire _w3509_ ;
	wire _w3510_ ;
	wire _w3511_ ;
	wire _w3512_ ;
	wire _w3513_ ;
	wire _w3514_ ;
	wire _w3515_ ;
	wire _w3516_ ;
	wire _w3517_ ;
	wire _w3518_ ;
	wire _w3519_ ;
	wire _w3520_ ;
	wire _w3521_ ;
	wire _w3522_ ;
	wire _w3523_ ;
	wire _w3524_ ;
	wire _w3525_ ;
	wire _w3526_ ;
	wire _w3527_ ;
	wire _w3528_ ;
	wire _w3529_ ;
	wire _w3530_ ;
	wire _w3531_ ;
	wire _w3532_ ;
	wire _w3533_ ;
	wire _w3534_ ;
	wire _w3535_ ;
	wire _w3536_ ;
	wire _w3537_ ;
	wire _w3538_ ;
	wire _w3539_ ;
	wire _w3540_ ;
	wire _w3541_ ;
	wire _w3542_ ;
	wire _w3543_ ;
	wire _w3544_ ;
	wire _w3545_ ;
	wire _w3546_ ;
	wire _w3547_ ;
	wire _w3548_ ;
	wire _w3549_ ;
	wire _w3550_ ;
	wire _w3551_ ;
	wire _w3552_ ;
	wire _w3553_ ;
	wire _w3554_ ;
	wire _w3555_ ;
	wire _w3556_ ;
	wire _w3557_ ;
	wire _w3558_ ;
	wire _w3559_ ;
	wire _w3560_ ;
	wire _w3561_ ;
	wire _w3562_ ;
	wire _w3563_ ;
	wire _w3564_ ;
	wire _w3565_ ;
	wire _w3566_ ;
	wire _w3567_ ;
	wire _w3568_ ;
	wire _w3569_ ;
	wire _w3570_ ;
	wire _w3571_ ;
	wire _w3572_ ;
	wire _w3573_ ;
	wire _w3574_ ;
	wire _w3575_ ;
	wire _w3576_ ;
	wire _w3577_ ;
	wire _w3578_ ;
	wire _w3579_ ;
	wire _w3580_ ;
	wire _w3581_ ;
	wire _w3582_ ;
	wire _w3583_ ;
	wire _w3584_ ;
	wire _w3585_ ;
	wire _w3586_ ;
	wire _w3587_ ;
	wire _w3588_ ;
	wire _w3589_ ;
	wire _w3590_ ;
	wire _w3591_ ;
	wire _w3592_ ;
	wire _w3593_ ;
	wire _w3594_ ;
	wire _w3595_ ;
	wire _w3596_ ;
	wire _w3597_ ;
	wire _w3598_ ;
	wire _w3599_ ;
	wire _w3600_ ;
	wire _w3601_ ;
	wire _w3602_ ;
	wire _w3603_ ;
	wire _w3604_ ;
	wire _w3605_ ;
	wire _w3606_ ;
	wire _w3607_ ;
	wire _w3608_ ;
	wire _w3609_ ;
	wire _w3610_ ;
	wire _w3611_ ;
	wire _w3612_ ;
	wire _w3613_ ;
	wire _w3614_ ;
	wire _w3615_ ;
	wire _w3616_ ;
	wire _w3617_ ;
	wire _w3618_ ;
	wire _w3619_ ;
	wire _w3620_ ;
	wire _w3621_ ;
	wire _w3622_ ;
	wire _w3623_ ;
	wire _w3624_ ;
	wire _w3625_ ;
	wire _w3626_ ;
	wire _w3627_ ;
	wire _w3628_ ;
	wire _w3629_ ;
	wire _w3630_ ;
	wire _w3631_ ;
	wire _w3632_ ;
	wire _w3633_ ;
	wire _w3634_ ;
	wire _w3635_ ;
	wire _w3636_ ;
	wire _w3637_ ;
	wire _w3638_ ;
	wire _w3639_ ;
	wire _w3640_ ;
	wire _w3641_ ;
	wire _w3642_ ;
	wire _w3643_ ;
	wire _w3644_ ;
	wire _w3645_ ;
	wire _w3646_ ;
	wire _w3647_ ;
	wire _w3648_ ;
	wire _w3649_ ;
	wire _w3650_ ;
	wire _w3651_ ;
	wire _w3652_ ;
	wire _w3653_ ;
	wire _w3654_ ;
	wire _w3655_ ;
	wire _w3656_ ;
	wire _w3657_ ;
	wire _w3658_ ;
	wire _w3659_ ;
	wire _w3660_ ;
	wire _w3661_ ;
	wire _w3662_ ;
	wire _w3663_ ;
	wire _w3664_ ;
	wire _w3665_ ;
	wire _w3666_ ;
	wire _w3667_ ;
	wire _w3668_ ;
	wire _w3669_ ;
	wire _w3670_ ;
	wire _w3671_ ;
	wire _w3672_ ;
	wire _w3673_ ;
	wire _w3674_ ;
	wire _w3675_ ;
	wire _w3676_ ;
	wire _w3677_ ;
	wire _w3678_ ;
	wire _w3679_ ;
	wire _w3680_ ;
	wire _w3681_ ;
	wire _w3682_ ;
	wire _w3683_ ;
	wire _w3684_ ;
	wire _w3685_ ;
	wire _w3686_ ;
	wire _w3687_ ;
	wire _w3688_ ;
	wire _w3689_ ;
	wire _w3690_ ;
	wire _w3691_ ;
	wire _w3692_ ;
	wire _w3693_ ;
	wire _w3694_ ;
	wire _w3695_ ;
	wire _w3696_ ;
	wire _w3697_ ;
	wire _w3698_ ;
	wire _w3699_ ;
	wire _w3700_ ;
	wire _w3701_ ;
	wire _w3702_ ;
	wire _w3703_ ;
	wire _w3704_ ;
	wire _w3705_ ;
	wire _w3706_ ;
	wire _w3707_ ;
	wire _w3708_ ;
	wire _w3709_ ;
	wire _w3710_ ;
	wire _w3711_ ;
	wire _w3712_ ;
	wire _w3713_ ;
	wire _w3714_ ;
	wire _w3715_ ;
	wire _w3716_ ;
	wire _w3717_ ;
	wire _w3718_ ;
	wire _w3719_ ;
	wire _w3720_ ;
	wire _w3721_ ;
	wire _w3722_ ;
	wire _w3723_ ;
	wire _w3724_ ;
	wire _w3725_ ;
	wire _w3726_ ;
	wire _w3727_ ;
	wire _w3728_ ;
	wire _w3729_ ;
	wire _w3730_ ;
	wire _w3731_ ;
	wire _w3732_ ;
	wire _w3733_ ;
	wire _w3734_ ;
	wire _w3735_ ;
	wire _w3736_ ;
	wire _w3737_ ;
	wire _w3738_ ;
	wire _w3739_ ;
	wire _w3740_ ;
	wire _w3741_ ;
	wire _w3742_ ;
	wire _w3743_ ;
	wire _w3744_ ;
	wire _w3745_ ;
	wire _w3746_ ;
	wire _w3747_ ;
	wire _w3748_ ;
	wire _w3749_ ;
	wire _w3750_ ;
	wire _w3751_ ;
	wire _w3752_ ;
	wire _w3753_ ;
	wire _w3754_ ;
	wire _w3755_ ;
	wire _w3756_ ;
	wire _w3757_ ;
	wire _w3758_ ;
	wire _w3759_ ;
	wire _w3760_ ;
	wire _w3761_ ;
	wire _w3762_ ;
	wire _w3763_ ;
	wire _w3764_ ;
	wire _w3765_ ;
	wire _w3766_ ;
	wire _w3767_ ;
	wire _w3768_ ;
	wire _w3769_ ;
	wire _w3770_ ;
	wire _w3771_ ;
	wire _w3772_ ;
	wire _w3773_ ;
	wire _w3774_ ;
	wire _w3775_ ;
	wire _w3776_ ;
	wire _w3777_ ;
	wire _w3778_ ;
	wire _w3779_ ;
	wire _w3780_ ;
	wire _w3781_ ;
	wire _w3782_ ;
	wire _w3783_ ;
	wire _w3784_ ;
	wire _w3785_ ;
	wire _w3786_ ;
	wire _w3787_ ;
	wire _w3788_ ;
	wire _w3789_ ;
	wire _w3790_ ;
	wire _w3791_ ;
	wire _w3792_ ;
	wire _w3793_ ;
	wire _w3794_ ;
	wire _w3795_ ;
	wire _w3796_ ;
	wire _w3797_ ;
	wire _w3798_ ;
	wire _w3799_ ;
	wire _w3800_ ;
	wire _w3801_ ;
	wire _w3802_ ;
	wire _w3803_ ;
	wire _w3804_ ;
	wire _w3805_ ;
	wire _w3806_ ;
	wire _w3807_ ;
	wire _w3808_ ;
	wire _w3809_ ;
	wire _w3810_ ;
	wire _w3811_ ;
	wire _w3812_ ;
	wire _w3813_ ;
	wire _w3814_ ;
	wire _w3815_ ;
	wire _w3816_ ;
	wire _w3817_ ;
	wire _w3818_ ;
	wire _w3819_ ;
	wire _w3820_ ;
	wire _w3821_ ;
	wire _w3822_ ;
	wire _w3823_ ;
	wire _w3824_ ;
	wire _w3825_ ;
	wire _w3826_ ;
	wire _w3827_ ;
	wire _w3828_ ;
	wire _w3829_ ;
	wire _w3830_ ;
	wire _w3831_ ;
	wire _w3832_ ;
	wire _w3833_ ;
	wire _w3834_ ;
	wire _w3835_ ;
	wire _w3836_ ;
	wire _w3837_ ;
	wire _w3838_ ;
	wire _w3839_ ;
	wire _w3840_ ;
	wire _w3841_ ;
	wire _w3842_ ;
	wire _w3843_ ;
	wire _w3844_ ;
	wire _w3845_ ;
	wire _w3846_ ;
	wire _w3847_ ;
	wire _w3848_ ;
	wire _w3849_ ;
	wire _w3850_ ;
	wire _w3851_ ;
	wire _w3852_ ;
	wire _w3853_ ;
	wire _w3854_ ;
	wire _w3855_ ;
	wire _w3856_ ;
	wire _w3857_ ;
	wire _w3858_ ;
	wire _w3859_ ;
	wire _w3860_ ;
	wire _w3861_ ;
	wire _w3862_ ;
	wire _w3863_ ;
	wire _w3864_ ;
	wire _w3865_ ;
	wire _w3866_ ;
	wire _w3867_ ;
	wire _w3868_ ;
	wire _w3869_ ;
	wire _w3870_ ;
	wire _w3871_ ;
	wire _w3872_ ;
	wire _w3873_ ;
	wire _w3874_ ;
	wire _w3875_ ;
	wire _w3876_ ;
	wire _w3877_ ;
	wire _w3878_ ;
	wire _w3879_ ;
	wire _w3880_ ;
	wire _w3881_ ;
	wire _w3882_ ;
	wire _w3883_ ;
	wire _w3884_ ;
	wire _w3885_ ;
	wire _w3886_ ;
	wire _w3887_ ;
	wire _w3888_ ;
	wire _w3889_ ;
	wire _w3890_ ;
	wire _w3891_ ;
	wire _w3892_ ;
	wire _w3893_ ;
	wire _w3894_ ;
	wire _w3895_ ;
	wire _w3896_ ;
	wire _w3897_ ;
	wire _w3898_ ;
	wire _w3899_ ;
	wire _w3900_ ;
	wire _w3901_ ;
	wire _w3902_ ;
	wire _w3903_ ;
	wire _w3904_ ;
	wire _w3905_ ;
	wire _w3906_ ;
	wire _w3907_ ;
	wire _w3908_ ;
	wire _w3909_ ;
	wire _w3910_ ;
	wire _w3911_ ;
	wire _w3912_ ;
	wire _w3913_ ;
	wire _w3914_ ;
	wire _w3915_ ;
	wire _w3916_ ;
	wire _w3917_ ;
	wire _w3918_ ;
	wire _w3919_ ;
	wire _w3920_ ;
	wire _w3921_ ;
	wire _w3922_ ;
	wire _w3923_ ;
	wire _w3924_ ;
	wire _w3925_ ;
	wire _w3926_ ;
	wire _w3927_ ;
	wire _w3928_ ;
	wire _w3929_ ;
	wire _w3930_ ;
	wire _w3931_ ;
	wire _w3932_ ;
	wire _w3933_ ;
	wire _w3934_ ;
	wire _w3935_ ;
	wire _w3936_ ;
	wire _w3937_ ;
	wire _w3938_ ;
	wire _w3939_ ;
	wire _w3940_ ;
	wire _w3941_ ;
	wire _w3942_ ;
	wire _w3943_ ;
	wire _w3944_ ;
	wire _w3945_ ;
	wire _w3946_ ;
	wire _w3947_ ;
	wire _w3948_ ;
	wire _w3949_ ;
	wire _w3950_ ;
	wire _w3951_ ;
	wire _w3952_ ;
	wire _w3953_ ;
	wire _w3954_ ;
	wire _w3955_ ;
	wire _w3956_ ;
	wire _w3957_ ;
	wire _w3958_ ;
	wire _w3959_ ;
	wire _w3960_ ;
	wire _w3961_ ;
	wire _w3962_ ;
	wire _w3963_ ;
	wire _w3964_ ;
	wire _w3965_ ;
	wire _w3966_ ;
	wire _w3967_ ;
	wire _w3968_ ;
	wire _w3969_ ;
	wire _w3970_ ;
	wire _w3971_ ;
	wire _w3972_ ;
	wire _w3973_ ;
	wire _w3974_ ;
	wire _w3975_ ;
	wire _w3976_ ;
	wire _w3977_ ;
	wire _w3978_ ;
	wire _w3979_ ;
	wire _w3980_ ;
	wire _w3981_ ;
	wire _w3982_ ;
	wire _w3983_ ;
	wire _w3984_ ;
	wire _w3985_ ;
	wire _w3986_ ;
	wire _w3987_ ;
	wire _w3988_ ;
	wire _w3989_ ;
	wire _w3990_ ;
	wire _w3991_ ;
	wire _w3992_ ;
	wire _w3993_ ;
	wire _w3994_ ;
	wire _w3995_ ;
	wire _w3996_ ;
	wire _w3997_ ;
	wire _w3998_ ;
	wire _w3999_ ;
	wire _w4000_ ;
	wire _w4001_ ;
	wire _w4002_ ;
	wire _w4003_ ;
	wire _w4004_ ;
	wire _w4005_ ;
	wire _w4006_ ;
	wire _w4007_ ;
	wire _w4008_ ;
	wire _w4009_ ;
	wire _w4010_ ;
	wire _w4011_ ;
	wire _w4012_ ;
	wire _w4013_ ;
	wire _w4014_ ;
	wire _w4015_ ;
	wire _w4016_ ;
	wire _w4017_ ;
	wire _w4018_ ;
	wire _w4019_ ;
	wire _w4020_ ;
	wire _w4021_ ;
	wire _w4022_ ;
	wire _w4023_ ;
	wire _w4024_ ;
	wire _w4025_ ;
	wire _w4026_ ;
	wire _w4027_ ;
	wire _w4028_ ;
	wire _w4029_ ;
	wire _w4030_ ;
	wire _w4031_ ;
	wire _w4032_ ;
	wire _w4033_ ;
	wire _w4034_ ;
	wire _w4035_ ;
	wire _w4036_ ;
	wire _w4037_ ;
	wire _w4038_ ;
	wire _w4039_ ;
	wire _w4040_ ;
	wire _w4041_ ;
	wire _w4042_ ;
	wire _w4043_ ;
	wire _w4044_ ;
	wire _w4045_ ;
	wire _w4046_ ;
	wire _w4047_ ;
	wire _w4048_ ;
	wire _w4049_ ;
	wire _w4050_ ;
	wire _w4051_ ;
	wire _w4052_ ;
	wire _w4053_ ;
	wire _w4054_ ;
	wire _w4055_ ;
	wire _w4056_ ;
	wire _w4057_ ;
	wire _w4058_ ;
	wire _w4059_ ;
	wire _w4060_ ;
	wire _w4061_ ;
	wire _w4062_ ;
	wire _w4063_ ;
	wire _w4064_ ;
	wire _w4065_ ;
	wire _w4066_ ;
	wire _w4067_ ;
	wire _w4068_ ;
	wire _w4069_ ;
	wire _w4070_ ;
	wire _w4071_ ;
	wire _w4072_ ;
	wire _w4073_ ;
	wire _w4074_ ;
	wire _w4075_ ;
	wire _w4076_ ;
	wire _w4077_ ;
	wire _w4078_ ;
	wire _w4079_ ;
	wire _w4080_ ;
	wire _w4081_ ;
	wire _w4082_ ;
	wire _w4083_ ;
	wire _w4084_ ;
	wire _w4085_ ;
	wire _w4086_ ;
	wire _w4087_ ;
	wire _w4088_ ;
	wire _w4089_ ;
	wire _w4090_ ;
	wire _w4091_ ;
	wire _w4092_ ;
	wire _w4093_ ;
	wire _w4094_ ;
	wire _w4095_ ;
	wire _w4096_ ;
	wire _w4097_ ;
	wire _w4098_ ;
	wire _w4099_ ;
	wire _w4100_ ;
	wire _w4101_ ;
	wire _w4102_ ;
	wire _w4103_ ;
	wire _w4104_ ;
	wire _w4105_ ;
	wire _w4106_ ;
	wire _w4107_ ;
	wire _w4108_ ;
	wire _w4109_ ;
	wire _w4110_ ;
	wire _w4111_ ;
	wire _w4112_ ;
	wire _w4113_ ;
	wire _w4114_ ;
	wire _w4115_ ;
	wire _w4116_ ;
	wire _w4117_ ;
	wire _w4118_ ;
	wire _w4119_ ;
	wire _w4120_ ;
	wire _w4121_ ;
	wire _w4122_ ;
	wire _w4123_ ;
	wire _w4124_ ;
	wire _w4125_ ;
	wire _w4126_ ;
	wire _w4127_ ;
	wire _w4128_ ;
	wire _w4129_ ;
	wire _w4130_ ;
	wire _w4131_ ;
	wire _w4132_ ;
	wire _w4133_ ;
	wire _w4134_ ;
	wire _w4135_ ;
	wire _w4136_ ;
	wire _w4137_ ;
	wire _w4138_ ;
	wire _w4139_ ;
	wire _w4140_ ;
	wire _w4141_ ;
	wire _w4142_ ;
	wire _w4143_ ;
	wire _w4144_ ;
	wire _w4145_ ;
	wire _w4146_ ;
	wire _w4147_ ;
	wire _w4148_ ;
	wire _w4149_ ;
	wire _w4150_ ;
	wire _w4151_ ;
	wire _w4152_ ;
	wire _w4153_ ;
	wire _w4154_ ;
	wire _w4155_ ;
	wire _w4156_ ;
	wire _w4157_ ;
	wire _w4158_ ;
	wire _w4159_ ;
	wire _w4160_ ;
	wire _w4161_ ;
	wire _w4162_ ;
	wire _w4163_ ;
	wire _w4164_ ;
	wire _w4165_ ;
	wire _w4166_ ;
	wire _w4167_ ;
	wire _w4168_ ;
	wire _w4169_ ;
	wire _w4170_ ;
	wire _w4171_ ;
	wire _w4172_ ;
	wire _w4173_ ;
	wire _w4174_ ;
	wire _w4175_ ;
	wire _w4176_ ;
	wire _w4177_ ;
	wire _w4178_ ;
	wire _w4179_ ;
	wire _w4180_ ;
	wire _w4181_ ;
	wire _w4182_ ;
	wire _w4183_ ;
	wire _w4184_ ;
	wire _w4185_ ;
	wire _w4186_ ;
	wire _w4187_ ;
	wire _w4188_ ;
	wire _w4189_ ;
	wire _w4190_ ;
	wire _w4191_ ;
	wire _w4192_ ;
	wire _w4193_ ;
	wire _w4194_ ;
	wire _w4195_ ;
	wire _w4196_ ;
	wire _w4197_ ;
	wire _w4198_ ;
	wire _w4199_ ;
	wire _w4200_ ;
	wire _w4201_ ;
	wire _w4202_ ;
	wire _w4203_ ;
	wire _w4204_ ;
	wire _w4205_ ;
	wire _w4206_ ;
	wire _w4207_ ;
	wire _w4208_ ;
	wire _w4209_ ;
	wire _w4210_ ;
	wire _w4211_ ;
	wire _w4212_ ;
	wire _w4213_ ;
	wire _w4214_ ;
	wire _w4215_ ;
	wire _w4216_ ;
	wire _w4217_ ;
	wire _w4218_ ;
	wire _w4219_ ;
	wire _w4220_ ;
	wire _w4221_ ;
	wire _w4222_ ;
	wire _w4223_ ;
	wire _w4224_ ;
	wire _w4225_ ;
	wire _w4226_ ;
	wire _w4227_ ;
	wire _w4228_ ;
	wire _w4229_ ;
	wire _w4230_ ;
	wire _w4231_ ;
	wire _w4232_ ;
	wire _w4233_ ;
	wire _w4234_ ;
	wire _w4235_ ;
	wire _w4236_ ;
	wire _w4237_ ;
	wire _w4238_ ;
	wire _w4239_ ;
	wire _w4240_ ;
	wire _w4241_ ;
	wire _w4242_ ;
	wire _w4243_ ;
	wire _w4244_ ;
	wire _w4245_ ;
	wire _w4246_ ;
	wire _w4247_ ;
	wire _w4248_ ;
	wire _w4249_ ;
	wire _w4250_ ;
	wire _w4251_ ;
	wire _w4252_ ;
	wire _w4253_ ;
	wire _w4254_ ;
	wire _w4255_ ;
	wire _w4256_ ;
	wire _w4257_ ;
	wire _w4258_ ;
	wire _w4259_ ;
	wire _w4260_ ;
	wire _w4261_ ;
	wire _w4262_ ;
	wire _w4263_ ;
	wire _w4264_ ;
	wire _w4265_ ;
	wire _w4266_ ;
	wire _w4267_ ;
	wire _w4268_ ;
	wire _w4269_ ;
	wire _w4270_ ;
	wire _w4271_ ;
	wire _w4272_ ;
	wire _w4273_ ;
	wire _w4274_ ;
	wire _w4275_ ;
	wire _w4276_ ;
	wire _w4277_ ;
	wire _w4278_ ;
	wire _w4279_ ;
	wire _w4280_ ;
	wire _w4281_ ;
	wire _w4282_ ;
	wire _w4283_ ;
	wire _w4284_ ;
	wire _w4285_ ;
	wire _w4286_ ;
	wire _w4287_ ;
	wire _w4288_ ;
	wire _w4289_ ;
	wire _w4290_ ;
	wire _w4291_ ;
	wire _w4292_ ;
	wire _w4293_ ;
	wire _w4294_ ;
	wire _w4295_ ;
	wire _w4296_ ;
	wire _w4297_ ;
	wire _w4298_ ;
	wire _w4299_ ;
	wire _w4300_ ;
	wire _w4301_ ;
	wire _w4302_ ;
	wire _w4303_ ;
	wire _w4304_ ;
	wire _w4305_ ;
	wire _w4306_ ;
	wire _w4307_ ;
	wire _w4308_ ;
	wire _w4309_ ;
	wire _w4310_ ;
	wire _w4311_ ;
	wire _w4312_ ;
	wire _w4313_ ;
	wire _w4314_ ;
	wire _w4315_ ;
	wire _w4316_ ;
	wire _w4317_ ;
	wire _w4318_ ;
	wire _w4319_ ;
	wire _w4320_ ;
	wire _w4321_ ;
	wire _w4322_ ;
	wire _w4323_ ;
	wire _w4324_ ;
	wire _w4325_ ;
	wire _w4326_ ;
	wire _w4327_ ;
	wire _w4328_ ;
	wire _w4329_ ;
	wire _w4330_ ;
	wire _w4331_ ;
	wire _w4332_ ;
	wire _w4333_ ;
	wire _w4334_ ;
	wire _w4335_ ;
	wire _w4336_ ;
	wire _w4337_ ;
	wire _w4338_ ;
	wire _w4339_ ;
	wire _w4340_ ;
	wire _w4341_ ;
	wire _w4342_ ;
	wire _w4343_ ;
	wire _w4344_ ;
	wire _w4345_ ;
	wire _w4346_ ;
	wire _w4347_ ;
	wire _w4348_ ;
	wire _w4349_ ;
	wire _w4350_ ;
	wire _w4351_ ;
	wire _w4352_ ;
	wire _w4353_ ;
	wire _w4354_ ;
	wire _w4355_ ;
	wire _w4356_ ;
	wire _w4357_ ;
	wire _w4358_ ;
	wire _w4359_ ;
	wire _w4360_ ;
	wire _w4361_ ;
	wire _w4362_ ;
	wire _w4363_ ;
	wire _w4364_ ;
	wire _w4365_ ;
	wire _w4366_ ;
	wire _w4367_ ;
	wire _w4368_ ;
	wire _w4369_ ;
	wire _w4370_ ;
	wire _w4371_ ;
	wire _w4372_ ;
	wire _w4373_ ;
	wire _w4374_ ;
	wire _w4375_ ;
	wire _w4376_ ;
	wire _w4377_ ;
	wire _w4378_ ;
	wire _w4379_ ;
	wire _w4380_ ;
	wire _w4381_ ;
	wire _w4382_ ;
	wire _w4383_ ;
	wire _w4384_ ;
	wire _w4385_ ;
	wire _w4386_ ;
	wire _w4387_ ;
	wire _w4388_ ;
	wire _w4389_ ;
	wire _w4390_ ;
	wire _w4391_ ;
	wire _w4392_ ;
	wire _w4393_ ;
	wire _w4394_ ;
	wire _w4395_ ;
	wire _w4396_ ;
	wire _w4397_ ;
	wire _w4398_ ;
	wire _w4399_ ;
	wire _w4400_ ;
	wire _w4401_ ;
	wire _w4402_ ;
	wire _w4403_ ;
	wire _w4404_ ;
	wire _w4405_ ;
	wire _w4406_ ;
	wire _w4407_ ;
	wire _w4408_ ;
	wire _w4409_ ;
	wire _w4410_ ;
	wire _w4411_ ;
	wire _w4412_ ;
	wire _w4413_ ;
	wire _w4414_ ;
	wire _w4415_ ;
	wire _w4416_ ;
	wire _w4417_ ;
	wire _w4418_ ;
	wire _w4419_ ;
	wire _w4420_ ;
	wire _w4421_ ;
	wire _w4422_ ;
	wire _w4423_ ;
	wire _w4424_ ;
	wire _w4425_ ;
	wire _w4426_ ;
	wire _w4427_ ;
	wire _w4428_ ;
	wire _w4429_ ;
	wire _w4430_ ;
	wire _w4431_ ;
	wire _w4432_ ;
	wire _w4433_ ;
	wire _w4434_ ;
	wire _w4435_ ;
	wire _w4436_ ;
	wire _w4437_ ;
	wire _w4438_ ;
	wire _w4439_ ;
	wire _w4440_ ;
	wire _w4441_ ;
	wire _w4442_ ;
	wire _w4443_ ;
	wire _w4444_ ;
	wire _w4445_ ;
	wire _w4446_ ;
	wire _w4447_ ;
	wire _w4448_ ;
	wire _w4449_ ;
	wire _w4450_ ;
	wire _w4451_ ;
	wire _w4452_ ;
	wire _w4453_ ;
	wire _w4454_ ;
	wire _w4455_ ;
	wire _w4456_ ;
	wire _w4457_ ;
	wire _w4458_ ;
	wire _w4459_ ;
	wire _w4460_ ;
	wire _w4461_ ;
	wire _w4462_ ;
	wire _w4463_ ;
	wire _w4464_ ;
	wire _w4465_ ;
	wire _w4466_ ;
	wire _w4467_ ;
	wire _w4468_ ;
	wire _w4469_ ;
	wire _w4470_ ;
	wire _w4471_ ;
	wire _w4472_ ;
	wire _w4473_ ;
	wire _w4474_ ;
	wire _w4475_ ;
	wire _w4476_ ;
	wire _w4477_ ;
	wire _w4478_ ;
	wire _w4479_ ;
	wire _w4480_ ;
	wire _w4481_ ;
	wire _w4482_ ;
	wire _w4483_ ;
	wire _w4484_ ;
	wire _w4485_ ;
	wire _w4486_ ;
	wire _w4487_ ;
	wire _w4488_ ;
	wire _w4489_ ;
	wire _w4490_ ;
	wire _w4491_ ;
	wire _w4492_ ;
	wire _w4493_ ;
	wire _w4494_ ;
	wire _w4495_ ;
	wire _w4496_ ;
	wire _w4497_ ;
	wire _w4498_ ;
	wire _w4499_ ;
	wire _w4500_ ;
	wire _w4501_ ;
	wire _w4502_ ;
	wire _w4503_ ;
	LUT2 #(
		.INIT('h4)
	) name0 (
		\dma_ack_i[8]_pad ,
		\dma_req_o[8]_pad ,
		_w2147_
	);
	LUT4 #(
		.INIT('h0105)
	) name1 (
		\u11_status_reg[0]/P0001 ,
		\u11_status_reg[1]/P0001 ,
		\u13_icc_r_reg[20]/NET0131 ,
		\u13_icc_r_reg[21]/NET0131 ,
		_w2148_
	);
	LUT3 #(
		.INIT('h54)
	) name2 (
		\u11_full_reg/NET0131 ,
		\u11_status_reg[1]/P0001 ,
		\u13_icc_r_reg[21]/NET0131 ,
		_w2149_
	);
	LUT3 #(
		.INIT('h8a)
	) name3 (
		\u13_icc_r_reg[16]/NET0131 ,
		_w2148_,
		_w2149_,
		_w2150_
	);
	LUT2 #(
		.INIT('h4)
	) name4 (
		\dma_ack_i[8]_pad ,
		\u13_icc_r_reg[22]/NET0131 ,
		_w2151_
	);
	LUT4 #(
		.INIT('h8a00)
	) name5 (
		\u13_icc_r_reg[16]/NET0131 ,
		_w2148_,
		_w2149_,
		_w2151_,
		_w2152_
	);
	LUT3 #(
		.INIT('hec)
	) name6 (
		\u16_u8_dma_req_r1_reg/P0001 ,
		_w2147_,
		_w2152_,
		_w2153_
	);
	LUT2 #(
		.INIT('h8)
	) name7 (
		\u14_u5_en_out_l_reg/NET0131 ,
		\valid_s_reg/NET0131 ,
		_w2154_
	);
	LUT3 #(
		.INIT('h40)
	) name8 (
		\u14_u5_en_out_l2_reg/P0001 ,
		\u14_u5_en_out_l_reg/NET0131 ,
		\valid_s_reg/NET0131 ,
		_w2155_
	);
	LUT2 #(
		.INIT('h1)
	) name9 (
		\u13_occ1_r_reg[10]/NET0131 ,
		\u13_occ1_r_reg[11]/NET0131 ,
		_w2156_
	);
	LUT3 #(
		.INIT('h01)
	) name10 (
		\u13_occ1_r_reg[10]/NET0131 ,
		\u13_occ1_r_reg[11]/NET0131 ,
		\u8_rp_reg[0]/P0001 ,
		_w2157_
	);
	LUT2 #(
		.INIT('h8)
	) name11 (
		\u8_rp_reg[1]/NET0131 ,
		\u8_rp_reg[2]/NET0131 ,
		_w2158_
	);
	LUT3 #(
		.INIT('h20)
	) name12 (
		_w2155_,
		_w2157_,
		_w2158_,
		_w2159_
	);
	LUT3 #(
		.INIT('h28)
	) name13 (
		\u13_occ1_r_reg[8]/NET0131 ,
		\u8_rp_reg[3]/NET0131 ,
		_w2159_,
		_w2160_
	);
	LUT2 #(
		.INIT('h1)
	) name14 (
		\u0_slt0_r_reg[14]/P0001 ,
		\u2_ld_reg/P0001 ,
		_w2161_
	);
	LUT3 #(
		.INIT('h01)
	) name15 (
		\u14_u3_en_out_l_reg/NET0131 ,
		\u14_u4_en_out_l_reg/NET0131 ,
		\u14_u5_en_out_l_reg/NET0131 ,
		_w2162_
	);
	LUT2 #(
		.INIT('h4)
	) name16 (
		\u14_crac_wr_r_reg/P0001 ,
		\u2_ld_reg/P0001 ,
		_w2163_
	);
	LUT4 #(
		.INIT('h0001)
	) name17 (
		\u14_crac_valid_r_reg/P0001 ,
		\u14_u0_en_out_l_reg/NET0131 ,
		\u14_u1_en_out_l_reg/NET0131 ,
		\u14_u2_en_out_l_reg/NET0131 ,
		_w2164_
	);
	LUT4 #(
		.INIT('h1555)
	) name18 (
		_w2161_,
		_w2163_,
		_w2162_,
		_w2164_,
		_w2165_
	);
	LUT3 #(
		.INIT('hca)
	) name19 (
		\u0_slt0_r_reg[13]/P0001 ,
		\u14_crac_valid_r_reg/P0001 ,
		\u2_ld_reg/P0001 ,
		_w2166_
	);
	LUT3 #(
		.INIT('hca)
	) name20 (
		\u0_slt0_r_reg[12]/P0001 ,
		\u14_crac_wr_r_reg/P0001 ,
		\u2_ld_reg/P0001 ,
		_w2167_
	);
	LUT3 #(
		.INIT('hca)
	) name21 (
		\u0_slt0_r_reg[11]/P0001 ,
		\u14_u0_en_out_l_reg/NET0131 ,
		\u2_ld_reg/P0001 ,
		_w2168_
	);
	LUT3 #(
		.INIT('hca)
	) name22 (
		\u0_slt0_r_reg[10]/P0001 ,
		\u14_u1_en_out_l_reg/NET0131 ,
		\u2_ld_reg/P0001 ,
		_w2169_
	);
	LUT2 #(
		.INIT('h2)
	) name23 (
		\u0_slt0_r_reg[9]/P0001 ,
		\u2_ld_reg/P0001 ,
		_w2170_
	);
	LUT3 #(
		.INIT('hca)
	) name24 (
		\u0_slt0_r_reg[8]/P0001 ,
		\u14_u2_en_out_l_reg/NET0131 ,
		\u2_ld_reg/P0001 ,
		_w2171_
	);
	LUT3 #(
		.INIT('hca)
	) name25 (
		\u0_slt0_r_reg[7]/P0001 ,
		\u14_u3_en_out_l_reg/NET0131 ,
		\u2_ld_reg/P0001 ,
		_w2172_
	);
	LUT3 #(
		.INIT('hca)
	) name26 (
		\u0_slt0_r_reg[6]/P0001 ,
		\u14_u4_en_out_l_reg/NET0131 ,
		\u2_ld_reg/P0001 ,
		_w2173_
	);
	LUT3 #(
		.INIT('hca)
	) name27 (
		\u0_slt0_r_reg[5]/P0001 ,
		\u14_u5_en_out_l_reg/NET0131 ,
		\u2_ld_reg/P0001 ,
		_w2174_
	);
	LUT2 #(
		.INIT('h2)
	) name28 (
		\u0_slt0_r_reg[4]/P0001 ,
		\u2_ld_reg/P0001 ,
		_w2175_
	);
	LUT2 #(
		.INIT('h2)
	) name29 (
		\u0_slt0_r_reg[3]/P0001 ,
		\u2_ld_reg/P0001 ,
		_w2176_
	);
	LUT2 #(
		.INIT('h2)
	) name30 (
		\u0_slt0_r_reg[2]/P0001 ,
		\u2_ld_reg/P0001 ,
		_w2177_
	);
	LUT2 #(
		.INIT('h2)
	) name31 (
		\u0_slt0_r_reg[1]/P0001 ,
		\u2_ld_reg/P0001 ,
		_w2178_
	);
	LUT2 #(
		.INIT('h2)
	) name32 (
		\u0_slt0_r_reg[0]/P0001 ,
		\u2_ld_reg/P0001 ,
		_w2179_
	);
	LUT2 #(
		.INIT('h2)
	) name33 (
		\u0_slt1_r_reg[19]/P0001 ,
		\u2_ld_reg/P0001 ,
		_w2180_
	);
	LUT3 #(
		.INIT('hca)
	) name34 (
		\u0_slt1_r_reg[18]/P0001 ,
		\u13_crac_r_reg[7]/NET0131 ,
		\u2_ld_reg/P0001 ,
		_w2181_
	);
	LUT3 #(
		.INIT('hca)
	) name35 (
		\u0_slt1_r_reg[17]/P0001 ,
		\u13_crac_r_reg[6]/NET0131 ,
		\u2_ld_reg/P0001 ,
		_w2182_
	);
	LUT3 #(
		.INIT('hca)
	) name36 (
		\u0_slt1_r_reg[16]/P0001 ,
		\u13_crac_r_reg[5]/NET0131 ,
		\u2_ld_reg/P0001 ,
		_w2183_
	);
	LUT3 #(
		.INIT('hca)
	) name37 (
		\u0_slt1_r_reg[15]/P0001 ,
		\u13_crac_r_reg[4]/NET0131 ,
		\u2_ld_reg/P0001 ,
		_w2184_
	);
	LUT3 #(
		.INIT('hca)
	) name38 (
		\u0_slt1_r_reg[14]/P0001 ,
		\u13_crac_r_reg[3]/NET0131 ,
		\u2_ld_reg/P0001 ,
		_w2185_
	);
	LUT3 #(
		.INIT('hca)
	) name39 (
		\u0_slt1_r_reg[13]/P0001 ,
		\u13_crac_r_reg[2]/NET0131 ,
		\u2_ld_reg/P0001 ,
		_w2186_
	);
	LUT3 #(
		.INIT('hca)
	) name40 (
		\u0_slt1_r_reg[12]/P0001 ,
		\u13_crac_r_reg[1]/NET0131 ,
		\u2_ld_reg/P0001 ,
		_w2187_
	);
	LUT3 #(
		.INIT('hca)
	) name41 (
		\u0_slt1_r_reg[11]/P0001 ,
		\u13_crac_r_reg[0]/NET0131 ,
		\u2_ld_reg/P0001 ,
		_w2188_
	);
	LUT2 #(
		.INIT('h2)
	) name42 (
		\u0_slt1_r_reg[10]/P0001 ,
		\u2_ld_reg/P0001 ,
		_w2189_
	);
	LUT2 #(
		.INIT('h2)
	) name43 (
		\u0_slt1_r_reg[9]/P0001 ,
		\u2_ld_reg/P0001 ,
		_w2190_
	);
	LUT2 #(
		.INIT('h2)
	) name44 (
		\u0_slt1_r_reg[8]/P0001 ,
		\u2_ld_reg/P0001 ,
		_w2191_
	);
	LUT2 #(
		.INIT('h2)
	) name45 (
		\u0_slt1_r_reg[7]/P0001 ,
		\u2_ld_reg/P0001 ,
		_w2192_
	);
	LUT2 #(
		.INIT('h2)
	) name46 (
		\u0_slt1_r_reg[6]/P0001 ,
		\u2_ld_reg/P0001 ,
		_w2193_
	);
	LUT2 #(
		.INIT('h2)
	) name47 (
		\u0_slt1_r_reg[5]/P0001 ,
		\u2_ld_reg/P0001 ,
		_w2194_
	);
	LUT2 #(
		.INIT('h2)
	) name48 (
		\u0_slt1_r_reg[4]/P0001 ,
		\u2_ld_reg/P0001 ,
		_w2195_
	);
	LUT2 #(
		.INIT('h2)
	) name49 (
		\u0_slt1_r_reg[3]/P0001 ,
		\u2_ld_reg/P0001 ,
		_w2196_
	);
	LUT2 #(
		.INIT('h2)
	) name50 (
		\u0_slt1_r_reg[2]/P0001 ,
		\u2_ld_reg/P0001 ,
		_w2197_
	);
	LUT2 #(
		.INIT('h2)
	) name51 (
		\u0_slt1_r_reg[1]/P0001 ,
		\u2_ld_reg/P0001 ,
		_w2198_
	);
	LUT2 #(
		.INIT('h2)
	) name52 (
		\u0_slt1_r_reg[0]/P0001 ,
		\u2_ld_reg/P0001 ,
		_w2199_
	);
	LUT2 #(
		.INIT('h2)
	) name53 (
		\u0_slt2_r_reg[19]/P0001 ,
		\u2_ld_reg/P0001 ,
		_w2200_
	);
	LUT3 #(
		.INIT('hca)
	) name54 (
		\u0_slt2_r_reg[18]/P0001 ,
		\u13_crac_dout_r_reg[15]/P0001 ,
		\u2_ld_reg/P0001 ,
		_w2201_
	);
	LUT3 #(
		.INIT('hca)
	) name55 (
		\u0_slt2_r_reg[17]/P0001 ,
		\u13_crac_dout_r_reg[14]/P0001 ,
		\u2_ld_reg/P0001 ,
		_w2202_
	);
	LUT3 #(
		.INIT('hca)
	) name56 (
		\u0_slt2_r_reg[16]/P0001 ,
		\u13_crac_dout_r_reg[13]/P0001 ,
		\u2_ld_reg/P0001 ,
		_w2203_
	);
	LUT3 #(
		.INIT('hca)
	) name57 (
		\u0_slt2_r_reg[15]/P0001 ,
		\u13_crac_dout_r_reg[12]/P0001 ,
		\u2_ld_reg/P0001 ,
		_w2204_
	);
	LUT3 #(
		.INIT('hca)
	) name58 (
		\u0_slt2_r_reg[14]/P0001 ,
		\u13_crac_dout_r_reg[11]/P0001 ,
		\u2_ld_reg/P0001 ,
		_w2205_
	);
	LUT3 #(
		.INIT('hca)
	) name59 (
		\u0_slt2_r_reg[13]/P0001 ,
		\u13_crac_dout_r_reg[10]/P0001 ,
		\u2_ld_reg/P0001 ,
		_w2206_
	);
	LUT3 #(
		.INIT('hca)
	) name60 (
		\u0_slt2_r_reg[12]/P0001 ,
		\u13_crac_dout_r_reg[9]/P0001 ,
		\u2_ld_reg/P0001 ,
		_w2207_
	);
	LUT3 #(
		.INIT('hca)
	) name61 (
		\u0_slt2_r_reg[11]/P0001 ,
		\u13_crac_dout_r_reg[8]/P0001 ,
		\u2_ld_reg/P0001 ,
		_w2208_
	);
	LUT3 #(
		.INIT('hca)
	) name62 (
		\u0_slt2_r_reg[10]/P0001 ,
		\u13_crac_dout_r_reg[7]/P0001 ,
		\u2_ld_reg/P0001 ,
		_w2209_
	);
	LUT3 #(
		.INIT('hca)
	) name63 (
		\u0_slt2_r_reg[9]/P0001 ,
		\u13_crac_dout_r_reg[6]/P0001 ,
		\u2_ld_reg/P0001 ,
		_w2210_
	);
	LUT3 #(
		.INIT('hca)
	) name64 (
		\u0_slt2_r_reg[8]/P0001 ,
		\u13_crac_dout_r_reg[5]/P0001 ,
		\u2_ld_reg/P0001 ,
		_w2211_
	);
	LUT3 #(
		.INIT('hca)
	) name65 (
		\u0_slt2_r_reg[7]/P0001 ,
		\u13_crac_dout_r_reg[4]/P0001 ,
		\u2_ld_reg/P0001 ,
		_w2212_
	);
	LUT3 #(
		.INIT('hca)
	) name66 (
		\u0_slt2_r_reg[6]/P0001 ,
		\u13_crac_dout_r_reg[3]/P0001 ,
		\u2_ld_reg/P0001 ,
		_w2213_
	);
	LUT3 #(
		.INIT('hca)
	) name67 (
		\u0_slt2_r_reg[5]/P0001 ,
		\u13_crac_dout_r_reg[2]/P0001 ,
		\u2_ld_reg/P0001 ,
		_w2214_
	);
	LUT3 #(
		.INIT('hca)
	) name68 (
		\u0_slt2_r_reg[4]/P0001 ,
		\u13_crac_dout_r_reg[1]/P0001 ,
		\u2_ld_reg/P0001 ,
		_w2215_
	);
	LUT3 #(
		.INIT('hca)
	) name69 (
		\u0_slt2_r_reg[3]/P0001 ,
		\u13_crac_dout_r_reg[0]/P0001 ,
		\u2_ld_reg/P0001 ,
		_w2216_
	);
	LUT2 #(
		.INIT('h2)
	) name70 (
		\u0_slt2_r_reg[2]/P0001 ,
		\u2_ld_reg/P0001 ,
		_w2217_
	);
	LUT2 #(
		.INIT('h2)
	) name71 (
		\u0_slt2_r_reg[1]/P0001 ,
		\u2_ld_reg/P0001 ,
		_w2218_
	);
	LUT2 #(
		.INIT('h2)
	) name72 (
		\u0_slt2_r_reg[0]/P0001 ,
		\u2_ld_reg/P0001 ,
		_w2219_
	);
	LUT2 #(
		.INIT('h2)
	) name73 (
		\u0_slt3_r_reg[19]/P0001 ,
		\u2_ld_reg/P0001 ,
		_w2220_
	);
	LUT3 #(
		.INIT('he2)
	) name74 (
		\u0_slt3_r_reg[18]/P0001 ,
		\u2_ld_reg/P0001 ,
		\u3_dout_reg[19]/P0001 ,
		_w2221_
	);
	LUT3 #(
		.INIT('he2)
	) name75 (
		\u0_slt3_r_reg[17]/P0001 ,
		\u2_ld_reg/P0001 ,
		\u3_dout_reg[18]/P0001 ,
		_w2222_
	);
	LUT3 #(
		.INIT('he2)
	) name76 (
		\u0_slt3_r_reg[16]/P0001 ,
		\u2_ld_reg/P0001 ,
		\u3_dout_reg[17]/P0001 ,
		_w2223_
	);
	LUT3 #(
		.INIT('he2)
	) name77 (
		\u0_slt3_r_reg[15]/P0001 ,
		\u2_ld_reg/P0001 ,
		\u3_dout_reg[16]/P0001 ,
		_w2224_
	);
	LUT3 #(
		.INIT('he2)
	) name78 (
		\u0_slt3_r_reg[14]/P0001 ,
		\u2_ld_reg/P0001 ,
		\u3_dout_reg[15]/P0001 ,
		_w2225_
	);
	LUT3 #(
		.INIT('he2)
	) name79 (
		\u0_slt3_r_reg[13]/P0001 ,
		\u2_ld_reg/P0001 ,
		\u3_dout_reg[14]/P0001 ,
		_w2226_
	);
	LUT3 #(
		.INIT('he2)
	) name80 (
		\u0_slt3_r_reg[12]/P0001 ,
		\u2_ld_reg/P0001 ,
		\u3_dout_reg[13]/P0001 ,
		_w2227_
	);
	LUT3 #(
		.INIT('he2)
	) name81 (
		\u0_slt3_r_reg[11]/P0001 ,
		\u2_ld_reg/P0001 ,
		\u3_dout_reg[12]/P0001 ,
		_w2228_
	);
	LUT3 #(
		.INIT('he2)
	) name82 (
		\u0_slt3_r_reg[10]/P0001 ,
		\u2_ld_reg/P0001 ,
		\u3_dout_reg[11]/P0001 ,
		_w2229_
	);
	LUT3 #(
		.INIT('he2)
	) name83 (
		\u0_slt3_r_reg[9]/P0001 ,
		\u2_ld_reg/P0001 ,
		\u3_dout_reg[10]/P0001 ,
		_w2230_
	);
	LUT3 #(
		.INIT('he2)
	) name84 (
		\u0_slt3_r_reg[8]/P0001 ,
		\u2_ld_reg/P0001 ,
		\u3_dout_reg[9]/P0001 ,
		_w2231_
	);
	LUT3 #(
		.INIT('he2)
	) name85 (
		\u0_slt3_r_reg[7]/P0001 ,
		\u2_ld_reg/P0001 ,
		\u3_dout_reg[8]/P0001 ,
		_w2232_
	);
	LUT3 #(
		.INIT('he2)
	) name86 (
		\u0_slt3_r_reg[6]/P0001 ,
		\u2_ld_reg/P0001 ,
		\u3_dout_reg[7]/P0001 ,
		_w2233_
	);
	LUT3 #(
		.INIT('he2)
	) name87 (
		\u0_slt3_r_reg[5]/P0001 ,
		\u2_ld_reg/P0001 ,
		\u3_dout_reg[6]/P0001 ,
		_w2234_
	);
	LUT3 #(
		.INIT('he2)
	) name88 (
		\u0_slt3_r_reg[4]/P0001 ,
		\u2_ld_reg/P0001 ,
		\u3_dout_reg[5]/P0001 ,
		_w2235_
	);
	LUT3 #(
		.INIT('he2)
	) name89 (
		\u0_slt3_r_reg[3]/P0001 ,
		\u2_ld_reg/P0001 ,
		\u3_dout_reg[4]/P0001 ,
		_w2236_
	);
	LUT3 #(
		.INIT('he2)
	) name90 (
		\u0_slt3_r_reg[2]/P0001 ,
		\u2_ld_reg/P0001 ,
		\u3_dout_reg[3]/P0001 ,
		_w2237_
	);
	LUT3 #(
		.INIT('he2)
	) name91 (
		\u0_slt3_r_reg[1]/P0001 ,
		\u2_ld_reg/P0001 ,
		\u3_dout_reg[2]/P0001 ,
		_w2238_
	);
	LUT3 #(
		.INIT('he2)
	) name92 (
		\u0_slt3_r_reg[0]/P0001 ,
		\u2_ld_reg/P0001 ,
		\u3_dout_reg[1]/P0001 ,
		_w2239_
	);
	LUT3 #(
		.INIT('he2)
	) name93 (
		\u0_slt4_r_reg[19]/P0001 ,
		\u2_ld_reg/P0001 ,
		\u3_dout_reg[0]/P0001 ,
		_w2240_
	);
	LUT3 #(
		.INIT('he2)
	) name94 (
		\u0_slt4_r_reg[18]/P0001 ,
		\u2_ld_reg/P0001 ,
		\u4_dout_reg[19]/P0001 ,
		_w2241_
	);
	LUT3 #(
		.INIT('he2)
	) name95 (
		\u0_slt4_r_reg[17]/P0001 ,
		\u2_ld_reg/P0001 ,
		\u4_dout_reg[18]/P0001 ,
		_w2242_
	);
	LUT3 #(
		.INIT('he2)
	) name96 (
		\u0_slt4_r_reg[16]/P0001 ,
		\u2_ld_reg/P0001 ,
		\u4_dout_reg[17]/P0001 ,
		_w2243_
	);
	LUT3 #(
		.INIT('he2)
	) name97 (
		\u0_slt4_r_reg[15]/P0001 ,
		\u2_ld_reg/P0001 ,
		\u4_dout_reg[16]/P0001 ,
		_w2244_
	);
	LUT3 #(
		.INIT('he2)
	) name98 (
		\u0_slt4_r_reg[14]/P0001 ,
		\u2_ld_reg/P0001 ,
		\u4_dout_reg[15]/P0001 ,
		_w2245_
	);
	LUT3 #(
		.INIT('he2)
	) name99 (
		\u0_slt4_r_reg[13]/P0001 ,
		\u2_ld_reg/P0001 ,
		\u4_dout_reg[14]/P0001 ,
		_w2246_
	);
	LUT3 #(
		.INIT('he2)
	) name100 (
		\u0_slt4_r_reg[12]/P0001 ,
		\u2_ld_reg/P0001 ,
		\u4_dout_reg[13]/P0001 ,
		_w2247_
	);
	LUT3 #(
		.INIT('he2)
	) name101 (
		\u0_slt4_r_reg[11]/P0001 ,
		\u2_ld_reg/P0001 ,
		\u4_dout_reg[12]/P0001 ,
		_w2248_
	);
	LUT3 #(
		.INIT('he2)
	) name102 (
		\u0_slt4_r_reg[10]/P0001 ,
		\u2_ld_reg/P0001 ,
		\u4_dout_reg[11]/P0001 ,
		_w2249_
	);
	LUT3 #(
		.INIT('he2)
	) name103 (
		\u0_slt4_r_reg[9]/P0001 ,
		\u2_ld_reg/P0001 ,
		\u4_dout_reg[10]/P0001 ,
		_w2250_
	);
	LUT3 #(
		.INIT('he2)
	) name104 (
		\u0_slt4_r_reg[8]/P0001 ,
		\u2_ld_reg/P0001 ,
		\u4_dout_reg[9]/P0001 ,
		_w2251_
	);
	LUT3 #(
		.INIT('he2)
	) name105 (
		\u0_slt4_r_reg[7]/P0001 ,
		\u2_ld_reg/P0001 ,
		\u4_dout_reg[8]/P0001 ,
		_w2252_
	);
	LUT3 #(
		.INIT('he2)
	) name106 (
		\u0_slt4_r_reg[6]/P0001 ,
		\u2_ld_reg/P0001 ,
		\u4_dout_reg[7]/P0001 ,
		_w2253_
	);
	LUT3 #(
		.INIT('he2)
	) name107 (
		\u0_slt4_r_reg[5]/P0001 ,
		\u2_ld_reg/P0001 ,
		\u4_dout_reg[6]/P0001 ,
		_w2254_
	);
	LUT3 #(
		.INIT('he2)
	) name108 (
		\u0_slt4_r_reg[4]/P0001 ,
		\u2_ld_reg/P0001 ,
		\u4_dout_reg[5]/P0001 ,
		_w2255_
	);
	LUT3 #(
		.INIT('he2)
	) name109 (
		\u0_slt4_r_reg[3]/P0001 ,
		\u2_ld_reg/P0001 ,
		\u4_dout_reg[4]/P0001 ,
		_w2256_
	);
	LUT3 #(
		.INIT('he2)
	) name110 (
		\u0_slt4_r_reg[2]/P0001 ,
		\u2_ld_reg/P0001 ,
		\u4_dout_reg[3]/P0001 ,
		_w2257_
	);
	LUT3 #(
		.INIT('he2)
	) name111 (
		\u0_slt4_r_reg[1]/P0001 ,
		\u2_ld_reg/P0001 ,
		\u4_dout_reg[2]/P0001 ,
		_w2258_
	);
	LUT3 #(
		.INIT('he2)
	) name112 (
		\u0_slt4_r_reg[0]/P0001 ,
		\u2_ld_reg/P0001 ,
		\u4_dout_reg[1]/P0001 ,
		_w2259_
	);
	LUT3 #(
		.INIT('he2)
	) name113 (
		\u0_slt5_r_reg[19]/P0001 ,
		\u2_ld_reg/P0001 ,
		\u4_dout_reg[0]/P0001 ,
		_w2260_
	);
	LUT2 #(
		.INIT('h2)
	) name114 (
		\u0_slt5_r_reg[18]/P0001 ,
		\u2_ld_reg/P0001 ,
		_w2261_
	);
	LUT2 #(
		.INIT('h2)
	) name115 (
		\u0_slt5_r_reg[17]/P0001 ,
		\u2_ld_reg/P0001 ,
		_w2262_
	);
	LUT2 #(
		.INIT('h2)
	) name116 (
		\u0_slt5_r_reg[16]/P0001 ,
		\u2_ld_reg/P0001 ,
		_w2263_
	);
	LUT2 #(
		.INIT('h2)
	) name117 (
		\u0_slt5_r_reg[15]/P0001 ,
		\u2_ld_reg/P0001 ,
		_w2264_
	);
	LUT2 #(
		.INIT('h2)
	) name118 (
		\u0_slt5_r_reg[14]/P0001 ,
		\u2_ld_reg/P0001 ,
		_w2265_
	);
	LUT2 #(
		.INIT('h2)
	) name119 (
		\u0_slt5_r_reg[13]/P0001 ,
		\u2_ld_reg/P0001 ,
		_w2266_
	);
	LUT2 #(
		.INIT('h2)
	) name120 (
		\u0_slt5_r_reg[12]/P0001 ,
		\u2_ld_reg/P0001 ,
		_w2267_
	);
	LUT2 #(
		.INIT('h2)
	) name121 (
		\u0_slt5_r_reg[11]/P0001 ,
		\u2_ld_reg/P0001 ,
		_w2268_
	);
	LUT2 #(
		.INIT('h2)
	) name122 (
		\u0_slt5_r_reg[10]/P0001 ,
		\u2_ld_reg/P0001 ,
		_w2269_
	);
	LUT2 #(
		.INIT('h2)
	) name123 (
		\u0_slt5_r_reg[9]/P0001 ,
		\u2_ld_reg/P0001 ,
		_w2270_
	);
	LUT2 #(
		.INIT('h2)
	) name124 (
		\u0_slt5_r_reg[8]/P0001 ,
		\u2_ld_reg/P0001 ,
		_w2271_
	);
	LUT2 #(
		.INIT('h2)
	) name125 (
		\u0_slt5_r_reg[7]/P0001 ,
		\u2_ld_reg/P0001 ,
		_w2272_
	);
	LUT2 #(
		.INIT('h2)
	) name126 (
		\u0_slt5_r_reg[6]/P0001 ,
		\u2_ld_reg/P0001 ,
		_w2273_
	);
	LUT2 #(
		.INIT('h2)
	) name127 (
		\u0_slt5_r_reg[5]/P0001 ,
		\u2_ld_reg/P0001 ,
		_w2274_
	);
	LUT2 #(
		.INIT('h2)
	) name128 (
		\u0_slt5_r_reg[4]/P0001 ,
		\u2_ld_reg/P0001 ,
		_w2275_
	);
	LUT2 #(
		.INIT('h2)
	) name129 (
		\u0_slt5_r_reg[3]/P0001 ,
		\u2_ld_reg/P0001 ,
		_w2276_
	);
	LUT2 #(
		.INIT('h2)
	) name130 (
		\u0_slt5_r_reg[2]/P0001 ,
		\u2_ld_reg/P0001 ,
		_w2277_
	);
	LUT2 #(
		.INIT('h2)
	) name131 (
		\u0_slt5_r_reg[1]/P0001 ,
		\u2_ld_reg/P0001 ,
		_w2278_
	);
	LUT2 #(
		.INIT('h2)
	) name132 (
		\u0_slt5_r_reg[0]/P0001 ,
		\u2_ld_reg/P0001 ,
		_w2279_
	);
	LUT2 #(
		.INIT('h2)
	) name133 (
		\u0_slt6_r_reg[19]/P0001 ,
		\u2_ld_reg/P0001 ,
		_w2280_
	);
	LUT3 #(
		.INIT('he2)
	) name134 (
		\u0_slt6_r_reg[18]/P0001 ,
		\u2_ld_reg/P0001 ,
		\u5_dout_reg[19]/P0001 ,
		_w2281_
	);
	LUT3 #(
		.INIT('he2)
	) name135 (
		\u0_slt6_r_reg[17]/P0001 ,
		\u2_ld_reg/P0001 ,
		\u5_dout_reg[18]/P0001 ,
		_w2282_
	);
	LUT3 #(
		.INIT('he2)
	) name136 (
		\u0_slt6_r_reg[16]/P0001 ,
		\u2_ld_reg/P0001 ,
		\u5_dout_reg[17]/P0001 ,
		_w2283_
	);
	LUT3 #(
		.INIT('he2)
	) name137 (
		\u0_slt6_r_reg[15]/P0001 ,
		\u2_ld_reg/P0001 ,
		\u5_dout_reg[16]/P0001 ,
		_w2284_
	);
	LUT3 #(
		.INIT('he2)
	) name138 (
		\u0_slt6_r_reg[14]/P0001 ,
		\u2_ld_reg/P0001 ,
		\u5_dout_reg[15]/P0001 ,
		_w2285_
	);
	LUT3 #(
		.INIT('he2)
	) name139 (
		\u0_slt6_r_reg[13]/P0001 ,
		\u2_ld_reg/P0001 ,
		\u5_dout_reg[14]/P0001 ,
		_w2286_
	);
	LUT3 #(
		.INIT('he2)
	) name140 (
		\u0_slt6_r_reg[12]/P0001 ,
		\u2_ld_reg/P0001 ,
		\u5_dout_reg[13]/P0001 ,
		_w2287_
	);
	LUT3 #(
		.INIT('he2)
	) name141 (
		\u0_slt6_r_reg[11]/P0001 ,
		\u2_ld_reg/P0001 ,
		\u5_dout_reg[12]/P0001 ,
		_w2288_
	);
	LUT3 #(
		.INIT('he2)
	) name142 (
		\u0_slt6_r_reg[10]/P0001 ,
		\u2_ld_reg/P0001 ,
		\u5_dout_reg[11]/P0001 ,
		_w2289_
	);
	LUT3 #(
		.INIT('he2)
	) name143 (
		\u0_slt6_r_reg[9]/P0001 ,
		\u2_ld_reg/P0001 ,
		\u5_dout_reg[10]/P0001 ,
		_w2290_
	);
	LUT3 #(
		.INIT('he2)
	) name144 (
		\u0_slt6_r_reg[8]/P0001 ,
		\u2_ld_reg/P0001 ,
		\u5_dout_reg[9]/P0001 ,
		_w2291_
	);
	LUT3 #(
		.INIT('he2)
	) name145 (
		\u0_slt6_r_reg[7]/P0001 ,
		\u2_ld_reg/P0001 ,
		\u5_dout_reg[8]/P0001 ,
		_w2292_
	);
	LUT3 #(
		.INIT('he2)
	) name146 (
		\u0_slt6_r_reg[6]/P0001 ,
		\u2_ld_reg/P0001 ,
		\u5_dout_reg[7]/P0001 ,
		_w2293_
	);
	LUT3 #(
		.INIT('he2)
	) name147 (
		\u0_slt6_r_reg[5]/P0001 ,
		\u2_ld_reg/P0001 ,
		\u5_dout_reg[6]/P0001 ,
		_w2294_
	);
	LUT3 #(
		.INIT('he2)
	) name148 (
		\u0_slt6_r_reg[4]/P0001 ,
		\u2_ld_reg/P0001 ,
		\u5_dout_reg[5]/P0001 ,
		_w2295_
	);
	LUT3 #(
		.INIT('he2)
	) name149 (
		\u0_slt6_r_reg[3]/P0001 ,
		\u2_ld_reg/P0001 ,
		\u5_dout_reg[4]/P0001 ,
		_w2296_
	);
	LUT3 #(
		.INIT('he2)
	) name150 (
		\u0_slt6_r_reg[2]/P0001 ,
		\u2_ld_reg/P0001 ,
		\u5_dout_reg[3]/P0001 ,
		_w2297_
	);
	LUT3 #(
		.INIT('he2)
	) name151 (
		\u0_slt6_r_reg[1]/P0001 ,
		\u2_ld_reg/P0001 ,
		\u5_dout_reg[2]/P0001 ,
		_w2298_
	);
	LUT3 #(
		.INIT('he2)
	) name152 (
		\u0_slt6_r_reg[0]/P0001 ,
		\u2_ld_reg/P0001 ,
		\u5_dout_reg[1]/P0001 ,
		_w2299_
	);
	LUT3 #(
		.INIT('he2)
	) name153 (
		\u0_slt7_r_reg[19]/P0001 ,
		\u2_ld_reg/P0001 ,
		\u5_dout_reg[0]/P0001 ,
		_w2300_
	);
	LUT3 #(
		.INIT('he2)
	) name154 (
		\u0_slt7_r_reg[18]/P0001 ,
		\u2_ld_reg/P0001 ,
		\u6_dout_reg[19]/P0001 ,
		_w2301_
	);
	LUT3 #(
		.INIT('he2)
	) name155 (
		\u0_slt7_r_reg[17]/P0001 ,
		\u2_ld_reg/P0001 ,
		\u6_dout_reg[18]/P0001 ,
		_w2302_
	);
	LUT3 #(
		.INIT('he2)
	) name156 (
		\u0_slt7_r_reg[16]/P0001 ,
		\u2_ld_reg/P0001 ,
		\u6_dout_reg[17]/P0001 ,
		_w2303_
	);
	LUT3 #(
		.INIT('he2)
	) name157 (
		\u0_slt7_r_reg[15]/P0001 ,
		\u2_ld_reg/P0001 ,
		\u6_dout_reg[16]/P0001 ,
		_w2304_
	);
	LUT3 #(
		.INIT('he2)
	) name158 (
		\u0_slt7_r_reg[14]/P0001 ,
		\u2_ld_reg/P0001 ,
		\u6_dout_reg[15]/P0001 ,
		_w2305_
	);
	LUT3 #(
		.INIT('he2)
	) name159 (
		\u0_slt7_r_reg[13]/P0001 ,
		\u2_ld_reg/P0001 ,
		\u6_dout_reg[14]/P0001 ,
		_w2306_
	);
	LUT3 #(
		.INIT('he2)
	) name160 (
		\u0_slt7_r_reg[12]/P0001 ,
		\u2_ld_reg/P0001 ,
		\u6_dout_reg[13]/P0001 ,
		_w2307_
	);
	LUT3 #(
		.INIT('he2)
	) name161 (
		\u0_slt7_r_reg[11]/P0001 ,
		\u2_ld_reg/P0001 ,
		\u6_dout_reg[12]/P0001 ,
		_w2308_
	);
	LUT3 #(
		.INIT('he2)
	) name162 (
		\u0_slt7_r_reg[10]/P0001 ,
		\u2_ld_reg/P0001 ,
		\u6_dout_reg[11]/P0001 ,
		_w2309_
	);
	LUT3 #(
		.INIT('he2)
	) name163 (
		\u0_slt7_r_reg[9]/P0001 ,
		\u2_ld_reg/P0001 ,
		\u6_dout_reg[10]/P0001 ,
		_w2310_
	);
	LUT3 #(
		.INIT('he2)
	) name164 (
		\u0_slt7_r_reg[8]/P0001 ,
		\u2_ld_reg/P0001 ,
		\u6_dout_reg[9]/P0001 ,
		_w2311_
	);
	LUT3 #(
		.INIT('he2)
	) name165 (
		\u0_slt7_r_reg[7]/P0001 ,
		\u2_ld_reg/P0001 ,
		\u6_dout_reg[8]/P0001 ,
		_w2312_
	);
	LUT3 #(
		.INIT('he2)
	) name166 (
		\u0_slt7_r_reg[6]/P0001 ,
		\u2_ld_reg/P0001 ,
		\u6_dout_reg[7]/P0001 ,
		_w2313_
	);
	LUT3 #(
		.INIT('he2)
	) name167 (
		\u0_slt7_r_reg[5]/P0001 ,
		\u2_ld_reg/P0001 ,
		\u6_dout_reg[6]/P0001 ,
		_w2314_
	);
	LUT3 #(
		.INIT('he2)
	) name168 (
		\u0_slt7_r_reg[4]/P0001 ,
		\u2_ld_reg/P0001 ,
		\u6_dout_reg[5]/P0001 ,
		_w2315_
	);
	LUT3 #(
		.INIT('he2)
	) name169 (
		\u0_slt7_r_reg[3]/P0001 ,
		\u2_ld_reg/P0001 ,
		\u6_dout_reg[4]/P0001 ,
		_w2316_
	);
	LUT3 #(
		.INIT('he2)
	) name170 (
		\u0_slt7_r_reg[2]/P0001 ,
		\u2_ld_reg/P0001 ,
		\u6_dout_reg[3]/P0001 ,
		_w2317_
	);
	LUT3 #(
		.INIT('he2)
	) name171 (
		\u0_slt7_r_reg[1]/P0001 ,
		\u2_ld_reg/P0001 ,
		\u6_dout_reg[2]/P0001 ,
		_w2318_
	);
	LUT3 #(
		.INIT('he2)
	) name172 (
		\u0_slt7_r_reg[0]/P0001 ,
		\u2_ld_reg/P0001 ,
		\u6_dout_reg[1]/P0001 ,
		_w2319_
	);
	LUT3 #(
		.INIT('he2)
	) name173 (
		\u0_slt8_r_reg[19]/P0001 ,
		\u2_ld_reg/P0001 ,
		\u6_dout_reg[0]/P0001 ,
		_w2320_
	);
	LUT3 #(
		.INIT('he2)
	) name174 (
		\u0_slt8_r_reg[18]/P0001 ,
		\u2_ld_reg/P0001 ,
		\u7_dout_reg[19]/P0001 ,
		_w2321_
	);
	LUT3 #(
		.INIT('he2)
	) name175 (
		\u0_slt8_r_reg[17]/P0001 ,
		\u2_ld_reg/P0001 ,
		\u7_dout_reg[18]/P0001 ,
		_w2322_
	);
	LUT3 #(
		.INIT('he2)
	) name176 (
		\u0_slt8_r_reg[16]/P0001 ,
		\u2_ld_reg/P0001 ,
		\u7_dout_reg[17]/P0001 ,
		_w2323_
	);
	LUT3 #(
		.INIT('he2)
	) name177 (
		\u0_slt8_r_reg[15]/P0001 ,
		\u2_ld_reg/P0001 ,
		\u7_dout_reg[16]/P0001 ,
		_w2324_
	);
	LUT3 #(
		.INIT('he2)
	) name178 (
		\u0_slt8_r_reg[14]/P0001 ,
		\u2_ld_reg/P0001 ,
		\u7_dout_reg[15]/P0001 ,
		_w2325_
	);
	LUT3 #(
		.INIT('he2)
	) name179 (
		\u0_slt8_r_reg[13]/P0001 ,
		\u2_ld_reg/P0001 ,
		\u7_dout_reg[14]/P0001 ,
		_w2326_
	);
	LUT3 #(
		.INIT('he2)
	) name180 (
		\u0_slt8_r_reg[12]/P0001 ,
		\u2_ld_reg/P0001 ,
		\u7_dout_reg[13]/P0001 ,
		_w2327_
	);
	LUT3 #(
		.INIT('he2)
	) name181 (
		\u0_slt8_r_reg[11]/P0001 ,
		\u2_ld_reg/P0001 ,
		\u7_dout_reg[12]/P0001 ,
		_w2328_
	);
	LUT3 #(
		.INIT('he2)
	) name182 (
		\u0_slt8_r_reg[10]/P0001 ,
		\u2_ld_reg/P0001 ,
		\u7_dout_reg[11]/P0001 ,
		_w2329_
	);
	LUT3 #(
		.INIT('he2)
	) name183 (
		\u0_slt8_r_reg[9]/P0001 ,
		\u2_ld_reg/P0001 ,
		\u7_dout_reg[10]/P0001 ,
		_w2330_
	);
	LUT3 #(
		.INIT('he2)
	) name184 (
		\u0_slt8_r_reg[8]/P0001 ,
		\u2_ld_reg/P0001 ,
		\u7_dout_reg[9]/P0001 ,
		_w2331_
	);
	LUT3 #(
		.INIT('he2)
	) name185 (
		\u0_slt8_r_reg[7]/P0001 ,
		\u2_ld_reg/P0001 ,
		\u7_dout_reg[8]/P0001 ,
		_w2332_
	);
	LUT3 #(
		.INIT('he2)
	) name186 (
		\u0_slt8_r_reg[6]/P0001 ,
		\u2_ld_reg/P0001 ,
		\u7_dout_reg[7]/P0001 ,
		_w2333_
	);
	LUT3 #(
		.INIT('he2)
	) name187 (
		\u0_slt8_r_reg[5]/P0001 ,
		\u2_ld_reg/P0001 ,
		\u7_dout_reg[6]/P0001 ,
		_w2334_
	);
	LUT3 #(
		.INIT('he2)
	) name188 (
		\u0_slt8_r_reg[4]/P0001 ,
		\u2_ld_reg/P0001 ,
		\u7_dout_reg[5]/P0001 ,
		_w2335_
	);
	LUT3 #(
		.INIT('he2)
	) name189 (
		\u0_slt8_r_reg[3]/P0001 ,
		\u2_ld_reg/P0001 ,
		\u7_dout_reg[4]/P0001 ,
		_w2336_
	);
	LUT3 #(
		.INIT('he2)
	) name190 (
		\u0_slt8_r_reg[2]/P0001 ,
		\u2_ld_reg/P0001 ,
		\u7_dout_reg[3]/P0001 ,
		_w2337_
	);
	LUT3 #(
		.INIT('he2)
	) name191 (
		\u0_slt8_r_reg[1]/P0001 ,
		\u2_ld_reg/P0001 ,
		\u7_dout_reg[2]/P0001 ,
		_w2338_
	);
	LUT3 #(
		.INIT('he2)
	) name192 (
		\u0_slt8_r_reg[0]/P0001 ,
		\u2_ld_reg/P0001 ,
		\u7_dout_reg[1]/P0001 ,
		_w2339_
	);
	LUT3 #(
		.INIT('he2)
	) name193 (
		\u0_slt9_r_reg[19]/P0001 ,
		\u2_ld_reg/P0001 ,
		\u7_dout_reg[0]/P0001 ,
		_w2340_
	);
	LUT3 #(
		.INIT('he2)
	) name194 (
		\u0_slt9_r_reg[18]/P0001 ,
		\u2_ld_reg/P0001 ,
		\u8_dout_reg[19]/P0001 ,
		_w2341_
	);
	LUT3 #(
		.INIT('he2)
	) name195 (
		\u0_slt9_r_reg[17]/P0001 ,
		\u2_ld_reg/P0001 ,
		\u8_dout_reg[18]/P0001 ,
		_w2342_
	);
	LUT3 #(
		.INIT('he2)
	) name196 (
		\u0_slt9_r_reg[16]/P0001 ,
		\u2_ld_reg/P0001 ,
		\u8_dout_reg[17]/P0001 ,
		_w2343_
	);
	LUT3 #(
		.INIT('he2)
	) name197 (
		\u0_slt9_r_reg[15]/P0001 ,
		\u2_ld_reg/P0001 ,
		\u8_dout_reg[16]/P0001 ,
		_w2344_
	);
	LUT3 #(
		.INIT('he2)
	) name198 (
		\u0_slt9_r_reg[14]/P0001 ,
		\u2_ld_reg/P0001 ,
		\u8_dout_reg[15]/P0001 ,
		_w2345_
	);
	LUT3 #(
		.INIT('he2)
	) name199 (
		\u0_slt9_r_reg[13]/P0001 ,
		\u2_ld_reg/P0001 ,
		\u8_dout_reg[14]/P0001 ,
		_w2346_
	);
	LUT3 #(
		.INIT('he2)
	) name200 (
		\u0_slt9_r_reg[12]/P0001 ,
		\u2_ld_reg/P0001 ,
		\u8_dout_reg[13]/P0001 ,
		_w2347_
	);
	LUT3 #(
		.INIT('he2)
	) name201 (
		\u0_slt9_r_reg[11]/P0001 ,
		\u2_ld_reg/P0001 ,
		\u8_dout_reg[12]/P0001 ,
		_w2348_
	);
	LUT3 #(
		.INIT('he2)
	) name202 (
		\u0_slt9_r_reg[10]/P0001 ,
		\u2_ld_reg/P0001 ,
		\u8_dout_reg[11]/P0001 ,
		_w2349_
	);
	LUT3 #(
		.INIT('he2)
	) name203 (
		\u0_slt9_r_reg[9]/P0001 ,
		\u2_ld_reg/P0001 ,
		\u8_dout_reg[10]/P0001 ,
		_w2350_
	);
	LUT3 #(
		.INIT('he2)
	) name204 (
		\u0_slt9_r_reg[8]/P0001 ,
		\u2_ld_reg/P0001 ,
		\u8_dout_reg[9]/P0001 ,
		_w2351_
	);
	LUT3 #(
		.INIT('he2)
	) name205 (
		\u0_slt9_r_reg[7]/P0001 ,
		\u2_ld_reg/P0001 ,
		\u8_dout_reg[8]/P0001 ,
		_w2352_
	);
	LUT3 #(
		.INIT('he2)
	) name206 (
		\u0_slt9_r_reg[6]/P0001 ,
		\u2_ld_reg/P0001 ,
		\u8_dout_reg[7]/P0001 ,
		_w2353_
	);
	LUT3 #(
		.INIT('he2)
	) name207 (
		\u0_slt9_r_reg[5]/P0001 ,
		\u2_ld_reg/P0001 ,
		\u8_dout_reg[6]/P0001 ,
		_w2354_
	);
	LUT2 #(
		.INIT('h4)
	) name208 (
		\dma_ack_i[0]_pad ,
		\dma_req_o[0]_pad ,
		_w2355_
	);
	LUT4 #(
		.INIT('h0105)
	) name209 (
		\u13_occ0_r_reg[4]/NET0131 ,
		\u13_occ0_r_reg[5]/NET0131 ,
		\u3_status_reg[0]/P0001 ,
		\u3_status_reg[1]/P0001 ,
		_w2356_
	);
	LUT3 #(
		.INIT('h32)
	) name210 (
		\u13_occ0_r_reg[5]/NET0131 ,
		\u3_empty_reg/NET0131 ,
		\u3_status_reg[1]/P0001 ,
		_w2357_
	);
	LUT3 #(
		.INIT('h8a)
	) name211 (
		\u13_occ0_r_reg[0]/NET0131 ,
		_w2356_,
		_w2357_,
		_w2358_
	);
	LUT2 #(
		.INIT('h4)
	) name212 (
		\dma_ack_i[0]_pad ,
		\u13_occ0_r_reg[6]/NET0131 ,
		_w2359_
	);
	LUT4 #(
		.INIT('h8a00)
	) name213 (
		\u13_occ0_r_reg[0]/NET0131 ,
		_w2356_,
		_w2357_,
		_w2359_,
		_w2360_
	);
	LUT3 #(
		.INIT('hec)
	) name214 (
		\u16_u0_dma_req_r1_reg/P0001 ,
		_w2355_,
		_w2360_,
		_w2361_
	);
	LUT2 #(
		.INIT('h4)
	) name215 (
		\dma_ack_i[1]_pad ,
		\dma_req_o[1]_pad ,
		_w2362_
	);
	LUT4 #(
		.INIT('h0105)
	) name216 (
		\u13_occ0_r_reg[12]/NET0131 ,
		\u13_occ0_r_reg[13]/NET0131 ,
		\u4_status_reg[0]/P0001 ,
		\u4_status_reg[1]/P0001 ,
		_w2363_
	);
	LUT3 #(
		.INIT('h32)
	) name217 (
		\u13_occ0_r_reg[13]/NET0131 ,
		\u4_empty_reg/NET0131 ,
		\u4_status_reg[1]/P0001 ,
		_w2364_
	);
	LUT3 #(
		.INIT('h8a)
	) name218 (
		\u13_occ0_r_reg[8]/NET0131 ,
		_w2363_,
		_w2364_,
		_w2365_
	);
	LUT2 #(
		.INIT('h4)
	) name219 (
		\dma_ack_i[1]_pad ,
		\u13_occ0_r_reg[14]/NET0131 ,
		_w2366_
	);
	LUT4 #(
		.INIT('h8a00)
	) name220 (
		\u13_occ0_r_reg[8]/NET0131 ,
		_w2363_,
		_w2364_,
		_w2366_,
		_w2367_
	);
	LUT3 #(
		.INIT('hec)
	) name221 (
		\u16_u1_dma_req_r1_reg/P0001 ,
		_w2362_,
		_w2367_,
		_w2368_
	);
	LUT2 #(
		.INIT('h4)
	) name222 (
		\dma_ack_i[2]_pad ,
		\dma_req_o[2]_pad ,
		_w2369_
	);
	LUT4 #(
		.INIT('h0105)
	) name223 (
		\u13_occ0_r_reg[20]/NET0131 ,
		\u13_occ0_r_reg[21]/NET0131 ,
		\u5_status_reg[0]/P0001 ,
		\u5_status_reg[1]/P0001 ,
		_w2370_
	);
	LUT3 #(
		.INIT('h32)
	) name224 (
		\u13_occ0_r_reg[21]/NET0131 ,
		\u5_empty_reg/NET0131 ,
		\u5_status_reg[1]/P0001 ,
		_w2371_
	);
	LUT3 #(
		.INIT('h8a)
	) name225 (
		\u13_occ0_r_reg[16]/NET0131 ,
		_w2370_,
		_w2371_,
		_w2372_
	);
	LUT2 #(
		.INIT('h4)
	) name226 (
		\dma_ack_i[2]_pad ,
		\u13_occ0_r_reg[22]/NET0131 ,
		_w2373_
	);
	LUT4 #(
		.INIT('h8a00)
	) name227 (
		\u13_occ0_r_reg[16]/NET0131 ,
		_w2370_,
		_w2371_,
		_w2373_,
		_w2374_
	);
	LUT3 #(
		.INIT('hec)
	) name228 (
		\u16_u2_dma_req_r1_reg/P0001 ,
		_w2369_,
		_w2374_,
		_w2375_
	);
	LUT2 #(
		.INIT('h4)
	) name229 (
		\dma_ack_i[3]_pad ,
		\dma_req_o[3]_pad ,
		_w2376_
	);
	LUT4 #(
		.INIT('h0105)
	) name230 (
		\u13_occ0_r_reg[28]/NET0131 ,
		\u13_occ0_r_reg[29]/NET0131 ,
		\u6_status_reg[0]/P0001 ,
		\u6_status_reg[1]/P0001 ,
		_w2377_
	);
	LUT3 #(
		.INIT('h32)
	) name231 (
		\u13_occ0_r_reg[29]/NET0131 ,
		\u6_empty_reg/NET0131 ,
		\u6_status_reg[1]/P0001 ,
		_w2378_
	);
	LUT3 #(
		.INIT('h8a)
	) name232 (
		\u13_occ0_r_reg[24]/NET0131 ,
		_w2377_,
		_w2378_,
		_w2379_
	);
	LUT2 #(
		.INIT('h4)
	) name233 (
		\dma_ack_i[3]_pad ,
		\u13_occ0_r_reg[30]/NET0131 ,
		_w2380_
	);
	LUT4 #(
		.INIT('h8a00)
	) name234 (
		\u13_occ0_r_reg[24]/NET0131 ,
		_w2377_,
		_w2378_,
		_w2380_,
		_w2381_
	);
	LUT3 #(
		.INIT('hec)
	) name235 (
		\u16_u3_dma_req_r1_reg/P0001 ,
		_w2376_,
		_w2381_,
		_w2382_
	);
	LUT2 #(
		.INIT('h4)
	) name236 (
		\dma_ack_i[4]_pad ,
		\dma_req_o[4]_pad ,
		_w2383_
	);
	LUT4 #(
		.INIT('h0105)
	) name237 (
		\u13_occ1_r_reg[4]/NET0131 ,
		\u13_occ1_r_reg[5]/NET0131 ,
		\u7_status_reg[0]/P0001 ,
		\u7_status_reg[1]/P0001 ,
		_w2384_
	);
	LUT3 #(
		.INIT('h32)
	) name238 (
		\u13_occ1_r_reg[5]/NET0131 ,
		\u7_empty_reg/NET0131 ,
		\u7_status_reg[1]/P0001 ,
		_w2385_
	);
	LUT3 #(
		.INIT('h8a)
	) name239 (
		\u13_occ1_r_reg[0]/NET0131 ,
		_w2384_,
		_w2385_,
		_w2386_
	);
	LUT2 #(
		.INIT('h4)
	) name240 (
		\dma_ack_i[4]_pad ,
		\u13_occ1_r_reg[6]/NET0131 ,
		_w2387_
	);
	LUT4 #(
		.INIT('h8a00)
	) name241 (
		\u13_occ1_r_reg[0]/NET0131 ,
		_w2384_,
		_w2385_,
		_w2387_,
		_w2388_
	);
	LUT3 #(
		.INIT('hec)
	) name242 (
		\u16_u4_dma_req_r1_reg/P0001 ,
		_w2383_,
		_w2388_,
		_w2389_
	);
	LUT2 #(
		.INIT('h4)
	) name243 (
		\dma_ack_i[5]_pad ,
		\dma_req_o[5]_pad ,
		_w2390_
	);
	LUT4 #(
		.INIT('h0105)
	) name244 (
		\u13_occ1_r_reg[12]/NET0131 ,
		\u13_occ1_r_reg[13]/NET0131 ,
		\u8_status_reg[0]/P0001 ,
		\u8_status_reg[1]/P0001 ,
		_w2391_
	);
	LUT3 #(
		.INIT('h32)
	) name245 (
		\u13_occ1_r_reg[13]/NET0131 ,
		\u8_empty_reg/NET0131 ,
		\u8_status_reg[1]/P0001 ,
		_w2392_
	);
	LUT3 #(
		.INIT('h8a)
	) name246 (
		\u13_occ1_r_reg[8]/NET0131 ,
		_w2391_,
		_w2392_,
		_w2393_
	);
	LUT2 #(
		.INIT('h4)
	) name247 (
		\dma_ack_i[5]_pad ,
		\u13_occ1_r_reg[14]/NET0131 ,
		_w2394_
	);
	LUT4 #(
		.INIT('h8a00)
	) name248 (
		\u13_occ1_r_reg[8]/NET0131 ,
		_w2391_,
		_w2392_,
		_w2394_,
		_w2395_
	);
	LUT3 #(
		.INIT('hec)
	) name249 (
		\u16_u5_dma_req_r1_reg/P0001 ,
		_w2390_,
		_w2395_,
		_w2396_
	);
	LUT3 #(
		.INIT('he2)
	) name250 (
		\u0_slt9_r_reg[4]/P0001 ,
		\u2_ld_reg/P0001 ,
		\u8_dout_reg[5]/P0001 ,
		_w2397_
	);
	LUT2 #(
		.INIT('h1)
	) name251 (
		\u13_ints_r_reg[11]/NET0131 ,
		\u20_int_set_reg[0]/NET0131 ,
		_w2398_
	);
	LUT4 #(
		.INIT('h0040)
	) name252 (
		\u12_re2_reg/NET0131 ,
		wb_cyc_i_pad,
		wb_stb_i_pad,
		wb_we_i_pad,
		_w2399_
	);
	LUT2 #(
		.INIT('h8)
	) name253 (
		\u12_re1_reg/P0001 ,
		_w2399_,
		_w2400_
	);
	LUT2 #(
		.INIT('h1)
	) name254 (
		\wb_addr_i[5]_pad ,
		\wb_addr_i[6]_pad ,
		_w2401_
	);
	LUT3 #(
		.INIT('h40)
	) name255 (
		\wb_addr_i[2]_pad ,
		\wb_addr_i[3]_pad ,
		\wb_addr_i[4]_pad ,
		_w2402_
	);
	LUT4 #(
		.INIT('h8000)
	) name256 (
		\u12_re1_reg/P0001 ,
		_w2399_,
		_w2401_,
		_w2402_,
		_w2403_
	);
	LUT2 #(
		.INIT('h1)
	) name257 (
		_w2398_,
		_w2403_,
		_w2404_
	);
	LUT2 #(
		.INIT('h1)
	) name258 (
		\u13_ints_r_reg[14]/NET0131 ,
		\u21_int_set_reg[0]/NET0131 ,
		_w2405_
	);
	LUT2 #(
		.INIT('h1)
	) name259 (
		_w2403_,
		_w2405_,
		_w2406_
	);
	LUT2 #(
		.INIT('h1)
	) name260 (
		\u13_ints_r_reg[17]/NET0131 ,
		\u22_int_set_reg[0]/NET0131 ,
		_w2407_
	);
	LUT2 #(
		.INIT('h1)
	) name261 (
		_w2403_,
		_w2407_,
		_w2408_
	);
	LUT2 #(
		.INIT('h1)
	) name262 (
		\u13_ints_r_reg[2]/NET0131 ,
		\u17_int_set_reg[0]/NET0131 ,
		_w2409_
	);
	LUT2 #(
		.INIT('h1)
	) name263 (
		_w2403_,
		_w2409_,
		_w2410_
	);
	LUT2 #(
		.INIT('h1)
	) name264 (
		\u13_ints_r_reg[5]/NET0131 ,
		\u18_int_set_reg[0]/NET0131 ,
		_w2411_
	);
	LUT2 #(
		.INIT('h1)
	) name265 (
		_w2403_,
		_w2411_,
		_w2412_
	);
	LUT2 #(
		.INIT('h1)
	) name266 (
		\u13_ints_r_reg[8]/NET0131 ,
		\u19_int_set_reg[0]/NET0131 ,
		_w2413_
	);
	LUT2 #(
		.INIT('h1)
	) name267 (
		_w2403_,
		_w2413_,
		_w2414_
	);
	LUT3 #(
		.INIT('he2)
	) name268 (
		\u0_slt9_r_reg[3]/P0001 ,
		\u2_ld_reg/P0001 ,
		\u8_dout_reg[4]/P0001 ,
		_w2415_
	);
	LUT2 #(
		.INIT('h8)
	) name269 (
		\u14_u1_en_out_l_reg/NET0131 ,
		\valid_s_reg/NET0131 ,
		_w2416_
	);
	LUT3 #(
		.INIT('h40)
	) name270 (
		\u14_u1_en_out_l2_reg/P0001 ,
		\u14_u1_en_out_l_reg/NET0131 ,
		\valid_s_reg/NET0131 ,
		_w2417_
	);
	LUT2 #(
		.INIT('h1)
	) name271 (
		\u13_occ0_r_reg[10]/NET0131 ,
		\u13_occ0_r_reg[11]/NET0131 ,
		_w2418_
	);
	LUT3 #(
		.INIT('h01)
	) name272 (
		\u13_occ0_r_reg[10]/NET0131 ,
		\u13_occ0_r_reg[11]/NET0131 ,
		\u4_rp_reg[0]/P0001 ,
		_w2419_
	);
	LUT4 #(
		.INIT('h3313)
	) name273 (
		\u4_rp_reg[1]/NET0131 ,
		\u4_rp_reg[2]/NET0131 ,
		_w2417_,
		_w2419_,
		_w2420_
	);
	LUT2 #(
		.INIT('h8)
	) name274 (
		\u4_rp_reg[1]/NET0131 ,
		\u4_rp_reg[2]/NET0131 ,
		_w2421_
	);
	LUT3 #(
		.INIT('h20)
	) name275 (
		_w2417_,
		_w2419_,
		_w2421_,
		_w2422_
	);
	LUT4 #(
		.INIT('ha2aa)
	) name276 (
		\u13_occ0_r_reg[8]/NET0131 ,
		_w2417_,
		_w2419_,
		_w2421_,
		_w2423_
	);
	LUT2 #(
		.INIT('h4)
	) name277 (
		_w2420_,
		_w2423_,
		_w2424_
	);
	LUT2 #(
		.INIT('h8)
	) name278 (
		\u14_u2_en_out_l_reg/NET0131 ,
		\valid_s_reg/NET0131 ,
		_w2425_
	);
	LUT3 #(
		.INIT('h40)
	) name279 (
		\u14_u2_en_out_l2_reg/P0001 ,
		\u14_u2_en_out_l_reg/NET0131 ,
		\valid_s_reg/NET0131 ,
		_w2426_
	);
	LUT2 #(
		.INIT('h1)
	) name280 (
		\u13_occ0_r_reg[18]/NET0131 ,
		\u13_occ0_r_reg[19]/NET0131 ,
		_w2427_
	);
	LUT3 #(
		.INIT('h01)
	) name281 (
		\u13_occ0_r_reg[18]/NET0131 ,
		\u13_occ0_r_reg[19]/NET0131 ,
		\u5_rp_reg[0]/P0001 ,
		_w2428_
	);
	LUT4 #(
		.INIT('h3313)
	) name282 (
		\u5_rp_reg[1]/NET0131 ,
		\u5_rp_reg[2]/NET0131 ,
		_w2426_,
		_w2428_,
		_w2429_
	);
	LUT2 #(
		.INIT('h8)
	) name283 (
		\u5_rp_reg[1]/NET0131 ,
		\u5_rp_reg[2]/NET0131 ,
		_w2430_
	);
	LUT3 #(
		.INIT('h20)
	) name284 (
		_w2426_,
		_w2428_,
		_w2430_,
		_w2431_
	);
	LUT4 #(
		.INIT('ha2aa)
	) name285 (
		\u13_occ0_r_reg[16]/NET0131 ,
		_w2426_,
		_w2428_,
		_w2430_,
		_w2432_
	);
	LUT2 #(
		.INIT('h4)
	) name286 (
		_w2429_,
		_w2432_,
		_w2433_
	);
	LUT4 #(
		.INIT('h3313)
	) name287 (
		\u8_rp_reg[1]/NET0131 ,
		\u8_rp_reg[2]/NET0131 ,
		_w2155_,
		_w2157_,
		_w2434_
	);
	LUT4 #(
		.INIT('ha2aa)
	) name288 (
		\u13_occ1_r_reg[8]/NET0131 ,
		_w2155_,
		_w2157_,
		_w2158_,
		_w2435_
	);
	LUT2 #(
		.INIT('h4)
	) name289 (
		_w2434_,
		_w2435_,
		_w2436_
	);
	LUT2 #(
		.INIT('h1)
	) name290 (
		\u13_occ0_r_reg[2]/NET0131 ,
		\u13_occ0_r_reg[3]/NET0131 ,
		_w2437_
	);
	LUT3 #(
		.INIT('h01)
	) name291 (
		\u13_occ0_r_reg[2]/NET0131 ,
		\u13_occ0_r_reg[3]/NET0131 ,
		\u3_rp_reg[0]/P0001 ,
		_w2438_
	);
	LUT3 #(
		.INIT('h40)
	) name292 (
		\u14_u0_en_out_l2_reg/P0001 ,
		\u14_u0_en_out_l_reg/NET0131 ,
		\valid_s_reg/NET0131 ,
		_w2439_
	);
	LUT3 #(
		.INIT('h20)
	) name293 (
		\u3_rp_reg[1]/NET0131 ,
		_w2438_,
		_w2439_,
		_w2440_
	);
	LUT4 #(
		.INIT('h0800)
	) name294 (
		\u3_rp_reg[1]/NET0131 ,
		\u3_rp_reg[2]/NET0131 ,
		_w2438_,
		_w2439_,
		_w2441_
	);
	LUT3 #(
		.INIT('h28)
	) name295 (
		\u13_occ0_r_reg[0]/NET0131 ,
		\u3_rp_reg[2]/NET0131 ,
		_w2440_,
		_w2442_
	);
	LUT2 #(
		.INIT('h8)
	) name296 (
		\u14_u3_en_out_l_reg/NET0131 ,
		\valid_s_reg/NET0131 ,
		_w2443_
	);
	LUT3 #(
		.INIT('h40)
	) name297 (
		\u14_u3_en_out_l2_reg/P0001 ,
		\u14_u3_en_out_l_reg/NET0131 ,
		\valid_s_reg/NET0131 ,
		_w2444_
	);
	LUT2 #(
		.INIT('h1)
	) name298 (
		\u13_occ0_r_reg[26]/NET0131 ,
		\u13_occ0_r_reg[27]/NET0131 ,
		_w2445_
	);
	LUT3 #(
		.INIT('h01)
	) name299 (
		\u13_occ0_r_reg[26]/NET0131 ,
		\u13_occ0_r_reg[27]/NET0131 ,
		\u6_rp_reg[0]/P0001 ,
		_w2446_
	);
	LUT4 #(
		.INIT('h3313)
	) name300 (
		\u6_rp_reg[1]/NET0131 ,
		\u6_rp_reg[2]/NET0131 ,
		_w2444_,
		_w2446_,
		_w2447_
	);
	LUT2 #(
		.INIT('h8)
	) name301 (
		\u6_rp_reg[1]/NET0131 ,
		\u6_rp_reg[2]/NET0131 ,
		_w2448_
	);
	LUT3 #(
		.INIT('h20)
	) name302 (
		_w2444_,
		_w2446_,
		_w2448_,
		_w2449_
	);
	LUT4 #(
		.INIT('ha2aa)
	) name303 (
		\u13_occ0_r_reg[24]/NET0131 ,
		_w2444_,
		_w2446_,
		_w2448_,
		_w2450_
	);
	LUT2 #(
		.INIT('h4)
	) name304 (
		_w2447_,
		_w2450_,
		_w2451_
	);
	LUT2 #(
		.INIT('h1)
	) name305 (
		\u13_occ1_r_reg[2]/NET0131 ,
		\u13_occ1_r_reg[3]/NET0131 ,
		_w2452_
	);
	LUT3 #(
		.INIT('h01)
	) name306 (
		\u13_occ1_r_reg[2]/NET0131 ,
		\u13_occ1_r_reg[3]/NET0131 ,
		\u7_rp_reg[0]/P0001 ,
		_w2453_
	);
	LUT2 #(
		.INIT('h8)
	) name307 (
		\u14_u4_en_out_l_reg/NET0131 ,
		\valid_s_reg/NET0131 ,
		_w2454_
	);
	LUT3 #(
		.INIT('h40)
	) name308 (
		\u14_u4_en_out_l2_reg/P0001 ,
		\u14_u4_en_out_l_reg/NET0131 ,
		\valid_s_reg/NET0131 ,
		_w2455_
	);
	LUT3 #(
		.INIT('h20)
	) name309 (
		\u7_rp_reg[1]/NET0131 ,
		_w2453_,
		_w2455_,
		_w2456_
	);
	LUT4 #(
		.INIT('h0800)
	) name310 (
		\u7_rp_reg[1]/NET0131 ,
		\u7_rp_reg[2]/NET0131 ,
		_w2453_,
		_w2455_,
		_w2457_
	);
	LUT3 #(
		.INIT('h28)
	) name311 (
		\u13_occ1_r_reg[0]/NET0131 ,
		\u7_rp_reg[2]/NET0131 ,
		_w2456_,
		_w2458_
	);
	LUT3 #(
		.INIT('h28)
	) name312 (
		\u13_occ0_r_reg[0]/NET0131 ,
		\u3_rp_reg[3]/NET0131 ,
		_w2441_,
		_w2459_
	);
	LUT3 #(
		.INIT('h28)
	) name313 (
		\u13_occ0_r_reg[8]/NET0131 ,
		\u4_rp_reg[3]/NET0131 ,
		_w2422_,
		_w2460_
	);
	LUT2 #(
		.INIT('h1)
	) name314 (
		\u13_ints_r_reg[20]/NET0131 ,
		\u23_int_set_reg[0]/NET0131 ,
		_w2461_
	);
	LUT2 #(
		.INIT('h1)
	) name315 (
		_w2403_,
		_w2461_,
		_w2462_
	);
	LUT2 #(
		.INIT('h1)
	) name316 (
		\u13_ints_r_reg[23]/NET0131 ,
		\u24_int_set_reg[0]/NET0131 ,
		_w2463_
	);
	LUT2 #(
		.INIT('h1)
	) name317 (
		_w2403_,
		_w2463_,
		_w2464_
	);
	LUT2 #(
		.INIT('h1)
	) name318 (
		\u13_ints_r_reg[26]/NET0131 ,
		\u25_int_set_reg[0]/NET0131 ,
		_w2465_
	);
	LUT2 #(
		.INIT('h1)
	) name319 (
		_w2403_,
		_w2465_,
		_w2466_
	);
	LUT3 #(
		.INIT('h28)
	) name320 (
		\u13_occ0_r_reg[16]/NET0131 ,
		\u5_rp_reg[3]/NET0131 ,
		_w2431_,
		_w2467_
	);
	LUT3 #(
		.INIT('h28)
	) name321 (
		\u13_occ0_r_reg[24]/NET0131 ,
		\u6_rp_reg[3]/NET0131 ,
		_w2449_,
		_w2468_
	);
	LUT3 #(
		.INIT('h28)
	) name322 (
		\u13_occ1_r_reg[0]/NET0131 ,
		\u7_rp_reg[3]/NET0131 ,
		_w2457_,
		_w2469_
	);
	LUT4 #(
		.INIT('h8828)
	) name323 (
		\u13_occ1_r_reg[8]/NET0131 ,
		\u8_rp_reg[1]/NET0131 ,
		_w2155_,
		_w2157_,
		_w2470_
	);
	LUT4 #(
		.INIT('h8288)
	) name324 (
		\u13_occ0_r_reg[0]/NET0131 ,
		\u3_rp_reg[1]/NET0131 ,
		_w2438_,
		_w2439_,
		_w2471_
	);
	LUT4 #(
		.INIT('h8828)
	) name325 (
		\u13_occ0_r_reg[8]/NET0131 ,
		\u4_rp_reg[1]/NET0131 ,
		_w2417_,
		_w2419_,
		_w2472_
	);
	LUT4 #(
		.INIT('h8828)
	) name326 (
		\u13_occ0_r_reg[16]/NET0131 ,
		\u5_rp_reg[1]/NET0131 ,
		_w2426_,
		_w2428_,
		_w2473_
	);
	LUT4 #(
		.INIT('h8828)
	) name327 (
		\u13_occ0_r_reg[24]/NET0131 ,
		\u6_rp_reg[1]/NET0131 ,
		_w2444_,
		_w2446_,
		_w2474_
	);
	LUT4 #(
		.INIT('h8288)
	) name328 (
		\u13_occ1_r_reg[0]/NET0131 ,
		\u7_rp_reg[1]/NET0131 ,
		_w2453_,
		_w2455_,
		_w2475_
	);
	LUT3 #(
		.INIT('he2)
	) name329 (
		\u0_slt9_r_reg[2]/P0001 ,
		\u2_ld_reg/P0001 ,
		\u8_dout_reg[3]/P0001 ,
		_w2476_
	);
	LUT3 #(
		.INIT('h07)
	) name330 (
		suspended_o_pad,
		\u13_resume_req_reg/P0001 ,
		\u2_sync_resume_reg/NET0131 ,
		_w2477_
	);
	LUT4 #(
		.INIT('h0020)
	) name331 (
		\u2_res_cnt_reg[0]/P0001 ,
		\u2_res_cnt_reg[1]/P0001 ,
		\u2_res_cnt_reg[2]/P0001 ,
		\u2_res_cnt_reg[3]/P0001 ,
		_w2478_
	);
	LUT2 #(
		.INIT('h1)
	) name332 (
		_w2477_,
		_w2478_,
		_w2479_
	);
	LUT4 #(
		.INIT('h2888)
	) name333 (
		\u13_occ1_r_reg[8]/NET0131 ,
		\u8_rp_reg[0]/P0001 ,
		_w2155_,
		_w2156_,
		_w2480_
	);
	LUT4 #(
		.INIT('h2888)
	) name334 (
		\u13_occ0_r_reg[0]/NET0131 ,
		\u3_rp_reg[0]/P0001 ,
		_w2437_,
		_w2439_,
		_w2481_
	);
	LUT4 #(
		.INIT('h2888)
	) name335 (
		\u13_occ0_r_reg[8]/NET0131 ,
		\u4_rp_reg[0]/P0001 ,
		_w2417_,
		_w2418_,
		_w2482_
	);
	LUT4 #(
		.INIT('h2888)
	) name336 (
		\u13_occ0_r_reg[16]/NET0131 ,
		\u5_rp_reg[0]/P0001 ,
		_w2426_,
		_w2427_,
		_w2483_
	);
	LUT4 #(
		.INIT('h2888)
	) name337 (
		\u13_occ0_r_reg[24]/NET0131 ,
		\u6_rp_reg[0]/P0001 ,
		_w2444_,
		_w2445_,
		_w2484_
	);
	LUT4 #(
		.INIT('h2888)
	) name338 (
		\u13_occ1_r_reg[0]/NET0131 ,
		\u7_rp_reg[0]/P0001 ,
		_w2452_,
		_w2455_,
		_w2485_
	);
	LUT4 #(
		.INIT('h8aaa)
	) name339 (
		\u13_occ0_r_reg[8]/NET0131 ,
		\u14_u1_en_out_l2_reg/P0001 ,
		\u14_u1_en_out_l_reg/NET0131 ,
		\valid_s_reg/NET0131 ,
		_w2486_
	);
	LUT2 #(
		.INIT('h8)
	) name340 (
		\u4_dout_reg[0]/P0001 ,
		_w2486_,
		_w2487_
	);
	LUT4 #(
		.INIT('h35ff)
	) name341 (
		\u4_mem_reg[2][0]/NET0131 ,
		\u4_mem_reg[3][0]/NET0131 ,
		\u4_rp_reg[1]/NET0131 ,
		\u4_rp_reg[2]/NET0131 ,
		_w2488_
	);
	LUT4 #(
		.INIT('hff35)
	) name342 (
		\u4_mem_reg[0][0]/NET0131 ,
		\u4_mem_reg[1][0]/NET0131 ,
		\u4_rp_reg[1]/NET0131 ,
		\u4_rp_reg[2]/NET0131 ,
		_w2489_
	);
	LUT2 #(
		.INIT('h4)
	) name343 (
		\u13_occ0_r_reg[10]/NET0131 ,
		\u13_occ0_r_reg[11]/NET0131 ,
		_w2490_
	);
	LUT3 #(
		.INIT('h40)
	) name344 (
		\u13_occ0_r_reg[10]/NET0131 ,
		\u13_occ0_r_reg[11]/NET0131 ,
		\u13_occ0_r_reg[8]/NET0131 ,
		_w2491_
	);
	LUT4 #(
		.INIT('h2a00)
	) name345 (
		_w2417_,
		_w2488_,
		_w2489_,
		_w2491_,
		_w2492_
	);
	LUT2 #(
		.INIT('he)
	) name346 (
		_w2487_,
		_w2492_,
		_w2493_
	);
	LUT2 #(
		.INIT('h8)
	) name347 (
		\u4_dout_reg[1]/P0001 ,
		_w2486_,
		_w2494_
	);
	LUT4 #(
		.INIT('h35ff)
	) name348 (
		\u4_mem_reg[2][1]/NET0131 ,
		\u4_mem_reg[3][1]/NET0131 ,
		\u4_rp_reg[1]/NET0131 ,
		\u4_rp_reg[2]/NET0131 ,
		_w2495_
	);
	LUT4 #(
		.INIT('hff35)
	) name349 (
		\u4_mem_reg[0][1]/NET0131 ,
		\u4_mem_reg[1][1]/NET0131 ,
		\u4_rp_reg[1]/NET0131 ,
		\u4_rp_reg[2]/NET0131 ,
		_w2496_
	);
	LUT4 #(
		.INIT('h0888)
	) name350 (
		_w2417_,
		_w2491_,
		_w2495_,
		_w2496_,
		_w2497_
	);
	LUT2 #(
		.INIT('he)
	) name351 (
		_w2494_,
		_w2497_,
		_w2498_
	);
	LUT4 #(
		.INIT('h8aaa)
	) name352 (
		\u13_occ0_r_reg[16]/NET0131 ,
		\u14_u2_en_out_l2_reg/P0001 ,
		\u14_u2_en_out_l_reg/NET0131 ,
		\valid_s_reg/NET0131 ,
		_w2499_
	);
	LUT2 #(
		.INIT('h8)
	) name353 (
		\u5_dout_reg[0]/P0001 ,
		_w2499_,
		_w2500_
	);
	LUT4 #(
		.INIT('h3f5f)
	) name354 (
		\u5_mem_reg[1][0]/NET0131 ,
		\u5_mem_reg[3][0]/NET0131 ,
		\u5_rp_reg[1]/NET0131 ,
		\u5_rp_reg[2]/NET0131 ,
		_w2501_
	);
	LUT4 #(
		.INIT('hf3f5)
	) name355 (
		\u5_mem_reg[0][0]/NET0131 ,
		\u5_mem_reg[2][0]/NET0131 ,
		\u5_rp_reg[1]/NET0131 ,
		\u5_rp_reg[2]/NET0131 ,
		_w2502_
	);
	LUT2 #(
		.INIT('h4)
	) name356 (
		\u13_occ0_r_reg[18]/NET0131 ,
		\u13_occ0_r_reg[19]/NET0131 ,
		_w2503_
	);
	LUT3 #(
		.INIT('h20)
	) name357 (
		\u13_occ0_r_reg[16]/NET0131 ,
		\u13_occ0_r_reg[18]/NET0131 ,
		\u13_occ0_r_reg[19]/NET0131 ,
		_w2504_
	);
	LUT4 #(
		.INIT('h2a00)
	) name358 (
		_w2426_,
		_w2501_,
		_w2502_,
		_w2504_,
		_w2505_
	);
	LUT2 #(
		.INIT('he)
	) name359 (
		_w2500_,
		_w2505_,
		_w2506_
	);
	LUT2 #(
		.INIT('h8)
	) name360 (
		\u5_dout_reg[1]/P0001 ,
		_w2499_,
		_w2507_
	);
	LUT4 #(
		.INIT('h3f5f)
	) name361 (
		\u5_mem_reg[1][1]/NET0131 ,
		\u5_mem_reg[3][1]/NET0131 ,
		\u5_rp_reg[1]/NET0131 ,
		\u5_rp_reg[2]/NET0131 ,
		_w2508_
	);
	LUT4 #(
		.INIT('hf3f5)
	) name362 (
		\u5_mem_reg[0][1]/NET0131 ,
		\u5_mem_reg[2][1]/NET0131 ,
		\u5_rp_reg[1]/NET0131 ,
		\u5_rp_reg[2]/NET0131 ,
		_w2509_
	);
	LUT4 #(
		.INIT('h0888)
	) name363 (
		_w2426_,
		_w2504_,
		_w2508_,
		_w2509_,
		_w2510_
	);
	LUT2 #(
		.INIT('he)
	) name364 (
		_w2507_,
		_w2510_,
		_w2511_
	);
	LUT4 #(
		.INIT('h8aaa)
	) name365 (
		\u13_occ0_r_reg[24]/NET0131 ,
		\u14_u3_en_out_l2_reg/P0001 ,
		\u14_u3_en_out_l_reg/NET0131 ,
		\valid_s_reg/NET0131 ,
		_w2512_
	);
	LUT2 #(
		.INIT('h8)
	) name366 (
		\u6_dout_reg[0]/P0001 ,
		_w2512_,
		_w2513_
	);
	LUT4 #(
		.INIT('h35ff)
	) name367 (
		\u6_mem_reg[2][0]/NET0131 ,
		\u6_mem_reg[3][0]/NET0131 ,
		\u6_rp_reg[1]/NET0131 ,
		\u6_rp_reg[2]/NET0131 ,
		_w2514_
	);
	LUT4 #(
		.INIT('hff35)
	) name368 (
		\u6_mem_reg[0][0]/NET0131 ,
		\u6_mem_reg[1][0]/NET0131 ,
		\u6_rp_reg[1]/NET0131 ,
		\u6_rp_reg[2]/NET0131 ,
		_w2515_
	);
	LUT2 #(
		.INIT('h4)
	) name369 (
		\u13_occ0_r_reg[26]/NET0131 ,
		\u13_occ0_r_reg[27]/NET0131 ,
		_w2516_
	);
	LUT3 #(
		.INIT('h20)
	) name370 (
		\u13_occ0_r_reg[24]/NET0131 ,
		\u13_occ0_r_reg[26]/NET0131 ,
		\u13_occ0_r_reg[27]/NET0131 ,
		_w2517_
	);
	LUT4 #(
		.INIT('h2a00)
	) name371 (
		_w2444_,
		_w2514_,
		_w2515_,
		_w2517_,
		_w2518_
	);
	LUT2 #(
		.INIT('he)
	) name372 (
		_w2513_,
		_w2518_,
		_w2519_
	);
	LUT2 #(
		.INIT('h8)
	) name373 (
		\u6_dout_reg[1]/P0001 ,
		_w2512_,
		_w2520_
	);
	LUT4 #(
		.INIT('hf35f)
	) name374 (
		\u6_mem_reg[1][1]/NET0131 ,
		\u6_mem_reg[2][1]/NET0131 ,
		\u6_rp_reg[1]/NET0131 ,
		\u6_rp_reg[2]/NET0131 ,
		_w2521_
	);
	LUT4 #(
		.INIT('h3ff5)
	) name375 (
		\u6_mem_reg[0][1]/NET0131 ,
		\u6_mem_reg[3][1]/NET0131 ,
		\u6_rp_reg[1]/NET0131 ,
		\u6_rp_reg[2]/NET0131 ,
		_w2522_
	);
	LUT4 #(
		.INIT('h0888)
	) name376 (
		_w2444_,
		_w2517_,
		_w2521_,
		_w2522_,
		_w2523_
	);
	LUT2 #(
		.INIT('he)
	) name377 (
		_w2520_,
		_w2523_,
		_w2524_
	);
	LUT4 #(
		.INIT('h8aaa)
	) name378 (
		\u13_occ1_r_reg[0]/NET0131 ,
		\u14_u4_en_out_l2_reg/P0001 ,
		\u14_u4_en_out_l_reg/NET0131 ,
		\valid_s_reg/NET0131 ,
		_w2525_
	);
	LUT2 #(
		.INIT('h8)
	) name379 (
		\u7_dout_reg[0]/P0001 ,
		_w2525_,
		_w2526_
	);
	LUT4 #(
		.INIT('h35ff)
	) name380 (
		\u7_mem_reg[2][0]/NET0131 ,
		\u7_mem_reg[3][0]/NET0131 ,
		\u7_rp_reg[1]/NET0131 ,
		\u7_rp_reg[2]/NET0131 ,
		_w2527_
	);
	LUT4 #(
		.INIT('hff35)
	) name381 (
		\u7_mem_reg[0][0]/NET0131 ,
		\u7_mem_reg[1][0]/NET0131 ,
		\u7_rp_reg[1]/NET0131 ,
		\u7_rp_reg[2]/NET0131 ,
		_w2528_
	);
	LUT2 #(
		.INIT('h4)
	) name382 (
		\u13_occ1_r_reg[2]/NET0131 ,
		\u13_occ1_r_reg[3]/NET0131 ,
		_w2529_
	);
	LUT3 #(
		.INIT('h20)
	) name383 (
		\u13_occ1_r_reg[0]/NET0131 ,
		\u13_occ1_r_reg[2]/NET0131 ,
		\u13_occ1_r_reg[3]/NET0131 ,
		_w2530_
	);
	LUT4 #(
		.INIT('h2a00)
	) name384 (
		_w2455_,
		_w2527_,
		_w2528_,
		_w2530_,
		_w2531_
	);
	LUT2 #(
		.INIT('he)
	) name385 (
		_w2526_,
		_w2531_,
		_w2532_
	);
	LUT2 #(
		.INIT('h8)
	) name386 (
		\u7_dout_reg[1]/P0001 ,
		_w2525_,
		_w2533_
	);
	LUT4 #(
		.INIT('h35ff)
	) name387 (
		\u7_mem_reg[2][1]/NET0131 ,
		\u7_mem_reg[3][1]/NET0131 ,
		\u7_rp_reg[1]/NET0131 ,
		\u7_rp_reg[2]/NET0131 ,
		_w2534_
	);
	LUT4 #(
		.INIT('hff35)
	) name388 (
		\u7_mem_reg[0][1]/NET0131 ,
		\u7_mem_reg[1][1]/NET0131 ,
		\u7_rp_reg[1]/NET0131 ,
		\u7_rp_reg[2]/NET0131 ,
		_w2535_
	);
	LUT4 #(
		.INIT('h0888)
	) name389 (
		_w2455_,
		_w2530_,
		_w2534_,
		_w2535_,
		_w2536_
	);
	LUT2 #(
		.INIT('he)
	) name390 (
		_w2533_,
		_w2536_,
		_w2537_
	);
	LUT4 #(
		.INIT('h8aaa)
	) name391 (
		\u13_occ0_r_reg[0]/NET0131 ,
		\u14_u0_en_out_l2_reg/P0001 ,
		\u14_u0_en_out_l_reg/NET0131 ,
		\valid_s_reg/NET0131 ,
		_w2538_
	);
	LUT2 #(
		.INIT('h8)
	) name392 (
		\u3_dout_reg[0]/P0001 ,
		_w2538_,
		_w2539_
	);
	LUT4 #(
		.INIT('h35ff)
	) name393 (
		\u3_mem_reg[2][0]/NET0131 ,
		\u3_mem_reg[3][0]/NET0131 ,
		\u3_rp_reg[1]/NET0131 ,
		\u3_rp_reg[2]/NET0131 ,
		_w2540_
	);
	LUT4 #(
		.INIT('hff35)
	) name394 (
		\u3_mem_reg[0][0]/NET0131 ,
		\u3_mem_reg[1][0]/NET0131 ,
		\u3_rp_reg[1]/NET0131 ,
		\u3_rp_reg[2]/NET0131 ,
		_w2541_
	);
	LUT2 #(
		.INIT('h4)
	) name395 (
		\u13_occ0_r_reg[2]/NET0131 ,
		\u13_occ0_r_reg[3]/NET0131 ,
		_w2542_
	);
	LUT3 #(
		.INIT('h20)
	) name396 (
		\u13_occ0_r_reg[0]/NET0131 ,
		\u13_occ0_r_reg[2]/NET0131 ,
		\u13_occ0_r_reg[3]/NET0131 ,
		_w2543_
	);
	LUT4 #(
		.INIT('h2a00)
	) name397 (
		_w2439_,
		_w2540_,
		_w2541_,
		_w2543_,
		_w2544_
	);
	LUT2 #(
		.INIT('he)
	) name398 (
		_w2539_,
		_w2544_,
		_w2545_
	);
	LUT4 #(
		.INIT('h8aaa)
	) name399 (
		\u13_occ1_r_reg[8]/NET0131 ,
		\u14_u5_en_out_l2_reg/P0001 ,
		\u14_u5_en_out_l_reg/NET0131 ,
		\valid_s_reg/NET0131 ,
		_w2546_
	);
	LUT2 #(
		.INIT('h8)
	) name400 (
		\u8_dout_reg[0]/P0001 ,
		_w2546_,
		_w2547_
	);
	LUT4 #(
		.INIT('h35ff)
	) name401 (
		\u8_mem_reg[2][0]/NET0131 ,
		\u8_mem_reg[3][0]/NET0131 ,
		\u8_rp_reg[1]/NET0131 ,
		\u8_rp_reg[2]/NET0131 ,
		_w2548_
	);
	LUT4 #(
		.INIT('hff35)
	) name402 (
		\u8_mem_reg[0][0]/NET0131 ,
		\u8_mem_reg[1][0]/NET0131 ,
		\u8_rp_reg[1]/NET0131 ,
		\u8_rp_reg[2]/NET0131 ,
		_w2549_
	);
	LUT2 #(
		.INIT('h4)
	) name403 (
		\u13_occ1_r_reg[10]/NET0131 ,
		\u13_occ1_r_reg[11]/NET0131 ,
		_w2550_
	);
	LUT3 #(
		.INIT('h40)
	) name404 (
		\u13_occ1_r_reg[10]/NET0131 ,
		\u13_occ1_r_reg[11]/NET0131 ,
		\u13_occ1_r_reg[8]/NET0131 ,
		_w2551_
	);
	LUT4 #(
		.INIT('h2a00)
	) name405 (
		_w2155_,
		_w2548_,
		_w2549_,
		_w2551_,
		_w2552_
	);
	LUT2 #(
		.INIT('he)
	) name406 (
		_w2547_,
		_w2552_,
		_w2553_
	);
	LUT2 #(
		.INIT('h8)
	) name407 (
		\u3_dout_reg[1]/P0001 ,
		_w2538_,
		_w2554_
	);
	LUT4 #(
		.INIT('hf35f)
	) name408 (
		\u3_mem_reg[1][1]/NET0131 ,
		\u3_mem_reg[2][1]/NET0131 ,
		\u3_rp_reg[1]/NET0131 ,
		\u3_rp_reg[2]/NET0131 ,
		_w2555_
	);
	LUT4 #(
		.INIT('h3ff5)
	) name409 (
		\u3_mem_reg[0][1]/NET0131 ,
		\u3_mem_reg[3][1]/NET0131 ,
		\u3_rp_reg[1]/NET0131 ,
		\u3_rp_reg[2]/NET0131 ,
		_w2556_
	);
	LUT4 #(
		.INIT('h0888)
	) name410 (
		_w2439_,
		_w2543_,
		_w2555_,
		_w2556_,
		_w2557_
	);
	LUT2 #(
		.INIT('he)
	) name411 (
		_w2554_,
		_w2557_,
		_w2558_
	);
	LUT2 #(
		.INIT('h8)
	) name412 (
		\u8_dout_reg[1]/P0001 ,
		_w2546_,
		_w2559_
	);
	LUT4 #(
		.INIT('h35ff)
	) name413 (
		\u8_mem_reg[2][1]/NET0131 ,
		\u8_mem_reg[3][1]/NET0131 ,
		\u8_rp_reg[1]/NET0131 ,
		\u8_rp_reg[2]/NET0131 ,
		_w2560_
	);
	LUT4 #(
		.INIT('hff35)
	) name414 (
		\u8_mem_reg[0][1]/NET0131 ,
		\u8_mem_reg[1][1]/NET0131 ,
		\u8_rp_reg[1]/NET0131 ,
		\u8_rp_reg[2]/NET0131 ,
		_w2561_
	);
	LUT4 #(
		.INIT('h0888)
	) name415 (
		_w2155_,
		_w2551_,
		_w2560_,
		_w2561_,
		_w2562_
	);
	LUT2 #(
		.INIT('he)
	) name416 (
		_w2559_,
		_w2562_,
		_w2563_
	);
	LUT2 #(
		.INIT('h8)
	) name417 (
		\in_valid_s_reg[2]/NET0131 ,
		\u14_u8_en_out_l_reg/NET0131 ,
		_w2564_
	);
	LUT3 #(
		.INIT('h20)
	) name418 (
		\in_valid_s_reg[2]/NET0131 ,
		\u14_u8_en_out_l2_reg/P0001 ,
		\u14_u8_en_out_l_reg/NET0131 ,
		_w2565_
	);
	LUT2 #(
		.INIT('h1)
	) name419 (
		\u13_icc_r_reg[18]/NET0131 ,
		\u13_icc_r_reg[19]/NET0131 ,
		_w2566_
	);
	LUT3 #(
		.INIT('h01)
	) name420 (
		\u11_wp_reg[0]/NET0131 ,
		\u13_icc_r_reg[18]/NET0131 ,
		\u13_icc_r_reg[19]/NET0131 ,
		_w2567_
	);
	LUT2 #(
		.INIT('h2)
	) name421 (
		_w2565_,
		_w2567_,
		_w2568_
	);
	LUT3 #(
		.INIT('h08)
	) name422 (
		\u11_wp_reg[1]/P0001 ,
		_w2565_,
		_w2567_,
		_w2569_
	);
	LUT4 #(
		.INIT('h0080)
	) name423 (
		\u11_wp_reg[1]/P0001 ,
		\u11_wp_reg[2]/P0001 ,
		_w2565_,
		_w2567_,
		_w2570_
	);
	LUT3 #(
		.INIT('h48)
	) name424 (
		\u11_wp_reg[2]/P0001 ,
		\u13_icc_r_reg[16]/NET0131 ,
		_w2569_,
		_w2571_
	);
	LUT4 #(
		.INIT('hc4cc)
	) name425 (
		\u4_mem_reg[2][22]/NET0131 ,
		\u4_rp_reg[0]/P0001 ,
		\u4_rp_reg[1]/NET0131 ,
		\u4_rp_reg[2]/NET0131 ,
		_w2572_
	);
	LUT3 #(
		.INIT('h02)
	) name426 (
		\u4_mem_reg[0][22]/NET0131 ,
		\u4_rp_reg[1]/NET0131 ,
		\u4_rp_reg[2]/NET0131 ,
		_w2573_
	);
	LUT4 #(
		.INIT('h3f5f)
	) name427 (
		\u4_mem_reg[1][22]/NET0131 ,
		\u4_mem_reg[3][22]/NET0131 ,
		\u4_rp_reg[1]/NET0131 ,
		\u4_rp_reg[2]/NET0131 ,
		_w2574_
	);
	LUT3 #(
		.INIT('h40)
	) name428 (
		_w2573_,
		_w2572_,
		_w2574_,
		_w2575_
	);
	LUT4 #(
		.INIT('h35ff)
	) name429 (
		\u4_mem_reg[2][6]/NET0131 ,
		\u4_mem_reg[3][6]/NET0131 ,
		\u4_rp_reg[1]/NET0131 ,
		\u4_rp_reg[2]/NET0131 ,
		_w2576_
	);
	LUT4 #(
		.INIT('hff35)
	) name430 (
		\u4_mem_reg[0][6]/NET0131 ,
		\u4_mem_reg[1][6]/NET0131 ,
		\u4_rp_reg[1]/NET0131 ,
		\u4_rp_reg[2]/NET0131 ,
		_w2577_
	);
	LUT4 #(
		.INIT('h8ccc)
	) name431 (
		\u4_rp_reg[0]/P0001 ,
		_w2418_,
		_w2576_,
		_w2577_,
		_w2578_
	);
	LUT2 #(
		.INIT('h2)
	) name432 (
		\u13_occ0_r_reg[10]/NET0131 ,
		\u13_occ0_r_reg[11]/NET0131 ,
		_w2579_
	);
	LUT4 #(
		.INIT('h35ff)
	) name433 (
		\u4_mem_reg[2][8]/NET0131 ,
		\u4_mem_reg[3][8]/NET0131 ,
		\u4_rp_reg[1]/NET0131 ,
		\u4_rp_reg[2]/NET0131 ,
		_w2580_
	);
	LUT4 #(
		.INIT('hff35)
	) name434 (
		\u4_mem_reg[0][8]/NET0131 ,
		\u4_mem_reg[1][8]/NET0131 ,
		\u4_rp_reg[1]/NET0131 ,
		\u4_rp_reg[2]/NET0131 ,
		_w2581_
	);
	LUT3 #(
		.INIT('h2a)
	) name435 (
		_w2579_,
		_w2580_,
		_w2581_,
		_w2582_
	);
	LUT4 #(
		.INIT('h35ff)
	) name436 (
		\u4_mem_reg[2][10]/NET0131 ,
		\u4_mem_reg[3][10]/NET0131 ,
		\u4_rp_reg[1]/NET0131 ,
		\u4_rp_reg[2]/NET0131 ,
		_w2583_
	);
	LUT4 #(
		.INIT('hff35)
	) name437 (
		\u4_mem_reg[0][10]/NET0131 ,
		\u4_mem_reg[1][10]/NET0131 ,
		\u4_rp_reg[1]/NET0131 ,
		\u4_rp_reg[2]/NET0131 ,
		_w2584_
	);
	LUT4 #(
		.INIT('ha222)
	) name438 (
		_w2417_,
		_w2490_,
		_w2583_,
		_w2584_,
		_w2585_
	);
	LUT4 #(
		.INIT('h0b00)
	) name439 (
		_w2575_,
		_w2578_,
		_w2582_,
		_w2585_,
		_w2586_
	);
	LUT4 #(
		.INIT('h0b0f)
	) name440 (
		\u14_u1_en_out_l2_reg/P0001 ,
		\u14_u1_en_out_l_reg/NET0131 ,
		\u4_dout_reg[10]/P0001 ,
		\valid_s_reg/NET0131 ,
		_w2587_
	);
	LUT2 #(
		.INIT('h2)
	) name441 (
		\u13_occ0_r_reg[8]/NET0131 ,
		_w2587_,
		_w2588_
	);
	LUT2 #(
		.INIT('h4)
	) name442 (
		_w2586_,
		_w2588_,
		_w2589_
	);
	LUT4 #(
		.INIT('hc4cc)
	) name443 (
		\u4_mem_reg[2][23]/NET0131 ,
		\u4_rp_reg[0]/P0001 ,
		\u4_rp_reg[1]/NET0131 ,
		\u4_rp_reg[2]/NET0131 ,
		_w2590_
	);
	LUT3 #(
		.INIT('h02)
	) name444 (
		\u4_mem_reg[0][23]/NET0131 ,
		\u4_rp_reg[1]/NET0131 ,
		\u4_rp_reg[2]/NET0131 ,
		_w2591_
	);
	LUT4 #(
		.INIT('h3f5f)
	) name445 (
		\u4_mem_reg[1][23]/NET0131 ,
		\u4_mem_reg[3][23]/NET0131 ,
		\u4_rp_reg[1]/NET0131 ,
		\u4_rp_reg[2]/NET0131 ,
		_w2592_
	);
	LUT3 #(
		.INIT('h40)
	) name446 (
		_w2591_,
		_w2590_,
		_w2592_,
		_w2593_
	);
	LUT4 #(
		.INIT('hf35f)
	) name447 (
		\u4_mem_reg[1][7]/NET0131 ,
		\u4_mem_reg[2][7]/NET0131 ,
		\u4_rp_reg[1]/NET0131 ,
		\u4_rp_reg[2]/NET0131 ,
		_w2594_
	);
	LUT4 #(
		.INIT('h3ff5)
	) name448 (
		\u4_mem_reg[0][7]/NET0131 ,
		\u4_mem_reg[3][7]/NET0131 ,
		\u4_rp_reg[1]/NET0131 ,
		\u4_rp_reg[2]/NET0131 ,
		_w2595_
	);
	LUT4 #(
		.INIT('h8ccc)
	) name449 (
		\u4_rp_reg[0]/P0001 ,
		_w2418_,
		_w2594_,
		_w2595_,
		_w2596_
	);
	LUT4 #(
		.INIT('h3f5f)
	) name450 (
		\u4_mem_reg[1][9]/NET0131 ,
		\u4_mem_reg[3][9]/NET0131 ,
		\u4_rp_reg[1]/NET0131 ,
		\u4_rp_reg[2]/NET0131 ,
		_w2597_
	);
	LUT4 #(
		.INIT('hf3f5)
	) name451 (
		\u4_mem_reg[0][9]/NET0131 ,
		\u4_mem_reg[2][9]/NET0131 ,
		\u4_rp_reg[1]/NET0131 ,
		\u4_rp_reg[2]/NET0131 ,
		_w2598_
	);
	LUT3 #(
		.INIT('h2a)
	) name452 (
		_w2579_,
		_w2597_,
		_w2598_,
		_w2599_
	);
	LUT4 #(
		.INIT('h3f5f)
	) name453 (
		\u4_mem_reg[1][11]/NET0131 ,
		\u4_mem_reg[3][11]/NET0131 ,
		\u4_rp_reg[1]/NET0131 ,
		\u4_rp_reg[2]/NET0131 ,
		_w2600_
	);
	LUT4 #(
		.INIT('hf3f5)
	) name454 (
		\u4_mem_reg[0][11]/NET0131 ,
		\u4_mem_reg[2][11]/NET0131 ,
		\u4_rp_reg[1]/NET0131 ,
		\u4_rp_reg[2]/NET0131 ,
		_w2601_
	);
	LUT4 #(
		.INIT('ha222)
	) name455 (
		_w2417_,
		_w2490_,
		_w2600_,
		_w2601_,
		_w2602_
	);
	LUT4 #(
		.INIT('h0b00)
	) name456 (
		_w2593_,
		_w2596_,
		_w2599_,
		_w2602_,
		_w2603_
	);
	LUT4 #(
		.INIT('h0b0f)
	) name457 (
		\u14_u1_en_out_l2_reg/P0001 ,
		\u14_u1_en_out_l_reg/NET0131 ,
		\u4_dout_reg[11]/P0001 ,
		\valid_s_reg/NET0131 ,
		_w2604_
	);
	LUT2 #(
		.INIT('h2)
	) name458 (
		\u13_occ0_r_reg[8]/NET0131 ,
		_w2604_,
		_w2605_
	);
	LUT2 #(
		.INIT('h4)
	) name459 (
		_w2603_,
		_w2605_,
		_w2606_
	);
	LUT4 #(
		.INIT('hc4cc)
	) name460 (
		\u4_mem_reg[2][24]/NET0131 ,
		\u4_rp_reg[0]/P0001 ,
		\u4_rp_reg[1]/NET0131 ,
		\u4_rp_reg[2]/NET0131 ,
		_w2607_
	);
	LUT3 #(
		.INIT('h02)
	) name461 (
		\u4_mem_reg[0][24]/NET0131 ,
		\u4_rp_reg[1]/NET0131 ,
		\u4_rp_reg[2]/NET0131 ,
		_w2608_
	);
	LUT4 #(
		.INIT('h3f5f)
	) name462 (
		\u4_mem_reg[1][24]/NET0131 ,
		\u4_mem_reg[3][24]/NET0131 ,
		\u4_rp_reg[1]/NET0131 ,
		\u4_rp_reg[2]/NET0131 ,
		_w2609_
	);
	LUT3 #(
		.INIT('h40)
	) name463 (
		_w2608_,
		_w2607_,
		_w2609_,
		_w2610_
	);
	LUT4 #(
		.INIT('h8ccc)
	) name464 (
		\u4_rp_reg[0]/P0001 ,
		_w2418_,
		_w2580_,
		_w2581_,
		_w2611_
	);
	LUT3 #(
		.INIT('h70)
	) name465 (
		_w2583_,
		_w2584_,
		_w2579_,
		_w2612_
	);
	LUT4 #(
		.INIT('h35ff)
	) name466 (
		\u4_mem_reg[2][12]/NET0131 ,
		\u4_mem_reg[3][12]/NET0131 ,
		\u4_rp_reg[1]/NET0131 ,
		\u4_rp_reg[2]/NET0131 ,
		_w2613_
	);
	LUT4 #(
		.INIT('hff35)
	) name467 (
		\u4_mem_reg[0][12]/NET0131 ,
		\u4_mem_reg[1][12]/NET0131 ,
		\u4_rp_reg[1]/NET0131 ,
		\u4_rp_reg[2]/NET0131 ,
		_w2614_
	);
	LUT4 #(
		.INIT('ha222)
	) name468 (
		_w2417_,
		_w2490_,
		_w2613_,
		_w2614_,
		_w2615_
	);
	LUT4 #(
		.INIT('h0b00)
	) name469 (
		_w2610_,
		_w2611_,
		_w2612_,
		_w2615_,
		_w2616_
	);
	LUT4 #(
		.INIT('h0b0f)
	) name470 (
		\u14_u1_en_out_l2_reg/P0001 ,
		\u14_u1_en_out_l_reg/NET0131 ,
		\u4_dout_reg[12]/P0001 ,
		\valid_s_reg/NET0131 ,
		_w2617_
	);
	LUT2 #(
		.INIT('h2)
	) name471 (
		\u13_occ0_r_reg[8]/NET0131 ,
		_w2617_,
		_w2618_
	);
	LUT2 #(
		.INIT('h4)
	) name472 (
		_w2616_,
		_w2618_,
		_w2619_
	);
	LUT4 #(
		.INIT('hc4cc)
	) name473 (
		\u4_mem_reg[2][25]/NET0131 ,
		\u4_rp_reg[0]/P0001 ,
		\u4_rp_reg[1]/NET0131 ,
		\u4_rp_reg[2]/NET0131 ,
		_w2620_
	);
	LUT3 #(
		.INIT('h02)
	) name474 (
		\u4_mem_reg[0][25]/NET0131 ,
		\u4_rp_reg[1]/NET0131 ,
		\u4_rp_reg[2]/NET0131 ,
		_w2621_
	);
	LUT4 #(
		.INIT('h3f5f)
	) name475 (
		\u4_mem_reg[1][25]/NET0131 ,
		\u4_mem_reg[3][25]/NET0131 ,
		\u4_rp_reg[1]/NET0131 ,
		\u4_rp_reg[2]/NET0131 ,
		_w2622_
	);
	LUT3 #(
		.INIT('h40)
	) name476 (
		_w2621_,
		_w2620_,
		_w2622_,
		_w2623_
	);
	LUT4 #(
		.INIT('h8ccc)
	) name477 (
		\u4_rp_reg[0]/P0001 ,
		_w2418_,
		_w2597_,
		_w2598_,
		_w2624_
	);
	LUT3 #(
		.INIT('h2a)
	) name478 (
		_w2579_,
		_w2600_,
		_w2601_,
		_w2625_
	);
	LUT4 #(
		.INIT('h3f5f)
	) name479 (
		\u4_mem_reg[1][13]/NET0131 ,
		\u4_mem_reg[3][13]/NET0131 ,
		\u4_rp_reg[1]/NET0131 ,
		\u4_rp_reg[2]/NET0131 ,
		_w2626_
	);
	LUT4 #(
		.INIT('hf3f5)
	) name480 (
		\u4_mem_reg[0][13]/NET0131 ,
		\u4_mem_reg[2][13]/NET0131 ,
		\u4_rp_reg[1]/NET0131 ,
		\u4_rp_reg[2]/NET0131 ,
		_w2627_
	);
	LUT4 #(
		.INIT('ha222)
	) name481 (
		_w2417_,
		_w2490_,
		_w2626_,
		_w2627_,
		_w2628_
	);
	LUT4 #(
		.INIT('h0b00)
	) name482 (
		_w2623_,
		_w2624_,
		_w2625_,
		_w2628_,
		_w2629_
	);
	LUT4 #(
		.INIT('h0b0f)
	) name483 (
		\u14_u1_en_out_l2_reg/P0001 ,
		\u14_u1_en_out_l_reg/NET0131 ,
		\u4_dout_reg[13]/P0001 ,
		\valid_s_reg/NET0131 ,
		_w2630_
	);
	LUT2 #(
		.INIT('h2)
	) name484 (
		\u13_occ0_r_reg[8]/NET0131 ,
		_w2630_,
		_w2631_
	);
	LUT2 #(
		.INIT('h4)
	) name485 (
		_w2629_,
		_w2631_,
		_w2632_
	);
	LUT4 #(
		.INIT('hc4cc)
	) name486 (
		\u4_mem_reg[2][26]/NET0131 ,
		\u4_rp_reg[0]/P0001 ,
		\u4_rp_reg[1]/NET0131 ,
		\u4_rp_reg[2]/NET0131 ,
		_w2633_
	);
	LUT3 #(
		.INIT('h02)
	) name487 (
		\u4_mem_reg[0][26]/NET0131 ,
		\u4_rp_reg[1]/NET0131 ,
		\u4_rp_reg[2]/NET0131 ,
		_w2634_
	);
	LUT4 #(
		.INIT('h3f5f)
	) name488 (
		\u4_mem_reg[1][26]/NET0131 ,
		\u4_mem_reg[3][26]/NET0131 ,
		\u4_rp_reg[1]/NET0131 ,
		\u4_rp_reg[2]/NET0131 ,
		_w2635_
	);
	LUT3 #(
		.INIT('h40)
	) name489 (
		_w2634_,
		_w2633_,
		_w2635_,
		_w2636_
	);
	LUT4 #(
		.INIT('h8ccc)
	) name490 (
		\u4_rp_reg[0]/P0001 ,
		_w2418_,
		_w2583_,
		_w2584_,
		_w2637_
	);
	LUT3 #(
		.INIT('h2a)
	) name491 (
		_w2579_,
		_w2613_,
		_w2614_,
		_w2638_
	);
	LUT4 #(
		.INIT('hf35f)
	) name492 (
		\u4_mem_reg[1][14]/NET0131 ,
		\u4_mem_reg[2][14]/NET0131 ,
		\u4_rp_reg[1]/NET0131 ,
		\u4_rp_reg[2]/NET0131 ,
		_w2639_
	);
	LUT4 #(
		.INIT('h3ff5)
	) name493 (
		\u4_mem_reg[0][14]/NET0131 ,
		\u4_mem_reg[3][14]/NET0131 ,
		\u4_rp_reg[1]/NET0131 ,
		\u4_rp_reg[2]/NET0131 ,
		_w2640_
	);
	LUT4 #(
		.INIT('ha222)
	) name494 (
		_w2417_,
		_w2490_,
		_w2639_,
		_w2640_,
		_w2641_
	);
	LUT4 #(
		.INIT('h0b00)
	) name495 (
		_w2636_,
		_w2637_,
		_w2638_,
		_w2641_,
		_w2642_
	);
	LUT4 #(
		.INIT('h0b0f)
	) name496 (
		\u14_u1_en_out_l2_reg/P0001 ,
		\u14_u1_en_out_l_reg/NET0131 ,
		\u4_dout_reg[14]/P0001 ,
		\valid_s_reg/NET0131 ,
		_w2643_
	);
	LUT2 #(
		.INIT('h2)
	) name497 (
		\u13_occ0_r_reg[8]/NET0131 ,
		_w2643_,
		_w2644_
	);
	LUT2 #(
		.INIT('h4)
	) name498 (
		_w2642_,
		_w2644_,
		_w2645_
	);
	LUT4 #(
		.INIT('hc4cc)
	) name499 (
		\u4_mem_reg[2][27]/NET0131 ,
		\u4_rp_reg[0]/P0001 ,
		\u4_rp_reg[1]/NET0131 ,
		\u4_rp_reg[2]/NET0131 ,
		_w2646_
	);
	LUT3 #(
		.INIT('h02)
	) name500 (
		\u4_mem_reg[0][27]/NET0131 ,
		\u4_rp_reg[1]/NET0131 ,
		\u4_rp_reg[2]/NET0131 ,
		_w2647_
	);
	LUT4 #(
		.INIT('h3f5f)
	) name501 (
		\u4_mem_reg[1][27]/NET0131 ,
		\u4_mem_reg[3][27]/NET0131 ,
		\u4_rp_reg[1]/NET0131 ,
		\u4_rp_reg[2]/NET0131 ,
		_w2648_
	);
	LUT3 #(
		.INIT('h40)
	) name502 (
		_w2647_,
		_w2646_,
		_w2648_,
		_w2649_
	);
	LUT4 #(
		.INIT('h8ccc)
	) name503 (
		\u4_rp_reg[0]/P0001 ,
		_w2418_,
		_w2600_,
		_w2601_,
		_w2650_
	);
	LUT3 #(
		.INIT('h2a)
	) name504 (
		_w2579_,
		_w2626_,
		_w2627_,
		_w2651_
	);
	LUT4 #(
		.INIT('hf3f5)
	) name505 (
		\u4_mem_reg[0][15]/NET0131 ,
		\u4_mem_reg[2][15]/NET0131 ,
		\u4_rp_reg[1]/NET0131 ,
		\u4_rp_reg[2]/NET0131 ,
		_w2652_
	);
	LUT4 #(
		.INIT('h3f5f)
	) name506 (
		\u4_mem_reg[1][15]/NET0131 ,
		\u4_mem_reg[3][15]/NET0131 ,
		\u4_rp_reg[1]/NET0131 ,
		\u4_rp_reg[2]/NET0131 ,
		_w2653_
	);
	LUT4 #(
		.INIT('ha222)
	) name507 (
		_w2417_,
		_w2490_,
		_w2652_,
		_w2653_,
		_w2654_
	);
	LUT4 #(
		.INIT('h0b00)
	) name508 (
		_w2649_,
		_w2650_,
		_w2651_,
		_w2654_,
		_w2655_
	);
	LUT4 #(
		.INIT('h0b0f)
	) name509 (
		\u14_u1_en_out_l2_reg/P0001 ,
		\u14_u1_en_out_l_reg/NET0131 ,
		\u4_dout_reg[15]/P0001 ,
		\valid_s_reg/NET0131 ,
		_w2656_
	);
	LUT2 #(
		.INIT('h2)
	) name510 (
		\u13_occ0_r_reg[8]/NET0131 ,
		_w2656_,
		_w2657_
	);
	LUT2 #(
		.INIT('h4)
	) name511 (
		_w2655_,
		_w2657_,
		_w2658_
	);
	LUT4 #(
		.INIT('hc4cc)
	) name512 (
		\u4_mem_reg[2][28]/NET0131 ,
		\u4_rp_reg[0]/P0001 ,
		\u4_rp_reg[1]/NET0131 ,
		\u4_rp_reg[2]/NET0131 ,
		_w2659_
	);
	LUT3 #(
		.INIT('h02)
	) name513 (
		\u4_mem_reg[0][28]/NET0131 ,
		\u4_rp_reg[1]/NET0131 ,
		\u4_rp_reg[2]/NET0131 ,
		_w2660_
	);
	LUT4 #(
		.INIT('h3f5f)
	) name514 (
		\u4_mem_reg[1][28]/NET0131 ,
		\u4_mem_reg[3][28]/NET0131 ,
		\u4_rp_reg[1]/NET0131 ,
		\u4_rp_reg[2]/NET0131 ,
		_w2661_
	);
	LUT3 #(
		.INIT('h40)
	) name515 (
		_w2660_,
		_w2659_,
		_w2661_,
		_w2662_
	);
	LUT4 #(
		.INIT('h8ccc)
	) name516 (
		\u4_rp_reg[0]/P0001 ,
		_w2418_,
		_w2613_,
		_w2614_,
		_w2663_
	);
	LUT3 #(
		.INIT('h2a)
	) name517 (
		_w2579_,
		_w2639_,
		_w2640_,
		_w2664_
	);
	LUT4 #(
		.INIT('h35ff)
	) name518 (
		\u4_mem_reg[2][16]/NET0131 ,
		\u4_mem_reg[3][16]/NET0131 ,
		\u4_rp_reg[1]/NET0131 ,
		\u4_rp_reg[2]/NET0131 ,
		_w2665_
	);
	LUT4 #(
		.INIT('hff35)
	) name519 (
		\u4_mem_reg[0][16]/NET0131 ,
		\u4_mem_reg[1][16]/NET0131 ,
		\u4_rp_reg[1]/NET0131 ,
		\u4_rp_reg[2]/NET0131 ,
		_w2666_
	);
	LUT4 #(
		.INIT('ha222)
	) name520 (
		_w2417_,
		_w2490_,
		_w2665_,
		_w2666_,
		_w2667_
	);
	LUT4 #(
		.INIT('h0b00)
	) name521 (
		_w2662_,
		_w2663_,
		_w2664_,
		_w2667_,
		_w2668_
	);
	LUT4 #(
		.INIT('h0b0f)
	) name522 (
		\u14_u1_en_out_l2_reg/P0001 ,
		\u14_u1_en_out_l_reg/NET0131 ,
		\u4_dout_reg[16]/P0001 ,
		\valid_s_reg/NET0131 ,
		_w2669_
	);
	LUT2 #(
		.INIT('h2)
	) name523 (
		\u13_occ0_r_reg[8]/NET0131 ,
		_w2669_,
		_w2670_
	);
	LUT2 #(
		.INIT('h4)
	) name524 (
		_w2668_,
		_w2670_,
		_w2671_
	);
	LUT4 #(
		.INIT('hc4cc)
	) name525 (
		\u4_mem_reg[2][29]/NET0131 ,
		\u4_rp_reg[0]/P0001 ,
		\u4_rp_reg[1]/NET0131 ,
		\u4_rp_reg[2]/NET0131 ,
		_w2672_
	);
	LUT3 #(
		.INIT('h02)
	) name526 (
		\u4_mem_reg[0][29]/NET0131 ,
		\u4_rp_reg[1]/NET0131 ,
		\u4_rp_reg[2]/NET0131 ,
		_w2673_
	);
	LUT4 #(
		.INIT('h3f5f)
	) name527 (
		\u4_mem_reg[1][29]/NET0131 ,
		\u4_mem_reg[3][29]/NET0131 ,
		\u4_rp_reg[1]/NET0131 ,
		\u4_rp_reg[2]/NET0131 ,
		_w2674_
	);
	LUT3 #(
		.INIT('h40)
	) name528 (
		_w2673_,
		_w2672_,
		_w2674_,
		_w2675_
	);
	LUT4 #(
		.INIT('h8ccc)
	) name529 (
		\u4_rp_reg[0]/P0001 ,
		_w2418_,
		_w2626_,
		_w2627_,
		_w2676_
	);
	LUT3 #(
		.INIT('h2a)
	) name530 (
		_w2579_,
		_w2652_,
		_w2653_,
		_w2677_
	);
	LUT4 #(
		.INIT('h35ff)
	) name531 (
		\u4_mem_reg[2][17]/NET0131 ,
		\u4_mem_reg[3][17]/NET0131 ,
		\u4_rp_reg[1]/NET0131 ,
		\u4_rp_reg[2]/NET0131 ,
		_w2678_
	);
	LUT4 #(
		.INIT('hff35)
	) name532 (
		\u4_mem_reg[0][17]/NET0131 ,
		\u4_mem_reg[1][17]/NET0131 ,
		\u4_rp_reg[1]/NET0131 ,
		\u4_rp_reg[2]/NET0131 ,
		_w2679_
	);
	LUT4 #(
		.INIT('ha222)
	) name533 (
		_w2417_,
		_w2490_,
		_w2678_,
		_w2679_,
		_w2680_
	);
	LUT4 #(
		.INIT('h0b00)
	) name534 (
		_w2675_,
		_w2676_,
		_w2677_,
		_w2680_,
		_w2681_
	);
	LUT4 #(
		.INIT('h0b0f)
	) name535 (
		\u14_u1_en_out_l2_reg/P0001 ,
		\u14_u1_en_out_l_reg/NET0131 ,
		\u4_dout_reg[17]/P0001 ,
		\valid_s_reg/NET0131 ,
		_w2682_
	);
	LUT2 #(
		.INIT('h2)
	) name536 (
		\u13_occ0_r_reg[8]/NET0131 ,
		_w2682_,
		_w2683_
	);
	LUT2 #(
		.INIT('h4)
	) name537 (
		_w2681_,
		_w2683_,
		_w2684_
	);
	LUT2 #(
		.INIT('h8)
	) name538 (
		\in_valid_s_reg[0]/NET0131 ,
		\u14_u6_en_out_l_reg/NET0131 ,
		_w2685_
	);
	LUT3 #(
		.INIT('h20)
	) name539 (
		\in_valid_s_reg[0]/NET0131 ,
		\u14_u6_en_out_l2_reg/P0001 ,
		\u14_u6_en_out_l_reg/NET0131 ,
		_w2686_
	);
	LUT2 #(
		.INIT('h1)
	) name540 (
		\u13_icc_r_reg[2]/NET0131 ,
		\u13_icc_r_reg[3]/NET0131 ,
		_w2687_
	);
	LUT3 #(
		.INIT('h01)
	) name541 (
		\u13_icc_r_reg[2]/NET0131 ,
		\u13_icc_r_reg[3]/NET0131 ,
		\u9_wp_reg[0]/NET0131 ,
		_w2688_
	);
	LUT2 #(
		.INIT('h2)
	) name542 (
		_w2686_,
		_w2688_,
		_w2689_
	);
	LUT3 #(
		.INIT('h08)
	) name543 (
		\u9_wp_reg[1]/P0001 ,
		_w2686_,
		_w2688_,
		_w2690_
	);
	LUT4 #(
		.INIT('h0080)
	) name544 (
		\u9_wp_reg[1]/P0001 ,
		\u9_wp_reg[2]/P0001 ,
		_w2686_,
		_w2688_,
		_w2691_
	);
	LUT3 #(
		.INIT('h28)
	) name545 (
		\u13_icc_r_reg[0]/NET0131 ,
		\u9_wp_reg[2]/P0001 ,
		_w2690_,
		_w2692_
	);
	LUT4 #(
		.INIT('hc4cc)
	) name546 (
		\u4_mem_reg[2][30]/NET0131 ,
		\u4_rp_reg[0]/P0001 ,
		\u4_rp_reg[1]/NET0131 ,
		\u4_rp_reg[2]/NET0131 ,
		_w2693_
	);
	LUT3 #(
		.INIT('h02)
	) name547 (
		\u4_mem_reg[0][30]/NET0131 ,
		\u4_rp_reg[1]/NET0131 ,
		\u4_rp_reg[2]/NET0131 ,
		_w2694_
	);
	LUT4 #(
		.INIT('h3f5f)
	) name548 (
		\u4_mem_reg[1][30]/NET0131 ,
		\u4_mem_reg[3][30]/NET0131 ,
		\u4_rp_reg[1]/NET0131 ,
		\u4_rp_reg[2]/NET0131 ,
		_w2695_
	);
	LUT3 #(
		.INIT('h40)
	) name549 (
		_w2694_,
		_w2693_,
		_w2695_,
		_w2696_
	);
	LUT4 #(
		.INIT('h8ccc)
	) name550 (
		\u4_rp_reg[0]/P0001 ,
		_w2418_,
		_w2639_,
		_w2640_,
		_w2697_
	);
	LUT3 #(
		.INIT('h2a)
	) name551 (
		_w2579_,
		_w2665_,
		_w2666_,
		_w2698_
	);
	LUT4 #(
		.INIT('h3f5f)
	) name552 (
		\u4_mem_reg[1][18]/NET0131 ,
		\u4_mem_reg[3][18]/NET0131 ,
		\u4_rp_reg[1]/NET0131 ,
		\u4_rp_reg[2]/NET0131 ,
		_w2699_
	);
	LUT4 #(
		.INIT('hf3f5)
	) name553 (
		\u4_mem_reg[0][18]/NET0131 ,
		\u4_mem_reg[2][18]/NET0131 ,
		\u4_rp_reg[1]/NET0131 ,
		\u4_rp_reg[2]/NET0131 ,
		_w2700_
	);
	LUT4 #(
		.INIT('ha222)
	) name554 (
		_w2417_,
		_w2490_,
		_w2699_,
		_w2700_,
		_w2701_
	);
	LUT4 #(
		.INIT('h0b00)
	) name555 (
		_w2696_,
		_w2697_,
		_w2698_,
		_w2701_,
		_w2702_
	);
	LUT4 #(
		.INIT('h0b0f)
	) name556 (
		\u14_u1_en_out_l2_reg/P0001 ,
		\u14_u1_en_out_l_reg/NET0131 ,
		\u4_dout_reg[18]/P0001 ,
		\valid_s_reg/NET0131 ,
		_w2703_
	);
	LUT2 #(
		.INIT('h2)
	) name557 (
		\u13_occ0_r_reg[8]/NET0131 ,
		_w2703_,
		_w2704_
	);
	LUT2 #(
		.INIT('h4)
	) name558 (
		_w2702_,
		_w2704_,
		_w2705_
	);
	LUT4 #(
		.INIT('hc4cc)
	) name559 (
		\u4_mem_reg[2][31]/NET0131 ,
		\u4_rp_reg[0]/P0001 ,
		\u4_rp_reg[1]/NET0131 ,
		\u4_rp_reg[2]/NET0131 ,
		_w2706_
	);
	LUT3 #(
		.INIT('h02)
	) name560 (
		\u4_mem_reg[0][31]/NET0131 ,
		\u4_rp_reg[1]/NET0131 ,
		\u4_rp_reg[2]/NET0131 ,
		_w2707_
	);
	LUT4 #(
		.INIT('h3f5f)
	) name561 (
		\u4_mem_reg[1][31]/NET0131 ,
		\u4_mem_reg[3][31]/NET0131 ,
		\u4_rp_reg[1]/NET0131 ,
		\u4_rp_reg[2]/NET0131 ,
		_w2708_
	);
	LUT3 #(
		.INIT('h40)
	) name562 (
		_w2707_,
		_w2706_,
		_w2708_,
		_w2709_
	);
	LUT4 #(
		.INIT('h8ccc)
	) name563 (
		\u4_rp_reg[0]/P0001 ,
		_w2418_,
		_w2652_,
		_w2653_,
		_w2710_
	);
	LUT3 #(
		.INIT('h2a)
	) name564 (
		_w2579_,
		_w2678_,
		_w2679_,
		_w2711_
	);
	LUT4 #(
		.INIT('h35ff)
	) name565 (
		\u4_mem_reg[2][19]/NET0131 ,
		\u4_mem_reg[3][19]/NET0131 ,
		\u4_rp_reg[1]/NET0131 ,
		\u4_rp_reg[2]/NET0131 ,
		_w2712_
	);
	LUT4 #(
		.INIT('hff35)
	) name566 (
		\u4_mem_reg[0][19]/NET0131 ,
		\u4_mem_reg[1][19]/NET0131 ,
		\u4_rp_reg[1]/NET0131 ,
		\u4_rp_reg[2]/NET0131 ,
		_w2713_
	);
	LUT4 #(
		.INIT('ha222)
	) name567 (
		_w2417_,
		_w2490_,
		_w2712_,
		_w2713_,
		_w2714_
	);
	LUT4 #(
		.INIT('h0b00)
	) name568 (
		_w2709_,
		_w2710_,
		_w2711_,
		_w2714_,
		_w2715_
	);
	LUT4 #(
		.INIT('h0b0f)
	) name569 (
		\u14_u1_en_out_l2_reg/P0001 ,
		\u14_u1_en_out_l_reg/NET0131 ,
		\u4_dout_reg[19]/P0001 ,
		\valid_s_reg/NET0131 ,
		_w2716_
	);
	LUT2 #(
		.INIT('h2)
	) name570 (
		\u13_occ0_r_reg[8]/NET0131 ,
		_w2716_,
		_w2717_
	);
	LUT2 #(
		.INIT('h4)
	) name571 (
		_w2715_,
		_w2717_,
		_w2718_
	);
	LUT4 #(
		.INIT('hff35)
	) name572 (
		\u4_mem_reg[0][2]/NET0131 ,
		\u4_mem_reg[1][2]/NET0131 ,
		\u4_rp_reg[1]/NET0131 ,
		\u4_rp_reg[2]/NET0131 ,
		_w2719_
	);
	LUT4 #(
		.INIT('h35ff)
	) name573 (
		\u4_mem_reg[2][2]/NET0131 ,
		\u4_mem_reg[3][2]/NET0131 ,
		\u4_rp_reg[1]/NET0131 ,
		\u4_rp_reg[2]/NET0131 ,
		_w2720_
	);
	LUT3 #(
		.INIT('h2a)
	) name574 (
		_w2490_,
		_w2719_,
		_w2720_,
		_w2721_
	);
	LUT4 #(
		.INIT('h80aa)
	) name575 (
		_w2417_,
		_w2488_,
		_w2489_,
		_w2579_,
		_w2722_
	);
	LUT4 #(
		.INIT('h0b0f)
	) name576 (
		\u14_u1_en_out_l2_reg/P0001 ,
		\u14_u1_en_out_l_reg/NET0131 ,
		\u4_dout_reg[2]/P0001 ,
		\valid_s_reg/NET0131 ,
		_w2723_
	);
	LUT2 #(
		.INIT('h2)
	) name577 (
		\u13_occ0_r_reg[8]/NET0131 ,
		_w2723_,
		_w2724_
	);
	LUT3 #(
		.INIT('hb0)
	) name578 (
		_w2721_,
		_w2722_,
		_w2724_,
		_w2725_
	);
	LUT3 #(
		.INIT('h70)
	) name579 (
		_w2495_,
		_w2496_,
		_w2579_,
		_w2726_
	);
	LUT4 #(
		.INIT('h35ff)
	) name580 (
		\u4_mem_reg[2][3]/NET0131 ,
		\u4_mem_reg[3][3]/NET0131 ,
		\u4_rp_reg[1]/NET0131 ,
		\u4_rp_reg[2]/NET0131 ,
		_w2727_
	);
	LUT4 #(
		.INIT('hff35)
	) name581 (
		\u4_mem_reg[0][3]/NET0131 ,
		\u4_mem_reg[1][3]/NET0131 ,
		\u4_rp_reg[1]/NET0131 ,
		\u4_rp_reg[2]/NET0131 ,
		_w2728_
	);
	LUT4 #(
		.INIT('ha222)
	) name582 (
		_w2417_,
		_w2490_,
		_w2727_,
		_w2728_,
		_w2729_
	);
	LUT4 #(
		.INIT('h0b0f)
	) name583 (
		\u14_u1_en_out_l2_reg/P0001 ,
		\u14_u1_en_out_l_reg/NET0131 ,
		\u4_dout_reg[3]/P0001 ,
		\valid_s_reg/NET0131 ,
		_w2730_
	);
	LUT2 #(
		.INIT('h2)
	) name584 (
		\u13_occ0_r_reg[8]/NET0131 ,
		_w2730_,
		_w2731_
	);
	LUT3 #(
		.INIT('hb0)
	) name585 (
		_w2726_,
		_w2729_,
		_w2731_,
		_w2732_
	);
	LUT3 #(
		.INIT('h80)
	) name586 (
		\u4_rp_reg[0]/P0001 ,
		_w2665_,
		_w2666_,
		_w2733_
	);
	LUT4 #(
		.INIT('h8ccc)
	) name587 (
		\u4_rp_reg[0]/P0001 ,
		_w2418_,
		_w2488_,
		_w2489_,
		_w2734_
	);
	LUT3 #(
		.INIT('h2a)
	) name588 (
		_w2579_,
		_w2719_,
		_w2720_,
		_w2735_
	);
	LUT4 #(
		.INIT('h35ff)
	) name589 (
		\u4_mem_reg[2][4]/NET0131 ,
		\u4_mem_reg[3][4]/NET0131 ,
		\u4_rp_reg[1]/NET0131 ,
		\u4_rp_reg[2]/NET0131 ,
		_w2736_
	);
	LUT4 #(
		.INIT('hff35)
	) name590 (
		\u4_mem_reg[0][4]/NET0131 ,
		\u4_mem_reg[1][4]/NET0131 ,
		\u4_rp_reg[1]/NET0131 ,
		\u4_rp_reg[2]/NET0131 ,
		_w2737_
	);
	LUT4 #(
		.INIT('ha222)
	) name591 (
		_w2417_,
		_w2490_,
		_w2736_,
		_w2737_,
		_w2738_
	);
	LUT4 #(
		.INIT('h0b00)
	) name592 (
		_w2733_,
		_w2734_,
		_w2735_,
		_w2738_,
		_w2739_
	);
	LUT4 #(
		.INIT('h0b0f)
	) name593 (
		\u14_u1_en_out_l2_reg/P0001 ,
		\u14_u1_en_out_l_reg/NET0131 ,
		\u4_dout_reg[4]/P0001 ,
		\valid_s_reg/NET0131 ,
		_w2740_
	);
	LUT2 #(
		.INIT('h2)
	) name594 (
		\u13_occ0_r_reg[8]/NET0131 ,
		_w2740_,
		_w2741_
	);
	LUT2 #(
		.INIT('h4)
	) name595 (
		_w2739_,
		_w2741_,
		_w2742_
	);
	LUT3 #(
		.INIT('h80)
	) name596 (
		\u4_rp_reg[0]/P0001 ,
		_w2678_,
		_w2679_,
		_w2743_
	);
	LUT4 #(
		.INIT('h8ccc)
	) name597 (
		\u4_rp_reg[0]/P0001 ,
		_w2418_,
		_w2495_,
		_w2496_,
		_w2744_
	);
	LUT3 #(
		.INIT('h2a)
	) name598 (
		_w2579_,
		_w2727_,
		_w2728_,
		_w2745_
	);
	LUT4 #(
		.INIT('hf35f)
	) name599 (
		\u4_mem_reg[1][5]/NET0131 ,
		\u4_mem_reg[2][5]/NET0131 ,
		\u4_rp_reg[1]/NET0131 ,
		\u4_rp_reg[2]/NET0131 ,
		_w2746_
	);
	LUT4 #(
		.INIT('h3ff5)
	) name600 (
		\u4_mem_reg[0][5]/NET0131 ,
		\u4_mem_reg[3][5]/NET0131 ,
		\u4_rp_reg[1]/NET0131 ,
		\u4_rp_reg[2]/NET0131 ,
		_w2747_
	);
	LUT4 #(
		.INIT('ha222)
	) name601 (
		_w2417_,
		_w2490_,
		_w2746_,
		_w2747_,
		_w2748_
	);
	LUT4 #(
		.INIT('h0b00)
	) name602 (
		_w2743_,
		_w2744_,
		_w2745_,
		_w2748_,
		_w2749_
	);
	LUT4 #(
		.INIT('h0b0f)
	) name603 (
		\u14_u1_en_out_l2_reg/P0001 ,
		\u14_u1_en_out_l_reg/NET0131 ,
		\u4_dout_reg[5]/P0001 ,
		\valid_s_reg/NET0131 ,
		_w2750_
	);
	LUT2 #(
		.INIT('h2)
	) name604 (
		\u13_occ0_r_reg[8]/NET0131 ,
		_w2750_,
		_w2751_
	);
	LUT2 #(
		.INIT('h4)
	) name605 (
		_w2749_,
		_w2751_,
		_w2752_
	);
	LUT3 #(
		.INIT('h80)
	) name606 (
		\u4_rp_reg[0]/P0001 ,
		_w2699_,
		_w2700_,
		_w2753_
	);
	LUT4 #(
		.INIT('h8ccc)
	) name607 (
		\u4_rp_reg[0]/P0001 ,
		_w2418_,
		_w2719_,
		_w2720_,
		_w2754_
	);
	LUT3 #(
		.INIT('h2a)
	) name608 (
		_w2579_,
		_w2736_,
		_w2737_,
		_w2755_
	);
	LUT4 #(
		.INIT('ha222)
	) name609 (
		_w2417_,
		_w2490_,
		_w2576_,
		_w2577_,
		_w2756_
	);
	LUT4 #(
		.INIT('h0b00)
	) name610 (
		_w2753_,
		_w2754_,
		_w2755_,
		_w2756_,
		_w2757_
	);
	LUT4 #(
		.INIT('h0b0f)
	) name611 (
		\u14_u1_en_out_l2_reg/P0001 ,
		\u14_u1_en_out_l_reg/NET0131 ,
		\u4_dout_reg[6]/P0001 ,
		\valid_s_reg/NET0131 ,
		_w2758_
	);
	LUT2 #(
		.INIT('h2)
	) name612 (
		\u13_occ0_r_reg[8]/NET0131 ,
		_w2758_,
		_w2759_
	);
	LUT2 #(
		.INIT('h4)
	) name613 (
		_w2757_,
		_w2759_,
		_w2760_
	);
	LUT3 #(
		.INIT('h80)
	) name614 (
		\u4_rp_reg[0]/P0001 ,
		_w2712_,
		_w2713_,
		_w2761_
	);
	LUT4 #(
		.INIT('h8ccc)
	) name615 (
		\u4_rp_reg[0]/P0001 ,
		_w2418_,
		_w2727_,
		_w2728_,
		_w2762_
	);
	LUT3 #(
		.INIT('h2a)
	) name616 (
		_w2579_,
		_w2746_,
		_w2747_,
		_w2763_
	);
	LUT4 #(
		.INIT('ha222)
	) name617 (
		_w2417_,
		_w2490_,
		_w2594_,
		_w2595_,
		_w2764_
	);
	LUT4 #(
		.INIT('h0b00)
	) name618 (
		_w2761_,
		_w2762_,
		_w2763_,
		_w2764_,
		_w2765_
	);
	LUT4 #(
		.INIT('h0b0f)
	) name619 (
		\u14_u1_en_out_l2_reg/P0001 ,
		\u14_u1_en_out_l_reg/NET0131 ,
		\u4_dout_reg[7]/P0001 ,
		\valid_s_reg/NET0131 ,
		_w2766_
	);
	LUT2 #(
		.INIT('h2)
	) name620 (
		\u13_occ0_r_reg[8]/NET0131 ,
		_w2766_,
		_w2767_
	);
	LUT2 #(
		.INIT('h4)
	) name621 (
		_w2765_,
		_w2767_,
		_w2768_
	);
	LUT4 #(
		.INIT('hc4cc)
	) name622 (
		\u4_mem_reg[2][20]/NET0131 ,
		\u4_rp_reg[0]/P0001 ,
		\u4_rp_reg[1]/NET0131 ,
		\u4_rp_reg[2]/NET0131 ,
		_w2769_
	);
	LUT3 #(
		.INIT('h02)
	) name623 (
		\u4_mem_reg[0][20]/NET0131 ,
		\u4_rp_reg[1]/NET0131 ,
		\u4_rp_reg[2]/NET0131 ,
		_w2770_
	);
	LUT4 #(
		.INIT('h3f5f)
	) name624 (
		\u4_mem_reg[1][20]/NET0131 ,
		\u4_mem_reg[3][20]/NET0131 ,
		\u4_rp_reg[1]/NET0131 ,
		\u4_rp_reg[2]/NET0131 ,
		_w2771_
	);
	LUT3 #(
		.INIT('h40)
	) name625 (
		_w2770_,
		_w2769_,
		_w2771_,
		_w2772_
	);
	LUT4 #(
		.INIT('h8ccc)
	) name626 (
		\u4_rp_reg[0]/P0001 ,
		_w2418_,
		_w2736_,
		_w2737_,
		_w2773_
	);
	LUT3 #(
		.INIT('h70)
	) name627 (
		_w2576_,
		_w2577_,
		_w2579_,
		_w2774_
	);
	LUT4 #(
		.INIT('ha222)
	) name628 (
		_w2417_,
		_w2490_,
		_w2580_,
		_w2581_,
		_w2775_
	);
	LUT4 #(
		.INIT('h0b00)
	) name629 (
		_w2772_,
		_w2773_,
		_w2774_,
		_w2775_,
		_w2776_
	);
	LUT4 #(
		.INIT('h0b0f)
	) name630 (
		\u14_u1_en_out_l2_reg/P0001 ,
		\u14_u1_en_out_l_reg/NET0131 ,
		\u4_dout_reg[8]/P0001 ,
		\valid_s_reg/NET0131 ,
		_w2777_
	);
	LUT2 #(
		.INIT('h2)
	) name631 (
		\u13_occ0_r_reg[8]/NET0131 ,
		_w2777_,
		_w2778_
	);
	LUT2 #(
		.INIT('h4)
	) name632 (
		_w2776_,
		_w2778_,
		_w2779_
	);
	LUT4 #(
		.INIT('hc4cc)
	) name633 (
		\u4_mem_reg[2][21]/NET0131 ,
		\u4_rp_reg[0]/P0001 ,
		\u4_rp_reg[1]/NET0131 ,
		\u4_rp_reg[2]/NET0131 ,
		_w2780_
	);
	LUT3 #(
		.INIT('h02)
	) name634 (
		\u4_mem_reg[0][21]/NET0131 ,
		\u4_rp_reg[1]/NET0131 ,
		\u4_rp_reg[2]/NET0131 ,
		_w2781_
	);
	LUT4 #(
		.INIT('h3f5f)
	) name635 (
		\u4_mem_reg[1][21]/NET0131 ,
		\u4_mem_reg[3][21]/NET0131 ,
		\u4_rp_reg[1]/NET0131 ,
		\u4_rp_reg[2]/NET0131 ,
		_w2782_
	);
	LUT3 #(
		.INIT('h40)
	) name636 (
		_w2781_,
		_w2780_,
		_w2782_,
		_w2783_
	);
	LUT4 #(
		.INIT('h8ccc)
	) name637 (
		\u4_rp_reg[0]/P0001 ,
		_w2418_,
		_w2746_,
		_w2747_,
		_w2784_
	);
	LUT3 #(
		.INIT('h2a)
	) name638 (
		_w2579_,
		_w2594_,
		_w2595_,
		_w2785_
	);
	LUT4 #(
		.INIT('ha222)
	) name639 (
		_w2417_,
		_w2490_,
		_w2597_,
		_w2598_,
		_w2786_
	);
	LUT4 #(
		.INIT('h0b00)
	) name640 (
		_w2783_,
		_w2784_,
		_w2785_,
		_w2786_,
		_w2787_
	);
	LUT4 #(
		.INIT('h0b0f)
	) name641 (
		\u14_u1_en_out_l2_reg/P0001 ,
		\u14_u1_en_out_l_reg/NET0131 ,
		\u4_dout_reg[9]/P0001 ,
		\valid_s_reg/NET0131 ,
		_w2788_
	);
	LUT2 #(
		.INIT('h2)
	) name642 (
		\u13_occ0_r_reg[8]/NET0131 ,
		_w2788_,
		_w2789_
	);
	LUT2 #(
		.INIT('h4)
	) name643 (
		_w2787_,
		_w2789_,
		_w2790_
	);
	LUT2 #(
		.INIT('h8)
	) name644 (
		\in_valid_s_reg[1]/NET0131 ,
		\u14_u7_en_out_l_reg/NET0131 ,
		_w2791_
	);
	LUT3 #(
		.INIT('h20)
	) name645 (
		\in_valid_s_reg[1]/NET0131 ,
		\u14_u7_en_out_l2_reg/P0001 ,
		\u14_u7_en_out_l_reg/NET0131 ,
		_w2792_
	);
	LUT2 #(
		.INIT('h1)
	) name646 (
		\u13_icc_r_reg[10]/NET0131 ,
		\u13_icc_r_reg[11]/NET0131 ,
		_w2793_
	);
	LUT3 #(
		.INIT('h01)
	) name647 (
		\u10_wp_reg[0]/NET0131 ,
		\u13_icc_r_reg[10]/NET0131 ,
		\u13_icc_r_reg[11]/NET0131 ,
		_w2794_
	);
	LUT2 #(
		.INIT('h2)
	) name648 (
		_w2792_,
		_w2794_,
		_w2795_
	);
	LUT3 #(
		.INIT('h08)
	) name649 (
		\u10_wp_reg[1]/P0001 ,
		_w2792_,
		_w2794_,
		_w2796_
	);
	LUT4 #(
		.INIT('h0080)
	) name650 (
		\u10_wp_reg[1]/P0001 ,
		\u10_wp_reg[2]/P0001 ,
		_w2792_,
		_w2794_,
		_w2797_
	);
	LUT3 #(
		.INIT('h48)
	) name651 (
		\u10_wp_reg[2]/P0001 ,
		\u13_icc_r_reg[8]/NET0131 ,
		_w2796_,
		_w2798_
	);
	LUT4 #(
		.INIT('hc4cc)
	) name652 (
		\u5_mem_reg[2][22]/NET0131 ,
		\u5_rp_reg[0]/P0001 ,
		\u5_rp_reg[1]/NET0131 ,
		\u5_rp_reg[2]/NET0131 ,
		_w2799_
	);
	LUT3 #(
		.INIT('h02)
	) name653 (
		\u5_mem_reg[0][22]/NET0131 ,
		\u5_rp_reg[1]/NET0131 ,
		\u5_rp_reg[2]/NET0131 ,
		_w2800_
	);
	LUT4 #(
		.INIT('h3f5f)
	) name654 (
		\u5_mem_reg[1][22]/NET0131 ,
		\u5_mem_reg[3][22]/NET0131 ,
		\u5_rp_reg[1]/NET0131 ,
		\u5_rp_reg[2]/NET0131 ,
		_w2801_
	);
	LUT3 #(
		.INIT('h40)
	) name655 (
		_w2800_,
		_w2799_,
		_w2801_,
		_w2802_
	);
	LUT4 #(
		.INIT('hf35f)
	) name656 (
		\u5_mem_reg[1][6]/NET0131 ,
		\u5_mem_reg[2][6]/NET0131 ,
		\u5_rp_reg[1]/NET0131 ,
		\u5_rp_reg[2]/NET0131 ,
		_w2803_
	);
	LUT4 #(
		.INIT('h3ff5)
	) name657 (
		\u5_mem_reg[0][6]/NET0131 ,
		\u5_mem_reg[3][6]/NET0131 ,
		\u5_rp_reg[1]/NET0131 ,
		\u5_rp_reg[2]/NET0131 ,
		_w2804_
	);
	LUT4 #(
		.INIT('h8ccc)
	) name658 (
		\u5_rp_reg[0]/P0001 ,
		_w2427_,
		_w2803_,
		_w2804_,
		_w2805_
	);
	LUT2 #(
		.INIT('h2)
	) name659 (
		\u13_occ0_r_reg[18]/NET0131 ,
		\u13_occ0_r_reg[19]/NET0131 ,
		_w2806_
	);
	LUT4 #(
		.INIT('hf35f)
	) name660 (
		\u5_mem_reg[1][8]/NET0131 ,
		\u5_mem_reg[2][8]/NET0131 ,
		\u5_rp_reg[1]/NET0131 ,
		\u5_rp_reg[2]/NET0131 ,
		_w2807_
	);
	LUT4 #(
		.INIT('h3ff5)
	) name661 (
		\u5_mem_reg[0][8]/NET0131 ,
		\u5_mem_reg[3][8]/NET0131 ,
		\u5_rp_reg[1]/NET0131 ,
		\u5_rp_reg[2]/NET0131 ,
		_w2808_
	);
	LUT3 #(
		.INIT('h2a)
	) name662 (
		_w2806_,
		_w2807_,
		_w2808_,
		_w2809_
	);
	LUT4 #(
		.INIT('hf35f)
	) name663 (
		\u5_mem_reg[1][10]/NET0131 ,
		\u5_mem_reg[2][10]/NET0131 ,
		\u5_rp_reg[1]/NET0131 ,
		\u5_rp_reg[2]/NET0131 ,
		_w2810_
	);
	LUT4 #(
		.INIT('h3ff5)
	) name664 (
		\u5_mem_reg[0][10]/NET0131 ,
		\u5_mem_reg[3][10]/NET0131 ,
		\u5_rp_reg[1]/NET0131 ,
		\u5_rp_reg[2]/NET0131 ,
		_w2811_
	);
	LUT4 #(
		.INIT('ha222)
	) name665 (
		_w2426_,
		_w2503_,
		_w2810_,
		_w2811_,
		_w2812_
	);
	LUT4 #(
		.INIT('h0b00)
	) name666 (
		_w2802_,
		_w2805_,
		_w2809_,
		_w2812_,
		_w2813_
	);
	LUT4 #(
		.INIT('h0b0f)
	) name667 (
		\u14_u2_en_out_l2_reg/P0001 ,
		\u14_u2_en_out_l_reg/NET0131 ,
		\u5_dout_reg[10]/P0001 ,
		\valid_s_reg/NET0131 ,
		_w2814_
	);
	LUT2 #(
		.INIT('h2)
	) name668 (
		\u13_occ0_r_reg[16]/NET0131 ,
		_w2814_,
		_w2815_
	);
	LUT2 #(
		.INIT('h4)
	) name669 (
		_w2813_,
		_w2815_,
		_w2816_
	);
	LUT4 #(
		.INIT('hc4cc)
	) name670 (
		\u5_mem_reg[2][23]/NET0131 ,
		\u5_rp_reg[0]/P0001 ,
		\u5_rp_reg[1]/NET0131 ,
		\u5_rp_reg[2]/NET0131 ,
		_w2817_
	);
	LUT3 #(
		.INIT('h02)
	) name671 (
		\u5_mem_reg[0][23]/NET0131 ,
		\u5_rp_reg[1]/NET0131 ,
		\u5_rp_reg[2]/NET0131 ,
		_w2818_
	);
	LUT4 #(
		.INIT('h3f5f)
	) name672 (
		\u5_mem_reg[1][23]/NET0131 ,
		\u5_mem_reg[3][23]/NET0131 ,
		\u5_rp_reg[1]/NET0131 ,
		\u5_rp_reg[2]/NET0131 ,
		_w2819_
	);
	LUT3 #(
		.INIT('h40)
	) name673 (
		_w2818_,
		_w2817_,
		_w2819_,
		_w2820_
	);
	LUT4 #(
		.INIT('hf35f)
	) name674 (
		\u5_mem_reg[1][7]/NET0131 ,
		\u5_mem_reg[2][7]/NET0131 ,
		\u5_rp_reg[1]/NET0131 ,
		\u5_rp_reg[2]/NET0131 ,
		_w2821_
	);
	LUT4 #(
		.INIT('h3ff5)
	) name675 (
		\u5_mem_reg[0][7]/NET0131 ,
		\u5_mem_reg[3][7]/NET0131 ,
		\u5_rp_reg[1]/NET0131 ,
		\u5_rp_reg[2]/NET0131 ,
		_w2822_
	);
	LUT4 #(
		.INIT('h8ccc)
	) name676 (
		\u5_rp_reg[0]/P0001 ,
		_w2427_,
		_w2821_,
		_w2822_,
		_w2823_
	);
	LUT4 #(
		.INIT('hf35f)
	) name677 (
		\u5_mem_reg[1][9]/NET0131 ,
		\u5_mem_reg[2][9]/NET0131 ,
		\u5_rp_reg[1]/NET0131 ,
		\u5_rp_reg[2]/NET0131 ,
		_w2824_
	);
	LUT4 #(
		.INIT('h3ff5)
	) name678 (
		\u5_mem_reg[0][9]/NET0131 ,
		\u5_mem_reg[3][9]/NET0131 ,
		\u5_rp_reg[1]/NET0131 ,
		\u5_rp_reg[2]/NET0131 ,
		_w2825_
	);
	LUT3 #(
		.INIT('h2a)
	) name679 (
		_w2806_,
		_w2824_,
		_w2825_,
		_w2826_
	);
	LUT4 #(
		.INIT('hf35f)
	) name680 (
		\u5_mem_reg[1][11]/NET0131 ,
		\u5_mem_reg[2][11]/NET0131 ,
		\u5_rp_reg[1]/NET0131 ,
		\u5_rp_reg[2]/NET0131 ,
		_w2827_
	);
	LUT4 #(
		.INIT('h3ff5)
	) name681 (
		\u5_mem_reg[0][11]/NET0131 ,
		\u5_mem_reg[3][11]/NET0131 ,
		\u5_rp_reg[1]/NET0131 ,
		\u5_rp_reg[2]/NET0131 ,
		_w2828_
	);
	LUT4 #(
		.INIT('ha222)
	) name682 (
		_w2426_,
		_w2503_,
		_w2827_,
		_w2828_,
		_w2829_
	);
	LUT4 #(
		.INIT('h0b00)
	) name683 (
		_w2820_,
		_w2823_,
		_w2826_,
		_w2829_,
		_w2830_
	);
	LUT4 #(
		.INIT('h0b0f)
	) name684 (
		\u14_u2_en_out_l2_reg/P0001 ,
		\u14_u2_en_out_l_reg/NET0131 ,
		\u5_dout_reg[11]/P0001 ,
		\valid_s_reg/NET0131 ,
		_w2831_
	);
	LUT2 #(
		.INIT('h2)
	) name685 (
		\u13_occ0_r_reg[16]/NET0131 ,
		_w2831_,
		_w2832_
	);
	LUT2 #(
		.INIT('h4)
	) name686 (
		_w2830_,
		_w2832_,
		_w2833_
	);
	LUT4 #(
		.INIT('hc4cc)
	) name687 (
		\u5_mem_reg[2][24]/NET0131 ,
		\u5_rp_reg[0]/P0001 ,
		\u5_rp_reg[1]/NET0131 ,
		\u5_rp_reg[2]/NET0131 ,
		_w2834_
	);
	LUT3 #(
		.INIT('h02)
	) name688 (
		\u5_mem_reg[0][24]/NET0131 ,
		\u5_rp_reg[1]/NET0131 ,
		\u5_rp_reg[2]/NET0131 ,
		_w2835_
	);
	LUT4 #(
		.INIT('h3f5f)
	) name689 (
		\u5_mem_reg[1][24]/NET0131 ,
		\u5_mem_reg[3][24]/NET0131 ,
		\u5_rp_reg[1]/NET0131 ,
		\u5_rp_reg[2]/NET0131 ,
		_w2836_
	);
	LUT3 #(
		.INIT('h40)
	) name690 (
		_w2835_,
		_w2834_,
		_w2836_,
		_w2837_
	);
	LUT4 #(
		.INIT('h8ccc)
	) name691 (
		\u5_rp_reg[0]/P0001 ,
		_w2427_,
		_w2807_,
		_w2808_,
		_w2838_
	);
	LUT3 #(
		.INIT('h70)
	) name692 (
		_w2810_,
		_w2811_,
		_w2806_,
		_w2839_
	);
	LUT4 #(
		.INIT('hf35f)
	) name693 (
		\u5_mem_reg[1][12]/NET0131 ,
		\u5_mem_reg[2][12]/NET0131 ,
		\u5_rp_reg[1]/NET0131 ,
		\u5_rp_reg[2]/NET0131 ,
		_w2840_
	);
	LUT4 #(
		.INIT('h3ff5)
	) name694 (
		\u5_mem_reg[0][12]/NET0131 ,
		\u5_mem_reg[3][12]/NET0131 ,
		\u5_rp_reg[1]/NET0131 ,
		\u5_rp_reg[2]/NET0131 ,
		_w2841_
	);
	LUT4 #(
		.INIT('ha222)
	) name695 (
		_w2426_,
		_w2503_,
		_w2840_,
		_w2841_,
		_w2842_
	);
	LUT4 #(
		.INIT('h0b00)
	) name696 (
		_w2837_,
		_w2838_,
		_w2839_,
		_w2842_,
		_w2843_
	);
	LUT4 #(
		.INIT('h0b0f)
	) name697 (
		\u14_u2_en_out_l2_reg/P0001 ,
		\u14_u2_en_out_l_reg/NET0131 ,
		\u5_dout_reg[12]/P0001 ,
		\valid_s_reg/NET0131 ,
		_w2844_
	);
	LUT2 #(
		.INIT('h2)
	) name698 (
		\u13_occ0_r_reg[16]/NET0131 ,
		_w2844_,
		_w2845_
	);
	LUT2 #(
		.INIT('h4)
	) name699 (
		_w2843_,
		_w2845_,
		_w2846_
	);
	LUT4 #(
		.INIT('hc4cc)
	) name700 (
		\u5_mem_reg[2][25]/NET0131 ,
		\u5_rp_reg[0]/P0001 ,
		\u5_rp_reg[1]/NET0131 ,
		\u5_rp_reg[2]/NET0131 ,
		_w2847_
	);
	LUT3 #(
		.INIT('h02)
	) name701 (
		\u5_mem_reg[0][25]/NET0131 ,
		\u5_rp_reg[1]/NET0131 ,
		\u5_rp_reg[2]/NET0131 ,
		_w2848_
	);
	LUT4 #(
		.INIT('h3f5f)
	) name702 (
		\u5_mem_reg[1][25]/NET0131 ,
		\u5_mem_reg[3][25]/NET0131 ,
		\u5_rp_reg[1]/NET0131 ,
		\u5_rp_reg[2]/NET0131 ,
		_w2849_
	);
	LUT3 #(
		.INIT('h40)
	) name703 (
		_w2848_,
		_w2847_,
		_w2849_,
		_w2850_
	);
	LUT4 #(
		.INIT('h8ccc)
	) name704 (
		\u5_rp_reg[0]/P0001 ,
		_w2427_,
		_w2824_,
		_w2825_,
		_w2851_
	);
	LUT3 #(
		.INIT('h2a)
	) name705 (
		_w2806_,
		_w2827_,
		_w2828_,
		_w2852_
	);
	LUT4 #(
		.INIT('hf35f)
	) name706 (
		\u5_mem_reg[1][13]/NET0131 ,
		\u5_mem_reg[2][13]/NET0131 ,
		\u5_rp_reg[1]/NET0131 ,
		\u5_rp_reg[2]/NET0131 ,
		_w2853_
	);
	LUT4 #(
		.INIT('h3ff5)
	) name707 (
		\u5_mem_reg[0][13]/NET0131 ,
		\u5_mem_reg[3][13]/NET0131 ,
		\u5_rp_reg[1]/NET0131 ,
		\u5_rp_reg[2]/NET0131 ,
		_w2854_
	);
	LUT4 #(
		.INIT('ha222)
	) name708 (
		_w2426_,
		_w2503_,
		_w2853_,
		_w2854_,
		_w2855_
	);
	LUT4 #(
		.INIT('h0b00)
	) name709 (
		_w2850_,
		_w2851_,
		_w2852_,
		_w2855_,
		_w2856_
	);
	LUT4 #(
		.INIT('h0b0f)
	) name710 (
		\u14_u2_en_out_l2_reg/P0001 ,
		\u14_u2_en_out_l_reg/NET0131 ,
		\u5_dout_reg[13]/P0001 ,
		\valid_s_reg/NET0131 ,
		_w2857_
	);
	LUT2 #(
		.INIT('h2)
	) name711 (
		\u13_occ0_r_reg[16]/NET0131 ,
		_w2857_,
		_w2858_
	);
	LUT2 #(
		.INIT('h4)
	) name712 (
		_w2856_,
		_w2858_,
		_w2859_
	);
	LUT4 #(
		.INIT('hc4cc)
	) name713 (
		\u5_mem_reg[2][26]/NET0131 ,
		\u5_rp_reg[0]/P0001 ,
		\u5_rp_reg[1]/NET0131 ,
		\u5_rp_reg[2]/NET0131 ,
		_w2860_
	);
	LUT3 #(
		.INIT('h02)
	) name714 (
		\u5_mem_reg[0][26]/NET0131 ,
		\u5_rp_reg[1]/NET0131 ,
		\u5_rp_reg[2]/NET0131 ,
		_w2861_
	);
	LUT4 #(
		.INIT('h3f5f)
	) name715 (
		\u5_mem_reg[1][26]/NET0131 ,
		\u5_mem_reg[3][26]/NET0131 ,
		\u5_rp_reg[1]/NET0131 ,
		\u5_rp_reg[2]/NET0131 ,
		_w2862_
	);
	LUT3 #(
		.INIT('h40)
	) name716 (
		_w2861_,
		_w2860_,
		_w2862_,
		_w2863_
	);
	LUT4 #(
		.INIT('h8ccc)
	) name717 (
		\u5_rp_reg[0]/P0001 ,
		_w2427_,
		_w2810_,
		_w2811_,
		_w2864_
	);
	LUT3 #(
		.INIT('h2a)
	) name718 (
		_w2806_,
		_w2840_,
		_w2841_,
		_w2865_
	);
	LUT4 #(
		.INIT('h35ff)
	) name719 (
		\u5_mem_reg[2][14]/NET0131 ,
		\u5_mem_reg[3][14]/NET0131 ,
		\u5_rp_reg[1]/NET0131 ,
		\u5_rp_reg[2]/NET0131 ,
		_w2866_
	);
	LUT4 #(
		.INIT('hff35)
	) name720 (
		\u5_mem_reg[0][14]/NET0131 ,
		\u5_mem_reg[1][14]/NET0131 ,
		\u5_rp_reg[1]/NET0131 ,
		\u5_rp_reg[2]/NET0131 ,
		_w2867_
	);
	LUT4 #(
		.INIT('ha222)
	) name721 (
		_w2426_,
		_w2503_,
		_w2866_,
		_w2867_,
		_w2868_
	);
	LUT4 #(
		.INIT('h0b00)
	) name722 (
		_w2863_,
		_w2864_,
		_w2865_,
		_w2868_,
		_w2869_
	);
	LUT4 #(
		.INIT('h0b0f)
	) name723 (
		\u14_u2_en_out_l2_reg/P0001 ,
		\u14_u2_en_out_l_reg/NET0131 ,
		\u5_dout_reg[14]/P0001 ,
		\valid_s_reg/NET0131 ,
		_w2870_
	);
	LUT2 #(
		.INIT('h2)
	) name724 (
		\u13_occ0_r_reg[16]/NET0131 ,
		_w2870_,
		_w2871_
	);
	LUT2 #(
		.INIT('h4)
	) name725 (
		_w2869_,
		_w2871_,
		_w2872_
	);
	LUT4 #(
		.INIT('hc4cc)
	) name726 (
		\u5_mem_reg[2][27]/NET0131 ,
		\u5_rp_reg[0]/P0001 ,
		\u5_rp_reg[1]/NET0131 ,
		\u5_rp_reg[2]/NET0131 ,
		_w2873_
	);
	LUT3 #(
		.INIT('h02)
	) name727 (
		\u5_mem_reg[0][27]/NET0131 ,
		\u5_rp_reg[1]/NET0131 ,
		\u5_rp_reg[2]/NET0131 ,
		_w2874_
	);
	LUT4 #(
		.INIT('h3f5f)
	) name728 (
		\u5_mem_reg[1][27]/NET0131 ,
		\u5_mem_reg[3][27]/NET0131 ,
		\u5_rp_reg[1]/NET0131 ,
		\u5_rp_reg[2]/NET0131 ,
		_w2875_
	);
	LUT3 #(
		.INIT('h40)
	) name729 (
		_w2874_,
		_w2873_,
		_w2875_,
		_w2876_
	);
	LUT4 #(
		.INIT('h8ccc)
	) name730 (
		\u5_rp_reg[0]/P0001 ,
		_w2427_,
		_w2827_,
		_w2828_,
		_w2877_
	);
	LUT3 #(
		.INIT('h2a)
	) name731 (
		_w2806_,
		_w2853_,
		_w2854_,
		_w2878_
	);
	LUT4 #(
		.INIT('h3f5f)
	) name732 (
		\u5_mem_reg[1][15]/NET0131 ,
		\u5_mem_reg[3][15]/NET0131 ,
		\u5_rp_reg[1]/NET0131 ,
		\u5_rp_reg[2]/NET0131 ,
		_w2879_
	);
	LUT4 #(
		.INIT('hf3f5)
	) name733 (
		\u5_mem_reg[0][15]/NET0131 ,
		\u5_mem_reg[2][15]/NET0131 ,
		\u5_rp_reg[1]/NET0131 ,
		\u5_rp_reg[2]/NET0131 ,
		_w2880_
	);
	LUT4 #(
		.INIT('ha222)
	) name734 (
		_w2426_,
		_w2503_,
		_w2879_,
		_w2880_,
		_w2881_
	);
	LUT4 #(
		.INIT('h0b00)
	) name735 (
		_w2876_,
		_w2877_,
		_w2878_,
		_w2881_,
		_w2882_
	);
	LUT4 #(
		.INIT('h0b0f)
	) name736 (
		\u14_u2_en_out_l2_reg/P0001 ,
		\u14_u2_en_out_l_reg/NET0131 ,
		\u5_dout_reg[15]/P0001 ,
		\valid_s_reg/NET0131 ,
		_w2883_
	);
	LUT2 #(
		.INIT('h2)
	) name737 (
		\u13_occ0_r_reg[16]/NET0131 ,
		_w2883_,
		_w2884_
	);
	LUT2 #(
		.INIT('h4)
	) name738 (
		_w2882_,
		_w2884_,
		_w2885_
	);
	LUT4 #(
		.INIT('hc4cc)
	) name739 (
		\u5_mem_reg[2][28]/NET0131 ,
		\u5_rp_reg[0]/P0001 ,
		\u5_rp_reg[1]/NET0131 ,
		\u5_rp_reg[2]/NET0131 ,
		_w2886_
	);
	LUT3 #(
		.INIT('h02)
	) name740 (
		\u5_mem_reg[0][28]/NET0131 ,
		\u5_rp_reg[1]/NET0131 ,
		\u5_rp_reg[2]/NET0131 ,
		_w2887_
	);
	LUT4 #(
		.INIT('h3f5f)
	) name741 (
		\u5_mem_reg[1][28]/NET0131 ,
		\u5_mem_reg[3][28]/NET0131 ,
		\u5_rp_reg[1]/NET0131 ,
		\u5_rp_reg[2]/NET0131 ,
		_w2888_
	);
	LUT3 #(
		.INIT('h40)
	) name742 (
		_w2887_,
		_w2886_,
		_w2888_,
		_w2889_
	);
	LUT4 #(
		.INIT('h8ccc)
	) name743 (
		\u5_rp_reg[0]/P0001 ,
		_w2427_,
		_w2840_,
		_w2841_,
		_w2890_
	);
	LUT3 #(
		.INIT('h2a)
	) name744 (
		_w2806_,
		_w2866_,
		_w2867_,
		_w2891_
	);
	LUT4 #(
		.INIT('h3f5f)
	) name745 (
		\u5_mem_reg[1][16]/NET0131 ,
		\u5_mem_reg[3][16]/NET0131 ,
		\u5_rp_reg[1]/NET0131 ,
		\u5_rp_reg[2]/NET0131 ,
		_w2892_
	);
	LUT4 #(
		.INIT('hf3f5)
	) name746 (
		\u5_mem_reg[0][16]/NET0131 ,
		\u5_mem_reg[2][16]/NET0131 ,
		\u5_rp_reg[1]/NET0131 ,
		\u5_rp_reg[2]/NET0131 ,
		_w2893_
	);
	LUT4 #(
		.INIT('ha222)
	) name747 (
		_w2426_,
		_w2503_,
		_w2892_,
		_w2893_,
		_w2894_
	);
	LUT4 #(
		.INIT('h0b00)
	) name748 (
		_w2889_,
		_w2890_,
		_w2891_,
		_w2894_,
		_w2895_
	);
	LUT4 #(
		.INIT('h0b0f)
	) name749 (
		\u14_u2_en_out_l2_reg/P0001 ,
		\u14_u2_en_out_l_reg/NET0131 ,
		\u5_dout_reg[16]/P0001 ,
		\valid_s_reg/NET0131 ,
		_w2896_
	);
	LUT2 #(
		.INIT('h2)
	) name750 (
		\u13_occ0_r_reg[16]/NET0131 ,
		_w2896_,
		_w2897_
	);
	LUT2 #(
		.INIT('h4)
	) name751 (
		_w2895_,
		_w2897_,
		_w2898_
	);
	LUT4 #(
		.INIT('hc4cc)
	) name752 (
		\u5_mem_reg[2][29]/NET0131 ,
		\u5_rp_reg[0]/P0001 ,
		\u5_rp_reg[1]/NET0131 ,
		\u5_rp_reg[2]/NET0131 ,
		_w2899_
	);
	LUT3 #(
		.INIT('h02)
	) name753 (
		\u5_mem_reg[0][29]/NET0131 ,
		\u5_rp_reg[1]/NET0131 ,
		\u5_rp_reg[2]/NET0131 ,
		_w2900_
	);
	LUT4 #(
		.INIT('h3f5f)
	) name754 (
		\u5_mem_reg[1][29]/NET0131 ,
		\u5_mem_reg[3][29]/NET0131 ,
		\u5_rp_reg[1]/NET0131 ,
		\u5_rp_reg[2]/NET0131 ,
		_w2901_
	);
	LUT3 #(
		.INIT('h40)
	) name755 (
		_w2900_,
		_w2899_,
		_w2901_,
		_w2902_
	);
	LUT4 #(
		.INIT('h8ccc)
	) name756 (
		\u5_rp_reg[0]/P0001 ,
		_w2427_,
		_w2853_,
		_w2854_,
		_w2903_
	);
	LUT3 #(
		.INIT('h2a)
	) name757 (
		_w2806_,
		_w2879_,
		_w2880_,
		_w2904_
	);
	LUT4 #(
		.INIT('h35ff)
	) name758 (
		\u5_mem_reg[2][17]/NET0131 ,
		\u5_mem_reg[3][17]/NET0131 ,
		\u5_rp_reg[1]/NET0131 ,
		\u5_rp_reg[2]/NET0131 ,
		_w2905_
	);
	LUT4 #(
		.INIT('hff35)
	) name759 (
		\u5_mem_reg[0][17]/NET0131 ,
		\u5_mem_reg[1][17]/NET0131 ,
		\u5_rp_reg[1]/NET0131 ,
		\u5_rp_reg[2]/NET0131 ,
		_w2906_
	);
	LUT4 #(
		.INIT('ha222)
	) name760 (
		_w2426_,
		_w2503_,
		_w2905_,
		_w2906_,
		_w2907_
	);
	LUT4 #(
		.INIT('h0b00)
	) name761 (
		_w2902_,
		_w2903_,
		_w2904_,
		_w2907_,
		_w2908_
	);
	LUT4 #(
		.INIT('h0b0f)
	) name762 (
		\u14_u2_en_out_l2_reg/P0001 ,
		\u14_u2_en_out_l_reg/NET0131 ,
		\u5_dout_reg[17]/P0001 ,
		\valid_s_reg/NET0131 ,
		_w2909_
	);
	LUT2 #(
		.INIT('h2)
	) name763 (
		\u13_occ0_r_reg[16]/NET0131 ,
		_w2909_,
		_w2910_
	);
	LUT2 #(
		.INIT('h4)
	) name764 (
		_w2908_,
		_w2910_,
		_w2911_
	);
	LUT4 #(
		.INIT('hc4cc)
	) name765 (
		\u5_mem_reg[2][30]/NET0131 ,
		\u5_rp_reg[0]/P0001 ,
		\u5_rp_reg[1]/NET0131 ,
		\u5_rp_reg[2]/NET0131 ,
		_w2912_
	);
	LUT3 #(
		.INIT('h02)
	) name766 (
		\u5_mem_reg[0][30]/NET0131 ,
		\u5_rp_reg[1]/NET0131 ,
		\u5_rp_reg[2]/NET0131 ,
		_w2913_
	);
	LUT4 #(
		.INIT('h3f5f)
	) name767 (
		\u5_mem_reg[1][30]/NET0131 ,
		\u5_mem_reg[3][30]/NET0131 ,
		\u5_rp_reg[1]/NET0131 ,
		\u5_rp_reg[2]/NET0131 ,
		_w2914_
	);
	LUT3 #(
		.INIT('h40)
	) name768 (
		_w2913_,
		_w2912_,
		_w2914_,
		_w2915_
	);
	LUT4 #(
		.INIT('h8ccc)
	) name769 (
		\u5_rp_reg[0]/P0001 ,
		_w2427_,
		_w2866_,
		_w2867_,
		_w2916_
	);
	LUT3 #(
		.INIT('h2a)
	) name770 (
		_w2806_,
		_w2892_,
		_w2893_,
		_w2917_
	);
	LUT4 #(
		.INIT('hf35f)
	) name771 (
		\u5_mem_reg[1][18]/NET0131 ,
		\u5_mem_reg[2][18]/NET0131 ,
		\u5_rp_reg[1]/NET0131 ,
		\u5_rp_reg[2]/NET0131 ,
		_w2918_
	);
	LUT4 #(
		.INIT('h3ff5)
	) name772 (
		\u5_mem_reg[0][18]/NET0131 ,
		\u5_mem_reg[3][18]/NET0131 ,
		\u5_rp_reg[1]/NET0131 ,
		\u5_rp_reg[2]/NET0131 ,
		_w2919_
	);
	LUT4 #(
		.INIT('ha222)
	) name773 (
		_w2426_,
		_w2503_,
		_w2918_,
		_w2919_,
		_w2920_
	);
	LUT4 #(
		.INIT('h0b00)
	) name774 (
		_w2915_,
		_w2916_,
		_w2917_,
		_w2920_,
		_w2921_
	);
	LUT4 #(
		.INIT('h0b0f)
	) name775 (
		\u14_u2_en_out_l2_reg/P0001 ,
		\u14_u2_en_out_l_reg/NET0131 ,
		\u5_dout_reg[18]/P0001 ,
		\valid_s_reg/NET0131 ,
		_w2922_
	);
	LUT2 #(
		.INIT('h2)
	) name776 (
		\u13_occ0_r_reg[16]/NET0131 ,
		_w2922_,
		_w2923_
	);
	LUT2 #(
		.INIT('h4)
	) name777 (
		_w2921_,
		_w2923_,
		_w2924_
	);
	LUT4 #(
		.INIT('hc4cc)
	) name778 (
		\u5_mem_reg[2][31]/NET0131 ,
		\u5_rp_reg[0]/P0001 ,
		\u5_rp_reg[1]/NET0131 ,
		\u5_rp_reg[2]/NET0131 ,
		_w2925_
	);
	LUT3 #(
		.INIT('h02)
	) name779 (
		\u5_mem_reg[0][31]/NET0131 ,
		\u5_rp_reg[1]/NET0131 ,
		\u5_rp_reg[2]/NET0131 ,
		_w2926_
	);
	LUT4 #(
		.INIT('h3f5f)
	) name780 (
		\u5_mem_reg[1][31]/NET0131 ,
		\u5_mem_reg[3][31]/NET0131 ,
		\u5_rp_reg[1]/NET0131 ,
		\u5_rp_reg[2]/NET0131 ,
		_w2927_
	);
	LUT3 #(
		.INIT('h40)
	) name781 (
		_w2926_,
		_w2925_,
		_w2927_,
		_w2928_
	);
	LUT4 #(
		.INIT('h8ccc)
	) name782 (
		\u5_rp_reg[0]/P0001 ,
		_w2427_,
		_w2879_,
		_w2880_,
		_w2929_
	);
	LUT3 #(
		.INIT('h2a)
	) name783 (
		_w2806_,
		_w2905_,
		_w2906_,
		_w2930_
	);
	LUT4 #(
		.INIT('h35ff)
	) name784 (
		\u5_mem_reg[2][19]/NET0131 ,
		\u5_mem_reg[3][19]/NET0131 ,
		\u5_rp_reg[1]/NET0131 ,
		\u5_rp_reg[2]/NET0131 ,
		_w2931_
	);
	LUT4 #(
		.INIT('hff35)
	) name785 (
		\u5_mem_reg[0][19]/NET0131 ,
		\u5_mem_reg[1][19]/NET0131 ,
		\u5_rp_reg[1]/NET0131 ,
		\u5_rp_reg[2]/NET0131 ,
		_w2932_
	);
	LUT4 #(
		.INIT('ha222)
	) name786 (
		_w2426_,
		_w2503_,
		_w2931_,
		_w2932_,
		_w2933_
	);
	LUT4 #(
		.INIT('h0b00)
	) name787 (
		_w2928_,
		_w2929_,
		_w2930_,
		_w2933_,
		_w2934_
	);
	LUT4 #(
		.INIT('h0b0f)
	) name788 (
		\u14_u2_en_out_l2_reg/P0001 ,
		\u14_u2_en_out_l_reg/NET0131 ,
		\u5_dout_reg[19]/P0001 ,
		\valid_s_reg/NET0131 ,
		_w2935_
	);
	LUT2 #(
		.INIT('h2)
	) name789 (
		\u13_occ0_r_reg[16]/NET0131 ,
		_w2935_,
		_w2936_
	);
	LUT2 #(
		.INIT('h4)
	) name790 (
		_w2934_,
		_w2936_,
		_w2937_
	);
	LUT4 #(
		.INIT('hff35)
	) name791 (
		\u5_mem_reg[0][2]/NET0131 ,
		\u5_mem_reg[1][2]/NET0131 ,
		\u5_rp_reg[1]/NET0131 ,
		\u5_rp_reg[2]/NET0131 ,
		_w2938_
	);
	LUT4 #(
		.INIT('h35ff)
	) name792 (
		\u5_mem_reg[2][2]/NET0131 ,
		\u5_mem_reg[3][2]/NET0131 ,
		\u5_rp_reg[1]/NET0131 ,
		\u5_rp_reg[2]/NET0131 ,
		_w2939_
	);
	LUT3 #(
		.INIT('h2a)
	) name793 (
		_w2503_,
		_w2938_,
		_w2939_,
		_w2940_
	);
	LUT4 #(
		.INIT('h80aa)
	) name794 (
		_w2426_,
		_w2501_,
		_w2502_,
		_w2806_,
		_w2941_
	);
	LUT4 #(
		.INIT('h0b0f)
	) name795 (
		\u14_u2_en_out_l2_reg/P0001 ,
		\u14_u2_en_out_l_reg/NET0131 ,
		\u5_dout_reg[2]/P0001 ,
		\valid_s_reg/NET0131 ,
		_w2942_
	);
	LUT2 #(
		.INIT('h2)
	) name796 (
		\u13_occ0_r_reg[16]/NET0131 ,
		_w2942_,
		_w2943_
	);
	LUT3 #(
		.INIT('hb0)
	) name797 (
		_w2940_,
		_w2941_,
		_w2943_,
		_w2944_
	);
	LUT4 #(
		.INIT('h35ff)
	) name798 (
		\u5_mem_reg[2][3]/NET0131 ,
		\u5_mem_reg[3][3]/NET0131 ,
		\u5_rp_reg[1]/NET0131 ,
		\u5_rp_reg[2]/NET0131 ,
		_w2945_
	);
	LUT4 #(
		.INIT('hff35)
	) name799 (
		\u5_mem_reg[0][3]/NET0131 ,
		\u5_mem_reg[1][3]/NET0131 ,
		\u5_rp_reg[1]/NET0131 ,
		\u5_rp_reg[2]/NET0131 ,
		_w2946_
	);
	LUT3 #(
		.INIT('h2a)
	) name800 (
		_w2503_,
		_w2945_,
		_w2946_,
		_w2947_
	);
	LUT4 #(
		.INIT('h80aa)
	) name801 (
		_w2426_,
		_w2508_,
		_w2509_,
		_w2806_,
		_w2948_
	);
	LUT4 #(
		.INIT('h0b0f)
	) name802 (
		\u14_u2_en_out_l2_reg/P0001 ,
		\u14_u2_en_out_l_reg/NET0131 ,
		\u5_dout_reg[3]/P0001 ,
		\valid_s_reg/NET0131 ,
		_w2949_
	);
	LUT2 #(
		.INIT('h2)
	) name803 (
		\u13_occ0_r_reg[16]/NET0131 ,
		_w2949_,
		_w2950_
	);
	LUT3 #(
		.INIT('hb0)
	) name804 (
		_w2947_,
		_w2948_,
		_w2950_,
		_w2951_
	);
	LUT3 #(
		.INIT('h80)
	) name805 (
		\u5_rp_reg[0]/P0001 ,
		_w2892_,
		_w2893_,
		_w2952_
	);
	LUT4 #(
		.INIT('h8ccc)
	) name806 (
		\u5_rp_reg[0]/P0001 ,
		_w2427_,
		_w2501_,
		_w2502_,
		_w2953_
	);
	LUT3 #(
		.INIT('h2a)
	) name807 (
		_w2806_,
		_w2938_,
		_w2939_,
		_w2954_
	);
	LUT4 #(
		.INIT('h3f5f)
	) name808 (
		\u5_mem_reg[1][4]/NET0131 ,
		\u5_mem_reg[3][4]/NET0131 ,
		\u5_rp_reg[1]/NET0131 ,
		\u5_rp_reg[2]/NET0131 ,
		_w2955_
	);
	LUT4 #(
		.INIT('hf3f5)
	) name809 (
		\u5_mem_reg[0][4]/NET0131 ,
		\u5_mem_reg[2][4]/NET0131 ,
		\u5_rp_reg[1]/NET0131 ,
		\u5_rp_reg[2]/NET0131 ,
		_w2956_
	);
	LUT4 #(
		.INIT('ha222)
	) name810 (
		_w2426_,
		_w2503_,
		_w2955_,
		_w2956_,
		_w2957_
	);
	LUT4 #(
		.INIT('h0b00)
	) name811 (
		_w2952_,
		_w2953_,
		_w2954_,
		_w2957_,
		_w2958_
	);
	LUT4 #(
		.INIT('h0b0f)
	) name812 (
		\u14_u2_en_out_l2_reg/P0001 ,
		\u14_u2_en_out_l_reg/NET0131 ,
		\u5_dout_reg[4]/P0001 ,
		\valid_s_reg/NET0131 ,
		_w2959_
	);
	LUT2 #(
		.INIT('h2)
	) name813 (
		\u13_occ0_r_reg[16]/NET0131 ,
		_w2959_,
		_w2960_
	);
	LUT2 #(
		.INIT('h4)
	) name814 (
		_w2958_,
		_w2960_,
		_w2961_
	);
	LUT3 #(
		.INIT('h80)
	) name815 (
		\u5_rp_reg[0]/P0001 ,
		_w2905_,
		_w2906_,
		_w2962_
	);
	LUT4 #(
		.INIT('h8ccc)
	) name816 (
		\u5_rp_reg[0]/P0001 ,
		_w2427_,
		_w2508_,
		_w2509_,
		_w2963_
	);
	LUT3 #(
		.INIT('h2a)
	) name817 (
		_w2806_,
		_w2945_,
		_w2946_,
		_w2964_
	);
	LUT4 #(
		.INIT('hf35f)
	) name818 (
		\u5_mem_reg[1][5]/NET0131 ,
		\u5_mem_reg[2][5]/NET0131 ,
		\u5_rp_reg[1]/NET0131 ,
		\u5_rp_reg[2]/NET0131 ,
		_w2965_
	);
	LUT4 #(
		.INIT('h3ff5)
	) name819 (
		\u5_mem_reg[0][5]/NET0131 ,
		\u5_mem_reg[3][5]/NET0131 ,
		\u5_rp_reg[1]/NET0131 ,
		\u5_rp_reg[2]/NET0131 ,
		_w2966_
	);
	LUT4 #(
		.INIT('ha222)
	) name820 (
		_w2426_,
		_w2503_,
		_w2965_,
		_w2966_,
		_w2967_
	);
	LUT4 #(
		.INIT('h0b00)
	) name821 (
		_w2962_,
		_w2963_,
		_w2964_,
		_w2967_,
		_w2968_
	);
	LUT4 #(
		.INIT('h0b0f)
	) name822 (
		\u14_u2_en_out_l2_reg/P0001 ,
		\u14_u2_en_out_l_reg/NET0131 ,
		\u5_dout_reg[5]/P0001 ,
		\valid_s_reg/NET0131 ,
		_w2969_
	);
	LUT2 #(
		.INIT('h2)
	) name823 (
		\u13_occ0_r_reg[16]/NET0131 ,
		_w2969_,
		_w2970_
	);
	LUT2 #(
		.INIT('h4)
	) name824 (
		_w2968_,
		_w2970_,
		_w2971_
	);
	LUT3 #(
		.INIT('h80)
	) name825 (
		\u5_rp_reg[0]/P0001 ,
		_w2918_,
		_w2919_,
		_w2972_
	);
	LUT4 #(
		.INIT('h8ccc)
	) name826 (
		\u5_rp_reg[0]/P0001 ,
		_w2427_,
		_w2938_,
		_w2939_,
		_w2973_
	);
	LUT3 #(
		.INIT('h2a)
	) name827 (
		_w2806_,
		_w2955_,
		_w2956_,
		_w2974_
	);
	LUT4 #(
		.INIT('ha222)
	) name828 (
		_w2426_,
		_w2503_,
		_w2803_,
		_w2804_,
		_w2975_
	);
	LUT4 #(
		.INIT('h0b00)
	) name829 (
		_w2972_,
		_w2973_,
		_w2974_,
		_w2975_,
		_w2976_
	);
	LUT4 #(
		.INIT('h0b0f)
	) name830 (
		\u14_u2_en_out_l2_reg/P0001 ,
		\u14_u2_en_out_l_reg/NET0131 ,
		\u5_dout_reg[6]/P0001 ,
		\valid_s_reg/NET0131 ,
		_w2977_
	);
	LUT2 #(
		.INIT('h2)
	) name831 (
		\u13_occ0_r_reg[16]/NET0131 ,
		_w2977_,
		_w2978_
	);
	LUT2 #(
		.INIT('h4)
	) name832 (
		_w2976_,
		_w2978_,
		_w2979_
	);
	LUT3 #(
		.INIT('h80)
	) name833 (
		\u5_rp_reg[0]/P0001 ,
		_w2931_,
		_w2932_,
		_w2980_
	);
	LUT4 #(
		.INIT('h8ccc)
	) name834 (
		\u5_rp_reg[0]/P0001 ,
		_w2427_,
		_w2945_,
		_w2946_,
		_w2981_
	);
	LUT3 #(
		.INIT('h2a)
	) name835 (
		_w2806_,
		_w2965_,
		_w2966_,
		_w2982_
	);
	LUT4 #(
		.INIT('ha222)
	) name836 (
		_w2426_,
		_w2503_,
		_w2821_,
		_w2822_,
		_w2983_
	);
	LUT4 #(
		.INIT('h0b00)
	) name837 (
		_w2980_,
		_w2981_,
		_w2982_,
		_w2983_,
		_w2984_
	);
	LUT4 #(
		.INIT('h0b0f)
	) name838 (
		\u14_u2_en_out_l2_reg/P0001 ,
		\u14_u2_en_out_l_reg/NET0131 ,
		\u5_dout_reg[7]/P0001 ,
		\valid_s_reg/NET0131 ,
		_w2985_
	);
	LUT2 #(
		.INIT('h2)
	) name839 (
		\u13_occ0_r_reg[16]/NET0131 ,
		_w2985_,
		_w2986_
	);
	LUT2 #(
		.INIT('h4)
	) name840 (
		_w2984_,
		_w2986_,
		_w2987_
	);
	LUT4 #(
		.INIT('hc4cc)
	) name841 (
		\u5_mem_reg[2][20]/NET0131 ,
		\u5_rp_reg[0]/P0001 ,
		\u5_rp_reg[1]/NET0131 ,
		\u5_rp_reg[2]/NET0131 ,
		_w2988_
	);
	LUT3 #(
		.INIT('h02)
	) name842 (
		\u5_mem_reg[0][20]/NET0131 ,
		\u5_rp_reg[1]/NET0131 ,
		\u5_rp_reg[2]/NET0131 ,
		_w2989_
	);
	LUT4 #(
		.INIT('h3f5f)
	) name843 (
		\u5_mem_reg[1][20]/NET0131 ,
		\u5_mem_reg[3][20]/NET0131 ,
		\u5_rp_reg[1]/NET0131 ,
		\u5_rp_reg[2]/NET0131 ,
		_w2990_
	);
	LUT3 #(
		.INIT('h40)
	) name844 (
		_w2989_,
		_w2988_,
		_w2990_,
		_w2991_
	);
	LUT4 #(
		.INIT('h8ccc)
	) name845 (
		\u5_rp_reg[0]/P0001 ,
		_w2427_,
		_w2955_,
		_w2956_,
		_w2992_
	);
	LUT3 #(
		.INIT('h70)
	) name846 (
		_w2803_,
		_w2804_,
		_w2806_,
		_w2993_
	);
	LUT4 #(
		.INIT('ha222)
	) name847 (
		_w2426_,
		_w2503_,
		_w2807_,
		_w2808_,
		_w2994_
	);
	LUT4 #(
		.INIT('h0b00)
	) name848 (
		_w2991_,
		_w2992_,
		_w2993_,
		_w2994_,
		_w2995_
	);
	LUT4 #(
		.INIT('h0b0f)
	) name849 (
		\u14_u2_en_out_l2_reg/P0001 ,
		\u14_u2_en_out_l_reg/NET0131 ,
		\u5_dout_reg[8]/P0001 ,
		\valid_s_reg/NET0131 ,
		_w2996_
	);
	LUT2 #(
		.INIT('h2)
	) name850 (
		\u13_occ0_r_reg[16]/NET0131 ,
		_w2996_,
		_w2997_
	);
	LUT2 #(
		.INIT('h4)
	) name851 (
		_w2995_,
		_w2997_,
		_w2998_
	);
	LUT4 #(
		.INIT('hc4cc)
	) name852 (
		\u5_mem_reg[2][21]/NET0131 ,
		\u5_rp_reg[0]/P0001 ,
		\u5_rp_reg[1]/NET0131 ,
		\u5_rp_reg[2]/NET0131 ,
		_w2999_
	);
	LUT3 #(
		.INIT('h02)
	) name853 (
		\u5_mem_reg[0][21]/NET0131 ,
		\u5_rp_reg[1]/NET0131 ,
		\u5_rp_reg[2]/NET0131 ,
		_w3000_
	);
	LUT4 #(
		.INIT('h3f5f)
	) name854 (
		\u5_mem_reg[1][21]/NET0131 ,
		\u5_mem_reg[3][21]/NET0131 ,
		\u5_rp_reg[1]/NET0131 ,
		\u5_rp_reg[2]/NET0131 ,
		_w3001_
	);
	LUT3 #(
		.INIT('h40)
	) name855 (
		_w3000_,
		_w2999_,
		_w3001_,
		_w3002_
	);
	LUT4 #(
		.INIT('h8ccc)
	) name856 (
		\u5_rp_reg[0]/P0001 ,
		_w2427_,
		_w2965_,
		_w2966_,
		_w3003_
	);
	LUT3 #(
		.INIT('h2a)
	) name857 (
		_w2806_,
		_w2821_,
		_w2822_,
		_w3004_
	);
	LUT4 #(
		.INIT('ha222)
	) name858 (
		_w2426_,
		_w2503_,
		_w2824_,
		_w2825_,
		_w3005_
	);
	LUT4 #(
		.INIT('h0b00)
	) name859 (
		_w3002_,
		_w3003_,
		_w3004_,
		_w3005_,
		_w3006_
	);
	LUT4 #(
		.INIT('h0b0f)
	) name860 (
		\u14_u2_en_out_l2_reg/P0001 ,
		\u14_u2_en_out_l_reg/NET0131 ,
		\u5_dout_reg[9]/P0001 ,
		\valid_s_reg/NET0131 ,
		_w3007_
	);
	LUT2 #(
		.INIT('h2)
	) name861 (
		\u13_occ0_r_reg[16]/NET0131 ,
		_w3007_,
		_w3008_
	);
	LUT2 #(
		.INIT('h4)
	) name862 (
		_w3006_,
		_w3008_,
		_w3009_
	);
	LUT4 #(
		.INIT('hc4cc)
	) name863 (
		\u6_mem_reg[2][22]/NET0131 ,
		\u6_rp_reg[0]/P0001 ,
		\u6_rp_reg[1]/NET0131 ,
		\u6_rp_reg[2]/NET0131 ,
		_w3010_
	);
	LUT3 #(
		.INIT('h02)
	) name864 (
		\u6_mem_reg[0][22]/NET0131 ,
		\u6_rp_reg[1]/NET0131 ,
		\u6_rp_reg[2]/NET0131 ,
		_w3011_
	);
	LUT4 #(
		.INIT('h3f5f)
	) name865 (
		\u6_mem_reg[1][22]/NET0131 ,
		\u6_mem_reg[3][22]/NET0131 ,
		\u6_rp_reg[1]/NET0131 ,
		\u6_rp_reg[2]/NET0131 ,
		_w3012_
	);
	LUT3 #(
		.INIT('h40)
	) name866 (
		_w3011_,
		_w3010_,
		_w3012_,
		_w3013_
	);
	LUT4 #(
		.INIT('h35ff)
	) name867 (
		\u6_mem_reg[2][6]/NET0131 ,
		\u6_mem_reg[3][6]/NET0131 ,
		\u6_rp_reg[1]/NET0131 ,
		\u6_rp_reg[2]/NET0131 ,
		_w3014_
	);
	LUT4 #(
		.INIT('hff35)
	) name868 (
		\u6_mem_reg[0][6]/NET0131 ,
		\u6_mem_reg[1][6]/NET0131 ,
		\u6_rp_reg[1]/NET0131 ,
		\u6_rp_reg[2]/NET0131 ,
		_w3015_
	);
	LUT4 #(
		.INIT('h8ccc)
	) name869 (
		\u6_rp_reg[0]/P0001 ,
		_w2445_,
		_w3014_,
		_w3015_,
		_w3016_
	);
	LUT2 #(
		.INIT('h2)
	) name870 (
		\u13_occ0_r_reg[26]/NET0131 ,
		\u13_occ0_r_reg[27]/NET0131 ,
		_w3017_
	);
	LUT4 #(
		.INIT('h35ff)
	) name871 (
		\u6_mem_reg[2][8]/NET0131 ,
		\u6_mem_reg[3][8]/NET0131 ,
		\u6_rp_reg[1]/NET0131 ,
		\u6_rp_reg[2]/NET0131 ,
		_w3018_
	);
	LUT4 #(
		.INIT('hff35)
	) name872 (
		\u6_mem_reg[0][8]/NET0131 ,
		\u6_mem_reg[1][8]/NET0131 ,
		\u6_rp_reg[1]/NET0131 ,
		\u6_rp_reg[2]/NET0131 ,
		_w3019_
	);
	LUT3 #(
		.INIT('h2a)
	) name873 (
		_w3017_,
		_w3018_,
		_w3019_,
		_w3020_
	);
	LUT4 #(
		.INIT('h3f5f)
	) name874 (
		\u6_mem_reg[1][10]/NET0131 ,
		\u6_mem_reg[3][10]/NET0131 ,
		\u6_rp_reg[1]/NET0131 ,
		\u6_rp_reg[2]/NET0131 ,
		_w3021_
	);
	LUT4 #(
		.INIT('hf3f5)
	) name875 (
		\u6_mem_reg[0][10]/NET0131 ,
		\u6_mem_reg[2][10]/NET0131 ,
		\u6_rp_reg[1]/NET0131 ,
		\u6_rp_reg[2]/NET0131 ,
		_w3022_
	);
	LUT4 #(
		.INIT('ha222)
	) name876 (
		_w2444_,
		_w2516_,
		_w3021_,
		_w3022_,
		_w3023_
	);
	LUT4 #(
		.INIT('h0b00)
	) name877 (
		_w3013_,
		_w3016_,
		_w3020_,
		_w3023_,
		_w3024_
	);
	LUT4 #(
		.INIT('h0b0f)
	) name878 (
		\u14_u3_en_out_l2_reg/P0001 ,
		\u14_u3_en_out_l_reg/NET0131 ,
		\u6_dout_reg[10]/P0001 ,
		\valid_s_reg/NET0131 ,
		_w3025_
	);
	LUT2 #(
		.INIT('h2)
	) name879 (
		\u13_occ0_r_reg[24]/NET0131 ,
		_w3025_,
		_w3026_
	);
	LUT2 #(
		.INIT('h4)
	) name880 (
		_w3024_,
		_w3026_,
		_w3027_
	);
	LUT4 #(
		.INIT('hc4cc)
	) name881 (
		\u6_mem_reg[2][23]/NET0131 ,
		\u6_rp_reg[0]/P0001 ,
		\u6_rp_reg[1]/NET0131 ,
		\u6_rp_reg[2]/NET0131 ,
		_w3028_
	);
	LUT3 #(
		.INIT('h02)
	) name882 (
		\u6_mem_reg[0][23]/NET0131 ,
		\u6_rp_reg[1]/NET0131 ,
		\u6_rp_reg[2]/NET0131 ,
		_w3029_
	);
	LUT4 #(
		.INIT('h3f5f)
	) name883 (
		\u6_mem_reg[1][23]/NET0131 ,
		\u6_mem_reg[3][23]/NET0131 ,
		\u6_rp_reg[1]/NET0131 ,
		\u6_rp_reg[2]/NET0131 ,
		_w3030_
	);
	LUT3 #(
		.INIT('h40)
	) name884 (
		_w3029_,
		_w3028_,
		_w3030_,
		_w3031_
	);
	LUT4 #(
		.INIT('h35ff)
	) name885 (
		\u6_mem_reg[2][7]/NET0131 ,
		\u6_mem_reg[3][7]/NET0131 ,
		\u6_rp_reg[1]/NET0131 ,
		\u6_rp_reg[2]/NET0131 ,
		_w3032_
	);
	LUT4 #(
		.INIT('hff35)
	) name886 (
		\u6_mem_reg[0][7]/NET0131 ,
		\u6_mem_reg[1][7]/NET0131 ,
		\u6_rp_reg[1]/NET0131 ,
		\u6_rp_reg[2]/NET0131 ,
		_w3033_
	);
	LUT4 #(
		.INIT('h8ccc)
	) name887 (
		\u6_rp_reg[0]/P0001 ,
		_w2445_,
		_w3032_,
		_w3033_,
		_w3034_
	);
	LUT4 #(
		.INIT('h3f5f)
	) name888 (
		\u6_mem_reg[1][9]/NET0131 ,
		\u6_mem_reg[3][9]/NET0131 ,
		\u6_rp_reg[1]/NET0131 ,
		\u6_rp_reg[2]/NET0131 ,
		_w3035_
	);
	LUT4 #(
		.INIT('hf3f5)
	) name889 (
		\u6_mem_reg[0][9]/NET0131 ,
		\u6_mem_reg[2][9]/NET0131 ,
		\u6_rp_reg[1]/NET0131 ,
		\u6_rp_reg[2]/NET0131 ,
		_w3036_
	);
	LUT3 #(
		.INIT('h2a)
	) name890 (
		_w3017_,
		_w3035_,
		_w3036_,
		_w3037_
	);
	LUT4 #(
		.INIT('h35ff)
	) name891 (
		\u6_mem_reg[2][11]/NET0131 ,
		\u6_mem_reg[3][11]/NET0131 ,
		\u6_rp_reg[1]/NET0131 ,
		\u6_rp_reg[2]/NET0131 ,
		_w3038_
	);
	LUT4 #(
		.INIT('hff35)
	) name892 (
		\u6_mem_reg[0][11]/NET0131 ,
		\u6_mem_reg[1][11]/NET0131 ,
		\u6_rp_reg[1]/NET0131 ,
		\u6_rp_reg[2]/NET0131 ,
		_w3039_
	);
	LUT4 #(
		.INIT('ha222)
	) name893 (
		_w2444_,
		_w2516_,
		_w3038_,
		_w3039_,
		_w3040_
	);
	LUT4 #(
		.INIT('h0b00)
	) name894 (
		_w3031_,
		_w3034_,
		_w3037_,
		_w3040_,
		_w3041_
	);
	LUT4 #(
		.INIT('h0b0f)
	) name895 (
		\u14_u3_en_out_l2_reg/P0001 ,
		\u14_u3_en_out_l_reg/NET0131 ,
		\u6_dout_reg[11]/P0001 ,
		\valid_s_reg/NET0131 ,
		_w3042_
	);
	LUT2 #(
		.INIT('h2)
	) name896 (
		\u13_occ0_r_reg[24]/NET0131 ,
		_w3042_,
		_w3043_
	);
	LUT2 #(
		.INIT('h4)
	) name897 (
		_w3041_,
		_w3043_,
		_w3044_
	);
	LUT4 #(
		.INIT('hc4cc)
	) name898 (
		\u6_mem_reg[2][24]/NET0131 ,
		\u6_rp_reg[0]/P0001 ,
		\u6_rp_reg[1]/NET0131 ,
		\u6_rp_reg[2]/NET0131 ,
		_w3045_
	);
	LUT3 #(
		.INIT('h02)
	) name899 (
		\u6_mem_reg[0][24]/NET0131 ,
		\u6_rp_reg[1]/NET0131 ,
		\u6_rp_reg[2]/NET0131 ,
		_w3046_
	);
	LUT4 #(
		.INIT('h3f5f)
	) name900 (
		\u6_mem_reg[1][24]/NET0131 ,
		\u6_mem_reg[3][24]/NET0131 ,
		\u6_rp_reg[1]/NET0131 ,
		\u6_rp_reg[2]/NET0131 ,
		_w3047_
	);
	LUT3 #(
		.INIT('h40)
	) name901 (
		_w3046_,
		_w3045_,
		_w3047_,
		_w3048_
	);
	LUT4 #(
		.INIT('h8ccc)
	) name902 (
		\u6_rp_reg[0]/P0001 ,
		_w2445_,
		_w3018_,
		_w3019_,
		_w3049_
	);
	LUT3 #(
		.INIT('h70)
	) name903 (
		_w3021_,
		_w3022_,
		_w3017_,
		_w3050_
	);
	LUT4 #(
		.INIT('h3f5f)
	) name904 (
		\u6_mem_reg[1][12]/NET0131 ,
		\u6_mem_reg[3][12]/NET0131 ,
		\u6_rp_reg[1]/NET0131 ,
		\u6_rp_reg[2]/NET0131 ,
		_w3051_
	);
	LUT4 #(
		.INIT('hf3f5)
	) name905 (
		\u6_mem_reg[0][12]/NET0131 ,
		\u6_mem_reg[2][12]/NET0131 ,
		\u6_rp_reg[1]/NET0131 ,
		\u6_rp_reg[2]/NET0131 ,
		_w3052_
	);
	LUT4 #(
		.INIT('ha222)
	) name906 (
		_w2444_,
		_w2516_,
		_w3051_,
		_w3052_,
		_w3053_
	);
	LUT4 #(
		.INIT('h0b00)
	) name907 (
		_w3048_,
		_w3049_,
		_w3050_,
		_w3053_,
		_w3054_
	);
	LUT4 #(
		.INIT('h0b0f)
	) name908 (
		\u14_u3_en_out_l2_reg/P0001 ,
		\u14_u3_en_out_l_reg/NET0131 ,
		\u6_dout_reg[12]/P0001 ,
		\valid_s_reg/NET0131 ,
		_w3055_
	);
	LUT2 #(
		.INIT('h2)
	) name909 (
		\u13_occ0_r_reg[24]/NET0131 ,
		_w3055_,
		_w3056_
	);
	LUT2 #(
		.INIT('h4)
	) name910 (
		_w3054_,
		_w3056_,
		_w3057_
	);
	LUT4 #(
		.INIT('hc4cc)
	) name911 (
		\u6_mem_reg[2][25]/NET0131 ,
		\u6_rp_reg[0]/P0001 ,
		\u6_rp_reg[1]/NET0131 ,
		\u6_rp_reg[2]/NET0131 ,
		_w3058_
	);
	LUT3 #(
		.INIT('h02)
	) name912 (
		\u6_mem_reg[0][25]/NET0131 ,
		\u6_rp_reg[1]/NET0131 ,
		\u6_rp_reg[2]/NET0131 ,
		_w3059_
	);
	LUT4 #(
		.INIT('h3f5f)
	) name913 (
		\u6_mem_reg[1][25]/NET0131 ,
		\u6_mem_reg[3][25]/NET0131 ,
		\u6_rp_reg[1]/NET0131 ,
		\u6_rp_reg[2]/NET0131 ,
		_w3060_
	);
	LUT3 #(
		.INIT('h40)
	) name914 (
		_w3059_,
		_w3058_,
		_w3060_,
		_w3061_
	);
	LUT4 #(
		.INIT('h8ccc)
	) name915 (
		\u6_rp_reg[0]/P0001 ,
		_w2445_,
		_w3035_,
		_w3036_,
		_w3062_
	);
	LUT3 #(
		.INIT('h2a)
	) name916 (
		_w3017_,
		_w3038_,
		_w3039_,
		_w3063_
	);
	LUT4 #(
		.INIT('h35ff)
	) name917 (
		\u6_mem_reg[2][13]/NET0131 ,
		\u6_mem_reg[3][13]/NET0131 ,
		\u6_rp_reg[1]/NET0131 ,
		\u6_rp_reg[2]/NET0131 ,
		_w3064_
	);
	LUT4 #(
		.INIT('hff35)
	) name918 (
		\u6_mem_reg[0][13]/NET0131 ,
		\u6_mem_reg[1][13]/NET0131 ,
		\u6_rp_reg[1]/NET0131 ,
		\u6_rp_reg[2]/NET0131 ,
		_w3065_
	);
	LUT4 #(
		.INIT('ha222)
	) name919 (
		_w2444_,
		_w2516_,
		_w3064_,
		_w3065_,
		_w3066_
	);
	LUT4 #(
		.INIT('h0b00)
	) name920 (
		_w3061_,
		_w3062_,
		_w3063_,
		_w3066_,
		_w3067_
	);
	LUT4 #(
		.INIT('h0b0f)
	) name921 (
		\u14_u3_en_out_l2_reg/P0001 ,
		\u14_u3_en_out_l_reg/NET0131 ,
		\u6_dout_reg[13]/P0001 ,
		\valid_s_reg/NET0131 ,
		_w3068_
	);
	LUT2 #(
		.INIT('h2)
	) name922 (
		\u13_occ0_r_reg[24]/NET0131 ,
		_w3068_,
		_w3069_
	);
	LUT2 #(
		.INIT('h4)
	) name923 (
		_w3067_,
		_w3069_,
		_w3070_
	);
	LUT4 #(
		.INIT('hc4cc)
	) name924 (
		\u6_mem_reg[2][26]/NET0131 ,
		\u6_rp_reg[0]/P0001 ,
		\u6_rp_reg[1]/NET0131 ,
		\u6_rp_reg[2]/NET0131 ,
		_w3071_
	);
	LUT3 #(
		.INIT('h02)
	) name925 (
		\u6_mem_reg[0][26]/NET0131 ,
		\u6_rp_reg[1]/NET0131 ,
		\u6_rp_reg[2]/NET0131 ,
		_w3072_
	);
	LUT4 #(
		.INIT('h3f5f)
	) name926 (
		\u6_mem_reg[1][26]/NET0131 ,
		\u6_mem_reg[3][26]/NET0131 ,
		\u6_rp_reg[1]/NET0131 ,
		\u6_rp_reg[2]/NET0131 ,
		_w3073_
	);
	LUT3 #(
		.INIT('h40)
	) name927 (
		_w3072_,
		_w3071_,
		_w3073_,
		_w3074_
	);
	LUT4 #(
		.INIT('h8ccc)
	) name928 (
		\u6_rp_reg[0]/P0001 ,
		_w2445_,
		_w3021_,
		_w3022_,
		_w3075_
	);
	LUT3 #(
		.INIT('h2a)
	) name929 (
		_w3017_,
		_w3051_,
		_w3052_,
		_w3076_
	);
	LUT4 #(
		.INIT('hff35)
	) name930 (
		\u6_mem_reg[0][14]/NET0131 ,
		\u6_mem_reg[1][14]/NET0131 ,
		\u6_rp_reg[1]/NET0131 ,
		\u6_rp_reg[2]/NET0131 ,
		_w3077_
	);
	LUT4 #(
		.INIT('h35ff)
	) name931 (
		\u6_mem_reg[2][14]/NET0131 ,
		\u6_mem_reg[3][14]/NET0131 ,
		\u6_rp_reg[1]/NET0131 ,
		\u6_rp_reg[2]/NET0131 ,
		_w3078_
	);
	LUT4 #(
		.INIT('ha222)
	) name932 (
		_w2444_,
		_w2516_,
		_w3077_,
		_w3078_,
		_w3079_
	);
	LUT4 #(
		.INIT('h0b00)
	) name933 (
		_w3074_,
		_w3075_,
		_w3076_,
		_w3079_,
		_w3080_
	);
	LUT4 #(
		.INIT('h0b0f)
	) name934 (
		\u14_u3_en_out_l2_reg/P0001 ,
		\u14_u3_en_out_l_reg/NET0131 ,
		\u6_dout_reg[14]/P0001 ,
		\valid_s_reg/NET0131 ,
		_w3081_
	);
	LUT2 #(
		.INIT('h2)
	) name935 (
		\u13_occ0_r_reg[24]/NET0131 ,
		_w3081_,
		_w3082_
	);
	LUT2 #(
		.INIT('h4)
	) name936 (
		_w3080_,
		_w3082_,
		_w3083_
	);
	LUT4 #(
		.INIT('hc4cc)
	) name937 (
		\u6_mem_reg[2][27]/NET0131 ,
		\u6_rp_reg[0]/P0001 ,
		\u6_rp_reg[1]/NET0131 ,
		\u6_rp_reg[2]/NET0131 ,
		_w3084_
	);
	LUT3 #(
		.INIT('h02)
	) name938 (
		\u6_mem_reg[0][27]/NET0131 ,
		\u6_rp_reg[1]/NET0131 ,
		\u6_rp_reg[2]/NET0131 ,
		_w3085_
	);
	LUT4 #(
		.INIT('h3f5f)
	) name939 (
		\u6_mem_reg[1][27]/NET0131 ,
		\u6_mem_reg[3][27]/NET0131 ,
		\u6_rp_reg[1]/NET0131 ,
		\u6_rp_reg[2]/NET0131 ,
		_w3086_
	);
	LUT3 #(
		.INIT('h40)
	) name940 (
		_w3085_,
		_w3084_,
		_w3086_,
		_w3087_
	);
	LUT4 #(
		.INIT('h8ccc)
	) name941 (
		\u6_rp_reg[0]/P0001 ,
		_w2445_,
		_w3038_,
		_w3039_,
		_w3088_
	);
	LUT3 #(
		.INIT('h2a)
	) name942 (
		_w3017_,
		_w3064_,
		_w3065_,
		_w3089_
	);
	LUT4 #(
		.INIT('h35ff)
	) name943 (
		\u6_mem_reg[2][15]/NET0131 ,
		\u6_mem_reg[3][15]/NET0131 ,
		\u6_rp_reg[1]/NET0131 ,
		\u6_rp_reg[2]/NET0131 ,
		_w3090_
	);
	LUT4 #(
		.INIT('hff35)
	) name944 (
		\u6_mem_reg[0][15]/NET0131 ,
		\u6_mem_reg[1][15]/NET0131 ,
		\u6_rp_reg[1]/NET0131 ,
		\u6_rp_reg[2]/NET0131 ,
		_w3091_
	);
	LUT4 #(
		.INIT('ha222)
	) name945 (
		_w2444_,
		_w2516_,
		_w3090_,
		_w3091_,
		_w3092_
	);
	LUT4 #(
		.INIT('h0b00)
	) name946 (
		_w3087_,
		_w3088_,
		_w3089_,
		_w3092_,
		_w3093_
	);
	LUT4 #(
		.INIT('h0b0f)
	) name947 (
		\u14_u3_en_out_l2_reg/P0001 ,
		\u14_u3_en_out_l_reg/NET0131 ,
		\u6_dout_reg[15]/P0001 ,
		\valid_s_reg/NET0131 ,
		_w3094_
	);
	LUT2 #(
		.INIT('h2)
	) name948 (
		\u13_occ0_r_reg[24]/NET0131 ,
		_w3094_,
		_w3095_
	);
	LUT2 #(
		.INIT('h4)
	) name949 (
		_w3093_,
		_w3095_,
		_w3096_
	);
	LUT4 #(
		.INIT('hc4cc)
	) name950 (
		\u6_mem_reg[2][28]/NET0131 ,
		\u6_rp_reg[0]/P0001 ,
		\u6_rp_reg[1]/NET0131 ,
		\u6_rp_reg[2]/NET0131 ,
		_w3097_
	);
	LUT3 #(
		.INIT('h02)
	) name951 (
		\u6_mem_reg[0][28]/NET0131 ,
		\u6_rp_reg[1]/NET0131 ,
		\u6_rp_reg[2]/NET0131 ,
		_w3098_
	);
	LUT4 #(
		.INIT('h3f5f)
	) name952 (
		\u6_mem_reg[1][28]/NET0131 ,
		\u6_mem_reg[3][28]/NET0131 ,
		\u6_rp_reg[1]/NET0131 ,
		\u6_rp_reg[2]/NET0131 ,
		_w3099_
	);
	LUT3 #(
		.INIT('h40)
	) name953 (
		_w3098_,
		_w3097_,
		_w3099_,
		_w3100_
	);
	LUT4 #(
		.INIT('h8ccc)
	) name954 (
		\u6_rp_reg[0]/P0001 ,
		_w2445_,
		_w3051_,
		_w3052_,
		_w3101_
	);
	LUT3 #(
		.INIT('h2a)
	) name955 (
		_w3017_,
		_w3077_,
		_w3078_,
		_w3102_
	);
	LUT4 #(
		.INIT('hff35)
	) name956 (
		\u6_mem_reg[0][16]/NET0131 ,
		\u6_mem_reg[1][16]/NET0131 ,
		\u6_rp_reg[1]/NET0131 ,
		\u6_rp_reg[2]/NET0131 ,
		_w3103_
	);
	LUT4 #(
		.INIT('h35ff)
	) name957 (
		\u6_mem_reg[2][16]/NET0131 ,
		\u6_mem_reg[3][16]/NET0131 ,
		\u6_rp_reg[1]/NET0131 ,
		\u6_rp_reg[2]/NET0131 ,
		_w3104_
	);
	LUT4 #(
		.INIT('ha222)
	) name958 (
		_w2444_,
		_w2516_,
		_w3103_,
		_w3104_,
		_w3105_
	);
	LUT4 #(
		.INIT('h0b00)
	) name959 (
		_w3100_,
		_w3101_,
		_w3102_,
		_w3105_,
		_w3106_
	);
	LUT4 #(
		.INIT('h0b0f)
	) name960 (
		\u14_u3_en_out_l2_reg/P0001 ,
		\u14_u3_en_out_l_reg/NET0131 ,
		\u6_dout_reg[16]/P0001 ,
		\valid_s_reg/NET0131 ,
		_w3107_
	);
	LUT2 #(
		.INIT('h2)
	) name961 (
		\u13_occ0_r_reg[24]/NET0131 ,
		_w3107_,
		_w3108_
	);
	LUT2 #(
		.INIT('h4)
	) name962 (
		_w3106_,
		_w3108_,
		_w3109_
	);
	LUT4 #(
		.INIT('hc4cc)
	) name963 (
		\u6_mem_reg[2][29]/NET0131 ,
		\u6_rp_reg[0]/P0001 ,
		\u6_rp_reg[1]/NET0131 ,
		\u6_rp_reg[2]/NET0131 ,
		_w3110_
	);
	LUT3 #(
		.INIT('h02)
	) name964 (
		\u6_mem_reg[0][29]/NET0131 ,
		\u6_rp_reg[1]/NET0131 ,
		\u6_rp_reg[2]/NET0131 ,
		_w3111_
	);
	LUT4 #(
		.INIT('h3f5f)
	) name965 (
		\u6_mem_reg[1][29]/NET0131 ,
		\u6_mem_reg[3][29]/NET0131 ,
		\u6_rp_reg[1]/NET0131 ,
		\u6_rp_reg[2]/NET0131 ,
		_w3112_
	);
	LUT3 #(
		.INIT('h40)
	) name966 (
		_w3111_,
		_w3110_,
		_w3112_,
		_w3113_
	);
	LUT4 #(
		.INIT('h8ccc)
	) name967 (
		\u6_rp_reg[0]/P0001 ,
		_w2445_,
		_w3064_,
		_w3065_,
		_w3114_
	);
	LUT3 #(
		.INIT('h2a)
	) name968 (
		_w3017_,
		_w3090_,
		_w3091_,
		_w3115_
	);
	LUT4 #(
		.INIT('h3f5f)
	) name969 (
		\u6_mem_reg[1][17]/NET0131 ,
		\u6_mem_reg[3][17]/NET0131 ,
		\u6_rp_reg[1]/NET0131 ,
		\u6_rp_reg[2]/NET0131 ,
		_w3116_
	);
	LUT4 #(
		.INIT('hf3f5)
	) name970 (
		\u6_mem_reg[0][17]/NET0131 ,
		\u6_mem_reg[2][17]/NET0131 ,
		\u6_rp_reg[1]/NET0131 ,
		\u6_rp_reg[2]/NET0131 ,
		_w3117_
	);
	LUT4 #(
		.INIT('ha222)
	) name971 (
		_w2444_,
		_w2516_,
		_w3116_,
		_w3117_,
		_w3118_
	);
	LUT4 #(
		.INIT('h0b00)
	) name972 (
		_w3113_,
		_w3114_,
		_w3115_,
		_w3118_,
		_w3119_
	);
	LUT4 #(
		.INIT('h0b0f)
	) name973 (
		\u14_u3_en_out_l2_reg/P0001 ,
		\u14_u3_en_out_l_reg/NET0131 ,
		\u6_dout_reg[17]/P0001 ,
		\valid_s_reg/NET0131 ,
		_w3120_
	);
	LUT2 #(
		.INIT('h2)
	) name974 (
		\u13_occ0_r_reg[24]/NET0131 ,
		_w3120_,
		_w3121_
	);
	LUT2 #(
		.INIT('h4)
	) name975 (
		_w3119_,
		_w3121_,
		_w3122_
	);
	LUT4 #(
		.INIT('hc4cc)
	) name976 (
		\u6_mem_reg[2][30]/NET0131 ,
		\u6_rp_reg[0]/P0001 ,
		\u6_rp_reg[1]/NET0131 ,
		\u6_rp_reg[2]/NET0131 ,
		_w3123_
	);
	LUT3 #(
		.INIT('h02)
	) name977 (
		\u6_mem_reg[0][30]/NET0131 ,
		\u6_rp_reg[1]/NET0131 ,
		\u6_rp_reg[2]/NET0131 ,
		_w3124_
	);
	LUT4 #(
		.INIT('h3f5f)
	) name978 (
		\u6_mem_reg[1][30]/NET0131 ,
		\u6_mem_reg[3][30]/NET0131 ,
		\u6_rp_reg[1]/NET0131 ,
		\u6_rp_reg[2]/NET0131 ,
		_w3125_
	);
	LUT3 #(
		.INIT('h40)
	) name979 (
		_w3124_,
		_w3123_,
		_w3125_,
		_w3126_
	);
	LUT4 #(
		.INIT('h8ccc)
	) name980 (
		\u6_rp_reg[0]/P0001 ,
		_w2445_,
		_w3077_,
		_w3078_,
		_w3127_
	);
	LUT3 #(
		.INIT('h2a)
	) name981 (
		_w3017_,
		_w3103_,
		_w3104_,
		_w3128_
	);
	LUT4 #(
		.INIT('h3f5f)
	) name982 (
		\u6_mem_reg[1][18]/NET0131 ,
		\u6_mem_reg[3][18]/NET0131 ,
		\u6_rp_reg[1]/NET0131 ,
		\u6_rp_reg[2]/NET0131 ,
		_w3129_
	);
	LUT4 #(
		.INIT('hf3f5)
	) name983 (
		\u6_mem_reg[0][18]/NET0131 ,
		\u6_mem_reg[2][18]/NET0131 ,
		\u6_rp_reg[1]/NET0131 ,
		\u6_rp_reg[2]/NET0131 ,
		_w3130_
	);
	LUT4 #(
		.INIT('ha222)
	) name984 (
		_w2444_,
		_w2516_,
		_w3129_,
		_w3130_,
		_w3131_
	);
	LUT4 #(
		.INIT('h0b00)
	) name985 (
		_w3126_,
		_w3127_,
		_w3128_,
		_w3131_,
		_w3132_
	);
	LUT4 #(
		.INIT('h0b0f)
	) name986 (
		\u14_u3_en_out_l2_reg/P0001 ,
		\u14_u3_en_out_l_reg/NET0131 ,
		\u6_dout_reg[18]/P0001 ,
		\valid_s_reg/NET0131 ,
		_w3133_
	);
	LUT2 #(
		.INIT('h2)
	) name987 (
		\u13_occ0_r_reg[24]/NET0131 ,
		_w3133_,
		_w3134_
	);
	LUT2 #(
		.INIT('h4)
	) name988 (
		_w3132_,
		_w3134_,
		_w3135_
	);
	LUT4 #(
		.INIT('hc4cc)
	) name989 (
		\u6_mem_reg[2][31]/NET0131 ,
		\u6_rp_reg[0]/P0001 ,
		\u6_rp_reg[1]/NET0131 ,
		\u6_rp_reg[2]/NET0131 ,
		_w3136_
	);
	LUT3 #(
		.INIT('h02)
	) name990 (
		\u6_mem_reg[0][31]/NET0131 ,
		\u6_rp_reg[1]/NET0131 ,
		\u6_rp_reg[2]/NET0131 ,
		_w3137_
	);
	LUT4 #(
		.INIT('h3f5f)
	) name991 (
		\u6_mem_reg[1][31]/NET0131 ,
		\u6_mem_reg[3][31]/NET0131 ,
		\u6_rp_reg[1]/NET0131 ,
		\u6_rp_reg[2]/NET0131 ,
		_w3138_
	);
	LUT3 #(
		.INIT('h40)
	) name992 (
		_w3137_,
		_w3136_,
		_w3138_,
		_w3139_
	);
	LUT4 #(
		.INIT('h8ccc)
	) name993 (
		\u6_rp_reg[0]/P0001 ,
		_w2445_,
		_w3090_,
		_w3091_,
		_w3140_
	);
	LUT3 #(
		.INIT('h2a)
	) name994 (
		_w3017_,
		_w3116_,
		_w3117_,
		_w3141_
	);
	LUT4 #(
		.INIT('h35ff)
	) name995 (
		\u6_mem_reg[2][19]/NET0131 ,
		\u6_mem_reg[3][19]/NET0131 ,
		\u6_rp_reg[1]/NET0131 ,
		\u6_rp_reg[2]/NET0131 ,
		_w3142_
	);
	LUT4 #(
		.INIT('hff35)
	) name996 (
		\u6_mem_reg[0][19]/NET0131 ,
		\u6_mem_reg[1][19]/NET0131 ,
		\u6_rp_reg[1]/NET0131 ,
		\u6_rp_reg[2]/NET0131 ,
		_w3143_
	);
	LUT4 #(
		.INIT('ha222)
	) name997 (
		_w2444_,
		_w2516_,
		_w3142_,
		_w3143_,
		_w3144_
	);
	LUT4 #(
		.INIT('h0b00)
	) name998 (
		_w3139_,
		_w3140_,
		_w3141_,
		_w3144_,
		_w3145_
	);
	LUT4 #(
		.INIT('h0b0f)
	) name999 (
		\u14_u3_en_out_l2_reg/P0001 ,
		\u14_u3_en_out_l_reg/NET0131 ,
		\u6_dout_reg[19]/P0001 ,
		\valid_s_reg/NET0131 ,
		_w3146_
	);
	LUT2 #(
		.INIT('h2)
	) name1000 (
		\u13_occ0_r_reg[24]/NET0131 ,
		_w3146_,
		_w3147_
	);
	LUT2 #(
		.INIT('h4)
	) name1001 (
		_w3145_,
		_w3147_,
		_w3148_
	);
	LUT4 #(
		.INIT('h35ff)
	) name1002 (
		\u6_mem_reg[2][2]/NET0131 ,
		\u6_mem_reg[3][2]/NET0131 ,
		\u6_rp_reg[1]/NET0131 ,
		\u6_rp_reg[2]/NET0131 ,
		_w3149_
	);
	LUT4 #(
		.INIT('hff35)
	) name1003 (
		\u6_mem_reg[0][2]/NET0131 ,
		\u6_mem_reg[1][2]/NET0131 ,
		\u6_rp_reg[1]/NET0131 ,
		\u6_rp_reg[2]/NET0131 ,
		_w3150_
	);
	LUT3 #(
		.INIT('h2a)
	) name1004 (
		_w2516_,
		_w3149_,
		_w3150_,
		_w3151_
	);
	LUT4 #(
		.INIT('h80aa)
	) name1005 (
		_w2444_,
		_w2514_,
		_w2515_,
		_w3017_,
		_w3152_
	);
	LUT4 #(
		.INIT('h0b0f)
	) name1006 (
		\u14_u3_en_out_l2_reg/P0001 ,
		\u14_u3_en_out_l_reg/NET0131 ,
		\u6_dout_reg[2]/P0001 ,
		\valid_s_reg/NET0131 ,
		_w3153_
	);
	LUT2 #(
		.INIT('h2)
	) name1007 (
		\u13_occ0_r_reg[24]/NET0131 ,
		_w3153_,
		_w3154_
	);
	LUT3 #(
		.INIT('hb0)
	) name1008 (
		_w3151_,
		_w3152_,
		_w3154_,
		_w3155_
	);
	LUT4 #(
		.INIT('h3f5f)
	) name1009 (
		\u6_mem_reg[1][3]/NET0131 ,
		\u6_mem_reg[3][3]/NET0131 ,
		\u6_rp_reg[1]/NET0131 ,
		\u6_rp_reg[2]/NET0131 ,
		_w3156_
	);
	LUT4 #(
		.INIT('hf3f5)
	) name1010 (
		\u6_mem_reg[0][3]/NET0131 ,
		\u6_mem_reg[2][3]/NET0131 ,
		\u6_rp_reg[1]/NET0131 ,
		\u6_rp_reg[2]/NET0131 ,
		_w3157_
	);
	LUT3 #(
		.INIT('h2a)
	) name1011 (
		_w2516_,
		_w3156_,
		_w3157_,
		_w3158_
	);
	LUT4 #(
		.INIT('h80aa)
	) name1012 (
		_w2444_,
		_w2521_,
		_w2522_,
		_w3017_,
		_w3159_
	);
	LUT4 #(
		.INIT('h0b0f)
	) name1013 (
		\u14_u3_en_out_l2_reg/P0001 ,
		\u14_u3_en_out_l_reg/NET0131 ,
		\u6_dout_reg[3]/P0001 ,
		\valid_s_reg/NET0131 ,
		_w3160_
	);
	LUT2 #(
		.INIT('h2)
	) name1014 (
		\u13_occ0_r_reg[24]/NET0131 ,
		_w3160_,
		_w3161_
	);
	LUT3 #(
		.INIT('hb0)
	) name1015 (
		_w3158_,
		_w3159_,
		_w3161_,
		_w3162_
	);
	LUT3 #(
		.INIT('h80)
	) name1016 (
		\u6_rp_reg[0]/P0001 ,
		_w3103_,
		_w3104_,
		_w3163_
	);
	LUT4 #(
		.INIT('h8ccc)
	) name1017 (
		\u6_rp_reg[0]/P0001 ,
		_w2445_,
		_w2514_,
		_w2515_,
		_w3164_
	);
	LUT3 #(
		.INIT('h2a)
	) name1018 (
		_w3017_,
		_w3149_,
		_w3150_,
		_w3165_
	);
	LUT4 #(
		.INIT('h35ff)
	) name1019 (
		\u6_mem_reg[2][4]/NET0131 ,
		\u6_mem_reg[3][4]/NET0131 ,
		\u6_rp_reg[1]/NET0131 ,
		\u6_rp_reg[2]/NET0131 ,
		_w3166_
	);
	LUT4 #(
		.INIT('hff35)
	) name1020 (
		\u6_mem_reg[0][4]/NET0131 ,
		\u6_mem_reg[1][4]/NET0131 ,
		\u6_rp_reg[1]/NET0131 ,
		\u6_rp_reg[2]/NET0131 ,
		_w3167_
	);
	LUT4 #(
		.INIT('ha222)
	) name1021 (
		_w2444_,
		_w2516_,
		_w3166_,
		_w3167_,
		_w3168_
	);
	LUT4 #(
		.INIT('h0b00)
	) name1022 (
		_w3163_,
		_w3164_,
		_w3165_,
		_w3168_,
		_w3169_
	);
	LUT4 #(
		.INIT('h0b0f)
	) name1023 (
		\u14_u3_en_out_l2_reg/P0001 ,
		\u14_u3_en_out_l_reg/NET0131 ,
		\u6_dout_reg[4]/P0001 ,
		\valid_s_reg/NET0131 ,
		_w3170_
	);
	LUT2 #(
		.INIT('h2)
	) name1024 (
		\u13_occ0_r_reg[24]/NET0131 ,
		_w3170_,
		_w3171_
	);
	LUT2 #(
		.INIT('h4)
	) name1025 (
		_w3169_,
		_w3171_,
		_w3172_
	);
	LUT3 #(
		.INIT('h80)
	) name1026 (
		\u6_rp_reg[0]/P0001 ,
		_w3116_,
		_w3117_,
		_w3173_
	);
	LUT4 #(
		.INIT('h8ccc)
	) name1027 (
		\u6_rp_reg[0]/P0001 ,
		_w2445_,
		_w2521_,
		_w2522_,
		_w3174_
	);
	LUT3 #(
		.INIT('h2a)
	) name1028 (
		_w3017_,
		_w3156_,
		_w3157_,
		_w3175_
	);
	LUT4 #(
		.INIT('h35ff)
	) name1029 (
		\u6_mem_reg[2][5]/NET0131 ,
		\u6_mem_reg[3][5]/NET0131 ,
		\u6_rp_reg[1]/NET0131 ,
		\u6_rp_reg[2]/NET0131 ,
		_w3176_
	);
	LUT4 #(
		.INIT('hff35)
	) name1030 (
		\u6_mem_reg[0][5]/NET0131 ,
		\u6_mem_reg[1][5]/NET0131 ,
		\u6_rp_reg[1]/NET0131 ,
		\u6_rp_reg[2]/NET0131 ,
		_w3177_
	);
	LUT4 #(
		.INIT('ha222)
	) name1031 (
		_w2444_,
		_w2516_,
		_w3176_,
		_w3177_,
		_w3178_
	);
	LUT4 #(
		.INIT('h0b00)
	) name1032 (
		_w3173_,
		_w3174_,
		_w3175_,
		_w3178_,
		_w3179_
	);
	LUT4 #(
		.INIT('h0b0f)
	) name1033 (
		\u14_u3_en_out_l2_reg/P0001 ,
		\u14_u3_en_out_l_reg/NET0131 ,
		\u6_dout_reg[5]/P0001 ,
		\valid_s_reg/NET0131 ,
		_w3180_
	);
	LUT2 #(
		.INIT('h2)
	) name1034 (
		\u13_occ0_r_reg[24]/NET0131 ,
		_w3180_,
		_w3181_
	);
	LUT2 #(
		.INIT('h4)
	) name1035 (
		_w3179_,
		_w3181_,
		_w3182_
	);
	LUT3 #(
		.INIT('h80)
	) name1036 (
		\u6_rp_reg[0]/P0001 ,
		_w3129_,
		_w3130_,
		_w3183_
	);
	LUT4 #(
		.INIT('h8ccc)
	) name1037 (
		\u6_rp_reg[0]/P0001 ,
		_w2445_,
		_w3149_,
		_w3150_,
		_w3184_
	);
	LUT3 #(
		.INIT('h2a)
	) name1038 (
		_w3017_,
		_w3166_,
		_w3167_,
		_w3185_
	);
	LUT4 #(
		.INIT('ha222)
	) name1039 (
		_w2444_,
		_w2516_,
		_w3014_,
		_w3015_,
		_w3186_
	);
	LUT4 #(
		.INIT('h0b00)
	) name1040 (
		_w3183_,
		_w3184_,
		_w3185_,
		_w3186_,
		_w3187_
	);
	LUT4 #(
		.INIT('h0b0f)
	) name1041 (
		\u14_u3_en_out_l2_reg/P0001 ,
		\u14_u3_en_out_l_reg/NET0131 ,
		\u6_dout_reg[6]/P0001 ,
		\valid_s_reg/NET0131 ,
		_w3188_
	);
	LUT2 #(
		.INIT('h2)
	) name1042 (
		\u13_occ0_r_reg[24]/NET0131 ,
		_w3188_,
		_w3189_
	);
	LUT2 #(
		.INIT('h4)
	) name1043 (
		_w3187_,
		_w3189_,
		_w3190_
	);
	LUT3 #(
		.INIT('h80)
	) name1044 (
		\u6_rp_reg[0]/P0001 ,
		_w3142_,
		_w3143_,
		_w3191_
	);
	LUT4 #(
		.INIT('h8ccc)
	) name1045 (
		\u6_rp_reg[0]/P0001 ,
		_w2445_,
		_w3156_,
		_w3157_,
		_w3192_
	);
	LUT3 #(
		.INIT('h2a)
	) name1046 (
		_w3017_,
		_w3176_,
		_w3177_,
		_w3193_
	);
	LUT4 #(
		.INIT('ha222)
	) name1047 (
		_w2444_,
		_w2516_,
		_w3032_,
		_w3033_,
		_w3194_
	);
	LUT4 #(
		.INIT('h0b00)
	) name1048 (
		_w3191_,
		_w3192_,
		_w3193_,
		_w3194_,
		_w3195_
	);
	LUT4 #(
		.INIT('h0b0f)
	) name1049 (
		\u14_u3_en_out_l2_reg/P0001 ,
		\u14_u3_en_out_l_reg/NET0131 ,
		\u6_dout_reg[7]/P0001 ,
		\valid_s_reg/NET0131 ,
		_w3196_
	);
	LUT2 #(
		.INIT('h2)
	) name1050 (
		\u13_occ0_r_reg[24]/NET0131 ,
		_w3196_,
		_w3197_
	);
	LUT2 #(
		.INIT('h4)
	) name1051 (
		_w3195_,
		_w3197_,
		_w3198_
	);
	LUT4 #(
		.INIT('hc4cc)
	) name1052 (
		\u6_mem_reg[2][20]/NET0131 ,
		\u6_rp_reg[0]/P0001 ,
		\u6_rp_reg[1]/NET0131 ,
		\u6_rp_reg[2]/NET0131 ,
		_w3199_
	);
	LUT3 #(
		.INIT('h02)
	) name1053 (
		\u6_mem_reg[0][20]/NET0131 ,
		\u6_rp_reg[1]/NET0131 ,
		\u6_rp_reg[2]/NET0131 ,
		_w3200_
	);
	LUT4 #(
		.INIT('h3f5f)
	) name1054 (
		\u6_mem_reg[1][20]/NET0131 ,
		\u6_mem_reg[3][20]/NET0131 ,
		\u6_rp_reg[1]/NET0131 ,
		\u6_rp_reg[2]/NET0131 ,
		_w3201_
	);
	LUT3 #(
		.INIT('h40)
	) name1055 (
		_w3200_,
		_w3199_,
		_w3201_,
		_w3202_
	);
	LUT4 #(
		.INIT('h8ccc)
	) name1056 (
		\u6_rp_reg[0]/P0001 ,
		_w2445_,
		_w3166_,
		_w3167_,
		_w3203_
	);
	LUT3 #(
		.INIT('h70)
	) name1057 (
		_w3014_,
		_w3015_,
		_w3017_,
		_w3204_
	);
	LUT4 #(
		.INIT('ha222)
	) name1058 (
		_w2444_,
		_w2516_,
		_w3018_,
		_w3019_,
		_w3205_
	);
	LUT4 #(
		.INIT('h0b00)
	) name1059 (
		_w3202_,
		_w3203_,
		_w3204_,
		_w3205_,
		_w3206_
	);
	LUT4 #(
		.INIT('h0b0f)
	) name1060 (
		\u14_u3_en_out_l2_reg/P0001 ,
		\u14_u3_en_out_l_reg/NET0131 ,
		\u6_dout_reg[8]/P0001 ,
		\valid_s_reg/NET0131 ,
		_w3207_
	);
	LUT2 #(
		.INIT('h2)
	) name1061 (
		\u13_occ0_r_reg[24]/NET0131 ,
		_w3207_,
		_w3208_
	);
	LUT2 #(
		.INIT('h4)
	) name1062 (
		_w3206_,
		_w3208_,
		_w3209_
	);
	LUT4 #(
		.INIT('hc4cc)
	) name1063 (
		\u6_mem_reg[2][21]/NET0131 ,
		\u6_rp_reg[0]/P0001 ,
		\u6_rp_reg[1]/NET0131 ,
		\u6_rp_reg[2]/NET0131 ,
		_w3210_
	);
	LUT3 #(
		.INIT('h02)
	) name1064 (
		\u6_mem_reg[0][21]/NET0131 ,
		\u6_rp_reg[1]/NET0131 ,
		\u6_rp_reg[2]/NET0131 ,
		_w3211_
	);
	LUT4 #(
		.INIT('h3f5f)
	) name1065 (
		\u6_mem_reg[1][21]/NET0131 ,
		\u6_mem_reg[3][21]/NET0131 ,
		\u6_rp_reg[1]/NET0131 ,
		\u6_rp_reg[2]/NET0131 ,
		_w3212_
	);
	LUT3 #(
		.INIT('h40)
	) name1066 (
		_w3211_,
		_w3210_,
		_w3212_,
		_w3213_
	);
	LUT4 #(
		.INIT('h8ccc)
	) name1067 (
		\u6_rp_reg[0]/P0001 ,
		_w2445_,
		_w3176_,
		_w3177_,
		_w3214_
	);
	LUT3 #(
		.INIT('h2a)
	) name1068 (
		_w3017_,
		_w3032_,
		_w3033_,
		_w3215_
	);
	LUT4 #(
		.INIT('ha222)
	) name1069 (
		_w2444_,
		_w2516_,
		_w3035_,
		_w3036_,
		_w3216_
	);
	LUT4 #(
		.INIT('h0b00)
	) name1070 (
		_w3213_,
		_w3214_,
		_w3215_,
		_w3216_,
		_w3217_
	);
	LUT4 #(
		.INIT('h0b0f)
	) name1071 (
		\u14_u3_en_out_l2_reg/P0001 ,
		\u14_u3_en_out_l_reg/NET0131 ,
		\u6_dout_reg[9]/P0001 ,
		\valid_s_reg/NET0131 ,
		_w3218_
	);
	LUT2 #(
		.INIT('h2)
	) name1072 (
		\u13_occ0_r_reg[24]/NET0131 ,
		_w3218_,
		_w3219_
	);
	LUT2 #(
		.INIT('h4)
	) name1073 (
		_w3217_,
		_w3219_,
		_w3220_
	);
	LUT4 #(
		.INIT('h35ff)
	) name1074 (
		\u7_mem_reg[2][6]/NET0131 ,
		\u7_mem_reg[3][6]/NET0131 ,
		\u7_rp_reg[1]/NET0131 ,
		\u7_rp_reg[2]/NET0131 ,
		_w3221_
	);
	LUT4 #(
		.INIT('hff35)
	) name1075 (
		\u7_mem_reg[0][6]/NET0131 ,
		\u7_mem_reg[1][6]/NET0131 ,
		\u7_rp_reg[1]/NET0131 ,
		\u7_rp_reg[2]/NET0131 ,
		_w3222_
	);
	LUT4 #(
		.INIT('hc444)
	) name1076 (
		_w2453_,
		_w2455_,
		_w3221_,
		_w3222_,
		_w3223_
	);
	LUT4 #(
		.INIT('h35ff)
	) name1077 (
		\u7_mem_reg[2][10]/NET0131 ,
		\u7_mem_reg[3][10]/NET0131 ,
		\u7_rp_reg[1]/NET0131 ,
		\u7_rp_reg[2]/NET0131 ,
		_w3224_
	);
	LUT4 #(
		.INIT('hff35)
	) name1078 (
		\u7_mem_reg[0][10]/NET0131 ,
		\u7_mem_reg[1][10]/NET0131 ,
		\u7_rp_reg[1]/NET0131 ,
		\u7_rp_reg[2]/NET0131 ,
		_w3225_
	);
	LUT3 #(
		.INIT('h2a)
	) name1079 (
		_w2529_,
		_w3224_,
		_w3225_,
		_w3226_
	);
	LUT2 #(
		.INIT('h2)
	) name1080 (
		\u13_occ1_r_reg[2]/NET0131 ,
		\u13_occ1_r_reg[3]/NET0131 ,
		_w3227_
	);
	LUT4 #(
		.INIT('h35ff)
	) name1081 (
		\u7_mem_reg[2][8]/NET0131 ,
		\u7_mem_reg[3][8]/NET0131 ,
		\u7_rp_reg[1]/NET0131 ,
		\u7_rp_reg[2]/NET0131 ,
		_w3228_
	);
	LUT4 #(
		.INIT('hff35)
	) name1082 (
		\u7_mem_reg[0][8]/NET0131 ,
		\u7_mem_reg[1][8]/NET0131 ,
		\u7_rp_reg[1]/NET0131 ,
		\u7_rp_reg[2]/NET0131 ,
		_w3229_
	);
	LUT3 #(
		.INIT('h2a)
	) name1083 (
		_w3227_,
		_w3228_,
		_w3229_,
		_w3230_
	);
	LUT3 #(
		.INIT('h10)
	) name1084 (
		\u13_occ1_r_reg[2]/NET0131 ,
		\u13_occ1_r_reg[3]/NET0131 ,
		\u7_rp_reg[0]/P0001 ,
		_w3231_
	);
	LUT4 #(
		.INIT('h3ff5)
	) name1085 (
		\u7_mem_reg[0][22]/NET0131 ,
		\u7_mem_reg[3][22]/NET0131 ,
		\u7_rp_reg[1]/NET0131 ,
		\u7_rp_reg[2]/NET0131 ,
		_w3232_
	);
	LUT4 #(
		.INIT('hf35f)
	) name1086 (
		\u7_mem_reg[1][22]/NET0131 ,
		\u7_mem_reg[2][22]/NET0131 ,
		\u7_rp_reg[1]/NET0131 ,
		\u7_rp_reg[2]/NET0131 ,
		_w3233_
	);
	LUT3 #(
		.INIT('h2a)
	) name1087 (
		_w3231_,
		_w3232_,
		_w3233_,
		_w3234_
	);
	LUT4 #(
		.INIT('h0100)
	) name1088 (
		_w3230_,
		_w3234_,
		_w3226_,
		_w3223_,
		_w3235_
	);
	LUT4 #(
		.INIT('h0b0f)
	) name1089 (
		\u14_u4_en_out_l2_reg/P0001 ,
		\u14_u4_en_out_l_reg/NET0131 ,
		\u7_dout_reg[10]/P0001 ,
		\valid_s_reg/NET0131 ,
		_w3236_
	);
	LUT2 #(
		.INIT('h2)
	) name1090 (
		\u13_occ1_r_reg[0]/NET0131 ,
		_w3236_,
		_w3237_
	);
	LUT2 #(
		.INIT('h4)
	) name1091 (
		_w3235_,
		_w3237_,
		_w3238_
	);
	LUT4 #(
		.INIT('hf35f)
	) name1092 (
		\u7_mem_reg[1][11]/NET0131 ,
		\u7_mem_reg[2][11]/NET0131 ,
		\u7_rp_reg[1]/NET0131 ,
		\u7_rp_reg[2]/NET0131 ,
		_w3239_
	);
	LUT4 #(
		.INIT('h3ff5)
	) name1093 (
		\u7_mem_reg[0][11]/NET0131 ,
		\u7_mem_reg[3][11]/NET0131 ,
		\u7_rp_reg[1]/NET0131 ,
		\u7_rp_reg[2]/NET0131 ,
		_w3240_
	);
	LUT4 #(
		.INIT('ha222)
	) name1094 (
		_w2455_,
		_w2529_,
		_w3239_,
		_w3240_,
		_w3241_
	);
	LUT4 #(
		.INIT('h3ff5)
	) name1095 (
		\u7_mem_reg[0][9]/NET0131 ,
		\u7_mem_reg[3][9]/NET0131 ,
		\u7_rp_reg[1]/NET0131 ,
		\u7_rp_reg[2]/NET0131 ,
		_w3242_
	);
	LUT4 #(
		.INIT('hf35f)
	) name1096 (
		\u7_mem_reg[1][9]/NET0131 ,
		\u7_mem_reg[2][9]/NET0131 ,
		\u7_rp_reg[1]/NET0131 ,
		\u7_rp_reg[2]/NET0131 ,
		_w3243_
	);
	LUT3 #(
		.INIT('h2a)
	) name1097 (
		_w3227_,
		_w3242_,
		_w3243_,
		_w3244_
	);
	LUT4 #(
		.INIT('h3f5f)
	) name1098 (
		\u7_mem_reg[1][7]/NET0131 ,
		\u7_mem_reg[3][7]/NET0131 ,
		\u7_rp_reg[1]/NET0131 ,
		\u7_rp_reg[2]/NET0131 ,
		_w3245_
	);
	LUT4 #(
		.INIT('hf3f5)
	) name1099 (
		\u7_mem_reg[0][7]/NET0131 ,
		\u7_mem_reg[2][7]/NET0131 ,
		\u7_rp_reg[1]/NET0131 ,
		\u7_rp_reg[2]/NET0131 ,
		_w3246_
	);
	LUT3 #(
		.INIT('h2a)
	) name1100 (
		_w2453_,
		_w3245_,
		_w3246_,
		_w3247_
	);
	LUT4 #(
		.INIT('hf3f5)
	) name1101 (
		\u7_mem_reg[0][23]/NET0131 ,
		\u7_mem_reg[2][23]/NET0131 ,
		\u7_rp_reg[1]/NET0131 ,
		\u7_rp_reg[2]/NET0131 ,
		_w3248_
	);
	LUT4 #(
		.INIT('h3f5f)
	) name1102 (
		\u7_mem_reg[1][23]/NET0131 ,
		\u7_mem_reg[3][23]/NET0131 ,
		\u7_rp_reg[1]/NET0131 ,
		\u7_rp_reg[2]/NET0131 ,
		_w3249_
	);
	LUT3 #(
		.INIT('h2a)
	) name1103 (
		_w3231_,
		_w3248_,
		_w3249_,
		_w3250_
	);
	LUT4 #(
		.INIT('h0100)
	) name1104 (
		_w3247_,
		_w3250_,
		_w3244_,
		_w3241_,
		_w3251_
	);
	LUT4 #(
		.INIT('h0b0f)
	) name1105 (
		\u14_u4_en_out_l2_reg/P0001 ,
		\u14_u4_en_out_l_reg/NET0131 ,
		\u7_dout_reg[11]/P0001 ,
		\valid_s_reg/NET0131 ,
		_w3252_
	);
	LUT2 #(
		.INIT('h2)
	) name1106 (
		\u13_occ1_r_reg[0]/NET0131 ,
		_w3252_,
		_w3253_
	);
	LUT2 #(
		.INIT('h4)
	) name1107 (
		_w3251_,
		_w3253_,
		_w3254_
	);
	LUT4 #(
		.INIT('h0105)
	) name1108 (
		\u13_icc_r_reg[4]/NET0131 ,
		\u13_icc_r_reg[5]/NET0131 ,
		\u9_status_reg[0]/P0001 ,
		\u9_status_reg[1]/P0001 ,
		_w3255_
	);
	LUT3 #(
		.INIT('h32)
	) name1109 (
		\u13_icc_r_reg[5]/NET0131 ,
		\u9_full_reg/NET0131 ,
		\u9_status_reg[1]/P0001 ,
		_w3256_
	);
	LUT3 #(
		.INIT('h8a)
	) name1110 (
		\u13_icc_r_reg[0]/NET0131 ,
		_w3255_,
		_w3256_,
		_w3257_
	);
	LUT4 #(
		.INIT('hc4cc)
	) name1111 (
		\u7_mem_reg[2][24]/NET0131 ,
		\u7_rp_reg[0]/P0001 ,
		\u7_rp_reg[1]/NET0131 ,
		\u7_rp_reg[2]/NET0131 ,
		_w3258_
	);
	LUT3 #(
		.INIT('h02)
	) name1112 (
		\u7_mem_reg[0][24]/NET0131 ,
		\u7_rp_reg[1]/NET0131 ,
		\u7_rp_reg[2]/NET0131 ,
		_w3259_
	);
	LUT4 #(
		.INIT('h3f5f)
	) name1113 (
		\u7_mem_reg[1][24]/NET0131 ,
		\u7_mem_reg[3][24]/NET0131 ,
		\u7_rp_reg[1]/NET0131 ,
		\u7_rp_reg[2]/NET0131 ,
		_w3260_
	);
	LUT3 #(
		.INIT('h40)
	) name1114 (
		_w3259_,
		_w3258_,
		_w3260_,
		_w3261_
	);
	LUT4 #(
		.INIT('h8ccc)
	) name1115 (
		\u7_rp_reg[0]/P0001 ,
		_w2452_,
		_w3228_,
		_w3229_,
		_w3262_
	);
	LUT3 #(
		.INIT('h2a)
	) name1116 (
		_w3227_,
		_w3224_,
		_w3225_,
		_w3263_
	);
	LUT4 #(
		.INIT('h35ff)
	) name1117 (
		\u7_mem_reg[2][12]/NET0131 ,
		\u7_mem_reg[3][12]/NET0131 ,
		\u7_rp_reg[1]/NET0131 ,
		\u7_rp_reg[2]/NET0131 ,
		_w3264_
	);
	LUT4 #(
		.INIT('hff35)
	) name1118 (
		\u7_mem_reg[0][12]/NET0131 ,
		\u7_mem_reg[1][12]/NET0131 ,
		\u7_rp_reg[1]/NET0131 ,
		\u7_rp_reg[2]/NET0131 ,
		_w3265_
	);
	LUT4 #(
		.INIT('ha222)
	) name1119 (
		_w2455_,
		_w2529_,
		_w3264_,
		_w3265_,
		_w3266_
	);
	LUT4 #(
		.INIT('h0b00)
	) name1120 (
		_w3261_,
		_w3262_,
		_w3263_,
		_w3266_,
		_w3267_
	);
	LUT4 #(
		.INIT('h0b0f)
	) name1121 (
		\u14_u4_en_out_l2_reg/P0001 ,
		\u14_u4_en_out_l_reg/NET0131 ,
		\u7_dout_reg[12]/P0001 ,
		\valid_s_reg/NET0131 ,
		_w3268_
	);
	LUT2 #(
		.INIT('h2)
	) name1122 (
		\u13_occ1_r_reg[0]/NET0131 ,
		_w3268_,
		_w3269_
	);
	LUT2 #(
		.INIT('h4)
	) name1123 (
		_w3267_,
		_w3269_,
		_w3270_
	);
	LUT4 #(
		.INIT('h0105)
	) name1124 (
		\u10_status_reg[0]/P0001 ,
		\u10_status_reg[1]/P0001 ,
		\u13_icc_r_reg[12]/NET0131 ,
		\u13_icc_r_reg[13]/NET0131 ,
		_w3271_
	);
	LUT3 #(
		.INIT('h54)
	) name1125 (
		\u10_full_reg/NET0131 ,
		\u10_status_reg[1]/P0001 ,
		\u13_icc_r_reg[13]/NET0131 ,
		_w3272_
	);
	LUT3 #(
		.INIT('h8a)
	) name1126 (
		\u13_icc_r_reg[8]/NET0131 ,
		_w3271_,
		_w3272_,
		_w3273_
	);
	LUT4 #(
		.INIT('hc4cc)
	) name1127 (
		\u7_mem_reg[2][25]/NET0131 ,
		\u7_rp_reg[0]/P0001 ,
		\u7_rp_reg[1]/NET0131 ,
		\u7_rp_reg[2]/NET0131 ,
		_w3274_
	);
	LUT3 #(
		.INIT('h02)
	) name1128 (
		\u7_mem_reg[0][25]/NET0131 ,
		\u7_rp_reg[1]/NET0131 ,
		\u7_rp_reg[2]/NET0131 ,
		_w3275_
	);
	LUT4 #(
		.INIT('h3f5f)
	) name1129 (
		\u7_mem_reg[1][25]/NET0131 ,
		\u7_mem_reg[3][25]/NET0131 ,
		\u7_rp_reg[1]/NET0131 ,
		\u7_rp_reg[2]/NET0131 ,
		_w3276_
	);
	LUT3 #(
		.INIT('h40)
	) name1130 (
		_w3275_,
		_w3274_,
		_w3276_,
		_w3277_
	);
	LUT4 #(
		.INIT('h8ccc)
	) name1131 (
		\u7_rp_reg[0]/P0001 ,
		_w2452_,
		_w3242_,
		_w3243_,
		_w3278_
	);
	LUT4 #(
		.INIT('h35ff)
	) name1132 (
		\u7_mem_reg[2][13]/NET0131 ,
		\u7_mem_reg[3][13]/NET0131 ,
		\u7_rp_reg[1]/NET0131 ,
		\u7_rp_reg[2]/NET0131 ,
		_w3279_
	);
	LUT4 #(
		.INIT('hff35)
	) name1133 (
		\u7_mem_reg[0][13]/NET0131 ,
		\u7_mem_reg[1][13]/NET0131 ,
		\u7_rp_reg[1]/NET0131 ,
		\u7_rp_reg[2]/NET0131 ,
		_w3280_
	);
	LUT3 #(
		.INIT('h2a)
	) name1134 (
		_w2529_,
		_w3279_,
		_w3280_,
		_w3281_
	);
	LUT4 #(
		.INIT('ha222)
	) name1135 (
		_w2455_,
		_w3227_,
		_w3239_,
		_w3240_,
		_w3282_
	);
	LUT4 #(
		.INIT('h4500)
	) name1136 (
		_w3281_,
		_w3277_,
		_w3278_,
		_w3282_,
		_w3283_
	);
	LUT4 #(
		.INIT('h0b0f)
	) name1137 (
		\u14_u4_en_out_l2_reg/P0001 ,
		\u14_u4_en_out_l_reg/NET0131 ,
		\u7_dout_reg[13]/P0001 ,
		\valid_s_reg/NET0131 ,
		_w3284_
	);
	LUT2 #(
		.INIT('h2)
	) name1138 (
		\u13_occ1_r_reg[0]/NET0131 ,
		_w3284_,
		_w3285_
	);
	LUT2 #(
		.INIT('h4)
	) name1139 (
		_w3283_,
		_w3285_,
		_w3286_
	);
	LUT4 #(
		.INIT('hc4cc)
	) name1140 (
		\u7_mem_reg[2][26]/NET0131 ,
		\u7_rp_reg[0]/P0001 ,
		\u7_rp_reg[1]/NET0131 ,
		\u7_rp_reg[2]/NET0131 ,
		_w3287_
	);
	LUT3 #(
		.INIT('h02)
	) name1141 (
		\u7_mem_reg[0][26]/NET0131 ,
		\u7_rp_reg[1]/NET0131 ,
		\u7_rp_reg[2]/NET0131 ,
		_w3288_
	);
	LUT4 #(
		.INIT('h3f5f)
	) name1142 (
		\u7_mem_reg[1][26]/NET0131 ,
		\u7_mem_reg[3][26]/NET0131 ,
		\u7_rp_reg[1]/NET0131 ,
		\u7_rp_reg[2]/NET0131 ,
		_w3289_
	);
	LUT3 #(
		.INIT('h40)
	) name1143 (
		_w3288_,
		_w3287_,
		_w3289_,
		_w3290_
	);
	LUT4 #(
		.INIT('h8ccc)
	) name1144 (
		\u7_rp_reg[0]/P0001 ,
		_w2452_,
		_w3224_,
		_w3225_,
		_w3291_
	);
	LUT3 #(
		.INIT('h2a)
	) name1145 (
		_w3227_,
		_w3264_,
		_w3265_,
		_w3292_
	);
	LUT4 #(
		.INIT('h35ff)
	) name1146 (
		\u7_mem_reg[2][14]/NET0131 ,
		\u7_mem_reg[3][14]/NET0131 ,
		\u7_rp_reg[1]/NET0131 ,
		\u7_rp_reg[2]/NET0131 ,
		_w3293_
	);
	LUT4 #(
		.INIT('hff35)
	) name1147 (
		\u7_mem_reg[0][14]/NET0131 ,
		\u7_mem_reg[1][14]/NET0131 ,
		\u7_rp_reg[1]/NET0131 ,
		\u7_rp_reg[2]/NET0131 ,
		_w3294_
	);
	LUT4 #(
		.INIT('ha222)
	) name1148 (
		_w2455_,
		_w2529_,
		_w3293_,
		_w3294_,
		_w3295_
	);
	LUT4 #(
		.INIT('h0b00)
	) name1149 (
		_w3290_,
		_w3291_,
		_w3292_,
		_w3295_,
		_w3296_
	);
	LUT4 #(
		.INIT('h0b0f)
	) name1150 (
		\u14_u4_en_out_l2_reg/P0001 ,
		\u14_u4_en_out_l_reg/NET0131 ,
		\u7_dout_reg[14]/P0001 ,
		\valid_s_reg/NET0131 ,
		_w3297_
	);
	LUT2 #(
		.INIT('h2)
	) name1151 (
		\u13_occ1_r_reg[0]/NET0131 ,
		_w3297_,
		_w3298_
	);
	LUT2 #(
		.INIT('h4)
	) name1152 (
		_w3296_,
		_w3298_,
		_w3299_
	);
	LUT4 #(
		.INIT('hc444)
	) name1153 (
		_w2453_,
		_w2455_,
		_w3239_,
		_w3240_,
		_w3300_
	);
	LUT4 #(
		.INIT('h3f5f)
	) name1154 (
		\u7_mem_reg[1][15]/NET0131 ,
		\u7_mem_reg[3][15]/NET0131 ,
		\u7_rp_reg[1]/NET0131 ,
		\u7_rp_reg[2]/NET0131 ,
		_w3301_
	);
	LUT4 #(
		.INIT('hf3f5)
	) name1155 (
		\u7_mem_reg[0][15]/NET0131 ,
		\u7_mem_reg[2][15]/NET0131 ,
		\u7_rp_reg[1]/NET0131 ,
		\u7_rp_reg[2]/NET0131 ,
		_w3302_
	);
	LUT3 #(
		.INIT('h2a)
	) name1156 (
		_w2529_,
		_w3301_,
		_w3302_,
		_w3303_
	);
	LUT3 #(
		.INIT('h2a)
	) name1157 (
		_w3227_,
		_w3279_,
		_w3280_,
		_w3304_
	);
	LUT4 #(
		.INIT('hff35)
	) name1158 (
		\u7_mem_reg[0][27]/NET0131 ,
		\u7_mem_reg[1][27]/NET0131 ,
		\u7_rp_reg[1]/NET0131 ,
		\u7_rp_reg[2]/NET0131 ,
		_w3305_
	);
	LUT4 #(
		.INIT('h35ff)
	) name1159 (
		\u7_mem_reg[2][27]/NET0131 ,
		\u7_mem_reg[3][27]/NET0131 ,
		\u7_rp_reg[1]/NET0131 ,
		\u7_rp_reg[2]/NET0131 ,
		_w3306_
	);
	LUT3 #(
		.INIT('h2a)
	) name1160 (
		_w3231_,
		_w3305_,
		_w3306_,
		_w3307_
	);
	LUT4 #(
		.INIT('h0100)
	) name1161 (
		_w3304_,
		_w3307_,
		_w3303_,
		_w3300_,
		_w3308_
	);
	LUT4 #(
		.INIT('h0b0f)
	) name1162 (
		\u14_u4_en_out_l2_reg/P0001 ,
		\u14_u4_en_out_l_reg/NET0131 ,
		\u7_dout_reg[15]/P0001 ,
		\valid_s_reg/NET0131 ,
		_w3309_
	);
	LUT2 #(
		.INIT('h2)
	) name1163 (
		\u13_occ1_r_reg[0]/NET0131 ,
		_w3309_,
		_w3310_
	);
	LUT2 #(
		.INIT('h4)
	) name1164 (
		_w3308_,
		_w3310_,
		_w3311_
	);
	LUT4 #(
		.INIT('hc4cc)
	) name1165 (
		\u7_mem_reg[2][28]/NET0131 ,
		\u7_rp_reg[0]/P0001 ,
		\u7_rp_reg[1]/NET0131 ,
		\u7_rp_reg[2]/NET0131 ,
		_w3312_
	);
	LUT3 #(
		.INIT('h02)
	) name1166 (
		\u7_mem_reg[0][28]/NET0131 ,
		\u7_rp_reg[1]/NET0131 ,
		\u7_rp_reg[2]/NET0131 ,
		_w3313_
	);
	LUT4 #(
		.INIT('h3f5f)
	) name1167 (
		\u7_mem_reg[1][28]/NET0131 ,
		\u7_mem_reg[3][28]/NET0131 ,
		\u7_rp_reg[1]/NET0131 ,
		\u7_rp_reg[2]/NET0131 ,
		_w3314_
	);
	LUT3 #(
		.INIT('h40)
	) name1168 (
		_w3313_,
		_w3312_,
		_w3314_,
		_w3315_
	);
	LUT4 #(
		.INIT('h8ccc)
	) name1169 (
		\u7_rp_reg[0]/P0001 ,
		_w2452_,
		_w3264_,
		_w3265_,
		_w3316_
	);
	LUT3 #(
		.INIT('h2a)
	) name1170 (
		_w3227_,
		_w3293_,
		_w3294_,
		_w3317_
	);
	LUT4 #(
		.INIT('h35ff)
	) name1171 (
		\u7_mem_reg[2][16]/NET0131 ,
		\u7_mem_reg[3][16]/NET0131 ,
		\u7_rp_reg[1]/NET0131 ,
		\u7_rp_reg[2]/NET0131 ,
		_w3318_
	);
	LUT4 #(
		.INIT('hff35)
	) name1172 (
		\u7_mem_reg[0][16]/NET0131 ,
		\u7_mem_reg[1][16]/NET0131 ,
		\u7_rp_reg[1]/NET0131 ,
		\u7_rp_reg[2]/NET0131 ,
		_w3319_
	);
	LUT4 #(
		.INIT('ha222)
	) name1173 (
		_w2455_,
		_w2529_,
		_w3318_,
		_w3319_,
		_w3320_
	);
	LUT4 #(
		.INIT('h0b00)
	) name1174 (
		_w3315_,
		_w3316_,
		_w3317_,
		_w3320_,
		_w3321_
	);
	LUT4 #(
		.INIT('h0b0f)
	) name1175 (
		\u14_u4_en_out_l2_reg/P0001 ,
		\u14_u4_en_out_l_reg/NET0131 ,
		\u7_dout_reg[16]/P0001 ,
		\valid_s_reg/NET0131 ,
		_w3322_
	);
	LUT2 #(
		.INIT('h2)
	) name1176 (
		\u13_occ1_r_reg[0]/NET0131 ,
		_w3322_,
		_w3323_
	);
	LUT2 #(
		.INIT('h4)
	) name1177 (
		_w3321_,
		_w3323_,
		_w3324_
	);
	LUT4 #(
		.INIT('hc4cc)
	) name1178 (
		\u7_mem_reg[2][29]/NET0131 ,
		\u7_rp_reg[0]/P0001 ,
		\u7_rp_reg[1]/NET0131 ,
		\u7_rp_reg[2]/NET0131 ,
		_w3325_
	);
	LUT3 #(
		.INIT('h02)
	) name1179 (
		\u7_mem_reg[0][29]/NET0131 ,
		\u7_rp_reg[1]/NET0131 ,
		\u7_rp_reg[2]/NET0131 ,
		_w3326_
	);
	LUT4 #(
		.INIT('h3f5f)
	) name1180 (
		\u7_mem_reg[1][29]/NET0131 ,
		\u7_mem_reg[3][29]/NET0131 ,
		\u7_rp_reg[1]/NET0131 ,
		\u7_rp_reg[2]/NET0131 ,
		_w3327_
	);
	LUT3 #(
		.INIT('h40)
	) name1181 (
		_w3326_,
		_w3325_,
		_w3327_,
		_w3328_
	);
	LUT4 #(
		.INIT('h8ccc)
	) name1182 (
		\u7_rp_reg[0]/P0001 ,
		_w2452_,
		_w3279_,
		_w3280_,
		_w3329_
	);
	LUT3 #(
		.INIT('h2a)
	) name1183 (
		_w3227_,
		_w3301_,
		_w3302_,
		_w3330_
	);
	LUT4 #(
		.INIT('h3f5f)
	) name1184 (
		\u7_mem_reg[1][17]/NET0131 ,
		\u7_mem_reg[3][17]/NET0131 ,
		\u7_rp_reg[1]/NET0131 ,
		\u7_rp_reg[2]/NET0131 ,
		_w3331_
	);
	LUT4 #(
		.INIT('hf3f5)
	) name1185 (
		\u7_mem_reg[0][17]/NET0131 ,
		\u7_mem_reg[2][17]/NET0131 ,
		\u7_rp_reg[1]/NET0131 ,
		\u7_rp_reg[2]/NET0131 ,
		_w3332_
	);
	LUT4 #(
		.INIT('ha222)
	) name1186 (
		_w2455_,
		_w2529_,
		_w3331_,
		_w3332_,
		_w3333_
	);
	LUT4 #(
		.INIT('h0b00)
	) name1187 (
		_w3328_,
		_w3329_,
		_w3330_,
		_w3333_,
		_w3334_
	);
	LUT4 #(
		.INIT('h0b0f)
	) name1188 (
		\u14_u4_en_out_l2_reg/P0001 ,
		\u14_u4_en_out_l_reg/NET0131 ,
		\u7_dout_reg[17]/P0001 ,
		\valid_s_reg/NET0131 ,
		_w3335_
	);
	LUT2 #(
		.INIT('h2)
	) name1189 (
		\u13_occ1_r_reg[0]/NET0131 ,
		_w3335_,
		_w3336_
	);
	LUT2 #(
		.INIT('h4)
	) name1190 (
		_w3334_,
		_w3336_,
		_w3337_
	);
	LUT4 #(
		.INIT('hc4cc)
	) name1191 (
		\u7_mem_reg[2][30]/NET0131 ,
		\u7_rp_reg[0]/P0001 ,
		\u7_rp_reg[1]/NET0131 ,
		\u7_rp_reg[2]/NET0131 ,
		_w3338_
	);
	LUT3 #(
		.INIT('h02)
	) name1192 (
		\u7_mem_reg[0][30]/NET0131 ,
		\u7_rp_reg[1]/NET0131 ,
		\u7_rp_reg[2]/NET0131 ,
		_w3339_
	);
	LUT4 #(
		.INIT('h3f5f)
	) name1193 (
		\u7_mem_reg[1][30]/NET0131 ,
		\u7_mem_reg[3][30]/NET0131 ,
		\u7_rp_reg[1]/NET0131 ,
		\u7_rp_reg[2]/NET0131 ,
		_w3340_
	);
	LUT3 #(
		.INIT('h40)
	) name1194 (
		_w3339_,
		_w3338_,
		_w3340_,
		_w3341_
	);
	LUT4 #(
		.INIT('h8ccc)
	) name1195 (
		\u7_rp_reg[0]/P0001 ,
		_w2452_,
		_w3293_,
		_w3294_,
		_w3342_
	);
	LUT3 #(
		.INIT('h2a)
	) name1196 (
		_w3227_,
		_w3318_,
		_w3319_,
		_w3343_
	);
	LUT4 #(
		.INIT('hf35f)
	) name1197 (
		\u7_mem_reg[1][18]/NET0131 ,
		\u7_mem_reg[2][18]/NET0131 ,
		\u7_rp_reg[1]/NET0131 ,
		\u7_rp_reg[2]/NET0131 ,
		_w3344_
	);
	LUT4 #(
		.INIT('h3ff5)
	) name1198 (
		\u7_mem_reg[0][18]/NET0131 ,
		\u7_mem_reg[3][18]/NET0131 ,
		\u7_rp_reg[1]/NET0131 ,
		\u7_rp_reg[2]/NET0131 ,
		_w3345_
	);
	LUT4 #(
		.INIT('ha222)
	) name1199 (
		_w2455_,
		_w2529_,
		_w3344_,
		_w3345_,
		_w3346_
	);
	LUT4 #(
		.INIT('h0b00)
	) name1200 (
		_w3341_,
		_w3342_,
		_w3343_,
		_w3346_,
		_w3347_
	);
	LUT4 #(
		.INIT('h0b0f)
	) name1201 (
		\u14_u4_en_out_l2_reg/P0001 ,
		\u14_u4_en_out_l_reg/NET0131 ,
		\u7_dout_reg[18]/P0001 ,
		\valid_s_reg/NET0131 ,
		_w3348_
	);
	LUT2 #(
		.INIT('h2)
	) name1202 (
		\u13_occ1_r_reg[0]/NET0131 ,
		_w3348_,
		_w3349_
	);
	LUT2 #(
		.INIT('h4)
	) name1203 (
		_w3347_,
		_w3349_,
		_w3350_
	);
	LUT4 #(
		.INIT('hc4cc)
	) name1204 (
		\u7_mem_reg[2][31]/NET0131 ,
		\u7_rp_reg[0]/P0001 ,
		\u7_rp_reg[1]/NET0131 ,
		\u7_rp_reg[2]/NET0131 ,
		_w3351_
	);
	LUT3 #(
		.INIT('h02)
	) name1205 (
		\u7_mem_reg[0][31]/NET0131 ,
		\u7_rp_reg[1]/NET0131 ,
		\u7_rp_reg[2]/NET0131 ,
		_w3352_
	);
	LUT4 #(
		.INIT('h3f5f)
	) name1206 (
		\u7_mem_reg[1][31]/NET0131 ,
		\u7_mem_reg[3][31]/NET0131 ,
		\u7_rp_reg[1]/NET0131 ,
		\u7_rp_reg[2]/NET0131 ,
		_w3353_
	);
	LUT3 #(
		.INIT('h40)
	) name1207 (
		_w3352_,
		_w3351_,
		_w3353_,
		_w3354_
	);
	LUT4 #(
		.INIT('h8ccc)
	) name1208 (
		\u7_rp_reg[0]/P0001 ,
		_w2452_,
		_w3301_,
		_w3302_,
		_w3355_
	);
	LUT3 #(
		.INIT('h2a)
	) name1209 (
		_w3227_,
		_w3331_,
		_w3332_,
		_w3356_
	);
	LUT4 #(
		.INIT('h3ff5)
	) name1210 (
		\u7_mem_reg[0][19]/NET0131 ,
		\u7_mem_reg[3][19]/NET0131 ,
		\u7_rp_reg[1]/NET0131 ,
		\u7_rp_reg[2]/NET0131 ,
		_w3357_
	);
	LUT4 #(
		.INIT('hf35f)
	) name1211 (
		\u7_mem_reg[1][19]/NET0131 ,
		\u7_mem_reg[2][19]/NET0131 ,
		\u7_rp_reg[1]/NET0131 ,
		\u7_rp_reg[2]/NET0131 ,
		_w3358_
	);
	LUT4 #(
		.INIT('ha222)
	) name1212 (
		_w2455_,
		_w2529_,
		_w3357_,
		_w3358_,
		_w3359_
	);
	LUT4 #(
		.INIT('h0b00)
	) name1213 (
		_w3354_,
		_w3355_,
		_w3356_,
		_w3359_,
		_w3360_
	);
	LUT4 #(
		.INIT('h0b0f)
	) name1214 (
		\u14_u4_en_out_l2_reg/P0001 ,
		\u14_u4_en_out_l_reg/NET0131 ,
		\u7_dout_reg[19]/P0001 ,
		\valid_s_reg/NET0131 ,
		_w3361_
	);
	LUT2 #(
		.INIT('h2)
	) name1215 (
		\u13_occ1_r_reg[0]/NET0131 ,
		_w3361_,
		_w3362_
	);
	LUT2 #(
		.INIT('h4)
	) name1216 (
		_w3360_,
		_w3362_,
		_w3363_
	);
	LUT4 #(
		.INIT('h35ff)
	) name1217 (
		\u7_mem_reg[2][2]/NET0131 ,
		\u7_mem_reg[3][2]/NET0131 ,
		\u7_rp_reg[1]/NET0131 ,
		\u7_rp_reg[2]/NET0131 ,
		_w3364_
	);
	LUT4 #(
		.INIT('hff35)
	) name1218 (
		\u7_mem_reg[0][2]/NET0131 ,
		\u7_mem_reg[1][2]/NET0131 ,
		\u7_rp_reg[1]/NET0131 ,
		\u7_rp_reg[2]/NET0131 ,
		_w3365_
	);
	LUT3 #(
		.INIT('h2a)
	) name1219 (
		_w2529_,
		_w3364_,
		_w3365_,
		_w3366_
	);
	LUT4 #(
		.INIT('h80aa)
	) name1220 (
		_w2455_,
		_w2527_,
		_w2528_,
		_w3227_,
		_w3367_
	);
	LUT4 #(
		.INIT('h0b0f)
	) name1221 (
		\u14_u4_en_out_l2_reg/P0001 ,
		\u14_u4_en_out_l_reg/NET0131 ,
		\u7_dout_reg[2]/P0001 ,
		\valid_s_reg/NET0131 ,
		_w3368_
	);
	LUT2 #(
		.INIT('h2)
	) name1222 (
		\u13_occ1_r_reg[0]/NET0131 ,
		_w3368_,
		_w3369_
	);
	LUT3 #(
		.INIT('hb0)
	) name1223 (
		_w3366_,
		_w3367_,
		_w3369_,
		_w3370_
	);
	LUT3 #(
		.INIT('h70)
	) name1224 (
		_w2534_,
		_w2535_,
		_w3227_,
		_w3371_
	);
	LUT4 #(
		.INIT('h3f5f)
	) name1225 (
		\u7_mem_reg[1][3]/NET0131 ,
		\u7_mem_reg[3][3]/NET0131 ,
		\u7_rp_reg[1]/NET0131 ,
		\u7_rp_reg[2]/NET0131 ,
		_w3372_
	);
	LUT4 #(
		.INIT('hf3f5)
	) name1226 (
		\u7_mem_reg[0][3]/NET0131 ,
		\u7_mem_reg[2][3]/NET0131 ,
		\u7_rp_reg[1]/NET0131 ,
		\u7_rp_reg[2]/NET0131 ,
		_w3373_
	);
	LUT4 #(
		.INIT('ha222)
	) name1227 (
		_w2455_,
		_w2529_,
		_w3372_,
		_w3373_,
		_w3374_
	);
	LUT4 #(
		.INIT('h0b0f)
	) name1228 (
		\u14_u4_en_out_l2_reg/P0001 ,
		\u14_u4_en_out_l_reg/NET0131 ,
		\u7_dout_reg[3]/P0001 ,
		\valid_s_reg/NET0131 ,
		_w3375_
	);
	LUT2 #(
		.INIT('h2)
	) name1229 (
		\u13_occ1_r_reg[0]/NET0131 ,
		_w3375_,
		_w3376_
	);
	LUT3 #(
		.INIT('hb0)
	) name1230 (
		_w3371_,
		_w3374_,
		_w3376_,
		_w3377_
	);
	LUT3 #(
		.INIT('h80)
	) name1231 (
		\u7_rp_reg[0]/P0001 ,
		_w3318_,
		_w3319_,
		_w3378_
	);
	LUT4 #(
		.INIT('h8ccc)
	) name1232 (
		\u7_rp_reg[0]/P0001 ,
		_w2452_,
		_w2527_,
		_w2528_,
		_w3379_
	);
	LUT3 #(
		.INIT('h2a)
	) name1233 (
		_w3227_,
		_w3364_,
		_w3365_,
		_w3380_
	);
	LUT4 #(
		.INIT('hf35f)
	) name1234 (
		\u7_mem_reg[1][4]/NET0131 ,
		\u7_mem_reg[2][4]/NET0131 ,
		\u7_rp_reg[1]/NET0131 ,
		\u7_rp_reg[2]/NET0131 ,
		_w3381_
	);
	LUT4 #(
		.INIT('h3ff5)
	) name1235 (
		\u7_mem_reg[0][4]/NET0131 ,
		\u7_mem_reg[3][4]/NET0131 ,
		\u7_rp_reg[1]/NET0131 ,
		\u7_rp_reg[2]/NET0131 ,
		_w3382_
	);
	LUT4 #(
		.INIT('ha222)
	) name1236 (
		_w2455_,
		_w2529_,
		_w3381_,
		_w3382_,
		_w3383_
	);
	LUT4 #(
		.INIT('h0b00)
	) name1237 (
		_w3378_,
		_w3379_,
		_w3380_,
		_w3383_,
		_w3384_
	);
	LUT4 #(
		.INIT('h0b0f)
	) name1238 (
		\u14_u4_en_out_l2_reg/P0001 ,
		\u14_u4_en_out_l_reg/NET0131 ,
		\u7_dout_reg[4]/P0001 ,
		\valid_s_reg/NET0131 ,
		_w3385_
	);
	LUT2 #(
		.INIT('h2)
	) name1239 (
		\u13_occ1_r_reg[0]/NET0131 ,
		_w3385_,
		_w3386_
	);
	LUT2 #(
		.INIT('h4)
	) name1240 (
		_w3384_,
		_w3386_,
		_w3387_
	);
	LUT3 #(
		.INIT('h80)
	) name1241 (
		\u7_rp_reg[0]/P0001 ,
		_w3331_,
		_w3332_,
		_w3388_
	);
	LUT4 #(
		.INIT('h8ccc)
	) name1242 (
		\u7_rp_reg[0]/P0001 ,
		_w2452_,
		_w2534_,
		_w2535_,
		_w3389_
	);
	LUT3 #(
		.INIT('h2a)
	) name1243 (
		_w3227_,
		_w3372_,
		_w3373_,
		_w3390_
	);
	LUT4 #(
		.INIT('h3ff5)
	) name1244 (
		\u7_mem_reg[0][5]/NET0131 ,
		\u7_mem_reg[3][5]/NET0131 ,
		\u7_rp_reg[1]/NET0131 ,
		\u7_rp_reg[2]/NET0131 ,
		_w3391_
	);
	LUT4 #(
		.INIT('hf35f)
	) name1245 (
		\u7_mem_reg[1][5]/NET0131 ,
		\u7_mem_reg[2][5]/NET0131 ,
		\u7_rp_reg[1]/NET0131 ,
		\u7_rp_reg[2]/NET0131 ,
		_w3392_
	);
	LUT4 #(
		.INIT('ha222)
	) name1246 (
		_w2455_,
		_w2529_,
		_w3391_,
		_w3392_,
		_w3393_
	);
	LUT4 #(
		.INIT('h0b00)
	) name1247 (
		_w3388_,
		_w3389_,
		_w3390_,
		_w3393_,
		_w3394_
	);
	LUT4 #(
		.INIT('h0b0f)
	) name1248 (
		\u14_u4_en_out_l2_reg/P0001 ,
		\u14_u4_en_out_l_reg/NET0131 ,
		\u7_dout_reg[5]/P0001 ,
		\valid_s_reg/NET0131 ,
		_w3395_
	);
	LUT2 #(
		.INIT('h2)
	) name1249 (
		\u13_occ1_r_reg[0]/NET0131 ,
		_w3395_,
		_w3396_
	);
	LUT2 #(
		.INIT('h4)
	) name1250 (
		_w3394_,
		_w3396_,
		_w3397_
	);
	LUT3 #(
		.INIT('h80)
	) name1251 (
		\u7_rp_reg[0]/P0001 ,
		_w3344_,
		_w3345_,
		_w3398_
	);
	LUT4 #(
		.INIT('h8ccc)
	) name1252 (
		\u7_rp_reg[0]/P0001 ,
		_w2452_,
		_w3364_,
		_w3365_,
		_w3399_
	);
	LUT3 #(
		.INIT('h2a)
	) name1253 (
		_w3227_,
		_w3381_,
		_w3382_,
		_w3400_
	);
	LUT4 #(
		.INIT('ha222)
	) name1254 (
		_w2455_,
		_w2529_,
		_w3221_,
		_w3222_,
		_w3401_
	);
	LUT4 #(
		.INIT('h4500)
	) name1255 (
		_w3400_,
		_w3398_,
		_w3399_,
		_w3401_,
		_w3402_
	);
	LUT4 #(
		.INIT('h0b0f)
	) name1256 (
		\u14_u4_en_out_l2_reg/P0001 ,
		\u14_u4_en_out_l_reg/NET0131 ,
		\u7_dout_reg[6]/P0001 ,
		\valid_s_reg/NET0131 ,
		_w3403_
	);
	LUT2 #(
		.INIT('h2)
	) name1257 (
		\u13_occ1_r_reg[0]/NET0131 ,
		_w3403_,
		_w3404_
	);
	LUT2 #(
		.INIT('h4)
	) name1258 (
		_w3402_,
		_w3404_,
		_w3405_
	);
	LUT3 #(
		.INIT('h80)
	) name1259 (
		\u7_rp_reg[0]/P0001 ,
		_w3357_,
		_w3358_,
		_w3406_
	);
	LUT4 #(
		.INIT('h8ccc)
	) name1260 (
		\u7_rp_reg[0]/P0001 ,
		_w2452_,
		_w3372_,
		_w3373_,
		_w3407_
	);
	LUT3 #(
		.INIT('h2a)
	) name1261 (
		_w3227_,
		_w3391_,
		_w3392_,
		_w3408_
	);
	LUT4 #(
		.INIT('ha222)
	) name1262 (
		_w2455_,
		_w2529_,
		_w3245_,
		_w3246_,
		_w3409_
	);
	LUT4 #(
		.INIT('h4500)
	) name1263 (
		_w3408_,
		_w3406_,
		_w3407_,
		_w3409_,
		_w3410_
	);
	LUT4 #(
		.INIT('h0b0f)
	) name1264 (
		\u14_u4_en_out_l2_reg/P0001 ,
		\u14_u4_en_out_l_reg/NET0131 ,
		\u7_dout_reg[7]/P0001 ,
		\valid_s_reg/NET0131 ,
		_w3411_
	);
	LUT2 #(
		.INIT('h2)
	) name1265 (
		\u13_occ1_r_reg[0]/NET0131 ,
		_w3411_,
		_w3412_
	);
	LUT2 #(
		.INIT('h4)
	) name1266 (
		_w3410_,
		_w3412_,
		_w3413_
	);
	LUT4 #(
		.INIT('hc4cc)
	) name1267 (
		\u7_mem_reg[2][20]/NET0131 ,
		\u7_rp_reg[0]/P0001 ,
		\u7_rp_reg[1]/NET0131 ,
		\u7_rp_reg[2]/NET0131 ,
		_w3414_
	);
	LUT3 #(
		.INIT('h02)
	) name1268 (
		\u7_mem_reg[0][20]/NET0131 ,
		\u7_rp_reg[1]/NET0131 ,
		\u7_rp_reg[2]/NET0131 ,
		_w3415_
	);
	LUT4 #(
		.INIT('h3f5f)
	) name1269 (
		\u7_mem_reg[1][20]/NET0131 ,
		\u7_mem_reg[3][20]/NET0131 ,
		\u7_rp_reg[1]/NET0131 ,
		\u7_rp_reg[2]/NET0131 ,
		_w3416_
	);
	LUT3 #(
		.INIT('h40)
	) name1270 (
		_w3415_,
		_w3414_,
		_w3416_,
		_w3417_
	);
	LUT4 #(
		.INIT('h8ccc)
	) name1271 (
		\u7_rp_reg[0]/P0001 ,
		_w2452_,
		_w3381_,
		_w3382_,
		_w3418_
	);
	LUT3 #(
		.INIT('h2a)
	) name1272 (
		_w2529_,
		_w3228_,
		_w3229_,
		_w3419_
	);
	LUT4 #(
		.INIT('h80aa)
	) name1273 (
		_w2455_,
		_w3221_,
		_w3222_,
		_w3227_,
		_w3420_
	);
	LUT4 #(
		.INIT('h4500)
	) name1274 (
		_w3419_,
		_w3417_,
		_w3418_,
		_w3420_,
		_w3421_
	);
	LUT4 #(
		.INIT('h0b0f)
	) name1275 (
		\u14_u4_en_out_l2_reg/P0001 ,
		\u14_u4_en_out_l_reg/NET0131 ,
		\u7_dout_reg[8]/P0001 ,
		\valid_s_reg/NET0131 ,
		_w3422_
	);
	LUT2 #(
		.INIT('h2)
	) name1276 (
		\u13_occ1_r_reg[0]/NET0131 ,
		_w3422_,
		_w3423_
	);
	LUT2 #(
		.INIT('h4)
	) name1277 (
		_w3421_,
		_w3423_,
		_w3424_
	);
	LUT4 #(
		.INIT('hc4cc)
	) name1278 (
		\u7_mem_reg[2][21]/NET0131 ,
		\u7_rp_reg[0]/P0001 ,
		\u7_rp_reg[1]/NET0131 ,
		\u7_rp_reg[2]/NET0131 ,
		_w3425_
	);
	LUT3 #(
		.INIT('h02)
	) name1279 (
		\u7_mem_reg[0][21]/NET0131 ,
		\u7_rp_reg[1]/NET0131 ,
		\u7_rp_reg[2]/NET0131 ,
		_w3426_
	);
	LUT4 #(
		.INIT('h3f5f)
	) name1280 (
		\u7_mem_reg[1][21]/NET0131 ,
		\u7_mem_reg[3][21]/NET0131 ,
		\u7_rp_reg[1]/NET0131 ,
		\u7_rp_reg[2]/NET0131 ,
		_w3427_
	);
	LUT3 #(
		.INIT('h40)
	) name1281 (
		_w3426_,
		_w3425_,
		_w3427_,
		_w3428_
	);
	LUT4 #(
		.INIT('h8ccc)
	) name1282 (
		\u7_rp_reg[0]/P0001 ,
		_w2452_,
		_w3391_,
		_w3392_,
		_w3429_
	);
	LUT3 #(
		.INIT('h2a)
	) name1283 (
		_w2529_,
		_w3242_,
		_w3243_,
		_w3430_
	);
	LUT4 #(
		.INIT('ha222)
	) name1284 (
		_w2455_,
		_w3227_,
		_w3245_,
		_w3246_,
		_w3431_
	);
	LUT4 #(
		.INIT('h4500)
	) name1285 (
		_w3430_,
		_w3428_,
		_w3429_,
		_w3431_,
		_w3432_
	);
	LUT4 #(
		.INIT('h0b0f)
	) name1286 (
		\u14_u4_en_out_l2_reg/P0001 ,
		\u14_u4_en_out_l_reg/NET0131 ,
		\u7_dout_reg[9]/P0001 ,
		\valid_s_reg/NET0131 ,
		_w3433_
	);
	LUT2 #(
		.INIT('h2)
	) name1287 (
		\u13_occ1_r_reg[0]/NET0131 ,
		_w3433_,
		_w3434_
	);
	LUT2 #(
		.INIT('h4)
	) name1288 (
		_w3432_,
		_w3434_,
		_w3435_
	);
	LUT4 #(
		.INIT('hc4cc)
	) name1289 (
		\u3_mem_reg[2][22]/NET0131 ,
		\u3_rp_reg[0]/P0001 ,
		\u3_rp_reg[1]/NET0131 ,
		\u3_rp_reg[2]/NET0131 ,
		_w3436_
	);
	LUT3 #(
		.INIT('h02)
	) name1290 (
		\u3_mem_reg[0][22]/NET0131 ,
		\u3_rp_reg[1]/NET0131 ,
		\u3_rp_reg[2]/NET0131 ,
		_w3437_
	);
	LUT4 #(
		.INIT('h3f5f)
	) name1291 (
		\u3_mem_reg[1][22]/NET0131 ,
		\u3_mem_reg[3][22]/NET0131 ,
		\u3_rp_reg[1]/NET0131 ,
		\u3_rp_reg[2]/NET0131 ,
		_w3438_
	);
	LUT3 #(
		.INIT('h40)
	) name1292 (
		_w3437_,
		_w3436_,
		_w3438_,
		_w3439_
	);
	LUT4 #(
		.INIT('h35ff)
	) name1293 (
		\u3_mem_reg[2][6]/NET0131 ,
		\u3_mem_reg[3][6]/NET0131 ,
		\u3_rp_reg[1]/NET0131 ,
		\u3_rp_reg[2]/NET0131 ,
		_w3440_
	);
	LUT4 #(
		.INIT('hff35)
	) name1294 (
		\u3_mem_reg[0][6]/NET0131 ,
		\u3_mem_reg[1][6]/NET0131 ,
		\u3_rp_reg[1]/NET0131 ,
		\u3_rp_reg[2]/NET0131 ,
		_w3441_
	);
	LUT4 #(
		.INIT('h8ccc)
	) name1295 (
		\u3_rp_reg[0]/P0001 ,
		_w2437_,
		_w3440_,
		_w3441_,
		_w3442_
	);
	LUT2 #(
		.INIT('h2)
	) name1296 (
		\u13_occ0_r_reg[2]/NET0131 ,
		\u13_occ0_r_reg[3]/NET0131 ,
		_w3443_
	);
	LUT4 #(
		.INIT('h35ff)
	) name1297 (
		\u3_mem_reg[2][8]/NET0131 ,
		\u3_mem_reg[3][8]/NET0131 ,
		\u3_rp_reg[1]/NET0131 ,
		\u3_rp_reg[2]/NET0131 ,
		_w3444_
	);
	LUT4 #(
		.INIT('hff35)
	) name1298 (
		\u3_mem_reg[0][8]/NET0131 ,
		\u3_mem_reg[1][8]/NET0131 ,
		\u3_rp_reg[1]/NET0131 ,
		\u3_rp_reg[2]/NET0131 ,
		_w3445_
	);
	LUT3 #(
		.INIT('h2a)
	) name1299 (
		_w3443_,
		_w3444_,
		_w3445_,
		_w3446_
	);
	LUT4 #(
		.INIT('h35ff)
	) name1300 (
		\u3_mem_reg[2][10]/NET0131 ,
		\u3_mem_reg[3][10]/NET0131 ,
		\u3_rp_reg[1]/NET0131 ,
		\u3_rp_reg[2]/NET0131 ,
		_w3447_
	);
	LUT4 #(
		.INIT('hff35)
	) name1301 (
		\u3_mem_reg[0][10]/NET0131 ,
		\u3_mem_reg[1][10]/NET0131 ,
		\u3_rp_reg[1]/NET0131 ,
		\u3_rp_reg[2]/NET0131 ,
		_w3448_
	);
	LUT4 #(
		.INIT('ha222)
	) name1302 (
		_w2439_,
		_w2542_,
		_w3447_,
		_w3448_,
		_w3449_
	);
	LUT4 #(
		.INIT('h0b00)
	) name1303 (
		_w3439_,
		_w3442_,
		_w3446_,
		_w3449_,
		_w3450_
	);
	LUT4 #(
		.INIT('h0b0f)
	) name1304 (
		\u14_u0_en_out_l2_reg/P0001 ,
		\u14_u0_en_out_l_reg/NET0131 ,
		\u3_dout_reg[10]/P0001 ,
		\valid_s_reg/NET0131 ,
		_w3451_
	);
	LUT2 #(
		.INIT('h2)
	) name1305 (
		\u13_occ0_r_reg[0]/NET0131 ,
		_w3451_,
		_w3452_
	);
	LUT2 #(
		.INIT('h4)
	) name1306 (
		_w3450_,
		_w3452_,
		_w3453_
	);
	LUT4 #(
		.INIT('h35ff)
	) name1307 (
		\u3_mem_reg[2][9]/NET0131 ,
		\u3_mem_reg[3][9]/NET0131 ,
		\u3_rp_reg[1]/NET0131 ,
		\u3_rp_reg[2]/NET0131 ,
		_w3454_
	);
	LUT4 #(
		.INIT('hff35)
	) name1308 (
		\u3_mem_reg[0][9]/NET0131 ,
		\u3_mem_reg[1][9]/NET0131 ,
		\u3_rp_reg[1]/NET0131 ,
		\u3_rp_reg[2]/NET0131 ,
		_w3455_
	);
	LUT4 #(
		.INIT('ha222)
	) name1309 (
		_w2439_,
		_w3443_,
		_w3454_,
		_w3455_,
		_w3456_
	);
	LUT3 #(
		.INIT('h10)
	) name1310 (
		\u13_occ0_r_reg[2]/NET0131 ,
		\u13_occ0_r_reg[3]/NET0131 ,
		\u3_rp_reg[0]/P0001 ,
		_w3457_
	);
	LUT4 #(
		.INIT('hf3f5)
	) name1311 (
		\u3_mem_reg[0][23]/NET0131 ,
		\u3_mem_reg[2][23]/NET0131 ,
		\u3_rp_reg[1]/NET0131 ,
		\u3_rp_reg[2]/NET0131 ,
		_w3458_
	);
	LUT4 #(
		.INIT('h3f5f)
	) name1312 (
		\u3_mem_reg[1][23]/NET0131 ,
		\u3_mem_reg[3][23]/NET0131 ,
		\u3_rp_reg[1]/NET0131 ,
		\u3_rp_reg[2]/NET0131 ,
		_w3459_
	);
	LUT3 #(
		.INIT('h2a)
	) name1313 (
		_w3457_,
		_w3458_,
		_w3459_,
		_w3460_
	);
	LUT4 #(
		.INIT('h35ff)
	) name1314 (
		\u3_mem_reg[2][11]/NET0131 ,
		\u3_mem_reg[3][11]/NET0131 ,
		\u3_rp_reg[1]/NET0131 ,
		\u3_rp_reg[2]/NET0131 ,
		_w3461_
	);
	LUT4 #(
		.INIT('hff35)
	) name1315 (
		\u3_mem_reg[0][11]/NET0131 ,
		\u3_mem_reg[1][11]/NET0131 ,
		\u3_rp_reg[1]/NET0131 ,
		\u3_rp_reg[2]/NET0131 ,
		_w3462_
	);
	LUT3 #(
		.INIT('h2a)
	) name1316 (
		_w2542_,
		_w3461_,
		_w3462_,
		_w3463_
	);
	LUT4 #(
		.INIT('hf3f5)
	) name1317 (
		\u3_mem_reg[0][7]/NET0131 ,
		\u3_mem_reg[2][7]/NET0131 ,
		\u3_rp_reg[1]/NET0131 ,
		\u3_rp_reg[2]/NET0131 ,
		_w3464_
	);
	LUT4 #(
		.INIT('h3f5f)
	) name1318 (
		\u3_mem_reg[1][7]/NET0131 ,
		\u3_mem_reg[3][7]/NET0131 ,
		\u3_rp_reg[1]/NET0131 ,
		\u3_rp_reg[2]/NET0131 ,
		_w3465_
	);
	LUT3 #(
		.INIT('h2a)
	) name1319 (
		_w2438_,
		_w3464_,
		_w3465_,
		_w3466_
	);
	LUT4 #(
		.INIT('h0100)
	) name1320 (
		_w3463_,
		_w3466_,
		_w3460_,
		_w3456_,
		_w3467_
	);
	LUT4 #(
		.INIT('h0b0f)
	) name1321 (
		\u14_u0_en_out_l2_reg/P0001 ,
		\u14_u0_en_out_l_reg/NET0131 ,
		\u3_dout_reg[11]/P0001 ,
		\valid_s_reg/NET0131 ,
		_w3468_
	);
	LUT2 #(
		.INIT('h2)
	) name1322 (
		\u13_occ0_r_reg[0]/NET0131 ,
		_w3468_,
		_w3469_
	);
	LUT2 #(
		.INIT('h4)
	) name1323 (
		_w3467_,
		_w3469_,
		_w3470_
	);
	LUT4 #(
		.INIT('hc4cc)
	) name1324 (
		\u3_mem_reg[2][24]/NET0131 ,
		\u3_rp_reg[0]/P0001 ,
		\u3_rp_reg[1]/NET0131 ,
		\u3_rp_reg[2]/NET0131 ,
		_w3471_
	);
	LUT3 #(
		.INIT('h02)
	) name1325 (
		\u3_mem_reg[0][24]/NET0131 ,
		\u3_rp_reg[1]/NET0131 ,
		\u3_rp_reg[2]/NET0131 ,
		_w3472_
	);
	LUT4 #(
		.INIT('h3f5f)
	) name1326 (
		\u3_mem_reg[1][24]/NET0131 ,
		\u3_mem_reg[3][24]/NET0131 ,
		\u3_rp_reg[1]/NET0131 ,
		\u3_rp_reg[2]/NET0131 ,
		_w3473_
	);
	LUT3 #(
		.INIT('h40)
	) name1327 (
		_w3472_,
		_w3471_,
		_w3473_,
		_w3474_
	);
	LUT4 #(
		.INIT('h8ccc)
	) name1328 (
		\u3_rp_reg[0]/P0001 ,
		_w2437_,
		_w3444_,
		_w3445_,
		_w3475_
	);
	LUT3 #(
		.INIT('h70)
	) name1329 (
		_w3447_,
		_w3448_,
		_w3443_,
		_w3476_
	);
	LUT4 #(
		.INIT('h35ff)
	) name1330 (
		\u3_mem_reg[2][12]/NET0131 ,
		\u3_mem_reg[3][12]/NET0131 ,
		\u3_rp_reg[1]/NET0131 ,
		\u3_rp_reg[2]/NET0131 ,
		_w3477_
	);
	LUT4 #(
		.INIT('hff35)
	) name1331 (
		\u3_mem_reg[0][12]/NET0131 ,
		\u3_mem_reg[1][12]/NET0131 ,
		\u3_rp_reg[1]/NET0131 ,
		\u3_rp_reg[2]/NET0131 ,
		_w3478_
	);
	LUT4 #(
		.INIT('ha222)
	) name1332 (
		_w2439_,
		_w2542_,
		_w3477_,
		_w3478_,
		_w3479_
	);
	LUT4 #(
		.INIT('h0b00)
	) name1333 (
		_w3474_,
		_w3475_,
		_w3476_,
		_w3479_,
		_w3480_
	);
	LUT4 #(
		.INIT('h0b0f)
	) name1334 (
		\u14_u0_en_out_l2_reg/P0001 ,
		\u14_u0_en_out_l_reg/NET0131 ,
		\u3_dout_reg[12]/P0001 ,
		\valid_s_reg/NET0131 ,
		_w3481_
	);
	LUT2 #(
		.INIT('h2)
	) name1335 (
		\u13_occ0_r_reg[0]/NET0131 ,
		_w3481_,
		_w3482_
	);
	LUT2 #(
		.INIT('h4)
	) name1336 (
		_w3480_,
		_w3482_,
		_w3483_
	);
	LUT4 #(
		.INIT('hc444)
	) name1337 (
		_w2438_,
		_w2439_,
		_w3454_,
		_w3455_,
		_w3484_
	);
	LUT3 #(
		.INIT('h2a)
	) name1338 (
		_w3443_,
		_w3461_,
		_w3462_,
		_w3485_
	);
	LUT4 #(
		.INIT('h3f5f)
	) name1339 (
		\u3_mem_reg[1][13]/NET0131 ,
		\u3_mem_reg[3][13]/NET0131 ,
		\u3_rp_reg[1]/NET0131 ,
		\u3_rp_reg[2]/NET0131 ,
		_w3486_
	);
	LUT4 #(
		.INIT('hf3f5)
	) name1340 (
		\u3_mem_reg[0][13]/NET0131 ,
		\u3_mem_reg[2][13]/NET0131 ,
		\u3_rp_reg[1]/NET0131 ,
		\u3_rp_reg[2]/NET0131 ,
		_w3487_
	);
	LUT3 #(
		.INIT('h2a)
	) name1341 (
		_w2542_,
		_w3486_,
		_w3487_,
		_w3488_
	);
	LUT4 #(
		.INIT('h3f5f)
	) name1342 (
		\u3_mem_reg[1][25]/NET0131 ,
		\u3_mem_reg[3][25]/NET0131 ,
		\u3_rp_reg[1]/NET0131 ,
		\u3_rp_reg[2]/NET0131 ,
		_w3489_
	);
	LUT4 #(
		.INIT('hf3f5)
	) name1343 (
		\u3_mem_reg[0][25]/NET0131 ,
		\u3_mem_reg[2][25]/NET0131 ,
		\u3_rp_reg[1]/NET0131 ,
		\u3_rp_reg[2]/NET0131 ,
		_w3490_
	);
	LUT3 #(
		.INIT('h2a)
	) name1344 (
		_w3457_,
		_w3489_,
		_w3490_,
		_w3491_
	);
	LUT4 #(
		.INIT('h0100)
	) name1345 (
		_w3488_,
		_w3491_,
		_w3485_,
		_w3484_,
		_w3492_
	);
	LUT4 #(
		.INIT('h0b0f)
	) name1346 (
		\u14_u0_en_out_l2_reg/P0001 ,
		\u14_u0_en_out_l_reg/NET0131 ,
		\u3_dout_reg[13]/P0001 ,
		\valid_s_reg/NET0131 ,
		_w3493_
	);
	LUT2 #(
		.INIT('h2)
	) name1347 (
		\u13_occ0_r_reg[0]/NET0131 ,
		_w3493_,
		_w3494_
	);
	LUT2 #(
		.INIT('h4)
	) name1348 (
		_w3492_,
		_w3494_,
		_w3495_
	);
	LUT4 #(
		.INIT('hc4cc)
	) name1349 (
		\u3_mem_reg[2][26]/NET0131 ,
		\u3_rp_reg[0]/P0001 ,
		\u3_rp_reg[1]/NET0131 ,
		\u3_rp_reg[2]/NET0131 ,
		_w3496_
	);
	LUT3 #(
		.INIT('h02)
	) name1350 (
		\u3_mem_reg[0][26]/NET0131 ,
		\u3_rp_reg[1]/NET0131 ,
		\u3_rp_reg[2]/NET0131 ,
		_w3497_
	);
	LUT4 #(
		.INIT('h3f5f)
	) name1351 (
		\u3_mem_reg[1][26]/NET0131 ,
		\u3_mem_reg[3][26]/NET0131 ,
		\u3_rp_reg[1]/NET0131 ,
		\u3_rp_reg[2]/NET0131 ,
		_w3498_
	);
	LUT3 #(
		.INIT('h40)
	) name1352 (
		_w3497_,
		_w3496_,
		_w3498_,
		_w3499_
	);
	LUT4 #(
		.INIT('h8ccc)
	) name1353 (
		\u3_rp_reg[0]/P0001 ,
		_w2437_,
		_w3447_,
		_w3448_,
		_w3500_
	);
	LUT3 #(
		.INIT('h2a)
	) name1354 (
		_w3443_,
		_w3477_,
		_w3478_,
		_w3501_
	);
	LUT4 #(
		.INIT('h3f5f)
	) name1355 (
		\u3_mem_reg[1][14]/NET0131 ,
		\u3_mem_reg[3][14]/NET0131 ,
		\u3_rp_reg[1]/NET0131 ,
		\u3_rp_reg[2]/NET0131 ,
		_w3502_
	);
	LUT4 #(
		.INIT('hf3f5)
	) name1356 (
		\u3_mem_reg[0][14]/NET0131 ,
		\u3_mem_reg[2][14]/NET0131 ,
		\u3_rp_reg[1]/NET0131 ,
		\u3_rp_reg[2]/NET0131 ,
		_w3503_
	);
	LUT4 #(
		.INIT('ha222)
	) name1357 (
		_w2439_,
		_w2542_,
		_w3502_,
		_w3503_,
		_w3504_
	);
	LUT4 #(
		.INIT('h0b00)
	) name1358 (
		_w3499_,
		_w3500_,
		_w3501_,
		_w3504_,
		_w3505_
	);
	LUT4 #(
		.INIT('h0b0f)
	) name1359 (
		\u14_u0_en_out_l2_reg/P0001 ,
		\u14_u0_en_out_l_reg/NET0131 ,
		\u3_dout_reg[14]/P0001 ,
		\valid_s_reg/NET0131 ,
		_w3506_
	);
	LUT2 #(
		.INIT('h2)
	) name1360 (
		\u13_occ0_r_reg[0]/NET0131 ,
		_w3506_,
		_w3507_
	);
	LUT2 #(
		.INIT('h4)
	) name1361 (
		_w3505_,
		_w3507_,
		_w3508_
	);
	LUT4 #(
		.INIT('hc4cc)
	) name1362 (
		\u3_mem_reg[2][27]/NET0131 ,
		\u3_rp_reg[0]/P0001 ,
		\u3_rp_reg[1]/NET0131 ,
		\u3_rp_reg[2]/NET0131 ,
		_w3509_
	);
	LUT3 #(
		.INIT('h02)
	) name1363 (
		\u3_mem_reg[0][27]/NET0131 ,
		\u3_rp_reg[1]/NET0131 ,
		\u3_rp_reg[2]/NET0131 ,
		_w3510_
	);
	LUT4 #(
		.INIT('h3f5f)
	) name1364 (
		\u3_mem_reg[1][27]/NET0131 ,
		\u3_mem_reg[3][27]/NET0131 ,
		\u3_rp_reg[1]/NET0131 ,
		\u3_rp_reg[2]/NET0131 ,
		_w3511_
	);
	LUT3 #(
		.INIT('h40)
	) name1365 (
		_w3510_,
		_w3509_,
		_w3511_,
		_w3512_
	);
	LUT4 #(
		.INIT('h8ccc)
	) name1366 (
		\u3_rp_reg[0]/P0001 ,
		_w2437_,
		_w3461_,
		_w3462_,
		_w3513_
	);
	LUT4 #(
		.INIT('h35ff)
	) name1367 (
		\u3_mem_reg[2][15]/NET0131 ,
		\u3_mem_reg[3][15]/NET0131 ,
		\u3_rp_reg[1]/NET0131 ,
		\u3_rp_reg[2]/NET0131 ,
		_w3514_
	);
	LUT4 #(
		.INIT('hff35)
	) name1368 (
		\u3_mem_reg[0][15]/NET0131 ,
		\u3_mem_reg[1][15]/NET0131 ,
		\u3_rp_reg[1]/NET0131 ,
		\u3_rp_reg[2]/NET0131 ,
		_w3515_
	);
	LUT3 #(
		.INIT('h2a)
	) name1369 (
		_w2542_,
		_w3514_,
		_w3515_,
		_w3516_
	);
	LUT4 #(
		.INIT('ha222)
	) name1370 (
		_w2439_,
		_w3443_,
		_w3486_,
		_w3487_,
		_w3517_
	);
	LUT4 #(
		.INIT('h4500)
	) name1371 (
		_w3516_,
		_w3512_,
		_w3513_,
		_w3517_,
		_w3518_
	);
	LUT4 #(
		.INIT('h0b0f)
	) name1372 (
		\u14_u0_en_out_l2_reg/P0001 ,
		\u14_u0_en_out_l_reg/NET0131 ,
		\u3_dout_reg[15]/P0001 ,
		\valid_s_reg/NET0131 ,
		_w3519_
	);
	LUT2 #(
		.INIT('h2)
	) name1373 (
		\u13_occ0_r_reg[0]/NET0131 ,
		_w3519_,
		_w3520_
	);
	LUT2 #(
		.INIT('h4)
	) name1374 (
		_w3518_,
		_w3520_,
		_w3521_
	);
	LUT4 #(
		.INIT('hc4cc)
	) name1375 (
		\u3_mem_reg[2][28]/NET0131 ,
		\u3_rp_reg[0]/P0001 ,
		\u3_rp_reg[1]/NET0131 ,
		\u3_rp_reg[2]/NET0131 ,
		_w3522_
	);
	LUT3 #(
		.INIT('h02)
	) name1376 (
		\u3_mem_reg[0][28]/NET0131 ,
		\u3_rp_reg[1]/NET0131 ,
		\u3_rp_reg[2]/NET0131 ,
		_w3523_
	);
	LUT4 #(
		.INIT('h3f5f)
	) name1377 (
		\u3_mem_reg[1][28]/NET0131 ,
		\u3_mem_reg[3][28]/NET0131 ,
		\u3_rp_reg[1]/NET0131 ,
		\u3_rp_reg[2]/NET0131 ,
		_w3524_
	);
	LUT3 #(
		.INIT('h40)
	) name1378 (
		_w3523_,
		_w3522_,
		_w3524_,
		_w3525_
	);
	LUT4 #(
		.INIT('h8ccc)
	) name1379 (
		\u3_rp_reg[0]/P0001 ,
		_w2437_,
		_w3477_,
		_w3478_,
		_w3526_
	);
	LUT3 #(
		.INIT('h2a)
	) name1380 (
		_w3443_,
		_w3502_,
		_w3503_,
		_w3527_
	);
	LUT4 #(
		.INIT('h35ff)
	) name1381 (
		\u3_mem_reg[2][16]/NET0131 ,
		\u3_mem_reg[3][16]/NET0131 ,
		\u3_rp_reg[1]/NET0131 ,
		\u3_rp_reg[2]/NET0131 ,
		_w3528_
	);
	LUT4 #(
		.INIT('hff35)
	) name1382 (
		\u3_mem_reg[0][16]/NET0131 ,
		\u3_mem_reg[1][16]/NET0131 ,
		\u3_rp_reg[1]/NET0131 ,
		\u3_rp_reg[2]/NET0131 ,
		_w3529_
	);
	LUT4 #(
		.INIT('ha222)
	) name1383 (
		_w2439_,
		_w2542_,
		_w3528_,
		_w3529_,
		_w3530_
	);
	LUT4 #(
		.INIT('h0b00)
	) name1384 (
		_w3525_,
		_w3526_,
		_w3527_,
		_w3530_,
		_w3531_
	);
	LUT4 #(
		.INIT('h0b0f)
	) name1385 (
		\u14_u0_en_out_l2_reg/P0001 ,
		\u14_u0_en_out_l_reg/NET0131 ,
		\u3_dout_reg[16]/P0001 ,
		\valid_s_reg/NET0131 ,
		_w3532_
	);
	LUT2 #(
		.INIT('h2)
	) name1386 (
		\u13_occ0_r_reg[0]/NET0131 ,
		_w3532_,
		_w3533_
	);
	LUT2 #(
		.INIT('h4)
	) name1387 (
		_w3531_,
		_w3533_,
		_w3534_
	);
	LUT4 #(
		.INIT('ha222)
	) name1388 (
		_w2439_,
		_w3443_,
		_w3514_,
		_w3515_,
		_w3535_
	);
	LUT4 #(
		.INIT('h3f5f)
	) name1389 (
		\u3_mem_reg[1][17]/NET0131 ,
		\u3_mem_reg[3][17]/NET0131 ,
		\u3_rp_reg[1]/NET0131 ,
		\u3_rp_reg[2]/NET0131 ,
		_w3536_
	);
	LUT4 #(
		.INIT('hf3f5)
	) name1390 (
		\u3_mem_reg[0][17]/NET0131 ,
		\u3_mem_reg[2][17]/NET0131 ,
		\u3_rp_reg[1]/NET0131 ,
		\u3_rp_reg[2]/NET0131 ,
		_w3537_
	);
	LUT3 #(
		.INIT('h2a)
	) name1391 (
		_w2542_,
		_w3536_,
		_w3537_,
		_w3538_
	);
	LUT3 #(
		.INIT('h2a)
	) name1392 (
		_w2438_,
		_w3486_,
		_w3487_,
		_w3539_
	);
	LUT4 #(
		.INIT('h3ff5)
	) name1393 (
		\u3_mem_reg[0][29]/NET0131 ,
		\u3_mem_reg[3][29]/NET0131 ,
		\u3_rp_reg[1]/NET0131 ,
		\u3_rp_reg[2]/NET0131 ,
		_w3540_
	);
	LUT4 #(
		.INIT('hf35f)
	) name1394 (
		\u3_mem_reg[1][29]/NET0131 ,
		\u3_mem_reg[2][29]/NET0131 ,
		\u3_rp_reg[1]/NET0131 ,
		\u3_rp_reg[2]/NET0131 ,
		_w3541_
	);
	LUT3 #(
		.INIT('h2a)
	) name1395 (
		_w3457_,
		_w3540_,
		_w3541_,
		_w3542_
	);
	LUT4 #(
		.INIT('h0100)
	) name1396 (
		_w3539_,
		_w3542_,
		_w3538_,
		_w3535_,
		_w3543_
	);
	LUT4 #(
		.INIT('h0b0f)
	) name1397 (
		\u14_u0_en_out_l2_reg/P0001 ,
		\u14_u0_en_out_l_reg/NET0131 ,
		\u3_dout_reg[17]/P0001 ,
		\valid_s_reg/NET0131 ,
		_w3544_
	);
	LUT2 #(
		.INIT('h2)
	) name1398 (
		\u13_occ0_r_reg[0]/NET0131 ,
		_w3544_,
		_w3545_
	);
	LUT2 #(
		.INIT('h4)
	) name1399 (
		_w3543_,
		_w3545_,
		_w3546_
	);
	LUT4 #(
		.INIT('hc4cc)
	) name1400 (
		\u3_mem_reg[2][30]/NET0131 ,
		\u3_rp_reg[0]/P0001 ,
		\u3_rp_reg[1]/NET0131 ,
		\u3_rp_reg[2]/NET0131 ,
		_w3547_
	);
	LUT3 #(
		.INIT('h02)
	) name1401 (
		\u3_mem_reg[0][30]/NET0131 ,
		\u3_rp_reg[1]/NET0131 ,
		\u3_rp_reg[2]/NET0131 ,
		_w3548_
	);
	LUT4 #(
		.INIT('h3f5f)
	) name1402 (
		\u3_mem_reg[1][30]/NET0131 ,
		\u3_mem_reg[3][30]/NET0131 ,
		\u3_rp_reg[1]/NET0131 ,
		\u3_rp_reg[2]/NET0131 ,
		_w3549_
	);
	LUT3 #(
		.INIT('h40)
	) name1403 (
		_w3548_,
		_w3547_,
		_w3549_,
		_w3550_
	);
	LUT4 #(
		.INIT('h8ccc)
	) name1404 (
		\u3_rp_reg[0]/P0001 ,
		_w2437_,
		_w3502_,
		_w3503_,
		_w3551_
	);
	LUT3 #(
		.INIT('h2a)
	) name1405 (
		_w3443_,
		_w3528_,
		_w3529_,
		_w3552_
	);
	LUT4 #(
		.INIT('h3f5f)
	) name1406 (
		\u3_mem_reg[1][18]/NET0131 ,
		\u3_mem_reg[3][18]/NET0131 ,
		\u3_rp_reg[1]/NET0131 ,
		\u3_rp_reg[2]/NET0131 ,
		_w3553_
	);
	LUT4 #(
		.INIT('hf3f5)
	) name1407 (
		\u3_mem_reg[0][18]/NET0131 ,
		\u3_mem_reg[2][18]/NET0131 ,
		\u3_rp_reg[1]/NET0131 ,
		\u3_rp_reg[2]/NET0131 ,
		_w3554_
	);
	LUT4 #(
		.INIT('ha222)
	) name1408 (
		_w2439_,
		_w2542_,
		_w3553_,
		_w3554_,
		_w3555_
	);
	LUT4 #(
		.INIT('h0b00)
	) name1409 (
		_w3550_,
		_w3551_,
		_w3552_,
		_w3555_,
		_w3556_
	);
	LUT4 #(
		.INIT('h0b0f)
	) name1410 (
		\u14_u0_en_out_l2_reg/P0001 ,
		\u14_u0_en_out_l_reg/NET0131 ,
		\u3_dout_reg[18]/P0001 ,
		\valid_s_reg/NET0131 ,
		_w3557_
	);
	LUT2 #(
		.INIT('h2)
	) name1411 (
		\u13_occ0_r_reg[0]/NET0131 ,
		_w3557_,
		_w3558_
	);
	LUT2 #(
		.INIT('h4)
	) name1412 (
		_w3556_,
		_w3558_,
		_w3559_
	);
	LUT4 #(
		.INIT('hc4cc)
	) name1413 (
		\u8_mem_reg[2][22]/NET0131 ,
		\u8_rp_reg[0]/P0001 ,
		\u8_rp_reg[1]/NET0131 ,
		\u8_rp_reg[2]/NET0131 ,
		_w3560_
	);
	LUT3 #(
		.INIT('h02)
	) name1414 (
		\u8_mem_reg[0][22]/NET0131 ,
		\u8_rp_reg[1]/NET0131 ,
		\u8_rp_reg[2]/NET0131 ,
		_w3561_
	);
	LUT4 #(
		.INIT('h3f5f)
	) name1415 (
		\u8_mem_reg[1][22]/NET0131 ,
		\u8_mem_reg[3][22]/NET0131 ,
		\u8_rp_reg[1]/NET0131 ,
		\u8_rp_reg[2]/NET0131 ,
		_w3562_
	);
	LUT3 #(
		.INIT('h40)
	) name1416 (
		_w3561_,
		_w3560_,
		_w3562_,
		_w3563_
	);
	LUT4 #(
		.INIT('h35ff)
	) name1417 (
		\u8_mem_reg[2][6]/NET0131 ,
		\u8_mem_reg[3][6]/NET0131 ,
		\u8_rp_reg[1]/NET0131 ,
		\u8_rp_reg[2]/NET0131 ,
		_w3564_
	);
	LUT4 #(
		.INIT('hff35)
	) name1418 (
		\u8_mem_reg[0][6]/NET0131 ,
		\u8_mem_reg[1][6]/NET0131 ,
		\u8_rp_reg[1]/NET0131 ,
		\u8_rp_reg[2]/NET0131 ,
		_w3565_
	);
	LUT4 #(
		.INIT('h8ccc)
	) name1419 (
		\u8_rp_reg[0]/P0001 ,
		_w2156_,
		_w3564_,
		_w3565_,
		_w3566_
	);
	LUT2 #(
		.INIT('h2)
	) name1420 (
		\u13_occ1_r_reg[10]/NET0131 ,
		\u13_occ1_r_reg[11]/NET0131 ,
		_w3567_
	);
	LUT4 #(
		.INIT('h35ff)
	) name1421 (
		\u8_mem_reg[2][8]/NET0131 ,
		\u8_mem_reg[3][8]/NET0131 ,
		\u8_rp_reg[1]/NET0131 ,
		\u8_rp_reg[2]/NET0131 ,
		_w3568_
	);
	LUT4 #(
		.INIT('hff35)
	) name1422 (
		\u8_mem_reg[0][8]/NET0131 ,
		\u8_mem_reg[1][8]/NET0131 ,
		\u8_rp_reg[1]/NET0131 ,
		\u8_rp_reg[2]/NET0131 ,
		_w3569_
	);
	LUT3 #(
		.INIT('h2a)
	) name1423 (
		_w3567_,
		_w3568_,
		_w3569_,
		_w3570_
	);
	LUT4 #(
		.INIT('h35ff)
	) name1424 (
		\u8_mem_reg[2][10]/NET0131 ,
		\u8_mem_reg[3][10]/NET0131 ,
		\u8_rp_reg[1]/NET0131 ,
		\u8_rp_reg[2]/NET0131 ,
		_w3571_
	);
	LUT4 #(
		.INIT('hff35)
	) name1425 (
		\u8_mem_reg[0][10]/NET0131 ,
		\u8_mem_reg[1][10]/NET0131 ,
		\u8_rp_reg[1]/NET0131 ,
		\u8_rp_reg[2]/NET0131 ,
		_w3572_
	);
	LUT4 #(
		.INIT('ha222)
	) name1426 (
		_w2155_,
		_w2550_,
		_w3571_,
		_w3572_,
		_w3573_
	);
	LUT4 #(
		.INIT('h0b00)
	) name1427 (
		_w3563_,
		_w3566_,
		_w3570_,
		_w3573_,
		_w3574_
	);
	LUT4 #(
		.INIT('h0b0f)
	) name1428 (
		\u14_u5_en_out_l2_reg/P0001 ,
		\u14_u5_en_out_l_reg/NET0131 ,
		\u8_dout_reg[10]/P0001 ,
		\valid_s_reg/NET0131 ,
		_w3575_
	);
	LUT2 #(
		.INIT('h2)
	) name1429 (
		\u13_occ1_r_reg[8]/NET0131 ,
		_w3575_,
		_w3576_
	);
	LUT2 #(
		.INIT('h4)
	) name1430 (
		_w3574_,
		_w3576_,
		_w3577_
	);
	LUT4 #(
		.INIT('hc4cc)
	) name1431 (
		\u3_mem_reg[2][31]/NET0131 ,
		\u3_rp_reg[0]/P0001 ,
		\u3_rp_reg[1]/NET0131 ,
		\u3_rp_reg[2]/NET0131 ,
		_w3578_
	);
	LUT3 #(
		.INIT('h02)
	) name1432 (
		\u3_mem_reg[0][31]/NET0131 ,
		\u3_rp_reg[1]/NET0131 ,
		\u3_rp_reg[2]/NET0131 ,
		_w3579_
	);
	LUT4 #(
		.INIT('h3f5f)
	) name1433 (
		\u3_mem_reg[1][31]/NET0131 ,
		\u3_mem_reg[3][31]/NET0131 ,
		\u3_rp_reg[1]/NET0131 ,
		\u3_rp_reg[2]/NET0131 ,
		_w3580_
	);
	LUT3 #(
		.INIT('h40)
	) name1434 (
		_w3579_,
		_w3578_,
		_w3580_,
		_w3581_
	);
	LUT4 #(
		.INIT('h8ccc)
	) name1435 (
		\u3_rp_reg[0]/P0001 ,
		_w2437_,
		_w3514_,
		_w3515_,
		_w3582_
	);
	LUT3 #(
		.INIT('h2a)
	) name1436 (
		_w3443_,
		_w3536_,
		_w3537_,
		_w3583_
	);
	LUT4 #(
		.INIT('hf3f5)
	) name1437 (
		\u3_mem_reg[0][19]/NET0131 ,
		\u3_mem_reg[2][19]/NET0131 ,
		\u3_rp_reg[1]/NET0131 ,
		\u3_rp_reg[2]/NET0131 ,
		_w3584_
	);
	LUT4 #(
		.INIT('h3f5f)
	) name1438 (
		\u3_mem_reg[1][19]/NET0131 ,
		\u3_mem_reg[3][19]/NET0131 ,
		\u3_rp_reg[1]/NET0131 ,
		\u3_rp_reg[2]/NET0131 ,
		_w3585_
	);
	LUT4 #(
		.INIT('ha222)
	) name1439 (
		_w2439_,
		_w2542_,
		_w3584_,
		_w3585_,
		_w3586_
	);
	LUT4 #(
		.INIT('h0b00)
	) name1440 (
		_w3581_,
		_w3582_,
		_w3583_,
		_w3586_,
		_w3587_
	);
	LUT4 #(
		.INIT('h0b0f)
	) name1441 (
		\u14_u0_en_out_l2_reg/P0001 ,
		\u14_u0_en_out_l_reg/NET0131 ,
		\u3_dout_reg[19]/P0001 ,
		\valid_s_reg/NET0131 ,
		_w3588_
	);
	LUT2 #(
		.INIT('h2)
	) name1442 (
		\u13_occ0_r_reg[0]/NET0131 ,
		_w3588_,
		_w3589_
	);
	LUT2 #(
		.INIT('h4)
	) name1443 (
		_w3587_,
		_w3589_,
		_w3590_
	);
	LUT4 #(
		.INIT('hc4cc)
	) name1444 (
		\u8_mem_reg[2][23]/NET0131 ,
		\u8_rp_reg[0]/P0001 ,
		\u8_rp_reg[1]/NET0131 ,
		\u8_rp_reg[2]/NET0131 ,
		_w3591_
	);
	LUT3 #(
		.INIT('h02)
	) name1445 (
		\u8_mem_reg[0][23]/NET0131 ,
		\u8_rp_reg[1]/NET0131 ,
		\u8_rp_reg[2]/NET0131 ,
		_w3592_
	);
	LUT4 #(
		.INIT('h3f5f)
	) name1446 (
		\u8_mem_reg[1][23]/NET0131 ,
		\u8_mem_reg[3][23]/NET0131 ,
		\u8_rp_reg[1]/NET0131 ,
		\u8_rp_reg[2]/NET0131 ,
		_w3593_
	);
	LUT3 #(
		.INIT('h40)
	) name1447 (
		_w3592_,
		_w3591_,
		_w3593_,
		_w3594_
	);
	LUT4 #(
		.INIT('h35ff)
	) name1448 (
		\u8_mem_reg[2][7]/NET0131 ,
		\u8_mem_reg[3][7]/NET0131 ,
		\u8_rp_reg[1]/NET0131 ,
		\u8_rp_reg[2]/NET0131 ,
		_w3595_
	);
	LUT4 #(
		.INIT('hff35)
	) name1449 (
		\u8_mem_reg[0][7]/NET0131 ,
		\u8_mem_reg[1][7]/NET0131 ,
		\u8_rp_reg[1]/NET0131 ,
		\u8_rp_reg[2]/NET0131 ,
		_w3596_
	);
	LUT4 #(
		.INIT('h8ccc)
	) name1450 (
		\u8_rp_reg[0]/P0001 ,
		_w2156_,
		_w3595_,
		_w3596_,
		_w3597_
	);
	LUT4 #(
		.INIT('h3f5f)
	) name1451 (
		\u8_mem_reg[1][9]/NET0131 ,
		\u8_mem_reg[3][9]/NET0131 ,
		\u8_rp_reg[1]/NET0131 ,
		\u8_rp_reg[2]/NET0131 ,
		_w3598_
	);
	LUT4 #(
		.INIT('hf3f5)
	) name1452 (
		\u8_mem_reg[0][9]/NET0131 ,
		\u8_mem_reg[2][9]/NET0131 ,
		\u8_rp_reg[1]/NET0131 ,
		\u8_rp_reg[2]/NET0131 ,
		_w3599_
	);
	LUT3 #(
		.INIT('h2a)
	) name1453 (
		_w3567_,
		_w3598_,
		_w3599_,
		_w3600_
	);
	LUT4 #(
		.INIT('h35ff)
	) name1454 (
		\u8_mem_reg[2][11]/NET0131 ,
		\u8_mem_reg[3][11]/NET0131 ,
		\u8_rp_reg[1]/NET0131 ,
		\u8_rp_reg[2]/NET0131 ,
		_w3601_
	);
	LUT4 #(
		.INIT('hff35)
	) name1455 (
		\u8_mem_reg[0][11]/NET0131 ,
		\u8_mem_reg[1][11]/NET0131 ,
		\u8_rp_reg[1]/NET0131 ,
		\u8_rp_reg[2]/NET0131 ,
		_w3602_
	);
	LUT4 #(
		.INIT('ha222)
	) name1456 (
		_w2155_,
		_w2550_,
		_w3601_,
		_w3602_,
		_w3603_
	);
	LUT4 #(
		.INIT('h0b00)
	) name1457 (
		_w3594_,
		_w3597_,
		_w3600_,
		_w3603_,
		_w3604_
	);
	LUT4 #(
		.INIT('h0b0f)
	) name1458 (
		\u14_u5_en_out_l2_reg/P0001 ,
		\u14_u5_en_out_l_reg/NET0131 ,
		\u8_dout_reg[11]/P0001 ,
		\valid_s_reg/NET0131 ,
		_w3605_
	);
	LUT2 #(
		.INIT('h2)
	) name1459 (
		\u13_occ1_r_reg[8]/NET0131 ,
		_w3605_,
		_w3606_
	);
	LUT2 #(
		.INIT('h4)
	) name1460 (
		_w3604_,
		_w3606_,
		_w3607_
	);
	LUT4 #(
		.INIT('hc4cc)
	) name1461 (
		\u8_mem_reg[2][24]/NET0131 ,
		\u8_rp_reg[0]/P0001 ,
		\u8_rp_reg[1]/NET0131 ,
		\u8_rp_reg[2]/NET0131 ,
		_w3608_
	);
	LUT3 #(
		.INIT('h02)
	) name1462 (
		\u8_mem_reg[0][24]/NET0131 ,
		\u8_rp_reg[1]/NET0131 ,
		\u8_rp_reg[2]/NET0131 ,
		_w3609_
	);
	LUT4 #(
		.INIT('h3f5f)
	) name1463 (
		\u8_mem_reg[1][24]/NET0131 ,
		\u8_mem_reg[3][24]/NET0131 ,
		\u8_rp_reg[1]/NET0131 ,
		\u8_rp_reg[2]/NET0131 ,
		_w3610_
	);
	LUT3 #(
		.INIT('h40)
	) name1464 (
		_w3609_,
		_w3608_,
		_w3610_,
		_w3611_
	);
	LUT4 #(
		.INIT('h8ccc)
	) name1465 (
		\u8_rp_reg[0]/P0001 ,
		_w2156_,
		_w3568_,
		_w3569_,
		_w3612_
	);
	LUT3 #(
		.INIT('h70)
	) name1466 (
		_w3571_,
		_w3572_,
		_w3567_,
		_w3613_
	);
	LUT4 #(
		.INIT('h3f5f)
	) name1467 (
		\u8_mem_reg[1][12]/NET0131 ,
		\u8_mem_reg[3][12]/NET0131 ,
		\u8_rp_reg[1]/NET0131 ,
		\u8_rp_reg[2]/NET0131 ,
		_w3614_
	);
	LUT4 #(
		.INIT('hf3f5)
	) name1468 (
		\u8_mem_reg[0][12]/NET0131 ,
		\u8_mem_reg[2][12]/NET0131 ,
		\u8_rp_reg[1]/NET0131 ,
		\u8_rp_reg[2]/NET0131 ,
		_w3615_
	);
	LUT4 #(
		.INIT('ha222)
	) name1469 (
		_w2155_,
		_w2550_,
		_w3614_,
		_w3615_,
		_w3616_
	);
	LUT4 #(
		.INIT('h0b00)
	) name1470 (
		_w3611_,
		_w3612_,
		_w3613_,
		_w3616_,
		_w3617_
	);
	LUT4 #(
		.INIT('h0b0f)
	) name1471 (
		\u14_u5_en_out_l2_reg/P0001 ,
		\u14_u5_en_out_l_reg/NET0131 ,
		\u8_dout_reg[12]/P0001 ,
		\valid_s_reg/NET0131 ,
		_w3618_
	);
	LUT2 #(
		.INIT('h2)
	) name1472 (
		\u13_occ1_r_reg[8]/NET0131 ,
		_w3618_,
		_w3619_
	);
	LUT2 #(
		.INIT('h4)
	) name1473 (
		_w3617_,
		_w3619_,
		_w3620_
	);
	LUT4 #(
		.INIT('h35ff)
	) name1474 (
		\u3_mem_reg[2][2]/NET0131 ,
		\u3_mem_reg[3][2]/NET0131 ,
		\u3_rp_reg[1]/NET0131 ,
		\u3_rp_reg[2]/NET0131 ,
		_w3621_
	);
	LUT4 #(
		.INIT('hff35)
	) name1475 (
		\u3_mem_reg[0][2]/NET0131 ,
		\u3_mem_reg[1][2]/NET0131 ,
		\u3_rp_reg[1]/NET0131 ,
		\u3_rp_reg[2]/NET0131 ,
		_w3622_
	);
	LUT3 #(
		.INIT('h2a)
	) name1476 (
		_w2542_,
		_w3621_,
		_w3622_,
		_w3623_
	);
	LUT4 #(
		.INIT('h80aa)
	) name1477 (
		_w2439_,
		_w2540_,
		_w2541_,
		_w3443_,
		_w3624_
	);
	LUT4 #(
		.INIT('h0b0f)
	) name1478 (
		\u14_u0_en_out_l2_reg/P0001 ,
		\u14_u0_en_out_l_reg/NET0131 ,
		\u3_dout_reg[2]/P0001 ,
		\valid_s_reg/NET0131 ,
		_w3625_
	);
	LUT2 #(
		.INIT('h2)
	) name1479 (
		\u13_occ0_r_reg[0]/NET0131 ,
		_w3625_,
		_w3626_
	);
	LUT3 #(
		.INIT('hb0)
	) name1480 (
		_w3623_,
		_w3624_,
		_w3626_,
		_w3627_
	);
	LUT4 #(
		.INIT('hc4cc)
	) name1481 (
		\u8_mem_reg[2][25]/NET0131 ,
		\u8_rp_reg[0]/P0001 ,
		\u8_rp_reg[1]/NET0131 ,
		\u8_rp_reg[2]/NET0131 ,
		_w3628_
	);
	LUT3 #(
		.INIT('h02)
	) name1482 (
		\u8_mem_reg[0][25]/NET0131 ,
		\u8_rp_reg[1]/NET0131 ,
		\u8_rp_reg[2]/NET0131 ,
		_w3629_
	);
	LUT4 #(
		.INIT('h3f5f)
	) name1483 (
		\u8_mem_reg[1][25]/NET0131 ,
		\u8_mem_reg[3][25]/NET0131 ,
		\u8_rp_reg[1]/NET0131 ,
		\u8_rp_reg[2]/NET0131 ,
		_w3630_
	);
	LUT3 #(
		.INIT('h40)
	) name1484 (
		_w3629_,
		_w3628_,
		_w3630_,
		_w3631_
	);
	LUT4 #(
		.INIT('h8ccc)
	) name1485 (
		\u8_rp_reg[0]/P0001 ,
		_w2156_,
		_w3598_,
		_w3599_,
		_w3632_
	);
	LUT3 #(
		.INIT('h2a)
	) name1486 (
		_w3567_,
		_w3601_,
		_w3602_,
		_w3633_
	);
	LUT4 #(
		.INIT('h35ff)
	) name1487 (
		\u8_mem_reg[2][13]/NET0131 ,
		\u8_mem_reg[3][13]/NET0131 ,
		\u8_rp_reg[1]/NET0131 ,
		\u8_rp_reg[2]/NET0131 ,
		_w3634_
	);
	LUT4 #(
		.INIT('hff35)
	) name1488 (
		\u8_mem_reg[0][13]/NET0131 ,
		\u8_mem_reg[1][13]/NET0131 ,
		\u8_rp_reg[1]/NET0131 ,
		\u8_rp_reg[2]/NET0131 ,
		_w3635_
	);
	LUT4 #(
		.INIT('ha222)
	) name1489 (
		_w2155_,
		_w2550_,
		_w3634_,
		_w3635_,
		_w3636_
	);
	LUT4 #(
		.INIT('h0b00)
	) name1490 (
		_w3631_,
		_w3632_,
		_w3633_,
		_w3636_,
		_w3637_
	);
	LUT4 #(
		.INIT('h0b0f)
	) name1491 (
		\u14_u5_en_out_l2_reg/P0001 ,
		\u14_u5_en_out_l_reg/NET0131 ,
		\u8_dout_reg[13]/P0001 ,
		\valid_s_reg/NET0131 ,
		_w3638_
	);
	LUT2 #(
		.INIT('h2)
	) name1492 (
		\u13_occ1_r_reg[8]/NET0131 ,
		_w3638_,
		_w3639_
	);
	LUT2 #(
		.INIT('h4)
	) name1493 (
		_w3637_,
		_w3639_,
		_w3640_
	);
	LUT4 #(
		.INIT('h3f5f)
	) name1494 (
		\u3_mem_reg[1][3]/NET0131 ,
		\u3_mem_reg[3][3]/NET0131 ,
		\u3_rp_reg[1]/NET0131 ,
		\u3_rp_reg[2]/NET0131 ,
		_w3641_
	);
	LUT4 #(
		.INIT('hf3f5)
	) name1495 (
		\u3_mem_reg[0][3]/NET0131 ,
		\u3_mem_reg[2][3]/NET0131 ,
		\u3_rp_reg[1]/NET0131 ,
		\u3_rp_reg[2]/NET0131 ,
		_w3642_
	);
	LUT3 #(
		.INIT('h2a)
	) name1496 (
		_w2542_,
		_w3641_,
		_w3642_,
		_w3643_
	);
	LUT4 #(
		.INIT('h80aa)
	) name1497 (
		_w2439_,
		_w2555_,
		_w2556_,
		_w3443_,
		_w3644_
	);
	LUT4 #(
		.INIT('h0b0f)
	) name1498 (
		\u14_u0_en_out_l2_reg/P0001 ,
		\u14_u0_en_out_l_reg/NET0131 ,
		\u3_dout_reg[3]/P0001 ,
		\valid_s_reg/NET0131 ,
		_w3645_
	);
	LUT2 #(
		.INIT('h2)
	) name1499 (
		\u13_occ0_r_reg[0]/NET0131 ,
		_w3645_,
		_w3646_
	);
	LUT3 #(
		.INIT('hb0)
	) name1500 (
		_w3643_,
		_w3644_,
		_w3646_,
		_w3647_
	);
	LUT4 #(
		.INIT('hc4cc)
	) name1501 (
		\u8_mem_reg[2][26]/NET0131 ,
		\u8_rp_reg[0]/P0001 ,
		\u8_rp_reg[1]/NET0131 ,
		\u8_rp_reg[2]/NET0131 ,
		_w3648_
	);
	LUT3 #(
		.INIT('h02)
	) name1502 (
		\u8_mem_reg[0][26]/NET0131 ,
		\u8_rp_reg[1]/NET0131 ,
		\u8_rp_reg[2]/NET0131 ,
		_w3649_
	);
	LUT4 #(
		.INIT('h3f5f)
	) name1503 (
		\u8_mem_reg[1][26]/NET0131 ,
		\u8_mem_reg[3][26]/NET0131 ,
		\u8_rp_reg[1]/NET0131 ,
		\u8_rp_reg[2]/NET0131 ,
		_w3650_
	);
	LUT3 #(
		.INIT('h40)
	) name1504 (
		_w3649_,
		_w3648_,
		_w3650_,
		_w3651_
	);
	LUT4 #(
		.INIT('h8ccc)
	) name1505 (
		\u8_rp_reg[0]/P0001 ,
		_w2156_,
		_w3571_,
		_w3572_,
		_w3652_
	);
	LUT3 #(
		.INIT('h2a)
	) name1506 (
		_w3567_,
		_w3614_,
		_w3615_,
		_w3653_
	);
	LUT4 #(
		.INIT('h35ff)
	) name1507 (
		\u8_mem_reg[2][14]/NET0131 ,
		\u8_mem_reg[3][14]/NET0131 ,
		\u8_rp_reg[1]/NET0131 ,
		\u8_rp_reg[2]/NET0131 ,
		_w3654_
	);
	LUT4 #(
		.INIT('hff35)
	) name1508 (
		\u8_mem_reg[0][14]/NET0131 ,
		\u8_mem_reg[1][14]/NET0131 ,
		\u8_rp_reg[1]/NET0131 ,
		\u8_rp_reg[2]/NET0131 ,
		_w3655_
	);
	LUT4 #(
		.INIT('ha222)
	) name1509 (
		_w2155_,
		_w2550_,
		_w3654_,
		_w3655_,
		_w3656_
	);
	LUT4 #(
		.INIT('h0b00)
	) name1510 (
		_w3651_,
		_w3652_,
		_w3653_,
		_w3656_,
		_w3657_
	);
	LUT4 #(
		.INIT('h0b0f)
	) name1511 (
		\u14_u5_en_out_l2_reg/P0001 ,
		\u14_u5_en_out_l_reg/NET0131 ,
		\u8_dout_reg[14]/P0001 ,
		\valid_s_reg/NET0131 ,
		_w3658_
	);
	LUT2 #(
		.INIT('h2)
	) name1512 (
		\u13_occ1_r_reg[8]/NET0131 ,
		_w3658_,
		_w3659_
	);
	LUT2 #(
		.INIT('h4)
	) name1513 (
		_w3657_,
		_w3659_,
		_w3660_
	);
	LUT3 #(
		.INIT('h80)
	) name1514 (
		\u3_rp_reg[0]/P0001 ,
		_w3528_,
		_w3529_,
		_w3661_
	);
	LUT4 #(
		.INIT('h8ccc)
	) name1515 (
		\u3_rp_reg[0]/P0001 ,
		_w2437_,
		_w2540_,
		_w2541_,
		_w3662_
	);
	LUT3 #(
		.INIT('h2a)
	) name1516 (
		_w3443_,
		_w3621_,
		_w3622_,
		_w3663_
	);
	LUT4 #(
		.INIT('h35ff)
	) name1517 (
		\u3_mem_reg[2][4]/NET0131 ,
		\u3_mem_reg[3][4]/NET0131 ,
		\u3_rp_reg[1]/NET0131 ,
		\u3_rp_reg[2]/NET0131 ,
		_w3664_
	);
	LUT4 #(
		.INIT('hff35)
	) name1518 (
		\u3_mem_reg[0][4]/NET0131 ,
		\u3_mem_reg[1][4]/NET0131 ,
		\u3_rp_reg[1]/NET0131 ,
		\u3_rp_reg[2]/NET0131 ,
		_w3665_
	);
	LUT4 #(
		.INIT('ha222)
	) name1519 (
		_w2439_,
		_w2542_,
		_w3664_,
		_w3665_,
		_w3666_
	);
	LUT4 #(
		.INIT('h0b00)
	) name1520 (
		_w3661_,
		_w3662_,
		_w3663_,
		_w3666_,
		_w3667_
	);
	LUT4 #(
		.INIT('h0b0f)
	) name1521 (
		\u14_u0_en_out_l2_reg/P0001 ,
		\u14_u0_en_out_l_reg/NET0131 ,
		\u3_dout_reg[4]/P0001 ,
		\valid_s_reg/NET0131 ,
		_w3668_
	);
	LUT2 #(
		.INIT('h2)
	) name1522 (
		\u13_occ0_r_reg[0]/NET0131 ,
		_w3668_,
		_w3669_
	);
	LUT2 #(
		.INIT('h4)
	) name1523 (
		_w3667_,
		_w3669_,
		_w3670_
	);
	LUT4 #(
		.INIT('hc4cc)
	) name1524 (
		\u8_mem_reg[2][27]/NET0131 ,
		\u8_rp_reg[0]/P0001 ,
		\u8_rp_reg[1]/NET0131 ,
		\u8_rp_reg[2]/NET0131 ,
		_w3671_
	);
	LUT3 #(
		.INIT('h02)
	) name1525 (
		\u8_mem_reg[0][27]/NET0131 ,
		\u8_rp_reg[1]/NET0131 ,
		\u8_rp_reg[2]/NET0131 ,
		_w3672_
	);
	LUT4 #(
		.INIT('h3f5f)
	) name1526 (
		\u8_mem_reg[1][27]/NET0131 ,
		\u8_mem_reg[3][27]/NET0131 ,
		\u8_rp_reg[1]/NET0131 ,
		\u8_rp_reg[2]/NET0131 ,
		_w3673_
	);
	LUT3 #(
		.INIT('h40)
	) name1527 (
		_w3672_,
		_w3671_,
		_w3673_,
		_w3674_
	);
	LUT4 #(
		.INIT('h8ccc)
	) name1528 (
		\u8_rp_reg[0]/P0001 ,
		_w2156_,
		_w3601_,
		_w3602_,
		_w3675_
	);
	LUT3 #(
		.INIT('h2a)
	) name1529 (
		_w3567_,
		_w3634_,
		_w3635_,
		_w3676_
	);
	LUT4 #(
		.INIT('h35ff)
	) name1530 (
		\u8_mem_reg[2][15]/NET0131 ,
		\u8_mem_reg[3][15]/NET0131 ,
		\u8_rp_reg[1]/NET0131 ,
		\u8_rp_reg[2]/NET0131 ,
		_w3677_
	);
	LUT4 #(
		.INIT('hff35)
	) name1531 (
		\u8_mem_reg[0][15]/NET0131 ,
		\u8_mem_reg[1][15]/NET0131 ,
		\u8_rp_reg[1]/NET0131 ,
		\u8_rp_reg[2]/NET0131 ,
		_w3678_
	);
	LUT4 #(
		.INIT('ha222)
	) name1532 (
		_w2155_,
		_w2550_,
		_w3677_,
		_w3678_,
		_w3679_
	);
	LUT4 #(
		.INIT('h0b00)
	) name1533 (
		_w3674_,
		_w3675_,
		_w3676_,
		_w3679_,
		_w3680_
	);
	LUT4 #(
		.INIT('h0b0f)
	) name1534 (
		\u14_u5_en_out_l2_reg/P0001 ,
		\u14_u5_en_out_l_reg/NET0131 ,
		\u8_dout_reg[15]/P0001 ,
		\valid_s_reg/NET0131 ,
		_w3681_
	);
	LUT2 #(
		.INIT('h2)
	) name1535 (
		\u13_occ1_r_reg[8]/NET0131 ,
		_w3681_,
		_w3682_
	);
	LUT2 #(
		.INIT('h4)
	) name1536 (
		_w3680_,
		_w3682_,
		_w3683_
	);
	LUT3 #(
		.INIT('h80)
	) name1537 (
		\u3_rp_reg[0]/P0001 ,
		_w3536_,
		_w3537_,
		_w3684_
	);
	LUT4 #(
		.INIT('h8ccc)
	) name1538 (
		\u3_rp_reg[0]/P0001 ,
		_w2437_,
		_w2555_,
		_w2556_,
		_w3685_
	);
	LUT3 #(
		.INIT('h2a)
	) name1539 (
		_w3443_,
		_w3641_,
		_w3642_,
		_w3686_
	);
	LUT4 #(
		.INIT('h35ff)
	) name1540 (
		\u3_mem_reg[2][5]/NET0131 ,
		\u3_mem_reg[3][5]/NET0131 ,
		\u3_rp_reg[1]/NET0131 ,
		\u3_rp_reg[2]/NET0131 ,
		_w3687_
	);
	LUT4 #(
		.INIT('hff35)
	) name1541 (
		\u3_mem_reg[0][5]/NET0131 ,
		\u3_mem_reg[1][5]/NET0131 ,
		\u3_rp_reg[1]/NET0131 ,
		\u3_rp_reg[2]/NET0131 ,
		_w3688_
	);
	LUT4 #(
		.INIT('ha222)
	) name1542 (
		_w2439_,
		_w2542_,
		_w3687_,
		_w3688_,
		_w3689_
	);
	LUT4 #(
		.INIT('h0b00)
	) name1543 (
		_w3684_,
		_w3685_,
		_w3686_,
		_w3689_,
		_w3690_
	);
	LUT4 #(
		.INIT('h0b0f)
	) name1544 (
		\u14_u0_en_out_l2_reg/P0001 ,
		\u14_u0_en_out_l_reg/NET0131 ,
		\u3_dout_reg[5]/P0001 ,
		\valid_s_reg/NET0131 ,
		_w3691_
	);
	LUT2 #(
		.INIT('h2)
	) name1545 (
		\u13_occ0_r_reg[0]/NET0131 ,
		_w3691_,
		_w3692_
	);
	LUT2 #(
		.INIT('h4)
	) name1546 (
		_w3690_,
		_w3692_,
		_w3693_
	);
	LUT4 #(
		.INIT('hc4cc)
	) name1547 (
		\u8_mem_reg[2][28]/NET0131 ,
		\u8_rp_reg[0]/P0001 ,
		\u8_rp_reg[1]/NET0131 ,
		\u8_rp_reg[2]/NET0131 ,
		_w3694_
	);
	LUT3 #(
		.INIT('h02)
	) name1548 (
		\u8_mem_reg[0][28]/NET0131 ,
		\u8_rp_reg[1]/NET0131 ,
		\u8_rp_reg[2]/NET0131 ,
		_w3695_
	);
	LUT4 #(
		.INIT('h3f5f)
	) name1549 (
		\u8_mem_reg[1][28]/NET0131 ,
		\u8_mem_reg[3][28]/NET0131 ,
		\u8_rp_reg[1]/NET0131 ,
		\u8_rp_reg[2]/NET0131 ,
		_w3696_
	);
	LUT3 #(
		.INIT('h40)
	) name1550 (
		_w3695_,
		_w3694_,
		_w3696_,
		_w3697_
	);
	LUT4 #(
		.INIT('h8ccc)
	) name1551 (
		\u8_rp_reg[0]/P0001 ,
		_w2156_,
		_w3614_,
		_w3615_,
		_w3698_
	);
	LUT3 #(
		.INIT('h2a)
	) name1552 (
		_w3567_,
		_w3654_,
		_w3655_,
		_w3699_
	);
	LUT4 #(
		.INIT('hf3f5)
	) name1553 (
		\u8_mem_reg[0][16]/NET0131 ,
		\u8_mem_reg[2][16]/NET0131 ,
		\u8_rp_reg[1]/NET0131 ,
		\u8_rp_reg[2]/NET0131 ,
		_w3700_
	);
	LUT4 #(
		.INIT('h3f5f)
	) name1554 (
		\u8_mem_reg[1][16]/NET0131 ,
		\u8_mem_reg[3][16]/NET0131 ,
		\u8_rp_reg[1]/NET0131 ,
		\u8_rp_reg[2]/NET0131 ,
		_w3701_
	);
	LUT4 #(
		.INIT('ha222)
	) name1555 (
		_w2155_,
		_w2550_,
		_w3700_,
		_w3701_,
		_w3702_
	);
	LUT4 #(
		.INIT('h0b00)
	) name1556 (
		_w3697_,
		_w3698_,
		_w3699_,
		_w3702_,
		_w3703_
	);
	LUT4 #(
		.INIT('h0b0f)
	) name1557 (
		\u14_u5_en_out_l2_reg/P0001 ,
		\u14_u5_en_out_l_reg/NET0131 ,
		\u8_dout_reg[16]/P0001 ,
		\valid_s_reg/NET0131 ,
		_w3704_
	);
	LUT2 #(
		.INIT('h2)
	) name1558 (
		\u13_occ1_r_reg[8]/NET0131 ,
		_w3704_,
		_w3705_
	);
	LUT2 #(
		.INIT('h4)
	) name1559 (
		_w3703_,
		_w3705_,
		_w3706_
	);
	LUT4 #(
		.INIT('hc4cc)
	) name1560 (
		\u8_mem_reg[2][29]/NET0131 ,
		\u8_rp_reg[0]/P0001 ,
		\u8_rp_reg[1]/NET0131 ,
		\u8_rp_reg[2]/NET0131 ,
		_w3707_
	);
	LUT3 #(
		.INIT('h02)
	) name1561 (
		\u8_mem_reg[0][29]/NET0131 ,
		\u8_rp_reg[1]/NET0131 ,
		\u8_rp_reg[2]/NET0131 ,
		_w3708_
	);
	LUT4 #(
		.INIT('h3f5f)
	) name1562 (
		\u8_mem_reg[1][29]/NET0131 ,
		\u8_mem_reg[3][29]/NET0131 ,
		\u8_rp_reg[1]/NET0131 ,
		\u8_rp_reg[2]/NET0131 ,
		_w3709_
	);
	LUT3 #(
		.INIT('h40)
	) name1563 (
		_w3708_,
		_w3707_,
		_w3709_,
		_w3710_
	);
	LUT4 #(
		.INIT('h8ccc)
	) name1564 (
		\u8_rp_reg[0]/P0001 ,
		_w2156_,
		_w3634_,
		_w3635_,
		_w3711_
	);
	LUT3 #(
		.INIT('h2a)
	) name1565 (
		_w3567_,
		_w3677_,
		_w3678_,
		_w3712_
	);
	LUT4 #(
		.INIT('h35ff)
	) name1566 (
		\u8_mem_reg[2][17]/NET0131 ,
		\u8_mem_reg[3][17]/NET0131 ,
		\u8_rp_reg[1]/NET0131 ,
		\u8_rp_reg[2]/NET0131 ,
		_w3713_
	);
	LUT4 #(
		.INIT('hff35)
	) name1567 (
		\u8_mem_reg[0][17]/NET0131 ,
		\u8_mem_reg[1][17]/NET0131 ,
		\u8_rp_reg[1]/NET0131 ,
		\u8_rp_reg[2]/NET0131 ,
		_w3714_
	);
	LUT4 #(
		.INIT('ha222)
	) name1568 (
		_w2155_,
		_w2550_,
		_w3713_,
		_w3714_,
		_w3715_
	);
	LUT4 #(
		.INIT('h0b00)
	) name1569 (
		_w3710_,
		_w3711_,
		_w3712_,
		_w3715_,
		_w3716_
	);
	LUT4 #(
		.INIT('h0b0f)
	) name1570 (
		\u14_u5_en_out_l2_reg/P0001 ,
		\u14_u5_en_out_l_reg/NET0131 ,
		\u8_dout_reg[17]/P0001 ,
		\valid_s_reg/NET0131 ,
		_w3717_
	);
	LUT2 #(
		.INIT('h2)
	) name1571 (
		\u13_occ1_r_reg[8]/NET0131 ,
		_w3717_,
		_w3718_
	);
	LUT2 #(
		.INIT('h4)
	) name1572 (
		_w3716_,
		_w3718_,
		_w3719_
	);
	LUT3 #(
		.INIT('h80)
	) name1573 (
		\u3_rp_reg[0]/P0001 ,
		_w3553_,
		_w3554_,
		_w3720_
	);
	LUT4 #(
		.INIT('h8ccc)
	) name1574 (
		\u3_rp_reg[0]/P0001 ,
		_w2437_,
		_w3621_,
		_w3622_,
		_w3721_
	);
	LUT3 #(
		.INIT('h2a)
	) name1575 (
		_w3443_,
		_w3664_,
		_w3665_,
		_w3722_
	);
	LUT4 #(
		.INIT('ha222)
	) name1576 (
		_w2439_,
		_w2542_,
		_w3440_,
		_w3441_,
		_w3723_
	);
	LUT4 #(
		.INIT('h0b00)
	) name1577 (
		_w3720_,
		_w3721_,
		_w3722_,
		_w3723_,
		_w3724_
	);
	LUT4 #(
		.INIT('h0b0f)
	) name1578 (
		\u14_u0_en_out_l2_reg/P0001 ,
		\u14_u0_en_out_l_reg/NET0131 ,
		\u3_dout_reg[6]/P0001 ,
		\valid_s_reg/NET0131 ,
		_w3725_
	);
	LUT2 #(
		.INIT('h2)
	) name1579 (
		\u13_occ0_r_reg[0]/NET0131 ,
		_w3725_,
		_w3726_
	);
	LUT2 #(
		.INIT('h4)
	) name1580 (
		_w3724_,
		_w3726_,
		_w3727_
	);
	LUT3 #(
		.INIT('h80)
	) name1581 (
		\u3_rp_reg[0]/P0001 ,
		_w3584_,
		_w3585_,
		_w3728_
	);
	LUT4 #(
		.INIT('h8ccc)
	) name1582 (
		\u3_rp_reg[0]/P0001 ,
		_w2437_,
		_w3641_,
		_w3642_,
		_w3729_
	);
	LUT3 #(
		.INIT('h2a)
	) name1583 (
		_w3443_,
		_w3687_,
		_w3688_,
		_w3730_
	);
	LUT4 #(
		.INIT('ha222)
	) name1584 (
		_w2439_,
		_w2542_,
		_w3464_,
		_w3465_,
		_w3731_
	);
	LUT4 #(
		.INIT('h0b00)
	) name1585 (
		_w3728_,
		_w3729_,
		_w3730_,
		_w3731_,
		_w3732_
	);
	LUT4 #(
		.INIT('h0b0f)
	) name1586 (
		\u14_u0_en_out_l2_reg/P0001 ,
		\u14_u0_en_out_l_reg/NET0131 ,
		\u3_dout_reg[7]/P0001 ,
		\valid_s_reg/NET0131 ,
		_w3733_
	);
	LUT2 #(
		.INIT('h2)
	) name1587 (
		\u13_occ0_r_reg[0]/NET0131 ,
		_w3733_,
		_w3734_
	);
	LUT2 #(
		.INIT('h4)
	) name1588 (
		_w3732_,
		_w3734_,
		_w3735_
	);
	LUT4 #(
		.INIT('hc4cc)
	) name1589 (
		\u8_mem_reg[2][30]/NET0131 ,
		\u8_rp_reg[0]/P0001 ,
		\u8_rp_reg[1]/NET0131 ,
		\u8_rp_reg[2]/NET0131 ,
		_w3736_
	);
	LUT3 #(
		.INIT('h02)
	) name1590 (
		\u8_mem_reg[0][30]/NET0131 ,
		\u8_rp_reg[1]/NET0131 ,
		\u8_rp_reg[2]/NET0131 ,
		_w3737_
	);
	LUT4 #(
		.INIT('h3f5f)
	) name1591 (
		\u8_mem_reg[1][30]/NET0131 ,
		\u8_mem_reg[3][30]/NET0131 ,
		\u8_rp_reg[1]/NET0131 ,
		\u8_rp_reg[2]/NET0131 ,
		_w3738_
	);
	LUT3 #(
		.INIT('h40)
	) name1592 (
		_w3737_,
		_w3736_,
		_w3738_,
		_w3739_
	);
	LUT4 #(
		.INIT('h8ccc)
	) name1593 (
		\u8_rp_reg[0]/P0001 ,
		_w2156_,
		_w3654_,
		_w3655_,
		_w3740_
	);
	LUT3 #(
		.INIT('h2a)
	) name1594 (
		_w3567_,
		_w3700_,
		_w3701_,
		_w3741_
	);
	LUT4 #(
		.INIT('h35ff)
	) name1595 (
		\u8_mem_reg[2][18]/NET0131 ,
		\u8_mem_reg[3][18]/NET0131 ,
		\u8_rp_reg[1]/NET0131 ,
		\u8_rp_reg[2]/NET0131 ,
		_w3742_
	);
	LUT4 #(
		.INIT('hff35)
	) name1596 (
		\u8_mem_reg[0][18]/NET0131 ,
		\u8_mem_reg[1][18]/NET0131 ,
		\u8_rp_reg[1]/NET0131 ,
		\u8_rp_reg[2]/NET0131 ,
		_w3743_
	);
	LUT4 #(
		.INIT('ha222)
	) name1597 (
		_w2155_,
		_w2550_,
		_w3742_,
		_w3743_,
		_w3744_
	);
	LUT4 #(
		.INIT('h0b00)
	) name1598 (
		_w3739_,
		_w3740_,
		_w3741_,
		_w3744_,
		_w3745_
	);
	LUT4 #(
		.INIT('h0b0f)
	) name1599 (
		\u14_u5_en_out_l2_reg/P0001 ,
		\u14_u5_en_out_l_reg/NET0131 ,
		\u8_dout_reg[18]/P0001 ,
		\valid_s_reg/NET0131 ,
		_w3746_
	);
	LUT2 #(
		.INIT('h2)
	) name1600 (
		\u13_occ1_r_reg[8]/NET0131 ,
		_w3746_,
		_w3747_
	);
	LUT2 #(
		.INIT('h4)
	) name1601 (
		_w3745_,
		_w3747_,
		_w3748_
	);
	LUT4 #(
		.INIT('hc4cc)
	) name1602 (
		\u3_mem_reg[2][20]/NET0131 ,
		\u3_rp_reg[0]/P0001 ,
		\u3_rp_reg[1]/NET0131 ,
		\u3_rp_reg[2]/NET0131 ,
		_w3749_
	);
	LUT3 #(
		.INIT('h02)
	) name1603 (
		\u3_mem_reg[0][20]/NET0131 ,
		\u3_rp_reg[1]/NET0131 ,
		\u3_rp_reg[2]/NET0131 ,
		_w3750_
	);
	LUT4 #(
		.INIT('h3f5f)
	) name1604 (
		\u3_mem_reg[1][20]/NET0131 ,
		\u3_mem_reg[3][20]/NET0131 ,
		\u3_rp_reg[1]/NET0131 ,
		\u3_rp_reg[2]/NET0131 ,
		_w3751_
	);
	LUT3 #(
		.INIT('h40)
	) name1605 (
		_w3750_,
		_w3749_,
		_w3751_,
		_w3752_
	);
	LUT4 #(
		.INIT('h8ccc)
	) name1606 (
		\u3_rp_reg[0]/P0001 ,
		_w2437_,
		_w3664_,
		_w3665_,
		_w3753_
	);
	LUT3 #(
		.INIT('h70)
	) name1607 (
		_w3440_,
		_w3441_,
		_w3443_,
		_w3754_
	);
	LUT4 #(
		.INIT('ha222)
	) name1608 (
		_w2439_,
		_w2542_,
		_w3444_,
		_w3445_,
		_w3755_
	);
	LUT4 #(
		.INIT('h0b00)
	) name1609 (
		_w3752_,
		_w3753_,
		_w3754_,
		_w3755_,
		_w3756_
	);
	LUT4 #(
		.INIT('h0b0f)
	) name1610 (
		\u14_u0_en_out_l2_reg/P0001 ,
		\u14_u0_en_out_l_reg/NET0131 ,
		\u3_dout_reg[8]/P0001 ,
		\valid_s_reg/NET0131 ,
		_w3757_
	);
	LUT2 #(
		.INIT('h2)
	) name1611 (
		\u13_occ0_r_reg[0]/NET0131 ,
		_w3757_,
		_w3758_
	);
	LUT2 #(
		.INIT('h4)
	) name1612 (
		_w3756_,
		_w3758_,
		_w3759_
	);
	LUT4 #(
		.INIT('hc4cc)
	) name1613 (
		\u8_mem_reg[2][31]/NET0131 ,
		\u8_rp_reg[0]/P0001 ,
		\u8_rp_reg[1]/NET0131 ,
		\u8_rp_reg[2]/NET0131 ,
		_w3760_
	);
	LUT3 #(
		.INIT('h02)
	) name1614 (
		\u8_mem_reg[0][31]/NET0131 ,
		\u8_rp_reg[1]/NET0131 ,
		\u8_rp_reg[2]/NET0131 ,
		_w3761_
	);
	LUT4 #(
		.INIT('h3f5f)
	) name1615 (
		\u8_mem_reg[1][31]/NET0131 ,
		\u8_mem_reg[3][31]/NET0131 ,
		\u8_rp_reg[1]/NET0131 ,
		\u8_rp_reg[2]/NET0131 ,
		_w3762_
	);
	LUT3 #(
		.INIT('h40)
	) name1616 (
		_w3761_,
		_w3760_,
		_w3762_,
		_w3763_
	);
	LUT4 #(
		.INIT('h8ccc)
	) name1617 (
		\u8_rp_reg[0]/P0001 ,
		_w2156_,
		_w3677_,
		_w3678_,
		_w3764_
	);
	LUT3 #(
		.INIT('h2a)
	) name1618 (
		_w3567_,
		_w3713_,
		_w3714_,
		_w3765_
	);
	LUT4 #(
		.INIT('h3f5f)
	) name1619 (
		\u8_mem_reg[1][19]/NET0131 ,
		\u8_mem_reg[3][19]/NET0131 ,
		\u8_rp_reg[1]/NET0131 ,
		\u8_rp_reg[2]/NET0131 ,
		_w3766_
	);
	LUT4 #(
		.INIT('hf3f5)
	) name1620 (
		\u8_mem_reg[0][19]/NET0131 ,
		\u8_mem_reg[2][19]/NET0131 ,
		\u8_rp_reg[1]/NET0131 ,
		\u8_rp_reg[2]/NET0131 ,
		_w3767_
	);
	LUT4 #(
		.INIT('ha222)
	) name1621 (
		_w2155_,
		_w2550_,
		_w3766_,
		_w3767_,
		_w3768_
	);
	LUT4 #(
		.INIT('h0b00)
	) name1622 (
		_w3763_,
		_w3764_,
		_w3765_,
		_w3768_,
		_w3769_
	);
	LUT4 #(
		.INIT('h0b0f)
	) name1623 (
		\u14_u5_en_out_l2_reg/P0001 ,
		\u14_u5_en_out_l_reg/NET0131 ,
		\u8_dout_reg[19]/P0001 ,
		\valid_s_reg/NET0131 ,
		_w3770_
	);
	LUT2 #(
		.INIT('h2)
	) name1624 (
		\u13_occ1_r_reg[8]/NET0131 ,
		_w3770_,
		_w3771_
	);
	LUT2 #(
		.INIT('h4)
	) name1625 (
		_w3769_,
		_w3771_,
		_w3772_
	);
	LUT4 #(
		.INIT('hc4cc)
	) name1626 (
		\u3_mem_reg[2][21]/NET0131 ,
		\u3_rp_reg[0]/P0001 ,
		\u3_rp_reg[1]/NET0131 ,
		\u3_rp_reg[2]/NET0131 ,
		_w3773_
	);
	LUT3 #(
		.INIT('h02)
	) name1627 (
		\u3_mem_reg[0][21]/NET0131 ,
		\u3_rp_reg[1]/NET0131 ,
		\u3_rp_reg[2]/NET0131 ,
		_w3774_
	);
	LUT4 #(
		.INIT('h3f5f)
	) name1628 (
		\u3_mem_reg[1][21]/NET0131 ,
		\u3_mem_reg[3][21]/NET0131 ,
		\u3_rp_reg[1]/NET0131 ,
		\u3_rp_reg[2]/NET0131 ,
		_w3775_
	);
	LUT3 #(
		.INIT('h40)
	) name1629 (
		_w3774_,
		_w3773_,
		_w3775_,
		_w3776_
	);
	LUT4 #(
		.INIT('h8ccc)
	) name1630 (
		\u3_rp_reg[0]/P0001 ,
		_w2437_,
		_w3687_,
		_w3688_,
		_w3777_
	);
	LUT3 #(
		.INIT('h2a)
	) name1631 (
		_w3443_,
		_w3464_,
		_w3465_,
		_w3778_
	);
	LUT4 #(
		.INIT('ha222)
	) name1632 (
		_w2439_,
		_w2542_,
		_w3454_,
		_w3455_,
		_w3779_
	);
	LUT4 #(
		.INIT('h4500)
	) name1633 (
		_w3778_,
		_w3776_,
		_w3777_,
		_w3779_,
		_w3780_
	);
	LUT4 #(
		.INIT('h0b0f)
	) name1634 (
		\u14_u0_en_out_l2_reg/P0001 ,
		\u14_u0_en_out_l_reg/NET0131 ,
		\u3_dout_reg[9]/P0001 ,
		\valid_s_reg/NET0131 ,
		_w3781_
	);
	LUT2 #(
		.INIT('h2)
	) name1635 (
		\u13_occ0_r_reg[0]/NET0131 ,
		_w3781_,
		_w3782_
	);
	LUT2 #(
		.INIT('h4)
	) name1636 (
		_w3780_,
		_w3782_,
		_w3783_
	);
	LUT4 #(
		.INIT('h3ff5)
	) name1637 (
		\u8_mem_reg[0][2]/NET0131 ,
		\u8_mem_reg[3][2]/NET0131 ,
		\u8_rp_reg[1]/NET0131 ,
		\u8_rp_reg[2]/NET0131 ,
		_w3784_
	);
	LUT4 #(
		.INIT('hf35f)
	) name1638 (
		\u8_mem_reg[1][2]/NET0131 ,
		\u8_mem_reg[2][2]/NET0131 ,
		\u8_rp_reg[1]/NET0131 ,
		\u8_rp_reg[2]/NET0131 ,
		_w3785_
	);
	LUT3 #(
		.INIT('h2a)
	) name1639 (
		_w2550_,
		_w3784_,
		_w3785_,
		_w3786_
	);
	LUT4 #(
		.INIT('h80aa)
	) name1640 (
		_w2155_,
		_w2548_,
		_w2549_,
		_w3567_,
		_w3787_
	);
	LUT4 #(
		.INIT('h0b0f)
	) name1641 (
		\u14_u5_en_out_l2_reg/P0001 ,
		\u14_u5_en_out_l_reg/NET0131 ,
		\u8_dout_reg[2]/P0001 ,
		\valid_s_reg/NET0131 ,
		_w3788_
	);
	LUT2 #(
		.INIT('h2)
	) name1642 (
		\u13_occ1_r_reg[8]/NET0131 ,
		_w3788_,
		_w3789_
	);
	LUT3 #(
		.INIT('hb0)
	) name1643 (
		_w3786_,
		_w3787_,
		_w3789_,
		_w3790_
	);
	LUT4 #(
		.INIT('h3ff5)
	) name1644 (
		\u8_mem_reg[0][3]/NET0131 ,
		\u8_mem_reg[3][3]/NET0131 ,
		\u8_rp_reg[1]/NET0131 ,
		\u8_rp_reg[2]/NET0131 ,
		_w3791_
	);
	LUT4 #(
		.INIT('hf35f)
	) name1645 (
		\u8_mem_reg[1][3]/NET0131 ,
		\u8_mem_reg[2][3]/NET0131 ,
		\u8_rp_reg[1]/NET0131 ,
		\u8_rp_reg[2]/NET0131 ,
		_w3792_
	);
	LUT3 #(
		.INIT('h2a)
	) name1646 (
		_w2550_,
		_w3791_,
		_w3792_,
		_w3793_
	);
	LUT4 #(
		.INIT('h80aa)
	) name1647 (
		_w2155_,
		_w2560_,
		_w2561_,
		_w3567_,
		_w3794_
	);
	LUT4 #(
		.INIT('h0b0f)
	) name1648 (
		\u14_u5_en_out_l2_reg/P0001 ,
		\u14_u5_en_out_l_reg/NET0131 ,
		\u8_dout_reg[3]/P0001 ,
		\valid_s_reg/NET0131 ,
		_w3795_
	);
	LUT2 #(
		.INIT('h2)
	) name1649 (
		\u13_occ1_r_reg[8]/NET0131 ,
		_w3795_,
		_w3796_
	);
	LUT3 #(
		.INIT('hb0)
	) name1650 (
		_w3793_,
		_w3794_,
		_w3796_,
		_w3797_
	);
	LUT3 #(
		.INIT('h80)
	) name1651 (
		\u8_rp_reg[0]/P0001 ,
		_w3700_,
		_w3701_,
		_w3798_
	);
	LUT4 #(
		.INIT('h8ccc)
	) name1652 (
		\u8_rp_reg[0]/P0001 ,
		_w2156_,
		_w2548_,
		_w2549_,
		_w3799_
	);
	LUT3 #(
		.INIT('h2a)
	) name1653 (
		_w3567_,
		_w3784_,
		_w3785_,
		_w3800_
	);
	LUT4 #(
		.INIT('h35ff)
	) name1654 (
		\u8_mem_reg[2][4]/NET0131 ,
		\u8_mem_reg[3][4]/NET0131 ,
		\u8_rp_reg[1]/NET0131 ,
		\u8_rp_reg[2]/NET0131 ,
		_w3801_
	);
	LUT4 #(
		.INIT('hff35)
	) name1655 (
		\u8_mem_reg[0][4]/NET0131 ,
		\u8_mem_reg[1][4]/NET0131 ,
		\u8_rp_reg[1]/NET0131 ,
		\u8_rp_reg[2]/NET0131 ,
		_w3802_
	);
	LUT4 #(
		.INIT('ha222)
	) name1656 (
		_w2155_,
		_w2550_,
		_w3801_,
		_w3802_,
		_w3803_
	);
	LUT4 #(
		.INIT('h0b00)
	) name1657 (
		_w3798_,
		_w3799_,
		_w3800_,
		_w3803_,
		_w3804_
	);
	LUT4 #(
		.INIT('h0b0f)
	) name1658 (
		\u14_u5_en_out_l2_reg/P0001 ,
		\u14_u5_en_out_l_reg/NET0131 ,
		\u8_dout_reg[4]/P0001 ,
		\valid_s_reg/NET0131 ,
		_w3805_
	);
	LUT2 #(
		.INIT('h2)
	) name1659 (
		\u13_occ1_r_reg[8]/NET0131 ,
		_w3805_,
		_w3806_
	);
	LUT2 #(
		.INIT('h4)
	) name1660 (
		_w3804_,
		_w3806_,
		_w3807_
	);
	LUT3 #(
		.INIT('h80)
	) name1661 (
		\u8_rp_reg[0]/P0001 ,
		_w3713_,
		_w3714_,
		_w3808_
	);
	LUT4 #(
		.INIT('h8ccc)
	) name1662 (
		\u8_rp_reg[0]/P0001 ,
		_w2156_,
		_w2560_,
		_w2561_,
		_w3809_
	);
	LUT3 #(
		.INIT('h2a)
	) name1663 (
		_w3567_,
		_w3791_,
		_w3792_,
		_w3810_
	);
	LUT4 #(
		.INIT('h35ff)
	) name1664 (
		\u8_mem_reg[2][5]/NET0131 ,
		\u8_mem_reg[3][5]/NET0131 ,
		\u8_rp_reg[1]/NET0131 ,
		\u8_rp_reg[2]/NET0131 ,
		_w3811_
	);
	LUT4 #(
		.INIT('hff35)
	) name1665 (
		\u8_mem_reg[0][5]/NET0131 ,
		\u8_mem_reg[1][5]/NET0131 ,
		\u8_rp_reg[1]/NET0131 ,
		\u8_rp_reg[2]/NET0131 ,
		_w3812_
	);
	LUT4 #(
		.INIT('ha222)
	) name1666 (
		_w2155_,
		_w2550_,
		_w3811_,
		_w3812_,
		_w3813_
	);
	LUT4 #(
		.INIT('h0b00)
	) name1667 (
		_w3808_,
		_w3809_,
		_w3810_,
		_w3813_,
		_w3814_
	);
	LUT4 #(
		.INIT('h0b0f)
	) name1668 (
		\u14_u5_en_out_l2_reg/P0001 ,
		\u14_u5_en_out_l_reg/NET0131 ,
		\u8_dout_reg[5]/P0001 ,
		\valid_s_reg/NET0131 ,
		_w3815_
	);
	LUT2 #(
		.INIT('h2)
	) name1669 (
		\u13_occ1_r_reg[8]/NET0131 ,
		_w3815_,
		_w3816_
	);
	LUT2 #(
		.INIT('h4)
	) name1670 (
		_w3814_,
		_w3816_,
		_w3817_
	);
	LUT3 #(
		.INIT('h80)
	) name1671 (
		\u8_rp_reg[0]/P0001 ,
		_w3742_,
		_w3743_,
		_w3818_
	);
	LUT4 #(
		.INIT('h8ccc)
	) name1672 (
		\u8_rp_reg[0]/P0001 ,
		_w2156_,
		_w3784_,
		_w3785_,
		_w3819_
	);
	LUT3 #(
		.INIT('h2a)
	) name1673 (
		_w3567_,
		_w3801_,
		_w3802_,
		_w3820_
	);
	LUT4 #(
		.INIT('ha222)
	) name1674 (
		_w2155_,
		_w2550_,
		_w3564_,
		_w3565_,
		_w3821_
	);
	LUT4 #(
		.INIT('h0b00)
	) name1675 (
		_w3818_,
		_w3819_,
		_w3820_,
		_w3821_,
		_w3822_
	);
	LUT4 #(
		.INIT('h0b0f)
	) name1676 (
		\u14_u5_en_out_l2_reg/P0001 ,
		\u14_u5_en_out_l_reg/NET0131 ,
		\u8_dout_reg[6]/P0001 ,
		\valid_s_reg/NET0131 ,
		_w3823_
	);
	LUT2 #(
		.INIT('h2)
	) name1677 (
		\u13_occ1_r_reg[8]/NET0131 ,
		_w3823_,
		_w3824_
	);
	LUT2 #(
		.INIT('h4)
	) name1678 (
		_w3822_,
		_w3824_,
		_w3825_
	);
	LUT3 #(
		.INIT('h80)
	) name1679 (
		\u8_rp_reg[0]/P0001 ,
		_w3766_,
		_w3767_,
		_w3826_
	);
	LUT4 #(
		.INIT('h8ccc)
	) name1680 (
		\u8_rp_reg[0]/P0001 ,
		_w2156_,
		_w3791_,
		_w3792_,
		_w3827_
	);
	LUT3 #(
		.INIT('h2a)
	) name1681 (
		_w3567_,
		_w3811_,
		_w3812_,
		_w3828_
	);
	LUT4 #(
		.INIT('ha222)
	) name1682 (
		_w2155_,
		_w2550_,
		_w3595_,
		_w3596_,
		_w3829_
	);
	LUT4 #(
		.INIT('h0b00)
	) name1683 (
		_w3826_,
		_w3827_,
		_w3828_,
		_w3829_,
		_w3830_
	);
	LUT4 #(
		.INIT('h0b0f)
	) name1684 (
		\u14_u5_en_out_l2_reg/P0001 ,
		\u14_u5_en_out_l_reg/NET0131 ,
		\u8_dout_reg[7]/P0001 ,
		\valid_s_reg/NET0131 ,
		_w3831_
	);
	LUT2 #(
		.INIT('h2)
	) name1685 (
		\u13_occ1_r_reg[8]/NET0131 ,
		_w3831_,
		_w3832_
	);
	LUT2 #(
		.INIT('h4)
	) name1686 (
		_w3830_,
		_w3832_,
		_w3833_
	);
	LUT4 #(
		.INIT('hc4cc)
	) name1687 (
		\u8_mem_reg[2][20]/NET0131 ,
		\u8_rp_reg[0]/P0001 ,
		\u8_rp_reg[1]/NET0131 ,
		\u8_rp_reg[2]/NET0131 ,
		_w3834_
	);
	LUT3 #(
		.INIT('h02)
	) name1688 (
		\u8_mem_reg[0][20]/NET0131 ,
		\u8_rp_reg[1]/NET0131 ,
		\u8_rp_reg[2]/NET0131 ,
		_w3835_
	);
	LUT4 #(
		.INIT('h3f5f)
	) name1689 (
		\u8_mem_reg[1][20]/NET0131 ,
		\u8_mem_reg[3][20]/NET0131 ,
		\u8_rp_reg[1]/NET0131 ,
		\u8_rp_reg[2]/NET0131 ,
		_w3836_
	);
	LUT3 #(
		.INIT('h40)
	) name1690 (
		_w3835_,
		_w3834_,
		_w3836_,
		_w3837_
	);
	LUT4 #(
		.INIT('h8ccc)
	) name1691 (
		\u8_rp_reg[0]/P0001 ,
		_w2156_,
		_w3801_,
		_w3802_,
		_w3838_
	);
	LUT3 #(
		.INIT('h70)
	) name1692 (
		_w3564_,
		_w3565_,
		_w3567_,
		_w3839_
	);
	LUT4 #(
		.INIT('ha222)
	) name1693 (
		_w2155_,
		_w2550_,
		_w3568_,
		_w3569_,
		_w3840_
	);
	LUT4 #(
		.INIT('h0b00)
	) name1694 (
		_w3837_,
		_w3838_,
		_w3839_,
		_w3840_,
		_w3841_
	);
	LUT4 #(
		.INIT('h0b0f)
	) name1695 (
		\u14_u5_en_out_l2_reg/P0001 ,
		\u14_u5_en_out_l_reg/NET0131 ,
		\u8_dout_reg[8]/P0001 ,
		\valid_s_reg/NET0131 ,
		_w3842_
	);
	LUT2 #(
		.INIT('h2)
	) name1696 (
		\u13_occ1_r_reg[8]/NET0131 ,
		_w3842_,
		_w3843_
	);
	LUT2 #(
		.INIT('h4)
	) name1697 (
		_w3841_,
		_w3843_,
		_w3844_
	);
	LUT4 #(
		.INIT('hc4cc)
	) name1698 (
		\u8_mem_reg[2][21]/NET0131 ,
		\u8_rp_reg[0]/P0001 ,
		\u8_rp_reg[1]/NET0131 ,
		\u8_rp_reg[2]/NET0131 ,
		_w3845_
	);
	LUT3 #(
		.INIT('h02)
	) name1699 (
		\u8_mem_reg[0][21]/NET0131 ,
		\u8_rp_reg[1]/NET0131 ,
		\u8_rp_reg[2]/NET0131 ,
		_w3846_
	);
	LUT4 #(
		.INIT('h3f5f)
	) name1700 (
		\u8_mem_reg[1][21]/NET0131 ,
		\u8_mem_reg[3][21]/NET0131 ,
		\u8_rp_reg[1]/NET0131 ,
		\u8_rp_reg[2]/NET0131 ,
		_w3847_
	);
	LUT3 #(
		.INIT('h40)
	) name1701 (
		_w3846_,
		_w3845_,
		_w3847_,
		_w3848_
	);
	LUT4 #(
		.INIT('h8ccc)
	) name1702 (
		\u8_rp_reg[0]/P0001 ,
		_w2156_,
		_w3811_,
		_w3812_,
		_w3849_
	);
	LUT3 #(
		.INIT('h2a)
	) name1703 (
		_w3567_,
		_w3595_,
		_w3596_,
		_w3850_
	);
	LUT4 #(
		.INIT('ha222)
	) name1704 (
		_w2155_,
		_w2550_,
		_w3598_,
		_w3599_,
		_w3851_
	);
	LUT4 #(
		.INIT('h0b00)
	) name1705 (
		_w3848_,
		_w3849_,
		_w3850_,
		_w3851_,
		_w3852_
	);
	LUT4 #(
		.INIT('h0b0f)
	) name1706 (
		\u14_u5_en_out_l2_reg/P0001 ,
		\u14_u5_en_out_l_reg/NET0131 ,
		\u8_dout_reg[9]/P0001 ,
		\valid_s_reg/NET0131 ,
		_w3853_
	);
	LUT2 #(
		.INIT('h2)
	) name1707 (
		\u13_occ1_r_reg[8]/NET0131 ,
		_w3853_,
		_w3854_
	);
	LUT2 #(
		.INIT('h4)
	) name1708 (
		_w3852_,
		_w3854_,
		_w3855_
	);
	LUT4 #(
		.INIT('h8848)
	) name1709 (
		\u11_wp_reg[1]/P0001 ,
		\u13_icc_r_reg[16]/NET0131 ,
		_w2565_,
		_w2567_,
		_w3856_
	);
	LUT4 #(
		.INIT('h8828)
	) name1710 (
		\u13_icc_r_reg[0]/NET0131 ,
		\u9_wp_reg[1]/P0001 ,
		_w2686_,
		_w2688_,
		_w3857_
	);
	LUT4 #(
		.INIT('h8848)
	) name1711 (
		\u10_wp_reg[1]/P0001 ,
		\u13_icc_r_reg[8]/NET0131 ,
		_w2792_,
		_w2794_,
		_w3858_
	);
	LUT3 #(
		.INIT('h48)
	) name1712 (
		\u11_wp_reg[3]/P0001 ,
		\u13_icc_r_reg[16]/NET0131 ,
		_w2570_,
		_w3859_
	);
	LUT3 #(
		.INIT('h28)
	) name1713 (
		\u13_icc_r_reg[0]/NET0131 ,
		\u9_wp_reg[3]/P0001 ,
		_w2691_,
		_w3860_
	);
	LUT3 #(
		.INIT('h48)
	) name1714 (
		\u10_wp_reg[3]/P0001 ,
		\u13_icc_r_reg[8]/NET0131 ,
		_w2797_,
		_w3861_
	);
	LUT2 #(
		.INIT('h2)
	) name1715 (
		\u26_ps_cnt_reg[0]/NET0131 ,
		\u26_ps_cnt_reg[1]/NET0131 ,
		_w3862_
	);
	LUT4 #(
		.INIT('h1000)
	) name1716 (
		\u26_ps_cnt_reg[2]/NET0131 ,
		\u26_ps_cnt_reg[3]/NET0131 ,
		\u26_ps_cnt_reg[4]/NET0131 ,
		\u26_ps_cnt_reg[5]/NET0131 ,
		_w3863_
	);
	LUT3 #(
		.INIT('h15)
	) name1717 (
		\u13_ac97_rst_force_reg/P0001 ,
		_w3862_,
		_w3863_,
		_w3864_
	);
	LUT4 #(
		.INIT('h1111)
	) name1718 (
		\u13_ac97_rst_force_reg/P0001 ,
		\u26_ps_cnt_reg[0]/NET0131 ,
		\u26_ps_cnt_reg[1]/NET0131 ,
		_w3863_,
		_w3865_
	);
	LUT4 #(
		.INIT('h1014)
	) name1719 (
		\u13_ac97_rst_force_reg/P0001 ,
		\u26_ps_cnt_reg[0]/NET0131 ,
		\u26_ps_cnt_reg[1]/NET0131 ,
		_w3863_,
		_w3866_
	);
	LUT3 #(
		.INIT('h78)
	) name1720 (
		\u26_ps_cnt_reg[0]/NET0131 ,
		\u26_ps_cnt_reg[1]/NET0131 ,
		\u26_ps_cnt_reg[2]/NET0131 ,
		_w3867_
	);
	LUT4 #(
		.INIT('h1500)
	) name1721 (
		\u13_ac97_rst_force_reg/P0001 ,
		_w3862_,
		_w3863_,
		_w3867_,
		_w3868_
	);
	LUT4 #(
		.INIT('h8000)
	) name1722 (
		\u26_ps_cnt_reg[0]/NET0131 ,
		\u26_ps_cnt_reg[1]/NET0131 ,
		\u26_ps_cnt_reg[2]/NET0131 ,
		\u26_ps_cnt_reg[3]/NET0131 ,
		_w3869_
	);
	LUT4 #(
		.INIT('h7f80)
	) name1723 (
		\u26_ps_cnt_reg[0]/NET0131 ,
		\u26_ps_cnt_reg[1]/NET0131 ,
		\u26_ps_cnt_reg[2]/NET0131 ,
		\u26_ps_cnt_reg[3]/NET0131 ,
		_w3870_
	);
	LUT4 #(
		.INIT('h1500)
	) name1724 (
		\u13_ac97_rst_force_reg/P0001 ,
		_w3862_,
		_w3863_,
		_w3870_,
		_w3871_
	);
	LUT2 #(
		.INIT('h8)
	) name1725 (
		\u26_ps_cnt_reg[4]/NET0131 ,
		_w3869_,
		_w3872_
	);
	LUT3 #(
		.INIT('h48)
	) name1726 (
		\u26_ps_cnt_reg[4]/NET0131 ,
		_w3864_,
		_w3869_,
		_w3873_
	);
	LUT3 #(
		.INIT('h48)
	) name1727 (
		\u26_ps_cnt_reg[5]/NET0131 ,
		_w3864_,
		_w3872_,
		_w3874_
	);
	LUT4 #(
		.INIT('h4888)
	) name1728 (
		\u11_wp_reg[0]/NET0131 ,
		\u13_icc_r_reg[16]/NET0131 ,
		_w2565_,
		_w2566_,
		_w3875_
	);
	LUT4 #(
		.INIT('h2888)
	) name1729 (
		\u13_icc_r_reg[0]/NET0131 ,
		\u9_wp_reg[0]/NET0131 ,
		_w2686_,
		_w2687_,
		_w3876_
	);
	LUT4 #(
		.INIT('h4888)
	) name1730 (
		\u10_wp_reg[0]/NET0131 ,
		\u13_icc_r_reg[8]/NET0131 ,
		_w2792_,
		_w2793_,
		_w3877_
	);
	LUT2 #(
		.INIT('h4)
	) name1731 (
		\u10_wp_reg[1]/P0001 ,
		\u10_wp_reg[2]/P0001 ,
		_w3878_
	);
	LUT3 #(
		.INIT('h20)
	) name1732 (
		_w2792_,
		_w2794_,
		_w3878_,
		_w3879_
	);
	LUT4 #(
		.INIT('ha2aa)
	) name1733 (
		\u10_mem_reg[2][18]/P0001 ,
		_w2792_,
		_w2794_,
		_w3878_,
		_w3880_
	);
	LUT4 #(
		.INIT('haebf)
	) name1734 (
		\u13_icc_r_reg[10]/NET0131 ,
		\u13_icc_r_reg[11]/NET0131 ,
		\u1_slt4_reg[18]/P0001 ,
		\u1_slt4_reg[6]/P0001 ,
		_w3881_
	);
	LUT4 #(
		.INIT('h0020)
	) name1735 (
		_w2792_,
		_w2794_,
		_w3878_,
		_w3881_,
		_w3882_
	);
	LUT2 #(
		.INIT('he)
	) name1736 (
		_w3880_,
		_w3882_,
		_w3883_
	);
	LUT4 #(
		.INIT('ha2aa)
	) name1737 (
		\u10_mem_reg[2][19]/P0001 ,
		_w2792_,
		_w2794_,
		_w3878_,
		_w3884_
	);
	LUT4 #(
		.INIT('haebf)
	) name1738 (
		\u13_icc_r_reg[10]/NET0131 ,
		\u13_icc_r_reg[11]/NET0131 ,
		\u1_slt4_reg[19]/P0001 ,
		\u1_slt4_reg[7]/P0001 ,
		_w3885_
	);
	LUT4 #(
		.INIT('h0020)
	) name1739 (
		_w2792_,
		_w2794_,
		_w3878_,
		_w3885_,
		_w3886_
	);
	LUT2 #(
		.INIT('he)
	) name1740 (
		_w3884_,
		_w3886_,
		_w3887_
	);
	LUT4 #(
		.INIT('ha2aa)
	) name1741 (
		\u10_mem_reg[2][20]/P0001 ,
		_w2792_,
		_w2794_,
		_w3878_,
		_w3888_
	);
	LUT3 #(
		.INIT('h10)
	) name1742 (
		\u13_icc_r_reg[10]/NET0131 ,
		\u13_icc_r_reg[11]/NET0131 ,
		\u1_slt4_reg[8]/P0001 ,
		_w3889_
	);
	LUT4 #(
		.INIT('h2000)
	) name1743 (
		_w2792_,
		_w2794_,
		_w3878_,
		_w3889_,
		_w3890_
	);
	LUT2 #(
		.INIT('he)
	) name1744 (
		_w3888_,
		_w3890_,
		_w3891_
	);
	LUT4 #(
		.INIT('ha2aa)
	) name1745 (
		\u10_mem_reg[2][21]/P0001 ,
		_w2792_,
		_w2794_,
		_w3878_,
		_w3892_
	);
	LUT3 #(
		.INIT('h10)
	) name1746 (
		\u13_icc_r_reg[10]/NET0131 ,
		\u13_icc_r_reg[11]/NET0131 ,
		\u1_slt4_reg[9]/P0001 ,
		_w3893_
	);
	LUT4 #(
		.INIT('h2000)
	) name1747 (
		_w2792_,
		_w2794_,
		_w3878_,
		_w3893_,
		_w3894_
	);
	LUT2 #(
		.INIT('he)
	) name1748 (
		_w3892_,
		_w3894_,
		_w3895_
	);
	LUT4 #(
		.INIT('ha2aa)
	) name1749 (
		\u10_mem_reg[2][22]/P0001 ,
		_w2792_,
		_w2794_,
		_w3878_,
		_w3896_
	);
	LUT3 #(
		.INIT('h10)
	) name1750 (
		\u13_icc_r_reg[10]/NET0131 ,
		\u13_icc_r_reg[11]/NET0131 ,
		\u1_slt4_reg[10]/P0001 ,
		_w3897_
	);
	LUT4 #(
		.INIT('h2000)
	) name1751 (
		_w2792_,
		_w2794_,
		_w3878_,
		_w3897_,
		_w3898_
	);
	LUT2 #(
		.INIT('he)
	) name1752 (
		_w3896_,
		_w3898_,
		_w3899_
	);
	LUT4 #(
		.INIT('ha2aa)
	) name1753 (
		\u10_mem_reg[2][23]/P0001 ,
		_w2792_,
		_w2794_,
		_w3878_,
		_w3900_
	);
	LUT3 #(
		.INIT('h10)
	) name1754 (
		\u13_icc_r_reg[10]/NET0131 ,
		\u13_icc_r_reg[11]/NET0131 ,
		\u1_slt4_reg[11]/P0001 ,
		_w3901_
	);
	LUT4 #(
		.INIT('h2000)
	) name1755 (
		_w2792_,
		_w2794_,
		_w3878_,
		_w3901_,
		_w3902_
	);
	LUT2 #(
		.INIT('he)
	) name1756 (
		_w3900_,
		_w3902_,
		_w3903_
	);
	LUT2 #(
		.INIT('h1)
	) name1757 (
		\u9_wp_reg[1]/P0001 ,
		\u9_wp_reg[2]/P0001 ,
		_w3904_
	);
	LUT3 #(
		.INIT('h20)
	) name1758 (
		_w2686_,
		_w2688_,
		_w3904_,
		_w3905_
	);
	LUT4 #(
		.INIT('haebf)
	) name1759 (
		\u13_icc_r_reg[2]/NET0131 ,
		\u13_icc_r_reg[3]/NET0131 ,
		\u1_slt3_reg[18]/P0001 ,
		\u1_slt3_reg[6]/P0001 ,
		_w3906_
	);
	LUT4 #(
		.INIT('h0020)
	) name1760 (
		_w2686_,
		_w2688_,
		_w3904_,
		_w3906_,
		_w3907_
	);
	LUT4 #(
		.INIT('ha2aa)
	) name1761 (
		\u9_mem_reg[0][18]/P0001 ,
		_w2686_,
		_w2688_,
		_w3904_,
		_w3908_
	);
	LUT2 #(
		.INIT('he)
	) name1762 (
		_w3907_,
		_w3908_,
		_w3909_
	);
	LUT4 #(
		.INIT('haebf)
	) name1763 (
		\u13_icc_r_reg[2]/NET0131 ,
		\u13_icc_r_reg[3]/NET0131 ,
		\u1_slt3_reg[19]/P0001 ,
		\u1_slt3_reg[7]/P0001 ,
		_w3910_
	);
	LUT4 #(
		.INIT('h0020)
	) name1764 (
		_w2686_,
		_w2688_,
		_w3904_,
		_w3910_,
		_w3911_
	);
	LUT4 #(
		.INIT('ha2aa)
	) name1765 (
		\u9_mem_reg[0][19]/P0001 ,
		_w2686_,
		_w2688_,
		_w3904_,
		_w3912_
	);
	LUT2 #(
		.INIT('he)
	) name1766 (
		_w3911_,
		_w3912_,
		_w3913_
	);
	LUT4 #(
		.INIT('ha2aa)
	) name1767 (
		\u10_mem_reg[2][24]/P0001 ,
		_w2792_,
		_w2794_,
		_w3878_,
		_w3914_
	);
	LUT3 #(
		.INIT('h10)
	) name1768 (
		\u13_icc_r_reg[10]/NET0131 ,
		\u13_icc_r_reg[11]/NET0131 ,
		\u1_slt4_reg[12]/P0001 ,
		_w3915_
	);
	LUT4 #(
		.INIT('h2000)
	) name1769 (
		_w2792_,
		_w2794_,
		_w3878_,
		_w3915_,
		_w3916_
	);
	LUT2 #(
		.INIT('he)
	) name1770 (
		_w3914_,
		_w3916_,
		_w3917_
	);
	LUT4 #(
		.INIT('ha2aa)
	) name1771 (
		\u10_mem_reg[2][25]/P0001 ,
		_w2792_,
		_w2794_,
		_w3878_,
		_w3918_
	);
	LUT3 #(
		.INIT('h10)
	) name1772 (
		\u13_icc_r_reg[10]/NET0131 ,
		\u13_icc_r_reg[11]/NET0131 ,
		\u1_slt4_reg[13]/P0001 ,
		_w3919_
	);
	LUT4 #(
		.INIT('h2000)
	) name1773 (
		_w2792_,
		_w2794_,
		_w3878_,
		_w3919_,
		_w3920_
	);
	LUT2 #(
		.INIT('he)
	) name1774 (
		_w3918_,
		_w3920_,
		_w3921_
	);
	LUT4 #(
		.INIT('ha2aa)
	) name1775 (
		\u10_mem_reg[2][26]/P0001 ,
		_w2792_,
		_w2794_,
		_w3878_,
		_w3922_
	);
	LUT3 #(
		.INIT('h10)
	) name1776 (
		\u13_icc_r_reg[10]/NET0131 ,
		\u13_icc_r_reg[11]/NET0131 ,
		\u1_slt4_reg[14]/P0001 ,
		_w3923_
	);
	LUT4 #(
		.INIT('h2000)
	) name1777 (
		_w2792_,
		_w2794_,
		_w3878_,
		_w3923_,
		_w3924_
	);
	LUT2 #(
		.INIT('he)
	) name1778 (
		_w3922_,
		_w3924_,
		_w3925_
	);
	LUT4 #(
		.INIT('ha2aa)
	) name1779 (
		\u10_mem_reg[2][27]/P0001 ,
		_w2792_,
		_w2794_,
		_w3878_,
		_w3926_
	);
	LUT3 #(
		.INIT('h10)
	) name1780 (
		\u13_icc_r_reg[10]/NET0131 ,
		\u13_icc_r_reg[11]/NET0131 ,
		\u1_slt4_reg[15]/P0001 ,
		_w3927_
	);
	LUT4 #(
		.INIT('h2000)
	) name1781 (
		_w2792_,
		_w2794_,
		_w3878_,
		_w3927_,
		_w3928_
	);
	LUT2 #(
		.INIT('he)
	) name1782 (
		_w3926_,
		_w3928_,
		_w3929_
	);
	LUT4 #(
		.INIT('ha2aa)
	) name1783 (
		\u10_mem_reg[2][28]/P0001 ,
		_w2792_,
		_w2794_,
		_w3878_,
		_w3930_
	);
	LUT3 #(
		.INIT('h10)
	) name1784 (
		\u13_icc_r_reg[10]/NET0131 ,
		\u13_icc_r_reg[11]/NET0131 ,
		\u1_slt4_reg[16]/P0001 ,
		_w3931_
	);
	LUT4 #(
		.INIT('h2000)
	) name1785 (
		_w2792_,
		_w2794_,
		_w3878_,
		_w3931_,
		_w3932_
	);
	LUT2 #(
		.INIT('he)
	) name1786 (
		_w3930_,
		_w3932_,
		_w3933_
	);
	LUT4 #(
		.INIT('h0020)
	) name1787 (
		\u9_wp_reg[1]/P0001 ,
		\u9_wp_reg[2]/P0001 ,
		_w2686_,
		_w2688_,
		_w3934_
	);
	LUT3 #(
		.INIT('h3a)
	) name1788 (
		\u9_mem_reg[1][18]/P0001 ,
		_w3906_,
		_w3934_,
		_w3935_
	);
	LUT3 #(
		.INIT('h3a)
	) name1789 (
		\u9_mem_reg[1][19]/P0001 ,
		_w3910_,
		_w3934_,
		_w3936_
	);
	LUT3 #(
		.INIT('h10)
	) name1790 (
		\u13_icc_r_reg[2]/NET0131 ,
		\u13_icc_r_reg[3]/NET0131 ,
		\u1_slt3_reg[8]/P0001 ,
		_w3937_
	);
	LUT3 #(
		.INIT('he2)
	) name1791 (
		\u9_mem_reg[1][20]/P0001 ,
		_w3934_,
		_w3937_,
		_w3938_
	);
	LUT3 #(
		.INIT('h10)
	) name1792 (
		\u13_icc_r_reg[2]/NET0131 ,
		\u13_icc_r_reg[3]/NET0131 ,
		\u1_slt3_reg[9]/P0001 ,
		_w3939_
	);
	LUT3 #(
		.INIT('he2)
	) name1793 (
		\u9_mem_reg[1][21]/P0001 ,
		_w3934_,
		_w3939_,
		_w3940_
	);
	LUT4 #(
		.INIT('ha2aa)
	) name1794 (
		\u10_mem_reg[2][29]/P0001 ,
		_w2792_,
		_w2794_,
		_w3878_,
		_w3941_
	);
	LUT3 #(
		.INIT('h10)
	) name1795 (
		\u13_icc_r_reg[10]/NET0131 ,
		\u13_icc_r_reg[11]/NET0131 ,
		\u1_slt4_reg[17]/P0001 ,
		_w3942_
	);
	LUT4 #(
		.INIT('h2000)
	) name1796 (
		_w2792_,
		_w2794_,
		_w3878_,
		_w3942_,
		_w3943_
	);
	LUT2 #(
		.INIT('he)
	) name1797 (
		_w3941_,
		_w3943_,
		_w3944_
	);
	LUT3 #(
		.INIT('h10)
	) name1798 (
		\u13_icc_r_reg[2]/NET0131 ,
		\u13_icc_r_reg[3]/NET0131 ,
		\u1_slt3_reg[10]/P0001 ,
		_w3945_
	);
	LUT3 #(
		.INIT('he2)
	) name1799 (
		\u9_mem_reg[1][22]/P0001 ,
		_w3934_,
		_w3945_,
		_w3946_
	);
	LUT3 #(
		.INIT('h10)
	) name1800 (
		\u13_icc_r_reg[2]/NET0131 ,
		\u13_icc_r_reg[3]/NET0131 ,
		\u1_slt3_reg[11]/P0001 ,
		_w3947_
	);
	LUT3 #(
		.INIT('he2)
	) name1801 (
		\u9_mem_reg[1][23]/P0001 ,
		_w3934_,
		_w3947_,
		_w3948_
	);
	LUT3 #(
		.INIT('h10)
	) name1802 (
		\u13_icc_r_reg[2]/NET0131 ,
		\u13_icc_r_reg[3]/NET0131 ,
		\u1_slt3_reg[12]/P0001 ,
		_w3949_
	);
	LUT3 #(
		.INIT('he2)
	) name1803 (
		\u9_mem_reg[1][24]/P0001 ,
		_w3934_,
		_w3949_,
		_w3950_
	);
	LUT3 #(
		.INIT('h10)
	) name1804 (
		\u13_icc_r_reg[2]/NET0131 ,
		\u13_icc_r_reg[3]/NET0131 ,
		\u1_slt3_reg[13]/P0001 ,
		_w3951_
	);
	LUT3 #(
		.INIT('he2)
	) name1805 (
		\u9_mem_reg[1][25]/P0001 ,
		_w3934_,
		_w3951_,
		_w3952_
	);
	LUT3 #(
		.INIT('h10)
	) name1806 (
		\u13_icc_r_reg[2]/NET0131 ,
		\u13_icc_r_reg[3]/NET0131 ,
		\u1_slt3_reg[14]/P0001 ,
		_w3953_
	);
	LUT3 #(
		.INIT('he2)
	) name1807 (
		\u9_mem_reg[1][26]/P0001 ,
		_w3934_,
		_w3953_,
		_w3954_
	);
	LUT3 #(
		.INIT('h10)
	) name1808 (
		\u13_icc_r_reg[2]/NET0131 ,
		\u13_icc_r_reg[3]/NET0131 ,
		\u1_slt3_reg[15]/P0001 ,
		_w3955_
	);
	LUT3 #(
		.INIT('he2)
	) name1809 (
		\u9_mem_reg[1][27]/P0001 ,
		_w3934_,
		_w3955_,
		_w3956_
	);
	LUT3 #(
		.INIT('h10)
	) name1810 (
		\u13_icc_r_reg[2]/NET0131 ,
		\u13_icc_r_reg[3]/NET0131 ,
		\u1_slt3_reg[16]/P0001 ,
		_w3957_
	);
	LUT3 #(
		.INIT('he2)
	) name1811 (
		\u9_mem_reg[1][28]/P0001 ,
		_w3934_,
		_w3957_,
		_w3958_
	);
	LUT3 #(
		.INIT('h10)
	) name1812 (
		\u13_icc_r_reg[2]/NET0131 ,
		\u13_icc_r_reg[3]/NET0131 ,
		\u1_slt3_reg[17]/P0001 ,
		_w3959_
	);
	LUT3 #(
		.INIT('he2)
	) name1813 (
		\u9_mem_reg[1][29]/P0001 ,
		_w3934_,
		_w3959_,
		_w3960_
	);
	LUT3 #(
		.INIT('h10)
	) name1814 (
		\u13_icc_r_reg[2]/NET0131 ,
		\u13_icc_r_reg[3]/NET0131 ,
		\u1_slt3_reg[18]/P0001 ,
		_w3961_
	);
	LUT3 #(
		.INIT('he2)
	) name1815 (
		\u9_mem_reg[1][30]/P0001 ,
		_w3934_,
		_w3961_,
		_w3962_
	);
	LUT3 #(
		.INIT('h10)
	) name1816 (
		\u13_icc_r_reg[2]/NET0131 ,
		\u13_icc_r_reg[3]/NET0131 ,
		\u1_slt3_reg[19]/P0001 ,
		_w3963_
	);
	LUT3 #(
		.INIT('he2)
	) name1817 (
		\u9_mem_reg[1][31]/P0001 ,
		_w3934_,
		_w3963_,
		_w3964_
	);
	LUT4 #(
		.INIT('ha2aa)
	) name1818 (
		\u10_mem_reg[2][30]/P0001 ,
		_w2792_,
		_w2794_,
		_w3878_,
		_w3965_
	);
	LUT3 #(
		.INIT('h10)
	) name1819 (
		\u13_icc_r_reg[10]/NET0131 ,
		\u13_icc_r_reg[11]/NET0131 ,
		\u1_slt4_reg[18]/P0001 ,
		_w3966_
	);
	LUT4 #(
		.INIT('h2000)
	) name1820 (
		_w2792_,
		_w2794_,
		_w3878_,
		_w3966_,
		_w3967_
	);
	LUT2 #(
		.INIT('he)
	) name1821 (
		_w3965_,
		_w3967_,
		_w3968_
	);
	LUT4 #(
		.INIT('ha2aa)
	) name1822 (
		\u10_mem_reg[2][31]/P0001 ,
		_w2792_,
		_w2794_,
		_w3878_,
		_w3969_
	);
	LUT3 #(
		.INIT('h10)
	) name1823 (
		\u13_icc_r_reg[10]/NET0131 ,
		\u13_icc_r_reg[11]/NET0131 ,
		\u1_slt4_reg[19]/P0001 ,
		_w3970_
	);
	LUT4 #(
		.INIT('h2000)
	) name1824 (
		_w2792_,
		_w2794_,
		_w3878_,
		_w3970_,
		_w3971_
	);
	LUT2 #(
		.INIT('he)
	) name1825 (
		_w3969_,
		_w3971_,
		_w3972_
	);
	LUT2 #(
		.INIT('h4)
	) name1826 (
		\u9_wp_reg[1]/P0001 ,
		\u9_wp_reg[2]/P0001 ,
		_w3973_
	);
	LUT3 #(
		.INIT('h20)
	) name1827 (
		_w2686_,
		_w2688_,
		_w3973_,
		_w3974_
	);
	LUT4 #(
		.INIT('ha2aa)
	) name1828 (
		\u9_mem_reg[2][18]/P0001 ,
		_w2686_,
		_w2688_,
		_w3973_,
		_w3975_
	);
	LUT4 #(
		.INIT('h0200)
	) name1829 (
		_w2686_,
		_w2688_,
		_w3906_,
		_w3973_,
		_w3976_
	);
	LUT2 #(
		.INIT('he)
	) name1830 (
		_w3975_,
		_w3976_,
		_w3977_
	);
	LUT4 #(
		.INIT('ha2aa)
	) name1831 (
		\u9_mem_reg[2][19]/P0001 ,
		_w2686_,
		_w2688_,
		_w3973_,
		_w3978_
	);
	LUT4 #(
		.INIT('h0200)
	) name1832 (
		_w2686_,
		_w2688_,
		_w3910_,
		_w3973_,
		_w3979_
	);
	LUT2 #(
		.INIT('he)
	) name1833 (
		_w3978_,
		_w3979_,
		_w3980_
	);
	LUT4 #(
		.INIT('ha2aa)
	) name1834 (
		\u9_mem_reg[2][20]/P0001 ,
		_w2686_,
		_w2688_,
		_w3973_,
		_w3981_
	);
	LUT4 #(
		.INIT('h2000)
	) name1835 (
		_w2686_,
		_w2688_,
		_w3937_,
		_w3973_,
		_w3982_
	);
	LUT2 #(
		.INIT('he)
	) name1836 (
		_w3981_,
		_w3982_,
		_w3983_
	);
	LUT4 #(
		.INIT('ha2aa)
	) name1837 (
		\u9_mem_reg[2][21]/P0001 ,
		_w2686_,
		_w2688_,
		_w3973_,
		_w3984_
	);
	LUT4 #(
		.INIT('h2000)
	) name1838 (
		_w2686_,
		_w2688_,
		_w3939_,
		_w3973_,
		_w3985_
	);
	LUT2 #(
		.INIT('he)
	) name1839 (
		_w3984_,
		_w3985_,
		_w3986_
	);
	LUT4 #(
		.INIT('ha2aa)
	) name1840 (
		\u9_mem_reg[2][22]/P0001 ,
		_w2686_,
		_w2688_,
		_w3973_,
		_w3987_
	);
	LUT4 #(
		.INIT('h2000)
	) name1841 (
		_w2686_,
		_w2688_,
		_w3945_,
		_w3973_,
		_w3988_
	);
	LUT2 #(
		.INIT('he)
	) name1842 (
		_w3987_,
		_w3988_,
		_w3989_
	);
	LUT4 #(
		.INIT('ha2aa)
	) name1843 (
		\u9_mem_reg[2][23]/P0001 ,
		_w2686_,
		_w2688_,
		_w3973_,
		_w3990_
	);
	LUT4 #(
		.INIT('h2000)
	) name1844 (
		_w2686_,
		_w2688_,
		_w3947_,
		_w3973_,
		_w3991_
	);
	LUT2 #(
		.INIT('he)
	) name1845 (
		_w3990_,
		_w3991_,
		_w3992_
	);
	LUT4 #(
		.INIT('ha2aa)
	) name1846 (
		\u9_mem_reg[2][24]/P0001 ,
		_w2686_,
		_w2688_,
		_w3973_,
		_w3993_
	);
	LUT4 #(
		.INIT('h2000)
	) name1847 (
		_w2686_,
		_w2688_,
		_w3949_,
		_w3973_,
		_w3994_
	);
	LUT2 #(
		.INIT('he)
	) name1848 (
		_w3993_,
		_w3994_,
		_w3995_
	);
	LUT4 #(
		.INIT('ha2aa)
	) name1849 (
		\u9_mem_reg[2][25]/P0001 ,
		_w2686_,
		_w2688_,
		_w3973_,
		_w3996_
	);
	LUT4 #(
		.INIT('h2000)
	) name1850 (
		_w2686_,
		_w2688_,
		_w3951_,
		_w3973_,
		_w3997_
	);
	LUT2 #(
		.INIT('he)
	) name1851 (
		_w3996_,
		_w3997_,
		_w3998_
	);
	LUT4 #(
		.INIT('ha2aa)
	) name1852 (
		\u9_mem_reg[2][26]/P0001 ,
		_w2686_,
		_w2688_,
		_w3973_,
		_w3999_
	);
	LUT4 #(
		.INIT('h2000)
	) name1853 (
		_w2686_,
		_w2688_,
		_w3953_,
		_w3973_,
		_w4000_
	);
	LUT2 #(
		.INIT('he)
	) name1854 (
		_w3999_,
		_w4000_,
		_w4001_
	);
	LUT4 #(
		.INIT('ha2aa)
	) name1855 (
		\u9_mem_reg[2][27]/P0001 ,
		_w2686_,
		_w2688_,
		_w3973_,
		_w4002_
	);
	LUT4 #(
		.INIT('h2000)
	) name1856 (
		_w2686_,
		_w2688_,
		_w3955_,
		_w3973_,
		_w4003_
	);
	LUT2 #(
		.INIT('he)
	) name1857 (
		_w4002_,
		_w4003_,
		_w4004_
	);
	LUT4 #(
		.INIT('ha2aa)
	) name1858 (
		\u9_mem_reg[2][28]/P0001 ,
		_w2686_,
		_w2688_,
		_w3973_,
		_w4005_
	);
	LUT4 #(
		.INIT('h2000)
	) name1859 (
		_w2686_,
		_w2688_,
		_w3957_,
		_w3973_,
		_w4006_
	);
	LUT2 #(
		.INIT('he)
	) name1860 (
		_w4005_,
		_w4006_,
		_w4007_
	);
	LUT4 #(
		.INIT('ha2aa)
	) name1861 (
		\u9_mem_reg[2][29]/P0001 ,
		_w2686_,
		_w2688_,
		_w3973_,
		_w4008_
	);
	LUT4 #(
		.INIT('h2000)
	) name1862 (
		_w2686_,
		_w2688_,
		_w3959_,
		_w3973_,
		_w4009_
	);
	LUT2 #(
		.INIT('he)
	) name1863 (
		_w4008_,
		_w4009_,
		_w4010_
	);
	LUT4 #(
		.INIT('ha2aa)
	) name1864 (
		\u9_mem_reg[2][30]/P0001 ,
		_w2686_,
		_w2688_,
		_w3973_,
		_w4011_
	);
	LUT4 #(
		.INIT('h2000)
	) name1865 (
		_w2686_,
		_w2688_,
		_w3961_,
		_w3973_,
		_w4012_
	);
	LUT2 #(
		.INIT('he)
	) name1866 (
		_w4011_,
		_w4012_,
		_w4013_
	);
	LUT4 #(
		.INIT('ha2aa)
	) name1867 (
		\u9_mem_reg[2][31]/P0001 ,
		_w2686_,
		_w2688_,
		_w3973_,
		_w4014_
	);
	LUT4 #(
		.INIT('h2000)
	) name1868 (
		_w2686_,
		_w2688_,
		_w3963_,
		_w3973_,
		_w4015_
	);
	LUT2 #(
		.INIT('he)
	) name1869 (
		_w4014_,
		_w4015_,
		_w4016_
	);
	LUT3 #(
		.INIT('h2e)
	) name1870 (
		\u9_mem_reg[3][18]/P0001 ,
		_w2691_,
		_w3906_,
		_w4017_
	);
	LUT3 #(
		.INIT('h2e)
	) name1871 (
		\u9_mem_reg[3][19]/P0001 ,
		_w2691_,
		_w3910_,
		_w4018_
	);
	LUT3 #(
		.INIT('he2)
	) name1872 (
		\u9_mem_reg[3][20]/P0001 ,
		_w2691_,
		_w3937_,
		_w4019_
	);
	LUT3 #(
		.INIT('he2)
	) name1873 (
		\u9_mem_reg[3][21]/P0001 ,
		_w2691_,
		_w3939_,
		_w4020_
	);
	LUT3 #(
		.INIT('he2)
	) name1874 (
		\u9_mem_reg[3][22]/P0001 ,
		_w2691_,
		_w3945_,
		_w4021_
	);
	LUT3 #(
		.INIT('he2)
	) name1875 (
		\u9_mem_reg[3][23]/P0001 ,
		_w2691_,
		_w3947_,
		_w4022_
	);
	LUT3 #(
		.INIT('he2)
	) name1876 (
		\u9_mem_reg[3][24]/P0001 ,
		_w2691_,
		_w3949_,
		_w4023_
	);
	LUT3 #(
		.INIT('he2)
	) name1877 (
		\u9_mem_reg[3][25]/P0001 ,
		_w2691_,
		_w3951_,
		_w4024_
	);
	LUT3 #(
		.INIT('he2)
	) name1878 (
		\u9_mem_reg[3][26]/P0001 ,
		_w2691_,
		_w3953_,
		_w4025_
	);
	LUT3 #(
		.INIT('he2)
	) name1879 (
		\u9_mem_reg[3][27]/P0001 ,
		_w2691_,
		_w3955_,
		_w4026_
	);
	LUT3 #(
		.INIT('he2)
	) name1880 (
		\u9_mem_reg[3][28]/P0001 ,
		_w2691_,
		_w3957_,
		_w4027_
	);
	LUT3 #(
		.INIT('he2)
	) name1881 (
		\u9_mem_reg[3][29]/P0001 ,
		_w2691_,
		_w3959_,
		_w4028_
	);
	LUT3 #(
		.INIT('he2)
	) name1882 (
		\u9_mem_reg[3][30]/P0001 ,
		_w2691_,
		_w3961_,
		_w4029_
	);
	LUT3 #(
		.INIT('he2)
	) name1883 (
		\u9_mem_reg[3][31]/P0001 ,
		_w2691_,
		_w3963_,
		_w4030_
	);
	LUT3 #(
		.INIT('h2e)
	) name1884 (
		\u10_mem_reg[3][18]/P0001 ,
		_w2797_,
		_w3881_,
		_w4031_
	);
	LUT3 #(
		.INIT('h2e)
	) name1885 (
		\u10_mem_reg[3][19]/P0001 ,
		_w2797_,
		_w3885_,
		_w4032_
	);
	LUT3 #(
		.INIT('he2)
	) name1886 (
		\u10_mem_reg[3][20]/P0001 ,
		_w2797_,
		_w3889_,
		_w4033_
	);
	LUT3 #(
		.INIT('he2)
	) name1887 (
		\u10_mem_reg[3][21]/P0001 ,
		_w2797_,
		_w3893_,
		_w4034_
	);
	LUT3 #(
		.INIT('he2)
	) name1888 (
		\u10_mem_reg[3][22]/P0001 ,
		_w2797_,
		_w3897_,
		_w4035_
	);
	LUT3 #(
		.INIT('he2)
	) name1889 (
		\u10_mem_reg[3][23]/P0001 ,
		_w2797_,
		_w3901_,
		_w4036_
	);
	LUT3 #(
		.INIT('he2)
	) name1890 (
		\u10_mem_reg[3][24]/P0001 ,
		_w2797_,
		_w3915_,
		_w4037_
	);
	LUT3 #(
		.INIT('he2)
	) name1891 (
		\u10_mem_reg[3][25]/P0001 ,
		_w2797_,
		_w3919_,
		_w4038_
	);
	LUT3 #(
		.INIT('he2)
	) name1892 (
		\u10_mem_reg[3][26]/P0001 ,
		_w2797_,
		_w3923_,
		_w4039_
	);
	LUT3 #(
		.INIT('he2)
	) name1893 (
		\u10_mem_reg[3][27]/P0001 ,
		_w2797_,
		_w3927_,
		_w4040_
	);
	LUT3 #(
		.INIT('he2)
	) name1894 (
		\u10_mem_reg[3][28]/P0001 ,
		_w2797_,
		_w3931_,
		_w4041_
	);
	LUT3 #(
		.INIT('he2)
	) name1895 (
		\u10_mem_reg[3][29]/P0001 ,
		_w2797_,
		_w3942_,
		_w4042_
	);
	LUT3 #(
		.INIT('he2)
	) name1896 (
		\u10_mem_reg[3][30]/P0001 ,
		_w2797_,
		_w3966_,
		_w4043_
	);
	LUT3 #(
		.INIT('he2)
	) name1897 (
		\u10_mem_reg[3][31]/P0001 ,
		_w2797_,
		_w3970_,
		_w4044_
	);
	LUT2 #(
		.INIT('h1)
	) name1898 (
		\u10_wp_reg[1]/P0001 ,
		\u10_wp_reg[2]/P0001 ,
		_w4045_
	);
	LUT3 #(
		.INIT('h20)
	) name1899 (
		_w2792_,
		_w2794_,
		_w4045_,
		_w4046_
	);
	LUT4 #(
		.INIT('ha2aa)
	) name1900 (
		\u10_mem_reg[0][18]/P0001 ,
		_w2792_,
		_w2794_,
		_w4045_,
		_w4047_
	);
	LUT4 #(
		.INIT('h0200)
	) name1901 (
		_w2792_,
		_w2794_,
		_w3881_,
		_w4045_,
		_w4048_
	);
	LUT2 #(
		.INIT('he)
	) name1902 (
		_w4047_,
		_w4048_,
		_w4049_
	);
	LUT2 #(
		.INIT('h1)
	) name1903 (
		\u11_wp_reg[1]/P0001 ,
		\u11_wp_reg[2]/P0001 ,
		_w4050_
	);
	LUT3 #(
		.INIT('h20)
	) name1904 (
		_w2565_,
		_w2567_,
		_w4050_,
		_w4051_
	);
	LUT4 #(
		.INIT('haebf)
	) name1905 (
		\u13_icc_r_reg[18]/NET0131 ,
		\u13_icc_r_reg[19]/NET0131 ,
		\u1_slt6_reg[18]/P0001 ,
		\u1_slt6_reg[6]/P0001 ,
		_w4052_
	);
	LUT4 #(
		.INIT('h0020)
	) name1906 (
		_w2565_,
		_w2567_,
		_w4050_,
		_w4052_,
		_w4053_
	);
	LUT4 #(
		.INIT('ha2aa)
	) name1907 (
		\u11_mem_reg[0][18]/P0001 ,
		_w2565_,
		_w2567_,
		_w4050_,
		_w4054_
	);
	LUT2 #(
		.INIT('he)
	) name1908 (
		_w4053_,
		_w4054_,
		_w4055_
	);
	LUT4 #(
		.INIT('haebf)
	) name1909 (
		\u13_icc_r_reg[18]/NET0131 ,
		\u13_icc_r_reg[19]/NET0131 ,
		\u1_slt6_reg[19]/P0001 ,
		\u1_slt6_reg[7]/P0001 ,
		_w4056_
	);
	LUT4 #(
		.INIT('h0020)
	) name1910 (
		_w2565_,
		_w2567_,
		_w4050_,
		_w4056_,
		_w4057_
	);
	LUT4 #(
		.INIT('ha2aa)
	) name1911 (
		\u11_mem_reg[0][19]/P0001 ,
		_w2565_,
		_w2567_,
		_w4050_,
		_w4058_
	);
	LUT2 #(
		.INIT('he)
	) name1912 (
		_w4057_,
		_w4058_,
		_w4059_
	);
	LUT4 #(
		.INIT('ha2aa)
	) name1913 (
		\u10_mem_reg[0][19]/P0001 ,
		_w2792_,
		_w2794_,
		_w4045_,
		_w4060_
	);
	LUT4 #(
		.INIT('h0200)
	) name1914 (
		_w2792_,
		_w2794_,
		_w3885_,
		_w4045_,
		_w4061_
	);
	LUT2 #(
		.INIT('he)
	) name1915 (
		_w4060_,
		_w4061_,
		_w4062_
	);
	LUT4 #(
		.INIT('h0020)
	) name1916 (
		\u11_wp_reg[1]/P0001 ,
		\u11_wp_reg[2]/P0001 ,
		_w2565_,
		_w2567_,
		_w4063_
	);
	LUT3 #(
		.INIT('h3a)
	) name1917 (
		\u11_mem_reg[1][18]/P0001 ,
		_w4052_,
		_w4063_,
		_w4064_
	);
	LUT3 #(
		.INIT('h3a)
	) name1918 (
		\u11_mem_reg[1][19]/P0001 ,
		_w4056_,
		_w4063_,
		_w4065_
	);
	LUT3 #(
		.INIT('h10)
	) name1919 (
		\u13_icc_r_reg[18]/NET0131 ,
		\u13_icc_r_reg[19]/NET0131 ,
		\u1_slt6_reg[8]/P0001 ,
		_w4066_
	);
	LUT3 #(
		.INIT('he2)
	) name1920 (
		\u11_mem_reg[1][20]/P0001 ,
		_w4063_,
		_w4066_,
		_w4067_
	);
	LUT3 #(
		.INIT('h10)
	) name1921 (
		\u13_icc_r_reg[18]/NET0131 ,
		\u13_icc_r_reg[19]/NET0131 ,
		\u1_slt6_reg[9]/P0001 ,
		_w4068_
	);
	LUT3 #(
		.INIT('he2)
	) name1922 (
		\u11_mem_reg[1][21]/P0001 ,
		_w4063_,
		_w4068_,
		_w4069_
	);
	LUT3 #(
		.INIT('h10)
	) name1923 (
		\u13_icc_r_reg[18]/NET0131 ,
		\u13_icc_r_reg[19]/NET0131 ,
		\u1_slt6_reg[10]/P0001 ,
		_w4070_
	);
	LUT3 #(
		.INIT('he2)
	) name1924 (
		\u11_mem_reg[1][22]/P0001 ,
		_w4063_,
		_w4070_,
		_w4071_
	);
	LUT3 #(
		.INIT('h10)
	) name1925 (
		\u13_icc_r_reg[18]/NET0131 ,
		\u13_icc_r_reg[19]/NET0131 ,
		\u1_slt6_reg[11]/P0001 ,
		_w4072_
	);
	LUT3 #(
		.INIT('he2)
	) name1926 (
		\u11_mem_reg[1][23]/P0001 ,
		_w4063_,
		_w4072_,
		_w4073_
	);
	LUT3 #(
		.INIT('h10)
	) name1927 (
		\u13_icc_r_reg[18]/NET0131 ,
		\u13_icc_r_reg[19]/NET0131 ,
		\u1_slt6_reg[12]/P0001 ,
		_w4074_
	);
	LUT3 #(
		.INIT('he2)
	) name1928 (
		\u11_mem_reg[1][24]/P0001 ,
		_w4063_,
		_w4074_,
		_w4075_
	);
	LUT3 #(
		.INIT('h10)
	) name1929 (
		\u13_icc_r_reg[18]/NET0131 ,
		\u13_icc_r_reg[19]/NET0131 ,
		\u1_slt6_reg[13]/P0001 ,
		_w4076_
	);
	LUT3 #(
		.INIT('he2)
	) name1930 (
		\u11_mem_reg[1][25]/P0001 ,
		_w4063_,
		_w4076_,
		_w4077_
	);
	LUT3 #(
		.INIT('h10)
	) name1931 (
		\u13_icc_r_reg[18]/NET0131 ,
		\u13_icc_r_reg[19]/NET0131 ,
		\u1_slt6_reg[14]/P0001 ,
		_w4078_
	);
	LUT3 #(
		.INIT('he2)
	) name1932 (
		\u11_mem_reg[1][26]/P0001 ,
		_w4063_,
		_w4078_,
		_w4079_
	);
	LUT3 #(
		.INIT('h10)
	) name1933 (
		\u13_icc_r_reg[18]/NET0131 ,
		\u13_icc_r_reg[19]/NET0131 ,
		\u1_slt6_reg[15]/P0001 ,
		_w4080_
	);
	LUT3 #(
		.INIT('he2)
	) name1934 (
		\u11_mem_reg[1][27]/P0001 ,
		_w4063_,
		_w4080_,
		_w4081_
	);
	LUT3 #(
		.INIT('h10)
	) name1935 (
		\u13_icc_r_reg[18]/NET0131 ,
		\u13_icc_r_reg[19]/NET0131 ,
		\u1_slt6_reg[16]/P0001 ,
		_w4082_
	);
	LUT3 #(
		.INIT('he2)
	) name1936 (
		\u11_mem_reg[1][28]/P0001 ,
		_w4063_,
		_w4082_,
		_w4083_
	);
	LUT3 #(
		.INIT('h10)
	) name1937 (
		\u13_icc_r_reg[18]/NET0131 ,
		\u13_icc_r_reg[19]/NET0131 ,
		\u1_slt6_reg[17]/P0001 ,
		_w4084_
	);
	LUT3 #(
		.INIT('he2)
	) name1938 (
		\u11_mem_reg[1][29]/P0001 ,
		_w4063_,
		_w4084_,
		_w4085_
	);
	LUT3 #(
		.INIT('h10)
	) name1939 (
		\u13_icc_r_reg[18]/NET0131 ,
		\u13_icc_r_reg[19]/NET0131 ,
		\u1_slt6_reg[18]/P0001 ,
		_w4086_
	);
	LUT3 #(
		.INIT('he2)
	) name1940 (
		\u11_mem_reg[1][30]/P0001 ,
		_w4063_,
		_w4086_,
		_w4087_
	);
	LUT3 #(
		.INIT('h10)
	) name1941 (
		\u13_icc_r_reg[18]/NET0131 ,
		\u13_icc_r_reg[19]/NET0131 ,
		\u1_slt6_reg[19]/P0001 ,
		_w4088_
	);
	LUT3 #(
		.INIT('he2)
	) name1942 (
		\u11_mem_reg[1][31]/P0001 ,
		_w4063_,
		_w4088_,
		_w4089_
	);
	LUT2 #(
		.INIT('h4)
	) name1943 (
		\u11_wp_reg[1]/P0001 ,
		\u11_wp_reg[2]/P0001 ,
		_w4090_
	);
	LUT3 #(
		.INIT('h20)
	) name1944 (
		_w2565_,
		_w2567_,
		_w4090_,
		_w4091_
	);
	LUT4 #(
		.INIT('ha2aa)
	) name1945 (
		\u11_mem_reg[2][18]/P0001 ,
		_w2565_,
		_w2567_,
		_w4090_,
		_w4092_
	);
	LUT4 #(
		.INIT('h0200)
	) name1946 (
		_w2565_,
		_w2567_,
		_w4052_,
		_w4090_,
		_w4093_
	);
	LUT2 #(
		.INIT('he)
	) name1947 (
		_w4092_,
		_w4093_,
		_w4094_
	);
	LUT4 #(
		.INIT('ha2aa)
	) name1948 (
		\u11_mem_reg[2][19]/P0001 ,
		_w2565_,
		_w2567_,
		_w4090_,
		_w4095_
	);
	LUT4 #(
		.INIT('h0200)
	) name1949 (
		_w2565_,
		_w2567_,
		_w4056_,
		_w4090_,
		_w4096_
	);
	LUT2 #(
		.INIT('he)
	) name1950 (
		_w4095_,
		_w4096_,
		_w4097_
	);
	LUT4 #(
		.INIT('ha2aa)
	) name1951 (
		\u11_mem_reg[2][20]/P0001 ,
		_w2565_,
		_w2567_,
		_w4090_,
		_w4098_
	);
	LUT4 #(
		.INIT('h2000)
	) name1952 (
		_w2565_,
		_w2567_,
		_w4066_,
		_w4090_,
		_w4099_
	);
	LUT2 #(
		.INIT('he)
	) name1953 (
		_w4098_,
		_w4099_,
		_w4100_
	);
	LUT4 #(
		.INIT('ha2aa)
	) name1954 (
		\u11_mem_reg[2][21]/P0001 ,
		_w2565_,
		_w2567_,
		_w4090_,
		_w4101_
	);
	LUT4 #(
		.INIT('h2000)
	) name1955 (
		_w2565_,
		_w2567_,
		_w4068_,
		_w4090_,
		_w4102_
	);
	LUT2 #(
		.INIT('he)
	) name1956 (
		_w4101_,
		_w4102_,
		_w4103_
	);
	LUT4 #(
		.INIT('ha2aa)
	) name1957 (
		\u11_mem_reg[2][22]/P0001 ,
		_w2565_,
		_w2567_,
		_w4090_,
		_w4104_
	);
	LUT4 #(
		.INIT('h2000)
	) name1958 (
		_w2565_,
		_w2567_,
		_w4070_,
		_w4090_,
		_w4105_
	);
	LUT2 #(
		.INIT('he)
	) name1959 (
		_w4104_,
		_w4105_,
		_w4106_
	);
	LUT4 #(
		.INIT('ha2aa)
	) name1960 (
		\u11_mem_reg[2][23]/P0001 ,
		_w2565_,
		_w2567_,
		_w4090_,
		_w4107_
	);
	LUT4 #(
		.INIT('h2000)
	) name1961 (
		_w2565_,
		_w2567_,
		_w4072_,
		_w4090_,
		_w4108_
	);
	LUT2 #(
		.INIT('he)
	) name1962 (
		_w4107_,
		_w4108_,
		_w4109_
	);
	LUT4 #(
		.INIT('ha2aa)
	) name1963 (
		\u11_mem_reg[2][24]/P0001 ,
		_w2565_,
		_w2567_,
		_w4090_,
		_w4110_
	);
	LUT4 #(
		.INIT('h2000)
	) name1964 (
		_w2565_,
		_w2567_,
		_w4074_,
		_w4090_,
		_w4111_
	);
	LUT2 #(
		.INIT('he)
	) name1965 (
		_w4110_,
		_w4111_,
		_w4112_
	);
	LUT4 #(
		.INIT('ha2aa)
	) name1966 (
		\u11_mem_reg[2][25]/P0001 ,
		_w2565_,
		_w2567_,
		_w4090_,
		_w4113_
	);
	LUT4 #(
		.INIT('h2000)
	) name1967 (
		_w2565_,
		_w2567_,
		_w4076_,
		_w4090_,
		_w4114_
	);
	LUT2 #(
		.INIT('he)
	) name1968 (
		_w4113_,
		_w4114_,
		_w4115_
	);
	LUT4 #(
		.INIT('h0020)
	) name1969 (
		\u10_wp_reg[1]/P0001 ,
		\u10_wp_reg[2]/P0001 ,
		_w2792_,
		_w2794_,
		_w4116_
	);
	LUT3 #(
		.INIT('h3a)
	) name1970 (
		\u10_mem_reg[1][18]/P0001 ,
		_w3881_,
		_w4116_,
		_w4117_
	);
	LUT4 #(
		.INIT('ha2aa)
	) name1971 (
		\u11_mem_reg[2][26]/P0001 ,
		_w2565_,
		_w2567_,
		_w4090_,
		_w4118_
	);
	LUT4 #(
		.INIT('h2000)
	) name1972 (
		_w2565_,
		_w2567_,
		_w4078_,
		_w4090_,
		_w4119_
	);
	LUT2 #(
		.INIT('he)
	) name1973 (
		_w4118_,
		_w4119_,
		_w4120_
	);
	LUT4 #(
		.INIT('ha2aa)
	) name1974 (
		\u11_mem_reg[2][27]/P0001 ,
		_w2565_,
		_w2567_,
		_w4090_,
		_w4121_
	);
	LUT4 #(
		.INIT('h2000)
	) name1975 (
		_w2565_,
		_w2567_,
		_w4080_,
		_w4090_,
		_w4122_
	);
	LUT2 #(
		.INIT('he)
	) name1976 (
		_w4121_,
		_w4122_,
		_w4123_
	);
	LUT3 #(
		.INIT('h3a)
	) name1977 (
		\u10_mem_reg[1][19]/P0001 ,
		_w3885_,
		_w4116_,
		_w4124_
	);
	LUT4 #(
		.INIT('ha2aa)
	) name1978 (
		\u11_mem_reg[2][28]/P0001 ,
		_w2565_,
		_w2567_,
		_w4090_,
		_w4125_
	);
	LUT4 #(
		.INIT('h2000)
	) name1979 (
		_w2565_,
		_w2567_,
		_w4082_,
		_w4090_,
		_w4126_
	);
	LUT2 #(
		.INIT('he)
	) name1980 (
		_w4125_,
		_w4126_,
		_w4127_
	);
	LUT4 #(
		.INIT('ha2aa)
	) name1981 (
		\u11_mem_reg[2][29]/P0001 ,
		_w2565_,
		_w2567_,
		_w4090_,
		_w4128_
	);
	LUT4 #(
		.INIT('h2000)
	) name1982 (
		_w2565_,
		_w2567_,
		_w4084_,
		_w4090_,
		_w4129_
	);
	LUT2 #(
		.INIT('he)
	) name1983 (
		_w4128_,
		_w4129_,
		_w4130_
	);
	LUT4 #(
		.INIT('ha2aa)
	) name1984 (
		\u11_mem_reg[2][30]/P0001 ,
		_w2565_,
		_w2567_,
		_w4090_,
		_w4131_
	);
	LUT4 #(
		.INIT('h2000)
	) name1985 (
		_w2565_,
		_w2567_,
		_w4086_,
		_w4090_,
		_w4132_
	);
	LUT2 #(
		.INIT('he)
	) name1986 (
		_w4131_,
		_w4132_,
		_w4133_
	);
	LUT3 #(
		.INIT('hca)
	) name1987 (
		\u10_mem_reg[1][20]/P0001 ,
		_w3889_,
		_w4116_,
		_w4134_
	);
	LUT4 #(
		.INIT('ha2aa)
	) name1988 (
		\u11_mem_reg[2][31]/P0001 ,
		_w2565_,
		_w2567_,
		_w4090_,
		_w4135_
	);
	LUT4 #(
		.INIT('h2000)
	) name1989 (
		_w2565_,
		_w2567_,
		_w4088_,
		_w4090_,
		_w4136_
	);
	LUT2 #(
		.INIT('he)
	) name1990 (
		_w4135_,
		_w4136_,
		_w4137_
	);
	LUT3 #(
		.INIT('hca)
	) name1991 (
		\u10_mem_reg[1][21]/P0001 ,
		_w3893_,
		_w4116_,
		_w4138_
	);
	LUT3 #(
		.INIT('hca)
	) name1992 (
		\u10_mem_reg[1][22]/P0001 ,
		_w3897_,
		_w4116_,
		_w4139_
	);
	LUT3 #(
		.INIT('hca)
	) name1993 (
		\u10_mem_reg[1][23]/P0001 ,
		_w3901_,
		_w4116_,
		_w4140_
	);
	LUT3 #(
		.INIT('hca)
	) name1994 (
		\u10_mem_reg[1][24]/P0001 ,
		_w3915_,
		_w4116_,
		_w4141_
	);
	LUT3 #(
		.INIT('hca)
	) name1995 (
		\u10_mem_reg[1][25]/P0001 ,
		_w3919_,
		_w4116_,
		_w4142_
	);
	LUT3 #(
		.INIT('hca)
	) name1996 (
		\u10_mem_reg[1][26]/P0001 ,
		_w3923_,
		_w4116_,
		_w4143_
	);
	LUT3 #(
		.INIT('hca)
	) name1997 (
		\u10_mem_reg[1][27]/P0001 ,
		_w3927_,
		_w4116_,
		_w4144_
	);
	LUT3 #(
		.INIT('hca)
	) name1998 (
		\u10_mem_reg[1][28]/P0001 ,
		_w3931_,
		_w4116_,
		_w4145_
	);
	LUT3 #(
		.INIT('hca)
	) name1999 (
		\u10_mem_reg[1][29]/P0001 ,
		_w3942_,
		_w4116_,
		_w4146_
	);
	LUT3 #(
		.INIT('h2e)
	) name2000 (
		\u11_mem_reg[3][18]/P0001 ,
		_w2570_,
		_w4052_,
		_w4147_
	);
	LUT3 #(
		.INIT('h2e)
	) name2001 (
		\u11_mem_reg[3][19]/P0001 ,
		_w2570_,
		_w4056_,
		_w4148_
	);
	LUT3 #(
		.INIT('he2)
	) name2002 (
		\u11_mem_reg[3][20]/P0001 ,
		_w2570_,
		_w4066_,
		_w4149_
	);
	LUT3 #(
		.INIT('hca)
	) name2003 (
		\u10_mem_reg[1][30]/P0001 ,
		_w3966_,
		_w4116_,
		_w4150_
	);
	LUT3 #(
		.INIT('he2)
	) name2004 (
		\u11_mem_reg[3][21]/P0001 ,
		_w2570_,
		_w4068_,
		_w4151_
	);
	LUT3 #(
		.INIT('he2)
	) name2005 (
		\u11_mem_reg[3][22]/P0001 ,
		_w2570_,
		_w4070_,
		_w4152_
	);
	LUT3 #(
		.INIT('hca)
	) name2006 (
		\u10_mem_reg[1][31]/P0001 ,
		_w3970_,
		_w4116_,
		_w4153_
	);
	LUT3 #(
		.INIT('he2)
	) name2007 (
		\u11_mem_reg[3][23]/P0001 ,
		_w2570_,
		_w4072_,
		_w4154_
	);
	LUT3 #(
		.INIT('he2)
	) name2008 (
		\u11_mem_reg[3][24]/P0001 ,
		_w2570_,
		_w4074_,
		_w4155_
	);
	LUT3 #(
		.INIT('he2)
	) name2009 (
		\u11_mem_reg[3][25]/P0001 ,
		_w2570_,
		_w4076_,
		_w4156_
	);
	LUT3 #(
		.INIT('he2)
	) name2010 (
		\u11_mem_reg[3][26]/P0001 ,
		_w2570_,
		_w4078_,
		_w4157_
	);
	LUT3 #(
		.INIT('he2)
	) name2011 (
		\u11_mem_reg[3][27]/P0001 ,
		_w2570_,
		_w4080_,
		_w4158_
	);
	LUT3 #(
		.INIT('he2)
	) name2012 (
		\u11_mem_reg[3][28]/P0001 ,
		_w2570_,
		_w4082_,
		_w4159_
	);
	LUT3 #(
		.INIT('he2)
	) name2013 (
		\u11_mem_reg[3][29]/P0001 ,
		_w2570_,
		_w4084_,
		_w4160_
	);
	LUT3 #(
		.INIT('he2)
	) name2014 (
		\u11_mem_reg[3][30]/P0001 ,
		_w2570_,
		_w4086_,
		_w4161_
	);
	LUT3 #(
		.INIT('he2)
	) name2015 (
		\u11_mem_reg[3][31]/P0001 ,
		_w2570_,
		_w4088_,
		_w4162_
	);
	LUT4 #(
		.INIT('h5515)
	) name2016 (
		\u13_ints_r_reg[1]/NET0131 ,
		\u15_crac_wr_reg/NET0131 ,
		\u15_valid_r_reg/P0001 ,
		\valid_s_reg/NET0131 ,
		_w4163_
	);
	LUT2 #(
		.INIT('h1)
	) name2017 (
		_w2403_,
		_w4163_,
		_w4164_
	);
	LUT2 #(
		.INIT('h2)
	) name2018 (
		\wb_addr_i[5]_pad ,
		\wb_addr_i[6]_pad ,
		_w4165_
	);
	LUT4 #(
		.INIT('h0080)
	) name2019 (
		\wb_addr_i[3]_pad ,
		\wb_addr_i[4]_pad ,
		\wb_addr_i[5]_pad ,
		\wb_addr_i[6]_pad ,
		_w4166_
	);
	LUT3 #(
		.INIT('h01)
	) name2020 (
		\wb_addr_i[2]_pad ,
		\wb_addr_i[3]_pad ,
		\wb_addr_i[4]_pad ,
		_w4167_
	);
	LUT2 #(
		.INIT('h4)
	) name2021 (
		\wb_addr_i[5]_pad ,
		\wb_addr_i[6]_pad ,
		_w4168_
	);
	LUT3 #(
		.INIT('h15)
	) name2022 (
		_w4166_,
		_w4167_,
		_w4168_,
		_w4169_
	);
	LUT3 #(
		.INIT('h10)
	) name2023 (
		\wb_addr_i[2]_pad ,
		\wb_addr_i[3]_pad ,
		\wb_addr_i[4]_pad ,
		_w4170_
	);
	LUT4 #(
		.INIT('h0200)
	) name2024 (
		\u15_crac_din_reg[1]/NET0131 ,
		\wb_addr_i[2]_pad ,
		\wb_addr_i[3]_pad ,
		\wb_addr_i[4]_pad ,
		_w4171_
	);
	LUT4 #(
		.INIT('h0002)
	) name2025 (
		suspended_o_pad,
		\wb_addr_i[2]_pad ,
		\wb_addr_i[3]_pad ,
		\wb_addr_i[4]_pad ,
		_w4172_
	);
	LUT3 #(
		.INIT('h08)
	) name2026 (
		\wb_addr_i[2]_pad ,
		\wb_addr_i[3]_pad ,
		\wb_addr_i[4]_pad ,
		_w4173_
	);
	LUT4 #(
		.INIT('h0080)
	) name2027 (
		\u13_icc_r_reg[1]/NET0131 ,
		\wb_addr_i[2]_pad ,
		\wb_addr_i[3]_pad ,
		\wb_addr_i[4]_pad ,
		_w4174_
	);
	LUT3 #(
		.INIT('h01)
	) name2028 (
		_w4172_,
		_w4174_,
		_w4171_,
		_w4175_
	);
	LUT3 #(
		.INIT('h04)
	) name2029 (
		\wb_addr_i[2]_pad ,
		\wb_addr_i[3]_pad ,
		\wb_addr_i[4]_pad ,
		_w4176_
	);
	LUT4 #(
		.INIT('h0020)
	) name2030 (
		\u13_occ1_r_reg[1]/NET0131 ,
		\wb_addr_i[2]_pad ,
		\wb_addr_i[3]_pad ,
		\wb_addr_i[4]_pad ,
		_w4177_
	);
	LUT4 #(
		.INIT('h2000)
	) name2031 (
		\u13_ints_r_reg[1]/NET0131 ,
		\wb_addr_i[2]_pad ,
		\wb_addr_i[3]_pad ,
		\wb_addr_i[4]_pad ,
		_w4178_
	);
	LUT3 #(
		.INIT('h02)
	) name2032 (
		\wb_addr_i[2]_pad ,
		\wb_addr_i[3]_pad ,
		\wb_addr_i[4]_pad ,
		_w4179_
	);
	LUT4 #(
		.INIT('h0008)
	) name2033 (
		\u13_occ0_r_reg[1]/NET0131 ,
		\wb_addr_i[2]_pad ,
		\wb_addr_i[3]_pad ,
		\wb_addr_i[4]_pad ,
		_w4180_
	);
	LUT3 #(
		.INIT('h20)
	) name2034 (
		\wb_addr_i[2]_pad ,
		\wb_addr_i[3]_pad ,
		\wb_addr_i[4]_pad ,
		_w4181_
	);
	LUT4 #(
		.INIT('h0800)
	) name2035 (
		\u13_intm_r_reg[1]/NET0131 ,
		\wb_addr_i[2]_pad ,
		\wb_addr_i[3]_pad ,
		\wb_addr_i[4]_pad ,
		_w4182_
	);
	LUT4 #(
		.INIT('h0001)
	) name2036 (
		_w4177_,
		_w4178_,
		_w4180_,
		_w4182_,
		_w4183_
	);
	LUT3 #(
		.INIT('h2a)
	) name2037 (
		_w4169_,
		_w4175_,
		_w4183_,
		_w4184_
	);
	LUT3 #(
		.INIT('h80)
	) name2038 (
		\u11_dout_reg[1]/P0001 ,
		_w4167_,
		_w4168_,
		_w4185_
	);
	LUT4 #(
		.INIT('h53ff)
	) name2039 (
		\u10_dout_reg[1]/P0001 ,
		\u9_dout_reg[1]/P0001 ,
		\wb_addr_i[2]_pad ,
		_w4166_,
		_w4186_
	);
	LUT2 #(
		.INIT('h4)
	) name2040 (
		_w4185_,
		_w4186_,
		_w4187_
	);
	LUT2 #(
		.INIT('hb)
	) name2041 (
		_w4184_,
		_w4187_,
		_w4188_
	);
	LUT3 #(
		.INIT('h10)
	) name2042 (
		\u26_cnt_reg[0]/NET0131 ,
		\u26_cnt_reg[1]/NET0131 ,
		\u26_cnt_reg[2]/NET0131 ,
		_w4189_
	);
	LUT4 #(
		.INIT('h5515)
	) name2043 (
		\u26_cnt_reg[0]/NET0131 ,
		_w3862_,
		_w3863_,
		_w4189_,
		_w4190_
	);
	LUT3 #(
		.INIT('h80)
	) name2044 (
		\u26_cnt_reg[0]/NET0131 ,
		_w3862_,
		_w3863_,
		_w4191_
	);
	LUT4 #(
		.INIT('h1555)
	) name2045 (
		\u13_ac97_rst_force_reg/P0001 ,
		\u26_cnt_reg[0]/NET0131 ,
		_w3862_,
		_w3863_,
		_w4192_
	);
	LUT2 #(
		.INIT('h4)
	) name2046 (
		_w4190_,
		_w4192_,
		_w4193_
	);
	LUT4 #(
		.INIT('h8000)
	) name2047 (
		\u26_cnt_reg[0]/NET0131 ,
		\u26_cnt_reg[1]/NET0131 ,
		_w3862_,
		_w3863_,
		_w4194_
	);
	LUT3 #(
		.INIT('h14)
	) name2048 (
		\u13_ac97_rst_force_reg/P0001 ,
		\u26_cnt_reg[1]/NET0131 ,
		_w4191_,
		_w4195_
	);
	LUT3 #(
		.INIT('h14)
	) name2049 (
		\u13_ac97_rst_force_reg/P0001 ,
		\u26_cnt_reg[2]/NET0131 ,
		_w4194_,
		_w4196_
	);
	LUT4 #(
		.INIT('h4000)
	) name2050 (
		\u14_u0_en_out_l2_reg/P0001 ,
		\u14_u0_en_out_l_reg/NET0131 ,
		\u3_empty_reg/NET0131 ,
		\valid_s_reg/NET0131 ,
		_w4197_
	);
	LUT2 #(
		.INIT('he)
	) name2051 (
		\u17_int_set_reg[1]/NET0131 ,
		_w4197_,
		_w4198_
	);
	LUT4 #(
		.INIT('h4000)
	) name2052 (
		\u14_u1_en_out_l2_reg/P0001 ,
		\u14_u1_en_out_l_reg/NET0131 ,
		\u4_empty_reg/NET0131 ,
		\valid_s_reg/NET0131 ,
		_w4199_
	);
	LUT2 #(
		.INIT('he)
	) name2053 (
		\u18_int_set_reg[1]/NET0131 ,
		_w4199_,
		_w4200_
	);
	LUT4 #(
		.INIT('h4000)
	) name2054 (
		\u14_u2_en_out_l2_reg/P0001 ,
		\u14_u2_en_out_l_reg/NET0131 ,
		\u5_empty_reg/NET0131 ,
		\valid_s_reg/NET0131 ,
		_w4201_
	);
	LUT2 #(
		.INIT('he)
	) name2055 (
		\u19_int_set_reg[1]/NET0131 ,
		_w4201_,
		_w4202_
	);
	LUT4 #(
		.INIT('h4000)
	) name2056 (
		\u14_u3_en_out_l2_reg/P0001 ,
		\u14_u3_en_out_l_reg/NET0131 ,
		\u6_empty_reg/NET0131 ,
		\valid_s_reg/NET0131 ,
		_w4203_
	);
	LUT2 #(
		.INIT('he)
	) name2057 (
		\u20_int_set_reg[1]/NET0131 ,
		_w4203_,
		_w4204_
	);
	LUT4 #(
		.INIT('h4000)
	) name2058 (
		\u14_u4_en_out_l2_reg/P0001 ,
		\u14_u4_en_out_l_reg/NET0131 ,
		\u7_empty_reg/NET0131 ,
		\valid_s_reg/NET0131 ,
		_w4205_
	);
	LUT2 #(
		.INIT('he)
	) name2059 (
		\u21_int_set_reg[1]/NET0131 ,
		_w4205_,
		_w4206_
	);
	LUT4 #(
		.INIT('h4000)
	) name2060 (
		\u14_u5_en_out_l2_reg/P0001 ,
		\u14_u5_en_out_l_reg/NET0131 ,
		\u8_empty_reg/NET0131 ,
		\valid_s_reg/NET0131 ,
		_w4207_
	);
	LUT2 #(
		.INIT('he)
	) name2061 (
		\u22_int_set_reg[1]/NET0131 ,
		_w4207_,
		_w4208_
	);
	LUT4 #(
		.INIT('h2000)
	) name2062 (
		\in_valid_s_reg[0]/NET0131 ,
		\u14_u6_en_out_l2_reg/P0001 ,
		\u14_u6_en_out_l_reg/NET0131 ,
		\u9_full_reg/NET0131 ,
		_w4209_
	);
	LUT2 #(
		.INIT('he)
	) name2063 (
		\u23_int_set_reg[2]/NET0131 ,
		_w4209_,
		_w4210_
	);
	LUT4 #(
		.INIT('h0800)
	) name2064 (
		\in_valid_s_reg[1]/NET0131 ,
		\u10_full_reg/NET0131 ,
		\u14_u7_en_out_l2_reg/P0001 ,
		\u14_u7_en_out_l_reg/NET0131 ,
		_w4211_
	);
	LUT2 #(
		.INIT('he)
	) name2065 (
		\u24_int_set_reg[2]/NET0131 ,
		_w4211_,
		_w4212_
	);
	LUT4 #(
		.INIT('h0800)
	) name2066 (
		\in_valid_s_reg[2]/NET0131 ,
		\u11_full_reg/NET0131 ,
		\u14_u8_en_out_l2_reg/P0001 ,
		\u14_u8_en_out_l_reg/NET0131 ,
		_w4213_
	);
	LUT2 #(
		.INIT('he)
	) name2067 (
		\u25_int_set_reg[2]/NET0131 ,
		_w4213_,
		_w4214_
	);
	LUT4 #(
		.INIT('h5455)
	) name2068 (
		\ac97_reset_pad_o__pad ,
		\u26_cnt_reg[0]/NET0131 ,
		\u26_cnt_reg[1]/NET0131 ,
		\u26_cnt_reg[2]/NET0131 ,
		_w4215_
	);
	LUT2 #(
		.INIT('h1)
	) name2069 (
		\u13_ac97_rst_force_reg/P0001 ,
		_w4215_,
		_w4216_
	);
	LUT2 #(
		.INIT('h4)
	) name2070 (
		\u13_crac_r_reg[7]/NET0131 ,
		\u15_crac_we_r_reg/P0001 ,
		_w4217_
	);
	LUT3 #(
		.INIT('ha2)
	) name2071 (
		\u15_crac_wr_reg/NET0131 ,
		\u15_valid_r_reg/P0001 ,
		\valid_s_reg/NET0131 ,
		_w4218_
	);
	LUT2 #(
		.INIT('he)
	) name2072 (
		_w4217_,
		_w4218_,
		_w4219_
	);
	LUT2 #(
		.INIT('h8)
	) name2073 (
		\u13_crac_r_reg[7]/NET0131 ,
		\u15_crac_we_r_reg/P0001 ,
		_w4220_
	);
	LUT4 #(
		.INIT('ha2aa)
	) name2074 (
		\u15_crac_rd_reg/NET0131 ,
		\u15_rdd1_reg/NET0131 ,
		\u15_valid_r_reg/P0001 ,
		\valid_s_reg/NET0131 ,
		_w4221_
	);
	LUT2 #(
		.INIT('he)
	) name2075 (
		_w4220_,
		_w4221_,
		_w4222_
	);
	LUT3 #(
		.INIT('he2)
	) name2076 (
		\u0_slt9_r_reg[1]/P0001 ,
		\u2_ld_reg/P0001 ,
		\u8_dout_reg[2]/P0001 ,
		_w4223_
	);
	LUT4 #(
		.INIT('h8c23)
	) name2077 (
		\u3_rp_reg[1]/NET0131 ,
		\u3_rp_reg[2]/NET0131 ,
		\u3_wp_reg[0]/P0001 ,
		\u3_wp_reg[1]/NET0131 ,
		_w4224_
	);
	LUT2 #(
		.INIT('h6)
	) name2078 (
		\u3_rp_reg[3]/NET0131 ,
		\u3_wp_reg[2]/P0001 ,
		_w4225_
	);
	LUT3 #(
		.INIT('ha2)
	) name2079 (
		\u12_o3_we_reg/P0001 ,
		\u3_rp_reg[1]/NET0131 ,
		\u3_wp_reg[0]/P0001 ,
		_w4226_
	);
	LUT4 #(
		.INIT('heaaa)
	) name2080 (
		\u17_int_set_reg[2]/NET0131 ,
		_w4225_,
		_w4224_,
		_w4226_,
		_w4227_
	);
	LUT4 #(
		.INIT('h8c23)
	) name2081 (
		\u4_rp_reg[1]/NET0131 ,
		\u4_rp_reg[2]/NET0131 ,
		\u4_wp_reg[0]/P0001 ,
		\u4_wp_reg[1]/NET0131 ,
		_w4228_
	);
	LUT2 #(
		.INIT('h6)
	) name2082 (
		\u4_rp_reg[3]/NET0131 ,
		\u4_wp_reg[2]/P0001 ,
		_w4229_
	);
	LUT3 #(
		.INIT('ha2)
	) name2083 (
		\u12_o4_we_reg/P0001 ,
		\u4_rp_reg[1]/NET0131 ,
		\u4_wp_reg[0]/P0001 ,
		_w4230_
	);
	LUT4 #(
		.INIT('heaaa)
	) name2084 (
		\u18_int_set_reg[2]/NET0131 ,
		_w4228_,
		_w4229_,
		_w4230_,
		_w4231_
	);
	LUT4 #(
		.INIT('h8c23)
	) name2085 (
		\u5_rp_reg[1]/NET0131 ,
		\u5_rp_reg[2]/NET0131 ,
		\u5_wp_reg[0]/P0001 ,
		\u5_wp_reg[1]/NET0131 ,
		_w4232_
	);
	LUT2 #(
		.INIT('h6)
	) name2086 (
		\u5_rp_reg[3]/NET0131 ,
		\u5_wp_reg[2]/P0001 ,
		_w4233_
	);
	LUT3 #(
		.INIT('ha2)
	) name2087 (
		\u12_o6_we_reg/P0001 ,
		\u5_rp_reg[1]/NET0131 ,
		\u5_wp_reg[0]/P0001 ,
		_w4234_
	);
	LUT4 #(
		.INIT('heaaa)
	) name2088 (
		\u19_int_set_reg[2]/NET0131 ,
		_w4232_,
		_w4233_,
		_w4234_,
		_w4235_
	);
	LUT2 #(
		.INIT('h9)
	) name2089 (
		\u6_rp_reg[1]/NET0131 ,
		\u6_wp_reg[0]/P0001 ,
		_w4236_
	);
	LUT4 #(
		.INIT('h8421)
	) name2090 (
		\u6_rp_reg[1]/NET0131 ,
		\u6_rp_reg[2]/NET0131 ,
		\u6_wp_reg[0]/P0001 ,
		\u6_wp_reg[1]/NET0131 ,
		_w4237_
	);
	LUT2 #(
		.INIT('h6)
	) name2091 (
		\u6_rp_reg[3]/NET0131 ,
		\u6_wp_reg[2]/P0001 ,
		_w4238_
	);
	LUT3 #(
		.INIT('h28)
	) name2092 (
		\u12_o7_we_reg/P0001 ,
		\u6_rp_reg[3]/NET0131 ,
		\u6_wp_reg[2]/P0001 ,
		_w4239_
	);
	LUT3 #(
		.INIT('hea)
	) name2093 (
		\u20_int_set_reg[2]/NET0131 ,
		_w4237_,
		_w4239_,
		_w4240_
	);
	LUT4 #(
		.INIT('h8c23)
	) name2094 (
		\u7_rp_reg[1]/NET0131 ,
		\u7_rp_reg[2]/NET0131 ,
		\u7_wp_reg[0]/P0001 ,
		\u7_wp_reg[1]/NET0131 ,
		_w4241_
	);
	LUT2 #(
		.INIT('h6)
	) name2095 (
		\u7_rp_reg[3]/NET0131 ,
		\u7_wp_reg[2]/P0001 ,
		_w4242_
	);
	LUT3 #(
		.INIT('ha2)
	) name2096 (
		\u12_o8_we_reg/P0001 ,
		\u7_rp_reg[1]/NET0131 ,
		\u7_wp_reg[0]/P0001 ,
		_w4243_
	);
	LUT4 #(
		.INIT('heaaa)
	) name2097 (
		\u21_int_set_reg[2]/NET0131 ,
		_w4242_,
		_w4241_,
		_w4243_,
		_w4244_
	);
	LUT2 #(
		.INIT('h9)
	) name2098 (
		\u8_rp_reg[1]/NET0131 ,
		\u8_wp_reg[0]/P0001 ,
		_w4245_
	);
	LUT4 #(
		.INIT('h8421)
	) name2099 (
		\u8_rp_reg[1]/NET0131 ,
		\u8_rp_reg[2]/NET0131 ,
		\u8_wp_reg[0]/P0001 ,
		\u8_wp_reg[1]/NET0131 ,
		_w4246_
	);
	LUT2 #(
		.INIT('h6)
	) name2100 (
		\u8_rp_reg[3]/NET0131 ,
		\u8_wp_reg[2]/P0001 ,
		_w4247_
	);
	LUT3 #(
		.INIT('h28)
	) name2101 (
		\u12_o9_we_reg/P0001 ,
		\u8_rp_reg[3]/NET0131 ,
		\u8_wp_reg[2]/P0001 ,
		_w4248_
	);
	LUT3 #(
		.INIT('hea)
	) name2102 (
		\u22_int_set_reg[2]/NET0131 ,
		_w4246_,
		_w4248_,
		_w4249_
	);
	LUT3 #(
		.INIT('h80)
	) name2103 (
		\u12_o9_we_reg/P0001 ,
		\u8_wp_reg[0]/P0001 ,
		\u8_wp_reg[1]/NET0131 ,
		_w4250_
	);
	LUT3 #(
		.INIT('h28)
	) name2104 (
		\u13_occ1_r_reg[8]/NET0131 ,
		\u8_wp_reg[2]/P0001 ,
		_w4250_,
		_w4251_
	);
	LUT3 #(
		.INIT('h80)
	) name2105 (
		\u12_o4_we_reg/P0001 ,
		\u4_wp_reg[0]/P0001 ,
		\u4_wp_reg[1]/NET0131 ,
		_w4252_
	);
	LUT3 #(
		.INIT('h28)
	) name2106 (
		\u13_occ0_r_reg[8]/NET0131 ,
		\u4_wp_reg[2]/P0001 ,
		_w4252_,
		_w4253_
	);
	LUT3 #(
		.INIT('h80)
	) name2107 (
		\u12_o6_we_reg/P0001 ,
		\u5_wp_reg[0]/P0001 ,
		\u5_wp_reg[1]/NET0131 ,
		_w4254_
	);
	LUT3 #(
		.INIT('h28)
	) name2108 (
		\u13_occ0_r_reg[16]/NET0131 ,
		\u5_wp_reg[2]/P0001 ,
		_w4254_,
		_w4255_
	);
	LUT3 #(
		.INIT('h80)
	) name2109 (
		\u12_o3_we_reg/P0001 ,
		\u3_wp_reg[0]/P0001 ,
		\u3_wp_reg[1]/NET0131 ,
		_w4256_
	);
	LUT3 #(
		.INIT('h28)
	) name2110 (
		\u13_occ0_r_reg[0]/NET0131 ,
		\u3_wp_reg[2]/P0001 ,
		_w4256_,
		_w4257_
	);
	LUT3 #(
		.INIT('h80)
	) name2111 (
		\u12_o7_we_reg/P0001 ,
		\u6_wp_reg[0]/P0001 ,
		\u6_wp_reg[1]/NET0131 ,
		_w4258_
	);
	LUT3 #(
		.INIT('h28)
	) name2112 (
		\u13_occ0_r_reg[24]/NET0131 ,
		\u6_wp_reg[2]/P0001 ,
		_w4258_,
		_w4259_
	);
	LUT3 #(
		.INIT('h80)
	) name2113 (
		\u12_o8_we_reg/P0001 ,
		\u7_wp_reg[0]/P0001 ,
		\u7_wp_reg[1]/NET0131 ,
		_w4260_
	);
	LUT3 #(
		.INIT('h28)
	) name2114 (
		\u13_occ1_r_reg[0]/NET0131 ,
		\u7_wp_reg[2]/P0001 ,
		_w4260_,
		_w4261_
	);
	LUT4 #(
		.INIT('h0200)
	) name2115 (
		\in_valid_s_reg[2]/NET0131 ,
		\u11_wp_reg[0]/NET0131 ,
		\u14_u8_en_out_l2_reg/P0001 ,
		\u14_u8_en_out_l_reg/NET0131 ,
		_w4262_
	);
	LUT4 #(
		.INIT('h0020)
	) name2116 (
		\in_valid_s_reg[0]/NET0131 ,
		\u14_u6_en_out_l2_reg/P0001 ,
		\u14_u6_en_out_l_reg/NET0131 ,
		\u9_wp_reg[0]/NET0131 ,
		_w4263_
	);
	LUT4 #(
		.INIT('h0200)
	) name2117 (
		\in_valid_s_reg[1]/NET0131 ,
		\u10_wp_reg[0]/NET0131 ,
		\u14_u7_en_out_l2_reg/P0001 ,
		\u14_u7_en_out_l_reg/NET0131 ,
		_w4264_
	);
	LUT2 #(
		.INIT('h8)
	) name2118 (
		\u14_u0_en_out_l_reg/NET0131 ,
		\valid_s_reg/NET0131 ,
		_w4265_
	);
	LUT3 #(
		.INIT('h20)
	) name2119 (
		\u13_occ0_r_reg[0]/NET0131 ,
		\u14_u0_full_empty_r_reg/P0001 ,
		\u1_slt0_reg[15]/P0001 ,
		_w4266_
	);
	LUT4 #(
		.INIT('h5f4c)
	) name2120 (
		\u13_occ0_r_reg[1]/NET0131 ,
		\u14_u0_en_out_l_reg/NET0131 ,
		\u1_slt1_reg[11]/P0001 ,
		\valid_s_reg/NET0131 ,
		_w4267_
	);
	LUT3 #(
		.INIT('hea)
	) name2121 (
		_w4265_,
		_w4266_,
		_w4267_,
		_w4268_
	);
	LUT3 #(
		.INIT('h20)
	) name2122 (
		\u13_occ0_r_reg[8]/NET0131 ,
		\u14_u1_full_empty_r_reg/P0001 ,
		\u1_slt0_reg[15]/P0001 ,
		_w4269_
	);
	LUT4 #(
		.INIT('h5f4c)
	) name2123 (
		\u13_occ0_r_reg[9]/NET0131 ,
		\u14_u1_en_out_l_reg/NET0131 ,
		\u1_slt1_reg[10]/P0001 ,
		\valid_s_reg/NET0131 ,
		_w4270_
	);
	LUT3 #(
		.INIT('hea)
	) name2124 (
		_w2416_,
		_w4269_,
		_w4270_,
		_w4271_
	);
	LUT3 #(
		.INIT('h20)
	) name2125 (
		\u13_occ0_r_reg[16]/NET0131 ,
		\u14_u2_full_empty_r_reg/P0001 ,
		\u1_slt0_reg[15]/P0001 ,
		_w4272_
	);
	LUT4 #(
		.INIT('h5f4c)
	) name2126 (
		\u13_occ0_r_reg[17]/NET0131 ,
		\u14_u2_en_out_l_reg/NET0131 ,
		\u1_slt1_reg[8]/P0001 ,
		\valid_s_reg/NET0131 ,
		_w4273_
	);
	LUT3 #(
		.INIT('hea)
	) name2127 (
		_w2425_,
		_w4272_,
		_w4273_,
		_w4274_
	);
	LUT3 #(
		.INIT('h20)
	) name2128 (
		\u13_occ0_r_reg[24]/NET0131 ,
		\u14_u3_full_empty_r_reg/P0001 ,
		\u1_slt0_reg[15]/P0001 ,
		_w4275_
	);
	LUT4 #(
		.INIT('h5f4c)
	) name2129 (
		\u13_occ0_r_reg[25]/NET0131 ,
		\u14_u3_en_out_l_reg/NET0131 ,
		\u1_slt1_reg[7]/P0001 ,
		\valid_s_reg/NET0131 ,
		_w4276_
	);
	LUT3 #(
		.INIT('hea)
	) name2130 (
		_w2443_,
		_w4275_,
		_w4276_,
		_w4277_
	);
	LUT3 #(
		.INIT('h20)
	) name2131 (
		\u13_occ1_r_reg[0]/NET0131 ,
		\u14_u4_full_empty_r_reg/P0001 ,
		\u1_slt0_reg[15]/P0001 ,
		_w4278_
	);
	LUT4 #(
		.INIT('h5f4c)
	) name2132 (
		\u13_occ1_r_reg[1]/NET0131 ,
		\u14_u4_en_out_l_reg/NET0131 ,
		\u1_slt1_reg[6]/P0001 ,
		\valid_s_reg/NET0131 ,
		_w4279_
	);
	LUT3 #(
		.INIT('hea)
	) name2133 (
		_w2454_,
		_w4278_,
		_w4279_,
		_w4280_
	);
	LUT3 #(
		.INIT('h20)
	) name2134 (
		\u13_occ1_r_reg[8]/NET0131 ,
		\u14_u5_full_empty_r_reg/P0001 ,
		\u1_slt0_reg[15]/P0001 ,
		_w4281_
	);
	LUT4 #(
		.INIT('h5f4c)
	) name2135 (
		\u13_occ1_r_reg[9]/NET0131 ,
		\u14_u5_en_out_l_reg/NET0131 ,
		\u1_slt1_reg[5]/P0001 ,
		\valid_s_reg/NET0131 ,
		_w4282_
	);
	LUT3 #(
		.INIT('hea)
	) name2136 (
		_w2154_,
		_w4281_,
		_w4282_,
		_w4283_
	);
	LUT3 #(
		.INIT('h20)
	) name2137 (
		\u13_icc_r_reg[0]/NET0131 ,
		\u14_u6_full_empty_r_reg/P0001 ,
		\u1_slt0_reg[15]/P0001 ,
		_w4284_
	);
	LUT4 #(
		.INIT('hfa32)
	) name2138 (
		\in_valid_s_reg[0]/NET0131 ,
		\u13_icc_r_reg[1]/NET0131 ,
		\u14_u6_en_out_l_reg/NET0131 ,
		\u1_slt0_reg[12]/P0001 ,
		_w4285_
	);
	LUT3 #(
		.INIT('hea)
	) name2139 (
		_w2685_,
		_w4284_,
		_w4285_,
		_w4286_
	);
	LUT3 #(
		.INIT('h20)
	) name2140 (
		\u13_icc_r_reg[8]/NET0131 ,
		\u14_u7_full_empty_r_reg/P0001 ,
		\u1_slt0_reg[15]/P0001 ,
		_w4287_
	);
	LUT4 #(
		.INIT('hfa32)
	) name2141 (
		\in_valid_s_reg[1]/NET0131 ,
		\u13_icc_r_reg[9]/NET0131 ,
		\u14_u7_en_out_l_reg/NET0131 ,
		\u1_slt0_reg[11]/P0001 ,
		_w4288_
	);
	LUT3 #(
		.INIT('hea)
	) name2142 (
		_w2791_,
		_w4287_,
		_w4288_,
		_w4289_
	);
	LUT3 #(
		.INIT('h20)
	) name2143 (
		\u13_icc_r_reg[16]/NET0131 ,
		\u14_u8_full_empty_r_reg/P0001 ,
		\u1_slt0_reg[15]/P0001 ,
		_w4290_
	);
	LUT4 #(
		.INIT('hfa32)
	) name2144 (
		\in_valid_s_reg[2]/NET0131 ,
		\u13_icc_r_reg[17]/NET0131 ,
		\u14_u8_en_out_l_reg/NET0131 ,
		\u1_slt0_reg[9]/P0001 ,
		_w4291_
	);
	LUT3 #(
		.INIT('hea)
	) name2145 (
		_w2564_,
		_w4290_,
		_w4291_,
		_w4292_
	);
	LUT3 #(
		.INIT('h48)
	) name2146 (
		\u12_o9_we_reg/P0001 ,
		\u13_occ1_r_reg[8]/NET0131 ,
		\u8_wp_reg[0]/P0001 ,
		_w4293_
	);
	LUT3 #(
		.INIT('h48)
	) name2147 (
		\u12_o3_we_reg/P0001 ,
		\u13_occ0_r_reg[0]/NET0131 ,
		\u3_wp_reg[0]/P0001 ,
		_w4294_
	);
	LUT3 #(
		.INIT('h48)
	) name2148 (
		\u12_o4_we_reg/P0001 ,
		\u13_occ0_r_reg[8]/NET0131 ,
		\u4_wp_reg[0]/P0001 ,
		_w4295_
	);
	LUT3 #(
		.INIT('h48)
	) name2149 (
		\u12_o6_we_reg/P0001 ,
		\u13_occ0_r_reg[16]/NET0131 ,
		\u5_wp_reg[0]/P0001 ,
		_w4296_
	);
	LUT3 #(
		.INIT('h48)
	) name2150 (
		\u12_o7_we_reg/P0001 ,
		\u13_occ0_r_reg[24]/NET0131 ,
		\u6_wp_reg[0]/P0001 ,
		_w4297_
	);
	LUT3 #(
		.INIT('h48)
	) name2151 (
		\u12_o8_we_reg/P0001 ,
		\u13_occ1_r_reg[0]/NET0131 ,
		\u7_wp_reg[0]/P0001 ,
		_w4298_
	);
	LUT4 #(
		.INIT('h4c80)
	) name2152 (
		\u12_o9_we_reg/P0001 ,
		\u13_occ1_r_reg[8]/NET0131 ,
		\u8_wp_reg[0]/P0001 ,
		\u8_wp_reg[1]/NET0131 ,
		_w4299_
	);
	LUT4 #(
		.INIT('h4c80)
	) name2153 (
		\u12_o4_we_reg/P0001 ,
		\u13_occ0_r_reg[8]/NET0131 ,
		\u4_wp_reg[0]/P0001 ,
		\u4_wp_reg[1]/NET0131 ,
		_w4300_
	);
	LUT4 #(
		.INIT('h4c80)
	) name2154 (
		\u12_o6_we_reg/P0001 ,
		\u13_occ0_r_reg[16]/NET0131 ,
		\u5_wp_reg[0]/P0001 ,
		\u5_wp_reg[1]/NET0131 ,
		_w4301_
	);
	LUT4 #(
		.INIT('h4c80)
	) name2155 (
		\u12_o3_we_reg/P0001 ,
		\u13_occ0_r_reg[0]/NET0131 ,
		\u3_wp_reg[0]/P0001 ,
		\u3_wp_reg[1]/NET0131 ,
		_w4302_
	);
	LUT4 #(
		.INIT('h4c80)
	) name2156 (
		\u12_o7_we_reg/P0001 ,
		\u13_occ0_r_reg[24]/NET0131 ,
		\u6_wp_reg[0]/P0001 ,
		\u6_wp_reg[1]/NET0131 ,
		_w4303_
	);
	LUT4 #(
		.INIT('h4c80)
	) name2157 (
		\u12_o8_we_reg/P0001 ,
		\u13_occ1_r_reg[0]/NET0131 ,
		\u7_wp_reg[0]/P0001 ,
		\u7_wp_reg[1]/NET0131 ,
		_w4304_
	);
	LUT4 #(
		.INIT('h88a8)
	) name2158 (
		\u15_crac_rd_reg/NET0131 ,
		\u15_rdd1_reg/NET0131 ,
		\u15_valid_r_reg/P0001 ,
		\valid_s_reg/NET0131 ,
		_w4305_
	);
	LUT3 #(
		.INIT('h08)
	) name2159 (
		\u15_crac_rd_reg/NET0131 ,
		\u15_valid_r_reg/P0001 ,
		\valid_s_reg/NET0131 ,
		_w4306_
	);
	LUT3 #(
		.INIT('h4c)
	) name2160 (
		\u15_crac_rd_done_reg/P0001 ,
		\u15_rdd2_reg/NET0131 ,
		\u15_rdd3_reg/NET0131 ,
		_w4307_
	);
	LUT2 #(
		.INIT('he)
	) name2161 (
		_w4306_,
		_w4307_,
		_w4308_
	);
	LUT3 #(
		.INIT('h20)
	) name2162 (
		\u15_rdd2_reg/NET0131 ,
		\u15_valid_r_reg/P0001 ,
		\valid_s_reg/NET0131 ,
		_w4309_
	);
	LUT2 #(
		.INIT('h4)
	) name2163 (
		\u15_crac_rd_done_reg/P0001 ,
		\u15_rdd3_reg/NET0131 ,
		_w4310_
	);
	LUT2 #(
		.INIT('he)
	) name2164 (
		_w4309_,
		_w4310_,
		_w4311_
	);
	LUT3 #(
		.INIT('h80)
	) name2165 (
		\u2_res_cnt_reg[0]/P0001 ,
		_w3862_,
		_w3863_,
		_w4312_
	);
	LUT4 #(
		.INIT('h8000)
	) name2166 (
		\u2_res_cnt_reg[0]/P0001 ,
		\u2_res_cnt_reg[1]/P0001 ,
		_w3862_,
		_w3863_,
		_w4313_
	);
	LUT4 #(
		.INIT('h60c0)
	) name2167 (
		\u2_res_cnt_reg[2]/P0001 ,
		\u2_res_cnt_reg[3]/P0001 ,
		\u2_sync_resume_reg/NET0131 ,
		_w4313_,
		_w4314_
	);
	LUT4 #(
		.INIT('h0002)
	) name2168 (
		\u12_rf_we_reg/P0001 ,
		\wb_addr_i[2]_pad ,
		\wb_addr_i[3]_pad ,
		\wb_addr_i[4]_pad ,
		_w4315_
	);
	LUT2 #(
		.INIT('h8)
	) name2169 (
		\u12_dout_reg[0]/P0001 ,
		_w4315_,
		_w4316_
	);
	LUT2 #(
		.INIT('h8)
	) name2170 (
		\u12_dout_reg[1]/P0001 ,
		_w4315_,
		_w4317_
	);
	LUT4 #(
		.INIT('hfcaa)
	) name2171 (
		\u14_crac_valid_r_reg/P0001 ,
		\u15_crac_rd_reg/NET0131 ,
		\u15_crac_wr_reg/NET0131 ,
		\valid_s_reg/NET0131 ,
		_w4318_
	);
	LUT3 #(
		.INIT('h20)
	) name2172 (
		\u15_rdd3_reg/NET0131 ,
		\u15_valid_r_reg/P0001 ,
		\valid_s_reg/NET0131 ,
		_w4319_
	);
	LUT4 #(
		.INIT('h8000)
	) name2173 (
		\u2_cnt_reg[0]/NET0131 ,
		\u2_cnt_reg[1]/NET0131 ,
		\u2_cnt_reg[2]/NET0131 ,
		\u2_cnt_reg[3]/NET0131 ,
		_w4320_
	);
	LUT2 #(
		.INIT('h8)
	) name2174 (
		\u2_cnt_reg[5]/NET0131 ,
		\u2_cnt_reg[6]/NET0131 ,
		_w4321_
	);
	LUT3 #(
		.INIT('h80)
	) name2175 (
		\u2_cnt_reg[4]/NET0131 ,
		_w4320_,
		_w4321_,
		_w4322_
	);
	LUT3 #(
		.INIT('hbe)
	) name2176 (
		suspended_o_pad,
		\u2_cnt_reg[7]/NET0131 ,
		_w4322_,
		_w4323_
	);
	LUT3 #(
		.INIT('h80)
	) name2177 (
		\u2_to_cnt_reg[0]/NET0131 ,
		\u2_to_cnt_reg[1]/NET0131 ,
		\u2_to_cnt_reg[2]/NET0131 ,
		_w4324_
	);
	LUT4 #(
		.INIT('h8000)
	) name2178 (
		\u2_to_cnt_reg[0]/NET0131 ,
		\u2_to_cnt_reg[1]/NET0131 ,
		\u2_to_cnt_reg[2]/NET0131 ,
		\u2_to_cnt_reg[3]/NET0131 ,
		_w4325_
	);
	LUT3 #(
		.INIT('h14)
	) name2179 (
		\u2_bit_clk_e_reg/P0001 ,
		\u2_to_cnt_reg[3]/NET0131 ,
		_w4324_,
		_w4326_
	);
	LUT4 #(
		.INIT('hc4cc)
	) name2180 (
		\u12_o9_we_reg/P0001 ,
		\u8_mem_reg[2][5]/NET0131 ,
		\u8_wp_reg[0]/P0001 ,
		\u8_wp_reg[1]/NET0131 ,
		_w4327_
	);
	LUT4 #(
		.INIT('h0800)
	) name2181 (
		\u12_dout_reg[5]/P0001 ,
		\u12_o9_we_reg/P0001 ,
		\u8_wp_reg[0]/P0001 ,
		\u8_wp_reg[1]/NET0131 ,
		_w4328_
	);
	LUT2 #(
		.INIT('he)
	) name2182 (
		_w4327_,
		_w4328_,
		_w4329_
	);
	LUT4 #(
		.INIT('hcc4c)
	) name2183 (
		\u12_o3_we_reg/P0001 ,
		\u3_mem_reg[1][29]/NET0131 ,
		\u3_wp_reg[0]/P0001 ,
		\u3_wp_reg[1]/NET0131 ,
		_w4330_
	);
	LUT4 #(
		.INIT('h0080)
	) name2184 (
		\u12_dout_reg[29]/P0001 ,
		\u12_o3_we_reg/P0001 ,
		\u3_wp_reg[0]/P0001 ,
		\u3_wp_reg[1]/NET0131 ,
		_w4331_
	);
	LUT2 #(
		.INIT('he)
	) name2185 (
		_w4330_,
		_w4331_,
		_w4332_
	);
	LUT4 #(
		.INIT('hc4cc)
	) name2186 (
		\u12_o9_we_reg/P0001 ,
		\u8_mem_reg[2][6]/NET0131 ,
		\u8_wp_reg[0]/P0001 ,
		\u8_wp_reg[1]/NET0131 ,
		_w4333_
	);
	LUT4 #(
		.INIT('h0800)
	) name2187 (
		\u12_dout_reg[6]/P0001 ,
		\u12_o9_we_reg/P0001 ,
		\u8_wp_reg[0]/P0001 ,
		\u8_wp_reg[1]/NET0131 ,
		_w4334_
	);
	LUT2 #(
		.INIT('he)
	) name2188 (
		_w4333_,
		_w4334_,
		_w4335_
	);
	LUT4 #(
		.INIT('hc4cc)
	) name2189 (
		\u12_o9_we_reg/P0001 ,
		\u8_mem_reg[2][7]/NET0131 ,
		\u8_wp_reg[0]/P0001 ,
		\u8_wp_reg[1]/NET0131 ,
		_w4336_
	);
	LUT4 #(
		.INIT('h0800)
	) name2190 (
		\u12_dout_reg[7]/P0001 ,
		\u12_o9_we_reg/P0001 ,
		\u8_wp_reg[0]/P0001 ,
		\u8_wp_reg[1]/NET0131 ,
		_w4337_
	);
	LUT2 #(
		.INIT('he)
	) name2191 (
		_w4336_,
		_w4337_,
		_w4338_
	);
	LUT4 #(
		.INIT('hcc4c)
	) name2192 (
		\u12_o3_we_reg/P0001 ,
		\u3_mem_reg[1][2]/NET0131 ,
		\u3_wp_reg[0]/P0001 ,
		\u3_wp_reg[1]/NET0131 ,
		_w4339_
	);
	LUT4 #(
		.INIT('h0080)
	) name2193 (
		\u12_dout_reg[2]/P0001 ,
		\u12_o3_we_reg/P0001 ,
		\u3_wp_reg[0]/P0001 ,
		\u3_wp_reg[1]/NET0131 ,
		_w4340_
	);
	LUT2 #(
		.INIT('he)
	) name2194 (
		_w4339_,
		_w4340_,
		_w4341_
	);
	LUT4 #(
		.INIT('hc4cc)
	) name2195 (
		\u12_o9_we_reg/P0001 ,
		\u8_mem_reg[2][8]/NET0131 ,
		\u8_wp_reg[0]/P0001 ,
		\u8_wp_reg[1]/NET0131 ,
		_w4342_
	);
	LUT4 #(
		.INIT('h0800)
	) name2196 (
		\u12_dout_reg[8]/P0001 ,
		\u12_o9_we_reg/P0001 ,
		\u8_wp_reg[0]/P0001 ,
		\u8_wp_reg[1]/NET0131 ,
		_w4343_
	);
	LUT2 #(
		.INIT('he)
	) name2197 (
		_w4342_,
		_w4343_,
		_w4344_
	);
	LUT4 #(
		.INIT('hc4cc)
	) name2198 (
		\u12_o9_we_reg/P0001 ,
		\u8_mem_reg[2][9]/NET0131 ,
		\u8_wp_reg[0]/P0001 ,
		\u8_wp_reg[1]/NET0131 ,
		_w4345_
	);
	LUT4 #(
		.INIT('h0800)
	) name2199 (
		\u12_dout_reg[9]/P0001 ,
		\u12_o9_we_reg/P0001 ,
		\u8_wp_reg[0]/P0001 ,
		\u8_wp_reg[1]/NET0131 ,
		_w4346_
	);
	LUT2 #(
		.INIT('he)
	) name2200 (
		_w4345_,
		_w4346_,
		_w4347_
	);
	LUT4 #(
		.INIT('h4ccc)
	) name2201 (
		\u12_o9_we_reg/P0001 ,
		\u8_mem_reg[3][19]/NET0131 ,
		\u8_wp_reg[0]/P0001 ,
		\u8_wp_reg[1]/NET0131 ,
		_w4348_
	);
	LUT4 #(
		.INIT('h8000)
	) name2202 (
		\u12_dout_reg[19]/P0001 ,
		\u12_o9_we_reg/P0001 ,
		\u8_wp_reg[0]/P0001 ,
		\u8_wp_reg[1]/NET0131 ,
		_w4349_
	);
	LUT2 #(
		.INIT('he)
	) name2203 (
		_w4348_,
		_w4349_,
		_w4350_
	);
	LUT4 #(
		.INIT('h4ccc)
	) name2204 (
		\u12_o9_we_reg/P0001 ,
		\u8_mem_reg[3][0]/NET0131 ,
		\u8_wp_reg[0]/P0001 ,
		\u8_wp_reg[1]/NET0131 ,
		_w4351_
	);
	LUT4 #(
		.INIT('h8000)
	) name2205 (
		\u12_dout_reg[0]/P0001 ,
		\u12_o9_we_reg/P0001 ,
		\u8_wp_reg[0]/P0001 ,
		\u8_wp_reg[1]/NET0131 ,
		_w4352_
	);
	LUT2 #(
		.INIT('he)
	) name2206 (
		_w4351_,
		_w4352_,
		_w4353_
	);
	LUT4 #(
		.INIT('h4ccc)
	) name2207 (
		\u12_o9_we_reg/P0001 ,
		\u8_mem_reg[3][10]/NET0131 ,
		\u8_wp_reg[0]/P0001 ,
		\u8_wp_reg[1]/NET0131 ,
		_w4354_
	);
	LUT4 #(
		.INIT('h8000)
	) name2208 (
		\u12_dout_reg[10]/P0001 ,
		\u12_o9_we_reg/P0001 ,
		\u8_wp_reg[0]/P0001 ,
		\u8_wp_reg[1]/NET0131 ,
		_w4355_
	);
	LUT2 #(
		.INIT('he)
	) name2209 (
		_w4354_,
		_w4355_,
		_w4356_
	);
	LUT4 #(
		.INIT('hcc4c)
	) name2210 (
		\u12_o3_we_reg/P0001 ,
		\u3_mem_reg[1][31]/NET0131 ,
		\u3_wp_reg[0]/P0001 ,
		\u3_wp_reg[1]/NET0131 ,
		_w4357_
	);
	LUT4 #(
		.INIT('h0080)
	) name2211 (
		\u12_dout_reg[31]/P0001 ,
		\u12_o3_we_reg/P0001 ,
		\u3_wp_reg[0]/P0001 ,
		\u3_wp_reg[1]/NET0131 ,
		_w4358_
	);
	LUT2 #(
		.INIT('he)
	) name2212 (
		_w4357_,
		_w4358_,
		_w4359_
	);
	LUT4 #(
		.INIT('h4ccc)
	) name2213 (
		\u12_o9_we_reg/P0001 ,
		\u8_mem_reg[3][12]/NET0131 ,
		\u8_wp_reg[0]/P0001 ,
		\u8_wp_reg[1]/NET0131 ,
		_w4360_
	);
	LUT4 #(
		.INIT('h8000)
	) name2214 (
		\u12_dout_reg[12]/P0001 ,
		\u12_o9_we_reg/P0001 ,
		\u8_wp_reg[0]/P0001 ,
		\u8_wp_reg[1]/NET0131 ,
		_w4361_
	);
	LUT2 #(
		.INIT('he)
	) name2215 (
		_w4360_,
		_w4361_,
		_w4362_
	);
	LUT4 #(
		.INIT('hcc4c)
	) name2216 (
		\u12_o3_we_reg/P0001 ,
		\u3_mem_reg[1][3]/NET0131 ,
		\u3_wp_reg[0]/P0001 ,
		\u3_wp_reg[1]/NET0131 ,
		_w4363_
	);
	LUT4 #(
		.INIT('h0080)
	) name2217 (
		\u12_dout_reg[3]/P0001 ,
		\u12_o3_we_reg/P0001 ,
		\u3_wp_reg[0]/P0001 ,
		\u3_wp_reg[1]/NET0131 ,
		_w4364_
	);
	LUT2 #(
		.INIT('he)
	) name2218 (
		_w4363_,
		_w4364_,
		_w4365_
	);
	LUT4 #(
		.INIT('h4ccc)
	) name2219 (
		\u12_o9_we_reg/P0001 ,
		\u8_mem_reg[3][13]/NET0131 ,
		\u8_wp_reg[0]/P0001 ,
		\u8_wp_reg[1]/NET0131 ,
		_w4366_
	);
	LUT4 #(
		.INIT('h8000)
	) name2220 (
		\u12_dout_reg[13]/P0001 ,
		\u12_o9_we_reg/P0001 ,
		\u8_wp_reg[0]/P0001 ,
		\u8_wp_reg[1]/NET0131 ,
		_w4367_
	);
	LUT2 #(
		.INIT('he)
	) name2221 (
		_w4366_,
		_w4367_,
		_w4368_
	);
	LUT4 #(
		.INIT('h4ccc)
	) name2222 (
		\u12_o9_we_reg/P0001 ,
		\u8_mem_reg[3][14]/NET0131 ,
		\u8_wp_reg[0]/P0001 ,
		\u8_wp_reg[1]/NET0131 ,
		_w4369_
	);
	LUT4 #(
		.INIT('h8000)
	) name2223 (
		\u12_dout_reg[14]/P0001 ,
		\u12_o9_we_reg/P0001 ,
		\u8_wp_reg[0]/P0001 ,
		\u8_wp_reg[1]/NET0131 ,
		_w4370_
	);
	LUT2 #(
		.INIT('he)
	) name2224 (
		_w4369_,
		_w4370_,
		_w4371_
	);
	LUT4 #(
		.INIT('h4ccc)
	) name2225 (
		\u12_o9_we_reg/P0001 ,
		\u8_mem_reg[3][15]/NET0131 ,
		\u8_wp_reg[0]/P0001 ,
		\u8_wp_reg[1]/NET0131 ,
		_w4372_
	);
	LUT4 #(
		.INIT('h8000)
	) name2226 (
		\u12_dout_reg[15]/P0001 ,
		\u12_o9_we_reg/P0001 ,
		\u8_wp_reg[0]/P0001 ,
		\u8_wp_reg[1]/NET0131 ,
		_w4373_
	);
	LUT2 #(
		.INIT('he)
	) name2227 (
		_w4372_,
		_w4373_,
		_w4374_
	);
	LUT4 #(
		.INIT('hcc4c)
	) name2228 (
		\u12_o3_we_reg/P0001 ,
		\u3_mem_reg[1][4]/NET0131 ,
		\u3_wp_reg[0]/P0001 ,
		\u3_wp_reg[1]/NET0131 ,
		_w4375_
	);
	LUT4 #(
		.INIT('h0080)
	) name2229 (
		\u12_dout_reg[4]/P0001 ,
		\u12_o3_we_reg/P0001 ,
		\u3_wp_reg[0]/P0001 ,
		\u3_wp_reg[1]/NET0131 ,
		_w4376_
	);
	LUT2 #(
		.INIT('he)
	) name2230 (
		_w4375_,
		_w4376_,
		_w4377_
	);
	LUT4 #(
		.INIT('h4ccc)
	) name2231 (
		\u12_o9_we_reg/P0001 ,
		\u8_mem_reg[3][16]/NET0131 ,
		\u8_wp_reg[0]/P0001 ,
		\u8_wp_reg[1]/NET0131 ,
		_w4378_
	);
	LUT4 #(
		.INIT('h8000)
	) name2232 (
		\u12_dout_reg[16]/P0001 ,
		\u12_o9_we_reg/P0001 ,
		\u8_wp_reg[0]/P0001 ,
		\u8_wp_reg[1]/NET0131 ,
		_w4379_
	);
	LUT2 #(
		.INIT('he)
	) name2233 (
		_w4378_,
		_w4379_,
		_w4380_
	);
	LUT4 #(
		.INIT('hcc4c)
	) name2234 (
		\u12_o3_we_reg/P0001 ,
		\u3_mem_reg[1][5]/NET0131 ,
		\u3_wp_reg[0]/P0001 ,
		\u3_wp_reg[1]/NET0131 ,
		_w4381_
	);
	LUT4 #(
		.INIT('h0080)
	) name2235 (
		\u12_dout_reg[5]/P0001 ,
		\u12_o3_we_reg/P0001 ,
		\u3_wp_reg[0]/P0001 ,
		\u3_wp_reg[1]/NET0131 ,
		_w4382_
	);
	LUT2 #(
		.INIT('he)
	) name2236 (
		_w4381_,
		_w4382_,
		_w4383_
	);
	LUT4 #(
		.INIT('h4ccc)
	) name2237 (
		\u12_o9_we_reg/P0001 ,
		\u8_mem_reg[3][17]/NET0131 ,
		\u8_wp_reg[0]/P0001 ,
		\u8_wp_reg[1]/NET0131 ,
		_w4384_
	);
	LUT4 #(
		.INIT('h8000)
	) name2238 (
		\u12_dout_reg[17]/P0001 ,
		\u12_o9_we_reg/P0001 ,
		\u8_wp_reg[0]/P0001 ,
		\u8_wp_reg[1]/NET0131 ,
		_w4385_
	);
	LUT2 #(
		.INIT('he)
	) name2239 (
		_w4384_,
		_w4385_,
		_w4386_
	);
	LUT4 #(
		.INIT('h4ccc)
	) name2240 (
		\u12_o9_we_reg/P0001 ,
		\u8_mem_reg[3][18]/NET0131 ,
		\u8_wp_reg[0]/P0001 ,
		\u8_wp_reg[1]/NET0131 ,
		_w4387_
	);
	LUT4 #(
		.INIT('h8000)
	) name2241 (
		\u12_dout_reg[18]/P0001 ,
		\u12_o9_we_reg/P0001 ,
		\u8_wp_reg[0]/P0001 ,
		\u8_wp_reg[1]/NET0131 ,
		_w4388_
	);
	LUT2 #(
		.INIT('he)
	) name2242 (
		_w4387_,
		_w4388_,
		_w4389_
	);
	LUT4 #(
		.INIT('hcc4c)
	) name2243 (
		\u12_o3_we_reg/P0001 ,
		\u3_mem_reg[1][6]/NET0131 ,
		\u3_wp_reg[0]/P0001 ,
		\u3_wp_reg[1]/NET0131 ,
		_w4390_
	);
	LUT4 #(
		.INIT('h0080)
	) name2244 (
		\u12_dout_reg[6]/P0001 ,
		\u12_o3_we_reg/P0001 ,
		\u3_wp_reg[0]/P0001 ,
		\u3_wp_reg[1]/NET0131 ,
		_w4391_
	);
	LUT2 #(
		.INIT('he)
	) name2245 (
		_w4390_,
		_w4391_,
		_w4392_
	);
	LUT4 #(
		.INIT('h4ccc)
	) name2246 (
		\u12_o9_we_reg/P0001 ,
		\u8_mem_reg[3][1]/NET0131 ,
		\u8_wp_reg[0]/P0001 ,
		\u8_wp_reg[1]/NET0131 ,
		_w4393_
	);
	LUT4 #(
		.INIT('h8000)
	) name2247 (
		\u12_dout_reg[1]/P0001 ,
		\u12_o9_we_reg/P0001 ,
		\u8_wp_reg[0]/P0001 ,
		\u8_wp_reg[1]/NET0131 ,
		_w4394_
	);
	LUT2 #(
		.INIT('he)
	) name2248 (
		_w4393_,
		_w4394_,
		_w4395_
	);
	LUT4 #(
		.INIT('hcc4c)
	) name2249 (
		\u12_o3_we_reg/P0001 ,
		\u3_mem_reg[1][7]/NET0131 ,
		\u3_wp_reg[0]/P0001 ,
		\u3_wp_reg[1]/NET0131 ,
		_w4396_
	);
	LUT4 #(
		.INIT('h0080)
	) name2250 (
		\u12_dout_reg[7]/P0001 ,
		\u12_o3_we_reg/P0001 ,
		\u3_wp_reg[0]/P0001 ,
		\u3_wp_reg[1]/NET0131 ,
		_w4397_
	);
	LUT2 #(
		.INIT('he)
	) name2251 (
		_w4396_,
		_w4397_,
		_w4398_
	);
	LUT4 #(
		.INIT('h4ccc)
	) name2252 (
		\u12_o9_we_reg/P0001 ,
		\u8_mem_reg[3][20]/NET0131 ,
		\u8_wp_reg[0]/P0001 ,
		\u8_wp_reg[1]/NET0131 ,
		_w4399_
	);
	LUT4 #(
		.INIT('h8000)
	) name2253 (
		\u12_dout_reg[20]/P0001 ,
		\u12_o9_we_reg/P0001 ,
		\u8_wp_reg[0]/P0001 ,
		\u8_wp_reg[1]/NET0131 ,
		_w4400_
	);
	LUT2 #(
		.INIT('he)
	) name2254 (
		_w4399_,
		_w4400_,
		_w4401_
	);
	LUT4 #(
		.INIT('h4ccc)
	) name2255 (
		\u12_o9_we_reg/P0001 ,
		\u8_mem_reg[3][21]/NET0131 ,
		\u8_wp_reg[0]/P0001 ,
		\u8_wp_reg[1]/NET0131 ,
		_w4402_
	);
	LUT4 #(
		.INIT('h8000)
	) name2256 (
		\u12_dout_reg[21]/P0001 ,
		\u12_o9_we_reg/P0001 ,
		\u8_wp_reg[0]/P0001 ,
		\u8_wp_reg[1]/NET0131 ,
		_w4403_
	);
	LUT2 #(
		.INIT('he)
	) name2257 (
		_w4402_,
		_w4403_,
		_w4404_
	);
	LUT4 #(
		.INIT('hcc4c)
	) name2258 (
		\u12_o3_we_reg/P0001 ,
		\u3_mem_reg[1][8]/NET0131 ,
		\u3_wp_reg[0]/P0001 ,
		\u3_wp_reg[1]/NET0131 ,
		_w4405_
	);
	LUT4 #(
		.INIT('h0080)
	) name2259 (
		\u12_dout_reg[8]/P0001 ,
		\u12_o3_we_reg/P0001 ,
		\u3_wp_reg[0]/P0001 ,
		\u3_wp_reg[1]/NET0131 ,
		_w4406_
	);
	LUT2 #(
		.INIT('he)
	) name2260 (
		_w4405_,
		_w4406_,
		_w4407_
	);
	LUT4 #(
		.INIT('h4ccc)
	) name2261 (
		\u12_o9_we_reg/P0001 ,
		\u8_mem_reg[3][22]/NET0131 ,
		\u8_wp_reg[0]/P0001 ,
		\u8_wp_reg[1]/NET0131 ,
		_w4408_
	);
	LUT4 #(
		.INIT('h8000)
	) name2262 (
		\u12_dout_reg[22]/P0001 ,
		\u12_o9_we_reg/P0001 ,
		\u8_wp_reg[0]/P0001 ,
		\u8_wp_reg[1]/NET0131 ,
		_w4409_
	);
	LUT2 #(
		.INIT('he)
	) name2263 (
		_w4408_,
		_w4409_,
		_w4410_
	);
	LUT4 #(
		.INIT('h4ccc)
	) name2264 (
		\u12_o9_we_reg/P0001 ,
		\u8_mem_reg[3][23]/NET0131 ,
		\u8_wp_reg[0]/P0001 ,
		\u8_wp_reg[1]/NET0131 ,
		_w4411_
	);
	LUT4 #(
		.INIT('h8000)
	) name2265 (
		\u12_dout_reg[23]/P0001 ,
		\u12_o9_we_reg/P0001 ,
		\u8_wp_reg[0]/P0001 ,
		\u8_wp_reg[1]/NET0131 ,
		_w4412_
	);
	LUT2 #(
		.INIT('he)
	) name2266 (
		_w4411_,
		_w4412_,
		_w4413_
	);
	LUT4 #(
		.INIT('hcc4c)
	) name2267 (
		\u12_o3_we_reg/P0001 ,
		\u3_mem_reg[1][9]/NET0131 ,
		\u3_wp_reg[0]/P0001 ,
		\u3_wp_reg[1]/NET0131 ,
		_w4414_
	);
	LUT4 #(
		.INIT('h0080)
	) name2268 (
		\u12_dout_reg[9]/P0001 ,
		\u12_o3_we_reg/P0001 ,
		\u3_wp_reg[0]/P0001 ,
		\u3_wp_reg[1]/NET0131 ,
		_w4415_
	);
	LUT2 #(
		.INIT('he)
	) name2269 (
		_w4414_,
		_w4415_,
		_w4416_
	);
	LUT4 #(
		.INIT('h4ccc)
	) name2270 (
		\u12_o9_we_reg/P0001 ,
		\u8_mem_reg[3][24]/NET0131 ,
		\u8_wp_reg[0]/P0001 ,
		\u8_wp_reg[1]/NET0131 ,
		_w4417_
	);
	LUT4 #(
		.INIT('h8000)
	) name2271 (
		\u12_dout_reg[24]/P0001 ,
		\u12_o9_we_reg/P0001 ,
		\u8_wp_reg[0]/P0001 ,
		\u8_wp_reg[1]/NET0131 ,
		_w4418_
	);
	LUT2 #(
		.INIT('he)
	) name2272 (
		_w4417_,
		_w4418_,
		_w4419_
	);
	LUT4 #(
		.INIT('h4ccc)
	) name2273 (
		\u12_o9_we_reg/P0001 ,
		\u8_mem_reg[3][25]/NET0131 ,
		\u8_wp_reg[0]/P0001 ,
		\u8_wp_reg[1]/NET0131 ,
		_w4420_
	);
	LUT4 #(
		.INIT('h8000)
	) name2274 (
		\u12_dout_reg[25]/P0001 ,
		\u12_o9_we_reg/P0001 ,
		\u8_wp_reg[0]/P0001 ,
		\u8_wp_reg[1]/NET0131 ,
		_w4421_
	);
	LUT2 #(
		.INIT('he)
	) name2275 (
		_w4420_,
		_w4421_,
		_w4422_
	);
	LUT4 #(
		.INIT('hc4cc)
	) name2276 (
		\u12_o3_we_reg/P0001 ,
		\u3_mem_reg[2][0]/NET0131 ,
		\u3_wp_reg[0]/P0001 ,
		\u3_wp_reg[1]/NET0131 ,
		_w4423_
	);
	LUT4 #(
		.INIT('h0800)
	) name2277 (
		\u12_dout_reg[0]/P0001 ,
		\u12_o3_we_reg/P0001 ,
		\u3_wp_reg[0]/P0001 ,
		\u3_wp_reg[1]/NET0131 ,
		_w4424_
	);
	LUT2 #(
		.INIT('he)
	) name2278 (
		_w4423_,
		_w4424_,
		_w4425_
	);
	LUT4 #(
		.INIT('h4ccc)
	) name2279 (
		\u12_o9_we_reg/P0001 ,
		\u8_mem_reg[3][27]/NET0131 ,
		\u8_wp_reg[0]/P0001 ,
		\u8_wp_reg[1]/NET0131 ,
		_w4426_
	);
	LUT4 #(
		.INIT('h8000)
	) name2280 (
		\u12_dout_reg[27]/P0001 ,
		\u12_o9_we_reg/P0001 ,
		\u8_wp_reg[0]/P0001 ,
		\u8_wp_reg[1]/NET0131 ,
		_w4427_
	);
	LUT2 #(
		.INIT('he)
	) name2281 (
		_w4426_,
		_w4427_,
		_w4428_
	);
	LUT4 #(
		.INIT('hc4cc)
	) name2282 (
		\u12_o3_we_reg/P0001 ,
		\u3_mem_reg[2][10]/NET0131 ,
		\u3_wp_reg[0]/P0001 ,
		\u3_wp_reg[1]/NET0131 ,
		_w4429_
	);
	LUT4 #(
		.INIT('h0800)
	) name2283 (
		\u12_dout_reg[10]/P0001 ,
		\u12_o3_we_reg/P0001 ,
		\u3_wp_reg[0]/P0001 ,
		\u3_wp_reg[1]/NET0131 ,
		_w4430_
	);
	LUT2 #(
		.INIT('he)
	) name2284 (
		_w4429_,
		_w4430_,
		_w4431_
	);
	LUT4 #(
		.INIT('h4ccc)
	) name2285 (
		\u12_o9_we_reg/P0001 ,
		\u8_mem_reg[3][29]/NET0131 ,
		\u8_wp_reg[0]/P0001 ,
		\u8_wp_reg[1]/NET0131 ,
		_w4432_
	);
	LUT4 #(
		.INIT('h8000)
	) name2286 (
		\u12_dout_reg[29]/P0001 ,
		\u12_o9_we_reg/P0001 ,
		\u8_wp_reg[0]/P0001 ,
		\u8_wp_reg[1]/NET0131 ,
		_w4433_
	);
	LUT2 #(
		.INIT('he)
	) name2287 (
		_w4432_,
		_w4433_,
		_w4434_
	);
	LUT4 #(
		.INIT('hc4cc)
	) name2288 (
		\u12_o3_we_reg/P0001 ,
		\u3_mem_reg[2][11]/NET0131 ,
		\u3_wp_reg[0]/P0001 ,
		\u3_wp_reg[1]/NET0131 ,
		_w4435_
	);
	LUT4 #(
		.INIT('h0800)
	) name2289 (
		\u12_dout_reg[11]/P0001 ,
		\u12_o3_we_reg/P0001 ,
		\u3_wp_reg[0]/P0001 ,
		\u3_wp_reg[1]/NET0131 ,
		_w4436_
	);
	LUT2 #(
		.INIT('he)
	) name2290 (
		_w4435_,
		_w4436_,
		_w4437_
	);
	LUT4 #(
		.INIT('h4ccc)
	) name2291 (
		\u12_o9_we_reg/P0001 ,
		\u8_mem_reg[3][2]/NET0131 ,
		\u8_wp_reg[0]/P0001 ,
		\u8_wp_reg[1]/NET0131 ,
		_w4438_
	);
	LUT4 #(
		.INIT('h8000)
	) name2292 (
		\u12_dout_reg[2]/P0001 ,
		\u12_o9_we_reg/P0001 ,
		\u8_wp_reg[0]/P0001 ,
		\u8_wp_reg[1]/NET0131 ,
		_w4439_
	);
	LUT2 #(
		.INIT('he)
	) name2293 (
		_w4438_,
		_w4439_,
		_w4440_
	);
	LUT4 #(
		.INIT('h4ccc)
	) name2294 (
		\u12_o9_we_reg/P0001 ,
		\u8_mem_reg[3][30]/NET0131 ,
		\u8_wp_reg[0]/P0001 ,
		\u8_wp_reg[1]/NET0131 ,
		_w4441_
	);
	LUT4 #(
		.INIT('h8000)
	) name2295 (
		\u12_dout_reg[30]/P0001 ,
		\u12_o9_we_reg/P0001 ,
		\u8_wp_reg[0]/P0001 ,
		\u8_wp_reg[1]/NET0131 ,
		_w4442_
	);
	LUT2 #(
		.INIT('he)
	) name2296 (
		_w4441_,
		_w4442_,
		_w4443_
	);
	LUT4 #(
		.INIT('hc4cc)
	) name2297 (
		\u12_o3_we_reg/P0001 ,
		\u3_mem_reg[2][12]/NET0131 ,
		\u3_wp_reg[0]/P0001 ,
		\u3_wp_reg[1]/NET0131 ,
		_w4444_
	);
	LUT4 #(
		.INIT('h0800)
	) name2298 (
		\u12_dout_reg[12]/P0001 ,
		\u12_o3_we_reg/P0001 ,
		\u3_wp_reg[0]/P0001 ,
		\u3_wp_reg[1]/NET0131 ,
		_w4445_
	);
	LUT2 #(
		.INIT('he)
	) name2299 (
		_w4444_,
		_w4445_,
		_w4446_
	);
	LUT4 #(
		.INIT('h4ccc)
	) name2300 (
		\u12_o9_we_reg/P0001 ,
		\u8_mem_reg[3][3]/NET0131 ,
		\u8_wp_reg[0]/P0001 ,
		\u8_wp_reg[1]/NET0131 ,
		_w4447_
	);
	LUT4 #(
		.INIT('h8000)
	) name2301 (
		\u12_dout_reg[3]/P0001 ,
		\u12_o9_we_reg/P0001 ,
		\u8_wp_reg[0]/P0001 ,
		\u8_wp_reg[1]/NET0131 ,
		_w4448_
	);
	LUT2 #(
		.INIT('he)
	) name2302 (
		_w4447_,
		_w4448_,
		_w4449_
	);
	LUT4 #(
		.INIT('hc4cc)
	) name2303 (
		\u12_o3_we_reg/P0001 ,
		\u3_mem_reg[2][13]/NET0131 ,
		\u3_wp_reg[0]/P0001 ,
		\u3_wp_reg[1]/NET0131 ,
		_w4450_
	);
	LUT4 #(
		.INIT('h0800)
	) name2304 (
		\u12_dout_reg[13]/P0001 ,
		\u12_o3_we_reg/P0001 ,
		\u3_wp_reg[0]/P0001 ,
		\u3_wp_reg[1]/NET0131 ,
		_w4451_
	);
	LUT2 #(
		.INIT('he)
	) name2305 (
		_w4450_,
		_w4451_,
		_w4452_
	);
	LUT4 #(
		.INIT('h4ccc)
	) name2306 (
		\u12_o9_we_reg/P0001 ,
		\u8_mem_reg[3][5]/NET0131 ,
		\u8_wp_reg[0]/P0001 ,
		\u8_wp_reg[1]/NET0131 ,
		_w4453_
	);
	LUT4 #(
		.INIT('h8000)
	) name2307 (
		\u12_dout_reg[5]/P0001 ,
		\u12_o9_we_reg/P0001 ,
		\u8_wp_reg[0]/P0001 ,
		\u8_wp_reg[1]/NET0131 ,
		_w4454_
	);
	LUT2 #(
		.INIT('he)
	) name2308 (
		_w4453_,
		_w4454_,
		_w4455_
	);
	LUT4 #(
		.INIT('h4ccc)
	) name2309 (
		\u12_o9_we_reg/P0001 ,
		\u8_mem_reg[3][7]/NET0131 ,
		\u8_wp_reg[0]/P0001 ,
		\u8_wp_reg[1]/NET0131 ,
		_w4456_
	);
	LUT4 #(
		.INIT('h8000)
	) name2310 (
		\u12_dout_reg[7]/P0001 ,
		\u12_o9_we_reg/P0001 ,
		\u8_wp_reg[0]/P0001 ,
		\u8_wp_reg[1]/NET0131 ,
		_w4457_
	);
	LUT2 #(
		.INIT('he)
	) name2311 (
		_w4456_,
		_w4457_,
		_w4458_
	);
	LUT4 #(
		.INIT('hc4cc)
	) name2312 (
		\u12_o3_we_reg/P0001 ,
		\u3_mem_reg[2][15]/NET0131 ,
		\u3_wp_reg[0]/P0001 ,
		\u3_wp_reg[1]/NET0131 ,
		_w4459_
	);
	LUT4 #(
		.INIT('h0800)
	) name2313 (
		\u12_dout_reg[15]/P0001 ,
		\u12_o3_we_reg/P0001 ,
		\u3_wp_reg[0]/P0001 ,
		\u3_wp_reg[1]/NET0131 ,
		_w4460_
	);
	LUT2 #(
		.INIT('he)
	) name2314 (
		_w4459_,
		_w4460_,
		_w4461_
	);
	LUT4 #(
		.INIT('h4ccc)
	) name2315 (
		\u12_o9_we_reg/P0001 ,
		\u8_mem_reg[3][9]/NET0131 ,
		\u8_wp_reg[0]/P0001 ,
		\u8_wp_reg[1]/NET0131 ,
		_w4462_
	);
	LUT4 #(
		.INIT('h8000)
	) name2316 (
		\u12_dout_reg[9]/P0001 ,
		\u12_o9_we_reg/P0001 ,
		\u8_wp_reg[0]/P0001 ,
		\u8_wp_reg[1]/NET0131 ,
		_w4463_
	);
	LUT2 #(
		.INIT('he)
	) name2317 (
		_w4462_,
		_w4463_,
		_w4464_
	);
	LUT4 #(
		.INIT('hc4cc)
	) name2318 (
		\u12_o3_we_reg/P0001 ,
		\u3_mem_reg[2][16]/NET0131 ,
		\u3_wp_reg[0]/P0001 ,
		\u3_wp_reg[1]/NET0131 ,
		_w4465_
	);
	LUT4 #(
		.INIT('h0800)
	) name2319 (
		\u12_dout_reg[16]/P0001 ,
		\u12_o3_we_reg/P0001 ,
		\u3_wp_reg[0]/P0001 ,
		\u3_wp_reg[1]/NET0131 ,
		_w4466_
	);
	LUT2 #(
		.INIT('he)
	) name2320 (
		_w4465_,
		_w4466_,
		_w4467_
	);
	LUT4 #(
		.INIT('hcc4c)
	) name2321 (
		\u12_o9_we_reg/P0001 ,
		\u8_mem_reg[1][4]/NET0131 ,
		\u8_wp_reg[0]/P0001 ,
		\u8_wp_reg[1]/NET0131 ,
		_w4468_
	);
	LUT4 #(
		.INIT('h0080)
	) name2322 (
		\u12_dout_reg[4]/P0001 ,
		\u12_o9_we_reg/P0001 ,
		\u8_wp_reg[0]/P0001 ,
		\u8_wp_reg[1]/NET0131 ,
		_w4469_
	);
	LUT2 #(
		.INIT('he)
	) name2323 (
		_w4468_,
		_w4469_,
		_w4470_
	);
	LUT4 #(
		.INIT('hc4cc)
	) name2324 (
		\u12_o3_we_reg/P0001 ,
		\u3_mem_reg[2][18]/NET0131 ,
		\u3_wp_reg[0]/P0001 ,
		\u3_wp_reg[1]/NET0131 ,
		_w4471_
	);
	LUT4 #(
		.INIT('h0800)
	) name2325 (
		\u12_dout_reg[18]/P0001 ,
		\u12_o3_we_reg/P0001 ,
		\u3_wp_reg[0]/P0001 ,
		\u3_wp_reg[1]/NET0131 ,
		_w4472_
	);
	LUT2 #(
		.INIT('he)
	) name2326 (
		_w4471_,
		_w4472_,
		_w4473_
	);
	LUT4 #(
		.INIT('hc4cc)
	) name2327 (
		\u12_o3_we_reg/P0001 ,
		\u3_mem_reg[2][19]/NET0131 ,
		\u3_wp_reg[0]/P0001 ,
		\u3_wp_reg[1]/NET0131 ,
		_w4474_
	);
	LUT4 #(
		.INIT('h0800)
	) name2328 (
		\u12_dout_reg[19]/P0001 ,
		\u12_o3_we_reg/P0001 ,
		\u3_wp_reg[0]/P0001 ,
		\u3_wp_reg[1]/NET0131 ,
		_w4475_
	);
	LUT2 #(
		.INIT('he)
	) name2329 (
		_w4474_,
		_w4475_,
		_w4476_
	);
	LUT4 #(
		.INIT('hc4cc)
	) name2330 (
		\u12_o3_we_reg/P0001 ,
		\u3_mem_reg[2][1]/NET0131 ,
		\u3_wp_reg[0]/P0001 ,
		\u3_wp_reg[1]/NET0131 ,
		_w4477_
	);
	LUT4 #(
		.INIT('h0800)
	) name2331 (
		\u12_dout_reg[1]/P0001 ,
		\u12_o3_we_reg/P0001 ,
		\u3_wp_reg[0]/P0001 ,
		\u3_wp_reg[1]/NET0131 ,
		_w4478_
	);
	LUT2 #(
		.INIT('he)
	) name2332 (
		_w4477_,
		_w4478_,
		_w4479_
	);
	LUT4 #(
		.INIT('hcc4c)
	) name2333 (
		\u12_o3_we_reg/P0001 ,
		\u3_mem_reg[1][30]/NET0131 ,
		\u3_wp_reg[0]/P0001 ,
		\u3_wp_reg[1]/NET0131 ,
		_w4480_
	);
	LUT4 #(
		.INIT('h0080)
	) name2334 (
		\u12_dout_reg[30]/P0001 ,
		\u12_o3_we_reg/P0001 ,
		\u3_wp_reg[0]/P0001 ,
		\u3_wp_reg[1]/NET0131 ,
		_w4481_
	);
	LUT2 #(
		.INIT('he)
	) name2335 (
		_w4480_,
		_w4481_,
		_w4482_
	);
	LUT4 #(
		.INIT('hc4cc)
	) name2336 (
		\u12_o3_we_reg/P0001 ,
		\u3_mem_reg[2][21]/NET0131 ,
		\u3_wp_reg[0]/P0001 ,
		\u3_wp_reg[1]/NET0131 ,
		_w4483_
	);
	LUT4 #(
		.INIT('h0800)
	) name2337 (
		\u12_dout_reg[21]/P0001 ,
		\u12_o3_we_reg/P0001 ,
		\u3_wp_reg[0]/P0001 ,
		\u3_wp_reg[1]/NET0131 ,
		_w4484_
	);
	LUT2 #(
		.INIT('he)
	) name2338 (
		_w4483_,
		_w4484_,
		_w4485_
	);
	LUT4 #(
		.INIT('hc4cc)
	) name2339 (
		\u12_o3_we_reg/P0001 ,
		\u3_mem_reg[2][22]/NET0131 ,
		\u3_wp_reg[0]/P0001 ,
		\u3_wp_reg[1]/NET0131 ,
		_w4486_
	);
	LUT4 #(
		.INIT('h0800)
	) name2340 (
		\u12_dout_reg[22]/P0001 ,
		\u12_o3_we_reg/P0001 ,
		\u3_wp_reg[0]/P0001 ,
		\u3_wp_reg[1]/NET0131 ,
		_w4487_
	);
	LUT2 #(
		.INIT('he)
	) name2341 (
		_w4486_,
		_w4487_,
		_w4488_
	);
	LUT4 #(
		.INIT('hc4cc)
	) name2342 (
		\u12_o3_we_reg/P0001 ,
		\u3_mem_reg[2][24]/NET0131 ,
		\u3_wp_reg[0]/P0001 ,
		\u3_wp_reg[1]/NET0131 ,
		_w4489_
	);
	LUT4 #(
		.INIT('h0800)
	) name2343 (
		\u12_dout_reg[24]/P0001 ,
		\u12_o3_we_reg/P0001 ,
		\u3_wp_reg[0]/P0001 ,
		\u3_wp_reg[1]/NET0131 ,
		_w4490_
	);
	LUT2 #(
		.INIT('he)
	) name2344 (
		_w4489_,
		_w4490_,
		_w4491_
	);
	LUT4 #(
		.INIT('hc4cc)
	) name2345 (
		\u12_o3_we_reg/P0001 ,
		\u3_mem_reg[2][26]/NET0131 ,
		\u3_wp_reg[0]/P0001 ,
		\u3_wp_reg[1]/NET0131 ,
		_w4492_
	);
	LUT4 #(
		.INIT('h0800)
	) name2346 (
		\u12_dout_reg[26]/P0001 ,
		\u12_o3_we_reg/P0001 ,
		\u3_wp_reg[0]/P0001 ,
		\u3_wp_reg[1]/NET0131 ,
		_w4493_
	);
	LUT2 #(
		.INIT('he)
	) name2347 (
		_w4492_,
		_w4493_,
		_w4494_
	);
	LUT4 #(
		.INIT('hc4cc)
	) name2348 (
		\u12_o3_we_reg/P0001 ,
		\u3_mem_reg[2][27]/NET0131 ,
		\u3_wp_reg[0]/P0001 ,
		\u3_wp_reg[1]/NET0131 ,
		_w4495_
	);
	LUT4 #(
		.INIT('h0800)
	) name2349 (
		\u12_dout_reg[27]/P0001 ,
		\u12_o3_we_reg/P0001 ,
		\u3_wp_reg[0]/P0001 ,
		\u3_wp_reg[1]/NET0131 ,
		_w4496_
	);
	LUT2 #(
		.INIT('he)
	) name2350 (
		_w4495_,
		_w4496_,
		_w4497_
	);
	LUT4 #(
		.INIT('hc4cc)
	) name2351 (
		\u12_o3_we_reg/P0001 ,
		\u3_mem_reg[2][28]/NET0131 ,
		\u3_wp_reg[0]/P0001 ,
		\u3_wp_reg[1]/NET0131 ,
		_w4498_
	);
	LUT4 #(
		.INIT('h0800)
	) name2352 (
		\u12_dout_reg[28]/P0001 ,
		\u12_o3_we_reg/P0001 ,
		\u3_wp_reg[0]/P0001 ,
		\u3_wp_reg[1]/NET0131 ,
		_w4499_
	);
	LUT2 #(
		.INIT('he)
	) name2353 (
		_w4498_,
		_w4499_,
		_w4500_
	);
	LUT4 #(
		.INIT('hc4cc)
	) name2354 (
		\u12_o3_we_reg/P0001 ,
		\u3_mem_reg[2][29]/NET0131 ,
		\u3_wp_reg[0]/P0001 ,
		\u3_wp_reg[1]/NET0131 ,
		_w4501_
	);
	LUT4 #(
		.INIT('h0800)
	) name2355 (
		\u12_dout_reg[29]/P0001 ,
		\u12_o3_we_reg/P0001 ,
		\u3_wp_reg[0]/P0001 ,
		\u3_wp_reg[1]/NET0131 ,
		_w4502_
	);
	LUT2 #(
		.INIT('he)
	) name2356 (
		_w4501_,
		_w4502_,
		_w4503_
	);
	LUT4 #(
		.INIT('hc4cc)
	) name2357 (
		\u12_o3_we_reg/P0001 ,
		\u3_mem_reg[2][2]/NET0131 ,
		\u3_wp_reg[0]/P0001 ,
		\u3_wp_reg[1]/NET0131 ,
		_w4504_
	);
	LUT4 #(
		.INIT('h0800)
	) name2358 (
		\u12_dout_reg[2]/P0001 ,
		\u12_o3_we_reg/P0001 ,
		\u3_wp_reg[0]/P0001 ,
		\u3_wp_reg[1]/NET0131 ,
		_w4505_
	);
	LUT2 #(
		.INIT('he)
	) name2359 (
		_w4504_,
		_w4505_,
		_w4506_
	);
	LUT4 #(
		.INIT('hc4cc)
	) name2360 (
		\u12_o3_we_reg/P0001 ,
		\u3_mem_reg[2][30]/NET0131 ,
		\u3_wp_reg[0]/P0001 ,
		\u3_wp_reg[1]/NET0131 ,
		_w4507_
	);
	LUT4 #(
		.INIT('h0800)
	) name2361 (
		\u12_dout_reg[30]/P0001 ,
		\u12_o3_we_reg/P0001 ,
		\u3_wp_reg[0]/P0001 ,
		\u3_wp_reg[1]/NET0131 ,
		_w4508_
	);
	LUT2 #(
		.INIT('he)
	) name2362 (
		_w4507_,
		_w4508_,
		_w4509_
	);
	LUT4 #(
		.INIT('hc4cc)
	) name2363 (
		\u12_o3_we_reg/P0001 ,
		\u3_mem_reg[2][31]/NET0131 ,
		\u3_wp_reg[0]/P0001 ,
		\u3_wp_reg[1]/NET0131 ,
		_w4510_
	);
	LUT4 #(
		.INIT('h0800)
	) name2364 (
		\u12_dout_reg[31]/P0001 ,
		\u12_o3_we_reg/P0001 ,
		\u3_wp_reg[0]/P0001 ,
		\u3_wp_reg[1]/NET0131 ,
		_w4511_
	);
	LUT2 #(
		.INIT('he)
	) name2365 (
		_w4510_,
		_w4511_,
		_w4512_
	);
	LUT4 #(
		.INIT('hc4cc)
	) name2366 (
		\u12_o3_we_reg/P0001 ,
		\u3_mem_reg[2][3]/NET0131 ,
		\u3_wp_reg[0]/P0001 ,
		\u3_wp_reg[1]/NET0131 ,
		_w4513_
	);
	LUT4 #(
		.INIT('h0800)
	) name2367 (
		\u12_dout_reg[3]/P0001 ,
		\u12_o3_we_reg/P0001 ,
		\u3_wp_reg[0]/P0001 ,
		\u3_wp_reg[1]/NET0131 ,
		_w4514_
	);
	LUT2 #(
		.INIT('he)
	) name2368 (
		_w4513_,
		_w4514_,
		_w4515_
	);
	LUT4 #(
		.INIT('hc4cc)
	) name2369 (
		\u12_o3_we_reg/P0001 ,
		\u3_mem_reg[2][4]/NET0131 ,
		\u3_wp_reg[0]/P0001 ,
		\u3_wp_reg[1]/NET0131 ,
		_w4516_
	);
	LUT4 #(
		.INIT('h0800)
	) name2370 (
		\u12_dout_reg[4]/P0001 ,
		\u12_o3_we_reg/P0001 ,
		\u3_wp_reg[0]/P0001 ,
		\u3_wp_reg[1]/NET0131 ,
		_w4517_
	);
	LUT2 #(
		.INIT('he)
	) name2371 (
		_w4516_,
		_w4517_,
		_w4518_
	);
	LUT4 #(
		.INIT('hc4cc)
	) name2372 (
		\u12_o3_we_reg/P0001 ,
		\u3_mem_reg[2][5]/NET0131 ,
		\u3_wp_reg[0]/P0001 ,
		\u3_wp_reg[1]/NET0131 ,
		_w4519_
	);
	LUT4 #(
		.INIT('h0800)
	) name2373 (
		\u12_dout_reg[5]/P0001 ,
		\u12_o3_we_reg/P0001 ,
		\u3_wp_reg[0]/P0001 ,
		\u3_wp_reg[1]/NET0131 ,
		_w4520_
	);
	LUT2 #(
		.INIT('he)
	) name2374 (
		_w4519_,
		_w4520_,
		_w4521_
	);
	LUT4 #(
		.INIT('hc4cc)
	) name2375 (
		\u12_o3_we_reg/P0001 ,
		\u3_mem_reg[2][6]/NET0131 ,
		\u3_wp_reg[0]/P0001 ,
		\u3_wp_reg[1]/NET0131 ,
		_w4522_
	);
	LUT4 #(
		.INIT('h0800)
	) name2376 (
		\u12_dout_reg[6]/P0001 ,
		\u12_o3_we_reg/P0001 ,
		\u3_wp_reg[0]/P0001 ,
		\u3_wp_reg[1]/NET0131 ,
		_w4523_
	);
	LUT2 #(
		.INIT('he)
	) name2377 (
		_w4522_,
		_w4523_,
		_w4524_
	);
	LUT4 #(
		.INIT('hc4cc)
	) name2378 (
		\u12_o3_we_reg/P0001 ,
		\u3_mem_reg[2][7]/NET0131 ,
		\u3_wp_reg[0]/P0001 ,
		\u3_wp_reg[1]/NET0131 ,
		_w4525_
	);
	LUT4 #(
		.INIT('h0800)
	) name2379 (
		\u12_dout_reg[7]/P0001 ,
		\u12_o3_we_reg/P0001 ,
		\u3_wp_reg[0]/P0001 ,
		\u3_wp_reg[1]/NET0131 ,
		_w4526_
	);
	LUT2 #(
		.INIT('he)
	) name2380 (
		_w4525_,
		_w4526_,
		_w4527_
	);
	LUT4 #(
		.INIT('hc4cc)
	) name2381 (
		\u12_o3_we_reg/P0001 ,
		\u3_mem_reg[2][8]/NET0131 ,
		\u3_wp_reg[0]/P0001 ,
		\u3_wp_reg[1]/NET0131 ,
		_w4528_
	);
	LUT4 #(
		.INIT('h0800)
	) name2382 (
		\u12_dout_reg[8]/P0001 ,
		\u12_o3_we_reg/P0001 ,
		\u3_wp_reg[0]/P0001 ,
		\u3_wp_reg[1]/NET0131 ,
		_w4529_
	);
	LUT2 #(
		.INIT('he)
	) name2383 (
		_w4528_,
		_w4529_,
		_w4530_
	);
	LUT4 #(
		.INIT('hc4cc)
	) name2384 (
		\u12_o3_we_reg/P0001 ,
		\u3_mem_reg[2][9]/NET0131 ,
		\u3_wp_reg[0]/P0001 ,
		\u3_wp_reg[1]/NET0131 ,
		_w4531_
	);
	LUT4 #(
		.INIT('h0800)
	) name2385 (
		\u12_dout_reg[9]/P0001 ,
		\u12_o3_we_reg/P0001 ,
		\u3_wp_reg[0]/P0001 ,
		\u3_wp_reg[1]/NET0131 ,
		_w4532_
	);
	LUT2 #(
		.INIT('he)
	) name2386 (
		_w4531_,
		_w4532_,
		_w4533_
	);
	LUT4 #(
		.INIT('h4ccc)
	) name2387 (
		\u12_o3_we_reg/P0001 ,
		\u3_mem_reg[3][0]/NET0131 ,
		\u3_wp_reg[0]/P0001 ,
		\u3_wp_reg[1]/NET0131 ,
		_w4534_
	);
	LUT4 #(
		.INIT('h8000)
	) name2388 (
		\u12_dout_reg[0]/P0001 ,
		\u12_o3_we_reg/P0001 ,
		\u3_wp_reg[0]/P0001 ,
		\u3_wp_reg[1]/NET0131 ,
		_w4535_
	);
	LUT2 #(
		.INIT('he)
	) name2389 (
		_w4534_,
		_w4535_,
		_w4536_
	);
	LUT4 #(
		.INIT('h4ccc)
	) name2390 (
		\u12_o3_we_reg/P0001 ,
		\u3_mem_reg[3][10]/NET0131 ,
		\u3_wp_reg[0]/P0001 ,
		\u3_wp_reg[1]/NET0131 ,
		_w4537_
	);
	LUT4 #(
		.INIT('h8000)
	) name2391 (
		\u12_dout_reg[10]/P0001 ,
		\u12_o3_we_reg/P0001 ,
		\u3_wp_reg[0]/P0001 ,
		\u3_wp_reg[1]/NET0131 ,
		_w4538_
	);
	LUT2 #(
		.INIT('he)
	) name2392 (
		_w4537_,
		_w4538_,
		_w4539_
	);
	LUT4 #(
		.INIT('h4ccc)
	) name2393 (
		\u12_o3_we_reg/P0001 ,
		\u3_mem_reg[3][11]/NET0131 ,
		\u3_wp_reg[0]/P0001 ,
		\u3_wp_reg[1]/NET0131 ,
		_w4540_
	);
	LUT4 #(
		.INIT('h8000)
	) name2394 (
		\u12_dout_reg[11]/P0001 ,
		\u12_o3_we_reg/P0001 ,
		\u3_wp_reg[0]/P0001 ,
		\u3_wp_reg[1]/NET0131 ,
		_w4541_
	);
	LUT2 #(
		.INIT('he)
	) name2395 (
		_w4540_,
		_w4541_,
		_w4542_
	);
	LUT4 #(
		.INIT('h4ccc)
	) name2396 (
		\u12_o3_we_reg/P0001 ,
		\u3_mem_reg[3][12]/NET0131 ,
		\u3_wp_reg[0]/P0001 ,
		\u3_wp_reg[1]/NET0131 ,
		_w4543_
	);
	LUT4 #(
		.INIT('h8000)
	) name2397 (
		\u12_dout_reg[12]/P0001 ,
		\u12_o3_we_reg/P0001 ,
		\u3_wp_reg[0]/P0001 ,
		\u3_wp_reg[1]/NET0131 ,
		_w4544_
	);
	LUT2 #(
		.INIT('he)
	) name2398 (
		_w4543_,
		_w4544_,
		_w4545_
	);
	LUT4 #(
		.INIT('h4ccc)
	) name2399 (
		\u12_o3_we_reg/P0001 ,
		\u3_mem_reg[3][13]/NET0131 ,
		\u3_wp_reg[0]/P0001 ,
		\u3_wp_reg[1]/NET0131 ,
		_w4546_
	);
	LUT4 #(
		.INIT('h8000)
	) name2400 (
		\u12_dout_reg[13]/P0001 ,
		\u12_o3_we_reg/P0001 ,
		\u3_wp_reg[0]/P0001 ,
		\u3_wp_reg[1]/NET0131 ,
		_w4547_
	);
	LUT2 #(
		.INIT('he)
	) name2401 (
		_w4546_,
		_w4547_,
		_w4548_
	);
	LUT4 #(
		.INIT('h4ccc)
	) name2402 (
		\u12_o3_we_reg/P0001 ,
		\u3_mem_reg[3][14]/NET0131 ,
		\u3_wp_reg[0]/P0001 ,
		\u3_wp_reg[1]/NET0131 ,
		_w4549_
	);
	LUT4 #(
		.INIT('h8000)
	) name2403 (
		\u12_dout_reg[14]/P0001 ,
		\u12_o3_we_reg/P0001 ,
		\u3_wp_reg[0]/P0001 ,
		\u3_wp_reg[1]/NET0131 ,
		_w4550_
	);
	LUT2 #(
		.INIT('he)
	) name2404 (
		_w4549_,
		_w4550_,
		_w4551_
	);
	LUT4 #(
		.INIT('h4ccc)
	) name2405 (
		\u12_o3_we_reg/P0001 ,
		\u3_mem_reg[3][15]/NET0131 ,
		\u3_wp_reg[0]/P0001 ,
		\u3_wp_reg[1]/NET0131 ,
		_w4552_
	);
	LUT4 #(
		.INIT('h8000)
	) name2406 (
		\u12_dout_reg[15]/P0001 ,
		\u12_o3_we_reg/P0001 ,
		\u3_wp_reg[0]/P0001 ,
		\u3_wp_reg[1]/NET0131 ,
		_w4553_
	);
	LUT2 #(
		.INIT('he)
	) name2407 (
		_w4552_,
		_w4553_,
		_w4554_
	);
	LUT4 #(
		.INIT('h4ccc)
	) name2408 (
		\u12_o3_we_reg/P0001 ,
		\u3_mem_reg[3][16]/NET0131 ,
		\u3_wp_reg[0]/P0001 ,
		\u3_wp_reg[1]/NET0131 ,
		_w4555_
	);
	LUT4 #(
		.INIT('h8000)
	) name2409 (
		\u12_dout_reg[16]/P0001 ,
		\u12_o3_we_reg/P0001 ,
		\u3_wp_reg[0]/P0001 ,
		\u3_wp_reg[1]/NET0131 ,
		_w4556_
	);
	LUT2 #(
		.INIT('he)
	) name2410 (
		_w4555_,
		_w4556_,
		_w4557_
	);
	LUT4 #(
		.INIT('h4ccc)
	) name2411 (
		\u12_o3_we_reg/P0001 ,
		\u3_mem_reg[3][17]/NET0131 ,
		\u3_wp_reg[0]/P0001 ,
		\u3_wp_reg[1]/NET0131 ,
		_w4558_
	);
	LUT4 #(
		.INIT('h8000)
	) name2412 (
		\u12_dout_reg[17]/P0001 ,
		\u12_o3_we_reg/P0001 ,
		\u3_wp_reg[0]/P0001 ,
		\u3_wp_reg[1]/NET0131 ,
		_w4559_
	);
	LUT2 #(
		.INIT('he)
	) name2413 (
		_w4558_,
		_w4559_,
		_w4560_
	);
	LUT4 #(
		.INIT('h4ccc)
	) name2414 (
		\u12_o3_we_reg/P0001 ,
		\u3_mem_reg[3][18]/NET0131 ,
		\u3_wp_reg[0]/P0001 ,
		\u3_wp_reg[1]/NET0131 ,
		_w4561_
	);
	LUT4 #(
		.INIT('h8000)
	) name2415 (
		\u12_dout_reg[18]/P0001 ,
		\u12_o3_we_reg/P0001 ,
		\u3_wp_reg[0]/P0001 ,
		\u3_wp_reg[1]/NET0131 ,
		_w4562_
	);
	LUT2 #(
		.INIT('he)
	) name2416 (
		_w4561_,
		_w4562_,
		_w4563_
	);
	LUT4 #(
		.INIT('h4ccc)
	) name2417 (
		\u12_o3_we_reg/P0001 ,
		\u3_mem_reg[3][19]/NET0131 ,
		\u3_wp_reg[0]/P0001 ,
		\u3_wp_reg[1]/NET0131 ,
		_w4564_
	);
	LUT4 #(
		.INIT('h8000)
	) name2418 (
		\u12_dout_reg[19]/P0001 ,
		\u12_o3_we_reg/P0001 ,
		\u3_wp_reg[0]/P0001 ,
		\u3_wp_reg[1]/NET0131 ,
		_w4565_
	);
	LUT2 #(
		.INIT('he)
	) name2419 (
		_w4564_,
		_w4565_,
		_w4566_
	);
	LUT4 #(
		.INIT('h4ccc)
	) name2420 (
		\u12_o3_we_reg/P0001 ,
		\u3_mem_reg[3][1]/NET0131 ,
		\u3_wp_reg[0]/P0001 ,
		\u3_wp_reg[1]/NET0131 ,
		_w4567_
	);
	LUT4 #(
		.INIT('h8000)
	) name2421 (
		\u12_dout_reg[1]/P0001 ,
		\u12_o3_we_reg/P0001 ,
		\u3_wp_reg[0]/P0001 ,
		\u3_wp_reg[1]/NET0131 ,
		_w4568_
	);
	LUT2 #(
		.INIT('he)
	) name2422 (
		_w4567_,
		_w4568_,
		_w4569_
	);
	LUT4 #(
		.INIT('h4ccc)
	) name2423 (
		\u12_o3_we_reg/P0001 ,
		\u3_mem_reg[3][21]/NET0131 ,
		\u3_wp_reg[0]/P0001 ,
		\u3_wp_reg[1]/NET0131 ,
		_w4570_
	);
	LUT4 #(
		.INIT('h8000)
	) name2424 (
		\u12_dout_reg[21]/P0001 ,
		\u12_o3_we_reg/P0001 ,
		\u3_wp_reg[0]/P0001 ,
		\u3_wp_reg[1]/NET0131 ,
		_w4571_
	);
	LUT2 #(
		.INIT('he)
	) name2425 (
		_w4570_,
		_w4571_,
		_w4572_
	);
	LUT4 #(
		.INIT('h4ccc)
	) name2426 (
		\u12_o3_we_reg/P0001 ,
		\u3_mem_reg[3][22]/NET0131 ,
		\u3_wp_reg[0]/P0001 ,
		\u3_wp_reg[1]/NET0131 ,
		_w4573_
	);
	LUT4 #(
		.INIT('h8000)
	) name2427 (
		\u12_dout_reg[22]/P0001 ,
		\u12_o3_we_reg/P0001 ,
		\u3_wp_reg[0]/P0001 ,
		\u3_wp_reg[1]/NET0131 ,
		_w4574_
	);
	LUT2 #(
		.INIT('he)
	) name2428 (
		_w4573_,
		_w4574_,
		_w4575_
	);
	LUT4 #(
		.INIT('h4ccc)
	) name2429 (
		\u12_o3_we_reg/P0001 ,
		\u3_mem_reg[3][23]/NET0131 ,
		\u3_wp_reg[0]/P0001 ,
		\u3_wp_reg[1]/NET0131 ,
		_w4576_
	);
	LUT4 #(
		.INIT('h8000)
	) name2430 (
		\u12_dout_reg[23]/P0001 ,
		\u12_o3_we_reg/P0001 ,
		\u3_wp_reg[0]/P0001 ,
		\u3_wp_reg[1]/NET0131 ,
		_w4577_
	);
	LUT2 #(
		.INIT('he)
	) name2431 (
		_w4576_,
		_w4577_,
		_w4578_
	);
	LUT4 #(
		.INIT('h4ccc)
	) name2432 (
		\u12_o3_we_reg/P0001 ,
		\u3_mem_reg[3][24]/NET0131 ,
		\u3_wp_reg[0]/P0001 ,
		\u3_wp_reg[1]/NET0131 ,
		_w4579_
	);
	LUT4 #(
		.INIT('h8000)
	) name2433 (
		\u12_dout_reg[24]/P0001 ,
		\u12_o3_we_reg/P0001 ,
		\u3_wp_reg[0]/P0001 ,
		\u3_wp_reg[1]/NET0131 ,
		_w4580_
	);
	LUT2 #(
		.INIT('he)
	) name2434 (
		_w4579_,
		_w4580_,
		_w4581_
	);
	LUT4 #(
		.INIT('h4ccc)
	) name2435 (
		\u12_o3_we_reg/P0001 ,
		\u3_mem_reg[3][26]/NET0131 ,
		\u3_wp_reg[0]/P0001 ,
		\u3_wp_reg[1]/NET0131 ,
		_w4582_
	);
	LUT4 #(
		.INIT('h8000)
	) name2436 (
		\u12_dout_reg[26]/P0001 ,
		\u12_o3_we_reg/P0001 ,
		\u3_wp_reg[0]/P0001 ,
		\u3_wp_reg[1]/NET0131 ,
		_w4583_
	);
	LUT2 #(
		.INIT('he)
	) name2437 (
		_w4582_,
		_w4583_,
		_w4584_
	);
	LUT4 #(
		.INIT('h4ccc)
	) name2438 (
		\u12_o3_we_reg/P0001 ,
		\u3_mem_reg[3][27]/NET0131 ,
		\u3_wp_reg[0]/P0001 ,
		\u3_wp_reg[1]/NET0131 ,
		_w4585_
	);
	LUT4 #(
		.INIT('h8000)
	) name2439 (
		\u12_dout_reg[27]/P0001 ,
		\u12_o3_we_reg/P0001 ,
		\u3_wp_reg[0]/P0001 ,
		\u3_wp_reg[1]/NET0131 ,
		_w4586_
	);
	LUT2 #(
		.INIT('he)
	) name2440 (
		_w4585_,
		_w4586_,
		_w4587_
	);
	LUT4 #(
		.INIT('h4ccc)
	) name2441 (
		\u12_o9_we_reg/P0001 ,
		\u8_mem_reg[3][28]/NET0131 ,
		\u8_wp_reg[0]/P0001 ,
		\u8_wp_reg[1]/NET0131 ,
		_w4588_
	);
	LUT4 #(
		.INIT('h8000)
	) name2442 (
		\u12_dout_reg[28]/P0001 ,
		\u12_o9_we_reg/P0001 ,
		\u8_wp_reg[0]/P0001 ,
		\u8_wp_reg[1]/NET0131 ,
		_w4589_
	);
	LUT2 #(
		.INIT('he)
	) name2443 (
		_w4588_,
		_w4589_,
		_w4590_
	);
	LUT4 #(
		.INIT('h4ccc)
	) name2444 (
		\u12_o3_we_reg/P0001 ,
		\u3_mem_reg[3][28]/NET0131 ,
		\u3_wp_reg[0]/P0001 ,
		\u3_wp_reg[1]/NET0131 ,
		_w4591_
	);
	LUT4 #(
		.INIT('h8000)
	) name2445 (
		\u12_dout_reg[28]/P0001 ,
		\u12_o3_we_reg/P0001 ,
		\u3_wp_reg[0]/P0001 ,
		\u3_wp_reg[1]/NET0131 ,
		_w4592_
	);
	LUT2 #(
		.INIT('he)
	) name2446 (
		_w4591_,
		_w4592_,
		_w4593_
	);
	LUT4 #(
		.INIT('h4ccc)
	) name2447 (
		\u12_o3_we_reg/P0001 ,
		\u3_mem_reg[3][29]/NET0131 ,
		\u3_wp_reg[0]/P0001 ,
		\u3_wp_reg[1]/NET0131 ,
		_w4594_
	);
	LUT4 #(
		.INIT('h8000)
	) name2448 (
		\u12_dout_reg[29]/P0001 ,
		\u12_o3_we_reg/P0001 ,
		\u3_wp_reg[0]/P0001 ,
		\u3_wp_reg[1]/NET0131 ,
		_w4595_
	);
	LUT2 #(
		.INIT('he)
	) name2449 (
		_w4594_,
		_w4595_,
		_w4596_
	);
	LUT4 #(
		.INIT('h4ccc)
	) name2450 (
		\u12_o3_we_reg/P0001 ,
		\u3_mem_reg[3][2]/NET0131 ,
		\u3_wp_reg[0]/P0001 ,
		\u3_wp_reg[1]/NET0131 ,
		_w4597_
	);
	LUT4 #(
		.INIT('h8000)
	) name2451 (
		\u12_dout_reg[2]/P0001 ,
		\u12_o3_we_reg/P0001 ,
		\u3_wp_reg[0]/P0001 ,
		\u3_wp_reg[1]/NET0131 ,
		_w4598_
	);
	LUT2 #(
		.INIT('he)
	) name2452 (
		_w4597_,
		_w4598_,
		_w4599_
	);
	LUT4 #(
		.INIT('h4ccc)
	) name2453 (
		\u12_o3_we_reg/P0001 ,
		\u3_mem_reg[3][30]/NET0131 ,
		\u3_wp_reg[0]/P0001 ,
		\u3_wp_reg[1]/NET0131 ,
		_w4600_
	);
	LUT4 #(
		.INIT('h8000)
	) name2454 (
		\u12_dout_reg[30]/P0001 ,
		\u12_o3_we_reg/P0001 ,
		\u3_wp_reg[0]/P0001 ,
		\u3_wp_reg[1]/NET0131 ,
		_w4601_
	);
	LUT2 #(
		.INIT('he)
	) name2455 (
		_w4600_,
		_w4601_,
		_w4602_
	);
	LUT4 #(
		.INIT('h4ccc)
	) name2456 (
		\u12_o3_we_reg/P0001 ,
		\u3_mem_reg[3][31]/NET0131 ,
		\u3_wp_reg[0]/P0001 ,
		\u3_wp_reg[1]/NET0131 ,
		_w4603_
	);
	LUT4 #(
		.INIT('h8000)
	) name2457 (
		\u12_dout_reg[31]/P0001 ,
		\u12_o3_we_reg/P0001 ,
		\u3_wp_reg[0]/P0001 ,
		\u3_wp_reg[1]/NET0131 ,
		_w4604_
	);
	LUT2 #(
		.INIT('he)
	) name2458 (
		_w4603_,
		_w4604_,
		_w4605_
	);
	LUT4 #(
		.INIT('h4ccc)
	) name2459 (
		\u12_o3_we_reg/P0001 ,
		\u3_mem_reg[3][4]/NET0131 ,
		\u3_wp_reg[0]/P0001 ,
		\u3_wp_reg[1]/NET0131 ,
		_w4606_
	);
	LUT4 #(
		.INIT('h8000)
	) name2460 (
		\u12_dout_reg[4]/P0001 ,
		\u12_o3_we_reg/P0001 ,
		\u3_wp_reg[0]/P0001 ,
		\u3_wp_reg[1]/NET0131 ,
		_w4607_
	);
	LUT2 #(
		.INIT('he)
	) name2461 (
		_w4606_,
		_w4607_,
		_w4608_
	);
	LUT4 #(
		.INIT('h4ccc)
	) name2462 (
		\u12_o3_we_reg/P0001 ,
		\u3_mem_reg[3][5]/NET0131 ,
		\u3_wp_reg[0]/P0001 ,
		\u3_wp_reg[1]/NET0131 ,
		_w4609_
	);
	LUT4 #(
		.INIT('h8000)
	) name2463 (
		\u12_dout_reg[5]/P0001 ,
		\u12_o3_we_reg/P0001 ,
		\u3_wp_reg[0]/P0001 ,
		\u3_wp_reg[1]/NET0131 ,
		_w4610_
	);
	LUT2 #(
		.INIT('he)
	) name2464 (
		_w4609_,
		_w4610_,
		_w4611_
	);
	LUT4 #(
		.INIT('hcc4c)
	) name2465 (
		\u12_o3_we_reg/P0001 ,
		\u3_mem_reg[1][1]/NET0131 ,
		\u3_wp_reg[0]/P0001 ,
		\u3_wp_reg[1]/NET0131 ,
		_w4612_
	);
	LUT4 #(
		.INIT('h0080)
	) name2466 (
		\u12_dout_reg[1]/P0001 ,
		\u12_o3_we_reg/P0001 ,
		\u3_wp_reg[0]/P0001 ,
		\u3_wp_reg[1]/NET0131 ,
		_w4613_
	);
	LUT2 #(
		.INIT('he)
	) name2467 (
		_w4612_,
		_w4613_,
		_w4614_
	);
	LUT4 #(
		.INIT('h4ccc)
	) name2468 (
		\u12_o3_we_reg/P0001 ,
		\u3_mem_reg[3][6]/NET0131 ,
		\u3_wp_reg[0]/P0001 ,
		\u3_wp_reg[1]/NET0131 ,
		_w4615_
	);
	LUT4 #(
		.INIT('h8000)
	) name2469 (
		\u12_dout_reg[6]/P0001 ,
		\u12_o3_we_reg/P0001 ,
		\u3_wp_reg[0]/P0001 ,
		\u3_wp_reg[1]/NET0131 ,
		_w4616_
	);
	LUT2 #(
		.INIT('he)
	) name2470 (
		_w4615_,
		_w4616_,
		_w4617_
	);
	LUT4 #(
		.INIT('h4ccc)
	) name2471 (
		\u12_o3_we_reg/P0001 ,
		\u3_mem_reg[3][7]/NET0131 ,
		\u3_wp_reg[0]/P0001 ,
		\u3_wp_reg[1]/NET0131 ,
		_w4618_
	);
	LUT4 #(
		.INIT('h8000)
	) name2472 (
		\u12_dout_reg[7]/P0001 ,
		\u12_o3_we_reg/P0001 ,
		\u3_wp_reg[0]/P0001 ,
		\u3_wp_reg[1]/NET0131 ,
		_w4619_
	);
	LUT2 #(
		.INIT('he)
	) name2473 (
		_w4618_,
		_w4619_,
		_w4620_
	);
	LUT4 #(
		.INIT('h4ccc)
	) name2474 (
		\u12_o3_we_reg/P0001 ,
		\u3_mem_reg[3][8]/NET0131 ,
		\u3_wp_reg[0]/P0001 ,
		\u3_wp_reg[1]/NET0131 ,
		_w4621_
	);
	LUT4 #(
		.INIT('h8000)
	) name2475 (
		\u12_dout_reg[8]/P0001 ,
		\u12_o3_we_reg/P0001 ,
		\u3_wp_reg[0]/P0001 ,
		\u3_wp_reg[1]/NET0131 ,
		_w4622_
	);
	LUT2 #(
		.INIT('he)
	) name2476 (
		_w4621_,
		_w4622_,
		_w4623_
	);
	LUT4 #(
		.INIT('h4ccc)
	) name2477 (
		\u12_o3_we_reg/P0001 ,
		\u3_mem_reg[3][9]/NET0131 ,
		\u3_wp_reg[0]/P0001 ,
		\u3_wp_reg[1]/NET0131 ,
		_w4624_
	);
	LUT4 #(
		.INIT('h8000)
	) name2478 (
		\u12_dout_reg[9]/P0001 ,
		\u12_o3_we_reg/P0001 ,
		\u3_wp_reg[0]/P0001 ,
		\u3_wp_reg[1]/NET0131 ,
		_w4625_
	);
	LUT2 #(
		.INIT('he)
	) name2479 (
		_w4624_,
		_w4625_,
		_w4626_
	);
	LUT4 #(
		.INIT('hcc4c)
	) name2480 (
		\u12_o9_we_reg/P0001 ,
		\u8_mem_reg[1][31]/NET0131 ,
		\u8_wp_reg[0]/P0001 ,
		\u8_wp_reg[1]/NET0131 ,
		_w4627_
	);
	LUT4 #(
		.INIT('h0080)
	) name2481 (
		\u12_dout_reg[31]/P0001 ,
		\u12_o9_we_reg/P0001 ,
		\u8_wp_reg[0]/P0001 ,
		\u8_wp_reg[1]/NET0131 ,
		_w4628_
	);
	LUT2 #(
		.INIT('he)
	) name2482 (
		_w4627_,
		_w4628_,
		_w4629_
	);
	LUT4 #(
		.INIT('h4ccc)
	) name2483 (
		\u12_o9_we_reg/P0001 ,
		\u8_mem_reg[3][26]/NET0131 ,
		\u8_wp_reg[0]/P0001 ,
		\u8_wp_reg[1]/NET0131 ,
		_w4630_
	);
	LUT4 #(
		.INIT('h8000)
	) name2484 (
		\u12_dout_reg[26]/P0001 ,
		\u12_o9_we_reg/P0001 ,
		\u8_wp_reg[0]/P0001 ,
		\u8_wp_reg[1]/NET0131 ,
		_w4631_
	);
	LUT2 #(
		.INIT('he)
	) name2485 (
		_w4630_,
		_w4631_,
		_w4632_
	);
	LUT4 #(
		.INIT('hc4cc)
	) name2486 (
		\u12_o9_we_reg/P0001 ,
		\u8_mem_reg[2][3]/NET0131 ,
		\u8_wp_reg[0]/P0001 ,
		\u8_wp_reg[1]/NET0131 ,
		_w4633_
	);
	LUT4 #(
		.INIT('h0800)
	) name2487 (
		\u12_dout_reg[3]/P0001 ,
		\u12_o9_we_reg/P0001 ,
		\u8_wp_reg[0]/P0001 ,
		\u8_wp_reg[1]/NET0131 ,
		_w4634_
	);
	LUT2 #(
		.INIT('he)
	) name2488 (
		_w4633_,
		_w4634_,
		_w4635_
	);
	LUT4 #(
		.INIT('h4ccc)
	) name2489 (
		\u12_o3_we_reg/P0001 ,
		\u3_mem_reg[3][25]/NET0131 ,
		\u3_wp_reg[0]/P0001 ,
		\u3_wp_reg[1]/NET0131 ,
		_w4636_
	);
	LUT4 #(
		.INIT('h8000)
	) name2490 (
		\u12_dout_reg[25]/P0001 ,
		\u12_o3_we_reg/P0001 ,
		\u3_wp_reg[0]/P0001 ,
		\u3_wp_reg[1]/NET0131 ,
		_w4637_
	);
	LUT2 #(
		.INIT('he)
	) name2491 (
		_w4636_,
		_w4637_,
		_w4638_
	);
	LUT4 #(
		.INIT('hcc4c)
	) name2492 (
		\u12_o3_we_reg/P0001 ,
		\u3_mem_reg[1][27]/NET0131 ,
		\u3_wp_reg[0]/P0001 ,
		\u3_wp_reg[1]/NET0131 ,
		_w4639_
	);
	LUT4 #(
		.INIT('h0080)
	) name2493 (
		\u12_dout_reg[27]/P0001 ,
		\u12_o3_we_reg/P0001 ,
		\u3_wp_reg[0]/P0001 ,
		\u3_wp_reg[1]/NET0131 ,
		_w4640_
	);
	LUT2 #(
		.INIT('he)
	) name2494 (
		_w4639_,
		_w4640_,
		_w4641_
	);
	LUT4 #(
		.INIT('hc4cc)
	) name2495 (
		\u12_o3_we_reg/P0001 ,
		\u3_mem_reg[2][23]/NET0131 ,
		\u3_wp_reg[0]/P0001 ,
		\u3_wp_reg[1]/NET0131 ,
		_w4642_
	);
	LUT4 #(
		.INIT('h0800)
	) name2496 (
		\u12_dout_reg[23]/P0001 ,
		\u12_o3_we_reg/P0001 ,
		\u3_wp_reg[0]/P0001 ,
		\u3_wp_reg[1]/NET0131 ,
		_w4643_
	);
	LUT2 #(
		.INIT('he)
	) name2497 (
		_w4642_,
		_w4643_,
		_w4644_
	);
	LUT4 #(
		.INIT('hcc4c)
	) name2498 (
		\u12_o4_we_reg/P0001 ,
		\u4_mem_reg[1][0]/NET0131 ,
		\u4_wp_reg[0]/P0001 ,
		\u4_wp_reg[1]/NET0131 ,
		_w4645_
	);
	LUT4 #(
		.INIT('h0080)
	) name2499 (
		\u12_dout_reg[0]/P0001 ,
		\u12_o4_we_reg/P0001 ,
		\u4_wp_reg[0]/P0001 ,
		\u4_wp_reg[1]/NET0131 ,
		_w4646_
	);
	LUT2 #(
		.INIT('he)
	) name2500 (
		_w4645_,
		_w4646_,
		_w4647_
	);
	LUT4 #(
		.INIT('hcc4c)
	) name2501 (
		\u12_o4_we_reg/P0001 ,
		\u4_mem_reg[1][10]/NET0131 ,
		\u4_wp_reg[0]/P0001 ,
		\u4_wp_reg[1]/NET0131 ,
		_w4648_
	);
	LUT4 #(
		.INIT('h0080)
	) name2502 (
		\u12_dout_reg[10]/P0001 ,
		\u12_o4_we_reg/P0001 ,
		\u4_wp_reg[0]/P0001 ,
		\u4_wp_reg[1]/NET0131 ,
		_w4649_
	);
	LUT2 #(
		.INIT('he)
	) name2503 (
		_w4648_,
		_w4649_,
		_w4650_
	);
	LUT4 #(
		.INIT('hcc4c)
	) name2504 (
		\u12_o4_we_reg/P0001 ,
		\u4_mem_reg[1][11]/NET0131 ,
		\u4_wp_reg[0]/P0001 ,
		\u4_wp_reg[1]/NET0131 ,
		_w4651_
	);
	LUT4 #(
		.INIT('h0080)
	) name2505 (
		\u12_dout_reg[11]/P0001 ,
		\u12_o4_we_reg/P0001 ,
		\u4_wp_reg[0]/P0001 ,
		\u4_wp_reg[1]/NET0131 ,
		_w4652_
	);
	LUT2 #(
		.INIT('he)
	) name2506 (
		_w4651_,
		_w4652_,
		_w4653_
	);
	LUT4 #(
		.INIT('hcc4c)
	) name2507 (
		\u12_o4_we_reg/P0001 ,
		\u4_mem_reg[1][12]/NET0131 ,
		\u4_wp_reg[0]/P0001 ,
		\u4_wp_reg[1]/NET0131 ,
		_w4654_
	);
	LUT4 #(
		.INIT('h0080)
	) name2508 (
		\u12_dout_reg[12]/P0001 ,
		\u12_o4_we_reg/P0001 ,
		\u4_wp_reg[0]/P0001 ,
		\u4_wp_reg[1]/NET0131 ,
		_w4655_
	);
	LUT2 #(
		.INIT('he)
	) name2509 (
		_w4654_,
		_w4655_,
		_w4656_
	);
	LUT4 #(
		.INIT('hcc4c)
	) name2510 (
		\u12_o4_we_reg/P0001 ,
		\u4_mem_reg[1][13]/NET0131 ,
		\u4_wp_reg[0]/P0001 ,
		\u4_wp_reg[1]/NET0131 ,
		_w4657_
	);
	LUT4 #(
		.INIT('h0080)
	) name2511 (
		\u12_dout_reg[13]/P0001 ,
		\u12_o4_we_reg/P0001 ,
		\u4_wp_reg[0]/P0001 ,
		\u4_wp_reg[1]/NET0131 ,
		_w4658_
	);
	LUT2 #(
		.INIT('he)
	) name2512 (
		_w4657_,
		_w4658_,
		_w4659_
	);
	LUT4 #(
		.INIT('hcc4c)
	) name2513 (
		\u12_o4_we_reg/P0001 ,
		\u4_mem_reg[1][14]/NET0131 ,
		\u4_wp_reg[0]/P0001 ,
		\u4_wp_reg[1]/NET0131 ,
		_w4660_
	);
	LUT4 #(
		.INIT('h0080)
	) name2514 (
		\u12_dout_reg[14]/P0001 ,
		\u12_o4_we_reg/P0001 ,
		\u4_wp_reg[0]/P0001 ,
		\u4_wp_reg[1]/NET0131 ,
		_w4661_
	);
	LUT2 #(
		.INIT('he)
	) name2515 (
		_w4660_,
		_w4661_,
		_w4662_
	);
	LUT4 #(
		.INIT('hcc4c)
	) name2516 (
		\u12_o4_we_reg/P0001 ,
		\u4_mem_reg[1][15]/NET0131 ,
		\u4_wp_reg[0]/P0001 ,
		\u4_wp_reg[1]/NET0131 ,
		_w4663_
	);
	LUT4 #(
		.INIT('h0080)
	) name2517 (
		\u12_dout_reg[15]/P0001 ,
		\u12_o4_we_reg/P0001 ,
		\u4_wp_reg[0]/P0001 ,
		\u4_wp_reg[1]/NET0131 ,
		_w4664_
	);
	LUT2 #(
		.INIT('he)
	) name2518 (
		_w4663_,
		_w4664_,
		_w4665_
	);
	LUT4 #(
		.INIT('hcc4c)
	) name2519 (
		\u12_o4_we_reg/P0001 ,
		\u4_mem_reg[1][16]/NET0131 ,
		\u4_wp_reg[0]/P0001 ,
		\u4_wp_reg[1]/NET0131 ,
		_w4666_
	);
	LUT4 #(
		.INIT('h0080)
	) name2520 (
		\u12_dout_reg[16]/P0001 ,
		\u12_o4_we_reg/P0001 ,
		\u4_wp_reg[0]/P0001 ,
		\u4_wp_reg[1]/NET0131 ,
		_w4667_
	);
	LUT2 #(
		.INIT('he)
	) name2521 (
		_w4666_,
		_w4667_,
		_w4668_
	);
	LUT4 #(
		.INIT('hcc4c)
	) name2522 (
		\u12_o4_we_reg/P0001 ,
		\u4_mem_reg[1][17]/NET0131 ,
		\u4_wp_reg[0]/P0001 ,
		\u4_wp_reg[1]/NET0131 ,
		_w4669_
	);
	LUT4 #(
		.INIT('h0080)
	) name2523 (
		\u12_dout_reg[17]/P0001 ,
		\u12_o4_we_reg/P0001 ,
		\u4_wp_reg[0]/P0001 ,
		\u4_wp_reg[1]/NET0131 ,
		_w4670_
	);
	LUT2 #(
		.INIT('he)
	) name2524 (
		_w4669_,
		_w4670_,
		_w4671_
	);
	LUT4 #(
		.INIT('hcc4c)
	) name2525 (
		\u12_o4_we_reg/P0001 ,
		\u4_mem_reg[1][18]/NET0131 ,
		\u4_wp_reg[0]/P0001 ,
		\u4_wp_reg[1]/NET0131 ,
		_w4672_
	);
	LUT4 #(
		.INIT('h0080)
	) name2526 (
		\u12_dout_reg[18]/P0001 ,
		\u12_o4_we_reg/P0001 ,
		\u4_wp_reg[0]/P0001 ,
		\u4_wp_reg[1]/NET0131 ,
		_w4673_
	);
	LUT2 #(
		.INIT('he)
	) name2527 (
		_w4672_,
		_w4673_,
		_w4674_
	);
	LUT4 #(
		.INIT('hcc4c)
	) name2528 (
		\u12_o4_we_reg/P0001 ,
		\u4_mem_reg[1][19]/NET0131 ,
		\u4_wp_reg[0]/P0001 ,
		\u4_wp_reg[1]/NET0131 ,
		_w4675_
	);
	LUT4 #(
		.INIT('h0080)
	) name2529 (
		\u12_dout_reg[19]/P0001 ,
		\u12_o4_we_reg/P0001 ,
		\u4_wp_reg[0]/P0001 ,
		\u4_wp_reg[1]/NET0131 ,
		_w4676_
	);
	LUT2 #(
		.INIT('he)
	) name2530 (
		_w4675_,
		_w4676_,
		_w4677_
	);
	LUT4 #(
		.INIT('hcc4c)
	) name2531 (
		\u12_o4_we_reg/P0001 ,
		\u4_mem_reg[1][1]/NET0131 ,
		\u4_wp_reg[0]/P0001 ,
		\u4_wp_reg[1]/NET0131 ,
		_w4678_
	);
	LUT4 #(
		.INIT('h0080)
	) name2532 (
		\u12_dout_reg[1]/P0001 ,
		\u12_o4_we_reg/P0001 ,
		\u4_wp_reg[0]/P0001 ,
		\u4_wp_reg[1]/NET0131 ,
		_w4679_
	);
	LUT2 #(
		.INIT('he)
	) name2533 (
		_w4678_,
		_w4679_,
		_w4680_
	);
	LUT4 #(
		.INIT('hcc4c)
	) name2534 (
		\u12_o4_we_reg/P0001 ,
		\u4_mem_reg[1][20]/NET0131 ,
		\u4_wp_reg[0]/P0001 ,
		\u4_wp_reg[1]/NET0131 ,
		_w4681_
	);
	LUT4 #(
		.INIT('h0080)
	) name2535 (
		\u12_dout_reg[20]/P0001 ,
		\u12_o4_we_reg/P0001 ,
		\u4_wp_reg[0]/P0001 ,
		\u4_wp_reg[1]/NET0131 ,
		_w4682_
	);
	LUT2 #(
		.INIT('he)
	) name2536 (
		_w4681_,
		_w4682_,
		_w4683_
	);
	LUT4 #(
		.INIT('hcc4c)
	) name2537 (
		\u12_o4_we_reg/P0001 ,
		\u4_mem_reg[1][21]/NET0131 ,
		\u4_wp_reg[0]/P0001 ,
		\u4_wp_reg[1]/NET0131 ,
		_w4684_
	);
	LUT4 #(
		.INIT('h0080)
	) name2538 (
		\u12_dout_reg[21]/P0001 ,
		\u12_o4_we_reg/P0001 ,
		\u4_wp_reg[0]/P0001 ,
		\u4_wp_reg[1]/NET0131 ,
		_w4685_
	);
	LUT2 #(
		.INIT('he)
	) name2539 (
		_w4684_,
		_w4685_,
		_w4686_
	);
	LUT4 #(
		.INIT('hcc4c)
	) name2540 (
		\u12_o4_we_reg/P0001 ,
		\u4_mem_reg[1][22]/NET0131 ,
		\u4_wp_reg[0]/P0001 ,
		\u4_wp_reg[1]/NET0131 ,
		_w4687_
	);
	LUT4 #(
		.INIT('h0080)
	) name2541 (
		\u12_dout_reg[22]/P0001 ,
		\u12_o4_we_reg/P0001 ,
		\u4_wp_reg[0]/P0001 ,
		\u4_wp_reg[1]/NET0131 ,
		_w4688_
	);
	LUT2 #(
		.INIT('he)
	) name2542 (
		_w4687_,
		_w4688_,
		_w4689_
	);
	LUT4 #(
		.INIT('hcc4c)
	) name2543 (
		\u12_o4_we_reg/P0001 ,
		\u4_mem_reg[1][23]/NET0131 ,
		\u4_wp_reg[0]/P0001 ,
		\u4_wp_reg[1]/NET0131 ,
		_w4690_
	);
	LUT4 #(
		.INIT('h0080)
	) name2544 (
		\u12_dout_reg[23]/P0001 ,
		\u12_o4_we_reg/P0001 ,
		\u4_wp_reg[0]/P0001 ,
		\u4_wp_reg[1]/NET0131 ,
		_w4691_
	);
	LUT2 #(
		.INIT('he)
	) name2545 (
		_w4690_,
		_w4691_,
		_w4692_
	);
	LUT4 #(
		.INIT('hcc4c)
	) name2546 (
		\u12_o4_we_reg/P0001 ,
		\u4_mem_reg[1][24]/NET0131 ,
		\u4_wp_reg[0]/P0001 ,
		\u4_wp_reg[1]/NET0131 ,
		_w4693_
	);
	LUT4 #(
		.INIT('h0080)
	) name2547 (
		\u12_dout_reg[24]/P0001 ,
		\u12_o4_we_reg/P0001 ,
		\u4_wp_reg[0]/P0001 ,
		\u4_wp_reg[1]/NET0131 ,
		_w4694_
	);
	LUT2 #(
		.INIT('he)
	) name2548 (
		_w4693_,
		_w4694_,
		_w4695_
	);
	LUT4 #(
		.INIT('hcc4c)
	) name2549 (
		\u12_o4_we_reg/P0001 ,
		\u4_mem_reg[1][25]/NET0131 ,
		\u4_wp_reg[0]/P0001 ,
		\u4_wp_reg[1]/NET0131 ,
		_w4696_
	);
	LUT4 #(
		.INIT('h0080)
	) name2550 (
		\u12_dout_reg[25]/P0001 ,
		\u12_o4_we_reg/P0001 ,
		\u4_wp_reg[0]/P0001 ,
		\u4_wp_reg[1]/NET0131 ,
		_w4697_
	);
	LUT2 #(
		.INIT('he)
	) name2551 (
		_w4696_,
		_w4697_,
		_w4698_
	);
	LUT4 #(
		.INIT('hcc4c)
	) name2552 (
		\u12_o4_we_reg/P0001 ,
		\u4_mem_reg[1][26]/NET0131 ,
		\u4_wp_reg[0]/P0001 ,
		\u4_wp_reg[1]/NET0131 ,
		_w4699_
	);
	LUT4 #(
		.INIT('h0080)
	) name2553 (
		\u12_dout_reg[26]/P0001 ,
		\u12_o4_we_reg/P0001 ,
		\u4_wp_reg[0]/P0001 ,
		\u4_wp_reg[1]/NET0131 ,
		_w4700_
	);
	LUT2 #(
		.INIT('he)
	) name2554 (
		_w4699_,
		_w4700_,
		_w4701_
	);
	LUT4 #(
		.INIT('hcc4c)
	) name2555 (
		\u12_o4_we_reg/P0001 ,
		\u4_mem_reg[1][27]/NET0131 ,
		\u4_wp_reg[0]/P0001 ,
		\u4_wp_reg[1]/NET0131 ,
		_w4702_
	);
	LUT4 #(
		.INIT('h0080)
	) name2556 (
		\u12_dout_reg[27]/P0001 ,
		\u12_o4_we_reg/P0001 ,
		\u4_wp_reg[0]/P0001 ,
		\u4_wp_reg[1]/NET0131 ,
		_w4703_
	);
	LUT2 #(
		.INIT('he)
	) name2557 (
		_w4702_,
		_w4703_,
		_w4704_
	);
	LUT4 #(
		.INIT('hcc4c)
	) name2558 (
		\u12_o4_we_reg/P0001 ,
		\u4_mem_reg[1][28]/NET0131 ,
		\u4_wp_reg[0]/P0001 ,
		\u4_wp_reg[1]/NET0131 ,
		_w4705_
	);
	LUT4 #(
		.INIT('h0080)
	) name2559 (
		\u12_dout_reg[28]/P0001 ,
		\u12_o4_we_reg/P0001 ,
		\u4_wp_reg[0]/P0001 ,
		\u4_wp_reg[1]/NET0131 ,
		_w4706_
	);
	LUT2 #(
		.INIT('he)
	) name2560 (
		_w4705_,
		_w4706_,
		_w4707_
	);
	LUT4 #(
		.INIT('hcc4c)
	) name2561 (
		\u12_o4_we_reg/P0001 ,
		\u4_mem_reg[1][29]/NET0131 ,
		\u4_wp_reg[0]/P0001 ,
		\u4_wp_reg[1]/NET0131 ,
		_w4708_
	);
	LUT4 #(
		.INIT('h0080)
	) name2562 (
		\u12_dout_reg[29]/P0001 ,
		\u12_o4_we_reg/P0001 ,
		\u4_wp_reg[0]/P0001 ,
		\u4_wp_reg[1]/NET0131 ,
		_w4709_
	);
	LUT2 #(
		.INIT('he)
	) name2563 (
		_w4708_,
		_w4709_,
		_w4710_
	);
	LUT4 #(
		.INIT('hcc4c)
	) name2564 (
		\u12_o4_we_reg/P0001 ,
		\u4_mem_reg[1][2]/NET0131 ,
		\u4_wp_reg[0]/P0001 ,
		\u4_wp_reg[1]/NET0131 ,
		_w4711_
	);
	LUT4 #(
		.INIT('h0080)
	) name2565 (
		\u12_dout_reg[2]/P0001 ,
		\u12_o4_we_reg/P0001 ,
		\u4_wp_reg[0]/P0001 ,
		\u4_wp_reg[1]/NET0131 ,
		_w4712_
	);
	LUT2 #(
		.INIT('he)
	) name2566 (
		_w4711_,
		_w4712_,
		_w4713_
	);
	LUT4 #(
		.INIT('hcc4c)
	) name2567 (
		\u12_o4_we_reg/P0001 ,
		\u4_mem_reg[1][30]/NET0131 ,
		\u4_wp_reg[0]/P0001 ,
		\u4_wp_reg[1]/NET0131 ,
		_w4714_
	);
	LUT4 #(
		.INIT('h0080)
	) name2568 (
		\u12_dout_reg[30]/P0001 ,
		\u12_o4_we_reg/P0001 ,
		\u4_wp_reg[0]/P0001 ,
		\u4_wp_reg[1]/NET0131 ,
		_w4715_
	);
	LUT2 #(
		.INIT('he)
	) name2569 (
		_w4714_,
		_w4715_,
		_w4716_
	);
	LUT4 #(
		.INIT('hcc4c)
	) name2570 (
		\u12_o4_we_reg/P0001 ,
		\u4_mem_reg[1][31]/NET0131 ,
		\u4_wp_reg[0]/P0001 ,
		\u4_wp_reg[1]/NET0131 ,
		_w4717_
	);
	LUT4 #(
		.INIT('h0080)
	) name2571 (
		\u12_dout_reg[31]/P0001 ,
		\u12_o4_we_reg/P0001 ,
		\u4_wp_reg[0]/P0001 ,
		\u4_wp_reg[1]/NET0131 ,
		_w4718_
	);
	LUT2 #(
		.INIT('he)
	) name2572 (
		_w4717_,
		_w4718_,
		_w4719_
	);
	LUT4 #(
		.INIT('hcc4c)
	) name2573 (
		\u12_o4_we_reg/P0001 ,
		\u4_mem_reg[1][3]/NET0131 ,
		\u4_wp_reg[0]/P0001 ,
		\u4_wp_reg[1]/NET0131 ,
		_w4720_
	);
	LUT4 #(
		.INIT('h0080)
	) name2574 (
		\u12_dout_reg[3]/P0001 ,
		\u12_o4_we_reg/P0001 ,
		\u4_wp_reg[0]/P0001 ,
		\u4_wp_reg[1]/NET0131 ,
		_w4721_
	);
	LUT2 #(
		.INIT('he)
	) name2575 (
		_w4720_,
		_w4721_,
		_w4722_
	);
	LUT4 #(
		.INIT('hcc4c)
	) name2576 (
		\u12_o4_we_reg/P0001 ,
		\u4_mem_reg[1][4]/NET0131 ,
		\u4_wp_reg[0]/P0001 ,
		\u4_wp_reg[1]/NET0131 ,
		_w4723_
	);
	LUT4 #(
		.INIT('h0080)
	) name2577 (
		\u12_dout_reg[4]/P0001 ,
		\u12_o4_we_reg/P0001 ,
		\u4_wp_reg[0]/P0001 ,
		\u4_wp_reg[1]/NET0131 ,
		_w4724_
	);
	LUT2 #(
		.INIT('he)
	) name2578 (
		_w4723_,
		_w4724_,
		_w4725_
	);
	LUT4 #(
		.INIT('hcc4c)
	) name2579 (
		\u12_o4_we_reg/P0001 ,
		\u4_mem_reg[1][5]/NET0131 ,
		\u4_wp_reg[0]/P0001 ,
		\u4_wp_reg[1]/NET0131 ,
		_w4726_
	);
	LUT4 #(
		.INIT('h0080)
	) name2580 (
		\u12_dout_reg[5]/P0001 ,
		\u12_o4_we_reg/P0001 ,
		\u4_wp_reg[0]/P0001 ,
		\u4_wp_reg[1]/NET0131 ,
		_w4727_
	);
	LUT2 #(
		.INIT('he)
	) name2581 (
		_w4726_,
		_w4727_,
		_w4728_
	);
	LUT4 #(
		.INIT('hcc4c)
	) name2582 (
		\u12_o4_we_reg/P0001 ,
		\u4_mem_reg[1][6]/NET0131 ,
		\u4_wp_reg[0]/P0001 ,
		\u4_wp_reg[1]/NET0131 ,
		_w4729_
	);
	LUT4 #(
		.INIT('h0080)
	) name2583 (
		\u12_dout_reg[6]/P0001 ,
		\u12_o4_we_reg/P0001 ,
		\u4_wp_reg[0]/P0001 ,
		\u4_wp_reg[1]/NET0131 ,
		_w4730_
	);
	LUT2 #(
		.INIT('he)
	) name2584 (
		_w4729_,
		_w4730_,
		_w4731_
	);
	LUT4 #(
		.INIT('hcc4c)
	) name2585 (
		\u12_o4_we_reg/P0001 ,
		\u4_mem_reg[1][7]/NET0131 ,
		\u4_wp_reg[0]/P0001 ,
		\u4_wp_reg[1]/NET0131 ,
		_w4732_
	);
	LUT4 #(
		.INIT('h0080)
	) name2586 (
		\u12_dout_reg[7]/P0001 ,
		\u12_o4_we_reg/P0001 ,
		\u4_wp_reg[0]/P0001 ,
		\u4_wp_reg[1]/NET0131 ,
		_w4733_
	);
	LUT2 #(
		.INIT('he)
	) name2587 (
		_w4732_,
		_w4733_,
		_w4734_
	);
	LUT4 #(
		.INIT('hcc4c)
	) name2588 (
		\u12_o4_we_reg/P0001 ,
		\u4_mem_reg[1][8]/NET0131 ,
		\u4_wp_reg[0]/P0001 ,
		\u4_wp_reg[1]/NET0131 ,
		_w4735_
	);
	LUT4 #(
		.INIT('h0080)
	) name2589 (
		\u12_dout_reg[8]/P0001 ,
		\u12_o4_we_reg/P0001 ,
		\u4_wp_reg[0]/P0001 ,
		\u4_wp_reg[1]/NET0131 ,
		_w4736_
	);
	LUT2 #(
		.INIT('he)
	) name2590 (
		_w4735_,
		_w4736_,
		_w4737_
	);
	LUT4 #(
		.INIT('hcc4c)
	) name2591 (
		\u12_o4_we_reg/P0001 ,
		\u4_mem_reg[1][9]/NET0131 ,
		\u4_wp_reg[0]/P0001 ,
		\u4_wp_reg[1]/NET0131 ,
		_w4738_
	);
	LUT4 #(
		.INIT('h0080)
	) name2592 (
		\u12_dout_reg[9]/P0001 ,
		\u12_o4_we_reg/P0001 ,
		\u4_wp_reg[0]/P0001 ,
		\u4_wp_reg[1]/NET0131 ,
		_w4739_
	);
	LUT2 #(
		.INIT('he)
	) name2593 (
		_w4738_,
		_w4739_,
		_w4740_
	);
	LUT4 #(
		.INIT('hc4cc)
	) name2594 (
		\u12_o4_we_reg/P0001 ,
		\u4_mem_reg[2][0]/NET0131 ,
		\u4_wp_reg[0]/P0001 ,
		\u4_wp_reg[1]/NET0131 ,
		_w4741_
	);
	LUT4 #(
		.INIT('h0800)
	) name2595 (
		\u12_dout_reg[0]/P0001 ,
		\u12_o4_we_reg/P0001 ,
		\u4_wp_reg[0]/P0001 ,
		\u4_wp_reg[1]/NET0131 ,
		_w4742_
	);
	LUT2 #(
		.INIT('he)
	) name2596 (
		_w4741_,
		_w4742_,
		_w4743_
	);
	LUT4 #(
		.INIT('hc4cc)
	) name2597 (
		\u12_o4_we_reg/P0001 ,
		\u4_mem_reg[2][10]/NET0131 ,
		\u4_wp_reg[0]/P0001 ,
		\u4_wp_reg[1]/NET0131 ,
		_w4744_
	);
	LUT4 #(
		.INIT('h0800)
	) name2598 (
		\u12_dout_reg[10]/P0001 ,
		\u12_o4_we_reg/P0001 ,
		\u4_wp_reg[0]/P0001 ,
		\u4_wp_reg[1]/NET0131 ,
		_w4745_
	);
	LUT2 #(
		.INIT('he)
	) name2599 (
		_w4744_,
		_w4745_,
		_w4746_
	);
	LUT4 #(
		.INIT('hc4cc)
	) name2600 (
		\u12_o4_we_reg/P0001 ,
		\u4_mem_reg[2][11]/NET0131 ,
		\u4_wp_reg[0]/P0001 ,
		\u4_wp_reg[1]/NET0131 ,
		_w4747_
	);
	LUT4 #(
		.INIT('h0800)
	) name2601 (
		\u12_dout_reg[11]/P0001 ,
		\u12_o4_we_reg/P0001 ,
		\u4_wp_reg[0]/P0001 ,
		\u4_wp_reg[1]/NET0131 ,
		_w4748_
	);
	LUT2 #(
		.INIT('he)
	) name2602 (
		_w4747_,
		_w4748_,
		_w4749_
	);
	LUT4 #(
		.INIT('hc4cc)
	) name2603 (
		\u12_o4_we_reg/P0001 ,
		\u4_mem_reg[2][12]/NET0131 ,
		\u4_wp_reg[0]/P0001 ,
		\u4_wp_reg[1]/NET0131 ,
		_w4750_
	);
	LUT4 #(
		.INIT('h0800)
	) name2604 (
		\u12_dout_reg[12]/P0001 ,
		\u12_o4_we_reg/P0001 ,
		\u4_wp_reg[0]/P0001 ,
		\u4_wp_reg[1]/NET0131 ,
		_w4751_
	);
	LUT2 #(
		.INIT('he)
	) name2605 (
		_w4750_,
		_w4751_,
		_w4752_
	);
	LUT4 #(
		.INIT('hc4cc)
	) name2606 (
		\u12_o4_we_reg/P0001 ,
		\u4_mem_reg[2][13]/NET0131 ,
		\u4_wp_reg[0]/P0001 ,
		\u4_wp_reg[1]/NET0131 ,
		_w4753_
	);
	LUT4 #(
		.INIT('h0800)
	) name2607 (
		\u12_dout_reg[13]/P0001 ,
		\u12_o4_we_reg/P0001 ,
		\u4_wp_reg[0]/P0001 ,
		\u4_wp_reg[1]/NET0131 ,
		_w4754_
	);
	LUT2 #(
		.INIT('he)
	) name2608 (
		_w4753_,
		_w4754_,
		_w4755_
	);
	LUT4 #(
		.INIT('hc4cc)
	) name2609 (
		\u12_o4_we_reg/P0001 ,
		\u4_mem_reg[2][14]/NET0131 ,
		\u4_wp_reg[0]/P0001 ,
		\u4_wp_reg[1]/NET0131 ,
		_w4756_
	);
	LUT4 #(
		.INIT('h0800)
	) name2610 (
		\u12_dout_reg[14]/P0001 ,
		\u12_o4_we_reg/P0001 ,
		\u4_wp_reg[0]/P0001 ,
		\u4_wp_reg[1]/NET0131 ,
		_w4757_
	);
	LUT2 #(
		.INIT('he)
	) name2611 (
		_w4756_,
		_w4757_,
		_w4758_
	);
	LUT4 #(
		.INIT('hc4cc)
	) name2612 (
		\u12_o4_we_reg/P0001 ,
		\u4_mem_reg[2][15]/NET0131 ,
		\u4_wp_reg[0]/P0001 ,
		\u4_wp_reg[1]/NET0131 ,
		_w4759_
	);
	LUT4 #(
		.INIT('h0800)
	) name2613 (
		\u12_dout_reg[15]/P0001 ,
		\u12_o4_we_reg/P0001 ,
		\u4_wp_reg[0]/P0001 ,
		\u4_wp_reg[1]/NET0131 ,
		_w4760_
	);
	LUT2 #(
		.INIT('he)
	) name2614 (
		_w4759_,
		_w4760_,
		_w4761_
	);
	LUT4 #(
		.INIT('hc4cc)
	) name2615 (
		\u12_o4_we_reg/P0001 ,
		\u4_mem_reg[2][16]/NET0131 ,
		\u4_wp_reg[0]/P0001 ,
		\u4_wp_reg[1]/NET0131 ,
		_w4762_
	);
	LUT4 #(
		.INIT('h0800)
	) name2616 (
		\u12_dout_reg[16]/P0001 ,
		\u12_o4_we_reg/P0001 ,
		\u4_wp_reg[0]/P0001 ,
		\u4_wp_reg[1]/NET0131 ,
		_w4763_
	);
	LUT2 #(
		.INIT('he)
	) name2617 (
		_w4762_,
		_w4763_,
		_w4764_
	);
	LUT4 #(
		.INIT('hc4cc)
	) name2618 (
		\u12_o4_we_reg/P0001 ,
		\u4_mem_reg[2][17]/NET0131 ,
		\u4_wp_reg[0]/P0001 ,
		\u4_wp_reg[1]/NET0131 ,
		_w4765_
	);
	LUT4 #(
		.INIT('h0800)
	) name2619 (
		\u12_dout_reg[17]/P0001 ,
		\u12_o4_we_reg/P0001 ,
		\u4_wp_reg[0]/P0001 ,
		\u4_wp_reg[1]/NET0131 ,
		_w4766_
	);
	LUT2 #(
		.INIT('he)
	) name2620 (
		_w4765_,
		_w4766_,
		_w4767_
	);
	LUT4 #(
		.INIT('hc4cc)
	) name2621 (
		\u12_o4_we_reg/P0001 ,
		\u4_mem_reg[2][18]/NET0131 ,
		\u4_wp_reg[0]/P0001 ,
		\u4_wp_reg[1]/NET0131 ,
		_w4768_
	);
	LUT4 #(
		.INIT('h0800)
	) name2622 (
		\u12_dout_reg[18]/P0001 ,
		\u12_o4_we_reg/P0001 ,
		\u4_wp_reg[0]/P0001 ,
		\u4_wp_reg[1]/NET0131 ,
		_w4769_
	);
	LUT2 #(
		.INIT('he)
	) name2623 (
		_w4768_,
		_w4769_,
		_w4770_
	);
	LUT4 #(
		.INIT('hc4cc)
	) name2624 (
		\u12_o4_we_reg/P0001 ,
		\u4_mem_reg[2][19]/NET0131 ,
		\u4_wp_reg[0]/P0001 ,
		\u4_wp_reg[1]/NET0131 ,
		_w4771_
	);
	LUT4 #(
		.INIT('h0800)
	) name2625 (
		\u12_dout_reg[19]/P0001 ,
		\u12_o4_we_reg/P0001 ,
		\u4_wp_reg[0]/P0001 ,
		\u4_wp_reg[1]/NET0131 ,
		_w4772_
	);
	LUT2 #(
		.INIT('he)
	) name2626 (
		_w4771_,
		_w4772_,
		_w4773_
	);
	LUT4 #(
		.INIT('hc4cc)
	) name2627 (
		\u12_o4_we_reg/P0001 ,
		\u4_mem_reg[2][1]/NET0131 ,
		\u4_wp_reg[0]/P0001 ,
		\u4_wp_reg[1]/NET0131 ,
		_w4774_
	);
	LUT4 #(
		.INIT('h0800)
	) name2628 (
		\u12_dout_reg[1]/P0001 ,
		\u12_o4_we_reg/P0001 ,
		\u4_wp_reg[0]/P0001 ,
		\u4_wp_reg[1]/NET0131 ,
		_w4775_
	);
	LUT2 #(
		.INIT('he)
	) name2629 (
		_w4774_,
		_w4775_,
		_w4776_
	);
	LUT4 #(
		.INIT('hc4cc)
	) name2630 (
		\u12_o4_we_reg/P0001 ,
		\u4_mem_reg[2][20]/NET0131 ,
		\u4_wp_reg[0]/P0001 ,
		\u4_wp_reg[1]/NET0131 ,
		_w4777_
	);
	LUT4 #(
		.INIT('h0800)
	) name2631 (
		\u12_dout_reg[20]/P0001 ,
		\u12_o4_we_reg/P0001 ,
		\u4_wp_reg[0]/P0001 ,
		\u4_wp_reg[1]/NET0131 ,
		_w4778_
	);
	LUT2 #(
		.INIT('he)
	) name2632 (
		_w4777_,
		_w4778_,
		_w4779_
	);
	LUT4 #(
		.INIT('hc4cc)
	) name2633 (
		\u12_o4_we_reg/P0001 ,
		\u4_mem_reg[2][21]/NET0131 ,
		\u4_wp_reg[0]/P0001 ,
		\u4_wp_reg[1]/NET0131 ,
		_w4780_
	);
	LUT4 #(
		.INIT('h0800)
	) name2634 (
		\u12_dout_reg[21]/P0001 ,
		\u12_o4_we_reg/P0001 ,
		\u4_wp_reg[0]/P0001 ,
		\u4_wp_reg[1]/NET0131 ,
		_w4781_
	);
	LUT2 #(
		.INIT('he)
	) name2635 (
		_w4780_,
		_w4781_,
		_w4782_
	);
	LUT4 #(
		.INIT('hc4cc)
	) name2636 (
		\u12_o4_we_reg/P0001 ,
		\u4_mem_reg[2][22]/NET0131 ,
		\u4_wp_reg[0]/P0001 ,
		\u4_wp_reg[1]/NET0131 ,
		_w4783_
	);
	LUT4 #(
		.INIT('h0800)
	) name2637 (
		\u12_dout_reg[22]/P0001 ,
		\u12_o4_we_reg/P0001 ,
		\u4_wp_reg[0]/P0001 ,
		\u4_wp_reg[1]/NET0131 ,
		_w4784_
	);
	LUT2 #(
		.INIT('he)
	) name2638 (
		_w4783_,
		_w4784_,
		_w4785_
	);
	LUT4 #(
		.INIT('hc4cc)
	) name2639 (
		\u12_o4_we_reg/P0001 ,
		\u4_mem_reg[2][23]/NET0131 ,
		\u4_wp_reg[0]/P0001 ,
		\u4_wp_reg[1]/NET0131 ,
		_w4786_
	);
	LUT4 #(
		.INIT('h0800)
	) name2640 (
		\u12_dout_reg[23]/P0001 ,
		\u12_o4_we_reg/P0001 ,
		\u4_wp_reg[0]/P0001 ,
		\u4_wp_reg[1]/NET0131 ,
		_w4787_
	);
	LUT2 #(
		.INIT('he)
	) name2641 (
		_w4786_,
		_w4787_,
		_w4788_
	);
	LUT4 #(
		.INIT('hc4cc)
	) name2642 (
		\u12_o4_we_reg/P0001 ,
		\u4_mem_reg[2][24]/NET0131 ,
		\u4_wp_reg[0]/P0001 ,
		\u4_wp_reg[1]/NET0131 ,
		_w4789_
	);
	LUT4 #(
		.INIT('h0800)
	) name2643 (
		\u12_dout_reg[24]/P0001 ,
		\u12_o4_we_reg/P0001 ,
		\u4_wp_reg[0]/P0001 ,
		\u4_wp_reg[1]/NET0131 ,
		_w4790_
	);
	LUT2 #(
		.INIT('he)
	) name2644 (
		_w4789_,
		_w4790_,
		_w4791_
	);
	LUT4 #(
		.INIT('hc4cc)
	) name2645 (
		\u12_o4_we_reg/P0001 ,
		\u4_mem_reg[2][25]/NET0131 ,
		\u4_wp_reg[0]/P0001 ,
		\u4_wp_reg[1]/NET0131 ,
		_w4792_
	);
	LUT4 #(
		.INIT('h0800)
	) name2646 (
		\u12_dout_reg[25]/P0001 ,
		\u12_o4_we_reg/P0001 ,
		\u4_wp_reg[0]/P0001 ,
		\u4_wp_reg[1]/NET0131 ,
		_w4793_
	);
	LUT2 #(
		.INIT('he)
	) name2647 (
		_w4792_,
		_w4793_,
		_w4794_
	);
	LUT4 #(
		.INIT('hc4cc)
	) name2648 (
		\u12_o4_we_reg/P0001 ,
		\u4_mem_reg[2][26]/NET0131 ,
		\u4_wp_reg[0]/P0001 ,
		\u4_wp_reg[1]/NET0131 ,
		_w4795_
	);
	LUT4 #(
		.INIT('h0800)
	) name2649 (
		\u12_dout_reg[26]/P0001 ,
		\u12_o4_we_reg/P0001 ,
		\u4_wp_reg[0]/P0001 ,
		\u4_wp_reg[1]/NET0131 ,
		_w4796_
	);
	LUT2 #(
		.INIT('he)
	) name2650 (
		_w4795_,
		_w4796_,
		_w4797_
	);
	LUT4 #(
		.INIT('hc4cc)
	) name2651 (
		\u12_o4_we_reg/P0001 ,
		\u4_mem_reg[2][27]/NET0131 ,
		\u4_wp_reg[0]/P0001 ,
		\u4_wp_reg[1]/NET0131 ,
		_w4798_
	);
	LUT4 #(
		.INIT('h0800)
	) name2652 (
		\u12_dout_reg[27]/P0001 ,
		\u12_o4_we_reg/P0001 ,
		\u4_wp_reg[0]/P0001 ,
		\u4_wp_reg[1]/NET0131 ,
		_w4799_
	);
	LUT2 #(
		.INIT('he)
	) name2653 (
		_w4798_,
		_w4799_,
		_w4800_
	);
	LUT4 #(
		.INIT('hc4cc)
	) name2654 (
		\u12_o4_we_reg/P0001 ,
		\u4_mem_reg[2][28]/NET0131 ,
		\u4_wp_reg[0]/P0001 ,
		\u4_wp_reg[1]/NET0131 ,
		_w4801_
	);
	LUT4 #(
		.INIT('h0800)
	) name2655 (
		\u12_dout_reg[28]/P0001 ,
		\u12_o4_we_reg/P0001 ,
		\u4_wp_reg[0]/P0001 ,
		\u4_wp_reg[1]/NET0131 ,
		_w4802_
	);
	LUT2 #(
		.INIT('he)
	) name2656 (
		_w4801_,
		_w4802_,
		_w4803_
	);
	LUT4 #(
		.INIT('hc4cc)
	) name2657 (
		\u12_o4_we_reg/P0001 ,
		\u4_mem_reg[2][29]/NET0131 ,
		\u4_wp_reg[0]/P0001 ,
		\u4_wp_reg[1]/NET0131 ,
		_w4804_
	);
	LUT4 #(
		.INIT('h0800)
	) name2658 (
		\u12_dout_reg[29]/P0001 ,
		\u12_o4_we_reg/P0001 ,
		\u4_wp_reg[0]/P0001 ,
		\u4_wp_reg[1]/NET0131 ,
		_w4805_
	);
	LUT2 #(
		.INIT('he)
	) name2659 (
		_w4804_,
		_w4805_,
		_w4806_
	);
	LUT4 #(
		.INIT('hc4cc)
	) name2660 (
		\u12_o4_we_reg/P0001 ,
		\u4_mem_reg[2][2]/NET0131 ,
		\u4_wp_reg[0]/P0001 ,
		\u4_wp_reg[1]/NET0131 ,
		_w4807_
	);
	LUT4 #(
		.INIT('h0800)
	) name2661 (
		\u12_dout_reg[2]/P0001 ,
		\u12_o4_we_reg/P0001 ,
		\u4_wp_reg[0]/P0001 ,
		\u4_wp_reg[1]/NET0131 ,
		_w4808_
	);
	LUT2 #(
		.INIT('he)
	) name2662 (
		_w4807_,
		_w4808_,
		_w4809_
	);
	LUT4 #(
		.INIT('hc4cc)
	) name2663 (
		\u12_o4_we_reg/P0001 ,
		\u4_mem_reg[2][30]/NET0131 ,
		\u4_wp_reg[0]/P0001 ,
		\u4_wp_reg[1]/NET0131 ,
		_w4810_
	);
	LUT4 #(
		.INIT('h0800)
	) name2664 (
		\u12_dout_reg[30]/P0001 ,
		\u12_o4_we_reg/P0001 ,
		\u4_wp_reg[0]/P0001 ,
		\u4_wp_reg[1]/NET0131 ,
		_w4811_
	);
	LUT2 #(
		.INIT('he)
	) name2665 (
		_w4810_,
		_w4811_,
		_w4812_
	);
	LUT4 #(
		.INIT('hc4cc)
	) name2666 (
		\u12_o4_we_reg/P0001 ,
		\u4_mem_reg[2][31]/NET0131 ,
		\u4_wp_reg[0]/P0001 ,
		\u4_wp_reg[1]/NET0131 ,
		_w4813_
	);
	LUT4 #(
		.INIT('h0800)
	) name2667 (
		\u12_dout_reg[31]/P0001 ,
		\u12_o4_we_reg/P0001 ,
		\u4_wp_reg[0]/P0001 ,
		\u4_wp_reg[1]/NET0131 ,
		_w4814_
	);
	LUT2 #(
		.INIT('he)
	) name2668 (
		_w4813_,
		_w4814_,
		_w4815_
	);
	LUT4 #(
		.INIT('hc4cc)
	) name2669 (
		\u12_o4_we_reg/P0001 ,
		\u4_mem_reg[2][3]/NET0131 ,
		\u4_wp_reg[0]/P0001 ,
		\u4_wp_reg[1]/NET0131 ,
		_w4816_
	);
	LUT4 #(
		.INIT('h0800)
	) name2670 (
		\u12_dout_reg[3]/P0001 ,
		\u12_o4_we_reg/P0001 ,
		\u4_wp_reg[0]/P0001 ,
		\u4_wp_reg[1]/NET0131 ,
		_w4817_
	);
	LUT2 #(
		.INIT('he)
	) name2671 (
		_w4816_,
		_w4817_,
		_w4818_
	);
	LUT4 #(
		.INIT('hc4cc)
	) name2672 (
		\u12_o4_we_reg/P0001 ,
		\u4_mem_reg[2][4]/NET0131 ,
		\u4_wp_reg[0]/P0001 ,
		\u4_wp_reg[1]/NET0131 ,
		_w4819_
	);
	LUT4 #(
		.INIT('h0800)
	) name2673 (
		\u12_dout_reg[4]/P0001 ,
		\u12_o4_we_reg/P0001 ,
		\u4_wp_reg[0]/P0001 ,
		\u4_wp_reg[1]/NET0131 ,
		_w4820_
	);
	LUT2 #(
		.INIT('he)
	) name2674 (
		_w4819_,
		_w4820_,
		_w4821_
	);
	LUT4 #(
		.INIT('hc4cc)
	) name2675 (
		\u12_o4_we_reg/P0001 ,
		\u4_mem_reg[2][5]/NET0131 ,
		\u4_wp_reg[0]/P0001 ,
		\u4_wp_reg[1]/NET0131 ,
		_w4822_
	);
	LUT4 #(
		.INIT('h0800)
	) name2676 (
		\u12_dout_reg[5]/P0001 ,
		\u12_o4_we_reg/P0001 ,
		\u4_wp_reg[0]/P0001 ,
		\u4_wp_reg[1]/NET0131 ,
		_w4823_
	);
	LUT2 #(
		.INIT('he)
	) name2677 (
		_w4822_,
		_w4823_,
		_w4824_
	);
	LUT4 #(
		.INIT('hc4cc)
	) name2678 (
		\u12_o4_we_reg/P0001 ,
		\u4_mem_reg[2][6]/NET0131 ,
		\u4_wp_reg[0]/P0001 ,
		\u4_wp_reg[1]/NET0131 ,
		_w4825_
	);
	LUT4 #(
		.INIT('h0800)
	) name2679 (
		\u12_dout_reg[6]/P0001 ,
		\u12_o4_we_reg/P0001 ,
		\u4_wp_reg[0]/P0001 ,
		\u4_wp_reg[1]/NET0131 ,
		_w4826_
	);
	LUT2 #(
		.INIT('he)
	) name2680 (
		_w4825_,
		_w4826_,
		_w4827_
	);
	LUT4 #(
		.INIT('hc4cc)
	) name2681 (
		\u12_o4_we_reg/P0001 ,
		\u4_mem_reg[2][7]/NET0131 ,
		\u4_wp_reg[0]/P0001 ,
		\u4_wp_reg[1]/NET0131 ,
		_w4828_
	);
	LUT4 #(
		.INIT('h0800)
	) name2682 (
		\u12_dout_reg[7]/P0001 ,
		\u12_o4_we_reg/P0001 ,
		\u4_wp_reg[0]/P0001 ,
		\u4_wp_reg[1]/NET0131 ,
		_w4829_
	);
	LUT2 #(
		.INIT('he)
	) name2683 (
		_w4828_,
		_w4829_,
		_w4830_
	);
	LUT4 #(
		.INIT('hc4cc)
	) name2684 (
		\u12_o4_we_reg/P0001 ,
		\u4_mem_reg[2][8]/NET0131 ,
		\u4_wp_reg[0]/P0001 ,
		\u4_wp_reg[1]/NET0131 ,
		_w4831_
	);
	LUT4 #(
		.INIT('h0800)
	) name2685 (
		\u12_dout_reg[8]/P0001 ,
		\u12_o4_we_reg/P0001 ,
		\u4_wp_reg[0]/P0001 ,
		\u4_wp_reg[1]/NET0131 ,
		_w4832_
	);
	LUT2 #(
		.INIT('he)
	) name2686 (
		_w4831_,
		_w4832_,
		_w4833_
	);
	LUT4 #(
		.INIT('hc4cc)
	) name2687 (
		\u12_o4_we_reg/P0001 ,
		\u4_mem_reg[2][9]/NET0131 ,
		\u4_wp_reg[0]/P0001 ,
		\u4_wp_reg[1]/NET0131 ,
		_w4834_
	);
	LUT4 #(
		.INIT('h0800)
	) name2688 (
		\u12_dout_reg[9]/P0001 ,
		\u12_o4_we_reg/P0001 ,
		\u4_wp_reg[0]/P0001 ,
		\u4_wp_reg[1]/NET0131 ,
		_w4835_
	);
	LUT2 #(
		.INIT('he)
	) name2689 (
		_w4834_,
		_w4835_,
		_w4836_
	);
	LUT4 #(
		.INIT('h4ccc)
	) name2690 (
		\u12_o4_we_reg/P0001 ,
		\u4_mem_reg[3][0]/NET0131 ,
		\u4_wp_reg[0]/P0001 ,
		\u4_wp_reg[1]/NET0131 ,
		_w4837_
	);
	LUT4 #(
		.INIT('h8000)
	) name2691 (
		\u12_dout_reg[0]/P0001 ,
		\u12_o4_we_reg/P0001 ,
		\u4_wp_reg[0]/P0001 ,
		\u4_wp_reg[1]/NET0131 ,
		_w4838_
	);
	LUT2 #(
		.INIT('he)
	) name2692 (
		_w4837_,
		_w4838_,
		_w4839_
	);
	LUT4 #(
		.INIT('h4ccc)
	) name2693 (
		\u12_o4_we_reg/P0001 ,
		\u4_mem_reg[3][10]/NET0131 ,
		\u4_wp_reg[0]/P0001 ,
		\u4_wp_reg[1]/NET0131 ,
		_w4840_
	);
	LUT4 #(
		.INIT('h8000)
	) name2694 (
		\u12_dout_reg[10]/P0001 ,
		\u12_o4_we_reg/P0001 ,
		\u4_wp_reg[0]/P0001 ,
		\u4_wp_reg[1]/NET0131 ,
		_w4841_
	);
	LUT2 #(
		.INIT('he)
	) name2695 (
		_w4840_,
		_w4841_,
		_w4842_
	);
	LUT4 #(
		.INIT('h4ccc)
	) name2696 (
		\u12_o4_we_reg/P0001 ,
		\u4_mem_reg[3][11]/NET0131 ,
		\u4_wp_reg[0]/P0001 ,
		\u4_wp_reg[1]/NET0131 ,
		_w4843_
	);
	LUT4 #(
		.INIT('h8000)
	) name2697 (
		\u12_dout_reg[11]/P0001 ,
		\u12_o4_we_reg/P0001 ,
		\u4_wp_reg[0]/P0001 ,
		\u4_wp_reg[1]/NET0131 ,
		_w4844_
	);
	LUT2 #(
		.INIT('he)
	) name2698 (
		_w4843_,
		_w4844_,
		_w4845_
	);
	LUT4 #(
		.INIT('h4ccc)
	) name2699 (
		\u12_o4_we_reg/P0001 ,
		\u4_mem_reg[3][12]/NET0131 ,
		\u4_wp_reg[0]/P0001 ,
		\u4_wp_reg[1]/NET0131 ,
		_w4846_
	);
	LUT4 #(
		.INIT('h8000)
	) name2700 (
		\u12_dout_reg[12]/P0001 ,
		\u12_o4_we_reg/P0001 ,
		\u4_wp_reg[0]/P0001 ,
		\u4_wp_reg[1]/NET0131 ,
		_w4847_
	);
	LUT2 #(
		.INIT('he)
	) name2701 (
		_w4846_,
		_w4847_,
		_w4848_
	);
	LUT4 #(
		.INIT('h4ccc)
	) name2702 (
		\u12_o4_we_reg/P0001 ,
		\u4_mem_reg[3][13]/NET0131 ,
		\u4_wp_reg[0]/P0001 ,
		\u4_wp_reg[1]/NET0131 ,
		_w4849_
	);
	LUT4 #(
		.INIT('h8000)
	) name2703 (
		\u12_dout_reg[13]/P0001 ,
		\u12_o4_we_reg/P0001 ,
		\u4_wp_reg[0]/P0001 ,
		\u4_wp_reg[1]/NET0131 ,
		_w4850_
	);
	LUT2 #(
		.INIT('he)
	) name2704 (
		_w4849_,
		_w4850_,
		_w4851_
	);
	LUT4 #(
		.INIT('h4ccc)
	) name2705 (
		\u12_o4_we_reg/P0001 ,
		\u4_mem_reg[3][14]/NET0131 ,
		\u4_wp_reg[0]/P0001 ,
		\u4_wp_reg[1]/NET0131 ,
		_w4852_
	);
	LUT4 #(
		.INIT('h8000)
	) name2706 (
		\u12_dout_reg[14]/P0001 ,
		\u12_o4_we_reg/P0001 ,
		\u4_wp_reg[0]/P0001 ,
		\u4_wp_reg[1]/NET0131 ,
		_w4853_
	);
	LUT2 #(
		.INIT('he)
	) name2707 (
		_w4852_,
		_w4853_,
		_w4854_
	);
	LUT4 #(
		.INIT('h4ccc)
	) name2708 (
		\u12_o4_we_reg/P0001 ,
		\u4_mem_reg[3][15]/NET0131 ,
		\u4_wp_reg[0]/P0001 ,
		\u4_wp_reg[1]/NET0131 ,
		_w4855_
	);
	LUT4 #(
		.INIT('h8000)
	) name2709 (
		\u12_dout_reg[15]/P0001 ,
		\u12_o4_we_reg/P0001 ,
		\u4_wp_reg[0]/P0001 ,
		\u4_wp_reg[1]/NET0131 ,
		_w4856_
	);
	LUT2 #(
		.INIT('he)
	) name2710 (
		_w4855_,
		_w4856_,
		_w4857_
	);
	LUT4 #(
		.INIT('h4ccc)
	) name2711 (
		\u12_o4_we_reg/P0001 ,
		\u4_mem_reg[3][16]/NET0131 ,
		\u4_wp_reg[0]/P0001 ,
		\u4_wp_reg[1]/NET0131 ,
		_w4858_
	);
	LUT4 #(
		.INIT('h8000)
	) name2712 (
		\u12_dout_reg[16]/P0001 ,
		\u12_o4_we_reg/P0001 ,
		\u4_wp_reg[0]/P0001 ,
		\u4_wp_reg[1]/NET0131 ,
		_w4859_
	);
	LUT2 #(
		.INIT('he)
	) name2713 (
		_w4858_,
		_w4859_,
		_w4860_
	);
	LUT4 #(
		.INIT('h4ccc)
	) name2714 (
		\u12_o4_we_reg/P0001 ,
		\u4_mem_reg[3][17]/NET0131 ,
		\u4_wp_reg[0]/P0001 ,
		\u4_wp_reg[1]/NET0131 ,
		_w4861_
	);
	LUT4 #(
		.INIT('h8000)
	) name2715 (
		\u12_dout_reg[17]/P0001 ,
		\u12_o4_we_reg/P0001 ,
		\u4_wp_reg[0]/P0001 ,
		\u4_wp_reg[1]/NET0131 ,
		_w4862_
	);
	LUT2 #(
		.INIT('he)
	) name2716 (
		_w4861_,
		_w4862_,
		_w4863_
	);
	LUT4 #(
		.INIT('h4ccc)
	) name2717 (
		\u12_o4_we_reg/P0001 ,
		\u4_mem_reg[3][18]/NET0131 ,
		\u4_wp_reg[0]/P0001 ,
		\u4_wp_reg[1]/NET0131 ,
		_w4864_
	);
	LUT4 #(
		.INIT('h8000)
	) name2718 (
		\u12_dout_reg[18]/P0001 ,
		\u12_o4_we_reg/P0001 ,
		\u4_wp_reg[0]/P0001 ,
		\u4_wp_reg[1]/NET0131 ,
		_w4865_
	);
	LUT2 #(
		.INIT('he)
	) name2719 (
		_w4864_,
		_w4865_,
		_w4866_
	);
	LUT4 #(
		.INIT('h4ccc)
	) name2720 (
		\u12_o4_we_reg/P0001 ,
		\u4_mem_reg[3][19]/NET0131 ,
		\u4_wp_reg[0]/P0001 ,
		\u4_wp_reg[1]/NET0131 ,
		_w4867_
	);
	LUT4 #(
		.INIT('h8000)
	) name2721 (
		\u12_dout_reg[19]/P0001 ,
		\u12_o4_we_reg/P0001 ,
		\u4_wp_reg[0]/P0001 ,
		\u4_wp_reg[1]/NET0131 ,
		_w4868_
	);
	LUT2 #(
		.INIT('he)
	) name2722 (
		_w4867_,
		_w4868_,
		_w4869_
	);
	LUT4 #(
		.INIT('h4ccc)
	) name2723 (
		\u12_o4_we_reg/P0001 ,
		\u4_mem_reg[3][1]/NET0131 ,
		\u4_wp_reg[0]/P0001 ,
		\u4_wp_reg[1]/NET0131 ,
		_w4870_
	);
	LUT4 #(
		.INIT('h8000)
	) name2724 (
		\u12_dout_reg[1]/P0001 ,
		\u12_o4_we_reg/P0001 ,
		\u4_wp_reg[0]/P0001 ,
		\u4_wp_reg[1]/NET0131 ,
		_w4871_
	);
	LUT2 #(
		.INIT('he)
	) name2725 (
		_w4870_,
		_w4871_,
		_w4872_
	);
	LUT4 #(
		.INIT('h4ccc)
	) name2726 (
		\u12_o4_we_reg/P0001 ,
		\u4_mem_reg[3][20]/NET0131 ,
		\u4_wp_reg[0]/P0001 ,
		\u4_wp_reg[1]/NET0131 ,
		_w4873_
	);
	LUT4 #(
		.INIT('h8000)
	) name2727 (
		\u12_dout_reg[20]/P0001 ,
		\u12_o4_we_reg/P0001 ,
		\u4_wp_reg[0]/P0001 ,
		\u4_wp_reg[1]/NET0131 ,
		_w4874_
	);
	LUT2 #(
		.INIT('he)
	) name2728 (
		_w4873_,
		_w4874_,
		_w4875_
	);
	LUT4 #(
		.INIT('h4ccc)
	) name2729 (
		\u12_o4_we_reg/P0001 ,
		\u4_mem_reg[3][21]/NET0131 ,
		\u4_wp_reg[0]/P0001 ,
		\u4_wp_reg[1]/NET0131 ,
		_w4876_
	);
	LUT4 #(
		.INIT('h8000)
	) name2730 (
		\u12_dout_reg[21]/P0001 ,
		\u12_o4_we_reg/P0001 ,
		\u4_wp_reg[0]/P0001 ,
		\u4_wp_reg[1]/NET0131 ,
		_w4877_
	);
	LUT2 #(
		.INIT('he)
	) name2731 (
		_w4876_,
		_w4877_,
		_w4878_
	);
	LUT4 #(
		.INIT('h4ccc)
	) name2732 (
		\u12_o4_we_reg/P0001 ,
		\u4_mem_reg[3][22]/NET0131 ,
		\u4_wp_reg[0]/P0001 ,
		\u4_wp_reg[1]/NET0131 ,
		_w4879_
	);
	LUT4 #(
		.INIT('h8000)
	) name2733 (
		\u12_dout_reg[22]/P0001 ,
		\u12_o4_we_reg/P0001 ,
		\u4_wp_reg[0]/P0001 ,
		\u4_wp_reg[1]/NET0131 ,
		_w4880_
	);
	LUT2 #(
		.INIT('he)
	) name2734 (
		_w4879_,
		_w4880_,
		_w4881_
	);
	LUT4 #(
		.INIT('h4ccc)
	) name2735 (
		\u12_o4_we_reg/P0001 ,
		\u4_mem_reg[3][23]/NET0131 ,
		\u4_wp_reg[0]/P0001 ,
		\u4_wp_reg[1]/NET0131 ,
		_w4882_
	);
	LUT4 #(
		.INIT('h8000)
	) name2736 (
		\u12_dout_reg[23]/P0001 ,
		\u12_o4_we_reg/P0001 ,
		\u4_wp_reg[0]/P0001 ,
		\u4_wp_reg[1]/NET0131 ,
		_w4883_
	);
	LUT2 #(
		.INIT('he)
	) name2737 (
		_w4882_,
		_w4883_,
		_w4884_
	);
	LUT4 #(
		.INIT('h4ccc)
	) name2738 (
		\u12_o4_we_reg/P0001 ,
		\u4_mem_reg[3][24]/NET0131 ,
		\u4_wp_reg[0]/P0001 ,
		\u4_wp_reg[1]/NET0131 ,
		_w4885_
	);
	LUT4 #(
		.INIT('h8000)
	) name2739 (
		\u12_dout_reg[24]/P0001 ,
		\u12_o4_we_reg/P0001 ,
		\u4_wp_reg[0]/P0001 ,
		\u4_wp_reg[1]/NET0131 ,
		_w4886_
	);
	LUT2 #(
		.INIT('he)
	) name2740 (
		_w4885_,
		_w4886_,
		_w4887_
	);
	LUT4 #(
		.INIT('h4ccc)
	) name2741 (
		\u12_o4_we_reg/P0001 ,
		\u4_mem_reg[3][25]/NET0131 ,
		\u4_wp_reg[0]/P0001 ,
		\u4_wp_reg[1]/NET0131 ,
		_w4888_
	);
	LUT4 #(
		.INIT('h8000)
	) name2742 (
		\u12_dout_reg[25]/P0001 ,
		\u12_o4_we_reg/P0001 ,
		\u4_wp_reg[0]/P0001 ,
		\u4_wp_reg[1]/NET0131 ,
		_w4889_
	);
	LUT2 #(
		.INIT('he)
	) name2743 (
		_w4888_,
		_w4889_,
		_w4890_
	);
	LUT4 #(
		.INIT('h4ccc)
	) name2744 (
		\u12_o4_we_reg/P0001 ,
		\u4_mem_reg[3][26]/NET0131 ,
		\u4_wp_reg[0]/P0001 ,
		\u4_wp_reg[1]/NET0131 ,
		_w4891_
	);
	LUT4 #(
		.INIT('h8000)
	) name2745 (
		\u12_dout_reg[26]/P0001 ,
		\u12_o4_we_reg/P0001 ,
		\u4_wp_reg[0]/P0001 ,
		\u4_wp_reg[1]/NET0131 ,
		_w4892_
	);
	LUT2 #(
		.INIT('he)
	) name2746 (
		_w4891_,
		_w4892_,
		_w4893_
	);
	LUT4 #(
		.INIT('h4ccc)
	) name2747 (
		\u12_o4_we_reg/P0001 ,
		\u4_mem_reg[3][27]/NET0131 ,
		\u4_wp_reg[0]/P0001 ,
		\u4_wp_reg[1]/NET0131 ,
		_w4894_
	);
	LUT4 #(
		.INIT('h8000)
	) name2748 (
		\u12_dout_reg[27]/P0001 ,
		\u12_o4_we_reg/P0001 ,
		\u4_wp_reg[0]/P0001 ,
		\u4_wp_reg[1]/NET0131 ,
		_w4895_
	);
	LUT2 #(
		.INIT('he)
	) name2749 (
		_w4894_,
		_w4895_,
		_w4896_
	);
	LUT4 #(
		.INIT('h4ccc)
	) name2750 (
		\u12_o4_we_reg/P0001 ,
		\u4_mem_reg[3][28]/NET0131 ,
		\u4_wp_reg[0]/P0001 ,
		\u4_wp_reg[1]/NET0131 ,
		_w4897_
	);
	LUT4 #(
		.INIT('h8000)
	) name2751 (
		\u12_dout_reg[28]/P0001 ,
		\u12_o4_we_reg/P0001 ,
		\u4_wp_reg[0]/P0001 ,
		\u4_wp_reg[1]/NET0131 ,
		_w4898_
	);
	LUT2 #(
		.INIT('he)
	) name2752 (
		_w4897_,
		_w4898_,
		_w4899_
	);
	LUT4 #(
		.INIT('h4ccc)
	) name2753 (
		\u12_o4_we_reg/P0001 ,
		\u4_mem_reg[3][29]/NET0131 ,
		\u4_wp_reg[0]/P0001 ,
		\u4_wp_reg[1]/NET0131 ,
		_w4900_
	);
	LUT4 #(
		.INIT('h8000)
	) name2754 (
		\u12_dout_reg[29]/P0001 ,
		\u12_o4_we_reg/P0001 ,
		\u4_wp_reg[0]/P0001 ,
		\u4_wp_reg[1]/NET0131 ,
		_w4901_
	);
	LUT2 #(
		.INIT('he)
	) name2755 (
		_w4900_,
		_w4901_,
		_w4902_
	);
	LUT4 #(
		.INIT('h4ccc)
	) name2756 (
		\u12_o4_we_reg/P0001 ,
		\u4_mem_reg[3][2]/NET0131 ,
		\u4_wp_reg[0]/P0001 ,
		\u4_wp_reg[1]/NET0131 ,
		_w4903_
	);
	LUT4 #(
		.INIT('h8000)
	) name2757 (
		\u12_dout_reg[2]/P0001 ,
		\u12_o4_we_reg/P0001 ,
		\u4_wp_reg[0]/P0001 ,
		\u4_wp_reg[1]/NET0131 ,
		_w4904_
	);
	LUT2 #(
		.INIT('he)
	) name2758 (
		_w4903_,
		_w4904_,
		_w4905_
	);
	LUT4 #(
		.INIT('h4ccc)
	) name2759 (
		\u12_o4_we_reg/P0001 ,
		\u4_mem_reg[3][30]/NET0131 ,
		\u4_wp_reg[0]/P0001 ,
		\u4_wp_reg[1]/NET0131 ,
		_w4906_
	);
	LUT4 #(
		.INIT('h8000)
	) name2760 (
		\u12_dout_reg[30]/P0001 ,
		\u12_o4_we_reg/P0001 ,
		\u4_wp_reg[0]/P0001 ,
		\u4_wp_reg[1]/NET0131 ,
		_w4907_
	);
	LUT2 #(
		.INIT('he)
	) name2761 (
		_w4906_,
		_w4907_,
		_w4908_
	);
	LUT4 #(
		.INIT('h4ccc)
	) name2762 (
		\u12_o4_we_reg/P0001 ,
		\u4_mem_reg[3][31]/NET0131 ,
		\u4_wp_reg[0]/P0001 ,
		\u4_wp_reg[1]/NET0131 ,
		_w4909_
	);
	LUT4 #(
		.INIT('h8000)
	) name2763 (
		\u12_dout_reg[31]/P0001 ,
		\u12_o4_we_reg/P0001 ,
		\u4_wp_reg[0]/P0001 ,
		\u4_wp_reg[1]/NET0131 ,
		_w4910_
	);
	LUT2 #(
		.INIT('he)
	) name2764 (
		_w4909_,
		_w4910_,
		_w4911_
	);
	LUT4 #(
		.INIT('h4ccc)
	) name2765 (
		\u12_o4_we_reg/P0001 ,
		\u4_mem_reg[3][3]/NET0131 ,
		\u4_wp_reg[0]/P0001 ,
		\u4_wp_reg[1]/NET0131 ,
		_w4912_
	);
	LUT4 #(
		.INIT('h8000)
	) name2766 (
		\u12_dout_reg[3]/P0001 ,
		\u12_o4_we_reg/P0001 ,
		\u4_wp_reg[0]/P0001 ,
		\u4_wp_reg[1]/NET0131 ,
		_w4913_
	);
	LUT2 #(
		.INIT('he)
	) name2767 (
		_w4912_,
		_w4913_,
		_w4914_
	);
	LUT4 #(
		.INIT('h4ccc)
	) name2768 (
		\u12_o4_we_reg/P0001 ,
		\u4_mem_reg[3][4]/NET0131 ,
		\u4_wp_reg[0]/P0001 ,
		\u4_wp_reg[1]/NET0131 ,
		_w4915_
	);
	LUT4 #(
		.INIT('h8000)
	) name2769 (
		\u12_dout_reg[4]/P0001 ,
		\u12_o4_we_reg/P0001 ,
		\u4_wp_reg[0]/P0001 ,
		\u4_wp_reg[1]/NET0131 ,
		_w4916_
	);
	LUT2 #(
		.INIT('he)
	) name2770 (
		_w4915_,
		_w4916_,
		_w4917_
	);
	LUT4 #(
		.INIT('h4ccc)
	) name2771 (
		\u12_o4_we_reg/P0001 ,
		\u4_mem_reg[3][5]/NET0131 ,
		\u4_wp_reg[0]/P0001 ,
		\u4_wp_reg[1]/NET0131 ,
		_w4918_
	);
	LUT4 #(
		.INIT('h8000)
	) name2772 (
		\u12_dout_reg[5]/P0001 ,
		\u12_o4_we_reg/P0001 ,
		\u4_wp_reg[0]/P0001 ,
		\u4_wp_reg[1]/NET0131 ,
		_w4919_
	);
	LUT2 #(
		.INIT('he)
	) name2773 (
		_w4918_,
		_w4919_,
		_w4920_
	);
	LUT4 #(
		.INIT('h4ccc)
	) name2774 (
		\u12_o4_we_reg/P0001 ,
		\u4_mem_reg[3][6]/NET0131 ,
		\u4_wp_reg[0]/P0001 ,
		\u4_wp_reg[1]/NET0131 ,
		_w4921_
	);
	LUT4 #(
		.INIT('h8000)
	) name2775 (
		\u12_dout_reg[6]/P0001 ,
		\u12_o4_we_reg/P0001 ,
		\u4_wp_reg[0]/P0001 ,
		\u4_wp_reg[1]/NET0131 ,
		_w4922_
	);
	LUT2 #(
		.INIT('he)
	) name2776 (
		_w4921_,
		_w4922_,
		_w4923_
	);
	LUT4 #(
		.INIT('h4ccc)
	) name2777 (
		\u12_o4_we_reg/P0001 ,
		\u4_mem_reg[3][7]/NET0131 ,
		\u4_wp_reg[0]/P0001 ,
		\u4_wp_reg[1]/NET0131 ,
		_w4924_
	);
	LUT4 #(
		.INIT('h8000)
	) name2778 (
		\u12_dout_reg[7]/P0001 ,
		\u12_o4_we_reg/P0001 ,
		\u4_wp_reg[0]/P0001 ,
		\u4_wp_reg[1]/NET0131 ,
		_w4925_
	);
	LUT2 #(
		.INIT('he)
	) name2779 (
		_w4924_,
		_w4925_,
		_w4926_
	);
	LUT4 #(
		.INIT('h4ccc)
	) name2780 (
		\u12_o4_we_reg/P0001 ,
		\u4_mem_reg[3][8]/NET0131 ,
		\u4_wp_reg[0]/P0001 ,
		\u4_wp_reg[1]/NET0131 ,
		_w4927_
	);
	LUT4 #(
		.INIT('h8000)
	) name2781 (
		\u12_dout_reg[8]/P0001 ,
		\u12_o4_we_reg/P0001 ,
		\u4_wp_reg[0]/P0001 ,
		\u4_wp_reg[1]/NET0131 ,
		_w4928_
	);
	LUT2 #(
		.INIT('he)
	) name2782 (
		_w4927_,
		_w4928_,
		_w4929_
	);
	LUT4 #(
		.INIT('h4ccc)
	) name2783 (
		\u12_o4_we_reg/P0001 ,
		\u4_mem_reg[3][9]/NET0131 ,
		\u4_wp_reg[0]/P0001 ,
		\u4_wp_reg[1]/NET0131 ,
		_w4930_
	);
	LUT4 #(
		.INIT('h8000)
	) name2784 (
		\u12_dout_reg[9]/P0001 ,
		\u12_o4_we_reg/P0001 ,
		\u4_wp_reg[0]/P0001 ,
		\u4_wp_reg[1]/NET0131 ,
		_w4931_
	);
	LUT2 #(
		.INIT('he)
	) name2785 (
		_w4930_,
		_w4931_,
		_w4932_
	);
	LUT4 #(
		.INIT('hc4cc)
	) name2786 (
		\u12_o3_we_reg/P0001 ,
		\u3_mem_reg[2][14]/NET0131 ,
		\u3_wp_reg[0]/P0001 ,
		\u3_wp_reg[1]/NET0131 ,
		_w4933_
	);
	LUT4 #(
		.INIT('h0800)
	) name2787 (
		\u12_dout_reg[14]/P0001 ,
		\u12_o3_we_reg/P0001 ,
		\u3_wp_reg[0]/P0001 ,
		\u3_wp_reg[1]/NET0131 ,
		_w4934_
	);
	LUT2 #(
		.INIT('he)
	) name2788 (
		_w4933_,
		_w4934_,
		_w4935_
	);
	LUT4 #(
		.INIT('hcc4c)
	) name2789 (
		\u12_o6_we_reg/P0001 ,
		\u5_mem_reg[1][0]/NET0131 ,
		\u5_wp_reg[0]/P0001 ,
		\u5_wp_reg[1]/NET0131 ,
		_w4936_
	);
	LUT4 #(
		.INIT('h0080)
	) name2790 (
		\u12_dout_reg[0]/P0001 ,
		\u12_o6_we_reg/P0001 ,
		\u5_wp_reg[0]/P0001 ,
		\u5_wp_reg[1]/NET0131 ,
		_w4937_
	);
	LUT2 #(
		.INIT('he)
	) name2791 (
		_w4936_,
		_w4937_,
		_w4938_
	);
	LUT4 #(
		.INIT('hcc4c)
	) name2792 (
		\u12_o6_we_reg/P0001 ,
		\u5_mem_reg[1][10]/NET0131 ,
		\u5_wp_reg[0]/P0001 ,
		\u5_wp_reg[1]/NET0131 ,
		_w4939_
	);
	LUT4 #(
		.INIT('h0080)
	) name2793 (
		\u12_dout_reg[10]/P0001 ,
		\u12_o6_we_reg/P0001 ,
		\u5_wp_reg[0]/P0001 ,
		\u5_wp_reg[1]/NET0131 ,
		_w4940_
	);
	LUT2 #(
		.INIT('he)
	) name2794 (
		_w4939_,
		_w4940_,
		_w4941_
	);
	LUT4 #(
		.INIT('hcc4c)
	) name2795 (
		\u12_o6_we_reg/P0001 ,
		\u5_mem_reg[1][11]/NET0131 ,
		\u5_wp_reg[0]/P0001 ,
		\u5_wp_reg[1]/NET0131 ,
		_w4942_
	);
	LUT4 #(
		.INIT('h0080)
	) name2796 (
		\u12_dout_reg[11]/P0001 ,
		\u12_o6_we_reg/P0001 ,
		\u5_wp_reg[0]/P0001 ,
		\u5_wp_reg[1]/NET0131 ,
		_w4943_
	);
	LUT2 #(
		.INIT('he)
	) name2797 (
		_w4942_,
		_w4943_,
		_w4944_
	);
	LUT4 #(
		.INIT('hcc4c)
	) name2798 (
		\u12_o6_we_reg/P0001 ,
		\u5_mem_reg[1][12]/NET0131 ,
		\u5_wp_reg[0]/P0001 ,
		\u5_wp_reg[1]/NET0131 ,
		_w4945_
	);
	LUT4 #(
		.INIT('h0080)
	) name2799 (
		\u12_dout_reg[12]/P0001 ,
		\u12_o6_we_reg/P0001 ,
		\u5_wp_reg[0]/P0001 ,
		\u5_wp_reg[1]/NET0131 ,
		_w4946_
	);
	LUT2 #(
		.INIT('he)
	) name2800 (
		_w4945_,
		_w4946_,
		_w4947_
	);
	LUT4 #(
		.INIT('hcc4c)
	) name2801 (
		\u12_o6_we_reg/P0001 ,
		\u5_mem_reg[1][13]/NET0131 ,
		\u5_wp_reg[0]/P0001 ,
		\u5_wp_reg[1]/NET0131 ,
		_w4948_
	);
	LUT4 #(
		.INIT('h0080)
	) name2802 (
		\u12_dout_reg[13]/P0001 ,
		\u12_o6_we_reg/P0001 ,
		\u5_wp_reg[0]/P0001 ,
		\u5_wp_reg[1]/NET0131 ,
		_w4949_
	);
	LUT2 #(
		.INIT('he)
	) name2803 (
		_w4948_,
		_w4949_,
		_w4950_
	);
	LUT4 #(
		.INIT('hcc4c)
	) name2804 (
		\u12_o6_we_reg/P0001 ,
		\u5_mem_reg[1][14]/NET0131 ,
		\u5_wp_reg[0]/P0001 ,
		\u5_wp_reg[1]/NET0131 ,
		_w4951_
	);
	LUT4 #(
		.INIT('h0080)
	) name2805 (
		\u12_dout_reg[14]/P0001 ,
		\u12_o6_we_reg/P0001 ,
		\u5_wp_reg[0]/P0001 ,
		\u5_wp_reg[1]/NET0131 ,
		_w4952_
	);
	LUT2 #(
		.INIT('he)
	) name2806 (
		_w4951_,
		_w4952_,
		_w4953_
	);
	LUT4 #(
		.INIT('hcc4c)
	) name2807 (
		\u12_o6_we_reg/P0001 ,
		\u5_mem_reg[1][15]/NET0131 ,
		\u5_wp_reg[0]/P0001 ,
		\u5_wp_reg[1]/NET0131 ,
		_w4954_
	);
	LUT4 #(
		.INIT('h0080)
	) name2808 (
		\u12_dout_reg[15]/P0001 ,
		\u12_o6_we_reg/P0001 ,
		\u5_wp_reg[0]/P0001 ,
		\u5_wp_reg[1]/NET0131 ,
		_w4955_
	);
	LUT2 #(
		.INIT('he)
	) name2809 (
		_w4954_,
		_w4955_,
		_w4956_
	);
	LUT4 #(
		.INIT('hcc4c)
	) name2810 (
		\u12_o6_we_reg/P0001 ,
		\u5_mem_reg[1][16]/NET0131 ,
		\u5_wp_reg[0]/P0001 ,
		\u5_wp_reg[1]/NET0131 ,
		_w4957_
	);
	LUT4 #(
		.INIT('h0080)
	) name2811 (
		\u12_dout_reg[16]/P0001 ,
		\u12_o6_we_reg/P0001 ,
		\u5_wp_reg[0]/P0001 ,
		\u5_wp_reg[1]/NET0131 ,
		_w4958_
	);
	LUT2 #(
		.INIT('he)
	) name2812 (
		_w4957_,
		_w4958_,
		_w4959_
	);
	LUT4 #(
		.INIT('hcc4c)
	) name2813 (
		\u12_o6_we_reg/P0001 ,
		\u5_mem_reg[1][17]/NET0131 ,
		\u5_wp_reg[0]/P0001 ,
		\u5_wp_reg[1]/NET0131 ,
		_w4960_
	);
	LUT4 #(
		.INIT('h0080)
	) name2814 (
		\u12_dout_reg[17]/P0001 ,
		\u12_o6_we_reg/P0001 ,
		\u5_wp_reg[0]/P0001 ,
		\u5_wp_reg[1]/NET0131 ,
		_w4961_
	);
	LUT2 #(
		.INIT('he)
	) name2815 (
		_w4960_,
		_w4961_,
		_w4962_
	);
	LUT4 #(
		.INIT('hcc4c)
	) name2816 (
		\u12_o6_we_reg/P0001 ,
		\u5_mem_reg[1][18]/NET0131 ,
		\u5_wp_reg[0]/P0001 ,
		\u5_wp_reg[1]/NET0131 ,
		_w4963_
	);
	LUT4 #(
		.INIT('h0080)
	) name2817 (
		\u12_dout_reg[18]/P0001 ,
		\u12_o6_we_reg/P0001 ,
		\u5_wp_reg[0]/P0001 ,
		\u5_wp_reg[1]/NET0131 ,
		_w4964_
	);
	LUT2 #(
		.INIT('he)
	) name2818 (
		_w4963_,
		_w4964_,
		_w4965_
	);
	LUT4 #(
		.INIT('hcc4c)
	) name2819 (
		\u12_o6_we_reg/P0001 ,
		\u5_mem_reg[1][19]/NET0131 ,
		\u5_wp_reg[0]/P0001 ,
		\u5_wp_reg[1]/NET0131 ,
		_w4966_
	);
	LUT4 #(
		.INIT('h0080)
	) name2820 (
		\u12_dout_reg[19]/P0001 ,
		\u12_o6_we_reg/P0001 ,
		\u5_wp_reg[0]/P0001 ,
		\u5_wp_reg[1]/NET0131 ,
		_w4967_
	);
	LUT2 #(
		.INIT('he)
	) name2821 (
		_w4966_,
		_w4967_,
		_w4968_
	);
	LUT4 #(
		.INIT('hcc4c)
	) name2822 (
		\u12_o6_we_reg/P0001 ,
		\u5_mem_reg[1][1]/NET0131 ,
		\u5_wp_reg[0]/P0001 ,
		\u5_wp_reg[1]/NET0131 ,
		_w4969_
	);
	LUT4 #(
		.INIT('h0080)
	) name2823 (
		\u12_dout_reg[1]/P0001 ,
		\u12_o6_we_reg/P0001 ,
		\u5_wp_reg[0]/P0001 ,
		\u5_wp_reg[1]/NET0131 ,
		_w4970_
	);
	LUT2 #(
		.INIT('he)
	) name2824 (
		_w4969_,
		_w4970_,
		_w4971_
	);
	LUT4 #(
		.INIT('hcc4c)
	) name2825 (
		\u12_o6_we_reg/P0001 ,
		\u5_mem_reg[1][20]/NET0131 ,
		\u5_wp_reg[0]/P0001 ,
		\u5_wp_reg[1]/NET0131 ,
		_w4972_
	);
	LUT4 #(
		.INIT('h0080)
	) name2826 (
		\u12_dout_reg[20]/P0001 ,
		\u12_o6_we_reg/P0001 ,
		\u5_wp_reg[0]/P0001 ,
		\u5_wp_reg[1]/NET0131 ,
		_w4973_
	);
	LUT2 #(
		.INIT('he)
	) name2827 (
		_w4972_,
		_w4973_,
		_w4974_
	);
	LUT4 #(
		.INIT('hcc4c)
	) name2828 (
		\u12_o6_we_reg/P0001 ,
		\u5_mem_reg[1][21]/NET0131 ,
		\u5_wp_reg[0]/P0001 ,
		\u5_wp_reg[1]/NET0131 ,
		_w4975_
	);
	LUT4 #(
		.INIT('h0080)
	) name2829 (
		\u12_dout_reg[21]/P0001 ,
		\u12_o6_we_reg/P0001 ,
		\u5_wp_reg[0]/P0001 ,
		\u5_wp_reg[1]/NET0131 ,
		_w4976_
	);
	LUT2 #(
		.INIT('he)
	) name2830 (
		_w4975_,
		_w4976_,
		_w4977_
	);
	LUT4 #(
		.INIT('hcc4c)
	) name2831 (
		\u12_o6_we_reg/P0001 ,
		\u5_mem_reg[1][22]/NET0131 ,
		\u5_wp_reg[0]/P0001 ,
		\u5_wp_reg[1]/NET0131 ,
		_w4978_
	);
	LUT4 #(
		.INIT('h0080)
	) name2832 (
		\u12_dout_reg[22]/P0001 ,
		\u12_o6_we_reg/P0001 ,
		\u5_wp_reg[0]/P0001 ,
		\u5_wp_reg[1]/NET0131 ,
		_w4979_
	);
	LUT2 #(
		.INIT('he)
	) name2833 (
		_w4978_,
		_w4979_,
		_w4980_
	);
	LUT4 #(
		.INIT('hcc4c)
	) name2834 (
		\u12_o6_we_reg/P0001 ,
		\u5_mem_reg[1][23]/NET0131 ,
		\u5_wp_reg[0]/P0001 ,
		\u5_wp_reg[1]/NET0131 ,
		_w4981_
	);
	LUT4 #(
		.INIT('h0080)
	) name2835 (
		\u12_dout_reg[23]/P0001 ,
		\u12_o6_we_reg/P0001 ,
		\u5_wp_reg[0]/P0001 ,
		\u5_wp_reg[1]/NET0131 ,
		_w4982_
	);
	LUT2 #(
		.INIT('he)
	) name2836 (
		_w4981_,
		_w4982_,
		_w4983_
	);
	LUT4 #(
		.INIT('hcc4c)
	) name2837 (
		\u12_o6_we_reg/P0001 ,
		\u5_mem_reg[1][24]/NET0131 ,
		\u5_wp_reg[0]/P0001 ,
		\u5_wp_reg[1]/NET0131 ,
		_w4984_
	);
	LUT4 #(
		.INIT('h0080)
	) name2838 (
		\u12_dout_reg[24]/P0001 ,
		\u12_o6_we_reg/P0001 ,
		\u5_wp_reg[0]/P0001 ,
		\u5_wp_reg[1]/NET0131 ,
		_w4985_
	);
	LUT2 #(
		.INIT('he)
	) name2839 (
		_w4984_,
		_w4985_,
		_w4986_
	);
	LUT4 #(
		.INIT('hcc4c)
	) name2840 (
		\u12_o6_we_reg/P0001 ,
		\u5_mem_reg[1][25]/NET0131 ,
		\u5_wp_reg[0]/P0001 ,
		\u5_wp_reg[1]/NET0131 ,
		_w4987_
	);
	LUT4 #(
		.INIT('h0080)
	) name2841 (
		\u12_dout_reg[25]/P0001 ,
		\u12_o6_we_reg/P0001 ,
		\u5_wp_reg[0]/P0001 ,
		\u5_wp_reg[1]/NET0131 ,
		_w4988_
	);
	LUT2 #(
		.INIT('he)
	) name2842 (
		_w4987_,
		_w4988_,
		_w4989_
	);
	LUT4 #(
		.INIT('hcc4c)
	) name2843 (
		\u12_o6_we_reg/P0001 ,
		\u5_mem_reg[1][26]/NET0131 ,
		\u5_wp_reg[0]/P0001 ,
		\u5_wp_reg[1]/NET0131 ,
		_w4990_
	);
	LUT4 #(
		.INIT('h0080)
	) name2844 (
		\u12_dout_reg[26]/P0001 ,
		\u12_o6_we_reg/P0001 ,
		\u5_wp_reg[0]/P0001 ,
		\u5_wp_reg[1]/NET0131 ,
		_w4991_
	);
	LUT2 #(
		.INIT('he)
	) name2845 (
		_w4990_,
		_w4991_,
		_w4992_
	);
	LUT4 #(
		.INIT('hcc4c)
	) name2846 (
		\u12_o6_we_reg/P0001 ,
		\u5_mem_reg[1][27]/NET0131 ,
		\u5_wp_reg[0]/P0001 ,
		\u5_wp_reg[1]/NET0131 ,
		_w4993_
	);
	LUT4 #(
		.INIT('h0080)
	) name2847 (
		\u12_dout_reg[27]/P0001 ,
		\u12_o6_we_reg/P0001 ,
		\u5_wp_reg[0]/P0001 ,
		\u5_wp_reg[1]/NET0131 ,
		_w4994_
	);
	LUT2 #(
		.INIT('he)
	) name2848 (
		_w4993_,
		_w4994_,
		_w4995_
	);
	LUT4 #(
		.INIT('hcc4c)
	) name2849 (
		\u12_o6_we_reg/P0001 ,
		\u5_mem_reg[1][28]/NET0131 ,
		\u5_wp_reg[0]/P0001 ,
		\u5_wp_reg[1]/NET0131 ,
		_w4996_
	);
	LUT4 #(
		.INIT('h0080)
	) name2850 (
		\u12_dout_reg[28]/P0001 ,
		\u12_o6_we_reg/P0001 ,
		\u5_wp_reg[0]/P0001 ,
		\u5_wp_reg[1]/NET0131 ,
		_w4997_
	);
	LUT2 #(
		.INIT('he)
	) name2851 (
		_w4996_,
		_w4997_,
		_w4998_
	);
	LUT4 #(
		.INIT('hcc4c)
	) name2852 (
		\u12_o6_we_reg/P0001 ,
		\u5_mem_reg[1][29]/NET0131 ,
		\u5_wp_reg[0]/P0001 ,
		\u5_wp_reg[1]/NET0131 ,
		_w4999_
	);
	LUT4 #(
		.INIT('h0080)
	) name2853 (
		\u12_dout_reg[29]/P0001 ,
		\u12_o6_we_reg/P0001 ,
		\u5_wp_reg[0]/P0001 ,
		\u5_wp_reg[1]/NET0131 ,
		_w5000_
	);
	LUT2 #(
		.INIT('he)
	) name2854 (
		_w4999_,
		_w5000_,
		_w5001_
	);
	LUT4 #(
		.INIT('hcc4c)
	) name2855 (
		\u12_o6_we_reg/P0001 ,
		\u5_mem_reg[1][2]/NET0131 ,
		\u5_wp_reg[0]/P0001 ,
		\u5_wp_reg[1]/NET0131 ,
		_w5002_
	);
	LUT4 #(
		.INIT('h0080)
	) name2856 (
		\u12_dout_reg[2]/P0001 ,
		\u12_o6_we_reg/P0001 ,
		\u5_wp_reg[0]/P0001 ,
		\u5_wp_reg[1]/NET0131 ,
		_w5003_
	);
	LUT2 #(
		.INIT('he)
	) name2857 (
		_w5002_,
		_w5003_,
		_w5004_
	);
	LUT4 #(
		.INIT('hcc4c)
	) name2858 (
		\u12_o6_we_reg/P0001 ,
		\u5_mem_reg[1][30]/NET0131 ,
		\u5_wp_reg[0]/P0001 ,
		\u5_wp_reg[1]/NET0131 ,
		_w5005_
	);
	LUT4 #(
		.INIT('h0080)
	) name2859 (
		\u12_dout_reg[30]/P0001 ,
		\u12_o6_we_reg/P0001 ,
		\u5_wp_reg[0]/P0001 ,
		\u5_wp_reg[1]/NET0131 ,
		_w5006_
	);
	LUT2 #(
		.INIT('he)
	) name2860 (
		_w5005_,
		_w5006_,
		_w5007_
	);
	LUT4 #(
		.INIT('hcc4c)
	) name2861 (
		\u12_o6_we_reg/P0001 ,
		\u5_mem_reg[1][31]/NET0131 ,
		\u5_wp_reg[0]/P0001 ,
		\u5_wp_reg[1]/NET0131 ,
		_w5008_
	);
	LUT4 #(
		.INIT('h0080)
	) name2862 (
		\u12_dout_reg[31]/P0001 ,
		\u12_o6_we_reg/P0001 ,
		\u5_wp_reg[0]/P0001 ,
		\u5_wp_reg[1]/NET0131 ,
		_w5009_
	);
	LUT2 #(
		.INIT('he)
	) name2863 (
		_w5008_,
		_w5009_,
		_w5010_
	);
	LUT4 #(
		.INIT('hcc4c)
	) name2864 (
		\u12_o6_we_reg/P0001 ,
		\u5_mem_reg[1][3]/NET0131 ,
		\u5_wp_reg[0]/P0001 ,
		\u5_wp_reg[1]/NET0131 ,
		_w5011_
	);
	LUT4 #(
		.INIT('h0080)
	) name2865 (
		\u12_dout_reg[3]/P0001 ,
		\u12_o6_we_reg/P0001 ,
		\u5_wp_reg[0]/P0001 ,
		\u5_wp_reg[1]/NET0131 ,
		_w5012_
	);
	LUT2 #(
		.INIT('he)
	) name2866 (
		_w5011_,
		_w5012_,
		_w5013_
	);
	LUT4 #(
		.INIT('hcc4c)
	) name2867 (
		\u12_o6_we_reg/P0001 ,
		\u5_mem_reg[1][4]/NET0131 ,
		\u5_wp_reg[0]/P0001 ,
		\u5_wp_reg[1]/NET0131 ,
		_w5014_
	);
	LUT4 #(
		.INIT('h0080)
	) name2868 (
		\u12_dout_reg[4]/P0001 ,
		\u12_o6_we_reg/P0001 ,
		\u5_wp_reg[0]/P0001 ,
		\u5_wp_reg[1]/NET0131 ,
		_w5015_
	);
	LUT2 #(
		.INIT('he)
	) name2869 (
		_w5014_,
		_w5015_,
		_w5016_
	);
	LUT4 #(
		.INIT('hcc4c)
	) name2870 (
		\u12_o6_we_reg/P0001 ,
		\u5_mem_reg[1][5]/NET0131 ,
		\u5_wp_reg[0]/P0001 ,
		\u5_wp_reg[1]/NET0131 ,
		_w5017_
	);
	LUT4 #(
		.INIT('h0080)
	) name2871 (
		\u12_dout_reg[5]/P0001 ,
		\u12_o6_we_reg/P0001 ,
		\u5_wp_reg[0]/P0001 ,
		\u5_wp_reg[1]/NET0131 ,
		_w5018_
	);
	LUT2 #(
		.INIT('he)
	) name2872 (
		_w5017_,
		_w5018_,
		_w5019_
	);
	LUT4 #(
		.INIT('hcc4c)
	) name2873 (
		\u12_o6_we_reg/P0001 ,
		\u5_mem_reg[1][6]/NET0131 ,
		\u5_wp_reg[0]/P0001 ,
		\u5_wp_reg[1]/NET0131 ,
		_w5020_
	);
	LUT4 #(
		.INIT('h0080)
	) name2874 (
		\u12_dout_reg[6]/P0001 ,
		\u12_o6_we_reg/P0001 ,
		\u5_wp_reg[0]/P0001 ,
		\u5_wp_reg[1]/NET0131 ,
		_w5021_
	);
	LUT2 #(
		.INIT('he)
	) name2875 (
		_w5020_,
		_w5021_,
		_w5022_
	);
	LUT4 #(
		.INIT('hcc4c)
	) name2876 (
		\u12_o6_we_reg/P0001 ,
		\u5_mem_reg[1][7]/NET0131 ,
		\u5_wp_reg[0]/P0001 ,
		\u5_wp_reg[1]/NET0131 ,
		_w5023_
	);
	LUT4 #(
		.INIT('h0080)
	) name2877 (
		\u12_dout_reg[7]/P0001 ,
		\u12_o6_we_reg/P0001 ,
		\u5_wp_reg[0]/P0001 ,
		\u5_wp_reg[1]/NET0131 ,
		_w5024_
	);
	LUT2 #(
		.INIT('he)
	) name2878 (
		_w5023_,
		_w5024_,
		_w5025_
	);
	LUT4 #(
		.INIT('hcc4c)
	) name2879 (
		\u12_o6_we_reg/P0001 ,
		\u5_mem_reg[1][8]/NET0131 ,
		\u5_wp_reg[0]/P0001 ,
		\u5_wp_reg[1]/NET0131 ,
		_w5026_
	);
	LUT4 #(
		.INIT('h0080)
	) name2880 (
		\u12_dout_reg[8]/P0001 ,
		\u12_o6_we_reg/P0001 ,
		\u5_wp_reg[0]/P0001 ,
		\u5_wp_reg[1]/NET0131 ,
		_w5027_
	);
	LUT2 #(
		.INIT('he)
	) name2881 (
		_w5026_,
		_w5027_,
		_w5028_
	);
	LUT4 #(
		.INIT('hcc4c)
	) name2882 (
		\u12_o6_we_reg/P0001 ,
		\u5_mem_reg[1][9]/NET0131 ,
		\u5_wp_reg[0]/P0001 ,
		\u5_wp_reg[1]/NET0131 ,
		_w5029_
	);
	LUT4 #(
		.INIT('h0080)
	) name2883 (
		\u12_dout_reg[9]/P0001 ,
		\u12_o6_we_reg/P0001 ,
		\u5_wp_reg[0]/P0001 ,
		\u5_wp_reg[1]/NET0131 ,
		_w5030_
	);
	LUT2 #(
		.INIT('he)
	) name2884 (
		_w5029_,
		_w5030_,
		_w5031_
	);
	LUT4 #(
		.INIT('hc4cc)
	) name2885 (
		\u12_o6_we_reg/P0001 ,
		\u5_mem_reg[2][0]/NET0131 ,
		\u5_wp_reg[0]/P0001 ,
		\u5_wp_reg[1]/NET0131 ,
		_w5032_
	);
	LUT4 #(
		.INIT('h0800)
	) name2886 (
		\u12_dout_reg[0]/P0001 ,
		\u12_o6_we_reg/P0001 ,
		\u5_wp_reg[0]/P0001 ,
		\u5_wp_reg[1]/NET0131 ,
		_w5033_
	);
	LUT2 #(
		.INIT('he)
	) name2887 (
		_w5032_,
		_w5033_,
		_w5034_
	);
	LUT4 #(
		.INIT('hc4cc)
	) name2888 (
		\u12_o6_we_reg/P0001 ,
		\u5_mem_reg[2][10]/NET0131 ,
		\u5_wp_reg[0]/P0001 ,
		\u5_wp_reg[1]/NET0131 ,
		_w5035_
	);
	LUT4 #(
		.INIT('h0800)
	) name2889 (
		\u12_dout_reg[10]/P0001 ,
		\u12_o6_we_reg/P0001 ,
		\u5_wp_reg[0]/P0001 ,
		\u5_wp_reg[1]/NET0131 ,
		_w5036_
	);
	LUT2 #(
		.INIT('he)
	) name2890 (
		_w5035_,
		_w5036_,
		_w5037_
	);
	LUT4 #(
		.INIT('hc4cc)
	) name2891 (
		\u12_o6_we_reg/P0001 ,
		\u5_mem_reg[2][11]/NET0131 ,
		\u5_wp_reg[0]/P0001 ,
		\u5_wp_reg[1]/NET0131 ,
		_w5038_
	);
	LUT4 #(
		.INIT('h0800)
	) name2892 (
		\u12_dout_reg[11]/P0001 ,
		\u12_o6_we_reg/P0001 ,
		\u5_wp_reg[0]/P0001 ,
		\u5_wp_reg[1]/NET0131 ,
		_w5039_
	);
	LUT2 #(
		.INIT('he)
	) name2893 (
		_w5038_,
		_w5039_,
		_w5040_
	);
	LUT4 #(
		.INIT('hc4cc)
	) name2894 (
		\u12_o6_we_reg/P0001 ,
		\u5_mem_reg[2][12]/NET0131 ,
		\u5_wp_reg[0]/P0001 ,
		\u5_wp_reg[1]/NET0131 ,
		_w5041_
	);
	LUT4 #(
		.INIT('h0800)
	) name2895 (
		\u12_dout_reg[12]/P0001 ,
		\u12_o6_we_reg/P0001 ,
		\u5_wp_reg[0]/P0001 ,
		\u5_wp_reg[1]/NET0131 ,
		_w5042_
	);
	LUT2 #(
		.INIT('he)
	) name2896 (
		_w5041_,
		_w5042_,
		_w5043_
	);
	LUT4 #(
		.INIT('hc4cc)
	) name2897 (
		\u12_o6_we_reg/P0001 ,
		\u5_mem_reg[2][13]/NET0131 ,
		\u5_wp_reg[0]/P0001 ,
		\u5_wp_reg[1]/NET0131 ,
		_w5044_
	);
	LUT4 #(
		.INIT('h0800)
	) name2898 (
		\u12_dout_reg[13]/P0001 ,
		\u12_o6_we_reg/P0001 ,
		\u5_wp_reg[0]/P0001 ,
		\u5_wp_reg[1]/NET0131 ,
		_w5045_
	);
	LUT2 #(
		.INIT('he)
	) name2899 (
		_w5044_,
		_w5045_,
		_w5046_
	);
	LUT4 #(
		.INIT('hc4cc)
	) name2900 (
		\u12_o6_we_reg/P0001 ,
		\u5_mem_reg[2][14]/NET0131 ,
		\u5_wp_reg[0]/P0001 ,
		\u5_wp_reg[1]/NET0131 ,
		_w5047_
	);
	LUT4 #(
		.INIT('h0800)
	) name2901 (
		\u12_dout_reg[14]/P0001 ,
		\u12_o6_we_reg/P0001 ,
		\u5_wp_reg[0]/P0001 ,
		\u5_wp_reg[1]/NET0131 ,
		_w5048_
	);
	LUT2 #(
		.INIT('he)
	) name2902 (
		_w5047_,
		_w5048_,
		_w5049_
	);
	LUT4 #(
		.INIT('hc4cc)
	) name2903 (
		\u12_o6_we_reg/P0001 ,
		\u5_mem_reg[2][15]/NET0131 ,
		\u5_wp_reg[0]/P0001 ,
		\u5_wp_reg[1]/NET0131 ,
		_w5050_
	);
	LUT4 #(
		.INIT('h0800)
	) name2904 (
		\u12_dout_reg[15]/P0001 ,
		\u12_o6_we_reg/P0001 ,
		\u5_wp_reg[0]/P0001 ,
		\u5_wp_reg[1]/NET0131 ,
		_w5051_
	);
	LUT2 #(
		.INIT('he)
	) name2905 (
		_w5050_,
		_w5051_,
		_w5052_
	);
	LUT4 #(
		.INIT('hc4cc)
	) name2906 (
		\u12_o6_we_reg/P0001 ,
		\u5_mem_reg[2][16]/NET0131 ,
		\u5_wp_reg[0]/P0001 ,
		\u5_wp_reg[1]/NET0131 ,
		_w5053_
	);
	LUT4 #(
		.INIT('h0800)
	) name2907 (
		\u12_dout_reg[16]/P0001 ,
		\u12_o6_we_reg/P0001 ,
		\u5_wp_reg[0]/P0001 ,
		\u5_wp_reg[1]/NET0131 ,
		_w5054_
	);
	LUT2 #(
		.INIT('he)
	) name2908 (
		_w5053_,
		_w5054_,
		_w5055_
	);
	LUT4 #(
		.INIT('hc4cc)
	) name2909 (
		\u12_o6_we_reg/P0001 ,
		\u5_mem_reg[2][17]/NET0131 ,
		\u5_wp_reg[0]/P0001 ,
		\u5_wp_reg[1]/NET0131 ,
		_w5056_
	);
	LUT4 #(
		.INIT('h0800)
	) name2910 (
		\u12_dout_reg[17]/P0001 ,
		\u12_o6_we_reg/P0001 ,
		\u5_wp_reg[0]/P0001 ,
		\u5_wp_reg[1]/NET0131 ,
		_w5057_
	);
	LUT2 #(
		.INIT('he)
	) name2911 (
		_w5056_,
		_w5057_,
		_w5058_
	);
	LUT4 #(
		.INIT('hc4cc)
	) name2912 (
		\u12_o6_we_reg/P0001 ,
		\u5_mem_reg[2][18]/NET0131 ,
		\u5_wp_reg[0]/P0001 ,
		\u5_wp_reg[1]/NET0131 ,
		_w5059_
	);
	LUT4 #(
		.INIT('h0800)
	) name2913 (
		\u12_dout_reg[18]/P0001 ,
		\u12_o6_we_reg/P0001 ,
		\u5_wp_reg[0]/P0001 ,
		\u5_wp_reg[1]/NET0131 ,
		_w5060_
	);
	LUT2 #(
		.INIT('he)
	) name2914 (
		_w5059_,
		_w5060_,
		_w5061_
	);
	LUT4 #(
		.INIT('hc4cc)
	) name2915 (
		\u12_o6_we_reg/P0001 ,
		\u5_mem_reg[2][19]/NET0131 ,
		\u5_wp_reg[0]/P0001 ,
		\u5_wp_reg[1]/NET0131 ,
		_w5062_
	);
	LUT4 #(
		.INIT('h0800)
	) name2916 (
		\u12_dout_reg[19]/P0001 ,
		\u12_o6_we_reg/P0001 ,
		\u5_wp_reg[0]/P0001 ,
		\u5_wp_reg[1]/NET0131 ,
		_w5063_
	);
	LUT2 #(
		.INIT('he)
	) name2917 (
		_w5062_,
		_w5063_,
		_w5064_
	);
	LUT4 #(
		.INIT('hc4cc)
	) name2918 (
		\u12_o6_we_reg/P0001 ,
		\u5_mem_reg[2][1]/NET0131 ,
		\u5_wp_reg[0]/P0001 ,
		\u5_wp_reg[1]/NET0131 ,
		_w5065_
	);
	LUT4 #(
		.INIT('h0800)
	) name2919 (
		\u12_dout_reg[1]/P0001 ,
		\u12_o6_we_reg/P0001 ,
		\u5_wp_reg[0]/P0001 ,
		\u5_wp_reg[1]/NET0131 ,
		_w5066_
	);
	LUT2 #(
		.INIT('he)
	) name2920 (
		_w5065_,
		_w5066_,
		_w5067_
	);
	LUT4 #(
		.INIT('hc4cc)
	) name2921 (
		\u12_o6_we_reg/P0001 ,
		\u5_mem_reg[2][20]/NET0131 ,
		\u5_wp_reg[0]/P0001 ,
		\u5_wp_reg[1]/NET0131 ,
		_w5068_
	);
	LUT4 #(
		.INIT('h0800)
	) name2922 (
		\u12_dout_reg[20]/P0001 ,
		\u12_o6_we_reg/P0001 ,
		\u5_wp_reg[0]/P0001 ,
		\u5_wp_reg[1]/NET0131 ,
		_w5069_
	);
	LUT2 #(
		.INIT('he)
	) name2923 (
		_w5068_,
		_w5069_,
		_w5070_
	);
	LUT4 #(
		.INIT('hc4cc)
	) name2924 (
		\u12_o6_we_reg/P0001 ,
		\u5_mem_reg[2][21]/NET0131 ,
		\u5_wp_reg[0]/P0001 ,
		\u5_wp_reg[1]/NET0131 ,
		_w5071_
	);
	LUT4 #(
		.INIT('h0800)
	) name2925 (
		\u12_dout_reg[21]/P0001 ,
		\u12_o6_we_reg/P0001 ,
		\u5_wp_reg[0]/P0001 ,
		\u5_wp_reg[1]/NET0131 ,
		_w5072_
	);
	LUT2 #(
		.INIT('he)
	) name2926 (
		_w5071_,
		_w5072_,
		_w5073_
	);
	LUT4 #(
		.INIT('hc4cc)
	) name2927 (
		\u12_o6_we_reg/P0001 ,
		\u5_mem_reg[2][22]/NET0131 ,
		\u5_wp_reg[0]/P0001 ,
		\u5_wp_reg[1]/NET0131 ,
		_w5074_
	);
	LUT4 #(
		.INIT('h0800)
	) name2928 (
		\u12_dout_reg[22]/P0001 ,
		\u12_o6_we_reg/P0001 ,
		\u5_wp_reg[0]/P0001 ,
		\u5_wp_reg[1]/NET0131 ,
		_w5075_
	);
	LUT2 #(
		.INIT('he)
	) name2929 (
		_w5074_,
		_w5075_,
		_w5076_
	);
	LUT4 #(
		.INIT('hc4cc)
	) name2930 (
		\u12_o6_we_reg/P0001 ,
		\u5_mem_reg[2][23]/NET0131 ,
		\u5_wp_reg[0]/P0001 ,
		\u5_wp_reg[1]/NET0131 ,
		_w5077_
	);
	LUT4 #(
		.INIT('h0800)
	) name2931 (
		\u12_dout_reg[23]/P0001 ,
		\u12_o6_we_reg/P0001 ,
		\u5_wp_reg[0]/P0001 ,
		\u5_wp_reg[1]/NET0131 ,
		_w5078_
	);
	LUT2 #(
		.INIT('he)
	) name2932 (
		_w5077_,
		_w5078_,
		_w5079_
	);
	LUT4 #(
		.INIT('hc4cc)
	) name2933 (
		\u12_o6_we_reg/P0001 ,
		\u5_mem_reg[2][24]/NET0131 ,
		\u5_wp_reg[0]/P0001 ,
		\u5_wp_reg[1]/NET0131 ,
		_w5080_
	);
	LUT4 #(
		.INIT('h0800)
	) name2934 (
		\u12_dout_reg[24]/P0001 ,
		\u12_o6_we_reg/P0001 ,
		\u5_wp_reg[0]/P0001 ,
		\u5_wp_reg[1]/NET0131 ,
		_w5081_
	);
	LUT2 #(
		.INIT('he)
	) name2935 (
		_w5080_,
		_w5081_,
		_w5082_
	);
	LUT4 #(
		.INIT('hc4cc)
	) name2936 (
		\u12_o6_we_reg/P0001 ,
		\u5_mem_reg[2][25]/NET0131 ,
		\u5_wp_reg[0]/P0001 ,
		\u5_wp_reg[1]/NET0131 ,
		_w5083_
	);
	LUT4 #(
		.INIT('h0800)
	) name2937 (
		\u12_dout_reg[25]/P0001 ,
		\u12_o6_we_reg/P0001 ,
		\u5_wp_reg[0]/P0001 ,
		\u5_wp_reg[1]/NET0131 ,
		_w5084_
	);
	LUT2 #(
		.INIT('he)
	) name2938 (
		_w5083_,
		_w5084_,
		_w5085_
	);
	LUT4 #(
		.INIT('hc4cc)
	) name2939 (
		\u12_o6_we_reg/P0001 ,
		\u5_mem_reg[2][26]/NET0131 ,
		\u5_wp_reg[0]/P0001 ,
		\u5_wp_reg[1]/NET0131 ,
		_w5086_
	);
	LUT4 #(
		.INIT('h0800)
	) name2940 (
		\u12_dout_reg[26]/P0001 ,
		\u12_o6_we_reg/P0001 ,
		\u5_wp_reg[0]/P0001 ,
		\u5_wp_reg[1]/NET0131 ,
		_w5087_
	);
	LUT2 #(
		.INIT('he)
	) name2941 (
		_w5086_,
		_w5087_,
		_w5088_
	);
	LUT4 #(
		.INIT('hc4cc)
	) name2942 (
		\u12_o6_we_reg/P0001 ,
		\u5_mem_reg[2][27]/NET0131 ,
		\u5_wp_reg[0]/P0001 ,
		\u5_wp_reg[1]/NET0131 ,
		_w5089_
	);
	LUT4 #(
		.INIT('h0800)
	) name2943 (
		\u12_dout_reg[27]/P0001 ,
		\u12_o6_we_reg/P0001 ,
		\u5_wp_reg[0]/P0001 ,
		\u5_wp_reg[1]/NET0131 ,
		_w5090_
	);
	LUT2 #(
		.INIT('he)
	) name2944 (
		_w5089_,
		_w5090_,
		_w5091_
	);
	LUT4 #(
		.INIT('hc4cc)
	) name2945 (
		\u12_o6_we_reg/P0001 ,
		\u5_mem_reg[2][28]/NET0131 ,
		\u5_wp_reg[0]/P0001 ,
		\u5_wp_reg[1]/NET0131 ,
		_w5092_
	);
	LUT4 #(
		.INIT('h0800)
	) name2946 (
		\u12_dout_reg[28]/P0001 ,
		\u12_o6_we_reg/P0001 ,
		\u5_wp_reg[0]/P0001 ,
		\u5_wp_reg[1]/NET0131 ,
		_w5093_
	);
	LUT2 #(
		.INIT('he)
	) name2947 (
		_w5092_,
		_w5093_,
		_w5094_
	);
	LUT4 #(
		.INIT('hc4cc)
	) name2948 (
		\u12_o6_we_reg/P0001 ,
		\u5_mem_reg[2][29]/NET0131 ,
		\u5_wp_reg[0]/P0001 ,
		\u5_wp_reg[1]/NET0131 ,
		_w5095_
	);
	LUT4 #(
		.INIT('h0800)
	) name2949 (
		\u12_dout_reg[29]/P0001 ,
		\u12_o6_we_reg/P0001 ,
		\u5_wp_reg[0]/P0001 ,
		\u5_wp_reg[1]/NET0131 ,
		_w5096_
	);
	LUT2 #(
		.INIT('he)
	) name2950 (
		_w5095_,
		_w5096_,
		_w5097_
	);
	LUT4 #(
		.INIT('hc4cc)
	) name2951 (
		\u12_o6_we_reg/P0001 ,
		\u5_mem_reg[2][2]/NET0131 ,
		\u5_wp_reg[0]/P0001 ,
		\u5_wp_reg[1]/NET0131 ,
		_w5098_
	);
	LUT4 #(
		.INIT('h0800)
	) name2952 (
		\u12_dout_reg[2]/P0001 ,
		\u12_o6_we_reg/P0001 ,
		\u5_wp_reg[0]/P0001 ,
		\u5_wp_reg[1]/NET0131 ,
		_w5099_
	);
	LUT2 #(
		.INIT('he)
	) name2953 (
		_w5098_,
		_w5099_,
		_w5100_
	);
	LUT4 #(
		.INIT('hc4cc)
	) name2954 (
		\u12_o6_we_reg/P0001 ,
		\u5_mem_reg[2][30]/NET0131 ,
		\u5_wp_reg[0]/P0001 ,
		\u5_wp_reg[1]/NET0131 ,
		_w5101_
	);
	LUT4 #(
		.INIT('h0800)
	) name2955 (
		\u12_dout_reg[30]/P0001 ,
		\u12_o6_we_reg/P0001 ,
		\u5_wp_reg[0]/P0001 ,
		\u5_wp_reg[1]/NET0131 ,
		_w5102_
	);
	LUT2 #(
		.INIT('he)
	) name2956 (
		_w5101_,
		_w5102_,
		_w5103_
	);
	LUT4 #(
		.INIT('hc4cc)
	) name2957 (
		\u12_o6_we_reg/P0001 ,
		\u5_mem_reg[2][31]/NET0131 ,
		\u5_wp_reg[0]/P0001 ,
		\u5_wp_reg[1]/NET0131 ,
		_w5104_
	);
	LUT4 #(
		.INIT('h0800)
	) name2958 (
		\u12_dout_reg[31]/P0001 ,
		\u12_o6_we_reg/P0001 ,
		\u5_wp_reg[0]/P0001 ,
		\u5_wp_reg[1]/NET0131 ,
		_w5105_
	);
	LUT2 #(
		.INIT('he)
	) name2959 (
		_w5104_,
		_w5105_,
		_w5106_
	);
	LUT4 #(
		.INIT('hc4cc)
	) name2960 (
		\u12_o6_we_reg/P0001 ,
		\u5_mem_reg[2][3]/NET0131 ,
		\u5_wp_reg[0]/P0001 ,
		\u5_wp_reg[1]/NET0131 ,
		_w5107_
	);
	LUT4 #(
		.INIT('h0800)
	) name2961 (
		\u12_dout_reg[3]/P0001 ,
		\u12_o6_we_reg/P0001 ,
		\u5_wp_reg[0]/P0001 ,
		\u5_wp_reg[1]/NET0131 ,
		_w5108_
	);
	LUT2 #(
		.INIT('he)
	) name2962 (
		_w5107_,
		_w5108_,
		_w5109_
	);
	LUT4 #(
		.INIT('hc4cc)
	) name2963 (
		\u12_o6_we_reg/P0001 ,
		\u5_mem_reg[2][4]/NET0131 ,
		\u5_wp_reg[0]/P0001 ,
		\u5_wp_reg[1]/NET0131 ,
		_w5110_
	);
	LUT4 #(
		.INIT('h0800)
	) name2964 (
		\u12_dout_reg[4]/P0001 ,
		\u12_o6_we_reg/P0001 ,
		\u5_wp_reg[0]/P0001 ,
		\u5_wp_reg[1]/NET0131 ,
		_w5111_
	);
	LUT2 #(
		.INIT('he)
	) name2965 (
		_w5110_,
		_w5111_,
		_w5112_
	);
	LUT4 #(
		.INIT('hc4cc)
	) name2966 (
		\u12_o6_we_reg/P0001 ,
		\u5_mem_reg[2][5]/NET0131 ,
		\u5_wp_reg[0]/P0001 ,
		\u5_wp_reg[1]/NET0131 ,
		_w5113_
	);
	LUT4 #(
		.INIT('h0800)
	) name2967 (
		\u12_dout_reg[5]/P0001 ,
		\u12_o6_we_reg/P0001 ,
		\u5_wp_reg[0]/P0001 ,
		\u5_wp_reg[1]/NET0131 ,
		_w5114_
	);
	LUT2 #(
		.INIT('he)
	) name2968 (
		_w5113_,
		_w5114_,
		_w5115_
	);
	LUT4 #(
		.INIT('hc4cc)
	) name2969 (
		\u12_o6_we_reg/P0001 ,
		\u5_mem_reg[2][6]/NET0131 ,
		\u5_wp_reg[0]/P0001 ,
		\u5_wp_reg[1]/NET0131 ,
		_w5116_
	);
	LUT4 #(
		.INIT('h0800)
	) name2970 (
		\u12_dout_reg[6]/P0001 ,
		\u12_o6_we_reg/P0001 ,
		\u5_wp_reg[0]/P0001 ,
		\u5_wp_reg[1]/NET0131 ,
		_w5117_
	);
	LUT2 #(
		.INIT('he)
	) name2971 (
		_w5116_,
		_w5117_,
		_w5118_
	);
	LUT4 #(
		.INIT('hc4cc)
	) name2972 (
		\u12_o6_we_reg/P0001 ,
		\u5_mem_reg[2][7]/NET0131 ,
		\u5_wp_reg[0]/P0001 ,
		\u5_wp_reg[1]/NET0131 ,
		_w5119_
	);
	LUT4 #(
		.INIT('h0800)
	) name2973 (
		\u12_dout_reg[7]/P0001 ,
		\u12_o6_we_reg/P0001 ,
		\u5_wp_reg[0]/P0001 ,
		\u5_wp_reg[1]/NET0131 ,
		_w5120_
	);
	LUT2 #(
		.INIT('he)
	) name2974 (
		_w5119_,
		_w5120_,
		_w5121_
	);
	LUT4 #(
		.INIT('hc4cc)
	) name2975 (
		\u12_o6_we_reg/P0001 ,
		\u5_mem_reg[2][8]/NET0131 ,
		\u5_wp_reg[0]/P0001 ,
		\u5_wp_reg[1]/NET0131 ,
		_w5122_
	);
	LUT4 #(
		.INIT('h0800)
	) name2976 (
		\u12_dout_reg[8]/P0001 ,
		\u12_o6_we_reg/P0001 ,
		\u5_wp_reg[0]/P0001 ,
		\u5_wp_reg[1]/NET0131 ,
		_w5123_
	);
	LUT2 #(
		.INIT('he)
	) name2977 (
		_w5122_,
		_w5123_,
		_w5124_
	);
	LUT4 #(
		.INIT('hc4cc)
	) name2978 (
		\u12_o6_we_reg/P0001 ,
		\u5_mem_reg[2][9]/NET0131 ,
		\u5_wp_reg[0]/P0001 ,
		\u5_wp_reg[1]/NET0131 ,
		_w5125_
	);
	LUT4 #(
		.INIT('h0800)
	) name2979 (
		\u12_dout_reg[9]/P0001 ,
		\u12_o6_we_reg/P0001 ,
		\u5_wp_reg[0]/P0001 ,
		\u5_wp_reg[1]/NET0131 ,
		_w5126_
	);
	LUT2 #(
		.INIT('he)
	) name2980 (
		_w5125_,
		_w5126_,
		_w5127_
	);
	LUT4 #(
		.INIT('h4ccc)
	) name2981 (
		\u12_o6_we_reg/P0001 ,
		\u5_mem_reg[3][0]/NET0131 ,
		\u5_wp_reg[0]/P0001 ,
		\u5_wp_reg[1]/NET0131 ,
		_w5128_
	);
	LUT4 #(
		.INIT('h8000)
	) name2982 (
		\u12_dout_reg[0]/P0001 ,
		\u12_o6_we_reg/P0001 ,
		\u5_wp_reg[0]/P0001 ,
		\u5_wp_reg[1]/NET0131 ,
		_w5129_
	);
	LUT2 #(
		.INIT('he)
	) name2983 (
		_w5128_,
		_w5129_,
		_w5130_
	);
	LUT4 #(
		.INIT('h4ccc)
	) name2984 (
		\u12_o6_we_reg/P0001 ,
		\u5_mem_reg[3][10]/NET0131 ,
		\u5_wp_reg[0]/P0001 ,
		\u5_wp_reg[1]/NET0131 ,
		_w5131_
	);
	LUT4 #(
		.INIT('h8000)
	) name2985 (
		\u12_dout_reg[10]/P0001 ,
		\u12_o6_we_reg/P0001 ,
		\u5_wp_reg[0]/P0001 ,
		\u5_wp_reg[1]/NET0131 ,
		_w5132_
	);
	LUT2 #(
		.INIT('he)
	) name2986 (
		_w5131_,
		_w5132_,
		_w5133_
	);
	LUT4 #(
		.INIT('h4ccc)
	) name2987 (
		\u12_o6_we_reg/P0001 ,
		\u5_mem_reg[3][11]/NET0131 ,
		\u5_wp_reg[0]/P0001 ,
		\u5_wp_reg[1]/NET0131 ,
		_w5134_
	);
	LUT4 #(
		.INIT('h8000)
	) name2988 (
		\u12_dout_reg[11]/P0001 ,
		\u12_o6_we_reg/P0001 ,
		\u5_wp_reg[0]/P0001 ,
		\u5_wp_reg[1]/NET0131 ,
		_w5135_
	);
	LUT2 #(
		.INIT('he)
	) name2989 (
		_w5134_,
		_w5135_,
		_w5136_
	);
	LUT4 #(
		.INIT('h4ccc)
	) name2990 (
		\u12_o6_we_reg/P0001 ,
		\u5_mem_reg[3][12]/NET0131 ,
		\u5_wp_reg[0]/P0001 ,
		\u5_wp_reg[1]/NET0131 ,
		_w5137_
	);
	LUT4 #(
		.INIT('h8000)
	) name2991 (
		\u12_dout_reg[12]/P0001 ,
		\u12_o6_we_reg/P0001 ,
		\u5_wp_reg[0]/P0001 ,
		\u5_wp_reg[1]/NET0131 ,
		_w5138_
	);
	LUT2 #(
		.INIT('he)
	) name2992 (
		_w5137_,
		_w5138_,
		_w5139_
	);
	LUT4 #(
		.INIT('h4ccc)
	) name2993 (
		\u12_o6_we_reg/P0001 ,
		\u5_mem_reg[3][13]/NET0131 ,
		\u5_wp_reg[0]/P0001 ,
		\u5_wp_reg[1]/NET0131 ,
		_w5140_
	);
	LUT4 #(
		.INIT('h8000)
	) name2994 (
		\u12_dout_reg[13]/P0001 ,
		\u12_o6_we_reg/P0001 ,
		\u5_wp_reg[0]/P0001 ,
		\u5_wp_reg[1]/NET0131 ,
		_w5141_
	);
	LUT2 #(
		.INIT('he)
	) name2995 (
		_w5140_,
		_w5141_,
		_w5142_
	);
	LUT4 #(
		.INIT('h4ccc)
	) name2996 (
		\u12_o6_we_reg/P0001 ,
		\u5_mem_reg[3][14]/NET0131 ,
		\u5_wp_reg[0]/P0001 ,
		\u5_wp_reg[1]/NET0131 ,
		_w5143_
	);
	LUT4 #(
		.INIT('h8000)
	) name2997 (
		\u12_dout_reg[14]/P0001 ,
		\u12_o6_we_reg/P0001 ,
		\u5_wp_reg[0]/P0001 ,
		\u5_wp_reg[1]/NET0131 ,
		_w5144_
	);
	LUT2 #(
		.INIT('he)
	) name2998 (
		_w5143_,
		_w5144_,
		_w5145_
	);
	LUT4 #(
		.INIT('h4ccc)
	) name2999 (
		\u12_o6_we_reg/P0001 ,
		\u5_mem_reg[3][15]/NET0131 ,
		\u5_wp_reg[0]/P0001 ,
		\u5_wp_reg[1]/NET0131 ,
		_w5146_
	);
	LUT4 #(
		.INIT('h8000)
	) name3000 (
		\u12_dout_reg[15]/P0001 ,
		\u12_o6_we_reg/P0001 ,
		\u5_wp_reg[0]/P0001 ,
		\u5_wp_reg[1]/NET0131 ,
		_w5147_
	);
	LUT2 #(
		.INIT('he)
	) name3001 (
		_w5146_,
		_w5147_,
		_w5148_
	);
	LUT4 #(
		.INIT('h4ccc)
	) name3002 (
		\u12_o6_we_reg/P0001 ,
		\u5_mem_reg[3][16]/NET0131 ,
		\u5_wp_reg[0]/P0001 ,
		\u5_wp_reg[1]/NET0131 ,
		_w5149_
	);
	LUT4 #(
		.INIT('h8000)
	) name3003 (
		\u12_dout_reg[16]/P0001 ,
		\u12_o6_we_reg/P0001 ,
		\u5_wp_reg[0]/P0001 ,
		\u5_wp_reg[1]/NET0131 ,
		_w5150_
	);
	LUT2 #(
		.INIT('he)
	) name3004 (
		_w5149_,
		_w5150_,
		_w5151_
	);
	LUT4 #(
		.INIT('h4ccc)
	) name3005 (
		\u12_o6_we_reg/P0001 ,
		\u5_mem_reg[3][17]/NET0131 ,
		\u5_wp_reg[0]/P0001 ,
		\u5_wp_reg[1]/NET0131 ,
		_w5152_
	);
	LUT4 #(
		.INIT('h8000)
	) name3006 (
		\u12_dout_reg[17]/P0001 ,
		\u12_o6_we_reg/P0001 ,
		\u5_wp_reg[0]/P0001 ,
		\u5_wp_reg[1]/NET0131 ,
		_w5153_
	);
	LUT2 #(
		.INIT('he)
	) name3007 (
		_w5152_,
		_w5153_,
		_w5154_
	);
	LUT4 #(
		.INIT('h4ccc)
	) name3008 (
		\u12_o6_we_reg/P0001 ,
		\u5_mem_reg[3][18]/NET0131 ,
		\u5_wp_reg[0]/P0001 ,
		\u5_wp_reg[1]/NET0131 ,
		_w5155_
	);
	LUT4 #(
		.INIT('h8000)
	) name3009 (
		\u12_dout_reg[18]/P0001 ,
		\u12_o6_we_reg/P0001 ,
		\u5_wp_reg[0]/P0001 ,
		\u5_wp_reg[1]/NET0131 ,
		_w5156_
	);
	LUT2 #(
		.INIT('he)
	) name3010 (
		_w5155_,
		_w5156_,
		_w5157_
	);
	LUT4 #(
		.INIT('h4ccc)
	) name3011 (
		\u12_o6_we_reg/P0001 ,
		\u5_mem_reg[3][19]/NET0131 ,
		\u5_wp_reg[0]/P0001 ,
		\u5_wp_reg[1]/NET0131 ,
		_w5158_
	);
	LUT4 #(
		.INIT('h8000)
	) name3012 (
		\u12_dout_reg[19]/P0001 ,
		\u12_o6_we_reg/P0001 ,
		\u5_wp_reg[0]/P0001 ,
		\u5_wp_reg[1]/NET0131 ,
		_w5159_
	);
	LUT2 #(
		.INIT('he)
	) name3013 (
		_w5158_,
		_w5159_,
		_w5160_
	);
	LUT4 #(
		.INIT('h4ccc)
	) name3014 (
		\u12_o6_we_reg/P0001 ,
		\u5_mem_reg[3][1]/NET0131 ,
		\u5_wp_reg[0]/P0001 ,
		\u5_wp_reg[1]/NET0131 ,
		_w5161_
	);
	LUT4 #(
		.INIT('h8000)
	) name3015 (
		\u12_dout_reg[1]/P0001 ,
		\u12_o6_we_reg/P0001 ,
		\u5_wp_reg[0]/P0001 ,
		\u5_wp_reg[1]/NET0131 ,
		_w5162_
	);
	LUT2 #(
		.INIT('he)
	) name3016 (
		_w5161_,
		_w5162_,
		_w5163_
	);
	LUT4 #(
		.INIT('h4ccc)
	) name3017 (
		\u12_o6_we_reg/P0001 ,
		\u5_mem_reg[3][20]/NET0131 ,
		\u5_wp_reg[0]/P0001 ,
		\u5_wp_reg[1]/NET0131 ,
		_w5164_
	);
	LUT4 #(
		.INIT('h8000)
	) name3018 (
		\u12_dout_reg[20]/P0001 ,
		\u12_o6_we_reg/P0001 ,
		\u5_wp_reg[0]/P0001 ,
		\u5_wp_reg[1]/NET0131 ,
		_w5165_
	);
	LUT2 #(
		.INIT('he)
	) name3019 (
		_w5164_,
		_w5165_,
		_w5166_
	);
	LUT4 #(
		.INIT('h4ccc)
	) name3020 (
		\u12_o6_we_reg/P0001 ,
		\u5_mem_reg[3][21]/NET0131 ,
		\u5_wp_reg[0]/P0001 ,
		\u5_wp_reg[1]/NET0131 ,
		_w5167_
	);
	LUT4 #(
		.INIT('h8000)
	) name3021 (
		\u12_dout_reg[21]/P0001 ,
		\u12_o6_we_reg/P0001 ,
		\u5_wp_reg[0]/P0001 ,
		\u5_wp_reg[1]/NET0131 ,
		_w5168_
	);
	LUT2 #(
		.INIT('he)
	) name3022 (
		_w5167_,
		_w5168_,
		_w5169_
	);
	LUT4 #(
		.INIT('h4ccc)
	) name3023 (
		\u12_o6_we_reg/P0001 ,
		\u5_mem_reg[3][22]/NET0131 ,
		\u5_wp_reg[0]/P0001 ,
		\u5_wp_reg[1]/NET0131 ,
		_w5170_
	);
	LUT4 #(
		.INIT('h8000)
	) name3024 (
		\u12_dout_reg[22]/P0001 ,
		\u12_o6_we_reg/P0001 ,
		\u5_wp_reg[0]/P0001 ,
		\u5_wp_reg[1]/NET0131 ,
		_w5171_
	);
	LUT2 #(
		.INIT('he)
	) name3025 (
		_w5170_,
		_w5171_,
		_w5172_
	);
	LUT4 #(
		.INIT('h4ccc)
	) name3026 (
		\u12_o6_we_reg/P0001 ,
		\u5_mem_reg[3][23]/NET0131 ,
		\u5_wp_reg[0]/P0001 ,
		\u5_wp_reg[1]/NET0131 ,
		_w5173_
	);
	LUT4 #(
		.INIT('h8000)
	) name3027 (
		\u12_dout_reg[23]/P0001 ,
		\u12_o6_we_reg/P0001 ,
		\u5_wp_reg[0]/P0001 ,
		\u5_wp_reg[1]/NET0131 ,
		_w5174_
	);
	LUT2 #(
		.INIT('he)
	) name3028 (
		_w5173_,
		_w5174_,
		_w5175_
	);
	LUT4 #(
		.INIT('h4ccc)
	) name3029 (
		\u12_o6_we_reg/P0001 ,
		\u5_mem_reg[3][24]/NET0131 ,
		\u5_wp_reg[0]/P0001 ,
		\u5_wp_reg[1]/NET0131 ,
		_w5176_
	);
	LUT4 #(
		.INIT('h8000)
	) name3030 (
		\u12_dout_reg[24]/P0001 ,
		\u12_o6_we_reg/P0001 ,
		\u5_wp_reg[0]/P0001 ,
		\u5_wp_reg[1]/NET0131 ,
		_w5177_
	);
	LUT2 #(
		.INIT('he)
	) name3031 (
		_w5176_,
		_w5177_,
		_w5178_
	);
	LUT4 #(
		.INIT('h4ccc)
	) name3032 (
		\u12_o6_we_reg/P0001 ,
		\u5_mem_reg[3][25]/NET0131 ,
		\u5_wp_reg[0]/P0001 ,
		\u5_wp_reg[1]/NET0131 ,
		_w5179_
	);
	LUT4 #(
		.INIT('h8000)
	) name3033 (
		\u12_dout_reg[25]/P0001 ,
		\u12_o6_we_reg/P0001 ,
		\u5_wp_reg[0]/P0001 ,
		\u5_wp_reg[1]/NET0131 ,
		_w5180_
	);
	LUT2 #(
		.INIT('he)
	) name3034 (
		_w5179_,
		_w5180_,
		_w5181_
	);
	LUT4 #(
		.INIT('h4ccc)
	) name3035 (
		\u12_o6_we_reg/P0001 ,
		\u5_mem_reg[3][26]/NET0131 ,
		\u5_wp_reg[0]/P0001 ,
		\u5_wp_reg[1]/NET0131 ,
		_w5182_
	);
	LUT4 #(
		.INIT('h8000)
	) name3036 (
		\u12_dout_reg[26]/P0001 ,
		\u12_o6_we_reg/P0001 ,
		\u5_wp_reg[0]/P0001 ,
		\u5_wp_reg[1]/NET0131 ,
		_w5183_
	);
	LUT2 #(
		.INIT('he)
	) name3037 (
		_w5182_,
		_w5183_,
		_w5184_
	);
	LUT4 #(
		.INIT('h4ccc)
	) name3038 (
		\u12_o6_we_reg/P0001 ,
		\u5_mem_reg[3][27]/NET0131 ,
		\u5_wp_reg[0]/P0001 ,
		\u5_wp_reg[1]/NET0131 ,
		_w5185_
	);
	LUT4 #(
		.INIT('h8000)
	) name3039 (
		\u12_dout_reg[27]/P0001 ,
		\u12_o6_we_reg/P0001 ,
		\u5_wp_reg[0]/P0001 ,
		\u5_wp_reg[1]/NET0131 ,
		_w5186_
	);
	LUT2 #(
		.INIT('he)
	) name3040 (
		_w5185_,
		_w5186_,
		_w5187_
	);
	LUT4 #(
		.INIT('h4ccc)
	) name3041 (
		\u12_o6_we_reg/P0001 ,
		\u5_mem_reg[3][28]/NET0131 ,
		\u5_wp_reg[0]/P0001 ,
		\u5_wp_reg[1]/NET0131 ,
		_w5188_
	);
	LUT4 #(
		.INIT('h8000)
	) name3042 (
		\u12_dout_reg[28]/P0001 ,
		\u12_o6_we_reg/P0001 ,
		\u5_wp_reg[0]/P0001 ,
		\u5_wp_reg[1]/NET0131 ,
		_w5189_
	);
	LUT2 #(
		.INIT('he)
	) name3043 (
		_w5188_,
		_w5189_,
		_w5190_
	);
	LUT4 #(
		.INIT('h4ccc)
	) name3044 (
		\u12_o6_we_reg/P0001 ,
		\u5_mem_reg[3][29]/NET0131 ,
		\u5_wp_reg[0]/P0001 ,
		\u5_wp_reg[1]/NET0131 ,
		_w5191_
	);
	LUT4 #(
		.INIT('h8000)
	) name3045 (
		\u12_dout_reg[29]/P0001 ,
		\u12_o6_we_reg/P0001 ,
		\u5_wp_reg[0]/P0001 ,
		\u5_wp_reg[1]/NET0131 ,
		_w5192_
	);
	LUT2 #(
		.INIT('he)
	) name3046 (
		_w5191_,
		_w5192_,
		_w5193_
	);
	LUT4 #(
		.INIT('h4ccc)
	) name3047 (
		\u12_o6_we_reg/P0001 ,
		\u5_mem_reg[3][2]/NET0131 ,
		\u5_wp_reg[0]/P0001 ,
		\u5_wp_reg[1]/NET0131 ,
		_w5194_
	);
	LUT4 #(
		.INIT('h8000)
	) name3048 (
		\u12_dout_reg[2]/P0001 ,
		\u12_o6_we_reg/P0001 ,
		\u5_wp_reg[0]/P0001 ,
		\u5_wp_reg[1]/NET0131 ,
		_w5195_
	);
	LUT2 #(
		.INIT('he)
	) name3049 (
		_w5194_,
		_w5195_,
		_w5196_
	);
	LUT4 #(
		.INIT('h4ccc)
	) name3050 (
		\u12_o6_we_reg/P0001 ,
		\u5_mem_reg[3][30]/NET0131 ,
		\u5_wp_reg[0]/P0001 ,
		\u5_wp_reg[1]/NET0131 ,
		_w5197_
	);
	LUT4 #(
		.INIT('h8000)
	) name3051 (
		\u12_dout_reg[30]/P0001 ,
		\u12_o6_we_reg/P0001 ,
		\u5_wp_reg[0]/P0001 ,
		\u5_wp_reg[1]/NET0131 ,
		_w5198_
	);
	LUT2 #(
		.INIT('he)
	) name3052 (
		_w5197_,
		_w5198_,
		_w5199_
	);
	LUT4 #(
		.INIT('h4ccc)
	) name3053 (
		\u12_o6_we_reg/P0001 ,
		\u5_mem_reg[3][31]/NET0131 ,
		\u5_wp_reg[0]/P0001 ,
		\u5_wp_reg[1]/NET0131 ,
		_w5200_
	);
	LUT4 #(
		.INIT('h8000)
	) name3054 (
		\u12_dout_reg[31]/P0001 ,
		\u12_o6_we_reg/P0001 ,
		\u5_wp_reg[0]/P0001 ,
		\u5_wp_reg[1]/NET0131 ,
		_w5201_
	);
	LUT2 #(
		.INIT('he)
	) name3055 (
		_w5200_,
		_w5201_,
		_w5202_
	);
	LUT4 #(
		.INIT('h4ccc)
	) name3056 (
		\u12_o6_we_reg/P0001 ,
		\u5_mem_reg[3][3]/NET0131 ,
		\u5_wp_reg[0]/P0001 ,
		\u5_wp_reg[1]/NET0131 ,
		_w5203_
	);
	LUT4 #(
		.INIT('h8000)
	) name3057 (
		\u12_dout_reg[3]/P0001 ,
		\u12_o6_we_reg/P0001 ,
		\u5_wp_reg[0]/P0001 ,
		\u5_wp_reg[1]/NET0131 ,
		_w5204_
	);
	LUT2 #(
		.INIT('he)
	) name3058 (
		_w5203_,
		_w5204_,
		_w5205_
	);
	LUT4 #(
		.INIT('h4ccc)
	) name3059 (
		\u12_o6_we_reg/P0001 ,
		\u5_mem_reg[3][4]/NET0131 ,
		\u5_wp_reg[0]/P0001 ,
		\u5_wp_reg[1]/NET0131 ,
		_w5206_
	);
	LUT4 #(
		.INIT('h8000)
	) name3060 (
		\u12_dout_reg[4]/P0001 ,
		\u12_o6_we_reg/P0001 ,
		\u5_wp_reg[0]/P0001 ,
		\u5_wp_reg[1]/NET0131 ,
		_w5207_
	);
	LUT2 #(
		.INIT('he)
	) name3061 (
		_w5206_,
		_w5207_,
		_w5208_
	);
	LUT4 #(
		.INIT('h4ccc)
	) name3062 (
		\u12_o6_we_reg/P0001 ,
		\u5_mem_reg[3][5]/NET0131 ,
		\u5_wp_reg[0]/P0001 ,
		\u5_wp_reg[1]/NET0131 ,
		_w5209_
	);
	LUT4 #(
		.INIT('h8000)
	) name3063 (
		\u12_dout_reg[5]/P0001 ,
		\u12_o6_we_reg/P0001 ,
		\u5_wp_reg[0]/P0001 ,
		\u5_wp_reg[1]/NET0131 ,
		_w5210_
	);
	LUT2 #(
		.INIT('he)
	) name3064 (
		_w5209_,
		_w5210_,
		_w5211_
	);
	LUT4 #(
		.INIT('h4ccc)
	) name3065 (
		\u12_o6_we_reg/P0001 ,
		\u5_mem_reg[3][6]/NET0131 ,
		\u5_wp_reg[0]/P0001 ,
		\u5_wp_reg[1]/NET0131 ,
		_w5212_
	);
	LUT4 #(
		.INIT('h8000)
	) name3066 (
		\u12_dout_reg[6]/P0001 ,
		\u12_o6_we_reg/P0001 ,
		\u5_wp_reg[0]/P0001 ,
		\u5_wp_reg[1]/NET0131 ,
		_w5213_
	);
	LUT2 #(
		.INIT('he)
	) name3067 (
		_w5212_,
		_w5213_,
		_w5214_
	);
	LUT4 #(
		.INIT('h4ccc)
	) name3068 (
		\u12_o6_we_reg/P0001 ,
		\u5_mem_reg[3][7]/NET0131 ,
		\u5_wp_reg[0]/P0001 ,
		\u5_wp_reg[1]/NET0131 ,
		_w5215_
	);
	LUT4 #(
		.INIT('h8000)
	) name3069 (
		\u12_dout_reg[7]/P0001 ,
		\u12_o6_we_reg/P0001 ,
		\u5_wp_reg[0]/P0001 ,
		\u5_wp_reg[1]/NET0131 ,
		_w5216_
	);
	LUT2 #(
		.INIT('he)
	) name3070 (
		_w5215_,
		_w5216_,
		_w5217_
	);
	LUT4 #(
		.INIT('h4ccc)
	) name3071 (
		\u12_o6_we_reg/P0001 ,
		\u5_mem_reg[3][8]/NET0131 ,
		\u5_wp_reg[0]/P0001 ,
		\u5_wp_reg[1]/NET0131 ,
		_w5218_
	);
	LUT4 #(
		.INIT('h8000)
	) name3072 (
		\u12_dout_reg[8]/P0001 ,
		\u12_o6_we_reg/P0001 ,
		\u5_wp_reg[0]/P0001 ,
		\u5_wp_reg[1]/NET0131 ,
		_w5219_
	);
	LUT2 #(
		.INIT('he)
	) name3073 (
		_w5218_,
		_w5219_,
		_w5220_
	);
	LUT4 #(
		.INIT('h4ccc)
	) name3074 (
		\u12_o6_we_reg/P0001 ,
		\u5_mem_reg[3][9]/NET0131 ,
		\u5_wp_reg[0]/P0001 ,
		\u5_wp_reg[1]/NET0131 ,
		_w5221_
	);
	LUT4 #(
		.INIT('h8000)
	) name3075 (
		\u12_dout_reg[9]/P0001 ,
		\u12_o6_we_reg/P0001 ,
		\u5_wp_reg[0]/P0001 ,
		\u5_wp_reg[1]/NET0131 ,
		_w5222_
	);
	LUT2 #(
		.INIT('he)
	) name3076 (
		_w5221_,
		_w5222_,
		_w5223_
	);
	LUT4 #(
		.INIT('h4ccc)
	) name3077 (
		\u12_o9_we_reg/P0001 ,
		\u8_mem_reg[3][6]/NET0131 ,
		\u8_wp_reg[0]/P0001 ,
		\u8_wp_reg[1]/NET0131 ,
		_w5224_
	);
	LUT4 #(
		.INIT('h8000)
	) name3078 (
		\u12_dout_reg[6]/P0001 ,
		\u12_o9_we_reg/P0001 ,
		\u8_wp_reg[0]/P0001 ,
		\u8_wp_reg[1]/NET0131 ,
		_w5225_
	);
	LUT2 #(
		.INIT('he)
	) name3079 (
		_w5224_,
		_w5225_,
		_w5226_
	);
	LUT4 #(
		.INIT('hcc4c)
	) name3080 (
		\u12_o9_we_reg/P0001 ,
		\u8_mem_reg[1][28]/NET0131 ,
		\u8_wp_reg[0]/P0001 ,
		\u8_wp_reg[1]/NET0131 ,
		_w5227_
	);
	LUT4 #(
		.INIT('h0080)
	) name3081 (
		\u12_dout_reg[28]/P0001 ,
		\u12_o9_we_reg/P0001 ,
		\u8_wp_reg[0]/P0001 ,
		\u8_wp_reg[1]/NET0131 ,
		_w5228_
	);
	LUT2 #(
		.INIT('he)
	) name3082 (
		_w5227_,
		_w5228_,
		_w5229_
	);
	LUT4 #(
		.INIT('hc4cc)
	) name3083 (
		\u12_o3_we_reg/P0001 ,
		\u3_mem_reg[2][20]/NET0131 ,
		\u3_wp_reg[0]/P0001 ,
		\u3_wp_reg[1]/NET0131 ,
		_w5230_
	);
	LUT4 #(
		.INIT('h0800)
	) name3084 (
		\u12_dout_reg[20]/P0001 ,
		\u12_o3_we_reg/P0001 ,
		\u3_wp_reg[0]/P0001 ,
		\u3_wp_reg[1]/NET0131 ,
		_w5231_
	);
	LUT2 #(
		.INIT('he)
	) name3085 (
		_w5230_,
		_w5231_,
		_w5232_
	);
	LUT4 #(
		.INIT('h4ccc)
	) name3086 (
		\u12_o9_we_reg/P0001 ,
		\u8_mem_reg[3][31]/NET0131 ,
		\u8_wp_reg[0]/P0001 ,
		\u8_wp_reg[1]/NET0131 ,
		_w5233_
	);
	LUT4 #(
		.INIT('h8000)
	) name3087 (
		\u12_dout_reg[31]/P0001 ,
		\u12_o9_we_reg/P0001 ,
		\u8_wp_reg[0]/P0001 ,
		\u8_wp_reg[1]/NET0131 ,
		_w5234_
	);
	LUT2 #(
		.INIT('he)
	) name3088 (
		_w5233_,
		_w5234_,
		_w5235_
	);
	LUT4 #(
		.INIT('hcc4c)
	) name3089 (
		\u12_o7_we_reg/P0001 ,
		\u6_mem_reg[1][0]/NET0131 ,
		\u6_wp_reg[0]/P0001 ,
		\u6_wp_reg[1]/NET0131 ,
		_w5236_
	);
	LUT4 #(
		.INIT('h0080)
	) name3090 (
		\u12_dout_reg[0]/P0001 ,
		\u12_o7_we_reg/P0001 ,
		\u6_wp_reg[0]/P0001 ,
		\u6_wp_reg[1]/NET0131 ,
		_w5237_
	);
	LUT2 #(
		.INIT('he)
	) name3091 (
		_w5236_,
		_w5237_,
		_w5238_
	);
	LUT4 #(
		.INIT('hcc4c)
	) name3092 (
		\u12_o7_we_reg/P0001 ,
		\u6_mem_reg[1][10]/NET0131 ,
		\u6_wp_reg[0]/P0001 ,
		\u6_wp_reg[1]/NET0131 ,
		_w5239_
	);
	LUT4 #(
		.INIT('h0080)
	) name3093 (
		\u12_dout_reg[10]/P0001 ,
		\u12_o7_we_reg/P0001 ,
		\u6_wp_reg[0]/P0001 ,
		\u6_wp_reg[1]/NET0131 ,
		_w5240_
	);
	LUT2 #(
		.INIT('he)
	) name3094 (
		_w5239_,
		_w5240_,
		_w5241_
	);
	LUT4 #(
		.INIT('hcc4c)
	) name3095 (
		\u12_o7_we_reg/P0001 ,
		\u6_mem_reg[1][11]/NET0131 ,
		\u6_wp_reg[0]/P0001 ,
		\u6_wp_reg[1]/NET0131 ,
		_w5242_
	);
	LUT4 #(
		.INIT('h0080)
	) name3096 (
		\u12_dout_reg[11]/P0001 ,
		\u12_o7_we_reg/P0001 ,
		\u6_wp_reg[0]/P0001 ,
		\u6_wp_reg[1]/NET0131 ,
		_w5243_
	);
	LUT2 #(
		.INIT('he)
	) name3097 (
		_w5242_,
		_w5243_,
		_w5244_
	);
	LUT4 #(
		.INIT('hcc4c)
	) name3098 (
		\u12_o7_we_reg/P0001 ,
		\u6_mem_reg[1][12]/NET0131 ,
		\u6_wp_reg[0]/P0001 ,
		\u6_wp_reg[1]/NET0131 ,
		_w5245_
	);
	LUT4 #(
		.INIT('h0080)
	) name3099 (
		\u12_dout_reg[12]/P0001 ,
		\u12_o7_we_reg/P0001 ,
		\u6_wp_reg[0]/P0001 ,
		\u6_wp_reg[1]/NET0131 ,
		_w5246_
	);
	LUT2 #(
		.INIT('he)
	) name3100 (
		_w5245_,
		_w5246_,
		_w5247_
	);
	LUT4 #(
		.INIT('hcc4c)
	) name3101 (
		\u12_o7_we_reg/P0001 ,
		\u6_mem_reg[1][13]/NET0131 ,
		\u6_wp_reg[0]/P0001 ,
		\u6_wp_reg[1]/NET0131 ,
		_w5248_
	);
	LUT4 #(
		.INIT('h0080)
	) name3102 (
		\u12_dout_reg[13]/P0001 ,
		\u12_o7_we_reg/P0001 ,
		\u6_wp_reg[0]/P0001 ,
		\u6_wp_reg[1]/NET0131 ,
		_w5249_
	);
	LUT2 #(
		.INIT('he)
	) name3103 (
		_w5248_,
		_w5249_,
		_w5250_
	);
	LUT4 #(
		.INIT('hcc4c)
	) name3104 (
		\u12_o7_we_reg/P0001 ,
		\u6_mem_reg[1][14]/NET0131 ,
		\u6_wp_reg[0]/P0001 ,
		\u6_wp_reg[1]/NET0131 ,
		_w5251_
	);
	LUT4 #(
		.INIT('h0080)
	) name3105 (
		\u12_dout_reg[14]/P0001 ,
		\u12_o7_we_reg/P0001 ,
		\u6_wp_reg[0]/P0001 ,
		\u6_wp_reg[1]/NET0131 ,
		_w5252_
	);
	LUT2 #(
		.INIT('he)
	) name3106 (
		_w5251_,
		_w5252_,
		_w5253_
	);
	LUT4 #(
		.INIT('hcc4c)
	) name3107 (
		\u12_o7_we_reg/P0001 ,
		\u6_mem_reg[1][15]/NET0131 ,
		\u6_wp_reg[0]/P0001 ,
		\u6_wp_reg[1]/NET0131 ,
		_w5254_
	);
	LUT4 #(
		.INIT('h0080)
	) name3108 (
		\u12_dout_reg[15]/P0001 ,
		\u12_o7_we_reg/P0001 ,
		\u6_wp_reg[0]/P0001 ,
		\u6_wp_reg[1]/NET0131 ,
		_w5255_
	);
	LUT2 #(
		.INIT('he)
	) name3109 (
		_w5254_,
		_w5255_,
		_w5256_
	);
	LUT4 #(
		.INIT('hcc4c)
	) name3110 (
		\u12_o7_we_reg/P0001 ,
		\u6_mem_reg[1][16]/NET0131 ,
		\u6_wp_reg[0]/P0001 ,
		\u6_wp_reg[1]/NET0131 ,
		_w5257_
	);
	LUT4 #(
		.INIT('h0080)
	) name3111 (
		\u12_dout_reg[16]/P0001 ,
		\u12_o7_we_reg/P0001 ,
		\u6_wp_reg[0]/P0001 ,
		\u6_wp_reg[1]/NET0131 ,
		_w5258_
	);
	LUT2 #(
		.INIT('he)
	) name3112 (
		_w5257_,
		_w5258_,
		_w5259_
	);
	LUT4 #(
		.INIT('hcc4c)
	) name3113 (
		\u12_o7_we_reg/P0001 ,
		\u6_mem_reg[1][17]/NET0131 ,
		\u6_wp_reg[0]/P0001 ,
		\u6_wp_reg[1]/NET0131 ,
		_w5260_
	);
	LUT4 #(
		.INIT('h0080)
	) name3114 (
		\u12_dout_reg[17]/P0001 ,
		\u12_o7_we_reg/P0001 ,
		\u6_wp_reg[0]/P0001 ,
		\u6_wp_reg[1]/NET0131 ,
		_w5261_
	);
	LUT2 #(
		.INIT('he)
	) name3115 (
		_w5260_,
		_w5261_,
		_w5262_
	);
	LUT4 #(
		.INIT('hcc4c)
	) name3116 (
		\u12_o7_we_reg/P0001 ,
		\u6_mem_reg[1][18]/NET0131 ,
		\u6_wp_reg[0]/P0001 ,
		\u6_wp_reg[1]/NET0131 ,
		_w5263_
	);
	LUT4 #(
		.INIT('h0080)
	) name3117 (
		\u12_dout_reg[18]/P0001 ,
		\u12_o7_we_reg/P0001 ,
		\u6_wp_reg[0]/P0001 ,
		\u6_wp_reg[1]/NET0131 ,
		_w5264_
	);
	LUT2 #(
		.INIT('he)
	) name3118 (
		_w5263_,
		_w5264_,
		_w5265_
	);
	LUT4 #(
		.INIT('hcc4c)
	) name3119 (
		\u12_o7_we_reg/P0001 ,
		\u6_mem_reg[1][19]/NET0131 ,
		\u6_wp_reg[0]/P0001 ,
		\u6_wp_reg[1]/NET0131 ,
		_w5266_
	);
	LUT4 #(
		.INIT('h0080)
	) name3120 (
		\u12_dout_reg[19]/P0001 ,
		\u12_o7_we_reg/P0001 ,
		\u6_wp_reg[0]/P0001 ,
		\u6_wp_reg[1]/NET0131 ,
		_w5267_
	);
	LUT2 #(
		.INIT('he)
	) name3121 (
		_w5266_,
		_w5267_,
		_w5268_
	);
	LUT4 #(
		.INIT('hcc4c)
	) name3122 (
		\u12_o7_we_reg/P0001 ,
		\u6_mem_reg[1][1]/NET0131 ,
		\u6_wp_reg[0]/P0001 ,
		\u6_wp_reg[1]/NET0131 ,
		_w5269_
	);
	LUT4 #(
		.INIT('h0080)
	) name3123 (
		\u12_dout_reg[1]/P0001 ,
		\u12_o7_we_reg/P0001 ,
		\u6_wp_reg[0]/P0001 ,
		\u6_wp_reg[1]/NET0131 ,
		_w5270_
	);
	LUT2 #(
		.INIT('he)
	) name3124 (
		_w5269_,
		_w5270_,
		_w5271_
	);
	LUT4 #(
		.INIT('hcc4c)
	) name3125 (
		\u12_o7_we_reg/P0001 ,
		\u6_mem_reg[1][20]/NET0131 ,
		\u6_wp_reg[0]/P0001 ,
		\u6_wp_reg[1]/NET0131 ,
		_w5272_
	);
	LUT4 #(
		.INIT('h0080)
	) name3126 (
		\u12_dout_reg[20]/P0001 ,
		\u12_o7_we_reg/P0001 ,
		\u6_wp_reg[0]/P0001 ,
		\u6_wp_reg[1]/NET0131 ,
		_w5273_
	);
	LUT2 #(
		.INIT('he)
	) name3127 (
		_w5272_,
		_w5273_,
		_w5274_
	);
	LUT4 #(
		.INIT('hcc4c)
	) name3128 (
		\u12_o7_we_reg/P0001 ,
		\u6_mem_reg[1][21]/NET0131 ,
		\u6_wp_reg[0]/P0001 ,
		\u6_wp_reg[1]/NET0131 ,
		_w5275_
	);
	LUT4 #(
		.INIT('h0080)
	) name3129 (
		\u12_dout_reg[21]/P0001 ,
		\u12_o7_we_reg/P0001 ,
		\u6_wp_reg[0]/P0001 ,
		\u6_wp_reg[1]/NET0131 ,
		_w5276_
	);
	LUT2 #(
		.INIT('he)
	) name3130 (
		_w5275_,
		_w5276_,
		_w5277_
	);
	LUT4 #(
		.INIT('hcc4c)
	) name3131 (
		\u12_o7_we_reg/P0001 ,
		\u6_mem_reg[1][22]/NET0131 ,
		\u6_wp_reg[0]/P0001 ,
		\u6_wp_reg[1]/NET0131 ,
		_w5278_
	);
	LUT4 #(
		.INIT('h0080)
	) name3132 (
		\u12_dout_reg[22]/P0001 ,
		\u12_o7_we_reg/P0001 ,
		\u6_wp_reg[0]/P0001 ,
		\u6_wp_reg[1]/NET0131 ,
		_w5279_
	);
	LUT2 #(
		.INIT('he)
	) name3133 (
		_w5278_,
		_w5279_,
		_w5280_
	);
	LUT4 #(
		.INIT('hcc4c)
	) name3134 (
		\u12_o7_we_reg/P0001 ,
		\u6_mem_reg[1][23]/NET0131 ,
		\u6_wp_reg[0]/P0001 ,
		\u6_wp_reg[1]/NET0131 ,
		_w5281_
	);
	LUT4 #(
		.INIT('h0080)
	) name3135 (
		\u12_dout_reg[23]/P0001 ,
		\u12_o7_we_reg/P0001 ,
		\u6_wp_reg[0]/P0001 ,
		\u6_wp_reg[1]/NET0131 ,
		_w5282_
	);
	LUT2 #(
		.INIT('he)
	) name3136 (
		_w5281_,
		_w5282_,
		_w5283_
	);
	LUT4 #(
		.INIT('hcc4c)
	) name3137 (
		\u12_o7_we_reg/P0001 ,
		\u6_mem_reg[1][24]/NET0131 ,
		\u6_wp_reg[0]/P0001 ,
		\u6_wp_reg[1]/NET0131 ,
		_w5284_
	);
	LUT4 #(
		.INIT('h0080)
	) name3138 (
		\u12_dout_reg[24]/P0001 ,
		\u12_o7_we_reg/P0001 ,
		\u6_wp_reg[0]/P0001 ,
		\u6_wp_reg[1]/NET0131 ,
		_w5285_
	);
	LUT2 #(
		.INIT('he)
	) name3139 (
		_w5284_,
		_w5285_,
		_w5286_
	);
	LUT4 #(
		.INIT('hcc4c)
	) name3140 (
		\u12_o7_we_reg/P0001 ,
		\u6_mem_reg[1][25]/NET0131 ,
		\u6_wp_reg[0]/P0001 ,
		\u6_wp_reg[1]/NET0131 ,
		_w5287_
	);
	LUT4 #(
		.INIT('h0080)
	) name3141 (
		\u12_dout_reg[25]/P0001 ,
		\u12_o7_we_reg/P0001 ,
		\u6_wp_reg[0]/P0001 ,
		\u6_wp_reg[1]/NET0131 ,
		_w5288_
	);
	LUT2 #(
		.INIT('he)
	) name3142 (
		_w5287_,
		_w5288_,
		_w5289_
	);
	LUT4 #(
		.INIT('hcc4c)
	) name3143 (
		\u12_o7_we_reg/P0001 ,
		\u6_mem_reg[1][26]/NET0131 ,
		\u6_wp_reg[0]/P0001 ,
		\u6_wp_reg[1]/NET0131 ,
		_w5290_
	);
	LUT4 #(
		.INIT('h0080)
	) name3144 (
		\u12_dout_reg[26]/P0001 ,
		\u12_o7_we_reg/P0001 ,
		\u6_wp_reg[0]/P0001 ,
		\u6_wp_reg[1]/NET0131 ,
		_w5291_
	);
	LUT2 #(
		.INIT('he)
	) name3145 (
		_w5290_,
		_w5291_,
		_w5292_
	);
	LUT4 #(
		.INIT('hcc4c)
	) name3146 (
		\u12_o7_we_reg/P0001 ,
		\u6_mem_reg[1][27]/NET0131 ,
		\u6_wp_reg[0]/P0001 ,
		\u6_wp_reg[1]/NET0131 ,
		_w5293_
	);
	LUT4 #(
		.INIT('h0080)
	) name3147 (
		\u12_dout_reg[27]/P0001 ,
		\u12_o7_we_reg/P0001 ,
		\u6_wp_reg[0]/P0001 ,
		\u6_wp_reg[1]/NET0131 ,
		_w5294_
	);
	LUT2 #(
		.INIT('he)
	) name3148 (
		_w5293_,
		_w5294_,
		_w5295_
	);
	LUT4 #(
		.INIT('hcc4c)
	) name3149 (
		\u12_o7_we_reg/P0001 ,
		\u6_mem_reg[1][28]/NET0131 ,
		\u6_wp_reg[0]/P0001 ,
		\u6_wp_reg[1]/NET0131 ,
		_w5296_
	);
	LUT4 #(
		.INIT('h0080)
	) name3150 (
		\u12_dout_reg[28]/P0001 ,
		\u12_o7_we_reg/P0001 ,
		\u6_wp_reg[0]/P0001 ,
		\u6_wp_reg[1]/NET0131 ,
		_w5297_
	);
	LUT2 #(
		.INIT('he)
	) name3151 (
		_w5296_,
		_w5297_,
		_w5298_
	);
	LUT4 #(
		.INIT('hcc4c)
	) name3152 (
		\u12_o7_we_reg/P0001 ,
		\u6_mem_reg[1][29]/NET0131 ,
		\u6_wp_reg[0]/P0001 ,
		\u6_wp_reg[1]/NET0131 ,
		_w5299_
	);
	LUT4 #(
		.INIT('h0080)
	) name3153 (
		\u12_dout_reg[29]/P0001 ,
		\u12_o7_we_reg/P0001 ,
		\u6_wp_reg[0]/P0001 ,
		\u6_wp_reg[1]/NET0131 ,
		_w5300_
	);
	LUT2 #(
		.INIT('he)
	) name3154 (
		_w5299_,
		_w5300_,
		_w5301_
	);
	LUT4 #(
		.INIT('hcc4c)
	) name3155 (
		\u12_o7_we_reg/P0001 ,
		\u6_mem_reg[1][2]/NET0131 ,
		\u6_wp_reg[0]/P0001 ,
		\u6_wp_reg[1]/NET0131 ,
		_w5302_
	);
	LUT4 #(
		.INIT('h0080)
	) name3156 (
		\u12_dout_reg[2]/P0001 ,
		\u12_o7_we_reg/P0001 ,
		\u6_wp_reg[0]/P0001 ,
		\u6_wp_reg[1]/NET0131 ,
		_w5303_
	);
	LUT2 #(
		.INIT('he)
	) name3157 (
		_w5302_,
		_w5303_,
		_w5304_
	);
	LUT4 #(
		.INIT('hcc4c)
	) name3158 (
		\u12_o7_we_reg/P0001 ,
		\u6_mem_reg[1][30]/NET0131 ,
		\u6_wp_reg[0]/P0001 ,
		\u6_wp_reg[1]/NET0131 ,
		_w5305_
	);
	LUT4 #(
		.INIT('h0080)
	) name3159 (
		\u12_dout_reg[30]/P0001 ,
		\u12_o7_we_reg/P0001 ,
		\u6_wp_reg[0]/P0001 ,
		\u6_wp_reg[1]/NET0131 ,
		_w5306_
	);
	LUT2 #(
		.INIT('he)
	) name3160 (
		_w5305_,
		_w5306_,
		_w5307_
	);
	LUT4 #(
		.INIT('hcc4c)
	) name3161 (
		\u12_o7_we_reg/P0001 ,
		\u6_mem_reg[1][31]/NET0131 ,
		\u6_wp_reg[0]/P0001 ,
		\u6_wp_reg[1]/NET0131 ,
		_w5308_
	);
	LUT4 #(
		.INIT('h0080)
	) name3162 (
		\u12_dout_reg[31]/P0001 ,
		\u12_o7_we_reg/P0001 ,
		\u6_wp_reg[0]/P0001 ,
		\u6_wp_reg[1]/NET0131 ,
		_w5309_
	);
	LUT2 #(
		.INIT('he)
	) name3163 (
		_w5308_,
		_w5309_,
		_w5310_
	);
	LUT4 #(
		.INIT('hcc4c)
	) name3164 (
		\u12_o7_we_reg/P0001 ,
		\u6_mem_reg[1][3]/NET0131 ,
		\u6_wp_reg[0]/P0001 ,
		\u6_wp_reg[1]/NET0131 ,
		_w5311_
	);
	LUT4 #(
		.INIT('h0080)
	) name3165 (
		\u12_dout_reg[3]/P0001 ,
		\u12_o7_we_reg/P0001 ,
		\u6_wp_reg[0]/P0001 ,
		\u6_wp_reg[1]/NET0131 ,
		_w5312_
	);
	LUT2 #(
		.INIT('he)
	) name3166 (
		_w5311_,
		_w5312_,
		_w5313_
	);
	LUT4 #(
		.INIT('hcc4c)
	) name3167 (
		\u12_o7_we_reg/P0001 ,
		\u6_mem_reg[1][4]/NET0131 ,
		\u6_wp_reg[0]/P0001 ,
		\u6_wp_reg[1]/NET0131 ,
		_w5314_
	);
	LUT4 #(
		.INIT('h0080)
	) name3168 (
		\u12_dout_reg[4]/P0001 ,
		\u12_o7_we_reg/P0001 ,
		\u6_wp_reg[0]/P0001 ,
		\u6_wp_reg[1]/NET0131 ,
		_w5315_
	);
	LUT2 #(
		.INIT('he)
	) name3169 (
		_w5314_,
		_w5315_,
		_w5316_
	);
	LUT4 #(
		.INIT('hcc4c)
	) name3170 (
		\u12_o7_we_reg/P0001 ,
		\u6_mem_reg[1][5]/NET0131 ,
		\u6_wp_reg[0]/P0001 ,
		\u6_wp_reg[1]/NET0131 ,
		_w5317_
	);
	LUT4 #(
		.INIT('h0080)
	) name3171 (
		\u12_dout_reg[5]/P0001 ,
		\u12_o7_we_reg/P0001 ,
		\u6_wp_reg[0]/P0001 ,
		\u6_wp_reg[1]/NET0131 ,
		_w5318_
	);
	LUT2 #(
		.INIT('he)
	) name3172 (
		_w5317_,
		_w5318_,
		_w5319_
	);
	LUT4 #(
		.INIT('hcc4c)
	) name3173 (
		\u12_o7_we_reg/P0001 ,
		\u6_mem_reg[1][6]/NET0131 ,
		\u6_wp_reg[0]/P0001 ,
		\u6_wp_reg[1]/NET0131 ,
		_w5320_
	);
	LUT4 #(
		.INIT('h0080)
	) name3174 (
		\u12_dout_reg[6]/P0001 ,
		\u12_o7_we_reg/P0001 ,
		\u6_wp_reg[0]/P0001 ,
		\u6_wp_reg[1]/NET0131 ,
		_w5321_
	);
	LUT2 #(
		.INIT('he)
	) name3175 (
		_w5320_,
		_w5321_,
		_w5322_
	);
	LUT4 #(
		.INIT('hcc4c)
	) name3176 (
		\u12_o7_we_reg/P0001 ,
		\u6_mem_reg[1][7]/NET0131 ,
		\u6_wp_reg[0]/P0001 ,
		\u6_wp_reg[1]/NET0131 ,
		_w5323_
	);
	LUT4 #(
		.INIT('h0080)
	) name3177 (
		\u12_dout_reg[7]/P0001 ,
		\u12_o7_we_reg/P0001 ,
		\u6_wp_reg[0]/P0001 ,
		\u6_wp_reg[1]/NET0131 ,
		_w5324_
	);
	LUT2 #(
		.INIT('he)
	) name3178 (
		_w5323_,
		_w5324_,
		_w5325_
	);
	LUT4 #(
		.INIT('hcc4c)
	) name3179 (
		\u12_o7_we_reg/P0001 ,
		\u6_mem_reg[1][8]/NET0131 ,
		\u6_wp_reg[0]/P0001 ,
		\u6_wp_reg[1]/NET0131 ,
		_w5326_
	);
	LUT4 #(
		.INIT('h0080)
	) name3180 (
		\u12_dout_reg[8]/P0001 ,
		\u12_o7_we_reg/P0001 ,
		\u6_wp_reg[0]/P0001 ,
		\u6_wp_reg[1]/NET0131 ,
		_w5327_
	);
	LUT2 #(
		.INIT('he)
	) name3181 (
		_w5326_,
		_w5327_,
		_w5328_
	);
	LUT4 #(
		.INIT('hcc4c)
	) name3182 (
		\u12_o7_we_reg/P0001 ,
		\u6_mem_reg[1][9]/NET0131 ,
		\u6_wp_reg[0]/P0001 ,
		\u6_wp_reg[1]/NET0131 ,
		_w5329_
	);
	LUT4 #(
		.INIT('h0080)
	) name3183 (
		\u12_dout_reg[9]/P0001 ,
		\u12_o7_we_reg/P0001 ,
		\u6_wp_reg[0]/P0001 ,
		\u6_wp_reg[1]/NET0131 ,
		_w5330_
	);
	LUT2 #(
		.INIT('he)
	) name3184 (
		_w5329_,
		_w5330_,
		_w5331_
	);
	LUT4 #(
		.INIT('hc4cc)
	) name3185 (
		\u12_o7_we_reg/P0001 ,
		\u6_mem_reg[2][0]/NET0131 ,
		\u6_wp_reg[0]/P0001 ,
		\u6_wp_reg[1]/NET0131 ,
		_w5332_
	);
	LUT4 #(
		.INIT('h0800)
	) name3186 (
		\u12_dout_reg[0]/P0001 ,
		\u12_o7_we_reg/P0001 ,
		\u6_wp_reg[0]/P0001 ,
		\u6_wp_reg[1]/NET0131 ,
		_w5333_
	);
	LUT2 #(
		.INIT('he)
	) name3187 (
		_w5332_,
		_w5333_,
		_w5334_
	);
	LUT4 #(
		.INIT('hc4cc)
	) name3188 (
		\u12_o7_we_reg/P0001 ,
		\u6_mem_reg[2][10]/NET0131 ,
		\u6_wp_reg[0]/P0001 ,
		\u6_wp_reg[1]/NET0131 ,
		_w5335_
	);
	LUT4 #(
		.INIT('h0800)
	) name3189 (
		\u12_dout_reg[10]/P0001 ,
		\u12_o7_we_reg/P0001 ,
		\u6_wp_reg[0]/P0001 ,
		\u6_wp_reg[1]/NET0131 ,
		_w5336_
	);
	LUT2 #(
		.INIT('he)
	) name3190 (
		_w5335_,
		_w5336_,
		_w5337_
	);
	LUT4 #(
		.INIT('hc4cc)
	) name3191 (
		\u12_o7_we_reg/P0001 ,
		\u6_mem_reg[2][11]/NET0131 ,
		\u6_wp_reg[0]/P0001 ,
		\u6_wp_reg[1]/NET0131 ,
		_w5338_
	);
	LUT4 #(
		.INIT('h0800)
	) name3192 (
		\u12_dout_reg[11]/P0001 ,
		\u12_o7_we_reg/P0001 ,
		\u6_wp_reg[0]/P0001 ,
		\u6_wp_reg[1]/NET0131 ,
		_w5339_
	);
	LUT2 #(
		.INIT('he)
	) name3193 (
		_w5338_,
		_w5339_,
		_w5340_
	);
	LUT4 #(
		.INIT('hc4cc)
	) name3194 (
		\u12_o7_we_reg/P0001 ,
		\u6_mem_reg[2][12]/NET0131 ,
		\u6_wp_reg[0]/P0001 ,
		\u6_wp_reg[1]/NET0131 ,
		_w5341_
	);
	LUT4 #(
		.INIT('h0800)
	) name3195 (
		\u12_dout_reg[12]/P0001 ,
		\u12_o7_we_reg/P0001 ,
		\u6_wp_reg[0]/P0001 ,
		\u6_wp_reg[1]/NET0131 ,
		_w5342_
	);
	LUT2 #(
		.INIT('he)
	) name3196 (
		_w5341_,
		_w5342_,
		_w5343_
	);
	LUT4 #(
		.INIT('hc4cc)
	) name3197 (
		\u12_o7_we_reg/P0001 ,
		\u6_mem_reg[2][13]/NET0131 ,
		\u6_wp_reg[0]/P0001 ,
		\u6_wp_reg[1]/NET0131 ,
		_w5344_
	);
	LUT4 #(
		.INIT('h0800)
	) name3198 (
		\u12_dout_reg[13]/P0001 ,
		\u12_o7_we_reg/P0001 ,
		\u6_wp_reg[0]/P0001 ,
		\u6_wp_reg[1]/NET0131 ,
		_w5345_
	);
	LUT2 #(
		.INIT('he)
	) name3199 (
		_w5344_,
		_w5345_,
		_w5346_
	);
	LUT4 #(
		.INIT('hc4cc)
	) name3200 (
		\u12_o7_we_reg/P0001 ,
		\u6_mem_reg[2][14]/NET0131 ,
		\u6_wp_reg[0]/P0001 ,
		\u6_wp_reg[1]/NET0131 ,
		_w5347_
	);
	LUT4 #(
		.INIT('h0800)
	) name3201 (
		\u12_dout_reg[14]/P0001 ,
		\u12_o7_we_reg/P0001 ,
		\u6_wp_reg[0]/P0001 ,
		\u6_wp_reg[1]/NET0131 ,
		_w5348_
	);
	LUT2 #(
		.INIT('he)
	) name3202 (
		_w5347_,
		_w5348_,
		_w5349_
	);
	LUT4 #(
		.INIT('hc4cc)
	) name3203 (
		\u12_o7_we_reg/P0001 ,
		\u6_mem_reg[2][15]/NET0131 ,
		\u6_wp_reg[0]/P0001 ,
		\u6_wp_reg[1]/NET0131 ,
		_w5350_
	);
	LUT4 #(
		.INIT('h0800)
	) name3204 (
		\u12_dout_reg[15]/P0001 ,
		\u12_o7_we_reg/P0001 ,
		\u6_wp_reg[0]/P0001 ,
		\u6_wp_reg[1]/NET0131 ,
		_w5351_
	);
	LUT2 #(
		.INIT('he)
	) name3205 (
		_w5350_,
		_w5351_,
		_w5352_
	);
	LUT4 #(
		.INIT('hc4cc)
	) name3206 (
		\u12_o7_we_reg/P0001 ,
		\u6_mem_reg[2][16]/NET0131 ,
		\u6_wp_reg[0]/P0001 ,
		\u6_wp_reg[1]/NET0131 ,
		_w5353_
	);
	LUT4 #(
		.INIT('h0800)
	) name3207 (
		\u12_dout_reg[16]/P0001 ,
		\u12_o7_we_reg/P0001 ,
		\u6_wp_reg[0]/P0001 ,
		\u6_wp_reg[1]/NET0131 ,
		_w5354_
	);
	LUT2 #(
		.INIT('he)
	) name3208 (
		_w5353_,
		_w5354_,
		_w5355_
	);
	LUT4 #(
		.INIT('hc4cc)
	) name3209 (
		\u12_o7_we_reg/P0001 ,
		\u6_mem_reg[2][17]/NET0131 ,
		\u6_wp_reg[0]/P0001 ,
		\u6_wp_reg[1]/NET0131 ,
		_w5356_
	);
	LUT4 #(
		.INIT('h0800)
	) name3210 (
		\u12_dout_reg[17]/P0001 ,
		\u12_o7_we_reg/P0001 ,
		\u6_wp_reg[0]/P0001 ,
		\u6_wp_reg[1]/NET0131 ,
		_w5357_
	);
	LUT2 #(
		.INIT('he)
	) name3211 (
		_w5356_,
		_w5357_,
		_w5358_
	);
	LUT4 #(
		.INIT('hc4cc)
	) name3212 (
		\u12_o7_we_reg/P0001 ,
		\u6_mem_reg[2][18]/NET0131 ,
		\u6_wp_reg[0]/P0001 ,
		\u6_wp_reg[1]/NET0131 ,
		_w5359_
	);
	LUT4 #(
		.INIT('h0800)
	) name3213 (
		\u12_dout_reg[18]/P0001 ,
		\u12_o7_we_reg/P0001 ,
		\u6_wp_reg[0]/P0001 ,
		\u6_wp_reg[1]/NET0131 ,
		_w5360_
	);
	LUT2 #(
		.INIT('he)
	) name3214 (
		_w5359_,
		_w5360_,
		_w5361_
	);
	LUT4 #(
		.INIT('hc4cc)
	) name3215 (
		\u12_o7_we_reg/P0001 ,
		\u6_mem_reg[2][19]/NET0131 ,
		\u6_wp_reg[0]/P0001 ,
		\u6_wp_reg[1]/NET0131 ,
		_w5362_
	);
	LUT4 #(
		.INIT('h0800)
	) name3216 (
		\u12_dout_reg[19]/P0001 ,
		\u12_o7_we_reg/P0001 ,
		\u6_wp_reg[0]/P0001 ,
		\u6_wp_reg[1]/NET0131 ,
		_w5363_
	);
	LUT2 #(
		.INIT('he)
	) name3217 (
		_w5362_,
		_w5363_,
		_w5364_
	);
	LUT4 #(
		.INIT('hc4cc)
	) name3218 (
		\u12_o7_we_reg/P0001 ,
		\u6_mem_reg[2][1]/NET0131 ,
		\u6_wp_reg[0]/P0001 ,
		\u6_wp_reg[1]/NET0131 ,
		_w5365_
	);
	LUT4 #(
		.INIT('h0800)
	) name3219 (
		\u12_dout_reg[1]/P0001 ,
		\u12_o7_we_reg/P0001 ,
		\u6_wp_reg[0]/P0001 ,
		\u6_wp_reg[1]/NET0131 ,
		_w5366_
	);
	LUT2 #(
		.INIT('he)
	) name3220 (
		_w5365_,
		_w5366_,
		_w5367_
	);
	LUT4 #(
		.INIT('hc4cc)
	) name3221 (
		\u12_o7_we_reg/P0001 ,
		\u6_mem_reg[2][20]/NET0131 ,
		\u6_wp_reg[0]/P0001 ,
		\u6_wp_reg[1]/NET0131 ,
		_w5368_
	);
	LUT4 #(
		.INIT('h0800)
	) name3222 (
		\u12_dout_reg[20]/P0001 ,
		\u12_o7_we_reg/P0001 ,
		\u6_wp_reg[0]/P0001 ,
		\u6_wp_reg[1]/NET0131 ,
		_w5369_
	);
	LUT2 #(
		.INIT('he)
	) name3223 (
		_w5368_,
		_w5369_,
		_w5370_
	);
	LUT4 #(
		.INIT('hc4cc)
	) name3224 (
		\u12_o7_we_reg/P0001 ,
		\u6_mem_reg[2][21]/NET0131 ,
		\u6_wp_reg[0]/P0001 ,
		\u6_wp_reg[1]/NET0131 ,
		_w5371_
	);
	LUT4 #(
		.INIT('h0800)
	) name3225 (
		\u12_dout_reg[21]/P0001 ,
		\u12_o7_we_reg/P0001 ,
		\u6_wp_reg[0]/P0001 ,
		\u6_wp_reg[1]/NET0131 ,
		_w5372_
	);
	LUT2 #(
		.INIT('he)
	) name3226 (
		_w5371_,
		_w5372_,
		_w5373_
	);
	LUT4 #(
		.INIT('hc4cc)
	) name3227 (
		\u12_o7_we_reg/P0001 ,
		\u6_mem_reg[2][22]/NET0131 ,
		\u6_wp_reg[0]/P0001 ,
		\u6_wp_reg[1]/NET0131 ,
		_w5374_
	);
	LUT4 #(
		.INIT('h0800)
	) name3228 (
		\u12_dout_reg[22]/P0001 ,
		\u12_o7_we_reg/P0001 ,
		\u6_wp_reg[0]/P0001 ,
		\u6_wp_reg[1]/NET0131 ,
		_w5375_
	);
	LUT2 #(
		.INIT('he)
	) name3229 (
		_w5374_,
		_w5375_,
		_w5376_
	);
	LUT4 #(
		.INIT('hc4cc)
	) name3230 (
		\u12_o7_we_reg/P0001 ,
		\u6_mem_reg[2][23]/NET0131 ,
		\u6_wp_reg[0]/P0001 ,
		\u6_wp_reg[1]/NET0131 ,
		_w5377_
	);
	LUT4 #(
		.INIT('h0800)
	) name3231 (
		\u12_dout_reg[23]/P0001 ,
		\u12_o7_we_reg/P0001 ,
		\u6_wp_reg[0]/P0001 ,
		\u6_wp_reg[1]/NET0131 ,
		_w5378_
	);
	LUT2 #(
		.INIT('he)
	) name3232 (
		_w5377_,
		_w5378_,
		_w5379_
	);
	LUT4 #(
		.INIT('hc4cc)
	) name3233 (
		\u12_o7_we_reg/P0001 ,
		\u6_mem_reg[2][24]/NET0131 ,
		\u6_wp_reg[0]/P0001 ,
		\u6_wp_reg[1]/NET0131 ,
		_w5380_
	);
	LUT4 #(
		.INIT('h0800)
	) name3234 (
		\u12_dout_reg[24]/P0001 ,
		\u12_o7_we_reg/P0001 ,
		\u6_wp_reg[0]/P0001 ,
		\u6_wp_reg[1]/NET0131 ,
		_w5381_
	);
	LUT2 #(
		.INIT('he)
	) name3235 (
		_w5380_,
		_w5381_,
		_w5382_
	);
	LUT4 #(
		.INIT('hc4cc)
	) name3236 (
		\u12_o7_we_reg/P0001 ,
		\u6_mem_reg[2][25]/NET0131 ,
		\u6_wp_reg[0]/P0001 ,
		\u6_wp_reg[1]/NET0131 ,
		_w5383_
	);
	LUT4 #(
		.INIT('h0800)
	) name3237 (
		\u12_dout_reg[25]/P0001 ,
		\u12_o7_we_reg/P0001 ,
		\u6_wp_reg[0]/P0001 ,
		\u6_wp_reg[1]/NET0131 ,
		_w5384_
	);
	LUT2 #(
		.INIT('he)
	) name3238 (
		_w5383_,
		_w5384_,
		_w5385_
	);
	LUT4 #(
		.INIT('hc4cc)
	) name3239 (
		\u12_o7_we_reg/P0001 ,
		\u6_mem_reg[2][26]/NET0131 ,
		\u6_wp_reg[0]/P0001 ,
		\u6_wp_reg[1]/NET0131 ,
		_w5386_
	);
	LUT4 #(
		.INIT('h0800)
	) name3240 (
		\u12_dout_reg[26]/P0001 ,
		\u12_o7_we_reg/P0001 ,
		\u6_wp_reg[0]/P0001 ,
		\u6_wp_reg[1]/NET0131 ,
		_w5387_
	);
	LUT2 #(
		.INIT('he)
	) name3241 (
		_w5386_,
		_w5387_,
		_w5388_
	);
	LUT4 #(
		.INIT('hc4cc)
	) name3242 (
		\u12_o7_we_reg/P0001 ,
		\u6_mem_reg[2][27]/NET0131 ,
		\u6_wp_reg[0]/P0001 ,
		\u6_wp_reg[1]/NET0131 ,
		_w5389_
	);
	LUT4 #(
		.INIT('h0800)
	) name3243 (
		\u12_dout_reg[27]/P0001 ,
		\u12_o7_we_reg/P0001 ,
		\u6_wp_reg[0]/P0001 ,
		\u6_wp_reg[1]/NET0131 ,
		_w5390_
	);
	LUT2 #(
		.INIT('he)
	) name3244 (
		_w5389_,
		_w5390_,
		_w5391_
	);
	LUT4 #(
		.INIT('hc4cc)
	) name3245 (
		\u12_o7_we_reg/P0001 ,
		\u6_mem_reg[2][28]/NET0131 ,
		\u6_wp_reg[0]/P0001 ,
		\u6_wp_reg[1]/NET0131 ,
		_w5392_
	);
	LUT4 #(
		.INIT('h0800)
	) name3246 (
		\u12_dout_reg[28]/P0001 ,
		\u12_o7_we_reg/P0001 ,
		\u6_wp_reg[0]/P0001 ,
		\u6_wp_reg[1]/NET0131 ,
		_w5393_
	);
	LUT2 #(
		.INIT('he)
	) name3247 (
		_w5392_,
		_w5393_,
		_w5394_
	);
	LUT4 #(
		.INIT('hc4cc)
	) name3248 (
		\u12_o7_we_reg/P0001 ,
		\u6_mem_reg[2][29]/NET0131 ,
		\u6_wp_reg[0]/P0001 ,
		\u6_wp_reg[1]/NET0131 ,
		_w5395_
	);
	LUT4 #(
		.INIT('h0800)
	) name3249 (
		\u12_dout_reg[29]/P0001 ,
		\u12_o7_we_reg/P0001 ,
		\u6_wp_reg[0]/P0001 ,
		\u6_wp_reg[1]/NET0131 ,
		_w5396_
	);
	LUT2 #(
		.INIT('he)
	) name3250 (
		_w5395_,
		_w5396_,
		_w5397_
	);
	LUT4 #(
		.INIT('hc4cc)
	) name3251 (
		\u12_o7_we_reg/P0001 ,
		\u6_mem_reg[2][2]/NET0131 ,
		\u6_wp_reg[0]/P0001 ,
		\u6_wp_reg[1]/NET0131 ,
		_w5398_
	);
	LUT4 #(
		.INIT('h0800)
	) name3252 (
		\u12_dout_reg[2]/P0001 ,
		\u12_o7_we_reg/P0001 ,
		\u6_wp_reg[0]/P0001 ,
		\u6_wp_reg[1]/NET0131 ,
		_w5399_
	);
	LUT2 #(
		.INIT('he)
	) name3253 (
		_w5398_,
		_w5399_,
		_w5400_
	);
	LUT4 #(
		.INIT('hc4cc)
	) name3254 (
		\u12_o7_we_reg/P0001 ,
		\u6_mem_reg[2][30]/NET0131 ,
		\u6_wp_reg[0]/P0001 ,
		\u6_wp_reg[1]/NET0131 ,
		_w5401_
	);
	LUT4 #(
		.INIT('h0800)
	) name3255 (
		\u12_dout_reg[30]/P0001 ,
		\u12_o7_we_reg/P0001 ,
		\u6_wp_reg[0]/P0001 ,
		\u6_wp_reg[1]/NET0131 ,
		_w5402_
	);
	LUT2 #(
		.INIT('he)
	) name3256 (
		_w5401_,
		_w5402_,
		_w5403_
	);
	LUT4 #(
		.INIT('hc4cc)
	) name3257 (
		\u12_o7_we_reg/P0001 ,
		\u6_mem_reg[2][31]/NET0131 ,
		\u6_wp_reg[0]/P0001 ,
		\u6_wp_reg[1]/NET0131 ,
		_w5404_
	);
	LUT4 #(
		.INIT('h0800)
	) name3258 (
		\u12_dout_reg[31]/P0001 ,
		\u12_o7_we_reg/P0001 ,
		\u6_wp_reg[0]/P0001 ,
		\u6_wp_reg[1]/NET0131 ,
		_w5405_
	);
	LUT2 #(
		.INIT('he)
	) name3259 (
		_w5404_,
		_w5405_,
		_w5406_
	);
	LUT4 #(
		.INIT('hc4cc)
	) name3260 (
		\u12_o7_we_reg/P0001 ,
		\u6_mem_reg[2][3]/NET0131 ,
		\u6_wp_reg[0]/P0001 ,
		\u6_wp_reg[1]/NET0131 ,
		_w5407_
	);
	LUT4 #(
		.INIT('h0800)
	) name3261 (
		\u12_dout_reg[3]/P0001 ,
		\u12_o7_we_reg/P0001 ,
		\u6_wp_reg[0]/P0001 ,
		\u6_wp_reg[1]/NET0131 ,
		_w5408_
	);
	LUT2 #(
		.INIT('he)
	) name3262 (
		_w5407_,
		_w5408_,
		_w5409_
	);
	LUT4 #(
		.INIT('hc4cc)
	) name3263 (
		\u12_o7_we_reg/P0001 ,
		\u6_mem_reg[2][4]/NET0131 ,
		\u6_wp_reg[0]/P0001 ,
		\u6_wp_reg[1]/NET0131 ,
		_w5410_
	);
	LUT4 #(
		.INIT('h0800)
	) name3264 (
		\u12_dout_reg[4]/P0001 ,
		\u12_o7_we_reg/P0001 ,
		\u6_wp_reg[0]/P0001 ,
		\u6_wp_reg[1]/NET0131 ,
		_w5411_
	);
	LUT2 #(
		.INIT('he)
	) name3265 (
		_w5410_,
		_w5411_,
		_w5412_
	);
	LUT4 #(
		.INIT('hc4cc)
	) name3266 (
		\u12_o7_we_reg/P0001 ,
		\u6_mem_reg[2][5]/NET0131 ,
		\u6_wp_reg[0]/P0001 ,
		\u6_wp_reg[1]/NET0131 ,
		_w5413_
	);
	LUT4 #(
		.INIT('h0800)
	) name3267 (
		\u12_dout_reg[5]/P0001 ,
		\u12_o7_we_reg/P0001 ,
		\u6_wp_reg[0]/P0001 ,
		\u6_wp_reg[1]/NET0131 ,
		_w5414_
	);
	LUT2 #(
		.INIT('he)
	) name3268 (
		_w5413_,
		_w5414_,
		_w5415_
	);
	LUT4 #(
		.INIT('hc4cc)
	) name3269 (
		\u12_o7_we_reg/P0001 ,
		\u6_mem_reg[2][6]/NET0131 ,
		\u6_wp_reg[0]/P0001 ,
		\u6_wp_reg[1]/NET0131 ,
		_w5416_
	);
	LUT4 #(
		.INIT('h0800)
	) name3270 (
		\u12_dout_reg[6]/P0001 ,
		\u12_o7_we_reg/P0001 ,
		\u6_wp_reg[0]/P0001 ,
		\u6_wp_reg[1]/NET0131 ,
		_w5417_
	);
	LUT2 #(
		.INIT('he)
	) name3271 (
		_w5416_,
		_w5417_,
		_w5418_
	);
	LUT4 #(
		.INIT('hc4cc)
	) name3272 (
		\u12_o7_we_reg/P0001 ,
		\u6_mem_reg[2][7]/NET0131 ,
		\u6_wp_reg[0]/P0001 ,
		\u6_wp_reg[1]/NET0131 ,
		_w5419_
	);
	LUT4 #(
		.INIT('h0800)
	) name3273 (
		\u12_dout_reg[7]/P0001 ,
		\u12_o7_we_reg/P0001 ,
		\u6_wp_reg[0]/P0001 ,
		\u6_wp_reg[1]/NET0131 ,
		_w5420_
	);
	LUT2 #(
		.INIT('he)
	) name3274 (
		_w5419_,
		_w5420_,
		_w5421_
	);
	LUT4 #(
		.INIT('hc4cc)
	) name3275 (
		\u12_o7_we_reg/P0001 ,
		\u6_mem_reg[2][8]/NET0131 ,
		\u6_wp_reg[0]/P0001 ,
		\u6_wp_reg[1]/NET0131 ,
		_w5422_
	);
	LUT4 #(
		.INIT('h0800)
	) name3276 (
		\u12_dout_reg[8]/P0001 ,
		\u12_o7_we_reg/P0001 ,
		\u6_wp_reg[0]/P0001 ,
		\u6_wp_reg[1]/NET0131 ,
		_w5423_
	);
	LUT2 #(
		.INIT('he)
	) name3277 (
		_w5422_,
		_w5423_,
		_w5424_
	);
	LUT4 #(
		.INIT('hc4cc)
	) name3278 (
		\u12_o7_we_reg/P0001 ,
		\u6_mem_reg[2][9]/NET0131 ,
		\u6_wp_reg[0]/P0001 ,
		\u6_wp_reg[1]/NET0131 ,
		_w5425_
	);
	LUT4 #(
		.INIT('h0800)
	) name3279 (
		\u12_dout_reg[9]/P0001 ,
		\u12_o7_we_reg/P0001 ,
		\u6_wp_reg[0]/P0001 ,
		\u6_wp_reg[1]/NET0131 ,
		_w5426_
	);
	LUT2 #(
		.INIT('he)
	) name3280 (
		_w5425_,
		_w5426_,
		_w5427_
	);
	LUT4 #(
		.INIT('h4ccc)
	) name3281 (
		\u12_o7_we_reg/P0001 ,
		\u6_mem_reg[3][0]/NET0131 ,
		\u6_wp_reg[0]/P0001 ,
		\u6_wp_reg[1]/NET0131 ,
		_w5428_
	);
	LUT4 #(
		.INIT('h8000)
	) name3282 (
		\u12_dout_reg[0]/P0001 ,
		\u12_o7_we_reg/P0001 ,
		\u6_wp_reg[0]/P0001 ,
		\u6_wp_reg[1]/NET0131 ,
		_w5429_
	);
	LUT2 #(
		.INIT('he)
	) name3283 (
		_w5428_,
		_w5429_,
		_w5430_
	);
	LUT4 #(
		.INIT('h4ccc)
	) name3284 (
		\u12_o7_we_reg/P0001 ,
		\u6_mem_reg[3][10]/NET0131 ,
		\u6_wp_reg[0]/P0001 ,
		\u6_wp_reg[1]/NET0131 ,
		_w5431_
	);
	LUT4 #(
		.INIT('h8000)
	) name3285 (
		\u12_dout_reg[10]/P0001 ,
		\u12_o7_we_reg/P0001 ,
		\u6_wp_reg[0]/P0001 ,
		\u6_wp_reg[1]/NET0131 ,
		_w5432_
	);
	LUT2 #(
		.INIT('he)
	) name3286 (
		_w5431_,
		_w5432_,
		_w5433_
	);
	LUT4 #(
		.INIT('h4ccc)
	) name3287 (
		\u12_o7_we_reg/P0001 ,
		\u6_mem_reg[3][11]/NET0131 ,
		\u6_wp_reg[0]/P0001 ,
		\u6_wp_reg[1]/NET0131 ,
		_w5434_
	);
	LUT4 #(
		.INIT('h8000)
	) name3288 (
		\u12_dout_reg[11]/P0001 ,
		\u12_o7_we_reg/P0001 ,
		\u6_wp_reg[0]/P0001 ,
		\u6_wp_reg[1]/NET0131 ,
		_w5435_
	);
	LUT2 #(
		.INIT('he)
	) name3289 (
		_w5434_,
		_w5435_,
		_w5436_
	);
	LUT4 #(
		.INIT('h4ccc)
	) name3290 (
		\u12_o7_we_reg/P0001 ,
		\u6_mem_reg[3][12]/NET0131 ,
		\u6_wp_reg[0]/P0001 ,
		\u6_wp_reg[1]/NET0131 ,
		_w5437_
	);
	LUT4 #(
		.INIT('h8000)
	) name3291 (
		\u12_dout_reg[12]/P0001 ,
		\u12_o7_we_reg/P0001 ,
		\u6_wp_reg[0]/P0001 ,
		\u6_wp_reg[1]/NET0131 ,
		_w5438_
	);
	LUT2 #(
		.INIT('he)
	) name3292 (
		_w5437_,
		_w5438_,
		_w5439_
	);
	LUT4 #(
		.INIT('h4ccc)
	) name3293 (
		\u12_o7_we_reg/P0001 ,
		\u6_mem_reg[3][13]/NET0131 ,
		\u6_wp_reg[0]/P0001 ,
		\u6_wp_reg[1]/NET0131 ,
		_w5440_
	);
	LUT4 #(
		.INIT('h8000)
	) name3294 (
		\u12_dout_reg[13]/P0001 ,
		\u12_o7_we_reg/P0001 ,
		\u6_wp_reg[0]/P0001 ,
		\u6_wp_reg[1]/NET0131 ,
		_w5441_
	);
	LUT2 #(
		.INIT('he)
	) name3295 (
		_w5440_,
		_w5441_,
		_w5442_
	);
	LUT4 #(
		.INIT('h4ccc)
	) name3296 (
		\u12_o7_we_reg/P0001 ,
		\u6_mem_reg[3][14]/NET0131 ,
		\u6_wp_reg[0]/P0001 ,
		\u6_wp_reg[1]/NET0131 ,
		_w5443_
	);
	LUT4 #(
		.INIT('h8000)
	) name3297 (
		\u12_dout_reg[14]/P0001 ,
		\u12_o7_we_reg/P0001 ,
		\u6_wp_reg[0]/P0001 ,
		\u6_wp_reg[1]/NET0131 ,
		_w5444_
	);
	LUT2 #(
		.INIT('he)
	) name3298 (
		_w5443_,
		_w5444_,
		_w5445_
	);
	LUT4 #(
		.INIT('h4ccc)
	) name3299 (
		\u12_o7_we_reg/P0001 ,
		\u6_mem_reg[3][15]/NET0131 ,
		\u6_wp_reg[0]/P0001 ,
		\u6_wp_reg[1]/NET0131 ,
		_w5446_
	);
	LUT4 #(
		.INIT('h8000)
	) name3300 (
		\u12_dout_reg[15]/P0001 ,
		\u12_o7_we_reg/P0001 ,
		\u6_wp_reg[0]/P0001 ,
		\u6_wp_reg[1]/NET0131 ,
		_w5447_
	);
	LUT2 #(
		.INIT('he)
	) name3301 (
		_w5446_,
		_w5447_,
		_w5448_
	);
	LUT4 #(
		.INIT('h4ccc)
	) name3302 (
		\u12_o7_we_reg/P0001 ,
		\u6_mem_reg[3][16]/NET0131 ,
		\u6_wp_reg[0]/P0001 ,
		\u6_wp_reg[1]/NET0131 ,
		_w5449_
	);
	LUT4 #(
		.INIT('h8000)
	) name3303 (
		\u12_dout_reg[16]/P0001 ,
		\u12_o7_we_reg/P0001 ,
		\u6_wp_reg[0]/P0001 ,
		\u6_wp_reg[1]/NET0131 ,
		_w5450_
	);
	LUT2 #(
		.INIT('he)
	) name3304 (
		_w5449_,
		_w5450_,
		_w5451_
	);
	LUT4 #(
		.INIT('h4ccc)
	) name3305 (
		\u12_o7_we_reg/P0001 ,
		\u6_mem_reg[3][17]/NET0131 ,
		\u6_wp_reg[0]/P0001 ,
		\u6_wp_reg[1]/NET0131 ,
		_w5452_
	);
	LUT4 #(
		.INIT('h8000)
	) name3306 (
		\u12_dout_reg[17]/P0001 ,
		\u12_o7_we_reg/P0001 ,
		\u6_wp_reg[0]/P0001 ,
		\u6_wp_reg[1]/NET0131 ,
		_w5453_
	);
	LUT2 #(
		.INIT('he)
	) name3307 (
		_w5452_,
		_w5453_,
		_w5454_
	);
	LUT4 #(
		.INIT('h4ccc)
	) name3308 (
		\u12_o7_we_reg/P0001 ,
		\u6_mem_reg[3][18]/NET0131 ,
		\u6_wp_reg[0]/P0001 ,
		\u6_wp_reg[1]/NET0131 ,
		_w5455_
	);
	LUT4 #(
		.INIT('h8000)
	) name3309 (
		\u12_dout_reg[18]/P0001 ,
		\u12_o7_we_reg/P0001 ,
		\u6_wp_reg[0]/P0001 ,
		\u6_wp_reg[1]/NET0131 ,
		_w5456_
	);
	LUT2 #(
		.INIT('he)
	) name3310 (
		_w5455_,
		_w5456_,
		_w5457_
	);
	LUT4 #(
		.INIT('h4ccc)
	) name3311 (
		\u12_o7_we_reg/P0001 ,
		\u6_mem_reg[3][19]/NET0131 ,
		\u6_wp_reg[0]/P0001 ,
		\u6_wp_reg[1]/NET0131 ,
		_w5458_
	);
	LUT4 #(
		.INIT('h8000)
	) name3312 (
		\u12_dout_reg[19]/P0001 ,
		\u12_o7_we_reg/P0001 ,
		\u6_wp_reg[0]/P0001 ,
		\u6_wp_reg[1]/NET0131 ,
		_w5459_
	);
	LUT2 #(
		.INIT('he)
	) name3313 (
		_w5458_,
		_w5459_,
		_w5460_
	);
	LUT4 #(
		.INIT('h4ccc)
	) name3314 (
		\u12_o7_we_reg/P0001 ,
		\u6_mem_reg[3][1]/NET0131 ,
		\u6_wp_reg[0]/P0001 ,
		\u6_wp_reg[1]/NET0131 ,
		_w5461_
	);
	LUT4 #(
		.INIT('h8000)
	) name3315 (
		\u12_dout_reg[1]/P0001 ,
		\u12_o7_we_reg/P0001 ,
		\u6_wp_reg[0]/P0001 ,
		\u6_wp_reg[1]/NET0131 ,
		_w5462_
	);
	LUT2 #(
		.INIT('he)
	) name3316 (
		_w5461_,
		_w5462_,
		_w5463_
	);
	LUT4 #(
		.INIT('h4ccc)
	) name3317 (
		\u12_o7_we_reg/P0001 ,
		\u6_mem_reg[3][20]/NET0131 ,
		\u6_wp_reg[0]/P0001 ,
		\u6_wp_reg[1]/NET0131 ,
		_w5464_
	);
	LUT4 #(
		.INIT('h8000)
	) name3318 (
		\u12_dout_reg[20]/P0001 ,
		\u12_o7_we_reg/P0001 ,
		\u6_wp_reg[0]/P0001 ,
		\u6_wp_reg[1]/NET0131 ,
		_w5465_
	);
	LUT2 #(
		.INIT('he)
	) name3319 (
		_w5464_,
		_w5465_,
		_w5466_
	);
	LUT4 #(
		.INIT('h4ccc)
	) name3320 (
		\u12_o7_we_reg/P0001 ,
		\u6_mem_reg[3][21]/NET0131 ,
		\u6_wp_reg[0]/P0001 ,
		\u6_wp_reg[1]/NET0131 ,
		_w5467_
	);
	LUT4 #(
		.INIT('h8000)
	) name3321 (
		\u12_dout_reg[21]/P0001 ,
		\u12_o7_we_reg/P0001 ,
		\u6_wp_reg[0]/P0001 ,
		\u6_wp_reg[1]/NET0131 ,
		_w5468_
	);
	LUT2 #(
		.INIT('he)
	) name3322 (
		_w5467_,
		_w5468_,
		_w5469_
	);
	LUT4 #(
		.INIT('h4ccc)
	) name3323 (
		\u12_o7_we_reg/P0001 ,
		\u6_mem_reg[3][22]/NET0131 ,
		\u6_wp_reg[0]/P0001 ,
		\u6_wp_reg[1]/NET0131 ,
		_w5470_
	);
	LUT4 #(
		.INIT('h8000)
	) name3324 (
		\u12_dout_reg[22]/P0001 ,
		\u12_o7_we_reg/P0001 ,
		\u6_wp_reg[0]/P0001 ,
		\u6_wp_reg[1]/NET0131 ,
		_w5471_
	);
	LUT2 #(
		.INIT('he)
	) name3325 (
		_w5470_,
		_w5471_,
		_w5472_
	);
	LUT4 #(
		.INIT('h4ccc)
	) name3326 (
		\u12_o7_we_reg/P0001 ,
		\u6_mem_reg[3][23]/NET0131 ,
		\u6_wp_reg[0]/P0001 ,
		\u6_wp_reg[1]/NET0131 ,
		_w5473_
	);
	LUT4 #(
		.INIT('h8000)
	) name3327 (
		\u12_dout_reg[23]/P0001 ,
		\u12_o7_we_reg/P0001 ,
		\u6_wp_reg[0]/P0001 ,
		\u6_wp_reg[1]/NET0131 ,
		_w5474_
	);
	LUT2 #(
		.INIT('he)
	) name3328 (
		_w5473_,
		_w5474_,
		_w5475_
	);
	LUT4 #(
		.INIT('h4ccc)
	) name3329 (
		\u12_o7_we_reg/P0001 ,
		\u6_mem_reg[3][24]/NET0131 ,
		\u6_wp_reg[0]/P0001 ,
		\u6_wp_reg[1]/NET0131 ,
		_w5476_
	);
	LUT4 #(
		.INIT('h8000)
	) name3330 (
		\u12_dout_reg[24]/P0001 ,
		\u12_o7_we_reg/P0001 ,
		\u6_wp_reg[0]/P0001 ,
		\u6_wp_reg[1]/NET0131 ,
		_w5477_
	);
	LUT2 #(
		.INIT('he)
	) name3331 (
		_w5476_,
		_w5477_,
		_w5478_
	);
	LUT4 #(
		.INIT('h4ccc)
	) name3332 (
		\u12_o7_we_reg/P0001 ,
		\u6_mem_reg[3][25]/NET0131 ,
		\u6_wp_reg[0]/P0001 ,
		\u6_wp_reg[1]/NET0131 ,
		_w5479_
	);
	LUT4 #(
		.INIT('h8000)
	) name3333 (
		\u12_dout_reg[25]/P0001 ,
		\u12_o7_we_reg/P0001 ,
		\u6_wp_reg[0]/P0001 ,
		\u6_wp_reg[1]/NET0131 ,
		_w5480_
	);
	LUT2 #(
		.INIT('he)
	) name3334 (
		_w5479_,
		_w5480_,
		_w5481_
	);
	LUT4 #(
		.INIT('h4ccc)
	) name3335 (
		\u12_o7_we_reg/P0001 ,
		\u6_mem_reg[3][26]/NET0131 ,
		\u6_wp_reg[0]/P0001 ,
		\u6_wp_reg[1]/NET0131 ,
		_w5482_
	);
	LUT4 #(
		.INIT('h8000)
	) name3336 (
		\u12_dout_reg[26]/P0001 ,
		\u12_o7_we_reg/P0001 ,
		\u6_wp_reg[0]/P0001 ,
		\u6_wp_reg[1]/NET0131 ,
		_w5483_
	);
	LUT2 #(
		.INIT('he)
	) name3337 (
		_w5482_,
		_w5483_,
		_w5484_
	);
	LUT4 #(
		.INIT('h4ccc)
	) name3338 (
		\u12_o7_we_reg/P0001 ,
		\u6_mem_reg[3][27]/NET0131 ,
		\u6_wp_reg[0]/P0001 ,
		\u6_wp_reg[1]/NET0131 ,
		_w5485_
	);
	LUT4 #(
		.INIT('h8000)
	) name3339 (
		\u12_dout_reg[27]/P0001 ,
		\u12_o7_we_reg/P0001 ,
		\u6_wp_reg[0]/P0001 ,
		\u6_wp_reg[1]/NET0131 ,
		_w5486_
	);
	LUT2 #(
		.INIT('he)
	) name3340 (
		_w5485_,
		_w5486_,
		_w5487_
	);
	LUT4 #(
		.INIT('h4ccc)
	) name3341 (
		\u12_o7_we_reg/P0001 ,
		\u6_mem_reg[3][28]/NET0131 ,
		\u6_wp_reg[0]/P0001 ,
		\u6_wp_reg[1]/NET0131 ,
		_w5488_
	);
	LUT4 #(
		.INIT('h8000)
	) name3342 (
		\u12_dout_reg[28]/P0001 ,
		\u12_o7_we_reg/P0001 ,
		\u6_wp_reg[0]/P0001 ,
		\u6_wp_reg[1]/NET0131 ,
		_w5489_
	);
	LUT2 #(
		.INIT('he)
	) name3343 (
		_w5488_,
		_w5489_,
		_w5490_
	);
	LUT4 #(
		.INIT('h4ccc)
	) name3344 (
		\u12_o7_we_reg/P0001 ,
		\u6_mem_reg[3][29]/NET0131 ,
		\u6_wp_reg[0]/P0001 ,
		\u6_wp_reg[1]/NET0131 ,
		_w5491_
	);
	LUT4 #(
		.INIT('h8000)
	) name3345 (
		\u12_dout_reg[29]/P0001 ,
		\u12_o7_we_reg/P0001 ,
		\u6_wp_reg[0]/P0001 ,
		\u6_wp_reg[1]/NET0131 ,
		_w5492_
	);
	LUT2 #(
		.INIT('he)
	) name3346 (
		_w5491_,
		_w5492_,
		_w5493_
	);
	LUT4 #(
		.INIT('h4ccc)
	) name3347 (
		\u12_o7_we_reg/P0001 ,
		\u6_mem_reg[3][2]/NET0131 ,
		\u6_wp_reg[0]/P0001 ,
		\u6_wp_reg[1]/NET0131 ,
		_w5494_
	);
	LUT4 #(
		.INIT('h8000)
	) name3348 (
		\u12_dout_reg[2]/P0001 ,
		\u12_o7_we_reg/P0001 ,
		\u6_wp_reg[0]/P0001 ,
		\u6_wp_reg[1]/NET0131 ,
		_w5495_
	);
	LUT2 #(
		.INIT('he)
	) name3349 (
		_w5494_,
		_w5495_,
		_w5496_
	);
	LUT4 #(
		.INIT('h4ccc)
	) name3350 (
		\u12_o7_we_reg/P0001 ,
		\u6_mem_reg[3][30]/NET0131 ,
		\u6_wp_reg[0]/P0001 ,
		\u6_wp_reg[1]/NET0131 ,
		_w5497_
	);
	LUT4 #(
		.INIT('h8000)
	) name3351 (
		\u12_dout_reg[30]/P0001 ,
		\u12_o7_we_reg/P0001 ,
		\u6_wp_reg[0]/P0001 ,
		\u6_wp_reg[1]/NET0131 ,
		_w5498_
	);
	LUT2 #(
		.INIT('he)
	) name3352 (
		_w5497_,
		_w5498_,
		_w5499_
	);
	LUT4 #(
		.INIT('h4ccc)
	) name3353 (
		\u12_o7_we_reg/P0001 ,
		\u6_mem_reg[3][31]/NET0131 ,
		\u6_wp_reg[0]/P0001 ,
		\u6_wp_reg[1]/NET0131 ,
		_w5500_
	);
	LUT4 #(
		.INIT('h8000)
	) name3354 (
		\u12_dout_reg[31]/P0001 ,
		\u12_o7_we_reg/P0001 ,
		\u6_wp_reg[0]/P0001 ,
		\u6_wp_reg[1]/NET0131 ,
		_w5501_
	);
	LUT2 #(
		.INIT('he)
	) name3355 (
		_w5500_,
		_w5501_,
		_w5502_
	);
	LUT4 #(
		.INIT('h4ccc)
	) name3356 (
		\u12_o7_we_reg/P0001 ,
		\u6_mem_reg[3][3]/NET0131 ,
		\u6_wp_reg[0]/P0001 ,
		\u6_wp_reg[1]/NET0131 ,
		_w5503_
	);
	LUT4 #(
		.INIT('h8000)
	) name3357 (
		\u12_dout_reg[3]/P0001 ,
		\u12_o7_we_reg/P0001 ,
		\u6_wp_reg[0]/P0001 ,
		\u6_wp_reg[1]/NET0131 ,
		_w5504_
	);
	LUT2 #(
		.INIT('he)
	) name3358 (
		_w5503_,
		_w5504_,
		_w5505_
	);
	LUT4 #(
		.INIT('h4ccc)
	) name3359 (
		\u12_o7_we_reg/P0001 ,
		\u6_mem_reg[3][4]/NET0131 ,
		\u6_wp_reg[0]/P0001 ,
		\u6_wp_reg[1]/NET0131 ,
		_w5506_
	);
	LUT4 #(
		.INIT('h8000)
	) name3360 (
		\u12_dout_reg[4]/P0001 ,
		\u12_o7_we_reg/P0001 ,
		\u6_wp_reg[0]/P0001 ,
		\u6_wp_reg[1]/NET0131 ,
		_w5507_
	);
	LUT2 #(
		.INIT('he)
	) name3361 (
		_w5506_,
		_w5507_,
		_w5508_
	);
	LUT4 #(
		.INIT('h4ccc)
	) name3362 (
		\u12_o7_we_reg/P0001 ,
		\u6_mem_reg[3][5]/NET0131 ,
		\u6_wp_reg[0]/P0001 ,
		\u6_wp_reg[1]/NET0131 ,
		_w5509_
	);
	LUT4 #(
		.INIT('h8000)
	) name3363 (
		\u12_dout_reg[5]/P0001 ,
		\u12_o7_we_reg/P0001 ,
		\u6_wp_reg[0]/P0001 ,
		\u6_wp_reg[1]/NET0131 ,
		_w5510_
	);
	LUT2 #(
		.INIT('he)
	) name3364 (
		_w5509_,
		_w5510_,
		_w5511_
	);
	LUT4 #(
		.INIT('h4ccc)
	) name3365 (
		\u12_o7_we_reg/P0001 ,
		\u6_mem_reg[3][6]/NET0131 ,
		\u6_wp_reg[0]/P0001 ,
		\u6_wp_reg[1]/NET0131 ,
		_w5512_
	);
	LUT4 #(
		.INIT('h8000)
	) name3366 (
		\u12_dout_reg[6]/P0001 ,
		\u12_o7_we_reg/P0001 ,
		\u6_wp_reg[0]/P0001 ,
		\u6_wp_reg[1]/NET0131 ,
		_w5513_
	);
	LUT2 #(
		.INIT('he)
	) name3367 (
		_w5512_,
		_w5513_,
		_w5514_
	);
	LUT4 #(
		.INIT('h4ccc)
	) name3368 (
		\u12_o7_we_reg/P0001 ,
		\u6_mem_reg[3][7]/NET0131 ,
		\u6_wp_reg[0]/P0001 ,
		\u6_wp_reg[1]/NET0131 ,
		_w5515_
	);
	LUT4 #(
		.INIT('h8000)
	) name3369 (
		\u12_dout_reg[7]/P0001 ,
		\u12_o7_we_reg/P0001 ,
		\u6_wp_reg[0]/P0001 ,
		\u6_wp_reg[1]/NET0131 ,
		_w5516_
	);
	LUT2 #(
		.INIT('he)
	) name3370 (
		_w5515_,
		_w5516_,
		_w5517_
	);
	LUT4 #(
		.INIT('h4ccc)
	) name3371 (
		\u12_o7_we_reg/P0001 ,
		\u6_mem_reg[3][8]/NET0131 ,
		\u6_wp_reg[0]/P0001 ,
		\u6_wp_reg[1]/NET0131 ,
		_w5518_
	);
	LUT4 #(
		.INIT('h8000)
	) name3372 (
		\u12_dout_reg[8]/P0001 ,
		\u12_o7_we_reg/P0001 ,
		\u6_wp_reg[0]/P0001 ,
		\u6_wp_reg[1]/NET0131 ,
		_w5519_
	);
	LUT2 #(
		.INIT('he)
	) name3373 (
		_w5518_,
		_w5519_,
		_w5520_
	);
	LUT4 #(
		.INIT('h4ccc)
	) name3374 (
		\u12_o7_we_reg/P0001 ,
		\u6_mem_reg[3][9]/NET0131 ,
		\u6_wp_reg[0]/P0001 ,
		\u6_wp_reg[1]/NET0131 ,
		_w5521_
	);
	LUT4 #(
		.INIT('h8000)
	) name3375 (
		\u12_dout_reg[9]/P0001 ,
		\u12_o7_we_reg/P0001 ,
		\u6_wp_reg[0]/P0001 ,
		\u6_wp_reg[1]/NET0131 ,
		_w5522_
	);
	LUT2 #(
		.INIT('he)
	) name3376 (
		_w5521_,
		_w5522_,
		_w5523_
	);
	LUT4 #(
		.INIT('hcc4c)
	) name3377 (
		\u12_o9_we_reg/P0001 ,
		\u8_mem_reg[1][6]/NET0131 ,
		\u8_wp_reg[0]/P0001 ,
		\u8_wp_reg[1]/NET0131 ,
		_w5524_
	);
	LUT4 #(
		.INIT('h0080)
	) name3378 (
		\u12_dout_reg[6]/P0001 ,
		\u12_o9_we_reg/P0001 ,
		\u8_wp_reg[0]/P0001 ,
		\u8_wp_reg[1]/NET0131 ,
		_w5525_
	);
	LUT2 #(
		.INIT('he)
	) name3379 (
		_w5524_,
		_w5525_,
		_w5526_
	);
	LUT4 #(
		.INIT('hc4cc)
	) name3380 (
		\u12_o3_we_reg/P0001 ,
		\u3_mem_reg[2][25]/NET0131 ,
		\u3_wp_reg[0]/P0001 ,
		\u3_wp_reg[1]/NET0131 ,
		_w5527_
	);
	LUT4 #(
		.INIT('h0800)
	) name3381 (
		\u12_dout_reg[25]/P0001 ,
		\u12_o3_we_reg/P0001 ,
		\u3_wp_reg[0]/P0001 ,
		\u3_wp_reg[1]/NET0131 ,
		_w5528_
	);
	LUT2 #(
		.INIT('he)
	) name3382 (
		_w5527_,
		_w5528_,
		_w5529_
	);
	LUT4 #(
		.INIT('h4ccc)
	) name3383 (
		\u12_o9_we_reg/P0001 ,
		\u8_mem_reg[3][4]/NET0131 ,
		\u8_wp_reg[0]/P0001 ,
		\u8_wp_reg[1]/NET0131 ,
		_w5530_
	);
	LUT4 #(
		.INIT('h8000)
	) name3384 (
		\u12_dout_reg[4]/P0001 ,
		\u12_o9_we_reg/P0001 ,
		\u8_wp_reg[0]/P0001 ,
		\u8_wp_reg[1]/NET0131 ,
		_w5531_
	);
	LUT2 #(
		.INIT('he)
	) name3385 (
		_w5530_,
		_w5531_,
		_w5532_
	);
	LUT4 #(
		.INIT('h4ccc)
	) name3386 (
		\u12_o3_we_reg/P0001 ,
		\u3_mem_reg[3][3]/NET0131 ,
		\u3_wp_reg[0]/P0001 ,
		\u3_wp_reg[1]/NET0131 ,
		_w5533_
	);
	LUT4 #(
		.INIT('h8000)
	) name3387 (
		\u12_dout_reg[3]/P0001 ,
		\u12_o3_we_reg/P0001 ,
		\u3_wp_reg[0]/P0001 ,
		\u3_wp_reg[1]/NET0131 ,
		_w5534_
	);
	LUT2 #(
		.INIT('he)
	) name3388 (
		_w5533_,
		_w5534_,
		_w5535_
	);
	LUT4 #(
		.INIT('h4ccc)
	) name3389 (
		\u12_o9_we_reg/P0001 ,
		\u8_mem_reg[3][8]/NET0131 ,
		\u8_wp_reg[0]/P0001 ,
		\u8_wp_reg[1]/NET0131 ,
		_w5536_
	);
	LUT4 #(
		.INIT('h8000)
	) name3390 (
		\u12_dout_reg[8]/P0001 ,
		\u12_o9_we_reg/P0001 ,
		\u8_wp_reg[0]/P0001 ,
		\u8_wp_reg[1]/NET0131 ,
		_w5537_
	);
	LUT2 #(
		.INIT('he)
	) name3391 (
		_w5536_,
		_w5537_,
		_w5538_
	);
	LUT4 #(
		.INIT('hcc4c)
	) name3392 (
		\u12_o3_we_reg/P0001 ,
		\u3_mem_reg[1][14]/NET0131 ,
		\u3_wp_reg[0]/P0001 ,
		\u3_wp_reg[1]/NET0131 ,
		_w5539_
	);
	LUT4 #(
		.INIT('h0080)
	) name3393 (
		\u12_dout_reg[14]/P0001 ,
		\u12_o3_we_reg/P0001 ,
		\u3_wp_reg[0]/P0001 ,
		\u3_wp_reg[1]/NET0131 ,
		_w5540_
	);
	LUT2 #(
		.INIT('he)
	) name3394 (
		_w5539_,
		_w5540_,
		_w5541_
	);
	LUT4 #(
		.INIT('hcc4c)
	) name3395 (
		\u12_o8_we_reg/P0001 ,
		\u7_mem_reg[1][0]/NET0131 ,
		\u7_wp_reg[0]/P0001 ,
		\u7_wp_reg[1]/NET0131 ,
		_w5542_
	);
	LUT4 #(
		.INIT('h0080)
	) name3396 (
		\u12_dout_reg[0]/P0001 ,
		\u12_o8_we_reg/P0001 ,
		\u7_wp_reg[0]/P0001 ,
		\u7_wp_reg[1]/NET0131 ,
		_w5543_
	);
	LUT2 #(
		.INIT('he)
	) name3397 (
		_w5542_,
		_w5543_,
		_w5544_
	);
	LUT4 #(
		.INIT('hcc4c)
	) name3398 (
		\u12_o8_we_reg/P0001 ,
		\u7_mem_reg[1][10]/NET0131 ,
		\u7_wp_reg[0]/P0001 ,
		\u7_wp_reg[1]/NET0131 ,
		_w5545_
	);
	LUT4 #(
		.INIT('h0080)
	) name3399 (
		\u12_dout_reg[10]/P0001 ,
		\u12_o8_we_reg/P0001 ,
		\u7_wp_reg[0]/P0001 ,
		\u7_wp_reg[1]/NET0131 ,
		_w5546_
	);
	LUT2 #(
		.INIT('he)
	) name3400 (
		_w5545_,
		_w5546_,
		_w5547_
	);
	LUT4 #(
		.INIT('hcc4c)
	) name3401 (
		\u12_o8_we_reg/P0001 ,
		\u7_mem_reg[1][11]/NET0131 ,
		\u7_wp_reg[0]/P0001 ,
		\u7_wp_reg[1]/NET0131 ,
		_w5548_
	);
	LUT4 #(
		.INIT('h0080)
	) name3402 (
		\u12_dout_reg[11]/P0001 ,
		\u12_o8_we_reg/P0001 ,
		\u7_wp_reg[0]/P0001 ,
		\u7_wp_reg[1]/NET0131 ,
		_w5549_
	);
	LUT2 #(
		.INIT('he)
	) name3403 (
		_w5548_,
		_w5549_,
		_w5550_
	);
	LUT4 #(
		.INIT('hcc4c)
	) name3404 (
		\u12_o3_we_reg/P0001 ,
		\u3_mem_reg[1][23]/NET0131 ,
		\u3_wp_reg[0]/P0001 ,
		\u3_wp_reg[1]/NET0131 ,
		_w5551_
	);
	LUT4 #(
		.INIT('h0080)
	) name3405 (
		\u12_dout_reg[23]/P0001 ,
		\u12_o3_we_reg/P0001 ,
		\u3_wp_reg[0]/P0001 ,
		\u3_wp_reg[1]/NET0131 ,
		_w5552_
	);
	LUT2 #(
		.INIT('he)
	) name3406 (
		_w5551_,
		_w5552_,
		_w5553_
	);
	LUT4 #(
		.INIT('hcc4c)
	) name3407 (
		\u12_o8_we_reg/P0001 ,
		\u7_mem_reg[1][12]/NET0131 ,
		\u7_wp_reg[0]/P0001 ,
		\u7_wp_reg[1]/NET0131 ,
		_w5554_
	);
	LUT4 #(
		.INIT('h0080)
	) name3408 (
		\u12_dout_reg[12]/P0001 ,
		\u12_o8_we_reg/P0001 ,
		\u7_wp_reg[0]/P0001 ,
		\u7_wp_reg[1]/NET0131 ,
		_w5555_
	);
	LUT2 #(
		.INIT('he)
	) name3409 (
		_w5554_,
		_w5555_,
		_w5556_
	);
	LUT4 #(
		.INIT('hcc4c)
	) name3410 (
		\u12_o8_we_reg/P0001 ,
		\u7_mem_reg[1][13]/NET0131 ,
		\u7_wp_reg[0]/P0001 ,
		\u7_wp_reg[1]/NET0131 ,
		_w5557_
	);
	LUT4 #(
		.INIT('h0080)
	) name3411 (
		\u12_dout_reg[13]/P0001 ,
		\u12_o8_we_reg/P0001 ,
		\u7_wp_reg[0]/P0001 ,
		\u7_wp_reg[1]/NET0131 ,
		_w5558_
	);
	LUT2 #(
		.INIT('he)
	) name3412 (
		_w5557_,
		_w5558_,
		_w5559_
	);
	LUT4 #(
		.INIT('hcc4c)
	) name3413 (
		\u12_o8_we_reg/P0001 ,
		\u7_mem_reg[1][14]/NET0131 ,
		\u7_wp_reg[0]/P0001 ,
		\u7_wp_reg[1]/NET0131 ,
		_w5560_
	);
	LUT4 #(
		.INIT('h0080)
	) name3414 (
		\u12_dout_reg[14]/P0001 ,
		\u12_o8_we_reg/P0001 ,
		\u7_wp_reg[0]/P0001 ,
		\u7_wp_reg[1]/NET0131 ,
		_w5561_
	);
	LUT2 #(
		.INIT('he)
	) name3415 (
		_w5560_,
		_w5561_,
		_w5562_
	);
	LUT4 #(
		.INIT('hcc4c)
	) name3416 (
		\u12_o8_we_reg/P0001 ,
		\u7_mem_reg[1][15]/NET0131 ,
		\u7_wp_reg[0]/P0001 ,
		\u7_wp_reg[1]/NET0131 ,
		_w5563_
	);
	LUT4 #(
		.INIT('h0080)
	) name3417 (
		\u12_dout_reg[15]/P0001 ,
		\u12_o8_we_reg/P0001 ,
		\u7_wp_reg[0]/P0001 ,
		\u7_wp_reg[1]/NET0131 ,
		_w5564_
	);
	LUT2 #(
		.INIT('he)
	) name3418 (
		_w5563_,
		_w5564_,
		_w5565_
	);
	LUT4 #(
		.INIT('hcc4c)
	) name3419 (
		\u12_o8_we_reg/P0001 ,
		\u7_mem_reg[1][16]/NET0131 ,
		\u7_wp_reg[0]/P0001 ,
		\u7_wp_reg[1]/NET0131 ,
		_w5566_
	);
	LUT4 #(
		.INIT('h0080)
	) name3420 (
		\u12_dout_reg[16]/P0001 ,
		\u12_o8_we_reg/P0001 ,
		\u7_wp_reg[0]/P0001 ,
		\u7_wp_reg[1]/NET0131 ,
		_w5567_
	);
	LUT2 #(
		.INIT('he)
	) name3421 (
		_w5566_,
		_w5567_,
		_w5568_
	);
	LUT4 #(
		.INIT('hcc4c)
	) name3422 (
		\u12_o8_we_reg/P0001 ,
		\u7_mem_reg[1][17]/NET0131 ,
		\u7_wp_reg[0]/P0001 ,
		\u7_wp_reg[1]/NET0131 ,
		_w5569_
	);
	LUT4 #(
		.INIT('h0080)
	) name3423 (
		\u12_dout_reg[17]/P0001 ,
		\u12_o8_we_reg/P0001 ,
		\u7_wp_reg[0]/P0001 ,
		\u7_wp_reg[1]/NET0131 ,
		_w5570_
	);
	LUT2 #(
		.INIT('he)
	) name3424 (
		_w5569_,
		_w5570_,
		_w5571_
	);
	LUT4 #(
		.INIT('hcc4c)
	) name3425 (
		\u12_o8_we_reg/P0001 ,
		\u7_mem_reg[1][18]/NET0131 ,
		\u7_wp_reg[0]/P0001 ,
		\u7_wp_reg[1]/NET0131 ,
		_w5572_
	);
	LUT4 #(
		.INIT('h0080)
	) name3426 (
		\u12_dout_reg[18]/P0001 ,
		\u12_o8_we_reg/P0001 ,
		\u7_wp_reg[0]/P0001 ,
		\u7_wp_reg[1]/NET0131 ,
		_w5573_
	);
	LUT2 #(
		.INIT('he)
	) name3427 (
		_w5572_,
		_w5573_,
		_w5574_
	);
	LUT4 #(
		.INIT('hcc4c)
	) name3428 (
		\u12_o8_we_reg/P0001 ,
		\u7_mem_reg[1][19]/NET0131 ,
		\u7_wp_reg[0]/P0001 ,
		\u7_wp_reg[1]/NET0131 ,
		_w5575_
	);
	LUT4 #(
		.INIT('h0080)
	) name3429 (
		\u12_dout_reg[19]/P0001 ,
		\u12_o8_we_reg/P0001 ,
		\u7_wp_reg[0]/P0001 ,
		\u7_wp_reg[1]/NET0131 ,
		_w5576_
	);
	LUT2 #(
		.INIT('he)
	) name3430 (
		_w5575_,
		_w5576_,
		_w5577_
	);
	LUT4 #(
		.INIT('hcc4c)
	) name3431 (
		\u12_o8_we_reg/P0001 ,
		\u7_mem_reg[1][1]/NET0131 ,
		\u7_wp_reg[0]/P0001 ,
		\u7_wp_reg[1]/NET0131 ,
		_w5578_
	);
	LUT4 #(
		.INIT('h0080)
	) name3432 (
		\u12_dout_reg[1]/P0001 ,
		\u12_o8_we_reg/P0001 ,
		\u7_wp_reg[0]/P0001 ,
		\u7_wp_reg[1]/NET0131 ,
		_w5579_
	);
	LUT2 #(
		.INIT('he)
	) name3433 (
		_w5578_,
		_w5579_,
		_w5580_
	);
	LUT4 #(
		.INIT('hcc4c)
	) name3434 (
		\u12_o8_we_reg/P0001 ,
		\u7_mem_reg[1][20]/NET0131 ,
		\u7_wp_reg[0]/P0001 ,
		\u7_wp_reg[1]/NET0131 ,
		_w5581_
	);
	LUT4 #(
		.INIT('h0080)
	) name3435 (
		\u12_dout_reg[20]/P0001 ,
		\u12_o8_we_reg/P0001 ,
		\u7_wp_reg[0]/P0001 ,
		\u7_wp_reg[1]/NET0131 ,
		_w5582_
	);
	LUT2 #(
		.INIT('he)
	) name3436 (
		_w5581_,
		_w5582_,
		_w5583_
	);
	LUT4 #(
		.INIT('hcc4c)
	) name3437 (
		\u12_o8_we_reg/P0001 ,
		\u7_mem_reg[1][21]/NET0131 ,
		\u7_wp_reg[0]/P0001 ,
		\u7_wp_reg[1]/NET0131 ,
		_w5584_
	);
	LUT4 #(
		.INIT('h0080)
	) name3438 (
		\u12_dout_reg[21]/P0001 ,
		\u12_o8_we_reg/P0001 ,
		\u7_wp_reg[0]/P0001 ,
		\u7_wp_reg[1]/NET0131 ,
		_w5585_
	);
	LUT2 #(
		.INIT('he)
	) name3439 (
		_w5584_,
		_w5585_,
		_w5586_
	);
	LUT4 #(
		.INIT('hcc4c)
	) name3440 (
		\u12_o8_we_reg/P0001 ,
		\u7_mem_reg[1][22]/NET0131 ,
		\u7_wp_reg[0]/P0001 ,
		\u7_wp_reg[1]/NET0131 ,
		_w5587_
	);
	LUT4 #(
		.INIT('h0080)
	) name3441 (
		\u12_dout_reg[22]/P0001 ,
		\u12_o8_we_reg/P0001 ,
		\u7_wp_reg[0]/P0001 ,
		\u7_wp_reg[1]/NET0131 ,
		_w5588_
	);
	LUT2 #(
		.INIT('he)
	) name3442 (
		_w5587_,
		_w5588_,
		_w5589_
	);
	LUT4 #(
		.INIT('hcc4c)
	) name3443 (
		\u12_o8_we_reg/P0001 ,
		\u7_mem_reg[1][23]/NET0131 ,
		\u7_wp_reg[0]/P0001 ,
		\u7_wp_reg[1]/NET0131 ,
		_w5590_
	);
	LUT4 #(
		.INIT('h0080)
	) name3444 (
		\u12_dout_reg[23]/P0001 ,
		\u12_o8_we_reg/P0001 ,
		\u7_wp_reg[0]/P0001 ,
		\u7_wp_reg[1]/NET0131 ,
		_w5591_
	);
	LUT2 #(
		.INIT('he)
	) name3445 (
		_w5590_,
		_w5591_,
		_w5592_
	);
	LUT4 #(
		.INIT('hcc4c)
	) name3446 (
		\u12_o8_we_reg/P0001 ,
		\u7_mem_reg[1][24]/NET0131 ,
		\u7_wp_reg[0]/P0001 ,
		\u7_wp_reg[1]/NET0131 ,
		_w5593_
	);
	LUT4 #(
		.INIT('h0080)
	) name3447 (
		\u12_dout_reg[24]/P0001 ,
		\u12_o8_we_reg/P0001 ,
		\u7_wp_reg[0]/P0001 ,
		\u7_wp_reg[1]/NET0131 ,
		_w5594_
	);
	LUT2 #(
		.INIT('he)
	) name3448 (
		_w5593_,
		_w5594_,
		_w5595_
	);
	LUT4 #(
		.INIT('hcc4c)
	) name3449 (
		\u12_o8_we_reg/P0001 ,
		\u7_mem_reg[1][25]/NET0131 ,
		\u7_wp_reg[0]/P0001 ,
		\u7_wp_reg[1]/NET0131 ,
		_w5596_
	);
	LUT4 #(
		.INIT('h0080)
	) name3450 (
		\u12_dout_reg[25]/P0001 ,
		\u12_o8_we_reg/P0001 ,
		\u7_wp_reg[0]/P0001 ,
		\u7_wp_reg[1]/NET0131 ,
		_w5597_
	);
	LUT2 #(
		.INIT('he)
	) name3451 (
		_w5596_,
		_w5597_,
		_w5598_
	);
	LUT4 #(
		.INIT('hcc4c)
	) name3452 (
		\u12_o8_we_reg/P0001 ,
		\u7_mem_reg[1][26]/NET0131 ,
		\u7_wp_reg[0]/P0001 ,
		\u7_wp_reg[1]/NET0131 ,
		_w5599_
	);
	LUT4 #(
		.INIT('h0080)
	) name3453 (
		\u12_dout_reg[26]/P0001 ,
		\u12_o8_we_reg/P0001 ,
		\u7_wp_reg[0]/P0001 ,
		\u7_wp_reg[1]/NET0131 ,
		_w5600_
	);
	LUT2 #(
		.INIT('he)
	) name3454 (
		_w5599_,
		_w5600_,
		_w5601_
	);
	LUT4 #(
		.INIT('hcc4c)
	) name3455 (
		\u12_o8_we_reg/P0001 ,
		\u7_mem_reg[1][27]/NET0131 ,
		\u7_wp_reg[0]/P0001 ,
		\u7_wp_reg[1]/NET0131 ,
		_w5602_
	);
	LUT4 #(
		.INIT('h0080)
	) name3456 (
		\u12_dout_reg[27]/P0001 ,
		\u12_o8_we_reg/P0001 ,
		\u7_wp_reg[0]/P0001 ,
		\u7_wp_reg[1]/NET0131 ,
		_w5603_
	);
	LUT2 #(
		.INIT('he)
	) name3457 (
		_w5602_,
		_w5603_,
		_w5604_
	);
	LUT4 #(
		.INIT('hcc4c)
	) name3458 (
		\u12_o8_we_reg/P0001 ,
		\u7_mem_reg[1][28]/NET0131 ,
		\u7_wp_reg[0]/P0001 ,
		\u7_wp_reg[1]/NET0131 ,
		_w5605_
	);
	LUT4 #(
		.INIT('h0080)
	) name3459 (
		\u12_dout_reg[28]/P0001 ,
		\u12_o8_we_reg/P0001 ,
		\u7_wp_reg[0]/P0001 ,
		\u7_wp_reg[1]/NET0131 ,
		_w5606_
	);
	LUT2 #(
		.INIT('he)
	) name3460 (
		_w5605_,
		_w5606_,
		_w5607_
	);
	LUT4 #(
		.INIT('hcc4c)
	) name3461 (
		\u12_o8_we_reg/P0001 ,
		\u7_mem_reg[1][29]/NET0131 ,
		\u7_wp_reg[0]/P0001 ,
		\u7_wp_reg[1]/NET0131 ,
		_w5608_
	);
	LUT4 #(
		.INIT('h0080)
	) name3462 (
		\u12_dout_reg[29]/P0001 ,
		\u12_o8_we_reg/P0001 ,
		\u7_wp_reg[0]/P0001 ,
		\u7_wp_reg[1]/NET0131 ,
		_w5609_
	);
	LUT2 #(
		.INIT('he)
	) name3463 (
		_w5608_,
		_w5609_,
		_w5610_
	);
	LUT4 #(
		.INIT('hcc4c)
	) name3464 (
		\u12_o8_we_reg/P0001 ,
		\u7_mem_reg[1][2]/NET0131 ,
		\u7_wp_reg[0]/P0001 ,
		\u7_wp_reg[1]/NET0131 ,
		_w5611_
	);
	LUT4 #(
		.INIT('h0080)
	) name3465 (
		\u12_dout_reg[2]/P0001 ,
		\u12_o8_we_reg/P0001 ,
		\u7_wp_reg[0]/P0001 ,
		\u7_wp_reg[1]/NET0131 ,
		_w5612_
	);
	LUT2 #(
		.INIT('he)
	) name3466 (
		_w5611_,
		_w5612_,
		_w5613_
	);
	LUT4 #(
		.INIT('hcc4c)
	) name3467 (
		\u12_o8_we_reg/P0001 ,
		\u7_mem_reg[1][30]/NET0131 ,
		\u7_wp_reg[0]/P0001 ,
		\u7_wp_reg[1]/NET0131 ,
		_w5614_
	);
	LUT4 #(
		.INIT('h0080)
	) name3468 (
		\u12_dout_reg[30]/P0001 ,
		\u12_o8_we_reg/P0001 ,
		\u7_wp_reg[0]/P0001 ,
		\u7_wp_reg[1]/NET0131 ,
		_w5615_
	);
	LUT2 #(
		.INIT('he)
	) name3469 (
		_w5614_,
		_w5615_,
		_w5616_
	);
	LUT4 #(
		.INIT('hcc4c)
	) name3470 (
		\u12_o8_we_reg/P0001 ,
		\u7_mem_reg[1][31]/NET0131 ,
		\u7_wp_reg[0]/P0001 ,
		\u7_wp_reg[1]/NET0131 ,
		_w5617_
	);
	LUT4 #(
		.INIT('h0080)
	) name3471 (
		\u12_dout_reg[31]/P0001 ,
		\u12_o8_we_reg/P0001 ,
		\u7_wp_reg[0]/P0001 ,
		\u7_wp_reg[1]/NET0131 ,
		_w5618_
	);
	LUT2 #(
		.INIT('he)
	) name3472 (
		_w5617_,
		_w5618_,
		_w5619_
	);
	LUT4 #(
		.INIT('hcc4c)
	) name3473 (
		\u12_o8_we_reg/P0001 ,
		\u7_mem_reg[1][3]/NET0131 ,
		\u7_wp_reg[0]/P0001 ,
		\u7_wp_reg[1]/NET0131 ,
		_w5620_
	);
	LUT4 #(
		.INIT('h0080)
	) name3474 (
		\u12_dout_reg[3]/P0001 ,
		\u12_o8_we_reg/P0001 ,
		\u7_wp_reg[0]/P0001 ,
		\u7_wp_reg[1]/NET0131 ,
		_w5621_
	);
	LUT2 #(
		.INIT('he)
	) name3475 (
		_w5620_,
		_w5621_,
		_w5622_
	);
	LUT4 #(
		.INIT('hcc4c)
	) name3476 (
		\u12_o8_we_reg/P0001 ,
		\u7_mem_reg[1][4]/NET0131 ,
		\u7_wp_reg[0]/P0001 ,
		\u7_wp_reg[1]/NET0131 ,
		_w5623_
	);
	LUT4 #(
		.INIT('h0080)
	) name3477 (
		\u12_dout_reg[4]/P0001 ,
		\u12_o8_we_reg/P0001 ,
		\u7_wp_reg[0]/P0001 ,
		\u7_wp_reg[1]/NET0131 ,
		_w5624_
	);
	LUT2 #(
		.INIT('he)
	) name3478 (
		_w5623_,
		_w5624_,
		_w5625_
	);
	LUT4 #(
		.INIT('hcc4c)
	) name3479 (
		\u12_o8_we_reg/P0001 ,
		\u7_mem_reg[1][5]/NET0131 ,
		\u7_wp_reg[0]/P0001 ,
		\u7_wp_reg[1]/NET0131 ,
		_w5626_
	);
	LUT4 #(
		.INIT('h0080)
	) name3480 (
		\u12_dout_reg[5]/P0001 ,
		\u12_o8_we_reg/P0001 ,
		\u7_wp_reg[0]/P0001 ,
		\u7_wp_reg[1]/NET0131 ,
		_w5627_
	);
	LUT2 #(
		.INIT('he)
	) name3481 (
		_w5626_,
		_w5627_,
		_w5628_
	);
	LUT4 #(
		.INIT('hcc4c)
	) name3482 (
		\u12_o8_we_reg/P0001 ,
		\u7_mem_reg[1][6]/NET0131 ,
		\u7_wp_reg[0]/P0001 ,
		\u7_wp_reg[1]/NET0131 ,
		_w5629_
	);
	LUT4 #(
		.INIT('h0080)
	) name3483 (
		\u12_dout_reg[6]/P0001 ,
		\u12_o8_we_reg/P0001 ,
		\u7_wp_reg[0]/P0001 ,
		\u7_wp_reg[1]/NET0131 ,
		_w5630_
	);
	LUT2 #(
		.INIT('he)
	) name3484 (
		_w5629_,
		_w5630_,
		_w5631_
	);
	LUT4 #(
		.INIT('hcc4c)
	) name3485 (
		\u12_o8_we_reg/P0001 ,
		\u7_mem_reg[1][7]/NET0131 ,
		\u7_wp_reg[0]/P0001 ,
		\u7_wp_reg[1]/NET0131 ,
		_w5632_
	);
	LUT4 #(
		.INIT('h0080)
	) name3486 (
		\u12_dout_reg[7]/P0001 ,
		\u12_o8_we_reg/P0001 ,
		\u7_wp_reg[0]/P0001 ,
		\u7_wp_reg[1]/NET0131 ,
		_w5633_
	);
	LUT2 #(
		.INIT('he)
	) name3487 (
		_w5632_,
		_w5633_,
		_w5634_
	);
	LUT4 #(
		.INIT('hcc4c)
	) name3488 (
		\u12_o8_we_reg/P0001 ,
		\u7_mem_reg[1][8]/NET0131 ,
		\u7_wp_reg[0]/P0001 ,
		\u7_wp_reg[1]/NET0131 ,
		_w5635_
	);
	LUT4 #(
		.INIT('h0080)
	) name3489 (
		\u12_dout_reg[8]/P0001 ,
		\u12_o8_we_reg/P0001 ,
		\u7_wp_reg[0]/P0001 ,
		\u7_wp_reg[1]/NET0131 ,
		_w5636_
	);
	LUT2 #(
		.INIT('he)
	) name3490 (
		_w5635_,
		_w5636_,
		_w5637_
	);
	LUT4 #(
		.INIT('h4ccc)
	) name3491 (
		\u12_o3_we_reg/P0001 ,
		\u3_mem_reg[3][20]/NET0131 ,
		\u3_wp_reg[0]/P0001 ,
		\u3_wp_reg[1]/NET0131 ,
		_w5638_
	);
	LUT4 #(
		.INIT('h8000)
	) name3492 (
		\u12_dout_reg[20]/P0001 ,
		\u12_o3_we_reg/P0001 ,
		\u3_wp_reg[0]/P0001 ,
		\u3_wp_reg[1]/NET0131 ,
		_w5639_
	);
	LUT2 #(
		.INIT('he)
	) name3493 (
		_w5638_,
		_w5639_,
		_w5640_
	);
	LUT4 #(
		.INIT('hcc4c)
	) name3494 (
		\u12_o8_we_reg/P0001 ,
		\u7_mem_reg[1][9]/NET0131 ,
		\u7_wp_reg[0]/P0001 ,
		\u7_wp_reg[1]/NET0131 ,
		_w5641_
	);
	LUT4 #(
		.INIT('h0080)
	) name3495 (
		\u12_dout_reg[9]/P0001 ,
		\u12_o8_we_reg/P0001 ,
		\u7_wp_reg[0]/P0001 ,
		\u7_wp_reg[1]/NET0131 ,
		_w5642_
	);
	LUT2 #(
		.INIT('he)
	) name3496 (
		_w5641_,
		_w5642_,
		_w5643_
	);
	LUT4 #(
		.INIT('hc4cc)
	) name3497 (
		\u12_o8_we_reg/P0001 ,
		\u7_mem_reg[2][0]/NET0131 ,
		\u7_wp_reg[0]/P0001 ,
		\u7_wp_reg[1]/NET0131 ,
		_w5644_
	);
	LUT4 #(
		.INIT('h0800)
	) name3498 (
		\u12_dout_reg[0]/P0001 ,
		\u12_o8_we_reg/P0001 ,
		\u7_wp_reg[0]/P0001 ,
		\u7_wp_reg[1]/NET0131 ,
		_w5645_
	);
	LUT2 #(
		.INIT('he)
	) name3499 (
		_w5644_,
		_w5645_,
		_w5646_
	);
	LUT4 #(
		.INIT('hc4cc)
	) name3500 (
		\u12_o8_we_reg/P0001 ,
		\u7_mem_reg[2][10]/NET0131 ,
		\u7_wp_reg[0]/P0001 ,
		\u7_wp_reg[1]/NET0131 ,
		_w5647_
	);
	LUT4 #(
		.INIT('h0800)
	) name3501 (
		\u12_dout_reg[10]/P0001 ,
		\u12_o8_we_reg/P0001 ,
		\u7_wp_reg[0]/P0001 ,
		\u7_wp_reg[1]/NET0131 ,
		_w5648_
	);
	LUT2 #(
		.INIT('he)
	) name3502 (
		_w5647_,
		_w5648_,
		_w5649_
	);
	LUT4 #(
		.INIT('hc4cc)
	) name3503 (
		\u12_o8_we_reg/P0001 ,
		\u7_mem_reg[2][11]/NET0131 ,
		\u7_wp_reg[0]/P0001 ,
		\u7_wp_reg[1]/NET0131 ,
		_w5650_
	);
	LUT4 #(
		.INIT('h0800)
	) name3504 (
		\u12_dout_reg[11]/P0001 ,
		\u12_o8_we_reg/P0001 ,
		\u7_wp_reg[0]/P0001 ,
		\u7_wp_reg[1]/NET0131 ,
		_w5651_
	);
	LUT2 #(
		.INIT('he)
	) name3505 (
		_w5650_,
		_w5651_,
		_w5652_
	);
	LUT4 #(
		.INIT('hc4cc)
	) name3506 (
		\u12_o8_we_reg/P0001 ,
		\u7_mem_reg[2][12]/NET0131 ,
		\u7_wp_reg[0]/P0001 ,
		\u7_wp_reg[1]/NET0131 ,
		_w5653_
	);
	LUT4 #(
		.INIT('h0800)
	) name3507 (
		\u12_dout_reg[12]/P0001 ,
		\u12_o8_we_reg/P0001 ,
		\u7_wp_reg[0]/P0001 ,
		\u7_wp_reg[1]/NET0131 ,
		_w5654_
	);
	LUT2 #(
		.INIT('he)
	) name3508 (
		_w5653_,
		_w5654_,
		_w5655_
	);
	LUT4 #(
		.INIT('hc4cc)
	) name3509 (
		\u12_o8_we_reg/P0001 ,
		\u7_mem_reg[2][13]/NET0131 ,
		\u7_wp_reg[0]/P0001 ,
		\u7_wp_reg[1]/NET0131 ,
		_w5656_
	);
	LUT4 #(
		.INIT('h0800)
	) name3510 (
		\u12_dout_reg[13]/P0001 ,
		\u12_o8_we_reg/P0001 ,
		\u7_wp_reg[0]/P0001 ,
		\u7_wp_reg[1]/NET0131 ,
		_w5657_
	);
	LUT2 #(
		.INIT('he)
	) name3511 (
		_w5656_,
		_w5657_,
		_w5658_
	);
	LUT4 #(
		.INIT('hc4cc)
	) name3512 (
		\u12_o8_we_reg/P0001 ,
		\u7_mem_reg[2][14]/NET0131 ,
		\u7_wp_reg[0]/P0001 ,
		\u7_wp_reg[1]/NET0131 ,
		_w5659_
	);
	LUT4 #(
		.INIT('h0800)
	) name3513 (
		\u12_dout_reg[14]/P0001 ,
		\u12_o8_we_reg/P0001 ,
		\u7_wp_reg[0]/P0001 ,
		\u7_wp_reg[1]/NET0131 ,
		_w5660_
	);
	LUT2 #(
		.INIT('he)
	) name3514 (
		_w5659_,
		_w5660_,
		_w5661_
	);
	LUT4 #(
		.INIT('hc4cc)
	) name3515 (
		\u12_o8_we_reg/P0001 ,
		\u7_mem_reg[2][15]/NET0131 ,
		\u7_wp_reg[0]/P0001 ,
		\u7_wp_reg[1]/NET0131 ,
		_w5662_
	);
	LUT4 #(
		.INIT('h0800)
	) name3516 (
		\u12_dout_reg[15]/P0001 ,
		\u12_o8_we_reg/P0001 ,
		\u7_wp_reg[0]/P0001 ,
		\u7_wp_reg[1]/NET0131 ,
		_w5663_
	);
	LUT2 #(
		.INIT('he)
	) name3517 (
		_w5662_,
		_w5663_,
		_w5664_
	);
	LUT4 #(
		.INIT('hc4cc)
	) name3518 (
		\u12_o8_we_reg/P0001 ,
		\u7_mem_reg[2][16]/NET0131 ,
		\u7_wp_reg[0]/P0001 ,
		\u7_wp_reg[1]/NET0131 ,
		_w5665_
	);
	LUT4 #(
		.INIT('h0800)
	) name3519 (
		\u12_dout_reg[16]/P0001 ,
		\u12_o8_we_reg/P0001 ,
		\u7_wp_reg[0]/P0001 ,
		\u7_wp_reg[1]/NET0131 ,
		_w5666_
	);
	LUT2 #(
		.INIT('he)
	) name3520 (
		_w5665_,
		_w5666_,
		_w5667_
	);
	LUT4 #(
		.INIT('hc4cc)
	) name3521 (
		\u12_o8_we_reg/P0001 ,
		\u7_mem_reg[2][17]/NET0131 ,
		\u7_wp_reg[0]/P0001 ,
		\u7_wp_reg[1]/NET0131 ,
		_w5668_
	);
	LUT4 #(
		.INIT('h0800)
	) name3522 (
		\u12_dout_reg[17]/P0001 ,
		\u12_o8_we_reg/P0001 ,
		\u7_wp_reg[0]/P0001 ,
		\u7_wp_reg[1]/NET0131 ,
		_w5669_
	);
	LUT2 #(
		.INIT('he)
	) name3523 (
		_w5668_,
		_w5669_,
		_w5670_
	);
	LUT4 #(
		.INIT('hc4cc)
	) name3524 (
		\u12_o8_we_reg/P0001 ,
		\u7_mem_reg[2][18]/NET0131 ,
		\u7_wp_reg[0]/P0001 ,
		\u7_wp_reg[1]/NET0131 ,
		_w5671_
	);
	LUT4 #(
		.INIT('h0800)
	) name3525 (
		\u12_dout_reg[18]/P0001 ,
		\u12_o8_we_reg/P0001 ,
		\u7_wp_reg[0]/P0001 ,
		\u7_wp_reg[1]/NET0131 ,
		_w5672_
	);
	LUT2 #(
		.INIT('he)
	) name3526 (
		_w5671_,
		_w5672_,
		_w5673_
	);
	LUT4 #(
		.INIT('hc4cc)
	) name3527 (
		\u12_o8_we_reg/P0001 ,
		\u7_mem_reg[2][19]/NET0131 ,
		\u7_wp_reg[0]/P0001 ,
		\u7_wp_reg[1]/NET0131 ,
		_w5674_
	);
	LUT4 #(
		.INIT('h0800)
	) name3528 (
		\u12_dout_reg[19]/P0001 ,
		\u12_o8_we_reg/P0001 ,
		\u7_wp_reg[0]/P0001 ,
		\u7_wp_reg[1]/NET0131 ,
		_w5675_
	);
	LUT2 #(
		.INIT('he)
	) name3529 (
		_w5674_,
		_w5675_,
		_w5676_
	);
	LUT4 #(
		.INIT('hc4cc)
	) name3530 (
		\u12_o8_we_reg/P0001 ,
		\u7_mem_reg[2][1]/NET0131 ,
		\u7_wp_reg[0]/P0001 ,
		\u7_wp_reg[1]/NET0131 ,
		_w5677_
	);
	LUT4 #(
		.INIT('h0800)
	) name3531 (
		\u12_dout_reg[1]/P0001 ,
		\u12_o8_we_reg/P0001 ,
		\u7_wp_reg[0]/P0001 ,
		\u7_wp_reg[1]/NET0131 ,
		_w5678_
	);
	LUT2 #(
		.INIT('he)
	) name3532 (
		_w5677_,
		_w5678_,
		_w5679_
	);
	LUT4 #(
		.INIT('hc4cc)
	) name3533 (
		\u12_o8_we_reg/P0001 ,
		\u7_mem_reg[2][20]/NET0131 ,
		\u7_wp_reg[0]/P0001 ,
		\u7_wp_reg[1]/NET0131 ,
		_w5680_
	);
	LUT4 #(
		.INIT('h0800)
	) name3534 (
		\u12_dout_reg[20]/P0001 ,
		\u12_o8_we_reg/P0001 ,
		\u7_wp_reg[0]/P0001 ,
		\u7_wp_reg[1]/NET0131 ,
		_w5681_
	);
	LUT2 #(
		.INIT('he)
	) name3535 (
		_w5680_,
		_w5681_,
		_w5682_
	);
	LUT4 #(
		.INIT('hc4cc)
	) name3536 (
		\u12_o8_we_reg/P0001 ,
		\u7_mem_reg[2][21]/NET0131 ,
		\u7_wp_reg[0]/P0001 ,
		\u7_wp_reg[1]/NET0131 ,
		_w5683_
	);
	LUT4 #(
		.INIT('h0800)
	) name3537 (
		\u12_dout_reg[21]/P0001 ,
		\u12_o8_we_reg/P0001 ,
		\u7_wp_reg[0]/P0001 ,
		\u7_wp_reg[1]/NET0131 ,
		_w5684_
	);
	LUT2 #(
		.INIT('he)
	) name3538 (
		_w5683_,
		_w5684_,
		_w5685_
	);
	LUT4 #(
		.INIT('hc4cc)
	) name3539 (
		\u12_o8_we_reg/P0001 ,
		\u7_mem_reg[2][22]/NET0131 ,
		\u7_wp_reg[0]/P0001 ,
		\u7_wp_reg[1]/NET0131 ,
		_w5686_
	);
	LUT4 #(
		.INIT('h0800)
	) name3540 (
		\u12_dout_reg[22]/P0001 ,
		\u12_o8_we_reg/P0001 ,
		\u7_wp_reg[0]/P0001 ,
		\u7_wp_reg[1]/NET0131 ,
		_w5687_
	);
	LUT2 #(
		.INIT('he)
	) name3541 (
		_w5686_,
		_w5687_,
		_w5688_
	);
	LUT4 #(
		.INIT('hc4cc)
	) name3542 (
		\u12_o8_we_reg/P0001 ,
		\u7_mem_reg[2][23]/NET0131 ,
		\u7_wp_reg[0]/P0001 ,
		\u7_wp_reg[1]/NET0131 ,
		_w5689_
	);
	LUT4 #(
		.INIT('h0800)
	) name3543 (
		\u12_dout_reg[23]/P0001 ,
		\u12_o8_we_reg/P0001 ,
		\u7_wp_reg[0]/P0001 ,
		\u7_wp_reg[1]/NET0131 ,
		_w5690_
	);
	LUT2 #(
		.INIT('he)
	) name3544 (
		_w5689_,
		_w5690_,
		_w5691_
	);
	LUT4 #(
		.INIT('hc4cc)
	) name3545 (
		\u12_o8_we_reg/P0001 ,
		\u7_mem_reg[2][24]/NET0131 ,
		\u7_wp_reg[0]/P0001 ,
		\u7_wp_reg[1]/NET0131 ,
		_w5692_
	);
	LUT4 #(
		.INIT('h0800)
	) name3546 (
		\u12_dout_reg[24]/P0001 ,
		\u12_o8_we_reg/P0001 ,
		\u7_wp_reg[0]/P0001 ,
		\u7_wp_reg[1]/NET0131 ,
		_w5693_
	);
	LUT2 #(
		.INIT('he)
	) name3547 (
		_w5692_,
		_w5693_,
		_w5694_
	);
	LUT4 #(
		.INIT('hc4cc)
	) name3548 (
		\u12_o8_we_reg/P0001 ,
		\u7_mem_reg[2][25]/NET0131 ,
		\u7_wp_reg[0]/P0001 ,
		\u7_wp_reg[1]/NET0131 ,
		_w5695_
	);
	LUT4 #(
		.INIT('h0800)
	) name3549 (
		\u12_dout_reg[25]/P0001 ,
		\u12_o8_we_reg/P0001 ,
		\u7_wp_reg[0]/P0001 ,
		\u7_wp_reg[1]/NET0131 ,
		_w5696_
	);
	LUT2 #(
		.INIT('he)
	) name3550 (
		_w5695_,
		_w5696_,
		_w5697_
	);
	LUT4 #(
		.INIT('hc4cc)
	) name3551 (
		\u12_o8_we_reg/P0001 ,
		\u7_mem_reg[2][26]/NET0131 ,
		\u7_wp_reg[0]/P0001 ,
		\u7_wp_reg[1]/NET0131 ,
		_w5698_
	);
	LUT4 #(
		.INIT('h0800)
	) name3552 (
		\u12_dout_reg[26]/P0001 ,
		\u12_o8_we_reg/P0001 ,
		\u7_wp_reg[0]/P0001 ,
		\u7_wp_reg[1]/NET0131 ,
		_w5699_
	);
	LUT2 #(
		.INIT('he)
	) name3553 (
		_w5698_,
		_w5699_,
		_w5700_
	);
	LUT4 #(
		.INIT('hc4cc)
	) name3554 (
		\u12_o8_we_reg/P0001 ,
		\u7_mem_reg[2][27]/NET0131 ,
		\u7_wp_reg[0]/P0001 ,
		\u7_wp_reg[1]/NET0131 ,
		_w5701_
	);
	LUT4 #(
		.INIT('h0800)
	) name3555 (
		\u12_dout_reg[27]/P0001 ,
		\u12_o8_we_reg/P0001 ,
		\u7_wp_reg[0]/P0001 ,
		\u7_wp_reg[1]/NET0131 ,
		_w5702_
	);
	LUT2 #(
		.INIT('he)
	) name3556 (
		_w5701_,
		_w5702_,
		_w5703_
	);
	LUT4 #(
		.INIT('hc4cc)
	) name3557 (
		\u12_o8_we_reg/P0001 ,
		\u7_mem_reg[2][28]/NET0131 ,
		\u7_wp_reg[0]/P0001 ,
		\u7_wp_reg[1]/NET0131 ,
		_w5704_
	);
	LUT4 #(
		.INIT('h0800)
	) name3558 (
		\u12_dout_reg[28]/P0001 ,
		\u12_o8_we_reg/P0001 ,
		\u7_wp_reg[0]/P0001 ,
		\u7_wp_reg[1]/NET0131 ,
		_w5705_
	);
	LUT2 #(
		.INIT('he)
	) name3559 (
		_w5704_,
		_w5705_,
		_w5706_
	);
	LUT4 #(
		.INIT('hc4cc)
	) name3560 (
		\u12_o8_we_reg/P0001 ,
		\u7_mem_reg[2][29]/NET0131 ,
		\u7_wp_reg[0]/P0001 ,
		\u7_wp_reg[1]/NET0131 ,
		_w5707_
	);
	LUT4 #(
		.INIT('h0800)
	) name3561 (
		\u12_dout_reg[29]/P0001 ,
		\u12_o8_we_reg/P0001 ,
		\u7_wp_reg[0]/P0001 ,
		\u7_wp_reg[1]/NET0131 ,
		_w5708_
	);
	LUT2 #(
		.INIT('he)
	) name3562 (
		_w5707_,
		_w5708_,
		_w5709_
	);
	LUT4 #(
		.INIT('hc4cc)
	) name3563 (
		\u12_o8_we_reg/P0001 ,
		\u7_mem_reg[2][2]/NET0131 ,
		\u7_wp_reg[0]/P0001 ,
		\u7_wp_reg[1]/NET0131 ,
		_w5710_
	);
	LUT4 #(
		.INIT('h0800)
	) name3564 (
		\u12_dout_reg[2]/P0001 ,
		\u12_o8_we_reg/P0001 ,
		\u7_wp_reg[0]/P0001 ,
		\u7_wp_reg[1]/NET0131 ,
		_w5711_
	);
	LUT2 #(
		.INIT('he)
	) name3565 (
		_w5710_,
		_w5711_,
		_w5712_
	);
	LUT4 #(
		.INIT('hc4cc)
	) name3566 (
		\u12_o8_we_reg/P0001 ,
		\u7_mem_reg[2][30]/NET0131 ,
		\u7_wp_reg[0]/P0001 ,
		\u7_wp_reg[1]/NET0131 ,
		_w5713_
	);
	LUT4 #(
		.INIT('h0800)
	) name3567 (
		\u12_dout_reg[30]/P0001 ,
		\u12_o8_we_reg/P0001 ,
		\u7_wp_reg[0]/P0001 ,
		\u7_wp_reg[1]/NET0131 ,
		_w5714_
	);
	LUT2 #(
		.INIT('he)
	) name3568 (
		_w5713_,
		_w5714_,
		_w5715_
	);
	LUT4 #(
		.INIT('hc4cc)
	) name3569 (
		\u12_o8_we_reg/P0001 ,
		\u7_mem_reg[2][31]/NET0131 ,
		\u7_wp_reg[0]/P0001 ,
		\u7_wp_reg[1]/NET0131 ,
		_w5716_
	);
	LUT4 #(
		.INIT('h0800)
	) name3570 (
		\u12_dout_reg[31]/P0001 ,
		\u12_o8_we_reg/P0001 ,
		\u7_wp_reg[0]/P0001 ,
		\u7_wp_reg[1]/NET0131 ,
		_w5717_
	);
	LUT2 #(
		.INIT('he)
	) name3571 (
		_w5716_,
		_w5717_,
		_w5718_
	);
	LUT4 #(
		.INIT('hc4cc)
	) name3572 (
		\u12_o8_we_reg/P0001 ,
		\u7_mem_reg[2][3]/NET0131 ,
		\u7_wp_reg[0]/P0001 ,
		\u7_wp_reg[1]/NET0131 ,
		_w5719_
	);
	LUT4 #(
		.INIT('h0800)
	) name3573 (
		\u12_dout_reg[3]/P0001 ,
		\u12_o8_we_reg/P0001 ,
		\u7_wp_reg[0]/P0001 ,
		\u7_wp_reg[1]/NET0131 ,
		_w5720_
	);
	LUT2 #(
		.INIT('he)
	) name3574 (
		_w5719_,
		_w5720_,
		_w5721_
	);
	LUT4 #(
		.INIT('hc4cc)
	) name3575 (
		\u12_o8_we_reg/P0001 ,
		\u7_mem_reg[2][4]/NET0131 ,
		\u7_wp_reg[0]/P0001 ,
		\u7_wp_reg[1]/NET0131 ,
		_w5722_
	);
	LUT4 #(
		.INIT('h0800)
	) name3576 (
		\u12_dout_reg[4]/P0001 ,
		\u12_o8_we_reg/P0001 ,
		\u7_wp_reg[0]/P0001 ,
		\u7_wp_reg[1]/NET0131 ,
		_w5723_
	);
	LUT2 #(
		.INIT('he)
	) name3577 (
		_w5722_,
		_w5723_,
		_w5724_
	);
	LUT4 #(
		.INIT('hc4cc)
	) name3578 (
		\u12_o8_we_reg/P0001 ,
		\u7_mem_reg[2][5]/NET0131 ,
		\u7_wp_reg[0]/P0001 ,
		\u7_wp_reg[1]/NET0131 ,
		_w5725_
	);
	LUT4 #(
		.INIT('h0800)
	) name3579 (
		\u12_dout_reg[5]/P0001 ,
		\u12_o8_we_reg/P0001 ,
		\u7_wp_reg[0]/P0001 ,
		\u7_wp_reg[1]/NET0131 ,
		_w5726_
	);
	LUT2 #(
		.INIT('he)
	) name3580 (
		_w5725_,
		_w5726_,
		_w5727_
	);
	LUT4 #(
		.INIT('hc4cc)
	) name3581 (
		\u12_o8_we_reg/P0001 ,
		\u7_mem_reg[2][6]/NET0131 ,
		\u7_wp_reg[0]/P0001 ,
		\u7_wp_reg[1]/NET0131 ,
		_w5728_
	);
	LUT4 #(
		.INIT('h0800)
	) name3582 (
		\u12_dout_reg[6]/P0001 ,
		\u12_o8_we_reg/P0001 ,
		\u7_wp_reg[0]/P0001 ,
		\u7_wp_reg[1]/NET0131 ,
		_w5729_
	);
	LUT2 #(
		.INIT('he)
	) name3583 (
		_w5728_,
		_w5729_,
		_w5730_
	);
	LUT4 #(
		.INIT('hc4cc)
	) name3584 (
		\u12_o8_we_reg/P0001 ,
		\u7_mem_reg[2][7]/NET0131 ,
		\u7_wp_reg[0]/P0001 ,
		\u7_wp_reg[1]/NET0131 ,
		_w5731_
	);
	LUT4 #(
		.INIT('h0800)
	) name3585 (
		\u12_dout_reg[7]/P0001 ,
		\u12_o8_we_reg/P0001 ,
		\u7_wp_reg[0]/P0001 ,
		\u7_wp_reg[1]/NET0131 ,
		_w5732_
	);
	LUT2 #(
		.INIT('he)
	) name3586 (
		_w5731_,
		_w5732_,
		_w5733_
	);
	LUT4 #(
		.INIT('hc4cc)
	) name3587 (
		\u12_o8_we_reg/P0001 ,
		\u7_mem_reg[2][8]/NET0131 ,
		\u7_wp_reg[0]/P0001 ,
		\u7_wp_reg[1]/NET0131 ,
		_w5734_
	);
	LUT4 #(
		.INIT('h0800)
	) name3588 (
		\u12_dout_reg[8]/P0001 ,
		\u12_o8_we_reg/P0001 ,
		\u7_wp_reg[0]/P0001 ,
		\u7_wp_reg[1]/NET0131 ,
		_w5735_
	);
	LUT2 #(
		.INIT('he)
	) name3589 (
		_w5734_,
		_w5735_,
		_w5736_
	);
	LUT4 #(
		.INIT('hc4cc)
	) name3590 (
		\u12_o8_we_reg/P0001 ,
		\u7_mem_reg[2][9]/NET0131 ,
		\u7_wp_reg[0]/P0001 ,
		\u7_wp_reg[1]/NET0131 ,
		_w5737_
	);
	LUT4 #(
		.INIT('h0800)
	) name3591 (
		\u12_dout_reg[9]/P0001 ,
		\u12_o8_we_reg/P0001 ,
		\u7_wp_reg[0]/P0001 ,
		\u7_wp_reg[1]/NET0131 ,
		_w5738_
	);
	LUT2 #(
		.INIT('he)
	) name3592 (
		_w5737_,
		_w5738_,
		_w5739_
	);
	LUT4 #(
		.INIT('h4ccc)
	) name3593 (
		\u12_o8_we_reg/P0001 ,
		\u7_mem_reg[3][0]/NET0131 ,
		\u7_wp_reg[0]/P0001 ,
		\u7_wp_reg[1]/NET0131 ,
		_w5740_
	);
	LUT4 #(
		.INIT('h8000)
	) name3594 (
		\u12_dout_reg[0]/P0001 ,
		\u12_o8_we_reg/P0001 ,
		\u7_wp_reg[0]/P0001 ,
		\u7_wp_reg[1]/NET0131 ,
		_w5741_
	);
	LUT2 #(
		.INIT('he)
	) name3595 (
		_w5740_,
		_w5741_,
		_w5742_
	);
	LUT4 #(
		.INIT('h4ccc)
	) name3596 (
		\u12_o8_we_reg/P0001 ,
		\u7_mem_reg[3][10]/NET0131 ,
		\u7_wp_reg[0]/P0001 ,
		\u7_wp_reg[1]/NET0131 ,
		_w5743_
	);
	LUT4 #(
		.INIT('h8000)
	) name3597 (
		\u12_dout_reg[10]/P0001 ,
		\u12_o8_we_reg/P0001 ,
		\u7_wp_reg[0]/P0001 ,
		\u7_wp_reg[1]/NET0131 ,
		_w5744_
	);
	LUT2 #(
		.INIT('he)
	) name3598 (
		_w5743_,
		_w5744_,
		_w5745_
	);
	LUT4 #(
		.INIT('h4ccc)
	) name3599 (
		\u12_o8_we_reg/P0001 ,
		\u7_mem_reg[3][11]/NET0131 ,
		\u7_wp_reg[0]/P0001 ,
		\u7_wp_reg[1]/NET0131 ,
		_w5746_
	);
	LUT4 #(
		.INIT('h8000)
	) name3600 (
		\u12_dout_reg[11]/P0001 ,
		\u12_o8_we_reg/P0001 ,
		\u7_wp_reg[0]/P0001 ,
		\u7_wp_reg[1]/NET0131 ,
		_w5747_
	);
	LUT2 #(
		.INIT('he)
	) name3601 (
		_w5746_,
		_w5747_,
		_w5748_
	);
	LUT4 #(
		.INIT('h4ccc)
	) name3602 (
		\u12_o8_we_reg/P0001 ,
		\u7_mem_reg[3][12]/NET0131 ,
		\u7_wp_reg[0]/P0001 ,
		\u7_wp_reg[1]/NET0131 ,
		_w5749_
	);
	LUT4 #(
		.INIT('h8000)
	) name3603 (
		\u12_dout_reg[12]/P0001 ,
		\u12_o8_we_reg/P0001 ,
		\u7_wp_reg[0]/P0001 ,
		\u7_wp_reg[1]/NET0131 ,
		_w5750_
	);
	LUT2 #(
		.INIT('he)
	) name3604 (
		_w5749_,
		_w5750_,
		_w5751_
	);
	LUT4 #(
		.INIT('h4ccc)
	) name3605 (
		\u12_o8_we_reg/P0001 ,
		\u7_mem_reg[3][13]/NET0131 ,
		\u7_wp_reg[0]/P0001 ,
		\u7_wp_reg[1]/NET0131 ,
		_w5752_
	);
	LUT4 #(
		.INIT('h8000)
	) name3606 (
		\u12_dout_reg[13]/P0001 ,
		\u12_o8_we_reg/P0001 ,
		\u7_wp_reg[0]/P0001 ,
		\u7_wp_reg[1]/NET0131 ,
		_w5753_
	);
	LUT2 #(
		.INIT('he)
	) name3607 (
		_w5752_,
		_w5753_,
		_w5754_
	);
	LUT4 #(
		.INIT('h4ccc)
	) name3608 (
		\u12_o8_we_reg/P0001 ,
		\u7_mem_reg[3][14]/NET0131 ,
		\u7_wp_reg[0]/P0001 ,
		\u7_wp_reg[1]/NET0131 ,
		_w5755_
	);
	LUT4 #(
		.INIT('h8000)
	) name3609 (
		\u12_dout_reg[14]/P0001 ,
		\u12_o8_we_reg/P0001 ,
		\u7_wp_reg[0]/P0001 ,
		\u7_wp_reg[1]/NET0131 ,
		_w5756_
	);
	LUT2 #(
		.INIT('he)
	) name3610 (
		_w5755_,
		_w5756_,
		_w5757_
	);
	LUT4 #(
		.INIT('h4ccc)
	) name3611 (
		\u12_o8_we_reg/P0001 ,
		\u7_mem_reg[3][15]/NET0131 ,
		\u7_wp_reg[0]/P0001 ,
		\u7_wp_reg[1]/NET0131 ,
		_w5758_
	);
	LUT4 #(
		.INIT('h8000)
	) name3612 (
		\u12_dout_reg[15]/P0001 ,
		\u12_o8_we_reg/P0001 ,
		\u7_wp_reg[0]/P0001 ,
		\u7_wp_reg[1]/NET0131 ,
		_w5759_
	);
	LUT2 #(
		.INIT('he)
	) name3613 (
		_w5758_,
		_w5759_,
		_w5760_
	);
	LUT4 #(
		.INIT('h4ccc)
	) name3614 (
		\u12_o8_we_reg/P0001 ,
		\u7_mem_reg[3][16]/NET0131 ,
		\u7_wp_reg[0]/P0001 ,
		\u7_wp_reg[1]/NET0131 ,
		_w5761_
	);
	LUT4 #(
		.INIT('h8000)
	) name3615 (
		\u12_dout_reg[16]/P0001 ,
		\u12_o8_we_reg/P0001 ,
		\u7_wp_reg[0]/P0001 ,
		\u7_wp_reg[1]/NET0131 ,
		_w5762_
	);
	LUT2 #(
		.INIT('he)
	) name3616 (
		_w5761_,
		_w5762_,
		_w5763_
	);
	LUT4 #(
		.INIT('h4ccc)
	) name3617 (
		\u12_o8_we_reg/P0001 ,
		\u7_mem_reg[3][17]/NET0131 ,
		\u7_wp_reg[0]/P0001 ,
		\u7_wp_reg[1]/NET0131 ,
		_w5764_
	);
	LUT4 #(
		.INIT('h8000)
	) name3618 (
		\u12_dout_reg[17]/P0001 ,
		\u12_o8_we_reg/P0001 ,
		\u7_wp_reg[0]/P0001 ,
		\u7_wp_reg[1]/NET0131 ,
		_w5765_
	);
	LUT2 #(
		.INIT('he)
	) name3619 (
		_w5764_,
		_w5765_,
		_w5766_
	);
	LUT4 #(
		.INIT('h4ccc)
	) name3620 (
		\u12_o8_we_reg/P0001 ,
		\u7_mem_reg[3][18]/NET0131 ,
		\u7_wp_reg[0]/P0001 ,
		\u7_wp_reg[1]/NET0131 ,
		_w5767_
	);
	LUT4 #(
		.INIT('h8000)
	) name3621 (
		\u12_dout_reg[18]/P0001 ,
		\u12_o8_we_reg/P0001 ,
		\u7_wp_reg[0]/P0001 ,
		\u7_wp_reg[1]/NET0131 ,
		_w5768_
	);
	LUT2 #(
		.INIT('he)
	) name3622 (
		_w5767_,
		_w5768_,
		_w5769_
	);
	LUT4 #(
		.INIT('h4ccc)
	) name3623 (
		\u12_o8_we_reg/P0001 ,
		\u7_mem_reg[3][19]/NET0131 ,
		\u7_wp_reg[0]/P0001 ,
		\u7_wp_reg[1]/NET0131 ,
		_w5770_
	);
	LUT4 #(
		.INIT('h8000)
	) name3624 (
		\u12_dout_reg[19]/P0001 ,
		\u12_o8_we_reg/P0001 ,
		\u7_wp_reg[0]/P0001 ,
		\u7_wp_reg[1]/NET0131 ,
		_w5771_
	);
	LUT2 #(
		.INIT('he)
	) name3625 (
		_w5770_,
		_w5771_,
		_w5772_
	);
	LUT4 #(
		.INIT('h4ccc)
	) name3626 (
		\u12_o8_we_reg/P0001 ,
		\u7_mem_reg[3][1]/NET0131 ,
		\u7_wp_reg[0]/P0001 ,
		\u7_wp_reg[1]/NET0131 ,
		_w5773_
	);
	LUT4 #(
		.INIT('h8000)
	) name3627 (
		\u12_dout_reg[1]/P0001 ,
		\u12_o8_we_reg/P0001 ,
		\u7_wp_reg[0]/P0001 ,
		\u7_wp_reg[1]/NET0131 ,
		_w5774_
	);
	LUT2 #(
		.INIT('he)
	) name3628 (
		_w5773_,
		_w5774_,
		_w5775_
	);
	LUT4 #(
		.INIT('h4ccc)
	) name3629 (
		\u12_o8_we_reg/P0001 ,
		\u7_mem_reg[3][20]/NET0131 ,
		\u7_wp_reg[0]/P0001 ,
		\u7_wp_reg[1]/NET0131 ,
		_w5776_
	);
	LUT4 #(
		.INIT('h8000)
	) name3630 (
		\u12_dout_reg[20]/P0001 ,
		\u12_o8_we_reg/P0001 ,
		\u7_wp_reg[0]/P0001 ,
		\u7_wp_reg[1]/NET0131 ,
		_w5777_
	);
	LUT2 #(
		.INIT('he)
	) name3631 (
		_w5776_,
		_w5777_,
		_w5778_
	);
	LUT4 #(
		.INIT('h4ccc)
	) name3632 (
		\u12_o8_we_reg/P0001 ,
		\u7_mem_reg[3][21]/NET0131 ,
		\u7_wp_reg[0]/P0001 ,
		\u7_wp_reg[1]/NET0131 ,
		_w5779_
	);
	LUT4 #(
		.INIT('h8000)
	) name3633 (
		\u12_dout_reg[21]/P0001 ,
		\u12_o8_we_reg/P0001 ,
		\u7_wp_reg[0]/P0001 ,
		\u7_wp_reg[1]/NET0131 ,
		_w5780_
	);
	LUT2 #(
		.INIT('he)
	) name3634 (
		_w5779_,
		_w5780_,
		_w5781_
	);
	LUT4 #(
		.INIT('h4ccc)
	) name3635 (
		\u12_o8_we_reg/P0001 ,
		\u7_mem_reg[3][22]/NET0131 ,
		\u7_wp_reg[0]/P0001 ,
		\u7_wp_reg[1]/NET0131 ,
		_w5782_
	);
	LUT4 #(
		.INIT('h8000)
	) name3636 (
		\u12_dout_reg[22]/P0001 ,
		\u12_o8_we_reg/P0001 ,
		\u7_wp_reg[0]/P0001 ,
		\u7_wp_reg[1]/NET0131 ,
		_w5783_
	);
	LUT2 #(
		.INIT('he)
	) name3637 (
		_w5782_,
		_w5783_,
		_w5784_
	);
	LUT4 #(
		.INIT('h4ccc)
	) name3638 (
		\u12_o8_we_reg/P0001 ,
		\u7_mem_reg[3][23]/NET0131 ,
		\u7_wp_reg[0]/P0001 ,
		\u7_wp_reg[1]/NET0131 ,
		_w5785_
	);
	LUT4 #(
		.INIT('h8000)
	) name3639 (
		\u12_dout_reg[23]/P0001 ,
		\u12_o8_we_reg/P0001 ,
		\u7_wp_reg[0]/P0001 ,
		\u7_wp_reg[1]/NET0131 ,
		_w5786_
	);
	LUT2 #(
		.INIT('he)
	) name3640 (
		_w5785_,
		_w5786_,
		_w5787_
	);
	LUT4 #(
		.INIT('h4ccc)
	) name3641 (
		\u12_o8_we_reg/P0001 ,
		\u7_mem_reg[3][24]/NET0131 ,
		\u7_wp_reg[0]/P0001 ,
		\u7_wp_reg[1]/NET0131 ,
		_w5788_
	);
	LUT4 #(
		.INIT('h8000)
	) name3642 (
		\u12_dout_reg[24]/P0001 ,
		\u12_o8_we_reg/P0001 ,
		\u7_wp_reg[0]/P0001 ,
		\u7_wp_reg[1]/NET0131 ,
		_w5789_
	);
	LUT2 #(
		.INIT('he)
	) name3643 (
		_w5788_,
		_w5789_,
		_w5790_
	);
	LUT4 #(
		.INIT('h4ccc)
	) name3644 (
		\u12_o8_we_reg/P0001 ,
		\u7_mem_reg[3][25]/NET0131 ,
		\u7_wp_reg[0]/P0001 ,
		\u7_wp_reg[1]/NET0131 ,
		_w5791_
	);
	LUT4 #(
		.INIT('h8000)
	) name3645 (
		\u12_dout_reg[25]/P0001 ,
		\u12_o8_we_reg/P0001 ,
		\u7_wp_reg[0]/P0001 ,
		\u7_wp_reg[1]/NET0131 ,
		_w5792_
	);
	LUT2 #(
		.INIT('he)
	) name3646 (
		_w5791_,
		_w5792_,
		_w5793_
	);
	LUT4 #(
		.INIT('h4ccc)
	) name3647 (
		\u12_o8_we_reg/P0001 ,
		\u7_mem_reg[3][26]/NET0131 ,
		\u7_wp_reg[0]/P0001 ,
		\u7_wp_reg[1]/NET0131 ,
		_w5794_
	);
	LUT4 #(
		.INIT('h8000)
	) name3648 (
		\u12_dout_reg[26]/P0001 ,
		\u12_o8_we_reg/P0001 ,
		\u7_wp_reg[0]/P0001 ,
		\u7_wp_reg[1]/NET0131 ,
		_w5795_
	);
	LUT2 #(
		.INIT('he)
	) name3649 (
		_w5794_,
		_w5795_,
		_w5796_
	);
	LUT4 #(
		.INIT('h4ccc)
	) name3650 (
		\u12_o8_we_reg/P0001 ,
		\u7_mem_reg[3][27]/NET0131 ,
		\u7_wp_reg[0]/P0001 ,
		\u7_wp_reg[1]/NET0131 ,
		_w5797_
	);
	LUT4 #(
		.INIT('h8000)
	) name3651 (
		\u12_dout_reg[27]/P0001 ,
		\u12_o8_we_reg/P0001 ,
		\u7_wp_reg[0]/P0001 ,
		\u7_wp_reg[1]/NET0131 ,
		_w5798_
	);
	LUT2 #(
		.INIT('he)
	) name3652 (
		_w5797_,
		_w5798_,
		_w5799_
	);
	LUT4 #(
		.INIT('h4ccc)
	) name3653 (
		\u12_o8_we_reg/P0001 ,
		\u7_mem_reg[3][28]/NET0131 ,
		\u7_wp_reg[0]/P0001 ,
		\u7_wp_reg[1]/NET0131 ,
		_w5800_
	);
	LUT4 #(
		.INIT('h8000)
	) name3654 (
		\u12_dout_reg[28]/P0001 ,
		\u12_o8_we_reg/P0001 ,
		\u7_wp_reg[0]/P0001 ,
		\u7_wp_reg[1]/NET0131 ,
		_w5801_
	);
	LUT2 #(
		.INIT('he)
	) name3655 (
		_w5800_,
		_w5801_,
		_w5802_
	);
	LUT4 #(
		.INIT('h4ccc)
	) name3656 (
		\u12_o8_we_reg/P0001 ,
		\u7_mem_reg[3][29]/NET0131 ,
		\u7_wp_reg[0]/P0001 ,
		\u7_wp_reg[1]/NET0131 ,
		_w5803_
	);
	LUT4 #(
		.INIT('h8000)
	) name3657 (
		\u12_dout_reg[29]/P0001 ,
		\u12_o8_we_reg/P0001 ,
		\u7_wp_reg[0]/P0001 ,
		\u7_wp_reg[1]/NET0131 ,
		_w5804_
	);
	LUT2 #(
		.INIT('he)
	) name3658 (
		_w5803_,
		_w5804_,
		_w5805_
	);
	LUT4 #(
		.INIT('h4ccc)
	) name3659 (
		\u12_o8_we_reg/P0001 ,
		\u7_mem_reg[3][2]/NET0131 ,
		\u7_wp_reg[0]/P0001 ,
		\u7_wp_reg[1]/NET0131 ,
		_w5806_
	);
	LUT4 #(
		.INIT('h8000)
	) name3660 (
		\u12_dout_reg[2]/P0001 ,
		\u12_o8_we_reg/P0001 ,
		\u7_wp_reg[0]/P0001 ,
		\u7_wp_reg[1]/NET0131 ,
		_w5807_
	);
	LUT2 #(
		.INIT('he)
	) name3661 (
		_w5806_,
		_w5807_,
		_w5808_
	);
	LUT4 #(
		.INIT('h4ccc)
	) name3662 (
		\u12_o8_we_reg/P0001 ,
		\u7_mem_reg[3][30]/NET0131 ,
		\u7_wp_reg[0]/P0001 ,
		\u7_wp_reg[1]/NET0131 ,
		_w5809_
	);
	LUT4 #(
		.INIT('h8000)
	) name3663 (
		\u12_dout_reg[30]/P0001 ,
		\u12_o8_we_reg/P0001 ,
		\u7_wp_reg[0]/P0001 ,
		\u7_wp_reg[1]/NET0131 ,
		_w5810_
	);
	LUT2 #(
		.INIT('he)
	) name3664 (
		_w5809_,
		_w5810_,
		_w5811_
	);
	LUT4 #(
		.INIT('h4ccc)
	) name3665 (
		\u12_o8_we_reg/P0001 ,
		\u7_mem_reg[3][31]/NET0131 ,
		\u7_wp_reg[0]/P0001 ,
		\u7_wp_reg[1]/NET0131 ,
		_w5812_
	);
	LUT4 #(
		.INIT('h8000)
	) name3666 (
		\u12_dout_reg[31]/P0001 ,
		\u12_o8_we_reg/P0001 ,
		\u7_wp_reg[0]/P0001 ,
		\u7_wp_reg[1]/NET0131 ,
		_w5813_
	);
	LUT2 #(
		.INIT('he)
	) name3667 (
		_w5812_,
		_w5813_,
		_w5814_
	);
	LUT4 #(
		.INIT('h4ccc)
	) name3668 (
		\u12_o8_we_reg/P0001 ,
		\u7_mem_reg[3][3]/NET0131 ,
		\u7_wp_reg[0]/P0001 ,
		\u7_wp_reg[1]/NET0131 ,
		_w5815_
	);
	LUT4 #(
		.INIT('h8000)
	) name3669 (
		\u12_dout_reg[3]/P0001 ,
		\u12_o8_we_reg/P0001 ,
		\u7_wp_reg[0]/P0001 ,
		\u7_wp_reg[1]/NET0131 ,
		_w5816_
	);
	LUT2 #(
		.INIT('he)
	) name3670 (
		_w5815_,
		_w5816_,
		_w5817_
	);
	LUT4 #(
		.INIT('h4ccc)
	) name3671 (
		\u12_o8_we_reg/P0001 ,
		\u7_mem_reg[3][4]/NET0131 ,
		\u7_wp_reg[0]/P0001 ,
		\u7_wp_reg[1]/NET0131 ,
		_w5818_
	);
	LUT4 #(
		.INIT('h8000)
	) name3672 (
		\u12_dout_reg[4]/P0001 ,
		\u12_o8_we_reg/P0001 ,
		\u7_wp_reg[0]/P0001 ,
		\u7_wp_reg[1]/NET0131 ,
		_w5819_
	);
	LUT2 #(
		.INIT('he)
	) name3673 (
		_w5818_,
		_w5819_,
		_w5820_
	);
	LUT4 #(
		.INIT('h4ccc)
	) name3674 (
		\u12_o8_we_reg/P0001 ,
		\u7_mem_reg[3][5]/NET0131 ,
		\u7_wp_reg[0]/P0001 ,
		\u7_wp_reg[1]/NET0131 ,
		_w5821_
	);
	LUT4 #(
		.INIT('h8000)
	) name3675 (
		\u12_dout_reg[5]/P0001 ,
		\u12_o8_we_reg/P0001 ,
		\u7_wp_reg[0]/P0001 ,
		\u7_wp_reg[1]/NET0131 ,
		_w5822_
	);
	LUT2 #(
		.INIT('he)
	) name3676 (
		_w5821_,
		_w5822_,
		_w5823_
	);
	LUT4 #(
		.INIT('h4ccc)
	) name3677 (
		\u12_o8_we_reg/P0001 ,
		\u7_mem_reg[3][6]/NET0131 ,
		\u7_wp_reg[0]/P0001 ,
		\u7_wp_reg[1]/NET0131 ,
		_w5824_
	);
	LUT4 #(
		.INIT('h8000)
	) name3678 (
		\u12_dout_reg[6]/P0001 ,
		\u12_o8_we_reg/P0001 ,
		\u7_wp_reg[0]/P0001 ,
		\u7_wp_reg[1]/NET0131 ,
		_w5825_
	);
	LUT2 #(
		.INIT('he)
	) name3679 (
		_w5824_,
		_w5825_,
		_w5826_
	);
	LUT4 #(
		.INIT('h4ccc)
	) name3680 (
		\u12_o8_we_reg/P0001 ,
		\u7_mem_reg[3][7]/NET0131 ,
		\u7_wp_reg[0]/P0001 ,
		\u7_wp_reg[1]/NET0131 ,
		_w5827_
	);
	LUT4 #(
		.INIT('h8000)
	) name3681 (
		\u12_dout_reg[7]/P0001 ,
		\u12_o8_we_reg/P0001 ,
		\u7_wp_reg[0]/P0001 ,
		\u7_wp_reg[1]/NET0131 ,
		_w5828_
	);
	LUT2 #(
		.INIT('he)
	) name3682 (
		_w5827_,
		_w5828_,
		_w5829_
	);
	LUT4 #(
		.INIT('h4ccc)
	) name3683 (
		\u12_o8_we_reg/P0001 ,
		\u7_mem_reg[3][8]/NET0131 ,
		\u7_wp_reg[0]/P0001 ,
		\u7_wp_reg[1]/NET0131 ,
		_w5830_
	);
	LUT4 #(
		.INIT('h8000)
	) name3684 (
		\u12_dout_reg[8]/P0001 ,
		\u12_o8_we_reg/P0001 ,
		\u7_wp_reg[0]/P0001 ,
		\u7_wp_reg[1]/NET0131 ,
		_w5831_
	);
	LUT2 #(
		.INIT('he)
	) name3685 (
		_w5830_,
		_w5831_,
		_w5832_
	);
	LUT4 #(
		.INIT('h4ccc)
	) name3686 (
		\u12_o8_we_reg/P0001 ,
		\u7_mem_reg[3][9]/NET0131 ,
		\u7_wp_reg[0]/P0001 ,
		\u7_wp_reg[1]/NET0131 ,
		_w5833_
	);
	LUT4 #(
		.INIT('h8000)
	) name3687 (
		\u12_dout_reg[9]/P0001 ,
		\u12_o8_we_reg/P0001 ,
		\u7_wp_reg[0]/P0001 ,
		\u7_wp_reg[1]/NET0131 ,
		_w5834_
	);
	LUT2 #(
		.INIT('he)
	) name3688 (
		_w5833_,
		_w5834_,
		_w5835_
	);
	LUT4 #(
		.INIT('hc4cc)
	) name3689 (
		\u12_o3_we_reg/P0001 ,
		\u3_mem_reg[2][17]/NET0131 ,
		\u3_wp_reg[0]/P0001 ,
		\u3_wp_reg[1]/NET0131 ,
		_w5836_
	);
	LUT4 #(
		.INIT('h0800)
	) name3690 (
		\u12_dout_reg[17]/P0001 ,
		\u12_o3_we_reg/P0001 ,
		\u3_wp_reg[0]/P0001 ,
		\u3_wp_reg[1]/NET0131 ,
		_w5837_
	);
	LUT2 #(
		.INIT('he)
	) name3691 (
		_w5836_,
		_w5837_,
		_w5838_
	);
	LUT4 #(
		.INIT('hcc4c)
	) name3692 (
		\u12_o9_we_reg/P0001 ,
		\u8_mem_reg[1][0]/NET0131 ,
		\u8_wp_reg[0]/P0001 ,
		\u8_wp_reg[1]/NET0131 ,
		_w5839_
	);
	LUT4 #(
		.INIT('h0080)
	) name3693 (
		\u12_dout_reg[0]/P0001 ,
		\u12_o9_we_reg/P0001 ,
		\u8_wp_reg[0]/P0001 ,
		\u8_wp_reg[1]/NET0131 ,
		_w5840_
	);
	LUT2 #(
		.INIT('he)
	) name3694 (
		_w5839_,
		_w5840_,
		_w5841_
	);
	LUT4 #(
		.INIT('hcc4c)
	) name3695 (
		\u12_o9_we_reg/P0001 ,
		\u8_mem_reg[1][10]/NET0131 ,
		\u8_wp_reg[0]/P0001 ,
		\u8_wp_reg[1]/NET0131 ,
		_w5842_
	);
	LUT4 #(
		.INIT('h0080)
	) name3696 (
		\u12_dout_reg[10]/P0001 ,
		\u12_o9_we_reg/P0001 ,
		\u8_wp_reg[0]/P0001 ,
		\u8_wp_reg[1]/NET0131 ,
		_w5843_
	);
	LUT2 #(
		.INIT('he)
	) name3697 (
		_w5842_,
		_w5843_,
		_w5844_
	);
	LUT4 #(
		.INIT('hcc4c)
	) name3698 (
		\u12_o9_we_reg/P0001 ,
		\u8_mem_reg[1][11]/NET0131 ,
		\u8_wp_reg[0]/P0001 ,
		\u8_wp_reg[1]/NET0131 ,
		_w5845_
	);
	LUT4 #(
		.INIT('h0080)
	) name3699 (
		\u12_dout_reg[11]/P0001 ,
		\u12_o9_we_reg/P0001 ,
		\u8_wp_reg[0]/P0001 ,
		\u8_wp_reg[1]/NET0131 ,
		_w5846_
	);
	LUT2 #(
		.INIT('he)
	) name3700 (
		_w5845_,
		_w5846_,
		_w5847_
	);
	LUT4 #(
		.INIT('hcc4c)
	) name3701 (
		\u12_o9_we_reg/P0001 ,
		\u8_mem_reg[1][12]/NET0131 ,
		\u8_wp_reg[0]/P0001 ,
		\u8_wp_reg[1]/NET0131 ,
		_w5848_
	);
	LUT4 #(
		.INIT('h0080)
	) name3702 (
		\u12_dout_reg[12]/P0001 ,
		\u12_o9_we_reg/P0001 ,
		\u8_wp_reg[0]/P0001 ,
		\u8_wp_reg[1]/NET0131 ,
		_w5849_
	);
	LUT2 #(
		.INIT('he)
	) name3703 (
		_w5848_,
		_w5849_,
		_w5850_
	);
	LUT4 #(
		.INIT('hcc4c)
	) name3704 (
		\u12_o9_we_reg/P0001 ,
		\u8_mem_reg[1][13]/NET0131 ,
		\u8_wp_reg[0]/P0001 ,
		\u8_wp_reg[1]/NET0131 ,
		_w5851_
	);
	LUT4 #(
		.INIT('h0080)
	) name3705 (
		\u12_dout_reg[13]/P0001 ,
		\u12_o9_we_reg/P0001 ,
		\u8_wp_reg[0]/P0001 ,
		\u8_wp_reg[1]/NET0131 ,
		_w5852_
	);
	LUT2 #(
		.INIT('he)
	) name3706 (
		_w5851_,
		_w5852_,
		_w5853_
	);
	LUT4 #(
		.INIT('hcc4c)
	) name3707 (
		\u12_o9_we_reg/P0001 ,
		\u8_mem_reg[1][14]/NET0131 ,
		\u8_wp_reg[0]/P0001 ,
		\u8_wp_reg[1]/NET0131 ,
		_w5854_
	);
	LUT4 #(
		.INIT('h0080)
	) name3708 (
		\u12_dout_reg[14]/P0001 ,
		\u12_o9_we_reg/P0001 ,
		\u8_wp_reg[0]/P0001 ,
		\u8_wp_reg[1]/NET0131 ,
		_w5855_
	);
	LUT2 #(
		.INIT('he)
	) name3709 (
		_w5854_,
		_w5855_,
		_w5856_
	);
	LUT4 #(
		.INIT('hcc4c)
	) name3710 (
		\u12_o9_we_reg/P0001 ,
		\u8_mem_reg[1][15]/NET0131 ,
		\u8_wp_reg[0]/P0001 ,
		\u8_wp_reg[1]/NET0131 ,
		_w5857_
	);
	LUT4 #(
		.INIT('h0080)
	) name3711 (
		\u12_dout_reg[15]/P0001 ,
		\u12_o9_we_reg/P0001 ,
		\u8_wp_reg[0]/P0001 ,
		\u8_wp_reg[1]/NET0131 ,
		_w5858_
	);
	LUT2 #(
		.INIT('he)
	) name3712 (
		_w5857_,
		_w5858_,
		_w5859_
	);
	LUT4 #(
		.INIT('hcc4c)
	) name3713 (
		\u12_o9_we_reg/P0001 ,
		\u8_mem_reg[1][16]/NET0131 ,
		\u8_wp_reg[0]/P0001 ,
		\u8_wp_reg[1]/NET0131 ,
		_w5860_
	);
	LUT4 #(
		.INIT('h0080)
	) name3714 (
		\u12_dout_reg[16]/P0001 ,
		\u12_o9_we_reg/P0001 ,
		\u8_wp_reg[0]/P0001 ,
		\u8_wp_reg[1]/NET0131 ,
		_w5861_
	);
	LUT2 #(
		.INIT('he)
	) name3715 (
		_w5860_,
		_w5861_,
		_w5862_
	);
	LUT4 #(
		.INIT('hcc4c)
	) name3716 (
		\u12_o9_we_reg/P0001 ,
		\u8_mem_reg[1][17]/NET0131 ,
		\u8_wp_reg[0]/P0001 ,
		\u8_wp_reg[1]/NET0131 ,
		_w5863_
	);
	LUT4 #(
		.INIT('h0080)
	) name3717 (
		\u12_dout_reg[17]/P0001 ,
		\u12_o9_we_reg/P0001 ,
		\u8_wp_reg[0]/P0001 ,
		\u8_wp_reg[1]/NET0131 ,
		_w5864_
	);
	LUT2 #(
		.INIT('he)
	) name3718 (
		_w5863_,
		_w5864_,
		_w5865_
	);
	LUT4 #(
		.INIT('hcc4c)
	) name3719 (
		\u12_o9_we_reg/P0001 ,
		\u8_mem_reg[1][18]/NET0131 ,
		\u8_wp_reg[0]/P0001 ,
		\u8_wp_reg[1]/NET0131 ,
		_w5866_
	);
	LUT4 #(
		.INIT('h0080)
	) name3720 (
		\u12_dout_reg[18]/P0001 ,
		\u12_o9_we_reg/P0001 ,
		\u8_wp_reg[0]/P0001 ,
		\u8_wp_reg[1]/NET0131 ,
		_w5867_
	);
	LUT2 #(
		.INIT('he)
	) name3721 (
		_w5866_,
		_w5867_,
		_w5868_
	);
	LUT4 #(
		.INIT('hcc4c)
	) name3722 (
		\u12_o9_we_reg/P0001 ,
		\u8_mem_reg[1][19]/NET0131 ,
		\u8_wp_reg[0]/P0001 ,
		\u8_wp_reg[1]/NET0131 ,
		_w5869_
	);
	LUT4 #(
		.INIT('h0080)
	) name3723 (
		\u12_dout_reg[19]/P0001 ,
		\u12_o9_we_reg/P0001 ,
		\u8_wp_reg[0]/P0001 ,
		\u8_wp_reg[1]/NET0131 ,
		_w5870_
	);
	LUT2 #(
		.INIT('he)
	) name3724 (
		_w5869_,
		_w5870_,
		_w5871_
	);
	LUT4 #(
		.INIT('hcc4c)
	) name3725 (
		\u12_o9_we_reg/P0001 ,
		\u8_mem_reg[1][1]/NET0131 ,
		\u8_wp_reg[0]/P0001 ,
		\u8_wp_reg[1]/NET0131 ,
		_w5872_
	);
	LUT4 #(
		.INIT('h0080)
	) name3726 (
		\u12_dout_reg[1]/P0001 ,
		\u12_o9_we_reg/P0001 ,
		\u8_wp_reg[0]/P0001 ,
		\u8_wp_reg[1]/NET0131 ,
		_w5873_
	);
	LUT2 #(
		.INIT('he)
	) name3727 (
		_w5872_,
		_w5873_,
		_w5874_
	);
	LUT4 #(
		.INIT('hcc4c)
	) name3728 (
		\u12_o9_we_reg/P0001 ,
		\u8_mem_reg[1][20]/NET0131 ,
		\u8_wp_reg[0]/P0001 ,
		\u8_wp_reg[1]/NET0131 ,
		_w5875_
	);
	LUT4 #(
		.INIT('h0080)
	) name3729 (
		\u12_dout_reg[20]/P0001 ,
		\u12_o9_we_reg/P0001 ,
		\u8_wp_reg[0]/P0001 ,
		\u8_wp_reg[1]/NET0131 ,
		_w5876_
	);
	LUT2 #(
		.INIT('he)
	) name3730 (
		_w5875_,
		_w5876_,
		_w5877_
	);
	LUT4 #(
		.INIT('hcc4c)
	) name3731 (
		\u12_o9_we_reg/P0001 ,
		\u8_mem_reg[1][21]/NET0131 ,
		\u8_wp_reg[0]/P0001 ,
		\u8_wp_reg[1]/NET0131 ,
		_w5878_
	);
	LUT4 #(
		.INIT('h0080)
	) name3732 (
		\u12_dout_reg[21]/P0001 ,
		\u12_o9_we_reg/P0001 ,
		\u8_wp_reg[0]/P0001 ,
		\u8_wp_reg[1]/NET0131 ,
		_w5879_
	);
	LUT2 #(
		.INIT('he)
	) name3733 (
		_w5878_,
		_w5879_,
		_w5880_
	);
	LUT4 #(
		.INIT('hcc4c)
	) name3734 (
		\u12_o9_we_reg/P0001 ,
		\u8_mem_reg[1][22]/NET0131 ,
		\u8_wp_reg[0]/P0001 ,
		\u8_wp_reg[1]/NET0131 ,
		_w5881_
	);
	LUT4 #(
		.INIT('h0080)
	) name3735 (
		\u12_dout_reg[22]/P0001 ,
		\u12_o9_we_reg/P0001 ,
		\u8_wp_reg[0]/P0001 ,
		\u8_wp_reg[1]/NET0131 ,
		_w5882_
	);
	LUT2 #(
		.INIT('he)
	) name3736 (
		_w5881_,
		_w5882_,
		_w5883_
	);
	LUT4 #(
		.INIT('hcc4c)
	) name3737 (
		\u12_o9_we_reg/P0001 ,
		\u8_mem_reg[1][23]/NET0131 ,
		\u8_wp_reg[0]/P0001 ,
		\u8_wp_reg[1]/NET0131 ,
		_w5884_
	);
	LUT4 #(
		.INIT('h0080)
	) name3738 (
		\u12_dout_reg[23]/P0001 ,
		\u12_o9_we_reg/P0001 ,
		\u8_wp_reg[0]/P0001 ,
		\u8_wp_reg[1]/NET0131 ,
		_w5885_
	);
	LUT2 #(
		.INIT('he)
	) name3739 (
		_w5884_,
		_w5885_,
		_w5886_
	);
	LUT4 #(
		.INIT('hcc4c)
	) name3740 (
		\u12_o9_we_reg/P0001 ,
		\u8_mem_reg[1][24]/NET0131 ,
		\u8_wp_reg[0]/P0001 ,
		\u8_wp_reg[1]/NET0131 ,
		_w5887_
	);
	LUT4 #(
		.INIT('h0080)
	) name3741 (
		\u12_dout_reg[24]/P0001 ,
		\u12_o9_we_reg/P0001 ,
		\u8_wp_reg[0]/P0001 ,
		\u8_wp_reg[1]/NET0131 ,
		_w5888_
	);
	LUT2 #(
		.INIT('he)
	) name3742 (
		_w5887_,
		_w5888_,
		_w5889_
	);
	LUT4 #(
		.INIT('hcc4c)
	) name3743 (
		\u12_o9_we_reg/P0001 ,
		\u8_mem_reg[1][25]/NET0131 ,
		\u8_wp_reg[0]/P0001 ,
		\u8_wp_reg[1]/NET0131 ,
		_w5890_
	);
	LUT4 #(
		.INIT('h0080)
	) name3744 (
		\u12_dout_reg[25]/P0001 ,
		\u12_o9_we_reg/P0001 ,
		\u8_wp_reg[0]/P0001 ,
		\u8_wp_reg[1]/NET0131 ,
		_w5891_
	);
	LUT2 #(
		.INIT('he)
	) name3745 (
		_w5890_,
		_w5891_,
		_w5892_
	);
	LUT4 #(
		.INIT('hcc4c)
	) name3746 (
		\u12_o3_we_reg/P0001 ,
		\u3_mem_reg[1][0]/NET0131 ,
		\u3_wp_reg[0]/P0001 ,
		\u3_wp_reg[1]/NET0131 ,
		_w5893_
	);
	LUT4 #(
		.INIT('h0080)
	) name3747 (
		\u12_dout_reg[0]/P0001 ,
		\u12_o3_we_reg/P0001 ,
		\u3_wp_reg[0]/P0001 ,
		\u3_wp_reg[1]/NET0131 ,
		_w5894_
	);
	LUT2 #(
		.INIT('he)
	) name3748 (
		_w5893_,
		_w5894_,
		_w5895_
	);
	LUT4 #(
		.INIT('hcc4c)
	) name3749 (
		\u12_o9_we_reg/P0001 ,
		\u8_mem_reg[1][26]/NET0131 ,
		\u8_wp_reg[0]/P0001 ,
		\u8_wp_reg[1]/NET0131 ,
		_w5896_
	);
	LUT4 #(
		.INIT('h0080)
	) name3750 (
		\u12_dout_reg[26]/P0001 ,
		\u12_o9_we_reg/P0001 ,
		\u8_wp_reg[0]/P0001 ,
		\u8_wp_reg[1]/NET0131 ,
		_w5897_
	);
	LUT2 #(
		.INIT('he)
	) name3751 (
		_w5896_,
		_w5897_,
		_w5898_
	);
	LUT4 #(
		.INIT('hcc4c)
	) name3752 (
		\u12_o9_we_reg/P0001 ,
		\u8_mem_reg[1][27]/NET0131 ,
		\u8_wp_reg[0]/P0001 ,
		\u8_wp_reg[1]/NET0131 ,
		_w5899_
	);
	LUT4 #(
		.INIT('h0080)
	) name3753 (
		\u12_dout_reg[27]/P0001 ,
		\u12_o9_we_reg/P0001 ,
		\u8_wp_reg[0]/P0001 ,
		\u8_wp_reg[1]/NET0131 ,
		_w5900_
	);
	LUT2 #(
		.INIT('he)
	) name3754 (
		_w5899_,
		_w5900_,
		_w5901_
	);
	LUT4 #(
		.INIT('hcc4c)
	) name3755 (
		\u12_o3_we_reg/P0001 ,
		\u3_mem_reg[1][10]/NET0131 ,
		\u3_wp_reg[0]/P0001 ,
		\u3_wp_reg[1]/NET0131 ,
		_w5902_
	);
	LUT4 #(
		.INIT('h0080)
	) name3756 (
		\u12_dout_reg[10]/P0001 ,
		\u12_o3_we_reg/P0001 ,
		\u3_wp_reg[0]/P0001 ,
		\u3_wp_reg[1]/NET0131 ,
		_w5903_
	);
	LUT2 #(
		.INIT('he)
	) name3757 (
		_w5902_,
		_w5903_,
		_w5904_
	);
	LUT4 #(
		.INIT('hcc4c)
	) name3758 (
		\u12_o9_we_reg/P0001 ,
		\u8_mem_reg[1][29]/NET0131 ,
		\u8_wp_reg[0]/P0001 ,
		\u8_wp_reg[1]/NET0131 ,
		_w5905_
	);
	LUT4 #(
		.INIT('h0080)
	) name3759 (
		\u12_dout_reg[29]/P0001 ,
		\u12_o9_we_reg/P0001 ,
		\u8_wp_reg[0]/P0001 ,
		\u8_wp_reg[1]/NET0131 ,
		_w5906_
	);
	LUT2 #(
		.INIT('he)
	) name3760 (
		_w5905_,
		_w5906_,
		_w5907_
	);
	LUT4 #(
		.INIT('hcc4c)
	) name3761 (
		\u12_o3_we_reg/P0001 ,
		\u3_mem_reg[1][11]/NET0131 ,
		\u3_wp_reg[0]/P0001 ,
		\u3_wp_reg[1]/NET0131 ,
		_w5908_
	);
	LUT4 #(
		.INIT('h0080)
	) name3762 (
		\u12_dout_reg[11]/P0001 ,
		\u12_o3_we_reg/P0001 ,
		\u3_wp_reg[0]/P0001 ,
		\u3_wp_reg[1]/NET0131 ,
		_w5909_
	);
	LUT2 #(
		.INIT('he)
	) name3763 (
		_w5908_,
		_w5909_,
		_w5910_
	);
	LUT4 #(
		.INIT('hcc4c)
	) name3764 (
		\u12_o9_we_reg/P0001 ,
		\u8_mem_reg[1][2]/NET0131 ,
		\u8_wp_reg[0]/P0001 ,
		\u8_wp_reg[1]/NET0131 ,
		_w5911_
	);
	LUT4 #(
		.INIT('h0080)
	) name3765 (
		\u12_dout_reg[2]/P0001 ,
		\u12_o9_we_reg/P0001 ,
		\u8_wp_reg[0]/P0001 ,
		\u8_wp_reg[1]/NET0131 ,
		_w5912_
	);
	LUT2 #(
		.INIT('he)
	) name3766 (
		_w5911_,
		_w5912_,
		_w5913_
	);
	LUT4 #(
		.INIT('hcc4c)
	) name3767 (
		\u12_o9_we_reg/P0001 ,
		\u8_mem_reg[1][30]/NET0131 ,
		\u8_wp_reg[0]/P0001 ,
		\u8_wp_reg[1]/NET0131 ,
		_w5914_
	);
	LUT4 #(
		.INIT('h0080)
	) name3768 (
		\u12_dout_reg[30]/P0001 ,
		\u12_o9_we_reg/P0001 ,
		\u8_wp_reg[0]/P0001 ,
		\u8_wp_reg[1]/NET0131 ,
		_w5915_
	);
	LUT2 #(
		.INIT('he)
	) name3769 (
		_w5914_,
		_w5915_,
		_w5916_
	);
	LUT4 #(
		.INIT('hcc4c)
	) name3770 (
		\u12_o3_we_reg/P0001 ,
		\u3_mem_reg[1][12]/NET0131 ,
		\u3_wp_reg[0]/P0001 ,
		\u3_wp_reg[1]/NET0131 ,
		_w5917_
	);
	LUT4 #(
		.INIT('h0080)
	) name3771 (
		\u12_dout_reg[12]/P0001 ,
		\u12_o3_we_reg/P0001 ,
		\u3_wp_reg[0]/P0001 ,
		\u3_wp_reg[1]/NET0131 ,
		_w5918_
	);
	LUT2 #(
		.INIT('he)
	) name3772 (
		_w5917_,
		_w5918_,
		_w5919_
	);
	LUT4 #(
		.INIT('h4ccc)
	) name3773 (
		\u12_o9_we_reg/P0001 ,
		\u8_mem_reg[3][11]/NET0131 ,
		\u8_wp_reg[0]/P0001 ,
		\u8_wp_reg[1]/NET0131 ,
		_w5920_
	);
	LUT4 #(
		.INIT('h8000)
	) name3774 (
		\u12_dout_reg[11]/P0001 ,
		\u12_o9_we_reg/P0001 ,
		\u8_wp_reg[0]/P0001 ,
		\u8_wp_reg[1]/NET0131 ,
		_w5921_
	);
	LUT2 #(
		.INIT('he)
	) name3775 (
		_w5920_,
		_w5921_,
		_w5922_
	);
	LUT4 #(
		.INIT('hcc4c)
	) name3776 (
		\u12_o9_we_reg/P0001 ,
		\u8_mem_reg[1][3]/NET0131 ,
		\u8_wp_reg[0]/P0001 ,
		\u8_wp_reg[1]/NET0131 ,
		_w5923_
	);
	LUT4 #(
		.INIT('h0080)
	) name3777 (
		\u12_dout_reg[3]/P0001 ,
		\u12_o9_we_reg/P0001 ,
		\u8_wp_reg[0]/P0001 ,
		\u8_wp_reg[1]/NET0131 ,
		_w5924_
	);
	LUT2 #(
		.INIT('he)
	) name3778 (
		_w5923_,
		_w5924_,
		_w5925_
	);
	LUT4 #(
		.INIT('hcc4c)
	) name3779 (
		\u12_o3_we_reg/P0001 ,
		\u3_mem_reg[1][13]/NET0131 ,
		\u3_wp_reg[0]/P0001 ,
		\u3_wp_reg[1]/NET0131 ,
		_w5926_
	);
	LUT4 #(
		.INIT('h0080)
	) name3780 (
		\u12_dout_reg[13]/P0001 ,
		\u12_o3_we_reg/P0001 ,
		\u3_wp_reg[0]/P0001 ,
		\u3_wp_reg[1]/NET0131 ,
		_w5927_
	);
	LUT2 #(
		.INIT('he)
	) name3781 (
		_w5926_,
		_w5927_,
		_w5928_
	);
	LUT4 #(
		.INIT('hcc4c)
	) name3782 (
		\u12_o9_we_reg/P0001 ,
		\u8_mem_reg[1][5]/NET0131 ,
		\u8_wp_reg[0]/P0001 ,
		\u8_wp_reg[1]/NET0131 ,
		_w5929_
	);
	LUT4 #(
		.INIT('h0080)
	) name3783 (
		\u12_dout_reg[5]/P0001 ,
		\u12_o9_we_reg/P0001 ,
		\u8_wp_reg[0]/P0001 ,
		\u8_wp_reg[1]/NET0131 ,
		_w5930_
	);
	LUT2 #(
		.INIT('he)
	) name3784 (
		_w5929_,
		_w5930_,
		_w5931_
	);
	LUT4 #(
		.INIT('hcc4c)
	) name3785 (
		\u12_o9_we_reg/P0001 ,
		\u8_mem_reg[1][7]/NET0131 ,
		\u8_wp_reg[0]/P0001 ,
		\u8_wp_reg[1]/NET0131 ,
		_w5932_
	);
	LUT4 #(
		.INIT('h0080)
	) name3786 (
		\u12_dout_reg[7]/P0001 ,
		\u12_o9_we_reg/P0001 ,
		\u8_wp_reg[0]/P0001 ,
		\u8_wp_reg[1]/NET0131 ,
		_w5933_
	);
	LUT2 #(
		.INIT('he)
	) name3787 (
		_w5932_,
		_w5933_,
		_w5934_
	);
	LUT4 #(
		.INIT('hcc4c)
	) name3788 (
		\u12_o3_we_reg/P0001 ,
		\u3_mem_reg[1][15]/NET0131 ,
		\u3_wp_reg[0]/P0001 ,
		\u3_wp_reg[1]/NET0131 ,
		_w5935_
	);
	LUT4 #(
		.INIT('h0080)
	) name3789 (
		\u12_dout_reg[15]/P0001 ,
		\u12_o3_we_reg/P0001 ,
		\u3_wp_reg[0]/P0001 ,
		\u3_wp_reg[1]/NET0131 ,
		_w5936_
	);
	LUT2 #(
		.INIT('he)
	) name3790 (
		_w5935_,
		_w5936_,
		_w5937_
	);
	LUT4 #(
		.INIT('hcc4c)
	) name3791 (
		\u12_o9_we_reg/P0001 ,
		\u8_mem_reg[1][8]/NET0131 ,
		\u8_wp_reg[0]/P0001 ,
		\u8_wp_reg[1]/NET0131 ,
		_w5938_
	);
	LUT4 #(
		.INIT('h0080)
	) name3792 (
		\u12_dout_reg[8]/P0001 ,
		\u12_o9_we_reg/P0001 ,
		\u8_wp_reg[0]/P0001 ,
		\u8_wp_reg[1]/NET0131 ,
		_w5939_
	);
	LUT2 #(
		.INIT('he)
	) name3793 (
		_w5938_,
		_w5939_,
		_w5940_
	);
	LUT4 #(
		.INIT('hcc4c)
	) name3794 (
		\u12_o9_we_reg/P0001 ,
		\u8_mem_reg[1][9]/NET0131 ,
		\u8_wp_reg[0]/P0001 ,
		\u8_wp_reg[1]/NET0131 ,
		_w5941_
	);
	LUT4 #(
		.INIT('h0080)
	) name3795 (
		\u12_dout_reg[9]/P0001 ,
		\u12_o9_we_reg/P0001 ,
		\u8_wp_reg[0]/P0001 ,
		\u8_wp_reg[1]/NET0131 ,
		_w5942_
	);
	LUT2 #(
		.INIT('he)
	) name3796 (
		_w5941_,
		_w5942_,
		_w5943_
	);
	LUT4 #(
		.INIT('hcc4c)
	) name3797 (
		\u12_o3_we_reg/P0001 ,
		\u3_mem_reg[1][16]/NET0131 ,
		\u3_wp_reg[0]/P0001 ,
		\u3_wp_reg[1]/NET0131 ,
		_w5944_
	);
	LUT4 #(
		.INIT('h0080)
	) name3798 (
		\u12_dout_reg[16]/P0001 ,
		\u12_o3_we_reg/P0001 ,
		\u3_wp_reg[0]/P0001 ,
		\u3_wp_reg[1]/NET0131 ,
		_w5945_
	);
	LUT2 #(
		.INIT('he)
	) name3799 (
		_w5944_,
		_w5945_,
		_w5946_
	);
	LUT4 #(
		.INIT('hc4cc)
	) name3800 (
		\u12_o9_we_reg/P0001 ,
		\u8_mem_reg[2][0]/NET0131 ,
		\u8_wp_reg[0]/P0001 ,
		\u8_wp_reg[1]/NET0131 ,
		_w5947_
	);
	LUT4 #(
		.INIT('h0800)
	) name3801 (
		\u12_dout_reg[0]/P0001 ,
		\u12_o9_we_reg/P0001 ,
		\u8_wp_reg[0]/P0001 ,
		\u8_wp_reg[1]/NET0131 ,
		_w5948_
	);
	LUT2 #(
		.INIT('he)
	) name3802 (
		_w5947_,
		_w5948_,
		_w5949_
	);
	LUT4 #(
		.INIT('hc4cc)
	) name3803 (
		\u12_o9_we_reg/P0001 ,
		\u8_mem_reg[2][10]/NET0131 ,
		\u8_wp_reg[0]/P0001 ,
		\u8_wp_reg[1]/NET0131 ,
		_w5950_
	);
	LUT4 #(
		.INIT('h0800)
	) name3804 (
		\u12_dout_reg[10]/P0001 ,
		\u12_o9_we_reg/P0001 ,
		\u8_wp_reg[0]/P0001 ,
		\u8_wp_reg[1]/NET0131 ,
		_w5951_
	);
	LUT2 #(
		.INIT('he)
	) name3805 (
		_w5950_,
		_w5951_,
		_w5952_
	);
	LUT4 #(
		.INIT('hcc4c)
	) name3806 (
		\u12_o3_we_reg/P0001 ,
		\u3_mem_reg[1][17]/NET0131 ,
		\u3_wp_reg[0]/P0001 ,
		\u3_wp_reg[1]/NET0131 ,
		_w5953_
	);
	LUT4 #(
		.INIT('h0080)
	) name3807 (
		\u12_dout_reg[17]/P0001 ,
		\u12_o3_we_reg/P0001 ,
		\u3_wp_reg[0]/P0001 ,
		\u3_wp_reg[1]/NET0131 ,
		_w5954_
	);
	LUT2 #(
		.INIT('he)
	) name3808 (
		_w5953_,
		_w5954_,
		_w5955_
	);
	LUT4 #(
		.INIT('hc4cc)
	) name3809 (
		\u12_o9_we_reg/P0001 ,
		\u8_mem_reg[2][11]/NET0131 ,
		\u8_wp_reg[0]/P0001 ,
		\u8_wp_reg[1]/NET0131 ,
		_w5956_
	);
	LUT4 #(
		.INIT('h0800)
	) name3810 (
		\u12_dout_reg[11]/P0001 ,
		\u12_o9_we_reg/P0001 ,
		\u8_wp_reg[0]/P0001 ,
		\u8_wp_reg[1]/NET0131 ,
		_w5957_
	);
	LUT2 #(
		.INIT('he)
	) name3811 (
		_w5956_,
		_w5957_,
		_w5958_
	);
	LUT4 #(
		.INIT('hc4cc)
	) name3812 (
		\u12_o9_we_reg/P0001 ,
		\u8_mem_reg[2][12]/NET0131 ,
		\u8_wp_reg[0]/P0001 ,
		\u8_wp_reg[1]/NET0131 ,
		_w5959_
	);
	LUT4 #(
		.INIT('h0800)
	) name3813 (
		\u12_dout_reg[12]/P0001 ,
		\u12_o9_we_reg/P0001 ,
		\u8_wp_reg[0]/P0001 ,
		\u8_wp_reg[1]/NET0131 ,
		_w5960_
	);
	LUT2 #(
		.INIT('he)
	) name3814 (
		_w5959_,
		_w5960_,
		_w5961_
	);
	LUT4 #(
		.INIT('hcc4c)
	) name3815 (
		\u12_o3_we_reg/P0001 ,
		\u3_mem_reg[1][18]/NET0131 ,
		\u3_wp_reg[0]/P0001 ,
		\u3_wp_reg[1]/NET0131 ,
		_w5962_
	);
	LUT4 #(
		.INIT('h0080)
	) name3816 (
		\u12_dout_reg[18]/P0001 ,
		\u12_o3_we_reg/P0001 ,
		\u3_wp_reg[0]/P0001 ,
		\u3_wp_reg[1]/NET0131 ,
		_w5963_
	);
	LUT2 #(
		.INIT('he)
	) name3817 (
		_w5962_,
		_w5963_,
		_w5964_
	);
	LUT4 #(
		.INIT('hc4cc)
	) name3818 (
		\u12_o9_we_reg/P0001 ,
		\u8_mem_reg[2][13]/NET0131 ,
		\u8_wp_reg[0]/P0001 ,
		\u8_wp_reg[1]/NET0131 ,
		_w5965_
	);
	LUT4 #(
		.INIT('h0800)
	) name3819 (
		\u12_dout_reg[13]/P0001 ,
		\u12_o9_we_reg/P0001 ,
		\u8_wp_reg[0]/P0001 ,
		\u8_wp_reg[1]/NET0131 ,
		_w5966_
	);
	LUT2 #(
		.INIT('he)
	) name3820 (
		_w5965_,
		_w5966_,
		_w5967_
	);
	LUT4 #(
		.INIT('hc4cc)
	) name3821 (
		\u12_o9_we_reg/P0001 ,
		\u8_mem_reg[2][14]/NET0131 ,
		\u8_wp_reg[0]/P0001 ,
		\u8_wp_reg[1]/NET0131 ,
		_w5968_
	);
	LUT4 #(
		.INIT('h0800)
	) name3822 (
		\u12_dout_reg[14]/P0001 ,
		\u12_o9_we_reg/P0001 ,
		\u8_wp_reg[0]/P0001 ,
		\u8_wp_reg[1]/NET0131 ,
		_w5969_
	);
	LUT2 #(
		.INIT('he)
	) name3823 (
		_w5968_,
		_w5969_,
		_w5970_
	);
	LUT4 #(
		.INIT('hcc4c)
	) name3824 (
		\u12_o3_we_reg/P0001 ,
		\u3_mem_reg[1][19]/NET0131 ,
		\u3_wp_reg[0]/P0001 ,
		\u3_wp_reg[1]/NET0131 ,
		_w5971_
	);
	LUT4 #(
		.INIT('h0080)
	) name3825 (
		\u12_dout_reg[19]/P0001 ,
		\u12_o3_we_reg/P0001 ,
		\u3_wp_reg[0]/P0001 ,
		\u3_wp_reg[1]/NET0131 ,
		_w5972_
	);
	LUT2 #(
		.INIT('he)
	) name3826 (
		_w5971_,
		_w5972_,
		_w5973_
	);
	LUT4 #(
		.INIT('hc4cc)
	) name3827 (
		\u12_o9_we_reg/P0001 ,
		\u8_mem_reg[2][15]/NET0131 ,
		\u8_wp_reg[0]/P0001 ,
		\u8_wp_reg[1]/NET0131 ,
		_w5974_
	);
	LUT4 #(
		.INIT('h0800)
	) name3828 (
		\u12_dout_reg[15]/P0001 ,
		\u12_o9_we_reg/P0001 ,
		\u8_wp_reg[0]/P0001 ,
		\u8_wp_reg[1]/NET0131 ,
		_w5975_
	);
	LUT2 #(
		.INIT('he)
	) name3829 (
		_w5974_,
		_w5975_,
		_w5976_
	);
	LUT4 #(
		.INIT('hc4cc)
	) name3830 (
		\u12_o9_we_reg/P0001 ,
		\u8_mem_reg[2][16]/NET0131 ,
		\u8_wp_reg[0]/P0001 ,
		\u8_wp_reg[1]/NET0131 ,
		_w5977_
	);
	LUT4 #(
		.INIT('h0800)
	) name3831 (
		\u12_dout_reg[16]/P0001 ,
		\u12_o9_we_reg/P0001 ,
		\u8_wp_reg[0]/P0001 ,
		\u8_wp_reg[1]/NET0131 ,
		_w5978_
	);
	LUT2 #(
		.INIT('he)
	) name3832 (
		_w5977_,
		_w5978_,
		_w5979_
	);
	LUT4 #(
		.INIT('hc4cc)
	) name3833 (
		\u12_o9_we_reg/P0001 ,
		\u8_mem_reg[2][17]/NET0131 ,
		\u8_wp_reg[0]/P0001 ,
		\u8_wp_reg[1]/NET0131 ,
		_w5980_
	);
	LUT4 #(
		.INIT('h0800)
	) name3834 (
		\u12_dout_reg[17]/P0001 ,
		\u12_o9_we_reg/P0001 ,
		\u8_wp_reg[0]/P0001 ,
		\u8_wp_reg[1]/NET0131 ,
		_w5981_
	);
	LUT2 #(
		.INIT('he)
	) name3835 (
		_w5980_,
		_w5981_,
		_w5982_
	);
	LUT4 #(
		.INIT('hc4cc)
	) name3836 (
		\u12_o9_we_reg/P0001 ,
		\u8_mem_reg[2][18]/NET0131 ,
		\u8_wp_reg[0]/P0001 ,
		\u8_wp_reg[1]/NET0131 ,
		_w5983_
	);
	LUT4 #(
		.INIT('h0800)
	) name3837 (
		\u12_dout_reg[18]/P0001 ,
		\u12_o9_we_reg/P0001 ,
		\u8_wp_reg[0]/P0001 ,
		\u8_wp_reg[1]/NET0131 ,
		_w5984_
	);
	LUT2 #(
		.INIT('he)
	) name3838 (
		_w5983_,
		_w5984_,
		_w5985_
	);
	LUT4 #(
		.INIT('hcc4c)
	) name3839 (
		\u12_o3_we_reg/P0001 ,
		\u3_mem_reg[1][20]/NET0131 ,
		\u3_wp_reg[0]/P0001 ,
		\u3_wp_reg[1]/NET0131 ,
		_w5986_
	);
	LUT4 #(
		.INIT('h0080)
	) name3840 (
		\u12_dout_reg[20]/P0001 ,
		\u12_o3_we_reg/P0001 ,
		\u3_wp_reg[0]/P0001 ,
		\u3_wp_reg[1]/NET0131 ,
		_w5987_
	);
	LUT2 #(
		.INIT('he)
	) name3841 (
		_w5986_,
		_w5987_,
		_w5988_
	);
	LUT4 #(
		.INIT('hc4cc)
	) name3842 (
		\u12_o9_we_reg/P0001 ,
		\u8_mem_reg[2][19]/NET0131 ,
		\u8_wp_reg[0]/P0001 ,
		\u8_wp_reg[1]/NET0131 ,
		_w5989_
	);
	LUT4 #(
		.INIT('h0800)
	) name3843 (
		\u12_dout_reg[19]/P0001 ,
		\u12_o9_we_reg/P0001 ,
		\u8_wp_reg[0]/P0001 ,
		\u8_wp_reg[1]/NET0131 ,
		_w5990_
	);
	LUT2 #(
		.INIT('he)
	) name3844 (
		_w5989_,
		_w5990_,
		_w5991_
	);
	LUT4 #(
		.INIT('hc4cc)
	) name3845 (
		\u12_o9_we_reg/P0001 ,
		\u8_mem_reg[2][1]/NET0131 ,
		\u8_wp_reg[0]/P0001 ,
		\u8_wp_reg[1]/NET0131 ,
		_w5992_
	);
	LUT4 #(
		.INIT('h0800)
	) name3846 (
		\u12_dout_reg[1]/P0001 ,
		\u12_o9_we_reg/P0001 ,
		\u8_wp_reg[0]/P0001 ,
		\u8_wp_reg[1]/NET0131 ,
		_w5993_
	);
	LUT2 #(
		.INIT('he)
	) name3847 (
		_w5992_,
		_w5993_,
		_w5994_
	);
	LUT4 #(
		.INIT('hcc4c)
	) name3848 (
		\u12_o3_we_reg/P0001 ,
		\u3_mem_reg[1][21]/NET0131 ,
		\u3_wp_reg[0]/P0001 ,
		\u3_wp_reg[1]/NET0131 ,
		_w5995_
	);
	LUT4 #(
		.INIT('h0080)
	) name3849 (
		\u12_dout_reg[21]/P0001 ,
		\u12_o3_we_reg/P0001 ,
		\u3_wp_reg[0]/P0001 ,
		\u3_wp_reg[1]/NET0131 ,
		_w5996_
	);
	LUT2 #(
		.INIT('he)
	) name3850 (
		_w5995_,
		_w5996_,
		_w5997_
	);
	LUT4 #(
		.INIT('hc4cc)
	) name3851 (
		\u12_o9_we_reg/P0001 ,
		\u8_mem_reg[2][20]/NET0131 ,
		\u8_wp_reg[0]/P0001 ,
		\u8_wp_reg[1]/NET0131 ,
		_w5998_
	);
	LUT4 #(
		.INIT('h0800)
	) name3852 (
		\u12_dout_reg[20]/P0001 ,
		\u12_o9_we_reg/P0001 ,
		\u8_wp_reg[0]/P0001 ,
		\u8_wp_reg[1]/NET0131 ,
		_w5999_
	);
	LUT2 #(
		.INIT('he)
	) name3853 (
		_w5998_,
		_w5999_,
		_w6000_
	);
	LUT4 #(
		.INIT('hc4cc)
	) name3854 (
		\u12_o9_we_reg/P0001 ,
		\u8_mem_reg[2][21]/NET0131 ,
		\u8_wp_reg[0]/P0001 ,
		\u8_wp_reg[1]/NET0131 ,
		_w6001_
	);
	LUT4 #(
		.INIT('h0800)
	) name3855 (
		\u12_dout_reg[21]/P0001 ,
		\u12_o9_we_reg/P0001 ,
		\u8_wp_reg[0]/P0001 ,
		\u8_wp_reg[1]/NET0131 ,
		_w6002_
	);
	LUT2 #(
		.INIT('he)
	) name3856 (
		_w6001_,
		_w6002_,
		_w6003_
	);
	LUT4 #(
		.INIT('hcc4c)
	) name3857 (
		\u12_o3_we_reg/P0001 ,
		\u3_mem_reg[1][22]/NET0131 ,
		\u3_wp_reg[0]/P0001 ,
		\u3_wp_reg[1]/NET0131 ,
		_w6004_
	);
	LUT4 #(
		.INIT('h0080)
	) name3858 (
		\u12_dout_reg[22]/P0001 ,
		\u12_o3_we_reg/P0001 ,
		\u3_wp_reg[0]/P0001 ,
		\u3_wp_reg[1]/NET0131 ,
		_w6005_
	);
	LUT2 #(
		.INIT('he)
	) name3859 (
		_w6004_,
		_w6005_,
		_w6006_
	);
	LUT4 #(
		.INIT('hc4cc)
	) name3860 (
		\u12_o9_we_reg/P0001 ,
		\u8_mem_reg[2][22]/NET0131 ,
		\u8_wp_reg[0]/P0001 ,
		\u8_wp_reg[1]/NET0131 ,
		_w6007_
	);
	LUT4 #(
		.INIT('h0800)
	) name3861 (
		\u12_dout_reg[22]/P0001 ,
		\u12_o9_we_reg/P0001 ,
		\u8_wp_reg[0]/P0001 ,
		\u8_wp_reg[1]/NET0131 ,
		_w6008_
	);
	LUT2 #(
		.INIT('he)
	) name3862 (
		_w6007_,
		_w6008_,
		_w6009_
	);
	LUT4 #(
		.INIT('hc4cc)
	) name3863 (
		\u12_o9_we_reg/P0001 ,
		\u8_mem_reg[2][23]/NET0131 ,
		\u8_wp_reg[0]/P0001 ,
		\u8_wp_reg[1]/NET0131 ,
		_w6010_
	);
	LUT4 #(
		.INIT('h0800)
	) name3864 (
		\u12_dout_reg[23]/P0001 ,
		\u12_o9_we_reg/P0001 ,
		\u8_wp_reg[0]/P0001 ,
		\u8_wp_reg[1]/NET0131 ,
		_w6011_
	);
	LUT2 #(
		.INIT('he)
	) name3865 (
		_w6010_,
		_w6011_,
		_w6012_
	);
	LUT4 #(
		.INIT('hc4cc)
	) name3866 (
		\u12_o9_we_reg/P0001 ,
		\u8_mem_reg[2][24]/NET0131 ,
		\u8_wp_reg[0]/P0001 ,
		\u8_wp_reg[1]/NET0131 ,
		_w6013_
	);
	LUT4 #(
		.INIT('h0800)
	) name3867 (
		\u12_dout_reg[24]/P0001 ,
		\u12_o9_we_reg/P0001 ,
		\u8_wp_reg[0]/P0001 ,
		\u8_wp_reg[1]/NET0131 ,
		_w6014_
	);
	LUT2 #(
		.INIT('he)
	) name3868 (
		_w6013_,
		_w6014_,
		_w6015_
	);
	LUT4 #(
		.INIT('hc4cc)
	) name3869 (
		\u12_o9_we_reg/P0001 ,
		\u8_mem_reg[2][25]/NET0131 ,
		\u8_wp_reg[0]/P0001 ,
		\u8_wp_reg[1]/NET0131 ,
		_w6016_
	);
	LUT4 #(
		.INIT('h0800)
	) name3870 (
		\u12_dout_reg[25]/P0001 ,
		\u12_o9_we_reg/P0001 ,
		\u8_wp_reg[0]/P0001 ,
		\u8_wp_reg[1]/NET0131 ,
		_w6017_
	);
	LUT2 #(
		.INIT('he)
	) name3871 (
		_w6016_,
		_w6017_,
		_w6018_
	);
	LUT4 #(
		.INIT('hcc4c)
	) name3872 (
		\u12_o3_we_reg/P0001 ,
		\u3_mem_reg[1][24]/NET0131 ,
		\u3_wp_reg[0]/P0001 ,
		\u3_wp_reg[1]/NET0131 ,
		_w6019_
	);
	LUT4 #(
		.INIT('h0080)
	) name3873 (
		\u12_dout_reg[24]/P0001 ,
		\u12_o3_we_reg/P0001 ,
		\u3_wp_reg[0]/P0001 ,
		\u3_wp_reg[1]/NET0131 ,
		_w6020_
	);
	LUT2 #(
		.INIT('he)
	) name3874 (
		_w6019_,
		_w6020_,
		_w6021_
	);
	LUT4 #(
		.INIT('hc4cc)
	) name3875 (
		\u12_o9_we_reg/P0001 ,
		\u8_mem_reg[2][26]/NET0131 ,
		\u8_wp_reg[0]/P0001 ,
		\u8_wp_reg[1]/NET0131 ,
		_w6022_
	);
	LUT4 #(
		.INIT('h0800)
	) name3876 (
		\u12_dout_reg[26]/P0001 ,
		\u12_o9_we_reg/P0001 ,
		\u8_wp_reg[0]/P0001 ,
		\u8_wp_reg[1]/NET0131 ,
		_w6023_
	);
	LUT2 #(
		.INIT('he)
	) name3877 (
		_w6022_,
		_w6023_,
		_w6024_
	);
	LUT4 #(
		.INIT('hc4cc)
	) name3878 (
		\u12_o9_we_reg/P0001 ,
		\u8_mem_reg[2][27]/NET0131 ,
		\u8_wp_reg[0]/P0001 ,
		\u8_wp_reg[1]/NET0131 ,
		_w6025_
	);
	LUT4 #(
		.INIT('h0800)
	) name3879 (
		\u12_dout_reg[27]/P0001 ,
		\u12_o9_we_reg/P0001 ,
		\u8_wp_reg[0]/P0001 ,
		\u8_wp_reg[1]/NET0131 ,
		_w6026_
	);
	LUT2 #(
		.INIT('he)
	) name3880 (
		_w6025_,
		_w6026_,
		_w6027_
	);
	LUT4 #(
		.INIT('hcc4c)
	) name3881 (
		\u12_o3_we_reg/P0001 ,
		\u3_mem_reg[1][25]/NET0131 ,
		\u3_wp_reg[0]/P0001 ,
		\u3_wp_reg[1]/NET0131 ,
		_w6028_
	);
	LUT4 #(
		.INIT('h0080)
	) name3882 (
		\u12_dout_reg[25]/P0001 ,
		\u12_o3_we_reg/P0001 ,
		\u3_wp_reg[0]/P0001 ,
		\u3_wp_reg[1]/NET0131 ,
		_w6029_
	);
	LUT2 #(
		.INIT('he)
	) name3883 (
		_w6028_,
		_w6029_,
		_w6030_
	);
	LUT4 #(
		.INIT('hc4cc)
	) name3884 (
		\u12_o9_we_reg/P0001 ,
		\u8_mem_reg[2][28]/NET0131 ,
		\u8_wp_reg[0]/P0001 ,
		\u8_wp_reg[1]/NET0131 ,
		_w6031_
	);
	LUT4 #(
		.INIT('h0800)
	) name3885 (
		\u12_dout_reg[28]/P0001 ,
		\u12_o9_we_reg/P0001 ,
		\u8_wp_reg[0]/P0001 ,
		\u8_wp_reg[1]/NET0131 ,
		_w6032_
	);
	LUT2 #(
		.INIT('he)
	) name3886 (
		_w6031_,
		_w6032_,
		_w6033_
	);
	LUT4 #(
		.INIT('hc4cc)
	) name3887 (
		\u12_o9_we_reg/P0001 ,
		\u8_mem_reg[2][29]/NET0131 ,
		\u8_wp_reg[0]/P0001 ,
		\u8_wp_reg[1]/NET0131 ,
		_w6034_
	);
	LUT4 #(
		.INIT('h0800)
	) name3888 (
		\u12_dout_reg[29]/P0001 ,
		\u12_o9_we_reg/P0001 ,
		\u8_wp_reg[0]/P0001 ,
		\u8_wp_reg[1]/NET0131 ,
		_w6035_
	);
	LUT2 #(
		.INIT('he)
	) name3889 (
		_w6034_,
		_w6035_,
		_w6036_
	);
	LUT4 #(
		.INIT('hcc4c)
	) name3890 (
		\u12_o3_we_reg/P0001 ,
		\u3_mem_reg[1][26]/NET0131 ,
		\u3_wp_reg[0]/P0001 ,
		\u3_wp_reg[1]/NET0131 ,
		_w6037_
	);
	LUT4 #(
		.INIT('h0080)
	) name3891 (
		\u12_dout_reg[26]/P0001 ,
		\u12_o3_we_reg/P0001 ,
		\u3_wp_reg[0]/P0001 ,
		\u3_wp_reg[1]/NET0131 ,
		_w6038_
	);
	LUT2 #(
		.INIT('he)
	) name3892 (
		_w6037_,
		_w6038_,
		_w6039_
	);
	LUT4 #(
		.INIT('hc4cc)
	) name3893 (
		\u12_o9_we_reg/P0001 ,
		\u8_mem_reg[2][2]/NET0131 ,
		\u8_wp_reg[0]/P0001 ,
		\u8_wp_reg[1]/NET0131 ,
		_w6040_
	);
	LUT4 #(
		.INIT('h0800)
	) name3894 (
		\u12_dout_reg[2]/P0001 ,
		\u12_o9_we_reg/P0001 ,
		\u8_wp_reg[0]/P0001 ,
		\u8_wp_reg[1]/NET0131 ,
		_w6041_
	);
	LUT2 #(
		.INIT('he)
	) name3895 (
		_w6040_,
		_w6041_,
		_w6042_
	);
	LUT4 #(
		.INIT('hc4cc)
	) name3896 (
		\u12_o9_we_reg/P0001 ,
		\u8_mem_reg[2][30]/NET0131 ,
		\u8_wp_reg[0]/P0001 ,
		\u8_wp_reg[1]/NET0131 ,
		_w6043_
	);
	LUT4 #(
		.INIT('h0800)
	) name3897 (
		\u12_dout_reg[30]/P0001 ,
		\u12_o9_we_reg/P0001 ,
		\u8_wp_reg[0]/P0001 ,
		\u8_wp_reg[1]/NET0131 ,
		_w6044_
	);
	LUT2 #(
		.INIT('he)
	) name3898 (
		_w6043_,
		_w6044_,
		_w6045_
	);
	LUT4 #(
		.INIT('hc4cc)
	) name3899 (
		\u12_o9_we_reg/P0001 ,
		\u8_mem_reg[2][31]/NET0131 ,
		\u8_wp_reg[0]/P0001 ,
		\u8_wp_reg[1]/NET0131 ,
		_w6046_
	);
	LUT4 #(
		.INIT('h0800)
	) name3900 (
		\u12_dout_reg[31]/P0001 ,
		\u12_o9_we_reg/P0001 ,
		\u8_wp_reg[0]/P0001 ,
		\u8_wp_reg[1]/NET0131 ,
		_w6047_
	);
	LUT2 #(
		.INIT('he)
	) name3901 (
		_w6046_,
		_w6047_,
		_w6048_
	);
	LUT4 #(
		.INIT('hcc4c)
	) name3902 (
		\u12_o3_we_reg/P0001 ,
		\u3_mem_reg[1][28]/NET0131 ,
		\u3_wp_reg[0]/P0001 ,
		\u3_wp_reg[1]/NET0131 ,
		_w6049_
	);
	LUT4 #(
		.INIT('h0080)
	) name3903 (
		\u12_dout_reg[28]/P0001 ,
		\u12_o3_we_reg/P0001 ,
		\u3_wp_reg[0]/P0001 ,
		\u3_wp_reg[1]/NET0131 ,
		_w6050_
	);
	LUT2 #(
		.INIT('he)
	) name3904 (
		_w6049_,
		_w6050_,
		_w6051_
	);
	LUT4 #(
		.INIT('hc4cc)
	) name3905 (
		\u12_o9_we_reg/P0001 ,
		\u8_mem_reg[2][4]/NET0131 ,
		\u8_wp_reg[0]/P0001 ,
		\u8_wp_reg[1]/NET0131 ,
		_w6052_
	);
	LUT4 #(
		.INIT('h0800)
	) name3906 (
		\u12_dout_reg[4]/P0001 ,
		\u12_o9_we_reg/P0001 ,
		\u8_wp_reg[0]/P0001 ,
		\u8_wp_reg[1]/NET0131 ,
		_w6053_
	);
	LUT2 #(
		.INIT('he)
	) name3907 (
		_w6052_,
		_w6053_,
		_w6054_
	);
	LUT3 #(
		.INIT('h02)
	) name3908 (
		\u12_o3_we_reg/P0001 ,
		\u3_wp_reg[0]/P0001 ,
		\u3_wp_reg[1]/NET0131 ,
		_w6055_
	);
	LUT3 #(
		.INIT('h02)
	) name3909 (
		\u12_o4_we_reg/P0001 ,
		\u4_wp_reg[0]/P0001 ,
		\u4_wp_reg[1]/NET0131 ,
		_w6056_
	);
	LUT3 #(
		.INIT('h02)
	) name3910 (
		\u12_o6_we_reg/P0001 ,
		\u5_wp_reg[0]/P0001 ,
		\u5_wp_reg[1]/NET0131 ,
		_w6057_
	);
	LUT3 #(
		.INIT('h02)
	) name3911 (
		\u12_o7_we_reg/P0001 ,
		\u6_wp_reg[0]/P0001 ,
		\u6_wp_reg[1]/NET0131 ,
		_w6058_
	);
	LUT3 #(
		.INIT('h02)
	) name3912 (
		\u12_o8_we_reg/P0001 ,
		\u7_wp_reg[0]/P0001 ,
		\u7_wp_reg[1]/NET0131 ,
		_w6059_
	);
	LUT3 #(
		.INIT('h02)
	) name3913 (
		\u12_o9_we_reg/P0001 ,
		\u8_wp_reg[0]/P0001 ,
		\u8_wp_reg[1]/NET0131 ,
		_w6060_
	);
	LUT4 #(
		.INIT('h2000)
	) name3914 (
		\u13_ints_r_reg[0]/NET0131 ,
		\wb_addr_i[2]_pad ,
		\wb_addr_i[3]_pad ,
		\wb_addr_i[4]_pad ,
		_w6061_
	);
	LUT4 #(
		.INIT('h0008)
	) name3915 (
		\u13_occ0_r_reg[0]/NET0131 ,
		\wb_addr_i[2]_pad ,
		\wb_addr_i[3]_pad ,
		\wb_addr_i[4]_pad ,
		_w6062_
	);
	LUT2 #(
		.INIT('h1)
	) name3916 (
		_w6061_,
		_w6062_,
		_w6063_
	);
	LUT4 #(
		.INIT('h0800)
	) name3917 (
		\u13_intm_r_reg[0]/NET0131 ,
		\wb_addr_i[2]_pad ,
		\wb_addr_i[3]_pad ,
		\wb_addr_i[4]_pad ,
		_w6064_
	);
	LUT4 #(
		.INIT('h0080)
	) name3918 (
		\u13_icc_r_reg[0]/NET0131 ,
		\wb_addr_i[2]_pad ,
		\wb_addr_i[3]_pad ,
		\wb_addr_i[4]_pad ,
		_w6065_
	);
	LUT4 #(
		.INIT('h0020)
	) name3919 (
		\u13_occ1_r_reg[0]/NET0131 ,
		\wb_addr_i[2]_pad ,
		\wb_addr_i[3]_pad ,
		\wb_addr_i[4]_pad ,
		_w6066_
	);
	LUT4 #(
		.INIT('h0200)
	) name3920 (
		\u15_crac_din_reg[0]/NET0131 ,
		\wb_addr_i[2]_pad ,
		\wb_addr_i[3]_pad ,
		\wb_addr_i[4]_pad ,
		_w6067_
	);
	LUT4 #(
		.INIT('h0001)
	) name3921 (
		_w6064_,
		_w6065_,
		_w6066_,
		_w6067_,
		_w6068_
	);
	LUT3 #(
		.INIT('h2a)
	) name3922 (
		_w4169_,
		_w6063_,
		_w6068_,
		_w6069_
	);
	LUT3 #(
		.INIT('h80)
	) name3923 (
		\u11_dout_reg[0]/P0001 ,
		_w4167_,
		_w4168_,
		_w6070_
	);
	LUT4 #(
		.INIT('h53ff)
	) name3924 (
		\u10_dout_reg[0]/P0001 ,
		\u9_dout_reg[0]/P0001 ,
		\wb_addr_i[2]_pad ,
		_w4166_,
		_w6071_
	);
	LUT2 #(
		.INIT('h4)
	) name3925 (
		_w6070_,
		_w6071_,
		_w6072_
	);
	LUT2 #(
		.INIT('hb)
	) name3926 (
		_w6069_,
		_w6072_,
		_w6073_
	);
	LUT4 #(
		.INIT('h2000)
	) name3927 (
		\u13_ints_r_reg[10]/NET0131 ,
		\wb_addr_i[2]_pad ,
		\wb_addr_i[3]_pad ,
		\wb_addr_i[4]_pad ,
		_w6074_
	);
	LUT4 #(
		.INIT('h0008)
	) name3928 (
		\u13_occ0_r_reg[10]/NET0131 ,
		\wb_addr_i[2]_pad ,
		\wb_addr_i[3]_pad ,
		\wb_addr_i[4]_pad ,
		_w6075_
	);
	LUT2 #(
		.INIT('h1)
	) name3929 (
		_w6074_,
		_w6075_,
		_w6076_
	);
	LUT4 #(
		.INIT('h0800)
	) name3930 (
		\u13_intm_r_reg[10]/NET0131 ,
		\wb_addr_i[2]_pad ,
		\wb_addr_i[3]_pad ,
		\wb_addr_i[4]_pad ,
		_w6077_
	);
	LUT4 #(
		.INIT('h0080)
	) name3931 (
		\u13_icc_r_reg[10]/NET0131 ,
		\wb_addr_i[2]_pad ,
		\wb_addr_i[3]_pad ,
		\wb_addr_i[4]_pad ,
		_w6078_
	);
	LUT4 #(
		.INIT('h0020)
	) name3932 (
		\u13_occ1_r_reg[10]/NET0131 ,
		\wb_addr_i[2]_pad ,
		\wb_addr_i[3]_pad ,
		\wb_addr_i[4]_pad ,
		_w6079_
	);
	LUT4 #(
		.INIT('h0200)
	) name3933 (
		\u15_crac_din_reg[10]/NET0131 ,
		\wb_addr_i[2]_pad ,
		\wb_addr_i[3]_pad ,
		\wb_addr_i[4]_pad ,
		_w6080_
	);
	LUT4 #(
		.INIT('h0001)
	) name3934 (
		_w6077_,
		_w6078_,
		_w6079_,
		_w6080_,
		_w6081_
	);
	LUT3 #(
		.INIT('h2a)
	) name3935 (
		_w4169_,
		_w6076_,
		_w6081_,
		_w6082_
	);
	LUT3 #(
		.INIT('h80)
	) name3936 (
		\u11_dout_reg[10]/P0001 ,
		_w4167_,
		_w4168_,
		_w6083_
	);
	LUT4 #(
		.INIT('h53ff)
	) name3937 (
		\u10_dout_reg[10]/P0001 ,
		\u9_dout_reg[10]/P0001 ,
		\wb_addr_i[2]_pad ,
		_w4166_,
		_w6084_
	);
	LUT2 #(
		.INIT('h4)
	) name3938 (
		_w6083_,
		_w6084_,
		_w6085_
	);
	LUT2 #(
		.INIT('hb)
	) name3939 (
		_w6082_,
		_w6085_,
		_w6086_
	);
	LUT4 #(
		.INIT('h2000)
	) name3940 (
		\u13_ints_r_reg[11]/NET0131 ,
		\wb_addr_i[2]_pad ,
		\wb_addr_i[3]_pad ,
		\wb_addr_i[4]_pad ,
		_w6087_
	);
	LUT4 #(
		.INIT('h0008)
	) name3941 (
		\u13_occ0_r_reg[11]/NET0131 ,
		\wb_addr_i[2]_pad ,
		\wb_addr_i[3]_pad ,
		\wb_addr_i[4]_pad ,
		_w6088_
	);
	LUT2 #(
		.INIT('h1)
	) name3942 (
		_w6087_,
		_w6088_,
		_w6089_
	);
	LUT4 #(
		.INIT('h0800)
	) name3943 (
		\u13_intm_r_reg[11]/NET0131 ,
		\wb_addr_i[2]_pad ,
		\wb_addr_i[3]_pad ,
		\wb_addr_i[4]_pad ,
		_w6090_
	);
	LUT4 #(
		.INIT('h0080)
	) name3944 (
		\u13_icc_r_reg[11]/NET0131 ,
		\wb_addr_i[2]_pad ,
		\wb_addr_i[3]_pad ,
		\wb_addr_i[4]_pad ,
		_w6091_
	);
	LUT4 #(
		.INIT('h0020)
	) name3945 (
		\u13_occ1_r_reg[11]/NET0131 ,
		\wb_addr_i[2]_pad ,
		\wb_addr_i[3]_pad ,
		\wb_addr_i[4]_pad ,
		_w6092_
	);
	LUT4 #(
		.INIT('h0200)
	) name3946 (
		\u15_crac_din_reg[11]/NET0131 ,
		\wb_addr_i[2]_pad ,
		\wb_addr_i[3]_pad ,
		\wb_addr_i[4]_pad ,
		_w6093_
	);
	LUT4 #(
		.INIT('h0001)
	) name3947 (
		_w6090_,
		_w6091_,
		_w6092_,
		_w6093_,
		_w6094_
	);
	LUT3 #(
		.INIT('h2a)
	) name3948 (
		_w4169_,
		_w6089_,
		_w6094_,
		_w6095_
	);
	LUT3 #(
		.INIT('h80)
	) name3949 (
		\u11_dout_reg[11]/P0001 ,
		_w4167_,
		_w4168_,
		_w6096_
	);
	LUT4 #(
		.INIT('h53ff)
	) name3950 (
		\u10_dout_reg[11]/P0001 ,
		\u9_dout_reg[11]/P0001 ,
		\wb_addr_i[2]_pad ,
		_w4166_,
		_w6097_
	);
	LUT2 #(
		.INIT('h4)
	) name3951 (
		_w6096_,
		_w6097_,
		_w6098_
	);
	LUT2 #(
		.INIT('hb)
	) name3952 (
		_w6095_,
		_w6098_,
		_w6099_
	);
	LUT4 #(
		.INIT('h2000)
	) name3953 (
		\u13_ints_r_reg[12]/NET0131 ,
		\wb_addr_i[2]_pad ,
		\wb_addr_i[3]_pad ,
		\wb_addr_i[4]_pad ,
		_w6100_
	);
	LUT4 #(
		.INIT('h0008)
	) name3954 (
		\u13_occ0_r_reg[12]/NET0131 ,
		\wb_addr_i[2]_pad ,
		\wb_addr_i[3]_pad ,
		\wb_addr_i[4]_pad ,
		_w6101_
	);
	LUT2 #(
		.INIT('h1)
	) name3955 (
		_w6100_,
		_w6101_,
		_w6102_
	);
	LUT4 #(
		.INIT('h0800)
	) name3956 (
		\u13_intm_r_reg[12]/NET0131 ,
		\wb_addr_i[2]_pad ,
		\wb_addr_i[3]_pad ,
		\wb_addr_i[4]_pad ,
		_w6103_
	);
	LUT4 #(
		.INIT('h0080)
	) name3957 (
		\u13_icc_r_reg[12]/NET0131 ,
		\wb_addr_i[2]_pad ,
		\wb_addr_i[3]_pad ,
		\wb_addr_i[4]_pad ,
		_w6104_
	);
	LUT4 #(
		.INIT('h0020)
	) name3958 (
		\u13_occ1_r_reg[12]/NET0131 ,
		\wb_addr_i[2]_pad ,
		\wb_addr_i[3]_pad ,
		\wb_addr_i[4]_pad ,
		_w6105_
	);
	LUT4 #(
		.INIT('h0200)
	) name3959 (
		\u15_crac_din_reg[12]/NET0131 ,
		\wb_addr_i[2]_pad ,
		\wb_addr_i[3]_pad ,
		\wb_addr_i[4]_pad ,
		_w6106_
	);
	LUT4 #(
		.INIT('h0001)
	) name3960 (
		_w6103_,
		_w6104_,
		_w6105_,
		_w6106_,
		_w6107_
	);
	LUT3 #(
		.INIT('h2a)
	) name3961 (
		_w4169_,
		_w6102_,
		_w6107_,
		_w6108_
	);
	LUT3 #(
		.INIT('h80)
	) name3962 (
		\u11_dout_reg[12]/P0001 ,
		_w4167_,
		_w4168_,
		_w6109_
	);
	LUT4 #(
		.INIT('h53ff)
	) name3963 (
		\u10_dout_reg[12]/P0001 ,
		\u9_dout_reg[12]/P0001 ,
		\wb_addr_i[2]_pad ,
		_w4166_,
		_w6110_
	);
	LUT2 #(
		.INIT('h4)
	) name3964 (
		_w6109_,
		_w6110_,
		_w6111_
	);
	LUT2 #(
		.INIT('hb)
	) name3965 (
		_w6108_,
		_w6111_,
		_w6112_
	);
	LUT4 #(
		.INIT('h2000)
	) name3966 (
		\u13_ints_r_reg[13]/NET0131 ,
		\wb_addr_i[2]_pad ,
		\wb_addr_i[3]_pad ,
		\wb_addr_i[4]_pad ,
		_w6113_
	);
	LUT4 #(
		.INIT('h0008)
	) name3967 (
		\u13_occ0_r_reg[13]/NET0131 ,
		\wb_addr_i[2]_pad ,
		\wb_addr_i[3]_pad ,
		\wb_addr_i[4]_pad ,
		_w6114_
	);
	LUT2 #(
		.INIT('h1)
	) name3968 (
		_w6113_,
		_w6114_,
		_w6115_
	);
	LUT4 #(
		.INIT('h0800)
	) name3969 (
		\u13_intm_r_reg[13]/NET0131 ,
		\wb_addr_i[2]_pad ,
		\wb_addr_i[3]_pad ,
		\wb_addr_i[4]_pad ,
		_w6116_
	);
	LUT4 #(
		.INIT('h0080)
	) name3970 (
		\u13_icc_r_reg[13]/NET0131 ,
		\wb_addr_i[2]_pad ,
		\wb_addr_i[3]_pad ,
		\wb_addr_i[4]_pad ,
		_w6117_
	);
	LUT4 #(
		.INIT('h0020)
	) name3971 (
		\u13_occ1_r_reg[13]/NET0131 ,
		\wb_addr_i[2]_pad ,
		\wb_addr_i[3]_pad ,
		\wb_addr_i[4]_pad ,
		_w6118_
	);
	LUT4 #(
		.INIT('h0200)
	) name3972 (
		\u15_crac_din_reg[13]/NET0131 ,
		\wb_addr_i[2]_pad ,
		\wb_addr_i[3]_pad ,
		\wb_addr_i[4]_pad ,
		_w6119_
	);
	LUT4 #(
		.INIT('h0001)
	) name3973 (
		_w6116_,
		_w6117_,
		_w6118_,
		_w6119_,
		_w6120_
	);
	LUT3 #(
		.INIT('h2a)
	) name3974 (
		_w4169_,
		_w6115_,
		_w6120_,
		_w6121_
	);
	LUT3 #(
		.INIT('h80)
	) name3975 (
		\u11_dout_reg[13]/P0001 ,
		_w4167_,
		_w4168_,
		_w6122_
	);
	LUT4 #(
		.INIT('h53ff)
	) name3976 (
		\u10_dout_reg[13]/P0001 ,
		\u9_dout_reg[13]/P0001 ,
		\wb_addr_i[2]_pad ,
		_w4166_,
		_w6123_
	);
	LUT2 #(
		.INIT('h4)
	) name3977 (
		_w6122_,
		_w6123_,
		_w6124_
	);
	LUT2 #(
		.INIT('hb)
	) name3978 (
		_w6121_,
		_w6124_,
		_w6125_
	);
	LUT4 #(
		.INIT('h2000)
	) name3979 (
		\u13_ints_r_reg[14]/NET0131 ,
		\wb_addr_i[2]_pad ,
		\wb_addr_i[3]_pad ,
		\wb_addr_i[4]_pad ,
		_w6126_
	);
	LUT4 #(
		.INIT('h0008)
	) name3980 (
		\u13_occ0_r_reg[14]/NET0131 ,
		\wb_addr_i[2]_pad ,
		\wb_addr_i[3]_pad ,
		\wb_addr_i[4]_pad ,
		_w6127_
	);
	LUT2 #(
		.INIT('h1)
	) name3981 (
		_w6126_,
		_w6127_,
		_w6128_
	);
	LUT4 #(
		.INIT('h0800)
	) name3982 (
		\u13_intm_r_reg[14]/NET0131 ,
		\wb_addr_i[2]_pad ,
		\wb_addr_i[3]_pad ,
		\wb_addr_i[4]_pad ,
		_w6129_
	);
	LUT4 #(
		.INIT('h0080)
	) name3983 (
		\u13_icc_r_reg[14]/NET0131 ,
		\wb_addr_i[2]_pad ,
		\wb_addr_i[3]_pad ,
		\wb_addr_i[4]_pad ,
		_w6130_
	);
	LUT4 #(
		.INIT('h0020)
	) name3984 (
		\u13_occ1_r_reg[14]/NET0131 ,
		\wb_addr_i[2]_pad ,
		\wb_addr_i[3]_pad ,
		\wb_addr_i[4]_pad ,
		_w6131_
	);
	LUT4 #(
		.INIT('h0200)
	) name3985 (
		\u15_crac_din_reg[14]/NET0131 ,
		\wb_addr_i[2]_pad ,
		\wb_addr_i[3]_pad ,
		\wb_addr_i[4]_pad ,
		_w6132_
	);
	LUT4 #(
		.INIT('h0001)
	) name3986 (
		_w6129_,
		_w6130_,
		_w6131_,
		_w6132_,
		_w6133_
	);
	LUT3 #(
		.INIT('h2a)
	) name3987 (
		_w4169_,
		_w6128_,
		_w6133_,
		_w6134_
	);
	LUT3 #(
		.INIT('h80)
	) name3988 (
		\u11_dout_reg[14]/P0001 ,
		_w4167_,
		_w4168_,
		_w6135_
	);
	LUT4 #(
		.INIT('h53ff)
	) name3989 (
		\u10_dout_reg[14]/P0001 ,
		\u9_dout_reg[14]/P0001 ,
		\wb_addr_i[2]_pad ,
		_w4166_,
		_w6136_
	);
	LUT2 #(
		.INIT('h4)
	) name3990 (
		_w6135_,
		_w6136_,
		_w6137_
	);
	LUT2 #(
		.INIT('hb)
	) name3991 (
		_w6134_,
		_w6137_,
		_w6138_
	);
	LUT4 #(
		.INIT('h0800)
	) name3992 (
		\u13_intm_r_reg[15]/NET0131 ,
		\wb_addr_i[2]_pad ,
		\wb_addr_i[3]_pad ,
		\wb_addr_i[4]_pad ,
		_w6139_
	);
	LUT4 #(
		.INIT('h0020)
	) name3993 (
		\u13_occ1_r_reg[15]/NET0131 ,
		\wb_addr_i[2]_pad ,
		\wb_addr_i[3]_pad ,
		\wb_addr_i[4]_pad ,
		_w6140_
	);
	LUT2 #(
		.INIT('h1)
	) name3994 (
		_w6139_,
		_w6140_,
		_w6141_
	);
	LUT4 #(
		.INIT('h0008)
	) name3995 (
		\u13_occ0_r_reg[15]/NET0131 ,
		\wb_addr_i[2]_pad ,
		\wb_addr_i[3]_pad ,
		\wb_addr_i[4]_pad ,
		_w6142_
	);
	LUT4 #(
		.INIT('h0080)
	) name3996 (
		\u13_icc_r_reg[15]/NET0131 ,
		\wb_addr_i[2]_pad ,
		\wb_addr_i[3]_pad ,
		\wb_addr_i[4]_pad ,
		_w6143_
	);
	LUT4 #(
		.INIT('h2000)
	) name3997 (
		\u13_ints_r_reg[15]/NET0131 ,
		\wb_addr_i[2]_pad ,
		\wb_addr_i[3]_pad ,
		\wb_addr_i[4]_pad ,
		_w6144_
	);
	LUT4 #(
		.INIT('h0200)
	) name3998 (
		\u15_crac_din_reg[15]/NET0131 ,
		\wb_addr_i[2]_pad ,
		\wb_addr_i[3]_pad ,
		\wb_addr_i[4]_pad ,
		_w6145_
	);
	LUT4 #(
		.INIT('h0001)
	) name3999 (
		_w6142_,
		_w6143_,
		_w6144_,
		_w6145_,
		_w6146_
	);
	LUT3 #(
		.INIT('h2a)
	) name4000 (
		_w4169_,
		_w6141_,
		_w6146_,
		_w6147_
	);
	LUT3 #(
		.INIT('h80)
	) name4001 (
		\u11_dout_reg[15]/P0001 ,
		_w4167_,
		_w4168_,
		_w6148_
	);
	LUT4 #(
		.INIT('h53ff)
	) name4002 (
		\u10_dout_reg[15]/P0001 ,
		\u9_dout_reg[15]/P0001 ,
		\wb_addr_i[2]_pad ,
		_w4166_,
		_w6149_
	);
	LUT2 #(
		.INIT('h4)
	) name4003 (
		_w6148_,
		_w6149_,
		_w6150_
	);
	LUT2 #(
		.INIT('hb)
	) name4004 (
		_w6147_,
		_w6150_,
		_w6151_
	);
	LUT4 #(
		.INIT('h2000)
	) name4005 (
		\u13_ints_r_reg[2]/NET0131 ,
		\wb_addr_i[2]_pad ,
		\wb_addr_i[3]_pad ,
		\wb_addr_i[4]_pad ,
		_w6152_
	);
	LUT4 #(
		.INIT('h0008)
	) name4006 (
		\u13_occ0_r_reg[2]/NET0131 ,
		\wb_addr_i[2]_pad ,
		\wb_addr_i[3]_pad ,
		\wb_addr_i[4]_pad ,
		_w6153_
	);
	LUT2 #(
		.INIT('h1)
	) name4007 (
		_w6152_,
		_w6153_,
		_w6154_
	);
	LUT4 #(
		.INIT('h0800)
	) name4008 (
		\u13_intm_r_reg[2]/NET0131 ,
		\wb_addr_i[2]_pad ,
		\wb_addr_i[3]_pad ,
		\wb_addr_i[4]_pad ,
		_w6155_
	);
	LUT4 #(
		.INIT('h0080)
	) name4009 (
		\u13_icc_r_reg[2]/NET0131 ,
		\wb_addr_i[2]_pad ,
		\wb_addr_i[3]_pad ,
		\wb_addr_i[4]_pad ,
		_w6156_
	);
	LUT4 #(
		.INIT('h0020)
	) name4010 (
		\u13_occ1_r_reg[2]/NET0131 ,
		\wb_addr_i[2]_pad ,
		\wb_addr_i[3]_pad ,
		\wb_addr_i[4]_pad ,
		_w6157_
	);
	LUT4 #(
		.INIT('h0200)
	) name4011 (
		\u15_crac_din_reg[2]/NET0131 ,
		\wb_addr_i[2]_pad ,
		\wb_addr_i[3]_pad ,
		\wb_addr_i[4]_pad ,
		_w6158_
	);
	LUT4 #(
		.INIT('h0001)
	) name4012 (
		_w6155_,
		_w6156_,
		_w6157_,
		_w6158_,
		_w6159_
	);
	LUT3 #(
		.INIT('h2a)
	) name4013 (
		_w4169_,
		_w6154_,
		_w6159_,
		_w6160_
	);
	LUT3 #(
		.INIT('h80)
	) name4014 (
		\u11_dout_reg[2]/P0001 ,
		_w4167_,
		_w4168_,
		_w6161_
	);
	LUT4 #(
		.INIT('h53ff)
	) name4015 (
		\u10_dout_reg[2]/P0001 ,
		\u9_dout_reg[2]/P0001 ,
		\wb_addr_i[2]_pad ,
		_w4166_,
		_w6162_
	);
	LUT2 #(
		.INIT('h4)
	) name4016 (
		_w6161_,
		_w6162_,
		_w6163_
	);
	LUT2 #(
		.INIT('hb)
	) name4017 (
		_w6160_,
		_w6163_,
		_w6164_
	);
	LUT4 #(
		.INIT('h2000)
	) name4018 (
		\u13_ints_r_reg[3]/NET0131 ,
		\wb_addr_i[2]_pad ,
		\wb_addr_i[3]_pad ,
		\wb_addr_i[4]_pad ,
		_w6165_
	);
	LUT4 #(
		.INIT('h0008)
	) name4019 (
		\u13_occ0_r_reg[3]/NET0131 ,
		\wb_addr_i[2]_pad ,
		\wb_addr_i[3]_pad ,
		\wb_addr_i[4]_pad ,
		_w6166_
	);
	LUT2 #(
		.INIT('h1)
	) name4020 (
		_w6165_,
		_w6166_,
		_w6167_
	);
	LUT4 #(
		.INIT('h0800)
	) name4021 (
		\u13_intm_r_reg[3]/NET0131 ,
		\wb_addr_i[2]_pad ,
		\wb_addr_i[3]_pad ,
		\wb_addr_i[4]_pad ,
		_w6168_
	);
	LUT4 #(
		.INIT('h0080)
	) name4022 (
		\u13_icc_r_reg[3]/NET0131 ,
		\wb_addr_i[2]_pad ,
		\wb_addr_i[3]_pad ,
		\wb_addr_i[4]_pad ,
		_w6169_
	);
	LUT4 #(
		.INIT('h0020)
	) name4023 (
		\u13_occ1_r_reg[3]/NET0131 ,
		\wb_addr_i[2]_pad ,
		\wb_addr_i[3]_pad ,
		\wb_addr_i[4]_pad ,
		_w6170_
	);
	LUT4 #(
		.INIT('h0200)
	) name4024 (
		\u15_crac_din_reg[3]/NET0131 ,
		\wb_addr_i[2]_pad ,
		\wb_addr_i[3]_pad ,
		\wb_addr_i[4]_pad ,
		_w6171_
	);
	LUT4 #(
		.INIT('h0001)
	) name4025 (
		_w6168_,
		_w6169_,
		_w6170_,
		_w6171_,
		_w6172_
	);
	LUT3 #(
		.INIT('h2a)
	) name4026 (
		_w4169_,
		_w6167_,
		_w6172_,
		_w6173_
	);
	LUT3 #(
		.INIT('h80)
	) name4027 (
		\u11_dout_reg[3]/P0001 ,
		_w4167_,
		_w4168_,
		_w6174_
	);
	LUT4 #(
		.INIT('h53ff)
	) name4028 (
		\u10_dout_reg[3]/P0001 ,
		\u9_dout_reg[3]/P0001 ,
		\wb_addr_i[2]_pad ,
		_w4166_,
		_w6175_
	);
	LUT2 #(
		.INIT('h4)
	) name4029 (
		_w6174_,
		_w6175_,
		_w6176_
	);
	LUT2 #(
		.INIT('hb)
	) name4030 (
		_w6173_,
		_w6176_,
		_w6177_
	);
	LUT4 #(
		.INIT('h2000)
	) name4031 (
		\u13_ints_r_reg[4]/NET0131 ,
		\wb_addr_i[2]_pad ,
		\wb_addr_i[3]_pad ,
		\wb_addr_i[4]_pad ,
		_w6178_
	);
	LUT4 #(
		.INIT('h0008)
	) name4032 (
		\u13_occ0_r_reg[4]/NET0131 ,
		\wb_addr_i[2]_pad ,
		\wb_addr_i[3]_pad ,
		\wb_addr_i[4]_pad ,
		_w6179_
	);
	LUT2 #(
		.INIT('h1)
	) name4033 (
		_w6178_,
		_w6179_,
		_w6180_
	);
	LUT4 #(
		.INIT('h0800)
	) name4034 (
		\u13_intm_r_reg[4]/NET0131 ,
		\wb_addr_i[2]_pad ,
		\wb_addr_i[3]_pad ,
		\wb_addr_i[4]_pad ,
		_w6181_
	);
	LUT4 #(
		.INIT('h0080)
	) name4035 (
		\u13_icc_r_reg[4]/NET0131 ,
		\wb_addr_i[2]_pad ,
		\wb_addr_i[3]_pad ,
		\wb_addr_i[4]_pad ,
		_w6182_
	);
	LUT4 #(
		.INIT('h0020)
	) name4036 (
		\u13_occ1_r_reg[4]/NET0131 ,
		\wb_addr_i[2]_pad ,
		\wb_addr_i[3]_pad ,
		\wb_addr_i[4]_pad ,
		_w6183_
	);
	LUT4 #(
		.INIT('h0200)
	) name4037 (
		\u15_crac_din_reg[4]/NET0131 ,
		\wb_addr_i[2]_pad ,
		\wb_addr_i[3]_pad ,
		\wb_addr_i[4]_pad ,
		_w6184_
	);
	LUT4 #(
		.INIT('h0001)
	) name4038 (
		_w6181_,
		_w6182_,
		_w6183_,
		_w6184_,
		_w6185_
	);
	LUT3 #(
		.INIT('h2a)
	) name4039 (
		_w4169_,
		_w6180_,
		_w6185_,
		_w6186_
	);
	LUT3 #(
		.INIT('h80)
	) name4040 (
		\u11_dout_reg[4]/P0001 ,
		_w4167_,
		_w4168_,
		_w6187_
	);
	LUT4 #(
		.INIT('h53ff)
	) name4041 (
		\u10_dout_reg[4]/P0001 ,
		\u9_dout_reg[4]/P0001 ,
		\wb_addr_i[2]_pad ,
		_w4166_,
		_w6188_
	);
	LUT2 #(
		.INIT('h4)
	) name4042 (
		_w6187_,
		_w6188_,
		_w6189_
	);
	LUT2 #(
		.INIT('hb)
	) name4043 (
		_w6186_,
		_w6189_,
		_w6190_
	);
	LUT4 #(
		.INIT('h2000)
	) name4044 (
		\u13_ints_r_reg[5]/NET0131 ,
		\wb_addr_i[2]_pad ,
		\wb_addr_i[3]_pad ,
		\wb_addr_i[4]_pad ,
		_w6191_
	);
	LUT4 #(
		.INIT('h0008)
	) name4045 (
		\u13_occ0_r_reg[5]/NET0131 ,
		\wb_addr_i[2]_pad ,
		\wb_addr_i[3]_pad ,
		\wb_addr_i[4]_pad ,
		_w6192_
	);
	LUT2 #(
		.INIT('h1)
	) name4046 (
		_w6191_,
		_w6192_,
		_w6193_
	);
	LUT4 #(
		.INIT('h0800)
	) name4047 (
		\u13_intm_r_reg[5]/NET0131 ,
		\wb_addr_i[2]_pad ,
		\wb_addr_i[3]_pad ,
		\wb_addr_i[4]_pad ,
		_w6194_
	);
	LUT4 #(
		.INIT('h0080)
	) name4048 (
		\u13_icc_r_reg[5]/NET0131 ,
		\wb_addr_i[2]_pad ,
		\wb_addr_i[3]_pad ,
		\wb_addr_i[4]_pad ,
		_w6195_
	);
	LUT4 #(
		.INIT('h0020)
	) name4049 (
		\u13_occ1_r_reg[5]/NET0131 ,
		\wb_addr_i[2]_pad ,
		\wb_addr_i[3]_pad ,
		\wb_addr_i[4]_pad ,
		_w6196_
	);
	LUT4 #(
		.INIT('h0200)
	) name4050 (
		\u15_crac_din_reg[5]/NET0131 ,
		\wb_addr_i[2]_pad ,
		\wb_addr_i[3]_pad ,
		\wb_addr_i[4]_pad ,
		_w6197_
	);
	LUT4 #(
		.INIT('h0001)
	) name4051 (
		_w6194_,
		_w6195_,
		_w6196_,
		_w6197_,
		_w6198_
	);
	LUT3 #(
		.INIT('h2a)
	) name4052 (
		_w4169_,
		_w6193_,
		_w6198_,
		_w6199_
	);
	LUT3 #(
		.INIT('h80)
	) name4053 (
		\u11_dout_reg[5]/P0001 ,
		_w4167_,
		_w4168_,
		_w6200_
	);
	LUT4 #(
		.INIT('h53ff)
	) name4054 (
		\u10_dout_reg[5]/P0001 ,
		\u9_dout_reg[5]/P0001 ,
		\wb_addr_i[2]_pad ,
		_w4166_,
		_w6201_
	);
	LUT2 #(
		.INIT('h4)
	) name4055 (
		_w6200_,
		_w6201_,
		_w6202_
	);
	LUT2 #(
		.INIT('hb)
	) name4056 (
		_w6199_,
		_w6202_,
		_w6203_
	);
	LUT4 #(
		.INIT('h2000)
	) name4057 (
		\u13_ints_r_reg[6]/NET0131 ,
		\wb_addr_i[2]_pad ,
		\wb_addr_i[3]_pad ,
		\wb_addr_i[4]_pad ,
		_w6204_
	);
	LUT4 #(
		.INIT('h0008)
	) name4058 (
		\u13_occ0_r_reg[6]/NET0131 ,
		\wb_addr_i[2]_pad ,
		\wb_addr_i[3]_pad ,
		\wb_addr_i[4]_pad ,
		_w6205_
	);
	LUT2 #(
		.INIT('h1)
	) name4059 (
		_w6204_,
		_w6205_,
		_w6206_
	);
	LUT4 #(
		.INIT('h0800)
	) name4060 (
		\u13_intm_r_reg[6]/NET0131 ,
		\wb_addr_i[2]_pad ,
		\wb_addr_i[3]_pad ,
		\wb_addr_i[4]_pad ,
		_w6207_
	);
	LUT4 #(
		.INIT('h0080)
	) name4061 (
		\u13_icc_r_reg[6]/NET0131 ,
		\wb_addr_i[2]_pad ,
		\wb_addr_i[3]_pad ,
		\wb_addr_i[4]_pad ,
		_w6208_
	);
	LUT4 #(
		.INIT('h0020)
	) name4062 (
		\u13_occ1_r_reg[6]/NET0131 ,
		\wb_addr_i[2]_pad ,
		\wb_addr_i[3]_pad ,
		\wb_addr_i[4]_pad ,
		_w6209_
	);
	LUT4 #(
		.INIT('h0200)
	) name4063 (
		\u15_crac_din_reg[6]/NET0131 ,
		\wb_addr_i[2]_pad ,
		\wb_addr_i[3]_pad ,
		\wb_addr_i[4]_pad ,
		_w6210_
	);
	LUT4 #(
		.INIT('h0001)
	) name4064 (
		_w6207_,
		_w6208_,
		_w6209_,
		_w6210_,
		_w6211_
	);
	LUT3 #(
		.INIT('h2a)
	) name4065 (
		_w4169_,
		_w6206_,
		_w6211_,
		_w6212_
	);
	LUT3 #(
		.INIT('h80)
	) name4066 (
		\u11_dout_reg[6]/P0001 ,
		_w4167_,
		_w4168_,
		_w6213_
	);
	LUT4 #(
		.INIT('h53ff)
	) name4067 (
		\u10_dout_reg[6]/P0001 ,
		\u9_dout_reg[6]/P0001 ,
		\wb_addr_i[2]_pad ,
		_w4166_,
		_w6214_
	);
	LUT2 #(
		.INIT('h4)
	) name4068 (
		_w6213_,
		_w6214_,
		_w6215_
	);
	LUT2 #(
		.INIT('hb)
	) name4069 (
		_w6212_,
		_w6215_,
		_w6216_
	);
	LUT4 #(
		.INIT('h0800)
	) name4070 (
		\u13_intm_r_reg[7]/NET0131 ,
		\wb_addr_i[2]_pad ,
		\wb_addr_i[3]_pad ,
		\wb_addr_i[4]_pad ,
		_w6217_
	);
	LUT4 #(
		.INIT('h0020)
	) name4071 (
		\u13_occ1_r_reg[7]/NET0131 ,
		\wb_addr_i[2]_pad ,
		\wb_addr_i[3]_pad ,
		\wb_addr_i[4]_pad ,
		_w6218_
	);
	LUT2 #(
		.INIT('h1)
	) name4072 (
		_w6217_,
		_w6218_,
		_w6219_
	);
	LUT4 #(
		.INIT('h0008)
	) name4073 (
		\u13_occ0_r_reg[7]/NET0131 ,
		\wb_addr_i[2]_pad ,
		\wb_addr_i[3]_pad ,
		\wb_addr_i[4]_pad ,
		_w6220_
	);
	LUT4 #(
		.INIT('h0080)
	) name4074 (
		\u13_icc_r_reg[7]/NET0131 ,
		\wb_addr_i[2]_pad ,
		\wb_addr_i[3]_pad ,
		\wb_addr_i[4]_pad ,
		_w6221_
	);
	LUT4 #(
		.INIT('h2000)
	) name4075 (
		\u13_ints_r_reg[7]/NET0131 ,
		\wb_addr_i[2]_pad ,
		\wb_addr_i[3]_pad ,
		\wb_addr_i[4]_pad ,
		_w6222_
	);
	LUT4 #(
		.INIT('h0200)
	) name4076 (
		\u15_crac_din_reg[7]/NET0131 ,
		\wb_addr_i[2]_pad ,
		\wb_addr_i[3]_pad ,
		\wb_addr_i[4]_pad ,
		_w6223_
	);
	LUT4 #(
		.INIT('h0001)
	) name4077 (
		_w6220_,
		_w6221_,
		_w6222_,
		_w6223_,
		_w6224_
	);
	LUT3 #(
		.INIT('h2a)
	) name4078 (
		_w4169_,
		_w6219_,
		_w6224_,
		_w6225_
	);
	LUT3 #(
		.INIT('h80)
	) name4079 (
		\u11_dout_reg[7]/P0001 ,
		_w4167_,
		_w4168_,
		_w6226_
	);
	LUT4 #(
		.INIT('h53ff)
	) name4080 (
		\u10_dout_reg[7]/P0001 ,
		\u9_dout_reg[7]/P0001 ,
		\wb_addr_i[2]_pad ,
		_w4166_,
		_w6227_
	);
	LUT2 #(
		.INIT('h4)
	) name4081 (
		_w6226_,
		_w6227_,
		_w6228_
	);
	LUT2 #(
		.INIT('hb)
	) name4082 (
		_w6225_,
		_w6228_,
		_w6229_
	);
	LUT4 #(
		.INIT('h2000)
	) name4083 (
		\u13_ints_r_reg[8]/NET0131 ,
		\wb_addr_i[2]_pad ,
		\wb_addr_i[3]_pad ,
		\wb_addr_i[4]_pad ,
		_w6230_
	);
	LUT4 #(
		.INIT('h0008)
	) name4084 (
		\u13_occ0_r_reg[8]/NET0131 ,
		\wb_addr_i[2]_pad ,
		\wb_addr_i[3]_pad ,
		\wb_addr_i[4]_pad ,
		_w6231_
	);
	LUT2 #(
		.INIT('h1)
	) name4085 (
		_w6230_,
		_w6231_,
		_w6232_
	);
	LUT4 #(
		.INIT('h0800)
	) name4086 (
		\u13_intm_r_reg[8]/NET0131 ,
		\wb_addr_i[2]_pad ,
		\wb_addr_i[3]_pad ,
		\wb_addr_i[4]_pad ,
		_w6233_
	);
	LUT4 #(
		.INIT('h0080)
	) name4087 (
		\u13_icc_r_reg[8]/NET0131 ,
		\wb_addr_i[2]_pad ,
		\wb_addr_i[3]_pad ,
		\wb_addr_i[4]_pad ,
		_w6234_
	);
	LUT4 #(
		.INIT('h0020)
	) name4088 (
		\u13_occ1_r_reg[8]/NET0131 ,
		\wb_addr_i[2]_pad ,
		\wb_addr_i[3]_pad ,
		\wb_addr_i[4]_pad ,
		_w6235_
	);
	LUT4 #(
		.INIT('h0200)
	) name4089 (
		\u15_crac_din_reg[8]/NET0131 ,
		\wb_addr_i[2]_pad ,
		\wb_addr_i[3]_pad ,
		\wb_addr_i[4]_pad ,
		_w6236_
	);
	LUT4 #(
		.INIT('h0001)
	) name4090 (
		_w6233_,
		_w6234_,
		_w6235_,
		_w6236_,
		_w6237_
	);
	LUT3 #(
		.INIT('h2a)
	) name4091 (
		_w4169_,
		_w6232_,
		_w6237_,
		_w6238_
	);
	LUT3 #(
		.INIT('h80)
	) name4092 (
		\u11_dout_reg[8]/P0001 ,
		_w4167_,
		_w4168_,
		_w6239_
	);
	LUT4 #(
		.INIT('h53ff)
	) name4093 (
		\u10_dout_reg[8]/P0001 ,
		\u9_dout_reg[8]/P0001 ,
		\wb_addr_i[2]_pad ,
		_w4166_,
		_w6240_
	);
	LUT2 #(
		.INIT('h4)
	) name4094 (
		_w6239_,
		_w6240_,
		_w6241_
	);
	LUT2 #(
		.INIT('hb)
	) name4095 (
		_w6238_,
		_w6241_,
		_w6242_
	);
	LUT4 #(
		.INIT('h2000)
	) name4096 (
		\u13_ints_r_reg[9]/NET0131 ,
		\wb_addr_i[2]_pad ,
		\wb_addr_i[3]_pad ,
		\wb_addr_i[4]_pad ,
		_w6243_
	);
	LUT4 #(
		.INIT('h0008)
	) name4097 (
		\u13_occ0_r_reg[9]/NET0131 ,
		\wb_addr_i[2]_pad ,
		\wb_addr_i[3]_pad ,
		\wb_addr_i[4]_pad ,
		_w6244_
	);
	LUT2 #(
		.INIT('h1)
	) name4098 (
		_w6243_,
		_w6244_,
		_w6245_
	);
	LUT4 #(
		.INIT('h0800)
	) name4099 (
		\u13_intm_r_reg[9]/NET0131 ,
		\wb_addr_i[2]_pad ,
		\wb_addr_i[3]_pad ,
		\wb_addr_i[4]_pad ,
		_w6246_
	);
	LUT4 #(
		.INIT('h0080)
	) name4100 (
		\u13_icc_r_reg[9]/NET0131 ,
		\wb_addr_i[2]_pad ,
		\wb_addr_i[3]_pad ,
		\wb_addr_i[4]_pad ,
		_w6247_
	);
	LUT4 #(
		.INIT('h0020)
	) name4101 (
		\u13_occ1_r_reg[9]/NET0131 ,
		\wb_addr_i[2]_pad ,
		\wb_addr_i[3]_pad ,
		\wb_addr_i[4]_pad ,
		_w6248_
	);
	LUT4 #(
		.INIT('h0200)
	) name4102 (
		\u15_crac_din_reg[9]/NET0131 ,
		\wb_addr_i[2]_pad ,
		\wb_addr_i[3]_pad ,
		\wb_addr_i[4]_pad ,
		_w6249_
	);
	LUT4 #(
		.INIT('h0001)
	) name4103 (
		_w6246_,
		_w6247_,
		_w6248_,
		_w6249_,
		_w6250_
	);
	LUT3 #(
		.INIT('h2a)
	) name4104 (
		_w4169_,
		_w6245_,
		_w6250_,
		_w6251_
	);
	LUT3 #(
		.INIT('h80)
	) name4105 (
		\u11_dout_reg[9]/P0001 ,
		_w4167_,
		_w4168_,
		_w6252_
	);
	LUT4 #(
		.INIT('h53ff)
	) name4106 (
		\u10_dout_reg[9]/P0001 ,
		\u9_dout_reg[9]/P0001 ,
		\wb_addr_i[2]_pad ,
		_w4166_,
		_w6253_
	);
	LUT2 #(
		.INIT('h4)
	) name4107 (
		_w6252_,
		_w6253_,
		_w6254_
	);
	LUT2 #(
		.INIT('hb)
	) name4108 (
		_w6251_,
		_w6254_,
		_w6255_
	);
	LUT4 #(
		.INIT('h0200)
	) name4109 (
		\u12_rf_we_reg/P0001 ,
		\wb_addr_i[2]_pad ,
		\wb_addr_i[3]_pad ,
		\wb_addr_i[4]_pad ,
		_w6256_
	);
	LUT4 #(
		.INIT('h0080)
	) name4110 (
		\u12_rf_we_reg/P0001 ,
		\wb_addr_i[2]_pad ,
		\wb_addr_i[3]_pad ,
		\wb_addr_i[4]_pad ,
		_w6257_
	);
	LUT4 #(
		.INIT('h0800)
	) name4111 (
		\u12_rf_we_reg/P0001 ,
		\wb_addr_i[2]_pad ,
		\wb_addr_i[3]_pad ,
		\wb_addr_i[4]_pad ,
		_w6258_
	);
	LUT4 #(
		.INIT('h0008)
	) name4112 (
		\u12_rf_we_reg/P0001 ,
		\wb_addr_i[2]_pad ,
		\wb_addr_i[3]_pad ,
		\wb_addr_i[4]_pad ,
		_w6259_
	);
	LUT4 #(
		.INIT('h0020)
	) name4113 (
		\u12_rf_we_reg/P0001 ,
		\wb_addr_i[2]_pad ,
		\wb_addr_i[3]_pad ,
		\wb_addr_i[4]_pad ,
		_w6260_
	);
	LUT3 #(
		.INIT('hbe)
	) name4114 (
		suspended_o_pad,
		\u2_cnt_reg[4]/NET0131 ,
		_w4320_,
		_w6261_
	);
	LUT4 #(
		.INIT('h8008)
	) name4115 (
		\u4_rp_reg[1]/NET0131 ,
		\u4_rp_reg[2]/NET0131 ,
		\u4_rp_reg[3]/NET0131 ,
		\u4_wp_reg[2]/P0001 ,
		_w6262_
	);
	LUT4 #(
		.INIT('haaa8)
	) name4116 (
		\u4_rp_reg[0]/P0001 ,
		_w2418_,
		_w4228_,
		_w6262_,
		_w6263_
	);
	LUT4 #(
		.INIT('h31c4)
	) name4117 (
		\u4_rp_reg[1]/NET0131 ,
		\u4_rp_reg[2]/NET0131 ,
		\u4_wp_reg[0]/P0001 ,
		\u4_wp_reg[1]/NET0131 ,
		_w6264_
	);
	LUT2 #(
		.INIT('h9)
	) name4118 (
		\u4_rp_reg[1]/NET0131 ,
		\u4_wp_reg[0]/P0001 ,
		_w6265_
	);
	LUT3 #(
		.INIT('h14)
	) name4119 (
		\u4_rp_reg[0]/P0001 ,
		\u4_rp_reg[1]/NET0131 ,
		\u4_wp_reg[0]/P0001 ,
		_w6266_
	);
	LUT3 #(
		.INIT('h80)
	) name4120 (
		\u4_rp_reg[0]/P0001 ,
		\u4_rp_reg[1]/NET0131 ,
		\u4_rp_reg[2]/NET0131 ,
		_w6267_
	);
	LUT4 #(
		.INIT('h0031)
	) name4121 (
		_w4229_,
		_w6266_,
		_w6267_,
		_w6264_,
		_w6268_
	);
	LUT2 #(
		.INIT('h4)
	) name4122 (
		_w6263_,
		_w6268_,
		_w6269_
	);
	LUT4 #(
		.INIT('h8008)
	) name4123 (
		\u5_rp_reg[1]/NET0131 ,
		\u5_rp_reg[2]/NET0131 ,
		\u5_rp_reg[3]/NET0131 ,
		\u5_wp_reg[2]/P0001 ,
		_w6270_
	);
	LUT4 #(
		.INIT('haaa8)
	) name4124 (
		\u5_rp_reg[0]/P0001 ,
		_w2427_,
		_w4232_,
		_w6270_,
		_w6271_
	);
	LUT4 #(
		.INIT('h31c4)
	) name4125 (
		\u5_rp_reg[1]/NET0131 ,
		\u5_rp_reg[2]/NET0131 ,
		\u5_wp_reg[0]/P0001 ,
		\u5_wp_reg[1]/NET0131 ,
		_w6272_
	);
	LUT2 #(
		.INIT('h9)
	) name4126 (
		\u5_rp_reg[1]/NET0131 ,
		\u5_wp_reg[0]/P0001 ,
		_w6273_
	);
	LUT3 #(
		.INIT('h14)
	) name4127 (
		\u5_rp_reg[0]/P0001 ,
		\u5_rp_reg[1]/NET0131 ,
		\u5_wp_reg[0]/P0001 ,
		_w6274_
	);
	LUT3 #(
		.INIT('h80)
	) name4128 (
		\u5_rp_reg[0]/P0001 ,
		\u5_rp_reg[1]/NET0131 ,
		\u5_rp_reg[2]/NET0131 ,
		_w6275_
	);
	LUT4 #(
		.INIT('h0031)
	) name4129 (
		_w4233_,
		_w6274_,
		_w6275_,
		_w6272_,
		_w6276_
	);
	LUT2 #(
		.INIT('h4)
	) name4130 (
		_w6271_,
		_w6276_,
		_w6277_
	);
	LUT3 #(
		.INIT('hca)
	) name4131 (
		\u14_crac_wr_r_reg/P0001 ,
		\u15_crac_wr_reg/NET0131 ,
		\valid_s_reg/NET0131 ,
		_w6278_
	);
	LUT4 #(
		.INIT('hbde7)
	) name4132 (
		\u6_rp_reg[1]/NET0131 ,
		\u6_rp_reg[2]/NET0131 ,
		\u6_wp_reg[0]/P0001 ,
		\u6_wp_reg[1]/NET0131 ,
		_w6279_
	);
	LUT3 #(
		.INIT('ha8)
	) name4133 (
		\u6_rp_reg[0]/P0001 ,
		_w2445_,
		_w6279_,
		_w6280_
	);
	LUT4 #(
		.INIT('h8872)
	) name4134 (
		\u6_rp_reg[0]/P0001 ,
		_w2448_,
		_w4237_,
		_w4238_,
		_w6281_
	);
	LUT2 #(
		.INIT('h4)
	) name4135 (
		_w6280_,
		_w6281_,
		_w6282_
	);
	LUT2 #(
		.INIT('h9)
	) name4136 (
		\u7_rp_reg[1]/NET0131 ,
		\u7_wp_reg[0]/P0001 ,
		_w6283_
	);
	LUT4 #(
		.INIT('h2aa2)
	) name4137 (
		\u7_rp_reg[0]/P0001 ,
		\u7_rp_reg[1]/NET0131 ,
		\u7_rp_reg[2]/NET0131 ,
		\u7_wp_reg[1]/NET0131 ,
		_w6284_
	);
	LUT2 #(
		.INIT('h1)
	) name4138 (
		_w6283_,
		_w6284_,
		_w6285_
	);
	LUT4 #(
		.INIT('h0ee0)
	) name4139 (
		\u13_occ1_r_reg[2]/NET0131 ,
		\u13_occ1_r_reg[3]/NET0131 ,
		\u7_rp_reg[1]/NET0131 ,
		\u7_wp_reg[0]/P0001 ,
		_w6286_
	);
	LUT2 #(
		.INIT('h2)
	) name4140 (
		\u7_rp_reg[0]/P0001 ,
		_w6286_,
		_w6287_
	);
	LUT3 #(
		.INIT('h80)
	) name4141 (
		\u7_rp_reg[0]/P0001 ,
		\u7_rp_reg[1]/NET0131 ,
		\u7_rp_reg[2]/NET0131 ,
		_w6288_
	);
	LUT4 #(
		.INIT('h0770)
	) name4142 (
		\u7_rp_reg[0]/P0001 ,
		\u7_rp_reg[1]/NET0131 ,
		\u7_rp_reg[2]/NET0131 ,
		\u7_wp_reg[1]/NET0131 ,
		_w6289_
	);
	LUT3 #(
		.INIT('h09)
	) name4143 (
		_w4242_,
		_w6288_,
		_w6289_,
		_w6290_
	);
	LUT3 #(
		.INIT('h10)
	) name4144 (
		_w6285_,
		_w6287_,
		_w6290_,
		_w6291_
	);
	LUT2 #(
		.INIT('h9)
	) name4145 (
		\u3_rp_reg[1]/NET0131 ,
		\u3_wp_reg[0]/P0001 ,
		_w6292_
	);
	LUT4 #(
		.INIT('h2aa2)
	) name4146 (
		\u3_rp_reg[0]/P0001 ,
		\u3_rp_reg[1]/NET0131 ,
		\u3_rp_reg[2]/NET0131 ,
		\u3_wp_reg[1]/NET0131 ,
		_w6293_
	);
	LUT2 #(
		.INIT('h1)
	) name4147 (
		_w6292_,
		_w6293_,
		_w6294_
	);
	LUT4 #(
		.INIT('h0ee0)
	) name4148 (
		\u13_occ0_r_reg[2]/NET0131 ,
		\u13_occ0_r_reg[3]/NET0131 ,
		\u3_rp_reg[1]/NET0131 ,
		\u3_wp_reg[0]/P0001 ,
		_w6295_
	);
	LUT2 #(
		.INIT('h2)
	) name4149 (
		\u3_rp_reg[0]/P0001 ,
		_w6295_,
		_w6296_
	);
	LUT3 #(
		.INIT('h80)
	) name4150 (
		\u3_rp_reg[0]/P0001 ,
		\u3_rp_reg[1]/NET0131 ,
		\u3_rp_reg[2]/NET0131 ,
		_w6297_
	);
	LUT4 #(
		.INIT('h0770)
	) name4151 (
		\u3_rp_reg[0]/P0001 ,
		\u3_rp_reg[1]/NET0131 ,
		\u3_rp_reg[2]/NET0131 ,
		\u3_wp_reg[1]/NET0131 ,
		_w6298_
	);
	LUT3 #(
		.INIT('h09)
	) name4152 (
		_w4225_,
		_w6297_,
		_w6298_,
		_w6299_
	);
	LUT3 #(
		.INIT('h10)
	) name4153 (
		_w6294_,
		_w6296_,
		_w6299_,
		_w6300_
	);
	LUT4 #(
		.INIT('hbde7)
	) name4154 (
		\u8_rp_reg[1]/NET0131 ,
		\u8_rp_reg[2]/NET0131 ,
		\u8_wp_reg[0]/P0001 ,
		\u8_wp_reg[1]/NET0131 ,
		_w6301_
	);
	LUT3 #(
		.INIT('ha8)
	) name4155 (
		\u8_rp_reg[0]/P0001 ,
		_w2156_,
		_w6301_,
		_w6302_
	);
	LUT4 #(
		.INIT('h8872)
	) name4156 (
		\u8_rp_reg[0]/P0001 ,
		_w2158_,
		_w4246_,
		_w4247_,
		_w6303_
	);
	LUT2 #(
		.INIT('h4)
	) name4157 (
		_w6302_,
		_w6303_,
		_w6304_
	);
	LUT3 #(
		.INIT('he2)
	) name4158 (
		\u0_slt9_r_reg[0]/P0001 ,
		\u2_ld_reg/P0001 ,
		\u8_dout_reg[1]/P0001 ,
		_w6305_
	);
	LUT3 #(
		.INIT('h80)
	) name4159 (
		\u12_i3_re_reg/NET0131 ,
		\u9_rp_reg[0]/P0001 ,
		\u9_rp_reg[1]/P0001 ,
		_w6306_
	);
	LUT4 #(
		.INIT('h4c80)
	) name4160 (
		\u12_i3_re_reg/NET0131 ,
		\u13_icc_r_reg[0]/NET0131 ,
		\u9_rp_reg[0]/P0001 ,
		\u9_rp_reg[1]/P0001 ,
		_w6307_
	);
	LUT3 #(
		.INIT('h80)
	) name4161 (
		\u10_rp_reg[0]/P0001 ,
		\u10_rp_reg[1]/P0001 ,
		\u12_i4_re_reg/P0001 ,
		_w6308_
	);
	LUT4 #(
		.INIT('h6c00)
	) name4162 (
		\u10_rp_reg[0]/P0001 ,
		\u10_rp_reg[1]/P0001 ,
		\u12_i4_re_reg/P0001 ,
		\u13_icc_r_reg[8]/NET0131 ,
		_w6309_
	);
	LUT3 #(
		.INIT('h80)
	) name4163 (
		\u11_rp_reg[0]/P0001 ,
		\u11_rp_reg[1]/P0001 ,
		\u12_i6_re_reg/NET0131 ,
		_w6310_
	);
	LUT4 #(
		.INIT('h6c00)
	) name4164 (
		\u11_rp_reg[0]/P0001 ,
		\u11_rp_reg[1]/P0001 ,
		\u12_i6_re_reg/NET0131 ,
		\u13_icc_r_reg[16]/NET0131 ,
		_w6311_
	);
	LUT3 #(
		.INIT('h28)
	) name4165 (
		\u13_icc_r_reg[0]/NET0131 ,
		\u9_rp_reg[2]/P0001 ,
		_w6306_,
		_w6312_
	);
	LUT3 #(
		.INIT('h48)
	) name4166 (
		\u11_rp_reg[2]/P0001 ,
		\u13_icc_r_reg[16]/NET0131 ,
		_w6310_,
		_w6313_
	);
	LUT3 #(
		.INIT('h48)
	) name4167 (
		\u10_rp_reg[2]/P0001 ,
		\u13_icc_r_reg[8]/NET0131 ,
		_w6308_,
		_w6314_
	);
	LUT3 #(
		.INIT('h48)
	) name4168 (
		\u2_res_cnt_reg[2]/P0001 ,
		\u2_sync_resume_reg/NET0131 ,
		_w4313_,
		_w6315_
	);
	LUT3 #(
		.INIT('h60)
	) name4169 (
		\u11_rp_reg[0]/P0001 ,
		\u12_i6_re_reg/NET0131 ,
		\u13_icc_r_reg[16]/NET0131 ,
		_w6316_
	);
	LUT4 #(
		.INIT('h0200)
	) name4170 (
		\u13_crac_r_reg[0]/NET0131 ,
		\wb_addr_i[2]_pad ,
		\wb_addr_i[3]_pad ,
		\wb_addr_i[4]_pad ,
		_w6317_
	);
	LUT4 #(
		.INIT('h0800)
	) name4171 (
		\u13_intm_r_reg[16]/NET0131 ,
		\wb_addr_i[2]_pad ,
		\wb_addr_i[3]_pad ,
		\wb_addr_i[4]_pad ,
		_w6318_
	);
	LUT2 #(
		.INIT('h1)
	) name4172 (
		_w6317_,
		_w6318_,
		_w6319_
	);
	LUT4 #(
		.INIT('h2000)
	) name4173 (
		\u13_ints_r_reg[16]/NET0131 ,
		\wb_addr_i[2]_pad ,
		\wb_addr_i[3]_pad ,
		\wb_addr_i[4]_pad ,
		_w6320_
	);
	LUT4 #(
		.INIT('h0080)
	) name4174 (
		\u13_icc_r_reg[16]/NET0131 ,
		\wb_addr_i[2]_pad ,
		\wb_addr_i[3]_pad ,
		\wb_addr_i[4]_pad ,
		_w6321_
	);
	LUT4 #(
		.INIT('h0008)
	) name4175 (
		\u13_occ0_r_reg[16]/NET0131 ,
		\wb_addr_i[2]_pad ,
		\wb_addr_i[3]_pad ,
		\wb_addr_i[4]_pad ,
		_w6322_
	);
	LUT3 #(
		.INIT('h01)
	) name4176 (
		_w6321_,
		_w6322_,
		_w6320_,
		_w6323_
	);
	LUT3 #(
		.INIT('h2a)
	) name4177 (
		_w4169_,
		_w6319_,
		_w6323_,
		_w6324_
	);
	LUT3 #(
		.INIT('h80)
	) name4178 (
		\u11_dout_reg[16]/P0001 ,
		_w4167_,
		_w4168_,
		_w6325_
	);
	LUT4 #(
		.INIT('h53ff)
	) name4179 (
		\u10_dout_reg[16]/P0001 ,
		\u9_dout_reg[16]/P0001 ,
		\wb_addr_i[2]_pad ,
		_w4166_,
		_w6326_
	);
	LUT2 #(
		.INIT('h4)
	) name4180 (
		_w6325_,
		_w6326_,
		_w6327_
	);
	LUT2 #(
		.INIT('hb)
	) name4181 (
		_w6324_,
		_w6327_,
		_w6328_
	);
	LUT4 #(
		.INIT('h0080)
	) name4182 (
		\u13_icc_r_reg[17]/NET0131 ,
		\wb_addr_i[2]_pad ,
		\wb_addr_i[3]_pad ,
		\wb_addr_i[4]_pad ,
		_w6329_
	);
	LUT4 #(
		.INIT('h0800)
	) name4183 (
		\u13_intm_r_reg[17]/NET0131 ,
		\wb_addr_i[2]_pad ,
		\wb_addr_i[3]_pad ,
		\wb_addr_i[4]_pad ,
		_w6330_
	);
	LUT2 #(
		.INIT('h1)
	) name4184 (
		_w6329_,
		_w6330_,
		_w6331_
	);
	LUT4 #(
		.INIT('h2000)
	) name4185 (
		\u13_ints_r_reg[17]/NET0131 ,
		\wb_addr_i[2]_pad ,
		\wb_addr_i[3]_pad ,
		\wb_addr_i[4]_pad ,
		_w6332_
	);
	LUT4 #(
		.INIT('h0200)
	) name4186 (
		\u13_crac_r_reg[1]/NET0131 ,
		\wb_addr_i[2]_pad ,
		\wb_addr_i[3]_pad ,
		\wb_addr_i[4]_pad ,
		_w6333_
	);
	LUT4 #(
		.INIT('h0008)
	) name4187 (
		\u13_occ0_r_reg[17]/NET0131 ,
		\wb_addr_i[2]_pad ,
		\wb_addr_i[3]_pad ,
		\wb_addr_i[4]_pad ,
		_w6334_
	);
	LUT3 #(
		.INIT('h01)
	) name4188 (
		_w6333_,
		_w6334_,
		_w6332_,
		_w6335_
	);
	LUT3 #(
		.INIT('h2a)
	) name4189 (
		_w4169_,
		_w6331_,
		_w6335_,
		_w6336_
	);
	LUT3 #(
		.INIT('h80)
	) name4190 (
		\u11_dout_reg[17]/P0001 ,
		_w4167_,
		_w4168_,
		_w6337_
	);
	LUT4 #(
		.INIT('h53ff)
	) name4191 (
		\u10_dout_reg[17]/P0001 ,
		\u9_dout_reg[17]/P0001 ,
		\wb_addr_i[2]_pad ,
		_w4166_,
		_w6338_
	);
	LUT2 #(
		.INIT('h4)
	) name4192 (
		_w6337_,
		_w6338_,
		_w6339_
	);
	LUT2 #(
		.INIT('hb)
	) name4193 (
		_w6336_,
		_w6339_,
		_w6340_
	);
	LUT4 #(
		.INIT('h0200)
	) name4194 (
		\u13_crac_r_reg[3]/NET0131 ,
		\wb_addr_i[2]_pad ,
		\wb_addr_i[3]_pad ,
		\wb_addr_i[4]_pad ,
		_w6341_
	);
	LUT4 #(
		.INIT('h0800)
	) name4195 (
		\u13_intm_r_reg[19]/NET0131 ,
		\wb_addr_i[2]_pad ,
		\wb_addr_i[3]_pad ,
		\wb_addr_i[4]_pad ,
		_w6342_
	);
	LUT2 #(
		.INIT('h1)
	) name4196 (
		_w6341_,
		_w6342_,
		_w6343_
	);
	LUT4 #(
		.INIT('h2000)
	) name4197 (
		\u13_ints_r_reg[19]/NET0131 ,
		\wb_addr_i[2]_pad ,
		\wb_addr_i[3]_pad ,
		\wb_addr_i[4]_pad ,
		_w6344_
	);
	LUT4 #(
		.INIT('h0080)
	) name4198 (
		\u13_icc_r_reg[19]/NET0131 ,
		\wb_addr_i[2]_pad ,
		\wb_addr_i[3]_pad ,
		\wb_addr_i[4]_pad ,
		_w6345_
	);
	LUT4 #(
		.INIT('h0008)
	) name4199 (
		\u13_occ0_r_reg[19]/NET0131 ,
		\wb_addr_i[2]_pad ,
		\wb_addr_i[3]_pad ,
		\wb_addr_i[4]_pad ,
		_w6346_
	);
	LUT3 #(
		.INIT('h01)
	) name4200 (
		_w6345_,
		_w6346_,
		_w6344_,
		_w6347_
	);
	LUT3 #(
		.INIT('h2a)
	) name4201 (
		_w4169_,
		_w6343_,
		_w6347_,
		_w6348_
	);
	LUT3 #(
		.INIT('h80)
	) name4202 (
		\u11_dout_reg[19]/P0001 ,
		_w4167_,
		_w4168_,
		_w6349_
	);
	LUT4 #(
		.INIT('h53ff)
	) name4203 (
		\u10_dout_reg[19]/P0001 ,
		\u9_dout_reg[19]/P0001 ,
		\wb_addr_i[2]_pad ,
		_w4166_,
		_w6350_
	);
	LUT2 #(
		.INIT('h4)
	) name4204 (
		_w6349_,
		_w6350_,
		_w6351_
	);
	LUT2 #(
		.INIT('hb)
	) name4205 (
		_w6348_,
		_w6351_,
		_w6352_
	);
	LUT3 #(
		.INIT('h48)
	) name4206 (
		\u12_i3_re_reg/NET0131 ,
		\u13_icc_r_reg[0]/NET0131 ,
		\u9_rp_reg[0]/P0001 ,
		_w6353_
	);
	LUT4 #(
		.INIT('h0080)
	) name4207 (
		\u13_icc_r_reg[20]/NET0131 ,
		\wb_addr_i[2]_pad ,
		\wb_addr_i[3]_pad ,
		\wb_addr_i[4]_pad ,
		_w6354_
	);
	LUT4 #(
		.INIT('h0800)
	) name4208 (
		\u13_intm_r_reg[20]/NET0131 ,
		\wb_addr_i[2]_pad ,
		\wb_addr_i[3]_pad ,
		\wb_addr_i[4]_pad ,
		_w6355_
	);
	LUT2 #(
		.INIT('h1)
	) name4209 (
		_w6354_,
		_w6355_,
		_w6356_
	);
	LUT4 #(
		.INIT('h2000)
	) name4210 (
		\u13_ints_r_reg[20]/NET0131 ,
		\wb_addr_i[2]_pad ,
		\wb_addr_i[3]_pad ,
		\wb_addr_i[4]_pad ,
		_w6357_
	);
	LUT4 #(
		.INIT('h0200)
	) name4211 (
		\u13_crac_r_reg[4]/NET0131 ,
		\wb_addr_i[2]_pad ,
		\wb_addr_i[3]_pad ,
		\wb_addr_i[4]_pad ,
		_w6358_
	);
	LUT4 #(
		.INIT('h0008)
	) name4212 (
		\u13_occ0_r_reg[20]/NET0131 ,
		\wb_addr_i[2]_pad ,
		\wb_addr_i[3]_pad ,
		\wb_addr_i[4]_pad ,
		_w6359_
	);
	LUT3 #(
		.INIT('h01)
	) name4213 (
		_w6358_,
		_w6359_,
		_w6357_,
		_w6360_
	);
	LUT3 #(
		.INIT('h2a)
	) name4214 (
		_w4169_,
		_w6356_,
		_w6360_,
		_w6361_
	);
	LUT3 #(
		.INIT('h80)
	) name4215 (
		\u11_dout_reg[20]/P0001 ,
		_w4167_,
		_w4168_,
		_w6362_
	);
	LUT4 #(
		.INIT('h53ff)
	) name4216 (
		\u10_dout_reg[20]/P0001 ,
		\u9_dout_reg[20]/P0001 ,
		\wb_addr_i[2]_pad ,
		_w4166_,
		_w6363_
	);
	LUT2 #(
		.INIT('h4)
	) name4217 (
		_w6362_,
		_w6363_,
		_w6364_
	);
	LUT2 #(
		.INIT('hb)
	) name4218 (
		_w6361_,
		_w6364_,
		_w6365_
	);
	LUT4 #(
		.INIT('h0080)
	) name4219 (
		\u13_icc_r_reg[21]/NET0131 ,
		\wb_addr_i[2]_pad ,
		\wb_addr_i[3]_pad ,
		\wb_addr_i[4]_pad ,
		_w6366_
	);
	LUT4 #(
		.INIT('h0800)
	) name4220 (
		\u13_intm_r_reg[21]/NET0131 ,
		\wb_addr_i[2]_pad ,
		\wb_addr_i[3]_pad ,
		\wb_addr_i[4]_pad ,
		_w6367_
	);
	LUT2 #(
		.INIT('h1)
	) name4221 (
		_w6366_,
		_w6367_,
		_w6368_
	);
	LUT4 #(
		.INIT('h2000)
	) name4222 (
		\u13_ints_r_reg[21]/NET0131 ,
		\wb_addr_i[2]_pad ,
		\wb_addr_i[3]_pad ,
		\wb_addr_i[4]_pad ,
		_w6369_
	);
	LUT4 #(
		.INIT('h0200)
	) name4223 (
		\u13_crac_r_reg[5]/NET0131 ,
		\wb_addr_i[2]_pad ,
		\wb_addr_i[3]_pad ,
		\wb_addr_i[4]_pad ,
		_w6370_
	);
	LUT4 #(
		.INIT('h0008)
	) name4224 (
		\u13_occ0_r_reg[21]/NET0131 ,
		\wb_addr_i[2]_pad ,
		\wb_addr_i[3]_pad ,
		\wb_addr_i[4]_pad ,
		_w6371_
	);
	LUT3 #(
		.INIT('h01)
	) name4225 (
		_w6370_,
		_w6371_,
		_w6369_,
		_w6372_
	);
	LUT3 #(
		.INIT('h2a)
	) name4226 (
		_w4169_,
		_w6368_,
		_w6372_,
		_w6373_
	);
	LUT3 #(
		.INIT('h80)
	) name4227 (
		\u11_dout_reg[21]/P0001 ,
		_w4167_,
		_w4168_,
		_w6374_
	);
	LUT4 #(
		.INIT('h53ff)
	) name4228 (
		\u10_dout_reg[21]/P0001 ,
		\u9_dout_reg[21]/P0001 ,
		\wb_addr_i[2]_pad ,
		_w4166_,
		_w6375_
	);
	LUT2 #(
		.INIT('h4)
	) name4229 (
		_w6374_,
		_w6375_,
		_w6376_
	);
	LUT2 #(
		.INIT('hb)
	) name4230 (
		_w6373_,
		_w6376_,
		_w6377_
	);
	LUT4 #(
		.INIT('h0080)
	) name4231 (
		\u13_icc_r_reg[22]/NET0131 ,
		\wb_addr_i[2]_pad ,
		\wb_addr_i[3]_pad ,
		\wb_addr_i[4]_pad ,
		_w6378_
	);
	LUT4 #(
		.INIT('h0800)
	) name4232 (
		\u13_intm_r_reg[22]/NET0131 ,
		\wb_addr_i[2]_pad ,
		\wb_addr_i[3]_pad ,
		\wb_addr_i[4]_pad ,
		_w6379_
	);
	LUT2 #(
		.INIT('h1)
	) name4233 (
		_w6378_,
		_w6379_,
		_w6380_
	);
	LUT4 #(
		.INIT('h2000)
	) name4234 (
		\u13_ints_r_reg[22]/NET0131 ,
		\wb_addr_i[2]_pad ,
		\wb_addr_i[3]_pad ,
		\wb_addr_i[4]_pad ,
		_w6381_
	);
	LUT4 #(
		.INIT('h0200)
	) name4235 (
		\u13_crac_r_reg[6]/NET0131 ,
		\wb_addr_i[2]_pad ,
		\wb_addr_i[3]_pad ,
		\wb_addr_i[4]_pad ,
		_w6382_
	);
	LUT4 #(
		.INIT('h0008)
	) name4236 (
		\u13_occ0_r_reg[22]/NET0131 ,
		\wb_addr_i[2]_pad ,
		\wb_addr_i[3]_pad ,
		\wb_addr_i[4]_pad ,
		_w6383_
	);
	LUT3 #(
		.INIT('h01)
	) name4237 (
		_w6382_,
		_w6383_,
		_w6381_,
		_w6384_
	);
	LUT3 #(
		.INIT('h2a)
	) name4238 (
		_w4169_,
		_w6380_,
		_w6384_,
		_w6385_
	);
	LUT3 #(
		.INIT('h80)
	) name4239 (
		\u11_dout_reg[22]/P0001 ,
		_w4167_,
		_w4168_,
		_w6386_
	);
	LUT4 #(
		.INIT('h53ff)
	) name4240 (
		\u10_dout_reg[22]/P0001 ,
		\u9_dout_reg[22]/P0001 ,
		\wb_addr_i[2]_pad ,
		_w4166_,
		_w6387_
	);
	LUT2 #(
		.INIT('h4)
	) name4241 (
		_w6386_,
		_w6387_,
		_w6388_
	);
	LUT2 #(
		.INIT('hb)
	) name4242 (
		_w6385_,
		_w6388_,
		_w6389_
	);
	LUT4 #(
		.INIT('h2000)
	) name4243 (
		\u13_ints_r_reg[23]/NET0131 ,
		\wb_addr_i[2]_pad ,
		\wb_addr_i[3]_pad ,
		\wb_addr_i[4]_pad ,
		_w6390_
	);
	LUT4 #(
		.INIT('h0800)
	) name4244 (
		\u13_intm_r_reg[23]/NET0131 ,
		\wb_addr_i[2]_pad ,
		\wb_addr_i[3]_pad ,
		\wb_addr_i[4]_pad ,
		_w6391_
	);
	LUT4 #(
		.INIT('h0008)
	) name4245 (
		\u13_occ0_r_reg[23]/NET0131 ,
		\wb_addr_i[2]_pad ,
		\wb_addr_i[3]_pad ,
		\wb_addr_i[4]_pad ,
		_w6392_
	);
	LUT4 #(
		.INIT('h0080)
	) name4246 (
		\u13_icc_r_reg[23]/NET0131 ,
		\wb_addr_i[2]_pad ,
		\wb_addr_i[3]_pad ,
		\wb_addr_i[4]_pad ,
		_w6393_
	);
	LUT4 #(
		.INIT('h0001)
	) name4247 (
		_w6390_,
		_w6391_,
		_w6392_,
		_w6393_,
		_w6394_
	);
	LUT2 #(
		.INIT('h2)
	) name4248 (
		_w4169_,
		_w6394_,
		_w6395_
	);
	LUT3 #(
		.INIT('h80)
	) name4249 (
		\u10_dout_reg[23]/P0001 ,
		\wb_addr_i[2]_pad ,
		_w4166_,
		_w6396_
	);
	LUT3 #(
		.INIT('h20)
	) name4250 (
		\u9_dout_reg[23]/P0001 ,
		\wb_addr_i[2]_pad ,
		_w4166_,
		_w6397_
	);
	LUT3 #(
		.INIT('h80)
	) name4251 (
		\u11_dout_reg[23]/P0001 ,
		_w4167_,
		_w4168_,
		_w6398_
	);
	LUT3 #(
		.INIT('h01)
	) name4252 (
		_w6397_,
		_w6398_,
		_w6396_,
		_w6399_
	);
	LUT2 #(
		.INIT('hb)
	) name4253 (
		_w6395_,
		_w6399_,
		_w6400_
	);
	LUT3 #(
		.INIT('h60)
	) name4254 (
		\u10_rp_reg[0]/P0001 ,
		\u12_i4_re_reg/P0001 ,
		\u13_icc_r_reg[8]/NET0131 ,
		_w6401_
	);
	LUT4 #(
		.INIT('h0200)
	) name4255 (
		\u13_crac_r_reg[2]/NET0131 ,
		\wb_addr_i[2]_pad ,
		\wb_addr_i[3]_pad ,
		\wb_addr_i[4]_pad ,
		_w6402_
	);
	LUT4 #(
		.INIT('h0800)
	) name4256 (
		\u13_intm_r_reg[18]/NET0131 ,
		\wb_addr_i[2]_pad ,
		\wb_addr_i[3]_pad ,
		\wb_addr_i[4]_pad ,
		_w6403_
	);
	LUT2 #(
		.INIT('h1)
	) name4257 (
		_w6402_,
		_w6403_,
		_w6404_
	);
	LUT4 #(
		.INIT('h2000)
	) name4258 (
		\u13_ints_r_reg[18]/NET0131 ,
		\wb_addr_i[2]_pad ,
		\wb_addr_i[3]_pad ,
		\wb_addr_i[4]_pad ,
		_w6405_
	);
	LUT4 #(
		.INIT('h0080)
	) name4259 (
		\u13_icc_r_reg[18]/NET0131 ,
		\wb_addr_i[2]_pad ,
		\wb_addr_i[3]_pad ,
		\wb_addr_i[4]_pad ,
		_w6406_
	);
	LUT4 #(
		.INIT('h0008)
	) name4260 (
		\u13_occ0_r_reg[18]/NET0131 ,
		\wb_addr_i[2]_pad ,
		\wb_addr_i[3]_pad ,
		\wb_addr_i[4]_pad ,
		_w6407_
	);
	LUT3 #(
		.INIT('h01)
	) name4261 (
		_w6406_,
		_w6407_,
		_w6405_,
		_w6408_
	);
	LUT3 #(
		.INIT('h2a)
	) name4262 (
		_w4169_,
		_w6404_,
		_w6408_,
		_w6409_
	);
	LUT3 #(
		.INIT('h80)
	) name4263 (
		\u11_dout_reg[18]/P0001 ,
		_w4167_,
		_w4168_,
		_w6410_
	);
	LUT4 #(
		.INIT('h53ff)
	) name4264 (
		\u10_dout_reg[18]/P0001 ,
		\u9_dout_reg[18]/P0001 ,
		\wb_addr_i[2]_pad ,
		_w4166_,
		_w6411_
	);
	LUT2 #(
		.INIT('h4)
	) name4265 (
		_w6410_,
		_w6411_,
		_w6412_
	);
	LUT2 #(
		.INIT('hb)
	) name4266 (
		_w6409_,
		_w6412_,
		_w6413_
	);
	LUT3 #(
		.INIT('h14)
	) name4267 (
		\u2_bit_clk_e_reg/P0001 ,
		\u2_to_cnt_reg[4]/NET0131 ,
		_w4325_,
		_w6414_
	);
	LUT4 #(
		.INIT('h1450)
	) name4268 (
		\u2_bit_clk_e_reg/P0001 ,
		\u2_to_cnt_reg[4]/NET0131 ,
		\u2_to_cnt_reg[5]/NET0131 ,
		_w4325_,
		_w6415_
	);
	LUT4 #(
		.INIT('h1540)
	) name4269 (
		\u2_bit_clk_e_reg/P0001 ,
		\u2_to_cnt_reg[0]/NET0131 ,
		\u2_to_cnt_reg[1]/NET0131 ,
		\u2_to_cnt_reg[2]/NET0131 ,
		_w6416_
	);
	LUT3 #(
		.INIT('hec)
	) name4270 (
		\u12_i3_re_reg/NET0131 ,
		\u23_int_set_reg[1]/NET0131 ,
		\u9_empty_reg/P0001 ,
		_w6417_
	);
	LUT3 #(
		.INIT('hf8)
	) name4271 (
		\u10_empty_reg/P0001 ,
		\u12_i4_re_reg/P0001 ,
		\u24_int_set_reg[1]/NET0131 ,
		_w6418_
	);
	LUT3 #(
		.INIT('hf8)
	) name4272 (
		\u11_empty_reg/P0001 ,
		\u12_i6_re_reg/NET0131 ,
		\u25_int_set_reg[1]/NET0131 ,
		_w6419_
	);
	LUT4 #(
		.INIT('h4888)
	) name4273 (
		\u2_res_cnt_reg[0]/P0001 ,
		\u2_sync_resume_reg/NET0131 ,
		_w3862_,
		_w3863_,
		_w6420_
	);
	LUT3 #(
		.INIT('h80)
	) name4274 (
		wb_cyc_i_pad,
		wb_stb_i_pad,
		wb_we_i_pad,
		_w6421_
	);
	LUT4 #(
		.INIT('h8000)
	) name4275 (
		\u12_we1_reg/P0001 ,
		wb_cyc_i_pad,
		wb_stb_i_pad,
		wb_we_i_pad,
		_w6422_
	);
	LUT4 #(
		.INIT('h4000)
	) name4276 (
		\u12_we2_reg/P0001 ,
		_w4165_,
		_w4167_,
		_w6422_,
		_w6423_
	);
	LUT4 #(
		.INIT('h4000)
	) name4277 (
		\u12_we2_reg/P0001 ,
		_w4165_,
		_w4179_,
		_w6422_,
		_w6424_
	);
	LUT4 #(
		.INIT('h4000)
	) name4278 (
		\u12_we2_reg/P0001 ,
		_w4165_,
		_w4176_,
		_w6422_,
		_w6425_
	);
	LUT4 #(
		.INIT('h4000)
	) name4279 (
		\u12_we2_reg/P0001 ,
		_w4165_,
		_w4170_,
		_w6422_,
		_w6426_
	);
	LUT4 #(
		.INIT('h4000)
	) name4280 (
		\u12_we2_reg/P0001 ,
		_w4165_,
		_w4181_,
		_w6422_,
		_w6427_
	);
	LUT4 #(
		.INIT('h2000)
	) name4281 (
		\u13_ints_r_reg[24]/NET0131 ,
		\wb_addr_i[2]_pad ,
		\wb_addr_i[3]_pad ,
		\wb_addr_i[4]_pad ,
		_w6428_
	);
	LUT4 #(
		.INIT('h0008)
	) name4282 (
		\u13_occ0_r_reg[24]/NET0131 ,
		\wb_addr_i[2]_pad ,
		\wb_addr_i[3]_pad ,
		\wb_addr_i[4]_pad ,
		_w6429_
	);
	LUT4 #(
		.INIT('h0800)
	) name4283 (
		\u13_intm_r_reg[24]/NET0131 ,
		\wb_addr_i[2]_pad ,
		\wb_addr_i[3]_pad ,
		\wb_addr_i[4]_pad ,
		_w6430_
	);
	LUT3 #(
		.INIT('h01)
	) name4284 (
		_w6429_,
		_w6430_,
		_w6428_,
		_w6431_
	);
	LUT2 #(
		.INIT('h2)
	) name4285 (
		_w4169_,
		_w6431_,
		_w6432_
	);
	LUT3 #(
		.INIT('h80)
	) name4286 (
		\u10_dout_reg[24]/P0001 ,
		\wb_addr_i[2]_pad ,
		_w4166_,
		_w6433_
	);
	LUT3 #(
		.INIT('h20)
	) name4287 (
		\u9_dout_reg[24]/P0001 ,
		\wb_addr_i[2]_pad ,
		_w4166_,
		_w6434_
	);
	LUT3 #(
		.INIT('h80)
	) name4288 (
		\u11_dout_reg[24]/P0001 ,
		_w4167_,
		_w4168_,
		_w6435_
	);
	LUT3 #(
		.INIT('h01)
	) name4289 (
		_w6434_,
		_w6435_,
		_w6433_,
		_w6436_
	);
	LUT2 #(
		.INIT('hb)
	) name4290 (
		_w6432_,
		_w6436_,
		_w6437_
	);
	LUT4 #(
		.INIT('h2000)
	) name4291 (
		\u13_ints_r_reg[25]/NET0131 ,
		\wb_addr_i[2]_pad ,
		\wb_addr_i[3]_pad ,
		\wb_addr_i[4]_pad ,
		_w6438_
	);
	LUT4 #(
		.INIT('h0008)
	) name4292 (
		\u13_occ0_r_reg[25]/NET0131 ,
		\wb_addr_i[2]_pad ,
		\wb_addr_i[3]_pad ,
		\wb_addr_i[4]_pad ,
		_w6439_
	);
	LUT4 #(
		.INIT('h0800)
	) name4293 (
		\u13_intm_r_reg[25]/NET0131 ,
		\wb_addr_i[2]_pad ,
		\wb_addr_i[3]_pad ,
		\wb_addr_i[4]_pad ,
		_w6440_
	);
	LUT3 #(
		.INIT('h01)
	) name4294 (
		_w6439_,
		_w6440_,
		_w6438_,
		_w6441_
	);
	LUT2 #(
		.INIT('h2)
	) name4295 (
		_w4169_,
		_w6441_,
		_w6442_
	);
	LUT3 #(
		.INIT('h80)
	) name4296 (
		\u10_dout_reg[25]/P0001 ,
		\wb_addr_i[2]_pad ,
		_w4166_,
		_w6443_
	);
	LUT3 #(
		.INIT('h20)
	) name4297 (
		\u9_dout_reg[25]/P0001 ,
		\wb_addr_i[2]_pad ,
		_w4166_,
		_w6444_
	);
	LUT3 #(
		.INIT('h80)
	) name4298 (
		\u11_dout_reg[25]/P0001 ,
		_w4167_,
		_w4168_,
		_w6445_
	);
	LUT3 #(
		.INIT('h01)
	) name4299 (
		_w6444_,
		_w6445_,
		_w6443_,
		_w6446_
	);
	LUT2 #(
		.INIT('hb)
	) name4300 (
		_w6442_,
		_w6446_,
		_w6447_
	);
	LUT4 #(
		.INIT('h2000)
	) name4301 (
		\u13_ints_r_reg[26]/NET0131 ,
		\wb_addr_i[2]_pad ,
		\wb_addr_i[3]_pad ,
		\wb_addr_i[4]_pad ,
		_w6448_
	);
	LUT4 #(
		.INIT('h0008)
	) name4302 (
		\u13_occ0_r_reg[26]/NET0131 ,
		\wb_addr_i[2]_pad ,
		\wb_addr_i[3]_pad ,
		\wb_addr_i[4]_pad ,
		_w6449_
	);
	LUT4 #(
		.INIT('h0800)
	) name4303 (
		\u13_intm_r_reg[26]/NET0131 ,
		\wb_addr_i[2]_pad ,
		\wb_addr_i[3]_pad ,
		\wb_addr_i[4]_pad ,
		_w6450_
	);
	LUT3 #(
		.INIT('h01)
	) name4304 (
		_w6449_,
		_w6450_,
		_w6448_,
		_w6451_
	);
	LUT2 #(
		.INIT('h2)
	) name4305 (
		_w4169_,
		_w6451_,
		_w6452_
	);
	LUT3 #(
		.INIT('h80)
	) name4306 (
		\u10_dout_reg[26]/P0001 ,
		\wb_addr_i[2]_pad ,
		_w4166_,
		_w6453_
	);
	LUT3 #(
		.INIT('h20)
	) name4307 (
		\u9_dout_reg[26]/P0001 ,
		\wb_addr_i[2]_pad ,
		_w4166_,
		_w6454_
	);
	LUT3 #(
		.INIT('h80)
	) name4308 (
		\u11_dout_reg[26]/P0001 ,
		_w4167_,
		_w4168_,
		_w6455_
	);
	LUT3 #(
		.INIT('h01)
	) name4309 (
		_w6454_,
		_w6455_,
		_w6453_,
		_w6456_
	);
	LUT2 #(
		.INIT('hb)
	) name4310 (
		_w6452_,
		_w6456_,
		_w6457_
	);
	LUT4 #(
		.INIT('h2000)
	) name4311 (
		\u13_ints_r_reg[27]/NET0131 ,
		\wb_addr_i[2]_pad ,
		\wb_addr_i[3]_pad ,
		\wb_addr_i[4]_pad ,
		_w6458_
	);
	LUT4 #(
		.INIT('h0008)
	) name4312 (
		\u13_occ0_r_reg[27]/NET0131 ,
		\wb_addr_i[2]_pad ,
		\wb_addr_i[3]_pad ,
		\wb_addr_i[4]_pad ,
		_w6459_
	);
	LUT4 #(
		.INIT('h0800)
	) name4313 (
		\u13_intm_r_reg[27]/NET0131 ,
		\wb_addr_i[2]_pad ,
		\wb_addr_i[3]_pad ,
		\wb_addr_i[4]_pad ,
		_w6460_
	);
	LUT3 #(
		.INIT('h01)
	) name4314 (
		_w6459_,
		_w6460_,
		_w6458_,
		_w6461_
	);
	LUT2 #(
		.INIT('h2)
	) name4315 (
		_w4169_,
		_w6461_,
		_w6462_
	);
	LUT3 #(
		.INIT('h80)
	) name4316 (
		\u10_dout_reg[27]/P0001 ,
		\wb_addr_i[2]_pad ,
		_w4166_,
		_w6463_
	);
	LUT3 #(
		.INIT('h20)
	) name4317 (
		\u9_dout_reg[27]/P0001 ,
		\wb_addr_i[2]_pad ,
		_w4166_,
		_w6464_
	);
	LUT3 #(
		.INIT('h80)
	) name4318 (
		\u11_dout_reg[27]/P0001 ,
		_w4167_,
		_w4168_,
		_w6465_
	);
	LUT3 #(
		.INIT('h01)
	) name4319 (
		_w6464_,
		_w6465_,
		_w6463_,
		_w6466_
	);
	LUT2 #(
		.INIT('hb)
	) name4320 (
		_w6462_,
		_w6466_,
		_w6467_
	);
	LUT4 #(
		.INIT('h2000)
	) name4321 (
		\u13_ints_r_reg[28]/NET0131 ,
		\wb_addr_i[2]_pad ,
		\wb_addr_i[3]_pad ,
		\wb_addr_i[4]_pad ,
		_w6468_
	);
	LUT4 #(
		.INIT('h0008)
	) name4322 (
		\u13_occ0_r_reg[28]/NET0131 ,
		\wb_addr_i[2]_pad ,
		\wb_addr_i[3]_pad ,
		\wb_addr_i[4]_pad ,
		_w6469_
	);
	LUT4 #(
		.INIT('h0800)
	) name4323 (
		\u13_intm_r_reg[28]/NET0131 ,
		\wb_addr_i[2]_pad ,
		\wb_addr_i[3]_pad ,
		\wb_addr_i[4]_pad ,
		_w6470_
	);
	LUT3 #(
		.INIT('h01)
	) name4324 (
		_w6469_,
		_w6470_,
		_w6468_,
		_w6471_
	);
	LUT2 #(
		.INIT('h2)
	) name4325 (
		_w4169_,
		_w6471_,
		_w6472_
	);
	LUT3 #(
		.INIT('h80)
	) name4326 (
		\u10_dout_reg[28]/P0001 ,
		\wb_addr_i[2]_pad ,
		_w4166_,
		_w6473_
	);
	LUT3 #(
		.INIT('h20)
	) name4327 (
		\u9_dout_reg[28]/P0001 ,
		\wb_addr_i[2]_pad ,
		_w4166_,
		_w6474_
	);
	LUT3 #(
		.INIT('h80)
	) name4328 (
		\u11_dout_reg[28]/P0001 ,
		_w4167_,
		_w4168_,
		_w6475_
	);
	LUT3 #(
		.INIT('h01)
	) name4329 (
		_w6474_,
		_w6475_,
		_w6473_,
		_w6476_
	);
	LUT2 #(
		.INIT('hb)
	) name4330 (
		_w6472_,
		_w6476_,
		_w6477_
	);
	LUT4 #(
		.INIT('h0008)
	) name4331 (
		\u13_occ0_r_reg[29]/NET0131 ,
		\wb_addr_i[2]_pad ,
		\wb_addr_i[3]_pad ,
		\wb_addr_i[4]_pad ,
		_w6478_
	);
	LUT4 #(
		.INIT('h007f)
	) name4332 (
		\u11_dout_reg[29]/P0001 ,
		_w4167_,
		_w4168_,
		_w6478_,
		_w6479_
	);
	LUT4 #(
		.INIT('h53ff)
	) name4333 (
		\u10_dout_reg[29]/P0001 ,
		\u9_dout_reg[29]/P0001 ,
		\wb_addr_i[2]_pad ,
		_w4166_,
		_w6480_
	);
	LUT2 #(
		.INIT('h7)
	) name4334 (
		_w6479_,
		_w6480_,
		_w6481_
	);
	LUT4 #(
		.INIT('h0008)
	) name4335 (
		\u13_occ0_r_reg[30]/NET0131 ,
		\wb_addr_i[2]_pad ,
		\wb_addr_i[3]_pad ,
		\wb_addr_i[4]_pad ,
		_w6482_
	);
	LUT4 #(
		.INIT('h007f)
	) name4336 (
		\u11_dout_reg[30]/P0001 ,
		_w4167_,
		_w4168_,
		_w6482_,
		_w6483_
	);
	LUT4 #(
		.INIT('h53ff)
	) name4337 (
		\u10_dout_reg[30]/P0001 ,
		\u9_dout_reg[30]/P0001 ,
		\wb_addr_i[2]_pad ,
		_w4166_,
		_w6484_
	);
	LUT2 #(
		.INIT('h7)
	) name4338 (
		_w6483_,
		_w6484_,
		_w6485_
	);
	LUT3 #(
		.INIT('h80)
	) name4339 (
		\u10_dout_reg[31]/P0001 ,
		\wb_addr_i[2]_pad ,
		_w4166_,
		_w6486_
	);
	LUT4 #(
		.INIT('h0200)
	) name4340 (
		\u13_crac_r_reg[7]/NET0131 ,
		\wb_addr_i[2]_pad ,
		\wb_addr_i[3]_pad ,
		\wb_addr_i[4]_pad ,
		_w6487_
	);
	LUT4 #(
		.INIT('h0008)
	) name4341 (
		\u13_occ0_r_reg[31]/NET0131 ,
		\wb_addr_i[2]_pad ,
		\wb_addr_i[3]_pad ,
		\wb_addr_i[4]_pad ,
		_w6488_
	);
	LUT2 #(
		.INIT('h1)
	) name4342 (
		_w6487_,
		_w6488_,
		_w6489_
	);
	LUT3 #(
		.INIT('h80)
	) name4343 (
		\u11_dout_reg[31]/P0001 ,
		_w4167_,
		_w4168_,
		_w6490_
	);
	LUT3 #(
		.INIT('h20)
	) name4344 (
		\u9_dout_reg[31]/P0001 ,
		\wb_addr_i[2]_pad ,
		_w4166_,
		_w6491_
	);
	LUT4 #(
		.INIT('hfeff)
	) name4345 (
		_w6486_,
		_w6490_,
		_w6491_,
		_w6489_,
		_w6492_
	);
	LUT3 #(
		.INIT('h48)
	) name4346 (
		\u2_res_cnt_reg[1]/P0001 ,
		\u2_sync_resume_reg/NET0131 ,
		_w4312_,
		_w6493_
	);
	LUT4 #(
		.INIT('h7f80)
	) name4347 (
		\u2_cnt_reg[0]/NET0131 ,
		\u2_cnt_reg[1]/NET0131 ,
		\u2_cnt_reg[2]/NET0131 ,
		\u2_cnt_reg[3]/NET0131 ,
		_w6494_
	);
	LUT2 #(
		.INIT('he)
	) name4348 (
		suspended_o_pad,
		_w6494_,
		_w6495_
	);
	LUT4 #(
		.INIT('h135f)
	) name4349 (
		\u13_intm_r_reg[10]/NET0131 ,
		\u13_intm_r_reg[9]/NET0131 ,
		\u13_ints_r_reg[10]/NET0131 ,
		\u13_ints_r_reg[9]/NET0131 ,
		_w6496_
	);
	LUT4 #(
		.INIT('h135f)
	) name4350 (
		\u13_intm_r_reg[21]/NET0131 ,
		\u13_intm_r_reg[4]/NET0131 ,
		\u13_ints_r_reg[21]/NET0131 ,
		\u13_ints_r_reg[4]/NET0131 ,
		_w6497_
	);
	LUT4 #(
		.INIT('h135f)
	) name4351 (
		\u13_intm_r_reg[12]/NET0131 ,
		\u13_intm_r_reg[22]/NET0131 ,
		\u13_ints_r_reg[12]/NET0131 ,
		\u13_ints_r_reg[22]/NET0131 ,
		_w6498_
	);
	LUT4 #(
		.INIT('h135f)
	) name4352 (
		\u13_intm_r_reg[19]/NET0131 ,
		\u13_intm_r_reg[27]/NET0131 ,
		\u13_ints_r_reg[19]/NET0131 ,
		\u13_ints_r_reg[27]/NET0131 ,
		_w6499_
	);
	LUT4 #(
		.INIT('h8000)
	) name4353 (
		_w6498_,
		_w6499_,
		_w6496_,
		_w6497_,
		_w6500_
	);
	LUT2 #(
		.INIT('h8)
	) name4354 (
		\u13_intm_r_reg[3]/NET0131 ,
		\u13_ints_r_reg[3]/NET0131 ,
		_w6501_
	);
	LUT4 #(
		.INIT('h135f)
	) name4355 (
		\u13_intm_r_reg[18]/NET0131 ,
		\u13_intm_r_reg[25]/NET0131 ,
		\u13_ints_r_reg[18]/NET0131 ,
		\u13_ints_r_reg[25]/NET0131 ,
		_w6502_
	);
	LUT4 #(
		.INIT('h135f)
	) name4356 (
		\u13_intm_r_reg[16]/NET0131 ,
		\u13_intm_r_reg[17]/NET0131 ,
		\u13_ints_r_reg[16]/NET0131 ,
		\u13_ints_r_reg[17]/NET0131 ,
		_w6503_
	);
	LUT4 #(
		.INIT('h135f)
	) name4357 (
		\u13_intm_r_reg[20]/NET0131 ,
		\u13_intm_r_reg[2]/NET0131 ,
		\u13_ints_r_reg[20]/NET0131 ,
		\u13_ints_r_reg[2]/NET0131 ,
		_w6504_
	);
	LUT4 #(
		.INIT('h4000)
	) name4358 (
		_w6501_,
		_w6503_,
		_w6504_,
		_w6502_,
		_w6505_
	);
	LUT4 #(
		.INIT('h135f)
	) name4359 (
		\u13_intm_r_reg[15]/NET0131 ,
		\u13_intm_r_reg[26]/NET0131 ,
		\u13_ints_r_reg[15]/NET0131 ,
		\u13_ints_r_reg[26]/NET0131 ,
		_w6506_
	);
	LUT4 #(
		.INIT('h135f)
	) name4360 (
		\u13_intm_r_reg[0]/NET0131 ,
		\u13_intm_r_reg[28]/NET0131 ,
		\u13_ints_r_reg[0]/NET0131 ,
		\u13_ints_r_reg[28]/NET0131 ,
		_w6507_
	);
	LUT4 #(
		.INIT('h135f)
	) name4361 (
		\u13_intm_r_reg[13]/NET0131 ,
		\u13_intm_r_reg[1]/NET0131 ,
		\u13_ints_r_reg[13]/NET0131 ,
		\u13_ints_r_reg[1]/NET0131 ,
		_w6508_
	);
	LUT3 #(
		.INIT('h80)
	) name4362 (
		_w6506_,
		_w6507_,
		_w6508_,
		_w6509_
	);
	LUT4 #(
		.INIT('h135f)
	) name4363 (
		\u13_intm_r_reg[23]/NET0131 ,
		\u13_intm_r_reg[7]/NET0131 ,
		\u13_ints_r_reg[23]/NET0131 ,
		\u13_ints_r_reg[7]/NET0131 ,
		_w6510_
	);
	LUT4 #(
		.INIT('h135f)
	) name4364 (
		\u13_intm_r_reg[14]/NET0131 ,
		\u13_intm_r_reg[24]/NET0131 ,
		\u13_ints_r_reg[14]/NET0131 ,
		\u13_ints_r_reg[24]/NET0131 ,
		_w6511_
	);
	LUT4 #(
		.INIT('h135f)
	) name4365 (
		\u13_intm_r_reg[11]/NET0131 ,
		\u13_intm_r_reg[6]/NET0131 ,
		\u13_ints_r_reg[11]/NET0131 ,
		\u13_ints_r_reg[6]/NET0131 ,
		_w6512_
	);
	LUT4 #(
		.INIT('h135f)
	) name4366 (
		\u13_intm_r_reg[5]/NET0131 ,
		\u13_intm_r_reg[8]/NET0131 ,
		\u13_ints_r_reg[5]/NET0131 ,
		\u13_ints_r_reg[8]/NET0131 ,
		_w6513_
	);
	LUT4 #(
		.INIT('h8000)
	) name4367 (
		_w6512_,
		_w6513_,
		_w6510_,
		_w6511_,
		_w6514_
	);
	LUT4 #(
		.INIT('h7fff)
	) name4368 (
		_w6509_,
		_w6514_,
		_w6500_,
		_w6505_,
		_w6515_
	);
	LUT4 #(
		.INIT('h4000)
	) name4369 (
		\u12_we2_reg/P0001 ,
		_w4165_,
		_w4173_,
		_w6422_,
		_w6516_
	);
	LUT4 #(
		.INIT('h4c5f)
	) name4370 (
		\u12_re1_reg/P0001 ,
		\u12_we2_reg/P0001 ,
		_w2399_,
		_w6422_,
		_w6517_
	);
	LUT2 #(
		.INIT('h4)
	) name4371 (
		wb_ack_o_pad,
		wb_cyc_i_pad,
		_w6518_
	);
	LUT2 #(
		.INIT('h4)
	) name4372 (
		_w6517_,
		_w6518_,
		_w6519_
	);
	LUT4 #(
		.INIT('h9c63)
	) name4373 (
		\u8_rp_reg[1]/NET0131 ,
		\u8_rp_reg[2]/NET0131 ,
		\u8_wp_reg[0]/P0001 ,
		\u8_wp_reg[1]/NET0131 ,
		_w6520_
	);
	LUT4 #(
		.INIT('h9c63)
	) name4374 (
		\u3_rp_reg[1]/NET0131 ,
		\u3_rp_reg[2]/NET0131 ,
		\u3_wp_reg[0]/P0001 ,
		\u3_wp_reg[1]/NET0131 ,
		_w6521_
	);
	LUT4 #(
		.INIT('h9c63)
	) name4375 (
		\u4_rp_reg[1]/NET0131 ,
		\u4_rp_reg[2]/NET0131 ,
		\u4_wp_reg[0]/P0001 ,
		\u4_wp_reg[1]/NET0131 ,
		_w6522_
	);
	LUT4 #(
		.INIT('h9c63)
	) name4376 (
		\u5_rp_reg[1]/NET0131 ,
		\u5_rp_reg[2]/NET0131 ,
		\u5_wp_reg[0]/P0001 ,
		\u5_wp_reg[1]/NET0131 ,
		_w6523_
	);
	LUT4 #(
		.INIT('h9c63)
	) name4377 (
		\u6_rp_reg[1]/NET0131 ,
		\u6_rp_reg[2]/NET0131 ,
		\u6_wp_reg[0]/P0001 ,
		\u6_wp_reg[1]/NET0131 ,
		_w6524_
	);
	LUT4 #(
		.INIT('h9c63)
	) name4378 (
		\u7_rp_reg[1]/NET0131 ,
		\u7_rp_reg[2]/NET0131 ,
		\u7_wp_reg[0]/P0001 ,
		\u7_wp_reg[1]/NET0131 ,
		_w6525_
	);
	LUT3 #(
		.INIT('h40)
	) name4379 (
		\u12_we2_reg/P0001 ,
		_w2401_,
		_w6422_,
		_w6526_
	);
	LUT2 #(
		.INIT('h8)
	) name4380 (
		\u2_ld_reg/P0001 ,
		\u8_dout_reg[0]/P0001 ,
		_w6527_
	);
	LUT4 #(
		.INIT('hc639)
	) name4381 (
		\u11_rp_reg[0]/P0001 ,
		\u11_rp_reg[1]/P0001 ,
		\u11_wp_reg[1]/P0001 ,
		\u11_wp_reg[2]/P0001 ,
		_w6528_
	);
	LUT4 #(
		.INIT('hc639)
	) name4382 (
		\u9_rp_reg[0]/P0001 ,
		\u9_rp_reg[1]/P0001 ,
		\u9_wp_reg[1]/P0001 ,
		\u9_wp_reg[2]/P0001 ,
		_w6529_
	);
	LUT4 #(
		.INIT('hc639)
	) name4383 (
		\u10_rp_reg[0]/P0001 ,
		\u10_rp_reg[1]/P0001 ,
		\u10_wp_reg[1]/P0001 ,
		\u10_wp_reg[2]/P0001 ,
		_w6530_
	);
	LUT2 #(
		.INIT('h1)
	) name4384 (
		\u13_ints_r_reg[0]/NET0131 ,
		\u15_crac_rd_done_reg/P0001 ,
		_w6531_
	);
	LUT2 #(
		.INIT('h1)
	) name4385 (
		_w2403_,
		_w6531_,
		_w6532_
	);
	LUT2 #(
		.INIT('h1)
	) name4386 (
		\u13_ints_r_reg[10]/NET0131 ,
		\u19_int_set_reg[2]/NET0131 ,
		_w6533_
	);
	LUT2 #(
		.INIT('h1)
	) name4387 (
		_w2403_,
		_w6533_,
		_w6534_
	);
	LUT2 #(
		.INIT('h1)
	) name4388 (
		\u13_ints_r_reg[12]/NET0131 ,
		\u20_int_set_reg[1]/NET0131 ,
		_w6535_
	);
	LUT2 #(
		.INIT('h1)
	) name4389 (
		_w2403_,
		_w6535_,
		_w6536_
	);
	LUT2 #(
		.INIT('h1)
	) name4390 (
		\u13_ints_r_reg[13]/NET0131 ,
		\u20_int_set_reg[2]/NET0131 ,
		_w6537_
	);
	LUT2 #(
		.INIT('h1)
	) name4391 (
		_w2403_,
		_w6537_,
		_w6538_
	);
	LUT2 #(
		.INIT('h1)
	) name4392 (
		\u13_ints_r_reg[15]/NET0131 ,
		\u21_int_set_reg[1]/NET0131 ,
		_w6539_
	);
	LUT2 #(
		.INIT('h1)
	) name4393 (
		_w2403_,
		_w6539_,
		_w6540_
	);
	LUT2 #(
		.INIT('h1)
	) name4394 (
		\u13_ints_r_reg[16]/NET0131 ,
		\u21_int_set_reg[2]/NET0131 ,
		_w6541_
	);
	LUT2 #(
		.INIT('h1)
	) name4395 (
		_w2403_,
		_w6541_,
		_w6542_
	);
	LUT2 #(
		.INIT('h1)
	) name4396 (
		\u13_ints_r_reg[18]/NET0131 ,
		\u22_int_set_reg[1]/NET0131 ,
		_w6543_
	);
	LUT2 #(
		.INIT('h1)
	) name4397 (
		_w2403_,
		_w6543_,
		_w6544_
	);
	LUT2 #(
		.INIT('h1)
	) name4398 (
		\u13_ints_r_reg[19]/NET0131 ,
		\u22_int_set_reg[2]/NET0131 ,
		_w6545_
	);
	LUT2 #(
		.INIT('h1)
	) name4399 (
		_w2403_,
		_w6545_,
		_w6546_
	);
	LUT2 #(
		.INIT('h1)
	) name4400 (
		\u13_ints_r_reg[21]/NET0131 ,
		\u23_int_set_reg[1]/NET0131 ,
		_w6547_
	);
	LUT2 #(
		.INIT('h1)
	) name4401 (
		_w2403_,
		_w6547_,
		_w6548_
	);
	LUT2 #(
		.INIT('h1)
	) name4402 (
		\u13_ints_r_reg[22]/NET0131 ,
		\u23_int_set_reg[2]/NET0131 ,
		_w6549_
	);
	LUT2 #(
		.INIT('h1)
	) name4403 (
		_w2403_,
		_w6549_,
		_w6550_
	);
	LUT2 #(
		.INIT('h1)
	) name4404 (
		\u13_ints_r_reg[24]/NET0131 ,
		\u24_int_set_reg[1]/NET0131 ,
		_w6551_
	);
	LUT2 #(
		.INIT('h1)
	) name4405 (
		_w2403_,
		_w6551_,
		_w6552_
	);
	LUT2 #(
		.INIT('h1)
	) name4406 (
		\u13_ints_r_reg[25]/NET0131 ,
		\u24_int_set_reg[2]/NET0131 ,
		_w6553_
	);
	LUT2 #(
		.INIT('h1)
	) name4407 (
		_w2403_,
		_w6553_,
		_w6554_
	);
	LUT2 #(
		.INIT('h1)
	) name4408 (
		\u13_ints_r_reg[27]/NET0131 ,
		\u25_int_set_reg[1]/NET0131 ,
		_w6555_
	);
	LUT2 #(
		.INIT('h1)
	) name4409 (
		_w2403_,
		_w6555_,
		_w6556_
	);
	LUT2 #(
		.INIT('h1)
	) name4410 (
		\u13_ints_r_reg[28]/NET0131 ,
		\u25_int_set_reg[2]/NET0131 ,
		_w6557_
	);
	LUT2 #(
		.INIT('h1)
	) name4411 (
		_w2403_,
		_w6557_,
		_w6558_
	);
	LUT2 #(
		.INIT('h1)
	) name4412 (
		\u13_ints_r_reg[3]/NET0131 ,
		\u17_int_set_reg[1]/NET0131 ,
		_w6559_
	);
	LUT2 #(
		.INIT('h1)
	) name4413 (
		_w2403_,
		_w6559_,
		_w6560_
	);
	LUT2 #(
		.INIT('h1)
	) name4414 (
		\u13_ints_r_reg[4]/NET0131 ,
		\u17_int_set_reg[2]/NET0131 ,
		_w6561_
	);
	LUT2 #(
		.INIT('h1)
	) name4415 (
		_w2403_,
		_w6561_,
		_w6562_
	);
	LUT2 #(
		.INIT('h1)
	) name4416 (
		\u13_ints_r_reg[6]/NET0131 ,
		\u18_int_set_reg[1]/NET0131 ,
		_w6563_
	);
	LUT2 #(
		.INIT('h1)
	) name4417 (
		_w2403_,
		_w6563_,
		_w6564_
	);
	LUT2 #(
		.INIT('h1)
	) name4418 (
		\u13_ints_r_reg[7]/NET0131 ,
		\u18_int_set_reg[2]/NET0131 ,
		_w6565_
	);
	LUT2 #(
		.INIT('h1)
	) name4419 (
		_w2403_,
		_w6565_,
		_w6566_
	);
	LUT2 #(
		.INIT('h1)
	) name4420 (
		\u13_ints_r_reg[9]/NET0131 ,
		\u19_int_set_reg[1]/NET0131 ,
		_w6567_
	);
	LUT2 #(
		.INIT('h1)
	) name4421 (
		_w2403_,
		_w6567_,
		_w6568_
	);
	LUT2 #(
		.INIT('h9)
	) name4422 (
		\u9_rp_reg[0]/P0001 ,
		\u9_wp_reg[1]/P0001 ,
		_w6569_
	);
	LUT4 #(
		.INIT('h8421)
	) name4423 (
		\u9_rp_reg[0]/P0001 ,
		\u9_rp_reg[1]/P0001 ,
		\u9_wp_reg[1]/P0001 ,
		\u9_wp_reg[2]/P0001 ,
		_w6570_
	);
	LUT2 #(
		.INIT('h6)
	) name4424 (
		\u9_rp_reg[2]/P0001 ,
		\u9_wp_reg[3]/P0001 ,
		_w6571_
	);
	LUT3 #(
		.INIT('h20)
	) name4425 (
		_w2688_,
		_w6571_,
		_w6570_,
		_w6572_
	);
	LUT3 #(
		.INIT('h01)
	) name4426 (
		\wb_addr_i[29]_pad ,
		\wb_addr_i[30]_pad ,
		\wb_addr_i[31]_pad ,
		_w6573_
	);
	LUT4 #(
		.INIT('hd000)
	) name4427 (
		\u12_we1_reg/P0001 ,
		\u12_we2_reg/P0001 ,
		_w6421_,
		_w6573_,
		_w6574_
	);
	LUT4 #(
		.INIT('h0200)
	) name4428 (
		\u2_cnt_reg[0]/NET0131 ,
		\u2_cnt_reg[1]/NET0131 ,
		\u2_cnt_reg[4]/NET0131 ,
		\u2_cnt_reg[6]/NET0131 ,
		_w6575_
	);
	LUT4 #(
		.INIT('h0010)
	) name4429 (
		\u2_cnt_reg[2]/NET0131 ,
		\u2_cnt_reg[3]/NET0131 ,
		\u2_cnt_reg[5]/NET0131 ,
		\u2_cnt_reg[7]/NET0131 ,
		_w6576_
	);
	LUT2 #(
		.INIT('h8)
	) name4430 (
		_w6575_,
		_w6576_,
		_w6577_
	);
	LUT2 #(
		.INIT('h9)
	) name4431 (
		\u10_rp_reg[0]/P0001 ,
		\u10_wp_reg[1]/P0001 ,
		_w6578_
	);
	LUT4 #(
		.INIT('h8421)
	) name4432 (
		\u10_rp_reg[0]/P0001 ,
		\u10_rp_reg[1]/P0001 ,
		\u10_wp_reg[1]/P0001 ,
		\u10_wp_reg[2]/P0001 ,
		_w6579_
	);
	LUT2 #(
		.INIT('h6)
	) name4433 (
		\u10_rp_reg[2]/P0001 ,
		\u10_wp_reg[3]/P0001 ,
		_w6580_
	);
	LUT3 #(
		.INIT('h20)
	) name4434 (
		_w2794_,
		_w6580_,
		_w6579_,
		_w6581_
	);
	LUT2 #(
		.INIT('h9)
	) name4435 (
		\u11_rp_reg[0]/P0001 ,
		\u11_wp_reg[1]/P0001 ,
		_w6582_
	);
	LUT4 #(
		.INIT('h8421)
	) name4436 (
		\u11_rp_reg[0]/P0001 ,
		\u11_rp_reg[1]/P0001 ,
		\u11_wp_reg[1]/P0001 ,
		\u11_wp_reg[2]/P0001 ,
		_w6583_
	);
	LUT2 #(
		.INIT('h6)
	) name4437 (
		\u11_rp_reg[2]/P0001 ,
		\u11_wp_reg[3]/P0001 ,
		_w6584_
	);
	LUT3 #(
		.INIT('h20)
	) name4438 (
		_w2567_,
		_w6584_,
		_w6583_,
		_w6585_
	);
	LUT4 #(
		.INIT('hbefa)
	) name4439 (
		suspended_o_pad,
		\u2_cnt_reg[4]/NET0131 ,
		\u2_cnt_reg[5]/NET0131 ,
		_w4320_,
		_w6586_
	);
	LUT4 #(
		.INIT('h78f0)
	) name4440 (
		\u2_cnt_reg[4]/NET0131 ,
		\u2_cnt_reg[5]/NET0131 ,
		\u2_cnt_reg[6]/NET0131 ,
		_w4320_,
		_w6587_
	);
	LUT2 #(
		.INIT('he)
	) name4441 (
		suspended_o_pad,
		_w6587_,
		_w6588_
	);
	LUT2 #(
		.INIT('h1)
	) name4442 (
		\u2_cnt_reg[4]/NET0131 ,
		\u2_cnt_reg[5]/NET0131 ,
		_w6589_
	);
	LUT3 #(
		.INIT('h01)
	) name4443 (
		\u2_cnt_reg[4]/NET0131 ,
		\u2_cnt_reg[5]/NET0131 ,
		\u2_cnt_reg[6]/NET0131 ,
		_w6590_
	);
	LUT4 #(
		.INIT('h0200)
	) name4444 (
		\u2_cnt_reg[0]/NET0131 ,
		\u2_cnt_reg[1]/NET0131 ,
		\u2_cnt_reg[2]/NET0131 ,
		\u2_cnt_reg[3]/NET0131 ,
		_w6591_
	);
	LUT3 #(
		.INIT('h80)
	) name4445 (
		\u2_cnt_reg[7]/NET0131 ,
		_w6591_,
		_w6590_,
		_w6592_
	);
	LUT2 #(
		.INIT('h1)
	) name4446 (
		\u2_cnt_reg[6]/NET0131 ,
		\u2_cnt_reg[7]/NET0131 ,
		_w6593_
	);
	LUT4 #(
		.INIT('h0001)
	) name4447 (
		\u2_cnt_reg[4]/NET0131 ,
		\u2_cnt_reg[5]/NET0131 ,
		\u2_cnt_reg[6]/NET0131 ,
		\u2_cnt_reg[7]/NET0131 ,
		_w6594_
	);
	LUT4 #(
		.INIT('h0100)
	) name4448 (
		\u2_to_cnt_reg[2]/NET0131 ,
		\u2_to_cnt_reg[3]/NET0131 ,
		\u2_to_cnt_reg[4]/NET0131 ,
		\u2_to_cnt_reg[5]/NET0131 ,
		_w6595_
	);
	LUT2 #(
		.INIT('h2)
	) name4449 (
		\u2_to_cnt_reg[0]/NET0131 ,
		\u2_to_cnt_reg[1]/NET0131 ,
		_w6596_
	);
	LUT2 #(
		.INIT('h8)
	) name4450 (
		_w6595_,
		_w6596_,
		_w6597_
	);
	LUT4 #(
		.INIT('h1511)
	) name4451 (
		\u2_bit_clk_e_reg/P0001 ,
		\u2_to_cnt_reg[0]/NET0131 ,
		\u2_to_cnt_reg[1]/NET0131 ,
		_w6595_,
		_w6598_
	);
	LUT4 #(
		.INIT('h1014)
	) name4452 (
		\u2_bit_clk_e_reg/P0001 ,
		\u2_to_cnt_reg[0]/NET0131 ,
		\u2_to_cnt_reg[1]/NET0131 ,
		_w6595_,
		_w6599_
	);
	LUT2 #(
		.INIT('h8)
	) name4453 (
		_w6580_,
		_w6579_,
		_w6600_
	);
	LUT2 #(
		.INIT('h8)
	) name4454 (
		_w6584_,
		_w6583_,
		_w6601_
	);
	LUT4 #(
		.INIT('h0008)
	) name4455 (
		\u2_cnt_reg[2]/NET0131 ,
		\u2_cnt_reg[3]/NET0131 ,
		\u2_cnt_reg[5]/NET0131 ,
		\u2_cnt_reg[7]/NET0131 ,
		_w6602_
	);
	LUT2 #(
		.INIT('h8)
	) name4456 (
		_w6575_,
		_w6602_,
		_w6603_
	);
	LUT2 #(
		.INIT('h8)
	) name4457 (
		_w6571_,
		_w6570_,
		_w6604_
	);
	LUT3 #(
		.INIT('h01)
	) name4458 (
		\u2_cnt_reg[1]/NET0131 ,
		\u2_cnt_reg[2]/NET0131 ,
		\u2_cnt_reg[3]/NET0131 ,
		_w6605_
	);
	LUT4 #(
		.INIT('h0001)
	) name4459 (
		\u2_cnt_reg[1]/NET0131 ,
		\u2_cnt_reg[2]/NET0131 ,
		\u2_cnt_reg[3]/NET0131 ,
		\u2_cnt_reg[4]/NET0131 ,
		_w6606_
	);
	LUT3 #(
		.INIT('hae)
	) name4460 (
		\u2_cnt_reg[7]/NET0131 ,
		_w4321_,
		_w6606_,
		_w6607_
	);
	LUT4 #(
		.INIT('h2000)
	) name4461 (
		\u12_re1_reg/P0001 ,
		\wb_addr_i[2]_pad ,
		_w2399_,
		_w4166_,
		_w6608_
	);
	LUT4 #(
		.INIT('h8000)
	) name4462 (
		\u12_re1_reg/P0001 ,
		\wb_addr_i[2]_pad ,
		_w2399_,
		_w4166_,
		_w6609_
	);
	LUT3 #(
		.INIT('he0)
	) name4463 (
		\u2_cnt_reg[1]/NET0131 ,
		\u2_cnt_reg[2]/NET0131 ,
		\u2_cnt_reg[3]/NET0131 ,
		_w6610_
	);
	LUT2 #(
		.INIT('h8)
	) name4464 (
		\u2_cnt_reg[4]/NET0131 ,
		\u2_cnt_reg[5]/NET0131 ,
		_w6611_
	);
	LUT3 #(
		.INIT('hd5)
	) name4465 (
		_w6593_,
		_w6610_,
		_w6611_,
		_w6612_
	);
	LUT2 #(
		.INIT('hb)
	) name4466 (
		suspended_o_pad,
		\u2_cnt_reg[0]/NET0131 ,
		_w6613_
	);
	LUT3 #(
		.INIT('hbe)
	) name4467 (
		suspended_o_pad,
		\u2_cnt_reg[0]/NET0131 ,
		\u2_cnt_reg[1]/NET0131 ,
		_w6614_
	);
	LUT4 #(
		.INIT('hbfea)
	) name4468 (
		suspended_o_pad,
		\u2_cnt_reg[0]/NET0131 ,
		\u2_cnt_reg[1]/NET0131 ,
		\u2_cnt_reg[2]/NET0131 ,
		_w6615_
	);
	LUT3 #(
		.INIT('ha2)
	) name4469 (
		\u2_cnt_reg[7]/NET0131 ,
		_w6590_,
		_w6610_,
		_w6616_
	);
	LUT3 #(
		.INIT('h40)
	) name4470 (
		\u2_cnt_reg[0]/NET0131 ,
		_w6594_,
		_w6605_,
		_w6617_
	);
	LUT4 #(
		.INIT('h0800)
	) name4471 (
		\u2_cnt_reg[0]/NET0131 ,
		\u2_cnt_reg[2]/NET0131 ,
		\u2_cnt_reg[4]/NET0131 ,
		\u2_cnt_reg[5]/NET0131 ,
		_w6618_
	);
	LUT4 #(
		.INIT('h0001)
	) name4472 (
		\u2_cnt_reg[1]/NET0131 ,
		\u2_cnt_reg[3]/NET0131 ,
		\u2_cnt_reg[6]/NET0131 ,
		\u2_cnt_reg[7]/NET0131 ,
		_w6619_
	);
	LUT2 #(
		.INIT('h8)
	) name4473 (
		_w6618_,
		_w6619_,
		_w6620_
	);
	LUT4 #(
		.INIT('h8000)
	) name4474 (
		\u12_re1_reg/P0001 ,
		_w2399_,
		_w4167_,
		_w4168_,
		_w6621_
	);
	LUT3 #(
		.INIT('h80)
	) name4475 (
		\u2_cnt_reg[1]/NET0131 ,
		\u2_cnt_reg[2]/NET0131 ,
		\u2_cnt_reg[3]/NET0131 ,
		_w6622_
	);
	LUT4 #(
		.INIT('heece)
	) name4476 (
		\u2_cnt_reg[6]/NET0131 ,
		\u2_cnt_reg[7]/NET0131 ,
		_w6589_,
		_w6622_,
		_w6623_
	);
	LUT3 #(
		.INIT('h02)
	) name4477 (
		\u2_cnt_reg[4]/NET0131 ,
		\u2_cnt_reg[6]/NET0131 ,
		\u2_cnt_reg[7]/NET0131 ,
		_w6624_
	);
	LUT3 #(
		.INIT('h80)
	) name4478 (
		\u2_cnt_reg[5]/NET0131 ,
		_w6591_,
		_w6624_,
		_w6625_
	);
	LUT4 #(
		.INIT('hff35)
	) name4479 (
		\u9_mem_reg[0][0]/P0001 ,
		\u9_mem_reg[1][0]/P0001 ,
		\u9_rp_reg[0]/P0001 ,
		\u9_rp_reg[1]/P0001 ,
		_w6626_
	);
	LUT4 #(
		.INIT('h35ff)
	) name4480 (
		\u9_mem_reg[2][0]/P0001 ,
		\u9_mem_reg[3][0]/P0001 ,
		\u9_rp_reg[0]/P0001 ,
		\u9_rp_reg[1]/P0001 ,
		_w6627_
	);
	LUT2 #(
		.INIT('h7)
	) name4481 (
		_w6626_,
		_w6627_,
		_w6628_
	);
	LUT4 #(
		.INIT('hf3f5)
	) name4482 (
		\u9_mem_reg[0][10]/P0001 ,
		\u9_mem_reg[2][10]/P0001 ,
		\u9_rp_reg[0]/P0001 ,
		\u9_rp_reg[1]/P0001 ,
		_w6629_
	);
	LUT4 #(
		.INIT('h3f5f)
	) name4483 (
		\u9_mem_reg[1][10]/P0001 ,
		\u9_mem_reg[3][10]/P0001 ,
		\u9_rp_reg[0]/P0001 ,
		\u9_rp_reg[1]/P0001 ,
		_w6630_
	);
	LUT2 #(
		.INIT('h7)
	) name4484 (
		_w6629_,
		_w6630_,
		_w6631_
	);
	LUT4 #(
		.INIT('hff35)
	) name4485 (
		\u9_mem_reg[0][11]/P0001 ,
		\u9_mem_reg[1][11]/P0001 ,
		\u9_rp_reg[0]/P0001 ,
		\u9_rp_reg[1]/P0001 ,
		_w6632_
	);
	LUT4 #(
		.INIT('h35ff)
	) name4486 (
		\u9_mem_reg[2][11]/P0001 ,
		\u9_mem_reg[3][11]/P0001 ,
		\u9_rp_reg[0]/P0001 ,
		\u9_rp_reg[1]/P0001 ,
		_w6633_
	);
	LUT2 #(
		.INIT('h7)
	) name4487 (
		_w6632_,
		_w6633_,
		_w6634_
	);
	LUT4 #(
		.INIT('hff35)
	) name4488 (
		\u9_mem_reg[0][12]/P0001 ,
		\u9_mem_reg[1][12]/P0001 ,
		\u9_rp_reg[0]/P0001 ,
		\u9_rp_reg[1]/P0001 ,
		_w6635_
	);
	LUT4 #(
		.INIT('h35ff)
	) name4489 (
		\u9_mem_reg[2][12]/P0001 ,
		\u9_mem_reg[3][12]/P0001 ,
		\u9_rp_reg[0]/P0001 ,
		\u9_rp_reg[1]/P0001 ,
		_w6636_
	);
	LUT2 #(
		.INIT('h7)
	) name4490 (
		_w6635_,
		_w6636_,
		_w6637_
	);
	LUT4 #(
		.INIT('hff35)
	) name4491 (
		\u9_mem_reg[0][13]/P0001 ,
		\u9_mem_reg[1][13]/P0001 ,
		\u9_rp_reg[0]/P0001 ,
		\u9_rp_reg[1]/P0001 ,
		_w6638_
	);
	LUT4 #(
		.INIT('h35ff)
	) name4492 (
		\u9_mem_reg[2][13]/P0001 ,
		\u9_mem_reg[3][13]/P0001 ,
		\u9_rp_reg[0]/P0001 ,
		\u9_rp_reg[1]/P0001 ,
		_w6639_
	);
	LUT2 #(
		.INIT('h7)
	) name4493 (
		_w6638_,
		_w6639_,
		_w6640_
	);
	LUT4 #(
		.INIT('hff35)
	) name4494 (
		\u9_mem_reg[0][14]/P0001 ,
		\u9_mem_reg[1][14]/P0001 ,
		\u9_rp_reg[0]/P0001 ,
		\u9_rp_reg[1]/P0001 ,
		_w6641_
	);
	LUT4 #(
		.INIT('h35ff)
	) name4495 (
		\u9_mem_reg[2][14]/P0001 ,
		\u9_mem_reg[3][14]/P0001 ,
		\u9_rp_reg[0]/P0001 ,
		\u9_rp_reg[1]/P0001 ,
		_w6642_
	);
	LUT2 #(
		.INIT('h7)
	) name4496 (
		_w6641_,
		_w6642_,
		_w6643_
	);
	LUT4 #(
		.INIT('hff35)
	) name4497 (
		\u9_mem_reg[0][15]/P0001 ,
		\u9_mem_reg[1][15]/P0001 ,
		\u9_rp_reg[0]/P0001 ,
		\u9_rp_reg[1]/P0001 ,
		_w6644_
	);
	LUT4 #(
		.INIT('h35ff)
	) name4498 (
		\u9_mem_reg[2][15]/P0001 ,
		\u9_mem_reg[3][15]/P0001 ,
		\u9_rp_reg[0]/P0001 ,
		\u9_rp_reg[1]/P0001 ,
		_w6645_
	);
	LUT2 #(
		.INIT('h7)
	) name4499 (
		_w6644_,
		_w6645_,
		_w6646_
	);
	LUT4 #(
		.INIT('hf35f)
	) name4500 (
		\u9_mem_reg[1][16]/P0001 ,
		\u9_mem_reg[2][16]/P0001 ,
		\u9_rp_reg[0]/P0001 ,
		\u9_rp_reg[1]/P0001 ,
		_w6647_
	);
	LUT4 #(
		.INIT('h3ff5)
	) name4501 (
		\u9_mem_reg[0][16]/P0001 ,
		\u9_mem_reg[3][16]/P0001 ,
		\u9_rp_reg[0]/P0001 ,
		\u9_rp_reg[1]/P0001 ,
		_w6648_
	);
	LUT2 #(
		.INIT('h7)
	) name4502 (
		_w6647_,
		_w6648_,
		_w6649_
	);
	LUT4 #(
		.INIT('hff35)
	) name4503 (
		\u9_mem_reg[0][17]/P0001 ,
		\u9_mem_reg[1][17]/P0001 ,
		\u9_rp_reg[0]/P0001 ,
		\u9_rp_reg[1]/P0001 ,
		_w6650_
	);
	LUT4 #(
		.INIT('h35ff)
	) name4504 (
		\u9_mem_reg[2][17]/P0001 ,
		\u9_mem_reg[3][17]/P0001 ,
		\u9_rp_reg[0]/P0001 ,
		\u9_rp_reg[1]/P0001 ,
		_w6651_
	);
	LUT2 #(
		.INIT('h7)
	) name4505 (
		_w6650_,
		_w6651_,
		_w6652_
	);
	LUT4 #(
		.INIT('hf35f)
	) name4506 (
		\u9_mem_reg[1][18]/P0001 ,
		\u9_mem_reg[2][18]/P0001 ,
		\u9_rp_reg[0]/P0001 ,
		\u9_rp_reg[1]/P0001 ,
		_w6653_
	);
	LUT4 #(
		.INIT('h3ff5)
	) name4507 (
		\u9_mem_reg[0][18]/P0001 ,
		\u9_mem_reg[3][18]/P0001 ,
		\u9_rp_reg[0]/P0001 ,
		\u9_rp_reg[1]/P0001 ,
		_w6654_
	);
	LUT2 #(
		.INIT('h7)
	) name4508 (
		_w6653_,
		_w6654_,
		_w6655_
	);
	LUT4 #(
		.INIT('hf35f)
	) name4509 (
		\u9_mem_reg[1][19]/P0001 ,
		\u9_mem_reg[2][19]/P0001 ,
		\u9_rp_reg[0]/P0001 ,
		\u9_rp_reg[1]/P0001 ,
		_w6656_
	);
	LUT4 #(
		.INIT('h3ff5)
	) name4510 (
		\u9_mem_reg[0][19]/P0001 ,
		\u9_mem_reg[3][19]/P0001 ,
		\u9_rp_reg[0]/P0001 ,
		\u9_rp_reg[1]/P0001 ,
		_w6657_
	);
	LUT2 #(
		.INIT('h7)
	) name4511 (
		_w6656_,
		_w6657_,
		_w6658_
	);
	LUT4 #(
		.INIT('hff35)
	) name4512 (
		\u9_mem_reg[0][1]/P0001 ,
		\u9_mem_reg[1][1]/P0001 ,
		\u9_rp_reg[0]/P0001 ,
		\u9_rp_reg[1]/P0001 ,
		_w6659_
	);
	LUT4 #(
		.INIT('h35ff)
	) name4513 (
		\u9_mem_reg[2][1]/P0001 ,
		\u9_mem_reg[3][1]/P0001 ,
		\u9_rp_reg[0]/P0001 ,
		\u9_rp_reg[1]/P0001 ,
		_w6660_
	);
	LUT2 #(
		.INIT('h7)
	) name4514 (
		_w6659_,
		_w6660_,
		_w6661_
	);
	LUT4 #(
		.INIT('hf3f5)
	) name4515 (
		\u9_mem_reg[0][20]/P0001 ,
		\u9_mem_reg[2][20]/P0001 ,
		\u9_rp_reg[0]/P0001 ,
		\u9_rp_reg[1]/P0001 ,
		_w6662_
	);
	LUT4 #(
		.INIT('h3f5f)
	) name4516 (
		\u9_mem_reg[1][20]/P0001 ,
		\u9_mem_reg[3][20]/P0001 ,
		\u9_rp_reg[0]/P0001 ,
		\u9_rp_reg[1]/P0001 ,
		_w6663_
	);
	LUT2 #(
		.INIT('h7)
	) name4517 (
		_w6662_,
		_w6663_,
		_w6664_
	);
	LUT4 #(
		.INIT('hf35f)
	) name4518 (
		\u9_mem_reg[1][21]/P0001 ,
		\u9_mem_reg[2][21]/P0001 ,
		\u9_rp_reg[0]/P0001 ,
		\u9_rp_reg[1]/P0001 ,
		_w6665_
	);
	LUT4 #(
		.INIT('h3ff5)
	) name4519 (
		\u9_mem_reg[0][21]/P0001 ,
		\u9_mem_reg[3][21]/P0001 ,
		\u9_rp_reg[0]/P0001 ,
		\u9_rp_reg[1]/P0001 ,
		_w6666_
	);
	LUT2 #(
		.INIT('h7)
	) name4520 (
		_w6665_,
		_w6666_,
		_w6667_
	);
	LUT4 #(
		.INIT('hf35f)
	) name4521 (
		\u9_mem_reg[1][22]/P0001 ,
		\u9_mem_reg[2][22]/P0001 ,
		\u9_rp_reg[0]/P0001 ,
		\u9_rp_reg[1]/P0001 ,
		_w6668_
	);
	LUT4 #(
		.INIT('h3ff5)
	) name4522 (
		\u9_mem_reg[0][22]/P0001 ,
		\u9_mem_reg[3][22]/P0001 ,
		\u9_rp_reg[0]/P0001 ,
		\u9_rp_reg[1]/P0001 ,
		_w6669_
	);
	LUT2 #(
		.INIT('h7)
	) name4523 (
		_w6668_,
		_w6669_,
		_w6670_
	);
	LUT4 #(
		.INIT('hf35f)
	) name4524 (
		\u9_mem_reg[1][23]/P0001 ,
		\u9_mem_reg[2][23]/P0001 ,
		\u9_rp_reg[0]/P0001 ,
		\u9_rp_reg[1]/P0001 ,
		_w6671_
	);
	LUT4 #(
		.INIT('h3ff5)
	) name4525 (
		\u9_mem_reg[0][23]/P0001 ,
		\u9_mem_reg[3][23]/P0001 ,
		\u9_rp_reg[0]/P0001 ,
		\u9_rp_reg[1]/P0001 ,
		_w6672_
	);
	LUT2 #(
		.INIT('h7)
	) name4526 (
		_w6671_,
		_w6672_,
		_w6673_
	);
	LUT4 #(
		.INIT('hf35f)
	) name4527 (
		\u9_mem_reg[1][24]/P0001 ,
		\u9_mem_reg[2][24]/P0001 ,
		\u9_rp_reg[0]/P0001 ,
		\u9_rp_reg[1]/P0001 ,
		_w6674_
	);
	LUT4 #(
		.INIT('h3ff5)
	) name4528 (
		\u9_mem_reg[0][24]/P0001 ,
		\u9_mem_reg[3][24]/P0001 ,
		\u9_rp_reg[0]/P0001 ,
		\u9_rp_reg[1]/P0001 ,
		_w6675_
	);
	LUT2 #(
		.INIT('h7)
	) name4529 (
		_w6674_,
		_w6675_,
		_w6676_
	);
	LUT4 #(
		.INIT('hf35f)
	) name4530 (
		\u9_mem_reg[1][26]/P0001 ,
		\u9_mem_reg[2][26]/P0001 ,
		\u9_rp_reg[0]/P0001 ,
		\u9_rp_reg[1]/P0001 ,
		_w6677_
	);
	LUT4 #(
		.INIT('h3ff5)
	) name4531 (
		\u9_mem_reg[0][26]/P0001 ,
		\u9_mem_reg[3][26]/P0001 ,
		\u9_rp_reg[0]/P0001 ,
		\u9_rp_reg[1]/P0001 ,
		_w6678_
	);
	LUT2 #(
		.INIT('h7)
	) name4532 (
		_w6677_,
		_w6678_,
		_w6679_
	);
	LUT4 #(
		.INIT('hf35f)
	) name4533 (
		\u9_mem_reg[1][27]/P0001 ,
		\u9_mem_reg[2][27]/P0001 ,
		\u9_rp_reg[0]/P0001 ,
		\u9_rp_reg[1]/P0001 ,
		_w6680_
	);
	LUT4 #(
		.INIT('h3ff5)
	) name4534 (
		\u9_mem_reg[0][27]/P0001 ,
		\u9_mem_reg[3][27]/P0001 ,
		\u9_rp_reg[0]/P0001 ,
		\u9_rp_reg[1]/P0001 ,
		_w6681_
	);
	LUT2 #(
		.INIT('h7)
	) name4535 (
		_w6680_,
		_w6681_,
		_w6682_
	);
	LUT4 #(
		.INIT('hf35f)
	) name4536 (
		\u9_mem_reg[1][28]/P0001 ,
		\u9_mem_reg[2][28]/P0001 ,
		\u9_rp_reg[0]/P0001 ,
		\u9_rp_reg[1]/P0001 ,
		_w6683_
	);
	LUT4 #(
		.INIT('h3ff5)
	) name4537 (
		\u9_mem_reg[0][28]/P0001 ,
		\u9_mem_reg[3][28]/P0001 ,
		\u9_rp_reg[0]/P0001 ,
		\u9_rp_reg[1]/P0001 ,
		_w6684_
	);
	LUT2 #(
		.INIT('h7)
	) name4538 (
		_w6683_,
		_w6684_,
		_w6685_
	);
	LUT4 #(
		.INIT('hf35f)
	) name4539 (
		\u9_mem_reg[1][29]/P0001 ,
		\u9_mem_reg[2][29]/P0001 ,
		\u9_rp_reg[0]/P0001 ,
		\u9_rp_reg[1]/P0001 ,
		_w6686_
	);
	LUT4 #(
		.INIT('h3ff5)
	) name4540 (
		\u9_mem_reg[0][29]/P0001 ,
		\u9_mem_reg[3][29]/P0001 ,
		\u9_rp_reg[0]/P0001 ,
		\u9_rp_reg[1]/P0001 ,
		_w6687_
	);
	LUT2 #(
		.INIT('h7)
	) name4541 (
		_w6686_,
		_w6687_,
		_w6688_
	);
	LUT4 #(
		.INIT('hff35)
	) name4542 (
		\u9_mem_reg[0][2]/P0001 ,
		\u9_mem_reg[1][2]/P0001 ,
		\u9_rp_reg[0]/P0001 ,
		\u9_rp_reg[1]/P0001 ,
		_w6689_
	);
	LUT4 #(
		.INIT('h35ff)
	) name4543 (
		\u9_mem_reg[2][2]/P0001 ,
		\u9_mem_reg[3][2]/P0001 ,
		\u9_rp_reg[0]/P0001 ,
		\u9_rp_reg[1]/P0001 ,
		_w6690_
	);
	LUT2 #(
		.INIT('h7)
	) name4544 (
		_w6689_,
		_w6690_,
		_w6691_
	);
	LUT4 #(
		.INIT('hf35f)
	) name4545 (
		\u9_mem_reg[1][30]/P0001 ,
		\u9_mem_reg[2][30]/P0001 ,
		\u9_rp_reg[0]/P0001 ,
		\u9_rp_reg[1]/P0001 ,
		_w6692_
	);
	LUT4 #(
		.INIT('h3ff5)
	) name4546 (
		\u9_mem_reg[0][30]/P0001 ,
		\u9_mem_reg[3][30]/P0001 ,
		\u9_rp_reg[0]/P0001 ,
		\u9_rp_reg[1]/P0001 ,
		_w6693_
	);
	LUT2 #(
		.INIT('h7)
	) name4547 (
		_w6692_,
		_w6693_,
		_w6694_
	);
	LUT4 #(
		.INIT('hf35f)
	) name4548 (
		\u9_mem_reg[1][31]/P0001 ,
		\u9_mem_reg[2][31]/P0001 ,
		\u9_rp_reg[0]/P0001 ,
		\u9_rp_reg[1]/P0001 ,
		_w6695_
	);
	LUT4 #(
		.INIT('h3ff5)
	) name4549 (
		\u9_mem_reg[0][31]/P0001 ,
		\u9_mem_reg[3][31]/P0001 ,
		\u9_rp_reg[0]/P0001 ,
		\u9_rp_reg[1]/P0001 ,
		_w6696_
	);
	LUT2 #(
		.INIT('h7)
	) name4550 (
		_w6695_,
		_w6696_,
		_w6697_
	);
	LUT4 #(
		.INIT('hff35)
	) name4551 (
		\u9_mem_reg[0][3]/P0001 ,
		\u9_mem_reg[1][3]/P0001 ,
		\u9_rp_reg[0]/P0001 ,
		\u9_rp_reg[1]/P0001 ,
		_w6698_
	);
	LUT4 #(
		.INIT('h35ff)
	) name4552 (
		\u9_mem_reg[2][3]/P0001 ,
		\u9_mem_reg[3][3]/P0001 ,
		\u9_rp_reg[0]/P0001 ,
		\u9_rp_reg[1]/P0001 ,
		_w6699_
	);
	LUT2 #(
		.INIT('h7)
	) name4553 (
		_w6698_,
		_w6699_,
		_w6700_
	);
	LUT4 #(
		.INIT('hff35)
	) name4554 (
		\u9_mem_reg[0][5]/P0001 ,
		\u9_mem_reg[1][5]/P0001 ,
		\u9_rp_reg[0]/P0001 ,
		\u9_rp_reg[1]/P0001 ,
		_w6701_
	);
	LUT4 #(
		.INIT('h35ff)
	) name4555 (
		\u9_mem_reg[2][5]/P0001 ,
		\u9_mem_reg[3][5]/P0001 ,
		\u9_rp_reg[0]/P0001 ,
		\u9_rp_reg[1]/P0001 ,
		_w6702_
	);
	LUT2 #(
		.INIT('h7)
	) name4556 (
		_w6701_,
		_w6702_,
		_w6703_
	);
	LUT4 #(
		.INIT('hf35f)
	) name4557 (
		\u9_mem_reg[1][6]/P0001 ,
		\u9_mem_reg[2][6]/P0001 ,
		\u9_rp_reg[0]/P0001 ,
		\u9_rp_reg[1]/P0001 ,
		_w6704_
	);
	LUT4 #(
		.INIT('h3ff5)
	) name4558 (
		\u9_mem_reg[0][6]/P0001 ,
		\u9_mem_reg[3][6]/P0001 ,
		\u9_rp_reg[0]/P0001 ,
		\u9_rp_reg[1]/P0001 ,
		_w6705_
	);
	LUT2 #(
		.INIT('h7)
	) name4559 (
		_w6704_,
		_w6705_,
		_w6706_
	);
	LUT4 #(
		.INIT('hf3f5)
	) name4560 (
		\u9_mem_reg[0][7]/P0001 ,
		\u9_mem_reg[2][7]/P0001 ,
		\u9_rp_reg[0]/P0001 ,
		\u9_rp_reg[1]/P0001 ,
		_w6707_
	);
	LUT4 #(
		.INIT('h3f5f)
	) name4561 (
		\u9_mem_reg[1][7]/P0001 ,
		\u9_mem_reg[3][7]/P0001 ,
		\u9_rp_reg[0]/P0001 ,
		\u9_rp_reg[1]/P0001 ,
		_w6708_
	);
	LUT2 #(
		.INIT('h7)
	) name4562 (
		_w6707_,
		_w6708_,
		_w6709_
	);
	LUT4 #(
		.INIT('hf3f5)
	) name4563 (
		\u10_mem_reg[0][0]/P0001 ,
		\u10_mem_reg[2][0]/P0001 ,
		\u10_rp_reg[0]/P0001 ,
		\u10_rp_reg[1]/P0001 ,
		_w6710_
	);
	LUT4 #(
		.INIT('h3f5f)
	) name4564 (
		\u10_mem_reg[1][0]/P0001 ,
		\u10_mem_reg[3][0]/P0001 ,
		\u10_rp_reg[0]/P0001 ,
		\u10_rp_reg[1]/P0001 ,
		_w6711_
	);
	LUT2 #(
		.INIT('h7)
	) name4565 (
		_w6710_,
		_w6711_,
		_w6712_
	);
	LUT4 #(
		.INIT('hf35f)
	) name4566 (
		\u9_mem_reg[1][25]/P0001 ,
		\u9_mem_reg[2][25]/P0001 ,
		\u9_rp_reg[0]/P0001 ,
		\u9_rp_reg[1]/P0001 ,
		_w6713_
	);
	LUT4 #(
		.INIT('h3ff5)
	) name4567 (
		\u9_mem_reg[0][25]/P0001 ,
		\u9_mem_reg[3][25]/P0001 ,
		\u9_rp_reg[0]/P0001 ,
		\u9_rp_reg[1]/P0001 ,
		_w6714_
	);
	LUT2 #(
		.INIT('h7)
	) name4568 (
		_w6713_,
		_w6714_,
		_w6715_
	);
	LUT4 #(
		.INIT('hff35)
	) name4569 (
		\u10_mem_reg[0][11]/P0001 ,
		\u10_mem_reg[1][11]/P0001 ,
		\u10_rp_reg[0]/P0001 ,
		\u10_rp_reg[1]/P0001 ,
		_w6716_
	);
	LUT4 #(
		.INIT('h35ff)
	) name4570 (
		\u10_mem_reg[2][11]/P0001 ,
		\u10_mem_reg[3][11]/P0001 ,
		\u10_rp_reg[0]/P0001 ,
		\u10_rp_reg[1]/P0001 ,
		_w6717_
	);
	LUT2 #(
		.INIT('h7)
	) name4571 (
		_w6716_,
		_w6717_,
		_w6718_
	);
	LUT4 #(
		.INIT('hff35)
	) name4572 (
		\u10_mem_reg[0][12]/P0001 ,
		\u10_mem_reg[1][12]/P0001 ,
		\u10_rp_reg[0]/P0001 ,
		\u10_rp_reg[1]/P0001 ,
		_w6719_
	);
	LUT4 #(
		.INIT('h35ff)
	) name4573 (
		\u10_mem_reg[2][12]/P0001 ,
		\u10_mem_reg[3][12]/P0001 ,
		\u10_rp_reg[0]/P0001 ,
		\u10_rp_reg[1]/P0001 ,
		_w6720_
	);
	LUT2 #(
		.INIT('h7)
	) name4574 (
		_w6719_,
		_w6720_,
		_w6721_
	);
	LUT4 #(
		.INIT('hf3f5)
	) name4575 (
		\u10_mem_reg[0][13]/P0001 ,
		\u10_mem_reg[2][13]/P0001 ,
		\u10_rp_reg[0]/P0001 ,
		\u10_rp_reg[1]/P0001 ,
		_w6722_
	);
	LUT4 #(
		.INIT('h3f5f)
	) name4576 (
		\u10_mem_reg[1][13]/P0001 ,
		\u10_mem_reg[3][13]/P0001 ,
		\u10_rp_reg[0]/P0001 ,
		\u10_rp_reg[1]/P0001 ,
		_w6723_
	);
	LUT2 #(
		.INIT('h7)
	) name4577 (
		_w6722_,
		_w6723_,
		_w6724_
	);
	LUT4 #(
		.INIT('hf3f5)
	) name4578 (
		\u10_mem_reg[0][15]/P0001 ,
		\u10_mem_reg[2][15]/P0001 ,
		\u10_rp_reg[0]/P0001 ,
		\u10_rp_reg[1]/P0001 ,
		_w6725_
	);
	LUT4 #(
		.INIT('h3f5f)
	) name4579 (
		\u10_mem_reg[1][15]/P0001 ,
		\u10_mem_reg[3][15]/P0001 ,
		\u10_rp_reg[0]/P0001 ,
		\u10_rp_reg[1]/P0001 ,
		_w6726_
	);
	LUT2 #(
		.INIT('h7)
	) name4580 (
		_w6725_,
		_w6726_,
		_w6727_
	);
	LUT4 #(
		.INIT('hff35)
	) name4581 (
		\u10_mem_reg[0][16]/P0001 ,
		\u10_mem_reg[1][16]/P0001 ,
		\u10_rp_reg[0]/P0001 ,
		\u10_rp_reg[1]/P0001 ,
		_w6728_
	);
	LUT4 #(
		.INIT('h35ff)
	) name4582 (
		\u10_mem_reg[2][16]/P0001 ,
		\u10_mem_reg[3][16]/P0001 ,
		\u10_rp_reg[0]/P0001 ,
		\u10_rp_reg[1]/P0001 ,
		_w6729_
	);
	LUT2 #(
		.INIT('h7)
	) name4583 (
		_w6728_,
		_w6729_,
		_w6730_
	);
	LUT4 #(
		.INIT('hf35f)
	) name4584 (
		\u10_mem_reg[1][17]/P0001 ,
		\u10_mem_reg[2][17]/P0001 ,
		\u10_rp_reg[0]/P0001 ,
		\u10_rp_reg[1]/P0001 ,
		_w6731_
	);
	LUT4 #(
		.INIT('h3ff5)
	) name4585 (
		\u10_mem_reg[0][17]/P0001 ,
		\u10_mem_reg[3][17]/P0001 ,
		\u10_rp_reg[0]/P0001 ,
		\u10_rp_reg[1]/P0001 ,
		_w6732_
	);
	LUT2 #(
		.INIT('h7)
	) name4586 (
		_w6731_,
		_w6732_,
		_w6733_
	);
	LUT4 #(
		.INIT('hf35f)
	) name4587 (
		\u10_mem_reg[1][18]/P0001 ,
		\u10_mem_reg[2][18]/P0001 ,
		\u10_rp_reg[0]/P0001 ,
		\u10_rp_reg[1]/P0001 ,
		_w6734_
	);
	LUT4 #(
		.INIT('h3ff5)
	) name4588 (
		\u10_mem_reg[0][18]/P0001 ,
		\u10_mem_reg[3][18]/P0001 ,
		\u10_rp_reg[0]/P0001 ,
		\u10_rp_reg[1]/P0001 ,
		_w6735_
	);
	LUT2 #(
		.INIT('h7)
	) name4589 (
		_w6734_,
		_w6735_,
		_w6736_
	);
	LUT4 #(
		.INIT('hf3f5)
	) name4590 (
		\u10_mem_reg[0][19]/P0001 ,
		\u10_mem_reg[2][19]/P0001 ,
		\u10_rp_reg[0]/P0001 ,
		\u10_rp_reg[1]/P0001 ,
		_w6737_
	);
	LUT4 #(
		.INIT('h3f5f)
	) name4591 (
		\u10_mem_reg[1][19]/P0001 ,
		\u10_mem_reg[3][19]/P0001 ,
		\u10_rp_reg[0]/P0001 ,
		\u10_rp_reg[1]/P0001 ,
		_w6738_
	);
	LUT2 #(
		.INIT('h7)
	) name4592 (
		_w6737_,
		_w6738_,
		_w6739_
	);
	LUT4 #(
		.INIT('hf3f5)
	) name4593 (
		\u10_mem_reg[0][1]/P0001 ,
		\u10_mem_reg[2][1]/P0001 ,
		\u10_rp_reg[0]/P0001 ,
		\u10_rp_reg[1]/P0001 ,
		_w6740_
	);
	LUT4 #(
		.INIT('h3f5f)
	) name4594 (
		\u10_mem_reg[1][1]/P0001 ,
		\u10_mem_reg[3][1]/P0001 ,
		\u10_rp_reg[0]/P0001 ,
		\u10_rp_reg[1]/P0001 ,
		_w6741_
	);
	LUT2 #(
		.INIT('h7)
	) name4595 (
		_w6740_,
		_w6741_,
		_w6742_
	);
	LUT4 #(
		.INIT('hff35)
	) name4596 (
		\u11_mem_reg[0][6]/P0001 ,
		\u11_mem_reg[1][6]/P0001 ,
		\u11_rp_reg[0]/P0001 ,
		\u11_rp_reg[1]/P0001 ,
		_w6743_
	);
	LUT4 #(
		.INIT('h35ff)
	) name4597 (
		\u11_mem_reg[2][6]/P0001 ,
		\u11_mem_reg[3][6]/P0001 ,
		\u11_rp_reg[0]/P0001 ,
		\u11_rp_reg[1]/P0001 ,
		_w6744_
	);
	LUT2 #(
		.INIT('h7)
	) name4598 (
		_w6743_,
		_w6744_,
		_w6745_
	);
	LUT4 #(
		.INIT('hf3f5)
	) name4599 (
		\u10_mem_reg[0][20]/P0001 ,
		\u10_mem_reg[2][20]/P0001 ,
		\u10_rp_reg[0]/P0001 ,
		\u10_rp_reg[1]/P0001 ,
		_w6746_
	);
	LUT4 #(
		.INIT('h3f5f)
	) name4600 (
		\u10_mem_reg[1][20]/P0001 ,
		\u10_mem_reg[3][20]/P0001 ,
		\u10_rp_reg[0]/P0001 ,
		\u10_rp_reg[1]/P0001 ,
		_w6747_
	);
	LUT2 #(
		.INIT('h7)
	) name4601 (
		_w6746_,
		_w6747_,
		_w6748_
	);
	LUT4 #(
		.INIT('hf3f5)
	) name4602 (
		\u10_mem_reg[0][21]/P0001 ,
		\u10_mem_reg[2][21]/P0001 ,
		\u10_rp_reg[0]/P0001 ,
		\u10_rp_reg[1]/P0001 ,
		_w6749_
	);
	LUT4 #(
		.INIT('h3f5f)
	) name4603 (
		\u10_mem_reg[1][21]/P0001 ,
		\u10_mem_reg[3][21]/P0001 ,
		\u10_rp_reg[0]/P0001 ,
		\u10_rp_reg[1]/P0001 ,
		_w6750_
	);
	LUT2 #(
		.INIT('h7)
	) name4604 (
		_w6749_,
		_w6750_,
		_w6751_
	);
	LUT4 #(
		.INIT('hf35f)
	) name4605 (
		\u10_mem_reg[1][22]/P0001 ,
		\u10_mem_reg[2][22]/P0001 ,
		\u10_rp_reg[0]/P0001 ,
		\u10_rp_reg[1]/P0001 ,
		_w6752_
	);
	LUT4 #(
		.INIT('h3ff5)
	) name4606 (
		\u10_mem_reg[0][22]/P0001 ,
		\u10_mem_reg[3][22]/P0001 ,
		\u10_rp_reg[0]/P0001 ,
		\u10_rp_reg[1]/P0001 ,
		_w6753_
	);
	LUT2 #(
		.INIT('h7)
	) name4607 (
		_w6752_,
		_w6753_,
		_w6754_
	);
	LUT4 #(
		.INIT('hf3f5)
	) name4608 (
		\u10_mem_reg[0][23]/P0001 ,
		\u10_mem_reg[2][23]/P0001 ,
		\u10_rp_reg[0]/P0001 ,
		\u10_rp_reg[1]/P0001 ,
		_w6755_
	);
	LUT4 #(
		.INIT('h3f5f)
	) name4609 (
		\u10_mem_reg[1][23]/P0001 ,
		\u10_mem_reg[3][23]/P0001 ,
		\u10_rp_reg[0]/P0001 ,
		\u10_rp_reg[1]/P0001 ,
		_w6756_
	);
	LUT2 #(
		.INIT('h7)
	) name4610 (
		_w6755_,
		_w6756_,
		_w6757_
	);
	LUT4 #(
		.INIT('hf35f)
	) name4611 (
		\u10_mem_reg[1][24]/P0001 ,
		\u10_mem_reg[2][24]/P0001 ,
		\u10_rp_reg[0]/P0001 ,
		\u10_rp_reg[1]/P0001 ,
		_w6758_
	);
	LUT4 #(
		.INIT('h3ff5)
	) name4612 (
		\u10_mem_reg[0][24]/P0001 ,
		\u10_mem_reg[3][24]/P0001 ,
		\u10_rp_reg[0]/P0001 ,
		\u10_rp_reg[1]/P0001 ,
		_w6759_
	);
	LUT2 #(
		.INIT('h7)
	) name4613 (
		_w6758_,
		_w6759_,
		_w6760_
	);
	LUT4 #(
		.INIT('hf35f)
	) name4614 (
		\u10_mem_reg[1][25]/P0001 ,
		\u10_mem_reg[2][25]/P0001 ,
		\u10_rp_reg[0]/P0001 ,
		\u10_rp_reg[1]/P0001 ,
		_w6761_
	);
	LUT4 #(
		.INIT('h3ff5)
	) name4615 (
		\u10_mem_reg[0][25]/P0001 ,
		\u10_mem_reg[3][25]/P0001 ,
		\u10_rp_reg[0]/P0001 ,
		\u10_rp_reg[1]/P0001 ,
		_w6762_
	);
	LUT2 #(
		.INIT('h7)
	) name4616 (
		_w6761_,
		_w6762_,
		_w6763_
	);
	LUT4 #(
		.INIT('hf35f)
	) name4617 (
		\u10_mem_reg[1][26]/P0001 ,
		\u10_mem_reg[2][26]/P0001 ,
		\u10_rp_reg[0]/P0001 ,
		\u10_rp_reg[1]/P0001 ,
		_w6764_
	);
	LUT4 #(
		.INIT('h3ff5)
	) name4618 (
		\u10_mem_reg[0][26]/P0001 ,
		\u10_mem_reg[3][26]/P0001 ,
		\u10_rp_reg[0]/P0001 ,
		\u10_rp_reg[1]/P0001 ,
		_w6765_
	);
	LUT2 #(
		.INIT('h7)
	) name4619 (
		_w6764_,
		_w6765_,
		_w6766_
	);
	LUT4 #(
		.INIT('hf3f5)
	) name4620 (
		\u10_mem_reg[0][27]/P0001 ,
		\u10_mem_reg[2][27]/P0001 ,
		\u10_rp_reg[0]/P0001 ,
		\u10_rp_reg[1]/P0001 ,
		_w6767_
	);
	LUT4 #(
		.INIT('h3f5f)
	) name4621 (
		\u10_mem_reg[1][27]/P0001 ,
		\u10_mem_reg[3][27]/P0001 ,
		\u10_rp_reg[0]/P0001 ,
		\u10_rp_reg[1]/P0001 ,
		_w6768_
	);
	LUT2 #(
		.INIT('h7)
	) name4622 (
		_w6767_,
		_w6768_,
		_w6769_
	);
	LUT4 #(
		.INIT('hff35)
	) name4623 (
		\u9_mem_reg[0][4]/P0001 ,
		\u9_mem_reg[1][4]/P0001 ,
		\u9_rp_reg[0]/P0001 ,
		\u9_rp_reg[1]/P0001 ,
		_w6770_
	);
	LUT4 #(
		.INIT('h35ff)
	) name4624 (
		\u9_mem_reg[2][4]/P0001 ,
		\u9_mem_reg[3][4]/P0001 ,
		\u9_rp_reg[0]/P0001 ,
		\u9_rp_reg[1]/P0001 ,
		_w6771_
	);
	LUT2 #(
		.INIT('h7)
	) name4625 (
		_w6770_,
		_w6771_,
		_w6772_
	);
	LUT4 #(
		.INIT('hf3f5)
	) name4626 (
		\u10_mem_reg[0][28]/P0001 ,
		\u10_mem_reg[2][28]/P0001 ,
		\u10_rp_reg[0]/P0001 ,
		\u10_rp_reg[1]/P0001 ,
		_w6773_
	);
	LUT4 #(
		.INIT('h3f5f)
	) name4627 (
		\u10_mem_reg[1][28]/P0001 ,
		\u10_mem_reg[3][28]/P0001 ,
		\u10_rp_reg[0]/P0001 ,
		\u10_rp_reg[1]/P0001 ,
		_w6774_
	);
	LUT2 #(
		.INIT('h7)
	) name4628 (
		_w6773_,
		_w6774_,
		_w6775_
	);
	LUT4 #(
		.INIT('hf35f)
	) name4629 (
		\u10_mem_reg[1][29]/P0001 ,
		\u10_mem_reg[2][29]/P0001 ,
		\u10_rp_reg[0]/P0001 ,
		\u10_rp_reg[1]/P0001 ,
		_w6776_
	);
	LUT4 #(
		.INIT('h3ff5)
	) name4630 (
		\u10_mem_reg[0][29]/P0001 ,
		\u10_mem_reg[3][29]/P0001 ,
		\u10_rp_reg[0]/P0001 ,
		\u10_rp_reg[1]/P0001 ,
		_w6777_
	);
	LUT2 #(
		.INIT('h7)
	) name4631 (
		_w6776_,
		_w6777_,
		_w6778_
	);
	LUT4 #(
		.INIT('hff35)
	) name4632 (
		\u11_mem_reg[0][0]/P0001 ,
		\u11_mem_reg[1][0]/P0001 ,
		\u11_rp_reg[0]/P0001 ,
		\u11_rp_reg[1]/P0001 ,
		_w6779_
	);
	LUT4 #(
		.INIT('h35ff)
	) name4633 (
		\u11_mem_reg[2][0]/P0001 ,
		\u11_mem_reg[3][0]/P0001 ,
		\u11_rp_reg[0]/P0001 ,
		\u11_rp_reg[1]/P0001 ,
		_w6780_
	);
	LUT2 #(
		.INIT('h7)
	) name4634 (
		_w6779_,
		_w6780_,
		_w6781_
	);
	LUT4 #(
		.INIT('hff35)
	) name4635 (
		\u11_mem_reg[0][10]/P0001 ,
		\u11_mem_reg[1][10]/P0001 ,
		\u11_rp_reg[0]/P0001 ,
		\u11_rp_reg[1]/P0001 ,
		_w6782_
	);
	LUT4 #(
		.INIT('h35ff)
	) name4636 (
		\u11_mem_reg[2][10]/P0001 ,
		\u11_mem_reg[3][10]/P0001 ,
		\u11_rp_reg[0]/P0001 ,
		\u11_rp_reg[1]/P0001 ,
		_w6783_
	);
	LUT2 #(
		.INIT('h7)
	) name4637 (
		_w6782_,
		_w6783_,
		_w6784_
	);
	LUT4 #(
		.INIT('hf3f5)
	) name4638 (
		\u10_mem_reg[0][30]/P0001 ,
		\u10_mem_reg[2][30]/P0001 ,
		\u10_rp_reg[0]/P0001 ,
		\u10_rp_reg[1]/P0001 ,
		_w6785_
	);
	LUT4 #(
		.INIT('h3f5f)
	) name4639 (
		\u10_mem_reg[1][30]/P0001 ,
		\u10_mem_reg[3][30]/P0001 ,
		\u10_rp_reg[0]/P0001 ,
		\u10_rp_reg[1]/P0001 ,
		_w6786_
	);
	LUT2 #(
		.INIT('h7)
	) name4640 (
		_w6785_,
		_w6786_,
		_w6787_
	);
	LUT4 #(
		.INIT('hff35)
	) name4641 (
		\u11_mem_reg[0][11]/P0001 ,
		\u11_mem_reg[1][11]/P0001 ,
		\u11_rp_reg[0]/P0001 ,
		\u11_rp_reg[1]/P0001 ,
		_w6788_
	);
	LUT4 #(
		.INIT('h35ff)
	) name4642 (
		\u11_mem_reg[2][11]/P0001 ,
		\u11_mem_reg[3][11]/P0001 ,
		\u11_rp_reg[0]/P0001 ,
		\u11_rp_reg[1]/P0001 ,
		_w6789_
	);
	LUT2 #(
		.INIT('h7)
	) name4643 (
		_w6788_,
		_w6789_,
		_w6790_
	);
	LUT4 #(
		.INIT('hff35)
	) name4644 (
		\u11_mem_reg[0][12]/P0001 ,
		\u11_mem_reg[1][12]/P0001 ,
		\u11_rp_reg[0]/P0001 ,
		\u11_rp_reg[1]/P0001 ,
		_w6791_
	);
	LUT4 #(
		.INIT('h35ff)
	) name4645 (
		\u11_mem_reg[2][12]/P0001 ,
		\u11_mem_reg[3][12]/P0001 ,
		\u11_rp_reg[0]/P0001 ,
		\u11_rp_reg[1]/P0001 ,
		_w6792_
	);
	LUT2 #(
		.INIT('h7)
	) name4646 (
		_w6791_,
		_w6792_,
		_w6793_
	);
	LUT4 #(
		.INIT('hff35)
	) name4647 (
		\u11_mem_reg[0][13]/P0001 ,
		\u11_mem_reg[1][13]/P0001 ,
		\u11_rp_reg[0]/P0001 ,
		\u11_rp_reg[1]/P0001 ,
		_w6794_
	);
	LUT4 #(
		.INIT('h35ff)
	) name4648 (
		\u11_mem_reg[2][13]/P0001 ,
		\u11_mem_reg[3][13]/P0001 ,
		\u11_rp_reg[0]/P0001 ,
		\u11_rp_reg[1]/P0001 ,
		_w6795_
	);
	LUT2 #(
		.INIT('h7)
	) name4649 (
		_w6794_,
		_w6795_,
		_w6796_
	);
	LUT4 #(
		.INIT('hf3f5)
	) name4650 (
		\u11_mem_reg[0][14]/P0001 ,
		\u11_mem_reg[2][14]/P0001 ,
		\u11_rp_reg[0]/P0001 ,
		\u11_rp_reg[1]/P0001 ,
		_w6797_
	);
	LUT4 #(
		.INIT('h3f5f)
	) name4651 (
		\u11_mem_reg[1][14]/P0001 ,
		\u11_mem_reg[3][14]/P0001 ,
		\u11_rp_reg[0]/P0001 ,
		\u11_rp_reg[1]/P0001 ,
		_w6798_
	);
	LUT2 #(
		.INIT('h7)
	) name4652 (
		_w6797_,
		_w6798_,
		_w6799_
	);
	LUT4 #(
		.INIT('hf35f)
	) name4653 (
		\u10_mem_reg[1][3]/P0001 ,
		\u10_mem_reg[2][3]/P0001 ,
		\u10_rp_reg[0]/P0001 ,
		\u10_rp_reg[1]/P0001 ,
		_w6800_
	);
	LUT4 #(
		.INIT('h3ff5)
	) name4654 (
		\u10_mem_reg[0][3]/P0001 ,
		\u10_mem_reg[3][3]/P0001 ,
		\u10_rp_reg[0]/P0001 ,
		\u10_rp_reg[1]/P0001 ,
		_w6801_
	);
	LUT2 #(
		.INIT('h7)
	) name4655 (
		_w6800_,
		_w6801_,
		_w6802_
	);
	LUT4 #(
		.INIT('hff35)
	) name4656 (
		\u11_mem_reg[0][15]/P0001 ,
		\u11_mem_reg[1][15]/P0001 ,
		\u11_rp_reg[0]/P0001 ,
		\u11_rp_reg[1]/P0001 ,
		_w6803_
	);
	LUT4 #(
		.INIT('h35ff)
	) name4657 (
		\u11_mem_reg[2][15]/P0001 ,
		\u11_mem_reg[3][15]/P0001 ,
		\u11_rp_reg[0]/P0001 ,
		\u11_rp_reg[1]/P0001 ,
		_w6804_
	);
	LUT2 #(
		.INIT('h7)
	) name4658 (
		_w6803_,
		_w6804_,
		_w6805_
	);
	LUT4 #(
		.INIT('hff35)
	) name4659 (
		\u11_mem_reg[0][16]/P0001 ,
		\u11_mem_reg[1][16]/P0001 ,
		\u11_rp_reg[0]/P0001 ,
		\u11_rp_reg[1]/P0001 ,
		_w6806_
	);
	LUT4 #(
		.INIT('h35ff)
	) name4660 (
		\u11_mem_reg[2][16]/P0001 ,
		\u11_mem_reg[3][16]/P0001 ,
		\u11_rp_reg[0]/P0001 ,
		\u11_rp_reg[1]/P0001 ,
		_w6807_
	);
	LUT2 #(
		.INIT('h7)
	) name4661 (
		_w6806_,
		_w6807_,
		_w6808_
	);
	LUT4 #(
		.INIT('hf35f)
	) name4662 (
		\u10_mem_reg[1][4]/P0001 ,
		\u10_mem_reg[2][4]/P0001 ,
		\u10_rp_reg[0]/P0001 ,
		\u10_rp_reg[1]/P0001 ,
		_w6809_
	);
	LUT4 #(
		.INIT('h3ff5)
	) name4663 (
		\u10_mem_reg[0][4]/P0001 ,
		\u10_mem_reg[3][4]/P0001 ,
		\u10_rp_reg[0]/P0001 ,
		\u10_rp_reg[1]/P0001 ,
		_w6810_
	);
	LUT2 #(
		.INIT('h7)
	) name4664 (
		_w6809_,
		_w6810_,
		_w6811_
	);
	LUT4 #(
		.INIT('hff35)
	) name4665 (
		\u11_mem_reg[0][17]/P0001 ,
		\u11_mem_reg[1][17]/P0001 ,
		\u11_rp_reg[0]/P0001 ,
		\u11_rp_reg[1]/P0001 ,
		_w6812_
	);
	LUT4 #(
		.INIT('h35ff)
	) name4666 (
		\u11_mem_reg[2][17]/P0001 ,
		\u11_mem_reg[3][17]/P0001 ,
		\u11_rp_reg[0]/P0001 ,
		\u11_rp_reg[1]/P0001 ,
		_w6813_
	);
	LUT2 #(
		.INIT('h7)
	) name4667 (
		_w6812_,
		_w6813_,
		_w6814_
	);
	LUT4 #(
		.INIT('hf35f)
	) name4668 (
		\u11_mem_reg[1][18]/P0001 ,
		\u11_mem_reg[2][18]/P0001 ,
		\u11_rp_reg[0]/P0001 ,
		\u11_rp_reg[1]/P0001 ,
		_w6815_
	);
	LUT4 #(
		.INIT('h3ff5)
	) name4669 (
		\u11_mem_reg[0][18]/P0001 ,
		\u11_mem_reg[3][18]/P0001 ,
		\u11_rp_reg[0]/P0001 ,
		\u11_rp_reg[1]/P0001 ,
		_w6816_
	);
	LUT2 #(
		.INIT('h7)
	) name4670 (
		_w6815_,
		_w6816_,
		_w6817_
	);
	LUT4 #(
		.INIT('hf3f5)
	) name4671 (
		\u10_mem_reg[0][5]/P0001 ,
		\u10_mem_reg[2][5]/P0001 ,
		\u10_rp_reg[0]/P0001 ,
		\u10_rp_reg[1]/P0001 ,
		_w6818_
	);
	LUT4 #(
		.INIT('h3f5f)
	) name4672 (
		\u10_mem_reg[1][5]/P0001 ,
		\u10_mem_reg[3][5]/P0001 ,
		\u10_rp_reg[0]/P0001 ,
		\u10_rp_reg[1]/P0001 ,
		_w6819_
	);
	LUT2 #(
		.INIT('h7)
	) name4673 (
		_w6818_,
		_w6819_,
		_w6820_
	);
	LUT4 #(
		.INIT('hf35f)
	) name4674 (
		\u11_mem_reg[1][19]/P0001 ,
		\u11_mem_reg[2][19]/P0001 ,
		\u11_rp_reg[0]/P0001 ,
		\u11_rp_reg[1]/P0001 ,
		_w6821_
	);
	LUT4 #(
		.INIT('h3ff5)
	) name4675 (
		\u11_mem_reg[0][19]/P0001 ,
		\u11_mem_reg[3][19]/P0001 ,
		\u11_rp_reg[0]/P0001 ,
		\u11_rp_reg[1]/P0001 ,
		_w6822_
	);
	LUT2 #(
		.INIT('h7)
	) name4676 (
		_w6821_,
		_w6822_,
		_w6823_
	);
	LUT4 #(
		.INIT('hff35)
	) name4677 (
		\u11_mem_reg[0][1]/P0001 ,
		\u11_mem_reg[1][1]/P0001 ,
		\u11_rp_reg[0]/P0001 ,
		\u11_rp_reg[1]/P0001 ,
		_w6824_
	);
	LUT4 #(
		.INIT('h35ff)
	) name4678 (
		\u11_mem_reg[2][1]/P0001 ,
		\u11_mem_reg[3][1]/P0001 ,
		\u11_rp_reg[0]/P0001 ,
		\u11_rp_reg[1]/P0001 ,
		_w6825_
	);
	LUT2 #(
		.INIT('h7)
	) name4679 (
		_w6824_,
		_w6825_,
		_w6826_
	);
	LUT4 #(
		.INIT('hf35f)
	) name4680 (
		\u10_mem_reg[1][6]/P0001 ,
		\u10_mem_reg[2][6]/P0001 ,
		\u10_rp_reg[0]/P0001 ,
		\u10_rp_reg[1]/P0001 ,
		_w6827_
	);
	LUT4 #(
		.INIT('h3ff5)
	) name4681 (
		\u10_mem_reg[0][6]/P0001 ,
		\u10_mem_reg[3][6]/P0001 ,
		\u10_rp_reg[0]/P0001 ,
		\u10_rp_reg[1]/P0001 ,
		_w6828_
	);
	LUT2 #(
		.INIT('h7)
	) name4682 (
		_w6827_,
		_w6828_,
		_w6829_
	);
	LUT4 #(
		.INIT('hf35f)
	) name4683 (
		\u11_mem_reg[1][20]/P0001 ,
		\u11_mem_reg[2][20]/P0001 ,
		\u11_rp_reg[0]/P0001 ,
		\u11_rp_reg[1]/P0001 ,
		_w6830_
	);
	LUT4 #(
		.INIT('h3ff5)
	) name4684 (
		\u11_mem_reg[0][20]/P0001 ,
		\u11_mem_reg[3][20]/P0001 ,
		\u11_rp_reg[0]/P0001 ,
		\u11_rp_reg[1]/P0001 ,
		_w6831_
	);
	LUT2 #(
		.INIT('h7)
	) name4685 (
		_w6830_,
		_w6831_,
		_w6832_
	);
	LUT4 #(
		.INIT('hf35f)
	) name4686 (
		\u11_mem_reg[1][21]/P0001 ,
		\u11_mem_reg[2][21]/P0001 ,
		\u11_rp_reg[0]/P0001 ,
		\u11_rp_reg[1]/P0001 ,
		_w6833_
	);
	LUT4 #(
		.INIT('h3ff5)
	) name4687 (
		\u11_mem_reg[0][21]/P0001 ,
		\u11_mem_reg[3][21]/P0001 ,
		\u11_rp_reg[0]/P0001 ,
		\u11_rp_reg[1]/P0001 ,
		_w6834_
	);
	LUT2 #(
		.INIT('h7)
	) name4688 (
		_w6833_,
		_w6834_,
		_w6835_
	);
	LUT4 #(
		.INIT('hf35f)
	) name4689 (
		\u10_mem_reg[1][7]/P0001 ,
		\u10_mem_reg[2][7]/P0001 ,
		\u10_rp_reg[0]/P0001 ,
		\u10_rp_reg[1]/P0001 ,
		_w6836_
	);
	LUT4 #(
		.INIT('h3ff5)
	) name4690 (
		\u10_mem_reg[0][7]/P0001 ,
		\u10_mem_reg[3][7]/P0001 ,
		\u10_rp_reg[0]/P0001 ,
		\u10_rp_reg[1]/P0001 ,
		_w6837_
	);
	LUT2 #(
		.INIT('h7)
	) name4691 (
		_w6836_,
		_w6837_,
		_w6838_
	);
	LUT4 #(
		.INIT('hf35f)
	) name4692 (
		\u11_mem_reg[1][22]/P0001 ,
		\u11_mem_reg[2][22]/P0001 ,
		\u11_rp_reg[0]/P0001 ,
		\u11_rp_reg[1]/P0001 ,
		_w6839_
	);
	LUT4 #(
		.INIT('h3ff5)
	) name4693 (
		\u11_mem_reg[0][22]/P0001 ,
		\u11_mem_reg[3][22]/P0001 ,
		\u11_rp_reg[0]/P0001 ,
		\u11_rp_reg[1]/P0001 ,
		_w6840_
	);
	LUT2 #(
		.INIT('h7)
	) name4694 (
		_w6839_,
		_w6840_,
		_w6841_
	);
	LUT4 #(
		.INIT('hf35f)
	) name4695 (
		\u11_mem_reg[1][23]/P0001 ,
		\u11_mem_reg[2][23]/P0001 ,
		\u11_rp_reg[0]/P0001 ,
		\u11_rp_reg[1]/P0001 ,
		_w6842_
	);
	LUT4 #(
		.INIT('h3ff5)
	) name4696 (
		\u11_mem_reg[0][23]/P0001 ,
		\u11_mem_reg[3][23]/P0001 ,
		\u11_rp_reg[0]/P0001 ,
		\u11_rp_reg[1]/P0001 ,
		_w6843_
	);
	LUT2 #(
		.INIT('h7)
	) name4697 (
		_w6842_,
		_w6843_,
		_w6844_
	);
	LUT4 #(
		.INIT('hf3f5)
	) name4698 (
		\u10_mem_reg[0][8]/P0001 ,
		\u10_mem_reg[2][8]/P0001 ,
		\u10_rp_reg[0]/P0001 ,
		\u10_rp_reg[1]/P0001 ,
		_w6845_
	);
	LUT4 #(
		.INIT('h3f5f)
	) name4699 (
		\u10_mem_reg[1][8]/P0001 ,
		\u10_mem_reg[3][8]/P0001 ,
		\u10_rp_reg[0]/P0001 ,
		\u10_rp_reg[1]/P0001 ,
		_w6846_
	);
	LUT2 #(
		.INIT('h7)
	) name4700 (
		_w6845_,
		_w6846_,
		_w6847_
	);
	LUT4 #(
		.INIT('hf35f)
	) name4701 (
		\u11_mem_reg[1][24]/P0001 ,
		\u11_mem_reg[2][24]/P0001 ,
		\u11_rp_reg[0]/P0001 ,
		\u11_rp_reg[1]/P0001 ,
		_w6848_
	);
	LUT4 #(
		.INIT('h3ff5)
	) name4702 (
		\u11_mem_reg[0][24]/P0001 ,
		\u11_mem_reg[3][24]/P0001 ,
		\u11_rp_reg[0]/P0001 ,
		\u11_rp_reg[1]/P0001 ,
		_w6849_
	);
	LUT2 #(
		.INIT('h7)
	) name4703 (
		_w6848_,
		_w6849_,
		_w6850_
	);
	LUT4 #(
		.INIT('hf35f)
	) name4704 (
		\u11_mem_reg[1][25]/P0001 ,
		\u11_mem_reg[2][25]/P0001 ,
		\u11_rp_reg[0]/P0001 ,
		\u11_rp_reg[1]/P0001 ,
		_w6851_
	);
	LUT4 #(
		.INIT('h3ff5)
	) name4705 (
		\u11_mem_reg[0][25]/P0001 ,
		\u11_mem_reg[3][25]/P0001 ,
		\u11_rp_reg[0]/P0001 ,
		\u11_rp_reg[1]/P0001 ,
		_w6852_
	);
	LUT2 #(
		.INIT('h7)
	) name4706 (
		_w6851_,
		_w6852_,
		_w6853_
	);
	LUT4 #(
		.INIT('hff35)
	) name4707 (
		\u10_mem_reg[0][9]/P0001 ,
		\u10_mem_reg[1][9]/P0001 ,
		\u10_rp_reg[0]/P0001 ,
		\u10_rp_reg[1]/P0001 ,
		_w6854_
	);
	LUT4 #(
		.INIT('h35ff)
	) name4708 (
		\u10_mem_reg[2][9]/P0001 ,
		\u10_mem_reg[3][9]/P0001 ,
		\u10_rp_reg[0]/P0001 ,
		\u10_rp_reg[1]/P0001 ,
		_w6855_
	);
	LUT2 #(
		.INIT('h7)
	) name4709 (
		_w6854_,
		_w6855_,
		_w6856_
	);
	LUT4 #(
		.INIT('hf35f)
	) name4710 (
		\u11_mem_reg[1][26]/P0001 ,
		\u11_mem_reg[2][26]/P0001 ,
		\u11_rp_reg[0]/P0001 ,
		\u11_rp_reg[1]/P0001 ,
		_w6857_
	);
	LUT4 #(
		.INIT('h3ff5)
	) name4711 (
		\u11_mem_reg[0][26]/P0001 ,
		\u11_mem_reg[3][26]/P0001 ,
		\u11_rp_reg[0]/P0001 ,
		\u11_rp_reg[1]/P0001 ,
		_w6858_
	);
	LUT2 #(
		.INIT('h7)
	) name4712 (
		_w6857_,
		_w6858_,
		_w6859_
	);
	LUT4 #(
		.INIT('hf35f)
	) name4713 (
		\u11_mem_reg[1][27]/P0001 ,
		\u11_mem_reg[2][27]/P0001 ,
		\u11_rp_reg[0]/P0001 ,
		\u11_rp_reg[1]/P0001 ,
		_w6860_
	);
	LUT4 #(
		.INIT('h3ff5)
	) name4714 (
		\u11_mem_reg[0][27]/P0001 ,
		\u11_mem_reg[3][27]/P0001 ,
		\u11_rp_reg[0]/P0001 ,
		\u11_rp_reg[1]/P0001 ,
		_w6861_
	);
	LUT2 #(
		.INIT('h7)
	) name4715 (
		_w6860_,
		_w6861_,
		_w6862_
	);
	LUT4 #(
		.INIT('hf35f)
	) name4716 (
		\u11_mem_reg[1][28]/P0001 ,
		\u11_mem_reg[2][28]/P0001 ,
		\u11_rp_reg[0]/P0001 ,
		\u11_rp_reg[1]/P0001 ,
		_w6863_
	);
	LUT4 #(
		.INIT('h3ff5)
	) name4717 (
		\u11_mem_reg[0][28]/P0001 ,
		\u11_mem_reg[3][28]/P0001 ,
		\u11_rp_reg[0]/P0001 ,
		\u11_rp_reg[1]/P0001 ,
		_w6864_
	);
	LUT2 #(
		.INIT('h7)
	) name4718 (
		_w6863_,
		_w6864_,
		_w6865_
	);
	LUT4 #(
		.INIT('h35ff)
	) name4719 (
		\u10_mem_reg[2][14]/P0001 ,
		\u10_mem_reg[3][14]/P0001 ,
		\u10_rp_reg[0]/P0001 ,
		\u10_rp_reg[1]/P0001 ,
		_w6866_
	);
	LUT4 #(
		.INIT('hff35)
	) name4720 (
		\u10_mem_reg[0][14]/P0001 ,
		\u10_mem_reg[1][14]/P0001 ,
		\u10_rp_reg[0]/P0001 ,
		\u10_rp_reg[1]/P0001 ,
		_w6867_
	);
	LUT2 #(
		.INIT('h7)
	) name4721 (
		_w6866_,
		_w6867_,
		_w6868_
	);
	LUT4 #(
		.INIT('hf35f)
	) name4722 (
		\u11_mem_reg[1][29]/P0001 ,
		\u11_mem_reg[2][29]/P0001 ,
		\u11_rp_reg[0]/P0001 ,
		\u11_rp_reg[1]/P0001 ,
		_w6869_
	);
	LUT4 #(
		.INIT('h3ff5)
	) name4723 (
		\u11_mem_reg[0][29]/P0001 ,
		\u11_mem_reg[3][29]/P0001 ,
		\u11_rp_reg[0]/P0001 ,
		\u11_rp_reg[1]/P0001 ,
		_w6870_
	);
	LUT2 #(
		.INIT('h7)
	) name4724 (
		_w6869_,
		_w6870_,
		_w6871_
	);
	LUT4 #(
		.INIT('hff35)
	) name4725 (
		\u11_mem_reg[0][2]/P0001 ,
		\u11_mem_reg[1][2]/P0001 ,
		\u11_rp_reg[0]/P0001 ,
		\u11_rp_reg[1]/P0001 ,
		_w6872_
	);
	LUT4 #(
		.INIT('h35ff)
	) name4726 (
		\u11_mem_reg[2][2]/P0001 ,
		\u11_mem_reg[3][2]/P0001 ,
		\u11_rp_reg[0]/P0001 ,
		\u11_rp_reg[1]/P0001 ,
		_w6873_
	);
	LUT2 #(
		.INIT('h7)
	) name4727 (
		_w6872_,
		_w6873_,
		_w6874_
	);
	LUT4 #(
		.INIT('hf35f)
	) name4728 (
		\u11_mem_reg[1][30]/P0001 ,
		\u11_mem_reg[2][30]/P0001 ,
		\u11_rp_reg[0]/P0001 ,
		\u11_rp_reg[1]/P0001 ,
		_w6875_
	);
	LUT4 #(
		.INIT('h3ff5)
	) name4729 (
		\u11_mem_reg[0][30]/P0001 ,
		\u11_mem_reg[3][30]/P0001 ,
		\u11_rp_reg[0]/P0001 ,
		\u11_rp_reg[1]/P0001 ,
		_w6876_
	);
	LUT2 #(
		.INIT('h7)
	) name4730 (
		_w6875_,
		_w6876_,
		_w6877_
	);
	LUT4 #(
		.INIT('hf35f)
	) name4731 (
		\u11_mem_reg[1][31]/P0001 ,
		\u11_mem_reg[2][31]/P0001 ,
		\u11_rp_reg[0]/P0001 ,
		\u11_rp_reg[1]/P0001 ,
		_w6878_
	);
	LUT4 #(
		.INIT('h3ff5)
	) name4732 (
		\u11_mem_reg[0][31]/P0001 ,
		\u11_mem_reg[3][31]/P0001 ,
		\u11_rp_reg[0]/P0001 ,
		\u11_rp_reg[1]/P0001 ,
		_w6879_
	);
	LUT2 #(
		.INIT('h7)
	) name4733 (
		_w6878_,
		_w6879_,
		_w6880_
	);
	LUT4 #(
		.INIT('hff35)
	) name4734 (
		\u11_mem_reg[0][3]/P0001 ,
		\u11_mem_reg[1][3]/P0001 ,
		\u11_rp_reg[0]/P0001 ,
		\u11_rp_reg[1]/P0001 ,
		_w6881_
	);
	LUT4 #(
		.INIT('h35ff)
	) name4735 (
		\u11_mem_reg[2][3]/P0001 ,
		\u11_mem_reg[3][3]/P0001 ,
		\u11_rp_reg[0]/P0001 ,
		\u11_rp_reg[1]/P0001 ,
		_w6882_
	);
	LUT2 #(
		.INIT('h7)
	) name4736 (
		_w6881_,
		_w6882_,
		_w6883_
	);
	LUT4 #(
		.INIT('hff35)
	) name4737 (
		\u11_mem_reg[0][4]/P0001 ,
		\u11_mem_reg[1][4]/P0001 ,
		\u11_rp_reg[0]/P0001 ,
		\u11_rp_reg[1]/P0001 ,
		_w6884_
	);
	LUT4 #(
		.INIT('h35ff)
	) name4738 (
		\u11_mem_reg[2][4]/P0001 ,
		\u11_mem_reg[3][4]/P0001 ,
		\u11_rp_reg[0]/P0001 ,
		\u11_rp_reg[1]/P0001 ,
		_w6885_
	);
	LUT2 #(
		.INIT('h7)
	) name4739 (
		_w6884_,
		_w6885_,
		_w6886_
	);
	LUT4 #(
		.INIT('hff35)
	) name4740 (
		\u11_mem_reg[0][5]/P0001 ,
		\u11_mem_reg[1][5]/P0001 ,
		\u11_rp_reg[0]/P0001 ,
		\u11_rp_reg[1]/P0001 ,
		_w6887_
	);
	LUT4 #(
		.INIT('h35ff)
	) name4741 (
		\u11_mem_reg[2][5]/P0001 ,
		\u11_mem_reg[3][5]/P0001 ,
		\u11_rp_reg[0]/P0001 ,
		\u11_rp_reg[1]/P0001 ,
		_w6888_
	);
	LUT2 #(
		.INIT('h7)
	) name4742 (
		_w6887_,
		_w6888_,
		_w6889_
	);
	LUT4 #(
		.INIT('hf3f5)
	) name4743 (
		\u11_mem_reg[0][7]/P0001 ,
		\u11_mem_reg[2][7]/P0001 ,
		\u11_rp_reg[0]/P0001 ,
		\u11_rp_reg[1]/P0001 ,
		_w6890_
	);
	LUT4 #(
		.INIT('h3f5f)
	) name4744 (
		\u11_mem_reg[1][7]/P0001 ,
		\u11_mem_reg[3][7]/P0001 ,
		\u11_rp_reg[0]/P0001 ,
		\u11_rp_reg[1]/P0001 ,
		_w6891_
	);
	LUT2 #(
		.INIT('h7)
	) name4745 (
		_w6890_,
		_w6891_,
		_w6892_
	);
	LUT4 #(
		.INIT('hff35)
	) name4746 (
		\u11_mem_reg[0][8]/P0001 ,
		\u11_mem_reg[1][8]/P0001 ,
		\u11_rp_reg[0]/P0001 ,
		\u11_rp_reg[1]/P0001 ,
		_w6893_
	);
	LUT4 #(
		.INIT('h35ff)
	) name4747 (
		\u11_mem_reg[2][8]/P0001 ,
		\u11_mem_reg[3][8]/P0001 ,
		\u11_rp_reg[0]/P0001 ,
		\u11_rp_reg[1]/P0001 ,
		_w6894_
	);
	LUT2 #(
		.INIT('h7)
	) name4748 (
		_w6893_,
		_w6894_,
		_w6895_
	);
	LUT4 #(
		.INIT('hff35)
	) name4749 (
		\u11_mem_reg[0][9]/P0001 ,
		\u11_mem_reg[1][9]/P0001 ,
		\u11_rp_reg[0]/P0001 ,
		\u11_rp_reg[1]/P0001 ,
		_w6896_
	);
	LUT4 #(
		.INIT('h35ff)
	) name4750 (
		\u11_mem_reg[2][9]/P0001 ,
		\u11_mem_reg[3][9]/P0001 ,
		\u11_rp_reg[0]/P0001 ,
		\u11_rp_reg[1]/P0001 ,
		_w6897_
	);
	LUT2 #(
		.INIT('h7)
	) name4751 (
		_w6896_,
		_w6897_,
		_w6898_
	);
	LUT4 #(
		.INIT('hf3f5)
	) name4752 (
		\u10_mem_reg[0][10]/P0001 ,
		\u10_mem_reg[2][10]/P0001 ,
		\u10_rp_reg[0]/P0001 ,
		\u10_rp_reg[1]/P0001 ,
		_w6899_
	);
	LUT4 #(
		.INIT('h3f5f)
	) name4753 (
		\u10_mem_reg[1][10]/P0001 ,
		\u10_mem_reg[3][10]/P0001 ,
		\u10_rp_reg[0]/P0001 ,
		\u10_rp_reg[1]/P0001 ,
		_w6900_
	);
	LUT2 #(
		.INIT('h7)
	) name4754 (
		_w6899_,
		_w6900_,
		_w6901_
	);
	LUT4 #(
		.INIT('hf35f)
	) name4755 (
		\u10_mem_reg[1][2]/P0001 ,
		\u10_mem_reg[2][2]/P0001 ,
		\u10_rp_reg[0]/P0001 ,
		\u10_rp_reg[1]/P0001 ,
		_w6902_
	);
	LUT4 #(
		.INIT('h3ff5)
	) name4756 (
		\u10_mem_reg[0][2]/P0001 ,
		\u10_mem_reg[3][2]/P0001 ,
		\u10_rp_reg[0]/P0001 ,
		\u10_rp_reg[1]/P0001 ,
		_w6903_
	);
	LUT2 #(
		.INIT('h7)
	) name4757 (
		_w6902_,
		_w6903_,
		_w6904_
	);
	LUT4 #(
		.INIT('hff35)
	) name4758 (
		\u9_mem_reg[0][8]/P0001 ,
		\u9_mem_reg[1][8]/P0001 ,
		\u9_rp_reg[0]/P0001 ,
		\u9_rp_reg[1]/P0001 ,
		_w6905_
	);
	LUT4 #(
		.INIT('h35ff)
	) name4759 (
		\u9_mem_reg[2][8]/P0001 ,
		\u9_mem_reg[3][8]/P0001 ,
		\u9_rp_reg[0]/P0001 ,
		\u9_rp_reg[1]/P0001 ,
		_w6906_
	);
	LUT2 #(
		.INIT('h7)
	) name4760 (
		_w6905_,
		_w6906_,
		_w6907_
	);
	LUT4 #(
		.INIT('hf35f)
	) name4761 (
		\u10_mem_reg[1][31]/P0001 ,
		\u10_mem_reg[2][31]/P0001 ,
		\u10_rp_reg[0]/P0001 ,
		\u10_rp_reg[1]/P0001 ,
		_w6908_
	);
	LUT4 #(
		.INIT('h3ff5)
	) name4762 (
		\u10_mem_reg[0][31]/P0001 ,
		\u10_mem_reg[3][31]/P0001 ,
		\u10_rp_reg[0]/P0001 ,
		\u10_rp_reg[1]/P0001 ,
		_w6909_
	);
	LUT2 #(
		.INIT('h7)
	) name4763 (
		_w6908_,
		_w6909_,
		_w6910_
	);
	LUT4 #(
		.INIT('hff35)
	) name4764 (
		\u9_mem_reg[0][9]/P0001 ,
		\u9_mem_reg[1][9]/P0001 ,
		\u9_rp_reg[0]/P0001 ,
		\u9_rp_reg[1]/P0001 ,
		_w6911_
	);
	LUT4 #(
		.INIT('h35ff)
	) name4765 (
		\u9_mem_reg[2][9]/P0001 ,
		\u9_mem_reg[3][9]/P0001 ,
		\u9_rp_reg[0]/P0001 ,
		\u9_rp_reg[1]/P0001 ,
		_w6912_
	);
	LUT2 #(
		.INIT('h7)
	) name4766 (
		_w6911_,
		_w6912_,
		_w6913_
	);
	LUT3 #(
		.INIT('h02)
	) name4767 (
		\u10_din_tmp1_reg[3]/P0001 ,
		\u13_icc_r_reg[10]/NET0131 ,
		\u13_icc_r_reg[11]/NET0131 ,
		_w6914_
	);
	LUT4 #(
		.INIT('h9dbf)
	) name4768 (
		\u13_icc_r_reg[10]/NET0131 ,
		\u13_icc_r_reg[11]/NET0131 ,
		\u1_slt4_reg[3]/P0001 ,
		\u1_slt4_reg[5]/P0001 ,
		_w6915_
	);
	LUT2 #(
		.INIT('hb)
	) name4769 (
		_w6914_,
		_w6915_,
		_w6916_
	);
	LUT2 #(
		.INIT('h8)
	) name4770 (
		_w2399_,
		_w6573_,
		_w6917_
	);
	LUT3 #(
		.INIT('h10)
	) name4771 (
		\u13_icc_r_reg[2]/NET0131 ,
		\u13_icc_r_reg[3]/NET0131 ,
		\u9_din_tmp1_reg[1]/P0001 ,
		_w6918_
	);
	LUT4 #(
		.INIT('h9dbf)
	) name4772 (
		\u13_icc_r_reg[2]/NET0131 ,
		\u13_icc_r_reg[3]/NET0131 ,
		\u1_slt3_reg[1]/P0001 ,
		\u1_slt3_reg[3]/P0001 ,
		_w6919_
	);
	LUT2 #(
		.INIT('hb)
	) name4773 (
		_w6918_,
		_w6919_,
		_w6920_
	);
	LUT3 #(
		.INIT('h10)
	) name4774 (
		\u13_icc_r_reg[2]/NET0131 ,
		\u13_icc_r_reg[3]/NET0131 ,
		\u9_din_tmp1_reg[2]/P0001 ,
		_w6921_
	);
	LUT4 #(
		.INIT('h9dbf)
	) name4775 (
		\u13_icc_r_reg[2]/NET0131 ,
		\u13_icc_r_reg[3]/NET0131 ,
		\u1_slt3_reg[2]/P0001 ,
		\u1_slt3_reg[4]/P0001 ,
		_w6922_
	);
	LUT2 #(
		.INIT('hb)
	) name4776 (
		_w6921_,
		_w6922_,
		_w6923_
	);
	LUT3 #(
		.INIT('h10)
	) name4777 (
		\u13_icc_r_reg[2]/NET0131 ,
		\u13_icc_r_reg[3]/NET0131 ,
		\u9_din_tmp1_reg[8]/P0001 ,
		_w6924_
	);
	LUT4 #(
		.INIT('h9bdf)
	) name4778 (
		\u13_icc_r_reg[2]/NET0131 ,
		\u13_icc_r_reg[3]/NET0131 ,
		\u1_slt3_reg[10]/P0001 ,
		\u1_slt3_reg[8]/P0001 ,
		_w6925_
	);
	LUT2 #(
		.INIT('hb)
	) name4779 (
		_w6924_,
		_w6925_,
		_w6926_
	);
	LUT3 #(
		.INIT('h20)
	) name4780 (
		\u13_icc_r_reg[2]/NET0131 ,
		\u13_icc_r_reg[3]/NET0131 ,
		\u1_slt3_reg[19]/P0001 ,
		_w6927_
	);
	LUT4 #(
		.INIT('haebf)
	) name4781 (
		\u13_icc_r_reg[2]/NET0131 ,
		\u13_icc_r_reg[3]/NET0131 ,
		\u1_slt3_reg[17]/P0001 ,
		\u1_slt3_reg[5]/P0001 ,
		_w6928_
	);
	LUT2 #(
		.INIT('hb)
	) name4782 (
		_w6927_,
		_w6928_,
		_w6929_
	);
	LUT3 #(
		.INIT('h20)
	) name4783 (
		\u13_icc_r_reg[2]/NET0131 ,
		\u13_icc_r_reg[3]/NET0131 ,
		\u1_slt3_reg[18]/P0001 ,
		_w6930_
	);
	LUT4 #(
		.INIT('haebf)
	) name4784 (
		\u13_icc_r_reg[2]/NET0131 ,
		\u13_icc_r_reg[3]/NET0131 ,
		\u1_slt3_reg[16]/P0001 ,
		\u1_slt3_reg[4]/P0001 ,
		_w6931_
	);
	LUT2 #(
		.INIT('hb)
	) name4785 (
		_w6930_,
		_w6931_,
		_w6932_
	);
	LUT3 #(
		.INIT('h10)
	) name4786 (
		\u13_icc_r_reg[2]/NET0131 ,
		\u13_icc_r_reg[3]/NET0131 ,
		\u9_din_tmp1_reg[15]/P0001 ,
		_w6933_
	);
	LUT4 #(
		.INIT('h9dbf)
	) name4787 (
		\u13_icc_r_reg[2]/NET0131 ,
		\u13_icc_r_reg[3]/NET0131 ,
		\u1_slt3_reg[15]/P0001 ,
		\u1_slt3_reg[17]/P0001 ,
		_w6934_
	);
	LUT2 #(
		.INIT('hb)
	) name4788 (
		_w6933_,
		_w6934_,
		_w6935_
	);
	LUT3 #(
		.INIT('h10)
	) name4789 (
		\u13_icc_r_reg[2]/NET0131 ,
		\u13_icc_r_reg[3]/NET0131 ,
		\u9_din_tmp1_reg[14]/P0001 ,
		_w6936_
	);
	LUT4 #(
		.INIT('h9dbf)
	) name4790 (
		\u13_icc_r_reg[2]/NET0131 ,
		\u13_icc_r_reg[3]/NET0131 ,
		\u1_slt3_reg[14]/P0001 ,
		\u1_slt3_reg[16]/P0001 ,
		_w6937_
	);
	LUT2 #(
		.INIT('hb)
	) name4791 (
		_w6936_,
		_w6937_,
		_w6938_
	);
	LUT3 #(
		.INIT('h10)
	) name4792 (
		\u13_icc_r_reg[2]/NET0131 ,
		\u13_icc_r_reg[3]/NET0131 ,
		\u9_din_tmp1_reg[13]/P0001 ,
		_w6939_
	);
	LUT4 #(
		.INIT('h9dbf)
	) name4793 (
		\u13_icc_r_reg[2]/NET0131 ,
		\u13_icc_r_reg[3]/NET0131 ,
		\u1_slt3_reg[13]/P0001 ,
		\u1_slt3_reg[15]/P0001 ,
		_w6940_
	);
	LUT2 #(
		.INIT('hb)
	) name4794 (
		_w6939_,
		_w6940_,
		_w6941_
	);
	LUT3 #(
		.INIT('h10)
	) name4795 (
		\u13_icc_r_reg[2]/NET0131 ,
		\u13_icc_r_reg[3]/NET0131 ,
		\u9_din_tmp1_reg[12]/P0001 ,
		_w6942_
	);
	LUT4 #(
		.INIT('h9dbf)
	) name4796 (
		\u13_icc_r_reg[2]/NET0131 ,
		\u13_icc_r_reg[3]/NET0131 ,
		\u1_slt3_reg[12]/P0001 ,
		\u1_slt3_reg[14]/P0001 ,
		_w6943_
	);
	LUT2 #(
		.INIT('hb)
	) name4797 (
		_w6942_,
		_w6943_,
		_w6944_
	);
	LUT3 #(
		.INIT('h10)
	) name4798 (
		\u13_icc_r_reg[2]/NET0131 ,
		\u13_icc_r_reg[3]/NET0131 ,
		\u9_din_tmp1_reg[11]/P0001 ,
		_w6945_
	);
	LUT4 #(
		.INIT('h9dbf)
	) name4799 (
		\u13_icc_r_reg[2]/NET0131 ,
		\u13_icc_r_reg[3]/NET0131 ,
		\u1_slt3_reg[11]/P0001 ,
		\u1_slt3_reg[13]/P0001 ,
		_w6946_
	);
	LUT2 #(
		.INIT('hb)
	) name4800 (
		_w6945_,
		_w6946_,
		_w6947_
	);
	LUT3 #(
		.INIT('h10)
	) name4801 (
		\u13_icc_r_reg[2]/NET0131 ,
		\u13_icc_r_reg[3]/NET0131 ,
		\u9_din_tmp1_reg[9]/P0001 ,
		_w6948_
	);
	LUT4 #(
		.INIT('h9bdf)
	) name4802 (
		\u13_icc_r_reg[2]/NET0131 ,
		\u13_icc_r_reg[3]/NET0131 ,
		\u1_slt3_reg[11]/P0001 ,
		\u1_slt3_reg[9]/P0001 ,
		_w6949_
	);
	LUT2 #(
		.INIT('hb)
	) name4803 (
		_w6948_,
		_w6949_,
		_w6950_
	);
	LUT3 #(
		.INIT('h10)
	) name4804 (
		\u13_icc_r_reg[2]/NET0131 ,
		\u13_icc_r_reg[3]/NET0131 ,
		\u9_din_tmp1_reg[3]/P0001 ,
		_w6951_
	);
	LUT4 #(
		.INIT('h9dbf)
	) name4805 (
		\u13_icc_r_reg[2]/NET0131 ,
		\u13_icc_r_reg[3]/NET0131 ,
		\u1_slt3_reg[3]/P0001 ,
		\u1_slt3_reg[5]/P0001 ,
		_w6952_
	);
	LUT2 #(
		.INIT('hb)
	) name4806 (
		_w6951_,
		_w6952_,
		_w6953_
	);
	LUT3 #(
		.INIT('h10)
	) name4807 (
		\u13_icc_r_reg[2]/NET0131 ,
		\u13_icc_r_reg[3]/NET0131 ,
		\u9_din_tmp1_reg[10]/P0001 ,
		_w6954_
	);
	LUT4 #(
		.INIT('h9dbf)
	) name4808 (
		\u13_icc_r_reg[2]/NET0131 ,
		\u13_icc_r_reg[3]/NET0131 ,
		\u1_slt3_reg[10]/P0001 ,
		\u1_slt3_reg[12]/P0001 ,
		_w6955_
	);
	LUT2 #(
		.INIT('hb)
	) name4809 (
		_w6954_,
		_w6955_,
		_w6956_
	);
	LUT3 #(
		.INIT('h02)
	) name4810 (
		\u11_din_tmp1_reg[11]/P0001 ,
		\u13_icc_r_reg[18]/NET0131 ,
		\u13_icc_r_reg[19]/NET0131 ,
		_w6957_
	);
	LUT4 #(
		.INIT('h9dbf)
	) name4811 (
		\u13_icc_r_reg[18]/NET0131 ,
		\u13_icc_r_reg[19]/NET0131 ,
		\u1_slt6_reg[11]/P0001 ,
		\u1_slt6_reg[13]/P0001 ,
		_w6958_
	);
	LUT2 #(
		.INIT('hb)
	) name4812 (
		_w6957_,
		_w6958_,
		_w6959_
	);
	LUT3 #(
		.INIT('h02)
	) name4813 (
		\u10_din_tmp1_reg[9]/P0001 ,
		\u13_icc_r_reg[10]/NET0131 ,
		\u13_icc_r_reg[11]/NET0131 ,
		_w6960_
	);
	LUT4 #(
		.INIT('h9bdf)
	) name4814 (
		\u13_icc_r_reg[10]/NET0131 ,
		\u13_icc_r_reg[11]/NET0131 ,
		\u1_slt4_reg[11]/P0001 ,
		\u1_slt4_reg[9]/P0001 ,
		_w6961_
	);
	LUT2 #(
		.INIT('hb)
	) name4815 (
		_w6960_,
		_w6961_,
		_w6962_
	);
	LUT3 #(
		.INIT('h10)
	) name4816 (
		\u13_icc_r_reg[2]/NET0131 ,
		\u13_icc_r_reg[3]/NET0131 ,
		\u9_din_tmp1_reg[6]/P0001 ,
		_w6963_
	);
	LUT4 #(
		.INIT('h9dbf)
	) name4817 (
		\u13_icc_r_reg[2]/NET0131 ,
		\u13_icc_r_reg[3]/NET0131 ,
		\u1_slt3_reg[6]/P0001 ,
		\u1_slt3_reg[8]/P0001 ,
		_w6964_
	);
	LUT2 #(
		.INIT('hb)
	) name4818 (
		_w6963_,
		_w6964_,
		_w6965_
	);
	LUT3 #(
		.INIT('h02)
	) name4819 (
		\u10_din_tmp1_reg[0]/P0001 ,
		\u13_icc_r_reg[10]/NET0131 ,
		\u13_icc_r_reg[11]/NET0131 ,
		_w6966_
	);
	LUT4 #(
		.INIT('h9dbf)
	) name4820 (
		\u13_icc_r_reg[10]/NET0131 ,
		\u13_icc_r_reg[11]/NET0131 ,
		\u1_slt4_reg[0]/P0001 ,
		\u1_slt4_reg[2]/P0001 ,
		_w6967_
	);
	LUT2 #(
		.INIT('hb)
	) name4821 (
		_w6966_,
		_w6967_,
		_w6968_
	);
	LUT3 #(
		.INIT('h02)
	) name4822 (
		\u10_din_tmp1_reg[10]/P0001 ,
		\u13_icc_r_reg[10]/NET0131 ,
		\u13_icc_r_reg[11]/NET0131 ,
		_w6969_
	);
	LUT4 #(
		.INIT('h9dbf)
	) name4823 (
		\u13_icc_r_reg[10]/NET0131 ,
		\u13_icc_r_reg[11]/NET0131 ,
		\u1_slt4_reg[10]/P0001 ,
		\u1_slt4_reg[12]/P0001 ,
		_w6970_
	);
	LUT2 #(
		.INIT('hb)
	) name4824 (
		_w6969_,
		_w6970_,
		_w6971_
	);
	LUT3 #(
		.INIT('h02)
	) name4825 (
		\u10_din_tmp1_reg[11]/P0001 ,
		\u13_icc_r_reg[10]/NET0131 ,
		\u13_icc_r_reg[11]/NET0131 ,
		_w6972_
	);
	LUT4 #(
		.INIT('h9dbf)
	) name4826 (
		\u13_icc_r_reg[10]/NET0131 ,
		\u13_icc_r_reg[11]/NET0131 ,
		\u1_slt4_reg[11]/P0001 ,
		\u1_slt4_reg[13]/P0001 ,
		_w6973_
	);
	LUT2 #(
		.INIT('hb)
	) name4827 (
		_w6972_,
		_w6973_,
		_w6974_
	);
	LUT3 #(
		.INIT('h02)
	) name4828 (
		\u10_din_tmp1_reg[12]/P0001 ,
		\u13_icc_r_reg[10]/NET0131 ,
		\u13_icc_r_reg[11]/NET0131 ,
		_w6975_
	);
	LUT4 #(
		.INIT('h9dbf)
	) name4829 (
		\u13_icc_r_reg[10]/NET0131 ,
		\u13_icc_r_reg[11]/NET0131 ,
		\u1_slt4_reg[12]/P0001 ,
		\u1_slt4_reg[14]/P0001 ,
		_w6976_
	);
	LUT2 #(
		.INIT('hb)
	) name4830 (
		_w6975_,
		_w6976_,
		_w6977_
	);
	LUT3 #(
		.INIT('h10)
	) name4831 (
		\u13_icc_r_reg[2]/NET0131 ,
		\u13_icc_r_reg[3]/NET0131 ,
		\u9_din_tmp1_reg[7]/P0001 ,
		_w6978_
	);
	LUT4 #(
		.INIT('h9dbf)
	) name4832 (
		\u13_icc_r_reg[2]/NET0131 ,
		\u13_icc_r_reg[3]/NET0131 ,
		\u1_slt3_reg[7]/P0001 ,
		\u1_slt3_reg[9]/P0001 ,
		_w6979_
	);
	LUT2 #(
		.INIT('hb)
	) name4833 (
		_w6978_,
		_w6979_,
		_w6980_
	);
	LUT3 #(
		.INIT('h02)
	) name4834 (
		\u10_din_tmp1_reg[13]/P0001 ,
		\u13_icc_r_reg[10]/NET0131 ,
		\u13_icc_r_reg[11]/NET0131 ,
		_w6981_
	);
	LUT4 #(
		.INIT('h9dbf)
	) name4835 (
		\u13_icc_r_reg[10]/NET0131 ,
		\u13_icc_r_reg[11]/NET0131 ,
		\u1_slt4_reg[13]/P0001 ,
		\u1_slt4_reg[15]/P0001 ,
		_w6982_
	);
	LUT2 #(
		.INIT('hb)
	) name4836 (
		_w6981_,
		_w6982_,
		_w6983_
	);
	LUT3 #(
		.INIT('h10)
	) name4837 (
		\u13_icc_r_reg[2]/NET0131 ,
		\u13_icc_r_reg[3]/NET0131 ,
		\u9_din_tmp1_reg[5]/P0001 ,
		_w6984_
	);
	LUT4 #(
		.INIT('h9dbf)
	) name4838 (
		\u13_icc_r_reg[2]/NET0131 ,
		\u13_icc_r_reg[3]/NET0131 ,
		\u1_slt3_reg[5]/P0001 ,
		\u1_slt3_reg[7]/P0001 ,
		_w6985_
	);
	LUT2 #(
		.INIT('hb)
	) name4839 (
		_w6984_,
		_w6985_,
		_w6986_
	);
	LUT3 #(
		.INIT('h02)
	) name4840 (
		\u11_din_tmp1_reg[0]/P0001 ,
		\u13_icc_r_reg[18]/NET0131 ,
		\u13_icc_r_reg[19]/NET0131 ,
		_w6987_
	);
	LUT4 #(
		.INIT('h9dbf)
	) name4841 (
		\u13_icc_r_reg[18]/NET0131 ,
		\u13_icc_r_reg[19]/NET0131 ,
		\u1_slt6_reg[0]/P0001 ,
		\u1_slt6_reg[2]/P0001 ,
		_w6988_
	);
	LUT2 #(
		.INIT('hb)
	) name4842 (
		_w6987_,
		_w6988_,
		_w6989_
	);
	LUT3 #(
		.INIT('h02)
	) name4843 (
		\u11_din_tmp1_reg[10]/P0001 ,
		\u13_icc_r_reg[18]/NET0131 ,
		\u13_icc_r_reg[19]/NET0131 ,
		_w6990_
	);
	LUT4 #(
		.INIT('h9dbf)
	) name4844 (
		\u13_icc_r_reg[18]/NET0131 ,
		\u13_icc_r_reg[19]/NET0131 ,
		\u1_slt6_reg[10]/P0001 ,
		\u1_slt6_reg[12]/P0001 ,
		_w6991_
	);
	LUT2 #(
		.INIT('hb)
	) name4845 (
		_w6990_,
		_w6991_,
		_w6992_
	);
	LUT3 #(
		.INIT('h02)
	) name4846 (
		\u10_din_tmp1_reg[15]/P0001 ,
		\u13_icc_r_reg[10]/NET0131 ,
		\u13_icc_r_reg[11]/NET0131 ,
		_w6993_
	);
	LUT4 #(
		.INIT('h9dbf)
	) name4847 (
		\u13_icc_r_reg[10]/NET0131 ,
		\u13_icc_r_reg[11]/NET0131 ,
		\u1_slt4_reg[15]/P0001 ,
		\u1_slt4_reg[17]/P0001 ,
		_w6994_
	);
	LUT2 #(
		.INIT('hb)
	) name4848 (
		_w6993_,
		_w6994_,
		_w6995_
	);
	LUT3 #(
		.INIT('h02)
	) name4849 (
		\u11_din_tmp1_reg[12]/P0001 ,
		\u13_icc_r_reg[18]/NET0131 ,
		\u13_icc_r_reg[19]/NET0131 ,
		_w6996_
	);
	LUT4 #(
		.INIT('h9dbf)
	) name4850 (
		\u13_icc_r_reg[18]/NET0131 ,
		\u13_icc_r_reg[19]/NET0131 ,
		\u1_slt6_reg[12]/P0001 ,
		\u1_slt6_reg[14]/P0001 ,
		_w6997_
	);
	LUT2 #(
		.INIT('hb)
	) name4851 (
		_w6996_,
		_w6997_,
		_w6998_
	);
	LUT3 #(
		.INIT('h02)
	) name4852 (
		\u11_din_tmp1_reg[13]/P0001 ,
		\u13_icc_r_reg[18]/NET0131 ,
		\u13_icc_r_reg[19]/NET0131 ,
		_w6999_
	);
	LUT4 #(
		.INIT('h9dbf)
	) name4853 (
		\u13_icc_r_reg[18]/NET0131 ,
		\u13_icc_r_reg[19]/NET0131 ,
		\u1_slt6_reg[13]/P0001 ,
		\u1_slt6_reg[15]/P0001 ,
		_w7000_
	);
	LUT2 #(
		.INIT('hb)
	) name4854 (
		_w6999_,
		_w7000_,
		_w7001_
	);
	LUT3 #(
		.INIT('h40)
	) name4855 (
		\u13_icc_r_reg[10]/NET0131 ,
		\u13_icc_r_reg[11]/NET0131 ,
		\u1_slt4_reg[16]/P0001 ,
		_w7002_
	);
	LUT4 #(
		.INIT('hcedf)
	) name4856 (
		\u13_icc_r_reg[10]/NET0131 ,
		\u13_icc_r_reg[11]/NET0131 ,
		\u1_slt4_reg[18]/P0001 ,
		\u1_slt4_reg[4]/P0001 ,
		_w7003_
	);
	LUT2 #(
		.INIT('hb)
	) name4857 (
		_w7002_,
		_w7003_,
		_w7004_
	);
	LUT3 #(
		.INIT('h02)
	) name4858 (
		\u11_din_tmp1_reg[14]/P0001 ,
		\u13_icc_r_reg[18]/NET0131 ,
		\u13_icc_r_reg[19]/NET0131 ,
		_w7005_
	);
	LUT4 #(
		.INIT('h9dbf)
	) name4859 (
		\u13_icc_r_reg[18]/NET0131 ,
		\u13_icc_r_reg[19]/NET0131 ,
		\u1_slt6_reg[14]/P0001 ,
		\u1_slt6_reg[16]/P0001 ,
		_w7006_
	);
	LUT2 #(
		.INIT('hb)
	) name4860 (
		_w7005_,
		_w7006_,
		_w7007_
	);
	LUT3 #(
		.INIT('h40)
	) name4861 (
		\u13_icc_r_reg[10]/NET0131 ,
		\u13_icc_r_reg[11]/NET0131 ,
		\u1_slt4_reg[17]/P0001 ,
		_w7008_
	);
	LUT4 #(
		.INIT('hcedf)
	) name4862 (
		\u13_icc_r_reg[10]/NET0131 ,
		\u13_icc_r_reg[11]/NET0131 ,
		\u1_slt4_reg[19]/P0001 ,
		\u1_slt4_reg[5]/P0001 ,
		_w7009_
	);
	LUT2 #(
		.INIT('hb)
	) name4863 (
		_w7008_,
		_w7009_,
		_w7010_
	);
	LUT3 #(
		.INIT('h40)
	) name4864 (
		\u13_icc_r_reg[18]/NET0131 ,
		\u13_icc_r_reg[19]/NET0131 ,
		\u1_slt6_reg[17]/P0001 ,
		_w7011_
	);
	LUT4 #(
		.INIT('hcedf)
	) name4865 (
		\u13_icc_r_reg[18]/NET0131 ,
		\u13_icc_r_reg[19]/NET0131 ,
		\u1_slt6_reg[19]/P0001 ,
		\u1_slt6_reg[5]/P0001 ,
		_w7012_
	);
	LUT2 #(
		.INIT('hb)
	) name4866 (
		_w7011_,
		_w7012_,
		_w7013_
	);
	LUT3 #(
		.INIT('h02)
	) name4867 (
		\u11_din_tmp1_reg[1]/P0001 ,
		\u13_icc_r_reg[18]/NET0131 ,
		\u13_icc_r_reg[19]/NET0131 ,
		_w7014_
	);
	LUT4 #(
		.INIT('h9dbf)
	) name4868 (
		\u13_icc_r_reg[18]/NET0131 ,
		\u13_icc_r_reg[19]/NET0131 ,
		\u1_slt6_reg[1]/P0001 ,
		\u1_slt6_reg[3]/P0001 ,
		_w7015_
	);
	LUT2 #(
		.INIT('hb)
	) name4869 (
		_w7014_,
		_w7015_,
		_w7016_
	);
	LUT3 #(
		.INIT('h02)
	) name4870 (
		\u10_din_tmp1_reg[1]/P0001 ,
		\u13_icc_r_reg[10]/NET0131 ,
		\u13_icc_r_reg[11]/NET0131 ,
		_w7017_
	);
	LUT4 #(
		.INIT('h9dbf)
	) name4871 (
		\u13_icc_r_reg[10]/NET0131 ,
		\u13_icc_r_reg[11]/NET0131 ,
		\u1_slt4_reg[1]/P0001 ,
		\u1_slt4_reg[3]/P0001 ,
		_w7018_
	);
	LUT2 #(
		.INIT('hb)
	) name4872 (
		_w7017_,
		_w7018_,
		_w7019_
	);
	LUT3 #(
		.INIT('h02)
	) name4873 (
		\u10_din_tmp1_reg[14]/P0001 ,
		\u13_icc_r_reg[10]/NET0131 ,
		\u13_icc_r_reg[11]/NET0131 ,
		_w7020_
	);
	LUT4 #(
		.INIT('h9dbf)
	) name4874 (
		\u13_icc_r_reg[10]/NET0131 ,
		\u13_icc_r_reg[11]/NET0131 ,
		\u1_slt4_reg[14]/P0001 ,
		\u1_slt4_reg[16]/P0001 ,
		_w7021_
	);
	LUT2 #(
		.INIT('hb)
	) name4875 (
		_w7020_,
		_w7021_,
		_w7022_
	);
	LUT3 #(
		.INIT('h02)
	) name4876 (
		\u11_din_tmp1_reg[2]/P0001 ,
		\u13_icc_r_reg[18]/NET0131 ,
		\u13_icc_r_reg[19]/NET0131 ,
		_w7023_
	);
	LUT4 #(
		.INIT('h9dbf)
	) name4877 (
		\u13_icc_r_reg[18]/NET0131 ,
		\u13_icc_r_reg[19]/NET0131 ,
		\u1_slt6_reg[2]/P0001 ,
		\u1_slt6_reg[4]/P0001 ,
		_w7024_
	);
	LUT2 #(
		.INIT('hb)
	) name4878 (
		_w7023_,
		_w7024_,
		_w7025_
	);
	LUT3 #(
		.INIT('h40)
	) name4879 (
		\u13_icc_r_reg[18]/NET0131 ,
		\u13_icc_r_reg[19]/NET0131 ,
		\u1_slt6_reg[16]/P0001 ,
		_w7026_
	);
	LUT4 #(
		.INIT('hcedf)
	) name4880 (
		\u13_icc_r_reg[18]/NET0131 ,
		\u13_icc_r_reg[19]/NET0131 ,
		\u1_slt6_reg[18]/P0001 ,
		\u1_slt6_reg[4]/P0001 ,
		_w7027_
	);
	LUT2 #(
		.INIT('hb)
	) name4881 (
		_w7026_,
		_w7027_,
		_w7028_
	);
	LUT3 #(
		.INIT('h02)
	) name4882 (
		\u11_din_tmp1_reg[3]/P0001 ,
		\u13_icc_r_reg[18]/NET0131 ,
		\u13_icc_r_reg[19]/NET0131 ,
		_w7029_
	);
	LUT4 #(
		.INIT('h9dbf)
	) name4883 (
		\u13_icc_r_reg[18]/NET0131 ,
		\u13_icc_r_reg[19]/NET0131 ,
		\u1_slt6_reg[3]/P0001 ,
		\u1_slt6_reg[5]/P0001 ,
		_w7030_
	);
	LUT2 #(
		.INIT('hb)
	) name4884 (
		_w7029_,
		_w7030_,
		_w7031_
	);
	LUT3 #(
		.INIT('h02)
	) name4885 (
		\u11_din_tmp1_reg[4]/P0001 ,
		\u13_icc_r_reg[18]/NET0131 ,
		\u13_icc_r_reg[19]/NET0131 ,
		_w7032_
	);
	LUT4 #(
		.INIT('h9dbf)
	) name4886 (
		\u13_icc_r_reg[18]/NET0131 ,
		\u13_icc_r_reg[19]/NET0131 ,
		\u1_slt6_reg[4]/P0001 ,
		\u1_slt6_reg[6]/P0001 ,
		_w7033_
	);
	LUT2 #(
		.INIT('hb)
	) name4887 (
		_w7032_,
		_w7033_,
		_w7034_
	);
	LUT3 #(
		.INIT('h02)
	) name4888 (
		\u11_din_tmp1_reg[5]/P0001 ,
		\u13_icc_r_reg[18]/NET0131 ,
		\u13_icc_r_reg[19]/NET0131 ,
		_w7035_
	);
	LUT4 #(
		.INIT('h9dbf)
	) name4889 (
		\u13_icc_r_reg[18]/NET0131 ,
		\u13_icc_r_reg[19]/NET0131 ,
		\u1_slt6_reg[5]/P0001 ,
		\u1_slt6_reg[7]/P0001 ,
		_w7036_
	);
	LUT2 #(
		.INIT('hb)
	) name4890 (
		_w7035_,
		_w7036_,
		_w7037_
	);
	LUT3 #(
		.INIT('h02)
	) name4891 (
		\u11_din_tmp1_reg[6]/P0001 ,
		\u13_icc_r_reg[18]/NET0131 ,
		\u13_icc_r_reg[19]/NET0131 ,
		_w7038_
	);
	LUT4 #(
		.INIT('h9dbf)
	) name4892 (
		\u13_icc_r_reg[18]/NET0131 ,
		\u13_icc_r_reg[19]/NET0131 ,
		\u1_slt6_reg[6]/P0001 ,
		\u1_slt6_reg[8]/P0001 ,
		_w7039_
	);
	LUT2 #(
		.INIT('hb)
	) name4893 (
		_w7038_,
		_w7039_,
		_w7040_
	);
	LUT3 #(
		.INIT('h02)
	) name4894 (
		\u11_din_tmp1_reg[7]/P0001 ,
		\u13_icc_r_reg[18]/NET0131 ,
		\u13_icc_r_reg[19]/NET0131 ,
		_w7041_
	);
	LUT4 #(
		.INIT('h9dbf)
	) name4895 (
		\u13_icc_r_reg[18]/NET0131 ,
		\u13_icc_r_reg[19]/NET0131 ,
		\u1_slt6_reg[7]/P0001 ,
		\u1_slt6_reg[9]/P0001 ,
		_w7042_
	);
	LUT2 #(
		.INIT('hb)
	) name4896 (
		_w7041_,
		_w7042_,
		_w7043_
	);
	LUT3 #(
		.INIT('h02)
	) name4897 (
		\u11_din_tmp1_reg[8]/P0001 ,
		\u13_icc_r_reg[18]/NET0131 ,
		\u13_icc_r_reg[19]/NET0131 ,
		_w7044_
	);
	LUT4 #(
		.INIT('h9bdf)
	) name4898 (
		\u13_icc_r_reg[18]/NET0131 ,
		\u13_icc_r_reg[19]/NET0131 ,
		\u1_slt6_reg[10]/P0001 ,
		\u1_slt6_reg[8]/P0001 ,
		_w7045_
	);
	LUT2 #(
		.INIT('hb)
	) name4899 (
		_w7044_,
		_w7045_,
		_w7046_
	);
	LUT3 #(
		.INIT('h02)
	) name4900 (
		\u11_din_tmp1_reg[9]/P0001 ,
		\u13_icc_r_reg[18]/NET0131 ,
		\u13_icc_r_reg[19]/NET0131 ,
		_w7047_
	);
	LUT4 #(
		.INIT('h9bdf)
	) name4901 (
		\u13_icc_r_reg[18]/NET0131 ,
		\u13_icc_r_reg[19]/NET0131 ,
		\u1_slt6_reg[11]/P0001 ,
		\u1_slt6_reg[9]/P0001 ,
		_w7048_
	);
	LUT2 #(
		.INIT('hb)
	) name4902 (
		_w7047_,
		_w7048_,
		_w7049_
	);
	LUT3 #(
		.INIT('h02)
	) name4903 (
		\u10_din_tmp1_reg[2]/P0001 ,
		\u13_icc_r_reg[10]/NET0131 ,
		\u13_icc_r_reg[11]/NET0131 ,
		_w7050_
	);
	LUT4 #(
		.INIT('h9dbf)
	) name4904 (
		\u13_icc_r_reg[10]/NET0131 ,
		\u13_icc_r_reg[11]/NET0131 ,
		\u1_slt4_reg[2]/P0001 ,
		\u1_slt4_reg[4]/P0001 ,
		_w7051_
	);
	LUT2 #(
		.INIT('hb)
	) name4905 (
		_w7050_,
		_w7051_,
		_w7052_
	);
	LUT3 #(
		.INIT('h02)
	) name4906 (
		\u10_din_tmp1_reg[4]/P0001 ,
		\u13_icc_r_reg[10]/NET0131 ,
		\u13_icc_r_reg[11]/NET0131 ,
		_w7053_
	);
	LUT4 #(
		.INIT('h9dbf)
	) name4907 (
		\u13_icc_r_reg[10]/NET0131 ,
		\u13_icc_r_reg[11]/NET0131 ,
		\u1_slt4_reg[4]/P0001 ,
		\u1_slt4_reg[6]/P0001 ,
		_w7054_
	);
	LUT2 #(
		.INIT('hb)
	) name4908 (
		_w7053_,
		_w7054_,
		_w7055_
	);
	LUT3 #(
		.INIT('h02)
	) name4909 (
		\u10_din_tmp1_reg[5]/P0001 ,
		\u13_icc_r_reg[10]/NET0131 ,
		\u13_icc_r_reg[11]/NET0131 ,
		_w7056_
	);
	LUT4 #(
		.INIT('h9dbf)
	) name4910 (
		\u13_icc_r_reg[10]/NET0131 ,
		\u13_icc_r_reg[11]/NET0131 ,
		\u1_slt4_reg[5]/P0001 ,
		\u1_slt4_reg[7]/P0001 ,
		_w7057_
	);
	LUT2 #(
		.INIT('hb)
	) name4911 (
		_w7056_,
		_w7057_,
		_w7058_
	);
	LUT3 #(
		.INIT('h02)
	) name4912 (
		\u10_din_tmp1_reg[6]/P0001 ,
		\u13_icc_r_reg[10]/NET0131 ,
		\u13_icc_r_reg[11]/NET0131 ,
		_w7059_
	);
	LUT4 #(
		.INIT('h9dbf)
	) name4913 (
		\u13_icc_r_reg[10]/NET0131 ,
		\u13_icc_r_reg[11]/NET0131 ,
		\u1_slt4_reg[6]/P0001 ,
		\u1_slt4_reg[8]/P0001 ,
		_w7060_
	);
	LUT2 #(
		.INIT('hb)
	) name4914 (
		_w7059_,
		_w7060_,
		_w7061_
	);
	LUT3 #(
		.INIT('h02)
	) name4915 (
		\u10_din_tmp1_reg[7]/P0001 ,
		\u13_icc_r_reg[10]/NET0131 ,
		\u13_icc_r_reg[11]/NET0131 ,
		_w7062_
	);
	LUT4 #(
		.INIT('h9dbf)
	) name4916 (
		\u13_icc_r_reg[10]/NET0131 ,
		\u13_icc_r_reg[11]/NET0131 ,
		\u1_slt4_reg[7]/P0001 ,
		\u1_slt4_reg[9]/P0001 ,
		_w7063_
	);
	LUT2 #(
		.INIT('hb)
	) name4917 (
		_w7062_,
		_w7063_,
		_w7064_
	);
	LUT3 #(
		.INIT('h02)
	) name4918 (
		\u10_din_tmp1_reg[8]/P0001 ,
		\u13_icc_r_reg[10]/NET0131 ,
		\u13_icc_r_reg[11]/NET0131 ,
		_w7065_
	);
	LUT4 #(
		.INIT('h9bdf)
	) name4919 (
		\u13_icc_r_reg[10]/NET0131 ,
		\u13_icc_r_reg[11]/NET0131 ,
		\u1_slt4_reg[10]/P0001 ,
		\u1_slt4_reg[8]/P0001 ,
		_w7066_
	);
	LUT2 #(
		.INIT('hb)
	) name4920 (
		_w7065_,
		_w7066_,
		_w7067_
	);
	LUT3 #(
		.INIT('h02)
	) name4921 (
		\u11_din_tmp1_reg[15]/P0001 ,
		\u13_icc_r_reg[18]/NET0131 ,
		\u13_icc_r_reg[19]/NET0131 ,
		_w7068_
	);
	LUT4 #(
		.INIT('h9dbf)
	) name4922 (
		\u13_icc_r_reg[18]/NET0131 ,
		\u13_icc_r_reg[19]/NET0131 ,
		\u1_slt6_reg[15]/P0001 ,
		\u1_slt6_reg[17]/P0001 ,
		_w7069_
	);
	LUT2 #(
		.INIT('hb)
	) name4923 (
		_w7068_,
		_w7069_,
		_w7070_
	);
	LUT3 #(
		.INIT('h10)
	) name4924 (
		\u13_icc_r_reg[2]/NET0131 ,
		\u13_icc_r_reg[3]/NET0131 ,
		\u9_din_tmp1_reg[0]/P0001 ,
		_w7071_
	);
	LUT4 #(
		.INIT('h9dbf)
	) name4925 (
		\u13_icc_r_reg[2]/NET0131 ,
		\u13_icc_r_reg[3]/NET0131 ,
		\u1_slt3_reg[0]/P0001 ,
		\u1_slt3_reg[2]/P0001 ,
		_w7072_
	);
	LUT2 #(
		.INIT('hb)
	) name4926 (
		_w7071_,
		_w7072_,
		_w7073_
	);
	LUT3 #(
		.INIT('h10)
	) name4927 (
		\u13_icc_r_reg[2]/NET0131 ,
		\u13_icc_r_reg[3]/NET0131 ,
		\u9_din_tmp1_reg[4]/P0001 ,
		_w7074_
	);
	LUT4 #(
		.INIT('h9dbf)
	) name4928 (
		\u13_icc_r_reg[2]/NET0131 ,
		\u13_icc_r_reg[3]/NET0131 ,
		\u1_slt3_reg[4]/P0001 ,
		\u1_slt3_reg[6]/P0001 ,
		_w7075_
	);
	LUT2 #(
		.INIT('hb)
	) name4929 (
		_w7074_,
		_w7075_,
		_w7076_
	);
	LUT2 #(
		.INIT('h2)
	) name4930 (
		\u2_cnt_reg[0]/NET0131 ,
		\u2_cnt_reg[5]/NET0131 ,
		_w7077_
	);
	LUT3 #(
		.INIT('h80)
	) name4931 (
		_w6605_,
		_w6624_,
		_w7077_,
		_w7078_
	);
	LUT3 #(
		.INIT('he2)
	) name4932 (
		\u11_mem_reg[0][24]/P0001 ,
		_w4050_,
		_w4074_,
		_w7079_
	);
	LUT3 #(
		.INIT('hca)
	) name4933 (
		\u10_mem_reg[0][20]/P0001 ,
		_w3889_,
		_w4045_,
		_w7080_
	);
	LUT3 #(
		.INIT('he2)
	) name4934 (
		\u9_mem_reg[0][31]/P0001 ,
		_w3904_,
		_w3963_,
		_w7081_
	);
	LUT3 #(
		.INIT('he2)
	) name4935 (
		\u9_mem_reg[0][20]/P0001 ,
		_w3904_,
		_w3937_,
		_w7082_
	);
	LUT3 #(
		.INIT('he2)
	) name4936 (
		\u9_mem_reg[0][21]/P0001 ,
		_w3904_,
		_w3939_,
		_w7083_
	);
	LUT3 #(
		.INIT('he2)
	) name4937 (
		\u9_mem_reg[0][23]/P0001 ,
		_w3904_,
		_w3947_,
		_w7084_
	);
	LUT3 #(
		.INIT('he2)
	) name4938 (
		\u9_mem_reg[0][24]/P0001 ,
		_w3904_,
		_w3949_,
		_w7085_
	);
	LUT3 #(
		.INIT('he2)
	) name4939 (
		\u9_mem_reg[0][25]/P0001 ,
		_w3904_,
		_w3951_,
		_w7086_
	);
	LUT3 #(
		.INIT('he2)
	) name4940 (
		\u9_mem_reg[0][26]/P0001 ,
		_w3904_,
		_w3953_,
		_w7087_
	);
	LUT3 #(
		.INIT('he2)
	) name4941 (
		\u9_mem_reg[0][27]/P0001 ,
		_w3904_,
		_w3955_,
		_w7088_
	);
	LUT3 #(
		.INIT('he2)
	) name4942 (
		\u9_mem_reg[0][28]/P0001 ,
		_w3904_,
		_w3957_,
		_w7089_
	);
	LUT3 #(
		.INIT('he2)
	) name4943 (
		\u9_mem_reg[0][29]/P0001 ,
		_w3904_,
		_w3959_,
		_w7090_
	);
	LUT3 #(
		.INIT('he2)
	) name4944 (
		\u9_mem_reg[0][30]/P0001 ,
		_w3904_,
		_w3961_,
		_w7091_
	);
	LUT3 #(
		.INIT('he2)
	) name4945 (
		\u11_mem_reg[0][21]/P0001 ,
		_w4050_,
		_w4068_,
		_w7092_
	);
	LUT3 #(
		.INIT('hca)
	) name4946 (
		\u10_mem_reg[0][22]/P0001 ,
		_w3897_,
		_w4045_,
		_w7093_
	);
	LUT3 #(
		.INIT('he2)
	) name4947 (
		\u11_mem_reg[0][27]/P0001 ,
		_w4050_,
		_w4080_,
		_w7094_
	);
	LUT3 #(
		.INIT('he2)
	) name4948 (
		\u11_mem_reg[0][31]/P0001 ,
		_w4050_,
		_w4088_,
		_w7095_
	);
	LUT3 #(
		.INIT('he2)
	) name4949 (
		\u11_mem_reg[0][29]/P0001 ,
		_w4050_,
		_w4084_,
		_w7096_
	);
	LUT3 #(
		.INIT('he2)
	) name4950 (
		\u11_mem_reg[0][20]/P0001 ,
		_w4050_,
		_w4066_,
		_w7097_
	);
	LUT3 #(
		.INIT('he2)
	) name4951 (
		\u11_mem_reg[0][22]/P0001 ,
		_w4050_,
		_w4070_,
		_w7098_
	);
	LUT3 #(
		.INIT('he2)
	) name4952 (
		\u11_mem_reg[0][23]/P0001 ,
		_w4050_,
		_w4072_,
		_w7099_
	);
	LUT3 #(
		.INIT('he2)
	) name4953 (
		\u11_mem_reg[0][25]/P0001 ,
		_w4050_,
		_w4076_,
		_w7100_
	);
	LUT3 #(
		.INIT('hca)
	) name4954 (
		\u10_mem_reg[0][21]/P0001 ,
		_w3893_,
		_w4045_,
		_w7101_
	);
	LUT3 #(
		.INIT('he2)
	) name4955 (
		\u11_mem_reg[0][26]/P0001 ,
		_w4050_,
		_w4078_,
		_w7102_
	);
	LUT3 #(
		.INIT('hca)
	) name4956 (
		\u10_mem_reg[0][23]/P0001 ,
		_w3901_,
		_w4045_,
		_w7103_
	);
	LUT3 #(
		.INIT('he2)
	) name4957 (
		\u11_mem_reg[0][30]/P0001 ,
		_w4050_,
		_w4086_,
		_w7104_
	);
	LUT3 #(
		.INIT('hca)
	) name4958 (
		\u10_mem_reg[0][24]/P0001 ,
		_w3915_,
		_w4045_,
		_w7105_
	);
	LUT3 #(
		.INIT('hca)
	) name4959 (
		\u10_mem_reg[0][25]/P0001 ,
		_w3919_,
		_w4045_,
		_w7106_
	);
	LUT3 #(
		.INIT('hca)
	) name4960 (
		\u10_mem_reg[0][26]/P0001 ,
		_w3923_,
		_w4045_,
		_w7107_
	);
	LUT3 #(
		.INIT('hca)
	) name4961 (
		\u10_mem_reg[0][27]/P0001 ,
		_w3927_,
		_w4045_,
		_w7108_
	);
	LUT3 #(
		.INIT('hca)
	) name4962 (
		\u10_mem_reg[0][28]/P0001 ,
		_w3931_,
		_w4045_,
		_w7109_
	);
	LUT3 #(
		.INIT('he2)
	) name4963 (
		\u11_mem_reg[0][28]/P0001 ,
		_w4050_,
		_w4082_,
		_w7110_
	);
	LUT3 #(
		.INIT('hca)
	) name4964 (
		\u10_mem_reg[0][30]/P0001 ,
		_w3966_,
		_w4045_,
		_w7111_
	);
	LUT3 #(
		.INIT('hca)
	) name4965 (
		\u10_mem_reg[0][31]/P0001 ,
		_w3970_,
		_w4045_,
		_w7112_
	);
	LUT3 #(
		.INIT('hca)
	) name4966 (
		\u10_mem_reg[0][29]/P0001 ,
		_w3942_,
		_w4045_,
		_w7113_
	);
	LUT3 #(
		.INIT('he2)
	) name4967 (
		\u9_mem_reg[0][22]/P0001 ,
		_w3904_,
		_w3945_,
		_w7114_
	);
	LUT2 #(
		.INIT('h6)
	) name4968 (
		\u2_bit_clk_r1_reg/P0001 ,
		\u2_bit_clk_r_reg/P0001 ,
		_w7115_
	);
	LUT2 #(
		.INIT('h4)
	) name4969 (
		\dma_ack_i[6]_pad ,
		\dma_req_o[6]_pad ,
		_w7116_
	);
	LUT2 #(
		.INIT('h4)
	) name4970 (
		\dma_ack_i[6]_pad ,
		\u13_icc_r_reg[6]/NET0131 ,
		_w7117_
	);
	LUT4 #(
		.INIT('h8a00)
	) name4971 (
		\u13_icc_r_reg[0]/NET0131 ,
		_w3255_,
		_w3256_,
		_w7117_,
		_w7118_
	);
	LUT3 #(
		.INIT('hec)
	) name4972 (
		\u16_u6_dma_req_r1_reg/P0001 ,
		_w7116_,
		_w7118_,
		_w7119_
	);
	LUT2 #(
		.INIT('h4)
	) name4973 (
		\dma_ack_i[7]_pad ,
		\dma_req_o[7]_pad ,
		_w7120_
	);
	LUT2 #(
		.INIT('h4)
	) name4974 (
		\dma_ack_i[7]_pad ,
		\u13_icc_r_reg[14]/NET0131 ,
		_w7121_
	);
	LUT4 #(
		.INIT('h8a00)
	) name4975 (
		\u13_icc_r_reg[8]/NET0131 ,
		_w3271_,
		_w3272_,
		_w7121_,
		_w7122_
	);
	LUT3 #(
		.INIT('hec)
	) name4976 (
		\u16_u7_dma_req_r1_reg/P0001 ,
		_w7120_,
		_w7122_,
		_w7123_
	);
	LUT2 #(
		.INIT('he)
	) name4977 (
		\u2_sync_beat_reg/P0001 ,
		\u2_sync_resume_reg/NET0131 ,
		_w7124_
	);
	LUT3 #(
		.INIT('hac)
	) name4978 (
		\u14_u0_full_empty_r_reg/P0001 ,
		\u3_empty_reg/NET0131 ,
		\valid_s_reg/NET0131 ,
		_w7125_
	);
	LUT3 #(
		.INIT('hac)
	) name4979 (
		\u14_u1_full_empty_r_reg/P0001 ,
		\u4_empty_reg/NET0131 ,
		\valid_s_reg/NET0131 ,
		_w7126_
	);
	LUT3 #(
		.INIT('hac)
	) name4980 (
		\u14_u2_full_empty_r_reg/P0001 ,
		\u5_empty_reg/NET0131 ,
		\valid_s_reg/NET0131 ,
		_w7127_
	);
	LUT3 #(
		.INIT('hac)
	) name4981 (
		\u14_u3_full_empty_r_reg/P0001 ,
		\u6_empty_reg/NET0131 ,
		\valid_s_reg/NET0131 ,
		_w7128_
	);
	LUT3 #(
		.INIT('hac)
	) name4982 (
		\u14_u4_full_empty_r_reg/P0001 ,
		\u7_empty_reg/NET0131 ,
		\valid_s_reg/NET0131 ,
		_w7129_
	);
	LUT3 #(
		.INIT('hac)
	) name4983 (
		\u14_u5_full_empty_r_reg/P0001 ,
		\u8_empty_reg/NET0131 ,
		\valid_s_reg/NET0131 ,
		_w7130_
	);
	LUT3 #(
		.INIT('hd8)
	) name4984 (
		\in_valid_s_reg[0]/NET0131 ,
		\u14_u6_full_empty_r_reg/P0001 ,
		\u9_full_reg/NET0131 ,
		_w7131_
	);
	LUT3 #(
		.INIT('he4)
	) name4985 (
		\in_valid_s_reg[1]/NET0131 ,
		\u10_full_reg/NET0131 ,
		\u14_u7_full_empty_r_reg/P0001 ,
		_w7132_
	);
	LUT3 #(
		.INIT('he4)
	) name4986 (
		\in_valid_s_reg[2]/NET0131 ,
		\u11_full_reg/NET0131 ,
		\u14_u8_full_empty_r_reg/P0001 ,
		_w7133_
	);
	LUT3 #(
		.INIT('hca)
	) name4987 (
		\u1_slt0_reg[11]/P0001 ,
		\u1_sr_reg[11]/P0001 ,
		\u2_out_le_reg[0]/P0001 ,
		_w7134_
	);
	LUT3 #(
		.INIT('hca)
	) name4988 (
		\u1_slt0_reg[12]/P0001 ,
		\u1_sr_reg[12]/P0001 ,
		\u2_out_le_reg[0]/P0001 ,
		_w7135_
	);
	LUT3 #(
		.INIT('hca)
	) name4989 (
		\u1_slt0_reg[15]/P0001 ,
		\u1_sr_reg[15]/P0001 ,
		\u2_out_le_reg[0]/P0001 ,
		_w7136_
	);
	LUT3 #(
		.INIT('hca)
	) name4990 (
		\u1_slt0_reg[9]/P0001 ,
		\u1_sr_reg[9]/P0001 ,
		\u2_out_le_reg[0]/P0001 ,
		_w7137_
	);
	LUT3 #(
		.INIT('hca)
	) name4991 (
		\u1_slt1_reg[10]/P0001 ,
		\u1_sr_reg[10]/P0001 ,
		\u2_out_le_reg[1]/P0001 ,
		_w7138_
	);
	LUT3 #(
		.INIT('hca)
	) name4992 (
		\u1_slt1_reg[11]/P0001 ,
		\u1_sr_reg[11]/P0001 ,
		\u2_out_le_reg[1]/P0001 ,
		_w7139_
	);
	LUT3 #(
		.INIT('hca)
	) name4993 (
		\u1_slt1_reg[5]/P0001 ,
		\u1_sr_reg[5]/P0001 ,
		\u2_out_le_reg[1]/P0001 ,
		_w7140_
	);
	LUT3 #(
		.INIT('hca)
	) name4994 (
		\u1_slt1_reg[6]/P0001 ,
		\u1_sr_reg[6]/P0001 ,
		\u2_out_le_reg[1]/P0001 ,
		_w7141_
	);
	LUT3 #(
		.INIT('hca)
	) name4995 (
		\u1_slt1_reg[7]/P0001 ,
		\u1_sr_reg[7]/P0001 ,
		\u2_out_le_reg[1]/P0001 ,
		_w7142_
	);
	LUT3 #(
		.INIT('hca)
	) name4996 (
		\u1_slt1_reg[8]/P0001 ,
		\u1_sr_reg[8]/P0001 ,
		\u2_out_le_reg[1]/P0001 ,
		_w7143_
	);
	assign \_al_n1  = 1'b1;
	assign \g16/_0_  = _w2153_ ;
	assign \g23/_0_  = _w2160_ ;
	assign \g29500/_0_  = _w2165_ ;
	assign \g29503/_3_  = _w2166_ ;
	assign \g29505/_3_  = _w2167_ ;
	assign \g29507/_3_  = _w2168_ ;
	assign \g29509/_3_  = _w2169_ ;
	assign \g29511/_0_  = _w2170_ ;
	assign \g29513/_3_  = _w2171_ ;
	assign \g29515/_3_  = _w2172_ ;
	assign \g29517/_3_  = _w2173_ ;
	assign \g29519/_0_  = _w2174_ ;
	assign \g29522/_0_  = _w2175_ ;
	assign \g29524/_0_  = _w2176_ ;
	assign \g29526/_0_  = _w2177_ ;
	assign \g29528/_0_  = _w2178_ ;
	assign \g29530/_0_  = _w2179_ ;
	assign \g29532/_0_  = _w2180_ ;
	assign \g29534/_3_  = _w2181_ ;
	assign \g29536/_3_  = _w2182_ ;
	assign \g29538/_3_  = _w2183_ ;
	assign \g29540/_3_  = _w2184_ ;
	assign \g29542/_3_  = _w2185_ ;
	assign \g29544/_3_  = _w2186_ ;
	assign \g29546/_3_  = _w2187_ ;
	assign \g29548/_3_  = _w2188_ ;
	assign \g29550/_0_  = _w2189_ ;
	assign \g29552/_0_  = _w2190_ ;
	assign \g29554/_0_  = _w2191_ ;
	assign \g29556/_0_  = _w2192_ ;
	assign \g29558/_0_  = _w2193_ ;
	assign \g29560/_0_  = _w2194_ ;
	assign \g29562/_0_  = _w2195_ ;
	assign \g29564/_0_  = _w2196_ ;
	assign \g29566/_0_  = _w2197_ ;
	assign \g29568/_0_  = _w2198_ ;
	assign \g29570/_0_  = _w2199_ ;
	assign \g29572/_0_  = _w2200_ ;
	assign \g29574/_3_  = _w2201_ ;
	assign \g29576/_3_  = _w2202_ ;
	assign \g29578/_3_  = _w2203_ ;
	assign \g29580/_3_  = _w2204_ ;
	assign \g29582/_3_  = _w2205_ ;
	assign \g29584/_3_  = _w2206_ ;
	assign \g29586/_3_  = _w2207_ ;
	assign \g29588/_3_  = _w2208_ ;
	assign \g29590/_3_  = _w2209_ ;
	assign \g29592/_3_  = _w2210_ ;
	assign \g29594/_3_  = _w2211_ ;
	assign \g29596/_3_  = _w2212_ ;
	assign \g29598/_3_  = _w2213_ ;
	assign \g29600/_3_  = _w2214_ ;
	assign \g29602/_3_  = _w2215_ ;
	assign \g29604/_3_  = _w2216_ ;
	assign \g29606/_0_  = _w2217_ ;
	assign \g29608/_0_  = _w2218_ ;
	assign \g29610/_0_  = _w2219_ ;
	assign \g29612/_0_  = _w2220_ ;
	assign \g29614/_3_  = _w2221_ ;
	assign \g29616/_3_  = _w2222_ ;
	assign \g29618/_3_  = _w2223_ ;
	assign \g29620/_3_  = _w2224_ ;
	assign \g29622/_3_  = _w2225_ ;
	assign \g29624/_3_  = _w2226_ ;
	assign \g29626/_3_  = _w2227_ ;
	assign \g29628/_3_  = _w2228_ ;
	assign \g29630/_3_  = _w2229_ ;
	assign \g29632/_3_  = _w2230_ ;
	assign \g29634/_3_  = _w2231_ ;
	assign \g29636/_3_  = _w2232_ ;
	assign \g29638/_3_  = _w2233_ ;
	assign \g29640/_3_  = _w2234_ ;
	assign \g29642/_3_  = _w2235_ ;
	assign \g29644/_3_  = _w2236_ ;
	assign \g29646/_3_  = _w2237_ ;
	assign \g29648/_3_  = _w2238_ ;
	assign \g29650/_3_  = _w2239_ ;
	assign \g29652/_3_  = _w2240_ ;
	assign \g29654/_3_  = _w2241_ ;
	assign \g29656/_3_  = _w2242_ ;
	assign \g29658/_3_  = _w2243_ ;
	assign \g29660/_3_  = _w2244_ ;
	assign \g29662/_3_  = _w2245_ ;
	assign \g29664/_3_  = _w2246_ ;
	assign \g29666/_3_  = _w2247_ ;
	assign \g29668/_3_  = _w2248_ ;
	assign \g29670/_3_  = _w2249_ ;
	assign \g29672/_3_  = _w2250_ ;
	assign \g29674/_3_  = _w2251_ ;
	assign \g29676/_3_  = _w2252_ ;
	assign \g29678/_3_  = _w2253_ ;
	assign \g29680/_3_  = _w2254_ ;
	assign \g29682/_3_  = _w2255_ ;
	assign \g29684/_3_  = _w2256_ ;
	assign \g29686/_3_  = _w2257_ ;
	assign \g29688/_3_  = _w2258_ ;
	assign \g29690/_3_  = _w2259_ ;
	assign \g29692/_3_  = _w2260_ ;
	assign \g29694/_0_  = _w2261_ ;
	assign \g29696/_0_  = _w2262_ ;
	assign \g29698/_0_  = _w2263_ ;
	assign \g29700/_0_  = _w2264_ ;
	assign \g29702/_0_  = _w2265_ ;
	assign \g29704/_0_  = _w2266_ ;
	assign \g29706/_0_  = _w2267_ ;
	assign \g29708/_0_  = _w2268_ ;
	assign \g29710/_0_  = _w2269_ ;
	assign \g29712/_0_  = _w2270_ ;
	assign \g29714/_0_  = _w2271_ ;
	assign \g29716/_0_  = _w2272_ ;
	assign \g29718/_0_  = _w2273_ ;
	assign \g29720/_0_  = _w2274_ ;
	assign \g29722/_0_  = _w2275_ ;
	assign \g29724/_0_  = _w2276_ ;
	assign \g29726/_0_  = _w2277_ ;
	assign \g29728/_0_  = _w2278_ ;
	assign \g29730/_0_  = _w2279_ ;
	assign \g29732/_0_  = _w2280_ ;
	assign \g29734/_3_  = _w2281_ ;
	assign \g29736/_3_  = _w2282_ ;
	assign \g29738/_3_  = _w2283_ ;
	assign \g29740/_3_  = _w2284_ ;
	assign \g29742/_3_  = _w2285_ ;
	assign \g29744/_3_  = _w2286_ ;
	assign \g29746/_3_  = _w2287_ ;
	assign \g29748/_3_  = _w2288_ ;
	assign \g29750/_3_  = _w2289_ ;
	assign \g29752/_3_  = _w2290_ ;
	assign \g29754/_3_  = _w2291_ ;
	assign \g29756/_3_  = _w2292_ ;
	assign \g29758/_3_  = _w2293_ ;
	assign \g29760/_3_  = _w2294_ ;
	assign \g29762/_3_  = _w2295_ ;
	assign \g29764/_3_  = _w2296_ ;
	assign \g29766/_3_  = _w2297_ ;
	assign \g29768/_3_  = _w2298_ ;
	assign \g29770/_3_  = _w2299_ ;
	assign \g29772/_3_  = _w2300_ ;
	assign \g29774/_3_  = _w2301_ ;
	assign \g29776/_3_  = _w2302_ ;
	assign \g29778/_3_  = _w2303_ ;
	assign \g29780/_3_  = _w2304_ ;
	assign \g29782/_3_  = _w2305_ ;
	assign \g29784/_3_  = _w2306_ ;
	assign \g29786/_3_  = _w2307_ ;
	assign \g29788/_3_  = _w2308_ ;
	assign \g29790/_3_  = _w2309_ ;
	assign \g29792/_3_  = _w2310_ ;
	assign \g29794/_3_  = _w2311_ ;
	assign \g29796/_3_  = _w2312_ ;
	assign \g29798/_3_  = _w2313_ ;
	assign \g29800/_3_  = _w2314_ ;
	assign \g29802/_3_  = _w2315_ ;
	assign \g29804/_3_  = _w2316_ ;
	assign \g29806/_3_  = _w2317_ ;
	assign \g29808/_3_  = _w2318_ ;
	assign \g29810/_3_  = _w2319_ ;
	assign \g29812/_3_  = _w2320_ ;
	assign \g29814/_3_  = _w2321_ ;
	assign \g29816/_3_  = _w2322_ ;
	assign \g29818/_3_  = _w2323_ ;
	assign \g29820/_3_  = _w2324_ ;
	assign \g29822/_3_  = _w2325_ ;
	assign \g29824/_3_  = _w2326_ ;
	assign \g29826/_3_  = _w2327_ ;
	assign \g29828/_3_  = _w2328_ ;
	assign \g29830/_3_  = _w2329_ ;
	assign \g29832/_3_  = _w2330_ ;
	assign \g29834/_3_  = _w2331_ ;
	assign \g29836/_3_  = _w2332_ ;
	assign \g29838/_3_  = _w2333_ ;
	assign \g29840/_3_  = _w2334_ ;
	assign \g29842/_3_  = _w2335_ ;
	assign \g29844/_3_  = _w2336_ ;
	assign \g29846/_3_  = _w2337_ ;
	assign \g29848/_3_  = _w2338_ ;
	assign \g29850/_3_  = _w2339_ ;
	assign \g29852/_3_  = _w2340_ ;
	assign \g29854/_3_  = _w2341_ ;
	assign \g29856/_3_  = _w2342_ ;
	assign \g29858/_3_  = _w2343_ ;
	assign \g29860/_3_  = _w2344_ ;
	assign \g29862/_3_  = _w2345_ ;
	assign \g29864/_3_  = _w2346_ ;
	assign \g29866/_3_  = _w2347_ ;
	assign \g29868/_3_  = _w2348_ ;
	assign \g29870/_3_  = _w2349_ ;
	assign \g29872/_3_  = _w2350_ ;
	assign \g29874/_3_  = _w2351_ ;
	assign \g29876/_3_  = _w2352_ ;
	assign \g29878/_3_  = _w2353_ ;
	assign \g29880/_3_  = _w2354_ ;
	assign \g29904/_0_  = _w2361_ ;
	assign \g29905/_0_  = _w2368_ ;
	assign \g29906/_0_  = _w2375_ ;
	assign \g29907/_0_  = _w2382_ ;
	assign \g29908/_0_  = _w2389_ ;
	assign \g29909/_0_  = _w2396_ ;
	assign \g29914/_3_  = _w2397_ ;
	assign \g29952/_0_  = _w2404_ ;
	assign \g29953/_0_  = _w2406_ ;
	assign \g29954/_0_  = _w2408_ ;
	assign \g29955/_0_  = _w2410_ ;
	assign \g29956/_0_  = _w2412_ ;
	assign \g29957/_0_  = _w2414_ ;
	assign \g29975/_0_  = _w2360_ ;
	assign \g29976/_0_  = _w2367_ ;
	assign \g29977/_0_  = _w2374_ ;
	assign \g29978/_0_  = _w2381_ ;
	assign \g29979/_0_  = _w2388_ ;
	assign \g29980/_0_  = _w2395_ ;
	assign \g29989/_3_  = _w2415_ ;
	assign \g30020/_0_  = _w2424_ ;
	assign \g30021/_0_  = _w2433_ ;
	assign \g30045/_0_  = _w2436_ ;
	assign \g30046/_0_  = _w2442_ ;
	assign \g30047/_0_  = _w2451_ ;
	assign \g30048/_0_  = _w2458_ ;
	assign \g30049/_0_  = _w2358_ ;
	assign \g30050/_0_  = _w2365_ ;
	assign \g30051/_0_  = _w2372_ ;
	assign \g30052/_0_  = _w2379_ ;
	assign \g30053/_0_  = _w2386_ ;
	assign \g30054/_0_  = _w2393_ ;
	assign \g30062/_0_  = _w2459_ ;
	assign \g30063/_0_  = _w2460_ ;
	assign \g30064/_0_  = _w2462_ ;
	assign \g30065/_0_  = _w2464_ ;
	assign \g30066/_0_  = _w2466_ ;
	assign \g30067/_0_  = _w2467_ ;
	assign \g30068/_0_  = _w2468_ ;
	assign \g30069/_0_  = _w2469_ ;
	assign \g30070/_0_  = _w2470_ ;
	assign \g30071/_0_  = _w2471_ ;
	assign \g30072/_0_  = _w2472_ ;
	assign \g30073/_0_  = _w2473_ ;
	assign \g30074/_0_  = _w2474_ ;
	assign \g30075/_0_  = _w2475_ ;
	assign \g30136/_3_  = _w2476_ ;
	assign \g30707/_0_  = _w2479_ ;
	assign \g30708/_0_  = _w2480_ ;
	assign \g30711/_0_  = _w2481_ ;
	assign \g30714/_0_  = _w2482_ ;
	assign \g30715/_0_  = _w2483_ ;
	assign \g30720/_0_  = _w2484_ ;
	assign \g30725/_0_  = _w2485_ ;
	assign \g30741/_0_  = _w2493_ ;
	assign \g30742/_0_  = _w2498_ ;
	assign \g30743/_0_  = _w2506_ ;
	assign \g30744/_0_  = _w2511_ ;
	assign \g30745/_0_  = _w2519_ ;
	assign \g30746/_0_  = _w2524_ ;
	assign \g30747/_0_  = _w2532_ ;
	assign \g30748/_0_  = _w2537_ ;
	assign \g30749/_0_  = _w2545_ ;
	assign \g30750/_0_  = _w2553_ ;
	assign \g30751/_0_  = _w2558_ ;
	assign \g30752/_0_  = _w2563_ ;
	assign \g30789/_0_  = _w2571_ ;
	assign \g30790/_0_  = _w2589_ ;
	assign \g30791/_0_  = _w2606_ ;
	assign \g30792/_0_  = _w2619_ ;
	assign \g30793/_0_  = _w2632_ ;
	assign \g30794/_0_  = _w2645_ ;
	assign \g30795/_0_  = _w2658_ ;
	assign \g30796/_0_  = _w2671_ ;
	assign \g30797/_0_  = _w2684_ ;
	assign \g30798/_0_  = _w2692_ ;
	assign \g30799/_0_  = _w2705_ ;
	assign \g30800/_0_  = _w2718_ ;
	assign \g30801/_0_  = _w2725_ ;
	assign \g30802/_0_  = _w2732_ ;
	assign \g30803/_0_  = _w2742_ ;
	assign \g30804/_0_  = _w2752_ ;
	assign \g30805/_0_  = _w2760_ ;
	assign \g30806/_0_  = _w2768_ ;
	assign \g30807/_0_  = _w2779_ ;
	assign \g30808/_0_  = _w2790_ ;
	assign \g30809/_0_  = _w2798_ ;
	assign \g30810/_0_  = _w2816_ ;
	assign \g30811/_0_  = _w2833_ ;
	assign \g30812/_0_  = _w2846_ ;
	assign \g30813/_0_  = _w2859_ ;
	assign \g30814/_0_  = _w2872_ ;
	assign \g30815/_0_  = _w2885_ ;
	assign \g30816/_0_  = _w2898_ ;
	assign \g30817/_0_  = _w2911_ ;
	assign \g30818/_0_  = _w2924_ ;
	assign \g30819/_0_  = _w2937_ ;
	assign \g30820/_0_  = _w2944_ ;
	assign \g30821/_0_  = _w2951_ ;
	assign \g30822/_0_  = _w2961_ ;
	assign \g30823/_0_  = _w2971_ ;
	assign \g30824/_0_  = _w2979_ ;
	assign \g30825/_0_  = _w2987_ ;
	assign \g30826/_0_  = _w2998_ ;
	assign \g30827/_0_  = _w3009_ ;
	assign \g30828/_0_  = _w3027_ ;
	assign \g30829/_0_  = _w3044_ ;
	assign \g30830/_0_  = _w3057_ ;
	assign \g30831/_0_  = _w3070_ ;
	assign \g30832/_0_  = _w3083_ ;
	assign \g30833/_0_  = _w3096_ ;
	assign \g30834/_0_  = _w3109_ ;
	assign \g30835/_0_  = _w3122_ ;
	assign \g30836/_0_  = _w3135_ ;
	assign \g30837/_0_  = _w3148_ ;
	assign \g30838/_0_  = _w3155_ ;
	assign \g30839/_0_  = _w3162_ ;
	assign \g30840/_0_  = _w3172_ ;
	assign \g30841/_0_  = _w3182_ ;
	assign \g30842/_0_  = _w3190_ ;
	assign \g30843/_0_  = _w3198_ ;
	assign \g30844/_0_  = _w3209_ ;
	assign \g30845/_0_  = _w3220_ ;
	assign \g30846/_0_  = _w3238_ ;
	assign \g30847/_0_  = _w3254_ ;
	assign \g30848/_0_  = _w3257_ ;
	assign \g30849/_0_  = _w3270_ ;
	assign \g30850/_0_  = _w3273_ ;
	assign \g30851/_0_  = _w3286_ ;
	assign \g30852/_0_  = _w3299_ ;
	assign \g30853/_0_  = _w2150_ ;
	assign \g30854/_0_  = _w3311_ ;
	assign \g30855/_0_  = _w3324_ ;
	assign \g30856/_0_  = _w3337_ ;
	assign \g30857/_0_  = _w3350_ ;
	assign \g30858/_0_  = _w3363_ ;
	assign \g30859/_0_  = _w3370_ ;
	assign \g30860/_0_  = _w3377_ ;
	assign \g30861/_0_  = _w3387_ ;
	assign \g30862/_0_  = _w3397_ ;
	assign \g30863/_0_  = _w3405_ ;
	assign \g30864/_0_  = _w3413_ ;
	assign \g30865/_0_  = _w3424_ ;
	assign \g30866/_0_  = _w3435_ ;
	assign \g30867/_0_  = _w3453_ ;
	assign \g30868/_0_  = _w3470_ ;
	assign \g30869/_0_  = _w3483_ ;
	assign \g30870/_0_  = _w3495_ ;
	assign \g30871/_0_  = _w3508_ ;
	assign \g30872/_0_  = _w3521_ ;
	assign \g30873/_0_  = _w3534_ ;
	assign \g30874/_0_  = _w3546_ ;
	assign \g30875/_0_  = _w3559_ ;
	assign \g30876/_0_  = _w3577_ ;
	assign \g30877/_0_  = _w3590_ ;
	assign \g30878/_0_  = _w3607_ ;
	assign \g30879/_0_  = _w3620_ ;
	assign \g30880/_0_  = _w3627_ ;
	assign \g30881/_0_  = _w3640_ ;
	assign \g30882/_0_  = _w3647_ ;
	assign \g30883/_0_  = _w3660_ ;
	assign \g30884/_0_  = _w3670_ ;
	assign \g30885/_0_  = _w3683_ ;
	assign \g30886/_0_  = _w3693_ ;
	assign \g30887/_0_  = _w3706_ ;
	assign \g30888/_0_  = _w3719_ ;
	assign \g30889/_0_  = _w3727_ ;
	assign \g30890/_0_  = _w3735_ ;
	assign \g30891/_0_  = _w3748_ ;
	assign \g30892/_0_  = _w3759_ ;
	assign \g30893/_0_  = _w3772_ ;
	assign \g30894/_0_  = _w3783_ ;
	assign \g30895/_0_  = _w3790_ ;
	assign \g30896/_0_  = _w3797_ ;
	assign \g30897/_0_  = _w3807_ ;
	assign \g30898/_0_  = _w3817_ ;
	assign \g30899/_0_  = _w3825_ ;
	assign \g30900/_0_  = _w3833_ ;
	assign \g30901/_0_  = _w3844_ ;
	assign \g30902/_0_  = _w3855_ ;
	assign \g30906/_0_  = _w3856_ ;
	assign \g30907/_0_  = _w3857_ ;
	assign \g30908/_0_  = _w3858_ ;
	assign \g30909/_0_  = _w3859_ ;
	assign \g30910/_0_  = _w3860_ ;
	assign \g30911/_0_  = _w3861_ ;
	assign \g30918/_0_  = _w3865_ ;
	assign \g30919/_0_  = _w3866_ ;
	assign \g30920/_0_  = _w3868_ ;
	assign \g30921/_0_  = _w3871_ ;
	assign \g30922/_0_  = _w3873_ ;
	assign \g30923/_0_  = _w3874_ ;
	assign \g30924/_0_  = _w3875_ ;
	assign \g30925/_0_  = _w3876_ ;
	assign \g30926/_0_  = _w3877_ ;
	assign \g30946/_0_  = _w3883_ ;
	assign \g30947/_0_  = _w3887_ ;
	assign \g30948/_0_  = _w3891_ ;
	assign \g30949/_0_  = _w3895_ ;
	assign \g30950/_0_  = _w3899_ ;
	assign \g30951/_0_  = _w3903_ ;
	assign \g30952/_0_  = _w3909_ ;
	assign \g30953/_0_  = _w3913_ ;
	assign \g30954/_0_  = _w3917_ ;
	assign \g30955/_0_  = _w3921_ ;
	assign \g30956/_0_  = _w3925_ ;
	assign \g30957/_0_  = _w3929_ ;
	assign \g30958/_0_  = _w3933_ ;
	assign \g30959/_0_  = _w3935_ ;
	assign \g30960/_0_  = _w3936_ ;
	assign \g30961/_0_  = _w3938_ ;
	assign \g30962/_0_  = _w3940_ ;
	assign \g30963/_0_  = _w3944_ ;
	assign \g30964/_0_  = _w3946_ ;
	assign \g30965/_0_  = _w3948_ ;
	assign \g30966/_0_  = _w3950_ ;
	assign \g30967/_0_  = _w3952_ ;
	assign \g30968/_0_  = _w3954_ ;
	assign \g30969/_0_  = _w3956_ ;
	assign \g30970/_0_  = _w3958_ ;
	assign \g30971/_0_  = _w3960_ ;
	assign \g30972/_0_  = _w3962_ ;
	assign \g30973/_0_  = _w3964_ ;
	assign \g30974/_0_  = _w3968_ ;
	assign \g30975/_0_  = _w3972_ ;
	assign \g30976/_0_  = _w3977_ ;
	assign \g30977/_0_  = _w3980_ ;
	assign \g30978/_0_  = _w3983_ ;
	assign \g30979/_0_  = _w3986_ ;
	assign \g30980/_0_  = _w3989_ ;
	assign \g30981/_0_  = _w3992_ ;
	assign \g30982/_0_  = _w3995_ ;
	assign \g30983/_0_  = _w3998_ ;
	assign \g30984/_0_  = _w4001_ ;
	assign \g30985/_0_  = _w4004_ ;
	assign \g30986/_0_  = _w4007_ ;
	assign \g30987/_0_  = _w4010_ ;
	assign \g30988/_0_  = _w4013_ ;
	assign \g30989/_0_  = _w4016_ ;
	assign \g30990/_0_  = _w4017_ ;
	assign \g30991/_0_  = _w4018_ ;
	assign \g30992/_0_  = _w4019_ ;
	assign \g30993/_0_  = _w4020_ ;
	assign \g30994/_0_  = _w4021_ ;
	assign \g30995/_0_  = _w4022_ ;
	assign \g30996/_0_  = _w4023_ ;
	assign \g30997/_0_  = _w4024_ ;
	assign \g30998/_0_  = _w4025_ ;
	assign \g30999/_0_  = _w4026_ ;
	assign \g31000/_0_  = _w4027_ ;
	assign \g31001/_0_  = _w4028_ ;
	assign \g31002/_0_  = _w4029_ ;
	assign \g31003/_0_  = _w4030_ ;
	assign \g31004/_0_  = _w4031_ ;
	assign \g31005/_0_  = _w4032_ ;
	assign \g31006/_0_  = _w4033_ ;
	assign \g31007/_0_  = _w4034_ ;
	assign \g31008/_0_  = _w4035_ ;
	assign \g31009/_0_  = _w4036_ ;
	assign \g31010/_0_  = _w4037_ ;
	assign \g31011/_0_  = _w4038_ ;
	assign \g31012/_0_  = _w4039_ ;
	assign \g31013/_0_  = _w4040_ ;
	assign \g31014/_0_  = _w4041_ ;
	assign \g31015/_0_  = _w4042_ ;
	assign \g31016/_0_  = _w4043_ ;
	assign \g31017/_0_  = _w4044_ ;
	assign \g31018/_0_  = _w4049_ ;
	assign \g31019/_0_  = _w4055_ ;
	assign \g31020/_0_  = _w4059_ ;
	assign \g31021/_0_  = _w4062_ ;
	assign \g31022/_0_  = _w4064_ ;
	assign \g31023/_0_  = _w4065_ ;
	assign \g31024/_0_  = _w4067_ ;
	assign \g31025/_0_  = _w4069_ ;
	assign \g31026/_0_  = _w4071_ ;
	assign \g31027/_0_  = _w4073_ ;
	assign \g31028/_0_  = _w4075_ ;
	assign \g31029/_0_  = _w4077_ ;
	assign \g31030/_0_  = _w4079_ ;
	assign \g31031/_0_  = _w4081_ ;
	assign \g31032/_0_  = _w4083_ ;
	assign \g31033/_0_  = _w4085_ ;
	assign \g31034/_0_  = _w4087_ ;
	assign \g31035/_0_  = _w4089_ ;
	assign \g31036/_0_  = _w4094_ ;
	assign \g31037/_0_  = _w4097_ ;
	assign \g31038/_0_  = _w4100_ ;
	assign \g31039/_0_  = _w4103_ ;
	assign \g31040/_0_  = _w4106_ ;
	assign \g31041/_0_  = _w4109_ ;
	assign \g31042/_0_  = _w4112_ ;
	assign \g31043/_0_  = _w4115_ ;
	assign \g31044/_0_  = _w4117_ ;
	assign \g31045/_0_  = _w4120_ ;
	assign \g31046/_0_  = _w4123_ ;
	assign \g31047/_0_  = _w4124_ ;
	assign \g31048/_0_  = _w4127_ ;
	assign \g31049/_0_  = _w4130_ ;
	assign \g31050/_0_  = _w4133_ ;
	assign \g31051/_0_  = _w4134_ ;
	assign \g31052/_0_  = _w4137_ ;
	assign \g31053/_0_  = _w4138_ ;
	assign \g31054/_0_  = _w4139_ ;
	assign \g31055/_0_  = _w4140_ ;
	assign \g31056/_0_  = _w4141_ ;
	assign \g31057/_0_  = _w4142_ ;
	assign \g31058/_0_  = _w4143_ ;
	assign \g31059/_0_  = _w4144_ ;
	assign \g31060/_0_  = _w4145_ ;
	assign \g31061/_0_  = _w4146_ ;
	assign \g31062/_0_  = _w4147_ ;
	assign \g31063/_0_  = _w4148_ ;
	assign \g31064/_0_  = _w4149_ ;
	assign \g31065/_0_  = _w4150_ ;
	assign \g31066/_0_  = _w4151_ ;
	assign \g31067/_0_  = _w4152_ ;
	assign \g31068/_0_  = _w4153_ ;
	assign \g31069/_0_  = _w4154_ ;
	assign \g31070/_0_  = _w4155_ ;
	assign \g31071/_0_  = _w4156_ ;
	assign \g31072/_0_  = _w4157_ ;
	assign \g31073/_0_  = _w4158_ ;
	assign \g31074/_0_  = _w4159_ ;
	assign \g31075/_0_  = _w4160_ ;
	assign \g31076/_0_  = _w4161_ ;
	assign \g31077/_0_  = _w4162_ ;
	assign \g31084/u3_syn_4  = _w2570_ ;
	assign \g31085/u3_syn_4  = _w3879_ ;
	assign \g31096/u3_syn_4  = _w3934_ ;
	assign \g31115/u3_syn_4  = _w3974_ ;
	assign \g31136/u3_syn_4  = _w2691_ ;
	assign \g31158/u3_syn_4  = _w2797_ ;
	assign \g31176/u3_syn_4  = _w4063_ ;
	assign \g31193/u3_syn_4  = _w4116_ ;
	assign \g31195/u3_syn_4  = _w4091_ ;
	assign \g31247/u3_syn_4  = _w3905_ ;
	assign \g31280/u3_syn_4  = _w4046_ ;
	assign \g31285/u3_syn_4  = _w4051_ ;
	assign \g31568/_0_  = _w4164_ ;
	assign \g31631/_0_  = _w4188_ ;
	assign \g31672/_0_  = _w4193_ ;
	assign \g31731/_0_  = _w4195_ ;
	assign \g31732/_0_  = _w4196_ ;
	assign \g31742/_2_  = _w4198_ ;
	assign \g31744/_2_  = _w4200_ ;
	assign \g31746/_2_  = _w4202_ ;
	assign \g31748/_2_  = _w4204_ ;
	assign \g31751/_2_  = _w4206_ ;
	assign \g31754/_2_  = _w4208_ ;
	assign \g31756/_2_  = _w4210_ ;
	assign \g31758/_2_  = _w4212_ ;
	assign \g31760/_2_  = _w4214_ ;
	assign \g31761/_0_  = _w4216_ ;
	assign \g31789/_0_  = _w4219_ ;
	assign \g31807/_3_  = _w4222_ ;
	assign \g31825/_3_  = _w4223_ ;
	assign \g32607/_0_  = _w4227_ ;
	assign \g32608/_0_  = _w4231_ ;
	assign \g32609/_0_  = _w4235_ ;
	assign \g32610/_0_  = _w4240_ ;
	assign \g32611/_0_  = _w4244_ ;
	assign \g32612/_0_  = _w4249_ ;
	assign \g32613/_0_  = _w4251_ ;
	assign \g32614/_0_  = _w4253_ ;
	assign \g32615/_0_  = _w4255_ ;
	assign \g32616/_0_  = _w4257_ ;
	assign \g32617/_0_  = _w4259_ ;
	assign \g32618/_0_  = _w4261_ ;
	assign \g32645/_0__syn_2  = _w4262_ ;
	assign \g32687/_0__syn_2  = _w4263_ ;
	assign \g32749/_0__syn_2  = _w4264_ ;
	assign \g32757/_0_  = _w4268_ ;
	assign \g32758/_0_  = _w4271_ ;
	assign \g32759/_0_  = _w4274_ ;
	assign \g32760/_0_  = _w4277_ ;
	assign \g32761/_0_  = _w4280_ ;
	assign \g32762/_0_  = _w4283_ ;
	assign \g32763/_0_  = _w4286_ ;
	assign \g32764/_0_  = _w4289_ ;
	assign \g32765/_0_  = _w4292_ ;
	assign \g32769/_0_  = _w4293_ ;
	assign \g32835/_1_  = _w2689_ ;
	assign \g32839/_0_  = _w4294_ ;
	assign \g32844/_0_  = _w4295_ ;
	assign \g32901/_1_  = _w2795_ ;
	assign \g32902/_0_  = _w4296_ ;
	assign \g32963/_1_  = _w2568_ ;
	assign \g32972/_0_  = _w4297_ ;
	assign \g32977/_0_  = _w4298_ ;
	assign \g32979/_0_  = _w4299_ ;
	assign \g32980/_0_  = _w4300_ ;
	assign \g32981/_0_  = _w4301_ ;
	assign \g32982/_0_  = _w4302_ ;
	assign \g32983/_0_  = _w4303_ ;
	assign \g32987/_0_  = _w4304_ ;
	assign \g33018/_0_  = _w4305_ ;
	assign \g33019/_0_  = _w4308_ ;
	assign \g33088/_0_  = _w4311_ ;
	assign \g33261/_0_  = _w4314_ ;
	assign \g33264/_0_  = _w4316_ ;
	assign \g33275/_0_  = _w4317_ ;
	assign \g33276/_0_  = _w4318_ ;
	assign \g33277/_0_  = _w4319_ ;
	assign \g33371/_0_  = _w4323_ ;
	assign \g33382/_0_  = _w4326_ ;
	assign \g33401/_0_  = _w4329_ ;
	assign \g33402/_0_  = _w4332_ ;
	assign \g33403/_0_  = _w4335_ ;
	assign \g33404/_0_  = _w4338_ ;
	assign \g33405/_0_  = _w4341_ ;
	assign \g33406/_0_  = _w4344_ ;
	assign \g33407/_0_  = _w4347_ ;
	assign \g33408/_0_  = _w4350_ ;
	assign \g33409/_0_  = _w4353_ ;
	assign \g33410/_0_  = _w4356_ ;
	assign \g33411/_0_  = _w4359_ ;
	assign \g33412/_0_  = _w4362_ ;
	assign \g33413/_0_  = _w4365_ ;
	assign \g33414/_0_  = _w4368_ ;
	assign \g33415/_0_  = _w4371_ ;
	assign \g33416/_0_  = _w4374_ ;
	assign \g33417/_0_  = _w4377_ ;
	assign \g33418/_0_  = _w4380_ ;
	assign \g33419/_0_  = _w4383_ ;
	assign \g33420/_0_  = _w4386_ ;
	assign \g33421/_0_  = _w4389_ ;
	assign \g33422/_0_  = _w4392_ ;
	assign \g33423/_0_  = _w4395_ ;
	assign \g33424/_0_  = _w4398_ ;
	assign \g33425/_0_  = _w4401_ ;
	assign \g33426/_0_  = _w4404_ ;
	assign \g33427/_0_  = _w4407_ ;
	assign \g33428/_0_  = _w4410_ ;
	assign \g33429/_0_  = _w4413_ ;
	assign \g33430/_0_  = _w4416_ ;
	assign \g33431/_0_  = _w4419_ ;
	assign \g33432/_0_  = _w4422_ ;
	assign \g33433/_0_  = _w4425_ ;
	assign \g33434/_0_  = _w4428_ ;
	assign \g33435/_0_  = _w4431_ ;
	assign \g33436/_0_  = _w4434_ ;
	assign \g33437/_0_  = _w4437_ ;
	assign \g33438/_0_  = _w4440_ ;
	assign \g33439/_0_  = _w4443_ ;
	assign \g33440/_0_  = _w4446_ ;
	assign \g33441/_0_  = _w4449_ ;
	assign \g33442/_0_  = _w4452_ ;
	assign \g33443/_0_  = _w4455_ ;
	assign \g33444/_0_  = _w4458_ ;
	assign \g33445/_0_  = _w4461_ ;
	assign \g33446/_0_  = _w4464_ ;
	assign \g33447/_0_  = _w4467_ ;
	assign \g33448/_0_  = _w4470_ ;
	assign \g33449/_0_  = _w4473_ ;
	assign \g33450/_0_  = _w4476_ ;
	assign \g33451/_0_  = _w4479_ ;
	assign \g33452/_0_  = _w4482_ ;
	assign \g33453/_0_  = _w4485_ ;
	assign \g33454/_0_  = _w4488_ ;
	assign \g33455/_0_  = _w4491_ ;
	assign \g33456/_0_  = _w4494_ ;
	assign \g33457/_0_  = _w4497_ ;
	assign \g33458/_0_  = _w4500_ ;
	assign \g33459/_0_  = _w4503_ ;
	assign \g33460/_0_  = _w4506_ ;
	assign \g33461/_0_  = _w4509_ ;
	assign \g33462/_0_  = _w4512_ ;
	assign \g33463/_0_  = _w4515_ ;
	assign \g33464/_0_  = _w4518_ ;
	assign \g33465/_0_  = _w4521_ ;
	assign \g33466/_0_  = _w4524_ ;
	assign \g33467/_0_  = _w4527_ ;
	assign \g33468/_0_  = _w4530_ ;
	assign \g33469/_0_  = _w4533_ ;
	assign \g33470/_0_  = _w4536_ ;
	assign \g33471/_0_  = _w4539_ ;
	assign \g33472/_0_  = _w4542_ ;
	assign \g33473/_0_  = _w4545_ ;
	assign \g33474/_0_  = _w4548_ ;
	assign \g33475/_0_  = _w4551_ ;
	assign \g33476/_0_  = _w4554_ ;
	assign \g33477/_0_  = _w4557_ ;
	assign \g33478/_0_  = _w4560_ ;
	assign \g33479/_0_  = _w4563_ ;
	assign \g33480/_0_  = _w4566_ ;
	assign \g33481/_0_  = _w4569_ ;
	assign \g33482/_0_  = _w4572_ ;
	assign \g33483/_0_  = _w4575_ ;
	assign \g33484/_0_  = _w4578_ ;
	assign \g33485/_0_  = _w4581_ ;
	assign \g33486/_0_  = _w4584_ ;
	assign \g33487/_0_  = _w4587_ ;
	assign \g33488/_0_  = _w4590_ ;
	assign \g33489/_0_  = _w4593_ ;
	assign \g33490/_0_  = _w4596_ ;
	assign \g33491/_0_  = _w4599_ ;
	assign \g33492/_0_  = _w4602_ ;
	assign \g33493/_0_  = _w4605_ ;
	assign \g33494/_0_  = _w4608_ ;
	assign \g33495/_0_  = _w4611_ ;
	assign \g33496/_0_  = _w4614_ ;
	assign \g33497/_0_  = _w4617_ ;
	assign \g33498/_0_  = _w4620_ ;
	assign \g33499/_0_  = _w4623_ ;
	assign \g33500/_0_  = _w4626_ ;
	assign \g33501/_0_  = _w4629_ ;
	assign \g33502/_0_  = _w4632_ ;
	assign \g33503/_0_  = _w4635_ ;
	assign \g33504/_0_  = _w4638_ ;
	assign \g33505/_0_  = _w4641_ ;
	assign \g33506/_0_  = _w4644_ ;
	assign \g33507/_0_  = _w4647_ ;
	assign \g33508/_0_  = _w4650_ ;
	assign \g33509/_0_  = _w4653_ ;
	assign \g33510/_0_  = _w4656_ ;
	assign \g33511/_0_  = _w4659_ ;
	assign \g33512/_0_  = _w4662_ ;
	assign \g33513/_0_  = _w4665_ ;
	assign \g33514/_0_  = _w4668_ ;
	assign \g33515/_0_  = _w4671_ ;
	assign \g33516/_0_  = _w4674_ ;
	assign \g33517/_0_  = _w4677_ ;
	assign \g33518/_0_  = _w4680_ ;
	assign \g33519/_0_  = _w4683_ ;
	assign \g33520/_0_  = _w4686_ ;
	assign \g33521/_0_  = _w4689_ ;
	assign \g33522/_0_  = _w4692_ ;
	assign \g33523/_0_  = _w4695_ ;
	assign \g33524/_0_  = _w4698_ ;
	assign \g33525/_0_  = _w4701_ ;
	assign \g33526/_0_  = _w4704_ ;
	assign \g33527/_0_  = _w4707_ ;
	assign \g33528/_0_  = _w4710_ ;
	assign \g33529/_0_  = _w4713_ ;
	assign \g33530/_0_  = _w4716_ ;
	assign \g33531/_0_  = _w4719_ ;
	assign \g33532/_0_  = _w4722_ ;
	assign \g33533/_0_  = _w4725_ ;
	assign \g33534/_0_  = _w4728_ ;
	assign \g33535/_0_  = _w4731_ ;
	assign \g33536/_0_  = _w4734_ ;
	assign \g33537/_0_  = _w4737_ ;
	assign \g33538/_0_  = _w4740_ ;
	assign \g33539/_0_  = _w4743_ ;
	assign \g33540/_0_  = _w4746_ ;
	assign \g33541/_0_  = _w4749_ ;
	assign \g33542/_0_  = _w4752_ ;
	assign \g33543/_0_  = _w4755_ ;
	assign \g33544/_0_  = _w4758_ ;
	assign \g33545/_0_  = _w4761_ ;
	assign \g33546/_0_  = _w4764_ ;
	assign \g33547/_0_  = _w4767_ ;
	assign \g33548/_0_  = _w4770_ ;
	assign \g33549/_0_  = _w4773_ ;
	assign \g33550/_0_  = _w4776_ ;
	assign \g33551/_0_  = _w4779_ ;
	assign \g33552/_0_  = _w4782_ ;
	assign \g33553/_0_  = _w4785_ ;
	assign \g33554/_0_  = _w4788_ ;
	assign \g33555/_0_  = _w4791_ ;
	assign \g33556/_0_  = _w4794_ ;
	assign \g33557/_0_  = _w4797_ ;
	assign \g33558/_0_  = _w4800_ ;
	assign \g33559/_0_  = _w4803_ ;
	assign \g33560/_0_  = _w4806_ ;
	assign \g33561/_0_  = _w4809_ ;
	assign \g33562/_0_  = _w4812_ ;
	assign \g33563/_0_  = _w4815_ ;
	assign \g33564/_0_  = _w4818_ ;
	assign \g33565/_0_  = _w4821_ ;
	assign \g33566/_0_  = _w4824_ ;
	assign \g33567/_0_  = _w4827_ ;
	assign \g33568/_0_  = _w4830_ ;
	assign \g33569/_0_  = _w4833_ ;
	assign \g33570/_0_  = _w4836_ ;
	assign \g33571/_0_  = _w4839_ ;
	assign \g33572/_0_  = _w4842_ ;
	assign \g33573/_0_  = _w4845_ ;
	assign \g33574/_0_  = _w4848_ ;
	assign \g33575/_0_  = _w4851_ ;
	assign \g33576/_0_  = _w4854_ ;
	assign \g33577/_0_  = _w4857_ ;
	assign \g33578/_0_  = _w4860_ ;
	assign \g33579/_0_  = _w4863_ ;
	assign \g33580/_0_  = _w4866_ ;
	assign \g33581/_0_  = _w4869_ ;
	assign \g33582/_0_  = _w4872_ ;
	assign \g33583/_0_  = _w4875_ ;
	assign \g33584/_0_  = _w4878_ ;
	assign \g33585/_0_  = _w4881_ ;
	assign \g33586/_0_  = _w4884_ ;
	assign \g33587/_0_  = _w4887_ ;
	assign \g33588/_0_  = _w4890_ ;
	assign \g33589/_0_  = _w4893_ ;
	assign \g33590/_0_  = _w4896_ ;
	assign \g33591/_0_  = _w4899_ ;
	assign \g33592/_0_  = _w4902_ ;
	assign \g33593/_0_  = _w4905_ ;
	assign \g33594/_0_  = _w4908_ ;
	assign \g33595/_0_  = _w4911_ ;
	assign \g33596/_0_  = _w4914_ ;
	assign \g33597/_0_  = _w4917_ ;
	assign \g33598/_0_  = _w4920_ ;
	assign \g33599/_0_  = _w4923_ ;
	assign \g33600/_0_  = _w4926_ ;
	assign \g33601/_0_  = _w4929_ ;
	assign \g33602/_0_  = _w4932_ ;
	assign \g33603/_0_  = _w4935_ ;
	assign \g33604/_0_  = _w4938_ ;
	assign \g33605/_0_  = _w4941_ ;
	assign \g33606/_0_  = _w4944_ ;
	assign \g33607/_0_  = _w4947_ ;
	assign \g33608/_0_  = _w4950_ ;
	assign \g33609/_0_  = _w4953_ ;
	assign \g33610/_0_  = _w4956_ ;
	assign \g33611/_0_  = _w4959_ ;
	assign \g33612/_0_  = _w4962_ ;
	assign \g33613/_0_  = _w4965_ ;
	assign \g33614/_0_  = _w4968_ ;
	assign \g33615/_0_  = _w4971_ ;
	assign \g33616/_0_  = _w4974_ ;
	assign \g33617/_0_  = _w4977_ ;
	assign \g33618/_0_  = _w4980_ ;
	assign \g33619/_0_  = _w4983_ ;
	assign \g33620/_0_  = _w4986_ ;
	assign \g33621/_0_  = _w4989_ ;
	assign \g33622/_0_  = _w4992_ ;
	assign \g33623/_0_  = _w4995_ ;
	assign \g33624/_0_  = _w4998_ ;
	assign \g33625/_0_  = _w5001_ ;
	assign \g33626/_0_  = _w5004_ ;
	assign \g33627/_0_  = _w5007_ ;
	assign \g33628/_0_  = _w5010_ ;
	assign \g33629/_0_  = _w5013_ ;
	assign \g33630/_0_  = _w5016_ ;
	assign \g33631/_0_  = _w5019_ ;
	assign \g33632/_0_  = _w5022_ ;
	assign \g33633/_0_  = _w5025_ ;
	assign \g33634/_0_  = _w5028_ ;
	assign \g33635/_0_  = _w5031_ ;
	assign \g33636/_0_  = _w5034_ ;
	assign \g33637/_0_  = _w5037_ ;
	assign \g33638/_0_  = _w5040_ ;
	assign \g33639/_0_  = _w5043_ ;
	assign \g33640/_0_  = _w5046_ ;
	assign \g33641/_0_  = _w5049_ ;
	assign \g33642/_0_  = _w5052_ ;
	assign \g33643/_0_  = _w5055_ ;
	assign \g33644/_0_  = _w5058_ ;
	assign \g33645/_0_  = _w5061_ ;
	assign \g33646/_0_  = _w5064_ ;
	assign \g33647/_0_  = _w5067_ ;
	assign \g33648/_0_  = _w5070_ ;
	assign \g33649/_0_  = _w5073_ ;
	assign \g33650/_0_  = _w5076_ ;
	assign \g33651/_0_  = _w5079_ ;
	assign \g33652/_0_  = _w5082_ ;
	assign \g33653/_0_  = _w5085_ ;
	assign \g33654/_0_  = _w5088_ ;
	assign \g33655/_0_  = _w5091_ ;
	assign \g33656/_0_  = _w5094_ ;
	assign \g33657/_0_  = _w5097_ ;
	assign \g33658/_0_  = _w5100_ ;
	assign \g33659/_0_  = _w5103_ ;
	assign \g33660/_0_  = _w5106_ ;
	assign \g33661/_0_  = _w5109_ ;
	assign \g33662/_0_  = _w5112_ ;
	assign \g33663/_0_  = _w5115_ ;
	assign \g33664/_0_  = _w5118_ ;
	assign \g33665/_0_  = _w5121_ ;
	assign \g33666/_0_  = _w5124_ ;
	assign \g33667/_0_  = _w5127_ ;
	assign \g33668/_0_  = _w5130_ ;
	assign \g33669/_0_  = _w5133_ ;
	assign \g33670/_0_  = _w5136_ ;
	assign \g33671/_0_  = _w5139_ ;
	assign \g33672/_0_  = _w5142_ ;
	assign \g33673/_0_  = _w5145_ ;
	assign \g33674/_0_  = _w5148_ ;
	assign \g33675/_0_  = _w5151_ ;
	assign \g33676/_0_  = _w5154_ ;
	assign \g33677/_0_  = _w5157_ ;
	assign \g33678/_0_  = _w5160_ ;
	assign \g33679/_0_  = _w5163_ ;
	assign \g33680/_0_  = _w5166_ ;
	assign \g33681/_0_  = _w5169_ ;
	assign \g33682/_0_  = _w5172_ ;
	assign \g33683/_0_  = _w5175_ ;
	assign \g33684/_0_  = _w5178_ ;
	assign \g33685/_0_  = _w5181_ ;
	assign \g33686/_0_  = _w5184_ ;
	assign \g33687/_0_  = _w5187_ ;
	assign \g33688/_0_  = _w5190_ ;
	assign \g33689/_0_  = _w5193_ ;
	assign \g33690/_0_  = _w5196_ ;
	assign \g33691/_0_  = _w5199_ ;
	assign \g33692/_0_  = _w5202_ ;
	assign \g33693/_0_  = _w5205_ ;
	assign \g33694/_0_  = _w5208_ ;
	assign \g33695/_0_  = _w5211_ ;
	assign \g33696/_0_  = _w5214_ ;
	assign \g33697/_0_  = _w5217_ ;
	assign \g33698/_0_  = _w5220_ ;
	assign \g33699/_0_  = _w5223_ ;
	assign \g33700/_0_  = _w5226_ ;
	assign \g33701/_0_  = _w5229_ ;
	assign \g33702/_0_  = _w5232_ ;
	assign \g33703/_0_  = _w5235_ ;
	assign \g33704/_0_  = _w5238_ ;
	assign \g33705/_0_  = _w5241_ ;
	assign \g33706/_0_  = _w5244_ ;
	assign \g33707/_0_  = _w5247_ ;
	assign \g33708/_0_  = _w5250_ ;
	assign \g33709/_0_  = _w5253_ ;
	assign \g33710/_0_  = _w5256_ ;
	assign \g33711/_0_  = _w5259_ ;
	assign \g33712/_0_  = _w5262_ ;
	assign \g33713/_0_  = _w5265_ ;
	assign \g33714/_0_  = _w5268_ ;
	assign \g33715/_0_  = _w5271_ ;
	assign \g33716/_0_  = _w5274_ ;
	assign \g33717/_0_  = _w5277_ ;
	assign \g33718/_0_  = _w5280_ ;
	assign \g33719/_0_  = _w5283_ ;
	assign \g33720/_0_  = _w5286_ ;
	assign \g33721/_0_  = _w5289_ ;
	assign \g33722/_0_  = _w5292_ ;
	assign \g33723/_0_  = _w5295_ ;
	assign \g33724/_0_  = _w5298_ ;
	assign \g33725/_0_  = _w5301_ ;
	assign \g33726/_0_  = _w5304_ ;
	assign \g33727/_0_  = _w5307_ ;
	assign \g33728/_0_  = _w5310_ ;
	assign \g33729/_0_  = _w5313_ ;
	assign \g33730/_0_  = _w5316_ ;
	assign \g33731/_0_  = _w5319_ ;
	assign \g33732/_0_  = _w5322_ ;
	assign \g33733/_0_  = _w5325_ ;
	assign \g33734/_0_  = _w5328_ ;
	assign \g33735/_0_  = _w5331_ ;
	assign \g33736/_0_  = _w5334_ ;
	assign \g33737/_0_  = _w5337_ ;
	assign \g33738/_0_  = _w5340_ ;
	assign \g33739/_0_  = _w5343_ ;
	assign \g33740/_0_  = _w5346_ ;
	assign \g33741/_0_  = _w5349_ ;
	assign \g33742/_0_  = _w5352_ ;
	assign \g33743/_0_  = _w5355_ ;
	assign \g33744/_0_  = _w5358_ ;
	assign \g33745/_0_  = _w5361_ ;
	assign \g33746/_0_  = _w5364_ ;
	assign \g33747/_0_  = _w5367_ ;
	assign \g33748/_0_  = _w5370_ ;
	assign \g33749/_0_  = _w5373_ ;
	assign \g33750/_0_  = _w5376_ ;
	assign \g33751/_0_  = _w5379_ ;
	assign \g33752/_0_  = _w5382_ ;
	assign \g33753/_0_  = _w5385_ ;
	assign \g33754/_0_  = _w5388_ ;
	assign \g33755/_0_  = _w5391_ ;
	assign \g33756/_0_  = _w5394_ ;
	assign \g33757/_0_  = _w5397_ ;
	assign \g33758/_0_  = _w5400_ ;
	assign \g33759/_0_  = _w5403_ ;
	assign \g33760/_0_  = _w5406_ ;
	assign \g33761/_0_  = _w5409_ ;
	assign \g33762/_0_  = _w5412_ ;
	assign \g33763/_0_  = _w5415_ ;
	assign \g33764/_0_  = _w5418_ ;
	assign \g33765/_0_  = _w5421_ ;
	assign \g33766/_0_  = _w5424_ ;
	assign \g33767/_0_  = _w5427_ ;
	assign \g33768/_0_  = _w5430_ ;
	assign \g33769/_0_  = _w5433_ ;
	assign \g33770/_0_  = _w5436_ ;
	assign \g33771/_0_  = _w5439_ ;
	assign \g33772/_0_  = _w5442_ ;
	assign \g33773/_0_  = _w5445_ ;
	assign \g33774/_0_  = _w5448_ ;
	assign \g33775/_0_  = _w5451_ ;
	assign \g33776/_0_  = _w5454_ ;
	assign \g33777/_0_  = _w5457_ ;
	assign \g33778/_0_  = _w5460_ ;
	assign \g33779/_0_  = _w5463_ ;
	assign \g33780/_0_  = _w5466_ ;
	assign \g33781/_0_  = _w5469_ ;
	assign \g33782/_0_  = _w5472_ ;
	assign \g33783/_0_  = _w5475_ ;
	assign \g33784/_0_  = _w5478_ ;
	assign \g33785/_0_  = _w5481_ ;
	assign \g33786/_0_  = _w5484_ ;
	assign \g33787/_0_  = _w5487_ ;
	assign \g33788/_0_  = _w5490_ ;
	assign \g33789/_0_  = _w5493_ ;
	assign \g33790/_0_  = _w5496_ ;
	assign \g33791/_0_  = _w5499_ ;
	assign \g33792/_0_  = _w5502_ ;
	assign \g33793/_0_  = _w5505_ ;
	assign \g33794/_0_  = _w5508_ ;
	assign \g33795/_0_  = _w5511_ ;
	assign \g33796/_0_  = _w5514_ ;
	assign \g33797/_0_  = _w5517_ ;
	assign \g33798/_0_  = _w5520_ ;
	assign \g33799/_0_  = _w5523_ ;
	assign \g33800/_0_  = _w5526_ ;
	assign \g33801/_0_  = _w5529_ ;
	assign \g33802/_0_  = _w5532_ ;
	assign \g33803/_0_  = _w5535_ ;
	assign \g33804/_0_  = _w5538_ ;
	assign \g33805/_0_  = _w5541_ ;
	assign \g33806/_0_  = _w5544_ ;
	assign \g33807/_0_  = _w5547_ ;
	assign \g33808/_0_  = _w5550_ ;
	assign \g33809/_0_  = _w5553_ ;
	assign \g33810/_0_  = _w5556_ ;
	assign \g33811/_0_  = _w5559_ ;
	assign \g33812/_0_  = _w5562_ ;
	assign \g33813/_0_  = _w5565_ ;
	assign \g33814/_0_  = _w5568_ ;
	assign \g33815/_0_  = _w5571_ ;
	assign \g33816/_0_  = _w5574_ ;
	assign \g33817/_0_  = _w5577_ ;
	assign \g33818/_0_  = _w5580_ ;
	assign \g33819/_0_  = _w5583_ ;
	assign \g33820/_0_  = _w5586_ ;
	assign \g33821/_0_  = _w5589_ ;
	assign \g33822/_0_  = _w5592_ ;
	assign \g33823/_0_  = _w5595_ ;
	assign \g33824/_0_  = _w5598_ ;
	assign \g33825/_0_  = _w5601_ ;
	assign \g33826/_0_  = _w5604_ ;
	assign \g33827/_0_  = _w5607_ ;
	assign \g33828/_0_  = _w5610_ ;
	assign \g33829/_0_  = _w5613_ ;
	assign \g33830/_0_  = _w5616_ ;
	assign \g33831/_0_  = _w5619_ ;
	assign \g33832/_0_  = _w5622_ ;
	assign \g33833/_0_  = _w5625_ ;
	assign \g33834/_0_  = _w5628_ ;
	assign \g33835/_0_  = _w5631_ ;
	assign \g33836/_0_  = _w5634_ ;
	assign \g33837/_0_  = _w5637_ ;
	assign \g33838/_0_  = _w5640_ ;
	assign \g33839/_0_  = _w5643_ ;
	assign \g33840/_0_  = _w5646_ ;
	assign \g33841/_0_  = _w5649_ ;
	assign \g33842/_0_  = _w5652_ ;
	assign \g33843/_0_  = _w5655_ ;
	assign \g33844/_0_  = _w5658_ ;
	assign \g33845/_0_  = _w5661_ ;
	assign \g33846/_0_  = _w5664_ ;
	assign \g33847/_0_  = _w5667_ ;
	assign \g33848/_0_  = _w5670_ ;
	assign \g33849/_0_  = _w5673_ ;
	assign \g33850/_0_  = _w5676_ ;
	assign \g33851/_0_  = _w5679_ ;
	assign \g33852/_0_  = _w5682_ ;
	assign \g33853/_0_  = _w5685_ ;
	assign \g33854/_0_  = _w5688_ ;
	assign \g33855/_0_  = _w5691_ ;
	assign \g33856/_0_  = _w5694_ ;
	assign \g33857/_0_  = _w5697_ ;
	assign \g33858/_0_  = _w5700_ ;
	assign \g33859/_0_  = _w5703_ ;
	assign \g33860/_0_  = _w5706_ ;
	assign \g33861/_0_  = _w5709_ ;
	assign \g33862/_0_  = _w5712_ ;
	assign \g33863/_0_  = _w5715_ ;
	assign \g33864/_0_  = _w5718_ ;
	assign \g33865/_0_  = _w5721_ ;
	assign \g33866/_0_  = _w5724_ ;
	assign \g33867/_0_  = _w5727_ ;
	assign \g33868/_0_  = _w5730_ ;
	assign \g33869/_0_  = _w5733_ ;
	assign \g33870/_0_  = _w5736_ ;
	assign \g33871/_0_  = _w5739_ ;
	assign \g33872/_0_  = _w5742_ ;
	assign \g33873/_0_  = _w5745_ ;
	assign \g33874/_0_  = _w5748_ ;
	assign \g33875/_0_  = _w5751_ ;
	assign \g33876/_0_  = _w5754_ ;
	assign \g33877/_0_  = _w5757_ ;
	assign \g33878/_0_  = _w5760_ ;
	assign \g33879/_0_  = _w5763_ ;
	assign \g33880/_0_  = _w5766_ ;
	assign \g33881/_0_  = _w5769_ ;
	assign \g33882/_0_  = _w5772_ ;
	assign \g33883/_0_  = _w5775_ ;
	assign \g33884/_0_  = _w5778_ ;
	assign \g33885/_0_  = _w5781_ ;
	assign \g33886/_0_  = _w5784_ ;
	assign \g33887/_0_  = _w5787_ ;
	assign \g33888/_0_  = _w5790_ ;
	assign \g33889/_0_  = _w5793_ ;
	assign \g33890/_0_  = _w5796_ ;
	assign \g33891/_0_  = _w5799_ ;
	assign \g33892/_0_  = _w5802_ ;
	assign \g33893/_0_  = _w5805_ ;
	assign \g33894/_0_  = _w5808_ ;
	assign \g33895/_0_  = _w5811_ ;
	assign \g33896/_0_  = _w5814_ ;
	assign \g33897/_0_  = _w5817_ ;
	assign \g33898/_0_  = _w5820_ ;
	assign \g33899/_0_  = _w5823_ ;
	assign \g33900/_0_  = _w5826_ ;
	assign \g33901/_0_  = _w5829_ ;
	assign \g33902/_0_  = _w5832_ ;
	assign \g33903/_0_  = _w5835_ ;
	assign \g33904/_0_  = _w5838_ ;
	assign \g33905/_0_  = _w5841_ ;
	assign \g33906/_0_  = _w5844_ ;
	assign \g33907/_0_  = _w5847_ ;
	assign \g33908/_0_  = _w5850_ ;
	assign \g33909/_0_  = _w5853_ ;
	assign \g33910/_0_  = _w5856_ ;
	assign \g33911/_0_  = _w5859_ ;
	assign \g33912/_0_  = _w5862_ ;
	assign \g33913/_0_  = _w5865_ ;
	assign \g33914/_0_  = _w5868_ ;
	assign \g33915/_0_  = _w5871_ ;
	assign \g33916/_0_  = _w5874_ ;
	assign \g33917/_0_  = _w5877_ ;
	assign \g33918/_0_  = _w5880_ ;
	assign \g33919/_0_  = _w5883_ ;
	assign \g33920/_0_  = _w5886_ ;
	assign \g33921/_0_  = _w5889_ ;
	assign \g33922/_0_  = _w5892_ ;
	assign \g33923/_0_  = _w5895_ ;
	assign \g33924/_0_  = _w5898_ ;
	assign \g33925/_0_  = _w5901_ ;
	assign \g33926/_0_  = _w5904_ ;
	assign \g33927/_0_  = _w5907_ ;
	assign \g33928/_0_  = _w5910_ ;
	assign \g33929/_0_  = _w5913_ ;
	assign \g33930/_0_  = _w5916_ ;
	assign \g33931/_0_  = _w5919_ ;
	assign \g33932/_0_  = _w5922_ ;
	assign \g33933/_0_  = _w5925_ ;
	assign \g33934/_0_  = _w5928_ ;
	assign \g33935/_0_  = _w5931_ ;
	assign \g33936/_0_  = _w5934_ ;
	assign \g33937/_0_  = _w5937_ ;
	assign \g33938/_0_  = _w5940_ ;
	assign \g33939/_0_  = _w5943_ ;
	assign \g33940/_0_  = _w5946_ ;
	assign \g33941/_0_  = _w5949_ ;
	assign \g33942/_0_  = _w5952_ ;
	assign \g33943/_0_  = _w5955_ ;
	assign \g33944/_0_  = _w5958_ ;
	assign \g33945/_0_  = _w5961_ ;
	assign \g33946/_0_  = _w5964_ ;
	assign \g33947/_0_  = _w5967_ ;
	assign \g33948/_0_  = _w5970_ ;
	assign \g33949/_0_  = _w5973_ ;
	assign \g33950/_0_  = _w5976_ ;
	assign \g33951/_0_  = _w5979_ ;
	assign \g33952/_0_  = _w5982_ ;
	assign \g33953/_0_  = _w5985_ ;
	assign \g33954/_0_  = _w5988_ ;
	assign \g33955/_0_  = _w5991_ ;
	assign \g33956/_0_  = _w5994_ ;
	assign \g33957/_0_  = _w5997_ ;
	assign \g33958/_0_  = _w6000_ ;
	assign \g33959/_0_  = _w6003_ ;
	assign \g33960/_0_  = _w6006_ ;
	assign \g33961/_0_  = _w6009_ ;
	assign \g33962/_0_  = _w6012_ ;
	assign \g33963/_0_  = _w6015_ ;
	assign \g33964/_0_  = _w6018_ ;
	assign \g33965/_0_  = _w6021_ ;
	assign \g33966/_0_  = _w6024_ ;
	assign \g33967/_0_  = _w6027_ ;
	assign \g33968/_0_  = _w6030_ ;
	assign \g33969/_0_  = _w6033_ ;
	assign \g33970/_0_  = _w6036_ ;
	assign \g33971/_0_  = _w6039_ ;
	assign \g33972/_0_  = _w6042_ ;
	assign \g33973/_0_  = _w6045_ ;
	assign \g33974/_0_  = _w6048_ ;
	assign \g33975/_0_  = _w6051_ ;
	assign \g33976/_0_  = _w6054_ ;
	assign \g33977/u3_syn_4  = _w6055_ ;
	assign \g33981/u3_syn_4  = _w6056_ ;
	assign \g34014/u3_syn_4  = _w6057_ ;
	assign \g34047/u3_syn_4  = _w6058_ ;
	assign \g34084/u3_syn_4  = _w6059_ ;
	assign \g34123/u3_syn_4  = _w6060_ ;
	assign \g34306/_0_  = _w6073_ ;
	assign \g34316/_0_  = _w6086_ ;
	assign \g34324/_0_  = _w6099_ ;
	assign \g34326/_0_  = _w6112_ ;
	assign \g34328/_0_  = _w6125_ ;
	assign \g34331/_0_  = _w6138_ ;
	assign \g34333/_0_  = _w6151_ ;
	assign \g34344/_0_  = _w6164_ ;
	assign \g34347/_0_  = _w6177_ ;
	assign \g34351/_0_  = _w6190_ ;
	assign \g34361/_0_  = _w6203_ ;
	assign \g34368/_0_  = _w6216_ ;
	assign \g34377/_0_  = _w6229_ ;
	assign \g34385/_0_  = _w6242_ ;
	assign \g34393/_0_  = _w6255_ ;
	assign \g34414/_1_  = _w6256_ ;
	assign \g34451/_1_  = _w6257_ ;
	assign \g34476/_1_  = _w6258_ ;
	assign \g34487/_0_  = _w6259_ ;
	assign \g34490/_1_  = _w6260_ ;
	assign \g34715/_0_  = _w6261_ ;
	assign \g34878/_0_  = _w6269_ ;
	assign \g34882/_0_  = _w6277_ ;
	assign \g34883/_0_  = _w6278_ ;
	assign \g34893/_0_  = _w6282_ ;
	assign \g34896/_0_  = _w6291_ ;
	assign \g34898/_0_  = _w6300_ ;
	assign \g34899/_0_  = _w6304_ ;
	assign \g34916/_3_  = _w6305_ ;
	assign \g35264/_0_  = _w6307_ ;
	assign \g35265/_0_  = _w6309_ ;
	assign \g35266/_0_  = _w6311_ ;
	assign \g35267/_0_  = _w6312_ ;
	assign \g35268/_0_  = _w6313_ ;
	assign \g35269/_0_  = _w6314_ ;
	assign \g35270/_0_  = _w6315_ ;
	assign \g35271/_0_  = _w6316_ ;
	assign \g35272/_0_  = _w6328_ ;
	assign \g35273/_0_  = _w6340_ ;
	assign \g35274/_0_  = _w6352_ ;
	assign \g35275/_0_  = _w6353_ ;
	assign \g35276/_0_  = _w6365_ ;
	assign \g35277/_0_  = _w6377_ ;
	assign \g35278/_0_  = _w6389_ ;
	assign \g35279/_0_  = _w6400_ ;
	assign \g35283/_0_  = _w6401_ ;
	assign \g35287/_0_  = _w2564_ ;
	assign \g35294/_0_  = _w4265_ ;
	assign \g35300/_0_  = _w2416_ ;
	assign \g35304/_0_  = _w2425_ ;
	assign \g35308/_0_  = _w2443_ ;
	assign \g35312/_0_  = _w2454_ ;
	assign \g35316/_0_  = _w2154_ ;
	assign \g35318/_0_  = _w2685_ ;
	assign \g35326/_0_  = _w6413_ ;
	assign \g35334/_0_  = _w2791_ ;
	assign \g35336/_0_  = _w6414_ ;
	assign \g35337/_0_  = _w6415_ ;
	assign \g35338/_0_  = _w6416_ ;
	assign \g35357/_0_  = _w6417_ ;
	assign \g35358/_0_  = _w6418_ ;
	assign \g35359/_0_  = _w6419_ ;
	assign \g35419/_0_  = _w6420_ ;
	assign \g35438/_0_  = _w6423_ ;
	assign \g35439/_0_  = _w6424_ ;
	assign \g35440/_0_  = _w6425_ ;
	assign \g35441/_0_  = _w6426_ ;
	assign \g35442/_0_  = _w6427_ ;
	assign \g35444/_0_  = _w6437_ ;
	assign \g35445/_0_  = _w6447_ ;
	assign \g35446/_0_  = _w6457_ ;
	assign \g35447/_0_  = _w6467_ ;
	assign \g35448/_0_  = _w6477_ ;
	assign \g35449/_0_  = _w6481_ ;
	assign \g35450/_0_  = _w6485_ ;
	assign \g35451/_0_  = _w6492_ ;
	assign \g35452/_0_  = _w6493_ ;
	assign \g35463/_0_  = _w6495_ ;
	assign \g35464/_0_  = _w6515_ ;
	assign \g35466/_0_  = _w6516_ ;
	assign \g35485/_2_  = _w6519_ ;
	assign \g35495/_0_  = _w6520_ ;
	assign \g35496/_0_  = _w6521_ ;
	assign \g35499/_0_  = _w6522_ ;
	assign \g35500/_0_  = _w6523_ ;
	assign \g35501/_0_  = _w6524_ ;
	assign \g35502/_0_  = _w6525_ ;
	assign \g35563/_0_  = _w6526_ ;
	assign \g35633/_0_  = _w6527_ ;
	assign \g35717/_0_  = _w6528_ ;
	assign \g35718/_0_  = _w6529_ ;
	assign \g35719/_0_  = _w6530_ ;
	assign \g35809/_0_  = _w6532_ ;
	assign \g35810/_0_  = _w6534_ ;
	assign \g35811/_0_  = _w6536_ ;
	assign \g35812/_0_  = _w6538_ ;
	assign \g35813/_0_  = _w6540_ ;
	assign \g35814/_0_  = _w6542_ ;
	assign \g35815/_0_  = _w6544_ ;
	assign \g35816/_0_  = _w6546_ ;
	assign \g35817/_0_  = _w6548_ ;
	assign \g35818/_0_  = _w6550_ ;
	assign \g35819/_0_  = _w6552_ ;
	assign \g35820/_0_  = _w6554_ ;
	assign \g35821/_0_  = _w6556_ ;
	assign \g35822/_0_  = _w6558_ ;
	assign \g35823/_0_  = _w6560_ ;
	assign \g35824/_0_  = _w6562_ ;
	assign \g35825/_0_  = _w6564_ ;
	assign \g35826/_0_  = _w6566_ ;
	assign \g35827/_0_  = _w6568_ ;
	assign \g35830/_0_  = _w6572_ ;
	assign \g35833/_0_  = _w6574_ ;
	assign \g35835/_0_  = _w6577_ ;
	assign \g35836/_0_  = _w6581_ ;
	assign \g35837/_0_  = _w6585_ ;
	assign \g35839/_0_  = _w6586_ ;
	assign \g35840/_0_  = _w6588_ ;
	assign \g35841/_0_  = _w6592_ ;
	assign \g35843/_0_  = _w6594_ ;
	assign \g35844/_0_  = _w6598_ ;
	assign \g35845/_0_  = _w6599_ ;
	assign \g35853/_0_  = _w6600_ ;
	assign \g35854/_0_  = _w6601_ ;
	assign \g35855/_0_  = _w6603_ ;
	assign \g35856/_0_  = _w6604_ ;
	assign \g36306/_0_  = _w6607_ ;
	assign \g36414/_0_  = _w6608_ ;
	assign \g36415/_0_  = _w6609_ ;
	assign \g36449/_0_  = _w6612_ ;
	assign \g36550/_0_  = _w6613_ ;
	assign \g36551/_0_  = _w6614_ ;
	assign \g36553/_0_  = _w6615_ ;
	assign \g36560/_0_  = _w6616_ ;
	assign \g36562/_3_  = _w6617_ ;
	assign \g36563/_0_  = _w6620_ ;
	assign \g36612/_0_  = _w6621_ ;
	assign \g36614/_2_  = _w6623_ ;
	assign \g36695/_0_  = _w6625_ ;
	assign \g36784/_0_  = _w6628_ ;
	assign \g36785/_0_  = _w6631_ ;
	assign \g36786/_0_  = _w6634_ ;
	assign \g36787/_0_  = _w6637_ ;
	assign \g36788/_0_  = _w6640_ ;
	assign \g36789/_0_  = _w6643_ ;
	assign \g36790/_0_  = _w6646_ ;
	assign \g36791/_0_  = _w6649_ ;
	assign \g36792/_0_  = _w6652_ ;
	assign \g36793/_0_  = _w6655_ ;
	assign \g36794/_0_  = _w6658_ ;
	assign \g36796/_0_  = _w6661_ ;
	assign \g36797/_0_  = _w6664_ ;
	assign \g36798/_0_  = _w6667_ ;
	assign \g36799/_0_  = _w6670_ ;
	assign \g36800/_0_  = _w6673_ ;
	assign \g36801/_0_  = _w6676_ ;
	assign \g36802/_0_  = _w6679_ ;
	assign \g36803/_0_  = _w6682_ ;
	assign \g36804/_0_  = _w6685_ ;
	assign \g36805/_0_  = _w6688_ ;
	assign \g36806/_0_  = _w6691_ ;
	assign \g36807/_0_  = _w6694_ ;
	assign \g36808/_0_  = _w6697_ ;
	assign \g36809/_0_  = _w6700_ ;
	assign \g36810/_0_  = _w6703_ ;
	assign \g36811/_0_  = _w6706_ ;
	assign \g36813/_0_  = _w6709_ ;
	assign \g36814/_0_  = _w6712_ ;
	assign \g36815/_0_  = _w6715_ ;
	assign \g36820/_0_  = _w6718_ ;
	assign \g36825/_0_  = _w6721_ ;
	assign \g36832/_0_  = _w6724_ ;
	assign \g36846/_0_  = _w6727_ ;
	assign \g36855/_0_  = _w6730_ ;
	assign \g36857/_0_  = _w6733_ ;
	assign \g36859/_0_  = _w6736_ ;
	assign \g36860/_0_  = _w6739_ ;
	assign \g36861/_0_  = _w6742_ ;
	assign \g36862/_0_  = _w6745_ ;
	assign \g36863/_0_  = _w6748_ ;
	assign \g36864/_0_  = _w6751_ ;
	assign \g36867/_0_  = _w6754_ ;
	assign \g36870/_0_  = _w6757_ ;
	assign \g36871/_0_  = _w6760_ ;
	assign \g36877/_0_  = _w6763_ ;
	assign \g36879/_0_  = _w6766_ ;
	assign \g36892/_0_  = _w6769_ ;
	assign \g36893/_0_  = _w6772_ ;
	assign \g36901/_0_  = _w6775_ ;
	assign \g36909/_0_  = _w6778_ ;
	assign \g36914/_0_  = _w6781_ ;
	assign \g36919/_0_  = _w6784_ ;
	assign \g36922/_0_  = _w6787_ ;
	assign \g36923/_0_  = _w6790_ ;
	assign \g36927/_0_  = _w6793_ ;
	assign \g36930/_0_  = _w6796_ ;
	assign \g36931/_0_  = _w6799_ ;
	assign \g36933/_0_  = _w6802_ ;
	assign \g36934/_0_  = _w6805_ ;
	assign \g36935/_0_  = _w6808_ ;
	assign \g36936/_0_  = _w6811_ ;
	assign \g36937/_0_  = _w6814_ ;
	assign \g36938/_0_  = _w6817_ ;
	assign \g36939/_0_  = _w6820_ ;
	assign \g36940/_0_  = _w6823_ ;
	assign \g36941/_0_  = _w6826_ ;
	assign \g36943/_0_  = _w6829_ ;
	assign \g36944/_0_  = _w6832_ ;
	assign \g36945/_0_  = _w6835_ ;
	assign \g36946/_0_  = _w6838_ ;
	assign \g36947/_0_  = _w6841_ ;
	assign \g36948/_0_  = _w6844_ ;
	assign \g36949/_0_  = _w6847_ ;
	assign \g36950/_0_  = _w6850_ ;
	assign \g36951/_0_  = _w6853_ ;
	assign \g36952/_0_  = _w6856_ ;
	assign \g36953/_0_  = _w6859_ ;
	assign \g36954/_0_  = _w6862_ ;
	assign \g36957/_0_  = _w6865_ ;
	assign \g36958/_0_  = _w6868_ ;
	assign \g36959/_0_  = _w6871_ ;
	assign \g36960/_0_  = _w6874_ ;
	assign \g36961/_0_  = _w6877_ ;
	assign \g36962/_0_  = _w6880_ ;
	assign \g36963/_0_  = _w6883_ ;
	assign \g36970/_0_  = _w6886_ ;
	assign \g36977/_0_  = _w6889_ ;
	assign \g36986/_0_  = _w6892_ ;
	assign \g36991/_0_  = _w6895_ ;
	assign \g36994/_0_  = _w6898_ ;
	assign \g37015/_0_  = _w6901_ ;
	assign \g37057/_0_  = _w6904_ ;
	assign \g37073/_0_  = _w6907_ ;
	assign \g37128/_0_  = _w6910_ ;
	assign \g37129/_0_  = _w6913_ ;
	assign \g37138/_0_  = _w6916_ ;
	assign \g37139/_0_  = _w6917_ ;
	assign \g37140/_0_  = _w6920_ ;
	assign \g37141/_0_  = _w6923_ ;
	assign \g37142/_0_  = _w6926_ ;
	assign \g37143/_0_  = _w6929_ ;
	assign \g37144/_0_  = _w6932_ ;
	assign \g37145/_0_  = _w6935_ ;
	assign \g37146/_0_  = _w6938_ ;
	assign \g37147/_0_  = _w6941_ ;
	assign \g37148/_0_  = _w6944_ ;
	assign \g37149/_0_  = _w6947_ ;
	assign \g37150/_0_  = _w6950_ ;
	assign \g37151/_0_  = _w6953_ ;
	assign \g37152/_0_  = _w6956_ ;
	assign \g37153/_0_  = _w6959_ ;
	assign \g37154/_0_  = _w6962_ ;
	assign \g37155/_0_  = _w6965_ ;
	assign \g37156/_0_  = _w6968_ ;
	assign \g37157/_0_  = _w6971_ ;
	assign \g37158/_0_  = _w6974_ ;
	assign \g37159/_0_  = _w6977_ ;
	assign \g37160/_0_  = _w6980_ ;
	assign \g37161/_0_  = _w6983_ ;
	assign \g37162/_0_  = _w6986_ ;
	assign \g37163/_0_  = _w6989_ ;
	assign \g37164/_0_  = _w6992_ ;
	assign \g37165/_0_  = _w6995_ ;
	assign \g37166/_0_  = _w6998_ ;
	assign \g37167/_0_  = _w7001_ ;
	assign \g37168/_0_  = _w7004_ ;
	assign \g37169/_0_  = _w7007_ ;
	assign \g37170/_0_  = _w7010_ ;
	assign \g37171/_0_  = _w7013_ ;
	assign \g37172/_0_  = _w7016_ ;
	assign \g37173/_0_  = _w7019_ ;
	assign \g37174/_0_  = _w7022_ ;
	assign \g37175/_0_  = _w7025_ ;
	assign \g37176/_0_  = _w7028_ ;
	assign \g37177/_0_  = _w7031_ ;
	assign \g37178/_0_  = _w7034_ ;
	assign \g37179/_0_  = _w7037_ ;
	assign \g37180/_0_  = _w7040_ ;
	assign \g37181/_0_  = _w7043_ ;
	assign \g37182/_0_  = _w7046_ ;
	assign \g37183/_0_  = _w7049_ ;
	assign \g37184/_0_  = _w7052_ ;
	assign \g37185/_0_  = _w7055_ ;
	assign \g37187/_0_  = _w7058_ ;
	assign \g37188/_0_  = _w7061_ ;
	assign \g37190/_0_  = _w7064_ ;
	assign \g37191/_0_  = _w7067_ ;
	assign \g37192/_0_  = _w7070_ ;
	assign \g37193/_0_  = _w7073_ ;
	assign \g37194/_0_  = _w7076_ ;
	assign \g37372/_3_  = _w7078_ ;
	assign \g37377/_0_  = _w7079_ ;
	assign \g37378/_0_  = _w7080_ ;
	assign \g37379/_0_  = _w7081_ ;
	assign \g37380/_0_  = _w7082_ ;
	assign \g37381/_0_  = _w7083_ ;
	assign \g37382/_0_  = _w7084_ ;
	assign \g37383/_0_  = _w7085_ ;
	assign \g37384/_0_  = _w7086_ ;
	assign \g37385/_0_  = _w7087_ ;
	assign \g37386/_0_  = _w7088_ ;
	assign \g37387/_0_  = _w7089_ ;
	assign \g37388/_0_  = _w7090_ ;
	assign \g37389/_0_  = _w7091_ ;
	assign \g37390/_0_  = _w7092_ ;
	assign \g37391/_0_  = _w7093_ ;
	assign \g37392/_0_  = _w7094_ ;
	assign \g37393/_0_  = _w7095_ ;
	assign \g37394/_0_  = _w7096_ ;
	assign \g37395/_0_  = _w7097_ ;
	assign \g37396/_0_  = _w7098_ ;
	assign \g37397/_0_  = _w7099_ ;
	assign \g37398/_0_  = _w7100_ ;
	assign \g37399/_0_  = _w7101_ ;
	assign \g37400/_0_  = _w7102_ ;
	assign \g37401/_0_  = _w7103_ ;
	assign \g37402/_0_  = _w7104_ ;
	assign \g37403/_0_  = _w7105_ ;
	assign \g37404/_0_  = _w7106_ ;
	assign \g37405/_0_  = _w7107_ ;
	assign \g37406/_0_  = _w7108_ ;
	assign \g37407/_0_  = _w7109_ ;
	assign \g37408/_0_  = _w7110_ ;
	assign \g37409/_0_  = _w7111_ ;
	assign \g37410/_0_  = _w7112_ ;
	assign \g37411/_0_  = _w7113_ ;
	assign \g37412/_0_  = _w7114_ ;
	assign \g37413/_0_  = _w7115_ ;
	assign \g37576/_3_  = _w6597_ ;
	assign \g37590/_2_  = _w2400_ ;
	assign \g40278/_0_  = _w6422_ ;
	assign \g40379/_0_  = _w6273_ ;
	assign \g40389/_2_  = _w6569_ ;
	assign \g40390/_2_  = _w6578_ ;
	assign \g40391/_0_  = _w4245_ ;
	assign \g40393/_2_  = _w6582_ ;
	assign \g40395/_0_  = _w6283_ ;
	assign \g40397/_0_  = _w6265_ ;
	assign \g40400/_0_  = _w4236_ ;
	assign \g40402/_0_  = _w6292_ ;
	assign \g45458/_0_  = _w2152_ ;
	assign \g45675/_0_  = _w7119_ ;
	assign \g45677/_0_  = _w7118_ ;
	assign \g45678/_0_  = _w7123_ ;
	assign \g45682/_0_  = _w7122_ ;
	assign sync_pad_o_pad = _w7124_ ;
	assign \u14_u0_full_empty_r_reg/P0001_reg_syn_3  = _w7125_ ;
	assign \u14_u1_full_empty_r_reg/P0001_reg_syn_3  = _w7126_ ;
	assign \u14_u2_full_empty_r_reg/P0001_reg_syn_3  = _w7127_ ;
	assign \u14_u3_full_empty_r_reg/P0001_reg_syn_3  = _w7128_ ;
	assign \u14_u4_full_empty_r_reg/P0001_reg_syn_3  = _w7129_ ;
	assign \u14_u5_full_empty_r_reg/P0001_reg_syn_3  = _w7130_ ;
	assign \u14_u6_full_empty_r_reg/P0001_reg_syn_3  = _w7131_ ;
	assign \u14_u7_full_empty_r_reg/P0001_reg_syn_3  = _w7132_ ;
	assign \u14_u8_full_empty_r_reg/P0001_reg_syn_3  = _w7133_ ;
	assign \u1_slt0_reg[11]/P0001_reg_syn_3  = _w7134_ ;
	assign \u1_slt0_reg[12]/P0001_reg_syn_3  = _w7135_ ;
	assign \u1_slt0_reg[15]/P0001_reg_syn_3  = _w7136_ ;
	assign \u1_slt0_reg[9]/P0001_reg_syn_3  = _w7137_ ;
	assign \u1_slt1_reg[10]/P0001_reg_syn_3  = _w7138_ ;
	assign \u1_slt1_reg[11]/P0001_reg_syn_3  = _w7139_ ;
	assign \u1_slt1_reg[5]/P0001_reg_syn_3  = _w7140_ ;
	assign \u1_slt1_reg[6]/P0001_reg_syn_3  = _w7141_ ;
	assign \u1_slt1_reg[7]/P0001_reg_syn_3  = _w7142_ ;
	assign \u1_slt1_reg[8]/P0001_reg_syn_3  = _w7143_ ;
	assign wb_err_o_pad = 1'b0;
endmodule;